// Benchmark "top" written by ABC on Thu May 28 22:02:13 2020

module rf_sin ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    sin0 , sin1 , sin2 , sin3 , sin4 , sin5 , sin6 ,
    sin7 , sin8 , sin9 , sin10 , sin11 , sin12 ,
    sin13 , sin14 , sin15 , sin16 , sin17 , sin18 ,
    sin19 , sin20 , sin21 , sin22 , sin23 , sin24   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ;
  output sin0 , sin1 , sin2 , sin3 , sin4 , sin5 , sin6 ,
    sin7 , sin8 , sin9 , sin10 , sin11 , sin12 ,
    sin13 , sin14 , sin15 , sin16 , sin17 , sin18 ,
    sin19 , sin20 , sin21 , sin22 , sin23 , sin24 ;
  wire n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
    n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
    n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
    n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
    n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n792, n793, n794, n795, n796, n799, n800, n801, n802,
    n803, n804, n808, n810, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1057, n1058, n1059, n1060,
    n1061, n1063, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1147,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1704, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1821, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
    n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2272, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
    n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
    n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
    n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
    n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
    n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
    n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
    n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
    n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
    n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
    n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
    n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
    n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
    n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
    n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
    n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
    n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4606,
    n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
    n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
    n4667, n4668, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
    n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
    n4728, n4729, n4730, n4731, n4732, n4733, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
    n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
    n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
    n4942, n4943, n4944, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
    n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
    n5087, n5088, n5089, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5151,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160;
  jnot g0000(.din(a22 ), .dout(n49));
  jor  g0001(.dina(a2 ), .dinb(a1 ), .dout(n50));
  jor  g0002(.dina(n50), .dinb(a0 ), .dout(n51));
  jor  g0003(.dina(n51), .dinb(a3 ), .dout(n52));
  jor  g0004(.dina(n52), .dinb(a4 ), .dout(n53));
  jand g0005(.dina(n53), .dinb(n49), .dout(n54));
  jxor g0006(.dina(n54), .dinb(a5 ), .dout(n55));
  jnot g0007(.din(n55), .dout(n56));
  jand g0008(.dina(n51), .dinb(n49), .dout(n57));
  jxor g0009(.dina(n57), .dinb(a3 ), .dout(n58));
  jnot g0010(.din(n58), .dout(n59));
  jand g0011(.dina(a22 ), .dinb(a2 ), .dout(n60));
  jnot g0012(.din(a0 ), .dout(n61));
  jnot g0013(.din(a1 ), .dout(n62));
  jand g0014(.dina(n62), .dinb(n61), .dout(n63));
  jnot g0015(.din(n63), .dout(n64));
  jand g0016(.dina(n64), .dinb(a2 ), .dout(n65));
  jnot g0017(.din(n65), .dout(n66));
  jand g0018(.dina(n66), .dinb(n57), .dout(n67));
  jor  g0019(.dina(n67), .dinb(n60), .dout(n68));
  jxor g0020(.dina(n68), .dinb(n59), .dout(n69));
  jnot g0021(.din(n69), .dout(n70));
  jand g0022(.dina(a22 ), .dinb(a4 ), .dout(n71));
  jand g0023(.dina(n52), .dinb(a4 ), .dout(n72));
  jnot g0024(.din(n72), .dout(n73));
  jand g0025(.dina(n73), .dinb(n54), .dout(n74));
  jor  g0026(.dina(n74), .dinb(n71), .dout(n75));
  jxor g0027(.dina(n75), .dinb(n56), .dout(n76));
  jnot g0028(.din(n76), .dout(n77));
  jand g0029(.dina(n77), .dinb(n70), .dout(n78));
  jnot g0030(.din(n78), .dout(n79));
  jand g0031(.dina(a22 ), .dinb(a15 ), .dout(n80));
  jor  g0032(.dina(n53), .dinb(a5 ), .dout(n81));
  jor  g0033(.dina(n81), .dinb(a6 ), .dout(n82));
  jor  g0034(.dina(n82), .dinb(a7 ), .dout(n83));
  jor  g0035(.dina(n83), .dinb(a8 ), .dout(n84));
  jor  g0036(.dina(n84), .dinb(a9 ), .dout(n85));
  jor  g0037(.dina(n85), .dinb(a10 ), .dout(n86));
  jor  g0038(.dina(n86), .dinb(a11 ), .dout(n87));
  jor  g0039(.dina(n87), .dinb(a12 ), .dout(n88));
  jor  g0040(.dina(n88), .dinb(a13 ), .dout(n89));
  jor  g0041(.dina(n89), .dinb(a14 ), .dout(n90));
  jor  g0042(.dina(n90), .dinb(a15 ), .dout(n91));
  jand g0043(.dina(n91), .dinb(n49), .dout(n92));
  jand g0044(.dina(n90), .dinb(a15 ), .dout(n93));
  jnot g0045(.din(n93), .dout(n94));
  jand g0046(.dina(n94), .dinb(n92), .dout(n95));
  jor  g0047(.dina(n95), .dinb(n80), .dout(n96));
  jor  g0048(.dina(n91), .dinb(a16 ), .dout(n97));
  jor  g0049(.dina(n97), .dinb(a17 ), .dout(n98));
  jor  g0050(.dina(n98), .dinb(a18 ), .dout(n99));
  jor  g0051(.dina(n99), .dinb(a19 ), .dout(n100));
  jor  g0052(.dina(n100), .dinb(a20 ), .dout(n101));
  jand g0053(.dina(n101), .dinb(n49), .dout(n102));
  jxor g0054(.dina(n102), .dinb(a21 ), .dout(n103));
  jand g0055(.dina(a22 ), .dinb(a20 ), .dout(n104));
  jand g0056(.dina(n100), .dinb(a20 ), .dout(n105));
  jnot g0057(.din(n105), .dout(n106));
  jand g0058(.dina(n106), .dinb(n102), .dout(n107));
  jor  g0059(.dina(n107), .dinb(n104), .dout(n108));
  jand g0060(.dina(n108), .dinb(n103), .dout(n109));
  jand g0061(.dina(n109), .dinb(n96), .dout(n110));
  jand g0062(.dina(a22 ), .dinb(a18 ), .dout(n111));
  jand g0063(.dina(n99), .dinb(n49), .dout(n112));
  jand g0064(.dina(n98), .dinb(a18 ), .dout(n113));
  jnot g0065(.din(n113), .dout(n114));
  jand g0066(.dina(n114), .dinb(n112), .dout(n115));
  jor  g0067(.dina(n115), .dinb(n111), .dout(n116));
  jxor g0068(.dina(n112), .dinb(a19 ), .dout(n117));
  jnot g0069(.din(n117), .dout(n118));
  jor  g0070(.dina(n118), .dinb(n116), .dout(n119));
  jnot g0071(.din(n119), .dout(n120));
  jnot g0072(.din(a17 ), .dout(n121));
  jand g0073(.dina(n97), .dinb(n49), .dout(n122));
  jxor g0074(.dina(n122), .dinb(n121), .dout(n123));
  jnot g0075(.din(n123), .dout(n124));
  jxor g0076(.dina(n92), .dinb(a16 ), .dout(n125));
  jnot g0077(.din(n125), .dout(n126));
  jand g0078(.dina(n126), .dinb(n124), .dout(n127));
  jand g0079(.dina(n127), .dinb(n120), .dout(n128));
  jand g0080(.dina(n128), .dinb(n110), .dout(n129));
  jnot g0081(.din(n129), .dout(n130));
  jor  g0082(.dina(n126), .dinb(n123), .dout(n131));
  jnot g0083(.din(n131), .dout(n132));
  jnot g0084(.din(n116), .dout(n133));
  jand g0085(.dina(n118), .dinb(n133), .dout(n134));
  jand g0086(.dina(n134), .dinb(n132), .dout(n135));
  jand g0087(.dina(n135), .dinb(n109), .dout(n136));
  jand g0088(.dina(n136), .dinb(n96), .dout(n137));
  jnot g0089(.din(n137), .dout(n138));
  jand g0090(.dina(n117), .dinb(n116), .dout(n139));
  jand g0091(.dina(n125), .dinb(n123), .dout(n140));
  jand g0092(.dina(n140), .dinb(n139), .dout(n141));
  jnot g0093(.din(n141), .dout(n142));
  jnot g0094(.din(n96), .dout(n143));
  jnot g0095(.din(n103), .dout(n144));
  jor  g0096(.dina(n108), .dinb(n144), .dout(n145));
  jor  g0097(.dina(n145), .dinb(n143), .dout(n146));
  jor  g0098(.dina(n146), .dinb(n142), .dout(n147));
  jand g0099(.dina(n147), .dinb(n138), .dout(n148));
  jand g0100(.dina(n148), .dinb(n130), .dout(n149));
  jnot g0101(.din(n149), .dout(n150));
  jand g0102(.dina(n109), .dinb(n143), .dout(n151));
  jand g0103(.dina(n151), .dinb(n128), .dout(n152));
  jnot g0104(.din(n152), .dout(n153));
  jor  g0105(.dina(n131), .dinb(n119), .dout(n154));
  jnot g0106(.din(n154), .dout(n155));
  jand g0107(.dina(n155), .dinb(n151), .dout(n156));
  jnot g0108(.din(n156), .dout(n157));
  jand g0109(.dina(n157), .dinb(n153), .dout(n158));
  jnot g0110(.din(n158), .dout(n159));
  jand g0111(.dina(n136), .dinb(n143), .dout(n160));
  jnot g0112(.din(n146), .dout(n161));
  jand g0113(.dina(n126), .dinb(n123), .dout(n162));
  jand g0114(.dina(n162), .dinb(n139), .dout(n163));
  jand g0115(.dina(n163), .dinb(n161), .dout(n164));
  jor  g0116(.dina(n164), .dinb(n160), .dout(n165));
  jor  g0117(.dina(n165), .dinb(n159), .dout(n166));
  jor  g0118(.dina(n166), .dinb(n150), .dout(n167));
  jnot g0119(.din(n167), .dout(n168));
  jnot g0120(.din(n104), .dout(n169));
  jnot g0121(.din(a20 ), .dout(n170));
  jnot g0122(.din(a19 ), .dout(n171));
  jnot g0123(.din(a18 ), .dout(n172));
  jnot g0124(.din(a16 ), .dout(n173));
  jnot g0125(.din(a15 ), .dout(n174));
  jnot g0126(.din(a14 ), .dout(n175));
  jnot g0127(.din(a13 ), .dout(n176));
  jnot g0128(.din(a12 ), .dout(n177));
  jnot g0129(.din(a11 ), .dout(n178));
  jnot g0130(.din(a10 ), .dout(n179));
  jnot g0131(.din(a9 ), .dout(n180));
  jnot g0132(.din(a8 ), .dout(n181));
  jnot g0133(.din(a7 ), .dout(n182));
  jnot g0134(.din(a6 ), .dout(n183));
  jnot g0135(.din(a5 ), .dout(n184));
  jnot g0136(.din(a4 ), .dout(n185));
  jnot g0137(.din(a3 ), .dout(n186));
  jnot g0138(.din(a2 ), .dout(n187));
  jand g0139(.dina(n187), .dinb(n62), .dout(n188));
  jand g0140(.dina(n188), .dinb(n61), .dout(n189));
  jand g0141(.dina(n189), .dinb(n186), .dout(n190));
  jand g0142(.dina(n190), .dinb(n185), .dout(n191));
  jand g0143(.dina(n191), .dinb(n184), .dout(n192));
  jand g0144(.dina(n192), .dinb(n183), .dout(n193));
  jand g0145(.dina(n193), .dinb(n182), .dout(n194));
  jand g0146(.dina(n194), .dinb(n181), .dout(n195));
  jand g0147(.dina(n195), .dinb(n180), .dout(n196));
  jand g0148(.dina(n196), .dinb(n179), .dout(n197));
  jand g0149(.dina(n197), .dinb(n178), .dout(n198));
  jand g0150(.dina(n198), .dinb(n177), .dout(n199));
  jand g0151(.dina(n199), .dinb(n176), .dout(n200));
  jand g0152(.dina(n200), .dinb(n175), .dout(n201));
  jand g0153(.dina(n201), .dinb(n174), .dout(n202));
  jand g0154(.dina(n202), .dinb(n173), .dout(n203));
  jand g0155(.dina(n203), .dinb(n121), .dout(n204));
  jand g0156(.dina(n204), .dinb(n172), .dout(n205));
  jand g0157(.dina(n205), .dinb(n171), .dout(n206));
  jand g0158(.dina(n206), .dinb(n170), .dout(n207));
  jor  g0159(.dina(n207), .dinb(a22 ), .dout(n208));
  jor  g0160(.dina(n105), .dinb(n208), .dout(n209));
  jand g0161(.dina(n209), .dinb(n169), .dout(n210));
  jand g0162(.dina(n210), .dinb(n103), .dout(n211));
  jand g0163(.dina(n211), .dinb(n143), .dout(n212));
  jand g0164(.dina(n212), .dinb(n163), .dout(n213));
  jnot g0165(.din(n213), .dout(n214));
  jor  g0166(.dina(n145), .dinb(n96), .dout(n215));
  jor  g0167(.dina(n215), .dinb(n142), .dout(n216));
  jand g0168(.dina(n216), .dinb(n214), .dout(n217));
  jand g0169(.dina(n217), .dinb(n168), .dout(n218));
  jand g0170(.dina(n118), .dinb(n116), .dout(n219));
  jand g0171(.dina(n219), .dinb(n132), .dout(n220));
  jand g0172(.dina(n220), .dinb(n151), .dout(n221));
  jnot g0173(.din(n221), .dout(n222));
  jand g0174(.dina(n140), .dinb(n120), .dout(n223));
  jand g0175(.dina(n223), .dinb(n212), .dout(n224));
  jnot g0176(.din(n224), .dout(n225));
  jand g0177(.dina(n225), .dinb(n222), .dout(n226));
  jand g0178(.dina(n219), .dinb(n162), .dout(n227));
  jand g0179(.dina(n227), .dinb(n151), .dout(n228));
  jnot g0180(.din(n228), .dout(n229));
  jand g0181(.dina(n219), .dinb(n127), .dout(n230));
  jand g0182(.dina(n230), .dinb(n110), .dout(n231));
  jnot g0183(.din(n231), .dout(n232));
  jand g0184(.dina(n232), .dinb(n229), .dout(n233));
  jand g0185(.dina(n233), .dinb(n226), .dout(n234));
  jand g0186(.dina(n220), .dinb(n110), .dout(n235));
  jand g0187(.dina(n162), .dinb(n120), .dout(n236));
  jand g0188(.dina(n236), .dinb(n211), .dout(n237));
  jor  g0189(.dina(n237), .dinb(n235), .dout(n238));
  jnot g0190(.din(n238), .dout(n239));
  jand g0191(.dina(n227), .dinb(n110), .dout(n240));
  jnot g0192(.din(n240), .dout(n241));
  jnot g0193(.din(n223), .dout(n242));
  jor  g0194(.dina(n242), .dinb(n146), .dout(n243));
  jand g0195(.dina(n243), .dinb(n241), .dout(n244));
  jand g0196(.dina(n244), .dinb(n239), .dout(n245));
  jand g0197(.dina(n245), .dinb(n234), .dout(n246));
  jand g0198(.dina(n140), .dinb(n134), .dout(n247));
  jand g0199(.dina(n247), .dinb(n151), .dout(n248));
  jnot g0200(.din(n248), .dout(n249));
  jand g0201(.dina(n141), .dinb(n110), .dout(n250));
  jnot g0202(.din(n250), .dout(n251));
  jand g0203(.dina(n251), .dinb(n249), .dout(n252));
  jand g0204(.dina(n223), .dinb(n110), .dout(n253));
  jnot g0205(.din(n253), .dout(n254));
  jand g0206(.dina(n151), .dinb(n141), .dout(n255));
  jnot g0207(.din(n255), .dout(n256));
  jand g0208(.dina(n256), .dinb(n254), .dout(n257));
  jand g0209(.dina(n257), .dinb(n252), .dout(n258));
  jand g0210(.dina(n162), .dinb(n134), .dout(n259));
  jand g0211(.dina(n259), .dinb(n151), .dout(n260));
  jnot g0212(.din(n260), .dout(n261));
  jand g0213(.dina(n139), .dinb(n132), .dout(n262));
  jand g0214(.dina(n262), .dinb(n161), .dout(n263));
  jnot g0215(.din(n263), .dout(n264));
  jand g0216(.dina(n264), .dinb(n261), .dout(n265));
  jand g0217(.dina(n259), .dinb(n110), .dout(n266));
  jnot g0218(.din(n266), .dout(n267));
  jand g0219(.dina(n139), .dinb(n127), .dout(n268));
  jand g0220(.dina(n268), .dinb(n151), .dout(n269));
  jnot g0221(.din(n269), .dout(n270));
  jand g0222(.dina(n270), .dinb(n267), .dout(n271));
  jand g0223(.dina(n271), .dinb(n265), .dout(n272));
  jand g0224(.dina(n272), .dinb(n258), .dout(n273));
  jand g0225(.dina(n273), .dinb(n246), .dout(n274));
  jand g0226(.dina(n274), .dinb(n218), .dout(n275));
  jnot g0227(.din(n230), .dout(n276));
  jor  g0228(.dina(n276), .dinb(n146), .dout(n277));
  jand g0229(.dina(n220), .dinb(n212), .dout(n278));
  jnot g0230(.din(n278), .dout(n279));
  jand g0231(.dina(n279), .dinb(n277), .dout(n280));
  jnot g0232(.din(n220), .dout(n281));
  jor  g0233(.dina(n281), .dinb(n146), .dout(n282));
  jand g0234(.dina(n219), .dinb(n140), .dout(n283));
  jand g0235(.dina(n283), .dinb(n110), .dout(n284));
  jnot g0236(.din(n284), .dout(n285));
  jand g0237(.dina(n285), .dinb(n282), .dout(n286));
  jand g0238(.dina(n286), .dinb(n280), .dout(n287));
  jand g0239(.dina(n211), .dinb(n128), .dout(n288));
  jnot g0240(.din(n288), .dout(n289));
  jand g0241(.dina(n283), .dinb(n151), .dout(n290));
  jnot g0242(.din(n290), .dout(n291));
  jand g0243(.dina(n291), .dinb(n289), .dout(n292));
  jand g0244(.dina(n236), .dinb(n110), .dout(n293));
  jnot g0245(.din(n293), .dout(n294));
  jor  g0246(.dina(n154), .dinb(n146), .dout(n295));
  jand g0247(.dina(n295), .dinb(n294), .dout(n296));
  jand g0248(.dina(n296), .dinb(n292), .dout(n297));
  jand g0249(.dina(n223), .dinb(n151), .dout(n298));
  jand g0250(.dina(n230), .dinb(n151), .dout(n299));
  jor  g0251(.dina(n299), .dinb(n298), .dout(n300));
  jnot g0252(.din(n300), .dout(n301));
  jand g0253(.dina(n236), .dinb(n151), .dout(n302));
  jnot g0254(.din(n302), .dout(n303));
  jor  g0255(.dina(n215), .dinb(n154), .dout(n304));
  jand g0256(.dina(n304), .dinb(n303), .dout(n305));
  jand g0257(.dina(n305), .dinb(n301), .dout(n306));
  jand g0258(.dina(n306), .dinb(n297), .dout(n307));
  jand g0259(.dina(n307), .dinb(n287), .dout(n308));
  jand g0260(.dina(n262), .dinb(n212), .dout(n309));
  jnot g0261(.din(n309), .dout(n310));
  jand g0262(.dina(n155), .dinb(n110), .dout(n311));
  jnot g0263(.din(n311), .dout(n312));
  jnot g0264(.din(n268), .dout(n313));
  jor  g0265(.dina(n313), .dinb(n145), .dout(n314));
  jand g0266(.dina(n163), .dinb(n109), .dout(n315));
  jnot g0267(.din(n315), .dout(n316));
  jand g0268(.dina(n316), .dinb(n314), .dout(n317));
  jand g0269(.dina(n317), .dinb(n312), .dout(n318));
  jand g0270(.dina(n318), .dinb(n310), .dout(n319));
  jand g0271(.dina(n268), .dinb(n110), .dout(n320));
  jnot g0272(.din(n320), .dout(n321));
  jand g0273(.dina(n247), .dinb(n110), .dout(n322));
  jnot g0274(.din(n322), .dout(n323));
  jand g0275(.dina(n323), .dinb(n321), .dout(n324));
  jnot g0276(.din(n109), .dout(n325));
  jnot g0277(.din(n262), .dout(n326));
  jand g0278(.dina(n134), .dinb(n127), .dout(n327));
  jnot g0279(.din(n327), .dout(n328));
  jand g0280(.dina(n328), .dinb(n326), .dout(n329));
  jor  g0281(.dina(n329), .dinb(n325), .dout(n330));
  jand g0282(.dina(n330), .dinb(n324), .dout(n331));
  jand g0283(.dina(n331), .dinb(n319), .dout(n332));
  jand g0284(.dina(n332), .dinb(n308), .dout(n333));
  jand g0285(.dina(n333), .dinb(n275), .dout(n334));
  jnot g0286(.din(n334), .dout(n335));
  jand g0287(.dina(n82), .dinb(n49), .dout(n336));
  jxor g0288(.dina(n336), .dinb(a7 ), .dout(n337));
  jand g0289(.dina(n337), .dinb(n335), .dout(n338));
  jor  g0290(.dina(n108), .dinb(n103), .dout(n339));
  jor  g0291(.dina(n339), .dinb(n96), .dout(n340));
  jnot g0292(.din(n340), .dout(n341));
  jand g0293(.dina(n341), .dinb(n236), .dout(n342));
  jnot g0294(.din(n342), .dout(n343));
  jand g0295(.dina(n343), .dinb(n303), .dout(n344));
  jand g0296(.dina(n108), .dinb(n144), .dout(n345));
  jand g0297(.dina(n345), .dinb(n143), .dout(n346));
  jand g0298(.dina(n346), .dinb(n223), .dout(n347));
  jnot g0299(.din(n347), .dout(n348));
  jand g0300(.dina(n345), .dinb(n96), .dout(n349));
  jand g0301(.dina(n349), .dinb(n247), .dout(n350));
  jnot g0302(.din(n350), .dout(n351));
  jand g0303(.dina(n351), .dinb(n348), .dout(n352));
  jand g0304(.dina(n210), .dinb(n144), .dout(n353));
  jand g0305(.dina(n353), .dinb(n96), .dout(n354));
  jand g0306(.dina(n354), .dinb(n268), .dout(n355));
  jnot g0307(.din(n355), .dout(n356));
  jand g0308(.dina(n346), .dinb(n230), .dout(n357));
  jnot g0309(.din(n357), .dout(n358));
  jand g0310(.dina(n358), .dinb(n356), .dout(n359));
  jand g0311(.dina(n359), .dinb(n352), .dout(n360));
  jand g0312(.dina(n360), .dinb(n344), .dout(n361));
  jand g0313(.dina(n349), .dinb(n327), .dout(n362));
  jnot g0314(.din(n362), .dout(n363));
  jand g0315(.dina(n349), .dinb(n163), .dout(n364));
  jnot g0316(.din(n364), .dout(n365));
  jand g0317(.dina(n365), .dinb(n363), .dout(n366));
  jor  g0318(.dina(n339), .dinb(n143), .dout(n367));
  jor  g0319(.dina(n367), .dinb(n328), .dout(n368));
  jand g0320(.dina(n341), .dinb(n268), .dout(n369));
  jnot g0321(.din(n369), .dout(n370));
  jand g0322(.dina(n370), .dinb(n368), .dout(n371));
  jnot g0323(.din(n298), .dout(n372));
  jand g0324(.dina(n349), .dinb(n220), .dout(n373));
  jnot g0325(.din(n373), .dout(n374));
  jand g0326(.dina(n374), .dinb(n372), .dout(n375));
  jand g0327(.dina(n375), .dinb(n371), .dout(n376));
  jand g0328(.dina(n376), .dinb(n366), .dout(n377));
  jand g0329(.dina(n349), .dinb(n259), .dout(n378));
  jnot g0330(.din(n378), .dout(n379));
  jnot g0331(.din(n227), .dout(n380));
  jor  g0332(.dina(n380), .dinb(n146), .dout(n381));
  jnot g0333(.din(n283), .dout(n382));
  jor  g0334(.dina(n382), .dinb(n146), .dout(n383));
  jand g0335(.dina(n383), .dinb(n381), .dout(n384));
  jand g0336(.dina(n384), .dinb(n379), .dout(n385));
  jand g0337(.dina(n354), .dinb(n247), .dout(n386));
  jnot g0338(.din(n386), .dout(n387));
  jand g0339(.dina(n387), .dinb(n295), .dout(n388));
  jand g0340(.dina(n346), .dinb(n128), .dout(n389));
  jnot g0341(.din(n389), .dout(n390));
  jand g0342(.dina(n390), .dinb(n243), .dout(n391));
  jand g0343(.dina(n391), .dinb(n388), .dout(n392));
  jand g0344(.dina(n392), .dinb(n385), .dout(n393));
  jand g0345(.dina(n393), .dinb(n377), .dout(n394));
  jand g0346(.dina(n394), .dinb(n361), .dout(n395));
  jand g0347(.dina(n288), .dinb(n143), .dout(n396));
  jnot g0348(.din(n396), .dout(n397));
  jand g0349(.dina(n397), .dinb(n214), .dout(n398));
  jand g0350(.dina(n294), .dinb(n222), .dout(n399));
  jand g0351(.dina(n346), .dinb(n283), .dout(n400));
  jnot g0352(.din(n400), .dout(n401));
  jor  g0353(.dina(n276), .dinb(n215), .dout(n402));
  jand g0354(.dina(n402), .dinb(n401), .dout(n403));
  jand g0355(.dina(n403), .dinb(n399), .dout(n404));
  jand g0356(.dina(n404), .dinb(n398), .dout(n405));
  jand g0357(.dina(n341), .dinb(n220), .dout(n406));
  jor  g0358(.dina(n406), .dinb(n160), .dout(n407));
  jnot g0359(.din(n407), .dout(n408));
  jnot g0360(.din(n236), .dout(n409));
  jor  g0361(.dina(n409), .dinb(n215), .dout(n410));
  jand g0362(.dina(n346), .dinb(n268), .dout(n411));
  jnot g0363(.din(n411), .dout(n412));
  jand g0364(.dina(n412), .dinb(n410), .dout(n413));
  jand g0365(.dina(n354), .dinb(n230), .dout(n414));
  jand g0366(.dina(n349), .dinb(n236), .dout(n415));
  jor  g0367(.dina(n415), .dinb(n414), .dout(n416));
  jnot g0368(.din(n416), .dout(n417));
  jand g0369(.dina(n417), .dinb(n413), .dout(n418));
  jand g0370(.dina(n418), .dinb(n408), .dout(n419));
  jor  g0371(.dina(n380), .dinb(n215), .dout(n420));
  jor  g0372(.dina(n367), .dinb(n382), .dout(n421));
  jor  g0373(.dina(n367), .dinb(n380), .dout(n422));
  jand g0374(.dina(n422), .dinb(n421), .dout(n423));
  jand g0375(.dina(n423), .dinb(n420), .dout(n424));
  jand g0376(.dina(n349), .dinb(n262), .dout(n425));
  jnot g0377(.din(n425), .dout(n426));
  jor  g0378(.dina(n340), .dinb(n142), .dout(n427));
  jand g0379(.dina(n427), .dinb(n426), .dout(n428));
  jand g0380(.dina(n341), .dinb(n223), .dout(n429));
  jnot g0381(.din(n429), .dout(n430));
  jand g0382(.dina(n430), .dinb(n428), .dout(n431));
  jand g0383(.dina(n431), .dinb(n424), .dout(n432));
  jand g0384(.dina(n432), .dinb(n419), .dout(n433));
  jand g0385(.dina(n433), .dinb(n405), .dout(n434));
  jnot g0386(.din(n247), .dout(n435));
  jor  g0387(.dina(n435), .dinb(n215), .dout(n436));
  jor  g0388(.dina(n328), .dinb(n146), .dout(n437));
  jand g0389(.dina(n437), .dinb(n436), .dout(n438));
  jand g0390(.dina(n438), .dinb(n147), .dout(n439));
  jand g0391(.dina(n349), .dinb(n230), .dout(n440));
  jnot g0392(.din(n440), .dout(n441));
  jand g0393(.dina(n441), .dinb(n267), .dout(n442));
  jand g0394(.dina(n442), .dinb(n241), .dout(n443));
  jand g0395(.dina(n354), .dinb(n135), .dout(n444));
  jnot g0396(.din(n444), .dout(n445));
  jand g0397(.dina(n314), .dinb(n229), .dout(n446));
  jand g0398(.dina(n446), .dinb(n445), .dout(n447));
  jand g0399(.dina(n447), .dinb(n443), .dout(n448));
  jand g0400(.dina(n448), .dinb(n439), .dout(n449));
  jand g0401(.dina(n346), .dinb(n227), .dout(n450));
  jnot g0402(.din(n450), .dout(n451));
  jand g0403(.dina(n451), .dinb(n261), .dout(n452));
  jand g0404(.dina(n346), .dinb(n141), .dout(n453));
  jnot g0405(.din(n453), .dout(n454));
  jand g0406(.dina(n454), .dinb(n138), .dout(n455));
  jand g0407(.dina(n455), .dinb(n452), .dout(n456));
  jnot g0408(.din(n259), .dout(n457));
  jor  g0409(.dina(n367), .dinb(n457), .dout(n458));
  jand g0410(.dina(n458), .dinb(n249), .dout(n459));
  jand g0411(.dina(n341), .dinb(n128), .dout(n460));
  jnot g0412(.din(n460), .dout(n461));
  jnot g0413(.din(n163), .dout(n462));
  jor  g0414(.dina(n340), .dinb(n462), .dout(n463));
  jand g0415(.dina(n463), .dinb(n461), .dout(n464));
  jand g0416(.dina(n464), .dinb(n459), .dout(n465));
  jand g0417(.dina(n465), .dinb(n456), .dout(n466));
  jnot g0418(.din(n235), .dout(n467));
  jand g0419(.dina(n353), .dinb(n155), .dout(n468));
  jand g0420(.dina(n468), .dinb(n143), .dout(n469));
  jnot g0421(.din(n469), .dout(n470));
  jand g0422(.dina(n470), .dinb(n467), .dout(n471));
  jand g0423(.dina(n354), .dinb(n262), .dout(n472));
  jnot g0424(.din(n472), .dout(n473));
  jand g0425(.dina(n473), .dinb(n282), .dout(n474));
  jand g0426(.dina(n345), .dinb(n155), .dout(n475));
  jand g0427(.dina(n475), .dinb(n96), .dout(n476));
  jnot g0428(.din(n476), .dout(n477));
  jand g0429(.dina(n346), .dinb(n135), .dout(n478));
  jnot g0430(.din(n478), .dout(n479));
  jand g0431(.dina(n479), .dinb(n477), .dout(n480));
  jand g0432(.dina(n480), .dinb(n474), .dout(n481));
  jand g0433(.dina(n481), .dinb(n471), .dout(n482));
  jand g0434(.dina(n482), .dinb(n466), .dout(n483));
  jand g0435(.dina(n483), .dinb(n449), .dout(n484));
  jand g0436(.dina(n484), .dinb(n434), .dout(n485));
  jand g0437(.dina(n485), .dinb(n395), .dout(n486));
  jand g0438(.dina(n327), .dinb(n110), .dout(n487));
  jnot g0439(.din(n487), .dout(n488));
  jand g0440(.dina(n488), .dinb(n277), .dout(n489));
  jand g0441(.dina(n489), .dinb(n270), .dout(n490));
  jand g0442(.dina(n346), .dinb(n236), .dout(n491));
  jor  g0443(.dina(n491), .dinb(n478), .dout(n492));
  jnot g0444(.din(n492), .dout(n493));
  jand g0445(.dina(n426), .dinb(n310), .dout(n494));
  jand g0446(.dina(n494), .dinb(n286), .dout(n495));
  jand g0447(.dina(n495), .dinb(n493), .dout(n496));
  jand g0448(.dina(n496), .dinb(n490), .dout(n497));
  jnot g0449(.din(n497), .dout(n498));
  jnot g0450(.din(n406), .dout(n499));
  jor  g0451(.dina(n339), .dinb(n154), .dout(n500));
  jor  g0452(.dina(n500), .dinb(n143), .dout(n501));
  jand g0453(.dina(n501), .dinb(n368), .dout(n502));
  jand g0454(.dina(n502), .dinb(n499), .dout(n503));
  jand g0455(.dina(n412), .dinb(n256), .dout(n504));
  jand g0456(.dina(n259), .dinb(n161), .dout(n505));
  jnot g0457(.din(n505), .dout(n506));
  jand g0458(.dina(n506), .dinb(n454), .dout(n507));
  jand g0459(.dina(n507), .dinb(n504), .dout(n508));
  jand g0460(.dina(n508), .dinb(n503), .dout(n509));
  jnot g0461(.din(n509), .dout(n510));
  jand g0462(.dina(n463), .dinb(n304), .dout(n511));
  jand g0463(.dina(n511), .dinb(n397), .dout(n512));
  jand g0464(.dina(n512), .dinb(n459), .dout(n513));
  jnot g0465(.din(n513), .dout(n514));
  jor  g0466(.dina(n367), .dinb(n281), .dout(n515));
  jand g0467(.dina(n515), .dinb(n374), .dout(n516));
  jnot g0468(.din(n516), .dout(n517));
  jand g0469(.dina(n262), .dinb(n151), .dout(n518));
  jor  g0470(.dina(n518), .dinb(n164), .dout(n519));
  jor  g0471(.dina(n519), .dinb(n517), .dout(n520));
  jand g0472(.dina(n346), .dinb(n163), .dout(n521));
  jor  g0473(.dina(n521), .dinb(n440), .dout(n522));
  jnot g0474(.din(n522), .dout(n523));
  jand g0475(.dina(n351), .dinb(n157), .dout(n524));
  jand g0476(.dina(n524), .dinb(n523), .dout(n525));
  jnot g0477(.din(n525), .dout(n526));
  jor  g0478(.dina(n526), .dinb(n520), .dout(n527));
  jor  g0479(.dina(n527), .dinb(n514), .dout(n528));
  jor  g0480(.dina(n528), .dinb(n510), .dout(n529));
  jor  g0481(.dina(n529), .dinb(n498), .dout(n530));
  jand g0482(.dina(n341), .dinb(n262), .dout(n531));
  jnot g0483(.din(n531), .dout(n532));
  jand g0484(.dina(n532), .dinb(n390), .dout(n533));
  jand g0485(.dina(n341), .dinb(n135), .dout(n534));
  jnot g0486(.din(n534), .dout(n535));
  jand g0487(.dina(n535), .dinb(n130), .dout(n536));
  jand g0488(.dina(n536), .dinb(n533), .dout(n537));
  jand g0489(.dina(n537), .dinb(n239), .dout(n538));
  jnot g0490(.din(n538), .dout(n539));
  jand g0491(.dina(n401), .dinb(n138), .dout(n540));
  jand g0492(.dina(n540), .dinb(n225), .dout(n541));
  jnot g0493(.din(n541), .dout(n542));
  jand g0494(.dina(n348), .dinb(n251), .dout(n543));
  jnot g0495(.din(n543), .dout(n544));
  jor  g0496(.dina(n298), .dinb(n278), .dout(n545));
  jor  g0497(.dina(n545), .dinb(n544), .dout(n546));
  jor  g0498(.dina(n546), .dinb(n542), .dout(n547));
  jand g0499(.dina(n349), .dinb(n135), .dout(n548));
  jor  g0500(.dina(n548), .dinb(n444), .dout(n549));
  jor  g0501(.dina(n549), .dinb(n472), .dout(n550));
  jand g0502(.dina(n327), .dinb(n212), .dout(n551));
  jand g0503(.dina(n354), .dinb(n236), .dout(n552));
  jor  g0504(.dina(n552), .dinb(n551), .dout(n553));
  jand g0505(.dina(n346), .dinb(n262), .dout(n554));
  jor  g0506(.dina(n554), .dinb(n429), .dout(n555));
  jor  g0507(.dina(n555), .dinb(n553), .dout(n556));
  jor  g0508(.dina(n556), .dinb(n550), .dout(n557));
  jor  g0509(.dina(n557), .dinb(n547), .dout(n558));
  jor  g0510(.dina(n558), .dinb(n539), .dout(n559));
  jand g0511(.dina(n262), .dinb(n110), .dout(n560));
  jnot g0512(.din(n560), .dout(n561));
  jand g0513(.dina(n475), .dinb(n143), .dout(n562));
  jnot g0514(.din(n562), .dout(n563));
  jand g0515(.dina(n563), .dinb(n561), .dout(n564));
  jand g0516(.dina(n564), .dinb(n356), .dout(n565));
  jnot g0517(.din(n565), .dout(n566));
  jand g0518(.dina(n381), .dinb(n232), .dout(n567));
  jand g0519(.dina(n567), .dinb(n295), .dout(n568));
  jnot g0520(.din(n568), .dout(n569));
  jor  g0521(.dina(n342), .dinb(n320), .dout(n570));
  jor  g0522(.dina(n570), .dinb(n240), .dout(n571));
  jor  g0523(.dina(n571), .dinb(n569), .dout(n572));
  jor  g0524(.dina(n572), .dinb(n566), .dout(n573));
  jand g0525(.dina(n354), .dinb(n163), .dout(n574));
  jor  g0526(.dina(n574), .dinb(n266), .dout(n575));
  jor  g0527(.dina(n575), .dinb(n386), .dout(n576));
  jnot g0528(.din(n420), .dout(n577));
  jor  g0529(.dina(n577), .dinb(n213), .dout(n578));
  jor  g0530(.dina(n314), .dinb(n143), .dout(n579));
  jnot g0531(.din(n579), .dout(n580));
  jand g0532(.dina(n288), .dinb(n96), .dout(n581));
  jor  g0533(.dina(n581), .dinb(n580), .dout(n582));
  jor  g0534(.dina(n582), .dinb(n578), .dout(n583));
  jor  g0535(.dina(n583), .dinb(n576), .dout(n584));
  jnot g0536(.din(n437), .dout(n585));
  jand g0537(.dina(n341), .dinb(n327), .dout(n586));
  jor  g0538(.dina(n586), .dinb(n585), .dout(n587));
  jand g0539(.dina(n341), .dinb(n247), .dout(n588));
  jor  g0540(.dina(n588), .dinb(n263), .dout(n589));
  jor  g0541(.dina(n589), .dinb(n587), .dout(n590));
  jand g0542(.dina(n349), .dinb(n227), .dout(n591));
  jnot g0543(.din(n591), .dout(n592));
  jand g0544(.dina(n346), .dinb(n247), .dout(n593));
  jnot g0545(.din(n593), .dout(n594));
  jand g0546(.dina(n594), .dinb(n592), .dout(n595));
  jor  g0547(.dina(n340), .dinb(n457), .dout(n596));
  jand g0548(.dina(n596), .dinb(n243), .dout(n597));
  jand g0549(.dina(n597), .dinb(n595), .dout(n598));
  jnot g0550(.din(n598), .dout(n599));
  jor  g0551(.dina(n599), .dinb(n590), .dout(n600));
  jor  g0552(.dina(n600), .dinb(n584), .dout(n601));
  jor  g0553(.dina(n601), .dinb(n573), .dout(n602));
  jor  g0554(.dina(n602), .dinb(n559), .dout(n603));
  jor  g0555(.dina(n603), .dinb(n530), .dout(n604));
  jnot g0556(.din(n556), .dout(n605));
  jand g0557(.dina(n349), .dinb(n141), .dout(n606));
  jor  g0558(.dina(n606), .dinb(n518), .dout(n607));
  jand g0559(.dina(n315), .dinb(n143), .dout(n608));
  jor  g0560(.dina(n608), .dinb(n269), .dout(n609));
  jor  g0561(.dina(n609), .dinb(n607), .dout(n610));
  jnot g0562(.din(n610), .dout(n611));
  jor  g0563(.dina(n367), .dinb(n242), .dout(n612));
  jand g0564(.dina(n327), .dinb(n151), .dout(n613));
  jnot g0565(.din(n613), .dout(n614));
  jand g0566(.dina(n614), .dinb(n612), .dout(n615));
  jand g0567(.dina(n615), .dinb(n232), .dout(n616));
  jand g0568(.dina(n616), .dinb(n611), .dout(n617));
  jand g0569(.dina(n617), .dinb(n605), .dout(n618));
  jand g0570(.dina(n249), .dinb(n229), .dout(n619));
  jand g0571(.dina(n561), .dinb(n216), .dout(n620));
  jand g0572(.dina(n620), .dinb(n294), .dout(n621));
  jand g0573(.dina(n621), .dinb(n619), .dout(n622));
  jand g0574(.dina(n379), .dinb(n251), .dout(n623));
  jor  g0575(.dina(n314), .dinb(n96), .dout(n624));
  jand g0576(.dina(n624), .dinb(n454), .dout(n625));
  jand g0577(.dina(n436), .dinb(n264), .dout(n626));
  jand g0578(.dina(n626), .dinb(n625), .dout(n627));
  jand g0579(.dina(n627), .dinb(n623), .dout(n628));
  jand g0580(.dina(n628), .dinb(n622), .dout(n629));
  jand g0581(.dina(n629), .dinb(n618), .dout(n630));
  jand g0582(.dina(n315), .dinb(n96), .dout(n631));
  jnot g0583(.din(n631), .dout(n632));
  jand g0584(.dina(n632), .dinb(n303), .dout(n633));
  jand g0585(.dina(n499), .dinb(n343), .dout(n634));
  jand g0586(.dina(n634), .dinb(n633), .dout(n635));
  jand g0587(.dina(n635), .dinb(n630), .dout(n636));
  jor  g0588(.dina(n487), .dinb(n240), .dout(n637));
  jnot g0589(.din(n637), .dout(n638));
  jand g0590(.dina(n515), .dinb(n312), .dout(n639));
  jand g0591(.dina(n639), .dinb(n638), .dout(n640));
  jand g0592(.dina(n283), .dinb(n212), .dout(n641));
  jnot g0593(.din(n641), .dout(n642));
  jand g0594(.dina(n642), .dinb(n402), .dout(n643));
  jand g0595(.dina(n346), .dinb(n259), .dout(n644));
  jnot g0596(.din(n644), .dout(n645));
  jand g0597(.dina(n645), .dinb(n356), .dout(n646));
  jand g0598(.dina(n646), .dinb(n643), .dout(n647));
  jand g0599(.dina(n647), .dinb(n640), .dout(n648));
  jnot g0600(.din(n304), .dout(n649));
  jor  g0601(.dina(n562), .dinb(n440), .dout(n650));
  jor  g0602(.dina(n650), .dinb(n649), .dout(n651));
  jnot g0603(.din(n381), .dout(n652));
  jor  g0604(.dina(n469), .dinb(n652), .dout(n653));
  jor  g0605(.dina(n653), .dinb(n651), .dout(n654));
  jnot g0606(.din(n654), .dout(n655));
  jand g0607(.dina(n532), .dinb(n348), .dout(n656));
  jand g0608(.dina(n656), .dinb(n225), .dout(n657));
  jand g0609(.dina(n657), .dinb(n301), .dout(n658));
  jand g0610(.dina(n658), .dinb(n655), .dout(n659));
  jand g0611(.dina(n659), .dinb(n648), .dout(n660));
  jand g0612(.dina(n349), .dinb(n223), .dout(n661));
  jnot g0613(.din(n661), .dout(n662));
  jnot g0614(.din(n135), .dout(n663));
  jor  g0615(.dina(n145), .dinb(n663), .dout(n664));
  jor  g0616(.dina(n664), .dinb(n143), .dout(n665));
  jand g0617(.dina(n665), .dinb(n662), .dout(n666));
  jand g0618(.dina(n666), .dinb(n477), .dout(n667));
  jnot g0619(.din(n548), .dout(n668));
  jand g0620(.dina(n668), .dinb(n451), .dout(n669));
  jand g0621(.dina(n346), .dinb(n220), .dout(n670));
  jor  g0622(.dina(n670), .dinb(n320), .dout(n671));
  jnot g0623(.din(n671), .dout(n672));
  jand g0624(.dina(n672), .dinb(n398), .dout(n673));
  jand g0625(.dina(n673), .dinb(n669), .dout(n674));
  jand g0626(.dina(n674), .dinb(n667), .dout(n675));
  jand g0627(.dina(n579), .dinb(n410), .dout(n676));
  jand g0628(.dina(n676), .dinb(n461), .dout(n677));
  jand g0629(.dina(n354), .dinb(n128), .dout(n678));
  jnot g0630(.din(n678), .dout(n679));
  jand g0631(.dina(n679), .dinb(n473), .dout(n680));
  jand g0632(.dina(n506), .dinb(n256), .dout(n681));
  jand g0633(.dina(n479), .dinb(n279), .dout(n682));
  jand g0634(.dina(n682), .dinb(n681), .dout(n683));
  jand g0635(.dina(n683), .dinb(n680), .dout(n684));
  jand g0636(.dina(n684), .dinb(n677), .dout(n685));
  jand g0637(.dina(n685), .dinb(n675), .dout(n686));
  jand g0638(.dina(n686), .dinb(n660), .dout(n687));
  jand g0639(.dina(n687), .dinb(n636), .dout(n688));
  jnot g0640(.din(n688), .dout(n689));
  jand g0641(.dina(n689), .dinb(n604), .dout(n690));
  jor  g0642(.dina(n690), .dinb(n486), .dout(n691));
  jand g0643(.dina(n691), .dinb(n338), .dout(n692));
  jxor g0644(.dina(n691), .dinb(n338), .dout(n693));
  jand g0645(.dina(a22 ), .dinb(a8 ), .dout(n694));
  jand g0646(.dina(n84), .dinb(n49), .dout(n695));
  jand g0647(.dina(n83), .dinb(a8 ), .dout(n696));
  jnot g0648(.din(n696), .dout(n697));
  jand g0649(.dina(n697), .dinb(n695), .dout(n698));
  jor  g0650(.dina(n698), .dinb(n694), .dout(n699));
  jand g0651(.dina(n699), .dinb(n335), .dout(n700));
  jand g0652(.dina(n700), .dinb(n693), .dout(n701));
  jor  g0653(.dina(n701), .dinb(n692), .dout(n702));
  jand g0654(.dina(a22 ), .dinb(a10 ), .dout(n703));
  jand g0655(.dina(n86), .dinb(n49), .dout(n704));
  jand g0656(.dina(n85), .dinb(a10 ), .dout(n705));
  jnot g0657(.din(n705), .dout(n706));
  jand g0658(.dina(n706), .dinb(n704), .dout(n707));
  jor  g0659(.dina(n707), .dinb(n703), .dout(n708));
  jnot g0660(.din(n574), .dout(n709));
  jor  g0661(.dina(n367), .dinb(n142), .dout(n710));
  jand g0662(.dina(n710), .dinb(n709), .dout(n711));
  jand g0663(.dina(n642), .dinb(n420), .dout(n712));
  jand g0664(.dina(n532), .dinb(n427), .dout(n713));
  jand g0665(.dina(n713), .dinb(n712), .dout(n714));
  jand g0666(.dina(n714), .dinb(n711), .dout(n715));
  jand g0667(.dina(n473), .dinb(n370), .dout(n716));
  jand g0668(.dina(n716), .dinb(n646), .dout(n717));
  jand g0669(.dina(n717), .dinb(n385), .dout(n718));
  jand g0670(.dina(n718), .dinb(n715), .dout(n719));
  jand g0671(.dina(n500), .dinb(n463), .dout(n720));
  jand g0672(.dina(n720), .dinb(n679), .dout(n721));
  jand g0673(.dina(n721), .dinb(n719), .dout(n722));
  jand g0674(.dina(n259), .dinb(n212), .dout(n723));
  jnot g0675(.din(n723), .dout(n724));
  jand g0676(.dina(n211), .dinb(n135), .dout(n725));
  jand g0677(.dina(n725), .dinb(n96), .dout(n726));
  jor  g0678(.dina(n726), .dinb(n551), .dout(n727));
  jnot g0679(.din(n727), .dout(n728));
  jand g0680(.dina(n728), .dinb(n724), .dout(n729));
  jnot g0681(.din(n554), .dout(n730));
  jand g0682(.dina(n730), .dinb(n402), .dout(n731));
  jor  g0683(.dina(n435), .dinb(n146), .dout(n732));
  jand g0684(.dina(n732), .dinb(n437), .dout(n733));
  jnot g0685(.din(n521), .dout(n734));
  jand g0686(.dina(n734), .dinb(n506), .dout(n735));
  jand g0687(.dina(n735), .dinb(n733), .dout(n736));
  jand g0688(.dina(n736), .dinb(n731), .dout(n737));
  jand g0689(.dina(n737), .dinb(n729), .dout(n738));
  jnot g0690(.din(n606), .dout(n739));
  jand g0691(.dina(n739), .dinb(n365), .dout(n740));
  jand g0692(.dina(n740), .dinb(n454), .dout(n741));
  jnot g0693(.din(n475), .dout(n742));
  jand g0694(.dina(n349), .dinb(n268), .dout(n743));
  jnot g0695(.din(n743), .dout(n744));
  jand g0696(.dina(n744), .dinb(n742), .dout(n745));
  jand g0697(.dina(n745), .dinb(n741), .dout(n746));
  jand g0698(.dina(n436), .dinb(n412), .dout(n747));
  jand g0699(.dina(n725), .dinb(n143), .dout(n748));
  jnot g0700(.din(n748), .dout(n749));
  jand g0701(.dina(n349), .dinb(n128), .dout(n750));
  jnot g0702(.din(n750), .dout(n751));
  jand g0703(.dina(n751), .dinb(n426), .dout(n752));
  jand g0704(.dina(n752), .dinb(n749), .dout(n753));
  jand g0705(.dina(n753), .dinb(n747), .dout(n754));
  jand g0706(.dina(n754), .dinb(n746), .dout(n755));
  jand g0707(.dina(n755), .dinb(n738), .dout(n756));
  jnot g0708(.din(n552), .dout(n757));
  jand g0709(.dina(n612), .dinb(n757), .dout(n758));
  jand g0710(.dina(n461), .dinb(n430), .dout(n759));
  jand g0711(.dina(n759), .dinb(n758), .dout(n760));
  jand g0712(.dina(n760), .dinb(n756), .dout(n761));
  jand g0713(.dina(n761), .dinb(n722), .dout(n762));
  jnot g0714(.din(n670), .dout(n763));
  jand g0715(.dina(n349), .dinb(n283), .dout(n764));
  jnot g0716(.din(n764), .dout(n765));
  jand g0717(.dina(n765), .dinb(n763), .dout(n766));
  jand g0718(.dina(n766), .dinb(n358), .dout(n767));
  jnot g0719(.din(n415), .dout(n768));
  jand g0720(.dina(n662), .dinb(n441), .dout(n769));
  jand g0721(.dina(n769), .dinb(n768), .dout(n770));
  jand g0722(.dina(n390), .dinb(n374), .dout(n771));
  jnot g0723(.din(n491), .dout(n772));
  jand g0724(.dina(n772), .dinb(n348), .dout(n773));
  jand g0725(.dina(n773), .dinb(n771), .dout(n774));
  jand g0726(.dina(n774), .dinb(n770), .dout(n775));
  jand g0727(.dina(n775), .dinb(n767), .dout(n776));
  jand g0728(.dina(n712), .dinb(n384), .dout(n777));
  jand g0729(.dina(n777), .dinb(n776), .dout(n778));
  jand g0730(.dina(n778), .dinb(n756), .dout(n779));
  jand g0731(.dina(n346), .dinb(n327), .dout(n780));
  jnot g0732(.din(n780), .dout(n781));
  jand g0733(.dina(n781), .dinb(n479), .dout(n782));
  jand g0734(.dina(n782), .dinb(n351), .dout(n783));
  jand g0735(.dina(n783), .dinb(n595), .dout(n784));
  jand g0736(.dina(n669), .dinb(n363), .dout(n785));
  jand g0737(.dina(n785), .dinb(n784), .dout(n786));
  jand g0738(.dina(n786), .dinb(n401), .dout(n787));
  jand g0739(.dina(n787), .dinb(n779), .dout(n788));
  jxor g0740(.dina(n788), .dinb(n762), .dout(n789));
  jnot g0741(.din(n762), .dout(n790));
  jor  g0742(.dina(n790), .dinb(n789), .dout(n792));
  jand g0743(.dina(n792), .dinb(n708), .dout(n793));
  jnot g0744(.din(n708), .dout(n794));
  jnot g0745(.din(n789), .dout(n795));
  jor  g0746(.dina(n788), .dinb(n762), .dout(n796));
  jand g0747(.dina(n334), .dinb(n795), .dout(n799));
  jnot g0748(.din(n799), .dout(n800));
  jand g0749(.dina(n800), .dinb(n794), .dout(n801));
  jor  g0750(.dina(n801), .dinb(n793), .dout(n802));
  jxor g0751(.dina(n704), .dinb(a11 ), .dout(n803));
  jand g0752(.dina(n788), .dinb(n762), .dout(n804));
  jnot g0753(.din(n803), .dout(n808));
  jand g0754(.dina(n789), .dinb(n808), .dout(n810));
  jnot g0755(.din(n810), .dout(n812));
  jand g0756(.dina(n812), .dinb(n802), .dout(n813));
  jand g0757(.dina(n813), .dinb(n702), .dout(n814));
  jand g0758(.dina(a22 ), .dinb(a14 ), .dout(n815));
  jnot g0759(.din(n815), .dout(n816));
  jand g0760(.dina(n89), .dinb(a14 ), .dout(n817));
  jor  g0761(.dina(n817), .dinb(a22 ), .dout(n818));
  jor  g0762(.dina(n818), .dinb(n201), .dout(n819));
  jand g0763(.dina(n819), .dinb(n816), .dout(n820));
  jand g0764(.dina(n744), .dinb(n401), .dout(n821));
  jand g0765(.dina(n515), .dinb(n321), .dout(n822));
  jand g0766(.dina(n822), .dinb(n821), .dout(n823));
  jand g0767(.dina(n823), .dinb(n158), .dout(n824));
  jnot g0768(.din(n414), .dout(n825));
  jand g0769(.dina(n825), .dinb(n467), .dout(n826));
  jand g0770(.dina(n826), .dinb(n579), .dout(n827));
  jand g0771(.dina(n254), .dinb(n222), .dout(n828));
  jand g0772(.dina(n828), .dinb(n301), .dout(n829));
  jand g0773(.dina(n829), .dinb(n504), .dout(n830));
  jand g0774(.dina(n830), .dinb(n827), .dout(n831));
  jand g0775(.dina(n831), .dinb(n824), .dout(n832));
  jand g0776(.dina(n451), .dinb(n294), .dout(n833));
  jand g0777(.dina(n833), .dinb(n832), .dout(n834));
  jand g0778(.dina(n561), .dinb(n312), .dout(n835));
  jand g0779(.dina(n835), .dinb(n130), .dout(n836));
  jnot g0780(.din(n586), .dout(n837));
  jand g0781(.dina(n402), .dinb(n270), .dout(n838));
  jand g0782(.dina(n838), .dinb(n837), .dout(n839));
  jand g0783(.dina(n839), .dinb(n836), .dout(n840));
  jnot g0784(.din(n550), .dout(n841));
  jand g0785(.dina(n501), .dinb(n216), .dout(n842));
  jand g0786(.dina(n842), .dinb(n147), .dout(n843));
  jand g0787(.dina(n843), .dinb(n841), .dout(n844));
  jand g0788(.dina(n844), .dinb(n840), .dout(n845));
  jand g0789(.dina(n662), .dinb(n470), .dout(n846));
  jand g0790(.dina(n632), .dinb(n304), .dout(n847));
  jand g0791(.dina(n847), .dinb(n846), .dout(n848));
  jnot g0792(.din(n608), .dout(n849));
  jand g0793(.dina(n849), .dinb(n420), .dout(n850));
  jand g0794(.dina(n850), .dinb(n623), .dout(n851));
  jand g0795(.dina(n851), .dinb(n848), .dout(n852));
  jor  g0796(.dina(n340), .dinb(n276), .dout(n853));
  jand g0797(.dina(n853), .dinb(n368), .dout(n854));
  jand g0798(.dina(n854), .dinb(n532), .dout(n855));
  jand g0799(.dina(n283), .dinb(n109), .dout(n856));
  jnot g0800(.din(n856), .dout(n857));
  jand g0801(.dina(n857), .dinb(n855), .dout(n858));
  jand g0802(.dina(n858), .dinb(n852), .dout(n859));
  jand g0803(.dina(n859), .dinb(n845), .dout(n860));
  jor  g0804(.dina(n748), .dinb(n641), .dout(n861));
  jor  g0805(.dina(n606), .dinb(n213), .dout(n862));
  jor  g0806(.dina(n862), .dinb(n861), .dout(n863));
  jnot g0807(.din(n863), .dout(n864));
  jand g0808(.dina(n645), .dinb(n768), .dout(n865));
  jor  g0809(.dina(n554), .dinb(n406), .dout(n866));
  jnot g0810(.din(n866), .dout(n867));
  jnot g0811(.din(n164), .dout(n868));
  jand g0812(.dina(n535), .dinb(n868), .dout(n869));
  jand g0813(.dina(n869), .dinb(n867), .dout(n870));
  jand g0814(.dina(n870), .dinb(n865), .dout(n871));
  jand g0815(.dina(n871), .dinb(n864), .dout(n872));
  jand g0816(.dina(n463), .dinb(n303), .dout(n873));
  jand g0817(.dina(n665), .dinb(n426), .dout(n874));
  jand g0818(.dina(n874), .dinb(n873), .dout(n875));
  jand g0819(.dina(n875), .dinb(n568), .dout(n876));
  jand g0820(.dina(n390), .dinb(n383), .dout(n877));
  jnot g0821(.din(n581), .dout(n878));
  jand g0822(.dina(n624), .dinb(n878), .dout(n879));
  jand g0823(.dina(n879), .dinb(n343), .dout(n880));
  jand g0824(.dina(n880), .dinb(n877), .dout(n881));
  jnot g0825(.din(n518), .dout(n882));
  jand g0826(.dina(n592), .dinb(n882), .dout(n883));
  jand g0827(.dina(n883), .dinb(n679), .dout(n884));
  jand g0828(.dina(n884), .dinb(n773), .dout(n885));
  jand g0829(.dina(n885), .dinb(n881), .dout(n886));
  jand g0830(.dina(n886), .dinb(n876), .dout(n887));
  jand g0831(.dina(n887), .dinb(n872), .dout(n888));
  jand g0832(.dina(n888), .dinb(n860), .dout(n889));
  jand g0833(.dina(n889), .dinb(n834), .dout(n890));
  jand g0834(.dina(n763), .dinb(n383), .dout(n891));
  jand g0835(.dina(n891), .dinb(n158), .dout(n892));
  jand g0836(.dina(n341), .dinb(n283), .dout(n893));
  jor  g0837(.dina(n893), .dinb(n269), .dout(n894));
  jnot g0838(.din(n894), .dout(n895));
  jand g0839(.dina(n895), .dinb(n324), .dout(n896));
  jnot g0840(.din(n160), .dout(n897));
  jand g0841(.dina(n229), .dinb(n897), .dout(n898));
  jand g0842(.dina(n898), .dinb(n771), .dout(n899));
  jand g0843(.dina(n899), .dinb(n896), .dout(n900));
  jand g0844(.dina(n900), .dinb(n892), .dout(n901));
  jand g0845(.dina(n901), .dinb(n648), .dout(n902));
  jand g0846(.dina(n561), .dinb(n343), .dout(n903));
  jand g0847(.dina(n903), .dinb(n902), .dout(n904));
  jand g0848(.dina(n479), .dinb(n397), .dout(n905));
  jand g0849(.dina(n579), .dinb(n370), .dout(n906));
  jand g0850(.dina(n216), .dinb(n138), .dout(n907));
  jand g0851(.dina(n907), .dinb(n906), .dout(n908));
  jand g0852(.dina(n908), .dinb(n905), .dout(n909));
  jand g0853(.dina(n662), .dinb(n612), .dout(n910));
  jand g0854(.dina(n730), .dinb(n868), .dout(n911));
  jand g0855(.dina(n911), .dinb(n910), .dout(n912));
  jand g0856(.dina(n849), .dinb(n254), .dout(n913));
  jand g0857(.dina(n913), .dinb(n426), .dout(n914));
  jand g0858(.dina(n914), .dinb(n912), .dout(n915));
  jand g0859(.dina(n734), .dinb(n251), .dout(n916));
  jand g0860(.dina(n916), .dinb(n463), .dout(n917));
  jnot g0861(.din(n551), .dout(n918));
  jand g0862(.dina(n614), .dinb(n918), .dout(n919));
  jand g0863(.dina(n919), .dinb(n130), .dout(n920));
  jand g0864(.dina(n920), .dinb(n917), .dout(n921));
  jand g0865(.dina(n921), .dinb(n915), .dout(n922));
  jand g0866(.dina(n922), .dinb(n909), .dout(n923));
  jand g0867(.dina(n437), .dinb(n421), .dout(n924));
  jnot g0868(.din(n588), .dout(n925));
  jand g0869(.dina(n925), .dinb(n461), .dout(n926));
  jand g0870(.dina(n926), .dinb(n924), .dout(n927));
  jnot g0871(.din(n732), .dout(n928));
  jor  g0872(.dina(n928), .dinb(n534), .dout(n929));
  jnot g0873(.din(n929), .dout(n930));
  jand g0874(.dina(n930), .dinb(n821), .dout(n931));
  jand g0875(.dina(n931), .dinb(n927), .dout(n932));
  jand g0876(.dina(n932), .dinb(n366), .dout(n933));
  jand g0877(.dina(n632), .dinb(n243), .dout(n934));
  jor  g0878(.dina(n409), .dinb(n146), .dout(n935));
  jand g0879(.dina(n935), .dinb(n256), .dout(n936));
  jand g0880(.dina(n936), .dinb(n934), .dout(n937));
  jand g0881(.dina(n225), .dinb(n147), .dout(n938));
  jand g0882(.dina(n938), .dinb(n883), .dout(n939));
  jand g0883(.dina(n939), .dinb(n937), .dout(n940));
  jand g0884(.dina(n710), .dinb(n445), .dout(n941));
  jand g0885(.dina(n941), .dinb(n625), .dout(n942));
  jand g0886(.dina(n501), .dinb(n387), .dout(n943));
  jand g0887(.dina(n781), .dinb(n379), .dout(n944));
  jand g0888(.dina(n944), .dinb(n943), .dout(n945));
  jand g0889(.dina(n945), .dinb(n942), .dout(n946));
  jand g0890(.dina(n946), .dinb(n940), .dout(n947));
  jand g0891(.dina(n947), .dinb(n933), .dout(n948));
  jand g0892(.dina(n948), .dinb(n923), .dout(n949));
  jand g0893(.dina(n949), .dinb(n904), .dout(n950));
  jxor g0894(.dina(n950), .dinb(n486), .dout(n951));
  jand g0895(.dina(n951), .dinb(n890), .dout(n952));
  jand g0896(.dina(n952), .dinb(n820), .dout(n953));
  jnot g0897(.din(n820), .dout(n954));
  jnot g0898(.din(n890), .dout(n955));
  jand g0899(.dina(n951), .dinb(n955), .dout(n956));
  jand g0900(.dina(n956), .dinb(n954), .dout(n957));
  jor  g0901(.dina(n957), .dinb(n953), .dout(n958));
  jand g0902(.dina(n88), .dinb(n49), .dout(n959));
  jxor g0903(.dina(n959), .dinb(a13 ), .dout(n960));
  jnot g0904(.din(n960), .dout(n961));
  jnot g0905(.din(n951), .dout(n962));
  jor  g0906(.dina(n950), .dinb(n486), .dout(n963));
  jand g0907(.dina(n963), .dinb(n955), .dout(n964));
  jnot g0908(.din(n964), .dout(n965));
  jand g0909(.dina(n965), .dinb(n962), .dout(n966));
  jand g0910(.dina(n966), .dinb(n961), .dout(n967));
  jnot g0911(.din(n486), .dout(n968));
  jand g0912(.dina(n890), .dinb(n968), .dout(n969));
  jor  g0913(.dina(n969), .dinb(n951), .dout(n970));
  jnot g0914(.din(n970), .dout(n971));
  jand g0915(.dina(n971), .dinb(n960), .dout(n972));
  jor  g0916(.dina(n972), .dinb(n967), .dout(n973));
  jor  g0917(.dina(n973), .dinb(n958), .dout(n974));
  jnot g0918(.din(n974), .dout(n975));
  jand g0919(.dina(a22 ), .dinb(a12 ), .dout(n976));
  jand g0920(.dina(n87), .dinb(a12 ), .dout(n977));
  jnot g0921(.din(n977), .dout(n978));
  jand g0922(.dina(n978), .dinb(n959), .dout(n979));
  jor  g0923(.dina(n979), .dinb(n976), .dout(n980));
  jnot g0924(.din(n980), .dout(n981));
  jand g0925(.dina(n379), .dinb(n254), .dout(n982));
  jand g0926(.dina(n853), .dinb(n232), .dout(n983));
  jand g0927(.dina(n983), .dinb(n982), .dout(n984));
  jand g0928(.dina(n354), .dinb(n227), .dout(n985));
  jor  g0929(.dina(n985), .dinb(n369), .dout(n986));
  jnot g0930(.din(n986), .dout(n987));
  jand g0931(.dina(n768), .dinb(n358), .dout(n988));
  jand g0932(.dina(n988), .dinb(n301), .dout(n989));
  jand g0933(.dina(n989), .dinb(n987), .dout(n990));
  jand g0934(.dina(n990), .dinb(n984), .dout(n991));
  jand g0935(.dina(n749), .dinb(n709), .dout(n992));
  jor  g0936(.dina(n340), .dinb(n380), .dout(n993));
  jand g0937(.dina(n993), .dinb(n421), .dout(n994));
  jand g0938(.dina(n506), .dinb(n381), .dout(n995));
  jand g0939(.dina(n995), .dinb(n994), .dout(n996));
  jand g0940(.dina(n996), .dinb(n992), .dout(n997));
  jand g0941(.dina(n772), .dinb(n249), .dout(n998));
  jand g0942(.dina(n998), .dinb(n303), .dout(n999));
  jand g0943(.dina(n291), .dinb(n267), .dout(n1000));
  jand g0944(.dina(n662), .dinb(n467), .dout(n1001));
  jand g0945(.dina(n1001), .dinb(n1000), .dout(n1002));
  jand g0946(.dina(n1002), .dinb(n999), .dout(n1003));
  jand g0947(.dina(n1003), .dinb(n997), .dout(n1004));
  jand g0948(.dina(n1004), .dinb(n991), .dout(n1005));
  jand g0949(.dina(n1005), .dinb(n904), .dout(n1006));
  jand g0950(.dina(n473), .dinb(n825), .dout(n1007));
  jand g0951(.dina(n285), .dinb(n256), .dout(n1008));
  jand g0952(.dina(n1008), .dinb(n1007), .dout(n1009));
  jand g0953(.dina(n1009), .dinb(n626), .dout(n1010));
  jand g0954(.dina(n1010), .dinb(n920), .dout(n1011));
  jand g0955(.dina(n732), .dinb(n138), .dout(n1012));
  jand g0956(.dina(n1012), .dinb(n1011), .dout(n1013));
  jand g0957(.dina(n632), .dinb(n882), .dout(n1014));
  jand g0958(.dina(n441), .dinb(n437), .dout(n1015));
  jand g0959(.dina(n1015), .dinb(n1014), .dout(n1016));
  jor  g0960(.dina(n309), .dinb(n260), .dout(n1017));
  jnot g0961(.din(n1017), .dout(n1018));
  jand g0962(.dina(n1018), .dinb(n543), .dout(n1019));
  jand g0963(.dina(n1019), .dinb(n1016), .dout(n1020));
  jand g0964(.dina(n765), .dinb(n665), .dout(n1021));
  jand g0965(.dina(n532), .dinb(n420), .dout(n1022));
  jand g0966(.dina(n1022), .dinb(n499), .dout(n1023));
  jand g0967(.dina(n1023), .dinb(n1021), .dout(n1024));
  jand g0968(.dina(n724), .dinb(n427), .dout(n1025));
  jand g0969(.dina(n1025), .dinb(n849), .dout(n1026));
  jand g0970(.dina(n710), .dinb(n399), .dout(n1027));
  jand g0971(.dina(n1027), .dinb(n1026), .dout(n1028));
  jand g0972(.dina(n1028), .dinb(n1024), .dout(n1029));
  jand g0973(.dina(n1029), .dinb(n1020), .dout(n1030));
  jand g0974(.dina(n1030), .dinb(n1013), .dout(n1031));
  jand g0975(.dina(n1031), .dinb(n1006), .dout(n1032));
  jxor g0976(.dina(n1032), .dinb(n890), .dout(n1033));
  jand g0977(.dina(n1033), .dinb(n762), .dout(n1034));
  jnot g0978(.din(n1034), .dout(n1035));
  jand g0979(.dina(n1035), .dinb(n981), .dout(n1036));
  jand g0980(.dina(n1033), .dinb(n790), .dout(n1037));
  jnot g0981(.din(n1037), .dout(n1038));
  jand g0982(.dina(n1038), .dinb(n980), .dout(n1039));
  jor  g0983(.dina(n1039), .dinb(n1036), .dout(n1040));
  jand g0984(.dina(n955), .dinb(n762), .dout(n1041));
  jor  g0985(.dina(n1041), .dinb(n1033), .dout(n1042));
  jnot g0986(.din(n1042), .dout(n1043));
  jand g0987(.dina(n1043), .dinb(n803), .dout(n1044));
  jnot g0988(.din(n1033), .dout(n1045));
  jor  g0989(.dina(n1032), .dinb(n890), .dout(n1046));
  jand g0990(.dina(n1046), .dinb(n790), .dout(n1047));
  jnot g0991(.din(n1047), .dout(n1048));
  jand g0992(.dina(n1048), .dinb(n1045), .dout(n1049));
  jand g0993(.dina(n1049), .dinb(n808), .dout(n1050));
  jor  g0994(.dina(n1050), .dinb(n1044), .dout(n1051));
  jnot g0995(.din(n1051), .dout(n1052));
  jand g0996(.dina(n1052), .dinb(n1040), .dout(n1053));
  jand g0997(.dina(n1053), .dinb(n975), .dout(n1054));
  jxor g0998(.dina(n1053), .dinb(n975), .dout(n1055));
  jxor g0999(.dina(n695), .dinb(a9 ), .dout(n1057));
  jand g1000(.dina(n1057), .dinb(n804), .dout(n1058));
  jnot g1001(.din(n1057), .dout(n1059));
  jand g1002(.dina(n1059), .dinb(n799), .dout(n1060));
  jor  g1003(.dina(n1060), .dinb(n1058), .dout(n1061));
  jand g1004(.dina(n789), .dinb(n794), .dout(n1063));
  jor  g1005(.dina(n1063), .dinb(n1061), .dout(n1065));
  jnot g1006(.din(n1065), .dout(n1066));
  jand g1007(.dina(n1066), .dinb(n1055), .dout(n1067));
  jor  g1008(.dina(n1067), .dinb(n1054), .dout(n1068));
  jxor g1009(.dina(n813), .dinb(n702), .dout(n1069));
  jand g1010(.dina(n1069), .dinb(n1068), .dout(n1070));
  jor  g1011(.dina(n1070), .dinb(n814), .dout(n1071));
  jand g1012(.dina(n1057), .dinb(n335), .dout(n1072));
  jnot g1013(.din(n1072), .dout(n1073));
  jxor g1014(.dina(n1073), .dinb(n964), .dout(n1074));
  jand g1015(.dina(n708), .dinb(n335), .dout(n1075));
  jxor g1016(.dina(n1075), .dinb(n1074), .dout(n1076));
  jand g1017(.dina(n1076), .dinb(n1071), .dout(n1077));
  jxor g1018(.dina(n1076), .dinb(n1071), .dout(n1078));
  jand g1019(.dina(n962), .dinb(n954), .dout(n1079));
  jor  g1020(.dina(n1079), .dinb(n964), .dout(n1080));
  jand g1021(.dina(n971), .dinb(n954), .dout(n1081));
  jnot g1022(.din(n1081), .dout(n1082));
  jand g1023(.dina(n1082), .dinb(n1080), .dout(n1083));
  jand g1024(.dina(n1083), .dinb(n1073), .dout(n1084));
  jxor g1025(.dina(n1083), .dinb(n1073), .dout(n1085));
  jand g1026(.dina(n1037), .dinb(n960), .dout(n1086));
  jand g1027(.dina(n1034), .dinb(n961), .dout(n1087));
  jor  g1028(.dina(n1087), .dinb(n1086), .dout(n1088));
  jand g1029(.dina(n1043), .dinb(n980), .dout(n1089));
  jand g1030(.dina(n1049), .dinb(n981), .dout(n1090));
  jor  g1031(.dina(n1090), .dinb(n1089), .dout(n1091));
  jor  g1032(.dina(n1091), .dinb(n1088), .dout(n1092));
  jnot g1033(.din(n1092), .dout(n1093));
  jand g1034(.dina(n1093), .dinb(n1085), .dout(n1094));
  jor  g1035(.dina(n1094), .dinb(n1084), .dout(n1095));
  jand g1036(.dina(n803), .dinb(n804), .dout(n1096));
  jand g1037(.dina(n808), .dinb(n799), .dout(n1097));
  jor  g1038(.dina(n1097), .dinb(n1096), .dout(n1098));
  jand g1039(.dina(n981), .dinb(n789), .dout(n1100));
  jor  g1040(.dina(n1100), .dinb(n1098), .dout(n1102));
  jand g1041(.dina(n1034), .dinb(n820), .dout(n1103));
  jand g1042(.dina(n1037), .dinb(n954), .dout(n1104));
  jor  g1043(.dina(n1104), .dinb(n1103), .dout(n1105));
  jand g1044(.dina(n1049), .dinb(n961), .dout(n1106));
  jand g1045(.dina(n1043), .dinb(n960), .dout(n1107));
  jor  g1046(.dina(n1107), .dinb(n1106), .dout(n1108));
  jor  g1047(.dina(n1108), .dinb(n1105), .dout(n1109));
  jxor g1048(.dina(n1109), .dinb(n1102), .dout(n1110));
  jxor g1049(.dina(n1110), .dinb(n1095), .dout(n1111));
  jand g1050(.dina(n1111), .dinb(n1078), .dout(n1112));
  jor  g1051(.dina(n1112), .dinb(n1077), .dout(n1113));
  jand g1052(.dina(n803), .dinb(n335), .dout(n1114));
  jnot g1053(.din(n1114), .dout(n1115));
  jand g1054(.dina(n1045), .dinb(n954), .dout(n1116));
  jor  g1055(.dina(n1116), .dinb(n1047), .dout(n1117));
  jand g1056(.dina(n1043), .dinb(n954), .dout(n1118));
  jnot g1057(.din(n1118), .dout(n1119));
  jand g1058(.dina(n1119), .dinb(n1117), .dout(n1120));
  jxor g1059(.dina(n1120), .dinb(n1115), .dout(n1121));
  jand g1060(.dina(n981), .dinb(n799), .dout(n1122));
  jand g1061(.dina(n980), .dinb(n804), .dout(n1123));
  jor  g1062(.dina(n1123), .dinb(n1122), .dout(n1124));
  jand g1063(.dina(n961), .dinb(n789), .dout(n1125));
  jor  g1064(.dina(n1125), .dinb(n1124), .dout(n1128));
  jnot g1065(.din(n1128), .dout(n1129));
  jxor g1066(.dina(n1129), .dinb(n1121), .dout(n1130));
  jand g1067(.dina(n1072), .dinb(n965), .dout(n1131));
  jand g1068(.dina(n1075), .dinb(n1074), .dout(n1132));
  jor  g1069(.dina(n1132), .dinb(n1131), .dout(n1133));
  jnot g1070(.din(n1102), .dout(n1134));
  jnot g1071(.din(n1109), .dout(n1135));
  jand g1072(.dina(n1135), .dinb(n1134), .dout(n1136));
  jand g1073(.dina(n1110), .dinb(n1095), .dout(n1137));
  jor  g1074(.dina(n1137), .dinb(n1136), .dout(n1138));
  jxor g1075(.dina(n1138), .dinb(n1133), .dout(n1139));
  jxor g1076(.dina(n1139), .dinb(n1130), .dout(n1140));
  jand g1077(.dina(n1140), .dinb(n1113), .dout(n1141));
  jand g1078(.dina(n792), .dinb(n699), .dout(n1142));
  jnot g1079(.din(n699), .dout(n1143));
  jand g1080(.dina(n800), .dinb(n1143), .dout(n1144));
  jor  g1081(.dina(n1144), .dinb(n1142), .dout(n1145));
  jand g1082(.dina(n1059), .dinb(n789), .dout(n1147));
  jnot g1083(.din(n1147), .dout(n1149));
  jand g1084(.dina(n1149), .dinb(n1145), .dout(n1150));
  jand g1085(.dina(n1042), .dinb(n708), .dout(n1151));
  jnot g1086(.din(n1049), .dout(n1152));
  jand g1087(.dina(n1152), .dinb(n794), .dout(n1153));
  jor  g1088(.dina(n1153), .dinb(n1151), .dout(n1154));
  jand g1089(.dina(n1037), .dinb(n803), .dout(n1155));
  jand g1090(.dina(n1034), .dinb(n808), .dout(n1156));
  jor  g1091(.dina(n1156), .dinb(n1155), .dout(n1157));
  jnot g1092(.din(n1157), .dout(n1158));
  jand g1093(.dina(n1158), .dinb(n1154), .dout(n1159));
  jand g1094(.dina(n1159), .dinb(n1150), .dout(n1160));
  jnot g1095(.din(n1160), .dout(n1161));
  jxor g1096(.dina(n1159), .dinb(n1150), .dout(n1162));
  jnot g1097(.din(n1162), .dout(n1163));
  jnot g1098(.din(n519), .dout(n1164));
  jand g1099(.dina(n1164), .dinb(n516), .dout(n1165));
  jand g1100(.dina(n525), .dinb(n1165), .dout(n1166));
  jand g1101(.dina(n1166), .dinb(n513), .dout(n1167));
  jand g1102(.dina(n1167), .dinb(n509), .dout(n1168));
  jand g1103(.dina(n1168), .dinb(n497), .dout(n1169));
  jnot g1104(.din(n545), .dout(n1170));
  jand g1105(.dina(n1170), .dinb(n543), .dout(n1171));
  jand g1106(.dina(n1171), .dinb(n541), .dout(n1172));
  jnot g1107(.din(n557), .dout(n1173));
  jand g1108(.dina(n1173), .dinb(n1172), .dout(n1174));
  jand g1109(.dina(n1174), .dinb(n538), .dout(n1175));
  jnot g1110(.din(n571), .dout(n1176));
  jand g1111(.dina(n1176), .dinb(n568), .dout(n1177));
  jand g1112(.dina(n1177), .dinb(n565), .dout(n1178));
  jnot g1113(.din(n584), .dout(n1179));
  jnot g1114(.din(n590), .dout(n1180));
  jand g1115(.dina(n598), .dinb(n1180), .dout(n1181));
  jand g1116(.dina(n1181), .dinb(n1179), .dout(n1182));
  jand g1117(.dina(n1182), .dinb(n1178), .dout(n1183));
  jand g1118(.dina(n1183), .dinb(n1175), .dout(n1184));
  jand g1119(.dina(n1184), .dinb(n1169), .dout(n1185));
  jand g1120(.dina(n624), .dinb(n506), .dout(n1186));
  jand g1121(.dina(n1186), .dinb(n837), .dout(n1187));
  jand g1122(.dina(n402), .dinb(n351), .dout(n1188));
  jand g1123(.dina(n1188), .dinb(n594), .dout(n1189));
  jor  g1124(.dina(n748), .dinb(n631), .dout(n1190));
  jnot g1125(.din(n1190), .dout(n1191));
  jand g1126(.dina(n427), .dinb(n348), .dout(n1192));
  jand g1127(.dina(n1192), .dinb(n1191), .dout(n1193));
  jand g1128(.dina(n1193), .dinb(n1189), .dout(n1194));
  jand g1129(.dina(n1194), .dinb(n1187), .dout(n1195));
  jand g1130(.dina(n744), .dinb(n279), .dout(n1196));
  jand g1131(.dina(n882), .dinb(n426), .dout(n1197));
  jor  g1132(.dina(n678), .dinb(n400), .dout(n1198));
  jnot g1133(.din(n1198), .dout(n1199));
  jand g1134(.dina(n1199), .dinb(n1197), .dout(n1200));
  jand g1135(.dina(n1200), .dinb(n1196), .dout(n1201));
  jand g1136(.dina(n1201), .dinb(n622), .dout(n1202));
  jand g1137(.dina(n1202), .dinb(n1195), .dout(n1203));
  jand g1138(.dina(n993), .dinb(n612), .dout(n1204));
  jand g1139(.dina(n1204), .dinb(n638), .dout(n1205));
  jand g1140(.dina(n1205), .dinb(n408), .dout(n1206));
  jand g1141(.dina(n579), .dinb(n363), .dout(n1207));
  jand g1142(.dina(n1207), .dinb(n454), .dout(n1208));
  jnot g1143(.din(n299), .dout(n1209));
  jand g1144(.dina(n935), .dinb(n1209), .dout(n1210));
  jand g1145(.dina(n1210), .dinb(n597), .dout(n1211));
  jand g1146(.dina(n1211), .dinb(n1208), .dout(n1212));
  jand g1147(.dina(n1212), .dinb(n1206), .dout(n1213));
  jor  g1148(.dina(n355), .dinb(n288), .dout(n1214));
  jor  g1149(.dina(n750), .dinb(n591), .dout(n1215));
  jor  g1150(.dina(n1215), .dinb(n475), .dout(n1216));
  jor  g1151(.dina(n1216), .dinb(n1214), .dout(n1217));
  jnot g1152(.din(n1217), .dout(n1218));
  jand g1153(.dina(n1218), .dinb(n858), .dout(n1219));
  jand g1154(.dina(n1219), .dinb(n1213), .dout(n1220));
  jor  g1155(.dina(n415), .dinb(n224), .dout(n1221));
  jand g1156(.dina(n501), .dinb(n381), .dout(n1222));
  jnot g1157(.din(n1222), .dout(n1223));
  jor  g1158(.dina(n1223), .dinb(n1221), .dout(n1224));
  jnot g1159(.din(n1224), .dout(n1225));
  jand g1160(.dina(n924), .dinb(n523), .dout(n1226));
  jor  g1161(.dina(n364), .dinb(n235), .dout(n1227));
  jnot g1162(.din(n1227), .dout(n1228));
  jand g1163(.dina(n1228), .dinb(n850), .dout(n1229));
  jand g1164(.dina(n1229), .dinb(n1226), .dout(n1230));
  jand g1165(.dina(n1230), .dinb(n1225), .dout(n1231));
  jand g1166(.dina(n354), .dinb(n259), .dout(n1232));
  jor  g1167(.dina(n1232), .dinb(n213), .dout(n1233));
  jor  g1168(.dina(n1233), .dinb(n552), .dout(n1234));
  jor  g1169(.dina(n780), .dinb(n250), .dout(n1235));
  jor  g1170(.dina(n373), .dinb(n266), .dout(n1236));
  jor  g1171(.dina(n1236), .dinb(n1235), .dout(n1237));
  jor  g1172(.dina(n1237), .dinb(n727), .dout(n1238));
  jor  g1173(.dina(n1238), .dinb(n1234), .dout(n1239));
  jnot g1174(.din(n1239), .dout(n1240));
  jand g1175(.dina(n1240), .dinb(n1231), .dout(n1241));
  jand g1176(.dina(n1241), .dinb(n1220), .dout(n1242));
  jand g1177(.dina(n1242), .dinb(n1203), .dout(n1243));
  jand g1178(.dina(n1243), .dinb(n1185), .dout(n1244));
  jnot g1179(.din(n1244), .dout(n1245));
  jnot g1180(.din(n1187), .dout(n1246));
  jnot g1181(.din(n1189), .dout(n1247));
  jnot g1182(.din(n1192), .dout(n1248));
  jor  g1183(.dina(n1248), .dinb(n1190), .dout(n1249));
  jor  g1184(.dina(n1249), .dinb(n1247), .dout(n1250));
  jor  g1185(.dina(n1250), .dinb(n1246), .dout(n1251));
  jnot g1186(.din(n622), .dout(n1252));
  jnot g1187(.din(n1196), .dout(n1253));
  jnot g1188(.din(n1197), .dout(n1254));
  jor  g1189(.dina(n1198), .dinb(n1254), .dout(n1255));
  jor  g1190(.dina(n1255), .dinb(n1253), .dout(n1256));
  jor  g1191(.dina(n1256), .dinb(n1252), .dout(n1257));
  jor  g1192(.dina(n1257), .dinb(n1251), .dout(n1258));
  jnot g1193(.din(n1204), .dout(n1259));
  jor  g1194(.dina(n1259), .dinb(n637), .dout(n1260));
  jor  g1195(.dina(n1260), .dinb(n407), .dout(n1261));
  jor  g1196(.dina(n580), .dinb(n362), .dout(n1262));
  jor  g1197(.dina(n1262), .dinb(n453), .dout(n1263));
  jnot g1198(.din(n597), .dout(n1264));
  jnot g1199(.din(n935), .dout(n1265));
  jor  g1200(.dina(n1265), .dinb(n299), .dout(n1266));
  jor  g1201(.dina(n1266), .dinb(n1264), .dout(n1267));
  jor  g1202(.dina(n1267), .dinb(n1263), .dout(n1268));
  jor  g1203(.dina(n1268), .dinb(n1261), .dout(n1269));
  jnot g1204(.din(n854), .dout(n1270));
  jor  g1205(.dina(n1270), .dinb(n531), .dout(n1271));
  jor  g1206(.dina(n856), .dinb(n1271), .dout(n1272));
  jor  g1207(.dina(n1217), .dinb(n1272), .dout(n1273));
  jor  g1208(.dina(n1273), .dinb(n1269), .dout(n1274));
  jnot g1209(.din(n924), .dout(n1275));
  jor  g1210(.dina(n1275), .dinb(n522), .dout(n1276));
  jor  g1211(.dina(n608), .dinb(n577), .dout(n1277));
  jor  g1212(.dina(n1227), .dinb(n1277), .dout(n1278));
  jor  g1213(.dina(n1278), .dinb(n1276), .dout(n1279));
  jor  g1214(.dina(n1279), .dinb(n1224), .dout(n1280));
  jor  g1215(.dina(n1239), .dinb(n1280), .dout(n1281));
  jor  g1216(.dina(n1281), .dinb(n1274), .dout(n1282));
  jor  g1217(.dina(n1282), .dinb(n1258), .dout(n1283));
  jand g1218(.dina(n882), .dinb(n479), .dout(n1284));
  jand g1219(.dina(n1284), .dinb(n724), .dout(n1285));
  jand g1220(.dina(n1285), .dinb(n1176), .dout(n1286));
  jand g1221(.dina(n1286), .dinb(n1027), .dout(n1287));
  jor  g1222(.dina(n560), .dinb(n231), .dout(n1288));
  jnot g1223(.din(n1288), .dout(n1289));
  jand g1224(.dina(n1289), .dinb(n733), .dout(n1290));
  jand g1225(.dina(n1204), .dinb(n934), .dout(n1291));
  jand g1226(.dina(n1291), .dinb(n1290), .dout(n1292));
  jor  g1227(.dina(n661), .dinb(n152), .dout(n1293));
  jnot g1228(.din(n1293), .dout(n1294));
  jand g1229(.dina(n1294), .dinb(n286), .dout(n1295));
  jand g1230(.dina(n1295), .dinb(n895), .dout(n1296));
  jand g1231(.dina(n1296), .dinb(n1292), .dout(n1297));
  jand g1232(.dina(n1297), .dinb(n1218), .dout(n1298));
  jand g1233(.dina(n1298), .dinb(n1287), .dout(n1299));
  jor  g1234(.dina(n406), .dinb(n386), .dout(n1300));
  jor  g1235(.dina(n266), .dinb(n224), .dout(n1301));
  jor  g1236(.dina(n1301), .dinb(n1300), .dout(n1302));
  jnot g1237(.din(n1302), .dout(n1303));
  jand g1238(.dina(n402), .dinb(n323), .dout(n1304));
  jand g1239(.dina(n1304), .dinb(n511), .dout(n1305));
  jand g1240(.dina(n1305), .dinb(n1018), .dout(n1306));
  jand g1241(.dina(n1306), .dinb(n1303), .dout(n1307));
  jnot g1242(.din(n596), .dout(n1308));
  jor  g1243(.dina(n1308), .dinb(n588), .dout(n1309));
  jnot g1244(.din(n1309), .dout(n1310));
  jand g1245(.dina(n935), .dinb(n515), .dout(n1311));
  jand g1246(.dina(n1311), .dinb(n384), .dout(n1312));
  jand g1247(.dina(n1312), .dinb(n1310), .dout(n1313));
  jand g1248(.dina(n458), .dinb(n422), .dout(n1314));
  jand g1249(.dina(n1314), .dinb(n295), .dout(n1315));
  jand g1250(.dina(n1315), .dinb(n843), .dout(n1316));
  jand g1251(.dina(n1316), .dinb(n677), .dout(n1317));
  jand g1252(.dina(n1317), .dinb(n1313), .dout(n1318));
  jand g1253(.dina(n1318), .dinb(n1307), .dout(n1319));
  jor  g1254(.dina(n521), .dinb(n411), .dout(n1320));
  jor  g1255(.dina(n290), .dinb(n228), .dout(n1321));
  jor  g1256(.dina(n1321), .dinb(n1320), .dout(n1322));
  jor  g1257(.dina(n593), .dinb(n137), .dout(n1323));
  jor  g1258(.dina(n1323), .dinb(n156), .dout(n1324));
  jor  g1259(.dina(n1324), .dinb(n1322), .dout(n1325));
  jnot g1260(.din(n1325), .dout(n1326));
  jand g1261(.dina(n1326), .dinb(n741), .dout(n1327));
  jand g1262(.dina(n781), .dinb(n451), .dout(n1328));
  jor  g1263(.dina(n670), .dinb(n644), .dout(n1329));
  jnot g1264(.din(n1329), .dout(n1330));
  jand g1265(.dina(n1330), .dinb(n1021), .dout(n1331));
  jand g1266(.dina(n1331), .dinb(n1328), .dout(n1332));
  jand g1267(.dina(n428), .dinb(n301), .dout(n1333));
  jand g1268(.dina(n1333), .dinb(n771), .dout(n1334));
  jand g1269(.dina(n1334), .dinb(n1332), .dout(n1335));
  jand g1270(.dina(n1335), .dinb(n1327), .dout(n1336));
  jand g1271(.dina(n1336), .dinb(n1319), .dout(n1337));
  jand g1272(.dina(n1337), .dinb(n1299), .dout(n1338));
  jor  g1273(.dina(n1338), .dinb(n1243), .dout(n1339));
  jand g1274(.dina(n1339), .dinb(n604), .dout(n1340));
  jand g1275(.dina(n1340), .dinb(n1283), .dout(n1341));
  jnot g1276(.din(n1341), .dout(n1342));
  jand g1277(.dina(a22 ), .dinb(a6 ), .dout(n1343));
  jand g1278(.dina(n81), .dinb(a6 ), .dout(n1344));
  jnot g1279(.din(n1344), .dout(n1345));
  jand g1280(.dina(n1345), .dinb(n336), .dout(n1346));
  jor  g1281(.dina(n1346), .dinb(n1343), .dout(n1347));
  jand g1282(.dina(n1347), .dinb(n335), .dout(n1348));
  jand g1283(.dina(n1348), .dinb(n1342), .dout(n1349));
  jnot g1284(.din(n1349), .dout(n1350));
  jand g1285(.dina(n1350), .dinb(n1245), .dout(n1351));
  jor  g1286(.dina(n1351), .dinb(n1163), .dout(n1352));
  jand g1287(.dina(n1352), .dinb(n1161), .dout(n1353));
  jnot g1288(.din(n1353), .dout(n1354));
  jnot g1289(.din(n338), .dout(n1355));
  jxor g1290(.dina(n688), .dinb(n1185), .dout(n1356));
  jnot g1291(.din(n1356), .dout(n1357));
  jand g1292(.dina(n1357), .dinb(n954), .dout(n1358));
  jnot g1293(.din(n1358), .dout(n1359));
  jand g1294(.dina(n1359), .dinb(n691), .dout(n1360));
  jand g1295(.dina(n688), .dinb(n1185), .dout(n1361));
  jor  g1296(.dina(n1361), .dinb(n968), .dout(n1362));
  jand g1297(.dina(n1362), .dinb(n1358), .dout(n1363));
  jor  g1298(.dina(n1363), .dinb(n1360), .dout(n1364));
  jnot g1299(.din(n1364), .dout(n1365));
  jand g1300(.dina(n1365), .dinb(n1355), .dout(n1366));
  jxor g1301(.dina(n1364), .dinb(n338), .dout(n1367));
  jand g1302(.dina(n960), .dinb(n956), .dout(n1368));
  jand g1303(.dina(n961), .dinb(n952), .dout(n1369));
  jor  g1304(.dina(n1369), .dinb(n1368), .dout(n1370));
  jand g1305(.dina(n980), .dinb(n971), .dout(n1371));
  jand g1306(.dina(n981), .dinb(n966), .dout(n1372));
  jor  g1307(.dina(n1372), .dinb(n1371), .dout(n1373));
  jor  g1308(.dina(n1373), .dinb(n1370), .dout(n1374));
  jnot g1309(.din(n1374), .dout(n1375));
  jand g1310(.dina(n1375), .dinb(n1367), .dout(n1376));
  jor  g1311(.dina(n1376), .dinb(n1366), .dout(n1377));
  jand g1312(.dina(n1377), .dinb(n1354), .dout(n1378));
  jxor g1313(.dina(n700), .dinb(n693), .dout(n1379));
  jxor g1314(.dina(n1377), .dinb(n1354), .dout(n1380));
  jand g1315(.dina(n1380), .dinb(n1379), .dout(n1381));
  jor  g1316(.dina(n1381), .dinb(n1378), .dout(n1382));
  jxor g1317(.dina(n1093), .dinb(n1085), .dout(n1383));
  jand g1318(.dina(n1383), .dinb(n1382), .dout(n1384));
  jxor g1319(.dina(n1383), .dinb(n1382), .dout(n1385));
  jxor g1320(.dina(n1069), .dinb(n1068), .dout(n1386));
  jand g1321(.dina(n1386), .dinb(n1385), .dout(n1387));
  jor  g1322(.dina(n1387), .dinb(n1384), .dout(n1388));
  jxor g1323(.dina(n1111), .dinb(n1078), .dout(n1389));
  jand g1324(.dina(n1389), .dinb(n1388), .dout(n1390));
  jnot g1325(.din(n337), .dout(n1391));
  jand g1326(.dina(n799), .dinb(n1391), .dout(n1392));
  jnot g1327(.din(n1392), .dout(n1393));
  jand g1328(.dina(n804), .dinb(n337), .dout(n1394));
  jnot g1329(.din(n1394), .dout(n1395));
  jxor g1330(.dina(n1143), .dinb(n334), .dout(n1396));
  jor  g1331(.dina(n1396), .dinb(n795), .dout(n1397));
  jand g1332(.dina(n1397), .dinb(n1395), .dout(n1398));
  jand g1333(.dina(n1398), .dinb(n1393), .dout(n1399));
  jand g1334(.dina(n1035), .dinb(n794), .dout(n1400));
  jand g1335(.dina(n1038), .dinb(n708), .dout(n1401));
  jor  g1336(.dina(n1401), .dinb(n1400), .dout(n1402));
  jand g1337(.dina(n1057), .dinb(n1043), .dout(n1403));
  jand g1338(.dina(n1059), .dinb(n1049), .dout(n1404));
  jor  g1339(.dina(n1404), .dinb(n1403), .dout(n1405));
  jnot g1340(.din(n1405), .dout(n1406));
  jand g1341(.dina(n1406), .dinb(n1402), .dout(n1407));
  jand g1342(.dina(n1407), .dinb(n1399), .dout(n1408));
  jxor g1343(.dina(n1407), .dinb(n1399), .dout(n1409));
  jnot g1344(.din(n1362), .dout(n1410));
  jor  g1345(.dina(n1410), .dinb(n1356), .dout(n1411));
  jand g1346(.dina(n1411), .dinb(n960), .dout(n1412));
  jnot g1347(.din(n691), .dout(n1413));
  jor  g1348(.dina(n1356), .dinb(n1413), .dout(n1414));
  jand g1349(.dina(n1414), .dinb(n961), .dout(n1415));
  jor  g1350(.dina(n1415), .dinb(n1412), .dout(n1416));
  jor  g1351(.dina(n1361), .dinb(n691), .dout(n1417));
  jnot g1352(.din(n1417), .dout(n1418));
  jand g1353(.dina(n1418), .dinb(n954), .dout(n1419));
  jor  g1354(.dina(n1362), .dinb(n690), .dout(n1420));
  jnot g1355(.din(n1420), .dout(n1421));
  jand g1356(.dina(n1421), .dinb(n820), .dout(n1422));
  jor  g1357(.dina(n1422), .dinb(n1419), .dout(n1423));
  jnot g1358(.din(n1423), .dout(n1424));
  jand g1359(.dina(n1424), .dinb(n1416), .dout(n1425));
  jand g1360(.dina(n1425), .dinb(n1409), .dout(n1426));
  jor  g1361(.dina(n1426), .dinb(n1408), .dout(n1427));
  jxor g1362(.dina(n1375), .dinb(n1367), .dout(n1428));
  jand g1363(.dina(n1428), .dinb(n1427), .dout(n1429));
  jxor g1364(.dina(n1351), .dinb(n1163), .dout(n1430));
  jxor g1365(.dina(n1428), .dinb(n1427), .dout(n1431));
  jand g1366(.dina(n1431), .dinb(n1430), .dout(n1432));
  jor  g1367(.dina(n1432), .dinb(n1429), .dout(n1433));
  jxor g1368(.dina(n1066), .dinb(n1055), .dout(n1434));
  jand g1369(.dina(n1434), .dinb(n1433), .dout(n1435));
  jxor g1370(.dina(n1434), .dinb(n1433), .dout(n1436));
  jxor g1371(.dina(n1380), .dinb(n1379), .dout(n1437));
  jand g1372(.dina(n1437), .dinb(n1436), .dout(n1438));
  jor  g1373(.dina(n1438), .dinb(n1435), .dout(n1439));
  jxor g1374(.dina(n1386), .dinb(n1385), .dout(n1440));
  jand g1375(.dina(n1440), .dinb(n1439), .dout(n1441));
  jand g1376(.dina(n1342), .dinb(n1245), .dout(n1442));
  jnot g1377(.din(n1442), .dout(n1443));
  jand g1378(.dina(n1443), .dinb(n1348), .dout(n1444));
  jand g1379(.dina(n1442), .dinb(n1350), .dout(n1445));
  jor  g1380(.dina(n1445), .dinb(n1444), .dout(n1446));
  jand g1381(.dina(n981), .dinb(n952), .dout(n1447));
  jand g1382(.dina(n980), .dinb(n956), .dout(n1448));
  jor  g1383(.dina(n1448), .dinb(n1447), .dout(n1449));
  jand g1384(.dina(n966), .dinb(n808), .dout(n1450));
  jand g1385(.dina(n971), .dinb(n803), .dout(n1451));
  jor  g1386(.dina(n1451), .dinb(n1450), .dout(n1452));
  jor  g1387(.dina(n1452), .dinb(n1449), .dout(n1453));
  jnot g1388(.din(n1453), .dout(n1454));
  jand g1389(.dina(n1454), .dinb(n1446), .dout(n1455));
  jand g1390(.dina(n335), .dinb(n55), .dout(n1456));
  jand g1391(.dina(n1456), .dinb(n1283), .dout(n1457));
  jxor g1392(.dina(n1456), .dinb(n1283), .dout(n1458));
  jnot g1393(.din(n1027), .dout(n1459));
  jnot g1394(.din(n1285), .dout(n1460));
  jor  g1395(.dina(n1460), .dinb(n571), .dout(n1461));
  jor  g1396(.dina(n1461), .dinb(n1459), .dout(n1462));
  jnot g1397(.din(n733), .dout(n1463));
  jor  g1398(.dina(n1288), .dinb(n1463), .dout(n1464));
  jnot g1399(.din(n243), .dout(n1465));
  jor  g1400(.dina(n631), .dinb(n1465), .dout(n1466));
  jor  g1401(.dina(n1259), .dinb(n1466), .dout(n1467));
  jor  g1402(.dina(n1467), .dinb(n1464), .dout(n1468));
  jnot g1403(.din(n282), .dout(n1469));
  jor  g1404(.dina(n284), .dinb(n1469), .dout(n1470));
  jor  g1405(.dina(n1293), .dinb(n1470), .dout(n1471));
  jor  g1406(.dina(n1471), .dinb(n894), .dout(n1472));
  jor  g1407(.dina(n1472), .dinb(n1468), .dout(n1473));
  jor  g1408(.dina(n1473), .dinb(n1217), .dout(n1474));
  jor  g1409(.dina(n1474), .dinb(n1462), .dout(n1475));
  jnot g1410(.din(n511), .dout(n1476));
  jnot g1411(.din(n402), .dout(n1477));
  jor  g1412(.dina(n1477), .dinb(n322), .dout(n1478));
  jor  g1413(.dina(n1478), .dinb(n1476), .dout(n1479));
  jor  g1414(.dina(n1479), .dinb(n1017), .dout(n1480));
  jor  g1415(.dina(n1480), .dinb(n1302), .dout(n1481));
  jnot g1416(.din(n1312), .dout(n1482));
  jor  g1417(.dina(n1482), .dinb(n1309), .dout(n1483));
  jnot g1418(.din(n676), .dout(n1484));
  jor  g1419(.dina(n1484), .dinb(n460), .dout(n1485));
  jnot g1420(.din(n147), .dout(n1486));
  jand g1421(.dina(n212), .dinb(n141), .dout(n1487));
  jand g1422(.dina(n468), .dinb(n96), .dout(n1488));
  jor  g1423(.dina(n1488), .dinb(n1487), .dout(n1489));
  jor  g1424(.dina(n1489), .dinb(n1486), .dout(n1490));
  jnot g1425(.din(n295), .dout(n1491));
  jor  g1426(.dina(n1232), .dinb(n985), .dout(n1492));
  jor  g1427(.dina(n1492), .dinb(n1491), .dout(n1493));
  jor  g1428(.dina(n1493), .dinb(n1490), .dout(n1494));
  jor  g1429(.dina(n1494), .dinb(n1485), .dout(n1495));
  jor  g1430(.dina(n1495), .dinb(n1483), .dout(n1496));
  jor  g1431(.dina(n1496), .dinb(n1481), .dout(n1497));
  jnot g1432(.din(n741), .dout(n1498));
  jor  g1433(.dina(n1325), .dinb(n1498), .dout(n1499));
  jnot g1434(.din(n1328), .dout(n1500));
  jor  g1435(.dina(n764), .dinb(n726), .dout(n1501));
  jor  g1436(.dina(n1329), .dinb(n1501), .dout(n1502));
  jor  g1437(.dina(n1502), .dinb(n1500), .dout(n1503));
  jnot g1438(.din(n771), .dout(n1504));
  jnot g1439(.din(n427), .dout(n1505));
  jor  g1440(.dina(n1505), .dinb(n425), .dout(n1506));
  jor  g1441(.dina(n1506), .dinb(n300), .dout(n1507));
  jor  g1442(.dina(n1507), .dinb(n1504), .dout(n1508));
  jor  g1443(.dina(n1508), .dinb(n1503), .dout(n1509));
  jor  g1444(.dina(n1509), .dinb(n1499), .dout(n1510));
  jor  g1445(.dina(n1510), .dinb(n1497), .dout(n1511));
  jor  g1446(.dina(n1511), .dinb(n1475), .dout(n1512));
  jand g1447(.dina(n1512), .dinb(n1283), .dout(n1513));
  jor  g1448(.dina(n1513), .dinb(n1185), .dout(n1514));
  jxor g1449(.dina(n1338), .dinb(n1243), .dout(n1515));
  jnot g1450(.din(n1515), .dout(n1516));
  jand g1451(.dina(n1516), .dinb(n954), .dout(n1517));
  jnot g1452(.din(n1517), .dout(n1518));
  jand g1453(.dina(n1518), .dinb(n1514), .dout(n1519));
  jand g1454(.dina(n1338), .dinb(n1243), .dout(n1520));
  jor  g1455(.dina(n1520), .dinb(n604), .dout(n1521));
  jand g1456(.dina(n1521), .dinb(n1517), .dout(n1522));
  jor  g1457(.dina(n1522), .dinb(n1519), .dout(n1523));
  jnot g1458(.din(n1523), .dout(n1524));
  jand g1459(.dina(n1524), .dinb(n1458), .dout(n1525));
  jor  g1460(.dina(n1525), .dinb(n1457), .dout(n1526));
  jxor g1461(.dina(n1454), .dinb(n1446), .dout(n1527));
  jand g1462(.dina(n1527), .dinb(n1526), .dout(n1528));
  jor  g1463(.dina(n1528), .dinb(n1455), .dout(n1529));
  jand g1464(.dina(n1418), .dinb(n960), .dout(n1530));
  jand g1465(.dina(n1421), .dinb(n961), .dout(n1531));
  jor  g1466(.dina(n1531), .dinb(n1530), .dout(n1532));
  jnot g1467(.din(n1411), .dout(n1533));
  jand g1468(.dina(n1533), .dinb(n980), .dout(n1534));
  jnot g1469(.din(n1414), .dout(n1535));
  jand g1470(.dina(n1535), .dinb(n981), .dout(n1536));
  jor  g1471(.dina(n1536), .dinb(n1534), .dout(n1537));
  jor  g1472(.dina(n1537), .dinb(n1532), .dout(n1538));
  jnot g1473(.din(n1538), .dout(n1539));
  jand g1474(.dina(n970), .dinb(n708), .dout(n1540));
  jnot g1475(.din(n966), .dout(n1541));
  jand g1476(.dina(n1541), .dinb(n794), .dout(n1542));
  jor  g1477(.dina(n1542), .dinb(n1540), .dout(n1543));
  jand g1478(.dina(n956), .dinb(n803), .dout(n1544));
  jand g1479(.dina(n952), .dinb(n808), .dout(n1545));
  jor  g1480(.dina(n1545), .dinb(n1544), .dout(n1546));
  jnot g1481(.din(n1546), .dout(n1547));
  jand g1482(.dina(n1547), .dinb(n1543), .dout(n1548));
  jand g1483(.dina(n1548), .dinb(n1539), .dout(n1549));
  jxor g1484(.dina(n1548), .dinb(n1539), .dout(n1550));
  jand g1485(.dina(n1042), .dinb(n699), .dout(n1551));
  jand g1486(.dina(n1152), .dinb(n1143), .dout(n1552));
  jor  g1487(.dina(n1552), .dinb(n1551), .dout(n1553));
  jand g1488(.dina(n1057), .dinb(n1037), .dout(n1554));
  jand g1489(.dina(n1059), .dinb(n1034), .dout(n1555));
  jor  g1490(.dina(n1555), .dinb(n1554), .dout(n1556));
  jnot g1491(.din(n1556), .dout(n1557));
  jand g1492(.dina(n1557), .dinb(n1553), .dout(n1558));
  jand g1493(.dina(n1558), .dinb(n1550), .dout(n1559));
  jor  g1494(.dina(n1559), .dinb(n1549), .dout(n1560));
  jxor g1495(.dina(n1425), .dinb(n1409), .dout(n1561));
  jand g1496(.dina(n1561), .dinb(n1560), .dout(n1562));
  jand g1497(.dina(n335), .dinb(n75), .dout(n1563));
  jand g1498(.dina(n1563), .dinb(n1283), .dout(n1564));
  jxor g1499(.dina(n1563), .dinb(n1283), .dout(n1565));
  jor  g1500(.dina(n1521), .dinb(n1513), .dout(n1566));
  jand g1501(.dina(n1566), .dinb(n820), .dout(n1567));
  jor  g1502(.dina(n1520), .dinb(n1514), .dout(n1568));
  jand g1503(.dina(n1568), .dinb(n954), .dout(n1569));
  jor  g1504(.dina(n1569), .dinb(n1567), .dout(n1570));
  jor  g1505(.dina(n1515), .dinb(n1340), .dout(n1571));
  jnot g1506(.din(n1571), .dout(n1572));
  jand g1507(.dina(n1572), .dinb(n961), .dout(n1573));
  jnot g1508(.din(n1520), .dout(n1574));
  jor  g1509(.dina(n1339), .dinb(n1185), .dout(n1575));
  jand g1510(.dina(n1575), .dinb(n1574), .dout(n1576));
  jnot g1511(.din(n1576), .dout(n1577));
  jand g1512(.dina(n1577), .dinb(n960), .dout(n1578));
  jor  g1513(.dina(n1578), .dinb(n1573), .dout(n1579));
  jnot g1514(.din(n1579), .dout(n1580));
  jand g1515(.dina(n1580), .dinb(n1570), .dout(n1581));
  jand g1516(.dina(n1581), .dinb(n1565), .dout(n1582));
  jor  g1517(.dina(n1582), .dinb(n1564), .dout(n1583));
  jnot g1518(.din(n1347), .dout(n1584));
  jand g1519(.dina(n1584), .dinb(n799), .dout(n1585));
  jand g1520(.dina(n1347), .dinb(n804), .dout(n1586));
  jor  g1521(.dina(n1586), .dinb(n1585), .dout(n1587));
  jand g1522(.dina(n789), .dinb(n1391), .dout(n1588));
  jor  g1523(.dina(n1588), .dinb(n1587), .dout(n1591));
  jnot g1524(.din(n1591), .dout(n1592));
  jand g1525(.dina(n1592), .dinb(n1583), .dout(n1593));
  jxor g1526(.dina(n1592), .dinb(n1583), .dout(n1594));
  jnot g1527(.din(n952), .dout(n1595));
  jand g1528(.dina(n1595), .dinb(n794), .dout(n1596));
  jnot g1529(.din(n956), .dout(n1597));
  jand g1530(.dina(n1597), .dinb(n708), .dout(n1598));
  jor  g1531(.dina(n1598), .dinb(n1596), .dout(n1599));
  jand g1532(.dina(n1057), .dinb(n971), .dout(n1600));
  jand g1533(.dina(n1059), .dinb(n966), .dout(n1601));
  jor  g1534(.dina(n1601), .dinb(n1600), .dout(n1602));
  jnot g1535(.din(n1602), .dout(n1603));
  jand g1536(.dina(n1603), .dinb(n1599), .dout(n1604));
  jand g1537(.dina(n1411), .dinb(n803), .dout(n1605));
  jand g1538(.dina(n1414), .dinb(n808), .dout(n1606));
  jor  g1539(.dina(n1606), .dinb(n1605), .dout(n1607));
  jand g1540(.dina(n1418), .dinb(n980), .dout(n1608));
  jand g1541(.dina(n1421), .dinb(n981), .dout(n1609));
  jor  g1542(.dina(n1609), .dinb(n1608), .dout(n1610));
  jnot g1543(.din(n1610), .dout(n1611));
  jand g1544(.dina(n1611), .dinb(n1607), .dout(n1612));
  jand g1545(.dina(n1612), .dinb(n1604), .dout(n1613));
  jxor g1546(.dina(n1612), .dinb(n1604), .dout(n1614));
  jand g1547(.dina(n1035), .dinb(n1143), .dout(n1615));
  jand g1548(.dina(n1038), .dinb(n699), .dout(n1616));
  jor  g1549(.dina(n1616), .dinb(n1615), .dout(n1617));
  jand g1550(.dina(n1043), .dinb(n337), .dout(n1618));
  jand g1551(.dina(n1049), .dinb(n1391), .dout(n1619));
  jor  g1552(.dina(n1619), .dinb(n1618), .dout(n1620));
  jnot g1553(.din(n1620), .dout(n1621));
  jand g1554(.dina(n1621), .dinb(n1617), .dout(n1622));
  jand g1555(.dina(n1622), .dinb(n1614), .dout(n1623));
  jor  g1556(.dina(n1623), .dinb(n1613), .dout(n1624));
  jand g1557(.dina(n1624), .dinb(n1594), .dout(n1625));
  jor  g1558(.dina(n1625), .dinb(n1593), .dout(n1626));
  jxor g1559(.dina(n1561), .dinb(n1560), .dout(n1627));
  jand g1560(.dina(n1627), .dinb(n1626), .dout(n1628));
  jor  g1561(.dina(n1628), .dinb(n1562), .dout(n1629));
  jand g1562(.dina(n1629), .dinb(n1529), .dout(n1630));
  jxor g1563(.dina(n1431), .dinb(n1430), .dout(n1631));
  jxor g1564(.dina(n1629), .dinb(n1529), .dout(n1632));
  jand g1565(.dina(n1632), .dinb(n1631), .dout(n1633));
  jor  g1566(.dina(n1633), .dinb(n1630), .dout(n1634));
  jxor g1567(.dina(n1437), .dinb(n1436), .dout(n1635));
  jand g1568(.dina(n1635), .dinb(n1634), .dout(n1636));
  jxor g1569(.dina(n1524), .dinb(n1458), .dout(n1637));
  jxor g1570(.dina(n1558), .dinb(n1550), .dout(n1638));
  jand g1571(.dina(n1638), .dinb(n1637), .dout(n1639));
  jand g1572(.dina(n335), .dinb(n58), .dout(n1640));
  jand g1573(.dina(n724), .dinb(n267), .dout(n1641));
  jand g1574(.dina(n1641), .dinb(n324), .dout(n1642));
  jand g1575(.dina(n713), .dinb(n676), .dout(n1643));
  jand g1576(.dina(n1643), .dinb(n1642), .dout(n1644));
  jnot g1577(.din(n1644), .dout(n1645));
  jand g1578(.dina(n905), .dinb(n232), .dout(n1646));
  jnot g1579(.din(n1646), .dout(n1647));
  jand g1580(.dina(n668), .dinb(n303), .dout(n1648));
  jand g1581(.dina(n1648), .dinb(n216), .dout(n1649));
  jnot g1582(.din(n1649), .dout(n1650));
  jor  g1583(.dina(n1650), .dinb(n863), .dout(n1651));
  jor  g1584(.dina(n1651), .dinb(n1647), .dout(n1652));
  jor  g1585(.dina(n1652), .dinb(n1645), .dout(n1653));
  jand g1586(.dina(n592), .dinb(n291), .dout(n1654));
  jand g1587(.dina(n1654), .dinb(n849), .dout(n1655));
  jnot g1588(.din(n1655), .dout(n1656));
  jnot g1589(.din(n994), .dout(n1657));
  jor  g1590(.dina(n764), .dinb(n588), .dout(n1658));
  jor  g1591(.dina(n1658), .dinb(n1657), .dout(n1659));
  jor  g1592(.dina(n1659), .dinb(n986), .dout(n1660));
  jor  g1593(.dina(n1660), .dinb(n1656), .dout(n1661));
  jor  g1594(.dina(n1661), .dinb(n167), .dout(n1662));
  jand g1595(.dina(n285), .dinb(n243), .dout(n1663));
  jand g1596(.dina(n426), .dinb(n304), .dout(n1664));
  jand g1597(.dina(n1664), .dinb(n1663), .dout(n1665));
  jnot g1598(.din(n1665), .dout(n1666));
  jor  g1599(.dina(n929), .dinb(n587), .dout(n1667));
  jor  g1600(.dina(n1667), .dinb(n866), .dout(n1668));
  jor  g1601(.dina(n1668), .dinb(n1666), .dout(n1669));
  jand g1602(.dina(n596), .dinb(n515), .dout(n1670));
  jand g1603(.dina(n1670), .dinb(n665), .dout(n1671));
  jnot g1604(.din(n1671), .dout(n1672));
  jand g1605(.dina(n645), .dinb(n348), .dout(n1673));
  jnot g1606(.din(n1673), .dout(n1674));
  jor  g1607(.dina(n389), .dinb(n378), .dout(n1675));
  jor  g1608(.dina(n574), .dinb(n505), .dout(n1676));
  jor  g1609(.dina(n1676), .dinb(n1675), .dout(n1677));
  jor  g1610(.dina(n1677), .dinb(n1674), .dout(n1678));
  jor  g1611(.dina(n1678), .dinb(n1672), .dout(n1679));
  jor  g1612(.dina(n1679), .dinb(n1669), .dout(n1680));
  jor  g1613(.dina(n1680), .dinb(n1662), .dout(n1681));
  jor  g1614(.dina(n1681), .dinb(n1653), .dout(n1682));
  jand g1615(.dina(n1682), .dinb(n1283), .dout(n1683));
  jand g1616(.dina(n1283), .dinb(n820), .dout(n1684));
  jor  g1617(.dina(n1684), .dinb(n1683), .dout(n1685));
  jand g1618(.dina(n1685), .dinb(n1640), .dout(n1686));
  jxor g1619(.dina(n1685), .dinb(n1640), .dout(n1687));
  jnot g1620(.din(n1568), .dout(n1688));
  jand g1621(.dina(n1688), .dinb(n960), .dout(n1689));
  jnot g1622(.din(n1566), .dout(n1690));
  jand g1623(.dina(n1690), .dinb(n961), .dout(n1691));
  jor  g1624(.dina(n1691), .dinb(n1689), .dout(n1692));
  jand g1625(.dina(n1577), .dinb(n980), .dout(n1693));
  jand g1626(.dina(n1572), .dinb(n981), .dout(n1694));
  jor  g1627(.dina(n1694), .dinb(n1693), .dout(n1695));
  jor  g1628(.dina(n1695), .dinb(n1692), .dout(n1696));
  jnot g1629(.din(n1696), .dout(n1697));
  jand g1630(.dina(n1697), .dinb(n1687), .dout(n1698));
  jor  g1631(.dina(n1698), .dinb(n1686), .dout(n1699));
  jand g1632(.dina(n804), .dinb(n55), .dout(n1700));
  jand g1633(.dina(n799), .dinb(n56), .dout(n1701));
  jor  g1634(.dina(n1701), .dinb(n1700), .dout(n1702));
  jand g1635(.dina(n1584), .dinb(n789), .dout(n1704));
  jor  g1636(.dina(n1704), .dinb(n1702), .dout(n1706));
  jnot g1637(.din(n1706), .dout(n1707));
  jand g1638(.dina(n1707), .dinb(n1699), .dout(n1708));
  jxor g1639(.dina(n1707), .dinb(n1699), .dout(n1709));
  jand g1640(.dina(n970), .dinb(n699), .dout(n1710));
  jand g1641(.dina(n1541), .dinb(n1143), .dout(n1711));
  jor  g1642(.dina(n1711), .dinb(n1710), .dout(n1712));
  jand g1643(.dina(n1057), .dinb(n956), .dout(n1713));
  jand g1644(.dina(n1059), .dinb(n952), .dout(n1714));
  jor  g1645(.dina(n1714), .dinb(n1713), .dout(n1715));
  jnot g1646(.din(n1715), .dout(n1716));
  jand g1647(.dina(n1716), .dinb(n1712), .dout(n1717));
  jand g1648(.dina(n1418), .dinb(n803), .dout(n1718));
  jand g1649(.dina(n1421), .dinb(n808), .dout(n1719));
  jor  g1650(.dina(n1719), .dinb(n1718), .dout(n1720));
  jand g1651(.dina(n1533), .dinb(n708), .dout(n1721));
  jand g1652(.dina(n1535), .dinb(n794), .dout(n1722));
  jor  g1653(.dina(n1722), .dinb(n1721), .dout(n1723));
  jor  g1654(.dina(n1723), .dinb(n1720), .dout(n1724));
  jnot g1655(.din(n1724), .dout(n1725));
  jand g1656(.dina(n1725), .dinb(n1717), .dout(n1726));
  jxor g1657(.dina(n1725), .dinb(n1717), .dout(n1727));
  jand g1658(.dina(n1037), .dinb(n337), .dout(n1728));
  jand g1659(.dina(n1034), .dinb(n1391), .dout(n1729));
  jor  g1660(.dina(n1729), .dinb(n1728), .dout(n1730));
  jand g1661(.dina(n1347), .dinb(n1043), .dout(n1731));
  jand g1662(.dina(n1584), .dinb(n1049), .dout(n1732));
  jor  g1663(.dina(n1732), .dinb(n1731), .dout(n1733));
  jor  g1664(.dina(n1733), .dinb(n1730), .dout(n1734));
  jnot g1665(.din(n1734), .dout(n1735));
  jand g1666(.dina(n1735), .dinb(n1727), .dout(n1736));
  jor  g1667(.dina(n1736), .dinb(n1726), .dout(n1737));
  jand g1668(.dina(n1737), .dinb(n1709), .dout(n1738));
  jor  g1669(.dina(n1738), .dinb(n1708), .dout(n1739));
  jxor g1670(.dina(n1638), .dinb(n1637), .dout(n1740));
  jand g1671(.dina(n1740), .dinb(n1739), .dout(n1741));
  jor  g1672(.dina(n1741), .dinb(n1639), .dout(n1742));
  jxor g1673(.dina(n1527), .dinb(n1526), .dout(n1743));
  jand g1674(.dina(n1743), .dinb(n1742), .dout(n1744));
  jxor g1675(.dina(n1743), .dinb(n1742), .dout(n1745));
  jxor g1676(.dina(n1627), .dinb(n1626), .dout(n1746));
  jand g1677(.dina(n1746), .dinb(n1745), .dout(n1747));
  jor  g1678(.dina(n1747), .dinb(n1744), .dout(n1748));
  jxor g1679(.dina(n1632), .dinb(n1631), .dout(n1749));
  jand g1680(.dina(n1749), .dinb(n1748), .dout(n1750));
  jand g1681(.dina(n789), .dinb(n58), .dout(n1751));
  jand g1682(.dina(n1682), .dinb(n954), .dout(n1754));
  jand g1683(.dina(n1754), .dinb(n1283), .dout(n1755));
  jnot g1684(.din(n1755), .dout(n1756));
  jand g1685(.dina(n1283), .dinb(n961), .dout(n1757));
  jor  g1686(.dina(n1757), .dinb(n1754), .dout(n1758));
  jor  g1687(.dina(n1758), .dinb(n1683), .dout(n1759));
  jand g1688(.dina(n1759), .dinb(n1756), .dout(n1760));
  jand g1689(.dina(n1760), .dinb(n335), .dout(n1761));
  jnot g1690(.din(n75), .dout(n1762));
  jand g1691(.dina(n799), .dinb(n1762), .dout(n1763));
  jand g1692(.dina(n804), .dinb(n75), .dout(n1764));
  jor  g1693(.dina(n1764), .dinb(n1763), .dout(n1765));
  jand g1694(.dina(n789), .dinb(n56), .dout(n1766));
  jor  g1695(.dina(n1766), .dinb(n1765), .dout(n1769));
  jnot g1696(.din(n1769), .dout(n1770));
  jand g1697(.dina(n1770), .dinb(n1761), .dout(n1771));
  jand g1698(.dina(n1595), .dinb(n1143), .dout(n1772));
  jand g1699(.dina(n1597), .dinb(n699), .dout(n1773));
  jor  g1700(.dina(n1773), .dinb(n1772), .dout(n1774));
  jand g1701(.dina(n971), .dinb(n337), .dout(n1775));
  jand g1702(.dina(n966), .dinb(n1391), .dout(n1776));
  jor  g1703(.dina(n1776), .dinb(n1775), .dout(n1777));
  jnot g1704(.din(n1777), .dout(n1778));
  jand g1705(.dina(n1778), .dinb(n1774), .dout(n1779));
  jand g1706(.dina(n1584), .dinb(n1034), .dout(n1780));
  jand g1707(.dina(n1347), .dinb(n1037), .dout(n1781));
  jor  g1708(.dina(n1781), .dinb(n1780), .dout(n1782));
  jand g1709(.dina(n1049), .dinb(n56), .dout(n1783));
  jand g1710(.dina(n1043), .dinb(n55), .dout(n1784));
  jor  g1711(.dina(n1784), .dinb(n1783), .dout(n1785));
  jor  g1712(.dina(n1785), .dinb(n1782), .dout(n1786));
  jnot g1713(.din(n1786), .dout(n1787));
  jand g1714(.dina(n1787), .dinb(n1779), .dout(n1788));
  jxor g1715(.dina(n1787), .dinb(n1779), .dout(n1789));
  jand g1716(.dina(n1411), .dinb(n1057), .dout(n1790));
  jand g1717(.dina(n1414), .dinb(n1059), .dout(n1791));
  jor  g1718(.dina(n1791), .dinb(n1790), .dout(n1792));
  jand g1719(.dina(n1418), .dinb(n708), .dout(n1793));
  jand g1720(.dina(n1421), .dinb(n794), .dout(n1794));
  jor  g1721(.dina(n1794), .dinb(n1793), .dout(n1795));
  jnot g1722(.din(n1795), .dout(n1796));
  jand g1723(.dina(n1796), .dinb(n1792), .dout(n1797));
  jand g1724(.dina(n1797), .dinb(n1789), .dout(n1798));
  jor  g1725(.dina(n1798), .dinb(n1788), .dout(n1799));
  jxor g1726(.dina(n1770), .dinb(n1761), .dout(n1800));
  jand g1727(.dina(n1800), .dinb(n1799), .dout(n1801));
  jor  g1728(.dina(n1801), .dinb(n1771), .dout(n1802));
  jxor g1729(.dina(n1581), .dinb(n1565), .dout(n1803));
  jand g1730(.dina(n1803), .dinb(n1802), .dout(n1804));
  jxor g1731(.dina(n1803), .dinb(n1802), .dout(n1805));
  jxor g1732(.dina(n1622), .dinb(n1614), .dout(n1806));
  jand g1733(.dina(n1806), .dinb(n1805), .dout(n1807));
  jor  g1734(.dina(n1807), .dinb(n1804), .dout(n1808));
  jxor g1735(.dina(n1624), .dinb(n1594), .dout(n1809));
  jand g1736(.dina(n1809), .dinb(n1808), .dout(n1810));
  jxor g1737(.dina(n1809), .dinb(n1808), .dout(n1811));
  jxor g1738(.dina(n1740), .dinb(n1739), .dout(n1812));
  jand g1739(.dina(n1812), .dinb(n1811), .dout(n1813));
  jor  g1740(.dina(n1813), .dinb(n1810), .dout(n1814));
  jxor g1741(.dina(n1746), .dinb(n1745), .dout(n1815));
  jand g1742(.dina(n1815), .dinb(n1814), .dout(n1816));
  jand g1743(.dina(n804), .dinb(n58), .dout(n1817));
  jand g1744(.dina(n799), .dinb(n59), .dout(n1818));
  jor  g1745(.dina(n1818), .dinb(n1817), .dout(n1819));
  jand g1746(.dina(n789), .dinb(n1762), .dout(n1821));
  jor  g1747(.dina(n1821), .dinb(n1819), .dout(n1823));
  jnot g1748(.din(n1823), .dout(n1824));
  jand g1749(.dina(n1566), .dinb(n981), .dout(n1825));
  jand g1750(.dina(n1568), .dinb(n980), .dout(n1826));
  jor  g1751(.dina(n1826), .dinb(n1825), .dout(n1827));
  jand g1752(.dina(n1572), .dinb(n808), .dout(n1828));
  jand g1753(.dina(n1577), .dinb(n803), .dout(n1829));
  jor  g1754(.dina(n1829), .dinb(n1828), .dout(n1830));
  jnot g1755(.din(n1830), .dout(n1831));
  jand g1756(.dina(n1831), .dinb(n1827), .dout(n1832));
  jand g1757(.dina(n1832), .dinb(n1824), .dout(n1833));
  jxor g1758(.dina(n1760), .dinb(n335), .dout(n1834));
  jxor g1759(.dina(n1832), .dinb(n1824), .dout(n1835));
  jand g1760(.dina(n1835), .dinb(n1834), .dout(n1836));
  jor  g1761(.dina(n1836), .dinb(n1833), .dout(n1837));
  jxor g1762(.dina(n1697), .dinb(n1687), .dout(n1838));
  jand g1763(.dina(n1838), .dinb(n1837), .dout(n1839));
  jxor g1764(.dina(n1838), .dinb(n1837), .dout(n1840));
  jxor g1765(.dina(n1735), .dinb(n1727), .dout(n1841));
  jand g1766(.dina(n1841), .dinb(n1840), .dout(n1842));
  jor  g1767(.dina(n1842), .dinb(n1839), .dout(n1843));
  jxor g1768(.dina(n1737), .dinb(n1709), .dout(n1844));
  jand g1769(.dina(n1844), .dinb(n1843), .dout(n1845));
  jxor g1770(.dina(n1844), .dinb(n1843), .dout(n1846));
  jxor g1771(.dina(n1806), .dinb(n1805), .dout(n1847));
  jand g1772(.dina(n1847), .dinb(n1846), .dout(n1848));
  jor  g1773(.dina(n1848), .dinb(n1845), .dout(n1849));
  jxor g1774(.dina(n1812), .dinb(n1811), .dout(n1850));
  jand g1775(.dina(n1850), .dinb(n1849), .dout(n1851));
  jand g1776(.dina(n1418), .dinb(n1057), .dout(n1852));
  jand g1777(.dina(n1421), .dinb(n1059), .dout(n1853));
  jor  g1778(.dina(n1853), .dinb(n1852), .dout(n1854));
  jand g1779(.dina(n1533), .dinb(n699), .dout(n1855));
  jand g1780(.dina(n1535), .dinb(n1143), .dout(n1856));
  jor  g1781(.dina(n1856), .dinb(n1855), .dout(n1857));
  jor  g1782(.dina(n1857), .dinb(n1854), .dout(n1858));
  jnot g1783(.din(n1858), .dout(n1859));
  jand g1784(.dina(n956), .dinb(n337), .dout(n1860));
  jand g1785(.dina(n952), .dinb(n1391), .dout(n1861));
  jor  g1786(.dina(n1861), .dinb(n1860), .dout(n1862));
  jand g1787(.dina(n1347), .dinb(n971), .dout(n1863));
  jand g1788(.dina(n1584), .dinb(n966), .dout(n1864));
  jor  g1789(.dina(n1864), .dinb(n1863), .dout(n1865));
  jor  g1790(.dina(n1865), .dinb(n1862), .dout(n1866));
  jnot g1791(.din(n1866), .dout(n1867));
  jand g1792(.dina(n1867), .dinb(n1859), .dout(n1868));
  jand g1793(.dina(n1033), .dinb(n58), .dout(n1869));
  jnot g1794(.din(n1869), .dout(n1870));
  jand g1795(.dina(n1870), .dinb(n1047), .dout(n1871));
  jand g1796(.dina(n1682), .dinb(n980), .dout(n1872));
  jand g1797(.dina(n1872), .dinb(n1283), .dout(n1873));
  jnot g1798(.din(n1873), .dout(n1874));
  jand g1799(.dina(n1283), .dinb(n808), .dout(n1875));
  jor  g1800(.dina(n1875), .dinb(n1872), .dout(n1876));
  jor  g1801(.dina(n1876), .dinb(n1683), .dout(n1877));
  jand g1802(.dina(n1877), .dinb(n1874), .dout(n1878));
  jand g1803(.dina(n1878), .dinb(n1871), .dout(n1879));
  jxor g1804(.dina(n1866), .dinb(n1858), .dout(n1880));
  jand g1805(.dina(n1880), .dinb(n1879), .dout(n1881));
  jor  g1806(.dina(n1881), .dinb(n1868), .dout(n1882));
  jand g1807(.dina(n1682), .dinb(n960), .dout(n1883));
  jand g1808(.dina(n1883), .dinb(n1283), .dout(n1884));
  jnot g1809(.din(n1884), .dout(n1885));
  jand g1810(.dina(n1283), .dinb(n981), .dout(n1886));
  jor  g1811(.dina(n1886), .dinb(n1883), .dout(n1887));
  jor  g1812(.dina(n1887), .dinb(n1683), .dout(n1888));
  jand g1813(.dina(n1888), .dinb(n1885), .dout(n1889));
  jand g1814(.dina(n1688), .dinb(n803), .dout(n1890));
  jand g1815(.dina(n1690), .dinb(n808), .dout(n1891));
  jor  g1816(.dina(n1891), .dinb(n1890), .dout(n1892));
  jand g1817(.dina(n1577), .dinb(n708), .dout(n1893));
  jand g1818(.dina(n1572), .dinb(n794), .dout(n1894));
  jor  g1819(.dina(n1894), .dinb(n1893), .dout(n1895));
  jor  g1820(.dina(n1895), .dinb(n1892), .dout(n1896));
  jnot g1821(.din(n1896), .dout(n1897));
  jand g1822(.dina(n1897), .dinb(n1889), .dout(n1898));
  jxor g1823(.dina(n1897), .dinb(n1889), .dout(n1899));
  jand g1824(.dina(n1037), .dinb(n55), .dout(n1900));
  jand g1825(.dina(n1034), .dinb(n56), .dout(n1901));
  jor  g1826(.dina(n1901), .dinb(n1900), .dout(n1902));
  jand g1827(.dina(n1043), .dinb(n75), .dout(n1903));
  jand g1828(.dina(n1049), .dinb(n1762), .dout(n1904));
  jor  g1829(.dina(n1904), .dinb(n1903), .dout(n1905));
  jor  g1830(.dina(n1905), .dinb(n1902), .dout(n1906));
  jnot g1831(.din(n1906), .dout(n1907));
  jand g1832(.dina(n1907), .dinb(n1899), .dout(n1908));
  jor  g1833(.dina(n1908), .dinb(n1898), .dout(n1909));
  jand g1834(.dina(n1909), .dinb(n1882), .dout(n1910));
  jxor g1835(.dina(n1909), .dinb(n1882), .dout(n1911));
  jxor g1836(.dina(n1797), .dinb(n1789), .dout(n1912));
  jand g1837(.dina(n1912), .dinb(n1911), .dout(n1913));
  jor  g1838(.dina(n1913), .dinb(n1910), .dout(n1914));
  jxor g1839(.dina(n1800), .dinb(n1799), .dout(n1915));
  jand g1840(.dina(n1915), .dinb(n1914), .dout(n1916));
  jxor g1841(.dina(n1915), .dinb(n1914), .dout(n1917));
  jxor g1842(.dina(n1841), .dinb(n1840), .dout(n1918));
  jand g1843(.dina(n1918), .dinb(n1917), .dout(n1919));
  jor  g1844(.dina(n1919), .dinb(n1916), .dout(n1920));
  jxor g1845(.dina(n1847), .dinb(n1846), .dout(n1921));
  jand g1846(.dina(n1921), .dinb(n1920), .dout(n1922));
  jand g1847(.dina(n1566), .dinb(n794), .dout(n1923));
  jand g1848(.dina(n1568), .dinb(n708), .dout(n1924));
  jor  g1849(.dina(n1924), .dinb(n1923), .dout(n1925));
  jand g1850(.dina(n1572), .dinb(n1059), .dout(n1926));
  jand g1851(.dina(n1577), .dinb(n1057), .dout(n1927));
  jor  g1852(.dina(n1927), .dinb(n1926), .dout(n1928));
  jnot g1853(.din(n1928), .dout(n1929));
  jand g1854(.dina(n1929), .dinb(n1925), .dout(n1930));
  jand g1855(.dina(n1584), .dinb(n952), .dout(n1931));
  jand g1856(.dina(n1347), .dinb(n956), .dout(n1932));
  jor  g1857(.dina(n1932), .dinb(n1931), .dout(n1933));
  jand g1858(.dina(n966), .dinb(n56), .dout(n1934));
  jand g1859(.dina(n971), .dinb(n55), .dout(n1935));
  jor  g1860(.dina(n1935), .dinb(n1934), .dout(n1936));
  jor  g1861(.dina(n1936), .dinb(n1933), .dout(n1937));
  jnot g1862(.din(n1937), .dout(n1938));
  jand g1863(.dina(n1938), .dinb(n1930), .dout(n1939));
  jxor g1864(.dina(n1938), .dinb(n1930), .dout(n1940));
  jand g1865(.dina(n1411), .dinb(n337), .dout(n1941));
  jand g1866(.dina(n1414), .dinb(n1391), .dout(n1942));
  jor  g1867(.dina(n1942), .dinb(n1941), .dout(n1943));
  jand g1868(.dina(n1418), .dinb(n699), .dout(n1944));
  jand g1869(.dina(n1421), .dinb(n1143), .dout(n1945));
  jor  g1870(.dina(n1945), .dinb(n1944), .dout(n1946));
  jnot g1871(.din(n1946), .dout(n1947));
  jand g1872(.dina(n1947), .dinb(n1943), .dout(n1948));
  jand g1873(.dina(n1948), .dinb(n1940), .dout(n1949));
  jor  g1874(.dina(n1949), .dinb(n1939), .dout(n1950));
  jand g1875(.dina(n1950), .dinb(n1751), .dout(n1951));
  jxor g1876(.dina(n1880), .dinb(n1879), .dout(n1952));
  jxor g1877(.dina(n1950), .dinb(n1751), .dout(n1953));
  jand g1878(.dina(n1953), .dinb(n1952), .dout(n1954));
  jor  g1879(.dina(n1954), .dinb(n1951), .dout(n1955));
  jxor g1880(.dina(n1835), .dinb(n1834), .dout(n1956));
  jand g1881(.dina(n1956), .dinb(n1955), .dout(n1957));
  jxor g1882(.dina(n1956), .dinb(n1955), .dout(n1958));
  jxor g1883(.dina(n1912), .dinb(n1911), .dout(n1959));
  jand g1884(.dina(n1959), .dinb(n1958), .dout(n1960));
  jor  g1885(.dina(n1960), .dinb(n1957), .dout(n1961));
  jxor g1886(.dina(n1918), .dinb(n1917), .dout(n1962));
  jand g1887(.dina(n1962), .dinb(n1961), .dout(n1963));
  jxor g1888(.dina(n1962), .dinb(n1961), .dout(n1964));
  jxor g1889(.dina(n1878), .dinb(n1871), .dout(n1965));
  jand g1890(.dina(n1034), .dinb(n1762), .dout(n1966));
  jand g1891(.dina(n1037), .dinb(n75), .dout(n1967));
  jor  g1892(.dina(n1967), .dinb(n1966), .dout(n1968));
  jand g1893(.dina(n1049), .dinb(n59), .dout(n1969));
  jand g1894(.dina(n1043), .dinb(n58), .dout(n1970));
  jor  g1895(.dina(n1970), .dinb(n1969), .dout(n1971));
  jor  g1896(.dina(n1971), .dinb(n1968), .dout(n1972));
  jnot g1897(.din(n1972), .dout(n1973));
  jand g1898(.dina(n1973), .dinb(n1965), .dout(n1974));
  jand g1899(.dina(n1682), .dinb(n803), .dout(n1975));
  jand g1900(.dina(n1975), .dinb(n1283), .dout(n1976));
  jnot g1901(.din(n1976), .dout(n1977));
  jand g1902(.dina(n1283), .dinb(n794), .dout(n1978));
  jor  g1903(.dina(n1978), .dinb(n1975), .dout(n1979));
  jor  g1904(.dina(n1979), .dinb(n1683), .dout(n1980));
  jand g1905(.dina(n1980), .dinb(n1977), .dout(n1981));
  jand g1906(.dina(n1688), .dinb(n1057), .dout(n1982));
  jand g1907(.dina(n1690), .dinb(n1059), .dout(n1983));
  jor  g1908(.dina(n1983), .dinb(n1982), .dout(n1984));
  jand g1909(.dina(n1577), .dinb(n699), .dout(n1985));
  jand g1910(.dina(n1572), .dinb(n1143), .dout(n1986));
  jor  g1911(.dina(n1986), .dinb(n1985), .dout(n1987));
  jor  g1912(.dina(n1987), .dinb(n1984), .dout(n1988));
  jnot g1913(.din(n1988), .dout(n1989));
  jand g1914(.dina(n1989), .dinb(n1981), .dout(n1990));
  jxor g1915(.dina(n1989), .dinb(n1981), .dout(n1991));
  jand g1916(.dina(n1418), .dinb(n337), .dout(n1992));
  jand g1917(.dina(n1421), .dinb(n1391), .dout(n1993));
  jor  g1918(.dina(n1993), .dinb(n1992), .dout(n1994));
  jand g1919(.dina(n1533), .dinb(n1347), .dout(n1995));
  jand g1920(.dina(n1535), .dinb(n1584), .dout(n1996));
  jor  g1921(.dina(n1996), .dinb(n1995), .dout(n1997));
  jor  g1922(.dina(n1997), .dinb(n1994), .dout(n1998));
  jnot g1923(.din(n1998), .dout(n1999));
  jand g1924(.dina(n1999), .dinb(n1991), .dout(n2000));
  jor  g1925(.dina(n2000), .dinb(n1990), .dout(n2001));
  jxor g1926(.dina(n1973), .dinb(n1965), .dout(n2002));
  jand g1927(.dina(n2002), .dinb(n2001), .dout(n2003));
  jor  g1928(.dina(n2003), .dinb(n1974), .dout(n2004));
  jxor g1929(.dina(n1907), .dinb(n1899), .dout(n2005));
  jand g1930(.dina(n2005), .dinb(n2004), .dout(n2006));
  jxor g1931(.dina(n1953), .dinb(n1952), .dout(n2007));
  jxor g1932(.dina(n2005), .dinb(n2004), .dout(n2008));
  jand g1933(.dina(n2008), .dinb(n2007), .dout(n2009));
  jor  g1934(.dina(n2009), .dinb(n2006), .dout(n2010));
  jand g1935(.dina(n951), .dinb(n58), .dout(n2011));
  jnot g1936(.din(n2011), .dout(n2012));
  jand g1937(.dina(n2012), .dinb(n964), .dout(n2013));
  jand g1938(.dina(n1682), .dinb(n708), .dout(n2014));
  jand g1939(.dina(n2014), .dinb(n1283), .dout(n2015));
  jnot g1940(.din(n2015), .dout(n2016));
  jand g1941(.dina(n1283), .dinb(n1059), .dout(n2017));
  jor  g1942(.dina(n2017), .dinb(n2014), .dout(n2018));
  jor  g1943(.dina(n2018), .dinb(n1683), .dout(n2019));
  jand g1944(.dina(n2019), .dinb(n2016), .dout(n2020));
  jand g1945(.dina(n2020), .dinb(n2013), .dout(n2021));
  jand g1946(.dina(n956), .dinb(n55), .dout(n2022));
  jand g1947(.dina(n952), .dinb(n56), .dout(n2023));
  jor  g1948(.dina(n2023), .dinb(n2022), .dout(n2024));
  jand g1949(.dina(n971), .dinb(n75), .dout(n2025));
  jand g1950(.dina(n966), .dinb(n1762), .dout(n2026));
  jor  g1951(.dina(n2026), .dinb(n2025), .dout(n2027));
  jor  g1952(.dina(n2027), .dinb(n2024), .dout(n2028));
  jnot g1953(.din(n2028), .dout(n2029));
  jand g1954(.dina(n2029), .dinb(n2021), .dout(n2030));
  jxor g1955(.dina(n2029), .dinb(n2021), .dout(n2031));
  jand g1956(.dina(n2031), .dinb(n1869), .dout(n2032));
  jor  g1957(.dina(n2032), .dinb(n2030), .dout(n2033));
  jxor g1958(.dina(n1948), .dinb(n1940), .dout(n2034));
  jand g1959(.dina(n2034), .dinb(n2033), .dout(n2035));
  jxor g1960(.dina(n2034), .dinb(n2033), .dout(n2036));
  jxor g1961(.dina(n2002), .dinb(n2001), .dout(n2037));
  jand g1962(.dina(n2037), .dinb(n2036), .dout(n2038));
  jor  g1963(.dina(n2038), .dinb(n2035), .dout(n2039));
  jand g1964(.dina(n1566), .dinb(n1143), .dout(n2040));
  jand g1965(.dina(n1568), .dinb(n699), .dout(n2041));
  jor  g1966(.dina(n2041), .dinb(n2040), .dout(n2042));
  jand g1967(.dina(n1572), .dinb(n1391), .dout(n2043));
  jand g1968(.dina(n1577), .dinb(n337), .dout(n2044));
  jor  g1969(.dina(n2044), .dinb(n2043), .dout(n2045));
  jnot g1970(.din(n2045), .dout(n2046));
  jand g1971(.dina(n2046), .dinb(n2042), .dout(n2047));
  jand g1972(.dina(n1411), .dinb(n55), .dout(n2048));
  jand g1973(.dina(n1414), .dinb(n56), .dout(n2049));
  jor  g1974(.dina(n2049), .dinb(n2048), .dout(n2050));
  jand g1975(.dina(n1418), .dinb(n1347), .dout(n2051));
  jand g1976(.dina(n1421), .dinb(n1584), .dout(n2052));
  jor  g1977(.dina(n2052), .dinb(n2051), .dout(n2053));
  jnot g1978(.din(n2053), .dout(n2054));
  jand g1979(.dina(n2054), .dinb(n2050), .dout(n2055));
  jand g1980(.dina(n2055), .dinb(n2047), .dout(n2056));
  jxor g1981(.dina(n2055), .dinb(n2047), .dout(n2057));
  jand g1982(.dina(n952), .dinb(n1762), .dout(n2058));
  jand g1983(.dina(n956), .dinb(n75), .dout(n2059));
  jor  g1984(.dina(n2059), .dinb(n2058), .dout(n2060));
  jand g1985(.dina(n966), .dinb(n59), .dout(n2061));
  jand g1986(.dina(n971), .dinb(n58), .dout(n2062));
  jor  g1987(.dina(n2062), .dinb(n2061), .dout(n2063));
  jor  g1988(.dina(n2063), .dinb(n2060), .dout(n2064));
  jnot g1989(.din(n2064), .dout(n2065));
  jand g1990(.dina(n2065), .dinb(n2057), .dout(n2066));
  jor  g1991(.dina(n2066), .dinb(n2056), .dout(n2067));
  jxor g1992(.dina(n1999), .dinb(n1991), .dout(n2068));
  jand g1993(.dina(n2068), .dinb(n2067), .dout(n2069));
  jxor g1994(.dina(n2031), .dinb(n1869), .dout(n2070));
  jxor g1995(.dina(n2068), .dinb(n2067), .dout(n2071));
  jand g1996(.dina(n2071), .dinb(n2070), .dout(n2072));
  jor  g1997(.dina(n2072), .dinb(n2069), .dout(n2073));
  jxor g1998(.dina(n2020), .dinb(n2013), .dout(n2074));
  jand g1999(.dina(n1682), .dinb(n1057), .dout(n2075));
  jand g2000(.dina(n2075), .dinb(n1283), .dout(n2076));
  jnot g2001(.din(n2076), .dout(n2077));
  jand g2002(.dina(n1283), .dinb(n1143), .dout(n2078));
  jor  g2003(.dina(n2078), .dinb(n2075), .dout(n2079));
  jor  g2004(.dina(n2079), .dinb(n1683), .dout(n2080));
  jand g2005(.dina(n2080), .dinb(n2077), .dout(n2081));
  jand g2006(.dina(n1688), .dinb(n337), .dout(n2082));
  jand g2007(.dina(n1690), .dinb(n1391), .dout(n2083));
  jor  g2008(.dina(n2083), .dinb(n2082), .dout(n2084));
  jand g2009(.dina(n1577), .dinb(n1347), .dout(n2085));
  jand g2010(.dina(n1572), .dinb(n1584), .dout(n2086));
  jor  g2011(.dina(n2086), .dinb(n2085), .dout(n2087));
  jor  g2012(.dina(n2087), .dinb(n2084), .dout(n2088));
  jnot g2013(.din(n2088), .dout(n2089));
  jand g2014(.dina(n2089), .dinb(n2081), .dout(n2090));
  jxor g2015(.dina(n2089), .dinb(n2081), .dout(n2091));
  jand g2016(.dina(n1418), .dinb(n55), .dout(n2092));
  jand g2017(.dina(n1421), .dinb(n56), .dout(n2093));
  jor  g2018(.dina(n2093), .dinb(n2092), .dout(n2094));
  jand g2019(.dina(n1533), .dinb(n75), .dout(n2095));
  jand g2020(.dina(n1535), .dinb(n1762), .dout(n2096));
  jor  g2021(.dina(n2096), .dinb(n2095), .dout(n2097));
  jor  g2022(.dina(n2097), .dinb(n2094), .dout(n2098));
  jnot g2023(.din(n2098), .dout(n2099));
  jand g2024(.dina(n2099), .dinb(n2091), .dout(n2100));
  jor  g2025(.dina(n2100), .dinb(n2090), .dout(n2101));
  jand g2026(.dina(n2101), .dinb(n2074), .dout(n2102));
  jxor g2027(.dina(n2101), .dinb(n2074), .dout(n2103));
  jxor g2028(.dina(n2065), .dinb(n2057), .dout(n2104));
  jand g2029(.dina(n2104), .dinb(n2103), .dout(n2105));
  jor  g2030(.dina(n2105), .dinb(n2102), .dout(n2106));
  jand g2031(.dina(n1356), .dinb(n58), .dout(n2107));
  jnot g2032(.din(n2107), .dout(n2108));
  jand g2033(.dina(n2108), .dinb(n1413), .dout(n2109));
  jand g2034(.dina(n1682), .dinb(n699), .dout(n2110));
  jand g2035(.dina(n2110), .dinb(n1283), .dout(n2111));
  jnot g2036(.din(n2111), .dout(n2112));
  jand g2037(.dina(n1283), .dinb(n1391), .dout(n2113));
  jor  g2038(.dina(n2113), .dinb(n2110), .dout(n2114));
  jor  g2039(.dina(n2114), .dinb(n1683), .dout(n2115));
  jand g2040(.dina(n2115), .dinb(n2112), .dout(n2116));
  jand g2041(.dina(n2116), .dinb(n2109), .dout(n2117));
  jand g2042(.dina(n2117), .dinb(n2011), .dout(n2118));
  jand g2043(.dina(n1420), .dinb(n1762), .dout(n2119));
  jand g2044(.dina(n1417), .dinb(n75), .dout(n2120));
  jor  g2045(.dina(n2120), .dinb(n2119), .dout(n2121));
  jand g2046(.dina(n1411), .dinb(n58), .dout(n2122));
  jand g2047(.dina(n1414), .dinb(n59), .dout(n2123));
  jor  g2048(.dina(n2123), .dinb(n2122), .dout(n2124));
  jand g2049(.dina(n2124), .dinb(n2121), .dout(n2125));
  jand g2050(.dina(n1566), .dinb(n1584), .dout(n2126));
  jand g2051(.dina(n1568), .dinb(n1347), .dout(n2127));
  jor  g2052(.dina(n2127), .dinb(n2126), .dout(n2128));
  jor  g2053(.dina(n1571), .dinb(n55), .dout(n2129));
  jor  g2054(.dina(n1576), .dinb(n56), .dout(n2130));
  jand g2055(.dina(n2130), .dinb(n2129), .dout(n2131));
  jand g2056(.dina(n2131), .dinb(n2128), .dout(n2132));
  jand g2057(.dina(n2132), .dinb(n2125), .dout(n2133));
  jxor g2058(.dina(n2116), .dinb(n2109), .dout(n2134));
  jxor g2059(.dina(n2132), .dinb(n2125), .dout(n2135));
  jand g2060(.dina(n2135), .dinb(n2134), .dout(n2136));
  jor  g2061(.dina(n2136), .dinb(n2133), .dout(n2137));
  jxor g2062(.dina(n2117), .dinb(n2011), .dout(n2138));
  jand g2063(.dina(n2138), .dinb(n2137), .dout(n2139));
  jor  g2064(.dina(n2139), .dinb(n2118), .dout(n2140));
  jxor g2065(.dina(n2138), .dinb(n2137), .dout(n2141));
  jand g2066(.dina(n1682), .dinb(n337), .dout(n2142));
  jand g2067(.dina(n2142), .dinb(n1283), .dout(n2143));
  jnot g2068(.din(n2143), .dout(n2144));
  jand g2069(.dina(n1584), .dinb(n1283), .dout(n2145));
  jor  g2070(.dina(n2145), .dinb(n2142), .dout(n2146));
  jor  g2071(.dina(n2146), .dinb(n1683), .dout(n2147));
  jand g2072(.dina(n2147), .dinb(n2144), .dout(n2148));
  jor  g2073(.dina(n1568), .dinb(n56), .dout(n2149));
  jor  g2074(.dina(n1566), .dinb(n55), .dout(n2150));
  jand g2075(.dina(n2150), .dinb(n2149), .dout(n2151));
  jor  g2076(.dina(n1576), .dinb(n1762), .dout(n2152));
  jor  g2077(.dina(n1571), .dinb(n75), .dout(n2153));
  jand g2078(.dina(n2153), .dinb(n2152), .dout(n2154));
  jand g2079(.dina(n2154), .dinb(n2151), .dout(n2155));
  jand g2080(.dina(n2155), .dinb(n2148), .dout(n2156));
  jand g2081(.dina(n1574), .dinb(n58), .dout(n2157));
  jnot g2082(.din(n2157), .dout(n2158));
  jand g2083(.dina(n2158), .dinb(n1340), .dout(n2159));
  jand g2084(.dina(n1682), .dinb(n1347), .dout(n2160));
  jnot g2085(.din(n2160), .dout(n2161));
  jor  g2086(.dina(n2161), .dinb(n1243), .dout(n2162));
  jand g2087(.dina(n1283), .dinb(n56), .dout(n2163));
  jor  g2088(.dina(n2163), .dinb(n2160), .dout(n2164));
  jor  g2089(.dina(n2164), .dinb(n1683), .dout(n2165));
  jand g2090(.dina(n2165), .dinb(n2162), .dout(n2166));
  jand g2091(.dina(n2166), .dinb(n2159), .dout(n2167));
  jxor g2092(.dina(n2155), .dinb(n2148), .dout(n2168));
  jand g2093(.dina(n2168), .dinb(n2167), .dout(n2169));
  jor  g2094(.dina(n2169), .dinb(n2156), .dout(n2170));
  jxor g2095(.dina(n2135), .dinb(n2134), .dout(n2171));
  jor  g2096(.dina(n2171), .dinb(n2170), .dout(n2172));
  jand g2097(.dina(n2171), .dinb(n2170), .dout(n2173));
  jand g2098(.dina(n1682), .dinb(n55), .dout(n2174));
  jnot g2099(.din(n2174), .dout(n2175));
  jor  g2100(.dina(n2175), .dinb(n1243), .dout(n2176));
  jand g2101(.dina(n1283), .dinb(n1762), .dout(n2177));
  jor  g2102(.dina(n2177), .dinb(n2174), .dout(n2178));
  jor  g2103(.dina(n2178), .dinb(n1683), .dout(n2179));
  jand g2104(.dina(n2179), .dinb(n2176), .dout(n2180));
  jnot g2105(.din(n1682), .dout(n2181));
  jor  g2106(.dina(n2181), .dinb(n1762), .dout(n2182));
  jand g2107(.dina(n1283), .dinb(n59), .dout(n2183));
  jand g2108(.dina(n2183), .dinb(n2182), .dout(n2184));
  jor  g2109(.dina(n2184), .dinb(n2180), .dout(n2185));
  jand g2110(.dina(n2184), .dinb(n2180), .dout(n2186));
  jand g2111(.dina(n2157), .dinb(n1575), .dout(n2187));
  jand g2112(.dina(n2187), .dinb(n1339), .dout(n2188));
  jor  g2113(.dina(n2188), .dinb(n2186), .dout(n2189));
  jand g2114(.dina(n2189), .dinb(n2185), .dout(n2190));
  jxor g2115(.dina(n2166), .dinb(n2159), .dout(n2191));
  jand g2116(.dina(n1571), .dinb(n59), .dout(n2192));
  jor  g2117(.dina(n2192), .dinb(n2187), .dout(n2193));
  jor  g2118(.dina(n1568), .dinb(n1762), .dout(n2194));
  jor  g2119(.dina(n1566), .dinb(n75), .dout(n2195));
  jand g2120(.dina(n2195), .dinb(n2194), .dout(n2196));
  jand g2121(.dina(n2196), .dinb(n2193), .dout(n2197));
  jand g2122(.dina(n2197), .dinb(n2191), .dout(n2198));
  jor  g2123(.dina(n2198), .dinb(n2190), .dout(n2199));
  jor  g2124(.dina(n2197), .dinb(n2191), .dout(n2200));
  jand g2125(.dina(n2200), .dinb(n2199), .dout(n2201));
  jor  g2126(.dina(n2201), .dinb(n2107), .dout(n2202));
  jand g2127(.dina(n2201), .dinb(n2107), .dout(n2203));
  jxor g2128(.dina(n2168), .dinb(n2167), .dout(n2204));
  jor  g2129(.dina(n2204), .dinb(n2203), .dout(n2205));
  jand g2130(.dina(n2205), .dinb(n2202), .dout(n2206));
  jor  g2131(.dina(n2206), .dinb(n2173), .dout(n2207));
  jand g2132(.dina(n2207), .dinb(n2172), .dout(n2208));
  jor  g2133(.dina(n2208), .dinb(n2141), .dout(n2209));
  jand g2134(.dina(n2208), .dinb(n2141), .dout(n2210));
  jxor g2135(.dina(n2099), .dinb(n2091), .dout(n2211));
  jor  g2136(.dina(n2211), .dinb(n2210), .dout(n2212));
  jand g2137(.dina(n2212), .dinb(n2209), .dout(n2213));
  jor  g2138(.dina(n2213), .dinb(n2140), .dout(n2214));
  jand g2139(.dina(n2213), .dinb(n2140), .dout(n2215));
  jxor g2140(.dina(n2104), .dinb(n2103), .dout(n2216));
  jor  g2141(.dina(n2216), .dinb(n2215), .dout(n2217));
  jand g2142(.dina(n2217), .dinb(n2214), .dout(n2218));
  jor  g2143(.dina(n2218), .dinb(n2106), .dout(n2219));
  jand g2144(.dina(n2218), .dinb(n2106), .dout(n2220));
  jxor g2145(.dina(n2071), .dinb(n2070), .dout(n2221));
  jor  g2146(.dina(n2221), .dinb(n2220), .dout(n2222));
  jand g2147(.dina(n2222), .dinb(n2219), .dout(n2223));
  jor  g2148(.dina(n2223), .dinb(n2073), .dout(n2224));
  jand g2149(.dina(n2223), .dinb(n2073), .dout(n2225));
  jxor g2150(.dina(n2037), .dinb(n2036), .dout(n2226));
  jor  g2151(.dina(n2226), .dinb(n2225), .dout(n2227));
  jand g2152(.dina(n2227), .dinb(n2224), .dout(n2228));
  jor  g2153(.dina(n2228), .dinb(n2039), .dout(n2229));
  jand g2154(.dina(n2228), .dinb(n2039), .dout(n2230));
  jxor g2155(.dina(n2008), .dinb(n2007), .dout(n2231));
  jor  g2156(.dina(n2231), .dinb(n2230), .dout(n2232));
  jand g2157(.dina(n2232), .dinb(n2229), .dout(n2233));
  jor  g2158(.dina(n2233), .dinb(n2010), .dout(n2234));
  jand g2159(.dina(n2233), .dinb(n2010), .dout(n2235));
  jxor g2160(.dina(n1959), .dinb(n1958), .dout(n2236));
  jor  g2161(.dina(n2236), .dinb(n2235), .dout(n2237));
  jand g2162(.dina(n2237), .dinb(n2234), .dout(n2238));
  jand g2163(.dina(n2238), .dinb(n1964), .dout(n2239));
  jor  g2164(.dina(n2239), .dinb(n1963), .dout(n2240));
  jxor g2165(.dina(n1921), .dinb(n1920), .dout(n2241));
  jand g2166(.dina(n2241), .dinb(n2240), .dout(n2242));
  jor  g2167(.dina(n2242), .dinb(n1922), .dout(n2243));
  jxor g2168(.dina(n1850), .dinb(n1849), .dout(n2244));
  jand g2169(.dina(n2244), .dinb(n2243), .dout(n2245));
  jor  g2170(.dina(n2245), .dinb(n1851), .dout(n2246));
  jxor g2171(.dina(n1815), .dinb(n1814), .dout(n2247));
  jand g2172(.dina(n2247), .dinb(n2246), .dout(n2248));
  jor  g2173(.dina(n2248), .dinb(n1816), .dout(n2249));
  jxor g2174(.dina(n1749), .dinb(n1748), .dout(n2250));
  jand g2175(.dina(n2250), .dinb(n2249), .dout(n2251));
  jor  g2176(.dina(n2251), .dinb(n1750), .dout(n2252));
  jxor g2177(.dina(n1635), .dinb(n1634), .dout(n2253));
  jand g2178(.dina(n2253), .dinb(n2252), .dout(n2254));
  jor  g2179(.dina(n2254), .dinb(n1636), .dout(n2255));
  jxor g2180(.dina(n1440), .dinb(n1439), .dout(n2256));
  jand g2181(.dina(n2256), .dinb(n2255), .dout(n2257));
  jor  g2182(.dina(n2257), .dinb(n1441), .dout(n2258));
  jxor g2183(.dina(n1389), .dinb(n1388), .dout(n2259));
  jand g2184(.dina(n2259), .dinb(n2258), .dout(n2260));
  jor  g2185(.dina(n2260), .dinb(n1390), .dout(n2261));
  jxor g2186(.dina(n1140), .dinb(n1113), .dout(n2262));
  jand g2187(.dina(n2262), .dinb(n2261), .dout(n2263));
  jor  g2188(.dina(n2263), .dinb(n1141), .dout(n2264));
  jand g2189(.dina(n1138), .dinb(n1133), .dout(n2265));
  jand g2190(.dina(n1139), .dinb(n1130), .dout(n2266));
  jor  g2191(.dina(n2266), .dinb(n2265), .dout(n2267));
  jand g2192(.dina(n1120), .dinb(n1115), .dout(n2268));
  jand g2193(.dina(n1129), .dinb(n1121), .dout(n2269));
  jor  g2194(.dina(n2269), .dinb(n2268), .dout(n2270));
  jor  g2195(.dina(n954), .dinb(n795), .dout(n2272));
  jor  g2196(.dina(n960), .dinb(n800), .dout(n2275));
  jor  g2197(.dina(n961), .dinb(n792), .dout(n2276));
  jand g2198(.dina(n2276), .dinb(n2275), .dout(n2277));
  jand g2199(.dina(n2277), .dinb(n2272), .dout(n2278));
  jxor g2200(.dina(n2278), .dinb(n2270), .dout(n2279));
  jxor g2201(.dina(n1115), .dinb(n1047), .dout(n2280));
  jand g2202(.dina(n980), .dinb(n335), .dout(n2281));
  jxor g2203(.dina(n2281), .dinb(n2280), .dout(n2282));
  jxor g2204(.dina(n2282), .dinb(n2279), .dout(n2283));
  jxor g2205(.dina(n2283), .dinb(n2267), .dout(n2284));
  jxor g2206(.dina(n2284), .dinb(n2264), .dout(n2285));
  jand g2207(.dina(n645), .dinb(n261), .dout(n2286));
  jand g2208(.dina(n356), .dinb(n310), .dout(n2287));
  jand g2209(.dina(n2287), .dinb(n2286), .dout(n2288));
  jand g2210(.dina(n445), .dinb(n365), .dout(n2289));
  jand g2211(.dina(n2289), .dinb(n504), .dout(n2290));
  jand g2212(.dina(n2290), .dinb(n2288), .dout(n2291));
  jand g2213(.dina(n781), .dinb(n732), .dout(n2292));
  jand g2214(.dina(n2292), .dinb(n470), .dout(n2293));
  jand g2215(.dina(n2293), .dinb(n917), .dout(n2294));
  jand g2216(.dina(n490), .dinb(n392), .dout(n2295));
  jand g2217(.dina(n2295), .dinb(n2294), .dout(n2296));
  jand g2218(.dina(n2296), .dinb(n2291), .dout(n2297));
  jand g2219(.dina(n991), .dinb(n675), .dout(n2298));
  jand g2220(.dina(n2298), .dinb(n2297), .dout(n2299));
  jand g2221(.dina(n2299), .dinb(n1203), .dout(n2300));
  jor  g2222(.dina(n2300), .dinb(n2285), .dout(n2301));
  jxor g2223(.dina(n2262), .dinb(n2261), .dout(n2302));
  jand g2224(.dina(n477), .dinb(n401), .dout(n2303));
  jand g2225(.dina(n2303), .dinb(n436), .dout(n2304));
  jand g2226(.dina(n734), .dinb(n368), .dout(n2305));
  jand g2227(.dina(n2305), .dinb(n507), .dout(n2306));
  jand g2228(.dina(n2306), .dinb(n2304), .dout(n2307));
  jand g2229(.dina(n312), .dinb(n216), .dout(n2308));
  jand g2230(.dina(n387), .dinb(n243), .dout(n2309));
  jand g2231(.dina(n2309), .dinb(n2308), .dout(n2310));
  jand g2232(.dina(n2310), .dinb(n1002), .dout(n2311));
  jand g2233(.dina(n2311), .dinb(n885), .dout(n2312));
  jand g2234(.dina(n2312), .dinb(n2307), .dout(n2313));
  jand g2235(.dina(n765), .dinb(n412), .dout(n2314));
  jand g2236(.dina(n2314), .dinb(n676), .dout(n2315));
  jand g2237(.dina(n561), .dinb(n363), .dout(n2316));
  jand g2238(.dina(n285), .dinb(n147), .dout(n2317));
  jand g2239(.dina(n2317), .dinb(n2316), .dout(n2318));
  jand g2240(.dina(n2318), .dinb(n2315), .dout(n2319));
  jand g2241(.dina(n757), .dinb(n254), .dout(n2320));
  jand g2242(.dina(n2320), .dinb(n138), .dout(n2321));
  jand g2243(.dina(n642), .dinb(n264), .dout(n2322));
  jand g2244(.dina(n2322), .dinb(n614), .dout(n2323));
  jand g2245(.dina(n2323), .dinb(n2321), .dout(n2324));
  jand g2246(.dina(n2324), .dinb(n2319), .dout(n2325));
  jand g2247(.dina(n668), .dinb(n356), .dout(n2326));
  jand g2248(.dina(n2326), .dinb(n1018), .dout(n2327));
  jand g2249(.dina(n2327), .dinb(n924), .dout(n2328));
  jand g2250(.dina(n2328), .dinb(n881), .dout(n2329));
  jand g2251(.dina(n2329), .dinb(n2325), .dout(n2330));
  jand g2252(.dina(n430), .dinb(n282), .dout(n2331));
  jand g2253(.dina(n2331), .dinb(n441), .dout(n2332));
  jand g2254(.dina(n849), .dinb(n358), .dout(n2333));
  jand g2255(.dina(n2333), .dinb(n473), .dout(n2334));
  jand g2256(.dina(n935), .dinb(n709), .dout(n2335));
  jand g2257(.dina(n2335), .dinb(n710), .dout(n2336));
  jand g2258(.dina(n2336), .dinb(n2334), .dout(n2337));
  jand g2259(.dina(n2337), .dinb(n2332), .dout(n2338));
  jand g2260(.dina(n853), .dinb(n488), .dout(n2339));
  jand g2261(.dina(n1025), .dinb(n822), .dout(n2340));
  jand g2262(.dina(n2340), .dinb(n2339), .dout(n2341));
  jand g2263(.dina(n2341), .dinb(n876), .dout(n2342));
  jand g2264(.dina(n2342), .dinb(n2338), .dout(n2343));
  jand g2265(.dina(n2343), .dinb(n2330), .dout(n2344));
  jand g2266(.dina(n2344), .dinb(n2313), .dout(n2345));
  jor  g2267(.dina(n2345), .dinb(n2302), .dout(n2346));
  jxor g2268(.dina(n2259), .dinb(n2258), .dout(n2347));
  jand g2269(.dina(n501), .dinb(n157), .dout(n2348));
  jand g2270(.dina(n2348), .dinb(n422), .dout(n2349));
  jand g2271(.dina(n2349), .dinb(n2330), .dout(n2350));
  jand g2272(.dina(n594), .dinb(n897), .dout(n2351));
  jand g2273(.dina(n532), .dinb(n270), .dout(n2352));
  jand g2274(.dina(n2352), .dinb(n2351), .dout(n2353));
  jand g2275(.dina(n2353), .dinb(n305), .dout(n2354));
  jand g2276(.dina(n993), .dinb(n451), .dout(n2355));
  jand g2277(.dina(n2355), .dinb(n372), .dout(n2356));
  jand g2278(.dina(n2356), .dinb(n741), .dout(n2357));
  jand g2279(.dina(n2357), .dinb(n2334), .dout(n2358));
  jand g2280(.dina(n2358), .dinb(n2354), .dout(n2359));
  jand g2281(.dina(n401), .dinb(n225), .dout(n2360));
  jand g2282(.dina(n732), .dinb(n1209), .dout(n2361));
  jand g2283(.dina(n763), .dinb(n837), .dout(n2362));
  jand g2284(.dina(n2362), .dinb(n2361), .dout(n2363));
  jand g2285(.dina(n2363), .dinb(n2360), .dout(n2364));
  jand g2286(.dina(n2364), .dinb(n912), .dout(n2365));
  jand g2287(.dina(n664), .dinb(n295), .dout(n2366));
  jand g2288(.dina(n282), .dinb(n251), .dout(n2367));
  jand g2289(.dina(n2367), .dinb(n2366), .dout(n2368));
  jand g2290(.dina(n619), .dinb(n597), .dout(n2369));
  jand g2291(.dina(n2369), .dinb(n2368), .dout(n2370));
  jand g2292(.dina(n477), .dinb(n445), .dout(n2371));
  jand g2293(.dina(n2371), .dinb(n499), .dout(n2372));
  jand g2294(.dina(n2372), .dinb(n1646), .dout(n2373));
  jand g2295(.dina(n2373), .dinb(n2370), .dout(n2374));
  jand g2296(.dina(n2374), .dinb(n2365), .dout(n2375));
  jand g2297(.dina(n2375), .dinb(n2359), .dout(n2376));
  jand g2298(.dina(n2376), .dinb(n2350), .dout(n2377));
  jor  g2299(.dina(n2377), .dinb(n2347), .dout(n2378));
  jxor g2300(.dina(n2256), .dinb(n2255), .dout(n2379));
  jnot g2301(.din(n893), .dout(n2380));
  jand g2302(.dina(n2380), .dinb(n370), .dout(n2381));
  jand g2303(.dina(n2381), .dinb(n1169), .dout(n2382));
  jand g2304(.dina(n732), .dinb(n730), .dout(n2383));
  jand g2305(.dina(n2383), .dinb(n1204), .dout(n2384));
  jand g2306(.dina(n461), .dinb(n130), .dout(n2385));
  jand g2307(.dina(n2385), .dinb(n1025), .dout(n2386));
  jand g2308(.dina(n477), .dinb(n303), .dout(n2387));
  jand g2309(.dina(n2387), .dinb(n301), .dout(n2388));
  jand g2310(.dina(n2388), .dinb(n2386), .dout(n2389));
  jand g2311(.dina(n2389), .dinb(n2384), .dout(n2390));
  jand g2312(.dina(n2390), .dinb(n1179), .dout(n2391));
  jand g2313(.dina(n470), .dinb(n243), .dout(n2392));
  jand g2314(.dina(n668), .dinb(n222), .dout(n2393));
  jand g2315(.dina(n2393), .dinb(n2392), .dout(n2394));
  jnot g2316(.din(n1675), .dout(n2395));
  jand g2317(.dina(n763), .dinb(n312), .dout(n2396));
  jand g2318(.dina(n2396), .dinb(n2395), .dout(n2397));
  jand g2319(.dina(n2397), .dinb(n2394), .dout(n2398));
  jand g2320(.dina(n679), .dinb(n421), .dout(n2399));
  jand g2321(.dina(n744), .dinb(n294), .dout(n2400));
  jand g2322(.dina(n2400), .dinb(n383), .dout(n2401));
  jand g2323(.dina(n2401), .dinb(n2399), .dout(n2402));
  jand g2324(.dina(n614), .dinb(n138), .dout(n2403));
  jand g2325(.dina(n768), .dinb(n229), .dout(n2404));
  jand g2326(.dina(n2404), .dinb(n2403), .dout(n2405));
  jand g2327(.dina(n430), .dinb(n323), .dout(n2406));
  jand g2328(.dina(n2406), .dinb(n740), .dout(n2407));
  jand g2329(.dina(n2407), .dinb(n2405), .dout(n2408));
  jand g2330(.dina(n2408), .dinb(n2402), .dout(n2409));
  jand g2331(.dina(n2409), .dinb(n2398), .dout(n2410));
  jand g2332(.dina(n2410), .dinb(n2391), .dout(n2411));
  jand g2333(.dina(n2411), .dinb(n2382), .dout(n2412));
  jor  g2334(.dina(n2412), .dinb(n2379), .dout(n2413));
  jxor g2335(.dina(n2253), .dinb(n2252), .dout(n2414));
  jand g2336(.dina(n458), .dinb(n387), .dout(n2415));
  jand g2337(.dina(n2415), .dinb(n724), .dout(n2416));
  jand g2338(.dina(n2416), .dinb(n767), .dout(n2417));
  jand g2339(.dina(n992), .dinb(n524), .dout(n2418));
  jand g2340(.dina(n2418), .dinb(n286), .dout(n2419));
  jand g2341(.dina(n2419), .dinb(n2417), .dout(n2420));
  jand g2342(.dina(n2420), .dinb(n538), .dout(n2421));
  jand g2343(.dina(n662), .dinb(n772), .dout(n2422));
  jand g2344(.dina(n2422), .dinb(n523), .dout(n2423));
  jand g2345(.dina(n2380), .dinb(n679), .dout(n2424));
  jand g2346(.dina(n2424), .dinb(n1170), .dout(n2425));
  jand g2347(.dina(n2425), .dinb(n2423), .dout(n2426));
  jand g2348(.dina(n2426), .dinb(n424), .dout(n2427));
  jand g2349(.dina(n402), .dinb(n371), .dout(n2428));
  jand g2350(.dina(n744), .dinb(n222), .dout(n2429));
  jand g2351(.dina(n592), .dinb(n383), .dout(n2430));
  jand g2352(.dina(n2430), .dinb(n2429), .dout(n2431));
  jnot g2353(.din(n1214), .dout(n2432));
  jand g2354(.dina(n2432), .dinb(n324), .dout(n2433));
  jand g2355(.dina(n2433), .dinb(n2431), .dout(n2434));
  jand g2356(.dina(n2434), .dinb(n2428), .dout(n2435));
  jand g2357(.dina(n2435), .dinb(n2427), .dout(n2436));
  jand g2358(.dina(n2436), .dinb(n2421), .dout(n2437));
  jand g2359(.dina(n2437), .dinb(n630), .dout(n2438));
  jor  g2360(.dina(n2438), .dinb(n2414), .dout(n2439));
  jxor g2361(.dina(n2250), .dinb(n2249), .dout(n2440));
  jand g2362(.dina(n918), .dinb(n532), .dout(n2441));
  jand g2363(.dina(n2441), .dinb(n2385), .dout(n2442));
  jand g2364(.dina(n744), .dinb(n612), .dout(n2443));
  jand g2365(.dina(n579), .dinb(n304), .dout(n2444));
  jand g2366(.dina(n2444), .dinb(n2443), .dout(n2445));
  jand g2367(.dina(n2445), .dinb(n987), .dout(n2446));
  jand g2368(.dina(n2446), .dinb(n2442), .dout(n2447));
  jand g2369(.dina(n1332), .dinb(n881), .dout(n2448));
  jand g2370(.dina(n2448), .dinb(n2447), .dout(n2449));
  jand g2371(.dina(n822), .dinb(n397), .dout(n2450));
  jand g2372(.dina(n2450), .dinb(n2449), .dout(n2451));
  jand g2373(.dina(n853), .dinb(n264), .dout(n2452));
  jand g2374(.dina(n2452), .dinb(n739), .dout(n2453));
  jand g2375(.dina(n348), .dinb(n897), .dout(n2454));
  jand g2376(.dina(n2454), .dinb(n643), .dout(n2455));
  jand g2377(.dina(n445), .dinb(n323), .dout(n2456));
  jand g2378(.dina(n381), .dinb(n279), .dout(n2457));
  jand g2379(.dina(n2457), .dinb(n2456), .dout(n2458));
  jand g2380(.dina(n2458), .dinb(n2455), .dout(n2459));
  jand g2381(.dina(n2459), .dinb(n2453), .dout(n2460));
  jand g2382(.dina(n2460), .dinb(n509), .dout(n2461));
  jand g2383(.dina(n837), .dinb(n282), .dout(n2462));
  jand g2384(.dina(n751), .dinb(n216), .dout(n2463));
  jand g2385(.dina(n2463), .dinb(n2462), .dout(n2464));
  jand g2386(.dina(n2287), .dinb(n301), .dout(n2465));
  jand g2387(.dina(n2465), .dinb(n2464), .dout(n2466));
  jand g2388(.dina(n742), .dinb(n427), .dout(n2467));
  jand g2389(.dina(n295), .dinb(n285), .dout(n2468));
  jand g2390(.dina(n2468), .dinb(n2467), .dout(n2469));
  jnot g2391(.din(n346), .dout(n2470));
  jand g2392(.dina(n2470), .dinb(n325), .dout(n2471));
  jor  g2393(.dina(n2471), .dinb(n326), .dout(n2472));
  jand g2394(.dina(n2472), .dinb(n417), .dout(n2473));
  jand g2395(.dina(n2473), .dinb(n2469), .dout(n2474));
  jand g2396(.dina(n2474), .dinb(n2466), .dout(n2475));
  jand g2397(.dina(n2475), .dinb(n2461), .dout(n2476));
  jand g2398(.dina(n2476), .dinb(n2451), .dout(n2477));
  jor  g2399(.dina(n2477), .dinb(n2440), .dout(n2478));
  jxor g2400(.dina(n2247), .dinb(n2246), .dout(n2479));
  jand g2401(.dina(n2380), .dinb(n612), .dout(n2480));
  jand g2402(.dina(n665), .dinb(n772), .dout(n2481));
  jand g2403(.dina(n2481), .dinb(n2480), .dout(n2482));
  jand g2404(.dina(n2482), .dinb(n507), .dout(n2483));
  jand g2405(.dina(n2332), .dinb(n836), .dout(n2484));
  jand g2406(.dina(n2484), .dinb(n234), .dout(n2485));
  jand g2407(.dina(n2485), .dinb(n2483), .dout(n2486));
  jand g2408(.dina(n853), .dinb(n925), .dout(n2487));
  jand g2409(.dina(n2487), .dinb(n501), .dout(n2488));
  jand g2410(.dina(n668), .dinb(n138), .dout(n2489));
  jand g2411(.dina(n624), .dinb(n294), .dout(n2490));
  jand g2412(.dina(n2490), .dinb(n2489), .dout(n2491));
  jand g2413(.dina(n2491), .dinb(n2488), .dout(n2492));
  jand g2414(.dina(n2492), .dinb(n611), .dout(n2493));
  jnot g2415(.din(n1215), .dout(n2494));
  jand g2416(.dina(n642), .dinb(n768), .dout(n2495));
  jand g2417(.dina(n2495), .dinb(n2494), .dout(n2496));
  jand g2418(.dina(n1022), .dinb(n265), .dout(n2497));
  jand g2419(.dina(n2497), .dinb(n2496), .dout(n2498));
  jand g2420(.dina(n2335), .dinb(n821), .dout(n2499));
  jand g2421(.dina(n2499), .dinb(n869), .dout(n2500));
  jand g2422(.dina(n2500), .dinb(n2498), .dout(n2501));
  jand g2423(.dina(n2501), .dinb(n2493), .dout(n2502));
  jand g2424(.dina(n2502), .dinb(n2486), .dout(n2503));
  jand g2425(.dina(n2503), .dinb(n395), .dout(n2504));
  jor  g2426(.dina(n2504), .dinb(n2479), .dout(n2505));
  jxor g2427(.dina(n2244), .dinb(n2243), .dout(n2506));
  jand g2428(.dina(n612), .dinb(n427), .dout(n2507));
  jand g2429(.dina(n2507), .dinb(n987), .dout(n2508));
  jand g2430(.dina(n2508), .dinb(n605), .dout(n2509));
  jand g2431(.dina(n2509), .dinb(n2372), .dout(n2510));
  jand g2432(.dina(n993), .dinb(n837), .dout(n2511));
  jand g2433(.dina(n710), .dinb(n594), .dout(n2512));
  jand g2434(.dina(n2512), .dinb(n734), .dout(n2513));
  jand g2435(.dina(n2513), .dinb(n2511), .dout(n2514));
  jand g2436(.dina(n739), .dinb(n501), .dout(n2515));
  jand g2437(.dina(n2515), .dinb(n680), .dout(n2516));
  jand g2438(.dina(n2516), .dinb(n1328), .dout(n2517));
  jand g2439(.dina(n2517), .dinb(n2417), .dout(n2518));
  jand g2440(.dina(n2518), .dinb(n2514), .dout(n2519));
  jand g2441(.dina(n2519), .dinb(n2510), .dout(n2520));
  jand g2442(.dina(n374), .dinb(n343), .dout(n2521));
  jand g2443(.dina(n2521), .dinb(n597), .dout(n2522));
  jand g2444(.dina(n2522), .dinb(n938), .dout(n2523));
  jand g2445(.dina(n368), .dinb(n267), .dout(n2524));
  jand g2446(.dina(n2524), .dinb(n410), .dout(n2525));
  jand g2447(.dina(n665), .dinb(n614), .dout(n2526));
  jand g2448(.dina(n2526), .dinb(n305), .dout(n2527));
  jand g2449(.dina(n2527), .dinb(n2525), .dout(n2528));
  jand g2450(.dina(n2528), .dinb(n2523), .dout(n2529));
  jand g2451(.dina(n2498), .dinb(n622), .dout(n2530));
  jand g2452(.dina(n2530), .dinb(n2529), .dout(n2531));
  jand g2453(.dina(n2531), .dinb(n497), .dout(n2532));
  jand g2454(.dina(n2532), .dinb(n832), .dout(n2533));
  jand g2455(.dina(n2533), .dinb(n2520), .dout(n2534));
  jor  g2456(.dina(n2534), .dinb(n2506), .dout(n2535));
  jxor g2457(.dina(n2241), .dinb(n2240), .dout(n2536));
  jand g2458(.dina(n825), .dinb(n310), .dout(n2537));
  jand g2459(.dina(n765), .dinb(n251), .dout(n2538));
  jand g2460(.dina(n2538), .dinb(n918), .dout(n2539));
  jand g2461(.dina(n2539), .dinb(n2537), .dout(n2540));
  jand g2462(.dina(n1210), .dinb(n730), .dout(n2541));
  jand g2463(.dina(n853), .dinb(n312), .dout(n2542));
  jand g2464(.dina(n2542), .dinb(n157), .dout(n2543));
  jand g2465(.dina(n2543), .dinb(n2541), .dout(n2544));
  jand g2466(.dina(n353), .dinb(n220), .dout(n2545));
  jor  g2467(.dina(n2545), .dinb(n748), .dout(n2546));
  jnot g2468(.din(n2546), .dout(n2547));
  jand g2469(.dina(n732), .dinb(n451), .dout(n2548));
  jand g2470(.dina(n2548), .dinb(n2547), .dout(n2549));
  jand g2471(.dina(n2549), .dinb(n2544), .dout(n2550));
  jand g2472(.dina(n2550), .dinb(n2540), .dout(n2551));
  jand g2473(.dina(n291), .dinb(n254), .dout(n2552));
  jand g2474(.dina(n2552), .dinb(n2515), .dout(n2553));
  jand g2475(.dina(n2553), .dinb(n646), .dout(n2554));
  jand g2476(.dina(n878), .dinb(n243), .dout(n2555));
  jand g2477(.dina(n430), .dinb(n303), .dout(n2556));
  jand g2478(.dina(n2556), .dinb(n2555), .dout(n2557));
  jand g2479(.dina(n751), .dinb(n763), .dout(n2558));
  jand g2480(.dina(n2558), .dinb(n626), .dout(n2559));
  jand g2481(.dina(n2559), .dinb(n2557), .dout(n2560));
  jand g2482(.dina(n2560), .dinb(n942), .dout(n2561));
  jand g2483(.dina(n2561), .dinb(n2554), .dout(n2562));
  jand g2484(.dina(n2562), .dinb(n2427), .dout(n2563));
  jand g2485(.dina(n2563), .dinb(n2551), .dout(n2564));
  jor  g2486(.dina(n2564), .dinb(n2536), .dout(n2565));
  jxor g2487(.dina(n2238), .dinb(n1964), .dout(n2566));
  jand g2488(.dina(n1189), .dinb(n385), .dout(n2567));
  jand g2489(.dina(n2315), .dinb(n611), .dout(n2568));
  jand g2490(.dina(n2568), .dinb(n2567), .dout(n2569));
  jand g2491(.dina(n2286), .dinb(n365), .dout(n2570));
  jand g2492(.dina(n2570), .dinb(n1000), .dout(n2571));
  jand g2493(.dina(n854), .dinb(n515), .dout(n2572));
  jand g2494(.dina(n2572), .dinb(n417), .dout(n2573));
  jand g2495(.dina(n2573), .dinb(n2571), .dout(n2574));
  jand g2496(.dina(n2574), .dinb(n2569), .dout(n2575));
  jand g2497(.dina(n1193), .dinb(n439), .dout(n2576));
  jand g2498(.dina(n2576), .dinb(n392), .dout(n2577));
  jand g2499(.dina(n993), .dinb(n216), .dout(n2578));
  jand g2500(.dina(n2578), .dinb(n781), .dout(n2579));
  jand g2501(.dina(n878), .dinb(n563), .dout(n2580));
  jand g2502(.dina(n2580), .dinb(n987), .dout(n2581));
  jand g2503(.dina(n2581), .dinb(n2579), .dout(n2582));
  jand g2504(.dina(n2582), .dinb(n513), .dout(n2583));
  jand g2505(.dina(n2583), .dinb(n2577), .dout(n2584));
  jand g2506(.dina(n2584), .dinb(n2575), .dout(n2585));
  jand g2507(.dina(n2585), .dinb(n2486), .dout(n2586));
  jand g2508(.dina(n2586), .dinb(n2566), .dout(n2587));
  jnot g2509(.din(n2564), .dout(n2588));
  jxor g2510(.dina(n2588), .dinb(n2536), .dout(n2589));
  jor  g2511(.dina(n2589), .dinb(n2587), .dout(n2590));
  jand g2512(.dina(n2590), .dinb(n2565), .dout(n2591));
  jnot g2513(.din(n2534), .dout(n2592));
  jxor g2514(.dina(n2592), .dinb(n2506), .dout(n2593));
  jor  g2515(.dina(n2593), .dinb(n2591), .dout(n2594));
  jand g2516(.dina(n2594), .dinb(n2535), .dout(n2595));
  jnot g2517(.din(n2504), .dout(n2596));
  jxor g2518(.dina(n2596), .dinb(n2479), .dout(n2597));
  jor  g2519(.dina(n2597), .dinb(n2595), .dout(n2598));
  jand g2520(.dina(n2598), .dinb(n2505), .dout(n2599));
  jxor g2521(.dina(n2477), .dinb(n2440), .dout(n2600));
  jnot g2522(.din(n2600), .dout(n2601));
  jor  g2523(.dina(n2601), .dinb(n2599), .dout(n2602));
  jand g2524(.dina(n2602), .dinb(n2478), .dout(n2603));
  jxor g2525(.dina(n2438), .dinb(n2414), .dout(n2604));
  jnot g2526(.din(n2604), .dout(n2605));
  jor  g2527(.dina(n2605), .dinb(n2603), .dout(n2606));
  jand g2528(.dina(n2606), .dinb(n2439), .dout(n2607));
  jxor g2529(.dina(n2412), .dinb(n2379), .dout(n2608));
  jnot g2530(.din(n2608), .dout(n2609));
  jor  g2531(.dina(n2609), .dinb(n2607), .dout(n2610));
  jand g2532(.dina(n2610), .dinb(n2413), .dout(n2611));
  jxor g2533(.dina(n2377), .dinb(n2347), .dout(n2612));
  jnot g2534(.din(n2612), .dout(n2613));
  jor  g2535(.dina(n2613), .dinb(n2611), .dout(n2614));
  jand g2536(.dina(n2614), .dinb(n2378), .dout(n2615));
  jnot g2537(.din(n2615), .dout(n2616));
  jxor g2538(.dina(n2345), .dinb(n2302), .dout(n2617));
  jand g2539(.dina(n2617), .dinb(n2616), .dout(n2618));
  jnot g2540(.din(n2618), .dout(n2619));
  jand g2541(.dina(n2619), .dinb(n2346), .dout(n2620));
  jxor g2542(.dina(n2300), .dinb(n2285), .dout(n2621));
  jnot g2543(.din(n2621), .dout(n2622));
  jor  g2544(.dina(n2622), .dinb(n2620), .dout(n2623));
  jand g2545(.dina(n2623), .dinb(n2301), .dout(n2624));
  jand g2546(.dina(n2283), .dinb(n2267), .dout(n2625));
  jand g2547(.dina(n2284), .dinb(n2264), .dout(n2626));
  jor  g2548(.dina(n2626), .dinb(n2625), .dout(n2627));
  jand g2549(.dina(n2278), .dinb(n2270), .dout(n2628));
  jand g2550(.dina(n2282), .dinb(n2279), .dout(n2629));
  jor  g2551(.dina(n2629), .dinb(n2628), .dout(n2630));
  jand g2552(.dina(n2281), .dinb(n2280), .dout(n2632));
  jor  g2553(.dina(n2632), .dinb(n1114), .dout(n2633));
  jand g2554(.dina(n960), .dinb(n335), .dout(n2634));
  jand g2555(.dina(n954), .dinb(n795), .dout(n2635));
  jor  g2556(.dina(n2635), .dinb(n335), .dout(n2636));
  jand g2557(.dina(n954), .dinb(n804), .dout(n2637));
  jnot g2558(.din(n2637), .dout(n2638));
  jand g2559(.dina(n2638), .dinb(n2636), .dout(n2639));
  jnot g2560(.din(n2639), .dout(n2640));
  jxor g2561(.dina(n2640), .dinb(n2634), .dout(n2641));
  jxor g2562(.dina(n2641), .dinb(n2633), .dout(n2642));
  jxor g2563(.dina(n2642), .dinb(n2630), .dout(n2643));
  jxor g2564(.dina(n2643), .dinb(n2627), .dout(n2644));
  jand g2565(.dina(n936), .dinb(n158), .dout(n2645));
  jand g2566(.dina(n1022), .dinb(n280), .dout(n2646));
  jand g2567(.dina(n2646), .dinb(n2645), .dout(n2647));
  jand g2568(.dina(n614), .dinb(n422), .dout(n2648));
  jand g2569(.dina(n374), .dinb(n294), .dout(n2649));
  jand g2570(.dina(n2649), .dinb(n2648), .dout(n2650));
  jand g2571(.dina(n2650), .dinb(n2321), .dout(n2651));
  jand g2572(.dina(n2651), .dinb(n2647), .dout(n2652));
  jand g2573(.dina(n2652), .dinb(n482), .dout(n2653));
  jand g2574(.dina(n2653), .dinb(n2365), .dout(n2654));
  jand g2575(.dina(n781), .dinb(n709), .dout(n2655));
  jand g2576(.dina(n642), .dinb(n436), .dout(n2656));
  jand g2577(.dina(n2656), .dinb(n2380), .dout(n2657));
  jand g2578(.dina(n2657), .dinb(n2655), .dout(n2658));
  jand g2579(.dina(n624), .dinb(n535), .dout(n2659));
  jand g2580(.dina(n2659), .dinb(n563), .dout(n2660));
  jand g2581(.dina(n363), .dinb(n214), .dout(n2661));
  jand g2582(.dina(n2661), .dinb(n388), .dout(n2662));
  jand g2583(.dina(n2662), .dinb(n428), .dout(n2663));
  jand g2584(.dina(n2663), .dinb(n2660), .dout(n2664));
  jand g2585(.dina(n2664), .dinb(n2658), .dout(n2665));
  jand g2586(.dina(n2665), .dinb(n2575), .dout(n2666));
  jand g2587(.dina(n2666), .dinb(n2654), .dout(n2667));
  jxor g2588(.dina(n2667), .dinb(n2644), .dout(n2668));
  jxor g2589(.dina(n2668), .dinb(n2624), .dout(n2669));
  jnot g2590(.din(n2669), .dout(n2670));
  jxor g2591(.dina(n2621), .dinb(n2620), .dout(n2671));
  jnot g2592(.din(n2671), .dout(n2672));
  jand g2593(.dina(n2672), .dinb(n2670), .dout(n2673));
  jxor g2594(.dina(n2617), .dinb(n2615), .dout(n2674));
  jor  g2595(.dina(n2674), .dinb(n2671), .dout(n2675));
  jnot g2596(.din(n2675), .dout(n2676));
  jnot g2597(.din(n2674), .dout(n2677));
  jxor g2598(.dina(n2612), .dinb(n2611), .dout(n2678));
  jnot g2599(.din(n2678), .dout(n2679));
  jand g2600(.dina(n2679), .dinb(n2677), .dout(n2680));
  jxor g2601(.dina(n2608), .dinb(n2607), .dout(n2681));
  jor  g2602(.dina(n2681), .dinb(n2678), .dout(n2682));
  jnot g2603(.din(n2682), .dout(n2683));
  jnot g2604(.din(n2681), .dout(n2684));
  jxor g2605(.dina(n2605), .dinb(n2603), .dout(n2685));
  jand g2606(.dina(n2685), .dinb(n2684), .dout(n2686));
  jxor g2607(.dina(n2604), .dinb(n2603), .dout(n2687));
  jxor g2608(.dina(n2600), .dinb(n2599), .dout(n2688));
  jor  g2609(.dina(n2688), .dinb(n2687), .dout(n2689));
  jxor g2610(.dina(n2504), .dinb(n2479), .dout(n2690));
  jxor g2611(.dina(n2690), .dinb(n2595), .dout(n2691));
  jor  g2612(.dina(n2691), .dinb(n2688), .dout(n2692));
  jxor g2613(.dina(n2593), .dinb(n2591), .dout(n2693));
  jnot g2614(.din(n2693), .dout(n2694));
  jor  g2615(.dina(n2694), .dinb(n2691), .dout(n2695));
  jxor g2616(.dina(n2693), .dinb(n2691), .dout(n2696));
  jxor g2617(.dina(n2586), .dinb(n2566), .dout(n2697));
  jnot g2618(.din(n2697), .dout(n2698));
  jor  g2619(.dina(n2698), .dinb(n2693), .dout(n2699));
  jxor g2620(.dina(n2589), .dinb(n2587), .dout(n2700));
  jand g2621(.dina(n2700), .dinb(n2699), .dout(n2701));
  jnot g2622(.din(n2701), .dout(n2702));
  jor  g2623(.dina(n2702), .dinb(n2696), .dout(n2703));
  jand g2624(.dina(n2703), .dinb(n2695), .dout(n2704));
  jxor g2625(.dina(n2691), .dinb(n2688), .dout(n2705));
  jnot g2626(.din(n2705), .dout(n2706));
  jor  g2627(.dina(n2706), .dinb(n2704), .dout(n2707));
  jand g2628(.dina(n2707), .dinb(n2692), .dout(n2708));
  jxor g2629(.dina(n2688), .dinb(n2685), .dout(n2709));
  jor  g2630(.dina(n2709), .dinb(n2708), .dout(n2710));
  jand g2631(.dina(n2710), .dinb(n2689), .dout(n2711));
  jnot g2632(.din(n2711), .dout(n2712));
  jxor g2633(.dina(n2687), .dinb(n2681), .dout(n2713));
  jand g2634(.dina(n2713), .dinb(n2712), .dout(n2714));
  jor  g2635(.dina(n2714), .dinb(n2686), .dout(n2715));
  jxor g2636(.dina(n2681), .dinb(n2678), .dout(n2716));
  jand g2637(.dina(n2716), .dinb(n2715), .dout(n2717));
  jor  g2638(.dina(n2717), .dinb(n2683), .dout(n2718));
  jxor g2639(.dina(n2678), .dinb(n2674), .dout(n2719));
  jand g2640(.dina(n2719), .dinb(n2718), .dout(n2720));
  jor  g2641(.dina(n2720), .dinb(n2680), .dout(n2721));
  jxor g2642(.dina(n2674), .dinb(n2671), .dout(n2722));
  jand g2643(.dina(n2722), .dinb(n2721), .dout(n2723));
  jor  g2644(.dina(n2723), .dinb(n2676), .dout(n2724));
  jxor g2645(.dina(n2671), .dinb(n2669), .dout(n2725));
  jand g2646(.dina(n2725), .dinb(n2724), .dout(n2726));
  jor  g2647(.dina(n2726), .dinb(n2673), .dout(n2727));
  jnot g2648(.din(n2727), .dout(n2728));
  jor  g2649(.dina(n2667), .dinb(n2644), .dout(n2729));
  jnot g2650(.din(n2729), .dout(n2730));
  jnot g2651(.din(n2624), .dout(n2731));
  jand g2652(.dina(n2668), .dinb(n2731), .dout(n2732));
  jor  g2653(.dina(n2732), .dinb(n2730), .dout(n2733));
  jand g2654(.dina(n458), .dinb(n153), .dout(n2734));
  jand g2655(.dina(n2734), .dinb(n597), .dout(n2735));
  jand g2656(.dina(n925), .dinb(n410), .dout(n2736));
  jand g2657(.dina(n2736), .dinb(n731), .dout(n2737));
  jand g2658(.dina(n2552), .dinb(n992), .dout(n2738));
  jand g2659(.dina(n2738), .dinb(n2737), .dout(n2739));
  jand g2660(.dina(n2739), .dinb(n2735), .dout(n2740));
  jand g2661(.dina(n2380), .dinb(n279), .dout(n2741));
  jand g2662(.dina(n2741), .dinb(n470), .dout(n2742));
  jand g2663(.dina(n2742), .dinb(n2323), .dout(n2743));
  jand g2664(.dina(n935), .dinb(n633), .dout(n2744));
  jand g2665(.dina(n2744), .dinb(n2351), .dout(n2745));
  jand g2666(.dina(n2745), .dinb(n2743), .dout(n2746));
  jand g2667(.dina(n2746), .dinb(n2740), .dout(n2747));
  jand g2668(.dina(n1231), .dinb(n497), .dout(n2748));
  jand g2669(.dina(n2748), .dinb(n2747), .dout(n2749));
  jand g2670(.dina(n2749), .dinb(n2451), .dout(n2750));
  jxor g2671(.dina(n960), .dinb(n820), .dout(n2751));
  jnot g2672(.din(n2751), .dout(n2752));
  jand g2673(.dina(n2752), .dinb(n796), .dout(n2753));
  jnot g2674(.din(n2753), .dout(n2754));
  jand g2675(.dina(n335), .dinb(n2754), .dout(n2757));
  jand g2676(.dina(n2642), .dinb(n2630), .dout(n2758));
  jand g2677(.dina(n2643), .dinb(n2627), .dout(n2759));
  jor  g2678(.dina(n2759), .dinb(n2758), .dout(n2760));
  jor  g2679(.dina(n2640), .dinb(n2634), .dout(n2761));
  jnot g2680(.din(n2633), .dout(n2762));
  jnot g2681(.din(n2641), .dout(n2763));
  jor  g2682(.dina(n2763), .dinb(n2762), .dout(n2764));
  jand g2683(.dina(n2764), .dinb(n2761), .dout(n2765));
  jxor g2684(.dina(n2765), .dinb(n2760), .dout(n2766));
  jxor g2685(.dina(n2766), .dinb(n2757), .dout(n2767));
  jxor g2686(.dina(n2767), .dinb(n2750), .dout(n2768));
  jxor g2687(.dina(n2768), .dinb(n2733), .dout(n2769));
  jxor g2688(.dina(n2769), .dinb(n2670), .dout(n2770));
  jxor g2689(.dina(n2770), .dinb(n2728), .dout(n2771));
  jor  g2690(.dina(n2771), .dinb(n79), .dout(n2772));
  jnot g2691(.din(n2769), .dout(n2773));
  jand g2692(.dina(n76), .dinb(n70), .dout(n2774));
  jnot g2693(.din(n2774), .dout(n2775));
  jor  g2694(.dina(n2775), .dinb(n2773), .dout(n2776));
  jxor g2695(.dina(n75), .dinb(n59), .dout(n2777));
  jnot g2696(.din(n2777), .dout(n2778));
  jand g2697(.dina(n2778), .dinb(n69), .dout(n2779));
  jnot g2698(.din(n2779), .dout(n2780));
  jor  g2699(.dina(n2780), .dinb(n2669), .dout(n2781));
  jand g2700(.dina(n77), .dinb(n69), .dout(n2782));
  jand g2701(.dina(n2782), .dinb(n2777), .dout(n2783));
  jnot g2702(.din(n2783), .dout(n2784));
  jor  g2703(.dina(n2784), .dinb(n2671), .dout(n2785));
  jand g2704(.dina(n2785), .dinb(n2781), .dout(n2786));
  jand g2705(.dina(n2786), .dinb(n2776), .dout(n2787));
  jand g2706(.dina(n2787), .dinb(n2772), .dout(n2788));
  jxor g2707(.dina(n2788), .dinb(n56), .dout(n2789));
  jxor g2708(.dina(n1347), .dinb(n56), .dout(n2790));
  jnot g2709(.din(n2790), .dout(n2791));
  jxor g2710(.dina(n699), .dinb(n1391), .dout(n2792));
  jnot g2711(.din(n2792), .dout(n2793));
  jand g2712(.dina(n2793), .dinb(n2791), .dout(n2794));
  jnot g2713(.din(n2794), .dout(n2795));
  jxor g2714(.dina(n2684), .dinb(n2678), .dout(n2796));
  jxor g2715(.dina(n2796), .dinb(n2715), .dout(n2797));
  jor  g2716(.dina(n2797), .dinb(n2795), .dout(n2798));
  jand g2717(.dina(n2792), .dinb(n2791), .dout(n2799));
  jnot g2718(.din(n2799), .dout(n2800));
  jor  g2719(.dina(n2800), .dinb(n2678), .dout(n2801));
  jxor g2720(.dina(n1347), .dinb(n1391), .dout(n2802));
  jnot g2721(.din(n2802), .dout(n2803));
  jand g2722(.dina(n2803), .dinb(n2790), .dout(n2804));
  jnot g2723(.din(n2804), .dout(n2805));
  jor  g2724(.dina(n2805), .dinb(n2681), .dout(n2806));
  jand g2725(.dina(n2802), .dinb(n2790), .dout(n2807));
  jand g2726(.dina(n2807), .dinb(n2793), .dout(n2808));
  jnot g2727(.din(n2808), .dout(n2809));
  jor  g2728(.dina(n2809), .dinb(n2687), .dout(n2810));
  jand g2729(.dina(n2810), .dinb(n2806), .dout(n2811));
  jand g2730(.dina(n2811), .dinb(n2801), .dout(n2812));
  jand g2731(.dina(n2812), .dinb(n2798), .dout(n2813));
  jxor g2732(.dina(n2813), .dinb(n699), .dout(n2814));
  jnot g2733(.din(n2814), .dout(n2815));
  jxor g2734(.dina(n980), .dinb(n808), .dout(n2816));
  jnot g2735(.din(n2816), .dout(n2817));
  jand g2736(.dina(n2817), .dinb(n2698), .dout(n2818));
  jor  g2737(.dina(n2700), .dinb(n2697), .dout(n2819));
  jand g2738(.dina(n2697), .dinb(n2589), .dout(n2820));
  jnot g2739(.din(n2820), .dout(n2821));
  jand g2740(.dina(n2821), .dinb(n2819), .dout(n2822));
  jnot g2741(.din(n2822), .dout(n2823));
  jxor g2742(.dina(n1059), .dinb(n699), .dout(n2824));
  jnot g2743(.din(n2824), .dout(n2825));
  jxor g2744(.dina(n808), .dinb(n708), .dout(n2826));
  jnot g2745(.din(n2826), .dout(n2827));
  jand g2746(.dina(n2827), .dinb(n2825), .dout(n2828));
  jand g2747(.dina(n2828), .dinb(n2823), .dout(n2829));
  jxor g2748(.dina(n1059), .dinb(n708), .dout(n2830));
  jnot g2749(.din(n2830), .dout(n2831));
  jand g2750(.dina(n2831), .dinb(n2824), .dout(n2832));
  jand g2751(.dina(n2832), .dinb(n2698), .dout(n2833));
  jand g2752(.dina(n2826), .dinb(n2825), .dout(n2834));
  jand g2753(.dina(n2834), .dinb(n2700), .dout(n2835));
  jor  g2754(.dina(n2835), .dinb(n2833), .dout(n2836));
  jor  g2755(.dina(n2836), .dinb(n2829), .dout(n2837));
  jnot g2756(.din(n2837), .dout(n2838));
  jand g2757(.dina(n2825), .dinb(n2698), .dout(n2839));
  jnot g2758(.din(n2839), .dout(n2840));
  jand g2759(.dina(n2840), .dinb(n803), .dout(n2841));
  jand g2760(.dina(n2841), .dinb(n2838), .dout(n2842));
  jxor g2761(.dina(n2821), .dinb(n2693), .dout(n2843));
  jnot g2762(.din(n2843), .dout(n2844));
  jand g2763(.dina(n2844), .dinb(n2828), .dout(n2845));
  jand g2764(.dina(n2834), .dinb(n2693), .dout(n2846));
  jand g2765(.dina(n2830), .dinb(n2824), .dout(n2847));
  jand g2766(.dina(n2847), .dinb(n2827), .dout(n2848));
  jand g2767(.dina(n2848), .dinb(n2698), .dout(n2849));
  jand g2768(.dina(n2832), .dinb(n2700), .dout(n2850));
  jor  g2769(.dina(n2850), .dinb(n2849), .dout(n2851));
  jor  g2770(.dina(n2851), .dinb(n2846), .dout(n2852));
  jor  g2771(.dina(n2852), .dinb(n2845), .dout(n2853));
  jnot g2772(.din(n2853), .dout(n2854));
  jand g2773(.dina(n2854), .dinb(n2842), .dout(n2855));
  jand g2774(.dina(n2855), .dinb(n2818), .dout(n2856));
  jnot g2775(.din(n2828), .dout(n2857));
  jxor g2776(.dina(n2701), .dinb(n2696), .dout(n2858));
  jor  g2777(.dina(n2858), .dinb(n2857), .dout(n2859));
  jnot g2778(.din(n2834), .dout(n2860));
  jor  g2779(.dina(n2860), .dinb(n2691), .dout(n2861));
  jnot g2780(.din(n2700), .dout(n2862));
  jnot g2781(.din(n2848), .dout(n2863));
  jor  g2782(.dina(n2863), .dinb(n2862), .dout(n2864));
  jnot g2783(.din(n2832), .dout(n2865));
  jor  g2784(.dina(n2865), .dinb(n2694), .dout(n2866));
  jand g2785(.dina(n2866), .dinb(n2864), .dout(n2867));
  jand g2786(.dina(n2867), .dinb(n2861), .dout(n2868));
  jand g2787(.dina(n2868), .dinb(n2859), .dout(n2869));
  jxor g2788(.dina(n2869), .dinb(n808), .dout(n2870));
  jxor g2789(.dina(n2855), .dinb(n2818), .dout(n2871));
  jand g2790(.dina(n2871), .dinb(n2870), .dout(n2872));
  jor  g2791(.dina(n2872), .dinb(n2856), .dout(n2873));
  jxor g2792(.dina(n2705), .dinb(n2704), .dout(n2874));
  jor  g2793(.dina(n2874), .dinb(n2857), .dout(n2875));
  jor  g2794(.dina(n2860), .dinb(n2688), .dout(n2876));
  jor  g2795(.dina(n2865), .dinb(n2691), .dout(n2877));
  jor  g2796(.dina(n2863), .dinb(n2694), .dout(n2878));
  jand g2797(.dina(n2878), .dinb(n2877), .dout(n2879));
  jand g2798(.dina(n2879), .dinb(n2876), .dout(n2880));
  jand g2799(.dina(n2880), .dinb(n2875), .dout(n2881));
  jxor g2800(.dina(n2881), .dinb(n808), .dout(n2882));
  jand g2801(.dina(n2817), .dinb(n2752), .dout(n2883));
  jand g2802(.dina(n2883), .dinb(n2823), .dout(n2884));
  jxor g2803(.dina(n980), .dinb(n961), .dout(n2885));
  jnot g2804(.din(n2885), .dout(n2886));
  jand g2805(.dina(n2886), .dinb(n2816), .dout(n2887));
  jand g2806(.dina(n2887), .dinb(n2698), .dout(n2888));
  jand g2807(.dina(n2817), .dinb(n2751), .dout(n2889));
  jand g2808(.dina(n2889), .dinb(n2700), .dout(n2890));
  jor  g2809(.dina(n2890), .dinb(n2888), .dout(n2891));
  jor  g2810(.dina(n2891), .dinb(n2884), .dout(n2892));
  jand g2811(.dina(n2698), .dinb(n954), .dout(n2893));
  jand g2812(.dina(n2893), .dinb(n2817), .dout(n2894));
  jxor g2813(.dina(n2894), .dinb(n2892), .dout(n2895));
  jxor g2814(.dina(n2895), .dinb(n2882), .dout(n2896));
  jxor g2815(.dina(n2896), .dinb(n2873), .dout(n2897));
  jand g2816(.dina(n2897), .dinb(n2815), .dout(n2898));
  jxor g2817(.dina(n2713), .dinb(n2711), .dout(n2899));
  jor  g2818(.dina(n2899), .dinb(n2795), .dout(n2900));
  jor  g2819(.dina(n2800), .dinb(n2681), .dout(n2901));
  jor  g2820(.dina(n2805), .dinb(n2687), .dout(n2902));
  jor  g2821(.dina(n2809), .dinb(n2688), .dout(n2903));
  jand g2822(.dina(n2903), .dinb(n2902), .dout(n2904));
  jand g2823(.dina(n2904), .dinb(n2901), .dout(n2905));
  jand g2824(.dina(n2905), .dinb(n2900), .dout(n2906));
  jxor g2825(.dina(n2906), .dinb(n1143), .dout(n2907));
  jxor g2826(.dina(n2871), .dinb(n2870), .dout(n2908));
  jand g2827(.dina(n2908), .dinb(n2907), .dout(n2909));
  jxor g2828(.dina(n2688), .dinb(n2687), .dout(n2910));
  jxor g2829(.dina(n2910), .dinb(n2708), .dout(n2911));
  jor  g2830(.dina(n2911), .dinb(n2795), .dout(n2912));
  jor  g2831(.dina(n2800), .dinb(n2687), .dout(n2913));
  jor  g2832(.dina(n2805), .dinb(n2688), .dout(n2914));
  jor  g2833(.dina(n2809), .dinb(n2691), .dout(n2915));
  jand g2834(.dina(n2915), .dinb(n2914), .dout(n2916));
  jand g2835(.dina(n2916), .dinb(n2913), .dout(n2917));
  jand g2836(.dina(n2917), .dinb(n2912), .dout(n2918));
  jxor g2837(.dina(n2918), .dinb(n699), .dout(n2919));
  jnot g2838(.din(n2919), .dout(n2920));
  jor  g2839(.dina(n2842), .dinb(n808), .dout(n2921));
  jxor g2840(.dina(n2921), .dinb(n2854), .dout(n2922));
  jand g2841(.dina(n2922), .dinb(n2920), .dout(n2923));
  jor  g2842(.dina(n2874), .dinb(n2795), .dout(n2924));
  jor  g2843(.dina(n2800), .dinb(n2688), .dout(n2925));
  jor  g2844(.dina(n2805), .dinb(n2691), .dout(n2926));
  jor  g2845(.dina(n2809), .dinb(n2694), .dout(n2927));
  jand g2846(.dina(n2927), .dinb(n2926), .dout(n2928));
  jand g2847(.dina(n2928), .dinb(n2925), .dout(n2929));
  jand g2848(.dina(n2929), .dinb(n2924), .dout(n2930));
  jxor g2849(.dina(n2930), .dinb(n1143), .dout(n2931));
  jand g2850(.dina(n2839), .dinb(n803), .dout(n2932));
  jxor g2851(.dina(n2932), .dinb(n2837), .dout(n2933));
  jand g2852(.dina(n2933), .dinb(n2931), .dout(n2934));
  jand g2853(.dina(n2823), .dinb(n2794), .dout(n2935));
  jand g2854(.dina(n2804), .dinb(n2698), .dout(n2936));
  jand g2855(.dina(n2799), .dinb(n2700), .dout(n2937));
  jor  g2856(.dina(n2937), .dinb(n2936), .dout(n2938));
  jor  g2857(.dina(n2938), .dinb(n2935), .dout(n2939));
  jnot g2858(.din(n2939), .dout(n2940));
  jand g2859(.dina(n2791), .dinb(n2698), .dout(n2941));
  jnot g2860(.din(n2941), .dout(n2942));
  jand g2861(.dina(n2942), .dinb(n699), .dout(n2943));
  jand g2862(.dina(n2943), .dinb(n2940), .dout(n2944));
  jand g2863(.dina(n2844), .dinb(n2794), .dout(n2945));
  jand g2864(.dina(n2799), .dinb(n2693), .dout(n2946));
  jand g2865(.dina(n2808), .dinb(n2698), .dout(n2947));
  jand g2866(.dina(n2804), .dinb(n2700), .dout(n2948));
  jor  g2867(.dina(n2948), .dinb(n2947), .dout(n2949));
  jor  g2868(.dina(n2949), .dinb(n2946), .dout(n2950));
  jor  g2869(.dina(n2950), .dinb(n2945), .dout(n2951));
  jnot g2870(.din(n2951), .dout(n2952));
  jand g2871(.dina(n2952), .dinb(n2944), .dout(n2953));
  jand g2872(.dina(n2953), .dinb(n2839), .dout(n2954));
  jor  g2873(.dina(n2858), .dinb(n2795), .dout(n2955));
  jor  g2874(.dina(n2800), .dinb(n2691), .dout(n2956));
  jor  g2875(.dina(n2809), .dinb(n2862), .dout(n2957));
  jor  g2876(.dina(n2805), .dinb(n2694), .dout(n2958));
  jand g2877(.dina(n2958), .dinb(n2957), .dout(n2959));
  jand g2878(.dina(n2959), .dinb(n2956), .dout(n2960));
  jand g2879(.dina(n2960), .dinb(n2955), .dout(n2961));
  jxor g2880(.dina(n2961), .dinb(n699), .dout(n2962));
  jnot g2881(.din(n2962), .dout(n2963));
  jxor g2882(.dina(n2953), .dinb(n2839), .dout(n2964));
  jand g2883(.dina(n2964), .dinb(n2963), .dout(n2965));
  jor  g2884(.dina(n2965), .dinb(n2954), .dout(n2966));
  jxor g2885(.dina(n2933), .dinb(n2931), .dout(n2967));
  jand g2886(.dina(n2967), .dinb(n2966), .dout(n2968));
  jor  g2887(.dina(n2968), .dinb(n2934), .dout(n2969));
  jxor g2888(.dina(n2922), .dinb(n2920), .dout(n2970));
  jand g2889(.dina(n2970), .dinb(n2969), .dout(n2971));
  jor  g2890(.dina(n2971), .dinb(n2923), .dout(n2972));
  jxor g2891(.dina(n2908), .dinb(n2907), .dout(n2973));
  jand g2892(.dina(n2973), .dinb(n2972), .dout(n2974));
  jor  g2893(.dina(n2974), .dinb(n2909), .dout(n2975));
  jxor g2894(.dina(n2897), .dinb(n2815), .dout(n2976));
  jand g2895(.dina(n2976), .dinb(n2975), .dout(n2977));
  jor  g2896(.dina(n2977), .dinb(n2898), .dout(n2978));
  jand g2897(.dina(n2895), .dinb(n2882), .dout(n2979));
  jand g2898(.dina(n2896), .dinb(n2873), .dout(n2980));
  jor  g2899(.dina(n2980), .dinb(n2979), .dout(n2981));
  jor  g2900(.dina(n2911), .dinb(n2857), .dout(n2982));
  jor  g2901(.dina(n2860), .dinb(n2687), .dout(n2983));
  jor  g2902(.dina(n2865), .dinb(n2688), .dout(n2984));
  jor  g2903(.dina(n2863), .dinb(n2691), .dout(n2985));
  jand g2904(.dina(n2985), .dinb(n2984), .dout(n2986));
  jand g2905(.dina(n2986), .dinb(n2983), .dout(n2987));
  jand g2906(.dina(n2987), .dinb(n2982), .dout(n2988));
  jxor g2907(.dina(n2988), .dinb(n808), .dout(n2989));
  jor  g2908(.dina(n2892), .dinb(n2818), .dout(n2990));
  jand g2909(.dina(n2990), .dinb(n954), .dout(n2991));
  jand g2910(.dina(n2883), .dinb(n2844), .dout(n2992));
  jand g2911(.dina(n2889), .dinb(n2693), .dout(n2993));
  jand g2912(.dina(n2885), .dinb(n2816), .dout(n2994));
  jand g2913(.dina(n2994), .dinb(n2752), .dout(n2995));
  jand g2914(.dina(n2995), .dinb(n2698), .dout(n2996));
  jand g2915(.dina(n2887), .dinb(n2700), .dout(n2997));
  jor  g2916(.dina(n2997), .dinb(n2996), .dout(n2998));
  jor  g2917(.dina(n2998), .dinb(n2993), .dout(n2999));
  jor  g2918(.dina(n2999), .dinb(n2992), .dout(n3000));
  jxor g2919(.dina(n3000), .dinb(n2991), .dout(n3001));
  jxor g2920(.dina(n3001), .dinb(n2989), .dout(n3002));
  jxor g2921(.dina(n3002), .dinb(n2981), .dout(n3003));
  jxor g2922(.dina(n2719), .dinb(n2718), .dout(n3004));
  jand g2923(.dina(n3004), .dinb(n2794), .dout(n3005));
  jand g2924(.dina(n2799), .dinb(n2677), .dout(n3006));
  jand g2925(.dina(n2808), .dinb(n2684), .dout(n3007));
  jand g2926(.dina(n2804), .dinb(n2679), .dout(n3008));
  jor  g2927(.dina(n3008), .dinb(n3007), .dout(n3009));
  jor  g2928(.dina(n3009), .dinb(n3006), .dout(n3010));
  jor  g2929(.dina(n3010), .dinb(n3005), .dout(n3011));
  jxor g2930(.dina(n3011), .dinb(n699), .dout(n3012));
  jxor g2931(.dina(n3012), .dinb(n3003), .dout(n3013));
  jxor g2932(.dina(n3013), .dinb(n2978), .dout(n3014));
  jand g2933(.dina(n3014), .dinb(n2789), .dout(n3015));
  jxor g2934(.dina(n2725), .dinb(n2724), .dout(n3016));
  jand g2935(.dina(n3016), .dinb(n78), .dout(n3017));
  jand g2936(.dina(n2774), .dinb(n2670), .dout(n3018));
  jand g2937(.dina(n2783), .dinb(n2677), .dout(n3019));
  jand g2938(.dina(n2779), .dinb(n2672), .dout(n3020));
  jor  g2939(.dina(n3020), .dinb(n3019), .dout(n3021));
  jor  g2940(.dina(n3021), .dinb(n3018), .dout(n3022));
  jor  g2941(.dina(n3022), .dinb(n3017), .dout(n3023));
  jxor g2942(.dina(n3023), .dinb(n55), .dout(n3024));
  jxor g2943(.dina(n2976), .dinb(n2975), .dout(n3025));
  jand g2944(.dina(n3025), .dinb(n3024), .dout(n3026));
  jnot g2945(.din(n2721), .dout(n3027));
  jxor g2946(.dina(n2722), .dinb(n3027), .dout(n3028));
  jor  g2947(.dina(n3028), .dinb(n79), .dout(n3029));
  jor  g2948(.dina(n2775), .dinb(n2671), .dout(n3030));
  jor  g2949(.dina(n2780), .dinb(n2674), .dout(n3031));
  jor  g2950(.dina(n2784), .dinb(n2678), .dout(n3032));
  jand g2951(.dina(n3032), .dinb(n3031), .dout(n3033));
  jand g2952(.dina(n3033), .dinb(n3030), .dout(n3034));
  jand g2953(.dina(n3034), .dinb(n3029), .dout(n3035));
  jxor g2954(.dina(n3035), .dinb(n56), .dout(n3036));
  jxor g2955(.dina(n2973), .dinb(n2972), .dout(n3037));
  jand g2956(.dina(n3037), .dinb(n3036), .dout(n3038));
  jand g2957(.dina(n3004), .dinb(n78), .dout(n3039));
  jand g2958(.dina(n2774), .dinb(n2677), .dout(n3040));
  jand g2959(.dina(n2783), .dinb(n2684), .dout(n3041));
  jand g2960(.dina(n2779), .dinb(n2679), .dout(n3042));
  jor  g2961(.dina(n3042), .dinb(n3041), .dout(n3043));
  jor  g2962(.dina(n3043), .dinb(n3040), .dout(n3044));
  jor  g2963(.dina(n3044), .dinb(n3039), .dout(n3045));
  jxor g2964(.dina(n3045), .dinb(n55), .dout(n3046));
  jxor g2965(.dina(n2970), .dinb(n2969), .dout(n3047));
  jand g2966(.dina(n3047), .dinb(n3046), .dout(n3048));
  jor  g2967(.dina(n2797), .dinb(n79), .dout(n3049));
  jor  g2968(.dina(n2775), .dinb(n2678), .dout(n3050));
  jor  g2969(.dina(n2780), .dinb(n2681), .dout(n3051));
  jor  g2970(.dina(n2784), .dinb(n2687), .dout(n3052));
  jand g2971(.dina(n3052), .dinb(n3051), .dout(n3053));
  jand g2972(.dina(n3053), .dinb(n3050), .dout(n3054));
  jand g2973(.dina(n3054), .dinb(n3049), .dout(n3055));
  jxor g2974(.dina(n3055), .dinb(n56), .dout(n3056));
  jxor g2975(.dina(n2967), .dinb(n2966), .dout(n3057));
  jand g2976(.dina(n3057), .dinb(n3056), .dout(n3058));
  jor  g2977(.dina(n2899), .dinb(n79), .dout(n3059));
  jor  g2978(.dina(n2775), .dinb(n2681), .dout(n3060));
  jor  g2979(.dina(n2780), .dinb(n2687), .dout(n3061));
  jor  g2980(.dina(n2784), .dinb(n2688), .dout(n3062));
  jand g2981(.dina(n3062), .dinb(n3061), .dout(n3063));
  jand g2982(.dina(n3063), .dinb(n3060), .dout(n3064));
  jand g2983(.dina(n3064), .dinb(n3059), .dout(n3065));
  jxor g2984(.dina(n3065), .dinb(n56), .dout(n3066));
  jxor g2985(.dina(n2964), .dinb(n2963), .dout(n3067));
  jand g2986(.dina(n3067), .dinb(n3066), .dout(n3068));
  jor  g2987(.dina(n2911), .dinb(n79), .dout(n3069));
  jor  g2988(.dina(n2775), .dinb(n2687), .dout(n3070));
  jor  g2989(.dina(n2780), .dinb(n2688), .dout(n3071));
  jor  g2990(.dina(n2784), .dinb(n2691), .dout(n3072));
  jand g2991(.dina(n3072), .dinb(n3071), .dout(n3073));
  jand g2992(.dina(n3073), .dinb(n3070), .dout(n3074));
  jand g2993(.dina(n3074), .dinb(n3069), .dout(n3075));
  jxor g2994(.dina(n3075), .dinb(n56), .dout(n3076));
  jor  g2995(.dina(n2944), .dinb(n1143), .dout(n3077));
  jxor g2996(.dina(n3077), .dinb(n2952), .dout(n3078));
  jand g2997(.dina(n3078), .dinb(n3076), .dout(n3079));
  jor  g2998(.dina(n2874), .dinb(n79), .dout(n3080));
  jor  g2999(.dina(n2775), .dinb(n2688), .dout(n3081));
  jor  g3000(.dina(n2780), .dinb(n2691), .dout(n3082));
  jor  g3001(.dina(n2784), .dinb(n2694), .dout(n3083));
  jand g3002(.dina(n3083), .dinb(n3082), .dout(n3084));
  jand g3003(.dina(n3084), .dinb(n3081), .dout(n3085));
  jand g3004(.dina(n3085), .dinb(n3080), .dout(n3086));
  jxor g3005(.dina(n3086), .dinb(n56), .dout(n3087));
  jand g3006(.dina(n2941), .dinb(n699), .dout(n3088));
  jxor g3007(.dina(n3088), .dinb(n2939), .dout(n3089));
  jand g3008(.dina(n3089), .dinb(n3087), .dout(n3090));
  jand g3009(.dina(n2823), .dinb(n78), .dout(n3091));
  jand g3010(.dina(n2779), .dinb(n2698), .dout(n3092));
  jand g3011(.dina(n2774), .dinb(n2700), .dout(n3093));
  jor  g3012(.dina(n3093), .dinb(n3092), .dout(n3094));
  jor  g3013(.dina(n3094), .dinb(n3091), .dout(n3095));
  jnot g3014(.din(n3095), .dout(n3096));
  jand g3015(.dina(n2698), .dinb(n70), .dout(n3097));
  jnot g3016(.din(n3097), .dout(n3098));
  jand g3017(.dina(n3098), .dinb(n55), .dout(n3099));
  jand g3018(.dina(n3099), .dinb(n3096), .dout(n3100));
  jand g3019(.dina(n2844), .dinb(n78), .dout(n3101));
  jand g3020(.dina(n2774), .dinb(n2693), .dout(n3102));
  jand g3021(.dina(n2783), .dinb(n2698), .dout(n3103));
  jand g3022(.dina(n2779), .dinb(n2700), .dout(n3104));
  jor  g3023(.dina(n3104), .dinb(n3103), .dout(n3105));
  jor  g3024(.dina(n3105), .dinb(n3102), .dout(n3106));
  jor  g3025(.dina(n3106), .dinb(n3101), .dout(n3107));
  jnot g3026(.din(n3107), .dout(n3108));
  jand g3027(.dina(n3108), .dinb(n3100), .dout(n3109));
  jand g3028(.dina(n3109), .dinb(n2941), .dout(n3110));
  jor  g3029(.dina(n2858), .dinb(n79), .dout(n3111));
  jor  g3030(.dina(n2775), .dinb(n2691), .dout(n3112));
  jor  g3031(.dina(n2784), .dinb(n2862), .dout(n3113));
  jor  g3032(.dina(n2780), .dinb(n2694), .dout(n3114));
  jand g3033(.dina(n3114), .dinb(n3113), .dout(n3115));
  jand g3034(.dina(n3115), .dinb(n3112), .dout(n3116));
  jand g3035(.dina(n3116), .dinb(n3111), .dout(n3117));
  jxor g3036(.dina(n3117), .dinb(n56), .dout(n3118));
  jxor g3037(.dina(n3109), .dinb(n2941), .dout(n3119));
  jand g3038(.dina(n3119), .dinb(n3118), .dout(n3120));
  jor  g3039(.dina(n3120), .dinb(n3110), .dout(n3121));
  jxor g3040(.dina(n3089), .dinb(n3087), .dout(n3122));
  jand g3041(.dina(n3122), .dinb(n3121), .dout(n3123));
  jor  g3042(.dina(n3123), .dinb(n3090), .dout(n3124));
  jxor g3043(.dina(n3078), .dinb(n3076), .dout(n3125));
  jand g3044(.dina(n3125), .dinb(n3124), .dout(n3126));
  jor  g3045(.dina(n3126), .dinb(n3079), .dout(n3127));
  jxor g3046(.dina(n3067), .dinb(n3066), .dout(n3128));
  jand g3047(.dina(n3128), .dinb(n3127), .dout(n3129));
  jor  g3048(.dina(n3129), .dinb(n3068), .dout(n3130));
  jxor g3049(.dina(n3057), .dinb(n3056), .dout(n3131));
  jand g3050(.dina(n3131), .dinb(n3130), .dout(n3132));
  jor  g3051(.dina(n3132), .dinb(n3058), .dout(n3133));
  jxor g3052(.dina(n3047), .dinb(n3046), .dout(n3134));
  jand g3053(.dina(n3134), .dinb(n3133), .dout(n3135));
  jor  g3054(.dina(n3135), .dinb(n3048), .dout(n3136));
  jxor g3055(.dina(n3037), .dinb(n3036), .dout(n3137));
  jand g3056(.dina(n3137), .dinb(n3136), .dout(n3138));
  jor  g3057(.dina(n3138), .dinb(n3038), .dout(n3139));
  jxor g3058(.dina(n3025), .dinb(n3024), .dout(n3140));
  jand g3059(.dina(n3140), .dinb(n3139), .dout(n3141));
  jor  g3060(.dina(n3141), .dinb(n3026), .dout(n3142));
  jxor g3061(.dina(n3014), .dinb(n2789), .dout(n3143));
  jand g3062(.dina(n3143), .dinb(n3142), .dout(n3144));
  jor  g3063(.dina(n3144), .dinb(n3015), .dout(n3145));
  jand g3064(.dina(n2769), .dinb(n2670), .dout(n3146));
  jand g3065(.dina(n2770), .dinb(n2727), .dout(n3147));
  jor  g3066(.dina(n3147), .dinb(n3146), .dout(n3148));
  jor  g3067(.dina(n2767), .dinb(n2750), .dout(n3149));
  jnot g3068(.din(n3149), .dout(n3150));
  jand g3069(.dina(n2767), .dinb(n2750), .dout(n3151));
  jnot g3070(.din(n3151), .dout(n3152));
  jand g3071(.dina(n3152), .dinb(n2733), .dout(n3153));
  jor  g3072(.dina(n3153), .dinb(n3150), .dout(n3154));
  jnot g3073(.din(n1653), .dout(n3155));
  jand g3074(.dina(n461), .dinb(n312), .dout(n3156));
  jand g3075(.dina(n3156), .dinb(n304), .dout(n3157));
  jand g3076(.dina(n3157), .dinb(n898), .dout(n3158));
  jand g3077(.dina(n3158), .dinb(n914), .dout(n3159));
  jand g3078(.dina(n711), .dinb(n564), .dout(n3160));
  jand g3079(.dina(n3160), .dinb(n821), .dout(n3161));
  jand g3080(.dina(n612), .dinb(n499), .dout(n3162));
  jand g3081(.dina(n853), .dinb(n225), .dout(n3163));
  jand g3082(.dina(n3163), .dinb(n3162), .dout(n3164));
  jand g3083(.dina(n3164), .dinb(n1189), .dout(n3165));
  jand g3084(.dina(n3165), .dinb(n3161), .dout(n3166));
  jand g3085(.dina(n3166), .dinb(n3159), .dout(n3167));
  jand g3086(.dina(n2427), .dinb(n1011), .dout(n3168));
  jand g3087(.dina(n3168), .dinb(n3167), .dout(n3169));
  jand g3088(.dina(n3169), .dinb(n3155), .dout(n3170));
  jnot g3089(.din(n3170), .dout(n3171));
  jxor g3090(.dina(n3171), .dinb(n3154), .dout(n3172));
  jxor g3091(.dina(n3172), .dinb(n2773), .dout(n3173));
  jxor g3092(.dina(n3173), .dinb(n3148), .dout(n3174));
  jand g3093(.dina(n3174), .dinb(n78), .dout(n3175));
  jnot g3094(.din(n3172), .dout(n3176));
  jand g3095(.dina(n3176), .dinb(n2774), .dout(n3177));
  jand g3096(.dina(n2783), .dinb(n2670), .dout(n3178));
  jand g3097(.dina(n2779), .dinb(n2769), .dout(n3179));
  jor  g3098(.dina(n3179), .dinb(n3178), .dout(n3180));
  jor  g3099(.dina(n3180), .dinb(n3177), .dout(n3181));
  jor  g3100(.dina(n3181), .dinb(n3175), .dout(n3182));
  jxor g3101(.dina(n3182), .dinb(n55), .dout(n3183));
  jand g3102(.dina(n3012), .dinb(n3003), .dout(n3184));
  jand g3103(.dina(n3013), .dinb(n2978), .dout(n3185));
  jor  g3104(.dina(n3185), .dinb(n3184), .dout(n3186));
  jand g3105(.dina(n3001), .dinb(n2989), .dout(n3187));
  jand g3106(.dina(n3002), .dinb(n2981), .dout(n3188));
  jor  g3107(.dina(n3188), .dinb(n3187), .dout(n3189));
  jor  g3108(.dina(n2899), .dinb(n2857), .dout(n3190));
  jor  g3109(.dina(n2860), .dinb(n2681), .dout(n3191));
  jor  g3110(.dina(n2865), .dinb(n2687), .dout(n3192));
  jor  g3111(.dina(n2863), .dinb(n2688), .dout(n3193));
  jand g3112(.dina(n3193), .dinb(n3192), .dout(n3194));
  jand g3113(.dina(n3194), .dinb(n3191), .dout(n3195));
  jand g3114(.dina(n3195), .dinb(n3190), .dout(n3196));
  jxor g3115(.dina(n3196), .dinb(n808), .dout(n3197));
  jnot g3116(.din(n2883), .dout(n3198));
  jor  g3117(.dina(n3198), .dinb(n2858), .dout(n3199));
  jnot g3118(.din(n2889), .dout(n3200));
  jor  g3119(.dina(n3200), .dinb(n2691), .dout(n3201));
  jnot g3120(.din(n2995), .dout(n3202));
  jor  g3121(.dina(n3202), .dinb(n2862), .dout(n3203));
  jnot g3122(.din(n2887), .dout(n3204));
  jor  g3123(.dina(n3204), .dinb(n2694), .dout(n3205));
  jand g3124(.dina(n3205), .dinb(n3203), .dout(n3206));
  jand g3125(.dina(n3206), .dinb(n3201), .dout(n3207));
  jand g3126(.dina(n3207), .dinb(n3199), .dout(n3208));
  jxor g3127(.dina(n3208), .dinb(n954), .dout(n3209));
  jnot g3128(.din(n3209), .dout(n3210));
  jor  g3129(.dina(n3000), .dinb(n2990), .dout(n3211));
  jnot g3130(.din(n3211), .dout(n3212));
  jand g3131(.dina(n3212), .dinb(n954), .dout(n3213));
  jor  g3132(.dina(n3213), .dinb(n2893), .dout(n3214));
  jand g3133(.dina(n3212), .dinb(n2893), .dout(n3215));
  jnot g3134(.din(n3215), .dout(n3216));
  jand g3135(.dina(n3216), .dinb(n3214), .dout(n3217));
  jxor g3136(.dina(n3217), .dinb(n3210), .dout(n3218));
  jxor g3137(.dina(n3218), .dinb(n3197), .dout(n3219));
  jxor g3138(.dina(n3219), .dinb(n3189), .dout(n3220));
  jor  g3139(.dina(n3028), .dinb(n2795), .dout(n3221));
  jor  g3140(.dina(n2800), .dinb(n2671), .dout(n3222));
  jor  g3141(.dina(n2805), .dinb(n2674), .dout(n3223));
  jor  g3142(.dina(n2809), .dinb(n2678), .dout(n3224));
  jand g3143(.dina(n3224), .dinb(n3223), .dout(n3225));
  jand g3144(.dina(n3225), .dinb(n3222), .dout(n3226));
  jand g3145(.dina(n3226), .dinb(n3221), .dout(n3227));
  jxor g3146(.dina(n3227), .dinb(n1143), .dout(n3228));
  jxor g3147(.dina(n3228), .dinb(n3220), .dout(n3229));
  jxor g3148(.dina(n3229), .dinb(n3186), .dout(n3230));
  jxor g3149(.dina(n3230), .dinb(n3183), .dout(n3231));
  jxor g3150(.dina(n3231), .dinb(n3145), .dout(n3232));
  jnot g3151(.din(n68), .dout(n3233));
  jand g3152(.dina(n49), .dinb(a0 ), .dout(n3234));
  jxor g3153(.dina(n3234), .dinb(n62), .dout(n3235));
  jxor g3154(.dina(n3235), .dinb(n3233), .dout(n3236));
  jand g3155(.dina(n3236), .dinb(a0 ), .dout(n3237));
  jnot g3156(.din(n3237), .dout(n3238));
  jor  g3157(.dina(n3171), .dinb(n3154), .dout(n3239));
  jnot g3158(.din(n3239), .dout(n3240));
  jand g3159(.dina(n2380), .dinb(n437), .dout(n3241));
  jand g3160(.dina(n3241), .dinb(n936), .dout(n3242));
  jand g3161(.dina(n772), .dinb(n477), .dout(n3243));
  jand g3162(.dina(n624), .dinb(n261), .dout(n3244));
  jand g3163(.dina(n3244), .dinb(n3243), .dout(n3245));
  jand g3164(.dina(n3245), .dinb(n3242), .dout(n3246));
  jand g3165(.dina(n3246), .dinb(n2321), .dout(n3247));
  jand g3166(.dina(n882), .dinb(n323), .dout(n3248));
  jand g3167(.dina(n3248), .dinb(n381), .dout(n3249));
  jand g3168(.dina(n3249), .dinb(n2580), .dout(n3250));
  jand g3169(.dina(n724), .dinb(n918), .dout(n3251));
  jand g3170(.dina(n594), .dinb(n370), .dout(n3252));
  jand g3171(.dina(n3252), .dinb(n3251), .dout(n3253));
  jand g3172(.dina(n3253), .dinb(n2655), .dout(n3254));
  jand g3173(.dina(n3254), .dinb(n3250), .dout(n3255));
  jand g3174(.dina(n3255), .dinb(n3247), .dout(n3256));
  jand g3175(.dina(n363), .dinb(n291), .dout(n3257));
  jand g3176(.dina(n3257), .dinb(n277), .dout(n3258));
  jand g3177(.dina(n710), .dinb(n232), .dout(n3259));
  jand g3178(.dina(n3259), .dinb(n2538), .dout(n3260));
  jand g3179(.dina(n3260), .dinb(n3258), .dout(n3261));
  jand g3180(.dina(n3261), .dinb(n2453), .dout(n3262));
  jand g3181(.dina(n868), .dinb(n153), .dout(n3263));
  jand g3182(.dina(n506), .dinb(n312), .dout(n3264));
  jand g3183(.dina(n3264), .dinb(n3263), .dout(n3265));
  jand g3184(.dina(n3265), .dinb(n822), .dout(n3266));
  jand g3185(.dina(n3266), .dinb(n361), .dout(n3267));
  jand g3186(.dina(n3267), .dinb(n3262), .dout(n3268));
  jand g3187(.dina(n3268), .dinb(n3256), .dout(n3269));
  jand g3188(.dina(n3269), .dinb(n434), .dout(n3270));
  jand g3189(.dina(n3270), .dinb(n3240), .dout(n3271));
  jand g3190(.dina(n426), .dinb(n374), .dout(n3272));
  jand g3191(.dina(n3272), .dinb(n2289), .dout(n3273));
  jnot g3192(.din(n650), .dout(n3274));
  jand g3193(.dina(n1310), .dinb(n3274), .dout(n3275));
  jand g3194(.dina(n2511), .dinb(n930), .dout(n3276));
  jand g3195(.dina(n3276), .dinb(n3275), .dout(n3277));
  jand g3196(.dina(n3277), .dinb(n3273), .dout(n3278));
  jand g3197(.dina(n2417), .dinb(n2307), .dout(n3279));
  jand g3198(.dina(n3279), .dinb(n3278), .dout(n3280));
  jand g3199(.dina(n3280), .dinb(n719), .dout(n3281));
  jand g3200(.dina(n3281), .dinb(n275), .dout(n3282));
  jxor g3201(.dina(n3282), .dinb(n3271), .dout(n3283));
  jxor g3202(.dina(n3270), .dinb(n3240), .dout(n3284));
  jor  g3203(.dina(n3284), .dinb(n3283), .dout(n3285));
  jnot g3204(.din(n3285), .dout(n3286));
  jor  g3205(.dina(n3284), .dinb(n3172), .dout(n3287));
  jnot g3206(.din(n3287), .dout(n3288));
  jand g3207(.dina(n3176), .dinb(n2769), .dout(n3289));
  jand g3208(.dina(n3173), .dinb(n3148), .dout(n3290));
  jor  g3209(.dina(n3290), .dinb(n3289), .dout(n3291));
  jand g3210(.dina(n3270), .dinb(n3172), .dout(n3292));
  jnot g3211(.din(n3292), .dout(n3293));
  jand g3212(.dina(n3293), .dinb(n3287), .dout(n3294));
  jand g3213(.dina(n3294), .dinb(n3291), .dout(n3295));
  jor  g3214(.dina(n3295), .dinb(n3288), .dout(n3296));
  jand g3215(.dina(n3284), .dinb(n3282), .dout(n3297));
  jnot g3216(.din(n3297), .dout(n3298));
  jand g3217(.dina(n3298), .dinb(n3285), .dout(n3299));
  jand g3218(.dina(n3299), .dinb(n3296), .dout(n3300));
  jor  g3219(.dina(n3300), .dinb(n3286), .dout(n3301));
  jnot g3220(.din(n3283), .dout(n3302));
  jand g3221(.dina(n3282), .dinb(n3271), .dout(n3303));
  jnot g3222(.din(n1322), .dout(n3304));
  jand g3223(.dina(n3304), .dinb(n319), .dout(n3305));
  jand g3224(.dina(n3305), .dinb(n287), .dout(n3306));
  jand g3225(.dina(n254), .dinb(n241), .dout(n3307));
  jand g3226(.dina(n3307), .dinb(n1209), .dout(n3308));
  jand g3227(.dina(n3308), .dinb(n731), .dout(n3309));
  jand g3228(.dina(n3309), .dinb(n746), .dout(n3310));
  jand g3229(.dina(n3310), .dinb(n3306), .dout(n3311));
  jand g3230(.dina(n786), .dinb(n719), .dout(n3312));
  jand g3231(.dina(n3312), .dinb(n218), .dout(n3313));
  jand g3232(.dina(n3313), .dinb(n3311), .dout(n3314));
  jxor g3233(.dina(n3314), .dinb(n3303), .dout(n3315));
  jnot g3234(.din(n3315), .dout(n3316));
  jand g3235(.dina(n3316), .dinb(n3302), .dout(n3317));
  jand g3236(.dina(n3314), .dinb(n3283), .dout(n3318));
  jor  g3237(.dina(n3318), .dinb(n3317), .dout(n3319));
  jxor g3238(.dina(n3319), .dinb(n3301), .dout(n3320));
  jor  g3239(.dina(n3320), .dinb(n3238), .dout(n3321));
  jor  g3240(.dina(n3236), .dinb(n61), .dout(n3322));
  jor  g3241(.dina(n3322), .dinb(n3315), .dout(n3323));
  jand g3242(.dina(a1 ), .dinb(n61), .dout(n3324));
  jnot g3243(.din(n3324), .dout(n3325));
  jor  g3244(.dina(n3325), .dinb(n3283), .dout(n3326));
  jand g3245(.dina(n63), .dinb(a2 ), .dout(n3327));
  jnot g3246(.din(n3327), .dout(n3328));
  jor  g3247(.dina(n3328), .dinb(n3284), .dout(n3329));
  jand g3248(.dina(n3329), .dinb(n3326), .dout(n3330));
  jand g3249(.dina(n3330), .dinb(n3323), .dout(n3331));
  jand g3250(.dina(n3331), .dinb(n3321), .dout(n3332));
  jxor g3251(.dina(n3332), .dinb(n3233), .dout(n3333));
  jand g3252(.dina(n3333), .dinb(n3232), .dout(n3334));
  jxor g3253(.dina(n3143), .dinb(n3142), .dout(n3335));
  jnot g3254(.din(n3299), .dout(n3336));
  jxor g3255(.dina(n3336), .dinb(n3296), .dout(n3337));
  jor  g3256(.dina(n3337), .dinb(n3238), .dout(n3338));
  jor  g3257(.dina(n3322), .dinb(n3283), .dout(n3339));
  jor  g3258(.dina(n3325), .dinb(n3284), .dout(n3340));
  jor  g3259(.dina(n3328), .dinb(n3172), .dout(n3341));
  jand g3260(.dina(n3341), .dinb(n3340), .dout(n3342));
  jand g3261(.dina(n3342), .dinb(n3339), .dout(n3343));
  jand g3262(.dina(n3343), .dinb(n3338), .dout(n3344));
  jxor g3263(.dina(n3344), .dinb(n3233), .dout(n3345));
  jand g3264(.dina(n3345), .dinb(n3335), .dout(n3346));
  jxor g3265(.dina(n3345), .dinb(n3335), .dout(n3347));
  jxor g3266(.dina(n3140), .dinb(n3139), .dout(n3348));
  jxor g3267(.dina(n3137), .dinb(n3136), .dout(n3349));
  jxor g3268(.dina(n3134), .dinb(n3133), .dout(n3350));
  jxor g3269(.dina(n3131), .dinb(n3130), .dout(n3351));
  jxor g3270(.dina(n3128), .dinb(n3127), .dout(n3352));
  jxor g3271(.dina(n3125), .dinb(n3124), .dout(n3353));
  jxor g3272(.dina(n3122), .dinb(n3121), .dout(n3354));
  jor  g3273(.dina(n3238), .dinb(n2899), .dout(n3355));
  jor  g3274(.dina(n3322), .dinb(n2681), .dout(n3356));
  jor  g3275(.dina(n3325), .dinb(n2687), .dout(n3357));
  jor  g3276(.dina(n3328), .dinb(n2688), .dout(n3358));
  jand g3277(.dina(n3358), .dinb(n3357), .dout(n3359));
  jand g3278(.dina(n3359), .dinb(n3356), .dout(n3360));
  jand g3279(.dina(n3360), .dinb(n3355), .dout(n3361));
  jxor g3280(.dina(n3361), .dinb(n3233), .dout(n3362));
  jnot g3281(.din(n3100), .dout(n3363));
  jand g3282(.dina(n3363), .dinb(n55), .dout(n3364));
  jxor g3283(.dina(n3364), .dinb(n3107), .dout(n3365));
  jand g3284(.dina(n3097), .dinb(n55), .dout(n3366));
  jxor g3285(.dina(n3366), .dinb(n3095), .dout(n3367));
  jxor g3286(.dina(n2702), .dinb(n2696), .dout(n3368));
  jand g3287(.dina(n3237), .dinb(n3368), .dout(n3369));
  jor  g3288(.dina(n3322), .dinb(n2691), .dout(n3370));
  jand g3289(.dina(n3324), .dinb(n2693), .dout(n3371));
  jnot g3290(.din(n3371), .dout(n3372));
  jand g3291(.dina(n3372), .dinb(n3370), .dout(n3373));
  jnot g3292(.din(n3373), .dout(n3374));
  jor  g3293(.dina(n3374), .dinb(n3369), .dout(n3375));
  jand g3294(.dina(n2700), .dinb(n63), .dout(n3376));
  jor  g3295(.dina(n3376), .dinb(n3233), .dout(n3377));
  jnot g3296(.din(n3377), .dout(n3378));
  jor  g3297(.dina(n3378), .dinb(n3375), .dout(n3379));
  jor  g3298(.dina(n3238), .dinb(n2858), .dout(n3380));
  jand g3299(.dina(n3373), .dinb(n3380), .dout(n3381));
  jor  g3300(.dina(n3381), .dinb(n3233), .dout(n3382));
  jand g3301(.dina(n3238), .dinb(n2862), .dout(n3383));
  jand g3302(.dina(n3238), .dinb(n64), .dout(n3384));
  jnot g3303(.din(n3384), .dout(n3385));
  jand g3304(.dina(n3385), .dinb(n2822), .dout(n3386));
  jor  g3305(.dina(n3386), .dinb(n3383), .dout(n3387));
  jand g3306(.dina(n3387), .dinb(n2694), .dout(n3388));
  jor  g3307(.dina(n3235), .dinb(n2862), .dout(n3389));
  jand g3308(.dina(n3389), .dinb(n61), .dout(n3390));
  jor  g3309(.dina(n3390), .dinb(n3388), .dout(n3391));
  jand g3310(.dina(n2697), .dinb(n68), .dout(n3392));
  jand g3311(.dina(n3392), .dinb(n3391), .dout(n3393));
  jor  g3312(.dina(n3393), .dinb(n3097), .dout(n3394));
  jand g3313(.dina(n3394), .dinb(n3382), .dout(n3395));
  jand g3314(.dina(n3395), .dinb(n3379), .dout(n3396));
  jand g3315(.dina(n3396), .dinb(n3367), .dout(n3397));
  jor  g3316(.dina(n3396), .dinb(n3367), .dout(n3398));
  jor  g3317(.dina(n3238), .dinb(n2874), .dout(n3399));
  jor  g3318(.dina(n3322), .dinb(n2688), .dout(n3400));
  jor  g3319(.dina(n3325), .dinb(n2691), .dout(n3401));
  jor  g3320(.dina(n3328), .dinb(n2694), .dout(n3402));
  jand g3321(.dina(n3402), .dinb(n3401), .dout(n3403));
  jand g3322(.dina(n3403), .dinb(n3400), .dout(n3404));
  jand g3323(.dina(n3404), .dinb(n3399), .dout(n3405));
  jxor g3324(.dina(n3405), .dinb(n3233), .dout(n3406));
  jand g3325(.dina(n3406), .dinb(n3398), .dout(n3407));
  jor  g3326(.dina(n3407), .dinb(n3397), .dout(n3408));
  jor  g3327(.dina(n3408), .dinb(n3365), .dout(n3409));
  jand g3328(.dina(n3408), .dinb(n3365), .dout(n3410));
  jor  g3329(.dina(n3238), .dinb(n2911), .dout(n3411));
  jor  g3330(.dina(n3322), .dinb(n2687), .dout(n3412));
  jor  g3331(.dina(n3325), .dinb(n2688), .dout(n3413));
  jor  g3332(.dina(n3328), .dinb(n2691), .dout(n3414));
  jand g3333(.dina(n3414), .dinb(n3413), .dout(n3415));
  jand g3334(.dina(n3415), .dinb(n3412), .dout(n3416));
  jand g3335(.dina(n3416), .dinb(n3411), .dout(n3417));
  jxor g3336(.dina(n3417), .dinb(n3233), .dout(n3418));
  jor  g3337(.dina(n3418), .dinb(n3410), .dout(n3419));
  jand g3338(.dina(n3419), .dinb(n3409), .dout(n3420));
  jand g3339(.dina(n3420), .dinb(n3362), .dout(n3421));
  jor  g3340(.dina(n3420), .dinb(n3362), .dout(n3422));
  jxor g3341(.dina(n3119), .dinb(n3118), .dout(n3423));
  jand g3342(.dina(n3423), .dinb(n3422), .dout(n3424));
  jor  g3343(.dina(n3424), .dinb(n3421), .dout(n3425));
  jor  g3344(.dina(n3425), .dinb(n3354), .dout(n3426));
  jand g3345(.dina(n3425), .dinb(n3354), .dout(n3427));
  jor  g3346(.dina(n3238), .dinb(n2797), .dout(n3428));
  jor  g3347(.dina(n3322), .dinb(n2678), .dout(n3429));
  jor  g3348(.dina(n3325), .dinb(n2681), .dout(n3430));
  jor  g3349(.dina(n3328), .dinb(n2687), .dout(n3431));
  jand g3350(.dina(n3431), .dinb(n3430), .dout(n3432));
  jand g3351(.dina(n3432), .dinb(n3429), .dout(n3433));
  jand g3352(.dina(n3433), .dinb(n3428), .dout(n3434));
  jxor g3353(.dina(n3434), .dinb(n3233), .dout(n3435));
  jor  g3354(.dina(n3435), .dinb(n3427), .dout(n3436));
  jand g3355(.dina(n3436), .dinb(n3426), .dout(n3437));
  jand g3356(.dina(n3437), .dinb(n3353), .dout(n3438));
  jor  g3357(.dina(n3437), .dinb(n3353), .dout(n3439));
  jand g3358(.dina(n3237), .dinb(n3004), .dout(n3440));
  jor  g3359(.dina(n3322), .dinb(n2674), .dout(n3441));
  jand g3360(.dina(n3324), .dinb(n2679), .dout(n3442));
  jnot g3361(.din(n3442), .dout(n3443));
  jand g3362(.dina(n3443), .dinb(n3441), .dout(n3444));
  jnot g3363(.din(n3444), .dout(n3445));
  jor  g3364(.dina(n3445), .dinb(n3440), .dout(n3446));
  jand g3365(.dina(n3446), .dinb(n3233), .dout(n3447));
  jand g3366(.dina(n2684), .dinb(n63), .dout(n3448));
  jor  g3367(.dina(n3448), .dinb(n3233), .dout(n3449));
  jor  g3368(.dina(n3449), .dinb(n3446), .dout(n3450));
  jnot g3369(.din(n3450), .dout(n3451));
  jor  g3370(.dina(n3451), .dinb(n3447), .dout(n3452));
  jand g3371(.dina(n3452), .dinb(n3439), .dout(n3453));
  jor  g3372(.dina(n3453), .dinb(n3438), .dout(n3454));
  jand g3373(.dina(n3454), .dinb(n3352), .dout(n3455));
  jor  g3374(.dina(n3454), .dinb(n3352), .dout(n3456));
  jor  g3375(.dina(n3238), .dinb(n3028), .dout(n3457));
  jor  g3376(.dina(n3322), .dinb(n2671), .dout(n3458));
  jor  g3377(.dina(n3325), .dinb(n2674), .dout(n3459));
  jor  g3378(.dina(n3328), .dinb(n2678), .dout(n3460));
  jand g3379(.dina(n3460), .dinb(n3459), .dout(n3461));
  jand g3380(.dina(n3461), .dinb(n3458), .dout(n3462));
  jand g3381(.dina(n3462), .dinb(n3457), .dout(n3463));
  jxor g3382(.dina(n3463), .dinb(n3233), .dout(n3464));
  jand g3383(.dina(n3464), .dinb(n3456), .dout(n3465));
  jor  g3384(.dina(n3465), .dinb(n3455), .dout(n3466));
  jand g3385(.dina(n3466), .dinb(n3351), .dout(n3467));
  jor  g3386(.dina(n3466), .dinb(n3351), .dout(n3468));
  jand g3387(.dina(n3237), .dinb(n3016), .dout(n3469));
  jnot g3388(.din(n3469), .dout(n3470));
  jor  g3389(.dina(n3322), .dinb(n2669), .dout(n3471));
  jand g3390(.dina(n3324), .dinb(n2672), .dout(n3472));
  jnot g3391(.din(n3472), .dout(n3473));
  jand g3392(.dina(n3473), .dinb(n3471), .dout(n3474));
  jand g3393(.dina(n3474), .dinb(n3470), .dout(n3475));
  jnot g3394(.din(n3475), .dout(n3476));
  jand g3395(.dina(n3476), .dinb(n3233), .dout(n3477));
  jand g3396(.dina(n2677), .dinb(n63), .dout(n3478));
  jor  g3397(.dina(n3478), .dinb(n3233), .dout(n3479));
  jnot g3398(.din(n3479), .dout(n3480));
  jand g3399(.dina(n3480), .dinb(n3475), .dout(n3481));
  jor  g3400(.dina(n3481), .dinb(n3477), .dout(n3482));
  jand g3401(.dina(n3482), .dinb(n3468), .dout(n3483));
  jor  g3402(.dina(n3483), .dinb(n3467), .dout(n3484));
  jor  g3403(.dina(n3484), .dinb(n3350), .dout(n3485));
  jand g3404(.dina(n3484), .dinb(n3350), .dout(n3486));
  jor  g3405(.dina(n3238), .dinb(n2771), .dout(n3487));
  jor  g3406(.dina(n3322), .dinb(n2773), .dout(n3488));
  jor  g3407(.dina(n3325), .dinb(n2669), .dout(n3489));
  jor  g3408(.dina(n3328), .dinb(n2671), .dout(n3490));
  jand g3409(.dina(n3490), .dinb(n3489), .dout(n3491));
  jand g3410(.dina(n3491), .dinb(n3488), .dout(n3492));
  jand g3411(.dina(n3492), .dinb(n3487), .dout(n3493));
  jxor g3412(.dina(n3493), .dinb(n3233), .dout(n3494));
  jor  g3413(.dina(n3494), .dinb(n3486), .dout(n3495));
  jand g3414(.dina(n3495), .dinb(n3485), .dout(n3496));
  jand g3415(.dina(n3496), .dinb(n3349), .dout(n3497));
  jor  g3416(.dina(n3496), .dinb(n3349), .dout(n3498));
  jand g3417(.dina(n3237), .dinb(n3174), .dout(n3499));
  jnot g3418(.din(n3322), .dout(n3500));
  jand g3419(.dina(n3500), .dinb(n3176), .dout(n3501));
  jand g3420(.dina(n3324), .dinb(n2769), .dout(n3502));
  jor  g3421(.dina(n3502), .dinb(n3501), .dout(n3503));
  jor  g3422(.dina(n3503), .dinb(n3499), .dout(n3504));
  jand g3423(.dina(n3504), .dinb(n3233), .dout(n3505));
  jand g3424(.dina(n2670), .dinb(n63), .dout(n3506));
  jor  g3425(.dina(n3506), .dinb(n3233), .dout(n3507));
  jor  g3426(.dina(n3507), .dinb(n3504), .dout(n3508));
  jnot g3427(.din(n3508), .dout(n3509));
  jor  g3428(.dina(n3509), .dinb(n3505), .dout(n3510));
  jand g3429(.dina(n3510), .dinb(n3498), .dout(n3511));
  jor  g3430(.dina(n3511), .dinb(n3497), .dout(n3512));
  jor  g3431(.dina(n3512), .dinb(n3348), .dout(n3513));
  jand g3432(.dina(n3512), .dinb(n3348), .dout(n3514));
  jnot g3433(.din(n3291), .dout(n3515));
  jxor g3434(.dina(n3294), .dinb(n3515), .dout(n3516));
  jor  g3435(.dina(n3516), .dinb(n3238), .dout(n3517));
  jor  g3436(.dina(n3322), .dinb(n3284), .dout(n3518));
  jor  g3437(.dina(n3325), .dinb(n3172), .dout(n3519));
  jor  g3438(.dina(n3328), .dinb(n2773), .dout(n3520));
  jand g3439(.dina(n3520), .dinb(n3519), .dout(n3521));
  jand g3440(.dina(n3521), .dinb(n3518), .dout(n3522));
  jand g3441(.dina(n3522), .dinb(n3517), .dout(n3523));
  jxor g3442(.dina(n3523), .dinb(n68), .dout(n3524));
  jnot g3443(.din(n3524), .dout(n3525));
  jor  g3444(.dina(n3525), .dinb(n3514), .dout(n3526));
  jand g3445(.dina(n3526), .dinb(n3513), .dout(n3527));
  jand g3446(.dina(n3527), .dinb(n3347), .dout(n3528));
  jor  g3447(.dina(n3528), .dinb(n3346), .dout(n3529));
  jxor g3448(.dina(n3333), .dinb(n3232), .dout(n3530));
  jand g3449(.dina(n3530), .dinb(n3529), .dout(n3531));
  jor  g3450(.dina(n3531), .dinb(n3334), .dout(n3532));
  jand g3451(.dina(n3230), .dinb(n3183), .dout(n3533));
  jand g3452(.dina(n3231), .dinb(n3145), .dout(n3534));
  jor  g3453(.dina(n3534), .dinb(n3533), .dout(n3535));
  jor  g3454(.dina(n3516), .dinb(n79), .dout(n3536));
  jor  g3455(.dina(n3284), .dinb(n2775), .dout(n3537));
  jor  g3456(.dina(n3172), .dinb(n2780), .dout(n3538));
  jor  g3457(.dina(n2784), .dinb(n2773), .dout(n3539));
  jand g3458(.dina(n3539), .dinb(n3538), .dout(n3540));
  jand g3459(.dina(n3540), .dinb(n3537), .dout(n3541));
  jand g3460(.dina(n3541), .dinb(n3536), .dout(n3542));
  jxor g3461(.dina(n3542), .dinb(n56), .dout(n3543));
  jand g3462(.dina(n3228), .dinb(n3220), .dout(n3544));
  jand g3463(.dina(n3229), .dinb(n3186), .dout(n3545));
  jor  g3464(.dina(n3545), .dinb(n3544), .dout(n3546));
  jand g3465(.dina(n3016), .dinb(n2794), .dout(n3547));
  jand g3466(.dina(n2799), .dinb(n2670), .dout(n3548));
  jand g3467(.dina(n2808), .dinb(n2677), .dout(n3549));
  jand g3468(.dina(n2804), .dinb(n2672), .dout(n3550));
  jor  g3469(.dina(n3550), .dinb(n3549), .dout(n3551));
  jor  g3470(.dina(n3551), .dinb(n3548), .dout(n3552));
  jor  g3471(.dina(n3552), .dinb(n3547), .dout(n3553));
  jxor g3472(.dina(n3553), .dinb(n699), .dout(n3554));
  jand g3473(.dina(n3218), .dinb(n3197), .dout(n3555));
  jand g3474(.dina(n3219), .dinb(n3189), .dout(n3556));
  jor  g3475(.dina(n3556), .dinb(n3555), .dout(n3557));
  jor  g3476(.dina(n2857), .dinb(n2797), .dout(n3558));
  jor  g3477(.dina(n2860), .dinb(n2678), .dout(n3559));
  jor  g3478(.dina(n2865), .dinb(n2681), .dout(n3560));
  jor  g3479(.dina(n2863), .dinb(n2687), .dout(n3561));
  jand g3480(.dina(n3561), .dinb(n3560), .dout(n3562));
  jand g3481(.dina(n3562), .dinb(n3559), .dout(n3563));
  jand g3482(.dina(n3563), .dinb(n3558), .dout(n3564));
  jxor g3483(.dina(n3564), .dinb(n808), .dout(n3565));
  jand g3484(.dina(n3217), .dinb(n3210), .dout(n3566));
  jor  g3485(.dina(n3566), .dinb(n3215), .dout(n3567));
  jand g3486(.dina(n2862), .dinb(n954), .dout(n3568));
  jnot g3487(.din(n3568), .dout(n3569));
  jor  g3488(.dina(n3198), .dinb(n2874), .dout(n3570));
  jnot g3489(.din(n2688), .dout(n3571));
  jand g3490(.dina(n2889), .dinb(n3571), .dout(n3572));
  jnot g3491(.din(n2691), .dout(n3573));
  jand g3492(.dina(n2887), .dinb(n3573), .dout(n3574));
  jand g3493(.dina(n2995), .dinb(n2693), .dout(n3575));
  jor  g3494(.dina(n3575), .dinb(n3574), .dout(n3576));
  jor  g3495(.dina(n3576), .dinb(n3572), .dout(n3577));
  jnot g3496(.din(n3577), .dout(n3578));
  jand g3497(.dina(n3578), .dinb(n3570), .dout(n3579));
  jxor g3498(.dina(n3579), .dinb(n3569), .dout(n3580));
  jxor g3499(.dina(n3580), .dinb(n3567), .dout(n3581));
  jxor g3500(.dina(n3581), .dinb(n3565), .dout(n3582));
  jxor g3501(.dina(n3582), .dinb(n3557), .dout(n3583));
  jxor g3502(.dina(n3583), .dinb(n3554), .dout(n3584));
  jxor g3503(.dina(n3584), .dinb(n3546), .dout(n3585));
  jxor g3504(.dina(n3585), .dinb(n3543), .dout(n3586));
  jxor g3505(.dina(n3586), .dinb(n3535), .dout(n3587));
  jnot g3506(.din(n3319), .dout(n3588));
  jand g3507(.dina(n3588), .dinb(n3301), .dout(n3589));
  jor  g3508(.dina(n3589), .dinb(n3317), .dout(n3590));
  jand g3509(.dina(n3314), .dinb(n3303), .dout(n3591));
  jand g3510(.dina(n786), .dinb(n403), .dout(n3592));
  jnot g3511(.din(n136), .dout(n3593));
  jand g3512(.dina(n751), .dinb(n3593), .dout(n3594));
  jand g3513(.dina(n3594), .dinb(n246), .dout(n3595));
  jand g3514(.dina(n3595), .dinb(n776), .dout(n3596));
  jand g3515(.dina(n719), .dinb(n308), .dout(n3597));
  jand g3516(.dina(n3597), .dinb(n3596), .dout(n3598));
  jand g3517(.dina(n3598), .dinb(n3592), .dout(n3599));
  jxor g3518(.dina(n3599), .dinb(n3591), .dout(n3600));
  jnot g3519(.din(n3600), .dout(n3601));
  jand g3520(.dina(n3601), .dinb(n3316), .dout(n3602));
  jand g3521(.dina(n3599), .dinb(n3315), .dout(n3603));
  jor  g3522(.dina(n3603), .dinb(n3602), .dout(n3604));
  jxor g3523(.dina(n3604), .dinb(n3590), .dout(n3605));
  jor  g3524(.dina(n3605), .dinb(n3238), .dout(n3606));
  jor  g3525(.dina(n3600), .dinb(n3322), .dout(n3607));
  jor  g3526(.dina(n3325), .dinb(n3315), .dout(n3608));
  jor  g3527(.dina(n3328), .dinb(n3283), .dout(n3609));
  jand g3528(.dina(n3609), .dinb(n3608), .dout(n3610));
  jand g3529(.dina(n3610), .dinb(n3607), .dout(n3611));
  jand g3530(.dina(n3611), .dinb(n3606), .dout(n3612));
  jxor g3531(.dina(n3612), .dinb(n3233), .dout(n3613));
  jxor g3532(.dina(n3613), .dinb(n3587), .dout(n3614));
  jxor g3533(.dina(n3614), .dinb(n3532), .dout(n3615));
  jnot g3534(.din(n3615), .dout(n3616));
  jand g3535(.dina(n312), .dinb(n147), .dout(n3617));
  jand g3536(.dina(n751), .dinb(n612), .dout(n3618));
  jand g3537(.dina(n3618), .dinb(n3617), .dout(n3619));
  jand g3538(.dina(n3619), .dinb(n2490), .dout(n3620));
  jand g3539(.dina(n249), .dinb(n214), .dout(n3621));
  jand g3540(.dina(n422), .dinb(n232), .dout(n3622));
  jand g3541(.dina(n3622), .dinb(n3621), .dout(n3623));
  jand g3542(.dina(n445), .dinb(n368), .dout(n3624));
  jand g3543(.dina(n3624), .dinb(n877), .dout(n3625));
  jand g3544(.dina(n285), .dinb(n138), .dout(n3626));
  jand g3545(.dina(n3626), .dinb(n2326), .dout(n3627));
  jand g3546(.dina(n3627), .dinb(n3625), .dout(n3628));
  jand g3547(.dina(n3628), .dinb(n3623), .dout(n3629));
  jand g3548(.dina(n3629), .dinb(n3620), .dout(n3630));
  jand g3549(.dina(n426), .dinb(n421), .dout(n3631));
  jand g3550(.dina(n3631), .dinb(n1641), .dout(n3632));
  jand g3551(.dina(n3632), .dinb(n3630), .dout(n3633));
  jnot g3552(.din(n165), .dout(n3634));
  jand g3553(.dina(n454), .dinb(n295), .dout(n3635));
  jand g3554(.dina(n3635), .dinb(n3634), .dout(n3636));
  jand g3555(.dina(n3636), .dinb(n3250), .dout(n3637));
  jand g3556(.dina(n3637), .dinb(n852), .dout(n3638));
  jand g3557(.dina(n243), .dinb(n130), .dout(n3639));
  jand g3558(.dina(n592), .dinb(n270), .dout(n3640));
  jand g3559(.dina(n3640), .dinb(n3639), .dout(n3641));
  jand g3560(.dina(n2736), .dinb(n626), .dout(n3642));
  jand g3561(.dina(n3642), .dinb(n3641), .dout(n3643));
  jand g3562(.dina(n734), .dinb(n370), .dout(n3644));
  jand g3563(.dina(n3644), .dinb(n772), .dout(n3645));
  jand g3564(.dina(n3645), .dinb(n3258), .dout(n3646));
  jand g3565(.dina(n3646), .dinb(n3643), .dout(n3647));
  jand g3566(.dina(n3647), .dinb(n832), .dout(n3648));
  jand g3567(.dina(n3648), .dinb(n3638), .dout(n3649));
  jand g3568(.dina(n3649), .dinb(n3633), .dout(n3650));
  jor  g3569(.dina(n3650), .dinb(n3616), .dout(n3651));
  jxor g3570(.dina(n3650), .dinb(n3615), .dout(n3652));
  jnot g3571(.din(n3530), .dout(n3653));
  jxor g3572(.dina(n3653), .dinb(n3529), .dout(n3654));
  jand g3573(.dina(n837), .dinb(n264), .dout(n3655));
  jand g3574(.dina(n422), .dinb(n383), .dout(n3656));
  jand g3575(.dina(n3656), .dinb(n3655), .dout(n3657));
  jand g3576(.dina(n3657), .dinb(n771), .dout(n3658));
  jand g3577(.dina(n473), .dinb(n351), .dout(n3659));
  jand g3578(.dina(n3659), .dinb(n430), .dout(n3660));
  jand g3579(.dina(n3660), .dinb(n2442), .dout(n3661));
  jand g3580(.dina(n3661), .dinb(n3658), .dout(n3662));
  jand g3581(.dina(n3662), .dinb(n1292), .dout(n3663));
  jand g3582(.dina(n768), .dinb(n216), .dout(n3664));
  jand g3583(.dina(n3664), .dinb(n942), .dout(n3665));
  jand g3584(.dina(n3665), .dinb(n3663), .dout(n3666));
  jand g3585(.dina(n772), .dinb(n358), .dout(n3667));
  jand g3586(.dina(n3667), .dinb(n515), .dout(n3668));
  jand g3587(.dina(n3668), .dinb(n943), .dout(n3669));
  jand g3588(.dina(n412), .dinb(n372), .dout(n3670));
  jand g3589(.dina(n451), .dinb(n282), .dout(n3671));
  jand g3590(.dina(n3671), .dinb(n3670), .dout(n3672));
  jand g3591(.dina(n3263), .dinb(n906), .dout(n3673));
  jand g3592(.dina(n3673), .dinb(n938), .dout(n3674));
  jand g3593(.dina(n3674), .dinb(n3672), .dout(n3675));
  jand g3594(.dina(n3675), .dinb(n3669), .dout(n3676));
  jnot g3595(.din(n1676), .dout(n3677));
  jand g3596(.dina(n3677), .dinb(n463), .dout(n3678));
  jand g3597(.dina(n594), .dinb(n436), .dout(n3679));
  jand g3598(.dina(n3679), .dinb(n1228), .dout(n3680));
  jand g3599(.dina(n1196), .dinb(n619), .dout(n3681));
  jand g3600(.dina(n3681), .dinb(n3680), .dout(n3682));
  jand g3601(.dina(n3682), .dinb(n3678), .dout(n3683));
  jand g3602(.dina(n3683), .dinb(n2544), .dout(n3684));
  jand g3603(.dina(n3684), .dinb(n3676), .dout(n3685));
  jand g3604(.dina(n3685), .dinb(n3666), .dout(n3686));
  jand g3605(.dina(n3686), .dinb(n3654), .dout(n3687));
  jor  g3606(.dina(n3686), .dinb(n3654), .dout(n3688));
  jand g3607(.dina(n710), .dinb(n256), .dout(n3689));
  jand g3608(.dina(n3689), .dinb(n280), .dout(n3690));
  jand g3609(.dina(n3690), .dinb(n1673), .dout(n3691));
  jand g3610(.dina(n3691), .dinb(n2372), .dout(n3692));
  jand g3611(.dina(n3692), .dinb(n2398), .dout(n3693));
  jand g3612(.dina(n321), .dinb(n467), .dout(n3694));
  jand g3613(.dina(n3694), .dinb(n2745), .dout(n3695));
  jand g3614(.dina(n3695), .dinb(n932), .dout(n3696));
  jand g3615(.dina(n2515), .dinb(n992), .dout(n3697));
  jand g3616(.dina(n2521), .dinb(n728), .dout(n3698));
  jand g3617(.dina(n3698), .dinb(n3697), .dout(n3699));
  jand g3618(.dina(n214), .dinb(n138), .dout(n3700));
  jand g3619(.dina(n3700), .dinb(n153), .dout(n3701));
  jand g3620(.dina(n441), .dinb(n304), .dout(n3702));
  jand g3621(.dina(n488), .dinb(n261), .dout(n3703));
  jand g3622(.dina(n3703), .dinb(n3702), .dout(n3704));
  jand g3623(.dina(n3704), .dinb(n3701), .dout(n3705));
  jand g3624(.dina(n3705), .dinb(n3699), .dout(n3706));
  jand g3625(.dina(n3706), .dinb(n2466), .dout(n3707));
  jand g3626(.dina(n3707), .dinb(n3696), .dout(n3708));
  jand g3627(.dina(n3708), .dinb(n3693), .dout(n3709));
  jnot g3628(.din(n3347), .dout(n3710));
  jnot g3629(.din(n3513), .dout(n3711));
  jnot g3630(.din(n3348), .dout(n3712));
  jnot g3631(.din(n3497), .dout(n3713));
  jnot g3632(.din(n3349), .dout(n3714));
  jnot g3633(.din(n3485), .dout(n3715));
  jnot g3634(.din(n3350), .dout(n3716));
  jnot g3635(.din(n3467), .dout(n3717));
  jnot g3636(.din(n3351), .dout(n3718));
  jnot g3637(.din(n3455), .dout(n3719));
  jnot g3638(.din(n3352), .dout(n3720));
  jnot g3639(.din(n3438), .dout(n3721));
  jnot g3640(.din(n3353), .dout(n3722));
  jnot g3641(.din(n3426), .dout(n3723));
  jnot g3642(.din(n3354), .dout(n3724));
  jnot g3643(.din(n3421), .dout(n3725));
  jnot g3644(.din(n3362), .dout(n3726));
  jnot g3645(.din(n3409), .dout(n3727));
  jnot g3646(.din(n3365), .dout(n3728));
  jnot g3647(.din(n3397), .dout(n3729));
  jnot g3648(.din(n3367), .dout(n3730));
  jnot g3649(.din(n3379), .dout(n3731));
  jand g3650(.dina(n3375), .dinb(n68), .dout(n3732));
  jnot g3651(.din(n3394), .dout(n3733));
  jor  g3652(.dina(n3733), .dinb(n3732), .dout(n3734));
  jor  g3653(.dina(n3734), .dinb(n3731), .dout(n3735));
  jand g3654(.dina(n3735), .dinb(n3730), .dout(n3736));
  jnot g3655(.din(n3406), .dout(n3737));
  jor  g3656(.dina(n3737), .dinb(n3736), .dout(n3738));
  jand g3657(.dina(n3738), .dinb(n3729), .dout(n3739));
  jor  g3658(.dina(n3739), .dinb(n3728), .dout(n3740));
  jnot g3659(.din(n3418), .dout(n3741));
  jand g3660(.dina(n3741), .dinb(n3740), .dout(n3742));
  jor  g3661(.dina(n3742), .dinb(n3727), .dout(n3743));
  jand g3662(.dina(n3743), .dinb(n3726), .dout(n3744));
  jnot g3663(.din(n3423), .dout(n3745));
  jor  g3664(.dina(n3745), .dinb(n3744), .dout(n3746));
  jand g3665(.dina(n3746), .dinb(n3725), .dout(n3747));
  jor  g3666(.dina(n3747), .dinb(n3724), .dout(n3748));
  jnot g3667(.din(n3435), .dout(n3749));
  jand g3668(.dina(n3749), .dinb(n3748), .dout(n3750));
  jor  g3669(.dina(n3750), .dinb(n3723), .dout(n3751));
  jand g3670(.dina(n3751), .dinb(n3722), .dout(n3752));
  jnot g3671(.din(n3452), .dout(n3753));
  jor  g3672(.dina(n3753), .dinb(n3752), .dout(n3754));
  jand g3673(.dina(n3754), .dinb(n3721), .dout(n3755));
  jand g3674(.dina(n3755), .dinb(n3720), .dout(n3756));
  jnot g3675(.din(n3464), .dout(n3757));
  jor  g3676(.dina(n3757), .dinb(n3756), .dout(n3758));
  jand g3677(.dina(n3758), .dinb(n3719), .dout(n3759));
  jand g3678(.dina(n3759), .dinb(n3718), .dout(n3760));
  jnot g3679(.din(n3482), .dout(n3761));
  jor  g3680(.dina(n3761), .dinb(n3760), .dout(n3762));
  jand g3681(.dina(n3762), .dinb(n3717), .dout(n3763));
  jor  g3682(.dina(n3763), .dinb(n3716), .dout(n3764));
  jnot g3683(.din(n3494), .dout(n3765));
  jand g3684(.dina(n3765), .dinb(n3764), .dout(n3766));
  jor  g3685(.dina(n3766), .dinb(n3715), .dout(n3767));
  jand g3686(.dina(n3767), .dinb(n3714), .dout(n3768));
  jnot g3687(.din(n3510), .dout(n3769));
  jor  g3688(.dina(n3769), .dinb(n3768), .dout(n3770));
  jand g3689(.dina(n3770), .dinb(n3713), .dout(n3771));
  jor  g3690(.dina(n3771), .dinb(n3712), .dout(n3772));
  jand g3691(.dina(n3524), .dinb(n3772), .dout(n3773));
  jor  g3692(.dina(n3773), .dinb(n3711), .dout(n3774));
  jand g3693(.dina(n3774), .dinb(n3710), .dout(n3775));
  jor  g3694(.dina(n3775), .dinb(n3709), .dout(n3776));
  jor  g3695(.dina(n3776), .dinb(n3528), .dout(n3777));
  jand g3696(.dina(n3777), .dinb(n3688), .dout(n3778));
  jor  g3697(.dina(n3778), .dinb(n3687), .dout(n3779));
  jor  g3698(.dina(n3779), .dinb(n3652), .dout(n3780));
  jand g3699(.dina(n3780), .dinb(n3651), .dout(n3781));
  jand g3700(.dina(n3613), .dinb(n3587), .dout(n3782));
  jand g3701(.dina(n3614), .dinb(n3532), .dout(n3783));
  jor  g3702(.dina(n3783), .dinb(n3782), .dout(n3784));
  jnot g3703(.din(n3604), .dout(n3785));
  jand g3704(.dina(n3785), .dinb(n3590), .dout(n3786));
  jor  g3705(.dina(n3786), .dinb(n3602), .dout(n3787));
  jand g3706(.dina(n3599), .dinb(n3591), .dout(n3788));
  jand g3707(.dina(n397), .dinb(n243), .dout(n3789));
  jand g3708(.dina(n679), .dinb(n277), .dout(n3790));
  jand g3709(.dina(n3790), .dinb(n3789), .dout(n3791));
  jand g3710(.dina(n2331), .dinb(n869), .dout(n3792));
  jand g3711(.dina(n3792), .dinb(n3624), .dout(n3793));
  jand g3712(.dina(n3793), .dinb(n3791), .dout(n3794));
  jand g3713(.dina(n2511), .dinb(n758), .dout(n3795));
  jnot g3714(.din(n578), .dout(n3796));
  jand g3715(.dina(n2339), .dinb(n3796), .dout(n3797));
  jand g3716(.dina(n3797), .dinb(n3795), .dout(n3798));
  jand g3717(.dina(n825), .dinb(n249), .dout(n3799));
  jand g3718(.dina(n3799), .dinb(n421), .dout(n3800));
  jand g3719(.dina(n3800), .dinb(n880), .dout(n3801));
  jand g3720(.dina(n3801), .dinb(n3798), .dout(n3802));
  jand g3721(.dina(n3802), .dinb(n2743), .dout(n3803));
  jand g3722(.dina(n3803), .dinb(n3794), .dout(n3804));
  jand g3723(.dina(n3804), .dinb(n1319), .dout(n3805));
  jxor g3724(.dina(n3805), .dinb(n3788), .dout(n3806));
  jnot g3725(.din(n3806), .dout(n3807));
  jand g3726(.dina(n3807), .dinb(n3601), .dout(n3808));
  jand g3727(.dina(n3805), .dinb(n3600), .dout(n3809));
  jor  g3728(.dina(n3809), .dinb(n3808), .dout(n3810));
  jxor g3729(.dina(n3810), .dinb(n3787), .dout(n3811));
  jor  g3730(.dina(n3811), .dinb(n3238), .dout(n3812));
  jor  g3731(.dina(n3806), .dinb(n3322), .dout(n3813));
  jor  g3732(.dina(n3600), .dinb(n3325), .dout(n3814));
  jor  g3733(.dina(n3328), .dinb(n3315), .dout(n3815));
  jand g3734(.dina(n3815), .dinb(n3814), .dout(n3816));
  jand g3735(.dina(n3816), .dinb(n3813), .dout(n3817));
  jand g3736(.dina(n3817), .dinb(n3812), .dout(n3818));
  jxor g3737(.dina(n3818), .dinb(n68), .dout(n3819));
  jnot g3738(.din(n3819), .dout(n3820));
  jand g3739(.dina(n3585), .dinb(n3543), .dout(n3821));
  jand g3740(.dina(n3586), .dinb(n3535), .dout(n3822));
  jor  g3741(.dina(n3822), .dinb(n3821), .dout(n3823));
  jand g3742(.dina(n3583), .dinb(n3554), .dout(n3824));
  jand g3743(.dina(n3584), .dinb(n3546), .dout(n3825));
  jor  g3744(.dina(n3825), .dinb(n3824), .dout(n3826));
  jor  g3745(.dina(n2795), .dinb(n2771), .dout(n3827));
  jor  g3746(.dina(n2800), .dinb(n2773), .dout(n3828));
  jor  g3747(.dina(n2805), .dinb(n2669), .dout(n3829));
  jor  g3748(.dina(n2809), .dinb(n2671), .dout(n3830));
  jand g3749(.dina(n3830), .dinb(n3829), .dout(n3831));
  jand g3750(.dina(n3831), .dinb(n3828), .dout(n3832));
  jand g3751(.dina(n3832), .dinb(n3827), .dout(n3833));
  jxor g3752(.dina(n3833), .dinb(n699), .dout(n3834));
  jnot g3753(.din(n3834), .dout(n3835));
  jand g3754(.dina(n3581), .dinb(n3565), .dout(n3836));
  jand g3755(.dina(n3582), .dinb(n3557), .dout(n3837));
  jor  g3756(.dina(n3837), .dinb(n3836), .dout(n3838));
  jand g3757(.dina(n2694), .dinb(n954), .dout(n3839));
  jnot g3758(.din(n3839), .dout(n3840));
  jor  g3759(.dina(n2911), .dinb(n3198), .dout(n3841));
  jand g3760(.dina(n2889), .dinb(n2685), .dout(n3842));
  jand g3761(.dina(n2887), .dinb(n3571), .dout(n3843));
  jand g3762(.dina(n2995), .dinb(n3573), .dout(n3844));
  jor  g3763(.dina(n3844), .dinb(n3843), .dout(n3845));
  jor  g3764(.dina(n3845), .dinb(n3842), .dout(n3846));
  jnot g3765(.din(n3846), .dout(n3847));
  jand g3766(.dina(n3847), .dinb(n3841), .dout(n3848));
  jxor g3767(.dina(n3848), .dinb(n3840), .dout(n3849));
  jand g3768(.dina(n3580), .dinb(n3567), .dout(n3850));
  jand g3769(.dina(n2700), .dinb(n954), .dout(n3851));
  jand g3770(.dina(n3851), .dinb(n3579), .dout(n3852));
  jor  g3771(.dina(n3852), .dinb(n3850), .dout(n3853));
  jxor g3772(.dina(n3853), .dinb(n3849), .dout(n3854));
  jand g3773(.dina(n3004), .dinb(n2828), .dout(n3855));
  jand g3774(.dina(n2834), .dinb(n2677), .dout(n3856));
  jand g3775(.dina(n2848), .dinb(n2684), .dout(n3857));
  jand g3776(.dina(n2832), .dinb(n2679), .dout(n3858));
  jor  g3777(.dina(n3858), .dinb(n3857), .dout(n3859));
  jor  g3778(.dina(n3859), .dinb(n3856), .dout(n3860));
  jor  g3779(.dina(n3860), .dinb(n3855), .dout(n3861));
  jxor g3780(.dina(n3861), .dinb(n803), .dout(n3862));
  jxor g3781(.dina(n3862), .dinb(n3854), .dout(n3863));
  jxor g3782(.dina(n3863), .dinb(n3838), .dout(n3864));
  jxor g3783(.dina(n3864), .dinb(n3835), .dout(n3865));
  jxor g3784(.dina(n3865), .dinb(n3826), .dout(n3866));
  jor  g3785(.dina(n3337), .dinb(n79), .dout(n3867));
  jor  g3786(.dina(n3283), .dinb(n2775), .dout(n3868));
  jor  g3787(.dina(n3284), .dinb(n2780), .dout(n3869));
  jor  g3788(.dina(n3172), .dinb(n2784), .dout(n3870));
  jand g3789(.dina(n3870), .dinb(n3869), .dout(n3871));
  jand g3790(.dina(n3871), .dinb(n3868), .dout(n3872));
  jand g3791(.dina(n3872), .dinb(n3867), .dout(n3873));
  jxor g3792(.dina(n3873), .dinb(n56), .dout(n3874));
  jxor g3793(.dina(n3874), .dinb(n3866), .dout(n3875));
  jxor g3794(.dina(n3875), .dinb(n3823), .dout(n3876));
  jxor g3795(.dina(n3876), .dinb(n3820), .dout(n3877));
  jxor g3796(.dina(n3877), .dinb(n3784), .dout(n3878));
  jand g3797(.dina(n3258), .dinb(n1187), .dout(n3879));
  jand g3798(.dina(n3879), .dinb(n1646), .dout(n3880));
  jand g3799(.dina(n458), .dinb(n264), .dout(n3881));
  jand g3800(.dina(n3881), .dinb(n147), .dout(n3882));
  jand g3801(.dina(n3624), .dinb(n2360), .dout(n3883));
  jand g3802(.dina(n3883), .dinb(n3882), .dout(n3884));
  jand g3803(.dina(n3884), .dinb(n1020), .dout(n3885));
  jand g3804(.dina(n3885), .dinb(n3880), .dout(n3886));
  jand g3805(.dina(n3886), .dinb(n902), .dout(n3887));
  jand g3806(.dina(n3887), .dinb(n2391), .dout(n3888));
  jxor g3807(.dina(n3888), .dinb(n3878), .dout(n3889));
  jxor g3808(.dina(n3889), .dinb(n3781), .dout(n3890));
  jxor g3809(.dina(n3779), .dinb(n3652), .dout(n3891));
  jxor g3810(.dina(n3891), .dinb(n3890), .dout(sin0 ));
  jnot g3811(.din(n3878), .dout(n3893));
  jor  g3812(.dina(n3888), .dinb(n3893), .dout(n3894));
  jor  g3813(.dina(n3889), .dinb(n3781), .dout(n3895));
  jand g3814(.dina(n3895), .dinb(n3894), .dout(n3896));
  jand g3815(.dina(n3876), .dinb(n3820), .dout(n3897));
  jand g3816(.dina(n3877), .dinb(n3784), .dout(n3898));
  jor  g3817(.dina(n3898), .dinb(n3897), .dout(n3899));
  jnot g3818(.din(n3810), .dout(n3900));
  jand g3819(.dina(n3900), .dinb(n3787), .dout(n3901));
  jor  g3820(.dina(n3901), .dinb(n3808), .dout(n3902));
  jand g3821(.dina(n592), .dinb(n454), .dout(n3904));
  jand g3822(.dina(n3904), .dinb(n2326), .dout(n3905));
  jand g3823(.dina(n2521), .dinb(n417), .dout(n3906));
  jand g3824(.dina(n3906), .dinb(n846), .dout(n3907));
  jand g3825(.dina(n3907), .dinb(n3905), .dout(n3908));
  jand g3826(.dina(n3908), .dinb(n754), .dout(n3909));
  jnot g3827(.din(n1679), .dout(n3910));
  jand g3828(.dina(n3274), .dinb(n493), .dout(n3911));
  jand g3829(.dina(n463), .dinb(n351), .dout(n3912));
  jand g3830(.dina(n3912), .dinb(n2380), .dout(n3913));
  jand g3831(.dina(n3913), .dinb(n855), .dout(n3914));
  jand g3832(.dina(n3914), .dinb(n3911), .dout(n3915));
  jand g3833(.dina(n3915), .dinb(n3910), .dout(n3916));
  jand g3834(.dina(n3916), .dinb(n933), .dout(n3917));
  jand g3835(.dina(n3917), .dinb(n3909), .dout(n3918));
  jand g3836(.dina(n3918), .dinb(n2520), .dout(n3919));
  jnot g3837(.din(n3919), .dout(n3920));
  jand g3838(.dina(n3919), .dinb(n3807), .dout(n3923));
  jand g3839(.dina(n3920), .dinb(n3806), .dout(n3924));
  jor  g3840(.dina(n3924), .dinb(n3923), .dout(n3925));
  jnot g3841(.din(n3925), .dout(n3926));
  jxor g3842(.dina(n3926), .dinb(n3902), .dout(n3927));
  jor  g3843(.dina(n3927), .dinb(n3238), .dout(n3928));
  jor  g3844(.dina(n3919), .dinb(n3322), .dout(n3929));
  jor  g3845(.dina(n3806), .dinb(n3325), .dout(n3930));
  jor  g3846(.dina(n3600), .dinb(n3328), .dout(n3931));
  jand g3847(.dina(n3931), .dinb(n3930), .dout(n3932));
  jand g3848(.dina(n3932), .dinb(n3929), .dout(n3933));
  jand g3849(.dina(n3933), .dinb(n3928), .dout(n3934));
  jxor g3850(.dina(n3934), .dinb(n68), .dout(n3935));
  jnot g3851(.din(n3935), .dout(n3936));
  jand g3852(.dina(n3874), .dinb(n3866), .dout(n3937));
  jand g3853(.dina(n3875), .dinb(n3823), .dout(n3938));
  jor  g3854(.dina(n3938), .dinb(n3937), .dout(n3939));
  jand g3855(.dina(n3864), .dinb(n3835), .dout(n3940));
  jand g3856(.dina(n3865), .dinb(n3826), .dout(n3941));
  jor  g3857(.dina(n3941), .dinb(n3940), .dout(n3942));
  jand g3858(.dina(n3174), .dinb(n2794), .dout(n3943));
  jand g3859(.dina(n3176), .dinb(n2799), .dout(n3944));
  jand g3860(.dina(n2808), .dinb(n2670), .dout(n3945));
  jand g3861(.dina(n2804), .dinb(n2769), .dout(n3946));
  jor  g3862(.dina(n3946), .dinb(n3945), .dout(n3947));
  jor  g3863(.dina(n3947), .dinb(n3944), .dout(n3948));
  jor  g3864(.dina(n3948), .dinb(n3943), .dout(n3949));
  jxor g3865(.dina(n3949), .dinb(n1143), .dout(n3950));
  jnot g3866(.din(n3950), .dout(n3951));
  jand g3867(.dina(n3862), .dinb(n3854), .dout(n3952));
  jand g3868(.dina(n3863), .dinb(n3838), .dout(n3953));
  jor  g3869(.dina(n3953), .dinb(n3952), .dout(n3954));
  jor  g3870(.dina(n3028), .dinb(n2857), .dout(n3955));
  jor  g3871(.dina(n2860), .dinb(n2671), .dout(n3956));
  jor  g3872(.dina(n2865), .dinb(n2674), .dout(n3957));
  jor  g3873(.dina(n2863), .dinb(n2678), .dout(n3958));
  jand g3874(.dina(n3958), .dinb(n3957), .dout(n3959));
  jand g3875(.dina(n3959), .dinb(n3956), .dout(n3960));
  jand g3876(.dina(n3960), .dinb(n3955), .dout(n3961));
  jxor g3877(.dina(n3961), .dinb(n808), .dout(n3962));
  jand g3878(.dina(n2691), .dinb(n954), .dout(n3963));
  jnot g3879(.din(n3963), .dout(n3964));
  jor  g3880(.dina(n2899), .dinb(n3198), .dout(n3965));
  jand g3881(.dina(n2889), .dinb(n2684), .dout(n3966));
  jand g3882(.dina(n2887), .dinb(n2685), .dout(n3967));
  jand g3883(.dina(n2995), .dinb(n3571), .dout(n3968));
  jor  g3884(.dina(n3968), .dinb(n3967), .dout(n3969));
  jor  g3885(.dina(n3969), .dinb(n3966), .dout(n3970));
  jnot g3886(.din(n3970), .dout(n3971));
  jand g3887(.dina(n3971), .dinb(n3965), .dout(n3972));
  jxor g3888(.dina(n3972), .dinb(n3964), .dout(n3973));
  jand g3889(.dina(n3853), .dinb(n3849), .dout(n3974));
  jand g3890(.dina(n2693), .dinb(n954), .dout(n3975));
  jand g3891(.dina(n3975), .dinb(n3848), .dout(n3976));
  jor  g3892(.dina(n3976), .dinb(n3974), .dout(n3977));
  jxor g3893(.dina(n3977), .dinb(n3973), .dout(n3978));
  jxor g3894(.dina(n3978), .dinb(n3962), .dout(n3979));
  jxor g3895(.dina(n3979), .dinb(n3954), .dout(n3980));
  jxor g3896(.dina(n3980), .dinb(n3951), .dout(n3981));
  jxor g3897(.dina(n3981), .dinb(n3942), .dout(n3982));
  jor  g3898(.dina(n3320), .dinb(n79), .dout(n3983));
  jor  g3899(.dina(n3315), .dinb(n2775), .dout(n3984));
  jor  g3900(.dina(n3283), .dinb(n2780), .dout(n3985));
  jor  g3901(.dina(n3284), .dinb(n2784), .dout(n3986));
  jand g3902(.dina(n3986), .dinb(n3985), .dout(n3987));
  jand g3903(.dina(n3987), .dinb(n3984), .dout(n3988));
  jand g3904(.dina(n3988), .dinb(n3983), .dout(n3989));
  jxor g3905(.dina(n3989), .dinb(n56), .dout(n3990));
  jxor g3906(.dina(n3990), .dinb(n3982), .dout(n3991));
  jxor g3907(.dina(n3991), .dinb(n3939), .dout(n3992));
  jxor g3908(.dina(n3992), .dinb(n3936), .dout(n3993));
  jxor g3909(.dina(n3993), .dinb(n3899), .dout(n3994));
  jand g3910(.dina(n1018), .dinb(n417), .dout(n3995));
  jand g3911(.dina(n2457), .dinb(n2429), .dout(n3996));
  jand g3912(.dina(n3996), .dinb(n3995), .dout(n3997));
  jnot g3913(.din(n1658), .dout(n3998));
  jand g3914(.dina(n1209), .dinb(n241), .dout(n3999));
  jand g3915(.dina(n3999), .dinb(n3998), .dout(n4000));
  jand g3916(.dina(n592), .dinb(n430), .dout(n4001));
  jand g3917(.dina(n632), .dinb(n321), .dout(n4002));
  jand g3918(.dina(n4002), .dinb(n4001), .dout(n4003));
  jand g3919(.dina(n4003), .dinb(n4000), .dout(n4004));
  jand g3920(.dina(n3258), .dinb(n3242), .dout(n4005));
  jand g3921(.dina(n4005), .dinb(n4004), .dout(n4006));
  jand g3922(.dina(n4006), .dinb(n3997), .dout(n4007));
  jand g3923(.dina(n4007), .dinb(n3630), .dout(n4008));
  jand g3924(.dina(n4008), .dinb(n2359), .dout(n4009));
  jxor g3925(.dina(n4009), .dinb(n3994), .dout(n4010));
  jxor g3926(.dina(n4010), .dinb(n3896), .dout(n4011));
  jnot g3927(.din(n4011), .dout(n4012));
  jxor g3928(.dina(a23 ), .dinb(a22 ), .dout(n4013));
  jand g3929(.dina(n4013), .dinb(sin0 ), .dout(n4014));
  jand g3930(.dina(n4014), .dinb(n4012), .dout(n4015));
  jnot g3931(.din(n4014), .dout(n4016));
  jand g3932(.dina(n3891), .dinb(n3890), .dout(n4017));
  jxor g3933(.dina(n4011), .dinb(n4017), .dout(n4018));
  jand g3934(.dina(n4018), .dinb(n4016), .dout(n4019));
  jor  g3935(.dina(n4019), .dinb(n4015), .dout(sin1 ));
  jand g3936(.dina(n4011), .dinb(n4017), .dout(n4021));
  jnot g3937(.din(n3994), .dout(n4022));
  jor  g3938(.dina(n4009), .dinb(n4022), .dout(n4023));
  jor  g3939(.dina(n4010), .dinb(n3896), .dout(n4024));
  jand g3940(.dina(n4024), .dinb(n4023), .dout(n4025));
  jand g3941(.dina(n3992), .dinb(n3936), .dout(n4026));
  jand g3942(.dina(n3993), .dinb(n3899), .dout(n4027));
  jor  g3943(.dina(n4027), .dinb(n4026), .dout(n4028));
  jand g3944(.dina(n3990), .dinb(n3982), .dout(n4029));
  jand g3945(.dina(n3991), .dinb(n3939), .dout(n4030));
  jor  g3946(.dina(n4030), .dinb(n4029), .dout(n4031));
  jand g3947(.dina(n3980), .dinb(n3951), .dout(n4032));
  jand g3948(.dina(n3981), .dinb(n3942), .dout(n4033));
  jor  g3949(.dina(n4033), .dinb(n4032), .dout(n4034));
  jor  g3950(.dina(n3516), .dinb(n2795), .dout(n4035));
  jor  g3951(.dina(n3284), .dinb(n2800), .dout(n4036));
  jor  g3952(.dina(n3172), .dinb(n2805), .dout(n4037));
  jor  g3953(.dina(n2809), .dinb(n2773), .dout(n4038));
  jand g3954(.dina(n4038), .dinb(n4037), .dout(n4039));
  jand g3955(.dina(n4039), .dinb(n4036), .dout(n4040));
  jand g3956(.dina(n4040), .dinb(n4035), .dout(n4041));
  jxor g3957(.dina(n4041), .dinb(n699), .dout(n4042));
  jnot g3958(.din(n4042), .dout(n4043));
  jand g3959(.dina(n3978), .dinb(n3962), .dout(n4044));
  jand g3960(.dina(n3979), .dinb(n3954), .dout(n4045));
  jor  g3961(.dina(n4045), .dinb(n4044), .dout(n4046));
  jand g3962(.dina(n3016), .dinb(n2828), .dout(n4047));
  jand g3963(.dina(n2834), .dinb(n2670), .dout(n4048));
  jand g3964(.dina(n2848), .dinb(n2677), .dout(n4049));
  jand g3965(.dina(n2832), .dinb(n2672), .dout(n4050));
  jor  g3966(.dina(n4050), .dinb(n4049), .dout(n4051));
  jor  g3967(.dina(n4051), .dinb(n4048), .dout(n4052));
  jor  g3968(.dina(n4052), .dinb(n4047), .dout(n4053));
  jxor g3969(.dina(n4053), .dinb(n803), .dout(n4054));
  jand g3970(.dina(n2688), .dinb(n954), .dout(n4055));
  jnot g3971(.din(n4055), .dout(n4056));
  jor  g3972(.dina(n3198), .dinb(n2797), .dout(n4057));
  jand g3973(.dina(n2889), .dinb(n2679), .dout(n4058));
  jand g3974(.dina(n2887), .dinb(n2684), .dout(n4059));
  jand g3975(.dina(n2995), .dinb(n2685), .dout(n4060));
  jor  g3976(.dina(n4060), .dinb(n4059), .dout(n4061));
  jor  g3977(.dina(n4061), .dinb(n4058), .dout(n4062));
  jnot g3978(.din(n4062), .dout(n4063));
  jand g3979(.dina(n4063), .dinb(n4057), .dout(n4064));
  jxor g3980(.dina(n4064), .dinb(n4056), .dout(n4065));
  jand g3981(.dina(n3977), .dinb(n3973), .dout(n4066));
  jand g3982(.dina(n3573), .dinb(n954), .dout(n4067));
  jand g3983(.dina(n4067), .dinb(n3972), .dout(n4068));
  jor  g3984(.dina(n4068), .dinb(n4066), .dout(n4069));
  jxor g3985(.dina(n4069), .dinb(n4065), .dout(n4070));
  jxor g3986(.dina(n4070), .dinb(n4054), .dout(n4071));
  jxor g3987(.dina(n4071), .dinb(n4046), .dout(n4072));
  jxor g3988(.dina(n4072), .dinb(n4043), .dout(n4073));
  jxor g3989(.dina(n4073), .dinb(n4034), .dout(n4074));
  jor  g3990(.dina(n3605), .dinb(n79), .dout(n4075));
  jor  g3991(.dina(n3600), .dinb(n2775), .dout(n4076));
  jor  g3992(.dina(n3315), .dinb(n2780), .dout(n4077));
  jor  g3993(.dina(n3283), .dinb(n2784), .dout(n4078));
  jand g3994(.dina(n4078), .dinb(n4077), .dout(n4079));
  jand g3995(.dina(n4079), .dinb(n4076), .dout(n4080));
  jand g3996(.dina(n4080), .dinb(n4075), .dout(n4081));
  jxor g3997(.dina(n4081), .dinb(n56), .dout(n4082));
  jxor g3998(.dina(n4082), .dinb(n4074), .dout(n4083));
  jxor g3999(.dina(n4083), .dinb(n4031), .dout(n4084));
  jand g4000(.dina(n3920), .dinb(n3324), .dout(n4085));
  jand g4001(.dina(n3925), .dinb(n3902), .dout(n4086));
  jand g4002(.dina(n4086), .dinb(n3919), .dout(n4087));
  jnot g4003(.din(n4086), .dout(n4088));
  jand g4004(.dina(n4088), .dinb(n3924), .dout(n4089));
  jor  g4005(.dina(n4089), .dinb(n4087), .dout(n4090));
  jand g4006(.dina(n4090), .dinb(n3237), .dout(n4091));
  jor  g4007(.dina(n4091), .dinb(n4085), .dout(n4092));
  jand g4008(.dina(n3807), .dinb(n63), .dout(n4093));
  jor  g4009(.dina(n4093), .dinb(n3233), .dout(n4094));
  jnot g4010(.din(n4094), .dout(n4095));
  jor  g4011(.dina(n4095), .dinb(n4092), .dout(n4096));
  jnot g4012(.din(n4092), .dout(n4097));
  jor  g4013(.dina(n4097), .dinb(n3233), .dout(n4098));
  jand g4014(.dina(n4098), .dinb(n4096), .dout(n4099));
  jxor g4015(.dina(n4099), .dinb(n4084), .dout(n4100));
  jxor g4016(.dina(n4100), .dinb(n4028), .dout(n4101));
  jand g4017(.dina(n294), .dinb(n229), .dout(n4102));
  jand g4018(.dina(n4102), .dinb(n825), .dout(n4103));
  jand g4019(.dina(n412), .dinb(n270), .dout(n4104));
  jand g4020(.dina(n4104), .dinb(n2734), .dout(n4105));
  jand g4021(.dina(n4105), .dinb(n4103), .dout(n4106));
  jand g4022(.dina(n744), .dinb(n282), .dout(n4107));
  jand g4023(.dina(n4107), .dinb(n265), .dout(n4108));
  jand g4024(.dina(n4108), .dinb(n988), .dout(n4109));
  jand g4025(.dina(n2380), .dinb(n732), .dout(n4110));
  jand g4026(.dina(n4110), .dinb(n374), .dout(n4111));
  jand g4027(.dina(n4111), .dinb(n999), .dout(n4112));
  jand g4028(.dina(n4112), .dinb(n4109), .dout(n4113));
  jand g4029(.dina(n4113), .dinb(n4106), .dout(n4114));
  jand g4030(.dina(n4114), .dinb(n923), .dout(n4115));
  jand g4031(.dina(n4115), .dinb(n3693), .dout(n4116));
  jxor g4032(.dina(n4116), .dinb(n4101), .dout(n4117));
  jxor g4033(.dina(n4117), .dinb(n4025), .dout(n4118));
  jxor g4034(.dina(n4118), .dinb(n4021), .dout(n4119));
  jor  g4035(.dina(n4018), .dinb(sin0 ), .dout(n4120));
  jand g4036(.dina(n4120), .dinb(n4013), .dout(n4121));
  jxor g4037(.dina(n4121), .dinb(n4119), .dout(sin2 ));
  jor  g4038(.dina(n4120), .dinb(n4119), .dout(n4123));
  jand g4039(.dina(n4123), .dinb(n4013), .dout(n4124));
  jand g4040(.dina(n4118), .dinb(n4021), .dout(n4125));
  jnot g4041(.din(n4101), .dout(n4126));
  jor  g4042(.dina(n4116), .dinb(n4126), .dout(n4127));
  jor  g4043(.dina(n4117), .dinb(n4025), .dout(n4128));
  jand g4044(.dina(n4128), .dinb(n4127), .dout(n4129));
  jand g4045(.dina(n4099), .dinb(n4084), .dout(n4130));
  jand g4046(.dina(n4100), .dinb(n4028), .dout(n4131));
  jor  g4047(.dina(n4131), .dinb(n4130), .dout(n4132));
  jand g4048(.dina(n4082), .dinb(n4074), .dout(n4133));
  jand g4049(.dina(n4083), .dinb(n4031), .dout(n4134));
  jor  g4050(.dina(n4134), .dinb(n4133), .dout(n4135));
  jand g4051(.dina(n4088), .dinb(n3806), .dout(n4136));
  jor  g4052(.dina(n4136), .dinb(n3238), .dout(n4137));
  jand g4053(.dina(n4137), .dinb(n3328), .dout(n4138));
  jor  g4054(.dina(n4138), .dinb(n3919), .dout(n4139));
  jxor g4055(.dina(n4139), .dinb(n68), .dout(n4140));
  jnot g4056(.din(n4140), .dout(n4141));
  jand g4057(.dina(n4072), .dinb(n4043), .dout(n4142));
  jand g4058(.dina(n4073), .dinb(n4034), .dout(n4143));
  jor  g4059(.dina(n4143), .dinb(n4142), .dout(n4144));
  jor  g4060(.dina(n3337), .dinb(n2795), .dout(n4145));
  jor  g4061(.dina(n3283), .dinb(n2800), .dout(n4146));
  jor  g4062(.dina(n3284), .dinb(n2805), .dout(n4147));
  jor  g4063(.dina(n3172), .dinb(n2809), .dout(n4148));
  jand g4064(.dina(n4148), .dinb(n4147), .dout(n4149));
  jand g4065(.dina(n4149), .dinb(n4146), .dout(n4150));
  jand g4066(.dina(n4150), .dinb(n4145), .dout(n4151));
  jxor g4067(.dina(n4151), .dinb(n699), .dout(n4152));
  jnot g4068(.din(n4152), .dout(n4153));
  jand g4069(.dina(n4070), .dinb(n4054), .dout(n4154));
  jand g4070(.dina(n4071), .dinb(n4046), .dout(n4155));
  jor  g4071(.dina(n4155), .dinb(n4154), .dout(n4156));
  jor  g4072(.dina(n2857), .dinb(n2771), .dout(n4157));
  jor  g4073(.dina(n2860), .dinb(n2773), .dout(n4158));
  jor  g4074(.dina(n2865), .dinb(n2669), .dout(n4159));
  jor  g4075(.dina(n2863), .dinb(n2671), .dout(n4160));
  jand g4076(.dina(n4160), .dinb(n4159), .dout(n4161));
  jand g4077(.dina(n4161), .dinb(n4158), .dout(n4162));
  jand g4078(.dina(n4162), .dinb(n4157), .dout(n4163));
  jxor g4079(.dina(n4163), .dinb(n808), .dout(n4164));
  jand g4080(.dina(n2687), .dinb(n954), .dout(n4165));
  jand g4081(.dina(n3004), .dinb(n2883), .dout(n4166));
  jand g4082(.dina(n2889), .dinb(n2677), .dout(n4167));
  jand g4083(.dina(n2995), .dinb(n2684), .dout(n4168));
  jand g4084(.dina(n2887), .dinb(n2679), .dout(n4169));
  jor  g4085(.dina(n4169), .dinb(n4168), .dout(n4170));
  jor  g4086(.dina(n4170), .dinb(n4167), .dout(n4171));
  jor  g4087(.dina(n4171), .dinb(n4166), .dout(n4172));
  jxor g4088(.dina(n4172), .dinb(n4165), .dout(n4173));
  jand g4089(.dina(n4069), .dinb(n4065), .dout(n4174));
  jand g4090(.dina(n3571), .dinb(n954), .dout(n4175));
  jand g4091(.dina(n4175), .dinb(n4064), .dout(n4176));
  jor  g4092(.dina(n4176), .dinb(n4174), .dout(n4177));
  jxor g4093(.dina(n4177), .dinb(n4173), .dout(n4178));
  jxor g4094(.dina(n4178), .dinb(n4164), .dout(n4179));
  jxor g4095(.dina(n4179), .dinb(n4156), .dout(n4180));
  jxor g4096(.dina(n4180), .dinb(n4153), .dout(n4181));
  jxor g4097(.dina(n4181), .dinb(n4144), .dout(n4182));
  jor  g4098(.dina(n3811), .dinb(n79), .dout(n4183));
  jor  g4099(.dina(n3806), .dinb(n2775), .dout(n4184));
  jor  g4100(.dina(n3600), .dinb(n2780), .dout(n4185));
  jor  g4101(.dina(n3315), .dinb(n2784), .dout(n4186));
  jand g4102(.dina(n4186), .dinb(n4185), .dout(n4187));
  jand g4103(.dina(n4187), .dinb(n4184), .dout(n4188));
  jand g4104(.dina(n4188), .dinb(n4183), .dout(n4189));
  jxor g4105(.dina(n4189), .dinb(n56), .dout(n4190));
  jxor g4106(.dina(n4190), .dinb(n4182), .dout(n4191));
  jxor g4107(.dina(n4191), .dinb(n4141), .dout(n4192));
  jxor g4108(.dina(n4192), .dinb(n4135), .dout(n4193));
  jxor g4109(.dina(n4193), .dinb(n4132), .dout(n4194));
  jand g4110(.dina(n3669), .dinb(n466), .dout(n4195));
  jand g4111(.dina(n4195), .dinb(n881), .dout(n4196));
  jand g4112(.dina(n2429), .dinb(n2305), .dout(n4197));
  jand g4113(.dina(n4197), .dinb(n280), .dout(n4198));
  jand g4114(.dina(n925), .dinb(n918), .dout(n4199));
  jand g4115(.dina(n632), .dinb(n488), .dout(n4200));
  jand g4116(.dina(n4200), .dinb(n4199), .dout(n4201));
  jand g4117(.dina(n4201), .dinb(n565), .dout(n4202));
  jand g4118(.dina(n4202), .dinb(n4198), .dout(n4203));
  jand g4119(.dina(n4203), .dinb(n2365), .dout(n4204));
  jand g4120(.dina(n4204), .dinb(n4196), .dout(n4205));
  jand g4121(.dina(n4205), .dinb(n3155), .dout(n4206));
  jxor g4122(.dina(n4206), .dinb(n4194), .dout(n4207));
  jxor g4123(.dina(n4207), .dinb(n4129), .dout(n4208));
  jxor g4124(.dina(n4208), .dinb(n4125), .dout(n4209));
  jxor g4125(.dina(n4209), .dinb(n4124), .dout(sin3 ));
  jand g4126(.dina(n4208), .dinb(n4125), .dout(n4211));
  jnot g4127(.din(n4194), .dout(n4212));
  jor  g4128(.dina(n4206), .dinb(n4212), .dout(n4213));
  jor  g4129(.dina(n4207), .dinb(n4129), .dout(n4214));
  jand g4130(.dina(n4214), .dinb(n4213), .dout(n4215));
  jand g4131(.dina(n4192), .dinb(n4135), .dout(n4216));
  jand g4132(.dina(n4193), .dinb(n4132), .dout(n4217));
  jor  g4133(.dina(n4217), .dinb(n4216), .dout(n4218));
  jand g4134(.dina(n4190), .dinb(n4182), .dout(n4219));
  jand g4135(.dina(n4191), .dinb(n4141), .dout(n4220));
  jor  g4136(.dina(n4220), .dinb(n4219), .dout(n4221));
  jand g4137(.dina(n4180), .dinb(n4153), .dout(n4222));
  jand g4138(.dina(n4181), .dinb(n4144), .dout(n4223));
  jor  g4139(.dina(n4223), .dinb(n4222), .dout(n4224));
  jor  g4140(.dina(n3320), .dinb(n2795), .dout(n4225));
  jor  g4141(.dina(n3315), .dinb(n2800), .dout(n4226));
  jor  g4142(.dina(n3283), .dinb(n2805), .dout(n4227));
  jor  g4143(.dina(n3284), .dinb(n2809), .dout(n4228));
  jand g4144(.dina(n4228), .dinb(n4227), .dout(n4229));
  jand g4145(.dina(n4229), .dinb(n4226), .dout(n4230));
  jand g4146(.dina(n4230), .dinb(n4225), .dout(n4231));
  jxor g4147(.dina(n4231), .dinb(n699), .dout(n4232));
  jnot g4148(.din(n4232), .dout(n4233));
  jand g4149(.dina(n4178), .dinb(n4164), .dout(n4234));
  jand g4150(.dina(n4179), .dinb(n4156), .dout(n4235));
  jor  g4151(.dina(n4235), .dinb(n4234), .dout(n4236));
  jor  g4152(.dina(n3028), .dinb(n3198), .dout(n4237));
  jor  g4153(.dina(n3200), .dinb(n2671), .dout(n4238));
  jor  g4154(.dina(n3204), .dinb(n2674), .dout(n4239));
  jor  g4155(.dina(n3202), .dinb(n2678), .dout(n4240));
  jand g4156(.dina(n4240), .dinb(n4239), .dout(n4241));
  jand g4157(.dina(n4241), .dinb(n4238), .dout(n4242));
  jand g4158(.dina(n4242), .dinb(n4237), .dout(n4243));
  jxor g4159(.dina(n4243), .dinb(n954), .dout(n4244));
  jnot g4160(.din(n4244), .dout(n4245));
  jand g4161(.dina(n2684), .dinb(n954), .dout(n4246));
  jxor g4162(.dina(n4246), .dinb(n68), .dout(n4247));
  jxor g4163(.dina(n4247), .dinb(n4245), .dout(n4248));
  jand g4164(.dina(n4177), .dinb(n4173), .dout(n4249));
  jnot g4165(.din(n4172), .dout(n4250));
  jand g4166(.dina(n2685), .dinb(n954), .dout(n4251));
  jand g4167(.dina(n4251), .dinb(n4250), .dout(n4252));
  jor  g4168(.dina(n4252), .dinb(n4249), .dout(n4253));
  jxor g4169(.dina(n4253), .dinb(n4248), .dout(n4254));
  jand g4170(.dina(n3174), .dinb(n2828), .dout(n4255));
  jand g4171(.dina(n3176), .dinb(n2834), .dout(n4256));
  jand g4172(.dina(n2848), .dinb(n2670), .dout(n4257));
  jand g4173(.dina(n2832), .dinb(n2769), .dout(n4258));
  jor  g4174(.dina(n4258), .dinb(n4257), .dout(n4259));
  jor  g4175(.dina(n4259), .dinb(n4256), .dout(n4260));
  jor  g4176(.dina(n4260), .dinb(n4255), .dout(n4261));
  jxor g4177(.dina(n4261), .dinb(n803), .dout(n4262));
  jxor g4178(.dina(n4262), .dinb(n4254), .dout(n4263));
  jxor g4179(.dina(n4263), .dinb(n4236), .dout(n4264));
  jxor g4180(.dina(n4264), .dinb(n4233), .dout(n4265));
  jxor g4181(.dina(n4265), .dinb(n4224), .dout(n4266));
  jor  g4182(.dina(n3927), .dinb(n79), .dout(n4267));
  jor  g4183(.dina(n3919), .dinb(n2775), .dout(n4268));
  jor  g4184(.dina(n3806), .dinb(n2780), .dout(n4269));
  jor  g4185(.dina(n3600), .dinb(n2784), .dout(n4270));
  jand g4186(.dina(n4270), .dinb(n4269), .dout(n4271));
  jand g4187(.dina(n4271), .dinb(n4268), .dout(n4272));
  jand g4188(.dina(n4272), .dinb(n4267), .dout(n4273));
  jxor g4189(.dina(n4273), .dinb(n56), .dout(n4274));
  jxor g4190(.dina(n4274), .dinb(n4266), .dout(n4275));
  jxor g4191(.dina(n4275), .dinb(n4221), .dout(n4276));
  jxor g4192(.dina(n4276), .dinb(n4218), .dout(n4277));
  jand g4193(.dina(n2511), .dinb(n595), .dout(n4278));
  jand g4194(.dina(n4278), .dinb(n924), .dout(n4279));
  jand g4195(.dina(n535), .dinb(n323), .dout(n4280));
  jand g4196(.dina(n4280), .dinb(n2734), .dout(n4281));
  jand g4197(.dina(n4281), .dinb(n1026), .dout(n4282));
  jand g4198(.dina(n4282), .dinb(n4279), .dout(n4283));
  jand g4199(.dina(n4283), .dinb(n685), .dout(n4284));
  jand g4200(.dina(n4284), .dinb(n2551), .dout(n4285));
  jand g4201(.dina(n4285), .dinb(n395), .dout(n4286));
  jxor g4202(.dina(n4286), .dinb(n4277), .dout(n4287));
  jxor g4203(.dina(n4287), .dinb(n4215), .dout(n4288));
  jxor g4204(.dina(n4288), .dinb(n4211), .dout(n4289));
  jor  g4205(.dina(n4209), .dinb(n4123), .dout(n4290));
  jand g4206(.dina(n4290), .dinb(n4013), .dout(n4291));
  jxor g4207(.dina(n4291), .dinb(n4289), .dout(sin4 ));
  jand g4208(.dina(n4288), .dinb(n4211), .dout(n4293));
  jnot g4209(.din(n4277), .dout(n4294));
  jor  g4210(.dina(n4286), .dinb(n4294), .dout(n4295));
  jor  g4211(.dina(n4287), .dinb(n4215), .dout(n4296));
  jand g4212(.dina(n4296), .dinb(n4295), .dout(n4297));
  jand g4213(.dina(n4275), .dinb(n4221), .dout(n4298));
  jand g4214(.dina(n4276), .dinb(n4218), .dout(n4299));
  jor  g4215(.dina(n4299), .dinb(n4298), .dout(n4300));
  jand g4216(.dina(n4265), .dinb(n4224), .dout(n4301));
  jand g4217(.dina(n4274), .dinb(n4266), .dout(n4302));
  jor  g4218(.dina(n4302), .dinb(n4301), .dout(n4303));
  jand g4219(.dina(n4090), .dinb(n78), .dout(n4304));
  jand g4220(.dina(n3807), .dinb(n2783), .dout(n4305));
  jand g4221(.dina(n3920), .dinb(n2779), .dout(n4306));
  jor  g4222(.dina(n4306), .dinb(n4305), .dout(n4307));
  jor  g4223(.dina(n4307), .dinb(n4304), .dout(n4308));
  jxor g4224(.dina(n4308), .dinb(n55), .dout(n4309));
  jand g4225(.dina(n4263), .dinb(n4236), .dout(n4310));
  jand g4226(.dina(n4264), .dinb(n4233), .dout(n4311));
  jor  g4227(.dina(n4311), .dinb(n4310), .dout(n4312));
  jor  g4228(.dina(n3605), .dinb(n2795), .dout(n4313));
  jor  g4229(.dina(n3600), .dinb(n2800), .dout(n4314));
  jor  g4230(.dina(n3315), .dinb(n2805), .dout(n4315));
  jor  g4231(.dina(n3283), .dinb(n2809), .dout(n4316));
  jand g4232(.dina(n4316), .dinb(n4315), .dout(n4317));
  jand g4233(.dina(n4317), .dinb(n4314), .dout(n4318));
  jand g4234(.dina(n4318), .dinb(n4313), .dout(n4319));
  jxor g4235(.dina(n4319), .dinb(n699), .dout(n4320));
  jnot g4236(.din(n4320), .dout(n4321));
  jand g4237(.dina(n4253), .dinb(n4248), .dout(n4322));
  jand g4238(.dina(n4262), .dinb(n4254), .dout(n4323));
  jor  g4239(.dina(n4323), .dinb(n4322), .dout(n4324));
  jor  g4240(.dina(n3516), .dinb(n2857), .dout(n4325));
  jor  g4241(.dina(n3284), .dinb(n2860), .dout(n4326));
  jor  g4242(.dina(n3172), .dinb(n2865), .dout(n4327));
  jor  g4243(.dina(n2863), .dinb(n2773), .dout(n4328));
  jand g4244(.dina(n4328), .dinb(n4327), .dout(n4329));
  jand g4245(.dina(n4329), .dinb(n4326), .dout(n4330));
  jand g4246(.dina(n4330), .dinb(n4325), .dout(n4331));
  jxor g4247(.dina(n4331), .dinb(n808), .dout(n4332));
  jand g4248(.dina(n3016), .dinb(n2883), .dout(n4333));
  jand g4249(.dina(n2889), .dinb(n2670), .dout(n4334));
  jand g4250(.dina(n2995), .dinb(n2677), .dout(n4335));
  jand g4251(.dina(n2887), .dinb(n2672), .dout(n4336));
  jor  g4252(.dina(n4336), .dinb(n4335), .dout(n4337));
  jor  g4253(.dina(n4337), .dinb(n4334), .dout(n4338));
  jor  g4254(.dina(n4338), .dinb(n4333), .dout(n4339));
  jxor g4255(.dina(n4339), .dinb(n954), .dout(n4340));
  jand g4256(.dina(n4246), .dinb(n68), .dout(n4341));
  jand g4257(.dina(n4247), .dinb(n4245), .dout(n4342));
  jor  g4258(.dina(n4342), .dinb(n4341), .dout(n4343));
  jand g4259(.dina(n2679), .dinb(n954), .dout(n4344));
  jxor g4260(.dina(n4344), .dinb(n68), .dout(n4345));
  jxor g4261(.dina(n4345), .dinb(n4343), .dout(n4346));
  jxor g4262(.dina(n4346), .dinb(n4340), .dout(n4347));
  jxor g4263(.dina(n4347), .dinb(n4332), .dout(n4348));
  jxor g4264(.dina(n4348), .dinb(n4324), .dout(n4349));
  jxor g4265(.dina(n4349), .dinb(n4321), .dout(n4350));
  jxor g4266(.dina(n4350), .dinb(n4312), .dout(n4351));
  jxor g4267(.dina(n4351), .dinb(n4309), .dout(n4352));
  jxor g4268(.dina(n4352), .dinb(n4303), .dout(n4353));
  jxor g4269(.dina(n4353), .dinb(n4300), .dout(n4354));
  jand g4270(.dina(n2385), .dinb(n3634), .dout(n4355));
  jand g4271(.dina(n488), .dinb(n427), .dout(n4356));
  jand g4272(.dina(n4356), .dinb(n451), .dout(n4357));
  jand g4273(.dina(n4357), .dinb(n4355), .dout(n4358));
  jand g4274(.dina(n4358), .dinb(n4000), .dout(n4359));
  jand g4275(.dina(n849), .dinb(n216), .dout(n4360));
  jand g4276(.dina(n445), .dinb(n225), .dout(n4361));
  jand g4277(.dina(n4361), .dinb(n4360), .dout(n4362));
  jand g4278(.dina(n934), .dinb(n286), .dout(n4363));
  jand g4279(.dina(n4363), .dinb(n4362), .dout(n4364));
  jand g4280(.dina(n4364), .dinb(n2402), .dout(n4365));
  jand g4281(.dina(n4365), .dinb(n4359), .dout(n4366));
  jand g4282(.dina(n4366), .dinb(n3909), .dout(n4367));
  jand g4283(.dina(n4367), .dinb(n3256), .dout(n4368));
  jxor g4284(.dina(n4368), .dinb(n4354), .dout(n4369));
  jxor g4285(.dina(n4369), .dinb(n4297), .dout(n4370));
  jxor g4286(.dina(n4370), .dinb(n4293), .dout(n4371));
  jor  g4287(.dina(n4290), .dinb(n4289), .dout(n4372));
  jand g4288(.dina(n4372), .dinb(n4013), .dout(n4373));
  jxor g4289(.dina(n4373), .dinb(n4371), .dout(sin5 ));
  jand g4290(.dina(n4370), .dinb(n4293), .dout(n4375));
  jnot g4291(.din(n4354), .dout(n4376));
  jor  g4292(.dina(n4368), .dinb(n4376), .dout(n4377));
  jor  g4293(.dina(n4369), .dinb(n4297), .dout(n4378));
  jand g4294(.dina(n4378), .dinb(n4377), .dout(n4379));
  jand g4295(.dina(n4352), .dinb(n4303), .dout(n4380));
  jand g4296(.dina(n4353), .dinb(n4300), .dout(n4381));
  jor  g4297(.dina(n4381), .dinb(n4380), .dout(n4382));
  jand g4298(.dina(n4350), .dinb(n4312), .dout(n4383));
  jand g4299(.dina(n4351), .dinb(n4309), .dout(n4384));
  jor  g4300(.dina(n4384), .dinb(n4383), .dout(n4385));
  jand g4301(.dina(n4348), .dinb(n4324), .dout(n4386));
  jand g4302(.dina(n4349), .dinb(n4321), .dout(n4387));
  jor  g4303(.dina(n4387), .dinb(n4386), .dout(n4388));
  jnot g4304(.din(n4388), .dout(n4389));
  jor  g4305(.dina(n4136), .dinb(n79), .dout(n4390));
  jand g4306(.dina(n4390), .dinb(n2784), .dout(n4391));
  jor  g4307(.dina(n4391), .dinb(n3919), .dout(n4392));
  jxor g4308(.dina(n4392), .dinb(n55), .dout(n4393));
  jxor g4309(.dina(n4393), .dinb(n4389), .dout(n4394));
  jor  g4310(.dina(n3811), .dinb(n2795), .dout(n4395));
  jor  g4311(.dina(n3806), .dinb(n2800), .dout(n4396));
  jor  g4312(.dina(n3600), .dinb(n2805), .dout(n4397));
  jor  g4313(.dina(n3315), .dinb(n2809), .dout(n4398));
  jand g4314(.dina(n4398), .dinb(n4397), .dout(n4399));
  jand g4315(.dina(n4399), .dinb(n4396), .dout(n4400));
  jand g4316(.dina(n4400), .dinb(n4395), .dout(n4401));
  jxor g4317(.dina(n4401), .dinb(n699), .dout(n4402));
  jnot g4318(.din(n4402), .dout(n4403));
  jand g4319(.dina(n4346), .dinb(n4340), .dout(n4404));
  jand g4320(.dina(n4347), .dinb(n4332), .dout(n4405));
  jor  g4321(.dina(n4405), .dinb(n4404), .dout(n4406));
  jor  g4322(.dina(n3337), .dinb(n2857), .dout(n4407));
  jor  g4323(.dina(n3283), .dinb(n2860), .dout(n4408));
  jor  g4324(.dina(n3284), .dinb(n2865), .dout(n4409));
  jor  g4325(.dina(n3172), .dinb(n2863), .dout(n4410));
  jand g4326(.dina(n4410), .dinb(n4409), .dout(n4411));
  jand g4327(.dina(n4411), .dinb(n4408), .dout(n4412));
  jand g4328(.dina(n4412), .dinb(n4407), .dout(n4413));
  jxor g4329(.dina(n4413), .dinb(n808), .dout(n4414));
  jor  g4330(.dina(n3198), .dinb(n2771), .dout(n4415));
  jor  g4331(.dina(n3200), .dinb(n2773), .dout(n4416));
  jor  g4332(.dina(n3204), .dinb(n2669), .dout(n4417));
  jor  g4333(.dina(n3202), .dinb(n2671), .dout(n4418));
  jand g4334(.dina(n4418), .dinb(n4417), .dout(n4419));
  jand g4335(.dina(n4419), .dinb(n4416), .dout(n4420));
  jand g4336(.dina(n4420), .dinb(n4415), .dout(n4421));
  jxor g4337(.dina(n4421), .dinb(n820), .dout(n4422));
  jand g4338(.dina(n4344), .dinb(n68), .dout(n4423));
  jand g4339(.dina(n4345), .dinb(n4343), .dout(n4424));
  jor  g4340(.dina(n4424), .dinb(n4423), .dout(n4425));
  jand g4341(.dina(n2677), .dinb(n954), .dout(n4426));
  jxor g4342(.dina(n4426), .dinb(n68), .dout(n4427));
  jxor g4343(.dina(n4427), .dinb(n4425), .dout(n4428));
  jxor g4344(.dina(n4428), .dinb(n4422), .dout(n4429));
  jxor g4345(.dina(n4429), .dinb(n4414), .dout(n4430));
  jxor g4346(.dina(n4430), .dinb(n4406), .dout(n4431));
  jxor g4347(.dina(n4431), .dinb(n4403), .dout(n4432));
  jxor g4348(.dina(n4432), .dinb(n4394), .dout(n4433));
  jxor g4349(.dina(n4433), .dinb(n4385), .dout(n4434));
  jxor g4350(.dina(n4434), .dinb(n4382), .dout(n4435));
  jand g4351(.dina(n2429), .dinb(n763), .dout(n4436));
  jand g4352(.dina(n4436), .dinb(n3911), .dout(n4437));
  jand g4353(.dina(n4437), .dinb(n2541), .dout(n4438));
  jand g4354(.dina(n865), .dinb(n822), .dout(n4439));
  jand g4355(.dina(n4439), .dinb(n2385), .dout(n4440));
  jand g4356(.dina(n4440), .dinb(n2514), .dout(n4441));
  jand g4357(.dina(n4441), .dinb(n4438), .dout(n4442));
  jand g4358(.dina(n401), .dinb(n379), .dout(n4443));
  jand g4359(.dina(n4443), .dinb(n680), .dout(n4444));
  jand g4360(.dina(n3307), .dinb(n1294), .dout(n4445));
  jand g4361(.dina(n4445), .dinb(n2387), .dout(n4446));
  jand g4362(.dina(n4446), .dinb(n4444), .dout(n4447));
  jand g4363(.dina(n4447), .dinb(n2540), .dout(n4448));
  jand g4364(.dina(n4448), .dinb(n4442), .dout(n4449));
  jand g4365(.dina(n4449), .dinb(n3633), .dout(n4450));
  jxor g4366(.dina(n4450), .dinb(n4435), .dout(n4451));
  jxor g4367(.dina(n4451), .dinb(n4379), .dout(n4452));
  jxor g4368(.dina(n4452), .dinb(n4375), .dout(n4453));
  jor  g4369(.dina(n4372), .dinb(n4371), .dout(n4454));
  jand g4370(.dina(n4454), .dinb(n4013), .dout(n4455));
  jxor g4371(.dina(n4455), .dinb(n4453), .dout(sin6 ));
  jand g4372(.dina(n4452), .dinb(n4375), .dout(n4457));
  jnot g4373(.din(n4435), .dout(n4458));
  jor  g4374(.dina(n4450), .dinb(n4458), .dout(n4459));
  jor  g4375(.dina(n4451), .dinb(n4379), .dout(n4460));
  jand g4376(.dina(n4460), .dinb(n4459), .dout(n4461));
  jand g4377(.dina(n4433), .dinb(n4385), .dout(n4462));
  jand g4378(.dina(n4434), .dinb(n4382), .dout(n4463));
  jor  g4379(.dina(n4463), .dinb(n4462), .dout(n4464));
  jor  g4380(.dina(n4393), .dinb(n4389), .dout(n4465));
  jand g4381(.dina(n4432), .dinb(n4394), .dout(n4466));
  jnot g4382(.din(n4466), .dout(n4467));
  jand g4383(.dina(n4467), .dinb(n4465), .dout(n4468));
  jnot g4384(.din(n4468), .dout(n4469));
  jand g4385(.dina(n4430), .dinb(n4406), .dout(n4470));
  jand g4386(.dina(n4431), .dinb(n4403), .dout(n4471));
  jor  g4387(.dina(n4471), .dinb(n4470), .dout(n4472));
  jor  g4388(.dina(n3927), .dinb(n2795), .dout(n4473));
  jor  g4389(.dina(n3919), .dinb(n2800), .dout(n4474));
  jor  g4390(.dina(n3806), .dinb(n2805), .dout(n4475));
  jor  g4391(.dina(n3600), .dinb(n2809), .dout(n4476));
  jand g4392(.dina(n4476), .dinb(n4475), .dout(n4477));
  jand g4393(.dina(n4477), .dinb(n4474), .dout(n4478));
  jand g4394(.dina(n4478), .dinb(n4473), .dout(n4479));
  jxor g4395(.dina(n4479), .dinb(n1143), .dout(n4480));
  jxor g4396(.dina(n4480), .dinb(n4472), .dout(n4481));
  jand g4397(.dina(n4428), .dinb(n4422), .dout(n4482));
  jand g4398(.dina(n4429), .dinb(n4414), .dout(n4483));
  jor  g4399(.dina(n4483), .dinb(n4482), .dout(n4484));
  jand g4400(.dina(n4426), .dinb(n68), .dout(n4485));
  jand g4401(.dina(n4427), .dinb(n4425), .dout(n4486));
  jor  g4402(.dina(n4486), .dinb(n4485), .dout(n4487));
  jand g4403(.dina(n3174), .dinb(n2883), .dout(n4488));
  jand g4404(.dina(n3176), .dinb(n2889), .dout(n4489));
  jand g4405(.dina(n2995), .dinb(n2670), .dout(n4490));
  jand g4406(.dina(n2887), .dinb(n2769), .dout(n4491));
  jor  g4407(.dina(n4491), .dinb(n4490), .dout(n4492));
  jor  g4408(.dina(n4492), .dinb(n4489), .dout(n4493));
  jor  g4409(.dina(n4493), .dinb(n4488), .dout(n4494));
  jxor g4410(.dina(n4494), .dinb(n820), .dout(n4495));
  jnot g4411(.din(n4495), .dout(n4496));
  jand g4412(.dina(n2672), .dinb(n954), .dout(n4497));
  jxor g4413(.dina(n68), .dinb(n55), .dout(n4498));
  jxor g4414(.dina(n4498), .dinb(n4497), .dout(n4499));
  jxor g4415(.dina(n4499), .dinb(n4496), .dout(n4500));
  jxor g4416(.dina(n4500), .dinb(n4487), .dout(n4501));
  jor  g4417(.dina(n3320), .dinb(n2857), .dout(n4502));
  jor  g4418(.dina(n3315), .dinb(n2860), .dout(n4503));
  jor  g4419(.dina(n3283), .dinb(n2865), .dout(n4504));
  jor  g4420(.dina(n3284), .dinb(n2863), .dout(n4505));
  jand g4421(.dina(n4505), .dinb(n4504), .dout(n4506));
  jand g4422(.dina(n4506), .dinb(n4503), .dout(n4507));
  jand g4423(.dina(n4507), .dinb(n4502), .dout(n4508));
  jxor g4424(.dina(n4508), .dinb(n808), .dout(n4509));
  jxor g4425(.dina(n4509), .dinb(n4501), .dout(n4510));
  jxor g4426(.dina(n4510), .dinb(n4484), .dout(n4511));
  jxor g4427(.dina(n4511), .dinb(n4481), .dout(n4512));
  jxor g4428(.dina(n4512), .dinb(n4469), .dout(n4513));
  jxor g4429(.dina(n4513), .dinb(n4464), .dout(n4514));
  jand g4430(.dina(n1188), .dinb(n471), .dout(n4515));
  jand g4431(.dina(n2406), .dinb(n1170), .dout(n4516));
  jand g4432(.dina(n4516), .dinb(n4515), .dout(n4517));
  jand g4433(.dina(n270), .dinb(n214), .dout(n4518));
  jand g4434(.dina(n4518), .dinb(n930), .dout(n4519));
  jand g4435(.dina(n4519), .dinb(n4357), .dout(n4520));
  jand g4436(.dina(n4520), .dinb(n4517), .dout(n4521));
  jand g4437(.dina(n4521), .dinb(n4442), .dout(n4522));
  jand g4438(.dina(n4522), .dinb(n2350), .dout(n4523));
  jxor g4439(.dina(n4523), .dinb(n4514), .dout(n4524));
  jxor g4440(.dina(n4524), .dinb(n4461), .dout(n4525));
  jxor g4441(.dina(n4525), .dinb(n4457), .dout(n4526));
  jor  g4442(.dina(n4454), .dinb(n4453), .dout(n4527));
  jand g4443(.dina(n4527), .dinb(n4013), .dout(n4528));
  jxor g4444(.dina(n4528), .dinb(n4526), .dout(sin7 ));
  jand g4445(.dina(n4525), .dinb(n4457), .dout(n4530));
  jnot g4446(.din(n4514), .dout(n4531));
  jor  g4447(.dina(n4523), .dinb(n4531), .dout(n4532));
  jor  g4448(.dina(n4524), .dinb(n4461), .dout(n4533));
  jand g4449(.dina(n4533), .dinb(n4532), .dout(n4534));
  jand g4450(.dina(n4512), .dinb(n4469), .dout(n4535));
  jand g4451(.dina(n4513), .dinb(n4464), .dout(n4536));
  jor  g4452(.dina(n4536), .dinb(n4535), .dout(n4537));
  jand g4453(.dina(n4480), .dinb(n4472), .dout(n4538));
  jand g4454(.dina(n4511), .dinb(n4481), .dout(n4539));
  jor  g4455(.dina(n4539), .dinb(n4538), .dout(n4540));
  jand g4456(.dina(n4090), .dinb(n2794), .dout(n4541));
  jand g4457(.dina(n3807), .dinb(n2808), .dout(n4542));
  jand g4458(.dina(n3920), .dinb(n2804), .dout(n4543));
  jor  g4459(.dina(n4543), .dinb(n4542), .dout(n4544));
  jor  g4460(.dina(n4544), .dinb(n4541), .dout(n4545));
  jxor g4461(.dina(n4545), .dinb(n1143), .dout(n4546));
  jnot g4462(.din(n4546), .dout(n4547));
  jand g4463(.dina(n4509), .dinb(n4501), .dout(n4548));
  jand g4464(.dina(n4510), .dinb(n4484), .dout(n4549));
  jor  g4465(.dina(n4549), .dinb(n4548), .dout(n4550));
  jor  g4466(.dina(n3605), .dinb(n2857), .dout(n4551));
  jor  g4467(.dina(n3600), .dinb(n2860), .dout(n4552));
  jor  g4468(.dina(n3315), .dinb(n2865), .dout(n4553));
  jor  g4469(.dina(n3283), .dinb(n2863), .dout(n4554));
  jand g4470(.dina(n4554), .dinb(n4553), .dout(n4555));
  jand g4471(.dina(n4555), .dinb(n4552), .dout(n4556));
  jand g4472(.dina(n4556), .dinb(n4551), .dout(n4557));
  jxor g4473(.dina(n4557), .dinb(n808), .dout(n4558));
  jand g4474(.dina(n4499), .dinb(n4496), .dout(n4559));
  jand g4475(.dina(n4500), .dinb(n4487), .dout(n4560));
  jor  g4476(.dina(n4560), .dinb(n4559), .dout(n4561));
  jor  g4477(.dina(n3516), .dinb(n3198), .dout(n4562));
  jor  g4478(.dina(n3284), .dinb(n3200), .dout(n4563));
  jor  g4479(.dina(n3172), .dinb(n3204), .dout(n4564));
  jor  g4480(.dina(n3202), .dinb(n2773), .dout(n4565));
  jand g4481(.dina(n4565), .dinb(n4564), .dout(n4566));
  jand g4482(.dina(n4566), .dinb(n4563), .dout(n4567));
  jand g4483(.dina(n4567), .dinb(n4562), .dout(n4568));
  jxor g4484(.dina(n4568), .dinb(n820), .dout(n4569));
  jand g4485(.dina(n2670), .dinb(n954), .dout(n4570));
  jnot g4486(.din(n4570), .dout(n4571));
  jand g4487(.dina(n3233), .dinb(n56), .dout(n4572));
  jand g4488(.dina(n4498), .dinb(n4497), .dout(n4573));
  jor  g4489(.dina(n4573), .dinb(n4572), .dout(n4574));
  jxor g4490(.dina(n4574), .dinb(n4571), .dout(n4575));
  jxor g4491(.dina(n4575), .dinb(n4569), .dout(n4576));
  jxor g4492(.dina(n4576), .dinb(n4561), .dout(n4577));
  jxor g4493(.dina(n4577), .dinb(n4558), .dout(n4578));
  jxor g4494(.dina(n4578), .dinb(n4550), .dout(n4579));
  jxor g4495(.dina(n4579), .dinb(n4547), .dout(n4580));
  jxor g4496(.dina(n4580), .dinb(n4540), .dout(n4581));
  jxor g4497(.dina(n4581), .dinb(n4537), .dout(n4582));
  jand g4498(.dina(n421), .dinb(n147), .dout(n4583));
  jand g4499(.dina(n4583), .dinb(n295), .dout(n4584));
  jand g4500(.dina(n735), .dinb(n638), .dout(n4585));
  jand g4501(.dina(n4585), .dinb(n3626), .dout(n4586));
  jand g4502(.dina(n4586), .dinb(n4584), .dout(n4587));
  jand g4503(.dina(n4587), .dinb(n2571), .dout(n4588));
  jand g4504(.dina(n4588), .dinb(n832), .dout(n4589));
  jand g4505(.dina(n277), .dinb(n229), .dout(n4590));
  jand g4506(.dina(n4590), .dinb(n410), .dout(n4591));
  jand g4507(.dina(n765), .dinb(n751), .dout(n4592));
  jand g4508(.dina(n4592), .dinb(n2424), .dout(n4593));
  jand g4509(.dina(n4593), .dinb(n4591), .dout(n4594));
  jand g4510(.dina(n2428), .dinb(n667), .dout(n4595));
  jand g4511(.dina(n4595), .dinb(n4594), .dout(n4596));
  jand g4512(.dina(n4596), .dinb(n655), .dout(n4597));
  jand g4513(.dina(n4597), .dinb(n4589), .dout(n4598));
  jand g4514(.dina(n4598), .dinb(n3666), .dout(n4599));
  jxor g4515(.dina(n4599), .dinb(n4582), .dout(n4600));
  jxor g4516(.dina(n4600), .dinb(n4534), .dout(n4601));
  jxor g4517(.dina(n4601), .dinb(n4530), .dout(n4602));
  jor  g4518(.dina(n4527), .dinb(n4526), .dout(n4603));
  jand g4519(.dina(n4603), .dinb(n4013), .dout(n4604));
  jxor g4520(.dina(n4604), .dinb(n4602), .dout(sin8 ));
  jand g4521(.dina(n4601), .dinb(n4530), .dout(n4606));
  jnot g4522(.din(n4582), .dout(n4607));
  jor  g4523(.dina(n4599), .dinb(n4607), .dout(n4608));
  jor  g4524(.dina(n4600), .dinb(n4534), .dout(n4609));
  jand g4525(.dina(n4609), .dinb(n4608), .dout(n4610));
  jand g4526(.dina(n4580), .dinb(n4540), .dout(n4611));
  jand g4527(.dina(n4581), .dinb(n4537), .dout(n4612));
  jor  g4528(.dina(n4612), .dinb(n4611), .dout(n4613));
  jand g4529(.dina(n4578), .dinb(n4550), .dout(n4614));
  jand g4530(.dina(n4579), .dinb(n4547), .dout(n4615));
  jor  g4531(.dina(n4615), .dinb(n4614), .dout(n4616));
  jand g4532(.dina(n4576), .dinb(n4561), .dout(n4617));
  jand g4533(.dina(n4577), .dinb(n4558), .dout(n4618));
  jor  g4534(.dina(n4618), .dinb(n4617), .dout(n4619));
  jnot g4535(.din(n4619), .dout(n4620));
  jor  g4536(.dina(n4136), .dinb(n2795), .dout(n4621));
  jand g4537(.dina(n4621), .dinb(n2809), .dout(n4622));
  jor  g4538(.dina(n4622), .dinb(n3919), .dout(n4623));
  jxor g4539(.dina(n4623), .dinb(n699), .dout(n4624));
  jxor g4540(.dina(n4624), .dinb(n4620), .dout(n4625));
  jand g4541(.dina(n4574), .dinb(n4571), .dout(n4626));
  jand g4542(.dina(n4575), .dinb(n4569), .dout(n4627));
  jor  g4543(.dina(n4627), .dinb(n4626), .dout(n4628));
  jor  g4544(.dina(n3337), .dinb(n3198), .dout(n4629));
  jor  g4545(.dina(n3283), .dinb(n3200), .dout(n4630));
  jor  g4546(.dina(n3284), .dinb(n3204), .dout(n4631));
  jor  g4547(.dina(n3172), .dinb(n3202), .dout(n4632));
  jand g4548(.dina(n4632), .dinb(n4631), .dout(n4633));
  jand g4549(.dina(n4633), .dinb(n4630), .dout(n4634));
  jand g4550(.dina(n4634), .dinb(n4629), .dout(n4635));
  jxor g4551(.dina(n4635), .dinb(n954), .dout(n4636));
  jand g4552(.dina(n2770), .dinb(n954), .dout(n4637));
  jxor g4553(.dina(n4637), .dinb(n4636), .dout(n4638));
  jxor g4554(.dina(n4638), .dinb(n4628), .dout(n4639));
  jor  g4555(.dina(n3811), .dinb(n2857), .dout(n4640));
  jor  g4556(.dina(n3806), .dinb(n2860), .dout(n4641));
  jor  g4557(.dina(n3600), .dinb(n2865), .dout(n4642));
  jor  g4558(.dina(n3315), .dinb(n2863), .dout(n4643));
  jand g4559(.dina(n4643), .dinb(n4642), .dout(n4644));
  jand g4560(.dina(n4644), .dinb(n4641), .dout(n4645));
  jand g4561(.dina(n4645), .dinb(n4640), .dout(n4646));
  jxor g4562(.dina(n4646), .dinb(n808), .dout(n4647));
  jxor g4563(.dina(n4647), .dinb(n4639), .dout(n4648));
  jxor g4564(.dina(n4648), .dinb(n4625), .dout(n4649));
  jxor g4565(.dina(n4649), .dinb(n4616), .dout(n4650));
  jxor g4566(.dina(n4650), .dinb(n4613), .dout(n4651));
  jand g4567(.dina(n668), .dinb(n279), .dout(n4652));
  jand g4568(.dina(n645), .dinb(n147), .dout(n4653));
  jand g4569(.dina(n4653), .dinb(n4652), .dout(n4654));
  jand g4570(.dina(n3307), .dinb(n930), .dout(n4655));
  jand g4571(.dina(n4655), .dinb(n4654), .dout(n4656));
  jand g4572(.dina(n579), .dinb(n390), .dout(n4657));
  jand g4573(.dina(n4657), .dinb(n303), .dout(n4658));
  jand g4574(.dina(n4658), .dinb(n3242), .dout(n4659));
  jand g4575(.dina(n4659), .dinb(n4656), .dout(n4660));
  jand g4576(.dina(n4660), .dinb(n405), .dout(n4661));
  jand g4577(.dina(n4661), .dinb(n3638), .dout(n4662));
  jand g4578(.dina(n4662), .dinb(n2520), .dout(n4663));
  jxor g4579(.dina(n4663), .dinb(n4651), .dout(n4664));
  jxor g4580(.dina(n4664), .dinb(n4610), .dout(n4665));
  jxor g4581(.dina(n4665), .dinb(n4606), .dout(n4666));
  jor  g4582(.dina(n4603), .dinb(n4602), .dout(n4667));
  jand g4583(.dina(n4667), .dinb(n4013), .dout(n4668));
  jxor g4584(.dina(n4668), .dinb(n4666), .dout(sin9 ));
  jand g4585(.dina(n4665), .dinb(n4606), .dout(n4670));
  jnot g4586(.din(n4651), .dout(n4671));
  jor  g4587(.dina(n4663), .dinb(n4671), .dout(n4672));
  jor  g4588(.dina(n4664), .dinb(n4610), .dout(n4673));
  jand g4589(.dina(n4673), .dinb(n4672), .dout(n4674));
  jand g4590(.dina(n4649), .dinb(n4616), .dout(n4675));
  jand g4591(.dina(n4650), .dinb(n4613), .dout(n4676));
  jor  g4592(.dina(n4676), .dinb(n4675), .dout(n4677));
  jor  g4593(.dina(n4624), .dinb(n4620), .dout(n4678));
  jand g4594(.dina(n4648), .dinb(n4625), .dout(n4679));
  jnot g4595(.din(n4679), .dout(n4680));
  jand g4596(.dina(n4680), .dinb(n4678), .dout(n4681));
  jnot g4597(.din(n4681), .dout(n4682));
  jand g4598(.dina(n4638), .dinb(n4628), .dout(n4683));
  jand g4599(.dina(n4647), .dinb(n4639), .dout(n4684));
  jor  g4600(.dina(n4684), .dinb(n4683), .dout(n4685));
  jor  g4601(.dina(n3927), .dinb(n2857), .dout(n4686));
  jor  g4602(.dina(n3919), .dinb(n2860), .dout(n4687));
  jor  g4603(.dina(n3806), .dinb(n2865), .dout(n4688));
  jor  g4604(.dina(n3600), .dinb(n2863), .dout(n4689));
  jand g4605(.dina(n4689), .dinb(n4688), .dout(n4690));
  jand g4606(.dina(n4690), .dinb(n4687), .dout(n4691));
  jand g4607(.dina(n4691), .dinb(n4686), .dout(n4692));
  jxor g4608(.dina(n4692), .dinb(n808), .dout(n4693));
  jxor g4609(.dina(n4693), .dinb(n4685), .dout(n4694));
  jor  g4610(.dina(n3320), .dinb(n3198), .dout(n4695));
  jor  g4611(.dina(n3315), .dinb(n3200), .dout(n4696));
  jor  g4612(.dina(n3283), .dinb(n3204), .dout(n4697));
  jor  g4613(.dina(n3284), .dinb(n3202), .dout(n4698));
  jand g4614(.dina(n4698), .dinb(n4697), .dout(n4699));
  jand g4615(.dina(n4699), .dinb(n4696), .dout(n4700));
  jand g4616(.dina(n4700), .dinb(n4695), .dout(n4701));
  jxor g4617(.dina(n4701), .dinb(n954), .dout(n4702));
  jnot g4618(.din(n4702), .dout(n4703));
  jand g4619(.dina(n3176), .dinb(n954), .dout(n4704));
  jxor g4620(.dina(n4704), .dinb(n1143), .dout(n4705));
  jxor g4621(.dina(n4705), .dinb(n4571), .dout(n4706));
  jor  g4622(.dina(n4637), .dinb(n4636), .dout(n4707));
  jand g4623(.dina(n2669), .dinb(n954), .dout(n4708));
  jand g4624(.dina(n4708), .dinb(n2769), .dout(n4709));
  jnot g4625(.din(n4709), .dout(n4710));
  jand g4626(.dina(n4710), .dinb(n4707), .dout(n4711));
  jxor g4627(.dina(n4711), .dinb(n4706), .dout(n4712));
  jxor g4628(.dina(n4712), .dinb(n4703), .dout(n4713));
  jxor g4629(.dina(n4713), .dinb(n4694), .dout(n4714));
  jxor g4630(.dina(n4714), .dinb(n4682), .dout(n4715));
  jxor g4631(.dina(n4715), .dinb(n4677), .dout(n4716));
  jand g4632(.dina(n3307), .dinb(n2736), .dout(n4717));
  jand g4633(.dina(n4717), .dinb(n771), .dout(n4718));
  jand g4634(.dina(n878), .dinb(n310), .dout(n4719));
  jand g4635(.dina(n4719), .dinb(n479), .dout(n4720));
  jand g4636(.dina(n4720), .dinb(n385), .dout(n4721));
  jnot g4637(.din(n651), .dout(n4722));
  jand g4638(.dina(n3258), .dinb(n4722), .dout(n4723));
  jand g4639(.dina(n4723), .dinb(n4721), .dout(n4724));
  jand g4640(.dina(n4724), .dinb(n4718), .dout(n4725));
  jand g4641(.dina(n4725), .dinb(n1203), .dout(n4726));
  jand g4642(.dina(n3676), .dinb(n1013), .dout(n4727));
  jand g4643(.dina(n4727), .dinb(n4726), .dout(n4728));
  jxor g4644(.dina(n4728), .dinb(n4716), .dout(n4729));
  jxor g4645(.dina(n4729), .dinb(n4674), .dout(n4730));
  jxor g4646(.dina(n4730), .dinb(n4670), .dout(n4731));
  jor  g4647(.dina(n4667), .dinb(n4666), .dout(n4732));
  jand g4648(.dina(n4732), .dinb(n4013), .dout(n4733));
  jxor g4649(.dina(n4733), .dinb(n4731), .dout(sin10 ));
  jand g4650(.dina(n4730), .dinb(n4670), .dout(n4735));
  jnot g4651(.din(n4716), .dout(n4736));
  jor  g4652(.dina(n4728), .dinb(n4736), .dout(n4737));
  jor  g4653(.dina(n4729), .dinb(n4674), .dout(n4738));
  jand g4654(.dina(n4738), .dinb(n4737), .dout(n4739));
  jand g4655(.dina(n4714), .dinb(n4682), .dout(n4740));
  jand g4656(.dina(n4715), .dinb(n4677), .dout(n4741));
  jor  g4657(.dina(n4741), .dinb(n4740), .dout(n4742));
  jand g4658(.dina(n4693), .dinb(n4685), .dout(n4743));
  jand g4659(.dina(n4713), .dinb(n4694), .dout(n4744));
  jor  g4660(.dina(n4744), .dinb(n4743), .dout(n4745));
  jand g4661(.dina(n4090), .dinb(n2828), .dout(n4746));
  jand g4662(.dina(n3807), .dinb(n2848), .dout(n4747));
  jand g4663(.dina(n3920), .dinb(n2832), .dout(n4748));
  jor  g4664(.dina(n4748), .dinb(n4747), .dout(n4749));
  jor  g4665(.dina(n4749), .dinb(n4746), .dout(n4750));
  jxor g4666(.dina(n4750), .dinb(n803), .dout(n4751));
  jor  g4667(.dina(n3605), .dinb(n3198), .dout(n4752));
  jor  g4668(.dina(n3600), .dinb(n3200), .dout(n4753));
  jor  g4669(.dina(n3315), .dinb(n3204), .dout(n4754));
  jor  g4670(.dina(n3283), .dinb(n3202), .dout(n4755));
  jand g4671(.dina(n4755), .dinb(n4754), .dout(n4756));
  jand g4672(.dina(n4756), .dinb(n4753), .dout(n4757));
  jand g4673(.dina(n4757), .dinb(n4752), .dout(n4758));
  jxor g4674(.dina(n4758), .dinb(n820), .dout(n4759));
  jor  g4675(.dina(n3284), .dinb(n820), .dout(n4760));
  jnot g4676(.din(n4704), .dout(n4761));
  jand g4677(.dina(n4761), .dinb(n699), .dout(n4762));
  jnot g4678(.din(n4762), .dout(n4763));
  jand g4679(.dina(n4704), .dinb(n1143), .dout(n4764));
  jor  g4680(.dina(n4764), .dinb(n4570), .dout(n4765));
  jand g4681(.dina(n4765), .dinb(n4763), .dout(n4766));
  jxor g4682(.dina(n4766), .dinb(n4760), .dout(n4767));
  jxor g4683(.dina(n4767), .dinb(n4759), .dout(n4768));
  jand g4684(.dina(n4711), .dinb(n4706), .dout(n4769));
  jnot g4685(.din(n4769), .dout(n4770));
  jnot g4686(.din(n4706), .dout(n4771));
  jnot g4687(.din(n4711), .dout(n4772));
  jand g4688(.dina(n4772), .dinb(n4771), .dout(n4773));
  jor  g4689(.dina(n4773), .dinb(n4703), .dout(n4774));
  jand g4690(.dina(n4774), .dinb(n4770), .dout(n4775));
  jxor g4691(.dina(n4775), .dinb(n4768), .dout(n4776));
  jxor g4692(.dina(n4776), .dinb(n4751), .dout(n4777));
  jxor g4693(.dina(n4777), .dinb(n4745), .dout(n4778));
  jxor g4694(.dina(n4778), .dinb(n4742), .dout(n4779));
  jand g4695(.dina(n935), .dinb(n511), .dout(n4780));
  jand g4696(.dina(n4780), .dinb(n677), .dout(n4781));
  jand g4697(.dina(n4781), .dinb(n746), .dout(n4782));
  jand g4698(.dina(n4782), .dinb(n784), .dout(n4783));
  jand g4699(.dina(n4783), .dinb(n3794), .dout(n4784));
  jand g4700(.dina(n4784), .dinb(n1006), .dout(n4785));
  jxor g4701(.dina(n4785), .dinb(n4779), .dout(n4786));
  jxor g4702(.dina(n4786), .dinb(n4739), .dout(n4787));
  jxor g4703(.dina(n4787), .dinb(n4735), .dout(n4788));
  jor  g4704(.dina(n4732), .dinb(n4731), .dout(n4789));
  jand g4705(.dina(n4789), .dinb(n4013), .dout(n4790));
  jxor g4706(.dina(n4790), .dinb(n4788), .dout(sin11 ));
  jand g4707(.dina(n4787), .dinb(n4735), .dout(n4792));
  jnot g4708(.din(n4779), .dout(n4793));
  jor  g4709(.dina(n4785), .dinb(n4793), .dout(n4794));
  jor  g4710(.dina(n4786), .dinb(n4739), .dout(n4795));
  jand g4711(.dina(n4795), .dinb(n4794), .dout(n4796));
  jand g4712(.dina(n4777), .dinb(n4745), .dout(n4797));
  jand g4713(.dina(n4778), .dinb(n4742), .dout(n4798));
  jor  g4714(.dina(n4798), .dinb(n4797), .dout(n4799));
  jand g4715(.dina(n4775), .dinb(n4768), .dout(n4800));
  jand g4716(.dina(n4776), .dinb(n4751), .dout(n4801));
  jor  g4717(.dina(n4801), .dinb(n4800), .dout(n4802));
  jand g4718(.dina(n4766), .dinb(n4760), .dout(n4803));
  jand g4719(.dina(n4767), .dinb(n4759), .dout(n4804));
  jor  g4720(.dina(n4804), .dinb(n4803), .dout(n4805));
  jnot g4721(.din(n4805), .dout(n4806));
  jand g4722(.dina(n3299), .dinb(n954), .dout(n4807));
  jxor g4723(.dina(n4807), .dinb(n4806), .dout(n4808));
  jor  g4724(.dina(n3811), .dinb(n3198), .dout(n4809));
  jor  g4725(.dina(n3806), .dinb(n3200), .dout(n4810));
  jor  g4726(.dina(n3600), .dinb(n3204), .dout(n4811));
  jor  g4727(.dina(n3315), .dinb(n3202), .dout(n4812));
  jand g4728(.dina(n4812), .dinb(n4811), .dout(n4813));
  jand g4729(.dina(n4813), .dinb(n4810), .dout(n4814));
  jand g4730(.dina(n4814), .dinb(n4809), .dout(n4815));
  jxor g4731(.dina(n4815), .dinb(n954), .dout(n4816));
  jor  g4732(.dina(n4136), .dinb(n2857), .dout(n4817));
  jand g4733(.dina(n4817), .dinb(n2863), .dout(n4818));
  jor  g4734(.dina(n4818), .dinb(n3919), .dout(n4819));
  jxor g4735(.dina(n4819), .dinb(n803), .dout(n4820));
  jxor g4736(.dina(n4820), .dinb(n4816), .dout(n4821));
  jxor g4737(.dina(n4821), .dinb(n4808), .dout(n4822));
  jxor g4738(.dina(n4822), .dinb(n4802), .dout(n4823));
  jxor g4739(.dina(n4823), .dinb(n4799), .dout(n4824));
  jand g4740(.dina(n421), .dinb(n254), .dout(n4825));
  jand g4741(.dina(n4825), .dinb(n372), .dout(n4826));
  jand g4742(.dina(n4826), .dinb(n2456), .dout(n4827));
  jand g4743(.dina(n4827), .dinb(n565), .dout(n4828));
  jand g4744(.dina(n668), .dinb(n420), .dout(n4829));
  jand g4745(.dina(n594), .dinb(n868), .dout(n4830));
  jand g4746(.dina(n4830), .dinb(n277), .dout(n4831));
  jand g4747(.dina(n4831), .dinb(n4829), .dout(n4832));
  jand g4748(.dina(n4832), .dinb(n4106), .dout(n4833));
  jand g4749(.dina(n4833), .dinb(n4828), .dout(n4834));
  jand g4750(.dina(n4834), .dinb(n2449), .dout(n4835));
  jand g4751(.dina(n4835), .dinb(n2313), .dout(n4836));
  jxor g4752(.dina(n4836), .dinb(n4824), .dout(n4837));
  jxor g4753(.dina(n4837), .dinb(n4796), .dout(n4838));
  jxor g4754(.dina(n4838), .dinb(n4792), .dout(n4839));
  jor  g4755(.dina(n4789), .dinb(n4788), .dout(n4840));
  jand g4756(.dina(n4840), .dinb(n4013), .dout(n4841));
  jxor g4757(.dina(n4841), .dinb(n4839), .dout(sin12 ));
  jand g4758(.dina(n4838), .dinb(n4792), .dout(n4843));
  jnot g4759(.din(n4824), .dout(n4844));
  jor  g4760(.dina(n4836), .dinb(n4844), .dout(n4845));
  jor  g4761(.dina(n4837), .dinb(n4796), .dout(n4846));
  jand g4762(.dina(n4846), .dinb(n4845), .dout(n4847));
  jand g4763(.dina(n4822), .dinb(n4802), .dout(n4848));
  jand g4764(.dina(n4823), .dinb(n4799), .dout(n4849));
  jor  g4765(.dina(n4849), .dinb(n4848), .dout(n4850));
  jor  g4766(.dina(n4820), .dinb(n4816), .dout(n4851));
  jand g4767(.dina(n4821), .dinb(n4808), .dout(n4852));
  jnot g4768(.din(n4852), .dout(n4853));
  jand g4769(.dina(n4853), .dinb(n4851), .dout(n4854));
  jnot g4770(.din(n4854), .dout(n4855));
  jor  g4771(.dina(n4807), .dinb(n4806), .dout(n4856));
  jor  g4772(.dina(n4760), .dinb(n3302), .dout(n4857));
  jand g4773(.dina(n4857), .dinb(n4856), .dout(n4858));
  jnot g4774(.din(n4858), .dout(n4859));
  jor  g4775(.dina(n3927), .dinb(n3198), .dout(n4860));
  jor  g4776(.dina(n3919), .dinb(n3200), .dout(n4861));
  jor  g4777(.dina(n3806), .dinb(n3204), .dout(n4862));
  jor  g4778(.dina(n3600), .dinb(n3202), .dout(n4863));
  jand g4779(.dina(n4863), .dinb(n4862), .dout(n4864));
  jand g4780(.dina(n4864), .dinb(n4861), .dout(n4865));
  jand g4781(.dina(n4865), .dinb(n4860), .dout(n4866));
  jxor g4782(.dina(n4866), .dinb(n954), .dout(n4867));
  jnot g4783(.din(n4867), .dout(n4868));
  jand g4784(.dina(n3302), .dinb(n954), .dout(n4869));
  jxor g4785(.dina(n4869), .dinb(n808), .dout(n4870));
  jand g4786(.dina(n3316), .dinb(n954), .dout(n4871));
  jxor g4787(.dina(n4871), .dinb(n4870), .dout(n4872));
  jxor g4788(.dina(n4872), .dinb(n4868), .dout(n4873));
  jxor g4789(.dina(n4873), .dinb(n4859), .dout(n4874));
  jxor g4790(.dina(n4874), .dinb(n4855), .dout(n4875));
  jxor g4791(.dina(n4875), .dinb(n4850), .dout(n4876));
  jand g4792(.dina(n592), .dinb(n323), .dout(n4877));
  jand g4793(.dina(n665), .dinb(n561), .dout(n4878));
  jand g4794(.dina(n4878), .dinb(n264), .dout(n4879));
  jand g4795(.dina(n4879), .dinb(n4877), .dout(n4880));
  jand g4796(.dina(n662), .dinb(n463), .dout(n4881));
  jand g4797(.dina(n4881), .dinb(n619), .dout(n4882));
  jand g4798(.dina(n822), .dinb(n413), .dout(n4883));
  jand g4799(.dina(n4883), .dinb(n4882), .dout(n4884));
  jand g4800(.dina(n749), .dinb(n343), .dout(n4885));
  jand g4801(.dina(n4885), .dinb(n882), .dout(n4886));
  jand g4802(.dina(n4886), .dinb(n4000), .dout(n4887));
  jand g4803(.dina(n4887), .dinb(n4884), .dout(n4888));
  jand g4804(.dina(n4888), .dinb(n4880), .dout(n4889));
  jand g4805(.dina(n4889), .dinb(n1231), .dout(n4890));
  jand g4806(.dina(n3693), .dinb(n2665), .dout(n4891));
  jand g4807(.dina(n4891), .dinb(n4890), .dout(n4892));
  jxor g4808(.dina(n4892), .dinb(n4876), .dout(n4893));
  jxor g4809(.dina(n4893), .dinb(n4847), .dout(n4894));
  jxor g4810(.dina(n4894), .dinb(n4843), .dout(n4895));
  jor  g4811(.dina(n4840), .dinb(n4839), .dout(n4896));
  jand g4812(.dina(n4896), .dinb(n4013), .dout(n4897));
  jxor g4813(.dina(n4897), .dinb(n4895), .dout(sin13 ));
  jand g4814(.dina(n4894), .dinb(n4843), .dout(n4899));
  jnot g4815(.din(n4876), .dout(n4900));
  jor  g4816(.dina(n4892), .dinb(n4900), .dout(n4901));
  jor  g4817(.dina(n4893), .dinb(n4847), .dout(n4902));
  jand g4818(.dina(n4902), .dinb(n4901), .dout(n4903));
  jand g4819(.dina(n4874), .dinb(n4855), .dout(n4904));
  jand g4820(.dina(n4875), .dinb(n4850), .dout(n4905));
  jor  g4821(.dina(n4905), .dinb(n4904), .dout(n4906));
  jand g4822(.dina(n4872), .dinb(n4868), .dout(n4907));
  jand g4823(.dina(n4873), .dinb(n4859), .dout(n4908));
  jor  g4824(.dina(n4908), .dinb(n4907), .dout(n4909));
  jand g4825(.dina(n4090), .dinb(n2883), .dout(n4910));
  jand g4826(.dina(n3807), .dinb(n2995), .dout(n4911));
  jand g4827(.dina(n3920), .dinb(n2887), .dout(n4912));
  jor  g4828(.dina(n4912), .dinb(n4911), .dout(n4913));
  jor  g4829(.dina(n4913), .dinb(n4910), .dout(n4914));
  jxor g4830(.dina(n4914), .dinb(n954), .dout(n4915));
  jand g4831(.dina(n3601), .dinb(n954), .dout(n4916));
  jnot g4832(.din(n4916), .dout(n4917));
  jand g4833(.dina(n4869), .dinb(n808), .dout(n4918));
  jand g4834(.dina(n4871), .dinb(n4870), .dout(n4919));
  jor  g4835(.dina(n4919), .dinb(n4918), .dout(n4920));
  jxor g4836(.dina(n4920), .dinb(n4917), .dout(n4921));
  jxor g4837(.dina(n4921), .dinb(n4915), .dout(n4922));
  jxor g4838(.dina(n4922), .dinb(n4909), .dout(n4923));
  jxor g4839(.dina(n4923), .dinb(n4906), .dout(n4924));
  jand g4840(.dina(n2456), .dinb(n712), .dout(n4925));
  jand g4841(.dina(n3307), .dinb(n2521), .dout(n4926));
  jand g4842(.dina(n4926), .dinb(n4925), .dout(n4927));
  jand g4843(.dina(n749), .dinb(n222), .dout(n4928));
  jand g4844(.dina(n4928), .dinb(n918), .dout(n4929));
  jand g4845(.dina(n935), .dinb(n251), .dout(n4930));
  jand g4846(.dina(n358), .dinb(n130), .dout(n4931));
  jand g4847(.dina(n4931), .dinb(n4930), .dout(n4932));
  jand g4848(.dina(n4932), .dinb(n4929), .dout(n4933));
  jand g4849(.dina(n4933), .dinb(n4927), .dout(n4934));
  jand g4850(.dina(n4934), .dinb(n622), .dout(n4935));
  jnot g4851(.din(n1669), .dout(n4936));
  jand g4852(.dina(n4936), .dinb(n675), .dout(n4937));
  jand g4853(.dina(n4937), .dinb(n4935), .dout(n4938));
  jand g4854(.dina(n4938), .dinb(n2575), .dout(n4939));
  jxor g4855(.dina(n4939), .dinb(n4924), .dout(n4940));
  jxor g4856(.dina(n4940), .dinb(n4903), .dout(n4941));
  jxor g4857(.dina(n4941), .dinb(n4899), .dout(n4942));
  jor  g4858(.dina(n4896), .dinb(n4895), .dout(n4943));
  jand g4859(.dina(n4943), .dinb(n4013), .dout(n4944));
  jxor g4860(.dina(n4944), .dinb(n4942), .dout(sin14 ));
  jand g4861(.dina(n4941), .dinb(n4899), .dout(n4946));
  jnot g4862(.din(n4924), .dout(n4947));
  jor  g4863(.dina(n4939), .dinb(n4947), .dout(n4948));
  jor  g4864(.dina(n4940), .dinb(n4903), .dout(n4949));
  jand g4865(.dina(n4949), .dinb(n4948), .dout(n4950));
  jand g4866(.dina(n4920), .dinb(n4917), .dout(n4951));
  jand g4867(.dina(n4921), .dinb(n4915), .dout(n4952));
  jor  g4868(.dina(n4952), .dinb(n4951), .dout(n4953));
  jnot g4869(.din(n4136), .dout(n4954));
  jand g4870(.dina(n4954), .dinb(n2883), .dout(n4955));
  jor  g4871(.dina(n4955), .dinb(n2995), .dout(n4956));
  jand g4872(.dina(n4956), .dinb(n3920), .dout(n4957));
  jxor g4873(.dina(n4957), .dinb(n820), .dout(n4958));
  jand g4874(.dina(n3900), .dinb(n954), .dout(n4959));
  jor  g4875(.dina(n4959), .dinb(n4958), .dout(n4960));
  jnot g4876(.din(n4957), .dout(n4961));
  jnot g4877(.din(n4959), .dout(n4962));
  jor  g4878(.dina(n4962), .dinb(n4961), .dout(n4963));
  jand g4879(.dina(n4963), .dinb(n4960), .dout(n4964));
  jxor g4880(.dina(n4964), .dinb(n4953), .dout(n4965));
  jand g4881(.dina(n4922), .dinb(n4909), .dout(n4966));
  jand g4882(.dina(n4923), .dinb(n4906), .dout(n4967));
  jor  g4883(.dina(n4967), .dinb(n4966), .dout(n4968));
  jxor g4884(.dina(n4968), .dinb(n4965), .dout(n4969));
  jand g4885(.dina(n614), .dinb(n436), .dout(n4970));
  jand g4886(.dina(n4970), .dinb(n303), .dout(n4971));
  jand g4887(.dina(n4971), .dinb(n1299), .dout(n4972));
  jand g4888(.dina(n387), .dinb(n383), .dout(n4973));
  jand g4889(.dina(n4973), .dinb(n4931), .dout(n4974));
  jand g4890(.dina(n645), .dinb(n624), .dout(n4975));
  jand g4891(.dina(n4975), .dinb(n992), .dout(n4976));
  jand g4892(.dina(n4976), .dinb(n680), .dout(n4977));
  jand g4893(.dina(n4977), .dinb(n4974), .dout(n4978));
  jand g4894(.dina(n4978), .dinb(n4832), .dout(n4979));
  jand g4895(.dina(n4979), .dinb(n1240), .dout(n4980));
  jand g4896(.dina(n4980), .dinb(n2461), .dout(n4981));
  jand g4897(.dina(n4981), .dinb(n4972), .dout(n4982));
  jxor g4898(.dina(n4982), .dinb(n4969), .dout(n4983));
  jxor g4899(.dina(n4983), .dinb(n4950), .dout(n4984));
  jxor g4900(.dina(n4984), .dinb(n4946), .dout(n4985));
  jor  g4901(.dina(n4943), .dinb(n4942), .dout(n4986));
  jand g4902(.dina(n4986), .dinb(n4013), .dout(n4987));
  jxor g4903(.dina(n4987), .dinb(n4985), .dout(sin15 ));
  jand g4904(.dina(n4984), .dinb(n4946), .dout(n4989));
  jnot g4905(.din(n4969), .dout(n4990));
  jor  g4906(.dina(n4982), .dinb(n4990), .dout(n4991));
  jor  g4907(.dina(n4983), .dinb(n4950), .dout(n4992));
  jand g4908(.dina(n4992), .dinb(n4991), .dout(n4993));
  jnot g4909(.din(n4993), .dout(n4994));
  jand g4910(.dina(n477), .dinb(n291), .dout(n4995));
  jand g4911(.dina(n4995), .dinb(n710), .dout(n4996));
  jand g4912(.dina(n543), .dinb(n384), .dout(n4997));
  jand g4913(.dina(n4997), .dinb(n4996), .dout(n4998));
  jand g4914(.dina(n4998), .dinb(n2334), .dout(n4999));
  jand g4915(.dina(n4880), .dinb(n3620), .dout(n5000));
  jand g4916(.dina(n5000), .dinb(n4999), .dout(n5001));
  jand g4917(.dina(n5001), .dinb(n3696), .dout(n5002));
  jand g4918(.dina(n5002), .dinb(n2382), .dout(n5003));
  jand g4919(.dina(n3600), .dinb(n954), .dout(n5004));
  jand g4920(.dina(n5004), .dinb(n3807), .dout(n5005));
  jnot g4921(.din(n5005), .dout(n5006));
  jand g4922(.dina(n5006), .dinb(n4960), .dout(n5007));
  jnot g4923(.din(n5007), .dout(n5008));
  jand g4924(.dina(n4964), .dinb(n4953), .dout(n5009));
  jand g4925(.dina(n4968), .dinb(n4965), .dout(n5010));
  jor  g4926(.dina(n5010), .dinb(n5009), .dout(n5011));
  jor  g4927(.dina(n3920), .dinb(n3600), .dout(n5012));
  jor  g4928(.dina(n3919), .dinb(n3601), .dout(n5013));
  jand g4929(.dina(n5013), .dinb(n954), .dout(n5014));
  jand g4930(.dina(n5014), .dinb(n5012), .dout(n5015));
  jxor g4931(.dina(n5015), .dinb(n5011), .dout(n5016));
  jxor g4932(.dina(n5016), .dinb(n5008), .dout(n5017));
  jxor g4933(.dina(n5017), .dinb(n5003), .dout(n5018));
  jxor g4934(.dina(n5018), .dinb(n4994), .dout(n5019));
  jxor g4935(.dina(n5019), .dinb(n4989), .dout(n5020));
  jor  g4936(.dina(n4986), .dinb(n4985), .dout(n5021));
  jand g4937(.dina(n5021), .dinb(n4013), .dout(n5022));
  jxor g4938(.dina(n5022), .dinb(n5020), .dout(sin16 ));
  jor  g4939(.dina(n5021), .dinb(n5020), .dout(n5024));
  jand g4940(.dina(n5024), .dinb(n4013), .dout(n5025));
  jand g4941(.dina(n5019), .dinb(n4989), .dout(n5026));
  jor  g4942(.dina(n5017), .dinb(n5003), .dout(n5027));
  jxor g4943(.dina(n5016), .dinb(n5007), .dout(n5028));
  jxor g4944(.dina(n5028), .dinb(n5003), .dout(n5029));
  jor  g4945(.dina(n5029), .dinb(n4993), .dout(n5030));
  jand g4946(.dina(n5030), .dinb(n5027), .dout(n5031));
  jand g4947(.dina(n461), .dinb(n372), .dout(n5032));
  jand g4948(.dina(n5032), .dinb(n619), .dout(n5033));
  jand g4949(.dina(n2736), .dinb(n507), .dout(n5034));
  jand g4950(.dina(n5034), .dinb(n5033), .dout(n5035));
  jand g4951(.dina(n365), .dinb(n277), .dout(n5036));
  jand g4952(.dina(n5036), .dinb(n422), .dout(n5037));
  jand g4953(.dina(n5037), .dinb(n443), .dout(n5038));
  jand g4954(.dina(n5038), .dinb(n5035), .dout(n5039));
  jand g4955(.dina(n5039), .dinb(n824), .dout(n5040));
  jand g4956(.dina(n5040), .dinb(n3256), .dout(n5041));
  jand g4957(.dina(n5041), .dinb(n860), .dout(n5042));
  jxor g4958(.dina(n5042), .dinb(n5031), .dout(n5043));
  jxor g4959(.dina(n5043), .dinb(n5026), .dout(n5044));
  jxor g4960(.dina(n5044), .dinb(n5025), .dout(sin17 ));
  jnot g4961(.din(n4013), .dout(n5046));
  jnot g4962(.din(n5024), .dout(n5047));
  jnot g4963(.din(n5026), .dout(n5048));
  jxor g4964(.dina(n5043), .dinb(n5048), .dout(n5049));
  jand g4965(.dina(n5049), .dinb(n5047), .dout(n5050));
  jor  g4966(.dina(n5050), .dinb(n5046), .dout(n5051));
  jnot g4967(.din(n5027), .dout(n5052));
  jand g4968(.dina(n5018), .dinb(n4994), .dout(n5053));
  jor  g4969(.dina(n5053), .dinb(n5052), .dout(n5054));
  jnot g4970(.din(n5042), .dout(n5055));
  jand g4971(.dina(n5055), .dinb(n5054), .dout(n5056));
  jand g4972(.dina(n5043), .dinb(n5026), .dout(n5057));
  jor  g4973(.dina(n5057), .dinb(n5056), .dout(n5058));
  jand g4974(.dina(n277), .dinb(n251), .dout(n5059));
  jand g4975(.dina(n5059), .dinb(n368), .dout(n5060));
  jand g4976(.dina(n5060), .dinb(n2396), .dout(n5061));
  jand g4977(.dina(n999), .dinb(n611), .dout(n5062));
  jand g4978(.dina(n5062), .dinb(n5061), .dout(n5063));
  jand g4979(.dina(n2658), .dinb(n1218), .dout(n5064));
  jand g4980(.dina(n5064), .dinb(n5063), .dout(n5065));
  jand g4981(.dina(n5065), .dinb(n1307), .dout(n5066));
  jand g4982(.dina(n5066), .dinb(n3663), .dout(n5067));
  jand g4983(.dina(n5067), .dinb(n834), .dout(n5068));
  jxor g4984(.dina(n5068), .dinb(n5058), .dout(n5069));
  jxor g4985(.dina(n5069), .dinb(n5051), .dout(sin18 ));
  jor  g4986(.dina(n5042), .dinb(n5031), .dout(n5071));
  jor  g4987(.dina(n5068), .dinb(n5071), .dout(n5072));
  jand g4988(.dina(n3257), .dinb(n681), .dout(n5073));
  jand g4989(.dina(n5073), .dinb(n987), .dout(n5074));
  jand g4990(.dina(n768), .dinb(n157), .dout(n5075));
  jand g4991(.dina(n5075), .dinb(n1209), .dout(n5076));
  jand g4992(.dina(n5076), .dinb(n4357), .dout(n5077));
  jand g4993(.dina(n5077), .dinb(n5074), .dout(n5078));
  jand g4994(.dina(n5078), .dinb(n3159), .dout(n5079));
  jand g4995(.dina(n5079), .dinb(n1175), .dout(n5080));
  jand g4996(.dina(n5080), .dinb(n4972), .dout(n5081));
  jxor g4997(.dina(n5081), .dinb(n5072), .dout(n5082));
  jnot g4998(.din(n5068), .dout(n5083));
  jand g4999(.dina(n5083), .dinb(n5057), .dout(n5084));
  jxor g5000(.dina(n5084), .dinb(n5082), .dout(n5085));
  jor  g5001(.dina(n5044), .dinb(n5024), .dout(n5086));
  jxor g5002(.dina(n5083), .dinb(n5058), .dout(n5087));
  jor  g5003(.dina(n5087), .dinb(n5086), .dout(n5088));
  jand g5004(.dina(n5088), .dinb(n4013), .dout(n5089));
  jxor g5005(.dina(n5089), .dinb(n5085), .dout(sin19 ));
  jand g5006(.dina(n5083), .dinb(n5056), .dout(n5091));
  jxor g5007(.dina(n5081), .dinb(n5091), .dout(n5092));
  jxor g5008(.dina(n5084), .dinb(n5092), .dout(n5093));
  jand g5009(.dina(n5069), .dinb(n5050), .dout(n5094));
  jand g5010(.dina(n5094), .dinb(n5093), .dout(n5095));
  jor  g5011(.dina(n5095), .dinb(n5046), .dout(n5096));
  jnot g5012(.din(n5081), .dout(n5097));
  jand g5013(.dina(n5097), .dinb(n5091), .dout(n5098));
  jand g5014(.dina(n5084), .dinb(n5082), .dout(n5099));
  jor  g5015(.dina(n5099), .dinb(n5098), .dout(n5100));
  jand g5016(.dina(n733), .dinb(n494), .dout(n5101));
  jand g5017(.dina(n5101), .dinb(n2542), .dout(n5102));
  jand g5018(.dina(n724), .dinb(n323), .dout(n5103));
  jand g5019(.dina(n5103), .dinb(n214), .dout(n5104));
  jand g5020(.dina(n5104), .dinb(n4355), .dout(n5105));
  jand g5021(.dina(n5105), .dinb(n5102), .dout(n5106));
  jand g5022(.dina(n5106), .dinb(n786), .dout(n5107));
  jand g5023(.dina(n5107), .dinb(n4589), .dout(n5108));
  jand g5024(.dina(n5108), .dinb(n636), .dout(n5109));
  jxor g5025(.dina(n5109), .dinb(n5100), .dout(n5110));
  jxor g5026(.dina(n5110), .dinb(n5096), .dout(sin20 ));
  jnot g5027(.din(n5109), .dout(n5112));
  jand g5028(.dina(n5112), .dinb(n5098), .dout(n5113));
  jand g5029(.dina(n3592), .dinb(n664), .dout(n5114));
  jand g5030(.dina(n5114), .dinb(n722), .dout(n5115));
  jand g5031(.dina(n5115), .dinb(n334), .dout(n5116));
  jnot g5032(.din(n5116), .dout(n5117));
  jxor g5033(.dina(n5117), .dinb(n5113), .dout(n5118));
  jand g5034(.dina(n5112), .dinb(n5099), .dout(n5119));
  jxor g5035(.dina(n5119), .dinb(n5118), .dout(n5120));
  jor  g5036(.dina(n5088), .dinb(n5085), .dout(n5121));
  jxor g5037(.dina(n5112), .dinb(n5100), .dout(n5122));
  jor  g5038(.dina(n5122), .dinb(n5121), .dout(n5123));
  jand g5039(.dina(n5123), .dinb(n4013), .dout(n5124));
  jxor g5040(.dina(n5124), .dinb(n5120), .dout(sin21 ));
  jor  g5041(.dina(n5123), .dinb(n5120), .dout(n5126));
  jand g5042(.dina(n5126), .dinb(n4013), .dout(n5127));
  jand g5043(.dina(n779), .dinb(n334), .dout(n5128));
  jnot g5044(.din(n5128), .dout(n5129));
  jand g5045(.dina(n5117), .dinb(n5113), .dout(n5130));
  jand g5046(.dina(n5119), .dinb(n5118), .dout(n5131));
  jor  g5047(.dina(n5131), .dinb(n5130), .dout(n5132));
  jxor g5048(.dina(n5132), .dinb(n5129), .dout(n5133));
  jxor g5049(.dina(n5133), .dinb(n5127), .dout(sin22 ));
  jnot g5050(.din(a21 ), .dout(n5135));
  jand g5051(.dina(n49), .dinb(n5135), .dout(n5136));
  jand g5052(.dina(n5136), .dinb(n207), .dout(n5137));
  jor  g5053(.dina(n5133), .dinb(n5126), .dout(n5138));
  jand g5054(.dina(n5138), .dinb(n4013), .dout(n5139));
  jand g5055(.dina(n5132), .dinb(n5129), .dout(n5140));
  jnot g5056(.din(n5130), .dout(n5141));
  jxor g5057(.dina(n5116), .dinb(n5113), .dout(n5142));
  jxor g5058(.dina(n5042), .dinb(n5054), .dout(n5143));
  jor  g5059(.dina(n5143), .dinb(n5048), .dout(n5144));
  jor  g5060(.dina(n5068), .dinb(n5144), .dout(n5145));
  jor  g5061(.dina(n5145), .dinb(n5092), .dout(n5146));
  jor  g5062(.dina(n5109), .dinb(n5146), .dout(n5147));
  jor  g5063(.dina(n5147), .dinb(n5142), .dout(n5148));
  jor  g5064(.dina(n5148), .dinb(n5141), .dout(n5149));
  jxor g5065(.dina(n5140), .dinb(n5139), .dout(n5151));
  jor  g5066(.dina(n5151), .dinb(n5137), .dout(sin23 ));
  jor  g5067(.dina(n5149), .dinb(n5128), .dout(n5153));
  jand g5068(.dina(n5153), .dinb(n5138), .dout(n5154));
  jxor g5069(.dina(n5119), .dinb(n5142), .dout(n5155));
  jand g5070(.dina(n5110), .dinb(n5095), .dout(n5156));
  jand g5071(.dina(n5156), .dinb(n5155), .dout(n5157));
  jand g5072(.dina(n5140), .dinb(n5157), .dout(n5158));
  jor  g5073(.dina(n5158), .dinb(n5137), .dout(n5159));
  jor  g5074(.dina(n5159), .dinb(n5154), .dout(n5160));
  jand g5075(.dina(n5160), .dinb(n4013), .dout(sin24 ));
endmodule


