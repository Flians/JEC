module rf_c3540(G1698, G330, G326, G343, G317, G311, G303, G294, G2897, G274, G250, G244, G238, G232, G322, G226, G223, G270, G200, G257, G77, G20, G125, G116, G283, G143, G45, G190, G68, G1, G58, G132, G33, G150, G87, G128, G97, G107, G124, G329, G264, G222, G50, G137, G159, G41, G169, G13, G179, G213, G409, G407, G381, G375, G378, G393, G353, G361, G390, G396, G351, G372, G384, G405, G358, G355, G369, G399, G364, G367, G402, G387);
    input G1698, G330, G326, G343, G317, G311, G303, G294, G2897, G274, G250, G244, G238, G232, G322, G226, G223, G270, G200, G257, G77, G20, G125, G116, G283, G143, G45, G190, G68, G1, G58, G132, G33, G150, G87, G128, G97, G107, G124, G329, G264, G222, G50, G137, G159, G41, G169, G13, G179, G213;
    output G409, G407, G381, G375, G378, G393, G353, G361, G390, G396, G351, G372, G384, G405, G358, G355, G369, G399, G364, G367, G402, G387;
    wire n74;
    wire n77;
    wire n80;
    wire n83;
    wire n87;
    wire n91;
    wire n95;
    wire n98;
    wire n101;
    wire n105;
    wire n108;
    wire n112;
    wire n115;
    wire n119;
    wire n122;
    wire n126;
    wire n129;
    wire n133;
    wire n137;
    wire n140;
    wire n144;
    wire n147;
    wire n151;
    wire n155;
    wire n159;
    wire n162;
    wire n165;
    wire n169;
    wire n172;
    wire n176;
    wire n180;
    wire n183;
    wire n187;
    wire n190;
    wire n193;
    wire n197;
    wire n201;
    wire n205;
    wire n209;
    wire n213;
    wire n216;
    wire n219;
    wire n222;
    wire n226;
    wire n230;
    wire n233;
    wire n237;
    wire n240;
    wire n244;
    wire n248;
    wire n252;
    wire n255;
    wire n259;
    wire n263;
    wire n267;
    wire n271;
    wire n275;
    wire n279;
    wire n283;
    wire n287;
    wire n290;
    wire n294;
    wire n298;
    wire n302;
    wire n306;
    wire n310;
    wire n313;
    wire n317;
    wire n321;
    wire n324;
    wire n328;
    wire n332;
    wire n336;
    wire n340;
    wire n343;
    wire n347;
    wire n350;
    wire n353;
    wire n357;
    wire n361;
    wire n365;
    wire n369;
    wire n372;
    wire n376;
    wire n380;
    wire n384;
    wire n388;
    wire n392;
    wire n396;
    wire n399;
    wire n403;
    wire n407;
    wire n410;
    wire n414;
    wire n418;
    wire n422;
    wire n426;
    wire n430;
    wire n434;
    wire n438;
    wire n442;
    wire n446;
    wire n450;
    wire n454;
    wire n457;
    wire n461;
    wire n465;
    wire n469;
    wire n473;
    wire n477;
    wire n481;
    wire n485;
    wire n489;
    wire n493;
    wire n497;
    wire n500;
    wire n504;
    wire n508;
    wire n512;
    wire n516;
    wire n520;
    wire n524;
    wire n528;
    wire n532;
    wire n535;
    wire n539;
    wire n543;
    wire n547;
    wire n551;
    wire n554;
    wire n558;
    wire n562;
    wire n566;
    wire n569;
    wire n573;
    wire n577;
    wire n581;
    wire n585;
    wire n589;
    wire n593;
    wire n597;
    wire n601;
    wire n604;
    wire n608;
    wire n612;
    wire n616;
    wire n620;
    wire n624;
    wire n628;
    wire n632;
    wire n635;
    wire n639;
    wire n643;
    wire n647;
    wire n651;
    wire n655;
    wire n659;
    wire n663;
    wire n667;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n695;
    wire n699;
    wire n703;
    wire n707;
    wire n711;
    wire n715;
    wire n719;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n778;
    wire n782;
    wire n785;
    wire n788;
    wire n792;
    wire n795;
    wire n799;
    wire n803;
    wire n807;
    wire n811;
    wire n815;
    wire n819;
    wire n823;
    wire n827;
    wire n831;
    wire n835;
    wire n839;
    wire n843;
    wire n847;
    wire n851;
    wire n855;
    wire n859;
    wire n863;
    wire n867;
    wire n871;
    wire n875;
    wire n879;
    wire n883;
    wire n887;
    wire n891;
    wire n895;
    wire n899;
    wire n903;
    wire n907;
    wire n911;
    wire n915;
    wire n918;
    wire n922;
    wire n926;
    wire n929;
    wire n933;
    wire n936;
    wire n940;
    wire n944;
    wire n948;
    wire n952;
    wire n956;
    wire n959;
    wire n963;
    wire n967;
    wire n971;
    wire n975;
    wire n979;
    wire n983;
    wire n987;
    wire n991;
    wire n995;
    wire n999;
    wire n1003;
    wire n1006;
    wire n1010;
    wire n1014;
    wire n1018;
    wire n1022;
    wire n1026;
    wire n1030;
    wire n1034;
    wire n1038;
    wire n1042;
    wire n1046;
    wire n1050;
    wire n1054;
    wire n1058;
    wire n1062;
    wire n1066;
    wire n1070;
    wire n1074;
    wire n1077;
    wire n1081;
    wire n1085;
    wire n1089;
    wire n1093;
    wire n1096;
    wire n1100;
    wire n1104;
    wire n1108;
    wire n1112;
    wire n1116;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1148;
    wire n1152;
    wire n1156;
    wire n1160;
    wire n1164;
    wire n1168;
    wire n1172;
    wire n1176;
    wire n1180;
    wire n1184;
    wire n1188;
    wire n1192;
    wire n1196;
    wire n1200;
    wire n1204;
    wire n1208;
    wire n1212;
    wire n1216;
    wire n1220;
    wire n1224;
    wire n1228;
    wire n1232;
    wire n1236;
    wire n1240;
    wire n1244;
    wire n1248;
    wire n1252;
    wire n1256;
    wire n1260;
    wire n1264;
    wire n1268;
    wire n1271;
    wire n1275;
    wire n1279;
    wire n1283;
    wire n1287;
    wire n1290;
    wire n1294;
    wire n1298;
    wire n1302;
    wire n1306;
    wire n1310;
    wire n1314;
    wire n1318;
    wire n1322;
    wire n1326;
    wire n1330;
    wire n1334;
    wire n1338;
    wire n1342;
    wire n1346;
    wire n1350;
    wire n1353;
    wire n1357;
    wire n1360;
    wire n1364;
    wire n1367;
    wire n1371;
    wire n1375;
    wire n1379;
    wire n1383;
    wire n1387;
    wire n1391;
    wire n1395;
    wire n1399;
    wire n1403;
    wire n1407;
    wire n1411;
    wire n1415;
    wire n1418;
    wire n1422;
    wire n1426;
    wire n1430;
    wire n1433;
    wire n1437;
    wire n1441;
    wire n1445;
    wire n1449;
    wire n1453;
    wire n1457;
    wire n1461;
    wire n1465;
    wire n1469;
    wire n1473;
    wire n1477;
    wire n1481;
    wire n1485;
    wire n1488;
    wire n1492;
    wire n1496;
    wire n1499;
    wire n1503;
    wire n1507;
    wire n1511;
    wire n1515;
    wire n1519;
    wire n1523;
    wire n1527;
    wire n1531;
    wire n1535;
    wire n1539;
    wire n1543;
    wire n1547;
    wire n1551;
    wire n1555;
    wire n1558;
    wire n1562;
    wire n1566;
    wire n1569;
    wire n1573;
    wire n1576;
    wire n1580;
    wire n1584;
    wire n1588;
    wire n1591;
    wire n1595;
    wire n1599;
    wire n1603;
    wire n1607;
    wire n1610;
    wire n1614;
    wire n1618;
    wire n1621;
    wire n1625;
    wire n1629;
    wire n1633;
    wire n1636;
    wire n1640;
    wire n1644;
    wire n1648;
    wire n1652;
    wire n1656;
    wire n1660;
    wire n1664;
    wire n1668;
    wire n1672;
    wire n1676;
    wire n1680;
    wire n1684;
    wire n1688;
    wire n1692;
    wire n1696;
    wire n1699;
    wire n1703;
    wire n1707;
    wire n1711;
    wire n1715;
    wire n1719;
    wire n1722;
    wire n1726;
    wire n1730;
    wire n1734;
    wire n1737;
    wire n1741;
    wire n1745;
    wire n1748;
    wire n1752;
    wire n1756;
    wire n1760;
    wire n1763;
    wire n1767;
    wire n1771;
    wire n1775;
    wire n1779;
    wire n1783;
    wire n1787;
    wire n1791;
    wire n1795;
    wire n1799;
    wire n1803;
    wire n1807;
    wire n1811;
    wire n1815;
    wire n1819;
    wire n1823;
    wire n1827;
    wire n1831;
    wire n1835;
    wire n1839;
    wire n1842;
    wire n1846;
    wire n1850;
    wire n1854;
    wire n1858;
    wire n1862;
    wire n1866;
    wire n1870;
    wire n1874;
    wire n1877;
    wire n1880;
    wire n1884;
    wire n1888;
    wire n1892;
    wire n1896;
    wire n1900;
    wire n1904;
    wire n1908;
    wire n1912;
    wire n1916;
    wire n1920;
    wire n1924;
    wire n1927;
    wire n1931;
    wire n1935;
    wire n1939;
    wire n1942;
    wire n1946;
    wire n1950;
    wire n1954;
    wire n1958;
    wire n1962;
    wire n1965;
    wire n1968;
    wire n1971;
    wire n1975;
    wire n1978;
    wire n1982;
    wire n1986;
    wire n1990;
    wire n1994;
    wire n1998;
    wire n2001;
    wire n2005;
    wire n2009;
    wire n2013;
    wire n2017;
    wire n2021;
    wire n2025;
    wire n2029;
    wire n2033;
    wire n2037;
    wire n2041;
    wire n2045;
    wire n2049;
    wire n2053;
    wire n2057;
    wire n2061;
    wire n2065;
    wire n2069;
    wire n2072;
    wire n2076;
    wire n2080;
    wire n2084;
    wire n2088;
    wire n2092;
    wire n2096;
    wire n2100;
    wire n2103;
    wire n2107;
    wire n2111;
    wire n2114;
    wire n2118;
    wire n2121;
    wire n2125;
    wire n2129;
    wire n2133;
    wire n2137;
    wire n2140;
    wire n2144;
    wire n2148;
    wire n2152;
    wire n2155;
    wire n2159;
    wire n2163;
    wire n2167;
    wire n2171;
    wire n2175;
    wire n2178;
    wire n2182;
    wire n2185;
    wire n2189;
    wire n2193;
    wire n2196;
    wire n2200;
    wire n2204;
    wire n2208;
    wire n2212;
    wire n2216;
    wire n2220;
    wire n2224;
    wire n2228;
    wire n2232;
    wire n2236;
    wire n2240;
    wire n2244;
    wire n2248;
    wire n2252;
    wire n2256;
    wire n2260;
    wire n2264;
    wire n2268;
    wire n2272;
    wire n2276;
    wire n2280;
    wire n2284;
    wire n2288;
    wire n2292;
    wire n2296;
    wire n2300;
    wire n2304;
    wire n2307;
    wire n2311;
    wire n2314;
    wire n2318;
    wire n2322;
    wire n2326;
    wire n2330;
    wire n2334;
    wire n2338;
    wire n2342;
    wire n2346;
    wire n2349;
    wire n2353;
    wire n2357;
    wire n2360;
    wire n2364;
    wire n2368;
    wire n2371;
    wire n2375;
    wire n2378;
    wire n2382;
    wire n2386;
    wire n2390;
    wire n2393;
    wire n2397;
    wire n2401;
    wire n2405;
    wire n2409;
    wire n2413;
    wire n2417;
    wire n2420;
    wire n2424;
    wire n2428;
    wire n2432;
    wire n2436;
    wire n2440;
    wire n2444;
    wire n2447;
    wire n2450;
    wire n2454;
    wire n2458;
    wire n2462;
    wire n2465;
    wire n2469;
    wire n2473;
    wire n2476;
    wire n2480;
    wire n2484;
    wire n2488;
    wire n2491;
    wire n2495;
    wire n2498;
    wire n2502;
    wire n2506;
    wire n2510;
    wire n2514;
    wire n2518;
    wire n2522;
    wire n2526;
    wire n2530;
    wire n2534;
    wire n2538;
    wire n2542;
    wire n2546;
    wire n2550;
    wire n2554;
    wire n2558;
    wire n2562;
    wire n2566;
    wire n2570;
    wire n2574;
    wire n2578;
    wire n2582;
    wire n2585;
    wire n2589;
    wire n2592;
    wire n2596;
    wire n2600;
    wire n2604;
    wire n2608;
    wire n2612;
    wire n2616;
    wire n2620;
    wire n2623;
    wire n2627;
    wire n2631;
    wire n2634;
    wire n2638;
    wire n2642;
    wire n2646;
    wire n2650;
    wire n2654;
    wire n2657;
    wire n2661;
    wire n2665;
    wire n2668;
    wire n2672;
    wire n2675;
    wire n2678;
    wire n2682;
    wire n2686;
    wire n2689;
    wire n2693;
    wire n2697;
    wire n2701;
    wire n2705;
    wire n2709;
    wire n2712;
    wire n2716;
    wire n2720;
    wire n2724;
    wire n2728;
    wire n2732;
    wire n2736;
    wire n2740;
    wire n2744;
    wire n2748;
    wire n2752;
    wire n2755;
    wire n2759;
    wire n2763;
    wire n2767;
    wire n2771;
    wire n2775;
    wire n2779;
    wire n2783;
    wire n2786;
    wire n2790;
    wire n2794;
    wire n2797;
    wire n2801;
    wire n2805;
    wire n2809;
    wire n2813;
    wire n2817;
    wire n2821;
    wire n2825;
    wire n2829;
    wire n2832;
    wire n2836;
    wire n2840;
    wire n2844;
    wire n2848;
    wire n2852;
    wire n2855;
    wire n2859;
    wire n2863;
    wire n2867;
    wire n2870;
    wire n2874;
    wire n2877;
    wire n2881;
    wire n2885;
    wire n2889;
    wire n2893;
    wire n2897;
    wire n2901;
    wire n2905;
    wire n2909;
    wire n2913;
    wire n2917;
    wire n2921;
    wire n2925;
    wire n2929;
    wire n2933;
    wire n2937;
    wire n2941;
    wire n2945;
    wire n2948;
    wire n2952;
    wire n2955;
    wire n2959;
    wire n2962;
    wire n2966;
    wire n2970;
    wire n2974;
    wire n2978;
    wire n2982;
    wire n2986;
    wire n2990;
    wire n2994;
    wire n2998;
    wire n3002;
    wire n3006;
    wire n3010;
    wire n3013;
    wire n3017;
    wire n3020;
    wire n3024;
    wire n3028;
    wire n3032;
    wire n3036;
    wire n3040;
    wire n3044;
    wire n3048;
    wire n3052;
    wire n3056;
    wire n3059;
    wire n3063;
    wire n3067;
    wire n3070;
    wire n3074;
    wire n3077;
    wire n3081;
    wire n3085;
    wire n3089;
    wire n3092;
    wire n3096;
    wire n3100;
    wire n3104;
    wire n3108;
    wire n3112;
    wire n3116;
    wire n3120;
    wire n3124;
    wire n3127;
    wire n3131;
    wire n3135;
    wire n3139;
    wire n3143;
    wire n3147;
    wire n3150;
    wire n3154;
    wire n3158;
    wire n3162;
    wire n3166;
    wire n3170;
    wire n3174;
    wire n3178;
    wire n3182;
    wire n3186;
    wire n3190;
    wire n3194;
    wire n3198;
    wire n3202;
    wire n3206;
    wire n3210;
    wire n3214;
    wire n3218;
    wire n3222;
    wire n3226;
    wire n3230;
    wire n3234;
    wire n3238;
    wire n3242;
    wire n3246;
    wire n3250;
    wire n3254;
    wire n3258;
    wire n3262;
    wire n3266;
    wire n3270;
    wire n3274;
    wire n3278;
    wire n3282;
    wire n3286;
    wire n3290;
    wire n3294;
    wire n3298;
    wire n3302;
    wire n3306;
    wire n3310;
    wire n3314;
    wire n3318;
    wire n3321;
    wire n3325;
    wire n3329;
    wire n3333;
    wire n3337;
    wire n3341;
    wire n3345;
    wire n3349;
    wire n3352;
    wire n3356;
    wire n3360;
    wire n3363;
    wire n3367;
    wire n3371;
    wire n3375;
    wire n3379;
    wire n3382;
    wire n3386;
    wire n3390;
    wire n3394;
    wire n3397;
    wire n3400;
    wire n3403;
    wire n3407;
    wire n3411;
    wire n3415;
    wire n3419;
    wire n3423;
    wire n3426;
    wire n3430;
    wire n3434;
    wire n3438;
    wire n3442;
    wire n3446;
    wire n3450;
    wire n3454;
    wire n3458;
    wire n3462;
    wire n3466;
    wire n3470;
    wire n3474;
    wire n3478;
    wire n3482;
    wire n3486;
    wire n3490;
    wire n3494;
    wire n3498;
    wire n3502;
    wire n3506;
    wire n3510;
    wire n3514;
    wire n3518;
    wire n3522;
    wire n3526;
    wire n3530;
    wire n3534;
    wire n3538;
    wire n3542;
    wire n3546;
    wire n3550;
    wire n3554;
    wire n3558;
    wire n3562;
    wire n3566;
    wire n3570;
    wire n3574;
    wire n3578;
    wire n3582;
    wire n3585;
    wire n3589;
    wire n3593;
    wire n3596;
    wire n3599;
    wire n3603;
    wire n3607;
    wire n3611;
    wire n3615;
    wire n3619;
    wire n3623;
    wire n3627;
    wire n3631;
    wire n3634;
    wire n3638;
    wire n3642;
    wire n3646;
    wire n3650;
    wire n3653;
    wire n3657;
    wire n3661;
    wire n3665;
    wire n3669;
    wire n3673;
    wire n3676;
    wire n3680;
    wire n3684;
    wire n3688;
    wire n3692;
    wire n3696;
    wire n3700;
    wire n3704;
    wire n3708;
    wire n3712;
    wire n3716;
    wire n3720;
    wire n3724;
    wire n3728;
    wire n3732;
    wire n3736;
    wire n3740;
    wire n3744;
    wire n3748;
    wire n3752;
    wire n3756;
    wire n3760;
    wire n3764;
    wire n3768;
    wire n3772;
    wire n3776;
    wire n3780;
    wire n3784;
    wire n3788;
    wire n3792;
    wire n3796;
    wire n3800;
    wire n3804;
    wire n3808;
    wire n3811;
    wire n3815;
    wire n3819;
    wire n3822;
    wire n3826;
    wire n3830;
    wire n3833;
    wire n3837;
    wire n3841;
    wire n3844;
    wire n3848;
    wire n3852;
    wire n3856;
    wire n3859;
    wire n3863;
    wire n3867;
    wire n3871;
    wire n3874;
    wire n3878;
    wire n3882;
    wire n3886;
    wire n3890;
    wire n3893;
    wire n3897;
    wire n3901;
    wire n3905;
    wire n3909;
    wire n3913;
    wire n3916;
    wire n3920;
    wire n3923;
    wire n3927;
    wire n3931;
    wire n3935;
    wire n3939;
    wire n3943;
    wire n3947;
    wire n3951;
    wire n3955;
    wire n3959;
    wire n3962;
    wire n3966;
    wire n3970;
    wire n3974;
    wire n3978;
    wire n3982;
    wire n3986;
    wire n3990;
    wire n3993;
    wire n3997;
    wire n4000;
    wire n4004;
    wire n4008;
    wire n4012;
    wire n4016;
    wire n4020;
    wire n4024;
    wire n4028;
    wire n4031;
    wire n4035;
    wire n4039;
    wire n4043;
    wire n4047;
    wire n4051;
    wire n4055;
    wire n4059;
    wire n4063;
    wire n4067;
    wire n4071;
    wire n4075;
    wire n4079;
    wire n4082;
    wire n4086;
    wire n4089;
    wire n4093;
    wire n4097;
    wire n4100;
    wire n4104;
    wire n4108;
    wire n4111;
    wire n4115;
    wire n4119;
    wire n4123;
    wire n4127;
    wire n4131;
    wire n4135;
    wire n4139;
    wire n4143;
    wire n4147;
    wire n4151;
    wire n4155;
    wire n4159;
    wire n4163;
    wire n4167;
    wire n4171;
    wire n4175;
    wire n4179;
    wire n4183;
    wire n4187;
    wire n4191;
    wire n4195;
    wire n4199;
    wire n4203;
    wire n4207;
    wire n4211;
    wire n4215;
    wire n4219;
    wire n4223;
    wire n4227;
    wire n4231;
    wire n4235;
    wire n4239;
    wire n4243;
    wire n4246;
    wire n4250;
    wire n4254;
    wire n4257;
    wire n4261;
    wire n4265;
    wire n4268;
    wire n4272;
    wire n4275;
    wire n4278;
    wire n4282;
    wire n4286;
    wire n4290;
    wire n4294;
    wire n4298;
    wire n4302;
    wire n4305;
    wire n4308;
    wire n4311;
    wire n4315;
    wire n4319;
    wire n4327;
    wire n4331;
    wire n4335;
    wire n4339;
    wire n4343;
    wire n4347;
    wire n4350;
    wire n4354;
    wire n4358;
    wire n4362;
    wire n4366;
    wire n4374;
    wire n6419;
    wire n6422;
    wire n6425;
    wire n6427;
    wire n6430;
    wire n6433;
    wire n6437;
    wire n6440;
    wire n6443;
    wire n6446;
    wire n6449;
    wire n6452;
    wire n6455;
    wire n6458;
    wire n6461;
    wire n6464;
    wire n6467;
    wire n6470;
    wire n6473;
    wire n6476;
    wire n6479;
    wire n6482;
    wire n6485;
    wire n6488;
    wire n6491;
    wire n6494;
    wire n6497;
    wire n6500;
    wire n6503;
    wire n6506;
    wire n6509;
    wire n6512;
    wire n6515;
    wire n6518;
    wire n6521;
    wire n6524;
    wire n6527;
    wire n6530;
    wire n6533;
    wire n6536;
    wire n6539;
    wire n6542;
    wire n6545;
    wire n6548;
    wire n6551;
    wire n6554;
    wire n6557;
    wire n6560;
    wire n6563;
    wire n6566;
    wire n6569;
    wire n6572;
    wire n6575;
    wire n6578;
    wire n6581;
    wire n6583;
    wire n6586;
    wire n6590;
    wire n6592;
    wire n6596;
    wire n6598;
    wire n6602;
    wire n6605;
    wire n6608;
    wire n6611;
    wire n6614;
    wire n6617;
    wire n6620;
    wire n6623;
    wire n6626;
    wire n6629;
    wire n6632;
    wire n6635;
    wire n6638;
    wire n6641;
    wire n6644;
    wire n6647;
    wire n6650;
    wire n6653;
    wire n6656;
    wire n6659;
    wire n6662;
    wire n6665;
    wire n6668;
    wire n6671;
    wire n6674;
    wire n6677;
    wire n6679;
    wire n6683;
    wire n6686;
    wire n6689;
    wire n6692;
    wire n6695;
    wire n6698;
    wire n6701;
    wire n6704;
    wire n6707;
    wire n6710;
    wire n6713;
    wire n6716;
    wire n6719;
    wire n6722;
    wire n6725;
    wire n6728;
    wire n6731;
    wire n6734;
    wire n6737;
    wire n6740;
    wire n6743;
    wire n6746;
    wire n6749;
    wire n6752;
    wire n6755;
    wire n6758;
    wire n6761;
    wire n6764;
    wire n6766;
    wire n6769;
    wire n6772;
    wire n6775;
    wire n6778;
    wire n6781;
    wire n6784;
    wire n6787;
    wire n6790;
    wire n6793;
    wire n6796;
    wire n6799;
    wire n6802;
    wire n6805;
    wire n6808;
    wire n6811;
    wire n6814;
    wire n6817;
    wire n6820;
    wire n6823;
    wire n6826;
    wire n6829;
    wire n6832;
    wire n6835;
    wire n6838;
    wire n6841;
    wire n6844;
    wire n6847;
    wire n6850;
    wire n6853;
    wire n6856;
    wire n6859;
    wire n6862;
    wire n6865;
    wire n6868;
    wire n6871;
    wire n6874;
    wire n6877;
    wire n6880;
    wire n6883;
    wire n6886;
    wire n6889;
    wire n6892;
    wire n6895;
    wire n6898;
    wire n6901;
    wire n6904;
    wire n6907;
    wire n6910;
    wire n6913;
    wire n6917;
    wire n6920;
    wire n6923;
    wire n6926;
    wire n6929;
    wire n6932;
    wire n6935;
    wire n6938;
    wire n6941;
    wire n6944;
    wire n6947;
    wire n6950;
    wire n6953;
    wire n6956;
    wire n6959;
    wire n6962;
    wire n6965;
    wire n6968;
    wire n6971;
    wire n6974;
    wire n6977;
    wire n6980;
    wire n6983;
    wire n6986;
    wire n6989;
    wire n6992;
    wire n6995;
    wire n6998;
    wire n7001;
    wire n7004;
    wire n7007;
    wire n7010;
    wire n7013;
    wire n7016;
    wire n7019;
    wire n7022;
    wire n7025;
    wire n7028;
    wire n7031;
    wire n7034;
    wire n7037;
    wire n7040;
    wire n7043;
    wire n7046;
    wire n7049;
    wire n7052;
    wire n7055;
    wire n7058;
    wire n7061;
    wire n7064;
    wire n7067;
    wire n7070;
    wire n7073;
    wire n7076;
    wire n7079;
    wire n7082;
    wire n7085;
    wire n7088;
    wire n7091;
    wire n7094;
    wire n7096;
    wire n7099;
    wire n7102;
    wire n7105;
    wire n7108;
    wire n7111;
    wire n7115;
    wire n7118;
    wire n7121;
    wire n7124;
    wire n7127;
    wire n7130;
    wire n7132;
    wire n7135;
    wire n7138;
    wire n7142;
    wire n7145;
    wire n7148;
    wire n7151;
    wire n7154;
    wire n7157;
    wire n7160;
    wire n7163;
    wire n7165;
    wire n7168;
    wire n7171;
    wire n7174;
    wire n7178;
    wire n7181;
    wire n7184;
    wire n7187;
    wire n7190;
    wire n7193;
    wire n7196;
    wire n7199;
    wire n7202;
    wire n7205;
    wire n7208;
    wire n7211;
    wire n7214;
    wire n7217;
    wire n7220;
    wire n7223;
    wire n7226;
    wire n7229;
    wire n7232;
    wire n7235;
    wire n7238;
    wire n7241;
    wire n7244;
    wire n7246;
    wire n7250;
    wire n7253;
    wire n7256;
    wire n7258;
    wire n7261;
    wire n7264;
    wire n7267;
    wire n7270;
    wire n7273;
    wire n7276;
    wire n7280;
    wire n7283;
    wire n7286;
    wire n7289;
    wire n7291;
    wire n7294;
    wire n7297;
    wire n7301;
    wire n7304;
    wire n7307;
    wire n7310;
    wire n7313;
    wire n7315;
    wire n7318;
    wire n7321;
    wire n7325;
    wire n7328;
    wire n7331;
    wire n7334;
    wire n7337;
    wire n7340;
    wire n7343;
    wire n7346;
    wire n7349;
    wire n7352;
    wire n7355;
    wire n7357;
    wire n7361;
    wire n7364;
    wire n7367;
    wire n7370;
    wire n7373;
    wire n7376;
    wire n7378;
    wire n7381;
    wire n7384;
    wire n7387;
    wire n7390;
    wire n7393;
    wire n7396;
    wire n7399;
    wire n7402;
    wire n7405;
    wire n7409;
    wire n7411;
    wire n7415;
    wire n7418;
    wire n7421;
    wire n7424;
    wire n7427;
    wire n7430;
    wire n7432;
    wire n7435;
    wire n7438;
    wire n7442;
    wire n7445;
    wire n7448;
    wire n7451;
    wire n7454;
    wire n7457;
    wire n7460;
    wire n7463;
    wire n7466;
    wire n7469;
    wire n7472;
    wire n7475;
    wire n7478;
    wire n7481;
    wire n7483;
    wire n7486;
    wire n7489;
    wire n7492;
    wire n7496;
    wire n7499;
    wire n7502;
    wire n7505;
    wire n7507;
    wire n7510;
    wire n7513;
    wire n7516;
    wire n7520;
    wire n7523;
    wire n7526;
    wire n7529;
    wire n7532;
    wire n7535;
    wire n7538;
    wire n7541;
    wire n7544;
    wire n7547;
    wire n7550;
    wire n7553;
    wire n7555;
    wire n7559;
    wire n7562;
    wire n7565;
    wire n7568;
    wire n7571;
    wire n7574;
    wire n7577;
    wire n7580;
    wire n7583;
    wire n7586;
    wire n7589;
    wire n7592;
    wire n7595;
    wire n7598;
    wire n7601;
    wire n7603;
    wire n7606;
    wire n7609;
    wire n7612;
    wire n7615;
    wire n7619;
    wire n7622;
    wire n7624;
    wire n7628;
    wire n7631;
    wire n7634;
    wire n7637;
    wire n7640;
    wire n7643;
    wire n7646;
    wire n7649;
    wire n7652;
    wire n7655;
    wire n7657;
    wire n7660;
    wire n7664;
    wire n7667;
    wire n7670;
    wire n7673;
    wire n7676;
    wire n7678;
    wire n7681;
    wire n7684;
    wire n7687;
    wire n7690;
    wire n7693;
    wire n7696;
    wire n7699;
    wire n7702;
    wire n7706;
    wire n7708;
    wire n7711;
    wire n7714;
    wire n7717;
    wire n7721;
    wire n7724;
    wire n7727;
    wire n7730;
    wire n7732;
    wire n7735;
    wire n7739;
    wire n7742;
    wire n7744;
    wire n7747;
    wire n7750;
    wire n7754;
    wire n7757;
    wire n7759;
    wire n7762;
    wire n7765;
    wire n7768;
    wire n7771;
    wire n7774;
    wire n7778;
    wire n7781;
    wire n7784;
    wire n7787;
    wire n7789;
    wire n7792;
    wire n7795;
    wire n7799;
    wire n7802;
    wire n7805;
    wire n7808;
    wire n7811;
    wire n7814;
    wire n7817;
    wire n7820;
    wire n7823;
    wire n7826;
    wire n7828;
    wire n7831;
    wire n7834;
    wire n7837;
    wire n7840;
    wire n7843;
    wire n7847;
    wire n7850;
    wire n7853;
    wire n7856;
    wire n7859;
    wire n7862;
    wire n7865;
    wire n7868;
    wire n7871;
    wire n7874;
    wire n7876;
    wire n7880;
    wire n7883;
    wire n7886;
    wire n7888;
    wire n7892;
    wire n7895;
    wire n7898;
    wire n7901;
    wire n7904;
    wire n7907;
    wire n7910;
    wire n7913;
    wire n7915;
    wire n7918;
    wire n7921;
    wire n7924;
    wire n7927;
    wire n7931;
    wire n7934;
    wire n7936;
    wire n7940;
    wire n7943;
    wire n7946;
    wire n7948;
    wire n7951;
    wire n7954;
    wire n7957;
    wire n7960;
    wire n7963;
    wire n7966;
    wire n7969;
    wire n7972;
    wire n7975;
    wire n7978;
    wire n7981;
    wire n7984;
    wire n7987;
    wire n7990;
    wire n7993;
    wire n7996;
    wire n7999;
    wire n8002;
    wire n8005;
    wire n8008;
    wire n8011;
    wire n8014;
    wire n8017;
    wire n8020;
    wire n8023;
    wire n8026;
    wire n8029;
    wire n8032;
    wire n8035;
    wire n8038;
    wire n8041;
    wire n8044;
    wire n8047;
    wire n8050;
    wire n8053;
    wire n8056;
    wire n8059;
    wire n8062;
    wire n8065;
    wire n8068;
    wire n8071;
    wire n8074;
    wire n8077;
    wire n8080;
    wire n8083;
    wire n8086;
    wire n8089;
    wire n8092;
    wire n8095;
    wire n8098;
    wire n8101;
    wire n8105;
    wire n8108;
    wire n8111;
    wire n8114;
    wire n8117;
    wire n8119;
    wire n8122;
    wire n8125;
    wire n8128;
    wire n8131;
    wire n8134;
    wire n8137;
    wire n8140;
    wire n8144;
    wire n8147;
    wire n8150;
    wire n8153;
    wire n8156;
    wire n8159;
    wire n8162;
    wire n8165;
    wire n8168;
    wire n8171;
    wire n8174;
    wire n8177;
    wire n8180;
    wire n8182;
    wire n8186;
    wire n8189;
    wire n8192;
    wire n8195;
    wire n8198;
    wire n8201;
    wire n8204;
    wire n8207;
    wire n8210;
    wire n8213;
    wire n8216;
    wire n8219;
    wire n8222;
    wire n8225;
    wire n8228;
    wire n8230;
    wire n8233;
    wire n8236;
    wire n8239;
    wire n8242;
    wire n8245;
    wire n8248;
    wire n8251;
    wire n8254;
    wire n8257;
    wire n8260;
    wire n8263;
    wire n8266;
    wire n8269;
    wire n8272;
    wire n8275;
    wire n8278;
    wire n8281;
    wire n8284;
    wire n8287;
    wire n8291;
    wire n8294;
    wire n8297;
    wire n8300;
    wire n8302;
    wire n8305;
    wire n8308;
    wire n8312;
    wire n8315;
    wire n8318;
    wire n8321;
    wire n8324;
    wire n8326;
    wire n8329;
    wire n8332;
    wire n8335;
    wire n8338;
    wire n8341;
    wire n8344;
    wire n8347;
    wire n8350;
    wire n8353;
    wire n8356;
    wire n8360;
    wire n8363;
    wire n8366;
    wire n8369;
    wire n8371;
    wire n8375;
    wire n8378;
    wire n8381;
    wire n8384;
    wire n8387;
    wire n8389;
    wire n8392;
    wire n8395;
    wire n8398;
    wire n8401;
    wire n8404;
    wire n8407;
    wire n8410;
    wire n8413;
    wire n8416;
    wire n8420;
    wire n8423;
    wire n8425;
    wire n8429;
    wire n8432;
    wire n8435;
    wire n8438;
    wire n8441;
    wire n8443;
    wire n8446;
    wire n8450;
    wire n8453;
    wire n8455;
    wire n8458;
    wire n8462;
    wire n8465;
    wire n8468;
    wire n8471;
    wire n8474;
    wire n8477;
    wire n8480;
    wire n8483;
    wire n8486;
    wire n8489;
    wire n8491;
    wire n8494;
    wire n8498;
    wire n8501;
    wire n8503;
    wire n8506;
    wire n8509;
    wire n8512;
    wire n8516;
    wire n8518;
    wire n8521;
    wire n8524;
    wire n8527;
    wire n8530;
    wire n8533;
    wire n8537;
    wire n8540;
    wire n8543;
    wire n8545;
    wire n8549;
    wire n8551;
    wire n8554;
    wire n8557;
    wire n8561;
    wire n8564;
    wire n8567;
    wire n8570;
    wire n8573;
    wire n8576;
    wire n8579;
    wire n8581;
    wire n8585;
    wire n8588;
    wire n8591;
    wire n8593;
    wire n8596;
    wire n8599;
    wire n8602;
    wire n8605;
    wire n8608;
    wire n8611;
    wire n8614;
    wire n8617;
    wire n8620;
    wire n8623;
    wire n8626;
    wire n8629;
    wire n8632;
    wire n8635;
    wire n8638;
    wire n8641;
    wire n8644;
    wire n8647;
    wire n8650;
    wire n8653;
    wire n8656;
    wire n8659;
    wire n8662;
    wire n8665;
    wire n8668;
    wire n8671;
    wire n8674;
    wire n8677;
    wire n8680;
    wire n8683;
    wire n8686;
    wire n8689;
    wire n8693;
    wire n8696;
    wire n8699;
    wire n8702;
    wire n8705;
    wire n8708;
    wire n8711;
    wire n8714;
    wire n8717;
    wire n8719;
    wire n8722;
    wire n8725;
    wire n8728;
    wire n8731;
    wire n8734;
    wire n8737;
    wire n8740;
    wire n8743;
    wire n8746;
    wire n8749;
    wire n8752;
    wire n8756;
    wire n8759;
    wire n8762;
    wire n8765;
    wire n8768;
    wire n8771;
    wire n8773;
    wire n8776;
    wire n8779;
    wire n8782;
    wire n8785;
    wire n8788;
    wire n8791;
    wire n8794;
    wire n8797;
    wire n8801;
    wire n8804;
    wire n8806;
    wire n8810;
    wire n8813;
    wire n8816;
    wire n8819;
    wire n8822;
    wire n8825;
    wire n8828;
    wire n8830;
    wire n8833;
    wire n8836;
    wire n8839;
    wire n8842;
    wire n8845;
    wire n8849;
    wire n8852;
    wire n8855;
    wire n8858;
    wire n8861;
    wire n8864;
    wire n8866;
    wire n8869;
    wire n8872;
    wire n8875;
    wire n8878;
    wire n8881;
    wire n8885;
    wire n8888;
    wire n8890;
    wire n8893;
    wire n8896;
    wire n8899;
    wire n8902;
    wire n8905;
    wire n8908;
    wire n8911;
    wire n8914;
    wire n8917;
    wire n8920;
    wire n8923;
    wire n8926;
    wire n8929;
    wire n8932;
    wire n8935;
    wire n8938;
    wire n8941;
    wire n8944;
    wire n8947;
    wire n8950;
    wire n8953;
    wire n8956;
    wire n8959;
    wire n8962;
    wire n8965;
    wire n8968;
    wire n8971;
    wire n8974;
    wire n8978;
    wire n8981;
    wire n8983;
    wire n8986;
    wire n8989;
    wire n8992;
    wire n8995;
    wire n8998;
    wire n9001;
    wire n9004;
    wire n9007;
    wire n9010;
    wire n9013;
    wire n9016;
    wire n9019;
    wire n9022;
    wire n9025;
    wire n9028;
    wire n9031;
    wire n9034;
    wire n9037;
    wire n9040;
    wire n9043;
    wire n9046;
    wire n9049;
    wire n9052;
    wire n9055;
    wire n9058;
    wire n9061;
    wire n9064;
    wire n9067;
    wire n9070;
    wire n9073;
    wire n9077;
    wire n9080;
    wire n9083;
    wire n9085;
    wire n9088;
    wire n9091;
    wire n9094;
    wire n9097;
    wire n9100;
    wire n9103;
    wire n9106;
    wire n9109;
    wire n9112;
    wire n9115;
    wire n9118;
    wire n9121;
    wire n9124;
    wire n9127;
    wire n9130;
    wire n9133;
    wire n9136;
    wire n9139;
    wire n9142;
    wire n9145;
    wire n9148;
    wire n9151;
    wire n9154;
    wire n9157;
    wire n9160;
    wire n9163;
    wire n9166;
    wire n9169;
    wire n9172;
    wire n9175;
    wire n9178;
    wire n9181;
    wire n9184;
    wire n9187;
    wire n9190;
    wire n9193;
    wire n9196;
    wire n9199;
    wire n9202;
    wire n9205;
    wire n9208;
    wire n9211;
    wire n9214;
    wire n9217;
    wire n9220;
    wire n9223;
    wire n9226;
    wire n9229;
    wire n9232;
    wire n9235;
    wire n9238;
    wire n9241;
    wire n9244;
    wire n9247;
    wire n9250;
    wire n9253;
    wire n9256;
    wire n9259;
    wire n9262;
    wire n9265;
    wire n9268;
    wire n9271;
    wire n9274;
    wire n9277;
    wire n9280;
    wire n9283;
    wire n9286;
    wire n9289;
    wire n9292;
    wire n9295;
    wire n9298;
    wire n9301;
    wire n9304;
    wire n9307;
    wire n9310;
    wire n9313;
    wire n9316;
    wire n9319;
    wire n9322;
    wire n9325;
    wire n9328;
    wire n9331;
    wire n9334;
    wire n9337;
    wire n9340;
    wire n9343;
    wire n9346;
    wire n9349;
    wire n9352;
    wire n9355;
    wire n9358;
    wire n9361;
    wire n9364;
    wire n9367;
    wire n9371;
    wire n9373;
    wire n9376;
    wire n9379;
    wire n9382;
    wire n9385;
    wire n9388;
    wire n9391;
    wire n9394;
    wire n9397;
    wire n9400;
    wire n9403;
    wire n9406;
    wire n9409;
    wire n9412;
    wire n9415;
    wire n9418;
    wire n9421;
    wire n9424;
    wire n9427;
    wire n9430;
    wire n9433;
    wire n9436;
    wire n9439;
    wire n9442;
    wire n9445;
    wire n9448;
    wire n9451;
    wire n9454;
    wire n9457;
    wire n9460;
    wire n9463;
    wire n9466;
    wire n9469;
    wire n9472;
    wire n9475;
    wire n9478;
    wire n9481;
    wire n9484;
    wire n9487;
    wire n9490;
    wire n9493;
    wire n9496;
    wire n9499;
    wire n9502;
    wire n9505;
    wire n9508;
    wire n9511;
    wire n9514;
    wire n9517;
    wire n9520;
    wire n9523;
    wire n9526;
    wire n9529;
    wire n9532;
    wire n9535;
    wire n9538;
    wire n9541;
    wire n9544;
    wire n9547;
    wire n9550;
    wire n9553;
    wire n9556;
    wire n9559;
    wire n9562;
    wire n9565;
    wire n9568;
    wire n9571;
    wire n9574;
    wire n9577;
    wire n9580;
    wire n9583;
    wire n9586;
    wire n9589;
    wire n9592;
    wire n9595;
    wire n9598;
    wire n9601;
    wire n9604;
    wire n9607;
    wire n9610;
    wire n9613;
    wire n9616;
    wire n9619;
    wire n9622;
    wire n9625;
    wire n9628;
    wire n9631;
    wire n9634;
    wire n9637;
    wire n9640;
    wire n9643;
    wire n9646;
    wire n9649;
    wire n9652;
    wire n9655;
    wire n9658;
    wire n9661;
    wire n9664;
    wire n9667;
    wire n9670;
    wire n9673;
    wire n9676;
    wire n9679;
    wire n9682;
    wire n9685;
    wire n9688;
    wire n9691;
    wire n9694;
    wire n9697;
    wire n9700;
    wire n9703;
    wire n9706;
    wire n9709;
    wire n9712;
    wire n9715;
    wire n9718;
    wire n9721;
    wire n9724;
    wire n9727;
    wire n9730;
    wire n9733;
    wire n9736;
    wire n9739;
    wire n9742;
    wire n9745;
    wire n9748;
    wire n9751;
    wire n9754;
    wire n9757;
    wire n9760;
    wire n9764;
    wire n9766;
    wire n9769;
    wire n9772;
    wire n9775;
    wire n9779;
    wire n9782;
    wire n9785;
    wire n9787;
    wire n9790;
    wire n9793;
    wire n9796;
    wire n9799;
    wire n9802;
    wire n9805;
    wire n9808;
    wire n9812;
    wire n9815;
    wire n9818;
    wire n9821;
    wire n9824;
    wire n9827;
    wire n9829;
    wire n9832;
    wire n9835;
    wire n9838;
    wire n9841;
    wire n9845;
    wire n9847;
    wire n9850;
    wire n9853;
    wire n9856;
    wire n9859;
    wire n9862;
    wire n9865;
    wire n9868;
    wire n9871;
    wire n9874;
    wire n9877;
    wire n9880;
    wire n9883;
    wire n9886;
    wire n9889;
    wire n9892;
    wire n9895;
    wire n9898;
    wire n9902;
    wire n9905;
    wire n9907;
    wire n9910;
    wire n9913;
    wire n9916;
    wire n9919;
    wire n9922;
    wire n9925;
    wire n9928;
    wire n9931;
    wire n9934;
    wire n9938;
    wire n9940;
    wire n9943;
    wire n9946;
    wire n9949;
    wire n9952;
    wire n9955;
    wire n9958;
    wire n9961;
    wire n9964;
    wire n9968;
    wire n9970;
    wire n9974;
    wire n9976;
    wire n9979;
    wire n9982;
    wire n9985;
    wire n9989;
    wire n9992;
    wire n9995;
    wire n9997;
    wire n10000;
    wire n10003;
    wire n10006;
    wire n10009;
    wire n10012;
    wire n10015;
    wire n10018;
    wire n10021;
    wire n10024;
    wire n10027;
    wire n10031;
    wire n10034;
    wire n10036;
    wire n10039;
    wire n10042;
    wire n10045;
    wire n10048;
    wire n10051;
    wire n10054;
    wire n10057;
    wire n10060;
    wire n10063;
    wire n10066;
    wire n10069;
    wire n10072;
    wire n10075;
    wire n10078;
    wire n10081;
    wire n10084;
    wire n10087;
    wire n10090;
    wire n10093;
    wire n10096;
    wire n10099;
    wire n10102;
    wire n10105;
    wire n10108;
    wire n10111;
    wire n10114;
    wire n10117;
    wire n10120;
    wire n10123;
    wire n10126;
    wire n10129;
    wire n10132;
    wire n10135;
    wire n10138;
    wire n10141;
    wire n10144;
    wire n10147;
    wire n10150;
    wire n10153;
    wire n10156;
    wire n10159;
    wire n10162;
    wire n10165;
    wire n10168;
    wire n10171;
    wire n10174;
    wire n10177;
    wire n10180;
    wire n10183;
    wire n10186;
    wire n10189;
    wire n10192;
    wire n10195;
    wire n10198;
    wire n10201;
    wire n10204;
    wire n10207;
    wire n10210;
    wire n10213;
    wire n10216;
    wire n10219;
    wire n10222;
    wire n10225;
    wire n10228;
    wire n10231;
    wire n10234;
    wire n10237;
    wire n10240;
    wire n10243;
    wire n10246;
    wire n10249;
    wire n10252;
    wire n10255;
    wire n10259;
    wire n10262;
    wire n10265;
    wire n10267;
    wire n10270;
    wire n10273;
    wire n10276;
    wire n10279;
    wire n10282;
    wire n10285;
    wire n10288;
    wire n10291;
    wire n10294;
    wire n10297;
    wire n10300;
    wire n10303;
    wire n10306;
    wire n10310;
    wire n10312;
    wire n10315;
    wire n10319;
    wire n10321;
    wire n10324;
    wire n10328;
    wire n10331;
    wire n10333;
    wire n10336;
    wire n10339;
    wire n10342;
    wire n10345;
    wire n10348;
    wire n10351;
    wire n10354;
    wire n10357;
    wire n10360;
    wire n10363;
    wire n10366;
    wire n10369;
    wire n10372;
    wire n10376;
    wire n10379;
    wire n10381;
    wire n10385;
    wire n10387;
    wire n10390;
    wire n10393;
    wire n10396;
    wire n10399;
    wire n10402;
    wire n10405;
    wire n10408;
    wire n10411;
    wire n10414;
    wire n10417;
    wire n10420;
    wire n10423;
    wire n10426;
    wire n10429;
    wire n10432;
    wire n10435;
    wire n10438;
    wire n10441;
    wire n10444;
    wire n10447;
    wire n10450;
    wire n10453;
    wire n10456;
    wire n10459;
    wire n10462;
    wire n10465;
    wire n10468;
    wire n10471;
    wire n10474;
    wire n10477;
    wire n10480;
    wire n10483;
    wire n10486;
    wire n10489;
    wire n10492;
    wire n10495;
    wire n10498;
    wire n10501;
    wire n10505;
    wire n10507;
    wire n10510;
    wire n10513;
    wire n10516;
    wire n10519;
    wire n10522;
    wire n10525;
    wire n10528;
    wire n10531;
    wire n10534;
    wire n10537;
    wire n10540;
    wire n10543;
    wire n10546;
    wire n10549;
    wire n10552;
    wire n10555;
    wire n10558;
    wire n10561;
    wire n10564;
    wire n10567;
    wire n10570;
    wire n10574;
    wire n10576;
    wire n10579;
    wire n10583;
    wire n10585;
    wire n10588;
    wire n10591;
    wire n10594;
    wire n10597;
    wire n10600;
    wire n10603;
    wire n10606;
    wire n10609;
    wire n10613;
    wire n10616;
    wire n10618;
    wire n10621;
    wire n10624;
    wire n10627;
    wire n10630;
    wire n10633;
    wire n10636;
    wire n10639;
    wire n10642;
    wire n10645;
    wire n10648;
    wire n10652;
    wire n10655;
    wire n10657;
    wire n10660;
    wire n10663;
    wire n10666;
    wire n10669;
    wire n10672;
    wire n10675;
    wire n10679;
    wire n10682;
    wire n10684;
    wire n10687;
    wire n10690;
    wire n10693;
    wire n10696;
    wire n10699;
    wire n10702;
    wire n10705;
    wire n10708;
    wire n10711;
    wire n10714;
    wire n10717;
    wire n10720;
    wire n10723;
    wire n10726;
    wire n10729;
    wire n10732;
    wire n10735;
    wire n10738;
    wire n10741;
    wire n10744;
    wire n10747;
    wire n10750;
    wire n10753;
    wire n10756;
    wire n10759;
    wire n10762;
    wire n10765;
    wire n10768;
    wire n10771;
    wire n10774;
    wire n10777;
    wire n10780;
    wire n10783;
    wire n10786;
    wire n10789;
    wire n10792;
    wire n10796;
    wire n10798;
    wire n10801;
    wire n10804;
    wire n10807;
    wire n10810;
    wire n10813;
    wire n10816;
    wire n10819;
    wire n10822;
    wire n10825;
    wire n10828;
    wire n10831;
    wire n10834;
    wire n10837;
    wire n10840;
    wire n10843;
    wire n10846;
    wire n10849;
    wire n10852;
    wire n10855;
    wire n10858;
    wire n10861;
    wire n10864;
    wire n10867;
    wire n10870;
    wire n10873;
    wire n10876;
    wire n10879;
    wire n10882;
    wire n10886;
    wire n10888;
    wire n10891;
    wire n10894;
    wire n10897;
    wire n10900;
    wire n10903;
    wire n10906;
    wire n10910;
    wire n10913;
    wire n10916;
    wire n10919;
    wire n10922;
    wire n10924;
    wire n10927;
    wire n10930;
    wire n10933;
    wire n10936;
    wire n10939;
    wire n10942;
    wire n10945;
    wire n10948;
    wire n10951;
    wire n10954;
    wire n10957;
    wire n10960;
    wire n10963;
    wire n10966;
    wire n10969;
    wire n10972;
    wire n10975;
    wire n10978;
    wire n10981;
    wire n10984;
    wire n10988;
    wire n10990;
    wire n10993;
    wire n10996;
    wire n10999;
    wire n11002;
    wire n11005;
    wire n11008;
    wire n11011;
    wire n11014;
    wire n11017;
    wire n11020;
    wire n11023;
    wire n11026;
    wire n11029;
    wire n11032;
    wire n11035;
    wire n11038;
    wire n11041;
    wire n11044;
    wire n11047;
    wire n11050;
    wire n11053;
    wire n11056;
    wire n11059;
    wire n11062;
    wire n11065;
    wire n11068;
    wire n11071;
    wire n11074;
    wire n11077;
    wire n11080;
    wire n11083;
    wire n11086;
    wire n11089;
    wire n11092;
    wire n11095;
    wire n11098;
    wire n11101;
    wire n11104;
    wire n11107;
    wire n11110;
    wire n11113;
    wire n11116;
    wire n11119;
    wire n11122;
    wire n11125;
    wire n11128;
    wire n11131;
    wire n11134;
    wire n11137;
    wire n11140;
    wire n11143;
    wire n11146;
    wire n11149;
    wire n11152;
    wire n11155;
    wire n11158;
    wire n11161;
    wire n11164;
    wire n11168;
    wire n11171;
    wire n11173;
    wire n11176;
    wire n11179;
    wire n11182;
    wire n11185;
    wire n11188;
    wire n11191;
    wire n11194;
    wire n11197;
    wire n11200;
    wire n11203;
    wire n11206;
    wire n11209;
    wire n11212;
    wire n11216;
    wire n11218;
    wire n11221;
    wire n11224;
    wire n11227;
    wire n11230;
    wire n11233;
    wire n11237;
    wire n11239;
    wire n11242;
    wire n11245;
    wire n11248;
    wire n11251;
    wire n11254;
    wire n11257;
    wire n11260;
    wire n11263;
    wire n11266;
    wire n11269;
    wire n11272;
    wire n11275;
    wire n11278;
    wire n11281;
    wire n11284;
    wire n11287;
    wire n11290;
    wire n11293;
    wire n11296;
    wire n11299;
    wire n11302;
    wire n11306;
    wire n11308;
    wire n11311;
    wire n11314;
    wire n11317;
    wire n11320;
    wire n11323;
    wire n11326;
    wire n11329;
    wire n11332;
    wire n11335;
    wire n11338;
    wire n11341;
    wire n11344;
    wire n11347;
    wire n11350;
    wire n11353;
    wire n11356;
    wire n11359;
    wire n11362;
    wire n11365;
    wire n11368;
    wire n11371;
    wire n11374;
    wire n11377;
    wire n11380;
    wire n11383;
    wire n11386;
    wire n11389;
    wire n11392;
    wire n11395;
    wire n11398;
    wire n11401;
    wire n11404;
    wire n11407;
    wire n11410;
    wire n11413;
    wire n11416;
    wire n11419;
    wire n11422;
    wire n11425;
    wire n11428;
    wire n11431;
    wire n11434;
    wire n11437;
    wire n11440;
    wire n11443;
    wire n11446;
    wire n11449;
    wire n11452;
    wire n11455;
    wire n11458;
    wire n11461;
    wire n11464;
    wire n11467;
    wire n11470;
    wire n11473;
    wire n11476;
    wire n11479;
    wire n11482;
    wire n11485;
    wire n11488;
    wire n11491;
    wire n11494;
    wire n11497;
    wire n11500;
    wire n11503;
    wire n11506;
    wire n11509;
    wire n11512;
    wire n11515;
    wire n11518;
    wire n11521;
    wire n11524;
    wire n11527;
    wire n11530;
    wire n11533;
    wire n11536;
    wire n11539;
    wire n11542;
    wire n11545;
    wire n11548;
    wire n11551;
    wire n11554;
    wire n11557;
    wire n11560;
    wire n11563;
    wire n11566;
    wire n11569;
    wire n11572;
    wire n11575;
    wire n11578;
    wire n11581;
    wire n11584;
    wire n11587;
    wire n11590;
    wire n11593;
    wire n11596;
    wire n11599;
    wire n11602;
    wire n11605;
    wire n11608;
    wire n11611;
    wire n11614;
    wire n11617;
    wire n11620;
    wire n11623;
    wire n11626;
    wire n11629;
    wire n11632;
    wire n11635;
    wire n11638;
    wire n11641;
    wire n11644;
    wire n11647;
    wire n11653;
    wire n11656;
    wire n11659;
    wire n11662;
    wire n11665;
    wire n11668;
    wire n11671;
    wire n11674;
    wire n11677;
    wire n11680;
    wire n11683;
    wire n11686;
    wire n11689;
    wire n11692;
    wire n11695;
    wire n11698;
    wire n11701;
    wire n11704;
    wire n11707;
    wire n11710;
    wire n11713;
    wire n11716;
    wire n11719;
    wire n11725;
    wire n11728;
    wire n11731;
    wire n11734;
    wire n11737;
    wire n11740;
    wire n11743;
    wire n11746;
    wire n11749;
    wire n11752;
    wire n11755;
    wire n11758;
    wire n11761;
    wire n11764;
    wire n11767;
    wire n11770;
    wire n11773;
    wire n11776;
    wire n11779;
    wire n11782;
    wire n11788;
    wire n11791;
    wire n11794;
    wire n11797;
    wire n11800;
    wire n11803;
    wire n11806;
    wire n11809;
    wire n11812;
    wire n11815;
    wire n11818;
    wire n11821;
    wire n11824;
    wire n11827;
    wire n11830;
    wire n11833;
    wire n11836;
    wire n11839;
    wire n11842;
    wire n11845;
    wire n11848;
    wire n11851;
    wire n11854;
    wire n11860;
    wire n11863;
    wire n11866;
    wire n11869;
    wire n11872;
    wire n11875;
    wire n11878;
    wire n11881;
    wire n11884;
    wire n11887;
    wire n11890;
    wire n11893;
    wire n11896;
    wire n11899;
    wire n11902;
    wire n11905;
    wire n11908;
    wire n11911;
    wire n11914;
    wire n11917;
    wire n11920;
    wire n11923;
    wire n11926;
    wire n11932;
    wire n11935;
    wire n11938;
    wire n11941;
    wire n11944;
    wire n11947;
    wire n11950;
    wire n11953;
    wire n11956;
    wire n11959;
    wire n11962;
    wire n11965;
    wire n11968;
    wire n11974;
    wire n11977;
    wire n11980;
    wire n11983;
    wire n11986;
    wire n11989;
    wire n11992;
    wire n11995;
    wire n11998;
    wire n12001;
    wire n12004;
    wire n12010;
    wire n12013;
    wire n12016;
    wire n12019;
    wire n12022;
    wire n12025;
    wire n12028;
    wire n12031;
    wire n12034;
    wire n12037;
    wire n12043;
    wire n12046;
    wire n12049;
    wire n12052;
    wire n12055;
    wire n12058;
    wire n12061;
    wire n12064;
    wire n12067;
    wire n12070;
    wire n12076;
    wire n12079;
    wire n12082;
    wire n12085;
    wire n12088;
    wire n12091;
    wire n12094;
    wire n12097;
    wire n12100;
    wire n12103;
    wire n12109;
    wire n12112;
    wire n12115;
    wire n12118;
    wire n12121;
    wire n12124;
    wire n12127;
    wire n12133;
    wire n12136;
    wire n12139;
    wire n12142;
    wire n12148;
    wire n12151;
    wire n12154;
    wire n12157;
    wire n12163;
    wire n12166;
    wire n12169;
    wire n12172;
    wire n12175;
    wire n12178;
    wire n12184;
    wire n12187;
    wire n12190;
    wire n12193;
    wire n12196;
    wire n12202;
    wire n12205;
    wire n12208;
    wire n12211;
    wire n12217;
    wire n12220;
    wire n12226;
    wire n12229;
    wire n12232;
    wire n12235;
    jnot g0000(.din(G77), .dout(n74));
    jnot g0001(.din(G50), .dout(n77));
    jnot g0002(.din(G58), .dout(n80));
    jnot g0003(.din(G68), .dout(n83));
    jand g0004(.dinb(n80), .dina(n83), .dout(n87));
    jor g0005(.dinb(n8635), .dina(n87), .dout(n91));
    jand g0006(.dinb(n6427), .dina(n91), .dout(n95));
    jnot g0007(.din(G97), .dout(n98));
    jdff g0008(.din(G107), .dout(n101));
    jand g0009(.dinb(n98), .dina(n101), .dout(n105));
    jnot g0010(.din(n105), .dout(n108));
    jand g0011(.dinb(n11095), .dina(n108), .dout(n112));
    jnot g0012(.din(n112), .dout(n115));
    jand g0013(.dinb(G1), .dina(G20), .dout(n119));
    jnot g0014(.din(G226), .dout(n122));
    jor g0015(.dinb(n77), .dina(n122), .dout(n126));
    jnot g0016(.din(G264), .dout(n129));
    jor g0017(.dinb(n101), .dina(n129), .dout(n133));
    jand g0018(.dinb(n126), .dina(n133), .dout(n137));
    jnot g0019(.din(G257), .dout(n140));
    jor g0020(.dinb(n98), .dina(n140), .dout(n144));
    jnot g0021(.din(G238), .dout(n147));
    jor g0022(.dinb(n83), .dina(n147), .dout(n151));
    jand g0023(.dinb(n144), .dina(n151), .dout(n155));
    jand g0024(.dinb(n137), .dina(n155), .dout(n159));
    jnot g0025(.din(G87), .dout(n162));
    jnot g0026(.din(G250), .dout(n165));
    jor g0027(.dinb(n162), .dina(n165), .dout(n169));
    jnot g0028(.din(G232), .dout(n172));
    jor g0029(.dinb(n80), .dina(n172), .dout(n176));
    jand g0030(.dinb(n169), .dina(n176), .dout(n180));
    jnot g0031(.din(G244), .dout(n183));
    jor g0032(.dinb(n74), .dina(n183), .dout(n187));
    jnot g0033(.din(G116), .dout(n190));
    jnot g0034(.din(G270), .dout(n193));
    jor g0035(.dinb(n190), .dina(n193), .dout(n197));
    jand g0036(.dinb(n187), .dina(n197), .dout(n201));
    jand g0037(.dinb(n180), .dina(n201), .dout(n205));
    jand g0038(.dinb(n159), .dina(n205), .dout(n209));
    jor g0039(.dinb(n11008), .dina(n209), .dout(n213));
    jnot g0040(.din(G20), .dout(n216));
    jnot g0041(.din(G1), .dout(n219));
    jnot g0042(.din(G13), .dout(n222));
    jor g0043(.dinb(n219), .dina(n222), .dout(n226));
    jor g0044(.dinb(n11125), .dina(n226), .dout(n230));
    jnot g0045(.din(n87), .dout(n233));
    jand g0046(.dinb(n8647), .dina(n233), .dout(n237));
    jnot g0047(.din(n237), .dout(n240));
    jor g0048(.dinb(n6583), .dina(n240), .dout(n244));
    jand g0049(.dinb(n11473), .dina(n222), .dout(n248));
    jand g0050(.dinb(n11161), .dina(n248), .dout(n252));
    jnot g0051(.din(n252), .dout(n255));
    jand g0052(.dinb(n140), .dina(n129), .dout(n259));
    jor g0053(.dinb(n6433), .dina(n259), .dout(n263));
    jor g0054(.dinb(n255), .dina(n6425), .dout(n267));
    jand g0055(.dinb(n244), .dina(n6422), .dout(n271));
    jand g0056(.dinb(n6419), .dina(n271), .dout(n275));
    jxor g0057(.dinb(G264), .dina(G270), .dout(n279));
    jxor g0058(.dinb(n165), .dina(n10723), .dout(n283));
    jxor g0059(.dinb(n7559), .dina(n283), .dout(n287));
    jnot g0060(.din(n287), .dout(n290));
    jxor g0061(.dinb(G238), .dina(G244), .dout(n294));
    jxor g0062(.dinb(n122), .dina(n9946), .dout(n298));
    jxor g0063(.dinb(n7664), .dina(n298), .dout(n302));
    jxor g0064(.dinb(n290), .dina(n7660), .dout(n306));
    jxor g0065(.dinb(G58), .dina(G68), .dout(n310));
    jnot g0066(.din(n310), .dout(n313));
    jxor g0067(.dinb(G50), .dina(G77), .dout(n317));
    jxor g0068(.dinb(n313), .dina(n7826), .dout(n321));
    jnot g0069(.din(n321), .dout(n324));
    jxor g0070(.dinb(G107), .dina(G116), .dout(n328));
    jxor g0071(.dinb(n162), .dina(n11083), .dout(n332));
    jxor g0072(.dinb(n7364), .dina(n332), .dout(n336));
    jxor g0073(.dinb(n324), .dina(n7361), .dout(n340));
    jnot g0074(.din(G169), .dout(n343));
    jand g0075(.dinb(G1), .dina(G13), .dout(n347));
    jnot g0076(.din(G33), .dout(n350));
    jnot g0077(.din(G41), .dout(n353));
    jor g0078(.dinb(n350), .dina(n353), .dout(n357));
    jand g0079(.dinb(n11458), .dina(n357), .dout(n361));
    jand g0080(.dinb(n350), .dina(n11374), .dout(n365));
    jand g0081(.dinb(n11377), .dina(n365), .dout(n369));
    jnot g0082(.din(G1698), .dout(n372));
    jand g0083(.dinb(n350), .dina(n372), .dout(n376));
    jand g0084(.dinb(n11350), .dina(n376), .dout(n380));
    jand g0085(.dinb(G33), .dina(G116), .dout(n384));
    jor g0086(.dinb(n380), .dina(n11314), .dout(n388));
    jor g0087(.dinb(n11306), .dina(n388), .dout(n392));
    jand g0088(.dinb(n11401), .dina(n392), .dout(n396));
    jnot g0089(.din(G45), .dout(n399));
    jor g0090(.dinb(n11470), .dina(n399), .dout(n403));
    jand g0091(.dinb(n11290), .dina(n403), .dout(n407));
    jnot g0092(.din(n407), .dout(n410));
    jand g0093(.dinb(G33), .dina(G41), .dout(n414));
    jor g0094(.dinb(n226), .dina(n11237), .dout(n418));
    jor g0095(.dinb(n11227), .dina(n403), .dout(n422));
    jand g0096(.dinb(n418), .dina(n422), .dout(n426));
    jand g0097(.dinb(n410), .dina(n426), .dout(n430));
    jor g0098(.dinb(n396), .dina(n11216), .dout(n434));
    jand g0099(.dinb(n11497), .dina(n434), .dout(n438));
    jand g0100(.dinb(G33), .dina(G97), .dout(n442));
    jand g0101(.dinb(n350), .dina(n11137), .dout(n446));
    jor g0102(.dinb(n11161), .dina(n446), .dout(n450));
    jor g0103(.dinb(n11171), .dina(n450), .dout(n454));
    jnot g0104(.din(n454), .dout(n457));
    jor g0105(.dinb(n219), .dina(n216), .dout(n461));
    jor g0106(.dinb(n11155), .dina(n461), .dout(n465));
    jand g0107(.dinb(n11239), .dina(n465), .dout(n469));
    jand g0108(.dinb(n11089), .dina(n105), .dout(n473));
    jand g0109(.dinb(n11158), .dina(n473), .dout(n477));
    jor g0110(.dinb(n469), .dina(n477), .dout(n481));
    jor g0111(.dinb(n457), .dina(n481), .dout(n485));
    jand g0112(.dinb(n219), .dina(n11164), .dout(n489));
    jand g0113(.dinb(n11464), .dina(n489), .dout(n493));
    jand g0114(.dinb(n11086), .dina(n493), .dout(n497));
    jnot g0115(.din(n497), .dout(n500));
    jand g0116(.dinb(n11209), .dina(n119), .dout(n504));
    jor g0117(.dinb(n11455), .dina(n504), .dout(n508));
    jor g0118(.dinb(n508), .dina(n493), .dout(n512));
    jand g0119(.dinb(n219), .dina(n11206), .dout(n516));
    jor g0120(.dinb(n11089), .dina(n516), .dout(n520));
    jor g0121(.dinb(n512), .dina(n10988), .dout(n524));
    jand g0122(.dinb(n500), .dina(n524), .dout(n528));
    jand g0123(.dinb(n485), .dina(n528), .dout(n532));
    jnot g0124(.din(G179), .dout(n535));
    jor g0125(.dinb(n10891), .dina(n372), .dout(n539));
    jor g0126(.dinb(n10894), .dina(n539), .dout(n543));
    jor g0127(.dinb(G33), .dina(G1698), .dout(n547));
    jor g0128(.dinb(n147), .dina(n547), .dout(n551));
    jnot g0129(.din(n384), .dout(n554));
    jand g0130(.dinb(n551), .dina(n554), .dout(n558));
    jand g0131(.dinb(n543), .dina(n558), .dout(n562));
    jor g0132(.dinb(n11233), .dina(n562), .dout(n566));
    jnot g0133(.din(G274), .dout(n569));
    jand g0134(.dinb(n219), .dina(n11266), .dout(n573));
    jand g0135(.dinb(n10886), .dina(n573), .dout(n577));
    jor g0136(.dinb(n361), .dina(n577), .dout(n581));
    jor g0137(.dinb(n11248), .dina(n581), .dout(n585));
    jand g0138(.dinb(n566), .dina(n585), .dout(n589));
    jand g0139(.dinb(n10922), .dina(n589), .dout(n593));
    jor g0140(.dinb(n532), .dina(n593), .dout(n597));
    jor g0141(.dinb(n438), .dina(n597), .dout(n601));
    jnot g0142(.din(n532), .dout(n604));
    jand g0143(.dinb(n10846), .dina(n589), .dout(n608));
    jand g0144(.dinb(n10798), .dina(n434), .dout(n612));
    jor g0145(.dinb(n10796), .dina(n612), .dout(n616));
    jor g0146(.dinb(n10873), .dina(n616), .dout(n620));
    jand g0147(.dinb(n10876), .dina(n620), .dout(n624));
    jor g0148(.dinb(n11287), .dina(n539), .dout(n628));
    jand g0149(.dinb(G33), .dina(G283), .dout(n632));
    jnot g0150(.din(n632), .dout(n635));
    jor g0151(.dinb(n183), .dina(n547), .dout(n639));
    jand g0152(.dinb(n635), .dina(n639), .dout(n643));
    jand g0153(.dinb(n628), .dina(n643), .dout(n647));
    jor g0154(.dinb(n10792), .dina(n647), .dout(n651));
    jor g0155(.dinb(n10882), .dina(n361), .dout(n655));
    jor g0156(.dinb(n11431), .dina(n403), .dout(n659));
    jor g0157(.dinb(n655), .dina(n10738), .dout(n663));
    jand g0158(.dinb(n11425), .dina(n573), .dout(n667));
    jor g0159(.dinb(n361), .dina(n667), .dout(n671));
    jor g0160(.dinb(n10699), .dina(n671), .dout(n675));
    jand g0161(.dinb(n663), .dina(n675), .dout(n679));
    jand g0162(.dinb(n10682), .dina(n679), .dout(n683));
    jor g0163(.dinb(n11497), .dina(n683), .dout(n687));
    jand g0164(.dinb(n11299), .dina(n365), .dout(n691));
    jand g0165(.dinb(n11395), .dina(n376), .dout(n695));
    jor g0166(.dinb(n10747), .dina(n695), .dout(n699));
    jor g0167(.dinb(n10679), .dina(n699), .dout(n703));
    jand g0168(.dinb(n10693), .dina(n703), .dout(n707));
    jand g0169(.dinb(n11218), .dina(n418), .dout(n711));
    jand g0170(.dinb(n711), .dina(n10684), .dout(n715));
    jand g0171(.dinb(n418), .dina(n659), .dout(n719));
    jand g0172(.dinb(n10711), .dina(n719), .dout(n723));
    jor g0173(.dinb(n715), .dina(n723), .dout(n727));
    jor g0174(.dinb(n707), .dina(n727), .dout(n731));
    jor g0175(.dinb(n10900), .dina(n731), .dout(n735));
    jand g0176(.dinb(n687), .dina(n735), .dout(n739));
    jand g0177(.dinb(G33), .dina(G107), .dout(n743));
    jand g0178(.dinb(n350), .dina(n10636), .dout(n747));
    jor g0179(.dinb(n11023), .dina(n747), .dout(n751));
    jor g0180(.dinb(n10655), .dina(n751), .dout(n755));
    jand g0181(.dinb(G97), .dina(G107), .dout(n759));
    jor g0182(.dinb(n216), .dina(n759), .dout(n763));
    jor g0183(.dinb(n105), .dina(n763), .dout(n767));
    jand g0184(.dinb(n755), .dina(n10630), .dout(n771));
    jand g0185(.dinb(n10993), .dina(n771), .dout(n775));
    jnot g0186(.din(n775), .dout(n778));
    jand g0187(.dinb(n11077), .dina(n493), .dout(n782));
    jnot g0188(.din(n782), .dout(n785));
    jnot g0189(.din(n516), .dout(n788));
    jand g0190(.dinb(n11173), .dina(n788), .dout(n792));
    jnot g0191(.din(n792), .dout(n795));
    jor g0192(.dinb(n10990), .dina(n795), .dout(n799));
    jand g0193(.dinb(n10616), .dina(n799), .dout(n803));
    jand g0194(.dinb(n778), .dina(n803), .dout(n807));
    jor g0195(.dinb(n739), .dina(n10613), .dout(n811));
    jand g0196(.dinb(n10798), .dina(n731), .dout(n815));
    jor g0197(.dinb(n11476), .dina(n216), .dout(n819));
    jor g0198(.dinb(n11242), .dina(n819), .dout(n823));
    jand g0199(.dinb(n469), .dina(n10583), .dout(n827));
    jand g0200(.dinb(n827), .dina(n10618), .dout(n831));
    jor g0201(.dinb(n10621), .dina(n831), .dout(n835));
    jor g0202(.dinb(n10627), .dina(n835), .dout(n839));
    jand g0203(.dinb(n10843), .dina(n683), .dout(n843));
    jor g0204(.dinb(n839), .dina(n843), .dout(n847));
    jor g0205(.dinb(n10574), .dina(n847), .dout(n851));
    jand g0206(.dinb(n811), .dina(n851), .dout(n855));
    jand g0207(.dinb(n624), .dina(n855), .dout(n859));
    jand g0208(.dinb(n10567), .dina(n365), .dout(n863));
    jand g0209(.dinb(G33), .dina(G303), .dout(n867));
    jand g0210(.dinb(n10732), .dina(n376), .dout(n871));
    jor g0211(.dinb(n10507), .dina(n871), .dout(n875));
    jor g0212(.dinb(n10505), .dina(n875), .dout(n879));
    jand g0213(.dinb(n10687), .dina(n879), .dout(n883));
    jand g0214(.dinb(n10492), .dina(n719), .dout(n887));
    jor g0215(.dinb(n715), .dina(n887), .dout(n891));
    jor g0216(.dinb(n883), .dina(n891), .dout(n895));
    jand g0217(.dinb(n11497), .dina(n895), .dout(n899));
    jand g0218(.dinb(n350), .dina(n11203), .dout(n903));
    jor g0219(.dinb(n11020), .dina(n903), .dout(n907));
    jor g0220(.dinb(n10741), .dina(n907), .dout(n911));
    jand g0221(.dinb(n11164), .dina(n190), .dout(n915));
    jnot g0222(.din(n915), .dout(n918));
    jand g0223(.dinb(n508), .dina(n918), .dout(n922));
    jand g0224(.dinb(n911), .dina(n922), .dout(n926));
    jnot g0225(.din(n926), .dout(n929));
    jand g0226(.dinb(n10435), .dina(n493), .dout(n933));
    jnot g0227(.din(n933), .dout(n936));
    jor g0228(.dinb(n10444), .dina(n516), .dout(n940));
    jor g0229(.dinb(n512), .dina(n10417), .dout(n944));
    jand g0230(.dinb(n936), .dina(n944), .dout(n948));
    jand g0231(.dinb(n929), .dina(n948), .dout(n952));
    jor g0232(.dinb(n10405), .dina(n539), .dout(n956));
    jnot g0233(.din(n867), .dout(n959));
    jor g0234(.dinb(n140), .dina(n547), .dout(n963));
    jand g0235(.dinb(n959), .dina(n963), .dout(n967));
    jand g0236(.dinb(n956), .dina(n967), .dout(n971));
    jor g0237(.dinb(n10411), .dina(n971), .dout(n975));
    jor g0238(.dinb(n10387), .dina(n671), .dout(n979));
    jand g0239(.dinb(n663), .dina(n979), .dout(n983));
    jand g0240(.dinb(n10385), .dina(n983), .dout(n987));
    jand g0241(.dinb(n10897), .dina(n987), .dout(n991));
    jor g0242(.dinb(n10414), .dina(n991), .dout(n995));
    jor g0243(.dinb(n10379), .dina(n995), .dout(n999));
    jand g0244(.dinb(n10798), .dina(n895), .dout(n1003));
    jnot g0245(.din(n940), .dout(n1006));
    jand g0246(.dinb(n827), .dina(n10376), .dout(n1010));
    jor g0247(.dinb(n10420), .dina(n1010), .dout(n1014));
    jor g0248(.dinb(n10438), .dina(n1014), .dout(n1018));
    jand g0249(.dinb(n10354), .dina(n987), .dout(n1022));
    jor g0250(.dinb(n1018), .dina(n1022), .dout(n1026));
    jor g0251(.dinb(n10331), .dina(n1026), .dout(n1030));
    jand g0252(.dinb(n999), .dina(n1030), .dout(n1034));
    jor g0253(.dinb(n10675), .dina(n162), .dout(n1038));
    jand g0254(.dinb(n10597), .dina(n1038), .dout(n1042));
    jand g0255(.dinb(n10888), .dina(n1042), .dout(n1046));
    jor g0256(.dinb(n469), .dina(n1046), .dout(n1050));
    jor g0257(.dinb(n10459), .dina(n1050), .dout(n1054));
    jand g0258(.dinb(n10657), .dina(n1054), .dout(n1058));
    jand g0259(.dinb(n10579), .dina(n1050), .dout(n1062));
    jor g0260(.dinb(n1058), .dina(n10328), .dout(n1066));
    jand g0261(.dinb(n11068), .dina(n788), .dout(n1070));
    jand g0262(.dinb(n827), .dina(n10319), .dout(n1074));
    jnot g0263(.din(n1074), .dout(n1077));
    jand g0264(.dinb(n1066), .dina(n10310), .dout(n1081));
    jor g0265(.dinb(n10708), .dina(n539), .dout(n1085));
    jor g0266(.dinb(n165), .dina(n547), .dout(n1089));
    jand g0267(.dinb(G33), .dina(G294), .dout(n1093));
    jnot g0268(.din(n1093), .dout(n1096));
    jand g0269(.dinb(n1089), .dina(n1096), .dout(n1100));
    jand g0270(.dinb(n1085), .dina(n1100), .dout(n1104));
    jor g0271(.dinb(n10408), .dina(n1104), .dout(n1108));
    jor g0272(.dinb(n10396), .dina(n671), .dout(n1112));
    jand g0273(.dinb(n663), .dina(n1112), .dout(n1116));
    jand g0274(.dinb(n10265), .dina(n1116), .dout(n1120));
    jand g0275(.dinb(n10903), .dina(n1120), .dout(n1124));
    jand g0276(.dinb(n10726), .dina(n365), .dout(n1128));
    jand g0277(.dinb(n11293), .dina(n376), .dout(n1132));
    jor g0278(.dinb(n1132), .dina(n10267), .dout(n1136));
    jor g0279(.dinb(n10262), .dina(n1136), .dout(n1140));
    jand g0280(.dinb(n11419), .dina(n1140), .dout(n1144));
    jand g0281(.dinb(n10555), .dina(n719), .dout(n1148));
    jor g0282(.dinb(n715), .dina(n1148), .dout(n1152));
    jor g0283(.dinb(n1144), .dina(n1152), .dout(n1156));
    jand g0284(.dinb(n11479), .dina(n1156), .dout(n1160));
    jor g0285(.dinb(n1124), .dina(n1160), .dout(n1164));
    jor g0286(.dinb(n1081), .dina(n1164), .dout(n1168));
    jand g0287(.dinb(n350), .dina(n11092), .dout(n1172));
    jor g0288(.dinb(n10456), .dina(n1172), .dout(n1176));
    jor g0289(.dinb(n11308), .dina(n1176), .dout(n1180));
    jand g0290(.dinb(n10471), .dina(n1180), .dout(n1184));
    jand g0291(.dinb(n10585), .dina(n1184), .dout(n1188));
    jor g0292(.dinb(n11035), .dina(n1188), .dout(n1192));
    jor g0293(.dinb(n10426), .dina(n1184), .dout(n1196));
    jand g0294(.dinb(n1192), .dina(n10259), .dout(n1200));
    jor g0295(.dinb(n1200), .dina(n10312), .dout(n1204));
    jor g0296(.dinb(n10333), .dina(n1156), .dout(n1208));
    jor g0297(.dinb(n10822), .dina(n1120), .dout(n1212));
    jand g0298(.dinb(n1208), .dina(n1212), .dout(n1216));
    jor g0299(.dinb(n1204), .dina(n1216), .dout(n1220));
    jand g0300(.dinb(n1168), .dina(n1220), .dout(n1224));
    jand g0301(.dinb(n1034), .dina(n1224), .dout(n1228));
    jand g0302(.dinb(n859), .dina(n1228), .dout(n1232));
    jand g0303(.dinb(n9940), .dina(n376), .dout(n1236));
    jand g0304(.dinb(n11368), .dina(n365), .dout(n1240));
    jor g0305(.dinb(n10655), .dina(n1240), .dout(n1244));
    jor g0306(.dinb(n9938), .dina(n1244), .dout(n1248));
    jand g0307(.dinb(n11419), .dina(n1248), .dout(n1252));
    jand g0308(.dinb(n353), .dina(n399), .dout(n1256));
    jor g0309(.dinb(n10609), .dina(n1256), .dout(n1260));
    jand g0310(.dinb(n418), .dina(n1260), .dout(n1264));
    jand g0311(.dinb(n11383), .dina(n1264), .dout(n1268));
    jnot g0312(.din(n1260), .dout(n1271));
    jand g0313(.dinb(n711), .dina(n1271), .dout(n1275));
    jor g0314(.dinb(n1268), .dina(n1275), .dout(n1279));
    jor g0315(.dinb(n1252), .dina(n1279), .dout(n1283));
    jand g0316(.dinb(n11479), .dina(n1283), .dout(n1287));
    jnot g0317(.din(n1287), .dout(n1290));
    jand g0318(.dinb(G33), .dina(G87), .dout(n1294));
    jand g0319(.dinb(n350), .dina(n9865), .dout(n1298));
    jor g0320(.dinb(n9895), .dina(n1298), .dout(n1302));
    jor g0321(.dinb(n9905), .dina(n1302), .dout(n1306));
    jor g0322(.dinb(n216), .dina(n10636), .dout(n1310));
    jand g0323(.dinb(n508), .dina(n9845), .dout(n1314));
    jand g0324(.dinb(n1306), .dina(n1314), .dout(n1318));
    jand g0325(.dinb(n9838), .dina(n493), .dout(n1322));
    jand g0326(.dinb(n10633), .dina(n819), .dout(n1326));
    jand g0327(.dinb(n827), .dina(n9827), .dout(n1330));
    jor g0328(.dinb(n9821), .dina(n1330), .dout(n1334));
    jor g0329(.dinb(n9815), .dina(n1334), .dout(n1338));
    jor g0330(.dinb(n10945), .dina(n1283), .dout(n1342));
    jand g0331(.dinb(n1338), .dina(n1342), .dout(n1346));
    jand g0332(.dinb(n1290), .dina(n1346), .dout(n1350));
    jnot g0333(.din(n1350), .dout(n1353));
    jand g0334(.dinb(n10822), .dina(n1283), .dout(n1357));
    jnot g0335(.din(G190), .dout(n1360));
    jor g0336(.dinb(n9787), .dina(n1283), .dout(n1364));
    jnot g0337(.din(n1364), .dout(n1367));
    jor g0338(.dinb(n9808), .dina(n1367), .dout(n1371));
    jor g0339(.dinb(n9785), .dina(n1371), .dout(n1375));
    jand g0340(.dinb(n1353), .dina(n1375), .dout(n1379));
    jand g0341(.dinb(n8443), .dina(n376), .dout(n1383));
    jand g0342(.dinb(n9961), .dina(n365), .dout(n1387));
    jor g0343(.dinb(n11171), .dina(n1387), .dout(n1391));
    jor g0344(.dinb(n8441), .dina(n1391), .dout(n1395));
    jand g0345(.dinb(n11419), .dina(n1395), .dout(n1399));
    jand g0346(.dinb(n11356), .dina(n1264), .dout(n1403));
    jor g0347(.dinb(n1275), .dina(n1403), .dout(n1407));
    jor g0348(.dinb(n1399), .dina(n1407), .dout(n1411));
    jand g0349(.dinb(n11479), .dina(n1411), .dout(n1415));
    jnot g0350(.din(n1415), .dout(n1418));
    jand g0351(.dinb(n11134), .dina(n819), .dout(n1422));
    jand g0352(.dinb(n827), .dina(n8438), .dout(n1426));
    jand g0353(.dinb(n222), .dina(n350), .dout(n1430));
    jnot g0354(.din(n1430), .dout(n1433));
    jand g0355(.dinb(n11002), .dina(n1433), .dout(n1437));
    jor g0356(.dinb(n8581), .dina(n1437), .dout(n1441));
    jand g0357(.dinb(n8602), .dina(n1441), .dout(n1445));
    jand g0358(.dinb(G33), .dina(G77), .dout(n1449));
    jand g0359(.dinb(n350), .dina(n8665), .dout(n1453));
    jor g0360(.dinb(n8549), .dina(n1453), .dout(n1457));
    jand g0361(.dinb(n9853), .dina(n1457), .dout(n1461));
    jand g0362(.dinb(n10999), .dina(n1461), .dout(n1465));
    jor g0363(.dinb(n1445), .dina(n8432), .dout(n1469));
    jor g0364(.dinb(n8429), .dina(n1469), .dout(n1473));
    jor g0365(.dinb(n10924), .dina(n1411), .dout(n1477));
    jand g0366(.dinb(n1473), .dina(n1477), .dout(n1481));
    jand g0367(.dinb(n1418), .dina(n1481), .dout(n1485));
    jnot g0368(.din(n1485), .dout(n1488));
    jand g0369(.dinb(n10822), .dina(n1411), .dout(n1492));
    jor g0370(.dinb(n9787), .dina(n1411), .dout(n1496));
    jnot g0371(.din(n1496), .dout(n1499));
    jor g0372(.dinb(n8425), .dina(n1499), .dout(n1503));
    jor g0373(.dinb(n8423), .dina(n1503), .dout(n1507));
    jand g0374(.dinb(n1488), .dina(n1507), .dout(n1511));
    jand g0375(.dinb(n1379), .dina(n1511), .dout(n1515));
    jand g0376(.dinb(n8564), .dina(n365), .dout(n1519));
    jand g0377(.dinb(n8543), .dina(n376), .dout(n1523));
    jor g0378(.dinb(n8545), .dina(n1523), .dout(n1527));
    jor g0379(.dinb(n8537), .dina(n1527), .dout(n1531));
    jand g0380(.dinb(n11413), .dina(n1531), .dout(n1535));
    jand g0381(.dinb(n8524), .dina(n1264), .dout(n1539));
    jor g0382(.dinb(n1275), .dina(n1539), .dout(n1543));
    jor g0383(.dinb(n1535), .dina(n1543), .dout(n1547));
    jand g0384(.dinb(n9178), .dina(n1547), .dout(n1551));
    jand g0385(.dinb(n8662), .dina(n819), .dout(n1555));
    jnot g0386(.din(n1555), .dout(n1558));
    jor g0387(.dinb(n512), .dina(n1558), .dout(n1562));
    jor g0388(.dinb(n9847), .dina(n91), .dout(n1566));
    jnot g0389(.din(G150), .dout(n1569));
    jand g0390(.dinb(n216), .dina(n350), .dout(n1573));
    jnot g0391(.din(n1573), .dout(n1576));
    jor g0392(.dinb(n8591), .dina(n1576), .dout(n1580));
    jand g0393(.dinb(n216), .dina(n11452), .dout(n1584));
    jand g0394(.dinb(n9862), .dina(n1584), .dout(n1588));
    jnot g0395(.din(n1588), .dout(n1591));
    jand g0396(.dinb(n1580), .dina(n1591), .dout(n1595));
    jand g0397(.dinb(n8585), .dina(n1595), .dout(n1599));
    jor g0398(.dinb(n11119), .dina(n1599), .dout(n1603));
    jand g0399(.dinb(n8629), .dina(n493), .dout(n1607));
    jnot g0400(.din(n1607), .dout(n1610));
    jand g0401(.dinb(n1603), .dina(n8579), .dout(n1614));
    jand g0402(.dinb(n8573), .dina(n1614), .dout(n1618));
    jnot g0403(.din(n1547), .dout(n1621));
    jand g0404(.dinb(n10306), .dina(n1621), .dout(n1625));
    jor g0405(.dinb(n1618), .dina(n1625), .dout(n1629));
    jor g0406(.dinb(n8501), .dina(n1629), .dout(n1633));
    jnot g0407(.din(n1618), .dout(n1636));
    jand g0408(.dinb(n8905), .dina(n1621), .dout(n1640));
    jand g0409(.dinb(n9040), .dina(n1547), .dout(n1644));
    jor g0410(.dinb(n1640), .dina(n8516), .dout(n1648));
    jor g0411(.dinb(n1636), .dina(n1648), .dout(n1652));
    jand g0412(.dinb(n1633), .dina(n1652), .dout(n1656));
    jand g0413(.dinb(n8518), .dina(n365), .dout(n1660));
    jand g0414(.dinb(n8564), .dina(n376), .dout(n1664));
    jor g0415(.dinb(n9905), .dina(n1664), .dout(n1668));
    jor g0416(.dinb(n8465), .dina(n1668), .dout(n1672));
    jand g0417(.dinb(n11407), .dina(n1672), .dout(n1676));
    jand g0418(.dinb(n9949), .dina(n1264), .dout(n1680));
    jor g0419(.dinb(n1275), .dina(n1680), .dout(n1684));
    jor g0420(.dinb(n1676), .dina(n1684), .dout(n1688));
    jand g0421(.dinb(n9160), .dina(n1688), .dout(n1692));
    jand g0422(.dinb(n9859), .dina(n819), .dout(n1696));
    jnot g0423(.din(n1696), .dout(n1699));
    jor g0424(.dinb(n512), .dina(n1699), .dout(n1703));
    jor g0425(.dinb(n216), .dina(n310), .dout(n1707));
    jand g0426(.dinb(n8888), .dina(n1573), .dout(n1711));
    jand g0427(.dinb(n11131), .dina(n1584), .dout(n1715));
    jor g0428(.dinb(n1711), .dina(n1715), .dout(n1719));
    jnot g0429(.din(n1719), .dout(n1722));
    jand g0430(.dinb(n8489), .dina(n1722), .dout(n1726));
    jor g0431(.dinb(n11113), .dina(n1726), .dout(n1730));
    jand g0432(.dinb(n8623), .dina(n493), .dout(n1734));
    jnot g0433(.din(n1734), .dout(n1737));
    jand g0434(.dinb(n1730), .dina(n8480), .dout(n1741));
    jand g0435(.dinb(n8474), .dina(n1741), .dout(n1745));
    jnot g0436(.din(n1688), .dout(n1748));
    jand g0437(.dinb(n10303), .dina(n1748), .dout(n1752));
    jor g0438(.dinb(n1745), .dina(n1752), .dout(n1756));
    jor g0439(.dinb(n8453), .dina(n1756), .dout(n1760));
    jnot g0440(.din(n1745), .dout(n1763));
    jand g0441(.dinb(n8890), .dina(n1748), .dout(n1767));
    jand g0442(.dinb(n9019), .dina(n1688), .dout(n1771));
    jor g0443(.dinb(n1767), .dina(n8462), .dout(n1775));
    jor g0444(.dinb(n1763), .dina(n1775), .dout(n1779));
    jand g0445(.dinb(n1760), .dina(n1779), .dout(n1783));
    jand g0446(.dinb(n1656), .dina(n1783), .dout(n1787));
    jand g0447(.dinb(n1515), .dina(n1787), .dout(n1791));
    jand g0448(.dinb(n10255), .dina(n1791), .dout(n1795));
    jor g0449(.dinb(n10966), .dina(n1156), .dout(n1799));
    jor g0450(.dinb(n11515), .dina(n1120), .dout(n1803));
    jand g0451(.dinb(n1799), .dina(n1803), .dout(n1807));
    jand g0452(.dinb(n1204), .dina(n1807), .dout(n1811));
    jor g0453(.dinb(n11557), .dina(n987), .dout(n1815));
    jor g0454(.dinb(n10966), .dina(n895), .dout(n1819));
    jand g0455(.dinb(n1018), .dina(n1819), .dout(n1823));
    jand g0456(.dinb(n9974), .dina(n1823), .dout(n1827));
    jand g0457(.dinb(n1827), .dina(n1220), .dout(n1831));
    jor g0458(.dinb(n9976), .dina(n1831), .dout(n1835));
    jand g0459(.dinb(n859), .dina(n1835), .dout(n1839));
    jnot g0460(.din(n601), .dout(n1842));
    jand g0461(.dinb(n11536), .dina(n731), .dout(n1846));
    jand g0462(.dinb(n10966), .dina(n683), .dout(n1850));
    jor g0463(.dinb(n1846), .dina(n1850), .dout(n1854));
    jand g0464(.dinb(n1854), .dina(n10576), .dout(n1858));
    jand g0465(.dinb(n620), .dina(n1858), .dout(n1862));
    jor g0466(.dinb(n9970), .dina(n1862), .dout(n1866));
    jor g0467(.dinb(n1839), .dina(n9968), .dout(n1870));
    jand g0468(.dinb(n1791), .dina(n1870), .dout(n1874));
    jnot g0469(.din(n1633), .dout(n1877));
    jnot g0470(.din(n1760), .dout(n1880));
    jor g0471(.dinb(n1350), .dina(n1485), .dout(n1884));
    jand g0472(.dinb(n1507), .dina(n1884), .dout(n1888));
    jor g0473(.dinb(n1880), .dina(n1888), .dout(n1892));
    jand g0474(.dinb(n8455), .dina(n1892), .dout(n1896));
    jor g0475(.dinb(n8491), .dina(n1896), .dout(n1900));
    jand g0476(.dinb(n8503), .dina(n1900), .dout(n1904));
    jor g0477(.dinb(n6437), .dina(n1904), .dout(n1908));
    jand g0478(.dinb(n11461), .dina(n216), .dout(n1912));
    jand g0479(.dinb(n219), .dina(n10192), .dout(n1916));
    jand g0480(.dinb(n1912), .dina(n1916), .dout(n1920));
    jand g0481(.dinb(n10246), .dina(n1920), .dout(n1924));
    jnot g0482(.din(n1924), .dout(n1927));
    jand g0483(.dinb(n1811), .dina(n8134), .dout(n1931));
    jand g0484(.dinb(n1827), .dina(n8125), .dout(n1935));
    jand g0485(.dinb(n1204), .dina(n10102), .dout(n1939));
    jnot g0486(.din(n1939), .dout(n1942));
    jand g0487(.dinb(n1224), .dina(n1942), .dout(n1946));
    jand g0488(.dinb(n9979), .dina(n1939), .dout(n1950));
    jor g0489(.dinb(n1946), .dina(n7781), .dout(n1954));
    jand g0490(.dinb(n7787), .dina(n1954), .dout(n1958));
    jor g0491(.dinb(n7526), .dina(n1958), .dout(n1962));
    jnot g0492(.din(n1954), .dout(n1965));
    jnot g0493(.din(G330), .dout(n1968));
    jnot g0494(.din(n1034), .dout(n1971));
    jor g0495(.dinb(n952), .dina(n10034), .dout(n1975));
    jnot g0496(.din(n1975), .dout(n1978));
    jor g0497(.dinb(n1971), .dina(n8117), .dout(n1982));
    jor g0498(.dinb(n999), .dina(n8119), .dout(n1986));
    jand g0499(.dinb(n1982), .dina(n8108), .dout(n1990));
    jor g0500(.dinb(n8180), .dina(n1990), .dout(n1994));
    jor g0501(.dinb(n7750), .dina(n1994), .dout(n1998));
    jnot g0502(.din(n1998), .dout(n2001));
    jor g0503(.dinb(n7513), .dina(n2001), .dout(n2005));
    jand g0504(.dinb(n1870), .dina(n10000), .dout(n2009));
    jor g0505(.dinb(n1232), .dina(n10075), .dout(n2013));
    jand g0506(.dinb(n10879), .dina(n1120), .dout(n2017));
    jand g0507(.dinb(n10381), .dina(n2017), .dout(n2021));
    jand g0508(.dinb(n10036), .dina(n2021), .dout(n2025));
    jand g0509(.dinb(n10906), .dina(n895), .dout(n2029));
    jand g0510(.dinb(n731), .dina(n1156), .dout(n2033));
    jand g0511(.dinb(n11212), .dina(n2033), .dout(n2037));
    jand g0512(.dinb(n9995), .dina(n2037), .dout(n2041));
    jor g0513(.dinb(n9997), .dina(n2041), .dout(n2045));
    jor g0514(.dinb(n9992), .dina(n2045), .dout(n2049));
    jand g0515(.dinb(n10039), .dina(n2049), .dout(n2053));
    jand g0516(.dinb(n2013), .dina(n9989), .dout(n2057));
    jor g0517(.dinb(n2009), .dina(n2057), .dout(n2061));
    jand g0518(.dinb(n10201), .dina(n2061), .dout(n2065));
    jand g0519(.dinb(n9931), .dina(n252), .dout(n2069));
    jnot g0520(.din(n2069), .dout(n2072));
    jand g0521(.dinb(n10432), .dina(n473), .dout(n2076));
    jand g0522(.dinb(n10600), .dina(n2076), .dout(n2080));
    jand g0523(.dinb(n2072), .dina(n2080), .dout(n2084));
    jand g0524(.dinb(n237), .dina(n2069), .dout(n2088));
    jor g0525(.dinb(n2084), .dina(n6470), .dout(n2092));
    jor g0526(.dinb(n2065), .dina(n6467), .dout(n2096));
    jand g0527(.dinb(n8180), .dina(n1990), .dout(n2100));
    jnot g0528(.din(n2100), .dout(n2103));
    jand g0529(.dinb(n11260), .dina(n1912), .dout(n2107));
    jor g0530(.dinb(n10195), .dina(n2107), .dout(n2111));
    jnot g0531(.din(n2111), .dout(n2114));
    jand g0532(.dinb(n2072), .dina(n2114), .dout(n2118));
    jnot g0533(.din(n2118), .dout(n2121));
    jand g0534(.dinb(n1994), .dina(n8719), .dout(n2125));
    jand g0535(.dinb(n2103), .dina(n2125), .dout(n2129));
    jand g0536(.dinb(n11245), .dina(n1573), .dout(n2133));
    jand g0537(.dinb(n1990), .dina(n8005), .dout(n2137));
    jnot g0538(.din(n2137), .dout(n2140));
    jand g0539(.dinb(n9892), .dina(n343), .dout(n2144));
    jor g0540(.dinb(n226), .dina(n2144), .dout(n2148));
    jand g0541(.dinb(G20), .dina(G179), .dout(n2152));
    jnot g0542(.din(n2152), .dout(n2155));
    jand g0543(.dinb(G20), .dina(G200), .dout(n2159));
    jand g0544(.dinb(n2155), .dina(n9016), .dout(n2163));
    jand g0545(.dinb(n10864), .dina(n2163), .dout(n2167));
    jand g0546(.dinb(n10522), .dina(n2167), .dout(n2171));
    jand g0547(.dinb(n11128), .dina(n1360), .dout(n2175));
    jnot g0548(.din(n2175), .dout(n2178));
    jor g0549(.dinb(n2152), .dina(n2159), .dout(n2182));
    jnot g0550(.din(n2182), .dout(n2185));
    jand g0551(.dinb(n2178), .dina(n2185), .dout(n2189));
    jand g0552(.dinb(n10273), .dina(n2189), .dout(n2193));
    jnot g0553(.din(G200), .dout(n2196));
    jand g0554(.dinb(n2196), .dina(n2152), .dout(n2200));
    jand g0555(.dinb(n10858), .dina(n2200), .dout(n2204));
    jand g0556(.dinb(n7946), .dina(n2204), .dout(n2208));
    jor g0557(.dinb(n2193), .dina(n7934), .dout(n2212));
    jor g0558(.dinb(n7931), .dina(n2212), .dout(n2216));
    jand g0559(.dinb(n9061), .dina(n2185), .dout(n2220));
    jand g0560(.dinb(n7913), .dina(n2220), .dout(n2224));
    jor g0561(.dinb(n7924), .dina(n2224), .dout(n2228));
    jand g0562(.dinb(n9067), .dina(n2163), .dout(n2232));
    jand g0563(.dinb(n10762), .dina(n2232), .dout(n2236));
    jand g0564(.dinb(n9064), .dina(n2200), .dout(n2240));
    jand g0565(.dinb(n8816), .dina(n2240), .dout(n2244));
    jor g0566(.dinb(n2236), .dina(n7901), .dout(n2248));
    jand g0567(.dinb(n10819), .dina(n2152), .dout(n2252));
    jand g0568(.dinb(n10858), .dina(n2252), .dout(n2256));
    jand g0569(.dinb(n7898), .dina(n2256), .dout(n2260));
    jand g0570(.dinb(n9805), .dina(n2252), .dout(n2264));
    jand g0571(.dinb(n7886), .dina(n2264), .dout(n2268));
    jor g0572(.dinb(n2260), .dina(n2268), .dout(n2272));
    jor g0573(.dinb(n2248), .dina(n7874), .dout(n2276));
    jor g0574(.dinb(n7871), .dina(n2276), .dout(n2280));
    jor g0575(.dinb(n7868), .dina(n2280), .dout(n2284));
    jand g0576(.dinb(n8869), .dina(n2220), .dout(n2288));
    jand g0577(.dinb(n8656), .dina(n2256), .dout(n2292));
    jand g0578(.dinb(n8839), .dina(n2264), .dout(n2296));
    jor g0579(.dinb(n2292), .dina(n2296), .dout(n2300));
    jor g0580(.dinb(n2288), .dina(n2300), .dout(n2304));
    jnot g0581(.din(n2304), .dout(n2307));
    jand g0582(.dinb(n9919), .dina(n2167), .dout(n2311));
    jnot g0583(.din(n2311), .dout(n2314));
    jand g0584(.dinb(n7915), .dina(n2314), .dout(n2318));
    jand g0585(.dinb(n10324), .dina(n2232), .dout(n2322));
    jand g0586(.dinb(n8551), .dina(n2240), .dout(n2326));
    jor g0587(.dinb(n2322), .dina(n7865), .dout(n2330));
    jand g0588(.dinb(n9883), .dina(n2204), .dout(n2334));
    jand g0589(.dinb(n10483), .dina(n2189), .dout(n2338));
    jor g0590(.dinb(n7862), .dina(n2338), .dout(n2342));
    jor g0591(.dinb(n2330), .dina(n2342), .dout(n2346));
    jnot g0592(.din(n2346), .dout(n2349));
    jand g0593(.dinb(n7859), .dina(n2349), .dout(n2353));
    jand g0594(.dinb(n7856), .dina(n2353), .dout(n2357));
    jnot g0595(.din(n2357), .dout(n2360));
    jand g0596(.dinb(n7850), .dina(n2360), .dout(n2364));
    jor g0597(.dinb(n7948), .dina(n2364), .dout(n2368));
    jnot g0598(.din(n2133), .dout(n2371));
    jand g0599(.dinb(n2371), .dina(n8326), .dout(n2375));
    jnot g0600(.din(n2375), .dout(n2378));
    jand g0601(.dinb(n11278), .dina(n321), .dout(n2382));
    jand g0602(.dinb(n11251), .dina(n237), .dout(n2386));
    jand g0603(.dinb(n8962), .dina(n252), .dout(n2390));
    jnot g0604(.din(n2390), .dout(n2393));
    jor g0605(.dinb(n2386), .dina(n2393), .dout(n2397));
    jor g0606(.dinb(n7823), .dina(n2397), .dout(n2401));
    jand g0607(.dinb(n10447), .dina(n255), .dout(n2405));
    jand g0608(.dinb(n9364), .dina(n252), .dout(n2409));
    jand g0609(.dinb(n115), .dina(n7817), .dout(n2413));
    jor g0610(.dinb(n7814), .dina(n2413), .dout(n2417));
    jnot g0611(.din(n2417), .dout(n2420));
    jand g0612(.dinb(n7811), .dina(n2420), .dout(n2424));
    jor g0613(.dinb(n7828), .dina(n2424), .dout(n2428));
    jand g0614(.dinb(n8743), .dina(n2428), .dout(n2432));
    jand g0615(.dinb(n2368), .dina(n7808), .dout(n2436));
    jand g0616(.dinb(n2140), .dina(n7802), .dout(n2440));
    jor g0617(.dinb(n2129), .dina(n2440), .dout(n2444));
    jnot g0618(.din(n2057), .dout(n2447));
    jnot g0619(.din(n1338), .dout(n2450));
    jor g0620(.dinb(n2450), .dina(n10024), .dout(n2454));
    jand g0621(.dinb(n1379), .dina(n9775), .dout(n2458));
    jor g0622(.dinb(n1353), .dina(n9779), .dout(n2462));
    jnot g0623(.din(n2462), .dout(n2465));
    jor g0624(.dinb(n2458), .dina(n2465), .dout(n2469));
    jxor g0625(.dinb(n2009), .dina(n9769), .dout(n2473));
    jnot g0626(.din(n2473), .dout(n2476));
    jand g0627(.dinb(n9764), .dina(n2476), .dout(n2480));
    jor g0628(.dinb(n9379), .dina(n3603), .dout(n2484));
    jor g0629(.dinb(n2480), .dina(n9371), .dout(n2488));
    jnot g0630(.din(n2469), .dout(n2491));
    jand g0631(.dinb(n9235), .dina(n2491), .dout(n2495));
    jnot g0632(.din(n2495), .dout(n2498));
    jand g0633(.dinb(n9073), .dina(n2220), .dout(n2502));
    jand g0634(.dinb(n9013), .dina(n2189), .dout(n2506));
    jand g0635(.dinb(n8983), .dina(n2264), .dout(n2510));
    jor g0636(.dinb(n2506), .dina(n8981), .dout(n2514));
    jor g0637(.dinb(n8978), .dina(n2514), .dout(n2518));
    jand g0638(.dinb(n8929), .dina(n2167), .dout(n2522));
    jor g0639(.dinb(n8950), .dina(n2522), .dout(n2526));
    jand g0640(.dinb(n8866), .dina(n2240), .dout(n2530));
    jand g0641(.dinb(n8864), .dina(n2204), .dout(n2534));
    jor g0642(.dinb(n2530), .dina(n2534), .dout(n2538));
    jand g0643(.dinb(n8855), .dina(n2256), .dout(n2542));
    jand g0644(.dinb(n8830), .dina(n2232), .dout(n2546));
    jor g0645(.dinb(n8828), .dina(n2546), .dout(n2550));
    jor g0646(.dinb(n8825), .dina(n2550), .dout(n2554));
    jor g0647(.dinb(n8822), .dina(n2554), .dout(n2558));
    jor g0648(.dinb(n8819), .dina(n2558), .dout(n2562));
    jand g0649(.dinb(n8806), .dina(n2220), .dout(n2566));
    jand g0650(.dinb(n10321), .dina(n2167), .dout(n2570));
    jand g0651(.dinb(n10753), .dina(n2264), .dout(n2574));
    jor g0652(.dinb(n2570), .dina(n8804), .dout(n2578));
    jor g0653(.dinb(n8801), .dina(n2578), .dout(n2582));
    jnot g0654(.din(n2582), .dout(n2585));
    jand g0655(.dinb(n9907), .dina(n2232), .dout(n2589));
    jnot g0656(.din(n2589), .dout(n2592));
    jand g0657(.dinb(n8794), .dina(n2592), .dout(n2596));
    jand g0658(.dinb(n8785), .dina(n2240), .dout(n2600));
    jand g0659(.dinb(n10294), .dina(n2204), .dout(n2604));
    jor g0660(.dinb(n2600), .dina(n2604), .dout(n2608));
    jand g0661(.dinb(n10513), .dina(n2256), .dout(n2612));
    jor g0662(.dinb(n2338), .dina(n8771), .dout(n2616));
    jor g0663(.dinb(n8768), .dina(n2616), .dout(n2620));
    jnot g0664(.din(n2620), .dout(n2623));
    jand g0665(.dinb(n8765), .dina(n2623), .dout(n2627));
    jand g0666(.dinb(n8762), .dina(n2627), .dout(n2631));
    jnot g0667(.din(n2631), .dout(n2634));
    jand g0668(.dinb(n8759), .dina(n2634), .dout(n2638));
    jor g0669(.dinb(n9112), .dina(n2638), .dout(n2642));
    jand g0670(.dinb(n1433), .dina(n2148), .dout(n2646));
    jand g0671(.dinb(n9829), .dina(n2646), .dout(n2650));
    jor g0672(.dinb(n2121), .dina(n8717), .dout(n2654));
    jnot g0673(.din(n2654), .dout(n2657));
    jand g0674(.dinb(n2642), .dina(n8711), .dout(n2661));
    jand g0675(.dinb(n2498), .dina(n8699), .dout(n2665));
    jnot g0676(.din(n2665), .dout(n2668));
    jand g0677(.dinb(n2488), .dina(n2668), .dout(n2672));
    jnot g0678(.din(n2672), .dout(n2675));
    jnot g0679(.din(n1920), .dout(n2678));
    jand g0680(.dinb(n1880), .dina(n7163), .dout(n2682));
    jand g0681(.dinb(n1763), .dina(n10168), .dout(n2686));
    jnot g0682(.din(n2686), .dout(n2689));
    jand g0683(.dinb(n1783), .dina(n2689), .dout(n2693));
    jand g0684(.dinb(n1880), .dina(n7276), .dout(n2697));
    jor g0685(.dinb(n2693), .dina(n2697), .dout(n2701));
    jand g0686(.dinb(n2009), .dina(n9766), .dout(n2705));
    jand g0687(.dinb(n1473), .dina(n10117), .dout(n2709));
    jnot g0688(.din(n2709), .dout(n2712));
    jand g0689(.dinb(n1511), .dina(n8369), .dout(n2716));
    jand g0690(.dinb(n1485), .dina(n8371), .dout(n2720));
    jor g0691(.dinb(n2716), .dina(n8363), .dout(n2724));
    jand g0692(.dinb(n2705), .dina(n7291), .dout(n2728));
    jor g0693(.dinb(n8407), .dina(n2724), .dout(n2732));
    jand g0694(.dinb(n1884), .dina(n8389), .dout(n2736));
    jand g0695(.dinb(n2732), .dina(n7289), .dout(n2740));
    jor g0696(.dinb(n2728), .dina(n7280), .dout(n2744));
    jand g0697(.dinb(n7132), .dina(n2744), .dout(n2748));
    jor g0698(.dinb(n7130), .dina(n2748), .dout(n2752));
    jnot g0699(.din(n2752), .dout(n2755));
    jand g0700(.dinb(n6598), .dina(n2009), .dout(n2759));
    jor g0701(.dinb(n1904), .dina(n2759), .dout(n2763));
    jand g0702(.dinb(n2469), .dina(n2724), .dout(n2767));
    jand g0703(.dinb(n7264), .dina(n2767), .dout(n2771));
    jxor g0704(.dinb(n8398), .dina(n2771), .dout(n2775));
    jand g0705(.dinb(n9982), .dina(n2775), .dout(n2779));
    jxor g0706(.dinb(n6596), .dina(n2779), .dout(n2783));
    jnot g0707(.din(n2783), .dout(n2786));
    jor g0708(.dinb(n2755), .dina(n6590), .dout(n2790));
    jor g0709(.dinb(n2752), .dina(n6592), .dout(n2794));
    jnot g0710(.din(n248), .dout(n2797));
    jand g0711(.dinb(n230), .dina(n2797), .dout(n2801));
    jand g0712(.dinb(n2794), .dina(n6581), .dout(n2805));
    jand g0713(.dinb(n2790), .dina(n2805), .dout(n2809));
    jand g0714(.dinb(G50), .dina(G77), .dout(n2813));
    jand g0715(.dinb(n310), .dina(n2813), .dout(n2817));
    jand g0716(.dinb(n77), .dina(n11152), .dout(n2821));
    jor g0717(.dinb(n2817), .dina(n2821), .dout(n2825));
    jand g0718(.dinb(n9760), .dina(n2825), .dout(n2829));
    jnot g0719(.din(n767), .dout(n2832));
    jand g0720(.dinb(n11347), .dina(n347), .dout(n2836));
    jand g0721(.dinb(n2832), .dina(n6530), .dout(n2840));
    jor g0722(.dinb(n6524), .dina(n2840), .dout(n2844));
    jor g0723(.dinb(n2809), .dina(n6521), .dout(n2848));
    jand g0724(.dinb(n604), .dina(n10117), .dout(n2852));
    jnot g0725(.din(n2852), .dout(n2855));
    jand g0726(.dinb(n624), .dina(n7622), .dout(n2859));
    jand g0727(.dinb(n1842), .dina(n7624), .dout(n2863));
    jor g0728(.dinb(n2859), .dina(n7619), .dout(n2867));
    jnot g0729(.din(n2867), .dout(n2870));
    jand g0730(.dinb(n7972), .dina(n2870), .dout(n2874));
    jnot g0731(.din(n2874), .dout(n2877));
    jand g0732(.dinb(n7876), .dina(n2220), .dout(n2881));
    jand g0733(.dinb(n7603), .dina(n2189), .dout(n2885));
    jand g0734(.dinb(n10294), .dina(n2264), .dout(n2889));
    jor g0735(.dinb(n2885), .dina(n7601), .dout(n2893));
    jor g0736(.dinb(n7598), .dina(n2893), .dout(n2897));
    jand g0737(.dinb(n8776), .dina(n2167), .dout(n2901));
    jor g0738(.dinb(n9352), .dina(n2901), .dout(n2905));
    jand g0739(.dinb(n10783), .dina(n2240), .dout(n2909));
    jand g0740(.dinb(n10534), .dina(n2204), .dout(n2913));
    jor g0741(.dinb(n2909), .dina(n2913), .dout(n2917));
    jand g0742(.dinb(n8816), .dina(n2256), .dout(n2921));
    jand g0743(.dinb(n10474), .dina(n2232), .dout(n2925));
    jor g0744(.dinb(n7595), .dina(n2925), .dout(n2929));
    jor g0745(.dinb(n7592), .dina(n2929), .dout(n2933));
    jor g0746(.dinb(n7589), .dina(n2933), .dout(n2937));
    jor g0747(.dinb(n7586), .dina(n2937), .dout(n2941));
    jand g0748(.dinb(n8845), .dina(n2220), .dout(n2945));
    jnot g0749(.din(n2945), .dout(n2948));
    jand g0750(.dinb(n7690), .dina(n2189), .dout(n2952));
    jnot g0751(.din(n2952), .dout(n2955));
    jand g0752(.dinb(n8251), .dina(n2232), .dout(n2959));
    jnot g0753(.din(n2959), .dout(n2962));
    jand g0754(.dinb(n2955), .dina(n2962), .dout(n2966));
    jand g0755(.dinb(n7583), .dina(n2966), .dout(n2970));
    jand g0756(.dinb(n8881), .dina(n2264), .dout(n2974));
    jor g0757(.dinb(n8968), .dina(n2974), .dout(n2978));
    jand g0758(.dinb(n8864), .dina(n2256), .dout(n2982));
    jand g0759(.dinb(n9001), .dina(n2204), .dout(n2986));
    jor g0760(.dinb(n2982), .dina(n2986), .dout(n2990));
    jand g0761(.dinb(n8920), .dina(n2240), .dout(n2994));
    jand g0762(.dinb(n9010), .dina(n2167), .dout(n2998));
    jor g0763(.dinb(n7580), .dina(n2998), .dout(n3002));
    jor g0764(.dinb(n7577), .dina(n3002), .dout(n3006));
    jor g0765(.dinb(n7574), .dina(n3006), .dout(n3010));
    jnot g0766(.din(n3010), .dout(n3013));
    jand g0767(.dinb(n7568), .dina(n3013), .dout(n3017));
    jnot g0768(.din(n3017), .dout(n3020));
    jand g0769(.dinb(n7565), .dina(n3020), .dout(n3024));
    jor g0770(.dinb(n9085), .dina(n3024), .dout(n3028));
    jand g0771(.dinb(n7555), .dina(n2390), .dout(n3032));
    jand g0772(.dinb(n8236), .dina(n255), .dout(n3036));
    jor g0773(.dinb(n2378), .dina(n7553), .dout(n3040));
    jor g0774(.dinb(n7550), .dina(n3040), .dout(n3044));
    jand g0775(.dinb(n9403), .dina(n3044), .dout(n3048));
    jand g0776(.dinb(n3028), .dina(n7544), .dout(n3052));
    jand g0777(.dinb(n2877), .dina(n7532), .dout(n3056));
    jnot g0778(.din(n2061), .dout(n3059));
    jxor g0779(.dinb(n7787), .dina(n1954), .dout(n3063));
    jxor g0780(.dinb(n1994), .dina(n7778), .dout(n3067));
    jnot g0781(.din(n3067), .dout(n3070));
    jand g0782(.dinb(n3059), .dina(n3070), .dout(n3074));
    jnot g0783(.din(n855), .dout(n3077));
    jand g0784(.dinb(n839), .dina(n10117), .dout(n3081));
    jor g0785(.dinb(n3077), .dina(n7505), .dout(n3085));
    jand g0786(.dinb(n1858), .dina(n10129), .dout(n3089));
    jnot g0787(.din(n3089), .dout(n3092));
    jand g0788(.dinb(n3085), .dina(n7496), .dout(n3096));
    jxor g0789(.dinb(n1998), .dina(n7483), .dout(n3100));
    jxor g0790(.dinb(n7507), .dina(n3100), .dout(n3104));
    jand g0791(.dinb(n3074), .dina(n3104), .dout(n3108));
    jor g0792(.dinb(n7759), .dina(n3108), .dout(n3112));
    jand g0793(.dinb(n9712), .dina(n3112), .dout(n3116));
    jor g0794(.dinb(n9529), .dina(n3116), .dout(n3120));
    jand g0795(.dinb(n1858), .dina(n10015), .dout(n3124));
    jnot g0796(.din(n3096), .dout(n3127));
    jand g0797(.dinb(n1962), .dina(n3127), .dout(n3131));
    jor g0798(.dinb(n7481), .dina(n3131), .dout(n3135));
    jor g0799(.dinb(n1998), .dina(n7489), .dout(n3139));
    jxor g0800(.dinb(n7606), .dina(n3139), .dout(n3143));
    jxor g0801(.dinb(n7466), .dina(n3143), .dout(n3147));
    jnot g0802(.din(n3147), .dout(n3150));
    jand g0803(.dinb(n3120), .dina(n7463), .dout(n3154));
    jor g0804(.dinb(n7457), .dina(n3154), .dout(n3158));
    jand g0805(.dinb(n2061), .dina(n3067), .dout(n3162));
    jor g0806(.dinb(n9580), .dina(n3074), .dout(n3166));
    jor g0807(.dinb(n7757), .dina(n3166), .dout(n3170));
    jor g0808(.dinb(n9415), .dina(n3067), .dout(n3174));
    jand g0809(.dinb(n1965), .dina(n8071), .dout(n3178));
    jand g0810(.dinb(n7888), .dina(n2220), .dout(n3182));
    jand g0811(.dinb(n7747), .dina(n2189), .dout(n3186));
    jand g0812(.dinb(n7886), .dina(n2204), .dout(n3190));
    jor g0813(.dinb(n3186), .dina(n7742), .dout(n3194));
    jor g0814(.dinb(n7739), .dina(n3194), .dout(n3198));
    jand g0815(.dinb(n8773), .dina(n2167), .dout(n3202));
    jor g0816(.dinb(n9352), .dina(n3202), .dout(n3206));
    jand g0817(.dinb(n7735), .dina(n2232), .dout(n3210));
    jand g0818(.dinb(n10534), .dina(n2240), .dout(n3214));
    jor g0819(.dinb(n3210), .dina(n7730), .dout(n3218));
    jand g0820(.dinb(n7946), .dina(n2256), .dout(n3222));
    jand g0821(.dinb(n8816), .dina(n2264), .dout(n3226));
    jor g0822(.dinb(n3222), .dina(n3226), .dout(n3230));
    jor g0823(.dinb(n3218), .dina(n7727), .dout(n3234));
    jor g0824(.dinb(n7724), .dina(n3234), .dout(n3238));
    jor g0825(.dinb(n7721), .dina(n3238), .dout(n3242));
    jand g0826(.dinb(n8233), .dina(n2189), .dout(n3246));
    jand g0827(.dinb(n7714), .dina(n2264), .dout(n3250));
    jor g0828(.dinb(n2925), .dina(n7706), .dout(n3254));
    jor g0829(.dinb(n8230), .dina(n3254), .dout(n3258));
    jand g0830(.dinb(n7702), .dina(n2220), .dout(n3262));
    jor g0831(.dinb(n8791), .dina(n3262), .dout(n3266));
    jand g0832(.dinb(n8881), .dina(n2256), .dout(n3270));
    jand g0833(.dinb(n7681), .dina(n2240), .dout(n3274));
    jor g0834(.dinb(n3270), .dina(n3274), .dout(n3278));
    jand g0835(.dinb(n8941), .dina(n2204), .dout(n3282));
    jand g0836(.dinb(n8239), .dina(n2167), .dout(n3286));
    jor g0837(.dinb(n7676), .dina(n3286), .dout(n3290));
    jor g0838(.dinb(n7673), .dina(n3290), .dout(n3294));
    jor g0839(.dinb(n7670), .dina(n3294), .dout(n3298));
    jor g0840(.dinb(n7667), .dina(n3298), .dout(n3302));
    jand g0841(.dinb(n3242), .dina(n3302), .dout(n3306));
    jor g0842(.dinb(n9139), .dina(n3306), .dout(n3310));
    jand g0843(.dinb(n11269), .dina(n302), .dout(n3314));
    jand g0844(.dinb(G68), .dina(G77), .dout(n3318));
    jnot g0845(.din(n3318), .dout(n3321));
    jand g0846(.dinb(n399), .dina(n9880), .dout(n3325));
    jand g0847(.dinb(n7657), .dina(n3325), .dout(n3329));
    jand g0848(.dinb(n7655), .dina(n3329), .dout(n3333));
    jand g0849(.dinb(n2076), .dina(n3333), .dout(n3337));
    jor g0850(.dinb(n2393), .dina(n3337), .dout(n3341));
    jor g0851(.dinb(n7652), .dina(n3341), .dout(n3345));
    jand g0852(.dinb(n11026), .dina(n255), .dout(n3349));
    jnot g0853(.din(n2076), .dout(n3352));
    jand g0854(.dinb(n3352), .dina(n7817), .dout(n3356));
    jor g0855(.dinb(n7646), .dina(n3356), .dout(n3360));
    jnot g0856(.din(n3360), .dout(n3363));
    jand g0857(.dinb(n7643), .dina(n3363), .dout(n3367));
    jor g0858(.dinb(n7837), .dina(n3367), .dout(n3371));
    jand g0859(.dinb(n9373), .dina(n3371), .dout(n3375));
    jand g0860(.dinb(n3310), .dina(n3375), .dout(n3379));
    jnot g0861(.din(n3379), .dout(n3382));
    jor g0862(.dinb(n3178), .dina(n7640), .dout(n3386));
    jand g0863(.dinb(n3174), .dina(n7634), .dout(n3390));
    jand g0864(.dinb(n3170), .dina(n7631), .dout(n3394));
    jnot g0865(.din(n3394), .dout(n3397));
    jnot g0866(.din(n3074), .dout(n3400));
    jnot g0867(.din(n3104), .dout(n3403));
    jand g0868(.dinb(n3400), .dina(n3403), .dout(n3407));
    jor g0869(.dinb(n7774), .dina(n3108), .dout(n3411));
    jor g0870(.dinb(n3407), .dina(n3411), .dout(n3415));
    jor g0871(.dinb(n9448), .dina(n3403), .dout(n3419));
    jand g0872(.dinb(n8038), .dina(n3096), .dout(n3423));
    jnot g0873(.din(n3423), .dout(n3426));
    jand g0874(.dinb(n7732), .dina(n2189), .dout(n3430));
    jand g0875(.dinb(n7744), .dina(n2167), .dout(n3434));
    jand g0876(.dinb(n10534), .dina(n2264), .dout(n3438));
    jor g0877(.dinb(n3434), .dina(n7430), .dout(n3442));
    jor g0878(.dinb(n7427), .dina(n3442), .dout(n3446));
    jand g0879(.dinb(n7936), .dina(n2220), .dout(n3450));
    jor g0880(.dinb(n9352), .dina(n3450), .dout(n3454));
    jand g0881(.dinb(n10285), .dina(n2240), .dout(n3458));
    jand g0882(.dinb(n8816), .dina(n2204), .dout(n3462));
    jor g0883(.dinb(n3458), .dina(n3462), .dout(n3466));
    jand g0884(.dinb(n7886), .dina(n2256), .dout(n3470));
    jor g0885(.dinb(n2322), .dina(n7424), .dout(n3474));
    jor g0886(.dinb(n7421), .dina(n3474), .dout(n3478));
    jor g0887(.dinb(n7418), .dina(n3478), .dout(n3482));
    jor g0888(.dinb(n7415), .dina(n3482), .dout(n3486));
    jand g0889(.dinb(n10639), .dina(n2189), .dout(n3490));
    jand g0890(.dinb(n11140), .dina(n2167), .dout(n3494));
    jand g0891(.dinb(n8941), .dina(n2264), .dout(n3498));
    jor g0892(.dinb(n3494), .dina(n7409), .dout(n3502));
    jor g0893(.dinb(n7411), .dina(n3502), .dout(n3506));
    jand g0894(.dinb(n7381), .dina(n2220), .dout(n3510));
    jor g0895(.dinb(n7396), .dina(n3510), .dout(n3514));
    jand g0896(.dinb(n7708), .dina(n2240), .dout(n3518));
    jand g0897(.dinb(n8881), .dina(n2204), .dout(n3522));
    jor g0898(.dinb(n3518), .dina(n3522), .dout(n3526));
    jand g0899(.dinb(n9001), .dina(n2256), .dout(n3530));
    jor g0900(.dinb(n2589), .dina(n7376), .dout(n3534));
    jor g0901(.dinb(n7373), .dina(n3534), .dout(n3538));
    jor g0902(.dinb(n7370), .dina(n3538), .dout(n3542));
    jor g0903(.dinb(n7367), .dina(n3542), .dout(n3546));
    jand g0904(.dinb(n3486), .dina(n3546), .dout(n3550));
    jor g0905(.dinb(n9139), .dina(n3550), .dout(n3554));
    jand g0906(.dinb(n7361), .dina(n2390), .dout(n3558));
    jand g0907(.dinb(n7357), .dina(n255), .dout(n3562));
    jor g0908(.dinb(n2378), .dina(n7355), .dout(n3566));
    jor g0909(.dinb(n7352), .dina(n3566), .dout(n3570));
    jand g0910(.dinb(n9409), .dina(n3570), .dout(n3574));
    jand g0911(.dinb(n3554), .dina(n7346), .dout(n3578));
    jand g0912(.dinb(n3426), .dina(n7340), .dout(n3582));
    jnot g0913(.din(n3582), .dout(n3585));
    jand g0914(.dinb(n3419), .dina(n7328), .dout(n3589));
    jand g0915(.dinb(n3415), .dina(n3589), .dout(n3593));
    jnot g0916(.din(n3593), .dout(n3596));
    jnot g0917(.din(n2701), .dout(n3599));
    jand g0918(.dinb(n2057), .dina(n9772), .dout(n3603));
    jand g0919(.dinb(n8353), .dina(n3603), .dout(n3607));
    jxor g0920(.dinb(n7258), .dina(n3607), .dout(n3611));
    jxor g0921(.dinb(n2744), .dina(n3611), .dout(n3615));
    jand g0922(.dinb(n8392), .dina(n2061), .dout(n3619));
    jor g0923(.dinb(n8404), .dina(n3619), .dout(n3623));
    jand g0924(.dinb(n1350), .dina(n10015), .dout(n3627));
    jor g0925(.dinb(n2705), .dina(n8387), .dout(n3631));
    jnot g0926(.din(n2724), .dout(n3634));
    jxor g0927(.dinb(n8350), .dina(n3603), .dout(n3638));
    jxor g0928(.dinb(n3631), .dina(n3638), .dout(n3642));
    jor g0929(.dinb(n3623), .dina(n3642), .dout(n3646));
    jor g0930(.dinb(n3615), .dina(n3646), .dout(n3650));
    jnot g0931(.din(n3650), .dout(n3653));
    jand g0932(.dinb(n3615), .dina(n3646), .dout(n3657));
    jor g0933(.dinb(n7768), .dina(n3657), .dout(n3661));
    jor g0934(.dinb(n3653), .dina(n3661), .dout(n3665));
    jor g0935(.dinb(n9448), .dina(n3615), .dout(n3669));
    jand g0936(.dinb(n9196), .dina(n3599), .dout(n3673));
    jnot g0937(.din(n3673), .dout(n3676));
    jand g0938(.dinb(n7246), .dina(n2220), .dout(n3680));
    jand g0939(.dinb(n8875), .dina(n2189), .dout(n3684));
    jand g0940(.dinb(n8855), .dina(n2264), .dout(n3688));
    jor g0941(.dinb(n3684), .dina(n7244), .dout(n3692));
    jor g0942(.dinb(n7241), .dina(n3692), .dout(n3696));
    jand g0943(.dinb(n8305), .dina(n2167), .dout(n3700));
    jor g0944(.dinb(n7384), .dina(n3700), .dout(n3704));
    jand g0945(.dinb(n8864), .dina(n2240), .dout(n3708));
    jand g0946(.dinb(n9083), .dina(n2204), .dout(n3712));
    jor g0947(.dinb(n3708), .dina(n3712), .dout(n3716));
    jand g0948(.dinb(n8318), .dina(n2256), .dout(n3720));
    jand g0949(.dinb(n7678), .dina(n2232), .dout(n3724));
    jor g0950(.dinb(n7238), .dina(n3724), .dout(n3728));
    jor g0951(.dinb(n7235), .dina(n3728), .dout(n3732));
    jor g0952(.dinb(n7232), .dina(n3732), .dout(n3736));
    jor g0953(.dinb(n7229), .dina(n3736), .dout(n3740));
    jand g0954(.dinb(n8287), .dina(n2220), .dout(n3744));
    jand g0955(.dinb(n11059), .dina(n2264), .dout(n3748));
    jor g0956(.dinb(n3490), .dina(n7226), .dout(n3752));
    jor g0957(.dinb(n7223), .dina(n3752), .dout(n3756));
    jand g0958(.dinb(n10774), .dina(n2256), .dout(n3760));
    jor g0959(.dinb(n8278), .dina(n3760), .dout(n3764));
    jand g0960(.dinb(n11194), .dina(n2240), .dout(n3768));
    jand g0961(.dinb(n11338), .dina(n2204), .dout(n3772));
    jor g0962(.dinb(n3768), .dina(n3772), .dout(n3776));
    jor g0963(.dinb(n2311), .dina(n2546), .dout(n3780));
    jor g0964(.dinb(n7220), .dina(n3780), .dout(n3784));
    jor g0965(.dinb(n7217), .dina(n3784), .dout(n3788));
    jor g0966(.dinb(n7211), .dina(n3788), .dout(n3792));
    jand g0967(.dinb(n3740), .dina(n3792), .dout(n3796));
    jor g0968(.dinb(n9139), .dina(n3796), .dout(n3800));
    jand g0969(.dinb(n8614), .dina(n2646), .dout(n3804));
    jor g0970(.dinb(n2121), .dina(n7208), .dout(n3808));
    jnot g0971(.din(n3808), .dout(n3811));
    jand g0972(.dinb(n3800), .dina(n7202), .dout(n3815));
    jand g0973(.dinb(n3676), .dina(n7196), .dout(n3819));
    jnot g0974(.din(n3819), .dout(n3822));
    jand g0975(.dinb(n3669), .dina(n7181), .dout(n3826));
    jand g0976(.dinb(n3665), .dina(n7178), .dout(n3830));
    jnot g0977(.din(n3830), .dout(n3833));
    jand g0978(.dinb(n7267), .dina(n3607), .dout(n3837));
    jand g0979(.dinb(n1636), .dina(n10147), .dout(n3841));
    jnot g0980(.din(n3841), .dout(n3844));
    jand g0981(.dinb(n1656), .dina(n3844), .dout(n3848));
    jand g0982(.dinb(n1877), .dina(n7111), .dout(n3852));
    jor g0983(.dinb(n3848), .dina(n3852), .dout(n3856));
    jnot g0984(.din(n3856), .dout(n3859));
    jxor g0985(.dinb(n2752), .dina(n7096), .dout(n3863));
    jxor g0986(.dinb(n7094), .dina(n3863), .dout(n3867));
    jor g0987(.dinb(n7432), .dina(n3867), .dout(n3871));
    jnot g0988(.din(n3623), .dout(n3874));
    jand g0989(.dinb(n7085), .dina(n3650), .dout(n3878));
    jor g0990(.dinb(n9619), .dina(n3878), .dout(n3882));
    jor g0991(.dinb(n3867), .dina(n3882), .dout(n3886));
    jand g0992(.dinb(n9313), .dina(n3859), .dout(n3890));
    jnot g0993(.din(n2148), .dout(n3893));
    jand g0994(.dinb(n9083), .dina(n2264), .dout(n3897));
    jand g0995(.dinb(n8318), .dina(n2204), .dout(n3901));
    jand g0996(.dinb(n8855), .dina(n2240), .dout(n3905));
    jor g0997(.dinb(n3901), .dina(n3905), .dout(n3909));
    jor g0998(.dinb(n7082), .dina(n3909), .dout(n3913));
    jnot g0999(.din(n3913), .dout(n3916));
    jand g1000(.dinb(n8302), .dina(n2189), .dout(n3920));
    jnot g1001(.din(n3920), .dout(n3923));
    jand g1002(.dinb(n350), .dina(n353), .dout(n3927));
    jand g1003(.dinb(n3923), .dina(n7079), .dout(n3931));
    jand g1004(.dinb(n7256), .dina(n2256), .dout(n3935));
    jand g1005(.dinb(n7378), .dina(n2167), .dout(n3939));
    jor g1006(.dinb(n7067), .dina(n3939), .dout(n3943));
    jand g1007(.dinb(n7064), .dina(n2220), .dout(n3947));
    jand g1008(.dinb(n8875), .dina(n2232), .dout(n3951));
    jor g1009(.dinb(n3947), .dina(n3951), .dout(n3955));
    jor g1010(.dinb(n3943), .dina(n3955), .dout(n3959));
    jnot g1011(.din(n3959), .dout(n3962));
    jand g1012(.dinb(n7052), .dina(n3962), .dout(n3966));
    jand g1013(.dinb(n7049), .dina(n3966), .dout(n3970));
    jand g1014(.dinb(n11059), .dina(n2204), .dout(n3974));
    jand g1015(.dinb(n9868), .dina(n2232), .dout(n3978));
    jand g1016(.dinb(n11104), .dina(n2240), .dout(n3982));
    jor g1017(.dinb(n3978), .dina(n7043), .dout(n3986));
    jor g1018(.dinb(n7040), .dina(n3986), .dout(n3990));
    jnot g1019(.din(n3990), .dout(n3993));
    jand g1020(.dinb(n11194), .dina(n2264), .dout(n3997));
    jnot g1021(.din(n3997), .dout(n4000));
    jand g1022(.dinb(n11452), .dina(n353), .dout(n4004));
    jand g1023(.dinb(n4000), .dina(n7034), .dout(n4008));
    jand g1024(.dinb(n8263), .dina(n2220), .dout(n4012));
    jor g1025(.dinb(n2952), .dina(n4012), .dout(n4016));
    jand g1026(.dinb(n11329), .dina(n2256), .dout(n4020));
    jor g1027(.dinb(n3286), .dina(n7025), .dout(n4024));
    jor g1028(.dinb(n4016), .dina(n4024), .dout(n4028));
    jnot g1029(.din(n4028), .dout(n4031));
    jand g1030(.dinb(n7022), .dina(n4031), .dout(n4035));
    jand g1031(.dinb(n7016), .dina(n4035), .dout(n4039));
    jand g1032(.dinb(n11428), .dina(n77), .dout(n4043));
    jor g1033(.dinb(n4039), .dina(n7013), .dout(n4047));
    jor g1034(.dinb(n6989), .dina(n4047), .dout(n4051));
    jand g1035(.dinb(n6986), .dina(n4051), .dout(n4055));
    jand g1036(.dinb(n8638), .dina(n2646), .dout(n4059));
    jor g1037(.dinb(n2121), .dina(n6962), .dout(n4063));
    jor g1038(.dinb(n4055), .dina(n6956), .dout(n4067));
    jor g1039(.dinb(n3890), .dina(n6941), .dout(n4071));
    jand g1040(.dinb(n3886), .dina(n6935), .dout(n4075));
    jand g1041(.dinb(n6917), .dina(n4075), .dout(n4079));
    jnot g1042(.din(n4079), .dout(n4082));
    jand g1043(.dinb(n3623), .dina(n3642), .dout(n4086));
    jnot g1044(.din(n4086), .dout(n4089));
    jand g1045(.dinb(n9667), .dina(n3646), .dout(n4093));
    jand g1046(.dinb(n4089), .dina(n4093), .dout(n4097));
    jnot g1047(.din(n4097), .dout(n4100));
    jor g1048(.dinb(n9490), .dina(n3642), .dout(n4104));
    jand g1049(.dinb(n9274), .dina(n3634), .dout(n4108));
    jnot g1050(.din(n4108), .dout(n4111));
    jand g1051(.dinb(n8668), .dina(n2189), .dout(n4115));
    jand g1052(.dinb(n8875), .dina(n2167), .dout(n4119));
    jand g1053(.dinb(n8864), .dina(n2264), .dout(n4123));
    jor g1054(.dinb(n4119), .dina(n8324), .dout(n4127));
    jor g1055(.dinb(n8321), .dina(n4127), .dout(n4131));
    jand g1056(.dinb(n8308), .dina(n2220), .dout(n4135));
    jor g1057(.dinb(n11437), .dina(n4135), .dout(n4139));
    jand g1058(.dinb(n8992), .dina(n2240), .dout(n4143));
    jand g1059(.dinb(n8855), .dina(n2204), .dout(n4147));
    jor g1060(.dinb(n4143), .dina(n4147), .dout(n4151));
    jand g1061(.dinb(n9083), .dina(n2256), .dout(n4155));
    jor g1062(.dinb(n3978), .dina(n8300), .dout(n4159));
    jor g1063(.dinb(n8297), .dina(n4159), .dout(n4163));
    jor g1064(.dinb(n8294), .dina(n4163), .dout(n4167));
    jor g1065(.dinb(n8291), .dina(n4167), .dout(n4171));
    jand g1066(.dinb(n11182), .dina(n2167), .dout(n4175));
    jand g1067(.dinb(n10285), .dina(n2256), .dout(n4179));
    jand g1068(.dinb(n11320), .dina(n2264), .dout(n4183));
    jor g1069(.dinb(n4179), .dina(n4183), .dout(n4187));
    jor g1070(.dinb(n4175), .dina(n4187), .dout(n4191));
    jand g1071(.dinb(n10543), .dina(n2220), .dout(n4195));
    jor g1072(.dinb(n8266), .dina(n4195), .dout(n4199));
    jand g1073(.dinb(n11050), .dina(n2240), .dout(n4203));
    jand g1074(.dinb(n10774), .dina(n2204), .dout(n4207));
    jor g1075(.dinb(n4203), .dina(n4207), .dout(n4211));
    jor g1076(.dinb(n2959), .dina(n3246), .dout(n4215));
    jor g1077(.dinb(n8228), .dina(n4215), .dout(n4219));
    jor g1078(.dinb(n8225), .dina(n4219), .dout(n4223));
    jor g1079(.dinb(n8222), .dina(n4223), .dout(n4227));
    jand g1080(.dinb(n4171), .dina(n4227), .dout(n4231));
    jor g1081(.dinb(n8329), .dina(n4231), .dout(n4235));
    jand g1082(.dinb(n8593), .dina(n2646), .dout(n4239));
    jor g1083(.dinb(n2121), .dina(n8216), .dout(n4243));
    jnot g1084(.din(n4243), .dout(n4246));
    jand g1085(.dinb(n4235), .dina(n8210), .dout(n4250));
    jand g1086(.dinb(n4111), .dina(n8204), .dout(n4254));
    jnot g1087(.din(n4254), .dout(n4257));
    jand g1088(.dinb(n4104), .dina(n4257), .dout(n4261));
    jand g1089(.dinb(n4100), .dina(n8189), .dout(n4265));
    jnot g1090(.din(n4265), .dout(n4268));
    jand g1091(.dinb(n7171), .dina(n4079), .dout(n4272));
    jnot g1092(.din(n3158), .dout(n4275));
    jnot g1093(.din(n2444), .dout(n4278));
    jand g1094(.dinb(n6686), .dina(n3394), .dout(n4282));
    jand g1095(.dinb(n8686), .dina(n4282), .dout(n4286));
    jand g1096(.dinb(n7321), .dina(n4286), .dout(n4290));
    jand g1097(.dinb(n8182), .dina(n4290), .dout(n4294));
    jand g1098(.dinb(n4275), .dina(n4294), .dout(n4298));
    jand g1099(.dinb(n4272), .dina(n4298), .dout(n4302));
    jnot g1100(.din(n4302), .dout(n4305));
    jnot g1101(.din(G213), .dout(n4308));
    jnot g1102(.din(G343), .dout(n4311));
    jand g1103(.dinb(n6838), .dina(n4272), .dout(n4315));
    jor g1104(.dinb(n6677), .dina(n4315), .dout(n4319));
    jor g1105(.dinb(n6679), .dina(n4319), .dout(G409));
    jxor g1106(.dinb(n8680), .dina(n4265), .dout(n4327));
    jxor g1107(.dinb(n7789), .dina(n3394), .dout(n4331));
    jxor g1108(.dinb(n3158), .dina(n7315), .dout(n4335));
    jxor g1109(.dinb(n7313), .dina(n4335), .dout(n4339));
    jxor g1110(.dinb(n7304), .dina(n4339), .dout(n4343));
    jand g1111(.dinb(n10189), .dina(n4311), .dout(n4347));
    jnot g1112(.din(n4347), .dout(n4350));
    jor g1113(.dinb(n6764), .dina(n4350), .dout(n4354));
    jxor g1114(.dinb(n7165), .dina(n4079), .dout(n4358));
    jor g1115(.dinb(n6766), .dina(n4358), .dout(n4362));
    jand g1116(.dinb(n6755), .dina(n4362), .dout(n4366));
    jxor g1117(.dinb(n7297), .dina(n4366), .dout(G405));
    jxor g1118(.dinb(n4343), .dina(n6913), .dout(n4374));
    jdff dff_A_ysFzlHig4_2(.din(n4374), .dout(G402));
    jdff dff_A_jCISqWYT9_1(.din(n4305), .dout(G407));
    jdff dff_A_UJV9lTxp4_0(.din(n12235), .dout(G381));
    jdff dff_A_FoPg98jD2_0(.din(n12232), .dout(n12235));
    jdff dff_A_Sp6VE8id9_0(.din(n12229), .dout(n12232));
    jdff dff_A_OYV2J0ds3_0(.din(n12226), .dout(n12229));
    jdff dff_A_BEk3hAnd8_1(.din(n4268), .dout(n12226));
    jdff dff_A_VKLgk1X27_0(.din(n12220), .dout(G375));
    jdff dff_A_CB5hT0D90_0(.din(n12217), .dout(n12220));
    jdff dff_A_ULxsSlua0_1(.din(n4082), .dout(n12217));
    jdff dff_A_RAOIGzOa2_0(.din(n12211), .dout(G378));
    jdff dff_A_KbweROGQ1_0(.din(n12208), .dout(n12211));
    jdff dff_A_Y34FfsEq6_0(.din(n12205), .dout(n12208));
    jdff dff_A_hCj3951Q9_0(.din(n12202), .dout(n12205));
    jdff dff_A_ywGiTRig5_1(.din(n3833), .dout(n12202));
    jdff dff_A_aUQ6yJFl6_0(.din(n12196), .dout(G390));
    jdff dff_A_Ev65jC9w8_0(.din(n12193), .dout(n12196));
    jdff dff_A_PDseqAHC6_0(.din(n12190), .dout(n12193));
    jdff dff_A_OSUarnG38_0(.din(n12187), .dout(n12190));
    jdff dff_A_h8B1FVzK0_0(.din(n12184), .dout(n12187));
    jdff dff_A_zmyyTuog8_1(.din(n3596), .dout(n12184));
    jdff dff_A_63rnxrt66_0(.din(n12178), .dout(G393));
    jdff dff_A_lGrXPsPf5_0(.din(n12175), .dout(n12178));
    jdff dff_A_7B7YrEgs1_0(.din(n12172), .dout(n12175));
    jdff dff_A_QDHzbLAS4_0(.din(n12169), .dout(n12172));
    jdff dff_A_EZIh7BOM0_0(.din(n12166), .dout(n12169));
    jdff dff_A_1wa6scRT4_0(.din(n12163), .dout(n12166));
    jdff dff_A_6AG3SgwF9_1(.din(n3397), .dout(n12163));
    jdff dff_A_C6v6yx9W8_0(.din(n12157), .dout(G387));
    jdff dff_A_lh9HrNeF8_0(.din(n12154), .dout(n12157));
    jdff dff_A_J8CYK0z98_0(.din(n12151), .dout(n12154));
    jdff dff_A_pePACUYr0_0(.din(n12148), .dout(n12151));
    jdff dff_A_gMbPIbhZ9_2(.din(n3158), .dout(n12148));
    jdff dff_A_1OsQOe6J0_0(.din(n12142), .dout(G367));
    jdff dff_A_VkvuCOeX2_0(.din(n12139), .dout(n12142));
    jdff dff_A_NuQSjE8t0_0(.din(n12136), .dout(n12139));
    jdff dff_A_kItvCpdm3_0(.din(n12133), .dout(n12136));
    jdff dff_A_OjXgsc6F9_2(.din(n2848), .dout(n12133));
    jdff dff_A_dwFfx8zJ1_0(.din(n12127), .dout(G384));
    jdff dff_A_KfbbFbyt7_0(.din(n12124), .dout(n12127));
    jdff dff_A_qeYaqAiR2_0(.din(n12121), .dout(n12124));
    jdff dff_A_Dz2LoSbI3_0(.din(n12118), .dout(n12121));
    jdff dff_A_pZuEXSwI3_0(.din(n12115), .dout(n12118));
    jdff dff_A_8GJ6RkPC8_0(.din(n12112), .dout(n12115));
    jdff dff_A_T3sTSkls0_0(.din(n12109), .dout(n12112));
    jdff dff_A_MK7puvqH4_1(.din(n2675), .dout(n12109));
    jdff dff_A_SdWRPurT6_0(.din(n12103), .dout(G396));
    jdff dff_A_yQqCGAVL5_0(.din(n12100), .dout(n12103));
    jdff dff_A_o6sNFGwq7_0(.din(n12097), .dout(n12100));
    jdff dff_A_idLnCTGo6_0(.din(n12094), .dout(n12097));
    jdff dff_A_KTddD5ff1_0(.din(n12091), .dout(n12094));
    jdff dff_A_hI41J0ac3_0(.din(n12088), .dout(n12091));
    jdff dff_A_LtUMQUBu0_0(.din(n12085), .dout(n12088));
    jdff dff_A_fgn35j2M0_0(.din(n12082), .dout(n12085));
    jdff dff_A_zJMLiDnG9_0(.din(n12079), .dout(n12082));
    jdff dff_A_7jU79r5T3_0(.din(n12076), .dout(n12079));
    jdff dff_A_JvhgudXb7_2(.din(n2444), .dout(n12076));
    jdff dff_A_eJhMTvLA1_0(.din(n12070), .dout(G364));
    jdff dff_A_x0zfNS5s1_0(.din(n12067), .dout(n12070));
    jdff dff_A_j3MvBzGw5_0(.din(n12064), .dout(n12067));
    jdff dff_A_iCJiOi5u8_0(.din(n12061), .dout(n12064));
    jdff dff_A_hblpjV0x7_0(.din(n12058), .dout(n12061));
    jdff dff_A_04fPKSR12_0(.din(n12055), .dout(n12058));
    jdff dff_A_WIolRQIE1_0(.din(n12052), .dout(n12055));
    jdff dff_A_nfIuEa7O8_0(.din(n12049), .dout(n12052));
    jdff dff_A_ipYufpMg8_0(.din(n12046), .dout(n12049));
    jdff dff_A_bjZscRO61_0(.din(n12043), .dout(n12046));
    jdff dff_A_0WVEvPGS5_2(.din(n2096), .dout(n12043));
    jdff dff_A_E7jguRXM1_0(.din(n12037), .dout(G399));
    jdff dff_A_hwO46wRc7_0(.din(n12034), .dout(n12037));
    jdff dff_A_kYLZHSdZ3_0(.din(n12031), .dout(n12034));
    jdff dff_A_wzJh5yps6_0(.din(n12028), .dout(n12031));
    jdff dff_A_IBhUu7Qm6_0(.din(n12025), .dout(n12028));
    jdff dff_A_bUqrFaCj4_0(.din(n12022), .dout(n12025));
    jdff dff_A_oYxdiuPb2_0(.din(n12019), .dout(n12022));
    jdff dff_A_dC2RTqVH5_0(.din(n12016), .dout(n12019));
    jdff dff_A_sZTAlPqr8_0(.din(n12013), .dout(n12016));
    jdff dff_A_40r01Umj8_0(.din(n12010), .dout(n12013));
    jdff dff_A_TMIQp7yB0_2(.din(n2005), .dout(n12010));
    jdff dff_A_SyK2xPPD8_0(.din(n12004), .dout(G369));
    jdff dff_A_Y7PXSUVf4_0(.din(n12001), .dout(n12004));
    jdff dff_A_On5sCEYo3_0(.din(n11998), .dout(n12001));
    jdff dff_A_Hsa47J9Y2_0(.din(n11995), .dout(n11998));
    jdff dff_A_EpvJVHbi5_0(.din(n11992), .dout(n11995));
    jdff dff_A_ohcL0so56_0(.din(n11989), .dout(n11992));
    jdff dff_A_Q5jFwPwD3_0(.din(n11986), .dout(n11989));
    jdff dff_A_LPvpTHiz2_0(.din(n11983), .dout(n11986));
    jdff dff_A_NE5UXxOC0_0(.din(n11980), .dout(n11983));
    jdff dff_A_VOcmU1MJ3_0(.din(n11977), .dout(n11980));
    jdff dff_A_ILl5k9cI5_0(.din(n11974), .dout(n11977));
    jdff dff_A_yKE6Pi2p6_2(.din(n1908), .dout(n11974));
    jdff dff_A_swsvL5td8_0(.din(n11968), .dout(G372));
    jdff dff_A_rPyJpGr71_0(.din(n11965), .dout(n11968));
    jdff dff_A_vj5vTeuW9_0(.din(n11962), .dout(n11965));
    jdff dff_A_zrjxHRTb1_0(.din(n11959), .dout(n11962));
    jdff dff_A_cAUmK5Mm7_0(.din(n11956), .dout(n11959));
    jdff dff_A_UU5ENAX71_0(.din(n11953), .dout(n11956));
    jdff dff_A_lMKux7055_0(.din(n11950), .dout(n11953));
    jdff dff_A_CHVGcIuR9_0(.din(n11947), .dout(n11950));
    jdff dff_A_issZT9NH3_0(.din(n11944), .dout(n11947));
    jdff dff_A_XnUb4Zlr3_0(.din(n11941), .dout(n11944));
    jdff dff_A_qyS5Wz0A7_0(.din(n11938), .dout(n11941));
    jdff dff_A_d1Py6wvc5_0(.din(n11935), .dout(n11938));
    jdff dff_A_3SRJIUlD6_0(.din(n11932), .dout(n11935));
    jdff dff_A_Fo7AjoZB3_2(.din(n1795), .dout(n11932));
    jdff dff_A_XBN2pRht0_0(.din(n11926), .dout(G351));
    jdff dff_A_dnWPRKXl7_0(.din(n11923), .dout(n11926));
    jdff dff_A_kqRTBoj71_0(.din(n11920), .dout(n11923));
    jdff dff_A_VK5lhS117_0(.din(n11917), .dout(n11920));
    jdff dff_A_hqzYHSbg0_0(.din(n11914), .dout(n11917));
    jdff dff_A_2w8vXaEC5_0(.din(n11911), .dout(n11914));
    jdff dff_A_OC9iKQH58_0(.din(n11908), .dout(n11911));
    jdff dff_A_eAyqwCzZ6_0(.din(n11905), .dout(n11908));
    jdff dff_A_bl42ncSb2_0(.din(n11902), .dout(n11905));
    jdff dff_A_Il4rDvRK9_0(.din(n11899), .dout(n11902));
    jdff dff_A_xyL8Gekh9_0(.din(n11896), .dout(n11899));
    jdff dff_A_o6u0Nn5F9_0(.din(n11893), .dout(n11896));
    jdff dff_A_k1fWSuVW4_0(.din(n11890), .dout(n11893));
    jdff dff_A_TOneLI254_0(.din(n11887), .dout(n11890));
    jdff dff_A_mgfaHL9H3_0(.din(n11884), .dout(n11887));
    jdff dff_A_egVfUnC77_0(.din(n11881), .dout(n11884));
    jdff dff_A_2S85BXrz9_0(.din(n11878), .dout(n11881));
    jdff dff_A_vXZQ5h5j9_0(.din(n11875), .dout(n11878));
    jdff dff_A_cBFbio7O4_0(.din(n11872), .dout(n11875));
    jdff dff_A_V7ZJnNfe1_0(.din(n11869), .dout(n11872));
    jdff dff_A_f4p5mze87_0(.din(n11866), .dout(n11869));
    jdff dff_A_u2pQx0fr2_0(.din(n11863), .dout(n11866));
    jdff dff_A_N4XF6Hnn0_0(.din(n11860), .dout(n11863));
    jdff dff_A_hm8XpUoB1_2(.din(n340), .dout(n11860));
    jdff dff_A_KNTDztRT6_0(.din(n11854), .dout(G358));
    jdff dff_A_fOdpVXOa1_0(.din(n11851), .dout(n11854));
    jdff dff_A_OcB7E4FS6_0(.din(n11848), .dout(n11851));
    jdff dff_A_dFuDFUHC4_0(.din(n11845), .dout(n11848));
    jdff dff_A_nyPwmjWf0_0(.din(n11842), .dout(n11845));
    jdff dff_A_oglXmj6O5_0(.din(n11839), .dout(n11842));
    jdff dff_A_f7inSK2C2_0(.din(n11836), .dout(n11839));
    jdff dff_A_GJc1JsfS1_0(.din(n11833), .dout(n11836));
    jdff dff_A_PrdI3O528_0(.din(n11830), .dout(n11833));
    jdff dff_A_XwkblzX26_0(.din(n11827), .dout(n11830));
    jdff dff_A_JxT0K3Sj4_0(.din(n11824), .dout(n11827));
    jdff dff_A_9JTme08A5_0(.din(n11821), .dout(n11824));
    jdff dff_A_Aw3cQnog9_0(.din(n11818), .dout(n11821));
    jdff dff_A_PSGaGukk8_0(.din(n11815), .dout(n11818));
    jdff dff_A_7xcccwWZ0_0(.din(n11812), .dout(n11815));
    jdff dff_A_kbFLxLLY1_0(.din(n11809), .dout(n11812));
    jdff dff_A_M1uryMSr8_0(.din(n11806), .dout(n11809));
    jdff dff_A_AJsGT4HC7_0(.din(n11803), .dout(n11806));
    jdff dff_A_S8gd0K6y9_0(.din(n11800), .dout(n11803));
    jdff dff_A_YLwcEg3v9_0(.din(n11797), .dout(n11800));
    jdff dff_A_b7GGSp3J5_0(.din(n11794), .dout(n11797));
    jdff dff_A_i5LiCjT30_0(.din(n11791), .dout(n11794));
    jdff dff_A_ETfMRraI8_0(.din(n11788), .dout(n11791));
    jdff dff_A_KxktjB0M1_2(.din(n306), .dout(n11788));
    jdff dff_A_hyFJq4Tp4_0(.din(n11782), .dout(G361));
    jdff dff_A_CLRBlX9P2_0(.din(n11779), .dout(n11782));
    jdff dff_A_h1nEpwY53_0(.din(n11776), .dout(n11779));
    jdff dff_A_6z13bnug1_0(.din(n11773), .dout(n11776));
    jdff dff_A_2j63eibE7_0(.din(n11770), .dout(n11773));
    jdff dff_A_igeNho1x0_0(.din(n11767), .dout(n11770));
    jdff dff_A_LCwPXFQN8_0(.din(n11764), .dout(n11767));
    jdff dff_A_F7PTQD1p0_0(.din(n11761), .dout(n11764));
    jdff dff_A_MUil1Pu22_0(.din(n11758), .dout(n11761));
    jdff dff_A_GgQZkZ8N0_0(.din(n11755), .dout(n11758));
    jdff dff_A_LSXYNV9I7_0(.din(n11752), .dout(n11755));
    jdff dff_A_gqOq2OKz3_0(.din(n11749), .dout(n11752));
    jdff dff_A_fLrCvENM3_0(.din(n11746), .dout(n11749));
    jdff dff_A_eFcD9XJe2_0(.din(n11743), .dout(n11746));
    jdff dff_A_rPmcsS9X7_0(.din(n11740), .dout(n11743));
    jdff dff_A_ypir7DjH3_0(.din(n11737), .dout(n11740));
    jdff dff_A_sMl3qcMf6_0(.din(n11734), .dout(n11737));
    jdff dff_A_mCSCtIhU9_0(.din(n11731), .dout(n11734));
    jdff dff_A_lGzCx7Df2_0(.din(n11728), .dout(n11731));
    jdff dff_A_bPEi8vwn8_0(.din(n11725), .dout(n11728));
    jdff dff_A_yu2mnwg27_2(.din(n275), .dout(n11725));
    jdff dff_A_yunia8tt0_0(.din(n11719), .dout(G355));
    jdff dff_A_gWKpw2w06_0(.din(n11716), .dout(n11719));
    jdff dff_A_oyZYblEz3_0(.din(n11713), .dout(n11716));
    jdff dff_A_JyflBbLh1_0(.din(n11710), .dout(n11713));
    jdff dff_A_k5zRfPFm4_0(.din(n11707), .dout(n11710));
    jdff dff_A_Hl1KhlD93_0(.din(n11704), .dout(n11707));
    jdff dff_A_GCl3sPpe3_0(.din(n11701), .dout(n11704));
    jdff dff_A_mHTJaAdx4_0(.din(n11698), .dout(n11701));
    jdff dff_A_A9gopoxK0_0(.din(n11695), .dout(n11698));
    jdff dff_A_uxR2QE8v0_0(.din(n11692), .dout(n11695));
    jdff dff_A_mzsI8NCp0_0(.din(n11689), .dout(n11692));
    jdff dff_A_XSxjnDbD9_0(.din(n11686), .dout(n11689));
    jdff dff_A_2VzzZEfu5_0(.din(n11683), .dout(n11686));
    jdff dff_A_2ewcdiOT9_0(.din(n11680), .dout(n11683));
    jdff dff_A_c60NlIbj0_0(.din(n11677), .dout(n11680));
    jdff dff_A_jsIA8eKB8_0(.din(n11674), .dout(n11677));
    jdff dff_A_XA72lHkS1_0(.din(n11671), .dout(n11674));
    jdff dff_A_aI3kkDP84_0(.din(n11668), .dout(n11671));
    jdff dff_A_wKJWkuGj9_0(.din(n11665), .dout(n11668));
    jdff dff_A_4ge9LgrV4_0(.din(n11662), .dout(n11665));
    jdff dff_A_0thdKQix0_0(.din(n11659), .dout(n11662));
    jdff dff_A_5nhhep6d9_0(.din(n11656), .dout(n11659));
    jdff dff_A_3D80Yf1i6_0(.din(n11653), .dout(n11656));
    jdff dff_A_b4JJi3Xo9_1(.din(n115), .dout(n11653));
    jdff dff_A_ihUofMly6_0(.din(n11647), .dout(G353));
    jdff dff_A_PFGQIOju3_0(.din(n11644), .dout(n11647));
    jdff dff_A_HGzp22941_0(.din(n11641), .dout(n11644));
    jdff dff_A_46Ybfo041_0(.din(n11638), .dout(n11641));
    jdff dff_A_mkE7Z8ts0_0(.din(n11635), .dout(n11638));
    jdff dff_A_LAqLvMI30_0(.din(n11632), .dout(n11635));
    jdff dff_A_MQoacw8Q9_0(.din(n11629), .dout(n11632));
    jdff dff_A_NbxblaA19_0(.din(n11626), .dout(n11629));
    jdff dff_A_W46RsyYx0_0(.din(n11623), .dout(n11626));
    jdff dff_A_XHUR7MiC5_0(.din(n11620), .dout(n11623));
    jdff dff_A_Py8YTI9G5_0(.din(n11617), .dout(n11620));
    jdff dff_A_sO0ezfUK2_0(.din(n11614), .dout(n11617));
    jdff dff_A_0TUAKMoS1_0(.din(n11611), .dout(n11614));
    jdff dff_A_Vdc5lXXl2_0(.din(n11608), .dout(n11611));
    jdff dff_A_FE7Sq7Tl2_0(.din(n11605), .dout(n11608));
    jdff dff_A_ja7F6qH94_0(.din(n11602), .dout(n11605));
    jdff dff_A_qtcryspU0_0(.din(n11599), .dout(n11602));
    jdff dff_A_ou87bcHz4_0(.din(n11596), .dout(n11599));
    jdff dff_A_04jcxYzU7_0(.din(n11593), .dout(n11596));
    jdff dff_A_XEUnkOtK1_0(.din(n11590), .dout(n11593));
    jdff dff_A_bPrcsCRS4_0(.din(n11587), .dout(n11590));
    jdff dff_A_8JwgpaaC9_0(.din(n11584), .dout(n11587));
    jdff dff_A_yTGtcVRg0_0(.din(n11581), .dout(n11584));
    jdff dff_A_oCeIctIc4_0(.din(n11578), .dout(n11581));
    jdff dff_A_jDDyjmOM9_2(.din(n95), .dout(n11578));
    jdff dff_A_QuWBZkPP5_2(.din(G169), .dout(n11575));
    jdff dff_A_YxIiNnCT8_2(.din(n11575), .dout(n11572));
    jdff dff_A_PWB9Dwhw3_2(.din(n11572), .dout(n11569));
    jdff dff_A_myXmhWVs2_2(.din(n11569), .dout(n11566));
    jdff dff_A_6mrcnqob9_2(.din(n11566), .dout(n11563));
    jdff dff_A_FLMG89st7_2(.din(n11563), .dout(n11560));
    jdff dff_A_jZlf7qoN7_2(.din(n11560), .dout(n11557));
    jdff dff_A_73xXv1qJ4_1(.din(G169), .dout(n11554));
    jdff dff_A_cNWazVGD3_1(.din(n11554), .dout(n11551));
    jdff dff_A_5YOTw2ai0_1(.din(n11551), .dout(n11548));
    jdff dff_A_gcq7ZLJ48_1(.din(n11548), .dout(n11545));
    jdff dff_A_SXKzKZXg9_1(.din(n11545), .dout(n11542));
    jdff dff_A_76qXpSFo4_1(.din(n11542), .dout(n11539));
    jdff dff_A_BTJJSqX32_1(.din(n11539), .dout(n11536));
    jdff dff_A_G6PyO8im8_0(.din(G169), .dout(n11533));
    jdff dff_A_Hn2rZI4c7_0(.din(n11533), .dout(n11530));
    jdff dff_A_6ZgD6zws4_0(.din(n11530), .dout(n11527));
    jdff dff_A_hdZFUim10_0(.din(n11527), .dout(n11524));
    jdff dff_A_sLGr2W334_0(.din(n11524), .dout(n11521));
    jdff dff_A_GM2LTRIx2_0(.din(n11521), .dout(n11518));
    jdff dff_A_SDNStn4c4_0(.din(n11518), .dout(n11515));
    jdff dff_A_fLtmlSke3_2(.din(n343), .dout(n11512));
    jdff dff_A_9tTkdQcL6_2(.din(n11512), .dout(n11509));
    jdff dff_A_VsF606or9_2(.din(n11509), .dout(n11506));
    jdff dff_A_PpQpP64P8_2(.din(n11506), .dout(n11503));
    jdff dff_A_awll7jxE2_2(.din(n11503), .dout(n11500));
    jdff dff_A_UBBdH3Pi7_2(.din(n11500), .dout(n11497));
    jdff dff_A_m8wv256D9_1(.din(n343), .dout(n11494));
    jdff dff_A_xsBHwhZ30_1(.din(n11494), .dout(n11491));
    jdff dff_A_quvSuv8u5_1(.din(n11491), .dout(n11488));
    jdff dff_A_l0bbccIh9_1(.din(n11488), .dout(n11485));
    jdff dff_A_EA9FYDxy9_1(.din(n11485), .dout(n11482));
    jdff dff_A_YK0gGx2Z1_1(.din(n11482), .dout(n11479));
    jdff dff_A_iAdXw7Hj8_0(.din(G1), .dout(n11476));
    jdff dff_A_O3PSfUPA3_2(.din(G1), .dout(n11473));
    jdff dff_A_3nvoBC4Z2_0(.din(G1), .dout(n11470));
    jdff dff_A_0eRuYOQO3_2(.din(G13), .dout(n11467));
    jdff dff_A_4bLfR68l3_2(.din(n11467), .dout(n11464));
    jdff dff_A_pLbnh99t5_1(.din(G13), .dout(n11461));
    jdff dff_A_PQfOk9nx5_2(.din(n347), .dout(n11458));
    jdff dff_A_slPEs5cW2_1(.din(n347), .dout(n11455));
    jdff dff_A_KPWEOBb32_0(.din(G33), .dout(n11452));
    jdff dff_A_8qgATIe62_2(.din(G33), .dout(n11449));
    jdff dff_A_a59X2VON1_2(.din(n11449), .dout(n11446));
    jdff dff_A_ogfXx8KF4_2(.din(n11446), .dout(n11443));
    jdff dff_A_inB6gsfz0_2(.din(n11443), .dout(n11440));
    jdff dff_A_a3mhyjEm2_2(.din(n11440), .dout(n11437));
    jdff dff_A_AH0KJFDU0_2(.din(G41), .dout(n11434));
    jdff dff_A_HgYY2dUb4_2(.din(n11434), .dout(n11431));
    jdff dff_A_eheZoAGo8_1(.din(G41), .dout(n11428));
    jdff dff_A_sgKsKajD0_0(.din(n353), .dout(n11425));
    jdff dff_A_bZl15ToZ9_1(.din(n361), .dout(n11422));
    jdff dff_A_FJazkNfU9_1(.din(n11422), .dout(n11419));
    jdff dff_A_EWytyrHp6_2(.din(n361), .dout(n11416));
    jdff dff_A_eRcHLr176_2(.din(n11416), .dout(n11413));
    jdff dff_A_kDyzheB88_1(.din(n361), .dout(n11410));
    jdff dff_A_rYRdCdk93_1(.din(n11410), .dout(n11407));
    jdff dff_A_upYG8lUr4_2(.din(n361), .dout(n11404));
    jdff dff_A_ppGTzq2G7_2(.din(n11404), .dout(n11401));
    jdff dff_A_bj6XxWiH2_2(.din(G244), .dout(n11398));
    jdff dff_A_4o0p8slk3_2(.din(n11398), .dout(n11395));
    jdff dff_A_iaPOG52y2_1(.din(G244), .dout(n11392));
    jdff dff_A_lJ3aMjpq8_1(.din(n11392), .dout(n11389));
    jdff dff_A_6nObsZ5H3_1(.din(n11389), .dout(n11386));
    jdff dff_A_06D0wKbJ5_1(.din(n11386), .dout(n11383));
    jdff dff_A_oHNNeNEI2_0(.din(G244), .dout(n11380));
    jdff dff_A_Z0cjFDHq7_0(.din(n11380), .dout(n11377));
    jdff dff_A_Mlfa3Jcp5_2(.din(G1698), .dout(n11374));
    jdff dff_A_9N91VHxD5_2(.din(G238), .dout(n11371));
    jdff dff_A_zPI9h0pG0_2(.din(n11371), .dout(n11368));
    jdff dff_A_pJc5Nymd0_1(.din(G238), .dout(n11365));
    jdff dff_A_XCrtveZf8_1(.din(n11365), .dout(n11362));
    jdff dff_A_f3QAmBdV4_1(.din(n11362), .dout(n11359));
    jdff dff_A_hukRPu1H1_1(.din(n11359), .dout(n11356));
    jdff dff_A_303rdBsU8_0(.din(G238), .dout(n11353));
    jdff dff_A_TBnhXvjT5_0(.din(n11353), .dout(n11350));
    jdff dff_A_JUzIhdWg1_2(.din(G116), .dout(n11347));
    jdff dff_A_6sEZr79Z9_1(.din(G116), .dout(n11344));
    jdff dff_A_UpmNlgzu2_1(.din(n11344), .dout(n11341));
    jdff dff_A_fglkHkid8_1(.din(n11341), .dout(n11338));
    jdff dff_A_pzus6SVP7_2(.din(G116), .dout(n11335));
    jdff dff_A_Ar3Xl1TE6_2(.din(n11335), .dout(n11332));
    jdff dff_A_ktoydHJt5_2(.din(n11332), .dout(n11329));
    jdff dff_A_raVhjKGT5_1(.din(G116), .dout(n11326));
    jdff dff_A_WHghHJm77_1(.din(n11326), .dout(n11323));
    jdff dff_A_ydHFQ62C3_1(.din(n11323), .dout(n11320));
    jdff dff_A_tcKA3BhQ5_2(.din(n384), .dout(n11317));
    jdff dff_A_DQKieqpc6_2(.din(n11317), .dout(n11314));
    jdff dff_A_GHAbKBh17_0(.din(n384), .dout(n11311));
    jdff dff_A_9ww3VlH63_0(.din(n11311), .dout(n11308));
    jdff dff_B_GRNElknY8_1(.din(n369), .dout(n11306));
    jdff dff_A_c67gaj6g8_1(.din(G250), .dout(n11302));
    jdff dff_A_rZmdm5qG0_1(.din(n11302), .dout(n11299));
    jdff dff_A_0Dr2K6jL4_0(.din(G250), .dout(n11296));
    jdff dff_A_LFyYcmB27_0(.din(n11296), .dout(n11293));
    jdff dff_A_KVIzA3Ct9_1(.din(n165), .dout(n11290));
    jdff dff_A_hEPKzEzv3_0(.din(n165), .dout(n11287));
    jdff dff_A_UYUfUEAd4_2(.din(G45), .dout(n11284));
    jdff dff_A_TRFGqDUJ8_2(.din(n11284), .dout(n11281));
    jdff dff_A_bV0VerXU7_2(.din(n11281), .dout(n11278));
    jdff dff_A_yQTxWFRA1_1(.din(G45), .dout(n11275));
    jdff dff_A_qrTS6Gwh7_1(.din(n11275), .dout(n11272));
    jdff dff_A_tEVBWGW62_1(.din(n11272), .dout(n11269));
    jdff dff_A_GFDKQ38K5_1(.din(G45), .dout(n11266));
    jdff dff_A_CO9EWdaC6_0(.din(G45), .dout(n11263));
    jdff dff_A_ZxELQh9I5_0(.din(n11263), .dout(n11260));
    jdff dff_A_pIExNAhw0_2(.din(n399), .dout(n11257));
    jdff dff_A_Xy8ZZeI59_2(.din(n11257), .dout(n11254));
    jdff dff_A_USztoXLK7_2(.din(n11254), .dout(n11251));
    jdff dff_A_hTYt0Sei3_0(.din(n407), .dout(n11248));
    jdff dff_A_FoBBaqwL2_1(.din(n222), .dout(n11245));
    jdff dff_A_NG8iqZFU6_0(.din(n222), .dout(n11242));
    jdff dff_A_vtqn6Ngn9_2(.din(n226), .dout(n11239));
    jdff dff_B_WYnzbP1T3_0(.din(n414), .dout(n11237));
    jdff dff_A_UAPhG3Vn9_0(.din(n418), .dout(n11233));
    jdff dff_A_5BzSVzfU8_2(.din(G274), .dout(n11230));
    jdff dff_A_0eV7BkGz8_2(.din(n11230), .dout(n11227));
    jdff dff_A_coUzNFjU0_0(.din(G274), .dout(n11224));
    jdff dff_A_YQsvCYYk7_0(.din(n11224), .dout(n11221));
    jdff dff_A_PoliPYxD4_0(.din(n11221), .dout(n11218));
    jdff dff_B_2Q9ieLS33_0(.din(n430), .dout(n11216));
    jdff dff_A_4Ouj8ThX9_0(.din(n434), .dout(n11212));
    jdff dff_A_uZz1fQBT7_1(.din(G33), .dout(n11209));
    jdff dff_A_fxc072rn5_0(.din(G33), .dout(n11206));
    jdff dff_A_8qEqV5IG1_2(.din(G97), .dout(n11203));
    jdff dff_A_C9em7tj81_1(.din(G97), .dout(n11200));
    jdff dff_A_ALhdn8qc6_1(.din(n11200), .dout(n11197));
    jdff dff_A_b8Aotwq21_1(.din(n11197), .dout(n11194));
    jdff dff_A_9oPM0F8E6_2(.din(G97), .dout(n11191));
    jdff dff_A_6TTriCEI5_2(.din(n11191), .dout(n11188));
    jdff dff_A_MERfyLJc9_2(.din(n11188), .dout(n11185));
    jdff dff_A_Afu5Kpga3_2(.din(n11185), .dout(n11182));
    jdff dff_A_uB9kAt2B0_0(.din(G97), .dout(n11179));
    jdff dff_A_VF4oUAvq4_0(.din(n11179), .dout(n11176));
    jdff dff_A_iGp4QjM17_0(.din(n11176), .dout(n11173));
    jdff dff_B_mCDef9Oe5_2(.din(n11168), .dout(n11171));
    jdff dff_B_dhtP6ddm7_2(.din(n442), .dout(n11168));
    jdff dff_A_nOj7S6af6_0(.din(G20), .dout(n11164));
    jdff dff_A_Ekx2lsgO5_2(.din(n11164), .dout(n11161));
    jdff dff_A_1hQTGFhM4_0(.din(n11161), .dout(n11158));
    jdff dff_A_1cQcbg208_1(.din(n350), .dout(n11155));
    jdff dff_A_si08ltWt9_2(.din(G68), .dout(n11152));
    jdff dff_A_aD3bYPsb3_2(.din(G68), .dout(n11149));
    jdff dff_A_h2tkC4do5_2(.din(n11149), .dout(n11146));
    jdff dff_A_0ztcYfpW6_2(.din(n11146), .dout(n11143));
    jdff dff_A_DxGsPXO13_2(.din(n11143), .dout(n11140));
    jdff dff_A_0corOKVj7_0(.din(G68), .dout(n11137));
    jdff dff_A_PJNWczpa1_1(.din(n11137), .dout(n11134));
    jdff dff_A_8wMjJHIG7_0(.din(n11137), .dout(n11131));
    jdff dff_A_Madlfysn3_1(.din(G20), .dout(n11128));
    jdff dff_A_VSlHQ9P36_2(.din(n216), .dout(n11125));
    jdff dff_A_F7j5jKl69_2(.din(n469), .dout(n11122));
    jdff dff_A_Vmkku8fN4_2(.din(n11122), .dout(n11119));
    jdff dff_A_jPwCkNEH8_1(.din(n469), .dout(n11116));
    jdff dff_A_w42ZATqo8_1(.din(n11116), .dout(n11113));
    jdff dff_A_yTyBwOZq2_0(.din(G87), .dout(n11110));
    jdff dff_A_vI1MDHPb8_0(.din(n11110), .dout(n11107));
    jdff dff_A_3AMTUf409_0(.din(n11107), .dout(n11104));
    jdff dff_A_c7vPv7cN1_2(.din(G87), .dout(n11101));
    jdff dff_A_oGYHcEpi4_2(.din(n11101), .dout(n11098));
    jdff dff_A_ZsQLVsqs3_2(.din(n11098), .dout(n11095));
    jdff dff_A_001aC8LN9_0(.din(G87), .dout(n11092));
    jdff dff_A_swqtA9sL9_0(.din(n162), .dout(n11089));
    jdff dff_A_AZl59P653_1(.din(n11089), .dout(n11086));
    jdff dff_A_GViDkCJD7_0(.din(G97), .dout(n11083));
    jdff dff_A_vIXjKMLs5_0(.din(n98), .dout(n11080));
    jdff dff_A_W52wfV0H7_0(.din(n11080), .dout(n11077));
    jdff dff_A_pw1EcozM1_2(.din(G107), .dout(n11074));
    jdff dff_A_fWt6MUaE7_2(.din(n11074), .dout(n11071));
    jdff dff_A_tsI1dVCL6_2(.din(n11071), .dout(n11068));
    jdff dff_A_FTkE7pQJ2_1(.din(G107), .dout(n11065));
    jdff dff_A_pd9Unxrj0_1(.din(n11065), .dout(n11062));
    jdff dff_A_31bST4RG1_1(.din(n11062), .dout(n11059));
    jdff dff_A_O1jHvSWP8_2(.din(G107), .dout(n11056));
    jdff dff_A_dmDIpHXg8_2(.din(n11056), .dout(n11053));
    jdff dff_A_NY5FChnJ6_2(.din(n11053), .dout(n11050));
    jdff dff_A_h6lmthOs1_2(.din(n101), .dout(n11047));
    jdff dff_A_Ilu1AmxG0_2(.din(n11047), .dout(n11044));
    jdff dff_A_lqG2rG0X8_2(.din(n11044), .dout(n11041));
    jdff dff_A_mnmkF3jC1_2(.din(n11041), .dout(n11038));
    jdff dff_A_6luVzNKG7_2(.din(n11038), .dout(n11035));
    jdff dff_A_ffrbgNc21_1(.din(n101), .dout(n11032));
    jdff dff_A_sasnW2SN5_1(.din(n11032), .dout(n11029));
    jdff dff_A_gHYXEe3V2_1(.din(n11029), .dout(n11026));
    jdff dff_A_J9rY81dQ7_1(.din(n11164), .dout(n11023));
    jdff dff_A_tnr0FCP54_0(.din(n11164), .dout(n11020));
    jdff dff_A_HZd2GatY8_2(.din(n119), .dout(n11017));
    jdff dff_A_VyS28cge1_2(.din(n11017), .dout(n11014));
    jdff dff_A_bDTE1pCU5_2(.din(n11014), .dout(n11011));
    jdff dff_A_UAB7M2MC5_2(.din(n11011), .dout(n11008));
    jdff dff_A_65zy7shZ0_0(.din(n119), .dout(n11005));
    jdff dff_A_tijpbY7D0_0(.din(n11005), .dout(n11002));
    jdff dff_A_ObhdSrtI1_2(.din(n508), .dout(n10999));
    jdff dff_A_bYTrrIyV4_0(.din(n508), .dout(n10996));
    jdff dff_A_NTvaMBSR8_0(.din(n10996), .dout(n10993));
    jdff dff_A_BhaIHiIi3_1(.din(n512), .dout(n10990));
    jdff dff_B_CTKC3q9z3_0(.din(n520), .dout(n10988));
    jdff dff_A_Dr0dLoVk1_0(.din(G179), .dout(n10984));
    jdff dff_A_f208jTEV9_0(.din(n10984), .dout(n10981));
    jdff dff_A_NS9sNu3e4_0(.din(n10981), .dout(n10978));
    jdff dff_A_WJoMVyUr7_0(.din(n10978), .dout(n10975));
    jdff dff_A_ZUQtZJlv5_0(.din(n10975), .dout(n10972));
    jdff dff_A_4SFMbZqQ6_0(.din(n10972), .dout(n10969));
    jdff dff_A_lF4JxzxQ2_0(.din(n10969), .dout(n10966));
    jdff dff_A_J1ih0qTn6_1(.din(G179), .dout(n10963));
    jdff dff_A_7k4l7qt24_1(.din(n10963), .dout(n10960));
    jdff dff_A_q1vMp6Xt8_1(.din(n10960), .dout(n10957));
    jdff dff_A_QzUOOnDj6_1(.din(n10957), .dout(n10954));
    jdff dff_A_q7JbCo8W6_1(.din(n10954), .dout(n10951));
    jdff dff_A_hJM2TBQB1_1(.din(n10951), .dout(n10948));
    jdff dff_A_DLUYiEM47_1(.din(n10948), .dout(n10945));
    jdff dff_A_suGe9WPO6_0(.din(G179), .dout(n10942));
    jdff dff_A_Fqlu81ZI1_0(.din(n10942), .dout(n10939));
    jdff dff_A_Ks2d8K442_0(.din(n10939), .dout(n10936));
    jdff dff_A_DE7AwlLp0_0(.din(n10936), .dout(n10933));
    jdff dff_A_e7tTGEca3_0(.din(n10933), .dout(n10930));
    jdff dff_A_XKSjJ5hH1_0(.din(n10930), .dout(n10927));
    jdff dff_A_xCs0uLOj3_0(.din(n10927), .dout(n10924));
    jdff dff_B_kIJv506o1_3(.din(n10919), .dout(n10922));
    jdff dff_B_vNKcW1C49_3(.din(n10916), .dout(n10919));
    jdff dff_B_uYtT4eQu5_3(.din(n10913), .dout(n10916));
    jdff dff_B_HskBRdxc1_3(.din(n10910), .dout(n10913));
    jdff dff_B_T99fJxNq5_3(.din(n535), .dout(n10910));
    jdff dff_A_JFjoZqRm7_2(.din(n10922), .dout(n10906));
    jdff dff_A_ZTcFboHJ9_0(.din(n10922), .dout(n10903));
    jdff dff_A_VCFA39Bw3_1(.din(n10922), .dout(n10900));
    jdff dff_A_PWuV5Axc5_0(.din(n10922), .dout(n10897));
    jdff dff_A_6k8eSR7l3_1(.din(n183), .dout(n10894));
    jdff dff_A_uzO5xhyl4_2(.din(G33), .dout(n10891));
    jdff dff_A_mVCFVMyS7_0(.din(n554), .dout(n10888));
    jdff dff_B_6KcOzGgC9_2(.din(n569), .dout(n10886));
    jdff dff_A_PbvQEbvw8_0(.din(n10886), .dout(n10882));
    jdff dff_A_hz48tvZj2_0(.din(n589), .dout(n10879));
    jdff dff_A_0M59mrjU1_1(.din(n601), .dout(n10876));
    jdff dff_A_4kFVSjYh8_1(.din(n604), .dout(n10873));
    jdff dff_A_wCBPIBH18_1(.din(G190), .dout(n10870));
    jdff dff_A_F0YiJfRp5_1(.din(n10870), .dout(n10867));
    jdff dff_A_Ac1t2Z0B9_1(.din(n10867), .dout(n10864));
    jdff dff_A_dVvesc1C1_0(.din(G190), .dout(n10861));
    jdff dff_A_MToV3uQi0_0(.din(n10861), .dout(n10858));
    jdff dff_A_tkwBkKGg1_0(.din(n10858), .dout(n10855));
    jdff dff_A_7rw9GJCL1_0(.din(n10855), .dout(n10852));
    jdff dff_A_eeXcb0LK1_0(.din(n10852), .dout(n10849));
    jdff dff_A_wAzwG5NF6_0(.din(n10849), .dout(n10846));
    jdff dff_A_qayL26XG4_0(.din(n10846), .dout(n10843));
    jdff dff_A_mJWlEdhi3_2(.din(G200), .dout(n10840));
    jdff dff_A_4Il5uod24_2(.din(n10840), .dout(n10837));
    jdff dff_A_sMpOPvSM9_2(.din(n10837), .dout(n10834));
    jdff dff_A_LPUcDJBS2_2(.din(n10834), .dout(n10831));
    jdff dff_A_bN7ldxU20_2(.din(n10831), .dout(n10828));
    jdff dff_A_I4W3GC0P2_2(.din(n10828), .dout(n10825));
    jdff dff_A_2nITGxT72_2(.din(n10825), .dout(n10822));
    jdff dff_A_2pTMC7fh9_1(.din(G200), .dout(n10819));
    jdff dff_A_bGE5KNDJ7_0(.din(G200), .dout(n10816));
    jdff dff_A_3FKnpT776_0(.din(n10816), .dout(n10813));
    jdff dff_A_mWcYaPyM8_0(.din(n10813), .dout(n10810));
    jdff dff_A_4CpzGqHi7_0(.din(n10810), .dout(n10807));
    jdff dff_A_lt9IHk169_0(.din(n10807), .dout(n10804));
    jdff dff_A_26xsE9xa2_0(.din(n10804), .dout(n10801));
    jdff dff_A_8yi5hHaE5_0(.din(n10801), .dout(n10798));
    jdff dff_B_suPl964r6_1(.din(n608), .dout(n10796));
    jdff dff_A_EhSyXoq93_2(.din(n418), .dout(n10792));
    jdff dff_A_zlfUFNxN7_1(.din(G283), .dout(n10789));
    jdff dff_A_M3EiS25C9_1(.din(n10789), .dout(n10786));
    jdff dff_A_32enTWEY8_1(.din(n10786), .dout(n10783));
    jdff dff_A_REC5uBRg6_0(.din(G283), .dout(n10780));
    jdff dff_A_m64AZkit3_0(.din(n10780), .dout(n10777));
    jdff dff_A_vc88hoFt9_0(.din(n10777), .dout(n10774));
    jdff dff_A_U3y76x5D0_1(.din(G283), .dout(n10771));
    jdff dff_A_RndfyFv52_1(.din(n10771), .dout(n10768));
    jdff dff_A_G3VZeg0G8_1(.din(n10768), .dout(n10765));
    jdff dff_A_KPDjnYZZ5_1(.din(n10765), .dout(n10762));
    jdff dff_A_8GO6iolU1_0(.din(G283), .dout(n10759));
    jdff dff_A_JnrTIHvl0_0(.din(n10759), .dout(n10756));
    jdff dff_A_e6fQA4aB6_0(.din(n10756), .dout(n10753));
    jdff dff_A_zzM06KLE7_1(.din(n632), .dout(n10750));
    jdff dff_A_wFYZV4pb7_1(.din(n10750), .dout(n10747));
    jdff dff_A_3xRNxzVm0_0(.din(n632), .dout(n10744));
    jdff dff_A_udrKFxna6_0(.din(n10744), .dout(n10741));
    jdff dff_A_DtA0yE6o6_1(.din(n659), .dout(n10738));
    jdff dff_A_irs9bHBr5_2(.din(G257), .dout(n10735));
    jdff dff_A_IbB9Taz62_2(.din(n10735), .dout(n10732));
    jdff dff_A_l4Toek0g7_1(.din(G257), .dout(n10729));
    jdff dff_A_B60DKuWp4_1(.din(n10729), .dout(n10726));
    jdff dff_A_TfyK3HW66_1(.din(G257), .dout(n10723));
    jdff dff_A_EcODS1TM6_0(.din(G257), .dout(n10720));
    jdff dff_A_llzU1GyE4_0(.din(n10720), .dout(n10717));
    jdff dff_A_OEyQfNX14_0(.din(n10717), .dout(n10714));
    jdff dff_A_FROdvvJx1_0(.din(n10714), .dout(n10711));
    jdff dff_A_PsGS15dS5_1(.din(n140), .dout(n10708));
    jdff dff_A_QS6hAFmE7_0(.din(n140), .dout(n10705));
    jdff dff_A_VcdHeGSe5_0(.din(n10705), .dout(n10702));
    jdff dff_A_Mc4qclDQ7_0(.din(n10702), .dout(n10699));
    jdff dff_A_H6Myhpd09_1(.din(n361), .dout(n10696));
    jdff dff_A_rT4nJnsx9_1(.din(n10696), .dout(n10693));
    jdff dff_A_HOvEmfsF0_0(.din(n361), .dout(n10690));
    jdff dff_A_eLh1wXtP2_0(.din(n10690), .dout(n10687));
    jdff dff_A_MjqUp2IV7_0(.din(n667), .dout(n10684));
    jdff dff_B_pauv6il10_1(.din(n651), .dout(n10682));
    jdff dff_B_HzC0cx2C7_1(.din(n691), .dout(n10679));
    jdff dff_A_PfzZNePP1_0(.din(G33), .dout(n10675));
    jdff dff_A_oJvYPEnJ3_0(.din(G107), .dout(n10672));
    jdff dff_A_wQjxCHQ43_0(.din(n10672), .dout(n10669));
    jdff dff_A_uORXY95T9_0(.din(n10669), .dout(n10666));
    jdff dff_A_iaCFZwZi5_0(.din(n10666), .dout(n10663));
    jdff dff_A_FREIkpu59_0(.din(n10663), .dout(n10660));
    jdff dff_A_xsnjI4353_0(.din(n10660), .dout(n10657));
    jdff dff_B_ZgjgcbpT5_2(.din(n10652), .dout(n10655));
    jdff dff_B_bwUjs0ls1_2(.din(n743), .dout(n10652));
    jdff dff_A_WUSlaZ817_2(.din(G77), .dout(n10648));
    jdff dff_A_oAMkPFud9_2(.din(n10648), .dout(n10645));
    jdff dff_A_7RCLjyTf9_2(.din(n10645), .dout(n10642));
    jdff dff_A_pllA2Bln3_2(.din(n10642), .dout(n10639));
    jdff dff_A_ByuNwsEG1_0(.din(G77), .dout(n10636));
    jdff dff_A_dfSf8Hys6_0(.din(n10636), .dout(n10633));
    jdff dff_A_DIxhcRxu7_1(.din(n767), .dout(n10630));
    jdff dff_A_Esk9FLPn0_0(.din(n775), .dout(n10627));
    jdff dff_A_v7wVNXzV8_0(.din(n782), .dout(n10624));
    jdff dff_A_EJ8QD03f7_0(.din(n10624), .dout(n10621));
    jdff dff_A_AribFjuc2_0(.din(n792), .dout(n10618));
    jdff dff_B_wdu0KqcM0_1(.din(n785), .dout(n10616));
    jdff dff_B_sT0q3vOJ5_0(.din(n807), .dout(n10613));
    jdff dff_A_nxOb1jX52_1(.din(n11476), .dout(n10609));
    jdff dff_A_ic6VYL2s1_0(.din(n11476), .dout(n10606));
    jdff dff_A_HhEUSmbu4_0(.din(n10606), .dout(n10603));
    jdff dff_A_VJNwAm6t4_0(.din(n10603), .dout(n10600));
    jdff dff_A_5pCyFonK3_1(.din(n216), .dout(n10597));
    jdff dff_A_TxZONEDW8_0(.din(n216), .dout(n10594));
    jdff dff_A_lAM3NFgD3_0(.din(n10594), .dout(n10591));
    jdff dff_A_qbX6Uqo06_0(.din(n10591), .dout(n10588));
    jdff dff_A_KlMvPo997_0(.din(n10588), .dout(n10585));
    jdff dff_B_SP53AS286_2(.din(n823), .dout(n10583));
    jdff dff_A_g5LRjXiN1_0(.din(n10583), .dout(n10579));
    jdff dff_A_Wl9EksWk0_1(.din(n839), .dout(n10576));
    jdff dff_B_E1mUxj7c0_1(.din(n815), .dout(n10574));
    jdff dff_A_iinwmgc79_2(.din(G264), .dout(n10570));
    jdff dff_A_nuy12LkE4_2(.din(n10570), .dout(n10567));
    jdff dff_A_MmzHCcUA0_1(.din(G264), .dout(n10564));
    jdff dff_A_h14eZX9o8_1(.din(n10564), .dout(n10561));
    jdff dff_B_ZbIvEJMZ1_1(.din(n213), .dout(n6419));
    jdff dff_B_RKYEFx1F2_0(.din(n267), .dout(n6422));
    jdff dff_B_XAQHaUNc9_0(.din(n263), .dout(n6425));
    jdff dff_A_35iZO2qL7_1(.din(n6430), .dout(n6427));
    jdff dff_A_vGw5cjWo7_1(.din(n74), .dout(n6430));
    jdff dff_A_QFqMBReo8_0(.din(n165), .dout(n6433));
    jdff dff_B_TiI7vb9P6_1(.din(n1874), .dout(n6437));
    jdff dff_B_57HSYb0W9_0(.din(n2092), .dout(n6440));
    jdff dff_B_gqmF82y40_0(.din(n6440), .dout(n6443));
    jdff dff_B_FqyPStGC8_0(.din(n6443), .dout(n6446));
    jdff dff_B_bR07qUFD3_0(.din(n6446), .dout(n6449));
    jdff dff_B_fekINiU85_0(.din(n6449), .dout(n6452));
    jdff dff_B_FfPOBCUt9_0(.din(n6452), .dout(n6455));
    jdff dff_B_Txu07bCc5_0(.din(n6455), .dout(n6458));
    jdff dff_B_oyBfdrSg1_0(.din(n6458), .dout(n6461));
    jdff dff_B_pnhV1Ahu7_0(.din(n6461), .dout(n6464));
    jdff dff_B_aW8cQsyk1_0(.din(n6464), .dout(n6467));
    jdff dff_B_30hQyZDl3_0(.din(n2088), .dout(n6470));
    jdff dff_B_z4aZpyvY0_0(.din(n2844), .dout(n6473));
    jdff dff_B_r7GeDUeT2_0(.din(n6473), .dout(n6476));
    jdff dff_B_eRMJhjTK0_0(.din(n6476), .dout(n6479));
    jdff dff_B_zRFfzQZT1_0(.din(n6479), .dout(n6482));
    jdff dff_B_GrKdLDr06_0(.din(n6482), .dout(n6485));
    jdff dff_B_wUJghsZH9_0(.din(n6485), .dout(n6488));
    jdff dff_B_KIZG7nLE8_0(.din(n6488), .dout(n6491));
    jdff dff_B_F9VlwxNV5_0(.din(n6491), .dout(n6494));
    jdff dff_B_0prqLHRs9_0(.din(n6494), .dout(n6497));
    jdff dff_B_3vzv6ll53_0(.din(n6497), .dout(n6500));
    jdff dff_B_1o8dJWyL5_0(.din(n6500), .dout(n6503));
    jdff dff_B_iS3n88y91_0(.din(n6503), .dout(n6506));
    jdff dff_B_gRaPGDVy3_0(.din(n6506), .dout(n6509));
    jdff dff_B_3ciAPUTD0_0(.din(n6509), .dout(n6512));
    jdff dff_B_abRt2R1v3_0(.din(n6512), .dout(n6515));
    jdff dff_B_7uld260A0_0(.din(n6515), .dout(n6518));
    jdff dff_B_iHgZDsFN1_0(.din(n6518), .dout(n6521));
    jdff dff_B_S17TyMTG2_1(.din(n2829), .dout(n6524));
    jdff dff_B_ucJF10Ej6_0(.din(n2836), .dout(n6527));
    jdff dff_B_oaMhJkbn7_0(.din(n6527), .dout(n6530));
    jdff dff_B_bgnk8CN45_0(.din(n2801), .dout(n6533));
    jdff dff_B_DiO322YL7_0(.din(n6533), .dout(n6536));
    jdff dff_B_QSAAz7sD6_0(.din(n6536), .dout(n6539));
    jdff dff_B_2phjyk4W1_0(.din(n6539), .dout(n6542));
    jdff dff_B_HKKGKKBb7_0(.din(n6542), .dout(n6545));
    jdff dff_B_slILIBFh7_0(.din(n6545), .dout(n6548));
    jdff dff_B_GnEZZa5h6_0(.din(n6548), .dout(n6551));
    jdff dff_B_2XRZcm3V8_0(.din(n6551), .dout(n6554));
    jdff dff_B_EFk3Y9Tt1_0(.din(n6554), .dout(n6557));
    jdff dff_B_zseAXeDE6_0(.din(n6557), .dout(n6560));
    jdff dff_B_9IuZgE8F7_0(.din(n6560), .dout(n6563));
    jdff dff_B_MpSWbReq4_0(.din(n6563), .dout(n6566));
    jdff dff_B_alibiwfi3_0(.din(n6566), .dout(n6569));
    jdff dff_B_L8rAT8m70_0(.din(n6569), .dout(n6572));
    jdff dff_B_39uXXub01_0(.din(n6572), .dout(n6575));
    jdff dff_B_bLDCNedl5_0(.din(n6575), .dout(n6578));
    jdff dff_B_Q1LIwqe58_0(.din(n6578), .dout(n6581));
    jdff dff_A_pq1kqkUf9_1(.din(n6586), .dout(n6583));
    jdff dff_A_76i7BKoX5_1(.din(n230), .dout(n6586));
    jdff dff_B_INXKO3Aj0_0(.din(n2786), .dout(n6590));
    jdff dff_A_3ErFUkCU3_0(.din(n2783), .dout(n6592));
    jdff dff_B_ismogaiY2_1(.din(n2763), .dout(n6596));
    jdff dff_A_Tqa4XRTQ6_0(.din(n1791), .dout(n6598));
    jdff dff_B_1lyPjolQ8_1(.din(n4308), .dout(n6602));
    jdff dff_B_STSgn9S99_1(.din(n6602), .dout(n6605));
    jdff dff_B_ksuYp0Ct0_1(.din(n6605), .dout(n6608));
    jdff dff_B_cUnlXmVH2_1(.din(n6608), .dout(n6611));
    jdff dff_B_7xWKsNru0_1(.din(n6611), .dout(n6614));
    jdff dff_B_OLwqOrq20_1(.din(n6614), .dout(n6617));
    jdff dff_B_j5kNHohR6_1(.din(n6617), .dout(n6620));
    jdff dff_B_av9rlSH53_1(.din(n6620), .dout(n6623));
    jdff dff_B_CQ4RFwI08_1(.din(n6623), .dout(n6626));
    jdff dff_B_EP064UMY9_1(.din(n6626), .dout(n6629));
    jdff dff_B_6wGLHJU34_1(.din(n6629), .dout(n6632));
    jdff dff_B_vckcHnIO7_1(.din(n6632), .dout(n6635));
    jdff dff_B_FYYw2jGJ6_1(.din(n6635), .dout(n6638));
    jdff dff_B_bIzB3b574_1(.din(n6638), .dout(n6641));
    jdff dff_B_GYgaBrU91_1(.din(n6641), .dout(n6644));
    jdff dff_B_m8yHHaLW0_1(.din(n6644), .dout(n6647));
    jdff dff_B_9dBhZNRm2_1(.din(n6647), .dout(n6650));
    jdff dff_B_ABL8aGuQ4_1(.din(n6650), .dout(n6653));
    jdff dff_B_oD7sEuKY4_1(.din(n6653), .dout(n6656));
    jdff dff_B_0cGMx41z6_1(.din(n6656), .dout(n6659));
    jdff dff_B_e8nhOBiv9_1(.din(n6659), .dout(n6662));
    jdff dff_B_7lWRFK0D9_1(.din(n6662), .dout(n6665));
    jdff dff_B_M7PXAHRb5_1(.din(n6665), .dout(n6668));
    jdff dff_B_PtNcMZnx7_1(.din(n6668), .dout(n6671));
    jdff dff_B_fVe4i1GS5_1(.din(n6671), .dout(n6674));
    jdff dff_B_Dkas4rHc5_1(.din(n6674), .dout(n6677));
    jdff dff_A_1gHWTp1M2_0(.din(n4302), .dout(n6679));
    jdff dff_B_d1iaAPKo4_1(.din(n4278), .dout(n6683));
    jdff dff_B_F6HiktET4_1(.din(n6683), .dout(n6686));
    jdff dff_B_Itre6EaQ7_1(.din(n4354), .dout(n6689));
    jdff dff_B_WPTFmLO94_1(.din(n6689), .dout(n6692));
    jdff dff_B_0KnA5P1y8_1(.din(n6692), .dout(n6695));
    jdff dff_B_qKV9czAu7_1(.din(n6695), .dout(n6698));
    jdff dff_B_S7POIotw4_1(.din(n6698), .dout(n6701));
    jdff dff_B_KGURSiXD8_1(.din(n6701), .dout(n6704));
    jdff dff_B_71sAdNul4_1(.din(n6704), .dout(n6707));
    jdff dff_B_oMD68yai7_1(.din(n6707), .dout(n6710));
    jdff dff_B_ow1ivQgc4_1(.din(n6710), .dout(n6713));
    jdff dff_B_Yw4TcDea7_1(.din(n6713), .dout(n6716));
    jdff dff_B_xRYm96vM2_1(.din(n6716), .dout(n6719));
    jdff dff_B_eUB6iv2E4_1(.din(n6719), .dout(n6722));
    jdff dff_B_cEsRtduB3_1(.din(n6722), .dout(n6725));
    jdff dff_B_8nXiF0Vw6_1(.din(n6725), .dout(n6728));
    jdff dff_B_srSpfLWX5_1(.din(n6728), .dout(n6731));
    jdff dff_B_aaCjEMMh1_1(.din(n6731), .dout(n6734));
    jdff dff_B_3XkVdb4L2_1(.din(n6734), .dout(n6737));
    jdff dff_B_haZlQY2K5_1(.din(n6737), .dout(n6740));
    jdff dff_B_eHtJxHqZ6_1(.din(n6740), .dout(n6743));
    jdff dff_B_atyYGVVP2_1(.din(n6743), .dout(n6746));
    jdff dff_B_GBCDlgHM7_1(.din(n6746), .dout(n6749));
    jdff dff_B_PNjCKbEy0_1(.din(n6749), .dout(n6752));
    jdff dff_B_nNzt09gq4_1(.din(n6752), .dout(n6755));
    jdff dff_B_nr9EUWKf8_1(.din(G2897), .dout(n6758));
    jdff dff_B_HoUtMLY20_1(.din(n6758), .dout(n6761));
    jdff dff_B_Tn5Dfvsh7_1(.din(n6761), .dout(n6764));
    jdff dff_A_FkrEWMOn2_0(.din(n6769), .dout(n6766));
    jdff dff_A_i13Nxk1d4_0(.din(n6772), .dout(n6769));
    jdff dff_A_wMshBjsY8_0(.din(n6775), .dout(n6772));
    jdff dff_A_elJ3kVjw5_0(.din(n6778), .dout(n6775));
    jdff dff_A_LXcfYMdX0_0(.din(n6781), .dout(n6778));
    jdff dff_A_0OlSHuzH1_0(.din(n6784), .dout(n6781));
    jdff dff_A_8XzyIIqw3_0(.din(n6787), .dout(n6784));
    jdff dff_A_7aIAM5uW5_0(.din(n6790), .dout(n6787));
    jdff dff_A_JX7QnrZu6_0(.din(n6793), .dout(n6790));
    jdff dff_A_YYX4gCcC9_0(.din(n6796), .dout(n6793));
    jdff dff_A_ezIhfjT26_0(.din(n6799), .dout(n6796));
    jdff dff_A_EinBL5jg3_0(.din(n6802), .dout(n6799));
    jdff dff_A_fWezhZQK1_0(.din(n6805), .dout(n6802));
    jdff dff_A_pyHyVM520_0(.din(n6808), .dout(n6805));
    jdff dff_A_uTB02lxm3_0(.din(n6811), .dout(n6808));
    jdff dff_A_Czfwup3U9_0(.din(n6814), .dout(n6811));
    jdff dff_A_s2qmCIG71_0(.din(n6817), .dout(n6814));
    jdff dff_A_fLRtkNEI5_0(.din(n6820), .dout(n6817));
    jdff dff_A_QiWqXZtD8_0(.din(n6823), .dout(n6820));
    jdff dff_A_hlIfiqL39_0(.din(n6826), .dout(n6823));
    jdff dff_A_wZ6b6fHU0_0(.din(n6829), .dout(n6826));
    jdff dff_A_0WDg3HZv0_0(.din(n6832), .dout(n6829));
    jdff dff_A_ED2r026o9_0(.din(n6835), .dout(n6832));
    jdff dff_A_2gFj4f353_0(.din(n4347), .dout(n6835));
    jdff dff_A_CUINI1G20_1(.din(n6841), .dout(n6838));
    jdff dff_A_qG5g4Kdt6_1(.din(n6844), .dout(n6841));
    jdff dff_A_VKYtCPlx4_1(.din(n6847), .dout(n6844));
    jdff dff_A_KWqK4jsg9_1(.din(n6850), .dout(n6847));
    jdff dff_A_fSoq5eSk9_1(.din(n6853), .dout(n6850));
    jdff dff_A_2RZGnjge1_1(.din(n6856), .dout(n6853));
    jdff dff_A_jlR3c4od4_1(.din(n6859), .dout(n6856));
    jdff dff_A_YbRQWkiM0_1(.din(n6862), .dout(n6859));
    jdff dff_A_LpgbsOwJ3_1(.din(n6865), .dout(n6862));
    jdff dff_A_HkHWyVHQ7_1(.din(n6868), .dout(n6865));
    jdff dff_A_bPrk78ai6_1(.din(n6871), .dout(n6868));
    jdff dff_A_RwyT5Put4_1(.din(n6874), .dout(n6871));
    jdff dff_A_BSkzwkY28_1(.din(n6877), .dout(n6874));
    jdff dff_A_GYfWShQb6_1(.din(n6880), .dout(n6877));
    jdff dff_A_9sO4ZTmB4_1(.din(n6883), .dout(n6880));
    jdff dff_A_EAUOJHMP3_1(.din(n6886), .dout(n6883));
    jdff dff_A_hjlqjJGa8_1(.din(n6889), .dout(n6886));
    jdff dff_A_WW1YB6Nx9_1(.din(n6892), .dout(n6889));
    jdff dff_A_6kQ4PVCa9_1(.din(n6895), .dout(n6892));
    jdff dff_A_UnE89SV35_1(.din(n6898), .dout(n6895));
    jdff dff_A_TwVIFBZk6_1(.din(n6901), .dout(n6898));
    jdff dff_A_BVhJRhXi2_1(.din(n6904), .dout(n6901));
    jdff dff_A_2P7m60Fo7_1(.din(n6907), .dout(n6904));
    jdff dff_A_TkG7pfVH7_1(.din(n6910), .dout(n6907));
    jdff dff_A_PBO6IMgf3_1(.din(n4311), .dout(n6910));
    jdff dff_A_75qdFNfU4_0(.din(n4358), .dout(n6913));
    jdff dff_B_DVFnj4U50_1(.din(n3871), .dout(n6917));
    jdff dff_B_kjZczfGZ9_0(.din(n4071), .dout(n6920));
    jdff dff_B_z9x0sSSx3_0(.din(n6920), .dout(n6923));
    jdff dff_B_mueMJx3S2_0(.din(n6923), .dout(n6926));
    jdff dff_B_krCILoBk6_0(.din(n6926), .dout(n6929));
    jdff dff_B_7VYOSbKx5_0(.din(n6929), .dout(n6932));
    jdff dff_B_H8cVUlWX9_0(.din(n6932), .dout(n6935));
    jdff dff_B_KyoqtR4A7_0(.din(n4067), .dout(n6938));
    jdff dff_B_92gJze930_0(.din(n6938), .dout(n6941));
    jdff dff_B_8BSMLYpj6_0(.din(n4063), .dout(n6944));
    jdff dff_B_9ILQ2W4v2_0(.din(n6944), .dout(n6947));
    jdff dff_B_S2QAhHBW2_0(.din(n6947), .dout(n6950));
    jdff dff_B_uRmScwGU2_0(.din(n6950), .dout(n6953));
    jdff dff_B_fS9LehUH7_0(.din(n6953), .dout(n6956));
    jdff dff_B_wBzgC1T75_0(.din(n4059), .dout(n6959));
    jdff dff_B_ROu9VDUx5_0(.din(n6959), .dout(n6962));
    jdff dff_B_2cDIwnZe2_1(.din(n3893), .dout(n6965));
    jdff dff_B_oF2J7WMc8_1(.din(n6965), .dout(n6968));
    jdff dff_B_SsjTCZ8P9_1(.din(n6968), .dout(n6971));
    jdff dff_B_bhAskbXh4_1(.din(n6971), .dout(n6974));
    jdff dff_B_BtmoNtxU2_1(.din(n6974), .dout(n6977));
    jdff dff_B_x9p7lb4a7_1(.din(n6977), .dout(n6980));
    jdff dff_B_IP1rCXvj1_1(.din(n6980), .dout(n6983));
    jdff dff_B_PeH7jio82_1(.din(n6983), .dout(n6986));
    jdff dff_B_VB52pyBY9_1(.din(n3970), .dout(n6989));
    jdff dff_B_qrhrT4zO7_0(.din(n4043), .dout(n6992));
    jdff dff_B_MQBvZFPF6_0(.din(n6992), .dout(n6995));
    jdff dff_B_LIftqJ252_0(.din(n6995), .dout(n6998));
    jdff dff_B_71J1ASuV1_0(.din(n6998), .dout(n7001));
    jdff dff_B_wH6kjyXK3_0(.din(n7001), .dout(n7004));
    jdff dff_B_snN3B2LV6_0(.din(n7004), .dout(n7007));
    jdff dff_B_LYXjIAr02_0(.din(n7007), .dout(n7010));
    jdff dff_B_7iHYmG9Z8_0(.din(n7010), .dout(n7013));
    jdff dff_B_l64JFMp40_1(.din(n3993), .dout(n7016));
    jdff dff_B_gLKpy3Be3_1(.din(n4008), .dout(n7019));
    jdff dff_B_NepKsP0S7_1(.din(n7019), .dout(n7022));
    jdff dff_B_hNlRGnM00_0(.din(n4020), .dout(n7025));
    jdff dff_B_W0sNcPpq6_0(.din(n4004), .dout(n7028));
    jdff dff_B_j0Bgs2dV7_0(.din(n7028), .dout(n7031));
    jdff dff_B_5S8Al6CO4_0(.din(n7031), .dout(n7034));
    jdff dff_B_NtJjTnVt0_1(.din(n3974), .dout(n7037));
    jdff dff_B_YsUganJu0_1(.din(n7037), .dout(n7040));
    jdff dff_B_HVAqcWer1_0(.din(n3982), .dout(n7043));
    jdff dff_B_TFXDdaWy7_1(.din(n3916), .dout(n7046));
    jdff dff_B_SFjiaPKT8_1(.din(n7046), .dout(n7049));
    jdff dff_B_ggGMsJUX2_1(.din(n3931), .dout(n7052));
    jdff dff_B_eJtHe2Jq2_1(.din(G124), .dout(n7055));
    jdff dff_B_10xCu5ic8_1(.din(n7055), .dout(n7058));
    jdff dff_B_9YDK52XL0_1(.din(n7058), .dout(n7061));
    jdff dff_B_vnVczlSn4_1(.din(n7061), .dout(n7064));
    jdff dff_B_EG6ARHJv1_1(.din(n3935), .dout(n7067));
    jdff dff_B_dYravbQS3_0(.din(n3927), .dout(n7070));
    jdff dff_B_7XdmRs1Y7_0(.din(n7070), .dout(n7073));
    jdff dff_B_AVUazYlt7_0(.din(n7073), .dout(n7076));
    jdff dff_B_dtJPXaif5_0(.din(n7076), .dout(n7079));
    jdff dff_B_9uif3c2I5_1(.din(n3897), .dout(n7082));
    jdff dff_B_qMUJgFx84_1(.din(n3874), .dout(n7085));
    jdff dff_B_MqphnD900_1(.din(n3837), .dout(n7088));
    jdff dff_B_XlWbM8QL0_1(.din(n7088), .dout(n7091));
    jdff dff_B_d1NIOL8X8_1(.din(n7091), .dout(n7094));
    jdff dff_A_RZtshrj92_1(.din(n7099), .dout(n7096));
    jdff dff_A_Xxqvm21W1_1(.din(n7102), .dout(n7099));
    jdff dff_A_j760mmVa3_1(.din(n7105), .dout(n7102));
    jdff dff_A_6aGBmUHX2_1(.din(n7108), .dout(n7105));
    jdff dff_A_gRcrxL502_1(.din(n3859), .dout(n7108));
    jdff dff_A_qQrMKb5R0_0(.din(n3841), .dout(n7111));
    jdff dff_B_1vL66lyp4_1(.din(n2682), .dout(n7115));
    jdff dff_B_C7ktbf3h3_1(.din(n7115), .dout(n7118));
    jdff dff_B_cRQJmgxW2_1(.din(n7118), .dout(n7121));
    jdff dff_B_66AscVry2_1(.din(n7121), .dout(n7124));
    jdff dff_B_tqzWkzFC0_1(.din(n7124), .dout(n7127));
    jdff dff_B_vGoV2cZb0_1(.din(n7127), .dout(n7130));
    jdff dff_A_5Tgp0F3a0_1(.din(n7135), .dout(n7132));
    jdff dff_A_kExtFxnH9_1(.din(n7138), .dout(n7135));
    jdff dff_A_XQEGH7Fg5_1(.din(n7264), .dout(n7138));
    jdff dff_B_tAnG3rFH9_0(.din(n2678), .dout(n7142));
    jdff dff_B_ROk0rJVR8_0(.din(n7142), .dout(n7145));
    jdff dff_B_sGAdXcQK9_0(.din(n7145), .dout(n7148));
    jdff dff_B_u9jzawup9_0(.din(n7148), .dout(n7151));
    jdff dff_B_ttQFE8Zp5_0(.din(n7151), .dout(n7154));
    jdff dff_B_OFsKvyEN6_0(.din(n7154), .dout(n7157));
    jdff dff_B_lsqKqCwg4_0(.din(n7157), .dout(n7160));
    jdff dff_B_Au4qUoU05_0(.din(n7160), .dout(n7163));
    jdff dff_A_WJXeNyEx8_0(.din(n7168), .dout(n7165));
    jdff dff_A_pbWzgCyS4_0(.din(n3830), .dout(n7168));
    jdff dff_A_pSs0Kn2T5_1(.din(n7174), .dout(n7171));
    jdff dff_A_qpemC9y70_1(.din(n3830), .dout(n7174));
    jdff dff_B_SWbG8yOW4_0(.din(n3826), .dout(n7178));
    jdff dff_B_Nrqi0ynE4_0(.din(n3822), .dout(n7181));
    jdff dff_B_tjgyHJ106_0(.din(n3815), .dout(n7184));
    jdff dff_B_DjOAi9Nd9_0(.din(n7184), .dout(n7187));
    jdff dff_B_QcnaCo5a3_0(.din(n7187), .dout(n7190));
    jdff dff_B_eAU6ZNs84_0(.din(n7190), .dout(n7193));
    jdff dff_B_VwXBFnol2_0(.din(n7193), .dout(n7196));
    jdff dff_B_2ViURvvM0_0(.din(n3811), .dout(n7199));
    jdff dff_B_v7qJ2qFU7_0(.din(n7199), .dout(n7202));
    jdff dff_B_l6gt4ru40_0(.din(n3804), .dout(n7205));
    jdff dff_B_LwLodLqI6_0(.din(n7205), .dout(n7208));
    jdff dff_B_Af0sdr0X2_1(.din(n3756), .dout(n7211));
    jdff dff_B_vXFnbtG86_1(.din(n3764), .dout(n7214));
    jdff dff_B_TQP1YUm59_1(.din(n7214), .dout(n7217));
    jdff dff_B_RP8VEQR27_1(.din(n3776), .dout(n7220));
    jdff dff_B_86zZpgHb2_1(.din(n3744), .dout(n7223));
    jdff dff_B_M3Zz5C7m8_0(.din(n3748), .dout(n7226));
    jdff dff_B_RFjhdhla7_1(.din(n3696), .dout(n7229));
    jdff dff_B_yGPfwFgA3_1(.din(n3704), .dout(n7232));
    jdff dff_B_wFxVZoM59_1(.din(n3716), .dout(n7235));
    jdff dff_B_0MkERJX76_1(.din(n3720), .dout(n7238));
    jdff dff_B_fUpwtMpE7_1(.din(n3680), .dout(n7241));
    jdff dff_B_UOaAKzrk5_0(.din(n3688), .dout(n7244));
    jdff dff_A_xsEWv84P2_1(.din(n7256), .dout(n7246));
    jdff dff_B_HHCElp5e4_2(.din(G125), .dout(n7250));
    jdff dff_B_G86RNpOp3_2(.din(n7250), .dout(n7253));
    jdff dff_B_p5Pr9xfC7_2(.din(n7253), .dout(n7256));
    jdff dff_A_slKm5Ewo6_1(.din(n7261), .dout(n7258));
    jdff dff_A_7FpSlnU95_1(.din(n3599), .dout(n7261));
    jdff dff_A_wMvQFKzl8_0(.din(n2701), .dout(n7264));
    jdff dff_A_hOWFdUb55_1(.din(n7270), .dout(n7267));
    jdff dff_A_MmctwkeV4_1(.din(n7273), .dout(n7270));
    jdff dff_A_qmBZvkLz6_1(.din(n2701), .dout(n7273));
    jdff dff_A_7ay8bsDi0_0(.din(n2686), .dout(n7276));
    jdff dff_B_BXD6qlQV4_0(.din(n2740), .dout(n7280));
    jdff dff_B_WgF3nB0b5_0(.din(n2736), .dout(n7283));
    jdff dff_B_gPf7eztG3_0(.din(n7283), .dout(n7286));
    jdff dff_B_YDYslqhf5_0(.din(n7286), .dout(n7289));
    jdff dff_A_pnr9ZWDy8_2(.din(n7294), .dout(n7291));
    jdff dff_A_FQjyNBXB6_2(.din(n2724), .dout(n7294));
    jdff dff_A_mU4FV3g02_1(.din(n4343), .dout(n7297));
    jdff dff_B_3exNftqn2_1(.din(n4327), .dout(n7301));
    jdff dff_B_mMffx1gt7_1(.din(n7301), .dout(n7304));
    jdff dff_B_sSNfvP074_1(.din(n4331), .dout(n7307));
    jdff dff_B_V1j9SyVP8_1(.din(n7307), .dout(n7310));
    jdff dff_B_nePEl5Xx0_1(.din(n7310), .dout(n7313));
    jdff dff_A_Cy2pFh2x2_0(.din(n7318), .dout(n7315));
    jdff dff_A_fyeVzkVI3_0(.din(n3593), .dout(n7318));
    jdff dff_A_O5BkJj945_1(.din(n3593), .dout(n7321));
    jdff dff_B_Cx17UkaA4_0(.din(n3585), .dout(n7325));
    jdff dff_B_fRdCpgyv1_0(.din(n7325), .dout(n7328));
    jdff dff_B_c6pRVtlX6_0(.din(n3578), .dout(n7331));
    jdff dff_B_2JuQXva06_0(.din(n7331), .dout(n7334));
    jdff dff_B_n3TuTuIJ8_0(.din(n7334), .dout(n7337));
    jdff dff_B_aNkwzhXz0_0(.din(n7337), .dout(n7340));
    jdff dff_B_M8nSWbet7_0(.din(n3574), .dout(n7343));
    jdff dff_B_rDa61NF65_0(.din(n7343), .dout(n7346));
    jdff dff_B_0avh9kPH0_1(.din(n3558), .dout(n7349));
    jdff dff_B_XvEe2tqO0_1(.din(n7349), .dout(n7352));
    jdff dff_B_Lb7neYNf5_0(.din(n3562), .dout(n7355));
    jdff dff_A_jQ6iCYFb7_2(.din(n11194), .dout(n7357));
    jdff dff_B_C5qcIsB09_2(.din(n336), .dout(n7361));
    jdff dff_B_MvjVfA9W0_1(.din(n328), .dout(n7364));
    jdff dff_B_ywj6lkni5_1(.din(n3506), .dout(n7367));
    jdff dff_B_whVeXqgD6_1(.din(n3514), .dout(n7370));
    jdff dff_B_WnjYk9sv3_1(.din(n3526), .dout(n7373));
    jdff dff_B_q2pNGgEz9_0(.din(n3530), .dout(n7376));
    jdff dff_A_PQFRbtVo2_0(.din(n8864), .dout(n7378));
    jdff dff_A_qQppqKnn2_2(.din(n8864), .dout(n7381));
    jdff dff_A_hfLMMskf5_1(.din(n7387), .dout(n7384));
    jdff dff_A_WWK0B2oo7_1(.din(n7390), .dout(n7387));
    jdff dff_A_FEpwPMUa3_1(.din(n7393), .dout(n7390));
    jdff dff_A_sVwYQHnY4_1(.din(n11452), .dout(n7393));
    jdff dff_A_mp6aKalC4_2(.din(n7399), .dout(n7396));
    jdff dff_A_gdXVBH7B5_2(.din(n7402), .dout(n7399));
    jdff dff_A_acilBIRd4_2(.din(n7405), .dout(n7402));
    jdff dff_A_yjpnAqiE4_2(.din(n11452), .dout(n7405));
    jdff dff_B_QnFifl5M3_0(.din(n3498), .dout(n7409));
    jdff dff_A_snOCCsqR1_1(.din(n3490), .dout(n7411));
    jdff dff_B_HzyL4HYi9_1(.din(n3446), .dout(n7415));
    jdff dff_B_OhcYGMIq1_1(.din(n3454), .dout(n7418));
    jdff dff_B_ByV9zlj97_1(.din(n3466), .dout(n7421));
    jdff dff_B_VJfuxWIR1_0(.din(n3470), .dout(n7424));
    jdff dff_B_AOeF9rv66_1(.din(n3430), .dout(n7427));
    jdff dff_B_8j7u9TlS3_0(.din(n3438), .dout(n7430));
    jdff dff_A_lgUsyUaz7_0(.din(n7435), .dout(n7432));
    jdff dff_A_Qfqo2AYs7_0(.din(n7438), .dout(n7435));
    jdff dff_A_P4ZigKiT8_0(.din(n9448), .dout(n7438));
    jdff dff_B_FStJrMIY0_1(.din(n3056), .dout(n7442));
    jdff dff_B_NmMHFuky2_1(.din(n7442), .dout(n7445));
    jdff dff_B_sHP7iWLK0_1(.din(n7445), .dout(n7448));
    jdff dff_B_Un1tSFFn9_1(.din(n7448), .dout(n7451));
    jdff dff_B_sdMd6HLu4_1(.din(n7451), .dout(n7454));
    jdff dff_B_eRk8zz767_1(.din(n7454), .dout(n7457));
    jdff dff_B_YYMkNhYA5_0(.din(n3150), .dout(n7460));
    jdff dff_B_roZoaxUK5_0(.din(n7460), .dout(n7463));
    jdff dff_B_6Fz6g5cU3_1(.din(n3135), .dout(n7466));
    jdff dff_B_xvuZQWgj8_1(.din(n3124), .dout(n7469));
    jdff dff_B_9rSm278z7_1(.din(n7469), .dout(n7472));
    jdff dff_B_Iti47Lbc7_1(.din(n7472), .dout(n7475));
    jdff dff_B_84D6kbgx2_1(.din(n7475), .dout(n7478));
    jdff dff_B_8swdFZdK9_1(.din(n7478), .dout(n7481));
    jdff dff_A_dgcepEnl3_1(.din(n7486), .dout(n7483));
    jdff dff_A_RyHrEmPo5_1(.din(n3096), .dout(n7486));
    jdff dff_A_rwQYYhjr9_2(.din(n7492), .dout(n7489));
    jdff dff_A_R0rFJcId8_2(.din(n3096), .dout(n7492));
    jdff dff_B_2jr7qtF45_0(.din(n3092), .dout(n7496));
    jdff dff_B_ZbbISUN88_0(.din(n3081), .dout(n7499));
    jdff dff_B_Sq1nVs155_0(.din(n7499), .dout(n7502));
    jdff dff_B_WuxO66pk5_0(.din(n7502), .dout(n7505));
    jdff dff_A_vBAbKGaa3_1(.din(n7510), .dout(n7507));
    jdff dff_A_phdcRowx4_1(.din(n1962), .dout(n7510));
    jdff dff_A_6IF8HUCr3_2(.din(n7516), .dout(n7513));
    jdff dff_A_qh0ueVTK0_2(.din(n1962), .dout(n7516));
    jdff dff_B_OEX3IkGW5_1(.din(n1931), .dout(n7520));
    jdff dff_B_O1xqApWe3_1(.din(n7520), .dout(n7523));
    jdff dff_B_76bfDyqF7_1(.din(n7523), .dout(n7526));
    jdff dff_B_mxVotttX4_0(.din(n3052), .dout(n7529));
    jdff dff_B_vakdpU0h4_0(.din(n7529), .dout(n7532));
    jdff dff_B_waiU3iPW9_0(.din(n3048), .dout(n7535));
    jdff dff_B_8GtkNEO43_0(.din(n7535), .dout(n7538));
    jdff dff_B_0dxtSe3b5_0(.din(n7538), .dout(n7541));
    jdff dff_B_XK9Rr1Md4_0(.din(n7541), .dout(n7544));
    jdff dff_B_HGegVXfg3_1(.din(n3032), .dout(n7547));
    jdff dff_B_EkAG2G5A5_1(.din(n7547), .dout(n7550));
    jdff dff_B_cNBDWlkf7_0(.din(n3036), .dout(n7553));
    jdff dff_A_6vLKW1ti3_0(.din(n287), .dout(n7555));
    jdff dff_B_dBwvH5b50_1(.din(n279), .dout(n7559));
    jdff dff_B_ZsphsNXi2_1(.din(n2941), .dout(n7562));
    jdff dff_B_9EpyEEZg7_1(.din(n7562), .dout(n7565));
    jdff dff_B_tafiDLO83_1(.din(n2970), .dout(n7568));
    jdff dff_B_E9q2u0Q57_1(.din(n2978), .dout(n7571));
    jdff dff_B_l1n21D5a6_1(.din(n7571), .dout(n7574));
    jdff dff_B_KfVTBMJA0_1(.din(n2990), .dout(n7577));
    jdff dff_B_GOaq4DFZ9_1(.din(n2994), .dout(n7580));
    jdff dff_B_Xkqgtt0R2_1(.din(n2948), .dout(n7583));
    jdff dff_B_qpC0aZAa8_1(.din(n2897), .dout(n7586));
    jdff dff_B_kG1WRgHS8_1(.din(n2905), .dout(n7589));
    jdff dff_B_TTOk1bak3_1(.din(n2917), .dout(n7592));
    jdff dff_B_LAJJ92v23_1(.din(n2921), .dout(n7595));
    jdff dff_B_liQ1UMAM7_1(.din(n2881), .dout(n7598));
    jdff dff_B_5f1pzdeI0_0(.din(n2889), .dout(n7601));
    jdff dff_A_bwpleDz36_2(.din(n11059), .dout(n7603));
    jdff dff_A_TdwTkyIG6_0(.din(n7609), .dout(n7606));
    jdff dff_A_eYQCiEqf0_0(.din(n7612), .dout(n7609));
    jdff dff_A_LTfKkiCi8_0(.din(n7615), .dout(n7612));
    jdff dff_A_4UiU7fNk1_0(.din(n2867), .dout(n7615));
    jdff dff_B_N4HDd12h4_0(.din(n2863), .dout(n7619));
    jdff dff_B_O0aVY1Bz7_0(.din(n2855), .dout(n7622));
    jdff dff_A_JPVkXb1c2_0(.din(n2852), .dout(n7624));
    jdff dff_B_SiD7b9u99_0(.din(n3390), .dout(n7628));
    jdff dff_B_afRYyTAp2_0(.din(n7628), .dout(n7631));
    jdff dff_B_VXjngd2T1_0(.din(n3386), .dout(n7634));
    jdff dff_B_ZNbBFqDO1_0(.din(n3382), .dout(n7637));
    jdff dff_B_Nw4q9f9k2_0(.din(n7637), .dout(n7640));
    jdff dff_B_lUDGU5Tm8_1(.din(n3345), .dout(n7643));
    jdff dff_B_l03SnlX31_1(.din(n3349), .dout(n7646));
    jdff dff_B_qd4Dr2xX7_1(.din(n3314), .dout(n7649));
    jdff dff_B_YfOZGs5a8_1(.din(n7649), .dout(n7652));
    jdff dff_B_1EorlipC6_1(.din(n3321), .dout(n7655));
    jdff dff_A_6VDFVZtn3_1(.din(n77), .dout(n7657));
    jdff dff_A_Eux4reDN6_1(.din(n302), .dout(n7660));
    jdff dff_B_hpJU5pAe0_1(.din(n294), .dout(n7664));
    jdff dff_B_y8ZMZmyl1_1(.din(n3258), .dout(n7667));
    jdff dff_B_dTs5iTOn6_1(.din(n3266), .dout(n7670));
    jdff dff_B_40pmEBcG8_1(.din(n3278), .dout(n7673));
    jdff dff_B_ywfEaQGJ9_1(.din(n3282), .dout(n7676));
    jdff dff_A_Atnr6eaZ2_0(.din(n8941), .dout(n7678));
    jdff dff_A_u6lMMEG02_1(.din(n7684), .dout(n7681));
    jdff dff_A_JEUNizrH2_1(.din(n7687), .dout(n7684));
    jdff dff_A_uiOC0J294_1(.din(G68), .dout(n7687));
    jdff dff_A_f2WoVYay3_2(.din(n7693), .dout(n7690));
    jdff dff_A_4ndtRwkk5_2(.din(n7696), .dout(n7693));
    jdff dff_A_YzKwCjno0_2(.din(n7699), .dout(n7696));
    jdff dff_A_6KVDIPDC3_2(.din(G68), .dout(n7699));
    jdff dff_A_UaieZtxF1_1(.din(n9001), .dout(n7702));
    jdff dff_B_fkrlfE7F9_0(.din(n3250), .dout(n7706));
    jdff dff_A_rBK6NEAD6_0(.din(n7711), .dout(n7708));
    jdff dff_A_n8CIkRW42_0(.din(n9880), .dout(n7711));
    jdff dff_A_05j5Fhvw0_2(.din(n7717), .dout(n7714));
    jdff dff_A_JtTPq6K41_2(.din(n9880), .dout(n7717));
    jdff dff_B_s3dYIOLe0_1(.din(n3198), .dout(n7721));
    jdff dff_B_t8HqBvIk0_1(.din(n3206), .dout(n7724));
    jdff dff_B_ijOsRv3d3_0(.din(n3230), .dout(n7727));
    jdff dff_B_oAB1G1BA4_0(.din(n3214), .dout(n7730));
    jdff dff_A_nFcxiCu25_1(.din(n11338), .dout(n7732));
    jdff dff_A_Ig1MTnX10_2(.din(n11338), .dout(n7735));
    jdff dff_B_C8F25GoX1_1(.din(n3182), .dout(n7739));
    jdff dff_B_ArWb2Guz8_0(.din(n3190), .dout(n7742));
    jdff dff_A_KSVncrO02_0(.din(n10783), .dout(n7744));
    jdff dff_A_cOYiOvKk8_1(.din(n10783), .dout(n7747));
    jdff dff_A_XSZpSyWq1_1(.din(n1965), .dout(n7750));
    jdff dff_B_GWUvgwss7_1(.din(n3162), .dout(n7754));
    jdff dff_B_CQS8NZev0_1(.din(n7754), .dout(n7757));
    jdff dff_A_TtFrPdwf5_0(.din(n7762), .dout(n7759));
    jdff dff_A_4OJKC0OR5_0(.din(n7765), .dout(n7762));
    jdff dff_A_0YiUR0Ss4_0(.din(n2061), .dout(n7765));
    jdff dff_A_PXFsuTRE2_0(.din(n7771), .dout(n7768));
    jdff dff_A_8VaEDlcY7_0(.din(n9580), .dout(n7771));
    jdff dff_A_Iq24XGYr3_1(.din(n9580), .dout(n7774));
    jdff dff_B_SYCE2BTn7_0(.din(n3063), .dout(n7778));
    jdff dff_B_IQmQYXWB0_0(.din(n1950), .dout(n7781));
    jdff dff_B_q1yVKbPA9_2(.din(n1935), .dout(n7784));
    jdff dff_B_6XuEDFwA5_2(.din(n7784), .dout(n7787));
    jdff dff_A_lRlMu4sD7_0(.din(n7792), .dout(n7789));
    jdff dff_A_M0tghYyO0_0(.din(n7795), .dout(n7792));
    jdff dff_A_i1S5ziKV7_0(.din(n2444), .dout(n7795));
    jdff dff_B_Ks7agVIe9_0(.din(n2436), .dout(n7799));
    jdff dff_B_pbid71fM7_0(.din(n7799), .dout(n7802));
    jdff dff_B_t2vIVQ5S6_0(.din(n2432), .dout(n7805));
    jdff dff_B_ijCClu5V1_0(.din(n7805), .dout(n7808));
    jdff dff_B_TgwTAz0T8_1(.din(n2401), .dout(n7811));
    jdff dff_B_PrSaw47k1_1(.din(n2405), .dout(n7814));
    jdff dff_B_wnaAccVc0_2(.din(n2409), .dout(n7817));
    jdff dff_B_tSC1lAtp1_1(.din(n2382), .dout(n7820));
    jdff dff_B_q8O96NZW0_1(.din(n7820), .dout(n7823));
    jdff dff_B_aPhNAm609_0(.din(n317), .dout(n7826));
    jdff dff_A_Hu6cMehe4_1(.din(n7831), .dout(n7828));
    jdff dff_A_lbvI5AZX7_1(.din(n7834), .dout(n7831));
    jdff dff_A_7SeFFzao1_1(.din(n2378), .dout(n7834));
    jdff dff_A_DMFkWSl72_2(.din(n7840), .dout(n7837));
    jdff dff_A_ndWtT0954_2(.din(n7843), .dout(n7840));
    jdff dff_A_s4K4jVzF7_2(.din(n2378), .dout(n7843));
    jdff dff_B_WR5Qgovz9_1(.din(n2284), .dout(n7847));
    jdff dff_B_SollERH45_1(.din(n7847), .dout(n7850));
    jdff dff_B_DUUwAbIW3_1(.din(n2307), .dout(n7853));
    jdff dff_B_JOmrejZn1_1(.din(n7853), .dout(n7856));
    jdff dff_B_NFw4p7kh4_1(.din(n2318), .dout(n7859));
    jdff dff_B_cnEI5OKQ2_1(.din(n2334), .dout(n7862));
    jdff dff_B_fNJBprkP0_0(.din(n2326), .dout(n7865));
    jdff dff_B_zytjr5lS4_1(.din(n2216), .dout(n7868));
    jdff dff_B_YeRo1S9M1_1(.din(n2228), .dout(n7871));
    jdff dff_B_xbbZLR3d2_0(.din(n2272), .dout(n7874));
    jdff dff_A_WorGWE6A7_0(.din(n7886), .dout(n7876));
    jdff dff_B_A1KkwWH95_3(.din(G317), .dout(n7880));
    jdff dff_B_3ApFXNkh1_3(.din(n7880), .dout(n7883));
    jdff dff_B_shLEtSI70_3(.din(n7883), .dout(n7886));
    jdff dff_A_U500Ob7a2_0(.din(n7898), .dout(n7888));
    jdff dff_B_8nMucfrd1_2(.din(G326), .dout(n7892));
    jdff dff_B_GGu0UJGT6_2(.din(n7892), .dout(n7895));
    jdff dff_B_uJt7CJLp2_2(.din(n7895), .dout(n7898));
    jdff dff_B_HZGkihJZ2_0(.din(n2244), .dout(n7901));
    jdff dff_B_gx73yGy73_1(.din(G329), .dout(n7904));
    jdff dff_B_HFEHj2gJ7_1(.din(n7904), .dout(n7907));
    jdff dff_B_ovBAT9NH3_1(.din(n7907), .dout(n7910));
    jdff dff_B_g3sqqxTD0_1(.din(n7910), .dout(n7913));
    jdff dff_A_zvJHdfOq5_1(.din(n7918), .dout(n7915));
    jdff dff_A_9QZE4nlL5_1(.din(n7921), .dout(n7918));
    jdff dff_A_Z4ls5wLR7_1(.din(n9364), .dout(n7921));
    jdff dff_A_dJDGDyOs2_2(.din(n7927), .dout(n7924));
    jdff dff_A_TLWREQpl6_2(.din(n9364), .dout(n7927));
    jdff dff_B_vPKyQSuR3_1(.din(n2171), .dout(n7931));
    jdff dff_B_luZy6lJH8_0(.din(n2208), .dout(n7934));
    jdff dff_A_2rrUxUIP9_0(.din(n7946), .dout(n7936));
    jdff dff_B_u0neskAZ0_3(.din(G322), .dout(n7940));
    jdff dff_B_bUL5dkCT3_3(.din(n7940), .dout(n7943));
    jdff dff_B_cWNoaYa40_3(.din(n7943), .dout(n7946));
    jdff dff_A_zP6meR3B7_1(.din(n7951), .dout(n7948));
    jdff dff_A_SvGabuyZ0_1(.din(n7954), .dout(n7951));
    jdff dff_A_v4aMslTG5_1(.din(n7957), .dout(n7954));
    jdff dff_A_mEvHV7Qt0_1(.din(n7960), .dout(n7957));
    jdff dff_A_fO1gaAU48_1(.din(n7963), .dout(n7960));
    jdff dff_A_pq2AYniU8_1(.din(n7966), .dout(n7963));
    jdff dff_A_tmTvCkbU6_1(.din(n7969), .dout(n7966));
    jdff dff_A_fKgJXFjY1_1(.din(n8326), .dout(n7969));
    jdff dff_A_YCzhrQoY5_0(.din(n7975), .dout(n7972));
    jdff dff_A_oHrPOyqK9_0(.din(n7978), .dout(n7975));
    jdff dff_A_D8WSjl5f6_0(.din(n7981), .dout(n7978));
    jdff dff_A_Pp5xVGwQ0_0(.din(n7984), .dout(n7981));
    jdff dff_A_SCHK0TrY7_0(.din(n7987), .dout(n7984));
    jdff dff_A_DEZNKbo81_0(.din(n7990), .dout(n7987));
    jdff dff_A_nBl04f0e9_0(.din(n7993), .dout(n7990));
    jdff dff_A_B0I6oQeg1_0(.din(n7996), .dout(n7993));
    jdff dff_A_w0rZFdYh7_0(.din(n7999), .dout(n7996));
    jdff dff_A_mLqKf1by0_0(.din(n8002), .dout(n7999));
    jdff dff_A_TGBdpbH83_0(.din(n2133), .dout(n8002));
    jdff dff_A_OSUnoYmz9_2(.din(n8008), .dout(n8005));
    jdff dff_A_dtUhY7JZ5_2(.din(n8011), .dout(n8008));
    jdff dff_A_tVr9P22h8_2(.din(n8014), .dout(n8011));
    jdff dff_A_6vPwiSX80_2(.din(n8017), .dout(n8014));
    jdff dff_A_iRk3bfpv5_2(.din(n8020), .dout(n8017));
    jdff dff_A_hO7d4Kf21_2(.din(n8023), .dout(n8020));
    jdff dff_A_gqzlGGGV6_2(.din(n8026), .dout(n8023));
    jdff dff_A_yKOyCE6l8_2(.din(n8029), .dout(n8026));
    jdff dff_A_zOV6tKue4_2(.din(n8032), .dout(n8029));
    jdff dff_A_duMeiHOw2_2(.din(n8035), .dout(n8032));
    jdff dff_A_VPwrvW8B8_2(.din(n2133), .dout(n8035));
    jdff dff_A_hmxa8FcC1_1(.din(n8041), .dout(n8038));
    jdff dff_A_vuWhESbr7_1(.din(n8044), .dout(n8041));
    jdff dff_A_9ANYxGzJ0_1(.din(n8047), .dout(n8044));
    jdff dff_A_4tFhnOGS8_1(.din(n8050), .dout(n8047));
    jdff dff_A_83D1z8j85_1(.din(n8053), .dout(n8050));
    jdff dff_A_qUKP8lz83_1(.din(n8056), .dout(n8053));
    jdff dff_A_DmbFSuqA3_1(.din(n8059), .dout(n8056));
    jdff dff_A_cZg4qVCH0_1(.din(n8062), .dout(n8059));
    jdff dff_A_Bgh0kV3x6_1(.din(n8065), .dout(n8062));
    jdff dff_A_Gs6Q1S7n4_1(.din(n8068), .dout(n8065));
    jdff dff_A_NoSDn8eT1_1(.din(n2133), .dout(n8068));
    jdff dff_A_C14hPYGJ7_2(.din(n8074), .dout(n8071));
    jdff dff_A_z19pZXV52_2(.din(n8077), .dout(n8074));
    jdff dff_A_hAhtHYXq4_2(.din(n8080), .dout(n8077));
    jdff dff_A_un2wKVAb1_2(.din(n8083), .dout(n8080));
    jdff dff_A_ym5MLrHo3_2(.din(n8086), .dout(n8083));
    jdff dff_A_38imtwwk0_2(.din(n8089), .dout(n8086));
    jdff dff_A_sCNAwjks1_2(.din(n8092), .dout(n8089));
    jdff dff_A_yXDZaVji8_2(.din(n8095), .dout(n8092));
    jdff dff_A_gzFbaoh53_2(.din(n8098), .dout(n8095));
    jdff dff_A_8VT3rPAv2_2(.din(n8101), .dout(n8098));
    jdff dff_A_BxA3UUOd6_2(.din(n2133), .dout(n8101));
    jdff dff_B_5JTB6iA73_0(.din(n1986), .dout(n8105));
    jdff dff_B_7Q94a7311_0(.din(n8105), .dout(n8108));
    jdff dff_B_ppoLYKA67_0(.din(n1978), .dout(n8111));
    jdff dff_B_jMsEwQnn4_0(.din(n8111), .dout(n8114));
    jdff dff_B_15lHvnoi4_0(.din(n8114), .dout(n8117));
    jdff dff_A_Z6UpHq8j9_0(.din(n8122), .dout(n8119));
    jdff dff_A_cJa5wY6U9_0(.din(n1975), .dout(n8122));
    jdff dff_A_zxUPhaMp4_1(.din(n8128), .dout(n8125));
    jdff dff_A_kgYENZ1Q6_1(.din(n8131), .dout(n8128));
    jdff dff_A_TXHv3qj30_1(.din(n10034), .dout(n8131));
    jdff dff_A_mqDiXdHA4_2(.din(n8137), .dout(n8134));
    jdff dff_A_bzLkRZRK6_2(.din(n8140), .dout(n8137));
    jdff dff_A_YFww9s9J9_2(.din(n10034), .dout(n8140));
    jdff dff_B_nX47N2lT6_2(.din(n1968), .dout(n8144));
    jdff dff_B_14nPjPx62_2(.din(n8144), .dout(n8147));
    jdff dff_B_DL4bW3ni6_2(.din(n8147), .dout(n8150));
    jdff dff_B_MAKAai9F3_2(.din(n8150), .dout(n8153));
    jdff dff_B_czCQDN6x0_2(.din(n8153), .dout(n8156));
    jdff dff_B_RNkarPww9_2(.din(n8156), .dout(n8159));
    jdff dff_B_habat80T5_2(.din(n8159), .dout(n8162));
    jdff dff_B_KsGKK0G76_2(.din(n8162), .dout(n8165));
    jdff dff_B_ZSSh2JVA7_2(.din(n8165), .dout(n8168));
    jdff dff_B_VDRNsdvG6_2(.din(n8168), .dout(n8171));
    jdff dff_B_AdqVhlJ89_2(.din(n8171), .dout(n8174));
    jdff dff_B_WXIz7OC84_2(.din(n8174), .dout(n8177));
    jdff dff_B_9D8UaAZR2_2(.din(n8177), .dout(n8180));
    jdff dff_A_5O7iKcwa2_1(.din(n4265), .dout(n8182));
    jdff dff_B_ozhs6JXt9_0(.din(n4261), .dout(n8186));
    jdff dff_B_CJNgHhWI8_0(.din(n8186), .dout(n8189));
    jdff dff_B_hsTIU0Cm3_0(.din(n4250), .dout(n8192));
    jdff dff_B_szGITtq51_0(.din(n8192), .dout(n8195));
    jdff dff_B_yb2WQYBS8_0(.din(n8195), .dout(n8198));
    jdff dff_B_J0Qggegj6_0(.din(n8198), .dout(n8201));
    jdff dff_B_kl4sFjwJ4_0(.din(n8201), .dout(n8204));
    jdff dff_B_Vkys7uUa8_0(.din(n4246), .dout(n8207));
    jdff dff_B_rHfN2sbM6_0(.din(n8207), .dout(n8210));
    jdff dff_B_fGBXe76r0_0(.din(n4239), .dout(n8213));
    jdff dff_B_QWgYZoqw4_0(.din(n8213), .dout(n8216));
    jdff dff_B_l531TE5W7_1(.din(n4191), .dout(n8219));
    jdff dff_B_gNhm7Jq30_1(.din(n8219), .dout(n8222));
    jdff dff_B_Vg4DbODl7_1(.din(n4199), .dout(n8225));
    jdff dff_B_txrUvoTl4_1(.din(n4211), .dout(n8228));
    jdff dff_A_aDjpHZsX8_1(.din(n3246), .dout(n8230));
    jdff dff_A_mKI2h6GU8_1(.din(n11104), .dout(n8233));
    jdff dff_A_d7F1LZsA6_2(.din(n11104), .dout(n8236));
    jdff dff_A_WKomwQt33_1(.din(n8242), .dout(n8239));
    jdff dff_A_pTgtjDkw0_1(.din(n8245), .dout(n8242));
    jdff dff_A_Jfle1PDM7_1(.din(n8248), .dout(n8245));
    jdff dff_A_qIt7Kmcb5_1(.din(G77), .dout(n8248));
    jdff dff_A_UUP4SJzO6_2(.din(n8254), .dout(n8251));
    jdff dff_A_mHDmsGcR5_2(.din(n8257), .dout(n8254));
    jdff dff_A_sZ8z3e048_2(.din(n8260), .dout(n8257));
    jdff dff_A_4vBQYFhr8_2(.din(G77), .dout(n8260));
    jdff dff_A_0gSbFn020_1(.din(n10774), .dout(n8263));
    jdff dff_A_KEt89Ekc1_0(.din(n8269), .dout(n8266));
    jdff dff_A_x3Kkhbnz1_0(.din(n8272), .dout(n8269));
    jdff dff_A_ih6rqG6O8_0(.din(n8275), .dout(n8272));
    jdff dff_A_U58CLjyT4_0(.din(n350), .dout(n8275));
    jdff dff_A_2wQ2Iwbd5_2(.din(n8281), .dout(n8278));
    jdff dff_A_h94jdN7j6_2(.din(n8284), .dout(n8281));
    jdff dff_A_bvHmkObR7_2(.din(n350), .dout(n8284));
    jdff dff_A_TtR7O4zu8_1(.din(n10285), .dout(n8287));
    jdff dff_B_tY6y2k0Q3_1(.din(n4131), .dout(n8291));
    jdff dff_B_2SeKlOP91_1(.din(n4139), .dout(n8294));
    jdff dff_B_Qnxe6shB7_1(.din(n4151), .dout(n8297));
    jdff dff_B_0c9EyVMM9_0(.din(n4155), .dout(n8300));
    jdff dff_A_pOidVMvc1_1(.din(n8992), .dout(n8302));
    jdff dff_A_oQWicbQb0_2(.din(n8992), .dout(n8305));
    jdff dff_A_SMHDbw023_0(.din(n8318), .dout(n8308));
    jdff dff_B_PFjQ1lNL0_3(.din(G128), .dout(n8312));
    jdff dff_B_ZdBjMDb04_3(.din(n8312), .dout(n8315));
    jdff dff_B_RnScCPeN8_3(.din(n8315), .dout(n8318));
    jdff dff_B_WXlW6o9w3_1(.din(n4115), .dout(n8321));
    jdff dff_B_fMJ8Nppx0_0(.din(n4123), .dout(n8324));
    jdff dff_A_sSARz3Q60_0(.din(n2148), .dout(n8326));
    jdff dff_A_zBlBIKOh8_1(.din(n8332), .dout(n8329));
    jdff dff_A_ApvMYCUy9_1(.din(n8335), .dout(n8332));
    jdff dff_A_CEa41W7O4_1(.din(n8338), .dout(n8335));
    jdff dff_A_hhva3E7w0_1(.din(n8341), .dout(n8338));
    jdff dff_A_NBZcib8g9_1(.din(n8344), .dout(n8341));
    jdff dff_A_kLq6bmX15_1(.din(n8347), .dout(n8344));
    jdff dff_A_qpAvnoHG2_1(.din(n2148), .dout(n8347));
    jdff dff_A_zVexCDq21_1(.din(n3634), .dout(n8350));
    jdff dff_A_ImVemRGn4_2(.din(n8356), .dout(n8353));
    jdff dff_A_Lohcljm11_2(.din(n2724), .dout(n8356));
    jdff dff_B_lTVgmxFJ7_0(.din(n2720), .dout(n8360));
    jdff dff_B_HkOfbMn44_0(.din(n8360), .dout(n8363));
    jdff dff_B_2kSKJuTH6_0(.din(n2712), .dout(n8366));
    jdff dff_B_0Jc9uF4g1_0(.din(n8366), .dout(n8369));
    jdff dff_A_3xcn83Zx7_0(.din(n2709), .dout(n8371));
    jdff dff_B_YExEAZQO6_0(.din(n3627), .dout(n8375));
    jdff dff_B_u4VORMBn5_0(.din(n8375), .dout(n8378));
    jdff dff_B_qKnH7FET3_0(.din(n8378), .dout(n8381));
    jdff dff_B_B7L1Bb4k5_0(.din(n8381), .dout(n8384));
    jdff dff_B_9Lpsubch3_0(.din(n8384), .dout(n8387));
    jdff dff_A_fzv4lvqZ5_2(.din(n10015), .dout(n8389));
    jdff dff_A_ObJL9Qaa6_1(.din(n8395), .dout(n8392));
    jdff dff_A_Qbg4QAcq7_1(.din(n1791), .dout(n8395));
    jdff dff_A_6kHp5xAf2_2(.din(n8401), .dout(n8398));
    jdff dff_A_tidmV6Lo7_2(.din(n1791), .dout(n8401));
    jdff dff_A_fjKKoOcc0_0(.din(n1904), .dout(n8404));
    jdff dff_A_ZCBBHjxo5_1(.din(n8410), .dout(n8407));
    jdff dff_A_RpbsJLj51_1(.din(n8413), .dout(n8410));
    jdff dff_A_bVqstwWx0_1(.din(n8416), .dout(n8413));
    jdff dff_A_Czkz7sXW1_1(.din(n1485), .dout(n8416));
    jdff dff_B_Z7Hernbb6_1(.din(n1492), .dout(n8420));
    jdff dff_B_ubAYFKGy2_1(.din(n8420), .dout(n8423));
    jdff dff_A_2IVlRPjg5_1(.din(n1473), .dout(n8425));
    jdff dff_B_3aaOt5mu4_1(.din(n1426), .dout(n8429));
    jdff dff_B_aqXTkkMr3_0(.din(n1465), .dout(n8432));
    jdff dff_B_VgwORNHx7_0(.din(n1422), .dout(n8435));
    jdff dff_B_Hn1TlILC1_0(.din(n8435), .dout(n8438));
    jdff dff_B_kXyk0Mo37_1(.din(n1383), .dout(n8441));
    jdff dff_A_0y4SqIvc2_0(.din(n8446), .dout(n8443));
    jdff dff_A_z5vuix598_0(.din(G226), .dout(n8446));
    jdff dff_B_Y6P4RbDG7_1(.din(n1692), .dout(n8450));
    jdff dff_B_tU88pgl64_1(.din(n8450), .dout(n8453));
    jdff dff_A_Mr7Yxxtc5_0(.din(n8458), .dout(n8455));
    jdff dff_A_Kv3wMfzj6_0(.din(n1779), .dout(n8458));
    jdff dff_B_mjwAJ0fu9_0(.din(n1771), .dout(n8462));
    jdff dff_B_pJ9vBfb10_1(.din(n1660), .dout(n8465));
    jdff dff_B_QBUlf6Y68_1(.din(n1703), .dout(n8468));
    jdff dff_B_fFkLKxll7_1(.din(n8468), .dout(n8471));
    jdff dff_B_E3nHGAMP2_1(.din(n8471), .dout(n8474));
    jdff dff_B_d1fElbSb7_0(.din(n1737), .dout(n8477));
    jdff dff_B_Qwl99s273_0(.din(n8477), .dout(n8480));
    jdff dff_B_Do6o7OWl5_1(.din(n1707), .dout(n8483));
    jdff dff_B_qsInAYaB2_1(.din(n8483), .dout(n8486));
    jdff dff_B_YL6HbYWE5_1(.din(n8486), .dout(n8489));
    jdff dff_A_iiFMhJsK0_1(.din(n8494), .dout(n8491));
    jdff dff_A_H2zRB4zY0_1(.din(n1877), .dout(n8494));
    jdff dff_B_ZtZugRSf2_1(.din(n1551), .dout(n8498));
    jdff dff_B_CaBe6qHK8_1(.din(n8498), .dout(n8501));
    jdff dff_A_yHGBWbls2_0(.din(n8506), .dout(n8503));
    jdff dff_A_JChnqbdl4_0(.din(n8509), .dout(n8506));
    jdff dff_A_kl66bIPt4_0(.din(n8512), .dout(n8509));
    jdff dff_A_OF2BZT4e7_0(.din(n1652), .dout(n8512));
    jdff dff_B_GpNB0XTN4_0(.din(n1644), .dout(n8516));
    jdff dff_A_eCFQ9eAD7_1(.din(n8521), .dout(n8518));
    jdff dff_A_khPh2FFN8_1(.din(G226), .dout(n8521));
    jdff dff_A_z5f1lVWD4_2(.din(n8527), .dout(n8524));
    jdff dff_A_6eS5xXQT3_2(.din(n8530), .dout(n8527));
    jdff dff_A_xE7CJdnU0_2(.din(n8533), .dout(n8530));
    jdff dff_A_K5vSNaX49_2(.din(G226), .dout(n8533));
    jdff dff_B_PusZ0kJy6_1(.din(n1519), .dout(n8537));
    jdff dff_B_Nv2GfN377_1(.din(G222), .dout(n8540));
    jdff dff_B_ymDCuxVv0_1(.din(n8540), .dout(n8543));
    jdff dff_A_JFeIDYY74_0(.din(n8549), .dout(n8545));
    jdff dff_B_C0Fl309u4_2(.din(n1449), .dout(n8549));
    jdff dff_A_TiB3qEKA3_1(.din(n8554), .dout(n8551));
    jdff dff_A_UVDxzX8X4_1(.din(n8557), .dout(n8554));
    jdff dff_A_O31Yevz94_1(.din(G77), .dout(n8557));
    jdff dff_B_ZA4Xncnc2_2(.din(G223), .dout(n8561));
    jdff dff_B_3TZf6n5G1_2(.din(n8561), .dout(n8564));
    jdff dff_B_5ysRGQcf9_1(.din(n1562), .dout(n8567));
    jdff dff_B_3Teu5xFQ4_1(.din(n8567), .dout(n8570));
    jdff dff_B_7vdPgLY42_1(.din(n8570), .dout(n8573));
    jdff dff_B_jWr6xEqu8_0(.din(n1610), .dout(n8576));
    jdff dff_B_7SgsIywN8_0(.din(n8576), .dout(n8579));
    jdff dff_A_Nwsjq0xo4_2(.din(n493), .dout(n8581));
    jdff dff_B_oW9LfIcp4_1(.din(n1566), .dout(n8585));
    jdff dff_B_3fcaVetG8_1(.din(n1569), .dout(n8588));
    jdff dff_B_6GLiXLf15_1(.din(n8588), .dout(n8591));
    jdff dff_A_OY2GCQl84_1(.din(n8596), .dout(n8593));
    jdff dff_A_iJX6d4KT1_1(.din(n8599), .dout(n8596));
    jdff dff_A_h1U14QZ20_1(.din(n83), .dout(n8599));
    jdff dff_A_cQXYitet4_2(.din(n8605), .dout(n8602));
    jdff dff_A_nBSbsODQ5_2(.din(n8608), .dout(n8605));
    jdff dff_A_sPbkiv5R3_2(.din(n8611), .dout(n8608));
    jdff dff_A_MwT9xHbC5_2(.din(n83), .dout(n8611));
    jdff dff_A_45ig0oRf4_1(.din(n8617), .dout(n8614));
    jdff dff_A_XNuT9Fvx8_1(.din(n8620), .dout(n8617));
    jdff dff_A_tPqs1ct78_1(.din(n80), .dout(n8620));
    jdff dff_A_JEStj55Q1_2(.din(n8626), .dout(n8623));
    jdff dff_A_efvVhaa88_2(.din(n80), .dout(n8626));
    jdff dff_A_DwRq8D7V4_0(.din(n8632), .dout(n8629));
    jdff dff_A_OzhMKkGv7_0(.din(n77), .dout(n8632));
    jdff dff_A_PVARDvkW4_2(.din(n77), .dout(n8635));
    jdff dff_A_puSTSz594_2(.din(n8641), .dout(n8638));
    jdff dff_A_EL2YGJlr6_2(.din(n8644), .dout(n8641));
    jdff dff_A_y6OI6irt9_2(.din(n77), .dout(n8644));
    jdff dff_A_ayd9RTX27_1(.din(n8650), .dout(n8647));
    jdff dff_A_0UwmGFFC3_1(.din(n8653), .dout(n8650));
    jdff dff_A_dc4sKXuE5_1(.din(G50), .dout(n8653));
    jdff dff_A_pJ3juYXa6_0(.din(n8659), .dout(n8656));
    jdff dff_A_UyoE6NVP6_0(.din(n8665), .dout(n8659));
    jdff dff_A_AEGITx9G9_1(.din(n8665), .dout(n8662));
    jdff dff_A_n01tZAbE4_0(.din(G50), .dout(n8665));
    jdff dff_A_scg5wolC8_2(.din(n8671), .dout(n8668));
    jdff dff_A_8FLMUrlX5_2(.din(n8674), .dout(n8671));
    jdff dff_A_0dGGcx4t0_2(.din(n8677), .dout(n8674));
    jdff dff_A_sQxHYeYf6_2(.din(G50), .dout(n8677));
    jdff dff_A_zwqU6G3F3_0(.din(n8683), .dout(n8680));
    jdff dff_A_ndypIZMF9_0(.din(n2675), .dout(n8683));
    jdff dff_A_Jz517UPj8_0(.din(n8689), .dout(n8686));
    jdff dff_A_cIUoVB911_0(.din(n2672), .dout(n8689));
    jdff dff_B_6Uzw4xNH4_0(.din(n2661), .dout(n8693));
    jdff dff_B_Oz0vXoYE2_0(.din(n8693), .dout(n8696));
    jdff dff_B_SfEUcmPy1_0(.din(n8696), .dout(n8699));
    jdff dff_B_3Tn9GTCJ1_0(.din(n2657), .dout(n8702));
    jdff dff_B_fwNpmsjn6_0(.din(n8702), .dout(n8705));
    jdff dff_B_ddHmRJrI4_0(.din(n8705), .dout(n8708));
    jdff dff_B_QLeR7zmG1_0(.din(n8708), .dout(n8711));
    jdff dff_B_kW1l0wiA6_0(.din(n2650), .dout(n8714));
    jdff dff_B_huqK92bP3_0(.din(n8714), .dout(n8717));
    jdff dff_A_kdtt9xD15_2(.din(n8722), .dout(n8719));
    jdff dff_A_sjnLsLoA7_2(.din(n8725), .dout(n8722));
    jdff dff_A_G4bUzfxV5_2(.din(n8728), .dout(n8725));
    jdff dff_A_SCpKaUiZ8_2(.din(n8731), .dout(n8728));
    jdff dff_A_W39ACTMm9_2(.din(n8734), .dout(n8731));
    jdff dff_A_AtOJHKKB4_2(.din(n8737), .dout(n8734));
    jdff dff_A_VIUQCjfj6_2(.din(n8740), .dout(n8737));
    jdff dff_A_a5wMNEEO6_2(.din(n2121), .dout(n8740));
    jdff dff_A_ZJcudOfX8_0(.din(n8746), .dout(n8743));
    jdff dff_A_OJPfcFCa2_0(.din(n8749), .dout(n8746));
    jdff dff_A_2EEPRluq6_0(.din(n8752), .dout(n8749));
    jdff dff_A_kKrqoSoW7_0(.din(n2118), .dout(n8752));
    jdff dff_B_3h42XZni7_1(.din(n2562), .dout(n8756));
    jdff dff_B_kltxwDtL7_1(.din(n8756), .dout(n8759));
    jdff dff_B_aEOYgQuj1_1(.din(n2585), .dout(n8762));
    jdff dff_B_iyLyyVWW7_1(.din(n2596), .dout(n8765));
    jdff dff_B_ZxTVggiG3_1(.din(n2608), .dout(n8768));
    jdff dff_B_ZNVwHKRe3_0(.din(n2612), .dout(n8771));
    jdff dff_A_dWwjfL9n6_0(.din(n10294), .dout(n8773));
    jdff dff_A_HaSaHwL92_0(.din(n8779), .dout(n8776));
    jdff dff_A_Au7l3aAv2_0(.din(n8782), .dout(n8779));
    jdff dff_A_gbf3SjqU5_0(.din(n11347), .dout(n8782));
    jdff dff_A_oXNKXIQd4_2(.din(n8788), .dout(n8785));
    jdff dff_A_RRAZWhbs1_2(.din(n11347), .dout(n8788));
    jdff dff_A_nByLp5Ye4_0(.din(n8968), .dout(n8791));
    jdff dff_A_vlp8hzqz8_2(.din(n8797), .dout(n8794));
    jdff dff_A_8G95VIjC4_2(.din(n8968), .dout(n8797));
    jdff dff_B_IAYrVm0P9_1(.din(n2566), .dout(n8801));
    jdff dff_B_kbc6CHlm6_0(.din(n2574), .dout(n8804));
    jdff dff_A_Rbqv7i2E2_1(.din(n8816), .dout(n8806));
    jdff dff_B_3Zls9Asu0_3(.din(G311), .dout(n8810));
    jdff dff_B_UKTj6RAy9_3(.din(n8810), .dout(n8813));
    jdff dff_B_mqa966gy6_3(.din(n8813), .dout(n8816));
    jdff dff_B_0Qpqs9IT5_1(.din(n2518), .dout(n8819));
    jdff dff_B_qOHNn4DT0_1(.din(n2526), .dout(n8822));
    jdff dff_B_mA1TS2tU5_1(.din(n2538), .dout(n8825));
    jdff dff_B_2WoV4lU33_1(.din(n2542), .dout(n8828));
    jdff dff_A_gYiziej66_1(.din(n8833), .dout(n8830));
    jdff dff_A_EuaQOspZ3_1(.din(n8836), .dout(n8833));
    jdff dff_A_2pHJVp7l8_1(.din(n11152), .dout(n8836));
    jdff dff_A_jZRrQYj11_2(.din(n8842), .dout(n8839));
    jdff dff_A_9JmFPU7u0_2(.din(n11152), .dout(n8842));
    jdff dff_A_36uqRPDS7_1(.din(n8855), .dout(n8845));
    jdff dff_B_aHADKo1m3_3(.din(G137), .dout(n8849));
    jdff dff_B_BfoOu98b4_3(.din(n8849), .dout(n8852));
    jdff dff_B_a8BNTn3r7_3(.din(n8852), .dout(n8855));
    jdff dff_B_HTpOZOSe8_3(.din(G143), .dout(n8858));
    jdff dff_B_e3iksa357_3(.din(n8858), .dout(n8861));
    jdff dff_B_9juV44ph8_3(.din(n8861), .dout(n8864));
    jdff dff_A_ZKbKDlC72_0(.din(n8888), .dout(n8866));
    jdff dff_A_hvwHxbc04_1(.din(n8872), .dout(n8869));
    jdff dff_A_Jkc8FQ2x6_1(.din(n8888), .dout(n8872));
    jdff dff_A_ML8Wsi7R7_0(.din(n8878), .dout(n8875));
    jdff dff_A_VmKgOIih9_0(.din(n8888), .dout(n8878));
    jdff dff_A_QZZj3G500_1(.din(n8888), .dout(n8881));
    jdff dff_B_qkfBigxd2_3(.din(G159), .dout(n8885));
    jdff dff_B_CuiEmr8G7_3(.din(n8885), .dout(n8888));
    jdff dff_A_SktWqd4B6_1(.din(n8893), .dout(n8890));
    jdff dff_A_ngQMY0wi1_1(.din(n8896), .dout(n8893));
    jdff dff_A_pnXBJf900_1(.din(n8899), .dout(n8896));
    jdff dff_A_HraerFyz3_1(.din(n8902), .dout(n8899));
    jdff dff_A_CAXAfBzv5_1(.din(n10864), .dout(n8902));
    jdff dff_A_qthwE6YC3_2(.din(n8908), .dout(n8905));
    jdff dff_A_sGBZWvyE2_2(.din(n8911), .dout(n8908));
    jdff dff_A_eSlwqHHA1_2(.din(n8914), .dout(n8911));
    jdff dff_A_X6IwQgEE1_2(.din(n8917), .dout(n8914));
    jdff dff_A_pNsegoOF1_2(.din(n10864), .dout(n8917));
    jdff dff_A_rPHqTFGY3_0(.din(n8923), .dout(n8920));
    jdff dff_A_QROsBE3b5_0(.din(n8926), .dout(n8923));
    jdff dff_A_o3YWIpC56_0(.din(G50), .dout(n8926));
    jdff dff_A_Babz9X3p5_2(.din(n8932), .dout(n8929));
    jdff dff_A_Y3f56pMO3_2(.din(n8935), .dout(n8932));
    jdff dff_A_xOecG1PY4_2(.din(n8938), .dout(n8935));
    jdff dff_A_r1HWMIYL7_2(.din(G50), .dout(n8938));
    jdff dff_A_3Dlfw6DB4_1(.din(n8944), .dout(n8941));
    jdff dff_A_8RbOiNs66_1(.din(n8947), .dout(n8944));
    jdff dff_A_ZukS50L22_1(.din(G50), .dout(n8947));
    jdff dff_A_DHGzt0N55_0(.din(n8953), .dout(n8950));
    jdff dff_A_RppjfKcu5_0(.din(n8956), .dout(n8953));
    jdff dff_A_hEyGmNLP2_0(.din(n8959), .dout(n8956));
    jdff dff_A_RACd9pjg9_0(.din(n11452), .dout(n8959));
    jdff dff_A_4PgoHSVp7_1(.din(n8965), .dout(n8962));
    jdff dff_A_oDlAgc7P2_1(.din(n11452), .dout(n8965));
    jdff dff_A_ybsNGNwS9_1(.din(n8971), .dout(n8968));
    jdff dff_A_uXXzrEnG6_1(.din(n8974), .dout(n8971));
    jdff dff_A_JkA8zOvk6_1(.din(n11452), .dout(n8974));
    jdff dff_B_y90EBVFx6_1(.din(n2502), .dout(n8978));
    jdff dff_B_h2dKfwho3_0(.din(n2510), .dout(n8981));
    jdff dff_A_aPGmUDHU2_0(.din(n8986), .dout(n8983));
    jdff dff_A_5v8xR5wt0_0(.din(n8989), .dout(n8986));
    jdff dff_A_wgMpoDW27_0(.din(G150), .dout(n8989));
    jdff dff_A_otD5R4BN9_0(.din(n8995), .dout(n8992));
    jdff dff_A_yX6ndfia3_0(.din(n8998), .dout(n8995));
    jdff dff_A_NQlKKxwd2_0(.din(G150), .dout(n8998));
    jdff dff_A_NkwA5IIM6_1(.din(n9004), .dout(n9001));
    jdff dff_A_8Xx64vZW0_1(.din(n9007), .dout(n9004));
    jdff dff_A_UpKDQn5S3_1(.din(G150), .dout(n9007));
    jdff dff_A_r5Tudtj48_0(.din(n9883), .dout(n9010));
    jdff dff_A_Rn3uLTyX2_1(.din(n9883), .dout(n9013));
    jdff dff_A_O0F2LtgJ8_1(.din(n2159), .dout(n9016));
    jdff dff_A_IlhzGVfX4_1(.din(n9022), .dout(n9019));
    jdff dff_A_WbvVSi4P5_1(.din(n9025), .dout(n9022));
    jdff dff_A_p9A7aHDN9_1(.din(n9028), .dout(n9025));
    jdff dff_A_U7BP3JGa3_1(.din(n9031), .dout(n9028));
    jdff dff_A_qmAdwVV27_1(.din(n9034), .dout(n9031));
    jdff dff_A_mz2Ma50S4_1(.din(n9037), .dout(n9034));
    jdff dff_A_3g9wCvOT0_1(.din(G200), .dout(n9037));
    jdff dff_A_im6BpvSm3_2(.din(n9043), .dout(n9040));
    jdff dff_A_37RYzBOf2_2(.din(n9046), .dout(n9043));
    jdff dff_A_Cd5N8OoT3_2(.din(n9049), .dout(n9046));
    jdff dff_A_ImJQOAUL9_2(.din(n9052), .dout(n9049));
    jdff dff_A_b7z7NBeM2_2(.din(n9055), .dout(n9052));
    jdff dff_A_vZuHoIeq9_2(.din(n9058), .dout(n9055));
    jdff dff_A_UHz0db1u2_2(.din(G200), .dout(n9058));
    jdff dff_A_V3ymdB0E2_0(.din(n2175), .dout(n9061));
    jdff dff_A_Zn9s1wEB5_0(.din(n1360), .dout(n9064));
    jdff dff_A_QvwrTc9j0_1(.din(n9070), .dout(n9067));
    jdff dff_A_ZwLwUUqu8_1(.din(n1360), .dout(n9070));
    jdff dff_A_BmJHWTNA3_1(.din(n9083), .dout(n9073));
    jdff dff_B_koyEFjA78_3(.din(G132), .dout(n9077));
    jdff dff_B_vdjU1Jx73_3(.din(n9077), .dout(n9080));
    jdff dff_B_9BanF2Hg6_3(.din(n9080), .dout(n9083));
    jdff dff_A_jXoD36EM4_0(.din(n9088), .dout(n9085));
    jdff dff_A_MJe5nHEv3_0(.din(n9091), .dout(n9088));
    jdff dff_A_z3nenk1G6_0(.din(n9094), .dout(n9091));
    jdff dff_A_b59GNd0f5_0(.din(n9097), .dout(n9094));
    jdff dff_A_x9e5xlAp3_0(.din(n9100), .dout(n9097));
    jdff dff_A_lTvxQf551_0(.din(n9103), .dout(n9100));
    jdff dff_A_y2vQ4Fxq2_0(.din(n9106), .dout(n9103));
    jdff dff_A_rVInVeyA9_0(.din(n9109), .dout(n9106));
    jdff dff_A_bOjiu0b69_0(.din(n2148), .dout(n9109));
    jdff dff_A_orL5Xhbm1_2(.din(n9115), .dout(n9112));
    jdff dff_A_6LUEUNu30_2(.din(n9118), .dout(n9115));
    jdff dff_A_p8SEAqju9_2(.din(n9121), .dout(n9118));
    jdff dff_A_A7y32vC20_2(.din(n9124), .dout(n9121));
    jdff dff_A_CWC3RigB3_2(.din(n9127), .dout(n9124));
    jdff dff_A_5arkXnx99_2(.din(n9130), .dout(n9127));
    jdff dff_A_Ul0QIhXY5_2(.din(n9133), .dout(n9130));
    jdff dff_A_O9EwWugZ5_2(.din(n9136), .dout(n9133));
    jdff dff_A_dBm7to3B0_2(.din(n2148), .dout(n9136));
    jdff dff_A_T7vBhMUj8_1(.din(n9142), .dout(n9139));
    jdff dff_A_aK57UsaL5_1(.din(n9145), .dout(n9142));
    jdff dff_A_9AWkHB5g3_1(.din(n9148), .dout(n9145));
    jdff dff_A_olxTOttA6_1(.din(n9151), .dout(n9148));
    jdff dff_A_gtx9BhxV3_1(.din(n9154), .dout(n9151));
    jdff dff_A_BwpN446w0_1(.din(n9157), .dout(n9154));
    jdff dff_A_UZVNZD1m5_1(.din(n2148), .dout(n9157));
    jdff dff_A_MfMg31SE1_1(.din(n9163), .dout(n9160));
    jdff dff_A_KVSAQB6x9_1(.din(n9166), .dout(n9163));
    jdff dff_A_wcuik72z9_1(.din(n9169), .dout(n9166));
    jdff dff_A_GWnmYwJh7_1(.din(n9172), .dout(n9169));
    jdff dff_A_lAyJxtep3_1(.din(n9175), .dout(n9172));
    jdff dff_A_pyxeLgzK9_1(.din(n343), .dout(n9175));
    jdff dff_A_REnI5YUr6_2(.din(n9181), .dout(n9178));
    jdff dff_A_wCBDH8kw1_2(.din(n9184), .dout(n9181));
    jdff dff_A_7cPEC6TA0_2(.din(n9187), .dout(n9184));
    jdff dff_A_Q2HUV31o5_2(.din(n9190), .dout(n9187));
    jdff dff_A_yCjTMs0C2_2(.din(n9193), .dout(n9190));
    jdff dff_A_o0x1YyjQ7_2(.din(n343), .dout(n9193));
    jdff dff_A_QFjLQ9A31_0(.din(n9199), .dout(n9196));
    jdff dff_A_Qj78QzEa8_0(.din(n9202), .dout(n9199));
    jdff dff_A_yz5Me03f0_0(.din(n9205), .dout(n9202));
    jdff dff_A_lo2DMc579_0(.din(n9208), .dout(n9205));
    jdff dff_A_pZgIn6Mn2_0(.din(n9211), .dout(n9208));
    jdff dff_A_9lcQDSgC5_0(.din(n9214), .dout(n9211));
    jdff dff_A_Y3zWFNcr3_0(.din(n9217), .dout(n9214));
    jdff dff_A_Q3jL4xQ95_0(.din(n9220), .dout(n9217));
    jdff dff_A_6y2D3p9b0_0(.din(n9223), .dout(n9220));
    jdff dff_A_YLSA4Nci2_0(.din(n9226), .dout(n9223));
    jdff dff_A_qyCW8pT93_0(.din(n9229), .dout(n9226));
    jdff dff_A_1rrweAxJ5_0(.din(n9232), .dout(n9229));
    jdff dff_A_U1nsvXFK9_0(.din(n1430), .dout(n9232));
    jdff dff_A_QlUl0lp24_1(.din(n9238), .dout(n9235));
    jdff dff_A_bir5F7eH1_1(.din(n9241), .dout(n9238));
    jdff dff_A_5sMzEO2c4_1(.din(n9244), .dout(n9241));
    jdff dff_A_EAuUh3eM7_1(.din(n9247), .dout(n9244));
    jdff dff_A_F2iBFrld3_1(.din(n9250), .dout(n9247));
    jdff dff_A_sfCHYGZB6_1(.din(n9253), .dout(n9250));
    jdff dff_A_HgWHZUp25_1(.din(n9256), .dout(n9253));
    jdff dff_A_BbBgQ5tH3_1(.din(n9259), .dout(n9256));
    jdff dff_A_x4Ctfyb41_1(.din(n9262), .dout(n9259));
    jdff dff_A_xW3tbapP7_1(.din(n9265), .dout(n9262));
    jdff dff_A_EoSQQ67C1_1(.din(n9268), .dout(n9265));
    jdff dff_A_frGaIkcL7_1(.din(n9271), .dout(n9268));
    jdff dff_A_01HEKiPv4_1(.din(n1430), .dout(n9271));
    jdff dff_A_apbNwcZG3_1(.din(n9277), .dout(n9274));
    jdff dff_A_bnQIZaMM6_1(.din(n9280), .dout(n9277));
    jdff dff_A_Iu4eF7L16_1(.din(n9283), .dout(n9280));
    jdff dff_A_gFnsGjdN1_1(.din(n9286), .dout(n9283));
    jdff dff_A_q46AWpcw8_1(.din(n9289), .dout(n9286));
    jdff dff_A_MZzf122x5_1(.din(n9292), .dout(n9289));
    jdff dff_A_3CMLQwKD1_1(.din(n9295), .dout(n9292));
    jdff dff_A_VmAgNmDG8_1(.din(n9298), .dout(n9295));
    jdff dff_A_fQNzXRoa0_1(.din(n9301), .dout(n9298));
    jdff dff_A_VYsKwuZb0_1(.din(n9304), .dout(n9301));
    jdff dff_A_xKz9M7fS3_1(.din(n9307), .dout(n9304));
    jdff dff_A_ubaIKEJ61_1(.din(n9310), .dout(n9307));
    jdff dff_A_juqvY5ge5_1(.din(n1430), .dout(n9310));
    jdff dff_A_Ieevp0XE1_2(.din(n9316), .dout(n9313));
    jdff dff_A_mcVKIyD40_2(.din(n9319), .dout(n9316));
    jdff dff_A_CL60yoVR8_2(.din(n9322), .dout(n9319));
    jdff dff_A_5yu8exKE4_2(.din(n9325), .dout(n9322));
    jdff dff_A_Uv0Xm1Bb8_2(.din(n9328), .dout(n9325));
    jdff dff_A_SX3EYtG92_2(.din(n9331), .dout(n9328));
    jdff dff_A_gfvpNFiO8_2(.din(n9334), .dout(n9331));
    jdff dff_A_7Y2f3YIX2_2(.din(n9337), .dout(n9334));
    jdff dff_A_6vzYT7Q89_2(.din(n9340), .dout(n9337));
    jdff dff_A_WXjVGyeo0_2(.din(n9343), .dout(n9340));
    jdff dff_A_icESleKK9_2(.din(n9346), .dout(n9343));
    jdff dff_A_9mB63LIe3_2(.din(n9349), .dout(n9346));
    jdff dff_A_Srm5kXMA6_2(.din(n1430), .dout(n9349));
    jdff dff_A_O64eRFnd9_0(.din(n9355), .dout(n9352));
    jdff dff_A_Zgm7zyNm4_0(.din(n9358), .dout(n9355));
    jdff dff_A_MY5eYnyZ8_0(.din(n9361), .dout(n9358));
    jdff dff_A_jQb7DLmM0_0(.din(n350), .dout(n9361));
    jdff dff_A_wbPRxEi36_1(.din(n9367), .dout(n9364));
    jdff dff_A_BYuIiKA37_1(.din(n350), .dout(n9367));
    jdff dff_B_ToFRmcGQ2_0(.din(n2484), .dout(n9371));
    jdff dff_A_2YbzKGby8_0(.din(n9376), .dout(n9373));
    jdff dff_A_i5Ds5bN29_0(.din(n9403), .dout(n9376));
    jdff dff_A_F0VobcyN5_2(.din(n9382), .dout(n9379));
    jdff dff_A_vjNhp4wO4_2(.din(n9385), .dout(n9382));
    jdff dff_A_f46lkmuH0_2(.din(n9388), .dout(n9385));
    jdff dff_A_LupTeA0c5_2(.din(n9391), .dout(n9388));
    jdff dff_A_BkhVbplY0_2(.din(n9394), .dout(n9391));
    jdff dff_A_ZEPqOYZy9_2(.din(n9397), .dout(n9394));
    jdff dff_A_cf21gQDV6_2(.din(n9400), .dout(n9397));
    jdff dff_A_OSkJvifp7_2(.din(n9403), .dout(n9400));
    jdff dff_A_igeVjMAd9_0(.din(n9406), .dout(n9403));
    jdff dff_A_DHZW8wk15_0(.din(n2118), .dout(n9406));
    jdff dff_A_wM0pIoMX7_2(.din(n9412), .dout(n9409));
    jdff dff_A_9f9VqMzN8_2(.din(n2118), .dout(n9412));
    jdff dff_A_RDucMg3G7_0(.din(n9418), .dout(n9415));
    jdff dff_A_8a8GQP3p1_0(.din(n9421), .dout(n9418));
    jdff dff_A_ZHy6qTz98_0(.din(n9424), .dout(n9421));
    jdff dff_A_eGnqnVtQ8_0(.din(n9427), .dout(n9424));
    jdff dff_A_MU4ralJA4_0(.din(n9430), .dout(n9427));
    jdff dff_A_xPo6llk43_0(.din(n9433), .dout(n9430));
    jdff dff_A_sitLDePJ2_0(.din(n9436), .dout(n9433));
    jdff dff_A_3HYZCYkx5_0(.din(n9439), .dout(n9436));
    jdff dff_A_0a75YB7r5_0(.din(n9442), .dout(n9439));
    jdff dff_A_yVn1imyF0_0(.din(n9445), .dout(n9442));
    jdff dff_A_UeTQRlg70_0(.din(n2114), .dout(n9445));
    jdff dff_A_qUiSdLMH8_0(.din(n9451), .dout(n9448));
    jdff dff_A_fpbiBcSI7_0(.din(n9454), .dout(n9451));
    jdff dff_A_tKvRylP32_0(.din(n9457), .dout(n9454));
    jdff dff_A_QcUlEmmC5_0(.din(n9460), .dout(n9457));
    jdff dff_A_ExKlLBAI1_0(.din(n9463), .dout(n9460));
    jdff dff_A_3ntxPuHO3_0(.din(n9466), .dout(n9463));
    jdff dff_A_8TwwIrNO1_0(.din(n9469), .dout(n9466));
    jdff dff_A_XSZ6sDf47_0(.din(n9472), .dout(n9469));
    jdff dff_A_f96h5L4Q5_0(.din(n9475), .dout(n9472));
    jdff dff_A_hr5bMELX1_0(.din(n9478), .dout(n9475));
    jdff dff_A_9B9zPNJo4_0(.din(n9481), .dout(n9478));
    jdff dff_A_OnG5Egny5_0(.din(n9484), .dout(n9481));
    jdff dff_A_67LEQ4PA8_0(.din(n9487), .dout(n9484));
    jdff dff_A_4RRiHoEs0_0(.din(n2114), .dout(n9487));
    jdff dff_A_hrOe6sHs6_2(.din(n9493), .dout(n9490));
    jdff dff_A_izinCztL5_2(.din(n9496), .dout(n9493));
    jdff dff_A_dh3MLIUd3_2(.din(n9499), .dout(n9496));
    jdff dff_A_mfRb8nQY3_2(.din(n9502), .dout(n9499));
    jdff dff_A_VqJR3Y8P5_2(.din(n9505), .dout(n9502));
    jdff dff_A_NQkrsk995_2(.din(n9508), .dout(n9505));
    jdff dff_A_h2SzWK0d5_2(.din(n9511), .dout(n9508));
    jdff dff_A_7cqMFiTh1_2(.din(n9514), .dout(n9511));
    jdff dff_A_4WHxmVZT4_2(.din(n9517), .dout(n9514));
    jdff dff_A_2RlqY59s8_2(.din(n9520), .dout(n9517));
    jdff dff_A_dzuvx9Vi0_2(.din(n9523), .dout(n9520));
    jdff dff_A_2eAAhsCk3_2(.din(n9526), .dout(n9523));
    jdff dff_A_NMzqwxXi2_2(.din(n2114), .dout(n9526));
    jdff dff_A_2KKKMxEO2_0(.din(n9532), .dout(n9529));
    jdff dff_A_kklXdGwp8_0(.din(n9535), .dout(n9532));
    jdff dff_A_kSUrakpl0_0(.din(n9538), .dout(n9535));
    jdff dff_A_Ze8pyVHu9_0(.din(n9541), .dout(n9538));
    jdff dff_A_Raxmyxn51_0(.din(n9544), .dout(n9541));
    jdff dff_A_uZI1uxxm9_0(.din(n9547), .dout(n9544));
    jdff dff_A_00EfuHWr5_0(.din(n9550), .dout(n9547));
    jdff dff_A_GMZfWSSF1_0(.din(n9553), .dout(n9550));
    jdff dff_A_ZdbF9i3h5_0(.din(n9556), .dout(n9553));
    jdff dff_A_TlThXpMa5_0(.din(n9559), .dout(n9556));
    jdff dff_A_IogcAiqi6_0(.din(n9562), .dout(n9559));
    jdff dff_A_KkVA1EWI4_0(.din(n9565), .dout(n9562));
    jdff dff_A_xqHPYubh0_0(.din(n9568), .dout(n9565));
    jdff dff_A_eZKsSnD04_0(.din(n9571), .dout(n9568));
    jdff dff_A_gETiBfap9_0(.din(n9574), .dout(n9571));
    jdff dff_A_bqP0hXwQ1_0(.din(n9577), .dout(n9574));
    jdff dff_A_hhWxJAtF1_0(.din(n2111), .dout(n9577));
    jdff dff_A_qJzcbsiQ5_0(.din(n9583), .dout(n9580));
    jdff dff_A_fm3xRMa22_0(.din(n9586), .dout(n9583));
    jdff dff_A_Bzdl7SUk7_0(.din(n9589), .dout(n9586));
    jdff dff_A_60nDHZ7A3_0(.din(n9592), .dout(n9589));
    jdff dff_A_r1a9DKN97_0(.din(n9595), .dout(n9592));
    jdff dff_A_twgUN3sy1_0(.din(n9598), .dout(n9595));
    jdff dff_A_EjT8DoTg4_0(.din(n9601), .dout(n9598));
    jdff dff_A_kC8sCidG6_0(.din(n9604), .dout(n9601));
    jdff dff_A_4EBPQli13_0(.din(n9607), .dout(n9604));
    jdff dff_A_w1Dw10HK4_0(.din(n9610), .dout(n9607));
    jdff dff_A_6X0v1u8U8_0(.din(n9613), .dout(n9610));
    jdff dff_A_8j4ASYBC0_0(.din(n9616), .dout(n9613));
    jdff dff_A_KNHB5mhX4_0(.din(n2072), .dout(n9616));
    jdff dff_A_tTRGCba08_2(.din(n9622), .dout(n9619));
    jdff dff_A_9XtKLYwL2_2(.din(n9625), .dout(n9622));
    jdff dff_A_mVGq03yY8_2(.din(n9628), .dout(n9625));
    jdff dff_A_l0g4ARMN5_2(.din(n9631), .dout(n9628));
    jdff dff_A_v63deK9y4_2(.din(n9634), .dout(n9631));
    jdff dff_A_sNeVUY8j4_2(.din(n9637), .dout(n9634));
    jdff dff_A_g4AOfy8l0_2(.din(n9640), .dout(n9637));
    jdff dff_A_vzpxu5bz9_2(.din(n9643), .dout(n9640));
    jdff dff_A_zifp6hnE8_2(.din(n9646), .dout(n9643));
    jdff dff_A_NM5hwlAr7_2(.din(n9649), .dout(n9646));
    jdff dff_A_bKRGQ5hY0_2(.din(n9652), .dout(n9649));
    jdff dff_A_3tXTZQie8_2(.din(n9655), .dout(n9652));
    jdff dff_A_8RFzvmkn8_2(.din(n9658), .dout(n9655));
    jdff dff_A_ImjYv5sH8_2(.din(n9661), .dout(n9658));
    jdff dff_A_vEtMHDQE6_2(.din(n9664), .dout(n9661));
    jdff dff_A_pbO59dpv8_2(.din(n2072), .dout(n9664));
    jdff dff_A_hXaqpHIU1_1(.din(n9670), .dout(n9667));
    jdff dff_A_q6PhK3IL6_1(.din(n9673), .dout(n9670));
    jdff dff_A_5XEw9YYy7_1(.din(n9676), .dout(n9673));
    jdff dff_A_ZuZ08gKE8_1(.din(n9679), .dout(n9676));
    jdff dff_A_QVJ07exF8_1(.din(n9682), .dout(n9679));
    jdff dff_A_0oqXYBeD5_1(.din(n9685), .dout(n9682));
    jdff dff_A_5QKhZG5x9_1(.din(n9688), .dout(n9685));
    jdff dff_A_rbymtoR63_1(.din(n9691), .dout(n9688));
    jdff dff_A_aVB2aesx0_1(.din(n9694), .dout(n9691));
    jdff dff_A_S5mYsdfC6_1(.din(n9697), .dout(n9694));
    jdff dff_A_kzp80mkF1_1(.din(n9700), .dout(n9697));
    jdff dff_A_ekH6s8rA2_1(.din(n9703), .dout(n9700));
    jdff dff_A_7UXBHXrr8_1(.din(n9706), .dout(n9703));
    jdff dff_A_hMqIvqxr9_1(.din(n9709), .dout(n9706));
    jdff dff_A_P99KkVrv0_1(.din(n2069), .dout(n9709));
    jdff dff_A_QdsBB7La3_2(.din(n9715), .dout(n9712));
    jdff dff_A_USn8cusi8_2(.din(n9718), .dout(n9715));
    jdff dff_A_aIuZPe2o1_2(.din(n9721), .dout(n9718));
    jdff dff_A_mH5eGrmt9_2(.din(n9724), .dout(n9721));
    jdff dff_A_319wHlOC7_2(.din(n9727), .dout(n9724));
    jdff dff_A_dz3mmXd33_2(.din(n9730), .dout(n9727));
    jdff dff_A_vDtdNpEu0_2(.din(n9733), .dout(n9730));
    jdff dff_A_msf1W9BA9_2(.din(n9736), .dout(n9733));
    jdff dff_A_gEkg5rZd3_2(.din(n9739), .dout(n9736));
    jdff dff_A_hcecLVZx0_2(.din(n9742), .dout(n9739));
    jdff dff_A_J7f9aLGS7_2(.din(n9745), .dout(n9742));
    jdff dff_A_FFiuvnBX3_2(.din(n9748), .dout(n9745));
    jdff dff_A_OcLCl1li7_2(.din(n9751), .dout(n9748));
    jdff dff_A_wOa8UGtJ2_2(.din(n9754), .dout(n9751));
    jdff dff_A_7Mf11hn86_2(.din(n9757), .dout(n9754));
    jdff dff_A_9oa9JSFi3_2(.din(n2069), .dout(n9757));
    jdff dff_A_o8jC3wy89_0(.din(n248), .dout(n9760));
    jdff dff_B_q5AGVv120_1(.din(n2447), .dout(n9764));
    jdff dff_A_FCrx7MFn5_0(.din(n2469), .dout(n9766));
    jdff dff_A_LzAARKpC1_2(.din(n2469), .dout(n9769));
    jdff dff_A_TBk7QCdd1_1(.din(n2469), .dout(n9772));
    jdff dff_A_Im8C63OO4_1(.din(n9779), .dout(n9775));
    jdff dff_B_cMsoc7sh1_2(.din(n2454), .dout(n9779));
    jdff dff_B_0IyZh3r87_1(.din(n1357), .dout(n9782));
    jdff dff_B_Ja2zN20d8_1(.din(n9782), .dout(n9785));
    jdff dff_A_QPOjnUF42_1(.din(n9790), .dout(n9787));
    jdff dff_A_CiMjb1I22_1(.din(n9793), .dout(n9790));
    jdff dff_A_e41t7c4X0_1(.din(n9796), .dout(n9793));
    jdff dff_A_fRyBsshg1_1(.din(n9799), .dout(n9796));
    jdff dff_A_RGq7ptNu3_1(.din(n9802), .dout(n9799));
    jdff dff_A_rM0bwNhF2_1(.din(n1360), .dout(n9802));
    jdff dff_A_iI3BAws32_2(.din(n1360), .dout(n9805));
    jdff dff_A_NuGbAMwL1_1(.din(n1338), .dout(n9808));
    jdff dff_B_ZH0hIGre5_1(.din(n1318), .dout(n9812));
    jdff dff_B_w8aVsJPu0_1(.din(n9812), .dout(n9815));
    jdff dff_B_7aS6B6hN6_1(.din(n1322), .dout(n9818));
    jdff dff_B_dP8ERMqf7_1(.din(n9818), .dout(n9821));
    jdff dff_B_AFu2vZVl4_0(.din(n1326), .dout(n9824));
    jdff dff_B_7Nb557uG9_0(.din(n9824), .dout(n9827));
    jdff dff_A_FZiDhw6C1_1(.din(n9832), .dout(n9829));
    jdff dff_A_GqESV7yA9_1(.din(n9835), .dout(n9832));
    jdff dff_A_S2bmOonB3_1(.din(n74), .dout(n9835));
    jdff dff_A_vLREaknN6_2(.din(n9841), .dout(n9838));
    jdff dff_A_FKNrCzj53_2(.din(n74), .dout(n9841));
    jdff dff_B_I3nt5hgZ5_0(.din(n1310), .dout(n9845));
    jdff dff_A_xzFq9UPv6_0(.din(n9850), .dout(n9847));
    jdff dff_A_XCiI2xG81_0(.din(n216), .dout(n9850));
    jdff dff_A_i59xcJY51_1(.din(n9856), .dout(n9853));
    jdff dff_A_63v7l7Vq9_1(.din(n216), .dout(n9856));
    jdff dff_A_QWWqCtkg0_0(.din(n9865), .dout(n9859));
    jdff dff_A_Mjh3b7UO7_1(.din(n9865), .dout(n9862));
    jdff dff_A_6m0bHzbb6_0(.din(G58), .dout(n9865));
    jdff dff_A_PrZhEze71_2(.din(n9871), .dout(n9868));
    jdff dff_A_Xg3pnDtJ4_2(.din(n9874), .dout(n9871));
    jdff dff_A_BtUpt0110_2(.din(n9877), .dout(n9874));
    jdff dff_A_pR8uKgO07_2(.din(G58), .dout(n9877));
    jdff dff_A_i85muIC40_1(.din(G58), .dout(n9880));
    jdff dff_A_vHIhuok02_2(.din(n9886), .dout(n9883));
    jdff dff_A_V3pXokVU0_2(.din(n9889), .dout(n9886));
    jdff dff_A_cxfkScNB3_2(.din(G58), .dout(n9889));
    jdff dff_A_Jgno6nkh7_1(.din(G20), .dout(n9892));
    jdff dff_A_igQewKez1_2(.din(n9898), .dout(n9895));
    jdff dff_A_7sF9HlrM6_2(.din(G20), .dout(n9898));
    jdff dff_B_NU60nkyg4_2(.din(n1294), .dout(n9902));
    jdff dff_B_MPLAYylK2_2(.din(n9902), .dout(n9905));
    jdff dff_A_yVgeO5789_0(.din(n9910), .dout(n9907));
    jdff dff_A_F2nHkO901_0(.din(n9913), .dout(n9910));
    jdff dff_A_pZJDfEC69_0(.din(n9916), .dout(n9913));
    jdff dff_A_aVsadp7V2_0(.din(G87), .dout(n9916));
    jdff dff_A_470PHLTQ0_1(.din(n9922), .dout(n9919));
    jdff dff_A_qq2etdfU1_1(.din(n9925), .dout(n9922));
    jdff dff_A_wcSOMHkc7_1(.din(n9928), .dout(n9925));
    jdff dff_A_rGYIVoJs5_1(.din(G87), .dout(n9928));
    jdff dff_A_UY8yXUs39_1(.din(n9934), .dout(n9931));
    jdff dff_A_nhFB6Wdy6_1(.din(n353), .dout(n9934));
    jdff dff_B_v9vq1SUv1_1(.din(n1236), .dout(n9938));
    jdff dff_A_qLHi8o0E6_0(.din(n9943), .dout(n9940));
    jdff dff_A_2sF6EAVe2_0(.din(G232), .dout(n9943));
    jdff dff_A_lwoF2VS19_1(.din(G232), .dout(n9946));
    jdff dff_A_3fRE8kKZ3_1(.din(n9952), .dout(n9949));
    jdff dff_A_PDBLOkoQ0_1(.din(n9955), .dout(n9952));
    jdff dff_A_rwJfIo3F3_1(.din(n9958), .dout(n9955));
    jdff dff_A_CZISefcV8_1(.din(G232), .dout(n9958));
    jdff dff_A_dfXod0py9_2(.din(n9964), .dout(n9961));
    jdff dff_A_wZ3zF3iC5_2(.din(G232), .dout(n9964));
    jdff dff_B_Yea19fe24_0(.din(n1866), .dout(n9968));
    jdff dff_A_lrS1MQPf1_1(.din(n1842), .dout(n9970));
    jdff dff_B_LzLWH8KM7_1(.din(n1815), .dout(n9974));
    jdff dff_A_IHmCwTyd5_1(.din(n1811), .dout(n9976));
    jdff dff_A_Uky4l53N4_0(.din(n1807), .dout(n9979));
    jdff dff_A_AdDCGg8T0_2(.din(n9985), .dout(n9982));
    jdff dff_A_ufRxWv6b1_2(.din(n2057), .dout(n9985));
    jdff dff_B_Ao6zYikO0_0(.din(n2053), .dout(n9989));
    jdff dff_B_2iHUmqcd2_1(.din(n2025), .dout(n9992));
    jdff dff_B_KdKHTE9v4_1(.din(n2029), .dout(n9995));
    jdff dff_A_bXVRJXjo6_1(.din(n10024), .dout(n9997));
    jdff dff_A_lE9FDNoY9_2(.din(n10003), .dout(n10000));
    jdff dff_A_SsxPyY0o6_2(.din(n10006), .dout(n10003));
    jdff dff_A_5zizEvxm1_2(.din(n10009), .dout(n10006));
    jdff dff_A_irrr2R7R5_2(.din(n10012), .dout(n10009));
    jdff dff_A_4iVzRieL8_2(.din(n10024), .dout(n10012));
    jdff dff_A_NINKWWWh6_0(.din(n10018), .dout(n10015));
    jdff dff_A_3ISqDeBM3_0(.din(n10021), .dout(n10018));
    jdff dff_A_P8mMtLYv0_0(.din(n10034), .dout(n10021));
    jdff dff_A_jwSb8tfs3_1(.din(n10027), .dout(n10024));
    jdff dff_A_hMeOEyx59_1(.din(n10034), .dout(n10027));
    jdff dff_B_URPYmcRE4_3(.din(n1927), .dout(n10031));
    jdff dff_B_4euaslRD6_3(.din(n10031), .dout(n10034));
    jdff dff_A_Ym3uFM6E0_0(.din(n1850), .dout(n10036));
    jdff dff_A_t7bUeRsk7_0(.din(n10042), .dout(n10039));
    jdff dff_A_xJcSlXtV9_0(.din(n10045), .dout(n10042));
    jdff dff_A_QZyOovr08_0(.din(n10048), .dout(n10045));
    jdff dff_A_Nai817tk0_0(.din(n10051), .dout(n10048));
    jdff dff_A_Ai49wWVh2_0(.din(n10054), .dout(n10051));
    jdff dff_A_Vbndpgai8_0(.din(n10057), .dout(n10054));
    jdff dff_A_pl2QGNfM2_0(.din(n10060), .dout(n10057));
    jdff dff_A_e30Kr4GF0_0(.din(n10063), .dout(n10060));
    jdff dff_A_dozsGobe8_0(.din(n10066), .dout(n10063));
    jdff dff_A_0JOd5oEu3_0(.din(n10069), .dout(n10066));
    jdff dff_A_L9d9XzyQ5_0(.din(n10072), .dout(n10069));
    jdff dff_A_slHywqOc0_0(.din(G330), .dout(n10072));
    jdff dff_A_FGocdD9N7_0(.din(n10078), .dout(n10075));
    jdff dff_A_A7wXq5rE3_0(.din(n10081), .dout(n10078));
    jdff dff_A_D6sZjnq76_0(.din(n10084), .dout(n10081));
    jdff dff_A_3cS0A53x5_0(.din(n10087), .dout(n10084));
    jdff dff_A_26Dzk5OR2_0(.din(n10090), .dout(n10087));
    jdff dff_A_82IQy6tX3_0(.din(n10093), .dout(n10090));
    jdff dff_A_96QSHZBZ9_0(.din(n10096), .dout(n10093));
    jdff dff_A_XTPuqfGv3_0(.din(n10099), .dout(n10096));
    jdff dff_A_1IoTyaGF1_0(.din(n1924), .dout(n10099));
    jdff dff_A_cuxQ11mA4_1(.din(n10105), .dout(n10102));
    jdff dff_A_fLATu3s21_1(.din(n10108), .dout(n10105));
    jdff dff_A_I1W9SNlC3_1(.din(n10111), .dout(n10108));
    jdff dff_A_LpwxVUGw7_1(.din(n10114), .dout(n10111));
    jdff dff_A_SgKpglzj9_1(.din(n1924), .dout(n10114));
    jdff dff_A_qcuyOwu73_0(.din(n10120), .dout(n10117));
    jdff dff_A_Nzq8A0ba9_0(.din(n10123), .dout(n10120));
    jdff dff_A_oRBHHkxw3_0(.din(n10126), .dout(n10123));
    jdff dff_A_TEJfY3zX3_0(.din(n1924), .dout(n10126));
    jdff dff_A_0yt1rV2I1_2(.din(n10132), .dout(n10129));
    jdff dff_A_sejDLEvb2_2(.din(n10135), .dout(n10132));
    jdff dff_A_jReJ0Rc02_2(.din(n10138), .dout(n10135));
    jdff dff_A_KbtCw2Be9_2(.din(n10141), .dout(n10138));
    jdff dff_A_uDb9li524_2(.din(n10144), .dout(n10141));
    jdff dff_A_sHrhhkQJ2_2(.din(n1924), .dout(n10144));
    jdff dff_A_CL3hdu101_1(.din(n10150), .dout(n10147));
    jdff dff_A_Uzp6K9k27_1(.din(n10153), .dout(n10150));
    jdff dff_A_ghBuExEe4_1(.din(n10156), .dout(n10153));
    jdff dff_A_P1pQTy2S6_1(.din(n10159), .dout(n10156));
    jdff dff_A_GfNU974E0_1(.din(n10162), .dout(n10159));
    jdff dff_A_G0TcI57k1_1(.din(n10165), .dout(n10162));
    jdff dff_A_YGVxfLki0_1(.din(n1920), .dout(n10165));
    jdff dff_A_VlSN2j3M8_2(.din(n10171), .dout(n10168));
    jdff dff_A_T0u8ZC016_2(.din(n10174), .dout(n10171));
    jdff dff_A_qZ6PRYIe3_2(.din(n10177), .dout(n10174));
    jdff dff_A_wYlX2dmG9_2(.din(n10180), .dout(n10177));
    jdff dff_A_KOyNZY7v0_2(.din(n10183), .dout(n10180));
    jdff dff_A_c7UUtwWp8_2(.din(n10186), .dout(n10183));
    jdff dff_A_q1KHmSbO4_2(.din(n1920), .dout(n10186));
    jdff dff_A_nj5ryxbi9_0(.din(G213), .dout(n10189));
    jdff dff_A_06UoBpWW4_2(.din(G213), .dout(n10192));
    jdff dff_A_G2iJTLxm5_0(.din(n10198), .dout(n10195));
    jdff dff_A_CoFQTjdU4_0(.din(n219), .dout(n10198));
    jdff dff_A_0FsblvdM4_1(.din(n10204), .dout(n10201));
    jdff dff_A_awiYCCAm5_1(.din(n10207), .dout(n10204));
    jdff dff_A_DvqUdaea1_1(.din(n10210), .dout(n10207));
    jdff dff_A_IVfs17j22_1(.din(n10213), .dout(n10210));
    jdff dff_A_L7dgG65K4_1(.din(n10216), .dout(n10213));
    jdff dff_A_yESD0x6O4_1(.din(n10219), .dout(n10216));
    jdff dff_A_275NIoSS5_1(.din(n10222), .dout(n10219));
    jdff dff_A_rhmi6y775_1(.din(n10225), .dout(n10222));
    jdff dff_A_Ihnghm883_1(.din(n10228), .dout(n10225));
    jdff dff_A_sjoCCasm5_1(.din(n10231), .dout(n10228));
    jdff dff_A_Q7ura78J7_1(.din(n10234), .dout(n10231));
    jdff dff_A_92H3T4840_1(.din(n10237), .dout(n10234));
    jdff dff_A_uDYQkja50_1(.din(n10240), .dout(n10237));
    jdff dff_A_umE1GkFi4_1(.din(n10243), .dout(n10240));
    jdff dff_A_BFcuhVbu6_1(.din(n219), .dout(n10243));
    jdff dff_A_k97hcDSh2_1(.din(n10249), .dout(n10246));
    jdff dff_A_aunUDTkh1_1(.din(n10252), .dout(n10249));
    jdff dff_A_Su7s7ao33_1(.din(G343), .dout(n10252));
    jdff dff_A_OLc4brm52_1(.din(n1232), .dout(n10255));
    jdff dff_B_nuHoV5pA2_0(.din(n1196), .dout(n10259));
    jdff dff_B_Dh2jux470_1(.din(n1128), .dout(n10262));
    jdff dff_B_0LuljrnG7_1(.din(n1108), .dout(n10265));
    jdff dff_A_c2WzAXFN8_0(.din(n10270), .dout(n10267));
    jdff dff_A_S9HSg5NO7_0(.din(n1093), .dout(n10270));
    jdff dff_A_7Og8lSIe5_0(.din(n10276), .dout(n10273));
    jdff dff_A_Bn0WMGDC3_0(.din(n10279), .dout(n10276));
    jdff dff_A_mMUfU7md6_0(.din(n10282), .dout(n10279));
    jdff dff_A_GsTMAoUY0_0(.din(G294), .dout(n10282));
    jdff dff_A_pnpF4iId6_0(.din(n10288), .dout(n10285));
    jdff dff_A_fjjXIW3l0_0(.din(n10291), .dout(n10288));
    jdff dff_A_IwzbsjN37_0(.din(G294), .dout(n10291));
    jdff dff_A_J5Js87zm5_1(.din(n10297), .dout(n10294));
    jdff dff_A_5N0sKK5d5_1(.din(n10300), .dout(n10297));
    jdff dff_A_KiT15BBB8_1(.din(G294), .dout(n10300));
    jdff dff_A_pH3RywLK4_0(.din(n10903), .dout(n10303));
    jdff dff_A_mgJE9RLR9_1(.din(n10903), .dout(n10306));
    jdff dff_B_xrpfOxV02_0(.din(n1077), .dout(n10310));
    jdff dff_A_i2aqhp5d0_0(.din(n10315), .dout(n10312));
    jdff dff_A_luOPKde94_0(.din(n1074), .dout(n10315));
    jdff dff_B_UDmTyMk91_0(.din(n1070), .dout(n10319));
    jdff dff_A_p2P0Q2Iy0_0(.din(n11068), .dout(n10321));
    jdff dff_A_HoFi2L3R1_1(.din(n11068), .dout(n10324));
    jdff dff_B_MNYOayjY1_0(.din(n1062), .dout(n10328));
    jdff dff_B_WMEaKdvL2_1(.din(n1003), .dout(n10331));
    jdff dff_A_PYEzkkyH2_1(.din(n10336), .dout(n10333));
    jdff dff_A_yvxDBaBU2_1(.din(n10339), .dout(n10336));
    jdff dff_A_SZozDlnA3_1(.din(n10342), .dout(n10339));
    jdff dff_A_5HCXgE3r5_1(.din(n10345), .dout(n10342));
    jdff dff_A_FDG7s6lR2_1(.din(n10348), .dout(n10345));
    jdff dff_A_C3p8AZF36_1(.din(n10351), .dout(n10348));
    jdff dff_A_XHC4JfNo2_1(.din(G190), .dout(n10351));
    jdff dff_A_Jks76VVu9_2(.din(n10357), .dout(n10354));
    jdff dff_A_JpmrROEI9_2(.din(n10360), .dout(n10357));
    jdff dff_A_htK27Vyk1_2(.din(n10363), .dout(n10360));
    jdff dff_A_MFiCQyL13_2(.din(n10366), .dout(n10363));
    jdff dff_A_mdaEY9wk8_2(.din(n10369), .dout(n10366));
    jdff dff_A_FpXd7hDV2_2(.din(n10372), .dout(n10369));
    jdff dff_A_59Z4Cv8n6_2(.din(G190), .dout(n10372));
    jdff dff_B_igReF1fn0_0(.din(n1006), .dout(n10376));
    jdff dff_B_IpaO9w8W7_1(.din(n899), .dout(n10379));
    jdff dff_A_kyk90hop2_1(.din(n987), .dout(n10381));
    jdff dff_B_xzNoOxiA6_1(.din(n975), .dout(n10385));
    jdff dff_A_v5uxyzdr9_0(.din(n10390), .dout(n10387));
    jdff dff_A_HZLZcV8W5_0(.din(n10393), .dout(n10390));
    jdff dff_A_kgIT8jEI1_0(.din(n193), .dout(n10393));
    jdff dff_A_YG7pT8e90_1(.din(n10399), .dout(n10396));
    jdff dff_A_9jxpiqiL7_1(.din(n10402), .dout(n10399));
    jdff dff_A_Q14htJgy1_1(.din(n129), .dout(n10402));
    jdff dff_A_UANVtvih1_2(.din(n129), .dout(n10405));
    jdff dff_A_oSJIeN5g9_1(.din(n418), .dout(n10408));
    jdff dff_A_0HjbQwMa6_2(.din(n418), .dout(n10411));
    jdff dff_A_O5qOvHQS3_1(.din(n952), .dout(n10414));
    jdff dff_A_8bu2HjsL3_1(.din(n940), .dout(n10417));
    jdff dff_A_stTYGT9I3_0(.din(n10423), .dout(n10420));
    jdff dff_A_gFIWSjUS3_0(.din(n933), .dout(n10423));
    jdff dff_A_mo8oFZxj4_1(.din(n10429), .dout(n10426));
    jdff dff_A_jBWtepp39_1(.din(n493), .dout(n10429));
    jdff dff_A_0cZKzsvq7_0(.din(n10444), .dout(n10432));
    jdff dff_A_1Sn75JW53_2(.din(n10444), .dout(n10435));
    jdff dff_A_GzRYhqYM5_0(.din(n10441), .dout(n10438));
    jdff dff_A_3zW65Z0I5_0(.din(n926), .dout(n10441));
    jdff dff_A_uDH37AKn4_0(.din(n190), .dout(n10444));
    jdff dff_A_ubeslu0t4_2(.din(n10450), .dout(n10447));
    jdff dff_A_iFfqgdzM0_2(.din(n10453), .dout(n10450));
    jdff dff_A_BWR7BzNB9_2(.din(n190), .dout(n10453));
    jdff dff_A_KXGCIGqG1_0(.din(n11164), .dout(n10456));
    jdff dff_A_zOSz57x41_1(.din(n10462), .dout(n10459));
    jdff dff_A_JBeus7uJ0_1(.din(n10465), .dout(n10462));
    jdff dff_A_7SAmofy49_1(.din(n10468), .dout(n10465));
    jdff dff_A_13G9R5bH5_1(.din(n11164), .dout(n10468));
    jdff dff_A_BAlsuDBm7_1(.din(n508), .dout(n10471));
    jdff dff_A_jfWcgGkF8_0(.din(n10477), .dout(n10474));
    jdff dff_A_hTVxTAEg9_0(.din(n10480), .dout(n10477));
    jdff dff_A_zgFStbQ32_0(.din(n11203), .dout(n10480));
    jdff dff_A_DyEtyjAH1_1(.din(n10486), .dout(n10483));
    jdff dff_A_Y612Y2Iu4_1(.din(n10489), .dout(n10486));
    jdff dff_A_ccuwuU1G7_1(.din(n11203), .dout(n10489));
    jdff dff_A_fhN7CvxK0_0(.din(n10495), .dout(n10492));
    jdff dff_A_5tAOFhHm9_0(.din(n10498), .dout(n10495));
    jdff dff_A_wltsfTSv8_0(.din(n10501), .dout(n10498));
    jdff dff_A_vbCK6CD48_0(.din(G270), .dout(n10501));
    jdff dff_B_TqeE9gwh0_1(.din(n863), .dout(n10505));
    jdff dff_A_mVRfsAVZ1_1(.din(n10510), .dout(n10507));
    jdff dff_A_1Aer3cB25_1(.din(n867), .dout(n10510));
    jdff dff_A_fsN6Eq2c3_0(.din(n10516), .dout(n10513));
    jdff dff_A_HmsmWUc61_0(.din(n10519), .dout(n10516));
    jdff dff_A_aqNT9f7j3_0(.din(G303), .dout(n10519));
    jdff dff_A_xeeYnU4x7_1(.din(n10525), .dout(n10522));
    jdff dff_A_xhzSbQc21_1(.din(n10528), .dout(n10525));
    jdff dff_A_x85Fx5Bk9_1(.din(n10531), .dout(n10528));
    jdff dff_A_pNIHpZ1O9_1(.din(G303), .dout(n10531));
    jdff dff_A_anOMJ07M0_0(.din(n10537), .dout(n10534));
    jdff dff_A_6Rvvtwnz2_0(.din(n10540), .dout(n10537));
    jdff dff_A_JSgvNSVS9_0(.din(G303), .dout(n10540));
    jdff dff_A_9pmlRJzT8_2(.din(n10546), .dout(n10543));
    jdff dff_A_I7DHatgn6_2(.din(n10549), .dout(n10546));
    jdff dff_A_AWdAOljJ4_2(.din(n10552), .dout(n10549));
    jdff dff_A_bKPcwFxw3_2(.din(G303), .dout(n10552));
    jdff dff_A_x2ult2f57_1(.din(n10558), .dout(n10555));
    jdff dff_A_BcTVejTc8_1(.din(n10561), .dout(n10558));
endmodule

