/*
rf_c880:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 1127
	jand: 153
	jor: 119

Summary:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 1127
	jand: 153
	jor: 119

The maximum logic level gap of any gate:
	rf_c880: 5
*/

module rf_c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n101;
	wire n102;
	wire n103;
	wire n105;
	wire n106;
	wire n107;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n118;
	wire n119;
	wire n121;
	wire n122;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [1:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [1:0] w_G159gat_2;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [1:0] w_G165gat_2;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [1:0] w_G171gat_2;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [1:0] w_G177gat_2;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [1:0] w_G183gat_2;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [2:0] w_G201gat_1;
	wire [2:0] w_G201gat_2;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [1:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [2:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n102_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n111_0;
	wire [2:0] w_n118_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n143_0;
	wire [1:0] w_n149_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n153_1;
	wire [2:0] w_n153_2;
	wire [1:0] w_n153_3;
	wire [1:0] w_n154_0;
	wire [1:0] w_n157_0;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [1:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [2:0] w_n165_0;
	wire [2:0] w_n165_1;
	wire [2:0] w_n167_0;
	wire [1:0] w_n167_1;
	wire [2:0] w_n168_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n181_2;
	wire [1:0] w_n181_3;
	wire [2:0] w_n193_0;
	wire [1:0] w_n193_1;
	wire [2:0] w_n194_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n213_0;
	wire [2:0] w_n217_0;
	wire [1:0] w_n217_1;
	wire [1:0] w_n218_0;
	wire [2:0] w_n222_0;
	wire [1:0] w_n222_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n230_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n236_0;
	wire [1:0] w_n238_0;
	wire [2:0] w_n252_0;
	wire [1:0] w_n255_0;
	wire [2:0] w_n273_0;
	wire [2:0] w_n292_0;
	wire [1:0] w_n292_1;
	wire [2:0] w_n296_0;
	wire [1:0] w_n296_1;
	wire [2:0] w_n299_0;
	wire [1:0] w_n299_1;
	wire [1:0] w_n302_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n305_0;
	wire [1:0] w_n305_1;
	wire [2:0] w_n312_0;
	wire [1:0] w_n312_1;
	wire [1:0] w_n315_0;
	wire [2:0] w_n321_0;
	wire [1:0] w_n321_1;
	wire [1:0] w_n322_0;
	wire [2:0] w_n328_0;
	wire [1:0] w_n328_1;
	wire [2:0] w_n329_0;
	wire [2:0] w_n330_0;
	wire [1:0] w_n331_0;
	wire [2:0] w_n335_0;
	wire [2:0] w_n337_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n340_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n346_1;
	wire [2:0] w_n347_0;
	wire [2:0] w_n367_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n405_0;
	wire w_dff_B_20dLN3zF8_2;
	wire w_dff_B_imBdP2hB7_1;
	wire w_dff_B_bSewn0At8_1;
	wire w_dff_A_HGAmaQlw0_1;
	wire w_dff_B_p1spw8vZ3_0;
	wire w_dff_B_0SVk7vvA0_1;
	wire w_dff_B_grGLpViM1_1;
	wire w_dff_B_Ph8WKAOg1_0;
	wire w_dff_B_rhfo69NT1_1;
	wire w_dff_B_B5B76rGU8_0;
	wire w_dff_B_0Ti6aoJG7_0;
	wire w_dff_B_qHOAPsD99_1;
	wire w_dff_B_gaEppACI8_0;
	wire w_dff_B_QgsYS31O1_2;
	wire w_dff_B_YGClbl2b5_0;
	wire w_dff_B_O4xtUkOQ4_0;
	wire w_dff_B_ybglk5AV2_0;
	wire w_dff_B_AzrEMCtS5_0;
	wire w_dff_B_p8U5SauZ6_0;
	wire w_dff_B_ixm5HORf2_0;
	wire w_dff_B_1Ckw5jTi5_0;
	wire w_dff_B_9ONUZyXy5_0;
	wire w_dff_B_5sfbu1df6_0;
	wire w_dff_B_gsRf9kRE5_0;
	wire w_dff_B_ay7CdLwp0_0;
	wire w_dff_B_lCubPa2y6_0;
	wire w_dff_B_e4tEbFwq7_0;
	wire w_dff_A_uyBtC1KM4_1;
	wire w_dff_A_d02kyb4O8_1;
	wire w_dff_A_zG0SrBk54_1;
	wire w_dff_A_NsjjrEY33_1;
	wire w_dff_A_BU2ztQuX6_1;
	wire w_dff_A_d5I7JrIA4_1;
	wire w_dff_A_y8SpNbTV6_1;
	wire w_dff_A_91NrIlWL9_1;
	wire w_dff_B_gLJK9rfG7_0;
	wire w_dff_B_wqovFkR87_0;
	wire w_dff_B_IFrpMZ5N0_0;
	wire w_dff_B_buhThgss7_0;
	wire w_dff_B_AHzH8W2L4_0;
	wire w_dff_B_T8PDaqa59_0;
	wire w_dff_B_GiovWExW0_0;
	wire w_dff_B_gbJbg8IZ7_0;
	wire w_dff_B_9pbRBZMr3_0;
	wire w_dff_B_5yE5FOPw1_0;
	wire w_dff_B_eny3aYSx1_0;
	wire w_dff_B_TBYpJrwa5_0;
	wire w_dff_B_LlKdc5LR6_0;
	wire w_dff_B_Lq3Kd2KJ5_0;
	wire w_dff_B_Rhy7Vwpy6_0;
	wire w_dff_B_0X2DTZyU9_0;
	wire w_dff_B_2KGvhXHX7_0;
	wire w_dff_B_PkuvAbhw4_0;
	wire w_dff_A_71SzKjgp3_0;
	wire w_dff_A_kMQa9KPt0_0;
	wire w_dff_A_r5yEQohJ0_0;
	wire w_dff_A_kfV1ScLC4_0;
	wire w_dff_B_ARNxSAtR9_1;
	wire w_dff_B_44Lon0vO1_1;
	wire w_dff_B_3aKBqgG15_1;
	wire w_dff_B_OnGJBMIS9_1;
	wire w_dff_A_dqYIZIoN4_1;
	wire w_dff_A_bPr74adn8_1;
	wire w_dff_A_2i2VcIGE8_1;
	wire w_dff_A_zrKGkpZa4_1;
	wire w_dff_A_3j60n8el0_0;
	wire w_dff_A_KjYrMeKG1_0;
	wire w_dff_A_U55PGDX44_0;
	wire w_dff_A_p6xXJuug1_0;
	wire w_dff_A_hHVkuQgB7_0;
	wire w_dff_A_aumyIOC68_0;
	wire w_dff_A_zlP5GoH65_0;
	wire w_dff_A_8UXupTrs7_0;
	wire w_dff_B_jKblZ1Io3_0;
	wire w_dff_B_4Oh6NWAF2_0;
	wire w_dff_B_K1mWKtft0_0;
	wire w_dff_B_AC8deFa16_0;
	wire w_dff_B_Azjf68mi8_0;
	wire w_dff_B_PwwxRCIU4_0;
	wire w_dff_B_PKOBX8gL3_0;
	wire w_dff_B_Z8JMqWBH9_0;
	wire w_dff_B_RGC0gZks6_0;
	wire w_dff_B_2ewSbTsW5_0;
	wire w_dff_B_MniE1BeU3_0;
	wire w_dff_B_MPxPuv9U3_0;
	wire w_dff_B_1B1che8B6_0;
	wire w_dff_B_utPzGWY18_0;
	wire w_dff_B_hM4RozQr3_0;
	wire w_dff_B_UNzA1csy7_0;
	wire w_dff_B_AHbSZy1E6_0;
	wire w_dff_B_jlP1OLvK8_1;
	wire w_dff_B_sCrphbuU2_1;
	wire w_dff_B_LSni4cBE7_1;
	wire w_dff_B_5g2hOEDC3_1;
	wire w_dff_A_GrPBqO918_1;
	wire w_dff_A_bnscJa248_1;
	wire w_dff_A_DxyktazZ8_1;
	wire w_dff_A_9rSqPCBT7_1;
	wire w_dff_B_e5bnfAO46_0;
	wire w_dff_B_bkPu8vnq1_0;
	wire w_dff_B_mXZ9OooB6_0;
	wire w_dff_B_Yf4oWFVd6_0;
	wire w_dff_B_7Nw6Hepr2_0;
	wire w_dff_B_mM67qCh82_0;
	wire w_dff_B_HOwL5CEw0_0;
	wire w_dff_B_ovZcmco80_0;
	wire w_dff_B_UbIOBVj62_0;
	wire w_dff_B_EDmjy9Uf2_0;
	wire w_dff_B_CKNTQsoL2_0;
	wire w_dff_B_BLQanJGl2_0;
	wire w_dff_B_XHEiAOyR0_0;
	wire w_dff_B_8BqY0Q968_0;
	wire w_dff_B_NLR683bv2_0;
	wire w_dff_B_4Uma8bE48_0;
	wire w_dff_B_htQwsgFs6_0;
	wire w_dff_A_HLvrnQlk3_1;
	wire w_dff_A_XRHeV7YM6_1;
	wire w_dff_B_9xZT2iRI4_1;
	wire w_dff_B_pHcCZFPs0_1;
	wire w_dff_B_vRnS05bD7_1;
	wire w_dff_B_nwHzjng78_1;
	wire w_dff_B_Zawc3RUZ2_1;
	wire w_dff_B_taifWXKy4_1;
	wire w_dff_B_aWax5gil0_1;
	wire w_dff_B_ekJRrZl70_1;
	wire w_dff_B_FJtONLbG5_1;
	wire w_dff_B_Vu62d98T6_1;
	wire w_dff_B_x8TNGM6s2_1;
	wire w_dff_B_bmBLbOZ03_1;
	wire w_dff_B_E54BZqYM6_1;
	wire w_dff_B_QG6DV6Jm6_1;
	wire w_dff_B_ZZklmh1s0_1;
	wire w_dff_B_ht8GZpwO0_1;
	wire w_dff_B_91k8CrMr2_1;
	wire w_dff_B_Gu84OHbr3_1;
	wire w_dff_B_bCNiqDY01_1;
	wire w_dff_A_zOBPkLcQ4_0;
	wire w_dff_A_MWDaFW5U3_0;
	wire w_dff_A_EH6Ydh4c5_0;
	wire w_dff_A_W3Rzjnlm1_0;
	wire w_dff_A_YUbiW5946_0;
	wire w_dff_A_QxkZQQRA3_0;
	wire w_dff_A_Gk5jogLs6_0;
	wire w_dff_B_8FQ52lYY8_0;
	wire w_dff_B_IX1kvsFC3_0;
	wire w_dff_B_RcHhDRc17_0;
	wire w_dff_B_l8StTNXe4_0;
	wire w_dff_B_pXwGRbk69_0;
	wire w_dff_B_hZSntnMI9_0;
	wire w_dff_B_WFQYmM1L3_0;
	wire w_dff_B_TaQMXKwf6_0;
	wire w_dff_B_QRwLWZYo2_0;
	wire w_dff_B_vwu3chqa7_0;
	wire w_dff_B_9JYDDdE36_0;
	wire w_dff_B_smpALfaa5_0;
	wire w_dff_B_iJ5QzUeg2_0;
	wire w_dff_B_XSfu6jy41_0;
	wire w_dff_B_iq5ceS9A8_0;
	wire w_dff_B_3I4pFtGl9_0;
	wire w_dff_B_bjeD6pub3_0;
	wire w_dff_B_7KXbOgVN3_0;
	wire w_dff_B_939bfeFA6_0;
	wire w_dff_A_qpejjR656_1;
	wire w_dff_A_ZGrPnzK36_2;
	wire w_dff_A_azNFpMhM8_0;
	wire w_dff_A_e7CKnUIu7_0;
	wire w_dff_A_T9jjpiEI2_0;
	wire w_dff_A_2ubPBvQG8_0;
	wire w_dff_A_dY5lbPeH2_2;
	wire w_dff_A_Y0KSzmJG1_2;
	wire w_dff_B_ocmLXuYB1_0;
	wire w_dff_B_QSNp8d8W0_0;
	wire w_dff_B_x1gLVjkK1_0;
	wire w_dff_B_8nRvfffo3_0;
	wire w_dff_B_UgI77JXC7_0;
	wire w_dff_B_8vVYtivF3_0;
	wire w_dff_B_ZATPpVoE5_0;
	wire w_dff_A_Hf4R2y4P9_1;
	wire w_dff_A_fnZaLzfw6_1;
	wire w_dff_A_iAJ93bts7_1;
	wire w_dff_A_izT8ZUpC3_1;
	wire w_dff_A_wUV9aZlo1_1;
	wire w_dff_A_7x4rsCSo3_1;
	wire w_dff_A_3Y6MdOJP6_1;
	wire w_dff_B_YP1ptw8m1_0;
	wire w_dff_B_qyAHTwhB0_0;
	wire w_dff_B_34uARqsn6_0;
	wire w_dff_B_vQMMS74M7_0;
	wire w_dff_B_6429jJEN6_0;
	wire w_dff_B_oC0b5SRv8_0;
	wire w_dff_B_hZWEU94y7_0;
	wire w_dff_B_AfRRtiyr7_0;
	wire w_dff_B_Fo1aHILk9_0;
	wire w_dff_B_Izf4783V0_0;
	wire w_dff_B_ym3pvic20_0;
	wire w_dff_B_MIHLAari6_0;
	wire w_dff_B_YtlP2FKE4_0;
	wire w_dff_B_Tcu6c5IJ4_0;
	wire w_dff_B_sgHWmJTp7_0;
	wire w_dff_B_jjcIAjEI9_0;
	wire w_dff_B_hgt6o9t34_0;
	wire w_dff_B_MlJi8swA5_0;
	wire w_dff_B_3DYU1nwt0_0;
	wire w_dff_B_utkHbiUL4_0;
	wire w_dff_B_Wh4Yu1TF4_0;
	wire w_dff_B_lQd04rdX2_0;
	wire w_dff_B_T9QDIIpq3_0;
	wire w_dff_B_sBvHmArP9_0;
	wire w_dff_B_1TRPL6zQ8_0;
	wire w_dff_B_2dDd7thp5_0;
	wire w_dff_B_cN5Fl1bl3_0;
	wire w_dff_B_lNQigljw6_0;
	wire w_dff_B_9qONROA47_0;
	wire w_dff_B_PNoVvop11_0;
	wire w_dff_A_GGqPTmaf8_1;
	wire w_dff_A_qJlR1Via2_1;
	wire w_dff_A_1c6f6JN29_1;
	wire w_dff_A_fYQhOLMb1_1;
	wire w_dff_A_PuEJQdU62_1;
	wire w_dff_A_glE6YjOI9_1;
	wire w_dff_A_DD5VzlQI2_1;
	wire w_dff_A_yLKQHjhw5_1;
	wire w_dff_A_zguWoSTU8_1;
	wire w_dff_B_Njars19K6_1;
	wire w_dff_B_T1w9DNB23_1;
	wire w_dff_B_nBOiScYI3_1;
	wire w_dff_A_3NFqrWk85_1;
	wire w_dff_A_XJ75fKMM1_1;
	wire w_dff_A_4sauANMr5_1;
	wire w_dff_A_5Rc1NTn82_1;
	wire w_dff_A_22EzaNRH2_1;
	wire w_dff_A_YFVx8Hve1_1;
	wire w_dff_A_3CXBDjGy9_1;
	wire w_dff_A_ONychntC1_2;
	wire w_dff_A_4GwYeHZU7_2;
	wire w_dff_A_rZWI63BR4_2;
	wire w_dff_A_rCHswxiA2_2;
	wire w_dff_A_4CYVFgmW9_2;
	wire w_dff_A_1b3pr0Eu8_2;
	wire w_dff_A_pFZYmTHO8_2;
	wire w_dff_A_7j1cYmm35_2;
	wire w_dff_A_7QNwRjLL8_2;
	wire w_dff_A_VALLlZDi7_2;
	wire w_dff_A_Y7MJgL9w2_2;
	wire w_dff_B_fI6OMezF4_0;
	wire w_dff_B_PUoCACqF5_0;
	wire w_dff_B_FCcmQtCQ5_0;
	wire w_dff_B_WjlhjVFz8_0;
	wire w_dff_A_L73bfKqD5_1;
	wire w_dff_A_QRSBxjvm0_1;
	wire w_dff_A_smHjJcy14_1;
	wire w_dff_A_AbClJDsC1_1;
	wire w_dff_B_JLFDRsbE1_1;
	wire w_dff_B_TI3tV9FD4_1;
	wire w_dff_B_6W5xi0fm4_1;
	wire w_dff_B_mLJ7Ql8H6_0;
	wire w_dff_B_7URkGVGW8_0;
	wire w_dff_B_EPuOvwon3_0;
	wire w_dff_B_LpuWcMhc0_0;
	wire w_dff_A_d5WapaAd8_1;
	wire w_dff_A_j39aCgnn3_1;
	wire w_dff_A_Aga2VbG81_1;
	wire w_dff_A_W22bFRvE6_1;
	wire w_dff_B_OJKZr1Pa1_1;
	wire w_dff_B_VE2PbU0n4_1;
	wire w_dff_B_PdEw4Pai8_1;
	wire w_dff_B_YbtlO2aU0_1;
	wire w_dff_B_U9yoAtHN1_1;
	wire w_dff_B_UsVqLjAM8_1;
	wire w_dff_B_pRJznE1q4_1;
	wire w_dff_B_CO0TEYyV5_0;
	wire w_dff_B_RfywZe636_0;
	wire w_dff_B_7q6IeY6F4_0;
	wire w_dff_B_R2TlDJIS9_0;
	wire w_dff_B_V8mtbQ7e9_0;
	wire w_dff_B_KiN71b3D9_0;
	wire w_dff_B_Feks7tyM3_0;
	wire w_dff_B_pD7DtAH65_0;
	wire w_dff_B_PxDM8Pdk2_0;
	wire w_dff_B_knFNQfaJ1_0;
	wire w_dff_B_TkBwFMYm3_0;
	wire w_dff_B_2spQn6sk2_0;
	wire w_dff_B_mKHVLYLl6_0;
	wire w_dff_B_r4tmjpNV0_0;
	wire w_dff_B_MBICdgy26_0;
	wire w_dff_B_qyXVzmYJ7_0;
	wire w_dff_A_hA9yRRx98_1;
	wire w_dff_A_EKF1ZGSF3_1;
	wire w_dff_A_hBLY9SOv4_1;
	wire w_dff_A_pBohs5H37_1;
	wire w_dff_A_6LWhfFPr7_1;
	wire w_dff_B_cB1AxH6V7_0;
	wire w_dff_B_KKaxXAic3_0;
	wire w_dff_B_CH4j4C5Y7_0;
	wire w_dff_B_ZAcBpBG22_0;
	wire w_dff_B_GJ3Zrlbj5_0;
	wire w_dff_B_t4CSkoIp3_1;
	wire w_dff_B_ow44jL611_1;
	wire w_dff_B_N35O9IcH8_1;
	wire w_dff_B_U8Jo871b9_1;
	wire w_dff_B_efg2qdYU1_1;
	wire w_dff_B_emH93ejM9_1;
	wire w_dff_B_mrW5kCZ85_1;
	wire w_dff_B_HQAup70o0_1;
	wire w_dff_B_OelSTeiU1_1;
	wire w_dff_B_mZuN47YQ3_1;
	wire w_dff_B_Jr5ZHMyQ0_1;
	wire w_dff_B_kn2ms3Rz5_1;
	wire w_dff_B_q4xEbWFW2_1;
	wire w_dff_B_QNGxCLSY9_1;
	wire w_dff_B_fkPCQbba7_1;
	wire w_dff_B_AlOKLYwV3_0;
	wire w_dff_B_FvY63EkL9_0;
	wire w_dff_B_fNYjGCB03_0;
	wire w_dff_B_f84puu9g0_0;
	wire w_dff_B_4z0SVa6o3_0;
	wire w_dff_B_3XQtlWSc7_0;
	wire w_dff_A_D5s9Hsp36_0;
	wire w_dff_A_3VFNgtBl1_0;
	wire w_dff_A_eiCg0iHe0_0;
	wire w_dff_A_YwyFruk58_0;
	wire w_dff_A_J8mq48JQ0_0;
	wire w_dff_A_dfDj8RWL9_0;
	wire w_dff_A_KbcVS7sh7_2;
	wire w_dff_A_KnGvYnNg0_0;
	wire w_dff_A_rIpQowp34_0;
	wire w_dff_A_qJKfoSUw4_0;
	wire w_dff_A_bPA3mF5m3_0;
	wire w_dff_A_90RkIKWw4_0;
	wire w_dff_A_wS7nXe1t7_0;
	wire w_dff_B_lkdbdiPE2_1;
	wire w_dff_A_Ko2xzVei3_0;
	wire w_dff_A_wuiXzE2p2_0;
	wire w_dff_A_5xkH4MHd4_0;
	wire w_dff_A_oLAu9PgN6_0;
	wire w_dff_A_DmMZkXHQ6_0;
	wire w_dff_A_UoymzHYZ3_0;
	wire w_dff_A_KPkjkTHf0_0;
	wire w_dff_A_iKnk4anM6_1;
	wire w_dff_A_ddbxkrov7_1;
	wire w_dff_A_Y1Bdosnl9_1;
	wire w_dff_A_diCDEsHX2_1;
	wire w_dff_A_RVw0n8sK9_1;
	wire w_dff_A_pndzv8ct0_1;
	wire w_dff_A_yMQ6iL6S3_1;
	wire w_dff_A_alIZJUzz0_1;
	wire w_dff_A_UJ7N9NOf9_1;
	wire w_dff_B_5CABIsTw2_0;
	wire w_dff_B_TjBTKXoi7_0;
	wire w_dff_B_i5cAmkLc7_0;
	wire w_dff_A_jvc0pF3Z5_1;
	wire w_dff_A_eJxtZOeL6_1;
	wire w_dff_A_j6aI7Icb3_1;
	wire w_dff_A_lTYqFZCO3_1;
	wire w_dff_A_TJCZ1xdI6_1;
	wire w_dff_A_WnLAxBC29_1;
	wire w_dff_A_jc7HTzSh1_1;
	wire w_dff_A_bsCysOS74_2;
	wire w_dff_A_vFormJ3P0_2;
	wire w_dff_A_jxuKexFD5_2;
	wire w_dff_A_pIJI1wR47_2;
	wire w_dff_A_sbFtc1u37_2;
	wire w_dff_A_VaX0XcJM4_2;
	wire w_dff_A_5KNPP9EU7_2;
	wire w_dff_A_eterAJUo3_2;
	wire w_dff_A_RYypYTir9_2;
	wire w_dff_A_7LdjYk5T4_2;
	wire w_dff_A_8XpGyw5C6_2;
	wire w_dff_B_zeyF7S7C6_0;
	wire w_dff_B_i6oBulh41_0;
	wire w_dff_B_EgtbQ1og3_0;
	wire w_dff_B_uGwKqtyq4_0;
	wire w_dff_B_ssY13juN7_0;
	wire w_dff_B_3ZBUr4P26_0;
	wire w_dff_B_pMpnmSFT7_0;
	wire w_dff_B_qMGeSdpT8_0;
	wire w_dff_B_xXJGaZgs1_0;
	wire w_dff_B_bBEt4ZWG5_0;
	wire w_dff_B_cYhKNdA75_0;
	wire w_dff_B_nBQKbeDD7_0;
	wire w_dff_B_LovpfXDU5_0;
	wire w_dff_B_ANnB8LUY2_0;
	wire w_dff_B_z0Aue9fS2_0;
	wire w_dff_B_Pv1yspMa9_0;
	wire w_dff_A_it6uYGN15_1;
	wire w_dff_A_N6o8wclS5_1;
	wire w_dff_A_F2bI8AQq9_1;
	wire w_dff_A_iKwxcC1S7_1;
	wire w_dff_A_98YQrYo79_1;
	wire w_dff_B_vTI34gNP8_1;
	wire w_dff_A_LxxNHobh5_0;
	wire w_dff_A_shD5mLGa3_0;
	wire w_dff_B_CrHvogc18_0;
	wire w_dff_B_k7j50dZ35_0;
	wire w_dff_B_lzpiCVSF1_0;
	wire w_dff_B_RckJwQxV6_0;
	wire w_dff_B_Gm0kNzhg3_0;
	wire w_dff_B_0gjBhWBg7_3;
	wire w_dff_A_JhAco3gd1_2;
	wire w_dff_B_yH1b8k1E3_3;
	wire w_dff_B_ZB59Gv4L7_3;
	wire w_dff_B_7sgX5yrC5_3;
	wire w_dff_B_OdRa28TU4_3;
	wire w_dff_B_Wy3Gey7V3_3;
	wire w_dff_B_T8GuwOpR6_3;
	wire w_dff_B_MSA3xcpb2_3;
	wire w_dff_B_cunaExpD1_3;
	wire w_dff_A_FWaJm0wq7_0;
	wire w_dff_A_s3hp9UnE5_0;
	wire w_dff_A_RcxMbyay4_0;
	wire w_dff_A_XopyLnzA5_0;
	wire w_dff_A_yvWTABtl4_0;
	wire w_dff_A_ViQqoSan2_0;
	wire w_dff_A_dL1MpdZe6_0;
	wire w_dff_A_2WeA3owF7_0;
	wire w_dff_A_WIADCNa01_1;
	wire w_dff_A_j2mV2HVv6_1;
	wire w_dff_B_LECh1TG46_3;
	wire w_dff_B_k2ACAfl64_3;
	wire w_dff_B_QAiyhTQn6_3;
	wire w_dff_B_hTK7h19Q7_3;
	wire w_dff_B_Wrja4ard4_3;
	wire w_dff_B_Zb8Mnr6N1_3;
	wire w_dff_B_JABA05kb4_3;
	wire w_dff_B_js1SSsc40_3;
	wire w_dff_B_iTMyeUSy8_3;
	wire w_dff_B_ZL8ZAyZh2_3;
	wire w_dff_B_NiV2AKPp7_1;
	wire w_dff_B_90CIGYAP8_1;
	wire w_dff_B_O7GIOyoc4_1;
	wire w_dff_B_MQ5HIeHj0_1;
	wire w_dff_B_ligpKIir9_1;
	wire w_dff_B_zy5x0kiP4_1;
	wire w_dff_B_VpozsdDg7_1;
	wire w_dff_B_2esykH8h4_1;
	wire w_dff_B_NLszNRtg2_1;
	wire w_dff_B_lYounoyC7_1;
	wire w_dff_B_fRQc0Ubi5_1;
	wire w_dff_B_PWsRhbmR1_1;
	wire w_dff_B_HVkZ9dnD0_1;
	wire w_dff_B_kHP8xzmV3_1;
	wire w_dff_B_0q7Y0Ifp9_1;
	wire w_dff_B_dvgKbKCL6_1;
	wire w_dff_B_QyXeecTJ0_1;
	wire w_dff_B_VLbt0aoS7_0;
	wire w_dff_B_tkk7Pp4Y7_0;
	wire w_dff_B_Fw2zGQ9u2_0;
	wire w_dff_B_u8LhLyL08_0;
	wire w_dff_B_3dK4KEEy6_0;
	wire w_dff_B_gorGpyFJ5_0;
	wire w_dff_B_L0320AkD2_0;
	wire w_dff_A_0lyqxPsZ5_0;
	wire w_dff_A_WzPbRMYu6_0;
	wire w_dff_A_tlvt9k2R0_0;
	wire w_dff_A_s3zgy9cj0_0;
	wire w_dff_A_OCJEHcr90_0;
	wire w_dff_A_burd5mjC4_0;
	wire w_dff_A_kScFJcsb4_0;
	wire w_dff_A_WK3aLGhH9_0;
	wire w_dff_A_jw1L4KQf4_0;
	wire w_dff_A_gF8O0kOx7_0;
	wire w_dff_A_h3AlJXLC9_0;
	wire w_dff_A_pX56OMCk2_0;
	wire w_dff_A_ZXyQHwlc3_0;
	wire w_dff_A_kPNf8Wh39_0;
	wire w_dff_B_M8u8lpIW6_1;
	wire w_dff_B_dfzaaTg61_1;
	wire w_dff_B_5JtSqqhk2_1;
	wire w_dff_B_XEQnazf80_1;
	wire w_dff_B_FxFBpVrk9_1;
	wire w_dff_B_wJ5ruUjE4_1;
	wire w_dff_B_NzKj01Qv2_1;
	wire w_dff_B_maYxTiIJ7_1;
	wire w_dff_B_BU8RXXAE6_1;
	wire w_dff_B_zCTWHUUc0_0;
	wire w_dff_A_U8VkxY2G1_0;
	wire w_dff_B_HJhhk2Za1_1;
	wire w_dff_A_yAdCop6Z3_0;
	wire w_dff_A_xMfnZn0I7_0;
	wire w_dff_A_C4oHFx8z8_0;
	wire w_dff_A_0UYYGZAd7_1;
	wire w_dff_A_dKYJ5aZf9_1;
	wire w_dff_A_aZn7jFaW6_1;
	wire w_dff_A_9LjsbrFf8_1;
	wire w_dff_A_pF2s8jJy7_1;
	wire w_dff_A_VB2fzTlZ8_1;
	wire w_dff_A_h6fWmWR07_1;
	wire w_dff_A_DTUD1R403_1;
	wire w_dff_A_JHMj1Keu4_2;
	wire w_dff_A_NaguskDQ5_2;
	wire w_dff_A_aZxjJvh80_2;
	wire w_dff_A_BjECwNAx5_2;
	wire w_dff_A_RqT43T9y2_2;
	wire w_dff_A_rCeAFLiN1_2;
	wire w_dff_A_Qv1SyCfy9_2;
	wire w_dff_A_fsxYyJjG3_2;
	wire w_dff_A_t2VKqC012_1;
	wire w_dff_A_rKur3qzb4_1;
	wire w_dff_A_6FlEJPGT6_1;
	wire w_dff_A_8s9P6lSF8_1;
	wire w_dff_A_ED5y1Mrd2_1;
	wire w_dff_A_rG8SlCZZ8_1;
	wire w_dff_A_jN2amZtz9_1;
	wire w_dff_A_Bk71gHeV9_1;
	wire w_dff_A_Ml3LPoRN6_2;
	wire w_dff_A_Cb2IXG5A8_2;
	wire w_dff_A_W7xMu0jm8_2;
	wire w_dff_A_U46mvkgj9_2;
	wire w_dff_A_KSUlxIVK5_2;
	wire w_dff_A_XkLLA4j06_2;
	wire w_dff_A_hMy2MXLM0_2;
	wire w_dff_A_ihUrwOyU2_2;
	wire w_dff_B_7A8CQ8wf1_0;
	wire w_dff_A_c2yYKDc01_0;
	wire w_dff_A_WkSOeeeh6_0;
	wire w_dff_A_EEBKWNz20_0;
	wire w_dff_B_rRvGpYtZ9_1;
	wire w_dff_A_v5nfyNWc3_0;
	wire w_dff_A_Eq6Muw3W5_0;
	wire w_dff_A_VQx0RyiS8_0;
	wire w_dff_A_OKECXWQi5_0;
	wire w_dff_A_fyBPgIOs4_0;
	wire w_dff_A_7WBawzON4_0;
	wire w_dff_A_QmSLiku04_0;
	wire w_dff_A_xFXitK0D6_0;
	wire w_dff_A_ksId0XEv9_0;
	wire w_dff_A_3C6fbs1i9_0;
	wire w_dff_A_FMfH9g317_0;
	wire w_dff_A_9XhzZTb43_0;
	wire w_dff_A_IpqDrjdh0_0;
	wire w_dff_A_HZkf69Kn8_2;
	wire w_dff_A_jrjUOp1I0_2;
	wire w_dff_A_vn9IGqtz7_2;
	wire w_dff_A_7tnFYHLD3_2;
	wire w_dff_B_HP1pRa9y2_1;
	wire w_dff_A_K4JB3bi80_1;
	wire w_dff_A_rLOPMm421_1;
	wire w_dff_A_O2Gy59Yd5_1;
	wire w_dff_A_eNwx5A8U0_1;
	wire w_dff_A_4J4xqKLW5_1;
	wire w_dff_A_kvfY68hY2_1;
	wire w_dff_B_g8xrYXn64_2;
	wire w_dff_B_ZDNC6rPy5_2;
	wire w_dff_B_LrlYXd8T1_2;
	wire w_dff_B_piD0i7Xt2_2;
	wire w_dff_A_avSQB05u4_0;
	wire w_dff_A_ohMpxTvy5_0;
	wire w_dff_A_18xIItvs4_0;
	wire w_dff_A_ZJEF9ZSQ7_0;
	wire w_dff_A_uLTmUqcE9_0;
	wire w_dff_A_gAhvSEBA2_0;
	wire w_dff_A_5MuUyKNx9_0;
	wire w_dff_A_PNmlGw7p8_0;
	wire w_dff_A_WKhiULLH2_2;
	wire w_dff_A_3evzTTmu8_2;
	wire w_dff_A_oqqOtPtr9_2;
	wire w_dff_A_7awGszEe9_2;
	wire w_dff_B_Bj9Xhqiq0_1;
	wire w_dff_B_YWJF9daW1_1;
	wire w_dff_B_0aZHIupd6_1;
	wire w_dff_B_zp8Q2MNX9_1;
	wire w_dff_B_Scid7VSd1_1;
	wire w_dff_B_6QO0Oz3U5_1;
	wire w_dff_B_kboDXVne9_1;
	wire w_dff_B_l3EjJiUZ8_1;
	wire w_dff_B_skd7gkZr8_1;
	wire w_dff_B_CRE4zai05_1;
	wire w_dff_B_aaNCrRes6_0;
	wire w_dff_B_teIs8hoA6_0;
	wire w_dff_B_F6Wksyvu4_1;
	wire w_dff_B_Ji6T9NuC1_1;
	wire w_dff_B_1maUqPPy8_1;
	wire w_dff_B_aGrgTfJx5_1;
	wire w_dff_B_308swCCT8_1;
	wire w_dff_B_WHqEB5UA4_1;
	wire w_dff_B_RgedzBox4_1;
	wire w_dff_B_zcWU9T686_1;
	wire w_dff_B_CEyhQme00_1;
	wire w_dff_B_OT2NGZCo5_2;
	wire w_dff_B_o62SLLAi8_2;
	wire w_dff_B_weoeNh1Z2_2;
	wire w_dff_B_QLqm9Rjl5_2;
	wire w_dff_B_fqdGfhSa0_2;
	wire w_dff_B_jlAjge222_2;
	wire w_dff_B_PNREf1H55_2;
	wire w_dff_B_O7IYYnW93_2;
	wire w_dff_B_W8buxaVQ2_2;
	wire w_dff_A_eI1hEaNQ3_0;
	wire w_dff_A_eEZuc3JX5_0;
	wire w_dff_A_gzGnGGAu2_0;
	wire w_dff_A_BXzaIjEq7_0;
	wire w_dff_A_6N9GaMhU6_0;
	wire w_dff_A_PqkO6H438_0;
	wire w_dff_A_MDCxWnEX0_0;
	wire w_dff_A_SkK6WUdn5_0;
	wire w_dff_A_EPD7r3wi6_0;
	wire w_dff_A_Zx2Dsoyo2_1;
	wire w_dff_A_xVZx3eOO5_1;
	wire w_dff_A_yy4Xcum80_1;
	wire w_dff_A_IKIePTK22_1;
	wire w_dff_A_xCoL9wn42_1;
	wire w_dff_A_ArIkvXv60_1;
	wire w_dff_A_xODEzUgS7_1;
	wire w_dff_A_gQitHaxw7_1;
	wire w_dff_A_fwjkoGRV6_1;
	wire w_dff_A_bSvZyBQD0_0;
	wire w_dff_A_WmCX4QAd4_1;
	wire w_dff_A_Ozb6AsFn9_0;
	wire w_dff_A_BZzvcps99_0;
	wire w_dff_A_NmSiOZAZ2_0;
	wire w_dff_A_9Q1Z28lf8_0;
	wire w_dff_A_WeingIaf9_0;
	wire w_dff_A_GWKmMSds5_1;
	wire w_dff_A_MZNSBQMW6_1;
	wire w_dff_A_dHCIQLS56_1;
	wire w_dff_A_CqfVyh1X8_1;
	wire w_dff_A_ZoFaf9jF1_1;
	wire w_dff_A_faiL1H6P0_1;
	wire w_dff_A_nbBr9Jmr4_1;
	wire w_dff_A_KCKcfahM1_1;
	wire w_dff_A_fqYz0gn91_2;
	wire w_dff_A_KkK22m7r8_2;
	wire w_dff_A_WyfH7fgS7_2;
	wire w_dff_A_bt1n3pah3_2;
	wire w_dff_A_nNciEC3p7_2;
	wire w_dff_A_Q4679qAd0_2;
	wire w_dff_A_f9bvKH217_2;
	wire w_dff_A_I0eyeOdC1_2;
	wire w_dff_A_V0DLYVtI8_2;
	wire w_dff_A_AWcbRMiQ4_2;
	wire w_dff_A_zpr6cEBJ4_2;
	wire w_dff_A_QZg04gcl8_2;
	wire w_dff_A_7PhRkVid1_1;
	wire w_dff_A_dr9yFtro2_1;
	wire w_dff_A_eXq9rgTs1_1;
	wire w_dff_A_yqcEP5M88_1;
	wire w_dff_A_d6UTlw6b8_1;
	wire w_dff_A_t1XsacIZ5_1;
	wire w_dff_A_VUDk8WcB1_1;
	wire w_dff_A_gKAnkFhG8_1;
	wire w_dff_A_YWGPJBXF6_1;
	wire w_dff_B_DGX4PC4T2_1;
	wire w_dff_A_HVyJZuJi9_1;
	wire w_dff_A_iAL4fUL74_1;
	wire w_dff_A_VWf8y2e67_1;
	wire w_dff_A_7RlY8bLN9_1;
	wire w_dff_A_uIjmtxar9_1;
	wire w_dff_A_tfwqjyyU3_1;
	wire w_dff_A_EftGHX5V2_1;
	wire w_dff_A_8oI9TO9J2_2;
	wire w_dff_A_vUIuLwci3_2;
	wire w_dff_A_ddvr60bq8_1;
	wire w_dff_A_rKyPGpVz7_1;
	wire w_dff_A_QlSQTq4C2_2;
	wire w_dff_A_w9FWJmsQ3_2;
	wire w_dff_B_8kWAgWBF9_0;
	wire w_dff_A_wI6DRQ022_0;
	wire w_dff_A_jds7d27L4_0;
	wire w_dff_A_Wzfu0KCD4_0;
	wire w_dff_A_XR9CSE6t7_1;
	wire w_dff_B_XOaP6XDE5_2;
	wire w_dff_B_ttmPs0EQ7_2;
	wire w_dff_B_zp4lH0lP0_2;
	wire w_dff_B_SKyVliyN8_2;
	wire w_dff_A_1W0H5qBI4_0;
	wire w_dff_A_wSAYqYIq6_0;
	wire w_dff_A_KTxNf5Mh6_0;
	wire w_dff_A_PomoBPfT4_0;
	wire w_dff_A_jMBcLWEX5_0;
	wire w_dff_A_ClVOk8HB2_0;
	wire w_dff_A_UztsRuXl7_0;
	wire w_dff_A_vSNtDbIa9_0;
	wire w_dff_A_jXmvuQg96_1;
	wire w_dff_A_pWHCK0eD6_1;
	wire w_dff_A_RE7WW2799_1;
	wire w_dff_A_M3JOp4nt7_1;
	wire w_dff_A_MAXA9IyN0_2;
	wire w_dff_A_bCaJ9rnB5_2;
	wire w_dff_A_iyvIJL261_2;
	wire w_dff_A_jKmKaN8m1_2;
	wire w_dff_A_i0ZiWJD53_2;
	wire w_dff_A_wjUNbkYd0_2;
	wire w_dff_A_NrRqS20P0_2;
	wire w_dff_A_bESZbtfo6_2;
	wire w_dff_A_mO5uSkrM3_0;
	wire w_dff_A_ZBKepXBW4_0;
	wire w_dff_A_iYAmN6LJ7_0;
	wire w_dff_A_yaXvQ9sw2_0;
	wire w_dff_A_hM2aoxTy5_0;
	wire w_dff_A_K8RBRrLP4_0;
	wire w_dff_A_PBBSU47T0_0;
	wire w_dff_A_AQyWoWVP1_0;
	wire w_dff_B_Ts3otrzS6_0;
	wire w_dff_B_6AipjvpJ7_0;
	wire w_dff_B_p6SyBldd6_0;
	wire w_dff_A_QTP6IFPs4_0;
	wire w_dff_A_d8ZqSQZm5_0;
	wire w_dff_A_wMZJN35v9_0;
	wire w_dff_A_X6eRaYX78_0;
	wire w_dff_A_HEsdDwwn8_2;
	wire w_dff_A_Jw8bTo2j2_2;
	wire w_dff_A_6pFHfPs42_2;
	wire w_dff_A_SVAwRhBm6_2;
	wire w_dff_A_qQHNDwii7_2;
	wire w_dff_A_yWMPujIT7_0;
	wire w_dff_A_AGG8RYi54_0;
	wire w_dff_A_ajWd8BSR1_0;
	wire w_dff_A_NUAbXkWe9_0;
	wire w_dff_A_7M8ANXzy7_0;
	wire w_dff_A_yD0VGvYK8_1;
	wire w_dff_A_FgeEyTeZ8_1;
	wire w_dff_A_1tBzBOUQ3_1;
	wire w_dff_A_j2xZuIC02_1;
	wire w_dff_A_yeHP93kZ5_1;
	wire w_dff_A_x3c0XfEU5_1;
	wire w_dff_A_m4k7EtwD6_1;
	wire w_dff_A_BdwHBUHD2_2;
	wire w_dff_A_KMn96lEg1_2;
	wire w_dff_A_CY8P0kfJ7_2;
	wire w_dff_A_WSKquXtZ5_2;
	wire w_dff_A_nNQ9DpNP8_2;
	wire w_dff_A_MTZAPu169_2;
	wire w_dff_A_szDrL2Wm8_2;
	wire w_dff_A_Z1jsBvNe5_2;
	wire w_dff_A_KmZYAzur6_2;
	wire w_dff_A_cHBGzICT0_2;
	wire w_dff_A_rP3rK1Vr4_2;
	wire w_dff_A_ECHHZQPu9_1;
	wire w_dff_A_XoYtyOy69_1;
	wire w_dff_A_a07NDFPc2_1;
	wire w_dff_A_FH4QgV1M8_1;
	wire w_dff_A_cM7tMsys0_1;
	wire w_dff_A_jvyYKYyr3_1;
	wire w_dff_A_qjnqF0wv6_1;
	wire w_dff_A_XaSQRJzn9_1;
	wire w_dff_A_t8uQFiOZ9_1;
	wire w_dff_B_zM4IdtOI4_0;
	wire w_dff_B_vUYxz9TH0_0;
	wire w_dff_B_yNPXiZOq1_0;
	wire w_dff_B_b3prPnl21_0;
	wire w_dff_A_LRt7OTZo0_0;
	wire w_dff_A_DFPhiLNs1_2;
	wire w_dff_A_yRtBaMq77_2;
	wire w_dff_A_v4FSawgS7_2;
	wire w_dff_A_nlkU6uhQ0_0;
	wire w_dff_A_A9E8vdJ38_2;
	wire w_dff_A_RDYRiz6I3_0;
	wire w_dff_A_bibeQP7Q3_0;
	wire w_dff_A_49kWzJ3N9_0;
	wire w_dff_A_vRztP4pg7_1;
	wire w_dff_A_QhYn5t4m1_1;
	wire w_dff_B_zvOTUrU43_2;
	wire w_dff_B_Zt7zWCQB8_2;
	wire w_dff_B_pL2mCnru0_2;
	wire w_dff_B_ds0xvXlA6_2;
	wire w_dff_B_ZRw0s8gv8_0;
	wire w_dff_A_jbDHMsX74_0;
	wire w_dff_A_WXECFDTI9_0;
	wire w_dff_B_7pT4tBQP9_0;
	wire w_dff_A_8DmXtU3j6_1;
	wire w_dff_A_iI9RsNaw6_1;
	wire w_dff_A_HavkOJJE6_1;
	wire w_dff_A_bywnkVAZ2_1;
	wire w_dff_A_i8iMz5ip7_1;
	wire w_dff_A_3vyI5rie3_1;
	wire w_dff_A_JzK7kycc4_1;
	wire w_dff_A_qtEIuVFu9_1;
	wire w_dff_A_EDqdme8J4_1;
	wire w_dff_A_oOBWseRU9_1;
	wire w_dff_A_be5oHboV7_1;
	wire w_dff_A_YZrrfRrS1_1;
	wire w_dff_A_nayQiYXK3_1;
	wire w_dff_A_9tSlHmkX2_1;
	wire w_dff_A_0OEzxPyU6_1;
	wire w_dff_A_Jr6sG1Ph8_1;
	wire w_dff_A_izl34Adi5_1;
	wire w_dff_A_RHfp2CIP1_1;
	wire w_dff_A_ryF2tkFQ7_1;
	wire w_dff_A_qRKbhJJt7_1;
	wire w_dff_A_1E524EgH1_2;
	wire w_dff_A_5DUnFiR40_2;
	wire w_dff_A_GkJHd3ou9_2;
	wire w_dff_A_zIU79f7v9_2;
	wire w_dff_A_AwXPWF3r1_2;
	wire w_dff_A_moQLh0bi9_2;
	wire w_dff_A_zDzKJnBE0_2;
	wire w_dff_A_wkhht0JW4_2;
	wire w_dff_A_zjRwJyqb7_2;
	wire w_dff_A_jtDD79jW1_2;
	wire w_dff_A_sBkbIeom1_2;
	wire w_dff_A_X0kHbAdb7_2;
	wire w_dff_A_GuAOCVhn2_0;
	wire w_dff_A_LKlLEh6J0_0;
	wire w_dff_A_QY1HNHBJ4_0;
	wire w_dff_A_aW2Db9OB6_0;
	wire w_dff_A_ppDEx3IG8_0;
	wire w_dff_A_hBXJmn1q4_0;
	wire w_dff_A_FcZzibNF5_0;
	wire w_dff_A_RjGobxKk6_0;
	wire w_dff_A_KLsQ9dIp4_0;
	wire w_dff_A_RvwfMsgN3_0;
	wire w_dff_A_7tU4sIsA9_0;
	wire w_dff_A_aZ6oFDTS2_0;
	wire w_dff_A_jrV05aOS6_0;
	wire w_dff_A_6q7s0qdu3_0;
	wire w_dff_A_nkt1lD8z7_0;
	wire w_dff_A_eNFRzgiG5_0;
	wire w_dff_A_ITEFn8wP3_0;
	wire w_dff_A_7i9jumX77_0;
	wire w_dff_A_Y1nK9cE15_2;
	wire w_dff_A_pxVP3Bml5_0;
	wire w_dff_A_uS7IE3Xd3_0;
	wire w_dff_A_xBieCWyF6_0;
	wire w_dff_A_vZnXxdw23_0;
	wire w_dff_A_DhjSzHIZ5_0;
	wire w_dff_A_q8JscRw53_0;
	wire w_dff_A_HT3gbkfU4_0;
	wire w_dff_A_qXGm286t0_0;
	wire w_dff_A_jO4U8LkB2_0;
	wire w_dff_A_HIBjT0qA1_0;
	wire w_dff_A_BtI0d3MF4_0;
	wire w_dff_A_S9KIXEaX7_0;
	wire w_dff_A_rlDvStwN0_0;
	wire w_dff_A_vUSHjRba9_0;
	wire w_dff_A_XySDXnhr5_0;
	wire w_dff_A_rchMZ7zR7_0;
	wire w_dff_A_52z0K9tC3_0;
	wire w_dff_A_8dNA4qOz6_0;
	wire w_dff_A_ZXpPQbxW2_2;
	wire w_dff_A_OTiqX9dw5_0;
	wire w_dff_A_pTDW5cen9_0;
	wire w_dff_A_zhlrvFaz9_0;
	wire w_dff_A_EKQQIoI42_0;
	wire w_dff_A_p3CTsA2X3_0;
	wire w_dff_A_0tBTn4xp7_0;
	wire w_dff_A_x4uE6wDa7_0;
	wire w_dff_A_188jnfxY0_0;
	wire w_dff_A_vfiaz7JC2_0;
	wire w_dff_A_0QEDlCjd3_0;
	wire w_dff_A_2CcnYQGP6_0;
	wire w_dff_A_M45ZyP6K8_0;
	wire w_dff_A_jy5KxXSS5_0;
	wire w_dff_A_AkCJCekU5_0;
	wire w_dff_A_vhmXD8te8_0;
	wire w_dff_A_5ntqW6Wo7_0;
	wire w_dff_A_f6hGMEQq3_0;
	wire w_dff_A_cJAURovK3_0;
	wire w_dff_A_SpizB91N3_2;
	wire w_dff_A_wFiDbO0J6_0;
	wire w_dff_A_k1Y13Y8V4_0;
	wire w_dff_A_b1VoSuUE0_0;
	wire w_dff_A_vWAO6IYk0_0;
	wire w_dff_A_1A2nlKG22_0;
	wire w_dff_A_IicdvabJ4_0;
	wire w_dff_A_I8ekCjS71_0;
	wire w_dff_A_peuVB3pl6_0;
	wire w_dff_A_UlI71KH61_0;
	wire w_dff_A_vauKkLvB3_0;
	wire w_dff_A_gZPnn3N70_0;
	wire w_dff_A_RmHT7Dty3_0;
	wire w_dff_A_zUP43K6b4_0;
	wire w_dff_A_7iflffAH3_0;
	wire w_dff_A_7qbnZ8U06_0;
	wire w_dff_A_8Soj1kAF1_0;
	wire w_dff_A_IZgVQmPA7_0;
	wire w_dff_A_jAQp9lAk2_0;
	wire w_dff_A_DTCDeFvN1_0;
	wire w_dff_A_DaA0Cm0b8_2;
	wire w_dff_A_kcvgynvC2_0;
	wire w_dff_A_pVzYYPWE4_0;
	wire w_dff_A_udigj5878_0;
	wire w_dff_A_AmwrHkzk7_0;
	wire w_dff_A_CpqIqHEB8_0;
	wire w_dff_A_gOD43Cmg6_0;
	wire w_dff_A_THoY87Un0_0;
	wire w_dff_A_kxVaw1Yf9_0;
	wire w_dff_A_X58358Id2_0;
	wire w_dff_A_321Hbrh97_0;
	wire w_dff_A_GVXUdRe55_0;
	wire w_dff_A_VCRxQNCe3_0;
	wire w_dff_A_Vtr8G3At1_0;
	wire w_dff_A_b8SS2enS3_0;
	wire w_dff_A_r9khn0Sj8_0;
	wire w_dff_A_kK4gBzNY9_0;
	wire w_dff_A_gm97eV5i6_0;
	wire w_dff_A_076S63OU4_0;
	wire w_dff_A_Q7Y9z1ZK3_2;
	wire w_dff_A_HzPxqt1Z6_0;
	wire w_dff_A_U6M9yE166_0;
	wire w_dff_A_YNdaR6bh9_0;
	wire w_dff_A_9Cy8yFQN2_0;
	wire w_dff_A_dQvVwmBJ9_0;
	wire w_dff_A_K9H0oYzO8_0;
	wire w_dff_A_XeIn005r7_0;
	wire w_dff_A_HRA0lOJY5_0;
	wire w_dff_A_ZnsDw7zE3_0;
	wire w_dff_A_HVRVC1VK8_0;
	wire w_dff_A_geW4UDfo4_0;
	wire w_dff_A_BKRIBCOx6_0;
	wire w_dff_A_7Tn18E0L6_0;
	wire w_dff_A_kHreSdkd2_0;
	wire w_dff_A_lkLcpaEg1_0;
	wire w_dff_A_uwCUJgbf2_0;
	wire w_dff_A_PC6qmYf30_2;
	wire w_dff_A_0FdV3wTW3_0;
	wire w_dff_A_Z8nbjcKD3_0;
	wire w_dff_A_z6pwVCWP5_0;
	wire w_dff_A_2ZC5W0XD0_0;
	wire w_dff_A_pDR1iKwO0_0;
	wire w_dff_A_uxUs2PCY8_0;
	wire w_dff_A_8I4fbpua4_0;
	wire w_dff_A_aTCXI97f2_0;
	wire w_dff_A_CR55BGBM5_0;
	wire w_dff_A_jSRamrSx0_0;
	wire w_dff_A_9hCgF8fD4_0;
	wire w_dff_A_qML2Jkjc9_0;
	wire w_dff_A_TCjHZf5d7_0;
	wire w_dff_A_kanGzhW38_0;
	wire w_dff_A_GEWHvxaL8_0;
	wire w_dff_A_52Fa1Yns7_0;
	wire w_dff_A_rLmSjeJg4_0;
	wire w_dff_A_KVpRZNKx4_2;
	wire w_dff_A_Rhynn9945_0;
	wire w_dff_A_wigCtVz05_0;
	wire w_dff_A_YKYRJEAY4_0;
	wire w_dff_A_RYjya74O8_0;
	wire w_dff_A_1caixoAE3_0;
	wire w_dff_A_gDP94gmv7_0;
	wire w_dff_A_rgVVfYiv7_0;
	wire w_dff_A_d2BtERMW8_0;
	wire w_dff_A_l7NK7DFj6_0;
	wire w_dff_A_iMxUOqYy0_0;
	wire w_dff_A_Ocz9z1wh1_0;
	wire w_dff_A_zj7HAygN9_0;
	wire w_dff_A_JBKPhhKh7_0;
	wire w_dff_A_jEc1bim20_0;
	wire w_dff_A_BFp5owVO5_0;
	wire w_dff_A_QNVKxMMM6_0;
	wire w_dff_A_yg0VlKrA6_0;
	wire w_dff_A_e8sPWf7F8_2;
	wire w_dff_A_SI057U6r4_0;
	wire w_dff_A_nA3S8Bqt0_0;
	wire w_dff_A_qdFba6oH0_0;
	wire w_dff_A_0kFxVnYG9_0;
	wire w_dff_A_dePyAu5j6_0;
	wire w_dff_A_0jL7wY0t2_0;
	wire w_dff_A_WDyrjHUh8_0;
	wire w_dff_A_HQy7LTtE8_0;
	wire w_dff_A_drtiOR7H3_0;
	wire w_dff_A_okes5AJ46_0;
	wire w_dff_A_OLSXyivU0_0;
	wire w_dff_A_zBpAOFK81_0;
	wire w_dff_A_xHrPpOCF5_0;
	wire w_dff_A_mPN3NODv5_0;
	wire w_dff_A_z7J8qGh39_0;
	wire w_dff_A_lmZZyiBz7_0;
	wire w_dff_A_aprmP46e1_0;
	wire w_dff_A_398D8Blp3_2;
	wire w_dff_A_9xtsT3pm2_0;
	wire w_dff_A_2t4rJmJw5_0;
	wire w_dff_A_iBunZqcK2_0;
	wire w_dff_A_IPn94Egd6_0;
	wire w_dff_A_EioGrX3Z4_0;
	wire w_dff_A_4rqMQxgh1_0;
	wire w_dff_A_lsF9shlh8_0;
	wire w_dff_A_Teh4GM4H0_0;
	wire w_dff_A_Un5Z3Ob27_0;
	wire w_dff_A_nCXLlWfk0_0;
	wire w_dff_A_ascmzqmL6_0;
	wire w_dff_A_PJrSBVSY8_0;
	wire w_dff_A_zN488CAe4_0;
	wire w_dff_A_I7IoKrtQ2_0;
	wire w_dff_A_SnGkx1gH4_0;
	wire w_dff_A_KRmvczNF6_0;
	wire w_dff_A_3qMyA9P25_0;
	wire w_dff_A_4EjUyHLf3_0;
	wire w_dff_A_K9PJEWpm2_2;
	wire w_dff_A_OjT0IQyU4_0;
	wire w_dff_A_Wo8dyX5s4_0;
	wire w_dff_A_QdI9JvV67_0;
	wire w_dff_A_F2VvoqcI3_0;
	wire w_dff_A_LDyGWqCN4_0;
	wire w_dff_A_VqeBgFVJ2_0;
	wire w_dff_A_9RROfpFx0_0;
	wire w_dff_A_7modmixP5_0;
	wire w_dff_A_6ngXizyP7_0;
	wire w_dff_A_SURhRANd5_0;
	wire w_dff_A_J99FjoF71_0;
	wire w_dff_A_r3vJIeo42_0;
	wire w_dff_A_GET4LZId2_0;
	wire w_dff_A_1dCwUPHy5_0;
	wire w_dff_A_RUQd7QgF4_0;
	wire w_dff_A_XNxCifA49_0;
	wire w_dff_A_4aE1HHNH6_1;
	wire w_dff_A_I9x3h4qN1_0;
	wire w_dff_A_5ibh62iE0_0;
	wire w_dff_A_1T43lxQM8_0;
	wire w_dff_A_dnb8rUiS2_0;
	wire w_dff_A_WPd6hMJ60_0;
	wire w_dff_A_k2fvyJjP1_0;
	wire w_dff_A_WgwIgCm09_0;
	wire w_dff_A_4RU2KqSQ4_0;
	wire w_dff_A_A9ztUOAT4_0;
	wire w_dff_A_Cr7eBnNh4_0;
	wire w_dff_A_wciQpmws5_0;
	wire w_dff_A_peBbtvtG6_0;
	wire w_dff_A_MSP2qFW88_0;
	wire w_dff_A_60hFFASs2_0;
	wire w_dff_A_mvOK2W9h7_0;
	wire w_dff_A_EKKJA5do1_0;
	wire w_dff_A_HGE1uK6W9_0;
	wire w_dff_A_zmegFpcB2_0;
	wire w_dff_A_up1EhJML0_2;
	wire w_dff_A_IjVS0GVL5_0;
	wire w_dff_A_aHk1J1aU1_0;
	wire w_dff_A_yXgFXQGu6_0;
	wire w_dff_A_iwvqaTI53_0;
	wire w_dff_A_xtUb4BHg8_0;
	wire w_dff_A_w33NIjZJ6_0;
	wire w_dff_A_aafD2M4u7_0;
	wire w_dff_A_UiTCakOA9_0;
	wire w_dff_A_7gVl9CFj9_0;
	wire w_dff_A_5SSV1iub4_0;
	wire w_dff_A_8LJkgOP54_0;
	wire w_dff_A_xgwledVq0_0;
	wire w_dff_A_rck1oucl5_0;
	wire w_dff_A_XweZXmXJ1_0;
	wire w_dff_A_W3dLmgUe1_0;
	wire w_dff_A_MkRBpyr40_0;
	wire w_dff_A_oaRMwzhY2_0;
	wire w_dff_A_csl3aRhX5_2;
	wire w_dff_A_mkY1nLu22_0;
	wire w_dff_A_XPMuzRkf4_0;
	wire w_dff_A_iySXuQF41_0;
	wire w_dff_A_1kUW6dBg2_0;
	wire w_dff_A_OjXFrgtr1_0;
	wire w_dff_A_864MDl3i8_0;
	wire w_dff_A_fEYCxMoo8_0;
	wire w_dff_A_dt74t9FM2_0;
	wire w_dff_A_JeZJ3xhm8_0;
	wire w_dff_A_EfRRtaOF5_0;
	wire w_dff_A_x9c69HAT5_0;
	wire w_dff_A_5zFJQRLR1_0;
	wire w_dff_A_UtEUmA5r4_0;
	wire w_dff_A_uVEAPLAS1_0;
	wire w_dff_A_niKJqv7r5_0;
	wire w_dff_A_2NM1ELsb7_0;
	wire w_dff_A_eRsuRZUc0_0;
	wire w_dff_A_CrUGfiSX7_2;
	wire w_dff_A_gQCgLpuQ3_0;
	wire w_dff_A_wp5znw2A7_0;
	wire w_dff_A_00R8rm1m6_0;
	wire w_dff_A_TFxh5nxS0_0;
	wire w_dff_A_IsILClwD4_0;
	wire w_dff_A_5HHzlktf9_0;
	wire w_dff_A_0O1rlOkM9_0;
	wire w_dff_A_1b1w5zwa7_0;
	wire w_dff_A_ZOeJBvtb0_0;
	wire w_dff_A_kEVaACIG0_0;
	wire w_dff_A_nlOkYiMg2_0;
	wire w_dff_A_oq6czHbW5_0;
	wire w_dff_A_08gBmKcK0_0;
	wire w_dff_A_f5aOjsHf0_0;
	wire w_dff_A_PHgt0RCM2_0;
	wire w_dff_A_nNZP1V5O0_0;
	wire w_dff_A_32HHgdDc0_0;
	wire w_dff_A_svC8UNFs8_0;
	wire w_dff_A_xsrmNVkq7_2;
	wire w_dff_A_uaor30g26_0;
	wire w_dff_A_Im3bDWIN7_0;
	wire w_dff_A_3G9WnZxV1_0;
	wire w_dff_A_JPLBFfI53_0;
	wire w_dff_A_QflP8YtV6_0;
	wire w_dff_A_fbfY82HE3_0;
	wire w_dff_A_IlpauXBo3_0;
	wire w_dff_A_viuvkxgk6_0;
	wire w_dff_A_QVyTf5I20_0;
	wire w_dff_A_aMpIvDcO3_0;
	wire w_dff_A_hV6sMuhr8_0;
	wire w_dff_A_20bCMobo8_0;
	wire w_dff_A_CugvgRr46_0;
	wire w_dff_A_sJmRVQDw9_0;
	wire w_dff_A_As6zZmd30_0;
	wire w_dff_A_0IlwTYZ81_0;
	wire w_dff_A_4vD5BJ2U0_2;
	wire w_dff_A_2Sfk8hZq5_0;
	wire w_dff_A_pWu2FU9w1_0;
	wire w_dff_A_0eEcsSck5_0;
	wire w_dff_A_DtIC18th4_0;
	wire w_dff_A_6Pw5vc0f1_0;
	wire w_dff_A_ZzdwRnFU3_0;
	wire w_dff_A_L6iLODd12_0;
	wire w_dff_A_4MpTUQrL9_0;
	wire w_dff_A_1QrvILdF1_0;
	wire w_dff_A_2SuZKbSr9_0;
	wire w_dff_A_Hzkem6hU8_0;
	wire w_dff_A_qUN49Yui5_0;
	wire w_dff_A_SC76EtqL9_0;
	wire w_dff_A_UEJG2x9F1_0;
	wire w_dff_A_CUal9O1N1_0;
	wire w_dff_A_ROsCN0oV9_0;
	wire w_dff_A_7W4PhO7b3_2;
	wire w_dff_A_gX40HpxM5_0;
	wire w_dff_A_aYieiXnk6_0;
	wire w_dff_A_J21VZuxz4_0;
	wire w_dff_A_YoqysCiO4_0;
	wire w_dff_A_ht8ABj3t4_0;
	wire w_dff_A_SCKs2Omb9_0;
	wire w_dff_A_EGj3SVRD2_0;
	wire w_dff_A_mgcnRDmm4_2;
	wire w_dff_A_y1E9JOjN1_0;
	wire w_dff_A_utUMXrRq9_0;
	wire w_dff_A_nO3QnoHq0_0;
	wire w_dff_A_VWu5r75i1_2;
	wire w_dff_A_wq0l5bdW9_0;
	wire w_dff_A_pTdiBhOH3_0;
	wire w_dff_A_j82oyDVy1_0;
	wire w_dff_A_yKfR0GGH1_2;
	wire w_dff_A_sworGvl53_0;
	wire w_dff_A_cUuhVVoP3_0;
	wire w_dff_A_z1oCuJhh8_0;
	wire w_dff_A_uqNWdzWx9_0;
	wire w_dff_A_NUrM0tWc5_0;
	wire w_dff_A_k24t8EOj8_2;
	wire w_dff_A_sr7IBH1k9_0;
	wire w_dff_A_4uviTJyN4_2;
	wire w_dff_A_bCGK6ity0_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_X0kHbAdb7_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_Y1nK9cE15_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_SpizB91N3_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_G17gat_2[2]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_n92_0[2]),.dout(w_dff_A_DaA0Cm0b8_2),.clk(gclk));
	jnot g009(.din(w_n93_0[0]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G1gat_1[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G26gat_0[1]),.dout(n97),.clk(gclk));
	jor g012(.dina(n97),.dinb(w_n96_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(w_n98_0[1]),.dinb(n95),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_Q7Y9z1ZK3_2),.clk(gclk));
	jnot g015(.din(w_G80gat_0[1]),.dout(n101),.clk(gclk));
	jand g016(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n102),.clk(gclk));
	jnot g017(.din(w_n102_0[1]),.dout(n103),.clk(gclk));
	jor g018(.dina(n103),.dinb(w_n101_0[1]),.dout(w_dff_A_PC6qmYf30_2),.clk(gclk));
	jnot g019(.din(w_G36gat_0[0]),.dout(n105),.clk(gclk));
	jnot g020(.din(w_G59gat_1[0]),.dout(n106),.clk(gclk));
	jor g021(.dina(w_n106_0[1]),.dinb(n105),.dout(n107),.clk(gclk));
	jor g022(.dina(w_n107_0[1]),.dinb(w_n101_0[0]),.dout(w_dff_A_KVpRZNKx4_2),.clk(gclk));
	jnot g023(.din(w_G42gat_1[2]),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n107_0[0]),.dinb(w_dff_B_imBdP2hB7_1),.dout(w_dff_A_e8sPWf7F8_2),.clk(gclk));
	jor g025(.dina(G88gat),.dinb(G87gat),.dout(n111),.clk(gclk));
	jand g026(.dina(w_n111_0[1]),.dinb(w_dff_B_bSewn0At8_1),.dout(w_dff_A_398D8Blp3_2),.clk(gclk));
	jnot g027(.din(w_G390gat_0[0]),.dout(n113),.clk(gclk));
	jor g028(.dina(w_n99_0[0]),.dinb(n113),.dout(w_dff_A_K9PJEWpm2_2),.clk(gclk));
	jand g029(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n115),.clk(gclk));
	jand g030(.dina(n115),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g031(.dina(w_G55gat_0[2]),.dinb(w_G13gat_0[0]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_n92_0[1]),.dout(n118),.clk(gclk));
	jand g033(.dina(w_G68gat_0[1]),.dinb(w_G29gat_0[0]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_dff_B_p1spw8vZ3_0),.dinb(w_n118_0[2]),.dout(w_dff_A_up1EhJML0_2),.clk(gclk));
	jand g035(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n121),.clk(gclk));
	jand g036(.dina(w_n121_0[1]),.dinb(w_dff_B_0SVk7vvA0_1),.dout(n122),.clk(gclk));
	jand g037(.dina(n122),.dinb(w_n118_0[1]),.dout(w_dff_A_csl3aRhX5_2),.clk(gclk));
	jand g038(.dina(w_n111_0[0]),.dinb(w_dff_B_grGLpViM1_1),.dout(w_dff_A_CrUGfiSX7_2),.clk(gclk));
	jxor g039(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n125),.clk(gclk));
	jxor g040(.dina(n125),.dinb(w_G130gat_0[1]),.dout(n126),.clk(gclk));
	jxor g041(.dina(w_G126gat_0[1]),.dinb(w_G121gat_0[2]),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_dff_B_B5B76rGU8_0),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g043(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n129),.clk(gclk));
	jxor g044(.dina(n129),.dinb(w_dff_B_rhfo69NT1_1),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(w_dff_B_Ph8WKAOg1_0),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n128),.dout(w_dff_A_xsrmNVkq7_2),.clk(gclk));
	jxor g048(.dina(w_G165gat_2[1]),.dinb(w_G159gat_2[1]),.dout(n134),.clk(gclk));
	jxor g049(.dina(n134),.dinb(w_G130gat_0[0]),.dout(n135),.clk(gclk));
	jxor g050(.dina(w_G201gat_2[2]),.dinb(w_G195gat_2[1]),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_dff_B_gaEppACI8_0),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g052(.dina(w_G189gat_2[1]),.dinb(w_G183gat_2[1]),.dout(n138),.clk(gclk));
	jxor g053(.dina(n138),.dinb(w_dff_B_qHOAPsD99_1),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G177gat_2[1]),.dinb(w_G171gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(w_dff_B_0Ti6aoJG7_0),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n137),.dout(w_dff_A_4vD5BJ2U0_2),.clk(gclk));
	jnot g057(.din(w_G261gat_0[2]),.dout(n143),.clk(gclk));
	jand g058(.dina(w_n102_0[0]),.dinb(w_G42gat_1[1]),.dout(n144),.clk(gclk));
	jnot g059(.din(n144),.dout(n145),.clk(gclk));
	jand g060(.dina(w_G51gat_1[0]),.dinb(w_G17gat_2[1]),.dout(n146),.clk(gclk));
	jand g061(.dina(n146),.dinb(w_n92_0[0]),.dout(n147),.clk(gclk));
	jand g062(.dina(w_dff_B_7pT4tBQP9_0),.dinb(n145),.dout(n148),.clk(gclk));
	jand g063(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n149),.clk(gclk));
	jxor g064(.dina(w_G42gat_1[0]),.dinb(w_G17gat_2[0]),.dout(n150),.clk(gclk));
	jand g065(.dina(n150),.dinb(w_n149_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(n151),.dinb(w_G447gat_1),.dout(n152),.clk(gclk));
	jor g067(.dina(w_dff_B_ZRw0s8gv8_0),.dinb(n148),.dout(n153),.clk(gclk));
	jand g068(.dina(w_n153_3[1]),.dinb(w_G126gat_0[0]),.dout(n154),.clk(gclk));
	jnot g069(.din(w_G156gat_0[0]),.dout(n155),.clk(gclk));
	jor g070(.dina(n155),.dinb(w_n106_0[0]),.dout(n156),.clk(gclk));
	jand g071(.dina(n156),.dinb(w_G447gat_0[2]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n157_0[1]),.dinb(w_G17gat_1[2]),.dout(n158),.clk(gclk));
	jor g073(.dina(n158),.dinb(w_n96_0[0]),.dout(n159),.clk(gclk));
	jand g074(.dina(w_n159_1[1]),.dinb(w_G153gat_0[2]),.dout(n160),.clk(gclk));
	jand g075(.dina(w_n86_0[0]),.dinb(w_G80gat_0[0]),.dout(n161),.clk(gclk));
	jand g076(.dina(n161),.dinb(w_G447gat_0[1]),.dout(n162),.clk(gclk));
	jnot g077(.din(w_G268gat_0[1]),.dout(n163),.clk(gclk));
	jand g078(.dina(w_n163_0[1]),.dinb(w_G55gat_0[1]),.dout(n164),.clk(gclk));
	jand g079(.dina(w_dff_B_8kWAgWBF9_0),.dinb(w_n162_0[1]),.dout(n165),.clk(gclk));
	jor g080(.dina(w_n165_1[2]),.dinb(n160),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n154_0[1]),.dout(n167),.clk(gclk));
	jxor g082(.dina(w_n167_1[1]),.dinb(w_G201gat_2[1]),.dout(n168),.clk(gclk));
	jnot g083(.din(w_n168_0[2]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n143_0[1]),.dout(n170),.clk(gclk));
	jor g085(.dina(w_n168_0[1]),.dinb(w_G261gat_0[1]),.dout(n171),.clk(gclk));
	jand g086(.dina(n171),.dinb(w_G219gat_3[1]),.dout(n172),.clk(gclk));
	jand g087(.dina(n172),.dinb(n170),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n168_0[0]),.dinb(w_G228gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_G237gat_3[1]),.dinb(w_G201gat_2[0]),.dout(n175),.clk(gclk));
	jor g090(.dina(n175),.dinb(w_G246gat_3[1]),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_e4tEbFwq7_0),.dinb(w_n167_1[0]),.dout(n177),.clk(gclk));
	jand g092(.dina(G72gat),.dinb(w_G42gat_0[2]),.dout(n178),.clk(gclk));
	jand g093(.dina(n178),.dinb(w_dff_B_vTI34gNP8_1),.dout(n179),.clk(gclk));
	jand g094(.dina(n179),.dinb(w_n121_0[0]),.dout(n180),.clk(gclk));
	jand g095(.dina(n180),.dinb(w_n118_0[0]),.dout(n181),.clk(gclk));
	jand g096(.dina(w_n181_3[1]),.dinb(w_G201gat_1[2]),.dout(n182),.clk(gclk));
	jand g097(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n183),.clk(gclk));
	jand g098(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(n184),.dinb(n183),.dout(n185),.clk(gclk));
	jor g100(.dina(w_dff_B_1Ckw5jTi5_0),.dinb(n182),.dout(n186),.clk(gclk));
	jor g101(.dina(w_dff_B_AzrEMCtS5_0),.dinb(n177),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(n174),.dout(n188),.clk(gclk));
	jor g103(.dina(w_dff_B_YGClbl2b5_0),.dinb(n173),.dout(w_dff_A_7W4PhO7b3_2),.clk(gclk));
	jand g104(.dina(w_n159_1[0]),.dinb(w_G143gat_0[1]),.dout(n190),.clk(gclk));
	jand g105(.dina(w_n153_3[0]),.dinb(w_G111gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(n191),.dinb(w_n165_1[1]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_dff_B_DGX4PC4T2_1),.dout(n193),.clk(gclk));
	jxor g108(.dina(w_n193_1[1]),.dinb(w_G183gat_2[0]),.dout(n194),.clk(gclk));
	jnot g109(.din(w_n194_0[2]),.dout(n195),.clk(gclk));
	jand g110(.dina(w_n167_0[2]),.dinb(w_G201gat_1[1]),.dout(n196),.clk(gclk));
	jnot g111(.din(w_n196_0[1]),.dout(n197),.clk(gclk));
	jnot g112(.din(w_G201gat_1[0]),.dout(n198),.clk(gclk));
	jnot g113(.din(w_n154_0[0]),.dout(n199),.clk(gclk));
	jnot g114(.din(w_G153gat_0[1]),.dout(n200),.clk(gclk));
	jnot g115(.din(w_G17gat_1[1]),.dout(n201),.clk(gclk));
	jnot g116(.din(w_G51gat_0[2]),.dout(n202),.clk(gclk));
	jor g117(.dina(w_n98_0[0]),.dinb(w_dff_B_CEyhQme00_1),.dout(n203),.clk(gclk));
	jor g118(.dina(w_n149_0[0]),.dinb(n203),.dout(n204),.clk(gclk));
	jor g119(.dina(n204),.dinb(w_dff_B_zcWU9T686_1),.dout(n205),.clk(gclk));
	jand g120(.dina(n205),.dinb(w_G1gat_0[1]),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_308swCCT8_1),.dout(n207),.clk(gclk));
	jnot g122(.din(w_n165_1[0]),.dout(n208),.clk(gclk));
	jand g123(.dina(w_dff_B_teIs8hoA6_0),.dinb(n207),.dout(n209),.clk(gclk));
	jand g124(.dina(n209),.dinb(w_dff_B_CRE4zai05_1),.dout(n210),.clk(gclk));
	jand g125(.dina(n210),.dinb(w_dff_B_skd7gkZr8_1),.dout(n211),.clk(gclk));
	jor g126(.dina(n211),.dinb(w_n143_0[0]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_Bj9Xhqiq0_1),.dout(n213),.clk(gclk));
	jand g128(.dina(w_n159_0[2]),.dinb(w_G146gat_0[1]),.dout(n214),.clk(gclk));
	jand g129(.dina(w_n153_2[2]),.dinb(w_G116gat_0[1]),.dout(n215),.clk(gclk));
	jor g130(.dina(n215),.dinb(w_n165_0[2]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_dff_B_HP1pRa9y2_1),.dout(n217),.clk(gclk));
	jor g132(.dina(w_n217_1[1]),.dinb(w_G189gat_2[0]),.dout(n218),.clk(gclk));
	jand g133(.dina(w_n159_0[1]),.dinb(w_G149gat_0[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n153_2[1]),.dinb(w_G121gat_0[0]),.dout(n220),.clk(gclk));
	jor g135(.dina(n220),.dinb(w_n165_0[1]),.dout(n221),.clk(gclk));
	jor g136(.dina(n221),.dinb(w_dff_B_rRvGpYtZ9_1),.dout(n222),.clk(gclk));
	jor g137(.dina(w_n222_1[1]),.dinb(w_G195gat_2[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n223_0[1]),.dinb(w_n218_0[1]),.dout(n224),.clk(gclk));
	jnot g139(.din(w_n224_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_7A8CQ8wf1_0),.dinb(w_n213_0[1]),.dout(n226),.clk(gclk));
	jand g141(.dina(w_n217_1[0]),.dinb(w_G189gat_1[2]),.dout(n227),.clk(gclk));
	jand g142(.dina(w_n222_1[0]),.dinb(w_G195gat_1[2]),.dout(n228),.clk(gclk));
	jand g143(.dina(w_n228_0[1]),.dinb(w_n218_0[0]),.dout(n229),.clk(gclk));
	jor g144(.dina(n229),.dinb(w_dff_B_HJhhk2Za1_1),.dout(n230),.clk(gclk));
	jnot g145(.din(w_n230_0[1]),.dout(n231),.clk(gclk));
	jand g146(.dina(w_dff_B_zCTWHUUc0_0),.dinb(n226),.dout(n232),.clk(gclk));
	jor g147(.dina(w_n232_0[1]),.dinb(w_dff_B_OnGJBMIS9_1),.dout(n233),.clk(gclk));
	jor g148(.dina(w_n167_0[1]),.dinb(w_G201gat_0[2]),.dout(n234),.clk(gclk));
	jand g149(.dina(n234),.dinb(w_G261gat_0[0]),.dout(n235),.clk(gclk));
	jor g150(.dina(n235),.dinb(w_n196_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n224_0[0]),.dinb(w_n236_0[2]),.dout(n237),.clk(gclk));
	jor g152(.dina(w_n230_0[0]),.dinb(n237),.dout(n238),.clk(gclk));
	jor g153(.dina(w_n238_0[1]),.dinb(w_n194_0[1]),.dout(n239),.clk(gclk));
	jand g154(.dina(n239),.dinb(w_G219gat_3[0]),.dout(n240),.clk(gclk));
	jand g155(.dina(n240),.dinb(n233),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n194_0[0]),.dinb(w_G228gat_3[0]),.dout(n242),.clk(gclk));
	jand g157(.dina(w_G237gat_3[0]),.dinb(w_G183gat_1[2]),.dout(n243),.clk(gclk));
	jor g158(.dina(n243),.dinb(w_G246gat_3[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(w_dff_B_PkuvAbhw4_0),.dinb(w_n193_1[0]),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n181_3[0]),.dinb(w_G183gat_1[1]),.dout(n246),.clk(gclk));
	jand g161(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n247),.clk(gclk));
	jor g162(.dina(w_dff_B_TBYpJrwa5_0),.dinb(n246),.dout(n248),.clk(gclk));
	jor g163(.dina(w_dff_B_gbJbg8IZ7_0),.dinb(n245),.dout(n249),.clk(gclk));
	jor g164(.dina(n249),.dinb(n242),.dout(n250),.clk(gclk));
	jor g165(.dina(w_dff_B_AHzH8W2L4_0),.dinb(n241),.dout(w_dff_A_mgcnRDmm4_2),.clk(gclk));
	jxor g166(.dina(w_n217_0[2]),.dinb(w_G189gat_1[1]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n252_0[2]),.dout(n253),.clk(gclk));
	jand g168(.dina(w_n223_0[0]),.dinb(w_n236_0[1]),.dout(n254),.clk(gclk));
	jor g169(.dina(n254),.dinb(w_n228_0[0]),.dout(n255),.clk(gclk));
	jnot g170(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jor g171(.dina(n256),.dinb(w_dff_B_5g2hOEDC3_1),.dout(n257),.clk(gclk));
	jor g172(.dina(w_n255_0[0]),.dinb(w_n252_0[1]),.dout(n258),.clk(gclk));
	jand g173(.dina(n258),.dinb(w_G219gat_2[2]),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(n257),.dout(n260),.clk(gclk));
	jand g175(.dina(w_n252_0[0]),.dinb(w_G228gat_2[2]),.dout(n261),.clk(gclk));
	jand g176(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n262),.clk(gclk));
	jor g177(.dina(n262),.dinb(w_G246gat_2[2]),.dout(n263),.clk(gclk));
	jand g178(.dina(w_dff_B_AHbSZy1E6_0),.dinb(w_n217_0[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(w_n181_2[2]),.dinb(w_G189gat_0[2]),.dout(n265),.clk(gclk));
	jand g180(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n266),.clk(gclk));
	jand g181(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n267),.clk(gclk));
	jor g182(.dina(n267),.dinb(n266),.dout(n268),.clk(gclk));
	jor g183(.dina(w_dff_B_MniE1BeU3_0),.dinb(n265),.dout(n269),.clk(gclk));
	jor g184(.dina(w_dff_B_Z8JMqWBH9_0),.dinb(n264),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(n261),.dout(n271),.clk(gclk));
	jor g186(.dina(w_dff_B_Azjf68mi8_0),.dinb(n260),.dout(w_dff_A_VWu5r75i1_2),.clk(gclk));
	jxor g187(.dina(w_n222_0[2]),.dinb(w_G195gat_1[1]),.dout(n273),.clk(gclk));
	jnot g188(.din(w_n273_0[2]),.dout(n274),.clk(gclk));
	jor g189(.dina(w_dff_B_htQwsgFs6_0),.dinb(w_n213_0[0]),.dout(n275),.clk(gclk));
	jor g190(.dina(w_n273_0[1]),.dinb(w_n236_0[0]),.dout(n276),.clk(gclk));
	jand g191(.dina(n276),.dinb(w_G219gat_2[1]),.dout(n277),.clk(gclk));
	jand g192(.dina(n277),.dinb(n275),.dout(n278),.clk(gclk));
	jand g193(.dina(w_n273_0[0]),.dinb(w_G228gat_2[1]),.dout(n279),.clk(gclk));
	jand g194(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(n280),.dinb(w_G246gat_2[1]),.dout(n281),.clk(gclk));
	jand g196(.dina(w_dff_B_NLR683bv2_0),.dinb(w_n222_0[1]),.dout(n282),.clk(gclk));
	jand g197(.dina(w_n181_2[1]),.dinb(w_G195gat_0[2]),.dout(n283),.clk(gclk));
	jand g198(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n284),.clk(gclk));
	jand g199(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n285),.clk(gclk));
	jor g200(.dina(n285),.dinb(n284),.dout(n286),.clk(gclk));
	jor g201(.dina(w_dff_B_UbIOBVj62_0),.dinb(n283),.dout(n287),.clk(gclk));
	jor g202(.dina(w_dff_B_mM67qCh82_0),.dinb(n282),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(n279),.dout(n289),.clk(gclk));
	jor g204(.dina(w_dff_B_mXZ9OooB6_0),.dinb(n278),.dout(w_dff_A_yKfR0GGH1_2),.clk(gclk));
	jand g205(.dina(w_n153_2[0]),.dinb(w_G91gat_0[1]),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n157_0[0]),.dinb(w_G55gat_0[0]),.dout(n292),.clk(gclk));
	jand g207(.dina(w_n292_1[1]),.dinb(w_G143gat_0[0]),.dout(n293),.clk(gclk));
	jand g208(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n294),.clk(gclk));
	jand g209(.dina(w_n163_0[0]),.dinb(w_G17gat_1[0]),.dout(n295),.clk(gclk));
	jand g210(.dina(w_dff_B_b3prPnl21_0),.dinb(w_n162_0[0]),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n296_1[1]),.dinb(w_dff_B_nBOiScYI3_1),.dout(n297),.clk(gclk));
	jor g212(.dina(n297),.dinb(n293),.dout(n298),.clk(gclk));
	jor g213(.dina(n298),.dinb(n291),.dout(n299),.clk(gclk));
	jand g214(.dina(w_n299_1[1]),.dinb(w_G159gat_2[0]),.dout(n300),.clk(gclk));
	jor g215(.dina(w_n299_1[0]),.dinb(w_G159gat_1[2]),.dout(n301),.clk(gclk));
	jand g216(.dina(w_n193_0[2]),.dinb(w_G183gat_1[0]),.dout(n302),.clk(gclk));
	jor g217(.dina(w_n193_0[1]),.dinb(w_G183gat_0[2]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n238_0[0]),.dinb(w_n303_0[1]),.dout(n304),.clk(gclk));
	jor g219(.dina(n304),.dinb(w_n302_0[1]),.dout(n305),.clk(gclk));
	jnot g220(.din(w_G165gat_2[0]),.dout(n306),.clk(gclk));
	jand g221(.dina(w_n153_1[2]),.dinb(w_G96gat_0[1]),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n292_1[0]),.dinb(w_G146gat_0[0]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_i5cAmkLc7_0),.dinb(w_n296_1[0]),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(n308),.dout(n311),.clk(gclk));
	jor g226(.dina(n311),.dinb(n307),.dout(n312),.clk(gclk));
	jnot g227(.din(w_n312_1[1]),.dout(n313),.clk(gclk));
	jand g228(.dina(n313),.dinb(w_dff_B_pRJznE1q4_1),.dout(n314),.clk(gclk));
	jnot g229(.din(n314),.dout(n315),.clk(gclk));
	jand g230(.dina(w_n153_1[1]),.dinb(w_G101gat_0[1]),.dout(n316),.clk(gclk));
	jand g231(.dina(w_n292_0[2]),.dinb(w_G149gat_0[0]),.dout(n317),.clk(gclk));
	jand g232(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n318),.clk(gclk));
	jor g233(.dina(w_dff_B_yNPXiZOq1_0),.dinb(w_n296_0[2]),.dout(n319),.clk(gclk));
	jor g234(.dina(n319),.dinb(n317),.dout(n320),.clk(gclk));
	jor g235(.dina(n320),.dinb(n316),.dout(n321),.clk(gclk));
	jor g236(.dina(w_n321_1[1]),.dinb(w_G171gat_2[0]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n153_1[0]),.dinb(w_G106gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_n292_0[1]),.dinb(w_G153gat_0[0]),.dout(n324),.clk(gclk));
	jand g239(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_p6SyBldd6_0),.dinb(w_n296_0[1]),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g242(.dina(n327),.dinb(n323),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n328_1[1]),.dinb(w_G177gat_2[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n329_0[2]),.dinb(w_n322_0[1]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n330_0[2]),.dinb(w_n315_0[1]),.dout(n331),.clk(gclk));
	jand g246(.dina(w_n331_0[1]),.dinb(w_n305_1[1]),.dout(n332),.clk(gclk));
	jand g247(.dina(w_n312_1[0]),.dinb(w_G165gat_1[2]),.dout(n333),.clk(gclk));
	jand g248(.dina(w_n321_1[0]),.dinb(w_G171gat_1[2]),.dout(n334),.clk(gclk));
	jand g249(.dina(w_n328_1[0]),.dinb(w_G177gat_1[2]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_0[2]),.dinb(w_n322_0[0]),.dout(n336),.clk(gclk));
	jor g251(.dina(n336),.dinb(w_dff_B_lkdbdiPE2_1),.dout(n337),.clk(gclk));
	jand g252(.dina(w_n337_0[2]),.dinb(w_n315_0[0]),.dout(n338),.clk(gclk));
	jor g253(.dina(n338),.dinb(w_dff_B_6W5xi0fm4_1),.dout(n339),.clk(gclk));
	jor g254(.dina(w_n339_0[1]),.dinb(n332),.dout(n340),.clk(gclk));
	jand g255(.dina(w_n340_0[1]),.dinb(w_dff_B_bCNiqDY01_1),.dout(n341),.clk(gclk));
	jor g256(.dina(n341),.dinb(w_dff_B_Vu62d98T6_1),.dout(w_dff_A_k24t8EOj8_2),.clk(gclk));
	jnot g257(.din(w_n302_0[0]),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n303_0[0]),.dout(n344),.clk(gclk));
	jor g259(.dina(w_n232_0[0]),.dinb(w_dff_B_BU8RXXAE6_1),.dout(n345),.clk(gclk));
	jand g260(.dina(n345),.dinb(w_dff_B_FxFBpVrk9_1),.dout(n346),.clk(gclk));
	jxor g261(.dina(w_n328_0[2]),.dinb(w_G177gat_1[1]),.dout(n347),.clk(gclk));
	jnot g262(.din(w_n347_0[2]),.dout(n348),.clk(gclk));
	jor g263(.dina(w_dff_B_ZATPpVoE5_0),.dinb(w_n346_1[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(w_n347_0[1]),.dinb(w_n305_1[0]),.dout(n350),.clk(gclk));
	jand g265(.dina(n350),.dinb(w_G219gat_2[0]),.dout(n351),.clk(gclk));
	jand g266(.dina(n351),.dinb(n349),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n347_0[0]),.dinb(w_G228gat_2[0]),.dout(n353),.clk(gclk));
	jand g268(.dina(w_G237gat_2[0]),.dinb(w_G177gat_1[0]),.dout(n354),.clk(gclk));
	jor g269(.dina(n354),.dinb(w_G246gat_2[0]),.dout(n355),.clk(gclk));
	jand g270(.dina(w_dff_B_939bfeFA6_0),.dinb(w_n328_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n181_2[0]),.dinb(w_G177gat_0[2]),.dout(n357),.clk(gclk));
	jand g272(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n358),.clk(gclk));
	jor g273(.dina(w_dff_B_XSfu6jy41_0),.dinb(n357),.dout(n359),.clk(gclk));
	jor g274(.dina(w_dff_B_vwu3chqa7_0),.dinb(n356),.dout(n360),.clk(gclk));
	jor g275(.dina(n360),.dinb(n353),.dout(n361),.clk(gclk));
	jor g276(.dina(w_dff_B_TaQMXKwf6_0),.dinb(n352),.dout(w_dff_A_4uviTJyN4_2),.clk(gclk));
	jnot g277(.din(w_n331_0[0]),.dout(n363),.clk(gclk));
	jor g278(.dina(w_dff_B_LpuWcMhc0_0),.dinb(w_n346_1[0]),.dout(n364),.clk(gclk));
	jnot g279(.din(w_n339_0[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_dff_B_WjlhjVFz8_0),.dinb(n364),.dout(n366),.clk(gclk));
	jxor g281(.dina(w_n299_0[2]),.dinb(w_G159gat_1[1]),.dout(n367),.clk(gclk));
	jnot g282(.din(w_n367_0[2]),.dout(n368),.clk(gclk));
	jor g283(.dina(w_dff_B_PNoVvop11_0),.dinb(n366),.dout(n369),.clk(gclk));
	jor g284(.dina(w_n367_0[1]),.dinb(w_n340_0[0]),.dout(n370),.clk(gclk));
	jand g285(.dina(n370),.dinb(w_G219gat_1[2]),.dout(n371),.clk(gclk));
	jand g286(.dina(n371),.dinb(n369),.dout(n372),.clk(gclk));
	jand g287(.dina(w_n367_0[0]),.dinb(w_G228gat_1[2]),.dout(n373),.clk(gclk));
	jand g288(.dina(w_G237gat_1[2]),.dinb(w_G159gat_1[0]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_G246gat_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(w_dff_B_Wh4Yu1TF4_0),.dinb(w_n299_0[1]),.dout(n376),.clk(gclk));
	jand g291(.dina(w_n181_1[2]),.dinb(w_G159gat_0[2]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n378),.clk(gclk));
	jor g293(.dina(w_dff_B_jjcIAjEI9_0),.dinb(n377),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_MIHLAari6_0),.dinb(n376),.dout(n380),.clk(gclk));
	jor g295(.dina(n380),.dinb(n373),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_Izf4783V0_0),.dinb(n372),.dout(G878gat),.clk(gclk));
	jxor g297(.dina(w_n312_0[2]),.dinb(w_G165gat_1[1]),.dout(n383),.clk(gclk));
	jnot g298(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n337_0[1]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n330_0[1]),.dout(n386),.clk(gclk));
	jor g301(.dina(w_dff_B_3XQtlWSc7_0),.dinb(w_n346_0[2]),.dout(n387),.clk(gclk));
	jand g302(.dina(n387),.dinb(w_dff_B_fkPCQbba7_1),.dout(n388),.clk(gclk));
	jor g303(.dina(n388),.dinb(w_dff_B_OelSTeiU1_1),.dout(n389),.clk(gclk));
	jand g304(.dina(w_n330_0[0]),.dinb(w_n305_0[2]),.dout(n390),.clk(gclk));
	jor g305(.dina(n390),.dinb(w_n337_0[0]),.dout(n391),.clk(gclk));
	jor g306(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_G219gat_1[1]),.dout(n393),.clk(gclk));
	jand g308(.dina(n393),.dinb(n389),.dout(n394),.clk(gclk));
	jand g309(.dina(w_n383_0[0]),.dinb(w_G228gat_1[1]),.dout(n395),.clk(gclk));
	jand g310(.dina(w_G237gat_1[1]),.dinb(w_G165gat_1[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(n396),.dinb(w_G246gat_1[1]),.dout(n397),.clk(gclk));
	jand g312(.dina(w_dff_B_GJ3Zrlbj5_0),.dinb(w_n312_0[1]),.dout(n398),.clk(gclk));
	jand g313(.dina(w_n181_1[1]),.dinb(w_G165gat_0[2]),.dout(n399),.clk(gclk));
	jand g314(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n400),.clk(gclk));
	jor g315(.dina(w_dff_B_qyXVzmYJ7_0),.dinb(n399),.dout(n401),.clk(gclk));
	jor g316(.dina(w_dff_B_2spQn6sk2_0),.dinb(n398),.dout(n402),.clk(gclk));
	jor g317(.dina(n402),.dinb(n395),.dout(n403),.clk(gclk));
	jor g318(.dina(w_dff_B_knFNQfaJ1_0),.dinb(n394),.dout(G879gat),.clk(gclk));
	jxor g319(.dina(w_n321_0[2]),.dinb(w_G171gat_1[1]),.dout(n405),.clk(gclk));
	jnot g320(.din(w_n405_0[2]),.dout(n406),.clk(gclk));
	jnot g321(.din(w_n335_0[1]),.dout(n407),.clk(gclk));
	jnot g322(.din(w_n329_0[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_L0320AkD2_0),.dinb(w_n346_0[1]),.dout(n409),.clk(gclk));
	jand g324(.dina(n409),.dinb(w_dff_B_QyXeecTJ0_1),.dout(n410),.clk(gclk));
	jor g325(.dina(n410),.dinb(w_dff_B_NLszNRtg2_1),.dout(n411),.clk(gclk));
	jand g326(.dina(w_n329_0[0]),.dinb(w_n305_0[1]),.dout(n412),.clk(gclk));
	jor g327(.dina(n412),.dinb(w_n335_0[0]),.dout(n413),.clk(gclk));
	jor g328(.dina(n413),.dinb(w_n405_0[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_G219gat_1[0]),.dout(n415),.clk(gclk));
	jand g330(.dina(n415),.dinb(n411),.dout(n416),.clk(gclk));
	jand g331(.dina(w_n405_0[0]),.dinb(w_G228gat_1[0]),.dout(n417),.clk(gclk));
	jand g332(.dina(w_G237gat_1[0]),.dinb(w_G171gat_1[0]),.dout(n418),.clk(gclk));
	jor g333(.dina(n418),.dinb(w_G246gat_1[0]),.dout(n419),.clk(gclk));
	jand g334(.dina(w_dff_B_Gm0kNzhg3_0),.dinb(w_n321_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n181_1[0]),.dinb(w_G171gat_0[2]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_Pv1yspMa9_0),.dinb(n421),.dout(n423),.clk(gclk));
	jor g338(.dina(w_dff_B_nBQKbeDD7_0),.dinb(n420),.dout(n424),.clk(gclk));
	jor g339(.dina(n424),.dinb(n417),.dout(n425),.clk(gclk));
	jor g340(.dina(w_dff_B_bBEt4ZWG5_0),.dinb(n416),.dout(G880gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_3vyI5rie3_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_G13gat_0[1]),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_LRt7OTZo0_0),.doutb(w_G17gat_1[1]),.doutc(w_dff_A_v4FSawgS7_2),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_G17gat_2[2]),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_G29gat_0[0]),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_qtEIuVFu9_1),.doutc(w_G42gat_0[2]),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_G42gat_1[0]),.doutb(w_dff_A_JzK7kycc4_1),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_8DmXtU3j6_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_49kWzJ3N9_0),.doutb(w_dff_A_vRztP4pg7_1),.doutc(w_G55gat_0[2]),.din(G55gat));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_G68gat_0[1]),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_nlkU6uhQ0_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_A9E8vdJ38_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_6LWhfFPr7_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_98YQrYo79_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_nayQiYXK3_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_7M8ANXzy7_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_uIjmtxar9_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_4J4xqKLW5_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_fyBPgIOs4_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl jspl_w_G126gat_0(.douta(w_dff_A_WeingIaf9_0),.doutb(w_G126gat_0[1]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_G130gat_0[1]),.din(w_dff_B_QgsYS31O1_2));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_XR9CSE6t7_1),.din(w_dff_B_SKyVliyN8_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_kvfY68hY2_1),.din(w_dff_B_piD0i7Xt2_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_QhYn5t4m1_1),.din(w_dff_B_ds0xvXlA6_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_X6eRaYX78_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_qQHNDwii7_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_G159gat_0[1]),.doutc(w_dff_A_Y7MJgL9w2_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_G159gat_1[0]),.doutb(w_dff_A_3CXBDjGy9_1),.doutc(w_dff_A_pFZYmTHO8_2),.din(w_G159gat_0[0]));
	jspl jspl_w_G159gat_2(.douta(w_dff_A_Gk5jogLs6_0),.doutb(w_G159gat_2[1]),.din(w_G159gat_0[1]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_G165gat_0[1]),.doutc(w_dff_A_8XpGyw5C6_2),.din(G165gat));
	jspl3 jspl3_w_G165gat_1(.douta(w_G165gat_1[0]),.doutb(w_dff_A_jc7HTzSh1_1),.doutc(w_dff_A_5KNPP9EU7_2),.din(w_G165gat_0[0]));
	jspl jspl_w_G165gat_2(.douta(w_G165gat_2[0]),.doutb(w_G165gat_2[1]),.din(w_G165gat_0[1]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_dff_A_sBkbIeom1_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_dff_A_qRKbhJJt7_1),.doutc(w_dff_A_zDzKJnBE0_2),.din(w_G171gat_0[0]));
	jspl jspl_w_G171gat_2(.douta(w_dff_A_KPkjkTHf0_0),.doutb(w_G171gat_2[1]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_G177gat_0[1]),.doutc(w_dff_A_rP3rK1Vr4_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_m4k7EtwD6_1),.doutc(w_dff_A_szDrL2Wm8_2),.din(w_G177gat_0[0]));
	jspl jspl_w_G177gat_2(.douta(w_dff_A_kPNf8Wh39_0),.doutb(w_G177gat_2[1]),.din(w_G177gat_0[1]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_bESZbtfo6_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_vSNtDbIa9_0),.doutb(w_dff_A_M3JOp4nt7_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl jspl_w_G183gat_2(.douta(w_dff_A_8UXupTrs7_0),.doutb(w_G183gat_2[1]),.din(w_G183gat_0[1]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_7awGszEe9_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_Bk71gHeV9_1),.doutc(w_dff_A_ihUrwOyU2_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_PNmlGw7p8_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_7tnFYHLD3_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_DTUD1R403_1),.doutc(w_dff_A_fsxYyJjG3_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_IpqDrjdh0_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_G201gat_0[1]),.doutc(w_dff_A_QZg04gcl8_2),.din(G201gat));
	jspl3 jspl3_w_G201gat_1(.douta(w_G201gat_1[0]),.doutb(w_dff_A_KCKcfahM1_1),.doutc(w_dff_A_bt1n3pah3_2),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G201gat_2(.douta(w_G201gat_2[0]),.doutb(w_dff_A_91NrIlWL9_1),.doutc(w_G201gat_2[2]),.din(w_G201gat_0[1]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_2WeA3owF7_0),.doutb(w_dff_A_j2mV2HVv6_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_ZL8ZAyZh2_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_G219gat_1[1]),.doutc(w_G219gat_1[2]),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_2ubPBvQG8_0),.doutb(w_G219gat_2[1]),.doutc(w_dff_A_Y0KSzmJG1_2),.din(w_G219gat_0[1]));
	jspl jspl_w_G219gat_3(.douta(w_dff_A_kfV1ScLC4_0),.doutb(w_G219gat_3[1]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.doutc(w_dff_A_JhAco3gd1_2),.din(w_dff_B_cunaExpD1_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_G228gat_2[0]),.doutb(w_dff_A_qpejjR656_1),.doutc(w_dff_A_ZGrPnzK36_2),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_G228gat_3[1]),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_G237gat_0[0]),.doutb(w_G237gat_0[1]),.doutc(w_G237gat_0[2]),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_G237gat_2[0]),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_G237gat_3[1]),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_G246gat_0[0]),.doutb(w_G246gat_0[1]),.doutc(w_G246gat_0[2]),.din(w_dff_B_0gjBhWBg7_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_G246gat_2[0]),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_G246gat_3[1]),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_EPD7r3wi6_0),.doutb(w_dff_A_fwjkoGRV6_1),.doutc(w_G261gat_0[2]),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_HGAmaQlw0_1),.doutc(w_dff_A_ZXpPQbxW2_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_G447gat_0[2]),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_4aE1HHNH6_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n96_0(.douta(w_dff_A_Wzfu0KCD4_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(w_dff_B_20dLN3zF8_2));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n118_0(.douta(w_dff_A_shD5mLGa3_0),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n121_0(.douta(w_dff_A_LxxNHobh5_0),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(w_dff_B_W8buxaVQ2_2));
	jspl jspl_w_n149_0(.douta(w_dff_A_WXECFDTI9_0),.doutb(w_n149_0[1]),.din(n149));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_n153_2[2]),.din(w_n153_0[1]));
	jspl jspl_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.din(w_n153_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_dff_A_WmCX4QAd4_1),.din(n154));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_rKyPGpVz7_1),.doutc(w_dff_A_w9FWJmsQ3_2),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_n165_1[0]),.doutb(w_dff_A_EftGHX5V2_1),.doutc(w_dff_A_vUIuLwci3_2),.din(w_n165_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n181_3(.douta(w_n181_3[0]),.doutb(w_n181_3[1]),.din(w_n181_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl jspl_w_n193_1(.douta(w_n193_1[0]),.doutb(w_n193_1[1]),.din(w_n193_0[0]));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_dff_A_zrKGkpZa4_1),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_dff_A_bSvZyBQD0_0),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl jspl_w_n217_1(.douta(w_n217_1[0]),.doutb(w_n217_1[1]),.din(w_n217_0[0]));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl jspl_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.din(w_n222_0[0]));
	jspl jspl_w_n223_0(.douta(w_dff_A_EEBKWNz20_0),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_dff_A_c2yYKDc01_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n228_0(.douta(w_dff_A_C4oHFx8z8_0),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_dff_A_U8VkxY2G1_0),.doutb(w_n230_0[1]),.din(n230));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.din(n238));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_9rSqPCBT7_1),.doutc(w_n252_0[2]),.din(n252));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_dff_A_XRHeV7YM6_1),.doutc(w_n273_0[2]),.din(n273));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n296_1(.douta(w_n296_1[0]),.doutb(w_n296_1[1]),.din(w_n296_0[0]));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl jspl_w_n299_1(.douta(w_n299_1[0]),.doutb(w_n299_1[1]),.din(w_n299_0[0]));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_dff_A_YWGPJBXF6_1),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_yqcEP5M88_1),.din(n303));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl jspl_w_n305_1(.douta(w_n305_1[0]),.doutb(w_n305_1[1]),.din(w_n305_0[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl jspl_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.din(w_n321_0[0]));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n328_1(.douta(w_n328_1[0]),.doutb(w_n328_1[1]),.din(w_n328_0[0]));
	jspl3 jspl3_w_n329_0(.douta(w_dff_A_kScFJcsb4_0),.doutb(w_n329_0[1]),.doutc(w_n329_0[2]),.din(n329));
	jspl3 jspl3_w_n330_0(.douta(w_dff_A_dfDj8RWL9_0),.doutb(w_n330_0[1]),.doutc(w_dff_A_KbcVS7sh7_2),.din(n330));
	jspl jspl_w_n331_0(.douta(w_n331_0[0]),.doutb(w_dff_A_W22bFRvE6_1),.din(n331));
	jspl3 jspl3_w_n335_0(.douta(w_dff_A_AQyWoWVP1_0),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n337_0(.douta(w_dff_A_wS7nXe1t7_0),.doutb(w_n337_0[1]),.doutc(w_n337_0[2]),.din(n337));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_dff_A_AbClJDsC1_1),.din(n339));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_3Y6MdOJP6_1),.doutc(w_n347_0[2]),.din(n347));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_dff_A_zguWoSTU8_1),.doutc(w_n367_0[2]),.din(n367));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_UJ7N9NOf9_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_dff_A_t8uQFiOZ9_1),.doutc(w_n405_0[2]),.din(n405));
	jdff dff_B_20dLN3zF8_2(.din(n101),.dout(w_dff_B_20dLN3zF8_2),.clk(gclk));
	jdff dff_B_imBdP2hB7_1(.din(n109),.dout(w_dff_B_imBdP2hB7_1),.clk(gclk));
	jdff dff_B_bSewn0At8_1(.din(G90gat),.dout(w_dff_B_bSewn0At8_1),.clk(gclk));
	jdff dff_A_HGAmaQlw0_1(.dout(w_G390gat_0[1]),.din(w_dff_A_HGAmaQlw0_1),.clk(gclk));
	jdff dff_B_p1spw8vZ3_0(.din(n119),.dout(w_dff_B_p1spw8vZ3_0),.clk(gclk));
	jdff dff_B_0SVk7vvA0_1(.din(G74gat),.dout(w_dff_B_0SVk7vvA0_1),.clk(gclk));
	jdff dff_B_grGLpViM1_1(.din(G89gat),.dout(w_dff_B_grGLpViM1_1),.clk(gclk));
	jdff dff_B_Ph8WKAOg1_0(.din(n131),.dout(w_dff_B_Ph8WKAOg1_0),.clk(gclk));
	jdff dff_B_rhfo69NT1_1(.din(G135gat),.dout(w_dff_B_rhfo69NT1_1),.clk(gclk));
	jdff dff_B_B5B76rGU8_0(.din(n127),.dout(w_dff_B_B5B76rGU8_0),.clk(gclk));
	jdff dff_B_0Ti6aoJG7_0(.din(n140),.dout(w_dff_B_0Ti6aoJG7_0),.clk(gclk));
	jdff dff_B_qHOAPsD99_1(.din(G207gat),.dout(w_dff_B_qHOAPsD99_1),.clk(gclk));
	jdff dff_B_gaEppACI8_0(.din(n136),.dout(w_dff_B_gaEppACI8_0),.clk(gclk));
	jdff dff_B_QgsYS31O1_2(.din(G130gat),.dout(w_dff_B_QgsYS31O1_2),.clk(gclk));
	jdff dff_B_YGClbl2b5_0(.din(n188),.dout(w_dff_B_YGClbl2b5_0),.clk(gclk));
	jdff dff_B_O4xtUkOQ4_0(.din(n186),.dout(w_dff_B_O4xtUkOQ4_0),.clk(gclk));
	jdff dff_B_ybglk5AV2_0(.din(w_dff_B_O4xtUkOQ4_0),.dout(w_dff_B_ybglk5AV2_0),.clk(gclk));
	jdff dff_B_AzrEMCtS5_0(.din(w_dff_B_ybglk5AV2_0),.dout(w_dff_B_AzrEMCtS5_0),.clk(gclk));
	jdff dff_B_p8U5SauZ6_0(.din(n185),.dout(w_dff_B_p8U5SauZ6_0),.clk(gclk));
	jdff dff_B_ixm5HORf2_0(.din(w_dff_B_p8U5SauZ6_0),.dout(w_dff_B_ixm5HORf2_0),.clk(gclk));
	jdff dff_B_1Ckw5jTi5_0(.din(w_dff_B_ixm5HORf2_0),.dout(w_dff_B_1Ckw5jTi5_0),.clk(gclk));
	jdff dff_B_9ONUZyXy5_0(.din(n176),.dout(w_dff_B_9ONUZyXy5_0),.clk(gclk));
	jdff dff_B_5sfbu1df6_0(.din(w_dff_B_9ONUZyXy5_0),.dout(w_dff_B_5sfbu1df6_0),.clk(gclk));
	jdff dff_B_gsRf9kRE5_0(.din(w_dff_B_5sfbu1df6_0),.dout(w_dff_B_gsRf9kRE5_0),.clk(gclk));
	jdff dff_B_ay7CdLwp0_0(.din(w_dff_B_gsRf9kRE5_0),.dout(w_dff_B_ay7CdLwp0_0),.clk(gclk));
	jdff dff_B_lCubPa2y6_0(.din(w_dff_B_ay7CdLwp0_0),.dout(w_dff_B_lCubPa2y6_0),.clk(gclk));
	jdff dff_B_e4tEbFwq7_0(.din(w_dff_B_lCubPa2y6_0),.dout(w_dff_B_e4tEbFwq7_0),.clk(gclk));
	jdff dff_A_uyBtC1KM4_1(.dout(w_G201gat_2[1]),.din(w_dff_A_uyBtC1KM4_1),.clk(gclk));
	jdff dff_A_d02kyb4O8_1(.dout(w_dff_A_uyBtC1KM4_1),.din(w_dff_A_d02kyb4O8_1),.clk(gclk));
	jdff dff_A_zG0SrBk54_1(.dout(w_dff_A_d02kyb4O8_1),.din(w_dff_A_zG0SrBk54_1),.clk(gclk));
	jdff dff_A_NsjjrEY33_1(.dout(w_dff_A_zG0SrBk54_1),.din(w_dff_A_NsjjrEY33_1),.clk(gclk));
	jdff dff_A_BU2ztQuX6_1(.dout(w_dff_A_NsjjrEY33_1),.din(w_dff_A_BU2ztQuX6_1),.clk(gclk));
	jdff dff_A_d5I7JrIA4_1(.dout(w_dff_A_BU2ztQuX6_1),.din(w_dff_A_d5I7JrIA4_1),.clk(gclk));
	jdff dff_A_y8SpNbTV6_1(.dout(w_dff_A_d5I7JrIA4_1),.din(w_dff_A_y8SpNbTV6_1),.clk(gclk));
	jdff dff_A_91NrIlWL9_1(.dout(w_dff_A_y8SpNbTV6_1),.din(w_dff_A_91NrIlWL9_1),.clk(gclk));
	jdff dff_B_gLJK9rfG7_0(.din(n250),.dout(w_dff_B_gLJK9rfG7_0),.clk(gclk));
	jdff dff_B_wqovFkR87_0(.din(w_dff_B_gLJK9rfG7_0),.dout(w_dff_B_wqovFkR87_0),.clk(gclk));
	jdff dff_B_IFrpMZ5N0_0(.din(w_dff_B_wqovFkR87_0),.dout(w_dff_B_IFrpMZ5N0_0),.clk(gclk));
	jdff dff_B_buhThgss7_0(.din(w_dff_B_IFrpMZ5N0_0),.dout(w_dff_B_buhThgss7_0),.clk(gclk));
	jdff dff_B_AHzH8W2L4_0(.din(w_dff_B_buhThgss7_0),.dout(w_dff_B_AHzH8W2L4_0),.clk(gclk));
	jdff dff_B_T8PDaqa59_0(.din(n248),.dout(w_dff_B_T8PDaqa59_0),.clk(gclk));
	jdff dff_B_GiovWExW0_0(.din(w_dff_B_T8PDaqa59_0),.dout(w_dff_B_GiovWExW0_0),.clk(gclk));
	jdff dff_B_gbJbg8IZ7_0(.din(w_dff_B_GiovWExW0_0),.dout(w_dff_B_gbJbg8IZ7_0),.clk(gclk));
	jdff dff_B_9pbRBZMr3_0(.din(n247),.dout(w_dff_B_9pbRBZMr3_0),.clk(gclk));
	jdff dff_B_5yE5FOPw1_0(.din(w_dff_B_9pbRBZMr3_0),.dout(w_dff_B_5yE5FOPw1_0),.clk(gclk));
	jdff dff_B_eny3aYSx1_0(.din(w_dff_B_5yE5FOPw1_0),.dout(w_dff_B_eny3aYSx1_0),.clk(gclk));
	jdff dff_B_TBYpJrwa5_0(.din(w_dff_B_eny3aYSx1_0),.dout(w_dff_B_TBYpJrwa5_0),.clk(gclk));
	jdff dff_B_LlKdc5LR6_0(.din(n244),.dout(w_dff_B_LlKdc5LR6_0),.clk(gclk));
	jdff dff_B_Lq3Kd2KJ5_0(.din(w_dff_B_LlKdc5LR6_0),.dout(w_dff_B_Lq3Kd2KJ5_0),.clk(gclk));
	jdff dff_B_Rhy7Vwpy6_0(.din(w_dff_B_Lq3Kd2KJ5_0),.dout(w_dff_B_Rhy7Vwpy6_0),.clk(gclk));
	jdff dff_B_0X2DTZyU9_0(.din(w_dff_B_Rhy7Vwpy6_0),.dout(w_dff_B_0X2DTZyU9_0),.clk(gclk));
	jdff dff_B_2KGvhXHX7_0(.din(w_dff_B_0X2DTZyU9_0),.dout(w_dff_B_2KGvhXHX7_0),.clk(gclk));
	jdff dff_B_PkuvAbhw4_0(.din(w_dff_B_2KGvhXHX7_0),.dout(w_dff_B_PkuvAbhw4_0),.clk(gclk));
	jdff dff_A_71SzKjgp3_0(.dout(w_G219gat_3[0]),.din(w_dff_A_71SzKjgp3_0),.clk(gclk));
	jdff dff_A_kMQa9KPt0_0(.dout(w_dff_A_71SzKjgp3_0),.din(w_dff_A_kMQa9KPt0_0),.clk(gclk));
	jdff dff_A_r5yEQohJ0_0(.dout(w_dff_A_kMQa9KPt0_0),.din(w_dff_A_r5yEQohJ0_0),.clk(gclk));
	jdff dff_A_kfV1ScLC4_0(.dout(w_dff_A_r5yEQohJ0_0),.din(w_dff_A_kfV1ScLC4_0),.clk(gclk));
	jdff dff_B_ARNxSAtR9_1(.din(n195),.dout(w_dff_B_ARNxSAtR9_1),.clk(gclk));
	jdff dff_B_44Lon0vO1_1(.din(w_dff_B_ARNxSAtR9_1),.dout(w_dff_B_44Lon0vO1_1),.clk(gclk));
	jdff dff_B_3aKBqgG15_1(.din(w_dff_B_44Lon0vO1_1),.dout(w_dff_B_3aKBqgG15_1),.clk(gclk));
	jdff dff_B_OnGJBMIS9_1(.din(w_dff_B_3aKBqgG15_1),.dout(w_dff_B_OnGJBMIS9_1),.clk(gclk));
	jdff dff_A_dqYIZIoN4_1(.dout(w_n194_0[1]),.din(w_dff_A_dqYIZIoN4_1),.clk(gclk));
	jdff dff_A_bPr74adn8_1(.dout(w_dff_A_dqYIZIoN4_1),.din(w_dff_A_bPr74adn8_1),.clk(gclk));
	jdff dff_A_2i2VcIGE8_1(.dout(w_dff_A_bPr74adn8_1),.din(w_dff_A_2i2VcIGE8_1),.clk(gclk));
	jdff dff_A_zrKGkpZa4_1(.dout(w_dff_A_2i2VcIGE8_1),.din(w_dff_A_zrKGkpZa4_1),.clk(gclk));
	jdff dff_A_3j60n8el0_0(.dout(w_G183gat_2[0]),.din(w_dff_A_3j60n8el0_0),.clk(gclk));
	jdff dff_A_KjYrMeKG1_0(.dout(w_dff_A_3j60n8el0_0),.din(w_dff_A_KjYrMeKG1_0),.clk(gclk));
	jdff dff_A_U55PGDX44_0(.dout(w_dff_A_KjYrMeKG1_0),.din(w_dff_A_U55PGDX44_0),.clk(gclk));
	jdff dff_A_p6xXJuug1_0(.dout(w_dff_A_U55PGDX44_0),.din(w_dff_A_p6xXJuug1_0),.clk(gclk));
	jdff dff_A_hHVkuQgB7_0(.dout(w_dff_A_p6xXJuug1_0),.din(w_dff_A_hHVkuQgB7_0),.clk(gclk));
	jdff dff_A_aumyIOC68_0(.dout(w_dff_A_hHVkuQgB7_0),.din(w_dff_A_aumyIOC68_0),.clk(gclk));
	jdff dff_A_zlP5GoH65_0(.dout(w_dff_A_aumyIOC68_0),.din(w_dff_A_zlP5GoH65_0),.clk(gclk));
	jdff dff_A_8UXupTrs7_0(.dout(w_dff_A_zlP5GoH65_0),.din(w_dff_A_8UXupTrs7_0),.clk(gclk));
	jdff dff_B_jKblZ1Io3_0(.din(n271),.dout(w_dff_B_jKblZ1Io3_0),.clk(gclk));
	jdff dff_B_4Oh6NWAF2_0(.din(w_dff_B_jKblZ1Io3_0),.dout(w_dff_B_4Oh6NWAF2_0),.clk(gclk));
	jdff dff_B_K1mWKtft0_0(.din(w_dff_B_4Oh6NWAF2_0),.dout(w_dff_B_K1mWKtft0_0),.clk(gclk));
	jdff dff_B_AC8deFa16_0(.din(w_dff_B_K1mWKtft0_0),.dout(w_dff_B_AC8deFa16_0),.clk(gclk));
	jdff dff_B_Azjf68mi8_0(.din(w_dff_B_AC8deFa16_0),.dout(w_dff_B_Azjf68mi8_0),.clk(gclk));
	jdff dff_B_PwwxRCIU4_0(.din(n269),.dout(w_dff_B_PwwxRCIU4_0),.clk(gclk));
	jdff dff_B_PKOBX8gL3_0(.din(w_dff_B_PwwxRCIU4_0),.dout(w_dff_B_PKOBX8gL3_0),.clk(gclk));
	jdff dff_B_Z8JMqWBH9_0(.din(w_dff_B_PKOBX8gL3_0),.dout(w_dff_B_Z8JMqWBH9_0),.clk(gclk));
	jdff dff_B_RGC0gZks6_0(.din(n268),.dout(w_dff_B_RGC0gZks6_0),.clk(gclk));
	jdff dff_B_2ewSbTsW5_0(.din(w_dff_B_RGC0gZks6_0),.dout(w_dff_B_2ewSbTsW5_0),.clk(gclk));
	jdff dff_B_MniE1BeU3_0(.din(w_dff_B_2ewSbTsW5_0),.dout(w_dff_B_MniE1BeU3_0),.clk(gclk));
	jdff dff_B_MPxPuv9U3_0(.din(n263),.dout(w_dff_B_MPxPuv9U3_0),.clk(gclk));
	jdff dff_B_1B1che8B6_0(.din(w_dff_B_MPxPuv9U3_0),.dout(w_dff_B_1B1che8B6_0),.clk(gclk));
	jdff dff_B_utPzGWY18_0(.din(w_dff_B_1B1che8B6_0),.dout(w_dff_B_utPzGWY18_0),.clk(gclk));
	jdff dff_B_hM4RozQr3_0(.din(w_dff_B_utPzGWY18_0),.dout(w_dff_B_hM4RozQr3_0),.clk(gclk));
	jdff dff_B_UNzA1csy7_0(.din(w_dff_B_hM4RozQr3_0),.dout(w_dff_B_UNzA1csy7_0),.clk(gclk));
	jdff dff_B_AHbSZy1E6_0(.din(w_dff_B_UNzA1csy7_0),.dout(w_dff_B_AHbSZy1E6_0),.clk(gclk));
	jdff dff_B_jlP1OLvK8_1(.din(n253),.dout(w_dff_B_jlP1OLvK8_1),.clk(gclk));
	jdff dff_B_sCrphbuU2_1(.din(w_dff_B_jlP1OLvK8_1),.dout(w_dff_B_sCrphbuU2_1),.clk(gclk));
	jdff dff_B_LSni4cBE7_1(.din(w_dff_B_sCrphbuU2_1),.dout(w_dff_B_LSni4cBE7_1),.clk(gclk));
	jdff dff_B_5g2hOEDC3_1(.din(w_dff_B_LSni4cBE7_1),.dout(w_dff_B_5g2hOEDC3_1),.clk(gclk));
	jdff dff_A_GrPBqO918_1(.dout(w_n252_0[1]),.din(w_dff_A_GrPBqO918_1),.clk(gclk));
	jdff dff_A_bnscJa248_1(.dout(w_dff_A_GrPBqO918_1),.din(w_dff_A_bnscJa248_1),.clk(gclk));
	jdff dff_A_DxyktazZ8_1(.dout(w_dff_A_bnscJa248_1),.din(w_dff_A_DxyktazZ8_1),.clk(gclk));
	jdff dff_A_9rSqPCBT7_1(.dout(w_dff_A_DxyktazZ8_1),.din(w_dff_A_9rSqPCBT7_1),.clk(gclk));
	jdff dff_B_e5bnfAO46_0(.din(n289),.dout(w_dff_B_e5bnfAO46_0),.clk(gclk));
	jdff dff_B_bkPu8vnq1_0(.din(w_dff_B_e5bnfAO46_0),.dout(w_dff_B_bkPu8vnq1_0),.clk(gclk));
	jdff dff_B_mXZ9OooB6_0(.din(w_dff_B_bkPu8vnq1_0),.dout(w_dff_B_mXZ9OooB6_0),.clk(gclk));
	jdff dff_B_Yf4oWFVd6_0(.din(n287),.dout(w_dff_B_Yf4oWFVd6_0),.clk(gclk));
	jdff dff_B_7Nw6Hepr2_0(.din(w_dff_B_Yf4oWFVd6_0),.dout(w_dff_B_7Nw6Hepr2_0),.clk(gclk));
	jdff dff_B_mM67qCh82_0(.din(w_dff_B_7Nw6Hepr2_0),.dout(w_dff_B_mM67qCh82_0),.clk(gclk));
	jdff dff_B_HOwL5CEw0_0(.din(n286),.dout(w_dff_B_HOwL5CEw0_0),.clk(gclk));
	jdff dff_B_ovZcmco80_0(.din(w_dff_B_HOwL5CEw0_0),.dout(w_dff_B_ovZcmco80_0),.clk(gclk));
	jdff dff_B_UbIOBVj62_0(.din(w_dff_B_ovZcmco80_0),.dout(w_dff_B_UbIOBVj62_0),.clk(gclk));
	jdff dff_B_EDmjy9Uf2_0(.din(n281),.dout(w_dff_B_EDmjy9Uf2_0),.clk(gclk));
	jdff dff_B_CKNTQsoL2_0(.din(w_dff_B_EDmjy9Uf2_0),.dout(w_dff_B_CKNTQsoL2_0),.clk(gclk));
	jdff dff_B_BLQanJGl2_0(.din(w_dff_B_CKNTQsoL2_0),.dout(w_dff_B_BLQanJGl2_0),.clk(gclk));
	jdff dff_B_XHEiAOyR0_0(.din(w_dff_B_BLQanJGl2_0),.dout(w_dff_B_XHEiAOyR0_0),.clk(gclk));
	jdff dff_B_8BqY0Q968_0(.din(w_dff_B_XHEiAOyR0_0),.dout(w_dff_B_8BqY0Q968_0),.clk(gclk));
	jdff dff_B_NLR683bv2_0(.din(w_dff_B_8BqY0Q968_0),.dout(w_dff_B_NLR683bv2_0),.clk(gclk));
	jdff dff_B_4Uma8bE48_0(.din(n274),.dout(w_dff_B_4Uma8bE48_0),.clk(gclk));
	jdff dff_B_htQwsgFs6_0(.din(w_dff_B_4Uma8bE48_0),.dout(w_dff_B_htQwsgFs6_0),.clk(gclk));
	jdff dff_A_HLvrnQlk3_1(.dout(w_n273_0[1]),.din(w_dff_A_HLvrnQlk3_1),.clk(gclk));
	jdff dff_A_XRHeV7YM6_1(.dout(w_dff_A_HLvrnQlk3_1),.din(w_dff_A_XRHeV7YM6_1),.clk(gclk));
	jdff dff_B_9xZT2iRI4_1(.din(n300),.dout(w_dff_B_9xZT2iRI4_1),.clk(gclk));
	jdff dff_B_pHcCZFPs0_1(.din(w_dff_B_9xZT2iRI4_1),.dout(w_dff_B_pHcCZFPs0_1),.clk(gclk));
	jdff dff_B_vRnS05bD7_1(.din(w_dff_B_pHcCZFPs0_1),.dout(w_dff_B_vRnS05bD7_1),.clk(gclk));
	jdff dff_B_nwHzjng78_1(.din(w_dff_B_vRnS05bD7_1),.dout(w_dff_B_nwHzjng78_1),.clk(gclk));
	jdff dff_B_Zawc3RUZ2_1(.din(w_dff_B_nwHzjng78_1),.dout(w_dff_B_Zawc3RUZ2_1),.clk(gclk));
	jdff dff_B_taifWXKy4_1(.din(w_dff_B_Zawc3RUZ2_1),.dout(w_dff_B_taifWXKy4_1),.clk(gclk));
	jdff dff_B_aWax5gil0_1(.din(w_dff_B_taifWXKy4_1),.dout(w_dff_B_aWax5gil0_1),.clk(gclk));
	jdff dff_B_ekJRrZl70_1(.din(w_dff_B_aWax5gil0_1),.dout(w_dff_B_ekJRrZl70_1),.clk(gclk));
	jdff dff_B_FJtONLbG5_1(.din(w_dff_B_ekJRrZl70_1),.dout(w_dff_B_FJtONLbG5_1),.clk(gclk));
	jdff dff_B_Vu62d98T6_1(.din(w_dff_B_FJtONLbG5_1),.dout(w_dff_B_Vu62d98T6_1),.clk(gclk));
	jdff dff_B_x8TNGM6s2_1(.din(n301),.dout(w_dff_B_x8TNGM6s2_1),.clk(gclk));
	jdff dff_B_bmBLbOZ03_1(.din(w_dff_B_x8TNGM6s2_1),.dout(w_dff_B_bmBLbOZ03_1),.clk(gclk));
	jdff dff_B_E54BZqYM6_1(.din(w_dff_B_bmBLbOZ03_1),.dout(w_dff_B_E54BZqYM6_1),.clk(gclk));
	jdff dff_B_QG6DV6Jm6_1(.din(w_dff_B_E54BZqYM6_1),.dout(w_dff_B_QG6DV6Jm6_1),.clk(gclk));
	jdff dff_B_ZZklmh1s0_1(.din(w_dff_B_QG6DV6Jm6_1),.dout(w_dff_B_ZZklmh1s0_1),.clk(gclk));
	jdff dff_B_ht8GZpwO0_1(.din(w_dff_B_ZZklmh1s0_1),.dout(w_dff_B_ht8GZpwO0_1),.clk(gclk));
	jdff dff_B_91k8CrMr2_1(.din(w_dff_B_ht8GZpwO0_1),.dout(w_dff_B_91k8CrMr2_1),.clk(gclk));
	jdff dff_B_Gu84OHbr3_1(.din(w_dff_B_91k8CrMr2_1),.dout(w_dff_B_Gu84OHbr3_1),.clk(gclk));
	jdff dff_B_bCNiqDY01_1(.din(w_dff_B_Gu84OHbr3_1),.dout(w_dff_B_bCNiqDY01_1),.clk(gclk));
	jdff dff_A_zOBPkLcQ4_0(.dout(w_G159gat_2[0]),.din(w_dff_A_zOBPkLcQ4_0),.clk(gclk));
	jdff dff_A_MWDaFW5U3_0(.dout(w_dff_A_zOBPkLcQ4_0),.din(w_dff_A_MWDaFW5U3_0),.clk(gclk));
	jdff dff_A_EH6Ydh4c5_0(.dout(w_dff_A_MWDaFW5U3_0),.din(w_dff_A_EH6Ydh4c5_0),.clk(gclk));
	jdff dff_A_W3Rzjnlm1_0(.dout(w_dff_A_EH6Ydh4c5_0),.din(w_dff_A_W3Rzjnlm1_0),.clk(gclk));
	jdff dff_A_YUbiW5946_0(.dout(w_dff_A_W3Rzjnlm1_0),.din(w_dff_A_YUbiW5946_0),.clk(gclk));
	jdff dff_A_QxkZQQRA3_0(.dout(w_dff_A_YUbiW5946_0),.din(w_dff_A_QxkZQQRA3_0),.clk(gclk));
	jdff dff_A_Gk5jogLs6_0(.dout(w_dff_A_QxkZQQRA3_0),.din(w_dff_A_Gk5jogLs6_0),.clk(gclk));
	jdff dff_B_8FQ52lYY8_0(.din(n361),.dout(w_dff_B_8FQ52lYY8_0),.clk(gclk));
	jdff dff_B_IX1kvsFC3_0(.din(w_dff_B_8FQ52lYY8_0),.dout(w_dff_B_IX1kvsFC3_0),.clk(gclk));
	jdff dff_B_RcHhDRc17_0(.din(w_dff_B_IX1kvsFC3_0),.dout(w_dff_B_RcHhDRc17_0),.clk(gclk));
	jdff dff_B_l8StTNXe4_0(.din(w_dff_B_RcHhDRc17_0),.dout(w_dff_B_l8StTNXe4_0),.clk(gclk));
	jdff dff_B_pXwGRbk69_0(.din(w_dff_B_l8StTNXe4_0),.dout(w_dff_B_pXwGRbk69_0),.clk(gclk));
	jdff dff_B_hZSntnMI9_0(.din(w_dff_B_pXwGRbk69_0),.dout(w_dff_B_hZSntnMI9_0),.clk(gclk));
	jdff dff_B_WFQYmM1L3_0(.din(w_dff_B_hZSntnMI9_0),.dout(w_dff_B_WFQYmM1L3_0),.clk(gclk));
	jdff dff_B_TaQMXKwf6_0(.din(w_dff_B_WFQYmM1L3_0),.dout(w_dff_B_TaQMXKwf6_0),.clk(gclk));
	jdff dff_B_QRwLWZYo2_0(.din(n359),.dout(w_dff_B_QRwLWZYo2_0),.clk(gclk));
	jdff dff_B_vwu3chqa7_0(.din(w_dff_B_QRwLWZYo2_0),.dout(w_dff_B_vwu3chqa7_0),.clk(gclk));
	jdff dff_B_9JYDDdE36_0(.din(n358),.dout(w_dff_B_9JYDDdE36_0),.clk(gclk));
	jdff dff_B_smpALfaa5_0(.din(w_dff_B_9JYDDdE36_0),.dout(w_dff_B_smpALfaa5_0),.clk(gclk));
	jdff dff_B_iJ5QzUeg2_0(.din(w_dff_B_smpALfaa5_0),.dout(w_dff_B_iJ5QzUeg2_0),.clk(gclk));
	jdff dff_B_XSfu6jy41_0(.din(w_dff_B_iJ5QzUeg2_0),.dout(w_dff_B_XSfu6jy41_0),.clk(gclk));
	jdff dff_B_iq5ceS9A8_0(.din(n355),.dout(w_dff_B_iq5ceS9A8_0),.clk(gclk));
	jdff dff_B_3I4pFtGl9_0(.din(w_dff_B_iq5ceS9A8_0),.dout(w_dff_B_3I4pFtGl9_0),.clk(gclk));
	jdff dff_B_bjeD6pub3_0(.din(w_dff_B_3I4pFtGl9_0),.dout(w_dff_B_bjeD6pub3_0),.clk(gclk));
	jdff dff_B_7KXbOgVN3_0(.din(w_dff_B_bjeD6pub3_0),.dout(w_dff_B_7KXbOgVN3_0),.clk(gclk));
	jdff dff_B_939bfeFA6_0(.din(w_dff_B_7KXbOgVN3_0),.dout(w_dff_B_939bfeFA6_0),.clk(gclk));
	jdff dff_A_qpejjR656_1(.dout(w_G228gat_2[1]),.din(w_dff_A_qpejjR656_1),.clk(gclk));
	jdff dff_A_ZGrPnzK36_2(.dout(w_G228gat_2[2]),.din(w_dff_A_ZGrPnzK36_2),.clk(gclk));
	jdff dff_A_azNFpMhM8_0(.dout(w_G219gat_2[0]),.din(w_dff_A_azNFpMhM8_0),.clk(gclk));
	jdff dff_A_e7CKnUIu7_0(.dout(w_dff_A_azNFpMhM8_0),.din(w_dff_A_e7CKnUIu7_0),.clk(gclk));
	jdff dff_A_T9jjpiEI2_0(.dout(w_dff_A_e7CKnUIu7_0),.din(w_dff_A_T9jjpiEI2_0),.clk(gclk));
	jdff dff_A_2ubPBvQG8_0(.dout(w_dff_A_T9jjpiEI2_0),.din(w_dff_A_2ubPBvQG8_0),.clk(gclk));
	jdff dff_A_dY5lbPeH2_2(.dout(w_G219gat_2[2]),.din(w_dff_A_dY5lbPeH2_2),.clk(gclk));
	jdff dff_A_Y0KSzmJG1_2(.dout(w_dff_A_dY5lbPeH2_2),.din(w_dff_A_Y0KSzmJG1_2),.clk(gclk));
	jdff dff_B_ocmLXuYB1_0(.din(n348),.dout(w_dff_B_ocmLXuYB1_0),.clk(gclk));
	jdff dff_B_QSNp8d8W0_0(.din(w_dff_B_ocmLXuYB1_0),.dout(w_dff_B_QSNp8d8W0_0),.clk(gclk));
	jdff dff_B_x1gLVjkK1_0(.din(w_dff_B_QSNp8d8W0_0),.dout(w_dff_B_x1gLVjkK1_0),.clk(gclk));
	jdff dff_B_8nRvfffo3_0(.din(w_dff_B_x1gLVjkK1_0),.dout(w_dff_B_8nRvfffo3_0),.clk(gclk));
	jdff dff_B_UgI77JXC7_0(.din(w_dff_B_8nRvfffo3_0),.dout(w_dff_B_UgI77JXC7_0),.clk(gclk));
	jdff dff_B_8vVYtivF3_0(.din(w_dff_B_UgI77JXC7_0),.dout(w_dff_B_8vVYtivF3_0),.clk(gclk));
	jdff dff_B_ZATPpVoE5_0(.din(w_dff_B_8vVYtivF3_0),.dout(w_dff_B_ZATPpVoE5_0),.clk(gclk));
	jdff dff_A_Hf4R2y4P9_1(.dout(w_n347_0[1]),.din(w_dff_A_Hf4R2y4P9_1),.clk(gclk));
	jdff dff_A_fnZaLzfw6_1(.dout(w_dff_A_Hf4R2y4P9_1),.din(w_dff_A_fnZaLzfw6_1),.clk(gclk));
	jdff dff_A_iAJ93bts7_1(.dout(w_dff_A_fnZaLzfw6_1),.din(w_dff_A_iAJ93bts7_1),.clk(gclk));
	jdff dff_A_izT8ZUpC3_1(.dout(w_dff_A_iAJ93bts7_1),.din(w_dff_A_izT8ZUpC3_1),.clk(gclk));
	jdff dff_A_wUV9aZlo1_1(.dout(w_dff_A_izT8ZUpC3_1),.din(w_dff_A_wUV9aZlo1_1),.clk(gclk));
	jdff dff_A_7x4rsCSo3_1(.dout(w_dff_A_wUV9aZlo1_1),.din(w_dff_A_7x4rsCSo3_1),.clk(gclk));
	jdff dff_A_3Y6MdOJP6_1(.dout(w_dff_A_7x4rsCSo3_1),.din(w_dff_A_3Y6MdOJP6_1),.clk(gclk));
	jdff dff_B_YP1ptw8m1_0(.din(n381),.dout(w_dff_B_YP1ptw8m1_0),.clk(gclk));
	jdff dff_B_qyAHTwhB0_0(.din(w_dff_B_YP1ptw8m1_0),.dout(w_dff_B_qyAHTwhB0_0),.clk(gclk));
	jdff dff_B_34uARqsn6_0(.din(w_dff_B_qyAHTwhB0_0),.dout(w_dff_B_34uARqsn6_0),.clk(gclk));
	jdff dff_B_vQMMS74M7_0(.din(w_dff_B_34uARqsn6_0),.dout(w_dff_B_vQMMS74M7_0),.clk(gclk));
	jdff dff_B_6429jJEN6_0(.din(w_dff_B_vQMMS74M7_0),.dout(w_dff_B_6429jJEN6_0),.clk(gclk));
	jdff dff_B_oC0b5SRv8_0(.din(w_dff_B_6429jJEN6_0),.dout(w_dff_B_oC0b5SRv8_0),.clk(gclk));
	jdff dff_B_hZWEU94y7_0(.din(w_dff_B_oC0b5SRv8_0),.dout(w_dff_B_hZWEU94y7_0),.clk(gclk));
	jdff dff_B_AfRRtiyr7_0(.din(w_dff_B_hZWEU94y7_0),.dout(w_dff_B_AfRRtiyr7_0),.clk(gclk));
	jdff dff_B_Fo1aHILk9_0(.din(w_dff_B_AfRRtiyr7_0),.dout(w_dff_B_Fo1aHILk9_0),.clk(gclk));
	jdff dff_B_Izf4783V0_0(.din(w_dff_B_Fo1aHILk9_0),.dout(w_dff_B_Izf4783V0_0),.clk(gclk));
	jdff dff_B_ym3pvic20_0(.din(n379),.dout(w_dff_B_ym3pvic20_0),.clk(gclk));
	jdff dff_B_MIHLAari6_0(.din(w_dff_B_ym3pvic20_0),.dout(w_dff_B_MIHLAari6_0),.clk(gclk));
	jdff dff_B_YtlP2FKE4_0(.din(n378),.dout(w_dff_B_YtlP2FKE4_0),.clk(gclk));
	jdff dff_B_Tcu6c5IJ4_0(.din(w_dff_B_YtlP2FKE4_0),.dout(w_dff_B_Tcu6c5IJ4_0),.clk(gclk));
	jdff dff_B_sgHWmJTp7_0(.din(w_dff_B_Tcu6c5IJ4_0),.dout(w_dff_B_sgHWmJTp7_0),.clk(gclk));
	jdff dff_B_jjcIAjEI9_0(.din(w_dff_B_sgHWmJTp7_0),.dout(w_dff_B_jjcIAjEI9_0),.clk(gclk));
	jdff dff_B_hgt6o9t34_0(.din(n375),.dout(w_dff_B_hgt6o9t34_0),.clk(gclk));
	jdff dff_B_MlJi8swA5_0(.din(w_dff_B_hgt6o9t34_0),.dout(w_dff_B_MlJi8swA5_0),.clk(gclk));
	jdff dff_B_3DYU1nwt0_0(.din(w_dff_B_MlJi8swA5_0),.dout(w_dff_B_3DYU1nwt0_0),.clk(gclk));
	jdff dff_B_utkHbiUL4_0(.din(w_dff_B_3DYU1nwt0_0),.dout(w_dff_B_utkHbiUL4_0),.clk(gclk));
	jdff dff_B_Wh4Yu1TF4_0(.din(w_dff_B_utkHbiUL4_0),.dout(w_dff_B_Wh4Yu1TF4_0),.clk(gclk));
	jdff dff_B_lQd04rdX2_0(.din(n368),.dout(w_dff_B_lQd04rdX2_0),.clk(gclk));
	jdff dff_B_T9QDIIpq3_0(.din(w_dff_B_lQd04rdX2_0),.dout(w_dff_B_T9QDIIpq3_0),.clk(gclk));
	jdff dff_B_sBvHmArP9_0(.din(w_dff_B_T9QDIIpq3_0),.dout(w_dff_B_sBvHmArP9_0),.clk(gclk));
	jdff dff_B_1TRPL6zQ8_0(.din(w_dff_B_sBvHmArP9_0),.dout(w_dff_B_1TRPL6zQ8_0),.clk(gclk));
	jdff dff_B_2dDd7thp5_0(.din(w_dff_B_1TRPL6zQ8_0),.dout(w_dff_B_2dDd7thp5_0),.clk(gclk));
	jdff dff_B_cN5Fl1bl3_0(.din(w_dff_B_2dDd7thp5_0),.dout(w_dff_B_cN5Fl1bl3_0),.clk(gclk));
	jdff dff_B_lNQigljw6_0(.din(w_dff_B_cN5Fl1bl3_0),.dout(w_dff_B_lNQigljw6_0),.clk(gclk));
	jdff dff_B_9qONROA47_0(.din(w_dff_B_lNQigljw6_0),.dout(w_dff_B_9qONROA47_0),.clk(gclk));
	jdff dff_B_PNoVvop11_0(.din(w_dff_B_9qONROA47_0),.dout(w_dff_B_PNoVvop11_0),.clk(gclk));
	jdff dff_A_GGqPTmaf8_1(.dout(w_n367_0[1]),.din(w_dff_A_GGqPTmaf8_1),.clk(gclk));
	jdff dff_A_qJlR1Via2_1(.dout(w_dff_A_GGqPTmaf8_1),.din(w_dff_A_qJlR1Via2_1),.clk(gclk));
	jdff dff_A_1c6f6JN29_1(.dout(w_dff_A_qJlR1Via2_1),.din(w_dff_A_1c6f6JN29_1),.clk(gclk));
	jdff dff_A_fYQhOLMb1_1(.dout(w_dff_A_1c6f6JN29_1),.din(w_dff_A_fYQhOLMb1_1),.clk(gclk));
	jdff dff_A_PuEJQdU62_1(.dout(w_dff_A_fYQhOLMb1_1),.din(w_dff_A_PuEJQdU62_1),.clk(gclk));
	jdff dff_A_glE6YjOI9_1(.dout(w_dff_A_PuEJQdU62_1),.din(w_dff_A_glE6YjOI9_1),.clk(gclk));
	jdff dff_A_DD5VzlQI2_1(.dout(w_dff_A_glE6YjOI9_1),.din(w_dff_A_DD5VzlQI2_1),.clk(gclk));
	jdff dff_A_yLKQHjhw5_1(.dout(w_dff_A_DD5VzlQI2_1),.din(w_dff_A_yLKQHjhw5_1),.clk(gclk));
	jdff dff_A_zguWoSTU8_1(.dout(w_dff_A_yLKQHjhw5_1),.din(w_dff_A_zguWoSTU8_1),.clk(gclk));
	jdff dff_B_Njars19K6_1(.din(n294),.dout(w_dff_B_Njars19K6_1),.clk(gclk));
	jdff dff_B_T1w9DNB23_1(.din(w_dff_B_Njars19K6_1),.dout(w_dff_B_T1w9DNB23_1),.clk(gclk));
	jdff dff_B_nBOiScYI3_1(.din(w_dff_B_T1w9DNB23_1),.dout(w_dff_B_nBOiScYI3_1),.clk(gclk));
	jdff dff_A_3NFqrWk85_1(.dout(w_G159gat_1[1]),.din(w_dff_A_3NFqrWk85_1),.clk(gclk));
	jdff dff_A_XJ75fKMM1_1(.dout(w_dff_A_3NFqrWk85_1),.din(w_dff_A_XJ75fKMM1_1),.clk(gclk));
	jdff dff_A_4sauANMr5_1(.dout(w_dff_A_XJ75fKMM1_1),.din(w_dff_A_4sauANMr5_1),.clk(gclk));
	jdff dff_A_5Rc1NTn82_1(.dout(w_dff_A_4sauANMr5_1),.din(w_dff_A_5Rc1NTn82_1),.clk(gclk));
	jdff dff_A_22EzaNRH2_1(.dout(w_dff_A_5Rc1NTn82_1),.din(w_dff_A_22EzaNRH2_1),.clk(gclk));
	jdff dff_A_YFVx8Hve1_1(.dout(w_dff_A_22EzaNRH2_1),.din(w_dff_A_YFVx8Hve1_1),.clk(gclk));
	jdff dff_A_3CXBDjGy9_1(.dout(w_dff_A_YFVx8Hve1_1),.din(w_dff_A_3CXBDjGy9_1),.clk(gclk));
	jdff dff_A_ONychntC1_2(.dout(w_G159gat_1[2]),.din(w_dff_A_ONychntC1_2),.clk(gclk));
	jdff dff_A_4GwYeHZU7_2(.dout(w_dff_A_ONychntC1_2),.din(w_dff_A_4GwYeHZU7_2),.clk(gclk));
	jdff dff_A_rZWI63BR4_2(.dout(w_dff_A_4GwYeHZU7_2),.din(w_dff_A_rZWI63BR4_2),.clk(gclk));
	jdff dff_A_rCHswxiA2_2(.dout(w_dff_A_rZWI63BR4_2),.din(w_dff_A_rCHswxiA2_2),.clk(gclk));
	jdff dff_A_4CYVFgmW9_2(.dout(w_dff_A_rCHswxiA2_2),.din(w_dff_A_4CYVFgmW9_2),.clk(gclk));
	jdff dff_A_1b3pr0Eu8_2(.dout(w_dff_A_4CYVFgmW9_2),.din(w_dff_A_1b3pr0Eu8_2),.clk(gclk));
	jdff dff_A_pFZYmTHO8_2(.dout(w_dff_A_1b3pr0Eu8_2),.din(w_dff_A_pFZYmTHO8_2),.clk(gclk));
	jdff dff_A_7j1cYmm35_2(.dout(w_G159gat_0[2]),.din(w_dff_A_7j1cYmm35_2),.clk(gclk));
	jdff dff_A_7QNwRjLL8_2(.dout(w_dff_A_7j1cYmm35_2),.din(w_dff_A_7QNwRjLL8_2),.clk(gclk));
	jdff dff_A_VALLlZDi7_2(.dout(w_dff_A_7QNwRjLL8_2),.din(w_dff_A_VALLlZDi7_2),.clk(gclk));
	jdff dff_A_Y7MJgL9w2_2(.dout(w_dff_A_VALLlZDi7_2),.din(w_dff_A_Y7MJgL9w2_2),.clk(gclk));
	jdff dff_B_fI6OMezF4_0(.din(n365),.dout(w_dff_B_fI6OMezF4_0),.clk(gclk));
	jdff dff_B_PUoCACqF5_0(.din(w_dff_B_fI6OMezF4_0),.dout(w_dff_B_PUoCACqF5_0),.clk(gclk));
	jdff dff_B_FCcmQtCQ5_0(.din(w_dff_B_PUoCACqF5_0),.dout(w_dff_B_FCcmQtCQ5_0),.clk(gclk));
	jdff dff_B_WjlhjVFz8_0(.din(w_dff_B_FCcmQtCQ5_0),.dout(w_dff_B_WjlhjVFz8_0),.clk(gclk));
	jdff dff_A_L73bfKqD5_1(.dout(w_n339_0[1]),.din(w_dff_A_L73bfKqD5_1),.clk(gclk));
	jdff dff_A_QRSBxjvm0_1(.dout(w_dff_A_L73bfKqD5_1),.din(w_dff_A_QRSBxjvm0_1),.clk(gclk));
	jdff dff_A_smHjJcy14_1(.dout(w_dff_A_QRSBxjvm0_1),.din(w_dff_A_smHjJcy14_1),.clk(gclk));
	jdff dff_A_AbClJDsC1_1(.dout(w_dff_A_smHjJcy14_1),.din(w_dff_A_AbClJDsC1_1),.clk(gclk));
	jdff dff_B_JLFDRsbE1_1(.din(n333),.dout(w_dff_B_JLFDRsbE1_1),.clk(gclk));
	jdff dff_B_TI3tV9FD4_1(.din(w_dff_B_JLFDRsbE1_1),.dout(w_dff_B_TI3tV9FD4_1),.clk(gclk));
	jdff dff_B_6W5xi0fm4_1(.din(w_dff_B_TI3tV9FD4_1),.dout(w_dff_B_6W5xi0fm4_1),.clk(gclk));
	jdff dff_B_mLJ7Ql8H6_0(.din(n363),.dout(w_dff_B_mLJ7Ql8H6_0),.clk(gclk));
	jdff dff_B_7URkGVGW8_0(.din(w_dff_B_mLJ7Ql8H6_0),.dout(w_dff_B_7URkGVGW8_0),.clk(gclk));
	jdff dff_B_EPuOvwon3_0(.din(w_dff_B_7URkGVGW8_0),.dout(w_dff_B_EPuOvwon3_0),.clk(gclk));
	jdff dff_B_LpuWcMhc0_0(.din(w_dff_B_EPuOvwon3_0),.dout(w_dff_B_LpuWcMhc0_0),.clk(gclk));
	jdff dff_A_d5WapaAd8_1(.dout(w_n331_0[1]),.din(w_dff_A_d5WapaAd8_1),.clk(gclk));
	jdff dff_A_j39aCgnn3_1(.dout(w_dff_A_d5WapaAd8_1),.din(w_dff_A_j39aCgnn3_1),.clk(gclk));
	jdff dff_A_Aga2VbG81_1(.dout(w_dff_A_j39aCgnn3_1),.din(w_dff_A_Aga2VbG81_1),.clk(gclk));
	jdff dff_A_W22bFRvE6_1(.dout(w_dff_A_Aga2VbG81_1),.din(w_dff_A_W22bFRvE6_1),.clk(gclk));
	jdff dff_B_OJKZr1Pa1_1(.din(n306),.dout(w_dff_B_OJKZr1Pa1_1),.clk(gclk));
	jdff dff_B_VE2PbU0n4_1(.din(w_dff_B_OJKZr1Pa1_1),.dout(w_dff_B_VE2PbU0n4_1),.clk(gclk));
	jdff dff_B_PdEw4Pai8_1(.din(w_dff_B_VE2PbU0n4_1),.dout(w_dff_B_PdEw4Pai8_1),.clk(gclk));
	jdff dff_B_YbtlO2aU0_1(.din(w_dff_B_PdEw4Pai8_1),.dout(w_dff_B_YbtlO2aU0_1),.clk(gclk));
	jdff dff_B_U9yoAtHN1_1(.din(w_dff_B_YbtlO2aU0_1),.dout(w_dff_B_U9yoAtHN1_1),.clk(gclk));
	jdff dff_B_UsVqLjAM8_1(.din(w_dff_B_U9yoAtHN1_1),.dout(w_dff_B_UsVqLjAM8_1),.clk(gclk));
	jdff dff_B_pRJznE1q4_1(.din(w_dff_B_UsVqLjAM8_1),.dout(w_dff_B_pRJznE1q4_1),.clk(gclk));
	jdff dff_B_CO0TEYyV5_0(.din(n403),.dout(w_dff_B_CO0TEYyV5_0),.clk(gclk));
	jdff dff_B_RfywZe636_0(.din(w_dff_B_CO0TEYyV5_0),.dout(w_dff_B_RfywZe636_0),.clk(gclk));
	jdff dff_B_7q6IeY6F4_0(.din(w_dff_B_RfywZe636_0),.dout(w_dff_B_7q6IeY6F4_0),.clk(gclk));
	jdff dff_B_R2TlDJIS9_0(.din(w_dff_B_7q6IeY6F4_0),.dout(w_dff_B_R2TlDJIS9_0),.clk(gclk));
	jdff dff_B_V8mtbQ7e9_0(.din(w_dff_B_R2TlDJIS9_0),.dout(w_dff_B_V8mtbQ7e9_0),.clk(gclk));
	jdff dff_B_KiN71b3D9_0(.din(w_dff_B_V8mtbQ7e9_0),.dout(w_dff_B_KiN71b3D9_0),.clk(gclk));
	jdff dff_B_Feks7tyM3_0(.din(w_dff_B_KiN71b3D9_0),.dout(w_dff_B_Feks7tyM3_0),.clk(gclk));
	jdff dff_B_pD7DtAH65_0(.din(w_dff_B_Feks7tyM3_0),.dout(w_dff_B_pD7DtAH65_0),.clk(gclk));
	jdff dff_B_PxDM8Pdk2_0(.din(w_dff_B_pD7DtAH65_0),.dout(w_dff_B_PxDM8Pdk2_0),.clk(gclk));
	jdff dff_B_knFNQfaJ1_0(.din(w_dff_B_PxDM8Pdk2_0),.dout(w_dff_B_knFNQfaJ1_0),.clk(gclk));
	jdff dff_B_TkBwFMYm3_0(.din(n401),.dout(w_dff_B_TkBwFMYm3_0),.clk(gclk));
	jdff dff_B_2spQn6sk2_0(.din(w_dff_B_TkBwFMYm3_0),.dout(w_dff_B_2spQn6sk2_0),.clk(gclk));
	jdff dff_B_mKHVLYLl6_0(.din(n400),.dout(w_dff_B_mKHVLYLl6_0),.clk(gclk));
	jdff dff_B_r4tmjpNV0_0(.din(w_dff_B_mKHVLYLl6_0),.dout(w_dff_B_r4tmjpNV0_0),.clk(gclk));
	jdff dff_B_MBICdgy26_0(.din(w_dff_B_r4tmjpNV0_0),.dout(w_dff_B_MBICdgy26_0),.clk(gclk));
	jdff dff_B_qyXVzmYJ7_0(.din(w_dff_B_MBICdgy26_0),.dout(w_dff_B_qyXVzmYJ7_0),.clk(gclk));
	jdff dff_A_hA9yRRx98_1(.dout(w_G91gat_0[1]),.din(w_dff_A_hA9yRRx98_1),.clk(gclk));
	jdff dff_A_EKF1ZGSF3_1(.dout(w_dff_A_hA9yRRx98_1),.din(w_dff_A_EKF1ZGSF3_1),.clk(gclk));
	jdff dff_A_hBLY9SOv4_1(.dout(w_dff_A_EKF1ZGSF3_1),.din(w_dff_A_hBLY9SOv4_1),.clk(gclk));
	jdff dff_A_pBohs5H37_1(.dout(w_dff_A_hBLY9SOv4_1),.din(w_dff_A_pBohs5H37_1),.clk(gclk));
	jdff dff_A_6LWhfFPr7_1(.dout(w_dff_A_pBohs5H37_1),.din(w_dff_A_6LWhfFPr7_1),.clk(gclk));
	jdff dff_B_cB1AxH6V7_0(.din(n397),.dout(w_dff_B_cB1AxH6V7_0),.clk(gclk));
	jdff dff_B_KKaxXAic3_0(.din(w_dff_B_cB1AxH6V7_0),.dout(w_dff_B_KKaxXAic3_0),.clk(gclk));
	jdff dff_B_CH4j4C5Y7_0(.din(w_dff_B_KKaxXAic3_0),.dout(w_dff_B_CH4j4C5Y7_0),.clk(gclk));
	jdff dff_B_ZAcBpBG22_0(.din(w_dff_B_CH4j4C5Y7_0),.dout(w_dff_B_ZAcBpBG22_0),.clk(gclk));
	jdff dff_B_GJ3Zrlbj5_0(.din(w_dff_B_ZAcBpBG22_0),.dout(w_dff_B_GJ3Zrlbj5_0),.clk(gclk));
	jdff dff_B_t4CSkoIp3_1(.din(n384),.dout(w_dff_B_t4CSkoIp3_1),.clk(gclk));
	jdff dff_B_ow44jL611_1(.din(w_dff_B_t4CSkoIp3_1),.dout(w_dff_B_ow44jL611_1),.clk(gclk));
	jdff dff_B_N35O9IcH8_1(.din(w_dff_B_ow44jL611_1),.dout(w_dff_B_N35O9IcH8_1),.clk(gclk));
	jdff dff_B_U8Jo871b9_1(.din(w_dff_B_N35O9IcH8_1),.dout(w_dff_B_U8Jo871b9_1),.clk(gclk));
	jdff dff_B_efg2qdYU1_1(.din(w_dff_B_U8Jo871b9_1),.dout(w_dff_B_efg2qdYU1_1),.clk(gclk));
	jdff dff_B_emH93ejM9_1(.din(w_dff_B_efg2qdYU1_1),.dout(w_dff_B_emH93ejM9_1),.clk(gclk));
	jdff dff_B_mrW5kCZ85_1(.din(w_dff_B_emH93ejM9_1),.dout(w_dff_B_mrW5kCZ85_1),.clk(gclk));
	jdff dff_B_HQAup70o0_1(.din(w_dff_B_mrW5kCZ85_1),.dout(w_dff_B_HQAup70o0_1),.clk(gclk));
	jdff dff_B_OelSTeiU1_1(.din(w_dff_B_HQAup70o0_1),.dout(w_dff_B_OelSTeiU1_1),.clk(gclk));
	jdff dff_B_mZuN47YQ3_1(.din(n385),.dout(w_dff_B_mZuN47YQ3_1),.clk(gclk));
	jdff dff_B_Jr5ZHMyQ0_1(.din(w_dff_B_mZuN47YQ3_1),.dout(w_dff_B_Jr5ZHMyQ0_1),.clk(gclk));
	jdff dff_B_kn2ms3Rz5_1(.din(w_dff_B_Jr5ZHMyQ0_1),.dout(w_dff_B_kn2ms3Rz5_1),.clk(gclk));
	jdff dff_B_q4xEbWFW2_1(.din(w_dff_B_kn2ms3Rz5_1),.dout(w_dff_B_q4xEbWFW2_1),.clk(gclk));
	jdff dff_B_QNGxCLSY9_1(.din(w_dff_B_q4xEbWFW2_1),.dout(w_dff_B_QNGxCLSY9_1),.clk(gclk));
	jdff dff_B_fkPCQbba7_1(.din(w_dff_B_QNGxCLSY9_1),.dout(w_dff_B_fkPCQbba7_1),.clk(gclk));
	jdff dff_B_AlOKLYwV3_0(.din(n386),.dout(w_dff_B_AlOKLYwV3_0),.clk(gclk));
	jdff dff_B_FvY63EkL9_0(.din(w_dff_B_AlOKLYwV3_0),.dout(w_dff_B_FvY63EkL9_0),.clk(gclk));
	jdff dff_B_fNYjGCB03_0(.din(w_dff_B_FvY63EkL9_0),.dout(w_dff_B_fNYjGCB03_0),.clk(gclk));
	jdff dff_B_f84puu9g0_0(.din(w_dff_B_fNYjGCB03_0),.dout(w_dff_B_f84puu9g0_0),.clk(gclk));
	jdff dff_B_4z0SVa6o3_0(.din(w_dff_B_f84puu9g0_0),.dout(w_dff_B_4z0SVa6o3_0),.clk(gclk));
	jdff dff_B_3XQtlWSc7_0(.din(w_dff_B_4z0SVa6o3_0),.dout(w_dff_B_3XQtlWSc7_0),.clk(gclk));
	jdff dff_A_D5s9Hsp36_0(.dout(w_n330_0[0]),.din(w_dff_A_D5s9Hsp36_0),.clk(gclk));
	jdff dff_A_3VFNgtBl1_0(.dout(w_dff_A_D5s9Hsp36_0),.din(w_dff_A_3VFNgtBl1_0),.clk(gclk));
	jdff dff_A_eiCg0iHe0_0(.dout(w_dff_A_3VFNgtBl1_0),.din(w_dff_A_eiCg0iHe0_0),.clk(gclk));
	jdff dff_A_YwyFruk58_0(.dout(w_dff_A_eiCg0iHe0_0),.din(w_dff_A_YwyFruk58_0),.clk(gclk));
	jdff dff_A_J8mq48JQ0_0(.dout(w_dff_A_YwyFruk58_0),.din(w_dff_A_J8mq48JQ0_0),.clk(gclk));
	jdff dff_A_dfDj8RWL9_0(.dout(w_dff_A_J8mq48JQ0_0),.din(w_dff_A_dfDj8RWL9_0),.clk(gclk));
	jdff dff_A_KbcVS7sh7_2(.dout(w_n330_0[2]),.din(w_dff_A_KbcVS7sh7_2),.clk(gclk));
	jdff dff_A_KnGvYnNg0_0(.dout(w_n337_0[0]),.din(w_dff_A_KnGvYnNg0_0),.clk(gclk));
	jdff dff_A_rIpQowp34_0(.dout(w_dff_A_KnGvYnNg0_0),.din(w_dff_A_rIpQowp34_0),.clk(gclk));
	jdff dff_A_qJKfoSUw4_0(.dout(w_dff_A_rIpQowp34_0),.din(w_dff_A_qJKfoSUw4_0),.clk(gclk));
	jdff dff_A_bPA3mF5m3_0(.dout(w_dff_A_qJKfoSUw4_0),.din(w_dff_A_bPA3mF5m3_0),.clk(gclk));
	jdff dff_A_90RkIKWw4_0(.dout(w_dff_A_bPA3mF5m3_0),.din(w_dff_A_90RkIKWw4_0),.clk(gclk));
	jdff dff_A_wS7nXe1t7_0(.dout(w_dff_A_90RkIKWw4_0),.din(w_dff_A_wS7nXe1t7_0),.clk(gclk));
	jdff dff_B_lkdbdiPE2_1(.din(n334),.dout(w_dff_B_lkdbdiPE2_1),.clk(gclk));
	jdff dff_A_Ko2xzVei3_0(.dout(w_G171gat_2[0]),.din(w_dff_A_Ko2xzVei3_0),.clk(gclk));
	jdff dff_A_wuiXzE2p2_0(.dout(w_dff_A_Ko2xzVei3_0),.din(w_dff_A_wuiXzE2p2_0),.clk(gclk));
	jdff dff_A_5xkH4MHd4_0(.dout(w_dff_A_wuiXzE2p2_0),.din(w_dff_A_5xkH4MHd4_0),.clk(gclk));
	jdff dff_A_oLAu9PgN6_0(.dout(w_dff_A_5xkH4MHd4_0),.din(w_dff_A_oLAu9PgN6_0),.clk(gclk));
	jdff dff_A_DmMZkXHQ6_0(.dout(w_dff_A_oLAu9PgN6_0),.din(w_dff_A_DmMZkXHQ6_0),.clk(gclk));
	jdff dff_A_UoymzHYZ3_0(.dout(w_dff_A_DmMZkXHQ6_0),.din(w_dff_A_UoymzHYZ3_0),.clk(gclk));
	jdff dff_A_KPkjkTHf0_0(.dout(w_dff_A_UoymzHYZ3_0),.din(w_dff_A_KPkjkTHf0_0),.clk(gclk));
	jdff dff_A_iKnk4anM6_1(.dout(w_n383_0[1]),.din(w_dff_A_iKnk4anM6_1),.clk(gclk));
	jdff dff_A_ddbxkrov7_1(.dout(w_dff_A_iKnk4anM6_1),.din(w_dff_A_ddbxkrov7_1),.clk(gclk));
	jdff dff_A_Y1Bdosnl9_1(.dout(w_dff_A_ddbxkrov7_1),.din(w_dff_A_Y1Bdosnl9_1),.clk(gclk));
	jdff dff_A_diCDEsHX2_1(.dout(w_dff_A_Y1Bdosnl9_1),.din(w_dff_A_diCDEsHX2_1),.clk(gclk));
	jdff dff_A_RVw0n8sK9_1(.dout(w_dff_A_diCDEsHX2_1),.din(w_dff_A_RVw0n8sK9_1),.clk(gclk));
	jdff dff_A_pndzv8ct0_1(.dout(w_dff_A_RVw0n8sK9_1),.din(w_dff_A_pndzv8ct0_1),.clk(gclk));
	jdff dff_A_yMQ6iL6S3_1(.dout(w_dff_A_pndzv8ct0_1),.din(w_dff_A_yMQ6iL6S3_1),.clk(gclk));
	jdff dff_A_alIZJUzz0_1(.dout(w_dff_A_yMQ6iL6S3_1),.din(w_dff_A_alIZJUzz0_1),.clk(gclk));
	jdff dff_A_UJ7N9NOf9_1(.dout(w_dff_A_alIZJUzz0_1),.din(w_dff_A_UJ7N9NOf9_1),.clk(gclk));
	jdff dff_B_5CABIsTw2_0(.din(n309),.dout(w_dff_B_5CABIsTw2_0),.clk(gclk));
	jdff dff_B_TjBTKXoi7_0(.din(w_dff_B_5CABIsTw2_0),.dout(w_dff_B_TjBTKXoi7_0),.clk(gclk));
	jdff dff_B_i5cAmkLc7_0(.din(w_dff_B_TjBTKXoi7_0),.dout(w_dff_B_i5cAmkLc7_0),.clk(gclk));
	jdff dff_A_jvc0pF3Z5_1(.dout(w_G165gat_1[1]),.din(w_dff_A_jvc0pF3Z5_1),.clk(gclk));
	jdff dff_A_eJxtZOeL6_1(.dout(w_dff_A_jvc0pF3Z5_1),.din(w_dff_A_eJxtZOeL6_1),.clk(gclk));
	jdff dff_A_j6aI7Icb3_1(.dout(w_dff_A_eJxtZOeL6_1),.din(w_dff_A_j6aI7Icb3_1),.clk(gclk));
	jdff dff_A_lTYqFZCO3_1(.dout(w_dff_A_j6aI7Icb3_1),.din(w_dff_A_lTYqFZCO3_1),.clk(gclk));
	jdff dff_A_TJCZ1xdI6_1(.dout(w_dff_A_lTYqFZCO3_1),.din(w_dff_A_TJCZ1xdI6_1),.clk(gclk));
	jdff dff_A_WnLAxBC29_1(.dout(w_dff_A_TJCZ1xdI6_1),.din(w_dff_A_WnLAxBC29_1),.clk(gclk));
	jdff dff_A_jc7HTzSh1_1(.dout(w_dff_A_WnLAxBC29_1),.din(w_dff_A_jc7HTzSh1_1),.clk(gclk));
	jdff dff_A_bsCysOS74_2(.dout(w_G165gat_1[2]),.din(w_dff_A_bsCysOS74_2),.clk(gclk));
	jdff dff_A_vFormJ3P0_2(.dout(w_dff_A_bsCysOS74_2),.din(w_dff_A_vFormJ3P0_2),.clk(gclk));
	jdff dff_A_jxuKexFD5_2(.dout(w_dff_A_vFormJ3P0_2),.din(w_dff_A_jxuKexFD5_2),.clk(gclk));
	jdff dff_A_pIJI1wR47_2(.dout(w_dff_A_jxuKexFD5_2),.din(w_dff_A_pIJI1wR47_2),.clk(gclk));
	jdff dff_A_sbFtc1u37_2(.dout(w_dff_A_pIJI1wR47_2),.din(w_dff_A_sbFtc1u37_2),.clk(gclk));
	jdff dff_A_VaX0XcJM4_2(.dout(w_dff_A_sbFtc1u37_2),.din(w_dff_A_VaX0XcJM4_2),.clk(gclk));
	jdff dff_A_5KNPP9EU7_2(.dout(w_dff_A_VaX0XcJM4_2),.din(w_dff_A_5KNPP9EU7_2),.clk(gclk));
	jdff dff_A_eterAJUo3_2(.dout(w_G165gat_0[2]),.din(w_dff_A_eterAJUo3_2),.clk(gclk));
	jdff dff_A_RYypYTir9_2(.dout(w_dff_A_eterAJUo3_2),.din(w_dff_A_RYypYTir9_2),.clk(gclk));
	jdff dff_A_7LdjYk5T4_2(.dout(w_dff_A_RYypYTir9_2),.din(w_dff_A_7LdjYk5T4_2),.clk(gclk));
	jdff dff_A_8XpGyw5C6_2(.dout(w_dff_A_7LdjYk5T4_2),.din(w_dff_A_8XpGyw5C6_2),.clk(gclk));
	jdff dff_B_zeyF7S7C6_0(.din(n425),.dout(w_dff_B_zeyF7S7C6_0),.clk(gclk));
	jdff dff_B_i6oBulh41_0(.din(w_dff_B_zeyF7S7C6_0),.dout(w_dff_B_i6oBulh41_0),.clk(gclk));
	jdff dff_B_EgtbQ1og3_0(.din(w_dff_B_i6oBulh41_0),.dout(w_dff_B_EgtbQ1og3_0),.clk(gclk));
	jdff dff_B_uGwKqtyq4_0(.din(w_dff_B_EgtbQ1og3_0),.dout(w_dff_B_uGwKqtyq4_0),.clk(gclk));
	jdff dff_B_ssY13juN7_0(.din(w_dff_B_uGwKqtyq4_0),.dout(w_dff_B_ssY13juN7_0),.clk(gclk));
	jdff dff_B_3ZBUr4P26_0(.din(w_dff_B_ssY13juN7_0),.dout(w_dff_B_3ZBUr4P26_0),.clk(gclk));
	jdff dff_B_pMpnmSFT7_0(.din(w_dff_B_3ZBUr4P26_0),.dout(w_dff_B_pMpnmSFT7_0),.clk(gclk));
	jdff dff_B_qMGeSdpT8_0(.din(w_dff_B_pMpnmSFT7_0),.dout(w_dff_B_qMGeSdpT8_0),.clk(gclk));
	jdff dff_B_xXJGaZgs1_0(.din(w_dff_B_qMGeSdpT8_0),.dout(w_dff_B_xXJGaZgs1_0),.clk(gclk));
	jdff dff_B_bBEt4ZWG5_0(.din(w_dff_B_xXJGaZgs1_0),.dout(w_dff_B_bBEt4ZWG5_0),.clk(gclk));
	jdff dff_B_cYhKNdA75_0(.din(n423),.dout(w_dff_B_cYhKNdA75_0),.clk(gclk));
	jdff dff_B_nBQKbeDD7_0(.din(w_dff_B_cYhKNdA75_0),.dout(w_dff_B_nBQKbeDD7_0),.clk(gclk));
	jdff dff_B_LovpfXDU5_0(.din(n422),.dout(w_dff_B_LovpfXDU5_0),.clk(gclk));
	jdff dff_B_ANnB8LUY2_0(.din(w_dff_B_LovpfXDU5_0),.dout(w_dff_B_ANnB8LUY2_0),.clk(gclk));
	jdff dff_B_z0Aue9fS2_0(.din(w_dff_B_ANnB8LUY2_0),.dout(w_dff_B_z0Aue9fS2_0),.clk(gclk));
	jdff dff_B_Pv1yspMa9_0(.din(w_dff_B_z0Aue9fS2_0),.dout(w_dff_B_Pv1yspMa9_0),.clk(gclk));
	jdff dff_A_it6uYGN15_1(.dout(w_G96gat_0[1]),.din(w_dff_A_it6uYGN15_1),.clk(gclk));
	jdff dff_A_N6o8wclS5_1(.dout(w_dff_A_it6uYGN15_1),.din(w_dff_A_N6o8wclS5_1),.clk(gclk));
	jdff dff_A_F2bI8AQq9_1(.dout(w_dff_A_N6o8wclS5_1),.din(w_dff_A_F2bI8AQq9_1),.clk(gclk));
	jdff dff_A_iKwxcC1S7_1(.dout(w_dff_A_F2bI8AQq9_1),.din(w_dff_A_iKwxcC1S7_1),.clk(gclk));
	jdff dff_A_98YQrYo79_1(.dout(w_dff_A_iKwxcC1S7_1),.din(w_dff_A_98YQrYo79_1),.clk(gclk));
	jdff dff_B_vTI34gNP8_1(.din(G73gat),.dout(w_dff_B_vTI34gNP8_1),.clk(gclk));
	jdff dff_A_LxxNHobh5_0(.dout(w_n121_0[0]),.din(w_dff_A_LxxNHobh5_0),.clk(gclk));
	jdff dff_A_shD5mLGa3_0(.dout(w_n118_0[0]),.din(w_dff_A_shD5mLGa3_0),.clk(gclk));
	jdff dff_B_CrHvogc18_0(.din(n419),.dout(w_dff_B_CrHvogc18_0),.clk(gclk));
	jdff dff_B_k7j50dZ35_0(.din(w_dff_B_CrHvogc18_0),.dout(w_dff_B_k7j50dZ35_0),.clk(gclk));
	jdff dff_B_lzpiCVSF1_0(.din(w_dff_B_k7j50dZ35_0),.dout(w_dff_B_lzpiCVSF1_0),.clk(gclk));
	jdff dff_B_RckJwQxV6_0(.din(w_dff_B_lzpiCVSF1_0),.dout(w_dff_B_RckJwQxV6_0),.clk(gclk));
	jdff dff_B_Gm0kNzhg3_0(.din(w_dff_B_RckJwQxV6_0),.dout(w_dff_B_Gm0kNzhg3_0),.clk(gclk));
	jdff dff_B_0gjBhWBg7_3(.din(G246gat),.dout(w_dff_B_0gjBhWBg7_3),.clk(gclk));
	jdff dff_A_JhAco3gd1_2(.dout(w_G228gat_0[2]),.din(w_dff_A_JhAco3gd1_2),.clk(gclk));
	jdff dff_B_yH1b8k1E3_3(.din(G228gat),.dout(w_dff_B_yH1b8k1E3_3),.clk(gclk));
	jdff dff_B_ZB59Gv4L7_3(.din(w_dff_B_yH1b8k1E3_3),.dout(w_dff_B_ZB59Gv4L7_3),.clk(gclk));
	jdff dff_B_7sgX5yrC5_3(.din(w_dff_B_ZB59Gv4L7_3),.dout(w_dff_B_7sgX5yrC5_3),.clk(gclk));
	jdff dff_B_OdRa28TU4_3(.din(w_dff_B_7sgX5yrC5_3),.dout(w_dff_B_OdRa28TU4_3),.clk(gclk));
	jdff dff_B_Wy3Gey7V3_3(.din(w_dff_B_OdRa28TU4_3),.dout(w_dff_B_Wy3Gey7V3_3),.clk(gclk));
	jdff dff_B_T8GuwOpR6_3(.din(w_dff_B_Wy3Gey7V3_3),.dout(w_dff_B_T8GuwOpR6_3),.clk(gclk));
	jdff dff_B_MSA3xcpb2_3(.din(w_dff_B_T8GuwOpR6_3),.dout(w_dff_B_MSA3xcpb2_3),.clk(gclk));
	jdff dff_B_cunaExpD1_3(.din(w_dff_B_MSA3xcpb2_3),.dout(w_dff_B_cunaExpD1_3),.clk(gclk));
	jdff dff_A_FWaJm0wq7_0(.dout(w_G219gat_0[0]),.din(w_dff_A_FWaJm0wq7_0),.clk(gclk));
	jdff dff_A_s3hp9UnE5_0(.dout(w_dff_A_FWaJm0wq7_0),.din(w_dff_A_s3hp9UnE5_0),.clk(gclk));
	jdff dff_A_RcxMbyay4_0(.dout(w_dff_A_s3hp9UnE5_0),.din(w_dff_A_RcxMbyay4_0),.clk(gclk));
	jdff dff_A_XopyLnzA5_0(.dout(w_dff_A_RcxMbyay4_0),.din(w_dff_A_XopyLnzA5_0),.clk(gclk));
	jdff dff_A_yvWTABtl4_0(.dout(w_dff_A_XopyLnzA5_0),.din(w_dff_A_yvWTABtl4_0),.clk(gclk));
	jdff dff_A_ViQqoSan2_0(.dout(w_dff_A_yvWTABtl4_0),.din(w_dff_A_ViQqoSan2_0),.clk(gclk));
	jdff dff_A_dL1MpdZe6_0(.dout(w_dff_A_ViQqoSan2_0),.din(w_dff_A_dL1MpdZe6_0),.clk(gclk));
	jdff dff_A_2WeA3owF7_0(.dout(w_dff_A_dL1MpdZe6_0),.din(w_dff_A_2WeA3owF7_0),.clk(gclk));
	jdff dff_A_WIADCNa01_1(.dout(w_G219gat_0[1]),.din(w_dff_A_WIADCNa01_1),.clk(gclk));
	jdff dff_A_j2mV2HVv6_1(.dout(w_dff_A_WIADCNa01_1),.din(w_dff_A_j2mV2HVv6_1),.clk(gclk));
	jdff dff_B_LECh1TG46_3(.din(G219gat),.dout(w_dff_B_LECh1TG46_3),.clk(gclk));
	jdff dff_B_k2ACAfl64_3(.din(w_dff_B_LECh1TG46_3),.dout(w_dff_B_k2ACAfl64_3),.clk(gclk));
	jdff dff_B_QAiyhTQn6_3(.din(w_dff_B_k2ACAfl64_3),.dout(w_dff_B_QAiyhTQn6_3),.clk(gclk));
	jdff dff_B_hTK7h19Q7_3(.din(w_dff_B_QAiyhTQn6_3),.dout(w_dff_B_hTK7h19Q7_3),.clk(gclk));
	jdff dff_B_Wrja4ard4_3(.din(w_dff_B_hTK7h19Q7_3),.dout(w_dff_B_Wrja4ard4_3),.clk(gclk));
	jdff dff_B_Zb8Mnr6N1_3(.din(w_dff_B_Wrja4ard4_3),.dout(w_dff_B_Zb8Mnr6N1_3),.clk(gclk));
	jdff dff_B_JABA05kb4_3(.din(w_dff_B_Zb8Mnr6N1_3),.dout(w_dff_B_JABA05kb4_3),.clk(gclk));
	jdff dff_B_js1SSsc40_3(.din(w_dff_B_JABA05kb4_3),.dout(w_dff_B_js1SSsc40_3),.clk(gclk));
	jdff dff_B_iTMyeUSy8_3(.din(w_dff_B_js1SSsc40_3),.dout(w_dff_B_iTMyeUSy8_3),.clk(gclk));
	jdff dff_B_ZL8ZAyZh2_3(.din(w_dff_B_iTMyeUSy8_3),.dout(w_dff_B_ZL8ZAyZh2_3),.clk(gclk));
	jdff dff_B_NiV2AKPp7_1(.din(n406),.dout(w_dff_B_NiV2AKPp7_1),.clk(gclk));
	jdff dff_B_90CIGYAP8_1(.din(w_dff_B_NiV2AKPp7_1),.dout(w_dff_B_90CIGYAP8_1),.clk(gclk));
	jdff dff_B_O7GIOyoc4_1(.din(w_dff_B_90CIGYAP8_1),.dout(w_dff_B_O7GIOyoc4_1),.clk(gclk));
	jdff dff_B_MQ5HIeHj0_1(.din(w_dff_B_O7GIOyoc4_1),.dout(w_dff_B_MQ5HIeHj0_1),.clk(gclk));
	jdff dff_B_ligpKIir9_1(.din(w_dff_B_MQ5HIeHj0_1),.dout(w_dff_B_ligpKIir9_1),.clk(gclk));
	jdff dff_B_zy5x0kiP4_1(.din(w_dff_B_ligpKIir9_1),.dout(w_dff_B_zy5x0kiP4_1),.clk(gclk));
	jdff dff_B_VpozsdDg7_1(.din(w_dff_B_zy5x0kiP4_1),.dout(w_dff_B_VpozsdDg7_1),.clk(gclk));
	jdff dff_B_2esykH8h4_1(.din(w_dff_B_VpozsdDg7_1),.dout(w_dff_B_2esykH8h4_1),.clk(gclk));
	jdff dff_B_NLszNRtg2_1(.din(w_dff_B_2esykH8h4_1),.dout(w_dff_B_NLszNRtg2_1),.clk(gclk));
	jdff dff_B_lYounoyC7_1(.din(n407),.dout(w_dff_B_lYounoyC7_1),.clk(gclk));
	jdff dff_B_fRQc0Ubi5_1(.din(w_dff_B_lYounoyC7_1),.dout(w_dff_B_fRQc0Ubi5_1),.clk(gclk));
	jdff dff_B_PWsRhbmR1_1(.din(w_dff_B_fRQc0Ubi5_1),.dout(w_dff_B_PWsRhbmR1_1),.clk(gclk));
	jdff dff_B_HVkZ9dnD0_1(.din(w_dff_B_PWsRhbmR1_1),.dout(w_dff_B_HVkZ9dnD0_1),.clk(gclk));
	jdff dff_B_kHP8xzmV3_1(.din(w_dff_B_HVkZ9dnD0_1),.dout(w_dff_B_kHP8xzmV3_1),.clk(gclk));
	jdff dff_B_0q7Y0Ifp9_1(.din(w_dff_B_kHP8xzmV3_1),.dout(w_dff_B_0q7Y0Ifp9_1),.clk(gclk));
	jdff dff_B_dvgKbKCL6_1(.din(w_dff_B_0q7Y0Ifp9_1),.dout(w_dff_B_dvgKbKCL6_1),.clk(gclk));
	jdff dff_B_QyXeecTJ0_1(.din(w_dff_B_dvgKbKCL6_1),.dout(w_dff_B_QyXeecTJ0_1),.clk(gclk));
	jdff dff_B_VLbt0aoS7_0(.din(n408),.dout(w_dff_B_VLbt0aoS7_0),.clk(gclk));
	jdff dff_B_tkk7Pp4Y7_0(.din(w_dff_B_VLbt0aoS7_0),.dout(w_dff_B_tkk7Pp4Y7_0),.clk(gclk));
	jdff dff_B_Fw2zGQ9u2_0(.din(w_dff_B_tkk7Pp4Y7_0),.dout(w_dff_B_Fw2zGQ9u2_0),.clk(gclk));
	jdff dff_B_u8LhLyL08_0(.din(w_dff_B_Fw2zGQ9u2_0),.dout(w_dff_B_u8LhLyL08_0),.clk(gclk));
	jdff dff_B_3dK4KEEy6_0(.din(w_dff_B_u8LhLyL08_0),.dout(w_dff_B_3dK4KEEy6_0),.clk(gclk));
	jdff dff_B_gorGpyFJ5_0(.din(w_dff_B_3dK4KEEy6_0),.dout(w_dff_B_gorGpyFJ5_0),.clk(gclk));
	jdff dff_B_L0320AkD2_0(.din(w_dff_B_gorGpyFJ5_0),.dout(w_dff_B_L0320AkD2_0),.clk(gclk));
	jdff dff_A_0lyqxPsZ5_0(.dout(w_n329_0[0]),.din(w_dff_A_0lyqxPsZ5_0),.clk(gclk));
	jdff dff_A_WzPbRMYu6_0(.dout(w_dff_A_0lyqxPsZ5_0),.din(w_dff_A_WzPbRMYu6_0),.clk(gclk));
	jdff dff_A_tlvt9k2R0_0(.dout(w_dff_A_WzPbRMYu6_0),.din(w_dff_A_tlvt9k2R0_0),.clk(gclk));
	jdff dff_A_s3zgy9cj0_0(.dout(w_dff_A_tlvt9k2R0_0),.din(w_dff_A_s3zgy9cj0_0),.clk(gclk));
	jdff dff_A_OCJEHcr90_0(.dout(w_dff_A_s3zgy9cj0_0),.din(w_dff_A_OCJEHcr90_0),.clk(gclk));
	jdff dff_A_burd5mjC4_0(.dout(w_dff_A_OCJEHcr90_0),.din(w_dff_A_burd5mjC4_0),.clk(gclk));
	jdff dff_A_kScFJcsb4_0(.dout(w_dff_A_burd5mjC4_0),.din(w_dff_A_kScFJcsb4_0),.clk(gclk));
	jdff dff_A_WK3aLGhH9_0(.dout(w_G177gat_2[0]),.din(w_dff_A_WK3aLGhH9_0),.clk(gclk));
	jdff dff_A_jw1L4KQf4_0(.dout(w_dff_A_WK3aLGhH9_0),.din(w_dff_A_jw1L4KQf4_0),.clk(gclk));
	jdff dff_A_gF8O0kOx7_0(.dout(w_dff_A_jw1L4KQf4_0),.din(w_dff_A_gF8O0kOx7_0),.clk(gclk));
	jdff dff_A_h3AlJXLC9_0(.dout(w_dff_A_gF8O0kOx7_0),.din(w_dff_A_h3AlJXLC9_0),.clk(gclk));
	jdff dff_A_pX56OMCk2_0(.dout(w_dff_A_h3AlJXLC9_0),.din(w_dff_A_pX56OMCk2_0),.clk(gclk));
	jdff dff_A_ZXyQHwlc3_0(.dout(w_dff_A_pX56OMCk2_0),.din(w_dff_A_ZXyQHwlc3_0),.clk(gclk));
	jdff dff_A_kPNf8Wh39_0(.dout(w_dff_A_ZXyQHwlc3_0),.din(w_dff_A_kPNf8Wh39_0),.clk(gclk));
	jdff dff_B_M8u8lpIW6_1(.din(n343),.dout(w_dff_B_M8u8lpIW6_1),.clk(gclk));
	jdff dff_B_dfzaaTg61_1(.din(w_dff_B_M8u8lpIW6_1),.dout(w_dff_B_dfzaaTg61_1),.clk(gclk));
	jdff dff_B_5JtSqqhk2_1(.din(w_dff_B_dfzaaTg61_1),.dout(w_dff_B_5JtSqqhk2_1),.clk(gclk));
	jdff dff_B_XEQnazf80_1(.din(w_dff_B_5JtSqqhk2_1),.dout(w_dff_B_XEQnazf80_1),.clk(gclk));
	jdff dff_B_FxFBpVrk9_1(.din(w_dff_B_XEQnazf80_1),.dout(w_dff_B_FxFBpVrk9_1),.clk(gclk));
	jdff dff_B_wJ5ruUjE4_1(.din(n344),.dout(w_dff_B_wJ5ruUjE4_1),.clk(gclk));
	jdff dff_B_NzKj01Qv2_1(.din(w_dff_B_wJ5ruUjE4_1),.dout(w_dff_B_NzKj01Qv2_1),.clk(gclk));
	jdff dff_B_maYxTiIJ7_1(.din(w_dff_B_NzKj01Qv2_1),.dout(w_dff_B_maYxTiIJ7_1),.clk(gclk));
	jdff dff_B_BU8RXXAE6_1(.din(w_dff_B_maYxTiIJ7_1),.dout(w_dff_B_BU8RXXAE6_1),.clk(gclk));
	jdff dff_B_zCTWHUUc0_0(.din(n231),.dout(w_dff_B_zCTWHUUc0_0),.clk(gclk));
	jdff dff_A_U8VkxY2G1_0(.dout(w_n230_0[0]),.din(w_dff_A_U8VkxY2G1_0),.clk(gclk));
	jdff dff_B_HJhhk2Za1_1(.din(n227),.dout(w_dff_B_HJhhk2Za1_1),.clk(gclk));
	jdff dff_A_yAdCop6Z3_0(.dout(w_n228_0[0]),.din(w_dff_A_yAdCop6Z3_0),.clk(gclk));
	jdff dff_A_xMfnZn0I7_0(.dout(w_dff_A_yAdCop6Z3_0),.din(w_dff_A_xMfnZn0I7_0),.clk(gclk));
	jdff dff_A_C4oHFx8z8_0(.dout(w_dff_A_xMfnZn0I7_0),.din(w_dff_A_C4oHFx8z8_0),.clk(gclk));
	jdff dff_A_0UYYGZAd7_1(.dout(w_G195gat_1[1]),.din(w_dff_A_0UYYGZAd7_1),.clk(gclk));
	jdff dff_A_dKYJ5aZf9_1(.dout(w_dff_A_0UYYGZAd7_1),.din(w_dff_A_dKYJ5aZf9_1),.clk(gclk));
	jdff dff_A_aZn7jFaW6_1(.dout(w_dff_A_dKYJ5aZf9_1),.din(w_dff_A_aZn7jFaW6_1),.clk(gclk));
	jdff dff_A_9LjsbrFf8_1(.dout(w_dff_A_aZn7jFaW6_1),.din(w_dff_A_9LjsbrFf8_1),.clk(gclk));
	jdff dff_A_pF2s8jJy7_1(.dout(w_dff_A_9LjsbrFf8_1),.din(w_dff_A_pF2s8jJy7_1),.clk(gclk));
	jdff dff_A_VB2fzTlZ8_1(.dout(w_dff_A_pF2s8jJy7_1),.din(w_dff_A_VB2fzTlZ8_1),.clk(gclk));
	jdff dff_A_h6fWmWR07_1(.dout(w_dff_A_VB2fzTlZ8_1),.din(w_dff_A_h6fWmWR07_1),.clk(gclk));
	jdff dff_A_DTUD1R403_1(.dout(w_dff_A_h6fWmWR07_1),.din(w_dff_A_DTUD1R403_1),.clk(gclk));
	jdff dff_A_JHMj1Keu4_2(.dout(w_G195gat_1[2]),.din(w_dff_A_JHMj1Keu4_2),.clk(gclk));
	jdff dff_A_NaguskDQ5_2(.dout(w_dff_A_JHMj1Keu4_2),.din(w_dff_A_NaguskDQ5_2),.clk(gclk));
	jdff dff_A_aZxjJvh80_2(.dout(w_dff_A_NaguskDQ5_2),.din(w_dff_A_aZxjJvh80_2),.clk(gclk));
	jdff dff_A_BjECwNAx5_2(.dout(w_dff_A_aZxjJvh80_2),.din(w_dff_A_BjECwNAx5_2),.clk(gclk));
	jdff dff_A_RqT43T9y2_2(.dout(w_dff_A_BjECwNAx5_2),.din(w_dff_A_RqT43T9y2_2),.clk(gclk));
	jdff dff_A_rCeAFLiN1_2(.dout(w_dff_A_RqT43T9y2_2),.din(w_dff_A_rCeAFLiN1_2),.clk(gclk));
	jdff dff_A_Qv1SyCfy9_2(.dout(w_dff_A_rCeAFLiN1_2),.din(w_dff_A_Qv1SyCfy9_2),.clk(gclk));
	jdff dff_A_fsxYyJjG3_2(.dout(w_dff_A_Qv1SyCfy9_2),.din(w_dff_A_fsxYyJjG3_2),.clk(gclk));
	jdff dff_A_t2VKqC012_1(.dout(w_G189gat_1[1]),.din(w_dff_A_t2VKqC012_1),.clk(gclk));
	jdff dff_A_rKur3qzb4_1(.dout(w_dff_A_t2VKqC012_1),.din(w_dff_A_rKur3qzb4_1),.clk(gclk));
	jdff dff_A_6FlEJPGT6_1(.dout(w_dff_A_rKur3qzb4_1),.din(w_dff_A_6FlEJPGT6_1),.clk(gclk));
	jdff dff_A_8s9P6lSF8_1(.dout(w_dff_A_6FlEJPGT6_1),.din(w_dff_A_8s9P6lSF8_1),.clk(gclk));
	jdff dff_A_ED5y1Mrd2_1(.dout(w_dff_A_8s9P6lSF8_1),.din(w_dff_A_ED5y1Mrd2_1),.clk(gclk));
	jdff dff_A_rG8SlCZZ8_1(.dout(w_dff_A_ED5y1Mrd2_1),.din(w_dff_A_rG8SlCZZ8_1),.clk(gclk));
	jdff dff_A_jN2amZtz9_1(.dout(w_dff_A_rG8SlCZZ8_1),.din(w_dff_A_jN2amZtz9_1),.clk(gclk));
	jdff dff_A_Bk71gHeV9_1(.dout(w_dff_A_jN2amZtz9_1),.din(w_dff_A_Bk71gHeV9_1),.clk(gclk));
	jdff dff_A_Ml3LPoRN6_2(.dout(w_G189gat_1[2]),.din(w_dff_A_Ml3LPoRN6_2),.clk(gclk));
	jdff dff_A_Cb2IXG5A8_2(.dout(w_dff_A_Ml3LPoRN6_2),.din(w_dff_A_Cb2IXG5A8_2),.clk(gclk));
	jdff dff_A_W7xMu0jm8_2(.dout(w_dff_A_Cb2IXG5A8_2),.din(w_dff_A_W7xMu0jm8_2),.clk(gclk));
	jdff dff_A_U46mvkgj9_2(.dout(w_dff_A_W7xMu0jm8_2),.din(w_dff_A_U46mvkgj9_2),.clk(gclk));
	jdff dff_A_KSUlxIVK5_2(.dout(w_dff_A_U46mvkgj9_2),.din(w_dff_A_KSUlxIVK5_2),.clk(gclk));
	jdff dff_A_XkLLA4j06_2(.dout(w_dff_A_KSUlxIVK5_2),.din(w_dff_A_XkLLA4j06_2),.clk(gclk));
	jdff dff_A_hMy2MXLM0_2(.dout(w_dff_A_XkLLA4j06_2),.din(w_dff_A_hMy2MXLM0_2),.clk(gclk));
	jdff dff_A_ihUrwOyU2_2(.dout(w_dff_A_hMy2MXLM0_2),.din(w_dff_A_ihUrwOyU2_2),.clk(gclk));
	jdff dff_B_7A8CQ8wf1_0(.din(n225),.dout(w_dff_B_7A8CQ8wf1_0),.clk(gclk));
	jdff dff_A_c2yYKDc01_0(.dout(w_n224_0[0]),.din(w_dff_A_c2yYKDc01_0),.clk(gclk));
	jdff dff_A_WkSOeeeh6_0(.dout(w_n223_0[0]),.din(w_dff_A_WkSOeeeh6_0),.clk(gclk));
	jdff dff_A_EEBKWNz20_0(.dout(w_dff_A_WkSOeeeh6_0),.din(w_dff_A_EEBKWNz20_0),.clk(gclk));
	jdff dff_B_rRvGpYtZ9_1(.din(n219),.dout(w_dff_B_rRvGpYtZ9_1),.clk(gclk));
	jdff dff_A_v5nfyNWc3_0(.dout(w_G121gat_0[0]),.din(w_dff_A_v5nfyNWc3_0),.clk(gclk));
	jdff dff_A_Eq6Muw3W5_0(.dout(w_dff_A_v5nfyNWc3_0),.din(w_dff_A_Eq6Muw3W5_0),.clk(gclk));
	jdff dff_A_VQx0RyiS8_0(.dout(w_dff_A_Eq6Muw3W5_0),.din(w_dff_A_VQx0RyiS8_0),.clk(gclk));
	jdff dff_A_OKECXWQi5_0(.dout(w_dff_A_VQx0RyiS8_0),.din(w_dff_A_OKECXWQi5_0),.clk(gclk));
	jdff dff_A_fyBPgIOs4_0(.dout(w_dff_A_OKECXWQi5_0),.din(w_dff_A_fyBPgIOs4_0),.clk(gclk));
	jdff dff_A_7WBawzON4_0(.dout(w_G195gat_2[0]),.din(w_dff_A_7WBawzON4_0),.clk(gclk));
	jdff dff_A_QmSLiku04_0(.dout(w_dff_A_7WBawzON4_0),.din(w_dff_A_QmSLiku04_0),.clk(gclk));
	jdff dff_A_xFXitK0D6_0(.dout(w_dff_A_QmSLiku04_0),.din(w_dff_A_xFXitK0D6_0),.clk(gclk));
	jdff dff_A_ksId0XEv9_0(.dout(w_dff_A_xFXitK0D6_0),.din(w_dff_A_ksId0XEv9_0),.clk(gclk));
	jdff dff_A_3C6fbs1i9_0(.dout(w_dff_A_ksId0XEv9_0),.din(w_dff_A_3C6fbs1i9_0),.clk(gclk));
	jdff dff_A_FMfH9g317_0(.dout(w_dff_A_3C6fbs1i9_0),.din(w_dff_A_FMfH9g317_0),.clk(gclk));
	jdff dff_A_9XhzZTb43_0(.dout(w_dff_A_FMfH9g317_0),.din(w_dff_A_9XhzZTb43_0),.clk(gclk));
	jdff dff_A_IpqDrjdh0_0(.dout(w_dff_A_9XhzZTb43_0),.din(w_dff_A_IpqDrjdh0_0),.clk(gclk));
	jdff dff_A_HZkf69Kn8_2(.dout(w_G195gat_0[2]),.din(w_dff_A_HZkf69Kn8_2),.clk(gclk));
	jdff dff_A_jrjUOp1I0_2(.dout(w_dff_A_HZkf69Kn8_2),.din(w_dff_A_jrjUOp1I0_2),.clk(gclk));
	jdff dff_A_vn9IGqtz7_2(.dout(w_dff_A_jrjUOp1I0_2),.din(w_dff_A_vn9IGqtz7_2),.clk(gclk));
	jdff dff_A_7tnFYHLD3_2(.dout(w_dff_A_vn9IGqtz7_2),.din(w_dff_A_7tnFYHLD3_2),.clk(gclk));
	jdff dff_B_HP1pRa9y2_1(.din(n214),.dout(w_dff_B_HP1pRa9y2_1),.clk(gclk));
	jdff dff_A_K4JB3bi80_1(.dout(w_G116gat_0[1]),.din(w_dff_A_K4JB3bi80_1),.clk(gclk));
	jdff dff_A_rLOPMm421_1(.dout(w_dff_A_K4JB3bi80_1),.din(w_dff_A_rLOPMm421_1),.clk(gclk));
	jdff dff_A_O2Gy59Yd5_1(.dout(w_dff_A_rLOPMm421_1),.din(w_dff_A_O2Gy59Yd5_1),.clk(gclk));
	jdff dff_A_eNwx5A8U0_1(.dout(w_dff_A_O2Gy59Yd5_1),.din(w_dff_A_eNwx5A8U0_1),.clk(gclk));
	jdff dff_A_4J4xqKLW5_1(.dout(w_dff_A_eNwx5A8U0_1),.din(w_dff_A_4J4xqKLW5_1),.clk(gclk));
	jdff dff_A_kvfY68hY2_1(.dout(w_G146gat_0[1]),.din(w_dff_A_kvfY68hY2_1),.clk(gclk));
	jdff dff_B_g8xrYXn64_2(.din(G146gat),.dout(w_dff_B_g8xrYXn64_2),.clk(gclk));
	jdff dff_B_ZDNC6rPy5_2(.din(w_dff_B_g8xrYXn64_2),.dout(w_dff_B_ZDNC6rPy5_2),.clk(gclk));
	jdff dff_B_LrlYXd8T1_2(.din(w_dff_B_ZDNC6rPy5_2),.dout(w_dff_B_LrlYXd8T1_2),.clk(gclk));
	jdff dff_B_piD0i7Xt2_2(.din(w_dff_B_LrlYXd8T1_2),.dout(w_dff_B_piD0i7Xt2_2),.clk(gclk));
	jdff dff_A_avSQB05u4_0(.dout(w_G189gat_2[0]),.din(w_dff_A_avSQB05u4_0),.clk(gclk));
	jdff dff_A_ohMpxTvy5_0(.dout(w_dff_A_avSQB05u4_0),.din(w_dff_A_ohMpxTvy5_0),.clk(gclk));
	jdff dff_A_18xIItvs4_0(.dout(w_dff_A_ohMpxTvy5_0),.din(w_dff_A_18xIItvs4_0),.clk(gclk));
	jdff dff_A_ZJEF9ZSQ7_0(.dout(w_dff_A_18xIItvs4_0),.din(w_dff_A_ZJEF9ZSQ7_0),.clk(gclk));
	jdff dff_A_uLTmUqcE9_0(.dout(w_dff_A_ZJEF9ZSQ7_0),.din(w_dff_A_uLTmUqcE9_0),.clk(gclk));
	jdff dff_A_gAhvSEBA2_0(.dout(w_dff_A_uLTmUqcE9_0),.din(w_dff_A_gAhvSEBA2_0),.clk(gclk));
	jdff dff_A_5MuUyKNx9_0(.dout(w_dff_A_gAhvSEBA2_0),.din(w_dff_A_5MuUyKNx9_0),.clk(gclk));
	jdff dff_A_PNmlGw7p8_0(.dout(w_dff_A_5MuUyKNx9_0),.din(w_dff_A_PNmlGw7p8_0),.clk(gclk));
	jdff dff_A_WKhiULLH2_2(.dout(w_G189gat_0[2]),.din(w_dff_A_WKhiULLH2_2),.clk(gclk));
	jdff dff_A_3evzTTmu8_2(.dout(w_dff_A_WKhiULLH2_2),.din(w_dff_A_3evzTTmu8_2),.clk(gclk));
	jdff dff_A_oqqOtPtr9_2(.dout(w_dff_A_3evzTTmu8_2),.din(w_dff_A_oqqOtPtr9_2),.clk(gclk));
	jdff dff_A_7awGszEe9_2(.dout(w_dff_A_oqqOtPtr9_2),.din(w_dff_A_7awGszEe9_2),.clk(gclk));
	jdff dff_B_Bj9Xhqiq0_1(.din(n197),.dout(w_dff_B_Bj9Xhqiq0_1),.clk(gclk));
	jdff dff_B_YWJF9daW1_1(.din(n198),.dout(w_dff_B_YWJF9daW1_1),.clk(gclk));
	jdff dff_B_0aZHIupd6_1(.din(w_dff_B_YWJF9daW1_1),.dout(w_dff_B_0aZHIupd6_1),.clk(gclk));
	jdff dff_B_zp8Q2MNX9_1(.din(w_dff_B_0aZHIupd6_1),.dout(w_dff_B_zp8Q2MNX9_1),.clk(gclk));
	jdff dff_B_Scid7VSd1_1(.din(w_dff_B_zp8Q2MNX9_1),.dout(w_dff_B_Scid7VSd1_1),.clk(gclk));
	jdff dff_B_6QO0Oz3U5_1(.din(w_dff_B_Scid7VSd1_1),.dout(w_dff_B_6QO0Oz3U5_1),.clk(gclk));
	jdff dff_B_kboDXVne9_1(.din(w_dff_B_6QO0Oz3U5_1),.dout(w_dff_B_kboDXVne9_1),.clk(gclk));
	jdff dff_B_l3EjJiUZ8_1(.din(w_dff_B_kboDXVne9_1),.dout(w_dff_B_l3EjJiUZ8_1),.clk(gclk));
	jdff dff_B_skd7gkZr8_1(.din(w_dff_B_l3EjJiUZ8_1),.dout(w_dff_B_skd7gkZr8_1),.clk(gclk));
	jdff dff_B_CRE4zai05_1(.din(n199),.dout(w_dff_B_CRE4zai05_1),.clk(gclk));
	jdff dff_B_aaNCrRes6_0(.din(n208),.dout(w_dff_B_aaNCrRes6_0),.clk(gclk));
	jdff dff_B_teIs8hoA6_0(.din(w_dff_B_aaNCrRes6_0),.dout(w_dff_B_teIs8hoA6_0),.clk(gclk));
	jdff dff_B_F6Wksyvu4_1(.din(n200),.dout(w_dff_B_F6Wksyvu4_1),.clk(gclk));
	jdff dff_B_Ji6T9NuC1_1(.din(w_dff_B_F6Wksyvu4_1),.dout(w_dff_B_Ji6T9NuC1_1),.clk(gclk));
	jdff dff_B_1maUqPPy8_1(.din(w_dff_B_Ji6T9NuC1_1),.dout(w_dff_B_1maUqPPy8_1),.clk(gclk));
	jdff dff_B_aGrgTfJx5_1(.din(w_dff_B_1maUqPPy8_1),.dout(w_dff_B_aGrgTfJx5_1),.clk(gclk));
	jdff dff_B_308swCCT8_1(.din(w_dff_B_aGrgTfJx5_1),.dout(w_dff_B_308swCCT8_1),.clk(gclk));
	jdff dff_B_WHqEB5UA4_1(.din(n201),.dout(w_dff_B_WHqEB5UA4_1),.clk(gclk));
	jdff dff_B_RgedzBox4_1(.din(w_dff_B_WHqEB5UA4_1),.dout(w_dff_B_RgedzBox4_1),.clk(gclk));
	jdff dff_B_zcWU9T686_1(.din(w_dff_B_RgedzBox4_1),.dout(w_dff_B_zcWU9T686_1),.clk(gclk));
	jdff dff_B_CEyhQme00_1(.din(n202),.dout(w_dff_B_CEyhQme00_1),.clk(gclk));
	jdff dff_B_OT2NGZCo5_2(.din(n143),.dout(w_dff_B_OT2NGZCo5_2),.clk(gclk));
	jdff dff_B_o62SLLAi8_2(.din(w_dff_B_OT2NGZCo5_2),.dout(w_dff_B_o62SLLAi8_2),.clk(gclk));
	jdff dff_B_weoeNh1Z2_2(.din(w_dff_B_o62SLLAi8_2),.dout(w_dff_B_weoeNh1Z2_2),.clk(gclk));
	jdff dff_B_QLqm9Rjl5_2(.din(w_dff_B_weoeNh1Z2_2),.dout(w_dff_B_QLqm9Rjl5_2),.clk(gclk));
	jdff dff_B_fqdGfhSa0_2(.din(w_dff_B_QLqm9Rjl5_2),.dout(w_dff_B_fqdGfhSa0_2),.clk(gclk));
	jdff dff_B_jlAjge222_2(.din(w_dff_B_fqdGfhSa0_2),.dout(w_dff_B_jlAjge222_2),.clk(gclk));
	jdff dff_B_PNREf1H55_2(.din(w_dff_B_jlAjge222_2),.dout(w_dff_B_PNREf1H55_2),.clk(gclk));
	jdff dff_B_O7IYYnW93_2(.din(w_dff_B_PNREf1H55_2),.dout(w_dff_B_O7IYYnW93_2),.clk(gclk));
	jdff dff_B_W8buxaVQ2_2(.din(w_dff_B_O7IYYnW93_2),.dout(w_dff_B_W8buxaVQ2_2),.clk(gclk));
	jdff dff_A_eI1hEaNQ3_0(.dout(w_G261gat_0[0]),.din(w_dff_A_eI1hEaNQ3_0),.clk(gclk));
	jdff dff_A_eEZuc3JX5_0(.dout(w_dff_A_eI1hEaNQ3_0),.din(w_dff_A_eEZuc3JX5_0),.clk(gclk));
	jdff dff_A_gzGnGGAu2_0(.dout(w_dff_A_eEZuc3JX5_0),.din(w_dff_A_gzGnGGAu2_0),.clk(gclk));
	jdff dff_A_BXzaIjEq7_0(.dout(w_dff_A_gzGnGGAu2_0),.din(w_dff_A_BXzaIjEq7_0),.clk(gclk));
	jdff dff_A_6N9GaMhU6_0(.dout(w_dff_A_BXzaIjEq7_0),.din(w_dff_A_6N9GaMhU6_0),.clk(gclk));
	jdff dff_A_PqkO6H438_0(.dout(w_dff_A_6N9GaMhU6_0),.din(w_dff_A_PqkO6H438_0),.clk(gclk));
	jdff dff_A_MDCxWnEX0_0(.dout(w_dff_A_PqkO6H438_0),.din(w_dff_A_MDCxWnEX0_0),.clk(gclk));
	jdff dff_A_SkK6WUdn5_0(.dout(w_dff_A_MDCxWnEX0_0),.din(w_dff_A_SkK6WUdn5_0),.clk(gclk));
	jdff dff_A_EPD7r3wi6_0(.dout(w_dff_A_SkK6WUdn5_0),.din(w_dff_A_EPD7r3wi6_0),.clk(gclk));
	jdff dff_A_Zx2Dsoyo2_1(.dout(w_G261gat_0[1]),.din(w_dff_A_Zx2Dsoyo2_1),.clk(gclk));
	jdff dff_A_xVZx3eOO5_1(.dout(w_dff_A_Zx2Dsoyo2_1),.din(w_dff_A_xVZx3eOO5_1),.clk(gclk));
	jdff dff_A_yy4Xcum80_1(.dout(w_dff_A_xVZx3eOO5_1),.din(w_dff_A_yy4Xcum80_1),.clk(gclk));
	jdff dff_A_IKIePTK22_1(.dout(w_dff_A_yy4Xcum80_1),.din(w_dff_A_IKIePTK22_1),.clk(gclk));
	jdff dff_A_xCoL9wn42_1(.dout(w_dff_A_IKIePTK22_1),.din(w_dff_A_xCoL9wn42_1),.clk(gclk));
	jdff dff_A_ArIkvXv60_1(.dout(w_dff_A_xCoL9wn42_1),.din(w_dff_A_ArIkvXv60_1),.clk(gclk));
	jdff dff_A_xODEzUgS7_1(.dout(w_dff_A_ArIkvXv60_1),.din(w_dff_A_xODEzUgS7_1),.clk(gclk));
	jdff dff_A_gQitHaxw7_1(.dout(w_dff_A_xODEzUgS7_1),.din(w_dff_A_gQitHaxw7_1),.clk(gclk));
	jdff dff_A_fwjkoGRV6_1(.dout(w_dff_A_gQitHaxw7_1),.din(w_dff_A_fwjkoGRV6_1),.clk(gclk));
	jdff dff_A_bSvZyBQD0_0(.dout(w_n196_0[0]),.din(w_dff_A_bSvZyBQD0_0),.clk(gclk));
	jdff dff_A_WmCX4QAd4_1(.dout(w_n154_0[1]),.din(w_dff_A_WmCX4QAd4_1),.clk(gclk));
	jdff dff_A_Ozb6AsFn9_0(.dout(w_G126gat_0[0]),.din(w_dff_A_Ozb6AsFn9_0),.clk(gclk));
	jdff dff_A_BZzvcps99_0(.dout(w_dff_A_Ozb6AsFn9_0),.din(w_dff_A_BZzvcps99_0),.clk(gclk));
	jdff dff_A_NmSiOZAZ2_0(.dout(w_dff_A_BZzvcps99_0),.din(w_dff_A_NmSiOZAZ2_0),.clk(gclk));
	jdff dff_A_9Q1Z28lf8_0(.dout(w_dff_A_NmSiOZAZ2_0),.din(w_dff_A_9Q1Z28lf8_0),.clk(gclk));
	jdff dff_A_WeingIaf9_0(.dout(w_dff_A_9Q1Z28lf8_0),.din(w_dff_A_WeingIaf9_0),.clk(gclk));
	jdff dff_A_GWKmMSds5_1(.dout(w_G201gat_1[1]),.din(w_dff_A_GWKmMSds5_1),.clk(gclk));
	jdff dff_A_MZNSBQMW6_1(.dout(w_dff_A_GWKmMSds5_1),.din(w_dff_A_MZNSBQMW6_1),.clk(gclk));
	jdff dff_A_dHCIQLS56_1(.dout(w_dff_A_MZNSBQMW6_1),.din(w_dff_A_dHCIQLS56_1),.clk(gclk));
	jdff dff_A_CqfVyh1X8_1(.dout(w_dff_A_dHCIQLS56_1),.din(w_dff_A_CqfVyh1X8_1),.clk(gclk));
	jdff dff_A_ZoFaf9jF1_1(.dout(w_dff_A_CqfVyh1X8_1),.din(w_dff_A_ZoFaf9jF1_1),.clk(gclk));
	jdff dff_A_faiL1H6P0_1(.dout(w_dff_A_ZoFaf9jF1_1),.din(w_dff_A_faiL1H6P0_1),.clk(gclk));
	jdff dff_A_nbBr9Jmr4_1(.dout(w_dff_A_faiL1H6P0_1),.din(w_dff_A_nbBr9Jmr4_1),.clk(gclk));
	jdff dff_A_KCKcfahM1_1(.dout(w_dff_A_nbBr9Jmr4_1),.din(w_dff_A_KCKcfahM1_1),.clk(gclk));
	jdff dff_A_fqYz0gn91_2(.dout(w_G201gat_1[2]),.din(w_dff_A_fqYz0gn91_2),.clk(gclk));
	jdff dff_A_KkK22m7r8_2(.dout(w_dff_A_fqYz0gn91_2),.din(w_dff_A_KkK22m7r8_2),.clk(gclk));
	jdff dff_A_WyfH7fgS7_2(.dout(w_dff_A_KkK22m7r8_2),.din(w_dff_A_WyfH7fgS7_2),.clk(gclk));
	jdff dff_A_bt1n3pah3_2(.dout(w_dff_A_WyfH7fgS7_2),.din(w_dff_A_bt1n3pah3_2),.clk(gclk));
	jdff dff_A_nNciEC3p7_2(.dout(w_G201gat_0[2]),.din(w_dff_A_nNciEC3p7_2),.clk(gclk));
	jdff dff_A_Q4679qAd0_2(.dout(w_dff_A_nNciEC3p7_2),.din(w_dff_A_Q4679qAd0_2),.clk(gclk));
	jdff dff_A_f9bvKH217_2(.dout(w_dff_A_Q4679qAd0_2),.din(w_dff_A_f9bvKH217_2),.clk(gclk));
	jdff dff_A_I0eyeOdC1_2(.dout(w_dff_A_f9bvKH217_2),.din(w_dff_A_I0eyeOdC1_2),.clk(gclk));
	jdff dff_A_V0DLYVtI8_2(.dout(w_dff_A_I0eyeOdC1_2),.din(w_dff_A_V0DLYVtI8_2),.clk(gclk));
	jdff dff_A_AWcbRMiQ4_2(.dout(w_dff_A_V0DLYVtI8_2),.din(w_dff_A_AWcbRMiQ4_2),.clk(gclk));
	jdff dff_A_zpr6cEBJ4_2(.dout(w_dff_A_AWcbRMiQ4_2),.din(w_dff_A_zpr6cEBJ4_2),.clk(gclk));
	jdff dff_A_QZg04gcl8_2(.dout(w_dff_A_zpr6cEBJ4_2),.din(w_dff_A_QZg04gcl8_2),.clk(gclk));
	jdff dff_A_7PhRkVid1_1(.dout(w_n303_0[1]),.din(w_dff_A_7PhRkVid1_1),.clk(gclk));
	jdff dff_A_dr9yFtro2_1(.dout(w_dff_A_7PhRkVid1_1),.din(w_dff_A_dr9yFtro2_1),.clk(gclk));
	jdff dff_A_eXq9rgTs1_1(.dout(w_dff_A_dr9yFtro2_1),.din(w_dff_A_eXq9rgTs1_1),.clk(gclk));
	jdff dff_A_yqcEP5M88_1(.dout(w_dff_A_eXq9rgTs1_1),.din(w_dff_A_yqcEP5M88_1),.clk(gclk));
	jdff dff_A_d6UTlw6b8_1(.dout(w_n302_0[1]),.din(w_dff_A_d6UTlw6b8_1),.clk(gclk));
	jdff dff_A_t1XsacIZ5_1(.dout(w_dff_A_d6UTlw6b8_1),.din(w_dff_A_t1XsacIZ5_1),.clk(gclk));
	jdff dff_A_VUDk8WcB1_1(.dout(w_dff_A_t1XsacIZ5_1),.din(w_dff_A_VUDk8WcB1_1),.clk(gclk));
	jdff dff_A_gKAnkFhG8_1(.dout(w_dff_A_VUDk8WcB1_1),.din(w_dff_A_gKAnkFhG8_1),.clk(gclk));
	jdff dff_A_YWGPJBXF6_1(.dout(w_dff_A_gKAnkFhG8_1),.din(w_dff_A_YWGPJBXF6_1),.clk(gclk));
	jdff dff_B_DGX4PC4T2_1(.din(n190),.dout(w_dff_B_DGX4PC4T2_1),.clk(gclk));
	jdff dff_A_HVyJZuJi9_1(.dout(w_G111gat_0[1]),.din(w_dff_A_HVyJZuJi9_1),.clk(gclk));
	jdff dff_A_iAL4fUL74_1(.dout(w_dff_A_HVyJZuJi9_1),.din(w_dff_A_iAL4fUL74_1),.clk(gclk));
	jdff dff_A_VWf8y2e67_1(.dout(w_dff_A_iAL4fUL74_1),.din(w_dff_A_VWf8y2e67_1),.clk(gclk));
	jdff dff_A_7RlY8bLN9_1(.dout(w_dff_A_VWf8y2e67_1),.din(w_dff_A_7RlY8bLN9_1),.clk(gclk));
	jdff dff_A_uIjmtxar9_1(.dout(w_dff_A_7RlY8bLN9_1),.din(w_dff_A_uIjmtxar9_1),.clk(gclk));
	jdff dff_A_tfwqjyyU3_1(.dout(w_n165_1[1]),.din(w_dff_A_tfwqjyyU3_1),.clk(gclk));
	jdff dff_A_EftGHX5V2_1(.dout(w_dff_A_tfwqjyyU3_1),.din(w_dff_A_EftGHX5V2_1),.clk(gclk));
	jdff dff_A_8oI9TO9J2_2(.dout(w_n165_1[2]),.din(w_dff_A_8oI9TO9J2_2),.clk(gclk));
	jdff dff_A_vUIuLwci3_2(.dout(w_dff_A_8oI9TO9J2_2),.din(w_dff_A_vUIuLwci3_2),.clk(gclk));
	jdff dff_A_ddvr60bq8_1(.dout(w_n165_0[1]),.din(w_dff_A_ddvr60bq8_1),.clk(gclk));
	jdff dff_A_rKyPGpVz7_1(.dout(w_dff_A_ddvr60bq8_1),.din(w_dff_A_rKyPGpVz7_1),.clk(gclk));
	jdff dff_A_QlSQTq4C2_2(.dout(w_n165_0[2]),.din(w_dff_A_QlSQTq4C2_2),.clk(gclk));
	jdff dff_A_w9FWJmsQ3_2(.dout(w_dff_A_QlSQTq4C2_2),.din(w_dff_A_w9FWJmsQ3_2),.clk(gclk));
	jdff dff_B_8kWAgWBF9_0(.din(n164),.dout(w_dff_B_8kWAgWBF9_0),.clk(gclk));
	jdff dff_A_wI6DRQ022_0(.dout(w_n96_0[0]),.din(w_dff_A_wI6DRQ022_0),.clk(gclk));
	jdff dff_A_jds7d27L4_0(.dout(w_dff_A_wI6DRQ022_0),.din(w_dff_A_jds7d27L4_0),.clk(gclk));
	jdff dff_A_Wzfu0KCD4_0(.dout(w_dff_A_jds7d27L4_0),.din(w_dff_A_Wzfu0KCD4_0),.clk(gclk));
	jdff dff_A_XR9CSE6t7_1(.dout(w_G143gat_0[1]),.din(w_dff_A_XR9CSE6t7_1),.clk(gclk));
	jdff dff_B_XOaP6XDE5_2(.din(G143gat),.dout(w_dff_B_XOaP6XDE5_2),.clk(gclk));
	jdff dff_B_ttmPs0EQ7_2(.din(w_dff_B_XOaP6XDE5_2),.dout(w_dff_B_ttmPs0EQ7_2),.clk(gclk));
	jdff dff_B_zp4lH0lP0_2(.din(w_dff_B_ttmPs0EQ7_2),.dout(w_dff_B_zp4lH0lP0_2),.clk(gclk));
	jdff dff_B_SKyVliyN8_2(.din(w_dff_B_zp4lH0lP0_2),.dout(w_dff_B_SKyVliyN8_2),.clk(gclk));
	jdff dff_A_1W0H5qBI4_0(.dout(w_G183gat_1[0]),.din(w_dff_A_1W0H5qBI4_0),.clk(gclk));
	jdff dff_A_wSAYqYIq6_0(.dout(w_dff_A_1W0H5qBI4_0),.din(w_dff_A_wSAYqYIq6_0),.clk(gclk));
	jdff dff_A_KTxNf5Mh6_0(.dout(w_dff_A_wSAYqYIq6_0),.din(w_dff_A_KTxNf5Mh6_0),.clk(gclk));
	jdff dff_A_PomoBPfT4_0(.dout(w_dff_A_KTxNf5Mh6_0),.din(w_dff_A_PomoBPfT4_0),.clk(gclk));
	jdff dff_A_jMBcLWEX5_0(.dout(w_dff_A_PomoBPfT4_0),.din(w_dff_A_jMBcLWEX5_0),.clk(gclk));
	jdff dff_A_ClVOk8HB2_0(.dout(w_dff_A_jMBcLWEX5_0),.din(w_dff_A_ClVOk8HB2_0),.clk(gclk));
	jdff dff_A_UztsRuXl7_0(.dout(w_dff_A_ClVOk8HB2_0),.din(w_dff_A_UztsRuXl7_0),.clk(gclk));
	jdff dff_A_vSNtDbIa9_0(.dout(w_dff_A_UztsRuXl7_0),.din(w_dff_A_vSNtDbIa9_0),.clk(gclk));
	jdff dff_A_jXmvuQg96_1(.dout(w_G183gat_1[1]),.din(w_dff_A_jXmvuQg96_1),.clk(gclk));
	jdff dff_A_pWHCK0eD6_1(.dout(w_dff_A_jXmvuQg96_1),.din(w_dff_A_pWHCK0eD6_1),.clk(gclk));
	jdff dff_A_RE7WW2799_1(.dout(w_dff_A_pWHCK0eD6_1),.din(w_dff_A_RE7WW2799_1),.clk(gclk));
	jdff dff_A_M3JOp4nt7_1(.dout(w_dff_A_RE7WW2799_1),.din(w_dff_A_M3JOp4nt7_1),.clk(gclk));
	jdff dff_A_MAXA9IyN0_2(.dout(w_G183gat_0[2]),.din(w_dff_A_MAXA9IyN0_2),.clk(gclk));
	jdff dff_A_bCaJ9rnB5_2(.dout(w_dff_A_MAXA9IyN0_2),.din(w_dff_A_bCaJ9rnB5_2),.clk(gclk));
	jdff dff_A_iyvIJL261_2(.dout(w_dff_A_bCaJ9rnB5_2),.din(w_dff_A_iyvIJL261_2),.clk(gclk));
	jdff dff_A_jKmKaN8m1_2(.dout(w_dff_A_iyvIJL261_2),.din(w_dff_A_jKmKaN8m1_2),.clk(gclk));
	jdff dff_A_i0ZiWJD53_2(.dout(w_dff_A_jKmKaN8m1_2),.din(w_dff_A_i0ZiWJD53_2),.clk(gclk));
	jdff dff_A_wjUNbkYd0_2(.dout(w_dff_A_i0ZiWJD53_2),.din(w_dff_A_wjUNbkYd0_2),.clk(gclk));
	jdff dff_A_NrRqS20P0_2(.dout(w_dff_A_wjUNbkYd0_2),.din(w_dff_A_NrRqS20P0_2),.clk(gclk));
	jdff dff_A_bESZbtfo6_2(.dout(w_dff_A_NrRqS20P0_2),.din(w_dff_A_bESZbtfo6_2),.clk(gclk));
	jdff dff_A_mO5uSkrM3_0(.dout(w_n335_0[0]),.din(w_dff_A_mO5uSkrM3_0),.clk(gclk));
	jdff dff_A_ZBKepXBW4_0(.dout(w_dff_A_mO5uSkrM3_0),.din(w_dff_A_ZBKepXBW4_0),.clk(gclk));
	jdff dff_A_iYAmN6LJ7_0(.dout(w_dff_A_ZBKepXBW4_0),.din(w_dff_A_iYAmN6LJ7_0),.clk(gclk));
	jdff dff_A_yaXvQ9sw2_0(.dout(w_dff_A_iYAmN6LJ7_0),.din(w_dff_A_yaXvQ9sw2_0),.clk(gclk));
	jdff dff_A_hM2aoxTy5_0(.dout(w_dff_A_yaXvQ9sw2_0),.din(w_dff_A_hM2aoxTy5_0),.clk(gclk));
	jdff dff_A_K8RBRrLP4_0(.dout(w_dff_A_hM2aoxTy5_0),.din(w_dff_A_K8RBRrLP4_0),.clk(gclk));
	jdff dff_A_PBBSU47T0_0(.dout(w_dff_A_K8RBRrLP4_0),.din(w_dff_A_PBBSU47T0_0),.clk(gclk));
	jdff dff_A_AQyWoWVP1_0(.dout(w_dff_A_PBBSU47T0_0),.din(w_dff_A_AQyWoWVP1_0),.clk(gclk));
	jdff dff_B_Ts3otrzS6_0(.din(n325),.dout(w_dff_B_Ts3otrzS6_0),.clk(gclk));
	jdff dff_B_6AipjvpJ7_0(.din(w_dff_B_Ts3otrzS6_0),.dout(w_dff_B_6AipjvpJ7_0),.clk(gclk));
	jdff dff_B_p6SyBldd6_0(.din(w_dff_B_6AipjvpJ7_0),.dout(w_dff_B_p6SyBldd6_0),.clk(gclk));
	jdff dff_A_QTP6IFPs4_0(.dout(w_G153gat_0[0]),.din(w_dff_A_QTP6IFPs4_0),.clk(gclk));
	jdff dff_A_d8ZqSQZm5_0(.dout(w_dff_A_QTP6IFPs4_0),.din(w_dff_A_d8ZqSQZm5_0),.clk(gclk));
	jdff dff_A_wMZJN35v9_0(.dout(w_dff_A_d8ZqSQZm5_0),.din(w_dff_A_wMZJN35v9_0),.clk(gclk));
	jdff dff_A_X6eRaYX78_0(.dout(w_dff_A_wMZJN35v9_0),.din(w_dff_A_X6eRaYX78_0),.clk(gclk));
	jdff dff_A_HEsdDwwn8_2(.dout(w_G153gat_0[2]),.din(w_dff_A_HEsdDwwn8_2),.clk(gclk));
	jdff dff_A_Jw8bTo2j2_2(.dout(w_dff_A_HEsdDwwn8_2),.din(w_dff_A_Jw8bTo2j2_2),.clk(gclk));
	jdff dff_A_6pFHfPs42_2(.dout(w_dff_A_Jw8bTo2j2_2),.din(w_dff_A_6pFHfPs42_2),.clk(gclk));
	jdff dff_A_SVAwRhBm6_2(.dout(w_dff_A_6pFHfPs42_2),.din(w_dff_A_SVAwRhBm6_2),.clk(gclk));
	jdff dff_A_qQHNDwii7_2(.dout(w_dff_A_SVAwRhBm6_2),.din(w_dff_A_qQHNDwii7_2),.clk(gclk));
	jdff dff_A_yWMPujIT7_0(.dout(w_G106gat_0[0]),.din(w_dff_A_yWMPujIT7_0),.clk(gclk));
	jdff dff_A_AGG8RYi54_0(.dout(w_dff_A_yWMPujIT7_0),.din(w_dff_A_AGG8RYi54_0),.clk(gclk));
	jdff dff_A_ajWd8BSR1_0(.dout(w_dff_A_AGG8RYi54_0),.din(w_dff_A_ajWd8BSR1_0),.clk(gclk));
	jdff dff_A_NUAbXkWe9_0(.dout(w_dff_A_ajWd8BSR1_0),.din(w_dff_A_NUAbXkWe9_0),.clk(gclk));
	jdff dff_A_7M8ANXzy7_0(.dout(w_dff_A_NUAbXkWe9_0),.din(w_dff_A_7M8ANXzy7_0),.clk(gclk));
	jdff dff_A_yD0VGvYK8_1(.dout(w_G177gat_1[1]),.din(w_dff_A_yD0VGvYK8_1),.clk(gclk));
	jdff dff_A_FgeEyTeZ8_1(.dout(w_dff_A_yD0VGvYK8_1),.din(w_dff_A_FgeEyTeZ8_1),.clk(gclk));
	jdff dff_A_1tBzBOUQ3_1(.dout(w_dff_A_FgeEyTeZ8_1),.din(w_dff_A_1tBzBOUQ3_1),.clk(gclk));
	jdff dff_A_j2xZuIC02_1(.dout(w_dff_A_1tBzBOUQ3_1),.din(w_dff_A_j2xZuIC02_1),.clk(gclk));
	jdff dff_A_yeHP93kZ5_1(.dout(w_dff_A_j2xZuIC02_1),.din(w_dff_A_yeHP93kZ5_1),.clk(gclk));
	jdff dff_A_x3c0XfEU5_1(.dout(w_dff_A_yeHP93kZ5_1),.din(w_dff_A_x3c0XfEU5_1),.clk(gclk));
	jdff dff_A_m4k7EtwD6_1(.dout(w_dff_A_x3c0XfEU5_1),.din(w_dff_A_m4k7EtwD6_1),.clk(gclk));
	jdff dff_A_BdwHBUHD2_2(.dout(w_G177gat_1[2]),.din(w_dff_A_BdwHBUHD2_2),.clk(gclk));
	jdff dff_A_KMn96lEg1_2(.dout(w_dff_A_BdwHBUHD2_2),.din(w_dff_A_KMn96lEg1_2),.clk(gclk));
	jdff dff_A_CY8P0kfJ7_2(.dout(w_dff_A_KMn96lEg1_2),.din(w_dff_A_CY8P0kfJ7_2),.clk(gclk));
	jdff dff_A_WSKquXtZ5_2(.dout(w_dff_A_CY8P0kfJ7_2),.din(w_dff_A_WSKquXtZ5_2),.clk(gclk));
	jdff dff_A_nNQ9DpNP8_2(.dout(w_dff_A_WSKquXtZ5_2),.din(w_dff_A_nNQ9DpNP8_2),.clk(gclk));
	jdff dff_A_MTZAPu169_2(.dout(w_dff_A_nNQ9DpNP8_2),.din(w_dff_A_MTZAPu169_2),.clk(gclk));
	jdff dff_A_szDrL2Wm8_2(.dout(w_dff_A_MTZAPu169_2),.din(w_dff_A_szDrL2Wm8_2),.clk(gclk));
	jdff dff_A_Z1jsBvNe5_2(.dout(w_G177gat_0[2]),.din(w_dff_A_Z1jsBvNe5_2),.clk(gclk));
	jdff dff_A_KmZYAzur6_2(.dout(w_dff_A_Z1jsBvNe5_2),.din(w_dff_A_KmZYAzur6_2),.clk(gclk));
	jdff dff_A_cHBGzICT0_2(.dout(w_dff_A_KmZYAzur6_2),.din(w_dff_A_cHBGzICT0_2),.clk(gclk));
	jdff dff_A_rP3rK1Vr4_2(.dout(w_dff_A_cHBGzICT0_2),.din(w_dff_A_rP3rK1Vr4_2),.clk(gclk));
	jdff dff_A_ECHHZQPu9_1(.dout(w_n405_0[1]),.din(w_dff_A_ECHHZQPu9_1),.clk(gclk));
	jdff dff_A_XoYtyOy69_1(.dout(w_dff_A_ECHHZQPu9_1),.din(w_dff_A_XoYtyOy69_1),.clk(gclk));
	jdff dff_A_a07NDFPc2_1(.dout(w_dff_A_XoYtyOy69_1),.din(w_dff_A_a07NDFPc2_1),.clk(gclk));
	jdff dff_A_FH4QgV1M8_1(.dout(w_dff_A_a07NDFPc2_1),.din(w_dff_A_FH4QgV1M8_1),.clk(gclk));
	jdff dff_A_cM7tMsys0_1(.dout(w_dff_A_FH4QgV1M8_1),.din(w_dff_A_cM7tMsys0_1),.clk(gclk));
	jdff dff_A_jvyYKYyr3_1(.dout(w_dff_A_cM7tMsys0_1),.din(w_dff_A_jvyYKYyr3_1),.clk(gclk));
	jdff dff_A_qjnqF0wv6_1(.dout(w_dff_A_jvyYKYyr3_1),.din(w_dff_A_qjnqF0wv6_1),.clk(gclk));
	jdff dff_A_XaSQRJzn9_1(.dout(w_dff_A_qjnqF0wv6_1),.din(w_dff_A_XaSQRJzn9_1),.clk(gclk));
	jdff dff_A_t8uQFiOZ9_1(.dout(w_dff_A_XaSQRJzn9_1),.din(w_dff_A_t8uQFiOZ9_1),.clk(gclk));
	jdff dff_B_zM4IdtOI4_0(.din(n318),.dout(w_dff_B_zM4IdtOI4_0),.clk(gclk));
	jdff dff_B_vUYxz9TH0_0(.din(w_dff_B_zM4IdtOI4_0),.dout(w_dff_B_vUYxz9TH0_0),.clk(gclk));
	jdff dff_B_yNPXiZOq1_0(.din(w_dff_B_vUYxz9TH0_0),.dout(w_dff_B_yNPXiZOq1_0),.clk(gclk));
	jdff dff_B_b3prPnl21_0(.din(n295),.dout(w_dff_B_b3prPnl21_0),.clk(gclk));
	jdff dff_A_LRt7OTZo0_0(.dout(w_G17gat_1[0]),.din(w_dff_A_LRt7OTZo0_0),.clk(gclk));
	jdff dff_A_DFPhiLNs1_2(.dout(w_G17gat_1[2]),.din(w_dff_A_DFPhiLNs1_2),.clk(gclk));
	jdff dff_A_yRtBaMq77_2(.dout(w_dff_A_DFPhiLNs1_2),.din(w_dff_A_yRtBaMq77_2),.clk(gclk));
	jdff dff_A_v4FSawgS7_2(.dout(w_dff_A_yRtBaMq77_2),.din(w_dff_A_v4FSawgS7_2),.clk(gclk));
	jdff dff_A_nlkU6uhQ0_0(.dout(w_G80gat_0[0]),.din(w_dff_A_nlkU6uhQ0_0),.clk(gclk));
	jdff dff_A_A9E8vdJ38_2(.dout(w_G80gat_0[2]),.din(w_dff_A_A9E8vdJ38_2),.clk(gclk));
	jdff dff_A_RDYRiz6I3_0(.dout(w_G55gat_0[0]),.din(w_dff_A_RDYRiz6I3_0),.clk(gclk));
	jdff dff_A_bibeQP7Q3_0(.dout(w_dff_A_RDYRiz6I3_0),.din(w_dff_A_bibeQP7Q3_0),.clk(gclk));
	jdff dff_A_49kWzJ3N9_0(.dout(w_dff_A_bibeQP7Q3_0),.din(w_dff_A_49kWzJ3N9_0),.clk(gclk));
	jdff dff_A_vRztP4pg7_1(.dout(w_G55gat_0[1]),.din(w_dff_A_vRztP4pg7_1),.clk(gclk));
	jdff dff_A_QhYn5t4m1_1(.dout(w_G149gat_0[1]),.din(w_dff_A_QhYn5t4m1_1),.clk(gclk));
	jdff dff_B_zvOTUrU43_2(.din(G149gat),.dout(w_dff_B_zvOTUrU43_2),.clk(gclk));
	jdff dff_B_Zt7zWCQB8_2(.din(w_dff_B_zvOTUrU43_2),.dout(w_dff_B_Zt7zWCQB8_2),.clk(gclk));
	jdff dff_B_pL2mCnru0_2(.din(w_dff_B_Zt7zWCQB8_2),.dout(w_dff_B_pL2mCnru0_2),.clk(gclk));
	jdff dff_B_ds0xvXlA6_2(.din(w_dff_B_pL2mCnru0_2),.dout(w_dff_B_ds0xvXlA6_2),.clk(gclk));
	jdff dff_B_ZRw0s8gv8_0(.din(n152),.dout(w_dff_B_ZRw0s8gv8_0),.clk(gclk));
	jdff dff_A_jbDHMsX74_0(.dout(w_n149_0[0]),.din(w_dff_A_jbDHMsX74_0),.clk(gclk));
	jdff dff_A_WXECFDTI9_0(.dout(w_dff_A_jbDHMsX74_0),.din(w_dff_A_WXECFDTI9_0),.clk(gclk));
	jdff dff_B_7pT4tBQP9_0(.din(n147),.dout(w_dff_B_7pT4tBQP9_0),.clk(gclk));
	jdff dff_A_8DmXtU3j6_1(.dout(w_G51gat_1[1]),.din(w_dff_A_8DmXtU3j6_1),.clk(gclk));
	jdff dff_A_iI9RsNaw6_1(.dout(w_G1gat_0[1]),.din(w_dff_A_iI9RsNaw6_1),.clk(gclk));
	jdff dff_A_HavkOJJE6_1(.dout(w_dff_A_iI9RsNaw6_1),.din(w_dff_A_HavkOJJE6_1),.clk(gclk));
	jdff dff_A_bywnkVAZ2_1(.dout(w_dff_A_HavkOJJE6_1),.din(w_dff_A_bywnkVAZ2_1),.clk(gclk));
	jdff dff_A_i8iMz5ip7_1(.dout(w_dff_A_bywnkVAZ2_1),.din(w_dff_A_i8iMz5ip7_1),.clk(gclk));
	jdff dff_A_3vyI5rie3_1(.dout(w_dff_A_i8iMz5ip7_1),.din(w_dff_A_3vyI5rie3_1),.clk(gclk));
	jdff dff_A_JzK7kycc4_1(.dout(w_G42gat_1[1]),.din(w_dff_A_JzK7kycc4_1),.clk(gclk));
	jdff dff_A_qtEIuVFu9_1(.dout(w_G42gat_0[1]),.din(w_dff_A_qtEIuVFu9_1),.clk(gclk));
	jdff dff_A_EDqdme8J4_1(.dout(w_G101gat_0[1]),.din(w_dff_A_EDqdme8J4_1),.clk(gclk));
	jdff dff_A_oOBWseRU9_1(.dout(w_dff_A_EDqdme8J4_1),.din(w_dff_A_oOBWseRU9_1),.clk(gclk));
	jdff dff_A_be5oHboV7_1(.dout(w_dff_A_oOBWseRU9_1),.din(w_dff_A_be5oHboV7_1),.clk(gclk));
	jdff dff_A_YZrrfRrS1_1(.dout(w_dff_A_be5oHboV7_1),.din(w_dff_A_YZrrfRrS1_1),.clk(gclk));
	jdff dff_A_nayQiYXK3_1(.dout(w_dff_A_YZrrfRrS1_1),.din(w_dff_A_nayQiYXK3_1),.clk(gclk));
	jdff dff_A_9tSlHmkX2_1(.dout(w_G171gat_1[1]),.din(w_dff_A_9tSlHmkX2_1),.clk(gclk));
	jdff dff_A_0OEzxPyU6_1(.dout(w_dff_A_9tSlHmkX2_1),.din(w_dff_A_0OEzxPyU6_1),.clk(gclk));
	jdff dff_A_Jr6sG1Ph8_1(.dout(w_dff_A_0OEzxPyU6_1),.din(w_dff_A_Jr6sG1Ph8_1),.clk(gclk));
	jdff dff_A_izl34Adi5_1(.dout(w_dff_A_Jr6sG1Ph8_1),.din(w_dff_A_izl34Adi5_1),.clk(gclk));
	jdff dff_A_RHfp2CIP1_1(.dout(w_dff_A_izl34Adi5_1),.din(w_dff_A_RHfp2CIP1_1),.clk(gclk));
	jdff dff_A_ryF2tkFQ7_1(.dout(w_dff_A_RHfp2CIP1_1),.din(w_dff_A_ryF2tkFQ7_1),.clk(gclk));
	jdff dff_A_qRKbhJJt7_1(.dout(w_dff_A_ryF2tkFQ7_1),.din(w_dff_A_qRKbhJJt7_1),.clk(gclk));
	jdff dff_A_1E524EgH1_2(.dout(w_G171gat_1[2]),.din(w_dff_A_1E524EgH1_2),.clk(gclk));
	jdff dff_A_5DUnFiR40_2(.dout(w_dff_A_1E524EgH1_2),.din(w_dff_A_5DUnFiR40_2),.clk(gclk));
	jdff dff_A_GkJHd3ou9_2(.dout(w_dff_A_5DUnFiR40_2),.din(w_dff_A_GkJHd3ou9_2),.clk(gclk));
	jdff dff_A_zIU79f7v9_2(.dout(w_dff_A_GkJHd3ou9_2),.din(w_dff_A_zIU79f7v9_2),.clk(gclk));
	jdff dff_A_AwXPWF3r1_2(.dout(w_dff_A_zIU79f7v9_2),.din(w_dff_A_AwXPWF3r1_2),.clk(gclk));
	jdff dff_A_moQLh0bi9_2(.dout(w_dff_A_AwXPWF3r1_2),.din(w_dff_A_moQLh0bi9_2),.clk(gclk));
	jdff dff_A_zDzKJnBE0_2(.dout(w_dff_A_moQLh0bi9_2),.din(w_dff_A_zDzKJnBE0_2),.clk(gclk));
	jdff dff_A_wkhht0JW4_2(.dout(w_G171gat_0[2]),.din(w_dff_A_wkhht0JW4_2),.clk(gclk));
	jdff dff_A_zjRwJyqb7_2(.dout(w_dff_A_wkhht0JW4_2),.din(w_dff_A_zjRwJyqb7_2),.clk(gclk));
	jdff dff_A_jtDD79jW1_2(.dout(w_dff_A_zjRwJyqb7_2),.din(w_dff_A_jtDD79jW1_2),.clk(gclk));
	jdff dff_A_sBkbIeom1_2(.dout(w_dff_A_jtDD79jW1_2),.din(w_dff_A_sBkbIeom1_2),.clk(gclk));
	jdff dff_A_X0kHbAdb7_2(.dout(w_dff_A_GuAOCVhn2_0),.din(w_dff_A_X0kHbAdb7_2),.clk(gclk));
	jdff dff_A_GuAOCVhn2_0(.dout(w_dff_A_LKlLEh6J0_0),.din(w_dff_A_GuAOCVhn2_0),.clk(gclk));
	jdff dff_A_LKlLEh6J0_0(.dout(w_dff_A_QY1HNHBJ4_0),.din(w_dff_A_LKlLEh6J0_0),.clk(gclk));
	jdff dff_A_QY1HNHBJ4_0(.dout(w_dff_A_aW2Db9OB6_0),.din(w_dff_A_QY1HNHBJ4_0),.clk(gclk));
	jdff dff_A_aW2Db9OB6_0(.dout(w_dff_A_ppDEx3IG8_0),.din(w_dff_A_aW2Db9OB6_0),.clk(gclk));
	jdff dff_A_ppDEx3IG8_0(.dout(w_dff_A_hBXJmn1q4_0),.din(w_dff_A_ppDEx3IG8_0),.clk(gclk));
	jdff dff_A_hBXJmn1q4_0(.dout(w_dff_A_FcZzibNF5_0),.din(w_dff_A_hBXJmn1q4_0),.clk(gclk));
	jdff dff_A_FcZzibNF5_0(.dout(w_dff_A_RjGobxKk6_0),.din(w_dff_A_FcZzibNF5_0),.clk(gclk));
	jdff dff_A_RjGobxKk6_0(.dout(w_dff_A_KLsQ9dIp4_0),.din(w_dff_A_RjGobxKk6_0),.clk(gclk));
	jdff dff_A_KLsQ9dIp4_0(.dout(w_dff_A_RvwfMsgN3_0),.din(w_dff_A_KLsQ9dIp4_0),.clk(gclk));
	jdff dff_A_RvwfMsgN3_0(.dout(w_dff_A_7tU4sIsA9_0),.din(w_dff_A_RvwfMsgN3_0),.clk(gclk));
	jdff dff_A_7tU4sIsA9_0(.dout(w_dff_A_aZ6oFDTS2_0),.din(w_dff_A_7tU4sIsA9_0),.clk(gclk));
	jdff dff_A_aZ6oFDTS2_0(.dout(w_dff_A_jrV05aOS6_0),.din(w_dff_A_aZ6oFDTS2_0),.clk(gclk));
	jdff dff_A_jrV05aOS6_0(.dout(w_dff_A_6q7s0qdu3_0),.din(w_dff_A_jrV05aOS6_0),.clk(gclk));
	jdff dff_A_6q7s0qdu3_0(.dout(w_dff_A_nkt1lD8z7_0),.din(w_dff_A_6q7s0qdu3_0),.clk(gclk));
	jdff dff_A_nkt1lD8z7_0(.dout(w_dff_A_eNFRzgiG5_0),.din(w_dff_A_nkt1lD8z7_0),.clk(gclk));
	jdff dff_A_eNFRzgiG5_0(.dout(w_dff_A_ITEFn8wP3_0),.din(w_dff_A_eNFRzgiG5_0),.clk(gclk));
	jdff dff_A_ITEFn8wP3_0(.dout(w_dff_A_7i9jumX77_0),.din(w_dff_A_ITEFn8wP3_0),.clk(gclk));
	jdff dff_A_7i9jumX77_0(.dout(G388gat),.din(w_dff_A_7i9jumX77_0),.clk(gclk));
	jdff dff_A_Y1nK9cE15_2(.dout(w_dff_A_pxVP3Bml5_0),.din(w_dff_A_Y1nK9cE15_2),.clk(gclk));
	jdff dff_A_pxVP3Bml5_0(.dout(w_dff_A_uS7IE3Xd3_0),.din(w_dff_A_pxVP3Bml5_0),.clk(gclk));
	jdff dff_A_uS7IE3Xd3_0(.dout(w_dff_A_xBieCWyF6_0),.din(w_dff_A_uS7IE3Xd3_0),.clk(gclk));
	jdff dff_A_xBieCWyF6_0(.dout(w_dff_A_vZnXxdw23_0),.din(w_dff_A_xBieCWyF6_0),.clk(gclk));
	jdff dff_A_vZnXxdw23_0(.dout(w_dff_A_DhjSzHIZ5_0),.din(w_dff_A_vZnXxdw23_0),.clk(gclk));
	jdff dff_A_DhjSzHIZ5_0(.dout(w_dff_A_q8JscRw53_0),.din(w_dff_A_DhjSzHIZ5_0),.clk(gclk));
	jdff dff_A_q8JscRw53_0(.dout(w_dff_A_HT3gbkfU4_0),.din(w_dff_A_q8JscRw53_0),.clk(gclk));
	jdff dff_A_HT3gbkfU4_0(.dout(w_dff_A_qXGm286t0_0),.din(w_dff_A_HT3gbkfU4_0),.clk(gclk));
	jdff dff_A_qXGm286t0_0(.dout(w_dff_A_jO4U8LkB2_0),.din(w_dff_A_qXGm286t0_0),.clk(gclk));
	jdff dff_A_jO4U8LkB2_0(.dout(w_dff_A_HIBjT0qA1_0),.din(w_dff_A_jO4U8LkB2_0),.clk(gclk));
	jdff dff_A_HIBjT0qA1_0(.dout(w_dff_A_BtI0d3MF4_0),.din(w_dff_A_HIBjT0qA1_0),.clk(gclk));
	jdff dff_A_BtI0d3MF4_0(.dout(w_dff_A_S9KIXEaX7_0),.din(w_dff_A_BtI0d3MF4_0),.clk(gclk));
	jdff dff_A_S9KIXEaX7_0(.dout(w_dff_A_rlDvStwN0_0),.din(w_dff_A_S9KIXEaX7_0),.clk(gclk));
	jdff dff_A_rlDvStwN0_0(.dout(w_dff_A_vUSHjRba9_0),.din(w_dff_A_rlDvStwN0_0),.clk(gclk));
	jdff dff_A_vUSHjRba9_0(.dout(w_dff_A_XySDXnhr5_0),.din(w_dff_A_vUSHjRba9_0),.clk(gclk));
	jdff dff_A_XySDXnhr5_0(.dout(w_dff_A_rchMZ7zR7_0),.din(w_dff_A_XySDXnhr5_0),.clk(gclk));
	jdff dff_A_rchMZ7zR7_0(.dout(w_dff_A_52z0K9tC3_0),.din(w_dff_A_rchMZ7zR7_0),.clk(gclk));
	jdff dff_A_52z0K9tC3_0(.dout(w_dff_A_8dNA4qOz6_0),.din(w_dff_A_52z0K9tC3_0),.clk(gclk));
	jdff dff_A_8dNA4qOz6_0(.dout(G389gat),.din(w_dff_A_8dNA4qOz6_0),.clk(gclk));
	jdff dff_A_ZXpPQbxW2_2(.dout(w_dff_A_OTiqX9dw5_0),.din(w_dff_A_ZXpPQbxW2_2),.clk(gclk));
	jdff dff_A_OTiqX9dw5_0(.dout(w_dff_A_pTDW5cen9_0),.din(w_dff_A_OTiqX9dw5_0),.clk(gclk));
	jdff dff_A_pTDW5cen9_0(.dout(w_dff_A_zhlrvFaz9_0),.din(w_dff_A_pTDW5cen9_0),.clk(gclk));
	jdff dff_A_zhlrvFaz9_0(.dout(w_dff_A_EKQQIoI42_0),.din(w_dff_A_zhlrvFaz9_0),.clk(gclk));
	jdff dff_A_EKQQIoI42_0(.dout(w_dff_A_p3CTsA2X3_0),.din(w_dff_A_EKQQIoI42_0),.clk(gclk));
	jdff dff_A_p3CTsA2X3_0(.dout(w_dff_A_0tBTn4xp7_0),.din(w_dff_A_p3CTsA2X3_0),.clk(gclk));
	jdff dff_A_0tBTn4xp7_0(.dout(w_dff_A_x4uE6wDa7_0),.din(w_dff_A_0tBTn4xp7_0),.clk(gclk));
	jdff dff_A_x4uE6wDa7_0(.dout(w_dff_A_188jnfxY0_0),.din(w_dff_A_x4uE6wDa7_0),.clk(gclk));
	jdff dff_A_188jnfxY0_0(.dout(w_dff_A_vfiaz7JC2_0),.din(w_dff_A_188jnfxY0_0),.clk(gclk));
	jdff dff_A_vfiaz7JC2_0(.dout(w_dff_A_0QEDlCjd3_0),.din(w_dff_A_vfiaz7JC2_0),.clk(gclk));
	jdff dff_A_0QEDlCjd3_0(.dout(w_dff_A_2CcnYQGP6_0),.din(w_dff_A_0QEDlCjd3_0),.clk(gclk));
	jdff dff_A_2CcnYQGP6_0(.dout(w_dff_A_M45ZyP6K8_0),.din(w_dff_A_2CcnYQGP6_0),.clk(gclk));
	jdff dff_A_M45ZyP6K8_0(.dout(w_dff_A_jy5KxXSS5_0),.din(w_dff_A_M45ZyP6K8_0),.clk(gclk));
	jdff dff_A_jy5KxXSS5_0(.dout(w_dff_A_AkCJCekU5_0),.din(w_dff_A_jy5KxXSS5_0),.clk(gclk));
	jdff dff_A_AkCJCekU5_0(.dout(w_dff_A_vhmXD8te8_0),.din(w_dff_A_AkCJCekU5_0),.clk(gclk));
	jdff dff_A_vhmXD8te8_0(.dout(w_dff_A_5ntqW6Wo7_0),.din(w_dff_A_vhmXD8te8_0),.clk(gclk));
	jdff dff_A_5ntqW6Wo7_0(.dout(w_dff_A_f6hGMEQq3_0),.din(w_dff_A_5ntqW6Wo7_0),.clk(gclk));
	jdff dff_A_f6hGMEQq3_0(.dout(w_dff_A_cJAURovK3_0),.din(w_dff_A_f6hGMEQq3_0),.clk(gclk));
	jdff dff_A_cJAURovK3_0(.dout(G390gat),.din(w_dff_A_cJAURovK3_0),.clk(gclk));
	jdff dff_A_SpizB91N3_2(.dout(w_dff_A_wFiDbO0J6_0),.din(w_dff_A_SpizB91N3_2),.clk(gclk));
	jdff dff_A_wFiDbO0J6_0(.dout(w_dff_A_k1Y13Y8V4_0),.din(w_dff_A_wFiDbO0J6_0),.clk(gclk));
	jdff dff_A_k1Y13Y8V4_0(.dout(w_dff_A_b1VoSuUE0_0),.din(w_dff_A_k1Y13Y8V4_0),.clk(gclk));
	jdff dff_A_b1VoSuUE0_0(.dout(w_dff_A_vWAO6IYk0_0),.din(w_dff_A_b1VoSuUE0_0),.clk(gclk));
	jdff dff_A_vWAO6IYk0_0(.dout(w_dff_A_1A2nlKG22_0),.din(w_dff_A_vWAO6IYk0_0),.clk(gclk));
	jdff dff_A_1A2nlKG22_0(.dout(w_dff_A_IicdvabJ4_0),.din(w_dff_A_1A2nlKG22_0),.clk(gclk));
	jdff dff_A_IicdvabJ4_0(.dout(w_dff_A_I8ekCjS71_0),.din(w_dff_A_IicdvabJ4_0),.clk(gclk));
	jdff dff_A_I8ekCjS71_0(.dout(w_dff_A_peuVB3pl6_0),.din(w_dff_A_I8ekCjS71_0),.clk(gclk));
	jdff dff_A_peuVB3pl6_0(.dout(w_dff_A_UlI71KH61_0),.din(w_dff_A_peuVB3pl6_0),.clk(gclk));
	jdff dff_A_UlI71KH61_0(.dout(w_dff_A_vauKkLvB3_0),.din(w_dff_A_UlI71KH61_0),.clk(gclk));
	jdff dff_A_vauKkLvB3_0(.dout(w_dff_A_gZPnn3N70_0),.din(w_dff_A_vauKkLvB3_0),.clk(gclk));
	jdff dff_A_gZPnn3N70_0(.dout(w_dff_A_RmHT7Dty3_0),.din(w_dff_A_gZPnn3N70_0),.clk(gclk));
	jdff dff_A_RmHT7Dty3_0(.dout(w_dff_A_zUP43K6b4_0),.din(w_dff_A_RmHT7Dty3_0),.clk(gclk));
	jdff dff_A_zUP43K6b4_0(.dout(w_dff_A_7iflffAH3_0),.din(w_dff_A_zUP43K6b4_0),.clk(gclk));
	jdff dff_A_7iflffAH3_0(.dout(w_dff_A_7qbnZ8U06_0),.din(w_dff_A_7iflffAH3_0),.clk(gclk));
	jdff dff_A_7qbnZ8U06_0(.dout(w_dff_A_8Soj1kAF1_0),.din(w_dff_A_7qbnZ8U06_0),.clk(gclk));
	jdff dff_A_8Soj1kAF1_0(.dout(w_dff_A_IZgVQmPA7_0),.din(w_dff_A_8Soj1kAF1_0),.clk(gclk));
	jdff dff_A_IZgVQmPA7_0(.dout(w_dff_A_jAQp9lAk2_0),.din(w_dff_A_IZgVQmPA7_0),.clk(gclk));
	jdff dff_A_jAQp9lAk2_0(.dout(w_dff_A_DTCDeFvN1_0),.din(w_dff_A_jAQp9lAk2_0),.clk(gclk));
	jdff dff_A_DTCDeFvN1_0(.dout(G391gat),.din(w_dff_A_DTCDeFvN1_0),.clk(gclk));
	jdff dff_A_DaA0Cm0b8_2(.dout(w_dff_A_kcvgynvC2_0),.din(w_dff_A_DaA0Cm0b8_2),.clk(gclk));
	jdff dff_A_kcvgynvC2_0(.dout(w_dff_A_pVzYYPWE4_0),.din(w_dff_A_kcvgynvC2_0),.clk(gclk));
	jdff dff_A_pVzYYPWE4_0(.dout(w_dff_A_udigj5878_0),.din(w_dff_A_pVzYYPWE4_0),.clk(gclk));
	jdff dff_A_udigj5878_0(.dout(w_dff_A_AmwrHkzk7_0),.din(w_dff_A_udigj5878_0),.clk(gclk));
	jdff dff_A_AmwrHkzk7_0(.dout(w_dff_A_CpqIqHEB8_0),.din(w_dff_A_AmwrHkzk7_0),.clk(gclk));
	jdff dff_A_CpqIqHEB8_0(.dout(w_dff_A_gOD43Cmg6_0),.din(w_dff_A_CpqIqHEB8_0),.clk(gclk));
	jdff dff_A_gOD43Cmg6_0(.dout(w_dff_A_THoY87Un0_0),.din(w_dff_A_gOD43Cmg6_0),.clk(gclk));
	jdff dff_A_THoY87Un0_0(.dout(w_dff_A_kxVaw1Yf9_0),.din(w_dff_A_THoY87Un0_0),.clk(gclk));
	jdff dff_A_kxVaw1Yf9_0(.dout(w_dff_A_X58358Id2_0),.din(w_dff_A_kxVaw1Yf9_0),.clk(gclk));
	jdff dff_A_X58358Id2_0(.dout(w_dff_A_321Hbrh97_0),.din(w_dff_A_X58358Id2_0),.clk(gclk));
	jdff dff_A_321Hbrh97_0(.dout(w_dff_A_GVXUdRe55_0),.din(w_dff_A_321Hbrh97_0),.clk(gclk));
	jdff dff_A_GVXUdRe55_0(.dout(w_dff_A_VCRxQNCe3_0),.din(w_dff_A_GVXUdRe55_0),.clk(gclk));
	jdff dff_A_VCRxQNCe3_0(.dout(w_dff_A_Vtr8G3At1_0),.din(w_dff_A_VCRxQNCe3_0),.clk(gclk));
	jdff dff_A_Vtr8G3At1_0(.dout(w_dff_A_b8SS2enS3_0),.din(w_dff_A_Vtr8G3At1_0),.clk(gclk));
	jdff dff_A_b8SS2enS3_0(.dout(w_dff_A_r9khn0Sj8_0),.din(w_dff_A_b8SS2enS3_0),.clk(gclk));
	jdff dff_A_r9khn0Sj8_0(.dout(w_dff_A_kK4gBzNY9_0),.din(w_dff_A_r9khn0Sj8_0),.clk(gclk));
	jdff dff_A_kK4gBzNY9_0(.dout(w_dff_A_gm97eV5i6_0),.din(w_dff_A_kK4gBzNY9_0),.clk(gclk));
	jdff dff_A_gm97eV5i6_0(.dout(w_dff_A_076S63OU4_0),.din(w_dff_A_gm97eV5i6_0),.clk(gclk));
	jdff dff_A_076S63OU4_0(.dout(G418gat),.din(w_dff_A_076S63OU4_0),.clk(gclk));
	jdff dff_A_Q7Y9z1ZK3_2(.dout(w_dff_A_HzPxqt1Z6_0),.din(w_dff_A_Q7Y9z1ZK3_2),.clk(gclk));
	jdff dff_A_HzPxqt1Z6_0(.dout(w_dff_A_U6M9yE166_0),.din(w_dff_A_HzPxqt1Z6_0),.clk(gclk));
	jdff dff_A_U6M9yE166_0(.dout(w_dff_A_YNdaR6bh9_0),.din(w_dff_A_U6M9yE166_0),.clk(gclk));
	jdff dff_A_YNdaR6bh9_0(.dout(w_dff_A_9Cy8yFQN2_0),.din(w_dff_A_YNdaR6bh9_0),.clk(gclk));
	jdff dff_A_9Cy8yFQN2_0(.dout(w_dff_A_dQvVwmBJ9_0),.din(w_dff_A_9Cy8yFQN2_0),.clk(gclk));
	jdff dff_A_dQvVwmBJ9_0(.dout(w_dff_A_K9H0oYzO8_0),.din(w_dff_A_dQvVwmBJ9_0),.clk(gclk));
	jdff dff_A_K9H0oYzO8_0(.dout(w_dff_A_XeIn005r7_0),.din(w_dff_A_K9H0oYzO8_0),.clk(gclk));
	jdff dff_A_XeIn005r7_0(.dout(w_dff_A_HRA0lOJY5_0),.din(w_dff_A_XeIn005r7_0),.clk(gclk));
	jdff dff_A_HRA0lOJY5_0(.dout(w_dff_A_ZnsDw7zE3_0),.din(w_dff_A_HRA0lOJY5_0),.clk(gclk));
	jdff dff_A_ZnsDw7zE3_0(.dout(w_dff_A_HVRVC1VK8_0),.din(w_dff_A_ZnsDw7zE3_0),.clk(gclk));
	jdff dff_A_HVRVC1VK8_0(.dout(w_dff_A_geW4UDfo4_0),.din(w_dff_A_HVRVC1VK8_0),.clk(gclk));
	jdff dff_A_geW4UDfo4_0(.dout(w_dff_A_BKRIBCOx6_0),.din(w_dff_A_geW4UDfo4_0),.clk(gclk));
	jdff dff_A_BKRIBCOx6_0(.dout(w_dff_A_7Tn18E0L6_0),.din(w_dff_A_BKRIBCOx6_0),.clk(gclk));
	jdff dff_A_7Tn18E0L6_0(.dout(w_dff_A_kHreSdkd2_0),.din(w_dff_A_7Tn18E0L6_0),.clk(gclk));
	jdff dff_A_kHreSdkd2_0(.dout(w_dff_A_lkLcpaEg1_0),.din(w_dff_A_kHreSdkd2_0),.clk(gclk));
	jdff dff_A_lkLcpaEg1_0(.dout(w_dff_A_uwCUJgbf2_0),.din(w_dff_A_lkLcpaEg1_0),.clk(gclk));
	jdff dff_A_uwCUJgbf2_0(.dout(G419gat),.din(w_dff_A_uwCUJgbf2_0),.clk(gclk));
	jdff dff_A_PC6qmYf30_2(.dout(w_dff_A_0FdV3wTW3_0),.din(w_dff_A_PC6qmYf30_2),.clk(gclk));
	jdff dff_A_0FdV3wTW3_0(.dout(w_dff_A_Z8nbjcKD3_0),.din(w_dff_A_0FdV3wTW3_0),.clk(gclk));
	jdff dff_A_Z8nbjcKD3_0(.dout(w_dff_A_z6pwVCWP5_0),.din(w_dff_A_Z8nbjcKD3_0),.clk(gclk));
	jdff dff_A_z6pwVCWP5_0(.dout(w_dff_A_2ZC5W0XD0_0),.din(w_dff_A_z6pwVCWP5_0),.clk(gclk));
	jdff dff_A_2ZC5W0XD0_0(.dout(w_dff_A_pDR1iKwO0_0),.din(w_dff_A_2ZC5W0XD0_0),.clk(gclk));
	jdff dff_A_pDR1iKwO0_0(.dout(w_dff_A_uxUs2PCY8_0),.din(w_dff_A_pDR1iKwO0_0),.clk(gclk));
	jdff dff_A_uxUs2PCY8_0(.dout(w_dff_A_8I4fbpua4_0),.din(w_dff_A_uxUs2PCY8_0),.clk(gclk));
	jdff dff_A_8I4fbpua4_0(.dout(w_dff_A_aTCXI97f2_0),.din(w_dff_A_8I4fbpua4_0),.clk(gclk));
	jdff dff_A_aTCXI97f2_0(.dout(w_dff_A_CR55BGBM5_0),.din(w_dff_A_aTCXI97f2_0),.clk(gclk));
	jdff dff_A_CR55BGBM5_0(.dout(w_dff_A_jSRamrSx0_0),.din(w_dff_A_CR55BGBM5_0),.clk(gclk));
	jdff dff_A_jSRamrSx0_0(.dout(w_dff_A_9hCgF8fD4_0),.din(w_dff_A_jSRamrSx0_0),.clk(gclk));
	jdff dff_A_9hCgF8fD4_0(.dout(w_dff_A_qML2Jkjc9_0),.din(w_dff_A_9hCgF8fD4_0),.clk(gclk));
	jdff dff_A_qML2Jkjc9_0(.dout(w_dff_A_TCjHZf5d7_0),.din(w_dff_A_qML2Jkjc9_0),.clk(gclk));
	jdff dff_A_TCjHZf5d7_0(.dout(w_dff_A_kanGzhW38_0),.din(w_dff_A_TCjHZf5d7_0),.clk(gclk));
	jdff dff_A_kanGzhW38_0(.dout(w_dff_A_GEWHvxaL8_0),.din(w_dff_A_kanGzhW38_0),.clk(gclk));
	jdff dff_A_GEWHvxaL8_0(.dout(w_dff_A_52Fa1Yns7_0),.din(w_dff_A_GEWHvxaL8_0),.clk(gclk));
	jdff dff_A_52Fa1Yns7_0(.dout(w_dff_A_rLmSjeJg4_0),.din(w_dff_A_52Fa1Yns7_0),.clk(gclk));
	jdff dff_A_rLmSjeJg4_0(.dout(G420gat),.din(w_dff_A_rLmSjeJg4_0),.clk(gclk));
	jdff dff_A_KVpRZNKx4_2(.dout(w_dff_A_Rhynn9945_0),.din(w_dff_A_KVpRZNKx4_2),.clk(gclk));
	jdff dff_A_Rhynn9945_0(.dout(w_dff_A_wigCtVz05_0),.din(w_dff_A_Rhynn9945_0),.clk(gclk));
	jdff dff_A_wigCtVz05_0(.dout(w_dff_A_YKYRJEAY4_0),.din(w_dff_A_wigCtVz05_0),.clk(gclk));
	jdff dff_A_YKYRJEAY4_0(.dout(w_dff_A_RYjya74O8_0),.din(w_dff_A_YKYRJEAY4_0),.clk(gclk));
	jdff dff_A_RYjya74O8_0(.dout(w_dff_A_1caixoAE3_0),.din(w_dff_A_RYjya74O8_0),.clk(gclk));
	jdff dff_A_1caixoAE3_0(.dout(w_dff_A_gDP94gmv7_0),.din(w_dff_A_1caixoAE3_0),.clk(gclk));
	jdff dff_A_gDP94gmv7_0(.dout(w_dff_A_rgVVfYiv7_0),.din(w_dff_A_gDP94gmv7_0),.clk(gclk));
	jdff dff_A_rgVVfYiv7_0(.dout(w_dff_A_d2BtERMW8_0),.din(w_dff_A_rgVVfYiv7_0),.clk(gclk));
	jdff dff_A_d2BtERMW8_0(.dout(w_dff_A_l7NK7DFj6_0),.din(w_dff_A_d2BtERMW8_0),.clk(gclk));
	jdff dff_A_l7NK7DFj6_0(.dout(w_dff_A_iMxUOqYy0_0),.din(w_dff_A_l7NK7DFj6_0),.clk(gclk));
	jdff dff_A_iMxUOqYy0_0(.dout(w_dff_A_Ocz9z1wh1_0),.din(w_dff_A_iMxUOqYy0_0),.clk(gclk));
	jdff dff_A_Ocz9z1wh1_0(.dout(w_dff_A_zj7HAygN9_0),.din(w_dff_A_Ocz9z1wh1_0),.clk(gclk));
	jdff dff_A_zj7HAygN9_0(.dout(w_dff_A_JBKPhhKh7_0),.din(w_dff_A_zj7HAygN9_0),.clk(gclk));
	jdff dff_A_JBKPhhKh7_0(.dout(w_dff_A_jEc1bim20_0),.din(w_dff_A_JBKPhhKh7_0),.clk(gclk));
	jdff dff_A_jEc1bim20_0(.dout(w_dff_A_BFp5owVO5_0),.din(w_dff_A_jEc1bim20_0),.clk(gclk));
	jdff dff_A_BFp5owVO5_0(.dout(w_dff_A_QNVKxMMM6_0),.din(w_dff_A_BFp5owVO5_0),.clk(gclk));
	jdff dff_A_QNVKxMMM6_0(.dout(w_dff_A_yg0VlKrA6_0),.din(w_dff_A_QNVKxMMM6_0),.clk(gclk));
	jdff dff_A_yg0VlKrA6_0(.dout(G421gat),.din(w_dff_A_yg0VlKrA6_0),.clk(gclk));
	jdff dff_A_e8sPWf7F8_2(.dout(w_dff_A_SI057U6r4_0),.din(w_dff_A_e8sPWf7F8_2),.clk(gclk));
	jdff dff_A_SI057U6r4_0(.dout(w_dff_A_nA3S8Bqt0_0),.din(w_dff_A_SI057U6r4_0),.clk(gclk));
	jdff dff_A_nA3S8Bqt0_0(.dout(w_dff_A_qdFba6oH0_0),.din(w_dff_A_nA3S8Bqt0_0),.clk(gclk));
	jdff dff_A_qdFba6oH0_0(.dout(w_dff_A_0kFxVnYG9_0),.din(w_dff_A_qdFba6oH0_0),.clk(gclk));
	jdff dff_A_0kFxVnYG9_0(.dout(w_dff_A_dePyAu5j6_0),.din(w_dff_A_0kFxVnYG9_0),.clk(gclk));
	jdff dff_A_dePyAu5j6_0(.dout(w_dff_A_0jL7wY0t2_0),.din(w_dff_A_dePyAu5j6_0),.clk(gclk));
	jdff dff_A_0jL7wY0t2_0(.dout(w_dff_A_WDyrjHUh8_0),.din(w_dff_A_0jL7wY0t2_0),.clk(gclk));
	jdff dff_A_WDyrjHUh8_0(.dout(w_dff_A_HQy7LTtE8_0),.din(w_dff_A_WDyrjHUh8_0),.clk(gclk));
	jdff dff_A_HQy7LTtE8_0(.dout(w_dff_A_drtiOR7H3_0),.din(w_dff_A_HQy7LTtE8_0),.clk(gclk));
	jdff dff_A_drtiOR7H3_0(.dout(w_dff_A_okes5AJ46_0),.din(w_dff_A_drtiOR7H3_0),.clk(gclk));
	jdff dff_A_okes5AJ46_0(.dout(w_dff_A_OLSXyivU0_0),.din(w_dff_A_okes5AJ46_0),.clk(gclk));
	jdff dff_A_OLSXyivU0_0(.dout(w_dff_A_zBpAOFK81_0),.din(w_dff_A_OLSXyivU0_0),.clk(gclk));
	jdff dff_A_zBpAOFK81_0(.dout(w_dff_A_xHrPpOCF5_0),.din(w_dff_A_zBpAOFK81_0),.clk(gclk));
	jdff dff_A_xHrPpOCF5_0(.dout(w_dff_A_mPN3NODv5_0),.din(w_dff_A_xHrPpOCF5_0),.clk(gclk));
	jdff dff_A_mPN3NODv5_0(.dout(w_dff_A_z7J8qGh39_0),.din(w_dff_A_mPN3NODv5_0),.clk(gclk));
	jdff dff_A_z7J8qGh39_0(.dout(w_dff_A_lmZZyiBz7_0),.din(w_dff_A_z7J8qGh39_0),.clk(gclk));
	jdff dff_A_lmZZyiBz7_0(.dout(w_dff_A_aprmP46e1_0),.din(w_dff_A_lmZZyiBz7_0),.clk(gclk));
	jdff dff_A_aprmP46e1_0(.dout(G422gat),.din(w_dff_A_aprmP46e1_0),.clk(gclk));
	jdff dff_A_398D8Blp3_2(.dout(w_dff_A_9xtsT3pm2_0),.din(w_dff_A_398D8Blp3_2),.clk(gclk));
	jdff dff_A_9xtsT3pm2_0(.dout(w_dff_A_2t4rJmJw5_0),.din(w_dff_A_9xtsT3pm2_0),.clk(gclk));
	jdff dff_A_2t4rJmJw5_0(.dout(w_dff_A_iBunZqcK2_0),.din(w_dff_A_2t4rJmJw5_0),.clk(gclk));
	jdff dff_A_iBunZqcK2_0(.dout(w_dff_A_IPn94Egd6_0),.din(w_dff_A_iBunZqcK2_0),.clk(gclk));
	jdff dff_A_IPn94Egd6_0(.dout(w_dff_A_EioGrX3Z4_0),.din(w_dff_A_IPn94Egd6_0),.clk(gclk));
	jdff dff_A_EioGrX3Z4_0(.dout(w_dff_A_4rqMQxgh1_0),.din(w_dff_A_EioGrX3Z4_0),.clk(gclk));
	jdff dff_A_4rqMQxgh1_0(.dout(w_dff_A_lsF9shlh8_0),.din(w_dff_A_4rqMQxgh1_0),.clk(gclk));
	jdff dff_A_lsF9shlh8_0(.dout(w_dff_A_Teh4GM4H0_0),.din(w_dff_A_lsF9shlh8_0),.clk(gclk));
	jdff dff_A_Teh4GM4H0_0(.dout(w_dff_A_Un5Z3Ob27_0),.din(w_dff_A_Teh4GM4H0_0),.clk(gclk));
	jdff dff_A_Un5Z3Ob27_0(.dout(w_dff_A_nCXLlWfk0_0),.din(w_dff_A_Un5Z3Ob27_0),.clk(gclk));
	jdff dff_A_nCXLlWfk0_0(.dout(w_dff_A_ascmzqmL6_0),.din(w_dff_A_nCXLlWfk0_0),.clk(gclk));
	jdff dff_A_ascmzqmL6_0(.dout(w_dff_A_PJrSBVSY8_0),.din(w_dff_A_ascmzqmL6_0),.clk(gclk));
	jdff dff_A_PJrSBVSY8_0(.dout(w_dff_A_zN488CAe4_0),.din(w_dff_A_PJrSBVSY8_0),.clk(gclk));
	jdff dff_A_zN488CAe4_0(.dout(w_dff_A_I7IoKrtQ2_0),.din(w_dff_A_zN488CAe4_0),.clk(gclk));
	jdff dff_A_I7IoKrtQ2_0(.dout(w_dff_A_SnGkx1gH4_0),.din(w_dff_A_I7IoKrtQ2_0),.clk(gclk));
	jdff dff_A_SnGkx1gH4_0(.dout(w_dff_A_KRmvczNF6_0),.din(w_dff_A_SnGkx1gH4_0),.clk(gclk));
	jdff dff_A_KRmvczNF6_0(.dout(w_dff_A_3qMyA9P25_0),.din(w_dff_A_KRmvczNF6_0),.clk(gclk));
	jdff dff_A_3qMyA9P25_0(.dout(w_dff_A_4EjUyHLf3_0),.din(w_dff_A_3qMyA9P25_0),.clk(gclk));
	jdff dff_A_4EjUyHLf3_0(.dout(G423gat),.din(w_dff_A_4EjUyHLf3_0),.clk(gclk));
	jdff dff_A_K9PJEWpm2_2(.dout(w_dff_A_OjT0IQyU4_0),.din(w_dff_A_K9PJEWpm2_2),.clk(gclk));
	jdff dff_A_OjT0IQyU4_0(.dout(w_dff_A_Wo8dyX5s4_0),.din(w_dff_A_OjT0IQyU4_0),.clk(gclk));
	jdff dff_A_Wo8dyX5s4_0(.dout(w_dff_A_QdI9JvV67_0),.din(w_dff_A_Wo8dyX5s4_0),.clk(gclk));
	jdff dff_A_QdI9JvV67_0(.dout(w_dff_A_F2VvoqcI3_0),.din(w_dff_A_QdI9JvV67_0),.clk(gclk));
	jdff dff_A_F2VvoqcI3_0(.dout(w_dff_A_LDyGWqCN4_0),.din(w_dff_A_F2VvoqcI3_0),.clk(gclk));
	jdff dff_A_LDyGWqCN4_0(.dout(w_dff_A_VqeBgFVJ2_0),.din(w_dff_A_LDyGWqCN4_0),.clk(gclk));
	jdff dff_A_VqeBgFVJ2_0(.dout(w_dff_A_9RROfpFx0_0),.din(w_dff_A_VqeBgFVJ2_0),.clk(gclk));
	jdff dff_A_9RROfpFx0_0(.dout(w_dff_A_7modmixP5_0),.din(w_dff_A_9RROfpFx0_0),.clk(gclk));
	jdff dff_A_7modmixP5_0(.dout(w_dff_A_6ngXizyP7_0),.din(w_dff_A_7modmixP5_0),.clk(gclk));
	jdff dff_A_6ngXizyP7_0(.dout(w_dff_A_SURhRANd5_0),.din(w_dff_A_6ngXizyP7_0),.clk(gclk));
	jdff dff_A_SURhRANd5_0(.dout(w_dff_A_J99FjoF71_0),.din(w_dff_A_SURhRANd5_0),.clk(gclk));
	jdff dff_A_J99FjoF71_0(.dout(w_dff_A_r3vJIeo42_0),.din(w_dff_A_J99FjoF71_0),.clk(gclk));
	jdff dff_A_r3vJIeo42_0(.dout(w_dff_A_GET4LZId2_0),.din(w_dff_A_r3vJIeo42_0),.clk(gclk));
	jdff dff_A_GET4LZId2_0(.dout(w_dff_A_1dCwUPHy5_0),.din(w_dff_A_GET4LZId2_0),.clk(gclk));
	jdff dff_A_1dCwUPHy5_0(.dout(w_dff_A_RUQd7QgF4_0),.din(w_dff_A_1dCwUPHy5_0),.clk(gclk));
	jdff dff_A_RUQd7QgF4_0(.dout(w_dff_A_XNxCifA49_0),.din(w_dff_A_RUQd7QgF4_0),.clk(gclk));
	jdff dff_A_XNxCifA49_0(.dout(G446gat),.din(w_dff_A_XNxCifA49_0),.clk(gclk));
	jdff dff_A_4aE1HHNH6_1(.dout(w_dff_A_I9x3h4qN1_0),.din(w_dff_A_4aE1HHNH6_1),.clk(gclk));
	jdff dff_A_I9x3h4qN1_0(.dout(w_dff_A_5ibh62iE0_0),.din(w_dff_A_I9x3h4qN1_0),.clk(gclk));
	jdff dff_A_5ibh62iE0_0(.dout(w_dff_A_1T43lxQM8_0),.din(w_dff_A_5ibh62iE0_0),.clk(gclk));
	jdff dff_A_1T43lxQM8_0(.dout(w_dff_A_dnb8rUiS2_0),.din(w_dff_A_1T43lxQM8_0),.clk(gclk));
	jdff dff_A_dnb8rUiS2_0(.dout(w_dff_A_WPd6hMJ60_0),.din(w_dff_A_dnb8rUiS2_0),.clk(gclk));
	jdff dff_A_WPd6hMJ60_0(.dout(w_dff_A_k2fvyJjP1_0),.din(w_dff_A_WPd6hMJ60_0),.clk(gclk));
	jdff dff_A_k2fvyJjP1_0(.dout(w_dff_A_WgwIgCm09_0),.din(w_dff_A_k2fvyJjP1_0),.clk(gclk));
	jdff dff_A_WgwIgCm09_0(.dout(w_dff_A_4RU2KqSQ4_0),.din(w_dff_A_WgwIgCm09_0),.clk(gclk));
	jdff dff_A_4RU2KqSQ4_0(.dout(w_dff_A_A9ztUOAT4_0),.din(w_dff_A_4RU2KqSQ4_0),.clk(gclk));
	jdff dff_A_A9ztUOAT4_0(.dout(w_dff_A_Cr7eBnNh4_0),.din(w_dff_A_A9ztUOAT4_0),.clk(gclk));
	jdff dff_A_Cr7eBnNh4_0(.dout(w_dff_A_wciQpmws5_0),.din(w_dff_A_Cr7eBnNh4_0),.clk(gclk));
	jdff dff_A_wciQpmws5_0(.dout(w_dff_A_peBbtvtG6_0),.din(w_dff_A_wciQpmws5_0),.clk(gclk));
	jdff dff_A_peBbtvtG6_0(.dout(w_dff_A_MSP2qFW88_0),.din(w_dff_A_peBbtvtG6_0),.clk(gclk));
	jdff dff_A_MSP2qFW88_0(.dout(w_dff_A_60hFFASs2_0),.din(w_dff_A_MSP2qFW88_0),.clk(gclk));
	jdff dff_A_60hFFASs2_0(.dout(w_dff_A_mvOK2W9h7_0),.din(w_dff_A_60hFFASs2_0),.clk(gclk));
	jdff dff_A_mvOK2W9h7_0(.dout(w_dff_A_EKKJA5do1_0),.din(w_dff_A_mvOK2W9h7_0),.clk(gclk));
	jdff dff_A_EKKJA5do1_0(.dout(w_dff_A_HGE1uK6W9_0),.din(w_dff_A_EKKJA5do1_0),.clk(gclk));
	jdff dff_A_HGE1uK6W9_0(.dout(w_dff_A_zmegFpcB2_0),.din(w_dff_A_HGE1uK6W9_0),.clk(gclk));
	jdff dff_A_zmegFpcB2_0(.dout(G447gat),.din(w_dff_A_zmegFpcB2_0),.clk(gclk));
	jdff dff_A_up1EhJML0_2(.dout(w_dff_A_IjVS0GVL5_0),.din(w_dff_A_up1EhJML0_2),.clk(gclk));
	jdff dff_A_IjVS0GVL5_0(.dout(w_dff_A_aHk1J1aU1_0),.din(w_dff_A_IjVS0GVL5_0),.clk(gclk));
	jdff dff_A_aHk1J1aU1_0(.dout(w_dff_A_yXgFXQGu6_0),.din(w_dff_A_aHk1J1aU1_0),.clk(gclk));
	jdff dff_A_yXgFXQGu6_0(.dout(w_dff_A_iwvqaTI53_0),.din(w_dff_A_yXgFXQGu6_0),.clk(gclk));
	jdff dff_A_iwvqaTI53_0(.dout(w_dff_A_xtUb4BHg8_0),.din(w_dff_A_iwvqaTI53_0),.clk(gclk));
	jdff dff_A_xtUb4BHg8_0(.dout(w_dff_A_w33NIjZJ6_0),.din(w_dff_A_xtUb4BHg8_0),.clk(gclk));
	jdff dff_A_w33NIjZJ6_0(.dout(w_dff_A_aafD2M4u7_0),.din(w_dff_A_w33NIjZJ6_0),.clk(gclk));
	jdff dff_A_aafD2M4u7_0(.dout(w_dff_A_UiTCakOA9_0),.din(w_dff_A_aafD2M4u7_0),.clk(gclk));
	jdff dff_A_UiTCakOA9_0(.dout(w_dff_A_7gVl9CFj9_0),.din(w_dff_A_UiTCakOA9_0),.clk(gclk));
	jdff dff_A_7gVl9CFj9_0(.dout(w_dff_A_5SSV1iub4_0),.din(w_dff_A_7gVl9CFj9_0),.clk(gclk));
	jdff dff_A_5SSV1iub4_0(.dout(w_dff_A_8LJkgOP54_0),.din(w_dff_A_5SSV1iub4_0),.clk(gclk));
	jdff dff_A_8LJkgOP54_0(.dout(w_dff_A_xgwledVq0_0),.din(w_dff_A_8LJkgOP54_0),.clk(gclk));
	jdff dff_A_xgwledVq0_0(.dout(w_dff_A_rck1oucl5_0),.din(w_dff_A_xgwledVq0_0),.clk(gclk));
	jdff dff_A_rck1oucl5_0(.dout(w_dff_A_XweZXmXJ1_0),.din(w_dff_A_rck1oucl5_0),.clk(gclk));
	jdff dff_A_XweZXmXJ1_0(.dout(w_dff_A_W3dLmgUe1_0),.din(w_dff_A_XweZXmXJ1_0),.clk(gclk));
	jdff dff_A_W3dLmgUe1_0(.dout(w_dff_A_MkRBpyr40_0),.din(w_dff_A_W3dLmgUe1_0),.clk(gclk));
	jdff dff_A_MkRBpyr40_0(.dout(w_dff_A_oaRMwzhY2_0),.din(w_dff_A_MkRBpyr40_0),.clk(gclk));
	jdff dff_A_oaRMwzhY2_0(.dout(G448gat),.din(w_dff_A_oaRMwzhY2_0),.clk(gclk));
	jdff dff_A_csl3aRhX5_2(.dout(w_dff_A_mkY1nLu22_0),.din(w_dff_A_csl3aRhX5_2),.clk(gclk));
	jdff dff_A_mkY1nLu22_0(.dout(w_dff_A_XPMuzRkf4_0),.din(w_dff_A_mkY1nLu22_0),.clk(gclk));
	jdff dff_A_XPMuzRkf4_0(.dout(w_dff_A_iySXuQF41_0),.din(w_dff_A_XPMuzRkf4_0),.clk(gclk));
	jdff dff_A_iySXuQF41_0(.dout(w_dff_A_1kUW6dBg2_0),.din(w_dff_A_iySXuQF41_0),.clk(gclk));
	jdff dff_A_1kUW6dBg2_0(.dout(w_dff_A_OjXFrgtr1_0),.din(w_dff_A_1kUW6dBg2_0),.clk(gclk));
	jdff dff_A_OjXFrgtr1_0(.dout(w_dff_A_864MDl3i8_0),.din(w_dff_A_OjXFrgtr1_0),.clk(gclk));
	jdff dff_A_864MDl3i8_0(.dout(w_dff_A_fEYCxMoo8_0),.din(w_dff_A_864MDl3i8_0),.clk(gclk));
	jdff dff_A_fEYCxMoo8_0(.dout(w_dff_A_dt74t9FM2_0),.din(w_dff_A_fEYCxMoo8_0),.clk(gclk));
	jdff dff_A_dt74t9FM2_0(.dout(w_dff_A_JeZJ3xhm8_0),.din(w_dff_A_dt74t9FM2_0),.clk(gclk));
	jdff dff_A_JeZJ3xhm8_0(.dout(w_dff_A_EfRRtaOF5_0),.din(w_dff_A_JeZJ3xhm8_0),.clk(gclk));
	jdff dff_A_EfRRtaOF5_0(.dout(w_dff_A_x9c69HAT5_0),.din(w_dff_A_EfRRtaOF5_0),.clk(gclk));
	jdff dff_A_x9c69HAT5_0(.dout(w_dff_A_5zFJQRLR1_0),.din(w_dff_A_x9c69HAT5_0),.clk(gclk));
	jdff dff_A_5zFJQRLR1_0(.dout(w_dff_A_UtEUmA5r4_0),.din(w_dff_A_5zFJQRLR1_0),.clk(gclk));
	jdff dff_A_UtEUmA5r4_0(.dout(w_dff_A_uVEAPLAS1_0),.din(w_dff_A_UtEUmA5r4_0),.clk(gclk));
	jdff dff_A_uVEAPLAS1_0(.dout(w_dff_A_niKJqv7r5_0),.din(w_dff_A_uVEAPLAS1_0),.clk(gclk));
	jdff dff_A_niKJqv7r5_0(.dout(w_dff_A_2NM1ELsb7_0),.din(w_dff_A_niKJqv7r5_0),.clk(gclk));
	jdff dff_A_2NM1ELsb7_0(.dout(w_dff_A_eRsuRZUc0_0),.din(w_dff_A_2NM1ELsb7_0),.clk(gclk));
	jdff dff_A_eRsuRZUc0_0(.dout(G449gat),.din(w_dff_A_eRsuRZUc0_0),.clk(gclk));
	jdff dff_A_CrUGfiSX7_2(.dout(w_dff_A_gQCgLpuQ3_0),.din(w_dff_A_CrUGfiSX7_2),.clk(gclk));
	jdff dff_A_gQCgLpuQ3_0(.dout(w_dff_A_wp5znw2A7_0),.din(w_dff_A_gQCgLpuQ3_0),.clk(gclk));
	jdff dff_A_wp5znw2A7_0(.dout(w_dff_A_00R8rm1m6_0),.din(w_dff_A_wp5znw2A7_0),.clk(gclk));
	jdff dff_A_00R8rm1m6_0(.dout(w_dff_A_TFxh5nxS0_0),.din(w_dff_A_00R8rm1m6_0),.clk(gclk));
	jdff dff_A_TFxh5nxS0_0(.dout(w_dff_A_IsILClwD4_0),.din(w_dff_A_TFxh5nxS0_0),.clk(gclk));
	jdff dff_A_IsILClwD4_0(.dout(w_dff_A_5HHzlktf9_0),.din(w_dff_A_IsILClwD4_0),.clk(gclk));
	jdff dff_A_5HHzlktf9_0(.dout(w_dff_A_0O1rlOkM9_0),.din(w_dff_A_5HHzlktf9_0),.clk(gclk));
	jdff dff_A_0O1rlOkM9_0(.dout(w_dff_A_1b1w5zwa7_0),.din(w_dff_A_0O1rlOkM9_0),.clk(gclk));
	jdff dff_A_1b1w5zwa7_0(.dout(w_dff_A_ZOeJBvtb0_0),.din(w_dff_A_1b1w5zwa7_0),.clk(gclk));
	jdff dff_A_ZOeJBvtb0_0(.dout(w_dff_A_kEVaACIG0_0),.din(w_dff_A_ZOeJBvtb0_0),.clk(gclk));
	jdff dff_A_kEVaACIG0_0(.dout(w_dff_A_nlOkYiMg2_0),.din(w_dff_A_kEVaACIG0_0),.clk(gclk));
	jdff dff_A_nlOkYiMg2_0(.dout(w_dff_A_oq6czHbW5_0),.din(w_dff_A_nlOkYiMg2_0),.clk(gclk));
	jdff dff_A_oq6czHbW5_0(.dout(w_dff_A_08gBmKcK0_0),.din(w_dff_A_oq6czHbW5_0),.clk(gclk));
	jdff dff_A_08gBmKcK0_0(.dout(w_dff_A_f5aOjsHf0_0),.din(w_dff_A_08gBmKcK0_0),.clk(gclk));
	jdff dff_A_f5aOjsHf0_0(.dout(w_dff_A_PHgt0RCM2_0),.din(w_dff_A_f5aOjsHf0_0),.clk(gclk));
	jdff dff_A_PHgt0RCM2_0(.dout(w_dff_A_nNZP1V5O0_0),.din(w_dff_A_PHgt0RCM2_0),.clk(gclk));
	jdff dff_A_nNZP1V5O0_0(.dout(w_dff_A_32HHgdDc0_0),.din(w_dff_A_nNZP1V5O0_0),.clk(gclk));
	jdff dff_A_32HHgdDc0_0(.dout(w_dff_A_svC8UNFs8_0),.din(w_dff_A_32HHgdDc0_0),.clk(gclk));
	jdff dff_A_svC8UNFs8_0(.dout(G450gat),.din(w_dff_A_svC8UNFs8_0),.clk(gclk));
	jdff dff_A_xsrmNVkq7_2(.dout(w_dff_A_uaor30g26_0),.din(w_dff_A_xsrmNVkq7_2),.clk(gclk));
	jdff dff_A_uaor30g26_0(.dout(w_dff_A_Im3bDWIN7_0),.din(w_dff_A_uaor30g26_0),.clk(gclk));
	jdff dff_A_Im3bDWIN7_0(.dout(w_dff_A_3G9WnZxV1_0),.din(w_dff_A_Im3bDWIN7_0),.clk(gclk));
	jdff dff_A_3G9WnZxV1_0(.dout(w_dff_A_JPLBFfI53_0),.din(w_dff_A_3G9WnZxV1_0),.clk(gclk));
	jdff dff_A_JPLBFfI53_0(.dout(w_dff_A_QflP8YtV6_0),.din(w_dff_A_JPLBFfI53_0),.clk(gclk));
	jdff dff_A_QflP8YtV6_0(.dout(w_dff_A_fbfY82HE3_0),.din(w_dff_A_QflP8YtV6_0),.clk(gclk));
	jdff dff_A_fbfY82HE3_0(.dout(w_dff_A_IlpauXBo3_0),.din(w_dff_A_fbfY82HE3_0),.clk(gclk));
	jdff dff_A_IlpauXBo3_0(.dout(w_dff_A_viuvkxgk6_0),.din(w_dff_A_IlpauXBo3_0),.clk(gclk));
	jdff dff_A_viuvkxgk6_0(.dout(w_dff_A_QVyTf5I20_0),.din(w_dff_A_viuvkxgk6_0),.clk(gclk));
	jdff dff_A_QVyTf5I20_0(.dout(w_dff_A_aMpIvDcO3_0),.din(w_dff_A_QVyTf5I20_0),.clk(gclk));
	jdff dff_A_aMpIvDcO3_0(.dout(w_dff_A_hV6sMuhr8_0),.din(w_dff_A_aMpIvDcO3_0),.clk(gclk));
	jdff dff_A_hV6sMuhr8_0(.dout(w_dff_A_20bCMobo8_0),.din(w_dff_A_hV6sMuhr8_0),.clk(gclk));
	jdff dff_A_20bCMobo8_0(.dout(w_dff_A_CugvgRr46_0),.din(w_dff_A_20bCMobo8_0),.clk(gclk));
	jdff dff_A_CugvgRr46_0(.dout(w_dff_A_sJmRVQDw9_0),.din(w_dff_A_CugvgRr46_0),.clk(gclk));
	jdff dff_A_sJmRVQDw9_0(.dout(w_dff_A_As6zZmd30_0),.din(w_dff_A_sJmRVQDw9_0),.clk(gclk));
	jdff dff_A_As6zZmd30_0(.dout(w_dff_A_0IlwTYZ81_0),.din(w_dff_A_As6zZmd30_0),.clk(gclk));
	jdff dff_A_0IlwTYZ81_0(.dout(G767gat),.din(w_dff_A_0IlwTYZ81_0),.clk(gclk));
	jdff dff_A_4vD5BJ2U0_2(.dout(w_dff_A_2Sfk8hZq5_0),.din(w_dff_A_4vD5BJ2U0_2),.clk(gclk));
	jdff dff_A_2Sfk8hZq5_0(.dout(w_dff_A_pWu2FU9w1_0),.din(w_dff_A_2Sfk8hZq5_0),.clk(gclk));
	jdff dff_A_pWu2FU9w1_0(.dout(w_dff_A_0eEcsSck5_0),.din(w_dff_A_pWu2FU9w1_0),.clk(gclk));
	jdff dff_A_0eEcsSck5_0(.dout(w_dff_A_DtIC18th4_0),.din(w_dff_A_0eEcsSck5_0),.clk(gclk));
	jdff dff_A_DtIC18th4_0(.dout(w_dff_A_6Pw5vc0f1_0),.din(w_dff_A_DtIC18th4_0),.clk(gclk));
	jdff dff_A_6Pw5vc0f1_0(.dout(w_dff_A_ZzdwRnFU3_0),.din(w_dff_A_6Pw5vc0f1_0),.clk(gclk));
	jdff dff_A_ZzdwRnFU3_0(.dout(w_dff_A_L6iLODd12_0),.din(w_dff_A_ZzdwRnFU3_0),.clk(gclk));
	jdff dff_A_L6iLODd12_0(.dout(w_dff_A_4MpTUQrL9_0),.din(w_dff_A_L6iLODd12_0),.clk(gclk));
	jdff dff_A_4MpTUQrL9_0(.dout(w_dff_A_1QrvILdF1_0),.din(w_dff_A_4MpTUQrL9_0),.clk(gclk));
	jdff dff_A_1QrvILdF1_0(.dout(w_dff_A_2SuZKbSr9_0),.din(w_dff_A_1QrvILdF1_0),.clk(gclk));
	jdff dff_A_2SuZKbSr9_0(.dout(w_dff_A_Hzkem6hU8_0),.din(w_dff_A_2SuZKbSr9_0),.clk(gclk));
	jdff dff_A_Hzkem6hU8_0(.dout(w_dff_A_qUN49Yui5_0),.din(w_dff_A_Hzkem6hU8_0),.clk(gclk));
	jdff dff_A_qUN49Yui5_0(.dout(w_dff_A_SC76EtqL9_0),.din(w_dff_A_qUN49Yui5_0),.clk(gclk));
	jdff dff_A_SC76EtqL9_0(.dout(w_dff_A_UEJG2x9F1_0),.din(w_dff_A_SC76EtqL9_0),.clk(gclk));
	jdff dff_A_UEJG2x9F1_0(.dout(w_dff_A_CUal9O1N1_0),.din(w_dff_A_UEJG2x9F1_0),.clk(gclk));
	jdff dff_A_CUal9O1N1_0(.dout(w_dff_A_ROsCN0oV9_0),.din(w_dff_A_CUal9O1N1_0),.clk(gclk));
	jdff dff_A_ROsCN0oV9_0(.dout(G768gat),.din(w_dff_A_ROsCN0oV9_0),.clk(gclk));
	jdff dff_A_7W4PhO7b3_2(.dout(w_dff_A_gX40HpxM5_0),.din(w_dff_A_7W4PhO7b3_2),.clk(gclk));
	jdff dff_A_gX40HpxM5_0(.dout(w_dff_A_aYieiXnk6_0),.din(w_dff_A_gX40HpxM5_0),.clk(gclk));
	jdff dff_A_aYieiXnk6_0(.dout(w_dff_A_J21VZuxz4_0),.din(w_dff_A_aYieiXnk6_0),.clk(gclk));
	jdff dff_A_J21VZuxz4_0(.dout(w_dff_A_YoqysCiO4_0),.din(w_dff_A_J21VZuxz4_0),.clk(gclk));
	jdff dff_A_YoqysCiO4_0(.dout(w_dff_A_ht8ABj3t4_0),.din(w_dff_A_YoqysCiO4_0),.clk(gclk));
	jdff dff_A_ht8ABj3t4_0(.dout(w_dff_A_SCKs2Omb9_0),.din(w_dff_A_ht8ABj3t4_0),.clk(gclk));
	jdff dff_A_SCKs2Omb9_0(.dout(w_dff_A_EGj3SVRD2_0),.din(w_dff_A_SCKs2Omb9_0),.clk(gclk));
	jdff dff_A_EGj3SVRD2_0(.dout(G850gat),.din(w_dff_A_EGj3SVRD2_0),.clk(gclk));
	jdff dff_A_mgcnRDmm4_2(.dout(w_dff_A_y1E9JOjN1_0),.din(w_dff_A_mgcnRDmm4_2),.clk(gclk));
	jdff dff_A_y1E9JOjN1_0(.dout(w_dff_A_utUMXrRq9_0),.din(w_dff_A_y1E9JOjN1_0),.clk(gclk));
	jdff dff_A_utUMXrRq9_0(.dout(w_dff_A_nO3QnoHq0_0),.din(w_dff_A_utUMXrRq9_0),.clk(gclk));
	jdff dff_A_nO3QnoHq0_0(.dout(G863gat),.din(w_dff_A_nO3QnoHq0_0),.clk(gclk));
	jdff dff_A_VWu5r75i1_2(.dout(w_dff_A_wq0l5bdW9_0),.din(w_dff_A_VWu5r75i1_2),.clk(gclk));
	jdff dff_A_wq0l5bdW9_0(.dout(w_dff_A_pTdiBhOH3_0),.din(w_dff_A_wq0l5bdW9_0),.clk(gclk));
	jdff dff_A_pTdiBhOH3_0(.dout(w_dff_A_j82oyDVy1_0),.din(w_dff_A_pTdiBhOH3_0),.clk(gclk));
	jdff dff_A_j82oyDVy1_0(.dout(G864gat),.din(w_dff_A_j82oyDVy1_0),.clk(gclk));
	jdff dff_A_yKfR0GGH1_2(.dout(w_dff_A_sworGvl53_0),.din(w_dff_A_yKfR0GGH1_2),.clk(gclk));
	jdff dff_A_sworGvl53_0(.dout(w_dff_A_cUuhVVoP3_0),.din(w_dff_A_sworGvl53_0),.clk(gclk));
	jdff dff_A_cUuhVVoP3_0(.dout(w_dff_A_z1oCuJhh8_0),.din(w_dff_A_cUuhVVoP3_0),.clk(gclk));
	jdff dff_A_z1oCuJhh8_0(.dout(w_dff_A_uqNWdzWx9_0),.din(w_dff_A_z1oCuJhh8_0),.clk(gclk));
	jdff dff_A_uqNWdzWx9_0(.dout(w_dff_A_NUrM0tWc5_0),.din(w_dff_A_uqNWdzWx9_0),.clk(gclk));
	jdff dff_A_NUrM0tWc5_0(.dout(G865gat),.din(w_dff_A_NUrM0tWc5_0),.clk(gclk));
	jdff dff_A_k24t8EOj8_2(.dout(w_dff_A_sr7IBH1k9_0),.din(w_dff_A_k24t8EOj8_2),.clk(gclk));
	jdff dff_A_sr7IBH1k9_0(.dout(G866gat),.din(w_dff_A_sr7IBH1k9_0),.clk(gclk));
	jdff dff_A_4uviTJyN4_2(.dout(w_dff_A_bCGK6ity0_0),.din(w_dff_A_4uviTJyN4_2),.clk(gclk));
	jdff dff_A_bCGK6ity0_0(.dout(G874gat),.din(w_dff_A_bCGK6ity0_0),.clk(gclk));
endmodule

