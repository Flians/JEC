/*
adder:
	jxor: 255
	jspl: 129
	jspl3: 254
	jcb: 254
	jdff: 32385
	jand: 255

Summary:
	jxor: 255
	jspl: 129
	jspl3: 254
	jcb: 254
	jdff: 32385
	jand: 255

The maximum logic level gap of any gate:
	adder: 127
*/

module adder(gclk, a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123, a124, a125, a126, a127, b0, b1, b2, b3, b4, b5, b6, b7, b8, b9, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b20, b21, b22, b23, b24, b25, b26, b27, b28, b29, b30, b31, b32, b33, b34, b35, b36, b37, b38, b39, b40, b41, b42, b43, b44, b45, b46, b47, b48, b49, b50, b51, b52, b53, b54, b55, b56, b57, b58, b59, b60, b61, b62, b63, b64, b65, b66, b67, b68, b69, b70, b71, b72, b73, b74, b75, b76, b77, b78, b79, b80, b81, b82, b83, b84, b85, b86, b87, b88, b89, b90, b91, b92, b93, b94, b95, b96, b97, b98, b99, b100, b101, b102, b103, b104, b105, b106, b107, b108, b109, b110, b111, b112, b113, b114, b115, b116, b117, b118, b119, b120, b121, b122, b123, b124, b125, b126, b127, f0, f1, f2, f3, f4, f5, f6, f7, f8, f9, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f20, f21, f22, f23, f24, f25, f26, f27, f28, f29, f30, f31, f32, f33, f34, f35, f36, f37, f38, f39, f40, f41, f42, f43, f44, f45, f46, f47, f48, f49, f50, f51, f52, f53, f54, f55, f56, f57, f58, f59, f60, f61, f62, f63, f64, f65, f66, f67, f68, f69, f70, f71, f72, f73, f74, f75, f76, f77, f78, f79, f80, f81, f82, f83, f84, f85, f86, f87, f88, f89, f90, f91, f92, f93, f94, f95, f96, f97, f98, f99, f100, f101, f102, f103, f104, f105, f106, f107, f108, f109, f110, f111, f112, f113, f114, f115, f116, f117, f118, f119, f120, f121, f122, f123, f124, f125, f126, f127, cOut);
	input gclk;
	input a0;
	input a1;
	input a2;
	input a3;
	input a4;
	input a5;
	input a6;
	input a7;
	input a8;
	input a9;
	input a10;
	input a11;
	input a12;
	input a13;
	input a14;
	input a15;
	input a16;
	input a17;
	input a18;
	input a19;
	input a20;
	input a21;
	input a22;
	input a23;
	input a24;
	input a25;
	input a26;
	input a27;
	input a28;
	input a29;
	input a30;
	input a31;
	input a32;
	input a33;
	input a34;
	input a35;
	input a36;
	input a37;
	input a38;
	input a39;
	input a40;
	input a41;
	input a42;
	input a43;
	input a44;
	input a45;
	input a46;
	input a47;
	input a48;
	input a49;
	input a50;
	input a51;
	input a52;
	input a53;
	input a54;
	input a55;
	input a56;
	input a57;
	input a58;
	input a59;
	input a60;
	input a61;
	input a62;
	input a63;
	input a64;
	input a65;
	input a66;
	input a67;
	input a68;
	input a69;
	input a70;
	input a71;
	input a72;
	input a73;
	input a74;
	input a75;
	input a76;
	input a77;
	input a78;
	input a79;
	input a80;
	input a81;
	input a82;
	input a83;
	input a84;
	input a85;
	input a86;
	input a87;
	input a88;
	input a89;
	input a90;
	input a91;
	input a92;
	input a93;
	input a94;
	input a95;
	input a96;
	input a97;
	input a98;
	input a99;
	input a100;
	input a101;
	input a102;
	input a103;
	input a104;
	input a105;
	input a106;
	input a107;
	input a108;
	input a109;
	input a110;
	input a111;
	input a112;
	input a113;
	input a114;
	input a115;
	input a116;
	input a117;
	input a118;
	input a119;
	input a120;
	input a121;
	input a122;
	input a123;
	input a124;
	input a125;
	input a126;
	input a127;
	input b0;
	input b1;
	input b2;
	input b3;
	input b4;
	input b5;
	input b6;
	input b7;
	input b8;
	input b9;
	input b10;
	input b11;
	input b12;
	input b13;
	input b14;
	input b15;
	input b16;
	input b17;
	input b18;
	input b19;
	input b20;
	input b21;
	input b22;
	input b23;
	input b24;
	input b25;
	input b26;
	input b27;
	input b28;
	input b29;
	input b30;
	input b31;
	input b32;
	input b33;
	input b34;
	input b35;
	input b36;
	input b37;
	input b38;
	input b39;
	input b40;
	input b41;
	input b42;
	input b43;
	input b44;
	input b45;
	input b46;
	input b47;
	input b48;
	input b49;
	input b50;
	input b51;
	input b52;
	input b53;
	input b54;
	input b55;
	input b56;
	input b57;
	input b58;
	input b59;
	input b60;
	input b61;
	input b62;
	input b63;
	input b64;
	input b65;
	input b66;
	input b67;
	input b68;
	input b69;
	input b70;
	input b71;
	input b72;
	input b73;
	input b74;
	input b75;
	input b76;
	input b77;
	input b78;
	input b79;
	input b80;
	input b81;
	input b82;
	input b83;
	input b84;
	input b85;
	input b86;
	input b87;
	input b88;
	input b89;
	input b90;
	input b91;
	input b92;
	input b93;
	input b94;
	input b95;
	input b96;
	input b97;
	input b98;
	input b99;
	input b100;
	input b101;
	input b102;
	input b103;
	input b104;
	input b105;
	input b106;
	input b107;
	input b108;
	input b109;
	input b110;
	input b111;
	input b112;
	input b113;
	input b114;
	input b115;
	input b116;
	input b117;
	input b118;
	input b119;
	input b120;
	input b121;
	input b122;
	input b123;
	input b124;
	input b125;
	input b126;
	input b127;
	output f0;
	output f1;
	output f2;
	output f3;
	output f4;
	output f5;
	output f6;
	output f7;
	output f8;
	output f9;
	output f10;
	output f11;
	output f12;
	output f13;
	output f14;
	output f15;
	output f16;
	output f17;
	output f18;
	output f19;
	output f20;
	output f21;
	output f22;
	output f23;
	output f24;
	output f25;
	output f26;
	output f27;
	output f28;
	output f29;
	output f30;
	output f31;
	output f32;
	output f33;
	output f34;
	output f35;
	output f36;
	output f37;
	output f38;
	output f39;
	output f40;
	output f41;
	output f42;
	output f43;
	output f44;
	output f45;
	output f46;
	output f47;
	output f48;
	output f49;
	output f50;
	output f51;
	output f52;
	output f53;
	output f54;
	output f55;
	output f56;
	output f57;
	output f58;
	output f59;
	output f60;
	output f61;
	output f62;
	output f63;
	output f64;
	output f65;
	output f66;
	output f67;
	output f68;
	output f69;
	output f70;
	output f71;
	output f72;
	output f73;
	output f74;
	output f75;
	output f76;
	output f77;
	output f78;
	output f79;
	output f80;
	output f81;
	output f82;
	output f83;
	output f84;
	output f85;
	output f86;
	output f87;
	output f88;
	output f89;
	output f90;
	output f91;
	output f92;
	output f93;
	output f94;
	output f95;
	output f96;
	output f97;
	output f98;
	output f99;
	output f100;
	output f101;
	output f102;
	output f103;
	output f104;
	output f105;
	output f106;
	output f107;
	output f108;
	output f109;
	output f110;
	output f111;
	output f112;
	output f113;
	output f114;
	output f115;
	output f116;
	output f117;
	output f118;
	output f119;
	output f120;
	output f121;
	output f122;
	output f123;
	output f124;
	output f125;
	output f126;
	output f127;
	output cOut;
	wire n387;
	wire n388;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1146;
	wire n1147;
	wire n1148;
	wire [1:0] w_a0_0;
	wire [2:0] w_a1_0;
	wire [2:0] w_a2_0;
	wire [2:0] w_a3_0;
	wire [2:0] w_a4_0;
	wire [2:0] w_a5_0;
	wire [2:0] w_a6_0;
	wire [2:0] w_a7_0;
	wire [2:0] w_a8_0;
	wire [2:0] w_a9_0;
	wire [2:0] w_a10_0;
	wire [2:0] w_a11_0;
	wire [2:0] w_a12_0;
	wire [2:0] w_a13_0;
	wire [2:0] w_a14_0;
	wire [2:0] w_a15_0;
	wire [2:0] w_a16_0;
	wire [2:0] w_a17_0;
	wire [2:0] w_a18_0;
	wire [2:0] w_a19_0;
	wire [2:0] w_a20_0;
	wire [2:0] w_a21_0;
	wire [2:0] w_a22_0;
	wire [2:0] w_a23_0;
	wire [2:0] w_a24_0;
	wire [2:0] w_a25_0;
	wire [2:0] w_a26_0;
	wire [2:0] w_a27_0;
	wire [2:0] w_a28_0;
	wire [2:0] w_a29_0;
	wire [2:0] w_a30_0;
	wire [2:0] w_a31_0;
	wire [2:0] w_a32_0;
	wire [2:0] w_a33_0;
	wire [2:0] w_a34_0;
	wire [2:0] w_a35_0;
	wire [2:0] w_a36_0;
	wire [2:0] w_a37_0;
	wire [2:0] w_a38_0;
	wire [2:0] w_a39_0;
	wire [2:0] w_a40_0;
	wire [2:0] w_a41_0;
	wire [2:0] w_a42_0;
	wire [2:0] w_a43_0;
	wire [2:0] w_a44_0;
	wire [2:0] w_a45_0;
	wire [2:0] w_a46_0;
	wire [2:0] w_a47_0;
	wire [2:0] w_a48_0;
	wire [2:0] w_a49_0;
	wire [2:0] w_a50_0;
	wire [2:0] w_a51_0;
	wire [2:0] w_a52_0;
	wire [2:0] w_a53_0;
	wire [2:0] w_a54_0;
	wire [2:0] w_a55_0;
	wire [2:0] w_a56_0;
	wire [2:0] w_a57_0;
	wire [2:0] w_a58_0;
	wire [2:0] w_a59_0;
	wire [2:0] w_a60_0;
	wire [2:0] w_a61_0;
	wire [2:0] w_a62_0;
	wire [2:0] w_a63_0;
	wire [2:0] w_a64_0;
	wire [2:0] w_a65_0;
	wire [2:0] w_a66_0;
	wire [2:0] w_a67_0;
	wire [2:0] w_a68_0;
	wire [2:0] w_a69_0;
	wire [2:0] w_a70_0;
	wire [2:0] w_a71_0;
	wire [2:0] w_a72_0;
	wire [2:0] w_a73_0;
	wire [2:0] w_a74_0;
	wire [2:0] w_a75_0;
	wire [2:0] w_a76_0;
	wire [2:0] w_a77_0;
	wire [2:0] w_a78_0;
	wire [2:0] w_a79_0;
	wire [2:0] w_a80_0;
	wire [2:0] w_a81_0;
	wire [2:0] w_a82_0;
	wire [2:0] w_a83_0;
	wire [2:0] w_a84_0;
	wire [2:0] w_a85_0;
	wire [2:0] w_a86_0;
	wire [2:0] w_a87_0;
	wire [2:0] w_a88_0;
	wire [2:0] w_a89_0;
	wire [2:0] w_a90_0;
	wire [2:0] w_a91_0;
	wire [2:0] w_a92_0;
	wire [2:0] w_a93_0;
	wire [2:0] w_a94_0;
	wire [2:0] w_a95_0;
	wire [2:0] w_a96_0;
	wire [2:0] w_a97_0;
	wire [2:0] w_a98_0;
	wire [2:0] w_a99_0;
	wire [2:0] w_a100_0;
	wire [2:0] w_a101_0;
	wire [2:0] w_a102_0;
	wire [2:0] w_a103_0;
	wire [2:0] w_a104_0;
	wire [2:0] w_a105_0;
	wire [2:0] w_a106_0;
	wire [2:0] w_a107_0;
	wire [2:0] w_a108_0;
	wire [2:0] w_a109_0;
	wire [2:0] w_a110_0;
	wire [2:0] w_a111_0;
	wire [2:0] w_a112_0;
	wire [2:0] w_a113_0;
	wire [2:0] w_a114_0;
	wire [2:0] w_a115_0;
	wire [2:0] w_a116_0;
	wire [2:0] w_a117_0;
	wire [2:0] w_a118_0;
	wire [2:0] w_a119_0;
	wire [2:0] w_a120_0;
	wire [2:0] w_a121_0;
	wire [2:0] w_a122_0;
	wire [2:0] w_a123_0;
	wire [2:0] w_a124_0;
	wire [2:0] w_a125_0;
	wire [2:0] w_a126_0;
	wire [2:0] w_a127_0;
	wire [1:0] w_b0_0;
	wire [2:0] w_b1_0;
	wire [2:0] w_b2_0;
	wire [2:0] w_b3_0;
	wire [2:0] w_b4_0;
	wire [2:0] w_b5_0;
	wire [2:0] w_b6_0;
	wire [2:0] w_b7_0;
	wire [2:0] w_b8_0;
	wire [2:0] w_b9_0;
	wire [2:0] w_b10_0;
	wire [2:0] w_b11_0;
	wire [2:0] w_b12_0;
	wire [2:0] w_b13_0;
	wire [2:0] w_b14_0;
	wire [2:0] w_b15_0;
	wire [2:0] w_b16_0;
	wire [2:0] w_b17_0;
	wire [2:0] w_b18_0;
	wire [2:0] w_b19_0;
	wire [2:0] w_b20_0;
	wire [2:0] w_b21_0;
	wire [2:0] w_b22_0;
	wire [2:0] w_b23_0;
	wire [2:0] w_b24_0;
	wire [2:0] w_b25_0;
	wire [2:0] w_b26_0;
	wire [2:0] w_b27_0;
	wire [2:0] w_b28_0;
	wire [2:0] w_b29_0;
	wire [2:0] w_b30_0;
	wire [2:0] w_b31_0;
	wire [2:0] w_b32_0;
	wire [2:0] w_b33_0;
	wire [2:0] w_b34_0;
	wire [2:0] w_b35_0;
	wire [2:0] w_b36_0;
	wire [2:0] w_b37_0;
	wire [2:0] w_b38_0;
	wire [2:0] w_b39_0;
	wire [2:0] w_b40_0;
	wire [2:0] w_b41_0;
	wire [2:0] w_b42_0;
	wire [2:0] w_b43_0;
	wire [2:0] w_b44_0;
	wire [2:0] w_b45_0;
	wire [2:0] w_b46_0;
	wire [2:0] w_b47_0;
	wire [2:0] w_b48_0;
	wire [2:0] w_b49_0;
	wire [2:0] w_b50_0;
	wire [2:0] w_b51_0;
	wire [2:0] w_b52_0;
	wire [2:0] w_b53_0;
	wire [2:0] w_b54_0;
	wire [2:0] w_b55_0;
	wire [2:0] w_b56_0;
	wire [2:0] w_b57_0;
	wire [2:0] w_b58_0;
	wire [2:0] w_b59_0;
	wire [2:0] w_b60_0;
	wire [2:0] w_b61_0;
	wire [2:0] w_b62_0;
	wire [2:0] w_b63_0;
	wire [2:0] w_b64_0;
	wire [2:0] w_b65_0;
	wire [2:0] w_b66_0;
	wire [2:0] w_b67_0;
	wire [2:0] w_b68_0;
	wire [2:0] w_b69_0;
	wire [2:0] w_b70_0;
	wire [2:0] w_b71_0;
	wire [2:0] w_b72_0;
	wire [2:0] w_b73_0;
	wire [2:0] w_b74_0;
	wire [2:0] w_b75_0;
	wire [2:0] w_b76_0;
	wire [2:0] w_b77_0;
	wire [2:0] w_b78_0;
	wire [2:0] w_b79_0;
	wire [2:0] w_b80_0;
	wire [2:0] w_b81_0;
	wire [2:0] w_b82_0;
	wire [2:0] w_b83_0;
	wire [2:0] w_b84_0;
	wire [2:0] w_b85_0;
	wire [2:0] w_b86_0;
	wire [2:0] w_b87_0;
	wire [2:0] w_b88_0;
	wire [2:0] w_b89_0;
	wire [2:0] w_b90_0;
	wire [2:0] w_b91_0;
	wire [2:0] w_b92_0;
	wire [2:0] w_b93_0;
	wire [2:0] w_b94_0;
	wire [2:0] w_b95_0;
	wire [2:0] w_b96_0;
	wire [2:0] w_b97_0;
	wire [2:0] w_b98_0;
	wire [2:0] w_b99_0;
	wire [2:0] w_b100_0;
	wire [2:0] w_b101_0;
	wire [2:0] w_b102_0;
	wire [2:0] w_b103_0;
	wire [2:0] w_b104_0;
	wire [2:0] w_b105_0;
	wire [2:0] w_b106_0;
	wire [2:0] w_b107_0;
	wire [2:0] w_b108_0;
	wire [2:0] w_b109_0;
	wire [2:0] w_b110_0;
	wire [2:0] w_b111_0;
	wire [2:0] w_b112_0;
	wire [2:0] w_b113_0;
	wire [2:0] w_b114_0;
	wire [2:0] w_b115_0;
	wire [2:0] w_b116_0;
	wire [2:0] w_b117_0;
	wire [2:0] w_b118_0;
	wire [2:0] w_b119_0;
	wire [2:0] w_b120_0;
	wire [2:0] w_b121_0;
	wire [2:0] w_b122_0;
	wire [2:0] w_b123_0;
	wire [2:0] w_b124_0;
	wire [2:0] w_b125_0;
	wire [2:0] w_b126_0;
	wire [2:0] w_b127_0;
	wire [1:0] w_n387_0;
	wire [1:0] w_n393_0;
	wire [1:0] w_n399_0;
	wire [1:0] w_n405_0;
	wire [1:0] w_n411_0;
	wire [1:0] w_n417_0;
	wire [1:0] w_n423_0;
	wire [1:0] w_n429_0;
	wire [1:0] w_n435_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n447_0;
	wire [1:0] w_n453_0;
	wire [1:0] w_n459_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n471_0;
	wire [1:0] w_n477_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n495_0;
	wire [1:0] w_n501_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n513_0;
	wire [1:0] w_n519_0;
	wire [1:0] w_n525_0;
	wire [1:0] w_n531_0;
	wire [1:0] w_n537_0;
	wire [1:0] w_n543_0;
	wire [1:0] w_n549_0;
	wire [1:0] w_n555_0;
	wire [1:0] w_n561_0;
	wire [1:0] w_n567_0;
	wire [1:0] w_n573_0;
	wire [1:0] w_n579_0;
	wire [1:0] w_n585_0;
	wire [1:0] w_n591_0;
	wire [1:0] w_n597_0;
	wire [1:0] w_n603_0;
	wire [1:0] w_n609_0;
	wire [1:0] w_n615_0;
	wire [1:0] w_n621_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n633_0;
	wire [1:0] w_n639_0;
	wire [1:0] w_n645_0;
	wire [1:0] w_n651_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n663_0;
	wire [1:0] w_n669_0;
	wire [1:0] w_n675_0;
	wire [1:0] w_n681_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n699_0;
	wire [1:0] w_n705_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n717_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n729_0;
	wire [1:0] w_n735_0;
	wire [1:0] w_n741_0;
	wire [1:0] w_n747_0;
	wire [1:0] w_n753_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n765_0;
	wire [1:0] w_n771_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n783_0;
	wire [1:0] w_n789_0;
	wire [1:0] w_n795_0;
	wire [1:0] w_n801_0;
	wire [1:0] w_n807_0;
	wire [1:0] w_n813_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n825_0;
	wire [1:0] w_n831_0;
	wire [1:0] w_n837_0;
	wire [1:0] w_n843_0;
	wire [1:0] w_n849_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n861_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n873_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n885_0;
	wire [1:0] w_n891_0;
	wire [1:0] w_n897_0;
	wire [1:0] w_n903_0;
	wire [1:0] w_n909_0;
	wire [1:0] w_n915_0;
	wire [1:0] w_n921_0;
	wire [1:0] w_n927_0;
	wire [1:0] w_n933_0;
	wire [1:0] w_n939_0;
	wire [1:0] w_n945_0;
	wire [1:0] w_n951_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n963_0;
	wire [1:0] w_n969_0;
	wire [1:0] w_n975_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n987_0;
	wire [1:0] w_n993_0;
	wire [1:0] w_n999_0;
	wire [1:0] w_n1005_0;
	wire [1:0] w_n1011_0;
	wire [1:0] w_n1017_0;
	wire [1:0] w_n1023_0;
	wire [1:0] w_n1029_0;
	wire [1:0] w_n1035_0;
	wire [1:0] w_n1041_0;
	wire [1:0] w_n1047_0;
	wire [1:0] w_n1053_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1065_0;
	wire [1:0] w_n1071_0;
	wire [1:0] w_n1077_0;
	wire [1:0] w_n1083_0;
	wire [1:0] w_n1089_0;
	wire [1:0] w_n1095_0;
	wire [1:0] w_n1101_0;
	wire [1:0] w_n1107_0;
	wire [1:0] w_n1113_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1125_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1137_0;
	wire [1:0] w_n1143_0;
	wire w_dff_B_y2pBBYfz5_0;
	wire w_dff_B_3J0ThVUc7_0;
	wire w_dff_B_S1pCGBH96_0;
	wire w_dff_B_mnbAlDI71_0;
	wire w_dff_B_NzAYujON5_0;
	wire w_dff_B_WlKsqUMj9_0;
	wire w_dff_B_Brc2L2JI6_0;
	wire w_dff_B_uhMTUALy6_0;
	wire w_dff_B_l3Z1Mo835_0;
	wire w_dff_B_Q6vqZJ6y8_0;
	wire w_dff_B_Vw0IBdke4_0;
	wire w_dff_B_VsIXMNjy6_0;
	wire w_dff_B_bSPwuxqp4_0;
	wire w_dff_B_s84U52Se8_0;
	wire w_dff_B_8jJ4BMCH1_0;
	wire w_dff_B_AEPIaLck4_0;
	wire w_dff_B_BPO87s3p9_0;
	wire w_dff_B_4zLuvkWy1_0;
	wire w_dff_B_Lyc0HPPJ1_0;
	wire w_dff_B_1hvRqtBe9_0;
	wire w_dff_B_7r08WE430_0;
	wire w_dff_B_xHIFgZia5_0;
	wire w_dff_B_ENitSJQy5_0;
	wire w_dff_B_HCc7mr6w4_0;
	wire w_dff_B_bd1c5jY57_0;
	wire w_dff_B_6C0ksYw72_0;
	wire w_dff_B_pgqcWTDx4_0;
	wire w_dff_B_i2DkyCua4_0;
	wire w_dff_B_mNcyzUcq1_0;
	wire w_dff_B_DbF5kOQi0_0;
	wire w_dff_B_DYOiTE2s7_0;
	wire w_dff_B_l0i7qBUN1_0;
	wire w_dff_B_FSyTsyEj6_0;
	wire w_dff_B_BR29qnUu8_0;
	wire w_dff_B_Qd56E6vg8_0;
	wire w_dff_B_xJonAAGK0_0;
	wire w_dff_B_BkDsgWbV3_0;
	wire w_dff_B_AnrW8w1J2_0;
	wire w_dff_B_b8mra9OC2_0;
	wire w_dff_B_AkNPTd1e7_0;
	wire w_dff_B_qhdODlqZ7_0;
	wire w_dff_B_Y5ecTrgg6_0;
	wire w_dff_B_VsdGWGmT1_0;
	wire w_dff_B_cXMlOdRu1_0;
	wire w_dff_B_KD70119c7_0;
	wire w_dff_B_SYcaX9bI7_0;
	wire w_dff_B_VgxfLs2T1_0;
	wire w_dff_B_X0F1zZE67_0;
	wire w_dff_B_cuC6wUPc7_0;
	wire w_dff_B_8191GAeV7_0;
	wire w_dff_B_YYa4o79w2_0;
	wire w_dff_B_GW7ply0u6_0;
	wire w_dff_B_8tl8GIG71_0;
	wire w_dff_B_u12WWdo53_0;
	wire w_dff_B_i8x4P8bS8_0;
	wire w_dff_B_TzFE9tjS7_0;
	wire w_dff_B_cU72aOqo1_0;
	wire w_dff_B_KZbuGsuV1_0;
	wire w_dff_B_LiAiLy0l0_0;
	wire w_dff_B_s5RweoEM8_0;
	wire w_dff_B_9v7STkiO0_0;
	wire w_dff_B_WmPJBbFW3_0;
	wire w_dff_B_lAaw1exA1_0;
	wire w_dff_B_DSniR09k7_0;
	wire w_dff_B_wsiOqmRM9_0;
	wire w_dff_B_bSj65Sek7_0;
	wire w_dff_B_utfAyrTF1_0;
	wire w_dff_B_TuXlM1jX9_0;
	wire w_dff_B_cLppZy5R6_0;
	wire w_dff_B_UuguPchZ9_0;
	wire w_dff_B_Nrl2Hk9v0_0;
	wire w_dff_B_mjt7gJjd2_0;
	wire w_dff_B_E3b75pyO2_0;
	wire w_dff_B_qoeeGdgd2_0;
	wire w_dff_B_sxe69lGc5_0;
	wire w_dff_B_2raBfihI9_0;
	wire w_dff_B_18la0t473_0;
	wire w_dff_B_YbutfiBd1_0;
	wire w_dff_B_6urZ322P0_0;
	wire w_dff_B_ShgIq1m37_0;
	wire w_dff_B_ETOlpfmb2_0;
	wire w_dff_B_CEUyN6ux6_0;
	wire w_dff_B_7C2MaevD6_0;
	wire w_dff_B_N6KhNZgu7_0;
	wire w_dff_B_pzJrvu0e1_0;
	wire w_dff_B_A6auZr8o3_0;
	wire w_dff_B_hBdeRio21_0;
	wire w_dff_B_TKSjOwA91_0;
	wire w_dff_B_ay9vxaw98_0;
	wire w_dff_B_13VDLqBe5_0;
	wire w_dff_B_yvhE8Xy08_0;
	wire w_dff_B_PTGcPJtE0_0;
	wire w_dff_B_JpC7cviR8_0;
	wire w_dff_B_H4c00HdU0_0;
	wire w_dff_B_upp86dzb0_0;
	wire w_dff_B_NDnEzvqu6_0;
	wire w_dff_B_RpVVfcSh6_0;
	wire w_dff_B_5jursZBQ8_0;
	wire w_dff_B_agPTNz1F6_0;
	wire w_dff_B_AvzbDx8H5_0;
	wire w_dff_B_014C95Vl8_0;
	wire w_dff_B_kJRmBb332_0;
	wire w_dff_B_tAQ3iZIB7_0;
	wire w_dff_B_cpH1PCxC9_0;
	wire w_dff_B_0CAb5BDY8_0;
	wire w_dff_B_CVnYksQq7_0;
	wire w_dff_B_LqmOP2qT4_0;
	wire w_dff_B_NgxMaCRH5_0;
	wire w_dff_B_gWx6oyEi2_0;
	wire w_dff_B_Mp1NdEXh5_0;
	wire w_dff_B_G9fjLTRe5_0;
	wire w_dff_B_axJqJbaM2_0;
	wire w_dff_B_IrnZEV9l1_0;
	wire w_dff_B_0mN764PL3_0;
	wire w_dff_B_SqhsNIcs4_0;
	wire w_dff_B_4OD9xZis8_0;
	wire w_dff_B_b0fr9tox6_0;
	wire w_dff_B_JxshsCdJ8_0;
	wire w_dff_B_qiG9o07C6_0;
	wire w_dff_B_M8i2g1ka6_0;
	wire w_dff_B_fV77TxYs1_0;
	wire w_dff_B_fksKxLpP4_0;
	wire w_dff_B_fCPoUfhW4_0;
	wire w_dff_B_pKQ0PvID3_0;
	wire w_dff_B_jk20wsIu8_0;
	wire w_dff_B_iGy5gPnm4_0;
	wire w_dff_B_ZRxQ7bzK9_0;
	wire w_dff_B_X5bNYZFd0_0;
	wire w_dff_B_VFOZkSK24_0;
	wire w_dff_B_QKU5NNEE8_0;
	wire w_dff_B_4ZHLJ0GC2_0;
	wire w_dff_B_H3qk8Ngk1_0;
	wire w_dff_B_sQQCfYEQ4_0;
	wire w_dff_B_JF1ZhYUE2_0;
	wire w_dff_B_F9X4gAYw8_0;
	wire w_dff_B_CPSxdA6Y0_0;
	wire w_dff_B_mMAUhrYt2_0;
	wire w_dff_B_2luq4joT1_0;
	wire w_dff_B_Pyt4EZZJ0_0;
	wire w_dff_B_Tt7ltl6B0_0;
	wire w_dff_B_eOOmDQhE2_0;
	wire w_dff_B_jEGVBdHU3_0;
	wire w_dff_B_sntaHEWZ2_0;
	wire w_dff_B_XXILh6AL2_0;
	wire w_dff_B_KwalMrsG6_0;
	wire w_dff_B_bp4Pi2yE2_0;
	wire w_dff_B_HfK1dh8X1_0;
	wire w_dff_B_zx6my8418_0;
	wire w_dff_B_4KOnpXUq5_0;
	wire w_dff_B_ZZOJ6x3S6_0;
	wire w_dff_B_vIxtPeBW1_0;
	wire w_dff_B_TRmgWZG88_0;
	wire w_dff_B_c7YZMJgL7_0;
	wire w_dff_B_6v93hQPr8_0;
	wire w_dff_B_4hKX96Vy7_0;
	wire w_dff_B_HHp5iX6Y7_0;
	wire w_dff_B_ESPc2d4a0_0;
	wire w_dff_B_fhX4SxUd6_0;
	wire w_dff_B_JPaywt4G5_0;
	wire w_dff_B_dvfpfhKU1_0;
	wire w_dff_B_jEeAVqY32_0;
	wire w_dff_B_cdEo1vsy4_0;
	wire w_dff_B_2wXLHRe55_0;
	wire w_dff_B_4Kc4XWH48_0;
	wire w_dff_B_nf5GK2AY6_0;
	wire w_dff_B_XnuqDCUM9_0;
	wire w_dff_B_xxgnqxpN8_0;
	wire w_dff_B_JbJSN1lV7_0;
	wire w_dff_B_RmSmdPOU2_0;
	wire w_dff_B_U67o42Lq5_0;
	wire w_dff_B_XC5aVfCd5_0;
	wire w_dff_B_G0S2GwZ09_0;
	wire w_dff_B_x62J4vje9_0;
	wire w_dff_B_SFRTN3Md5_0;
	wire w_dff_B_zkXuueZY3_0;
	wire w_dff_B_ogaTn6RF0_0;
	wire w_dff_B_E2Su59NV2_0;
	wire w_dff_B_fRq81AU46_0;
	wire w_dff_B_B8or83K73_0;
	wire w_dff_B_BQuR4S9t9_0;
	wire w_dff_B_dTVUfitb2_0;
	wire w_dff_B_eKoNYbty9_0;
	wire w_dff_B_jVgOMN7k5_0;
	wire w_dff_B_MVDz5b5o9_0;
	wire w_dff_B_R4DxsPjb8_0;
	wire w_dff_B_vDYeXq2q6_0;
	wire w_dff_B_R14b2tbL2_0;
	wire w_dff_B_SDeuqkeB9_0;
	wire w_dff_B_4GN11q8D0_0;
	wire w_dff_B_3Qs1UfWC8_0;
	wire w_dff_B_MnNDT1is2_0;
	wire w_dff_B_arKNd0oe8_0;
	wire w_dff_B_yF6uoUj18_0;
	wire w_dff_B_ncSfzHcb0_0;
	wire w_dff_B_NxB2xmNm4_0;
	wire w_dff_B_wW0WMAum1_0;
	wire w_dff_B_8bSlceo85_0;
	wire w_dff_B_VVBAFCbw6_0;
	wire w_dff_B_CfV4Qxud8_0;
	wire w_dff_B_ZUkx8TLO4_0;
	wire w_dff_B_8OWstOGa8_0;
	wire w_dff_B_mwc4vsM58_0;
	wire w_dff_B_LXCaRJJX6_0;
	wire w_dff_B_d9dzexGR9_0;
	wire w_dff_B_JSVYjlZ47_0;
	wire w_dff_B_8ttyBqZq6_0;
	wire w_dff_B_Ydoe6WSr2_0;
	wire w_dff_B_V3LACywI4_0;
	wire w_dff_B_fA6vTMAx9_0;
	wire w_dff_B_bBoBpv7g8_0;
	wire w_dff_B_kibI2Lsn7_0;
	wire w_dff_B_1i9E8opU8_0;
	wire w_dff_B_ZP0eLExa3_0;
	wire w_dff_B_69jMsuV44_0;
	wire w_dff_B_nGUovmCT4_0;
	wire w_dff_B_QO5EJtOg1_0;
	wire w_dff_B_C6xAknTs3_0;
	wire w_dff_B_UA952wVj9_0;
	wire w_dff_B_BB5baCUN0_0;
	wire w_dff_B_Vcl1IVhX3_0;
	wire w_dff_B_QyS5YQU86_0;
	wire w_dff_B_iZT3vNez4_0;
	wire w_dff_B_FmD0jpTl4_0;
	wire w_dff_B_4TmnnmTU3_0;
	wire w_dff_B_uI4p7ore3_0;
	wire w_dff_B_1sP5vJEI1_0;
	wire w_dff_B_4hDT4OW44_0;
	wire w_dff_B_DxtHLcJX3_0;
	wire w_dff_B_I3FRdpeY8_0;
	wire w_dff_B_LCjZqcA51_0;
	wire w_dff_B_3eiO5ewK6_0;
	wire w_dff_B_bZajaUav7_0;
	wire w_dff_B_2ywnCjrs2_0;
	wire w_dff_B_cakhkuZe6_0;
	wire w_dff_B_TxUsVKqT7_0;
	wire w_dff_B_nQWCc0GG1_0;
	wire w_dff_B_tjUf3Qkn1_0;
	wire w_dff_B_gl9iP9l19_0;
	wire w_dff_B_MZCl56Jb2_0;
	wire w_dff_B_XQG076hP3_0;
	wire w_dff_B_G7z5w1fs9_0;
	wire w_dff_B_EiYlgQFs2_0;
	wire w_dff_B_uqHn00Cu2_0;
	wire w_dff_B_KBlSjnf81_0;
	wire w_dff_B_qNnI4DkE3_0;
	wire w_dff_B_QTljKgdg2_0;
	wire w_dff_B_Gqcpt5RQ0_0;
	wire w_dff_B_Mt2LI6eB8_0;
	wire w_dff_B_RHnQ76dr0_0;
	wire w_dff_B_Gv1KoaIi9_0;
	wire w_dff_B_AxqivGkA1_0;
	wire w_dff_B_LEeGPhjq3_0;
	wire w_dff_B_tF6BKpIu3_0;
	wire w_dff_B_g4pazIHh5_0;
	wire w_dff_B_lpAuQVBB2_0;
	wire w_dff_B_ApCAiQzs9_0;
	wire w_dff_B_SpwoBTAt1_0;
	wire w_dff_B_U96RE8xy5_0;
	wire w_dff_B_eoBMukMa5_0;
	wire w_dff_B_4jXODQ3B9_0;
	wire w_dff_B_lZcoV0uk4_0;
	wire w_dff_B_OnmiEVf42_0;
	wire w_dff_B_UmPftrQi0_0;
	wire w_dff_B_lUONg07m6_0;
	wire w_dff_B_3y6SCpRw2_0;
	wire w_dff_B_zTvh3DqS2_0;
	wire w_dff_B_5ExXoyAL2_0;
	wire w_dff_B_jT9MDiMr0_0;
	wire w_dff_B_miyIiyMV2_0;
	wire w_dff_B_XvNxR3tj8_0;
	wire w_dff_B_i4DJRbcS1_0;
	wire w_dff_B_eDEzBdcY7_0;
	wire w_dff_B_oJonf9lR0_0;
	wire w_dff_B_9HpXUMLg0_0;
	wire w_dff_B_xCoyA7NO3_0;
	wire w_dff_B_IxLjw79f1_0;
	wire w_dff_B_4AYBlWCD3_0;
	wire w_dff_B_EVIdfRnr9_0;
	wire w_dff_B_M4gnDXts9_0;
	wire w_dff_B_iN37gDGy2_0;
	wire w_dff_B_9C8KmD8m6_0;
	wire w_dff_B_S5s5HRoI9_0;
	wire w_dff_B_jNAGm5og6_0;
	wire w_dff_B_VG20qrEr6_0;
	wire w_dff_B_EwOjsB8V3_0;
	wire w_dff_B_Zwux3rlQ9_0;
	wire w_dff_B_DbvO4vQO3_0;
	wire w_dff_B_xQjmoaY74_0;
	wire w_dff_B_6a5zADIs6_0;
	wire w_dff_B_k2Xd6nNb8_0;
	wire w_dff_B_ms8xh3EV8_0;
	wire w_dff_B_7kiHfSA64_0;
	wire w_dff_B_chBzimeL5_0;
	wire w_dff_B_mLe91Mmr8_0;
	wire w_dff_B_UeUg9eZ52_0;
	wire w_dff_B_wcqkNhM27_0;
	wire w_dff_B_81f8RSgK9_0;
	wire w_dff_B_4pW0pTNI6_0;
	wire w_dff_B_5IfrSx3F2_0;
	wire w_dff_B_poGlmfvO9_0;
	wire w_dff_B_PaeZgrzM0_0;
	wire w_dff_B_OEZ0XwQM3_0;
	wire w_dff_B_UvxWDdtn7_0;
	wire w_dff_B_0yzfU7hL0_0;
	wire w_dff_B_bkbGC4eG6_0;
	wire w_dff_B_3RIC7VLq9_0;
	wire w_dff_B_rksoprrK5_0;
	wire w_dff_B_ebRdoXBX5_0;
	wire w_dff_B_pKVnF7wr7_0;
	wire w_dff_B_tgSJ4YhL5_0;
	wire w_dff_B_tqmIASoO5_0;
	wire w_dff_B_1RIJh5oF4_0;
	wire w_dff_B_xAhqYGbf7_0;
	wire w_dff_B_0WEnK7gQ2_0;
	wire w_dff_B_BdA8GnSg2_0;
	wire w_dff_B_H8v9suBR8_0;
	wire w_dff_B_UriLMoYz8_0;
	wire w_dff_B_iL5oYczG6_0;
	wire w_dff_B_9HyMLtqN9_0;
	wire w_dff_B_GgaWNR6y0_0;
	wire w_dff_B_WE5q7h8v2_0;
	wire w_dff_B_6VKFKMrh4_0;
	wire w_dff_B_YKUCZU4c8_0;
	wire w_dff_B_DfmVt6Xm5_0;
	wire w_dff_B_aSGLFurX1_0;
	wire w_dff_B_RekwREfp2_0;
	wire w_dff_B_15CwFlLC1_0;
	wire w_dff_B_a8rEoPRG0_0;
	wire w_dff_B_vMYE1HsK1_0;
	wire w_dff_B_ovE2hrmu2_0;
	wire w_dff_B_4ZSnHJcP8_0;
	wire w_dff_B_zgD4yy7E3_0;
	wire w_dff_B_OYHF5RYQ2_0;
	wire w_dff_B_LLTdxF677_0;
	wire w_dff_B_eCj82QUd7_0;
	wire w_dff_B_DFtYZ7Vw7_0;
	wire w_dff_B_N6akSSGO5_0;
	wire w_dff_B_bGlP83Zj6_0;
	wire w_dff_B_XgB6zGjw4_0;
	wire w_dff_B_533bdWdP4_0;
	wire w_dff_B_GCW5oDqv4_0;
	wire w_dff_B_57lOSRw34_0;
	wire w_dff_B_CBBwr0FA9_0;
	wire w_dff_B_f1a1ZauG3_0;
	wire w_dff_B_ZpnRSzPu3_0;
	wire w_dff_B_7GqLJKET8_0;
	wire w_dff_B_HcuyY8As9_0;
	wire w_dff_B_vBhM5tQJ7_0;
	wire w_dff_B_uJBMCCFG4_0;
	wire w_dff_B_DbT98QkQ7_0;
	wire w_dff_B_0AYkSjrX9_0;
	wire w_dff_B_ZA1XkIpP0_0;
	wire w_dff_B_7Cg4vMHU1_0;
	wire w_dff_B_br3x518c5_0;
	wire w_dff_B_Go7xWMxR1_0;
	wire w_dff_B_sNH0JW9z6_0;
	wire w_dff_B_8moapIex2_0;
	wire w_dff_B_X3q3Tuf58_0;
	wire w_dff_B_uQpto6cv6_0;
	wire w_dff_B_QH7pv2fm3_0;
	wire w_dff_B_rudd1qJs9_0;
	wire w_dff_B_q9N0SUOT0_0;
	wire w_dff_B_c3kBIbUy9_0;
	wire w_dff_B_XWKrs8JL4_0;
	wire w_dff_B_XQAPy75b1_0;
	wire w_dff_B_3xRIeh9V5_0;
	wire w_dff_B_2CcKH1iZ1_0;
	wire w_dff_B_UFIj6DOr8_0;
	wire w_dff_B_ljBRYaAG6_0;
	wire w_dff_B_WShNyRcF1_0;
	wire w_dff_B_Ift2MArW2_0;
	wire w_dff_B_BnUgafsP1_0;
	wire w_dff_B_XqJZkZQq0_0;
	wire w_dff_B_8gmQCQmS9_0;
	wire w_dff_B_5C3W7TxS4_0;
	wire w_dff_B_74Scc9qY7_0;
	wire w_dff_B_mgwSIloA7_0;
	wire w_dff_B_bWpvlkFu0_0;
	wire w_dff_B_xk0VIGMy4_0;
	wire w_dff_B_OkRSIUZc4_0;
	wire w_dff_B_ZduKGcBM3_0;
	wire w_dff_B_A5WWflar5_0;
	wire w_dff_B_e1u8KWbN2_0;
	wire w_dff_B_Akd77nII6_0;
	wire w_dff_B_sci2xV2l0_0;
	wire w_dff_B_ArbpdaB97_0;
	wire w_dff_B_uZH9Vvxy2_0;
	wire w_dff_B_5thX7RJO0_0;
	wire w_dff_B_Ip28Qx8p6_0;
	wire w_dff_B_IBiIzxcM6_0;
	wire w_dff_B_p1vENyNf6_0;
	wire w_dff_B_e6e7Efdy7_0;
	wire w_dff_B_XgCxSUBy2_0;
	wire w_dff_B_4NoFRTwx4_0;
	wire w_dff_B_3QABQ9NP4_0;
	wire w_dff_B_vCI2geMr1_0;
	wire w_dff_B_gfbD7nhv5_0;
	wire w_dff_B_dqM3uZTx3_0;
	wire w_dff_B_tSAF1Htu7_0;
	wire w_dff_B_zdrtpEtz4_0;
	wire w_dff_B_gz9wlFdQ8_0;
	wire w_dff_B_zr26dsR85_0;
	wire w_dff_B_3xeDZl1F8_0;
	wire w_dff_B_UHpUPr7r5_0;
	wire w_dff_B_uaSvaVQI9_0;
	wire w_dff_B_OxgAFEkU9_0;
	wire w_dff_B_dkiH6k7t8_0;
	wire w_dff_B_z4Cbq2j73_0;
	wire w_dff_B_LPqaqJmf3_0;
	wire w_dff_B_GAEIV1Ke6_0;
	wire w_dff_B_ZBzNic8q8_0;
	wire w_dff_B_m43XMzew6_0;
	wire w_dff_B_6UDn0Zez6_0;
	wire w_dff_B_LCH7t6FF8_0;
	wire w_dff_B_PKAztZiL9_0;
	wire w_dff_B_IN3uvrr45_0;
	wire w_dff_B_zbrV0bNw3_0;
	wire w_dff_B_KO9pfjW92_0;
	wire w_dff_B_TTIbsp2K4_0;
	wire w_dff_B_72OJvSzO1_0;
	wire w_dff_B_54EoEQuC5_0;
	wire w_dff_B_lrZU6iDG3_0;
	wire w_dff_B_3GxWQUJx9_0;
	wire w_dff_B_0mxDNauX0_0;
	wire w_dff_B_OynKnJcY1_0;
	wire w_dff_B_uNe84uCH6_0;
	wire w_dff_B_Jho5xa795_0;
	wire w_dff_B_i7znTgNA4_0;
	wire w_dff_B_KhgyE6Vj7_0;
	wire w_dff_B_0zVq1WWZ9_0;
	wire w_dff_B_dZKk2RTS0_0;
	wire w_dff_B_n0Hq61xH4_0;
	wire w_dff_B_OOSrtPox1_0;
	wire w_dff_B_s93P21LQ8_0;
	wire w_dff_B_0NQGDTyH9_0;
	wire w_dff_B_CCeYgj5q7_0;
	wire w_dff_B_Gz5busOc2_0;
	wire w_dff_B_hMKQex3R8_0;
	wire w_dff_B_k4jQfFFP9_0;
	wire w_dff_B_A99Gj2sq0_0;
	wire w_dff_B_YrJgWPz39_0;
	wire w_dff_B_0hPskeWw2_0;
	wire w_dff_B_oN2xRZGe8_0;
	wire w_dff_B_ZXhiPTGj0_0;
	wire w_dff_B_aqCZpPbu3_0;
	wire w_dff_B_3KNPvgzG6_0;
	wire w_dff_B_tzFPXq6z6_0;
	wire w_dff_B_TYP5FPPc8_0;
	wire w_dff_B_vNHFGvCb7_0;
	wire w_dff_B_tnLjToGI0_0;
	wire w_dff_B_GowKRS1P7_0;
	wire w_dff_B_0Sxd84Kr2_0;
	wire w_dff_B_JJ5Bdcte9_0;
	wire w_dff_B_6OPNAG569_0;
	wire w_dff_B_DL50Llf17_0;
	wire w_dff_B_26ONQgce5_0;
	wire w_dff_B_hO1wFjem1_0;
	wire w_dff_B_uPgWI5GI7_0;
	wire w_dff_B_k9J5o1lq9_0;
	wire w_dff_B_NdhviSid4_0;
	wire w_dff_B_VuvCKVB06_0;
	wire w_dff_B_QoUC1qbN7_0;
	wire w_dff_B_wiC1SogH4_0;
	wire w_dff_B_rcaV8e814_0;
	wire w_dff_B_yCmWmTN77_0;
	wire w_dff_B_A1PhRP3d7_0;
	wire w_dff_B_4hgOkIVd0_0;
	wire w_dff_B_EVbbXczU0_0;
	wire w_dff_B_zQBLhk6e1_0;
	wire w_dff_B_083QX3LK8_0;
	wire w_dff_B_ApYemFwo3_0;
	wire w_dff_B_A8ANUUMb0_0;
	wire w_dff_B_Kme2bApf0_0;
	wire w_dff_B_s4c3ypYF6_0;
	wire w_dff_B_CsOBqpYH6_0;
	wire w_dff_B_2B8BQQnX5_0;
	wire w_dff_B_edRF8MSF4_0;
	wire w_dff_B_Qt58gf8K4_0;
	wire w_dff_B_aJnvWoRe3_0;
	wire w_dff_B_WgEnrC709_0;
	wire w_dff_B_MKaPkcfQ1_0;
	wire w_dff_B_7m3sKTyf9_0;
	wire w_dff_B_2abs3PCw6_0;
	wire w_dff_B_SJA6YXzi3_0;
	wire w_dff_B_pFTfDD0O2_0;
	wire w_dff_B_GOi7Ebvm7_0;
	wire w_dff_B_pFRLx8Ze0_0;
	wire w_dff_B_8TXVcxsV2_0;
	wire w_dff_B_NVZbxlKC0_0;
	wire w_dff_B_NmIm7Vs78_0;
	wire w_dff_B_gzUCBXVb7_0;
	wire w_dff_B_TYDZLs2Y9_0;
	wire w_dff_B_dbkJUWm80_0;
	wire w_dff_B_mLXkMxVF2_0;
	wire w_dff_B_h4lQj65l7_0;
	wire w_dff_B_FPJBFbiz2_0;
	wire w_dff_B_46awi8rt3_0;
	wire w_dff_B_YxVlzGpd7_0;
	wire w_dff_B_R1nitSyc6_0;
	wire w_dff_B_hqbYiICS9_0;
	wire w_dff_B_pg7DmpEf7_0;
	wire w_dff_B_pjKjhEQg4_0;
	wire w_dff_B_TVag2PWB0_0;
	wire w_dff_B_GnQcVHrg6_0;
	wire w_dff_B_tTV78Fti3_0;
	wire w_dff_B_gF7AmbBz8_0;
	wire w_dff_B_Z6KugE428_0;
	wire w_dff_B_JM0bsTRR3_0;
	wire w_dff_B_vBGMu0PG3_0;
	wire w_dff_B_6oNWWjBK6_0;
	wire w_dff_B_K4cteTvu4_0;
	wire w_dff_B_deVqox1S0_0;
	wire w_dff_B_HJ0VgJV42_0;
	wire w_dff_B_8vVQXlFI6_0;
	wire w_dff_B_j4zovaBD6_0;
	wire w_dff_B_jVByXBGy9_0;
	wire w_dff_B_axGXTgLD7_0;
	wire w_dff_B_WrhtyOD43_0;
	wire w_dff_B_ipdEi38z7_0;
	wire w_dff_B_FimWTP4Q8_0;
	wire w_dff_B_sB8PY9B63_0;
	wire w_dff_B_qmAnkWwJ9_0;
	wire w_dff_B_FLUg9zg23_0;
	wire w_dff_B_gsIXkc2A8_0;
	wire w_dff_B_PP7MsnfQ7_0;
	wire w_dff_B_grnNnAR75_0;
	wire w_dff_B_io49pKME4_0;
	wire w_dff_B_Qyetcsqv4_0;
	wire w_dff_B_6ACmcSqa9_0;
	wire w_dff_B_1MVci1aD8_0;
	wire w_dff_B_6wF6U1MK3_0;
	wire w_dff_B_ek9HuBVW9_0;
	wire w_dff_B_TG8No2tq9_0;
	wire w_dff_B_tLQdwva41_0;
	wire w_dff_B_vAlmn7XW9_0;
	wire w_dff_B_B1g3OnwJ8_0;
	wire w_dff_B_BpePRh142_0;
	wire w_dff_B_LIoqhgO00_0;
	wire w_dff_B_eRhkJaG89_0;
	wire w_dff_B_4dg2piZS6_0;
	wire w_dff_B_GLu4Oucg8_0;
	wire w_dff_B_jA4rHmDX3_0;
	wire w_dff_B_oCq0iOk96_0;
	wire w_dff_B_T9s7pZKK9_0;
	wire w_dff_B_4lrfvYUi3_0;
	wire w_dff_B_l30poSjP7_0;
	wire w_dff_B_M7lWWlfJ5_0;
	wire w_dff_B_BDK4HPd36_0;
	wire w_dff_B_3vTuy3Bk2_0;
	wire w_dff_B_OgM6eGew7_0;
	wire w_dff_B_5zcqJjUe4_0;
	wire w_dff_B_F9Dlndwv7_0;
	wire w_dff_B_yhUe41eF5_0;
	wire w_dff_B_TIbdHZ0n5_0;
	wire w_dff_B_pFCwMA4u9_0;
	wire w_dff_B_j67cCf9n0_0;
	wire w_dff_B_ZePjBeln3_0;
	wire w_dff_B_6lflNrwv4_0;
	wire w_dff_B_PxiUDOwK5_0;
	wire w_dff_B_2kvT58Jr3_0;
	wire w_dff_B_WbAXqjB88_0;
	wire w_dff_B_xAnXldkw5_0;
	wire w_dff_B_OWT8tJf08_0;
	wire w_dff_B_rGvlmkGX1_0;
	wire w_dff_B_coGLsrq49_0;
	wire w_dff_B_G9MmrI7b3_0;
	wire w_dff_B_S9MMtSVj8_0;
	wire w_dff_B_8tGXunFm6_0;
	wire w_dff_B_0A9VS7KY5_0;
	wire w_dff_B_rk3N94Bx3_0;
	wire w_dff_B_D8I1CfTd3_0;
	wire w_dff_B_7T9ullDj9_0;
	wire w_dff_B_Ek0OTX2n3_0;
	wire w_dff_B_HnEY1rzJ7_0;
	wire w_dff_B_Pioerm9g5_0;
	wire w_dff_B_3AUJECEi4_0;
	wire w_dff_B_2N4y2pWX4_0;
	wire w_dff_B_BA1I6UGy9_0;
	wire w_dff_B_F0uHJ1ep8_0;
	wire w_dff_B_42e3FdGp2_0;
	wire w_dff_B_0wKyjJXR3_0;
	wire w_dff_B_wyriGQ280_0;
	wire w_dff_B_7ZhPNr8I9_0;
	wire w_dff_B_v81X9vVW2_0;
	wire w_dff_B_oErTCF311_0;
	wire w_dff_B_VWYwBy3A1_0;
	wire w_dff_B_9zbAgTAq8_0;
	wire w_dff_B_aavi7VYB8_0;
	wire w_dff_B_4ufKLp5C0_0;
	wire w_dff_B_WYO79c0j5_0;
	wire w_dff_B_KvlHQr7L6_0;
	wire w_dff_B_UaQtGvqK4_0;
	wire w_dff_B_jkPkgNyK5_0;
	wire w_dff_B_iZCaN07y6_0;
	wire w_dff_B_tTqoaoGw3_0;
	wire w_dff_B_6CAW1Bi71_0;
	wire w_dff_B_EYQ4Ugbh9_0;
	wire w_dff_B_khqpYdj28_0;
	wire w_dff_B_BG4MiUsI7_0;
	wire w_dff_B_2ZdJIpg02_0;
	wire w_dff_B_LzvqDQab8_0;
	wire w_dff_B_bYQSosfp4_0;
	wire w_dff_B_vWFugr9c6_0;
	wire w_dff_B_cpzefdg00_0;
	wire w_dff_B_gTqNlWi62_0;
	wire w_dff_B_bAB7dH8h6_0;
	wire w_dff_B_tiKsYfsy3_0;
	wire w_dff_B_XwKEVTyN3_0;
	wire w_dff_B_lXZ4Dx5C8_0;
	wire w_dff_B_YxCaTOrB6_0;
	wire w_dff_B_5mJJ8JPY6_0;
	wire w_dff_B_FofErz5J6_0;
	wire w_dff_B_PguLnj7c1_0;
	wire w_dff_B_xTbGZsq29_0;
	wire w_dff_B_hsHJrtbC1_0;
	wire w_dff_B_uRsQPYt34_0;
	wire w_dff_B_sY4gQZYM2_0;
	wire w_dff_B_OGbwYld46_0;
	wire w_dff_B_qysdxons0_0;
	wire w_dff_B_6UlW1OEO3_0;
	wire w_dff_B_dXRCq7HD9_0;
	wire w_dff_B_TTTTHqOE9_0;
	wire w_dff_B_givM90s49_0;
	wire w_dff_B_1betfp328_0;
	wire w_dff_B_pJYiDME72_0;
	wire w_dff_B_noqs5PZE5_0;
	wire w_dff_B_SyUyvPfc1_0;
	wire w_dff_B_BaTwVzpv6_0;
	wire w_dff_B_9R7bTIZc0_0;
	wire w_dff_B_OVSEBGFt8_0;
	wire w_dff_B_lg7sDa4m3_0;
	wire w_dff_B_kIU5wzMk4_0;
	wire w_dff_B_oJ02hao28_0;
	wire w_dff_B_3s2YdROj7_0;
	wire w_dff_B_SCoeVMVN6_0;
	wire w_dff_B_cNZ24YRu3_0;
	wire w_dff_B_8ayMfOmq6_0;
	wire w_dff_B_hTGzDXm21_0;
	wire w_dff_B_DjEeqKiM9_0;
	wire w_dff_B_UbNdYlP46_0;
	wire w_dff_B_ryaiLADL4_0;
	wire w_dff_B_wocJxgUa1_0;
	wire w_dff_B_lZ6ownHW3_0;
	wire w_dff_B_zsLlWmoh9_0;
	wire w_dff_B_s6OFruit2_0;
	wire w_dff_B_jl4MHObG2_0;
	wire w_dff_B_lEiK5sDf6_0;
	wire w_dff_B_rleuJbWp1_0;
	wire w_dff_B_mT8kbtBw0_0;
	wire w_dff_B_xxSXxaR81_0;
	wire w_dff_B_sTanXs5T7_0;
	wire w_dff_B_D0J5w3ko0_0;
	wire w_dff_B_fTO4tuyx8_0;
	wire w_dff_B_sPbC4NKy2_0;
	wire w_dff_B_mUKvMdNk3_0;
	wire w_dff_B_5v9uNf036_0;
	wire w_dff_B_SUsZha0H6_0;
	wire w_dff_B_JNn35Cqb3_0;
	wire w_dff_B_govLfac43_0;
	wire w_dff_B_thHdjvLH8_0;
	wire w_dff_B_QvoA4r4r0_0;
	wire w_dff_B_e9IJL2vo2_0;
	wire w_dff_B_tNjfnhvM2_0;
	wire w_dff_B_zRB7IH6H0_0;
	wire w_dff_B_tXzk3lcN6_0;
	wire w_dff_B_hF6XnBIn6_0;
	wire w_dff_B_s6AOjeQ90_0;
	wire w_dff_B_L6wTZ6vD3_0;
	wire w_dff_B_QB9kMdMO7_0;
	wire w_dff_B_D3DqKLpZ9_0;
	wire w_dff_B_DUjdZrWQ9_0;
	wire w_dff_B_Q97YAQfT5_0;
	wire w_dff_B_ZS2tzXnP3_0;
	wire w_dff_B_SrYogtzg3_0;
	wire w_dff_B_pu9WYaR28_0;
	wire w_dff_B_z5QIV03e6_0;
	wire w_dff_B_U2tAN3m88_0;
	wire w_dff_B_3cS8tSB59_0;
	wire w_dff_B_ZxrXRBFu6_0;
	wire w_dff_B_7OInyd9t9_0;
	wire w_dff_B_GB4uq2sc2_0;
	wire w_dff_B_fnlH7jW21_0;
	wire w_dff_B_15OWADbF9_0;
	wire w_dff_B_g6s6WTRR0_0;
	wire w_dff_B_Qpf4OHly7_0;
	wire w_dff_B_CBdxbGoT2_0;
	wire w_dff_B_SBBc6YiC2_0;
	wire w_dff_B_fspb4EEp6_0;
	wire w_dff_B_iF5fgSvz1_0;
	wire w_dff_B_hs8zCiMD3_0;
	wire w_dff_B_HWWyhlvB1_0;
	wire w_dff_B_uc7qRFTA6_0;
	wire w_dff_B_k51Cr8G75_0;
	wire w_dff_B_xdCbxJwm1_0;
	wire w_dff_B_jWgQXuk67_0;
	wire w_dff_B_Y9NiFqeR8_0;
	wire w_dff_B_ZX8Ch3cj2_0;
	wire w_dff_B_KVHv0EiF7_0;
	wire w_dff_B_5g9D2yef7_0;
	wire w_dff_B_2UrH3rDD2_0;
	wire w_dff_B_rLtt4ApS1_0;
	wire w_dff_B_NHVH94YY0_0;
	wire w_dff_B_oTtWTlv49_0;
	wire w_dff_B_AYUTfkV56_0;
	wire w_dff_B_Jeqwa2rS2_0;
	wire w_dff_B_CmIIuVXd6_0;
	wire w_dff_B_qeBOZr342_0;
	wire w_dff_B_Cd4D5MsJ2_0;
	wire w_dff_B_iVKCevZj5_0;
	wire w_dff_B_40uHNE919_0;
	wire w_dff_B_vV7nwnsO8_0;
	wire w_dff_B_Bz1hKt9d8_0;
	wire w_dff_B_Lm9wk6Sc7_0;
	wire w_dff_B_4UU4N0og3_0;
	wire w_dff_B_xPZc4aF72_0;
	wire w_dff_B_uU69aT6S2_0;
	wire w_dff_B_e1LkrerN2_0;
	wire w_dff_B_0e0BqBiA0_0;
	wire w_dff_B_ax8tszjc8_0;
	wire w_dff_B_7tedKxfT2_0;
	wire w_dff_B_lhocc6gV7_0;
	wire w_dff_B_ufiuSoxG5_0;
	wire w_dff_B_lWQBwcZ00_0;
	wire w_dff_B_grNQbOGn0_0;
	wire w_dff_B_5OclPB0N7_0;
	wire w_dff_B_LSF7P0BU3_0;
	wire w_dff_B_W9ILXsuc8_0;
	wire w_dff_B_fdtXQixB2_0;
	wire w_dff_B_C0i8xH2k6_0;
	wire w_dff_B_C8IoAg1S2_0;
	wire w_dff_B_k0MTLwlW2_0;
	wire w_dff_B_Q3Cc1CiC7_0;
	wire w_dff_B_RyGgbFbM5_0;
	wire w_dff_B_qH2NRSqL8_0;
	wire w_dff_B_rAsMQhCl6_0;
	wire w_dff_B_BioZhb744_0;
	wire w_dff_B_teMkegph3_0;
	wire w_dff_B_adBxIslw7_0;
	wire w_dff_B_qD5TNK5w8_0;
	wire w_dff_B_6kPievLc6_0;
	wire w_dff_B_KlorpDbQ7_0;
	wire w_dff_B_XM4Wf54a0_0;
	wire w_dff_B_9S0qzORT2_0;
	wire w_dff_B_bxMgh0PH8_0;
	wire w_dff_B_PpbC8LTR0_0;
	wire w_dff_B_nBIJ4Egf1_0;
	wire w_dff_B_x49YZXhk0_0;
	wire w_dff_B_Vrk1oO4i9_0;
	wire w_dff_B_ZQ5NontA8_0;
	wire w_dff_B_8bGwQLNC7_0;
	wire w_dff_B_KlX3xzeC0_0;
	wire w_dff_B_Y76ycSQN8_0;
	wire w_dff_B_Ju8ucWYV8_0;
	wire w_dff_B_6ydS0C4u0_0;
	wire w_dff_B_FccqzLpO7_0;
	wire w_dff_B_ksDi6erO7_0;
	wire w_dff_B_AoPXskoG4_0;
	wire w_dff_B_LzZ7765N4_0;
	wire w_dff_B_19oxLLtM3_0;
	wire w_dff_B_SRRDBq9q4_0;
	wire w_dff_B_FMq2Bf1y1_0;
	wire w_dff_B_HUPcZtHT3_0;
	wire w_dff_B_21cZmwcf1_0;
	wire w_dff_B_G0Fah0Il8_0;
	wire w_dff_B_CeLIn9j27_0;
	wire w_dff_B_uCccFr792_0;
	wire w_dff_B_mecpBe8W0_0;
	wire w_dff_B_p6ieCHgl2_0;
	wire w_dff_B_2iccKVI69_0;
	wire w_dff_B_EHGcNkNL6_0;
	wire w_dff_B_FzDe7gxx2_0;
	wire w_dff_B_zYDVsHBR5_0;
	wire w_dff_B_K1QIor8x8_0;
	wire w_dff_B_U6bqcODq5_0;
	wire w_dff_B_YD1IGiht4_0;
	wire w_dff_B_bCQHAXsL2_0;
	wire w_dff_B_gQ14AX0l4_0;
	wire w_dff_B_oaSy403U7_0;
	wire w_dff_B_d7hK51g43_0;
	wire w_dff_B_eIHhFn8J8_0;
	wire w_dff_B_uzwh64ZQ1_0;
	wire w_dff_B_P26dG0r79_0;
	wire w_dff_B_YrIPbXsZ4_0;
	wire w_dff_B_xp16meGh1_0;
	wire w_dff_B_g0c7eyZI8_0;
	wire w_dff_B_lWtXOHqv1_0;
	wire w_dff_B_a2r6yoBS5_0;
	wire w_dff_B_0SgxtVVo5_0;
	wire w_dff_B_4f0Wic170_0;
	wire w_dff_B_GZ6Jq6qm9_0;
	wire w_dff_B_gsRdRIWq7_0;
	wire w_dff_B_XNNavWuD4_0;
	wire w_dff_B_XT8e6qB99_0;
	wire w_dff_B_eePq8pFt3_0;
	wire w_dff_B_SUABLWS71_0;
	wire w_dff_B_8BTAbnth5_0;
	wire w_dff_B_Ut2sz3us0_0;
	wire w_dff_B_Plic3a3j8_0;
	wire w_dff_B_MZEnoUNH3_0;
	wire w_dff_B_DTCGJKIN6_0;
	wire w_dff_B_K5u2vD9v1_0;
	wire w_dff_B_g3h6yE2P4_0;
	wire w_dff_B_sK0uWiil3_0;
	wire w_dff_B_kpCK9AYw5_0;
	wire w_dff_B_fKajguko2_0;
	wire w_dff_B_JHbXgzf36_0;
	wire w_dff_B_9DzzZAaj7_0;
	wire w_dff_B_WnC1ZTp31_0;
	wire w_dff_B_NTeej0HV4_0;
	wire w_dff_B_OoHRG8iE5_0;
	wire w_dff_B_fwQc2M8m5_0;
	wire w_dff_B_NKGDZyvl6_0;
	wire w_dff_B_7j9CpVE68_0;
	wire w_dff_B_f9MTalO10_0;
	wire w_dff_B_bdZ8XQ5Z6_0;
	wire w_dff_B_5Y14gjS09_0;
	wire w_dff_B_6Hws304o8_0;
	wire w_dff_B_Y0kU99sb4_0;
	wire w_dff_B_MCBIitm02_0;
	wire w_dff_B_HBMFIay39_0;
	wire w_dff_B_0shDgtgi6_0;
	wire w_dff_B_OwZF7A2q1_0;
	wire w_dff_B_Njp67Q9q1_0;
	wire w_dff_B_knggDeZI2_0;
	wire w_dff_B_bijPdv523_0;
	wire w_dff_B_lM6JNNjH4_0;
	wire w_dff_B_2zNi7IL35_0;
	wire w_dff_B_scuPywgt9_0;
	wire w_dff_B_hIgJRwBa4_0;
	wire w_dff_B_h2i7UkD71_0;
	wire w_dff_B_FhvbVRyo4_0;
	wire w_dff_B_XHuxvklI3_0;
	wire w_dff_B_G0qV8B3v2_0;
	wire w_dff_B_5cLs7z8c3_0;
	wire w_dff_B_NtOV4SLt6_0;
	wire w_dff_B_uryy4H9k8_0;
	wire w_dff_B_Au9BNQV14_0;
	wire w_dff_B_WfQJyuZA1_0;
	wire w_dff_B_jzsr3Afh1_0;
	wire w_dff_B_xwakBVa87_0;
	wire w_dff_B_8FeW9SoK2_0;
	wire w_dff_B_BOjsym2A9_0;
	wire w_dff_B_HcHVv9Zk6_0;
	wire w_dff_B_sRlJnjoU3_0;
	wire w_dff_B_dARBkwhE0_0;
	wire w_dff_B_u092cIuI7_0;
	wire w_dff_B_WznS65yE5_0;
	wire w_dff_B_K1bWBl5p3_0;
	wire w_dff_B_kw6iMMN12_0;
	wire w_dff_B_dZxlWiiz8_0;
	wire w_dff_B_Gq1zhtW23_0;
	wire w_dff_B_2dhpKj3Z5_0;
	wire w_dff_B_YN02L5Tb2_0;
	wire w_dff_B_nLXJy6dc4_0;
	wire w_dff_B_UNEo6wsu4_0;
	wire w_dff_B_tdOr23mj8_0;
	wire w_dff_B_4KUK3YVo4_0;
	wire w_dff_B_WPrisq2B5_0;
	wire w_dff_B_uohnTt1u7_0;
	wire w_dff_B_bPNl0kxX2_0;
	wire w_dff_B_UJ4VqMGy1_0;
	wire w_dff_B_Dw9LvKPt7_0;
	wire w_dff_B_F3HgZvHC3_0;
	wire w_dff_B_vpUc6sWw9_0;
	wire w_dff_B_MVoAxxd25_0;
	wire w_dff_B_bG5EeO7j0_0;
	wire w_dff_B_our3pX4s3_0;
	wire w_dff_B_SkbhW8q33_0;
	wire w_dff_B_LBl5ZMZc8_0;
	wire w_dff_B_DFK2HWJM3_0;
	wire w_dff_B_zoLJ1wL50_0;
	wire w_dff_B_uFCg0IJZ0_0;
	wire w_dff_B_aQlz3YYd5_0;
	wire w_dff_B_SlYUAo0z9_0;
	wire w_dff_B_sBBes0xc8_0;
	wire w_dff_B_5njRckK90_0;
	wire w_dff_B_85bgcXBo0_0;
	wire w_dff_B_XNJW62EU4_0;
	wire w_dff_B_rkaCF3Ll7_0;
	wire w_dff_B_O8h5cX5Y5_0;
	wire w_dff_B_n87STnP53_0;
	wire w_dff_B_aoEp5HyJ1_0;
	wire w_dff_B_vkl8CucJ7_0;
	wire w_dff_B_XSXQ0ndg2_0;
	wire w_dff_B_qOfmuQz04_0;
	wire w_dff_B_B6IwPksD0_0;
	wire w_dff_B_uYunf61j5_0;
	wire w_dff_B_ZMSEquwr8_0;
	wire w_dff_B_IMqFlEtW8_0;
	wire w_dff_B_fgI9Qkzi7_0;
	wire w_dff_B_RFb61G1o8_0;
	wire w_dff_B_GTjikBJ02_0;
	wire w_dff_B_k8qXUAkW5_0;
	wire w_dff_B_oI172RwO8_0;
	wire w_dff_B_rRnvMP1O8_0;
	wire w_dff_B_T255YwsT7_0;
	wire w_dff_B_42m6RJiu9_0;
	wire w_dff_B_3xcDFFQS6_0;
	wire w_dff_B_11p6Jy1p3_0;
	wire w_dff_B_WgaVymgg2_0;
	wire w_dff_B_rULrk60d0_0;
	wire w_dff_B_e5I5U3Sn2_0;
	wire w_dff_B_t6QLfecs2_0;
	wire w_dff_B_ipxo879F6_0;
	wire w_dff_B_LSskEnMJ6_0;
	wire w_dff_B_kSarhR290_0;
	wire w_dff_B_qwn9lQy21_0;
	wire w_dff_B_WKGrDndw1_0;
	wire w_dff_B_afJdtZAd7_0;
	wire w_dff_B_nNZZktFn6_0;
	wire w_dff_B_7MkIh2KA8_0;
	wire w_dff_B_2yQ49Zkb6_0;
	wire w_dff_B_cHmaKI156_0;
	wire w_dff_B_g6wJIYSG6_0;
	wire w_dff_B_8QVHYHU94_0;
	wire w_dff_B_OLFhO0Yd9_0;
	wire w_dff_B_PxB1hz0Q4_0;
	wire w_dff_B_oXVIDWno3_0;
	wire w_dff_B_PTTpeujz5_0;
	wire w_dff_B_Gwt3tcAo9_0;
	wire w_dff_B_GtQzg2ep8_0;
	wire w_dff_B_2n3G3H5L4_0;
	wire w_dff_B_tsECu0FY7_0;
	wire w_dff_B_VMRiwwx70_0;
	wire w_dff_B_XS0631CG3_0;
	wire w_dff_B_CCSelazc3_0;
	wire w_dff_B_Bsluvwhw1_0;
	wire w_dff_B_51VFRWtS5_0;
	wire w_dff_B_mTeLjdGv6_0;
	wire w_dff_B_yGur854F1_0;
	wire w_dff_B_QUUjOG627_0;
	wire w_dff_B_yoDLszcW6_0;
	wire w_dff_B_VIG8Z6DN4_0;
	wire w_dff_B_QJdXGEHe1_0;
	wire w_dff_B_N4Bt5eBE8_0;
	wire w_dff_B_e92iYarn4_0;
	wire w_dff_B_X76LfSTG3_0;
	wire w_dff_B_2xSQeiu16_0;
	wire w_dff_B_qvtBlUWO1_0;
	wire w_dff_B_YYkGdOSP9_0;
	wire w_dff_B_j3debmty7_0;
	wire w_dff_B_xs3cG4LX2_0;
	wire w_dff_B_x65iNM1F9_0;
	wire w_dff_B_EYuBOgii4_0;
	wire w_dff_B_wI3Cf3A44_0;
	wire w_dff_B_2nixnkQN6_0;
	wire w_dff_B_tGL8PZ947_0;
	wire w_dff_B_Xu7bofGJ3_0;
	wire w_dff_B_k1reFg2Z8_0;
	wire w_dff_B_wmCn36vi4_0;
	wire w_dff_B_tqXKCHTo3_0;
	wire w_dff_B_cIz092fC1_0;
	wire w_dff_B_Yb4ag7pK5_0;
	wire w_dff_B_IGfYsjbi7_0;
	wire w_dff_B_I9vqk8f01_0;
	wire w_dff_B_ZZ7QeuFW7_0;
	wire w_dff_B_RzKjdOXz7_0;
	wire w_dff_B_OTKGhE4w8_0;
	wire w_dff_B_2NqZLi6Q9_0;
	wire w_dff_B_tWOAFbuI2_0;
	wire w_dff_B_pmOHpTZh9_0;
	wire w_dff_B_VYgOSosZ4_0;
	wire w_dff_B_OcWz94yU5_0;
	wire w_dff_B_wfURwYwy5_0;
	wire w_dff_B_UEbPj2ex0_0;
	wire w_dff_B_7qf3MIVd5_0;
	wire w_dff_B_ZhpquE2L4_0;
	wire w_dff_B_Z1sEhCcS4_0;
	wire w_dff_B_aEU3q0Pn6_0;
	wire w_dff_B_49y7Vyes8_0;
	wire w_dff_B_7UwlhvjH8_0;
	wire w_dff_B_L8kWT1sg0_0;
	wire w_dff_B_XIehFfsR7_0;
	wire w_dff_B_3dWOH05e9_0;
	wire w_dff_B_p1G72ESf6_0;
	wire w_dff_B_1dMPIVHc7_0;
	wire w_dff_B_mgpiqFS94_0;
	wire w_dff_B_BIcdm2cr2_0;
	wire w_dff_B_M94wlmKC3_0;
	wire w_dff_B_vcvzEnob7_0;
	wire w_dff_B_JORzm03B9_0;
	wire w_dff_B_WDjfKekK6_0;
	wire w_dff_B_H3rIGwZJ9_0;
	wire w_dff_B_PataCVEL7_0;
	wire w_dff_B_rmNAAghH0_0;
	wire w_dff_B_Xyt7SfeP9_0;
	wire w_dff_B_RW7QdTNT6_0;
	wire w_dff_B_NOPjgN8E1_0;
	wire w_dff_B_t1FPDMuA6_0;
	wire w_dff_B_9PsGZFcP4_0;
	wire w_dff_B_trwb5HFP2_0;
	wire w_dff_B_MH85wwDq2_0;
	wire w_dff_B_TD8lqoHM9_0;
	wire w_dff_B_0zq07tCv1_0;
	wire w_dff_B_W8iGleAw0_0;
	wire w_dff_B_nEqsQrBN6_0;
	wire w_dff_B_pMmiKsav7_0;
	wire w_dff_B_SAq6hZza6_0;
	wire w_dff_B_jPIPrOSc4_0;
	wire w_dff_B_6ylCveDh5_0;
	wire w_dff_B_PvWvV6dw4_0;
	wire w_dff_B_TW2IQEPV5_0;
	wire w_dff_B_2QnUiGPM2_0;
	wire w_dff_B_W99afnE09_0;
	wire w_dff_B_vzjDST0P9_0;
	wire w_dff_B_4O0hpM4s0_0;
	wire w_dff_B_8xvFy2Pr7_0;
	wire w_dff_B_thDQF12t1_0;
	wire w_dff_B_wyMx9J7E2_0;
	wire w_dff_B_0kiQmwvd1_0;
	wire w_dff_B_Dpdunlgl8_0;
	wire w_dff_B_aZ0XF59r1_0;
	wire w_dff_B_iHqJpSWI3_0;
	wire w_dff_B_LO75H4Yn5_0;
	wire w_dff_B_x8z13wvt3_0;
	wire w_dff_B_hFi1hj1w5_0;
	wire w_dff_B_0QbxvLYk6_0;
	wire w_dff_B_Kpd8xOg80_0;
	wire w_dff_B_7pGZFqR42_0;
	wire w_dff_B_BoQxKRqO8_0;
	wire w_dff_B_nPhg2Y2v2_0;
	wire w_dff_B_WOwpDwsM4_0;
	wire w_dff_B_dTK5UeDT8_0;
	wire w_dff_B_Ta56FccG7_0;
	wire w_dff_B_JU7qH4C10_0;
	wire w_dff_B_kB4Q5G4N0_0;
	wire w_dff_B_bcYDuvh83_0;
	wire w_dff_B_8PQLi2Av1_0;
	wire w_dff_B_crRaYzpj9_0;
	wire w_dff_B_dAp8PLhJ4_0;
	wire w_dff_B_fQ7FwhEU7_0;
	wire w_dff_B_UnsEc2uE7_0;
	wire w_dff_B_pLQQcb9k9_0;
	wire w_dff_B_q1onKdbw1_0;
	wire w_dff_B_90EtCyrN6_0;
	wire w_dff_B_tOouyl232_0;
	wire w_dff_B_lFN408lB3_0;
	wire w_dff_B_45Df4SvE2_0;
	wire w_dff_B_U7sKnYuX5_0;
	wire w_dff_B_uwZdqMql6_0;
	wire w_dff_B_jKbNWyGV7_0;
	wire w_dff_B_YkeJOvbQ8_0;
	wire w_dff_B_OYCYOoLr7_0;
	wire w_dff_B_lO2m5XBt1_0;
	wire w_dff_B_wIqwPaG54_0;
	wire w_dff_B_eXa7IXzF1_0;
	wire w_dff_B_zaA4lWdO2_0;
	wire w_dff_B_ynd9DkOR4_0;
	wire w_dff_B_4HGp9GPk0_0;
	wire w_dff_B_OmdS5XFl0_0;
	wire w_dff_B_nba7JulH1_0;
	wire w_dff_B_veUelKvJ3_0;
	wire w_dff_B_tzpsxefS9_0;
	wire w_dff_B_QQFzepC22_0;
	wire w_dff_B_186BDbZ64_0;
	wire w_dff_B_5U3yHgHO5_0;
	wire w_dff_B_ZMD0PT6v8_0;
	wire w_dff_B_BlbrtC3g4_0;
	wire w_dff_B_n153tEVi8_0;
	wire w_dff_B_wfbTXZfQ7_0;
	wire w_dff_B_DsLZT1Gl4_0;
	wire w_dff_B_YSYKevg49_0;
	wire w_dff_B_B6OwF0Vk7_0;
	wire w_dff_B_eIv43cnw5_0;
	wire w_dff_B_FeesYoKp8_0;
	wire w_dff_B_Q2nhRqVk3_0;
	wire w_dff_B_6zUaJIuP2_0;
	wire w_dff_B_EfnJsW652_0;
	wire w_dff_B_TVOrJfM53_0;
	wire w_dff_B_lksUnRe12_0;
	wire w_dff_B_kpiv2kOJ0_0;
	wire w_dff_B_CJ4WeVhJ2_0;
	wire w_dff_B_tWfZRAvY2_0;
	wire w_dff_B_LCpV3k1U4_0;
	wire w_dff_B_Gc1eLvwX5_0;
	wire w_dff_B_ohQ0OD6A2_0;
	wire w_dff_B_dnOehzPz4_0;
	wire w_dff_B_h9TSedPf4_0;
	wire w_dff_B_fu6j3v8y6_0;
	wire w_dff_B_6wxPVSvQ2_0;
	wire w_dff_B_mkYl9cwU3_0;
	wire w_dff_B_sekaV9lY2_0;
	wire w_dff_B_s6xsKBGL4_0;
	wire w_dff_B_LztGLYxd8_0;
	wire w_dff_B_CiNhUuxW8_0;
	wire w_dff_B_k7BLmRYR0_0;
	wire w_dff_B_dk4YZXBy8_0;
	wire w_dff_B_PfP3E5vl4_0;
	wire w_dff_B_qFKiqkCl0_0;
	wire w_dff_B_8uBRtBl74_0;
	wire w_dff_B_Gw0bd02H8_0;
	wire w_dff_B_WidWbth75_0;
	wire w_dff_B_BSSA3qIB8_0;
	wire w_dff_B_SU53ty9J8_0;
	wire w_dff_B_7VIsqoqf7_0;
	wire w_dff_B_nMD9NL467_0;
	wire w_dff_B_yBvmhV2d6_0;
	wire w_dff_B_VNHljr520_0;
	wire w_dff_B_jeg0pcw54_0;
	wire w_dff_B_Ehnn5W3l9_0;
	wire w_dff_B_h6eZu3u20_0;
	wire w_dff_B_jJ915JOS1_0;
	wire w_dff_B_O7XTd4eo8_0;
	wire w_dff_B_TBg2fwns5_0;
	wire w_dff_B_Dvitz8RD4_0;
	wire w_dff_B_LWByTZ2Q6_0;
	wire w_dff_B_sxgDQVCz3_0;
	wire w_dff_B_OgDfNBaa0_0;
	wire w_dff_B_dJodql2R1_0;
	wire w_dff_B_MMcPhios7_0;
	wire w_dff_B_NnBTvtU18_0;
	wire w_dff_B_fpYlcgJ31_0;
	wire w_dff_B_aUWkSl9d9_0;
	wire w_dff_B_yAb9gPcI9_0;
	wire w_dff_B_PRneCuUS5_0;
	wire w_dff_B_4fwnKNCx5_0;
	wire w_dff_B_tMQ513e39_0;
	wire w_dff_B_RjS5uZ9V2_0;
	wire w_dff_B_S8ASuBaQ8_0;
	wire w_dff_B_OKgIkprX4_0;
	wire w_dff_B_we2ry5rk2_0;
	wire w_dff_B_tG45WYAK3_0;
	wire w_dff_B_ktByeRyp8_0;
	wire w_dff_B_OI0RpwXr6_0;
	wire w_dff_B_7SaVDecC8_0;
	wire w_dff_B_mP7mapQj4_0;
	wire w_dff_B_JcDN2b811_0;
	wire w_dff_B_BfaZkbuX5_0;
	wire w_dff_B_yxDNEeLM8_0;
	wire w_dff_B_57i6nzTN8_0;
	wire w_dff_B_2J8CZHmI3_0;
	wire w_dff_B_psDzKZjJ4_0;
	wire w_dff_B_0VddD8N92_0;
	wire w_dff_B_L1BV0WJ00_0;
	wire w_dff_B_WswSo2lL0_0;
	wire w_dff_B_CzFrxsGH7_0;
	wire w_dff_B_5KsNWqcz0_0;
	wire w_dff_B_8sICLYOY8_0;
	wire w_dff_B_p5pgjIrO1_0;
	wire w_dff_B_s7QCceE05_0;
	wire w_dff_B_Ywwt6kAd5_0;
	wire w_dff_B_IIKLaKLN3_0;
	wire w_dff_B_OXyTg80H4_0;
	wire w_dff_B_MSc4yDSg9_0;
	wire w_dff_B_pqJLXFQp1_0;
	wire w_dff_B_Vfx3pym31_0;
	wire w_dff_B_zt4I1oes2_0;
	wire w_dff_B_Yk6LgB6b9_0;
	wire w_dff_B_9aPdJM8K8_0;
	wire w_dff_B_SmsNyQ917_0;
	wire w_dff_B_Srpy44Sh5_0;
	wire w_dff_B_LW8epFDI1_0;
	wire w_dff_B_XtbzDpg11_0;
	wire w_dff_B_k2GTv2do1_0;
	wire w_dff_B_UBV3yPjF9_0;
	wire w_dff_B_nhWUOYV77_0;
	wire w_dff_B_OwAdHxPQ8_0;
	wire w_dff_B_fDafbnRY1_0;
	wire w_dff_B_RPwhy1YW9_0;
	wire w_dff_B_ILpazNn41_0;
	wire w_dff_B_JuZidfGR8_0;
	wire w_dff_B_TdQ3k8jt1_0;
	wire w_dff_B_TGMKnIs32_0;
	wire w_dff_B_3C1Z6RWy2_0;
	wire w_dff_B_ryw6tGTq3_0;
	wire w_dff_B_9LLEM4Rk9_0;
	wire w_dff_B_EutSCtWF0_0;
	wire w_dff_B_PQvP16zN4_0;
	wire w_dff_B_GPSvJbhD0_0;
	wire w_dff_B_6BttYcdu8_0;
	wire w_dff_B_169w74OF5_0;
	wire w_dff_B_v3tbDoey6_0;
	wire w_dff_B_uTo1T5Zm5_0;
	wire w_dff_B_gWZoEuR34_0;
	wire w_dff_B_E1wk1HtI2_0;
	wire w_dff_B_DruCwV8I3_0;
	wire w_dff_B_BUlLTBuT6_0;
	wire w_dff_B_oEbr8wJL8_0;
	wire w_dff_B_hiCdSWKo8_0;
	wire w_dff_B_rS70FZKg6_0;
	wire w_dff_B_eqquUWVM5_0;
	wire w_dff_B_AUaRWg5r2_0;
	wire w_dff_B_geFhxjpM3_0;
	wire w_dff_B_owMPRISI1_0;
	wire w_dff_B_6xRParBy0_0;
	wire w_dff_B_sdbroqEE6_0;
	wire w_dff_B_Be2uaERX3_0;
	wire w_dff_B_EmFoRkGX3_0;
	wire w_dff_B_6ViA2Bib7_0;
	wire w_dff_B_3eTgkbND3_0;
	wire w_dff_B_3OO8t8Jy7_0;
	wire w_dff_B_F2g8Hgm21_0;
	wire w_dff_B_wifpmEyU3_0;
	wire w_dff_B_Inu1hAM00_0;
	wire w_dff_B_MVkbOYWV6_0;
	wire w_dff_B_nYsC4c5E2_0;
	wire w_dff_B_c5HkVFLU9_0;
	wire w_dff_B_18VYH1cw3_0;
	wire w_dff_B_rSnRLbSs2_0;
	wire w_dff_B_eFeV68Nq8_0;
	wire w_dff_B_HW0oeEAb5_0;
	wire w_dff_B_K46a74sM1_0;
	wire w_dff_B_3dBMi0OY9_0;
	wire w_dff_B_9ev7klM63_0;
	wire w_dff_B_Rha8vPz39_0;
	wire w_dff_B_wKvtrW0a8_0;
	wire w_dff_B_1ruvJKk83_0;
	wire w_dff_B_rd7NC96t0_0;
	wire w_dff_B_q8LGSXAh2_0;
	wire w_dff_B_x44yHco41_0;
	wire w_dff_B_hI0h6frj6_0;
	wire w_dff_B_iP2nRo9t5_0;
	wire w_dff_B_i0z6fTE72_0;
	wire w_dff_B_Sz7SJ7zR9_0;
	wire w_dff_B_Nc7UXFJD6_0;
	wire w_dff_B_gJMLFpCx6_0;
	wire w_dff_B_Bei9iEcO9_0;
	wire w_dff_B_la3pvEnT1_0;
	wire w_dff_B_K4Cen4Yd5_0;
	wire w_dff_B_LQoFq0ky3_0;
	wire w_dff_B_ElBtdzJ98_0;
	wire w_dff_B_ZcFoxWzq4_0;
	wire w_dff_B_lXKQqJnz9_0;
	wire w_dff_B_kZJy5mzS5_0;
	wire w_dff_B_jmJiXT5P3_0;
	wire w_dff_B_sNAFJ17s9_0;
	wire w_dff_B_GY10BsD07_0;
	wire w_dff_B_4F7xIhH49_0;
	wire w_dff_B_40TwRlPe2_0;
	wire w_dff_B_cnw7ZXrt7_0;
	wire w_dff_B_5wGIlZSw0_0;
	wire w_dff_B_rUibQj4k7_0;
	wire w_dff_B_JVisCbx96_0;
	wire w_dff_B_K9bul2Ux1_0;
	wire w_dff_B_2K1zDfFj4_0;
	wire w_dff_B_LvzHN8Pt5_0;
	wire w_dff_B_IsZmvvDz7_0;
	wire w_dff_B_x6ZTmAG78_0;
	wire w_dff_B_Nnlu6zqz7_0;
	wire w_dff_B_fl2YKFxC3_0;
	wire w_dff_B_QafPK4mw6_0;
	wire w_dff_B_aY0s1SEW5_0;
	wire w_dff_B_dMpryHiW9_0;
	wire w_dff_B_8jpwtIwW6_0;
	wire w_dff_B_GGXDhljT5_0;
	wire w_dff_B_0JOcTsYA2_0;
	wire w_dff_B_zB6oGyAj9_0;
	wire w_dff_B_vBPOMeOQ3_0;
	wire w_dff_B_IapBKDmK5_0;
	wire w_dff_B_ODRXgujl5_0;
	wire w_dff_B_jKPXe0550_0;
	wire w_dff_B_Hd51AcOE8_0;
	wire w_dff_B_xBFkXBWB5_0;
	wire w_dff_B_dj7hx1W01_0;
	wire w_dff_B_S8AfUY190_0;
	wire w_dff_B_DXLQpCXf7_0;
	wire w_dff_B_JanyqvzG0_0;
	wire w_dff_B_TCmfaA4x9_0;
	wire w_dff_B_WvzYseF72_0;
	wire w_dff_B_6a4aBm4P1_0;
	wire w_dff_B_FtysMW8k5_0;
	wire w_dff_B_Uon6fcLy0_0;
	wire w_dff_B_9QZDgNNG5_0;
	wire w_dff_B_hbjWsio41_0;
	wire w_dff_B_OIsQTUTm0_0;
	wire w_dff_B_Yz3HFJhT3_0;
	wire w_dff_B_OqAbfmLI4_0;
	wire w_dff_B_MUt6SVHt2_0;
	wire w_dff_B_ibIrj1UC5_0;
	wire w_dff_B_IhYCeMkg9_0;
	wire w_dff_B_jZfDpBpZ8_0;
	wire w_dff_B_fdwWzORe9_0;
	wire w_dff_B_Lls6lBYm8_0;
	wire w_dff_B_3MewoJsf4_0;
	wire w_dff_B_V9qk1Xe17_0;
	wire w_dff_B_W0Q43Qoz4_0;
	wire w_dff_B_sQA8Q7vv4_0;
	wire w_dff_B_mCg4hTSy1_0;
	wire w_dff_B_BGPjhzNs0_0;
	wire w_dff_B_Z5d3liEd4_0;
	wire w_dff_B_JXBm3iQl2_0;
	wire w_dff_B_JA25AWF35_0;
	wire w_dff_B_BId30wwf6_0;
	wire w_dff_B_FqviFyMe3_0;
	wire w_dff_B_LiFn6f3S2_0;
	wire w_dff_B_XNuaHbLF9_0;
	wire w_dff_B_j4Dpw5Tz6_0;
	wire w_dff_B_uzC5qiMd1_0;
	wire w_dff_B_NmvSMw1S0_0;
	wire w_dff_B_FaiEpqTG7_0;
	wire w_dff_B_s6J6IifE4_0;
	wire w_dff_B_jkLhY60Q6_0;
	wire w_dff_B_plwjBdGt6_0;
	wire w_dff_B_SFfPXqUT8_0;
	wire w_dff_B_0OLCraVS5_0;
	wire w_dff_B_E2dnobgi5_0;
	wire w_dff_B_3tj5RSZx6_0;
	wire w_dff_B_zi1UCS4e0_0;
	wire w_dff_B_GS8UfAbF7_0;
	wire w_dff_B_by8f38tY4_0;
	wire w_dff_B_vvY2xB2h9_0;
	wire w_dff_B_r7R6QdA01_0;
	wire w_dff_B_eUBIbbcW0_0;
	wire w_dff_B_ZXBeAgIp8_0;
	wire w_dff_B_FhfD9a3Z4_0;
	wire w_dff_B_qefyVb0a7_0;
	wire w_dff_B_peEQAwoh9_0;
	wire w_dff_B_egXWiJTJ1_0;
	wire w_dff_B_2gX100wU4_0;
	wire w_dff_B_0cPouxdx1_0;
	wire w_dff_B_9ku9ANK83_0;
	wire w_dff_B_g3ddMMgx6_0;
	wire w_dff_B_R5L45zxX6_0;
	wire w_dff_B_tZgsYkFL5_0;
	wire w_dff_B_sSbbSwps5_0;
	wire w_dff_B_1PFFfEyj3_0;
	wire w_dff_B_vfGFsx5O2_0;
	wire w_dff_B_ziCdBN9y4_0;
	wire w_dff_B_MSvVpk5b0_0;
	wire w_dff_B_byECFDKU3_0;
	wire w_dff_B_nMB7fsea0_0;
	wire w_dff_B_bzCYf9Yo1_0;
	wire w_dff_B_5O7IJApJ7_0;
	wire w_dff_B_7HD4s21R5_0;
	wire w_dff_B_ZcwQEUZV8_0;
	wire w_dff_B_oLurYfyu7_0;
	wire w_dff_B_4fMJkTpw4_0;
	wire w_dff_B_3cbsogQI9_0;
	wire w_dff_B_Rbv02eXo8_0;
	wire w_dff_B_nR0Dmvzw8_0;
	wire w_dff_B_2bn6Tg174_0;
	wire w_dff_B_xyRRYFcf2_0;
	wire w_dff_B_Cp6X42IN4_0;
	wire w_dff_B_Vmi8WjnT2_0;
	wire w_dff_B_G17vDRnr2_0;
	wire w_dff_B_MvSJL1K94_0;
	wire w_dff_B_0cfnWS3U0_0;
	wire w_dff_B_Q5WprNHv7_0;
	wire w_dff_B_IKDT7cE84_0;
	wire w_dff_B_uxjXNiok6_0;
	wire w_dff_B_mIYGXKEz3_0;
	wire w_dff_B_zs3lhyZS7_0;
	wire w_dff_B_ulKpnZJN8_0;
	wire w_dff_B_O78II1793_0;
	wire w_dff_B_UkCQW7Wl2_0;
	wire w_dff_B_OwN5VRm39_0;
	wire w_dff_B_yxVi8SW62_0;
	wire w_dff_B_7YE2ABml3_0;
	wire w_dff_B_tu08v7UX3_0;
	wire w_dff_B_10M4d7Z52_0;
	wire w_dff_B_fRbqV2wy6_0;
	wire w_dff_B_NyJsLI0T3_0;
	wire w_dff_B_XbVtB5Mq2_0;
	wire w_dff_B_WAddHd7P2_0;
	wire w_dff_B_3sJIglB28_0;
	wire w_dff_B_rOaV7Ugv6_0;
	wire w_dff_B_bRfbUInS4_0;
	wire w_dff_B_nCKdcy2J1_0;
	wire w_dff_B_dRT6h8il9_0;
	wire w_dff_B_wSz2OSMi0_0;
	wire w_dff_B_96zrmQzl9_0;
	wire w_dff_B_ySTaNdRY2_0;
	wire w_dff_B_hcLJBzb28_0;
	wire w_dff_B_QmOxmh3e0_0;
	wire w_dff_B_RXgXFbQm8_0;
	wire w_dff_B_43y5TZ5D9_0;
	wire w_dff_B_O25vugCd0_0;
	wire w_dff_B_KbCjAkss5_0;
	wire w_dff_B_pZj7HHoE4_0;
	wire w_dff_B_cU8nlsz34_0;
	wire w_dff_B_uKfnj3hX2_0;
	wire w_dff_B_217awbSP8_0;
	wire w_dff_B_KjCxAh6I1_0;
	wire w_dff_B_enEOtW2b9_0;
	wire w_dff_B_9Qv9vLt90_0;
	wire w_dff_B_SfvNzWud0_0;
	wire w_dff_B_8Ckt47gu5_0;
	wire w_dff_B_pKa8yGRz6_0;
	wire w_dff_B_19ToeBs49_0;
	wire w_dff_B_IPTl48vD7_0;
	wire w_dff_B_HYG3fEyQ5_0;
	wire w_dff_B_U0anoE9b6_0;
	wire w_dff_B_IITT3hQl4_0;
	wire w_dff_B_zPfwqeM26_0;
	wire w_dff_B_dvk3k9Fa8_0;
	wire w_dff_B_1pp6wd6J6_0;
	wire w_dff_B_bLzcn3G90_0;
	wire w_dff_B_a332ttzI9_0;
	wire w_dff_B_xUiDCcYZ3_0;
	wire w_dff_B_R2YYj88I8_0;
	wire w_dff_B_GAwGDaAm2_0;
	wire w_dff_B_bKAolXuJ8_0;
	wire w_dff_B_5cKWBSSc4_0;
	wire w_dff_B_z6cMncOa4_0;
	wire w_dff_B_5oZj9Pw14_0;
	wire w_dff_B_0VtMN9ot0_0;
	wire w_dff_B_3oBs2ErA5_0;
	wire w_dff_B_CdHiS3wE8_0;
	wire w_dff_B_X7KQmGk40_0;
	wire w_dff_B_DA9hGyi26_0;
	wire w_dff_B_nrfe9TUa7_0;
	wire w_dff_B_qm4t8A883_0;
	wire w_dff_B_NIzJ9Xhw8_0;
	wire w_dff_B_uapVjAvX0_0;
	wire w_dff_B_nAQ4u5JI1_0;
	wire w_dff_B_Ibi5AWnv8_0;
	wire w_dff_B_nFoJi1rY6_0;
	wire w_dff_B_WFA7gEuT7_0;
	wire w_dff_B_s9thuebF3_0;
	wire w_dff_B_8Qi4DYt31_0;
	wire w_dff_B_WGWJJZAy6_0;
	wire w_dff_B_gFYySWJQ0_0;
	wire w_dff_B_6De8olHu6_0;
	wire w_dff_B_KajAw35f7_0;
	wire w_dff_B_MK6rQC9c3_0;
	wire w_dff_B_mSydxlTZ4_0;
	wire w_dff_B_LAF4lqFX7_0;
	wire w_dff_B_yJvNFCgN8_0;
	wire w_dff_B_cIJTFFrx3_0;
	wire w_dff_B_d8Xh6XLg9_0;
	wire w_dff_B_NDRUrUr44_0;
	wire w_dff_B_NJzcooRR5_0;
	wire w_dff_B_nI7y062u3_0;
	wire w_dff_B_VeDz4Sxq6_0;
	wire w_dff_B_oidi940U2_0;
	wire w_dff_B_jqYHvyuE2_0;
	wire w_dff_B_fiEW4LIG5_0;
	wire w_dff_B_un4q9vJO5_0;
	wire w_dff_B_4dsGElRY3_0;
	wire w_dff_B_PevDPDCH7_0;
	wire w_dff_B_U7KCbJ7j9_0;
	wire w_dff_B_5TuiCDz30_0;
	wire w_dff_B_QjdKY39e7_0;
	wire w_dff_B_g2siNU406_0;
	wire w_dff_B_XbFs8ObF9_0;
	wire w_dff_B_riJYA6HL1_0;
	wire w_dff_B_DN2eSvy50_0;
	wire w_dff_B_omRn9OPr4_0;
	wire w_dff_B_Q9hWcdLx1_0;
	wire w_dff_B_C4A8BV2D9_0;
	wire w_dff_B_jQlTkKXq3_0;
	wire w_dff_B_vzCeTABr8_0;
	wire w_dff_B_eyEC9i7o9_0;
	wire w_dff_B_Nu6GfRHJ2_0;
	wire w_dff_B_RoUAEUQC6_0;
	wire w_dff_B_V9WSAKDa9_0;
	wire w_dff_B_c19DGE9n1_0;
	wire w_dff_B_lETFpnV44_0;
	wire w_dff_B_oOk6Qdk90_0;
	wire w_dff_B_6O6Ff7HW3_0;
	wire w_dff_B_3E7xKsAN8_0;
	wire w_dff_B_qfXNonHn6_0;
	wire w_dff_B_HIHTiZ7C7_0;
	wire w_dff_B_U0xETE0X2_0;
	wire w_dff_B_s7O2DkFm3_0;
	wire w_dff_B_SVQM3aM76_0;
	wire w_dff_B_EJoxtvbF2_0;
	wire w_dff_B_gbeiSyXG1_0;
	wire w_dff_B_683DXW4G1_0;
	wire w_dff_B_BmhnnDgj4_0;
	wire w_dff_B_5bAtp4r32_0;
	wire w_dff_B_CjopLBoS1_0;
	wire w_dff_B_ttaQeut41_0;
	wire w_dff_B_xuig0HHX7_0;
	wire w_dff_B_McHRGvS39_0;
	wire w_dff_B_IDjDcG623_0;
	wire w_dff_B_XSeuToPy2_0;
	wire w_dff_B_PDpSigoa0_0;
	wire w_dff_B_34pJQqSm4_0;
	wire w_dff_B_ikr9acNu9_0;
	wire w_dff_B_UA4W1WE27_0;
	wire w_dff_B_iBHJO64Z5_0;
	wire w_dff_B_Rh4MhzGV0_0;
	wire w_dff_B_LQXrrTHw1_0;
	wire w_dff_B_ckVcF37S6_0;
	wire w_dff_B_yOJi19wI4_0;
	wire w_dff_B_5hWvwEST9_0;
	wire w_dff_B_5QJS6uLd2_0;
	wire w_dff_B_SnZrmw4R8_0;
	wire w_dff_B_ozoqehRA8_0;
	wire w_dff_B_g3SxB9Dm7_0;
	wire w_dff_B_jl9lQTkz5_0;
	wire w_dff_B_7gY3sxkf2_0;
	wire w_dff_B_bCXGpT5d5_0;
	wire w_dff_B_vinPkQyy1_0;
	wire w_dff_B_RZADuqLD0_0;
	wire w_dff_B_qMgMRE2O0_0;
	wire w_dff_B_DMyIg8314_0;
	wire w_dff_B_acXU7HXC4_0;
	wire w_dff_B_FugCq6a90_0;
	wire w_dff_B_xzgIeZa82_0;
	wire w_dff_B_AYtav6441_0;
	wire w_dff_B_H7tT1WGg7_0;
	wire w_dff_B_3OyFvk4g5_0;
	wire w_dff_B_4CNIiIZT6_0;
	wire w_dff_B_aoqb0R2S4_0;
	wire w_dff_B_xwJz2MHm6_0;
	wire w_dff_B_feSsaIf44_0;
	wire w_dff_B_SkkzHgmv3_0;
	wire w_dff_B_0vsm1U1t4_0;
	wire w_dff_B_Y7ZAL5IZ0_0;
	wire w_dff_B_1EBayVfX0_0;
	wire w_dff_B_XimjgfD55_0;
	wire w_dff_B_VLCqTYut9_0;
	wire w_dff_B_sARaI0Ke1_0;
	wire w_dff_B_CVZrcz8n5_0;
	wire w_dff_B_HyGs87ZG4_0;
	wire w_dff_B_kv9GIGkv4_0;
	wire w_dff_B_5zy633b08_0;
	wire w_dff_B_NaTYdP5T6_0;
	wire w_dff_B_QTy547KM6_0;
	wire w_dff_B_bwENjw0O5_0;
	wire w_dff_B_DONxhJQu0_0;
	wire w_dff_B_0KY7RqAv0_0;
	wire w_dff_B_v2XPfulv5_0;
	wire w_dff_B_iwOAdbGe8_0;
	wire w_dff_B_lj5oT0lg6_0;
	wire w_dff_B_b9TMSY913_0;
	wire w_dff_B_DTD5nbG36_0;
	wire w_dff_B_iTPMRVvg6_0;
	wire w_dff_B_tiske0pB1_0;
	wire w_dff_B_KUdz2CJa8_0;
	wire w_dff_B_X3NPnCiV5_0;
	wire w_dff_B_n0H4Z3Uk4_0;
	wire w_dff_B_cCLBdCMf8_0;
	wire w_dff_B_BVJmrVS73_0;
	wire w_dff_B_Hls79WUD8_0;
	wire w_dff_B_uma5x3EP1_0;
	wire w_dff_B_O4OgeXrX5_0;
	wire w_dff_B_XFvWNnpT5_0;
	wire w_dff_B_FdDuKjM23_0;
	wire w_dff_B_BpfTb8Mn0_0;
	wire w_dff_B_6YZ0MEFL6_0;
	wire w_dff_B_R9Rapnri9_0;
	wire w_dff_B_fjRGz4vp6_0;
	wire w_dff_B_tQF2amq15_0;
	wire w_dff_B_DexEJ0qv7_0;
	wire w_dff_B_iTGijb4G3_0;
	wire w_dff_B_OBMEBLRR5_0;
	wire w_dff_B_YzSXgHQL7_0;
	wire w_dff_B_iLhXKM2I1_0;
	wire w_dff_B_DF3UfJ7A4_0;
	wire w_dff_B_WBrmP0OL6_0;
	wire w_dff_B_M32JFkM21_0;
	wire w_dff_B_TbxqKTGH9_0;
	wire w_dff_B_NtFQpDHd1_0;
	wire w_dff_B_i2ZeriDB6_0;
	wire w_dff_B_Y0i3i1aI8_0;
	wire w_dff_B_kJ1OIEFu0_0;
	wire w_dff_B_515I7mq45_0;
	wire w_dff_B_Oeu12Ync6_0;
	wire w_dff_B_vW9kxOqW9_0;
	wire w_dff_B_cDVxcvt91_0;
	wire w_dff_B_pJtGYLR11_0;
	wire w_dff_B_q9r0iuA15_0;
	wire w_dff_B_xNHUsXCf0_0;
	wire w_dff_B_CTyWitmH7_0;
	wire w_dff_B_HbI5Xm1a1_0;
	wire w_dff_B_HvZTQnBa6_0;
	wire w_dff_B_GaY4qt4a6_0;
	wire w_dff_B_K3pQ5h3w7_0;
	wire w_dff_B_qo3EOGlQ0_0;
	wire w_dff_B_kMkBYx3G0_0;
	wire w_dff_B_3D7PmEZW1_0;
	wire w_dff_B_FRZFB3478_0;
	wire w_dff_B_vlaHuW2B7_0;
	wire w_dff_B_Gf76VPPs4_0;
	wire w_dff_B_BZFvn93D9_0;
	wire w_dff_B_fLKBBBCo5_0;
	wire w_dff_B_cjnZ9Qlu7_0;
	wire w_dff_B_0qILxkjt9_0;
	wire w_dff_B_FVAxEKMA6_0;
	wire w_dff_B_ER3waTSn2_0;
	wire w_dff_B_tjAPeAJ01_0;
	wire w_dff_B_na8ylLxA0_0;
	wire w_dff_B_fQentjdi1_0;
	wire w_dff_B_LPOgw3ob1_0;
	wire w_dff_B_1xwZuAru7_0;
	wire w_dff_B_rLkqJbTJ8_0;
	wire w_dff_B_4EazO7Zy9_0;
	wire w_dff_B_8qdQpabr3_0;
	wire w_dff_B_UWt7o4dv5_0;
	wire w_dff_B_eaMsKA4H0_0;
	wire w_dff_B_h4aUYj344_0;
	wire w_dff_B_oaTA7AA74_0;
	wire w_dff_B_AtWNkgKv1_0;
	wire w_dff_B_k6zCwV8k1_0;
	wire w_dff_B_O1KolSyU1_0;
	wire w_dff_B_3FVBTjde4_0;
	wire w_dff_B_Nn2pDx1S4_0;
	wire w_dff_B_jX7DVGGu5_0;
	wire w_dff_B_XeWl1wDu0_0;
	wire w_dff_B_vQLxsDKn6_0;
	wire w_dff_B_txjZgmlX0_0;
	wire w_dff_B_NYNGcIk41_0;
	wire w_dff_B_n1rpOmAn9_0;
	wire w_dff_B_NIhTncFp9_0;
	wire w_dff_B_HdqDu6U36_0;
	wire w_dff_B_RHJZsHOH9_0;
	wire w_dff_B_pMSCIz955_0;
	wire w_dff_B_My4ZOapN3_0;
	wire w_dff_B_gq6333Mh8_0;
	wire w_dff_B_ukokP1Kv3_0;
	wire w_dff_B_BXBwBDdk0_0;
	wire w_dff_B_sNvwIeOx5_0;
	wire w_dff_B_OcZ9YFZp5_0;
	wire w_dff_B_MJS4mRfO8_0;
	wire w_dff_B_MujxiHya4_0;
	wire w_dff_B_yhksFV181_0;
	wire w_dff_B_kyv3tfV22_0;
	wire w_dff_B_nP6cZpCl4_0;
	wire w_dff_B_l9xN2bV80_0;
	wire w_dff_B_Q7GsqJgO9_0;
	wire w_dff_B_Gy8x11xb5_0;
	wire w_dff_B_akCtNz9q8_0;
	wire w_dff_B_7bacJMT45_0;
	wire w_dff_B_Mu7xJ6494_0;
	wire w_dff_B_aiQujMYy4_0;
	wire w_dff_B_V54ZLEyd6_0;
	wire w_dff_B_OpDFoOTy1_0;
	wire w_dff_B_XJOIHvXK3_0;
	wire w_dff_B_cDh3cUFn2_0;
	wire w_dff_B_CWU2bbfI4_0;
	wire w_dff_B_k043bbsw9_0;
	wire w_dff_B_UPHwnOKn9_0;
	wire w_dff_B_Ursiat8U0_0;
	wire w_dff_B_WenzMoZn5_0;
	wire w_dff_B_Pedb5i9v1_0;
	wire w_dff_B_eGWiGWuv9_0;
	wire w_dff_B_Z6tMjP6B4_0;
	wire w_dff_B_hdhHwUwg1_0;
	wire w_dff_B_G6vSpW5m7_0;
	wire w_dff_B_xhUP7fvG0_0;
	wire w_dff_B_ICyfZ5Ai3_0;
	wire w_dff_B_5y4jQn4h6_0;
	wire w_dff_B_fPCg0bHC7_0;
	wire w_dff_B_a656EM6I6_0;
	wire w_dff_B_EKqKVKYc2_0;
	wire w_dff_B_UWRk1O027_0;
	wire w_dff_B_N7DmpM2p4_0;
	wire w_dff_B_xN4GSsOI9_0;
	wire w_dff_B_gOmI6URF1_0;
	wire w_dff_B_03uW9gTi8_0;
	wire w_dff_B_nqObvXTJ0_0;
	wire w_dff_B_qFUYtomk5_0;
	wire w_dff_B_myLaGLRL4_0;
	wire w_dff_B_Hdw3qxMg6_0;
	wire w_dff_B_TpAwsMsu0_0;
	wire w_dff_B_ZhA7BnFW3_0;
	wire w_dff_B_hL1I0h6t8_0;
	wire w_dff_B_2xYT2Nog2_0;
	wire w_dff_B_YiiTRArl1_0;
	wire w_dff_B_GE2mGqKL5_0;
	wire w_dff_B_chPYLgF62_0;
	wire w_dff_B_T2jR5Ota3_0;
	wire w_dff_B_jK2apygH2_0;
	wire w_dff_B_VBJFopmb1_0;
	wire w_dff_B_KAGUHmsE6_0;
	wire w_dff_B_qPCq6zoJ0_0;
	wire w_dff_B_dvXCZErz5_0;
	wire w_dff_B_bNn9kino5_0;
	wire w_dff_B_4AzEzqTM6_0;
	wire w_dff_B_xZm2pGyh8_0;
	wire w_dff_B_zUUlLEYb7_0;
	wire w_dff_B_sxSxIZwr7_0;
	wire w_dff_B_cV0tdWP02_0;
	wire w_dff_B_GoozpgYI0_0;
	wire w_dff_B_irIfkTAY9_0;
	wire w_dff_B_cRRE6kJz0_0;
	wire w_dff_B_S0hdnirW3_0;
	wire w_dff_B_AtBCkKkY5_0;
	wire w_dff_B_uOxYj7qZ1_0;
	wire w_dff_B_U4P79lTw3_0;
	wire w_dff_B_poqdFB3x7_0;
	wire w_dff_B_4vnyuzy01_0;
	wire w_dff_B_VuM2OjLO4_0;
	wire w_dff_B_oYUeOmx77_0;
	wire w_dff_B_uU8kckxO3_0;
	wire w_dff_B_mxiamplP9_0;
	wire w_dff_B_leaqwRHk4_0;
	wire w_dff_B_cZJonqiL8_0;
	wire w_dff_B_659s3U2q7_0;
	wire w_dff_B_9YaPMIhN0_0;
	wire w_dff_B_uMjB28FB9_0;
	wire w_dff_B_GG5sD3FW6_0;
	wire w_dff_B_f08spvnV0_0;
	wire w_dff_B_Rc1sRFHO8_0;
	wire w_dff_B_ZAgPOUSz7_0;
	wire w_dff_B_WRuwlgAp9_0;
	wire w_dff_B_pTDgQpyy0_0;
	wire w_dff_B_ZEx5grzP6_0;
	wire w_dff_B_WetPrXur0_0;
	wire w_dff_B_tG8aemG22_0;
	wire w_dff_B_lM0srbnz1_0;
	wire w_dff_B_c8cb8YR29_0;
	wire w_dff_B_QL4QL1ok3_0;
	wire w_dff_B_OvwJsaxy3_0;
	wire w_dff_B_qkyB8GPw3_0;
	wire w_dff_B_gcyrlYWI8_0;
	wire w_dff_B_utaX2tZo7_0;
	wire w_dff_B_3PY73daK5_0;
	wire w_dff_B_dtl0pjpD9_0;
	wire w_dff_B_wGd6jGjQ2_0;
	wire w_dff_B_W5O1D9Sp9_0;
	wire w_dff_B_FBhFPXnx9_0;
	wire w_dff_B_oc2VA5YM2_0;
	wire w_dff_B_EYo8R46K4_0;
	wire w_dff_B_jrRbyq497_0;
	wire w_dff_B_WiwTm3sF9_0;
	wire w_dff_B_98Tylq7e8_0;
	wire w_dff_B_UNX9CF5n9_0;
	wire w_dff_B_wmuF7Gyw8_0;
	wire w_dff_B_ixXLIgpD9_0;
	wire w_dff_B_RwcTgqMI0_0;
	wire w_dff_B_oYhZq91j9_0;
	wire w_dff_B_jg73UTkb8_0;
	wire w_dff_B_U6YufzZX2_0;
	wire w_dff_B_LGLrxn9n8_0;
	wire w_dff_B_nzVGwEhw3_0;
	wire w_dff_B_UsWbYh5u8_0;
	wire w_dff_B_mw3sseZp8_0;
	wire w_dff_B_6NZl6yYS6_0;
	wire w_dff_B_3gHD8I003_0;
	wire w_dff_B_9MSeXjVk6_0;
	wire w_dff_B_USJUgjM55_0;
	wire w_dff_B_CyOuxERh9_0;
	wire w_dff_B_V7Ib9fpJ1_0;
	wire w_dff_B_UNnD9opa5_0;
	wire w_dff_B_w4hhfaAA3_0;
	wire w_dff_B_RfnKpmUW5_0;
	wire w_dff_B_QFngED6z3_0;
	wire w_dff_B_zhUwLWLv2_0;
	wire w_dff_B_js52DzsR9_0;
	wire w_dff_B_cQv8lHFu4_0;
	wire w_dff_B_ASAy6Jg10_0;
	wire w_dff_B_fV5OmoIN2_0;
	wire w_dff_B_UTK9vC4t4_0;
	wire w_dff_B_U7zIeVLj4_0;
	wire w_dff_B_mdYh0M4r5_0;
	wire w_dff_B_PgRhADgl6_0;
	wire w_dff_B_ul48SBz97_0;
	wire w_dff_B_9p7xzlIp3_0;
	wire w_dff_B_CdeWzgM28_0;
	wire w_dff_B_5yBunGSQ8_0;
	wire w_dff_B_x0WdS5e65_0;
	wire w_dff_B_ZpqICiyX9_0;
	wire w_dff_B_otsDwvqB3_0;
	wire w_dff_B_eMqcbWqV4_0;
	wire w_dff_B_BnpiaI0O1_0;
	wire w_dff_B_FInMvcY67_0;
	wire w_dff_B_KQX3qftb1_0;
	wire w_dff_B_wR3EJoxe7_0;
	wire w_dff_B_57uY1CXv3_0;
	wire w_dff_B_1HRlSZAR2_0;
	wire w_dff_B_xnyzMUxu5_0;
	wire w_dff_B_8ubBVz866_0;
	wire w_dff_B_9EJx8tWJ3_0;
	wire w_dff_B_yjHX2iy78_0;
	wire w_dff_B_GDzeQc6Q8_0;
	wire w_dff_B_fUrlSf5P4_0;
	wire w_dff_B_ossniog09_0;
	wire w_dff_B_7UWCIscI1_0;
	wire w_dff_B_TYPlv2uD4_0;
	wire w_dff_B_X86le55n6_0;
	wire w_dff_B_DAC1g3TT6_0;
	wire w_dff_B_ZXJBwqzf4_0;
	wire w_dff_B_gWGVgIsu2_0;
	wire w_dff_B_EHBKLGB74_0;
	wire w_dff_B_SrGuoJOq9_0;
	wire w_dff_B_2Kzh4c4E2_0;
	wire w_dff_B_IS5Skb8y1_0;
	wire w_dff_B_ysJOZP5q0_0;
	wire w_dff_B_YbdqseU76_0;
	wire w_dff_B_gZ8DvZdn8_0;
	wire w_dff_B_uxmgcEOt7_0;
	wire w_dff_B_qEeD1Y121_0;
	wire w_dff_B_tGyFtL8g5_0;
	wire w_dff_B_ZMVjOfh13_0;
	wire w_dff_B_Yjq2hmXF0_0;
	wire w_dff_B_WieN8Xbb0_0;
	wire w_dff_B_HBpI1Stx1_0;
	wire w_dff_B_RnB35QRk1_0;
	wire w_dff_B_mPn94spR7_0;
	wire w_dff_B_G2fLqw7w0_0;
	wire w_dff_B_z7L8HmGP2_0;
	wire w_dff_B_bOYXgBcF0_0;
	wire w_dff_B_CKQVhFj62_0;
	wire w_dff_B_6ASsgS4d6_0;
	wire w_dff_B_AoWd7XVJ6_0;
	wire w_dff_B_mT6luw553_0;
	wire w_dff_B_RYyCr0Jl8_0;
	wire w_dff_B_VQHeG0RE9_0;
	wire w_dff_B_U1MaEUnW4_0;
	wire w_dff_B_7eW38oI83_0;
	wire w_dff_B_nMZ7Qmwa1_0;
	wire w_dff_B_pJdkeARO9_0;
	wire w_dff_B_RWqMEuI92_0;
	wire w_dff_B_PeohdI955_0;
	wire w_dff_B_W1uLlMar7_0;
	wire w_dff_B_nNlo2cPj5_0;
	wire w_dff_B_IQRe3tTm0_0;
	wire w_dff_B_002zxTFy5_0;
	wire w_dff_B_xX7EUYh51_0;
	wire w_dff_B_rxmp0ZJd1_0;
	wire w_dff_B_ZJKUfoRx0_0;
	wire w_dff_B_T0Aj8f960_0;
	wire w_dff_B_9irEKkA48_0;
	wire w_dff_B_Eztovppw0_0;
	wire w_dff_B_iTMTLhTL3_0;
	wire w_dff_B_ZwJF8mxF1_0;
	wire w_dff_B_4r5E3uWs9_0;
	wire w_dff_B_5l6h7VVR4_0;
	wire w_dff_B_Y3hWmEb72_0;
	wire w_dff_B_oK8jQHfj9_0;
	wire w_dff_B_E2MPlqZv8_0;
	wire w_dff_B_LPwPZoL92_0;
	wire w_dff_B_7eD41BBB2_0;
	wire w_dff_B_flSfCuIw5_0;
	wire w_dff_B_Xp9QBovF0_0;
	wire w_dff_B_CDZDHRbE1_0;
	wire w_dff_B_2LytpcSC1_0;
	wire w_dff_B_txdEc3XX4_0;
	wire w_dff_B_24N9Dxzp9_0;
	wire w_dff_B_xuLvqdrB8_0;
	wire w_dff_B_kmVvkjfY9_0;
	wire w_dff_B_vghfCz9w4_0;
	wire w_dff_B_cCrAwSXp4_0;
	wire w_dff_B_akSnWl4a4_0;
	wire w_dff_B_g8inP2hw8_0;
	wire w_dff_B_OOaMoRMD8_0;
	wire w_dff_B_N43TeiBD7_0;
	wire w_dff_B_LkDa6SzL3_0;
	wire w_dff_B_edGyBkYI7_0;
	wire w_dff_B_LFmc4WlW5_0;
	wire w_dff_B_dhV4u7s49_0;
	wire w_dff_B_ezBkCv0e7_0;
	wire w_dff_B_nTKJilRV1_0;
	wire w_dff_B_ac8co5MC9_0;
	wire w_dff_B_Ec9Nilic5_0;
	wire w_dff_B_FgwoQ8oz7_0;
	wire w_dff_B_5U9XJDKT8_0;
	wire w_dff_B_BHAwMt4x9_0;
	wire w_dff_B_HyKhLGrt0_0;
	wire w_dff_B_ahlsgZnF1_0;
	wire w_dff_B_dDsQNd3P2_0;
	wire w_dff_B_FtIWvVPE0_0;
	wire w_dff_B_rTIcnVp34_0;
	wire w_dff_B_skcRmArv1_0;
	wire w_dff_B_663jYFYu6_0;
	wire w_dff_B_DnYynrPR9_0;
	wire w_dff_B_DNRvwmFk7_0;
	wire w_dff_B_q2iQDC5i5_0;
	wire w_dff_B_FGpFsdqf2_0;
	wire w_dff_B_qJLgeLAP9_0;
	wire w_dff_B_DmqOkRzm7_0;
	wire w_dff_B_b182Fq3j2_0;
	wire w_dff_B_xN4tYXk49_0;
	wire w_dff_B_9xug5xDH5_0;
	wire w_dff_B_B7r84Fjh7_0;
	wire w_dff_B_6mQeXNux4_0;
	wire w_dff_B_vmjRRzfx6_0;
	wire w_dff_B_Q3Y7OAQm2_0;
	wire w_dff_B_5MvIazEW6_0;
	wire w_dff_B_pbzTpi4o4_0;
	wire w_dff_B_kmtiB6zx5_0;
	wire w_dff_B_Fx10VEcz9_0;
	wire w_dff_B_5wLAcNXb8_0;
	wire w_dff_B_2STa13D53_0;
	wire w_dff_B_uyOxNtuO5_0;
	wire w_dff_B_IrJaJ9z73_0;
	wire w_dff_B_bZqN31Th5_0;
	wire w_dff_B_0qqe029j5_0;
	wire w_dff_B_CmA98J3t2_0;
	wire w_dff_B_4OBh7iPL5_0;
	wire w_dff_B_XjSdbsaK1_0;
	wire w_dff_B_cUZt5DxM0_0;
	wire w_dff_B_Rh3ZUMp52_0;
	wire w_dff_B_bPqCWENT8_0;
	wire w_dff_B_6JwUP94n3_0;
	wire w_dff_B_mHpZ10hv2_0;
	wire w_dff_B_L1rg5cw88_0;
	wire w_dff_B_wneQG0uC7_0;
	wire w_dff_B_M5p0jvDy7_0;
	wire w_dff_B_DK1hHNJv9_0;
	wire w_dff_B_Ryw32P2a3_0;
	wire w_dff_B_BSSWA0AA3_0;
	wire w_dff_B_lVJ0xiQs5_0;
	wire w_dff_B_G2lXWRYT1_0;
	wire w_dff_B_LIAYzsse5_0;
	wire w_dff_B_f4nkdD6i2_0;
	wire w_dff_B_fMEyUaIT3_0;
	wire w_dff_B_MJOgI5Tc8_0;
	wire w_dff_B_l9494gur8_0;
	wire w_dff_B_0xgzJT2y1_0;
	wire w_dff_B_mnqrLOv22_0;
	wire w_dff_B_oXBcbJhl3_0;
	wire w_dff_B_3HCC4K1y4_0;
	wire w_dff_B_501avdZ33_0;
	wire w_dff_B_asE3GayY1_0;
	wire w_dff_B_iUDXFsaS3_0;
	wire w_dff_B_giK7g9yx2_0;
	wire w_dff_B_6R7Dh7px6_0;
	wire w_dff_B_Ifx59pLf6_0;
	wire w_dff_B_pimWYWdx2_0;
	wire w_dff_B_oIFulJes4_0;
	wire w_dff_B_WuPeaXXs8_0;
	wire w_dff_B_5xHWplqn2_0;
	wire w_dff_B_gC55LX6C2_0;
	wire w_dff_B_o64XK9bE4_0;
	wire w_dff_B_fCQBGIZ69_0;
	wire w_dff_B_0QA7Xj7o3_0;
	wire w_dff_B_Rt9HNFXs3_0;
	wire w_dff_B_DPB8dIwm2_0;
	wire w_dff_B_edIqXs2R6_0;
	wire w_dff_B_dBZ8UPtm0_0;
	wire w_dff_B_eoV108Gw8_0;
	wire w_dff_B_ZURMnqwx6_0;
	wire w_dff_B_bckQAAPB7_0;
	wire w_dff_B_AOn8vtPx9_0;
	wire w_dff_B_F2WvPzWR4_0;
	wire w_dff_B_UUF9AEbV8_0;
	wire w_dff_B_qKcTuZkc3_0;
	wire w_dff_B_PSBnQFqD2_0;
	wire w_dff_B_YwZPwZcG8_0;
	wire w_dff_B_y2YeFqmQ4_0;
	wire w_dff_B_RnW0Gm953_0;
	wire w_dff_B_RVI3Wf2a7_0;
	wire w_dff_B_Sf5gLHx05_0;
	wire w_dff_B_Ha4Boxhu5_0;
	wire w_dff_B_ZzaDVEjL2_0;
	wire w_dff_B_9Y3EJ03L8_0;
	wire w_dff_B_5F1KABog7_0;
	wire w_dff_B_kr0RBh2v6_0;
	wire w_dff_B_f6rVGAmV0_0;
	wire w_dff_B_o8aPkdjX8_0;
	wire w_dff_B_cEBpO5LL5_0;
	wire w_dff_B_G3IMKIUJ8_0;
	wire w_dff_B_XuPlBzz87_0;
	wire w_dff_B_DKD7axMF5_0;
	wire w_dff_B_73KFAbEP4_0;
	wire w_dff_B_62dTet6S2_0;
	wire w_dff_B_bKUQ5i801_0;
	wire w_dff_B_0Wk2wlyL4_0;
	wire w_dff_B_2OReU4Y06_0;
	wire w_dff_B_Lv8WuXOu5_0;
	wire w_dff_B_Af5Y2zzz6_0;
	wire w_dff_B_XkPvtMI32_0;
	wire w_dff_B_mJ1XUryB9_0;
	wire w_dff_B_gibCcTwN0_0;
	wire w_dff_B_79Vh9ZuL1_0;
	wire w_dff_B_JdGYQgyg8_0;
	wire w_dff_B_6VzbeitE7_0;
	wire w_dff_B_X8L8LwPo4_0;
	wire w_dff_B_cIvQSKz17_0;
	wire w_dff_B_bCDgvB6u8_0;
	wire w_dff_B_AZa3Ty4w1_0;
	wire w_dff_B_awCzRtA72_0;
	wire w_dff_B_MSTl2hYf1_0;
	wire w_dff_B_O9NJs6ZX4_0;
	wire w_dff_B_YRxR1LVA8_0;
	wire w_dff_B_G8PskRw15_0;
	wire w_dff_B_Z3WDt5Ih7_0;
	wire w_dff_B_lwby5Mh50_0;
	wire w_dff_B_eic3tLtR8_0;
	wire w_dff_B_cBEC74E59_0;
	wire w_dff_B_h9OvX51Z9_0;
	wire w_dff_B_OMdxyjmK4_0;
	wire w_dff_B_oGtPmaNF8_0;
	wire w_dff_B_kQsivHJf4_0;
	wire w_dff_B_Qf67nob83_0;
	wire w_dff_B_KoaiLJSL2_0;
	wire w_dff_B_5rTuTRhA7_0;
	wire w_dff_B_BgkCpQ985_0;
	wire w_dff_B_xW01B4j49_0;
	wire w_dff_B_mLA5TeLw9_0;
	wire w_dff_B_RtLE5QMn2_0;
	wire w_dff_B_1OZ8NVel5_0;
	wire w_dff_B_gGFcK9Yb2_0;
	wire w_dff_B_BEPcJJdl5_0;
	wire w_dff_B_OuqUwewK7_0;
	wire w_dff_B_LhWWmIhT3_0;
	wire w_dff_B_wrPEluAf3_0;
	wire w_dff_B_v2q8aYLY4_0;
	wire w_dff_B_gFOpIouM5_0;
	wire w_dff_B_n03IOPfk4_0;
	wire w_dff_B_lILpXwza7_0;
	wire w_dff_B_krrbxW3D4_0;
	wire w_dff_B_uz0YGazH1_0;
	wire w_dff_B_oeu2xniw1_0;
	wire w_dff_B_fwaYqs5M7_0;
	wire w_dff_B_WIdKIBsv3_0;
	wire w_dff_B_CixI2yI33_0;
	wire w_dff_B_ElNs0U4u4_0;
	wire w_dff_B_64VOXAXb8_0;
	wire w_dff_B_6OTmtGd90_0;
	wire w_dff_B_LV1iaPcs6_0;
	wire w_dff_B_C8mbCvAT8_0;
	wire w_dff_B_wBKYXJd46_0;
	wire w_dff_B_0cF1byO62_0;
	wire w_dff_B_7tBP0pSU8_0;
	wire w_dff_B_YFOvMl5c1_0;
	wire w_dff_B_OZSfx8AM0_0;
	wire w_dff_B_dUtt2DQQ5_0;
	wire w_dff_B_GEwKrSO94_0;
	wire w_dff_B_bU9DLaMx5_0;
	wire w_dff_B_XPR0PIQn0_0;
	wire w_dff_B_7rcaRNpq3_0;
	wire w_dff_B_BeQ7UtIn1_0;
	wire w_dff_B_snrQQy319_0;
	wire w_dff_B_97akbQ6i1_0;
	wire w_dff_B_6LC8AMi52_0;
	wire w_dff_B_oLV1RueZ1_0;
	wire w_dff_B_RdcO64tI8_0;
	wire w_dff_B_ou7AWJVb2_0;
	wire w_dff_B_qyexQIWU9_0;
	wire w_dff_B_9ivRqQdT2_0;
	wire w_dff_B_jk3ijHHm1_0;
	wire w_dff_B_H93DD0nF3_0;
	wire w_dff_B_8SXtvf059_0;
	wire w_dff_B_MYuLOHxF1_0;
	wire w_dff_B_0UMr1DXF2_0;
	wire w_dff_B_ByR9WVct7_0;
	wire w_dff_B_DFE8za0Y6_0;
	wire w_dff_B_eTO73Wi26_0;
	wire w_dff_B_UgDRVKEi3_0;
	wire w_dff_B_r9BUGi6K8_0;
	wire w_dff_B_ilVFZ8n37_0;
	wire w_dff_B_mUp05Keq0_0;
	wire w_dff_B_7mz2ApX05_0;
	wire w_dff_B_uvEu02rc7_0;
	wire w_dff_B_yA5JL2DC2_0;
	wire w_dff_B_oeXcKNM27_0;
	wire w_dff_B_4RqP3Tsd3_0;
	wire w_dff_B_UsHcIBFJ8_0;
	wire w_dff_B_ZXKcvya14_0;
	wire w_dff_B_tYyKXsSX6_0;
	wire w_dff_B_VQNZlPJU6_0;
	wire w_dff_B_H48w7ZK64_0;
	wire w_dff_B_84PtJf3j8_0;
	wire w_dff_B_6vGDRYsK8_0;
	wire w_dff_B_EmB0F3rz2_0;
	wire w_dff_B_YDxM8RvD9_0;
	wire w_dff_B_1bXMOldO3_0;
	wire w_dff_B_a9yFeR9J2_0;
	wire w_dff_B_yagBJeom2_0;
	wire w_dff_B_ZEFvyu3s1_0;
	wire w_dff_B_UDWZpxXx5_0;
	wire w_dff_B_S1OTrQt82_0;
	wire w_dff_B_eNp8XkoY1_0;
	wire w_dff_B_1X6NMZH98_0;
	wire w_dff_B_g3LEmZ0x0_0;
	wire w_dff_B_KevCz5qh3_0;
	wire w_dff_B_7gtftLoY5_0;
	wire w_dff_B_BMELB3022_0;
	wire w_dff_B_m2QO5VPj0_0;
	wire w_dff_B_B28S41fk9_0;
	wire w_dff_B_z5Dxn7683_0;
	wire w_dff_B_507vvQel3_0;
	wire w_dff_B_0LW7LDP95_0;
	wire w_dff_B_Nex9M55S9_0;
	wire w_dff_B_CEVq4Ild6_0;
	wire w_dff_B_Bj1gmevW8_0;
	wire w_dff_B_uMtHdGF47_0;
	wire w_dff_B_fYF9UXz07_0;
	wire w_dff_B_QAeX4v7Y2_0;
	wire w_dff_B_4f3IQ6te8_0;
	wire w_dff_B_PxVXR3hD0_0;
	wire w_dff_B_nsnTKwkU2_0;
	wire w_dff_B_6gGyzA4X6_0;
	wire w_dff_B_TaqQMqcn5_0;
	wire w_dff_B_qLRmuQ330_0;
	wire w_dff_B_mRnocC4A3_0;
	wire w_dff_B_wNzQNQMS8_0;
	wire w_dff_B_MWtU1QuQ8_0;
	wire w_dff_B_VkLYDPww2_0;
	wire w_dff_B_sZUtHWnX4_0;
	wire w_dff_B_z45pZN5j0_0;
	wire w_dff_B_EA39EuGF6_0;
	wire w_dff_B_U0kVPIme6_0;
	wire w_dff_B_zX9xjztb5_0;
	wire w_dff_B_GwwfIdIG0_0;
	wire w_dff_B_QSc3XySm2_0;
	wire w_dff_B_aOMPMwkk4_0;
	wire w_dff_B_82AmGAYp6_0;
	wire w_dff_B_fO2xFMpA9_0;
	wire w_dff_B_odjCbIQs7_0;
	wire w_dff_B_EK6QoiuF7_0;
	wire w_dff_B_0sPcfCEm5_0;
	wire w_dff_B_j74OIgf71_0;
	wire w_dff_B_giK3ZfKT3_0;
	wire w_dff_B_RqpnAtEb0_0;
	wire w_dff_B_RQQx7A414_0;
	wire w_dff_B_SCOroRu62_0;
	wire w_dff_B_2AT6RE5v8_0;
	wire w_dff_B_9GLbvQK51_0;
	wire w_dff_B_94ri8je74_0;
	wire w_dff_B_GHsgX6uq7_0;
	wire w_dff_B_9jQGw9qS3_0;
	wire w_dff_B_vRSFmdnY9_0;
	wire w_dff_B_0AFXUI3J1_0;
	wire w_dff_B_YbThWPGE9_0;
	wire w_dff_B_1JJ7VEFJ3_0;
	wire w_dff_B_ph4tuA5o9_0;
	wire w_dff_B_PXzo0FXR5_0;
	wire w_dff_B_EI6f7HZW0_0;
	wire w_dff_B_x4x6t1UZ5_0;
	wire w_dff_B_WQQyaq1I0_0;
	wire w_dff_B_LJlHrdKh4_0;
	wire w_dff_B_zpJzrBeX1_0;
	wire w_dff_B_w2OrBOlf7_0;
	wire w_dff_B_MLPgA7JX5_0;
	wire w_dff_B_PPrC5dsk9_0;
	wire w_dff_B_6E3PsTwz7_0;
	wire w_dff_B_MrDsvF7h6_0;
	wire w_dff_B_r5NccNIR1_0;
	wire w_dff_B_E4MrUu1v7_0;
	wire w_dff_B_nW1tMMwR7_0;
	wire w_dff_B_6RU7Wz3s6_0;
	wire w_dff_B_FBdmNrEp5_0;
	wire w_dff_B_dQqps2ge4_0;
	wire w_dff_B_u9VRLZr66_0;
	wire w_dff_B_P5Whr83Q3_0;
	wire w_dff_B_I4nuT0x68_0;
	wire w_dff_B_5BHPhDaZ7_0;
	wire w_dff_B_NZu8twoZ1_0;
	wire w_dff_B_s825yrPp4_0;
	wire w_dff_B_Z3uSCLx70_0;
	wire w_dff_B_g2A2f35Z6_0;
	wire w_dff_B_L36zlbqn7_0;
	wire w_dff_B_sFPFdYnj1_0;
	wire w_dff_B_uRJN2Z1S1_0;
	wire w_dff_B_UnriJoaA0_0;
	wire w_dff_B_V1rzDvpI3_0;
	wire w_dff_B_gbFJPRZS9_0;
	wire w_dff_B_r7owaA1L1_0;
	wire w_dff_B_NfOxH3mi8_0;
	wire w_dff_B_e57zDC3p4_0;
	wire w_dff_B_xiGkzxK49_0;
	wire w_dff_B_Jx6Mo8Vf4_0;
	wire w_dff_B_QeyU41Fr2_0;
	wire w_dff_B_Jo71CWFb7_0;
	wire w_dff_B_NMNHRPtb6_0;
	wire w_dff_B_lZIL4XvH3_0;
	wire w_dff_B_NQkDBRaw2_0;
	wire w_dff_B_wTQtsp8q0_0;
	wire w_dff_B_FD61d4J13_0;
	wire w_dff_B_xH71X5T02_0;
	wire w_dff_B_iOAzKUIi9_0;
	wire w_dff_B_mSkku9xs7_0;
	wire w_dff_B_AvPJCngU7_0;
	wire w_dff_B_yX0J0icS5_0;
	wire w_dff_B_a6NzBdXb7_0;
	wire w_dff_B_HdgOaw0K7_0;
	wire w_dff_B_FEODvdGk4_0;
	wire w_dff_B_FWlKx7Og0_0;
	wire w_dff_B_oksCqqwa4_0;
	wire w_dff_B_FCNovqwK4_0;
	wire w_dff_B_pCzqQPjj4_0;
	wire w_dff_B_20WcSLIP3_0;
	wire w_dff_B_h46I3nSG5_0;
	wire w_dff_B_gFNBuQyl4_0;
	wire w_dff_B_vqACgTsP6_0;
	wire w_dff_B_ifVNfQGj9_0;
	wire w_dff_B_b1SK9OI79_0;
	wire w_dff_B_aXx2AjZE0_0;
	wire w_dff_B_ISKEB67Q8_0;
	wire w_dff_B_rkRCeR1a7_0;
	wire w_dff_B_xW2c1SZ52_0;
	wire w_dff_B_nf3ri1wv4_0;
	wire w_dff_B_vF8SRzO08_0;
	wire w_dff_B_Ib2y6we34_0;
	wire w_dff_B_qnn6UrAm7_0;
	wire w_dff_B_1Va83HTI3_0;
	wire w_dff_B_m1DBBFnk4_0;
	wire w_dff_B_JePJUlNE8_0;
	wire w_dff_B_paCFAH7p6_0;
	wire w_dff_B_ZyYlB3Gf4_0;
	wire w_dff_B_BL0604YI1_0;
	wire w_dff_B_wQwXiO6k4_0;
	wire w_dff_B_mOc2EWeS7_0;
	wire w_dff_B_qg03r9Uq4_0;
	wire w_dff_B_dEPqaaQ91_0;
	wire w_dff_B_amyu1Ebk7_0;
	wire w_dff_B_oAZR17Pe4_0;
	wire w_dff_B_sXxPyr587_0;
	wire w_dff_B_K6HNtwHg0_0;
	wire w_dff_B_3orl7EEY8_0;
	wire w_dff_B_1YlJJ1RB6_0;
	wire w_dff_B_H4NY58EE0_0;
	wire w_dff_B_4mHE5FKx4_0;
	wire w_dff_B_YYw0Pgyg2_0;
	wire w_dff_B_Y9kCUqXx3_0;
	wire w_dff_B_Sm7os6q54_0;
	wire w_dff_B_XYV59m5b6_0;
	wire w_dff_B_vTZyJmn24_0;
	wire w_dff_B_qh3LR3EW9_0;
	wire w_dff_B_IBTJoY8s3_0;
	wire w_dff_B_iYBVjVoJ2_0;
	wire w_dff_B_MQB8pzWu9_0;
	wire w_dff_B_7Irxwdwa3_0;
	wire w_dff_B_A4gxXYeT5_0;
	wire w_dff_B_L5vEnBCe4_0;
	wire w_dff_B_kjqlBjnP7_0;
	wire w_dff_B_kdk7rieD3_0;
	wire w_dff_B_pz4y5f0W1_0;
	wire w_dff_B_nFSDgmgh7_0;
	wire w_dff_B_Ln5O11LD0_0;
	wire w_dff_B_gMj7s1Qq5_0;
	wire w_dff_B_AOs9NUAK2_0;
	wire w_dff_B_KqZIl82N4_0;
	wire w_dff_B_lE4zQQav5_0;
	wire w_dff_B_4R5fXsur6_0;
	wire w_dff_B_Xwf8NQiK3_0;
	wire w_dff_B_INcZZ9du1_0;
	wire w_dff_B_0ukkx5i97_0;
	wire w_dff_B_ejEwZdAO5_0;
	wire w_dff_B_gNkqF7ye2_0;
	wire w_dff_B_lOExTQCk0_0;
	wire w_dff_B_8ilnO7ao2_0;
	wire w_dff_B_mNhv8NzT0_0;
	wire w_dff_B_Vhsm7z3k9_0;
	wire w_dff_B_x1ZgcNBL8_0;
	wire w_dff_B_785CZbJD3_0;
	wire w_dff_B_NHxNd3fE4_0;
	wire w_dff_B_6oGj6A9X9_0;
	wire w_dff_B_6Ijlp6QV7_0;
	wire w_dff_B_mJqkvpO50_0;
	wire w_dff_B_RyDPoz1Z2_0;
	wire w_dff_B_EXwwDbRq0_0;
	wire w_dff_B_CUGELkob2_0;
	wire w_dff_B_5JXuxMkZ1_0;
	wire w_dff_B_yelkp9xh3_0;
	wire w_dff_B_MpLxlKvI0_0;
	wire w_dff_B_93Ub34Fw2_0;
	wire w_dff_B_kNmC3KVP8_0;
	wire w_dff_B_jZUSvEo03_0;
	wire w_dff_B_twT26NLx5_0;
	wire w_dff_B_ryAdrR3U8_0;
	wire w_dff_B_LnB9CBWC3_0;
	wire w_dff_B_1eFl5wzJ7_0;
	wire w_dff_B_rTyNG8fO2_0;
	wire w_dff_B_sGmwp9Yw9_0;
	wire w_dff_B_A7pKB0Tb8_0;
	wire w_dff_B_BvXOgf6L3_0;
	wire w_dff_B_MKfbWAlu6_0;
	wire w_dff_B_7rcRnx1W1_0;
	wire w_dff_B_cYQt0Qi32_0;
	wire w_dff_B_06iSBwe46_0;
	wire w_dff_B_wGijM75C1_0;
	wire w_dff_B_coNrT10v9_0;
	wire w_dff_B_uQ2KjSqG9_0;
	wire w_dff_B_cnhrdf764_0;
	wire w_dff_B_FVmLi4Tc9_0;
	wire w_dff_B_Sa0d1qbJ5_0;
	wire w_dff_B_7Ks559YV4_0;
	wire w_dff_B_xGLWstaY9_0;
	wire w_dff_B_QpfvsARL4_0;
	wire w_dff_B_30CG8MC89_0;
	wire w_dff_B_9nZW4qVC2_0;
	wire w_dff_B_UcgqJ7WF3_0;
	wire w_dff_B_KA9jg2v29_0;
	wire w_dff_B_YTgPN8Ci2_0;
	wire w_dff_B_iSPnGKGf4_0;
	wire w_dff_B_kZjuT8B68_0;
	wire w_dff_B_nr9LvYBe1_0;
	wire w_dff_B_17IgJkoN9_0;
	wire w_dff_B_LKs6pDE20_0;
	wire w_dff_B_e08V3hhG5_0;
	wire w_dff_B_ODV3X2tf2_0;
	wire w_dff_B_7jqXSN8o0_0;
	wire w_dff_B_zO1C5J2N3_0;
	wire w_dff_B_5vNkDRPz1_0;
	wire w_dff_B_yTDKng3N9_0;
	wire w_dff_B_gbTIqg2C1_0;
	wire w_dff_B_CgfxH41a9_0;
	wire w_dff_B_UW3Tmxwx5_0;
	wire w_dff_B_dAhtKta17_0;
	wire w_dff_B_svBcB5FP3_0;
	wire w_dff_B_VggTW5wC8_0;
	wire w_dff_B_aHBEsBAV9_0;
	wire w_dff_B_W2ekGea47_0;
	wire w_dff_B_pxRZbaAB5_0;
	wire w_dff_B_qKzm8EVx0_0;
	wire w_dff_B_FyKgAO4j8_0;
	wire w_dff_B_0al3Uir41_0;
	wire w_dff_B_U8CT8aKb0_0;
	wire w_dff_B_dwLqq59T8_0;
	wire w_dff_B_16sBN8mU4_0;
	wire w_dff_B_wIM70Lt96_0;
	wire w_dff_B_2Aa4akjp1_0;
	wire w_dff_B_IZLRc0Zq7_0;
	wire w_dff_B_GeiaIhpB2_0;
	wire w_dff_B_uTtxsdDb0_0;
	wire w_dff_B_YZ8kRwrG8_0;
	wire w_dff_B_bjK1uvg36_0;
	wire w_dff_B_Vm1jp9ST2_0;
	wire w_dff_B_1Xpydz3R9_0;
	wire w_dff_B_dIqU6Kl59_0;
	wire w_dff_B_DDZo36eF4_0;
	wire w_dff_B_93bkhjsh6_0;
	wire w_dff_B_YDXpRDLc6_0;
	wire w_dff_B_dkeCP9wb0_0;
	wire w_dff_B_IDIdyPVW1_0;
	wire w_dff_B_oBtENBKi1_0;
	wire w_dff_B_ukpxhzIT7_0;
	wire w_dff_B_ZLlHEj7f4_0;
	wire w_dff_B_cCMrRsyB5_0;
	wire w_dff_B_BHgpK55x7_0;
	wire w_dff_B_ahjKWMYI8_0;
	wire w_dff_B_ah2lFrXF4_0;
	wire w_dff_B_funlZuGw9_0;
	wire w_dff_B_vmV8GutO0_0;
	wire w_dff_B_CxiPEjsM7_0;
	wire w_dff_B_UqH2Lvhu9_0;
	wire w_dff_B_tegk8IxO0_0;
	wire w_dff_B_MfhyKy4s5_0;
	wire w_dff_B_USIgyRKd7_0;
	wire w_dff_B_TAMcDs7j9_0;
	wire w_dff_B_QmzSZcRl3_0;
	wire w_dff_B_YNSKKBuA8_0;
	wire w_dff_B_zoZMDuln1_0;
	wire w_dff_B_nuJIspEI8_0;
	wire w_dff_B_QvridlxU4_0;
	wire w_dff_B_21WICGu52_0;
	wire w_dff_B_4envusfo1_0;
	wire w_dff_B_QDFODqXv1_0;
	wire w_dff_B_5UXlMKaV7_0;
	wire w_dff_B_syJO6H2N9_0;
	wire w_dff_B_DlFk9U231_0;
	wire w_dff_B_zOsfWOV19_0;
	wire w_dff_B_8L6EIg5Q0_0;
	wire w_dff_B_mNOH6bvL0_0;
	wire w_dff_B_X6r5gaHs0_0;
	wire w_dff_B_ay0f40Es1_0;
	wire w_dff_B_aZdeldrI2_0;
	wire w_dff_B_4GGAXCGb2_0;
	wire w_dff_B_cCak4lRB8_0;
	wire w_dff_B_kY4vkloa9_0;
	wire w_dff_B_c1mXWdsp9_0;
	wire w_dff_B_f4L9FMuC6_0;
	wire w_dff_B_QrX5sXIn5_0;
	wire w_dff_B_sLEE0XhA0_0;
	wire w_dff_B_YTVe0hl81_0;
	wire w_dff_B_K7FBMU0B7_0;
	wire w_dff_B_Kh1u1Frr8_0;
	wire w_dff_B_IIZIbszu3_0;
	wire w_dff_B_0OENEO1i0_0;
	wire w_dff_B_nMUnz0Bg4_0;
	wire w_dff_B_OeAAUGJF9_0;
	wire w_dff_B_DjvEXiK80_0;
	wire w_dff_B_xn03Z1tL1_0;
	wire w_dff_B_QJLoltAD1_0;
	wire w_dff_B_Fb8SMVIa3_0;
	wire w_dff_B_P1VHCDv58_0;
	wire w_dff_B_PAFj1S6D1_0;
	wire w_dff_B_N2x4cjw34_0;
	wire w_dff_B_KnV2FWR59_0;
	wire w_dff_B_5kCbERLf3_0;
	wire w_dff_B_3JMxaSLI4_0;
	wire w_dff_B_ojhdoTNr5_0;
	wire w_dff_B_79hYDlnI2_0;
	wire w_dff_B_hv1CnjQo8_0;
	wire w_dff_B_kxzh6M3k2_0;
	wire w_dff_B_Nr5B1aJJ8_0;
	wire w_dff_B_5YtuNvVb7_0;
	wire w_dff_B_fTk6qELK8_0;
	wire w_dff_B_Y9GwHcLj4_0;
	wire w_dff_B_JHsTE69f6_0;
	wire w_dff_B_0yuJfA2i9_0;
	wire w_dff_B_sVYMKFjH8_0;
	wire w_dff_B_boqzDCTa7_0;
	wire w_dff_B_FlQP56M19_0;
	wire w_dff_B_pIvosuE11_0;
	wire w_dff_B_V1P11FnG5_0;
	wire w_dff_B_ZTPMJMoB1_0;
	wire w_dff_B_vsN6OyCu7_0;
	wire w_dff_B_RIiq7q8v4_0;
	wire w_dff_B_xxQqVvOs7_0;
	wire w_dff_B_VGi2UROn2_0;
	wire w_dff_B_LfbFJvMx6_0;
	wire w_dff_B_lzEq9KiS3_0;
	wire w_dff_B_51K0myhB2_0;
	wire w_dff_B_yVjpxSIL5_0;
	wire w_dff_B_u0mSMN5R4_0;
	wire w_dff_B_7Yx8Zfv35_0;
	wire w_dff_B_Edmle6YN9_0;
	wire w_dff_B_jh9DrEGX3_0;
	wire w_dff_B_uGz6KgcW3_0;
	wire w_dff_B_y4oDZyQ10_0;
	wire w_dff_B_TDBOi6gD3_0;
	wire w_dff_B_XvVdIYiY5_0;
	wire w_dff_B_EPxaUYP49_0;
	wire w_dff_B_irRoFLoY9_0;
	wire w_dff_B_EECg9nd90_0;
	wire w_dff_B_VgEzxSYs5_0;
	wire w_dff_B_7tkvVyl15_0;
	wire w_dff_B_aBm5XtYk9_0;
	wire w_dff_B_Go4FIk7g5_0;
	wire w_dff_B_RLqf8HKD8_0;
	wire w_dff_B_fvnQjbWl0_0;
	wire w_dff_B_TowlVJ0s3_0;
	wire w_dff_B_DDEY6Udx4_0;
	wire w_dff_B_DY0PG0Dn3_0;
	wire w_dff_B_zfqqG6SZ4_0;
	wire w_dff_B_MiIHbBHu4_0;
	wire w_dff_B_8BzBcwhQ4_0;
	wire w_dff_B_X8rmyqlc4_0;
	wire w_dff_B_8P2FhsK52_0;
	wire w_dff_B_ziWILxZA4_0;
	wire w_dff_B_jJoiKGuQ9_0;
	wire w_dff_B_sERyS6cS0_0;
	wire w_dff_B_7wHWZ19s7_0;
	wire w_dff_B_E2pvJraB9_0;
	wire w_dff_B_tHF5p0PX1_0;
	wire w_dff_B_ikvCzPGE3_0;
	wire w_dff_B_uTbkv3wM3_0;
	wire w_dff_B_nCrOTjUj5_0;
	wire w_dff_B_dWG8H5mb1_0;
	wire w_dff_B_FRzK9OWb5_0;
	wire w_dff_B_rG2duiSU8_0;
	wire w_dff_B_52EbAhTZ8_0;
	wire w_dff_B_iZ8uguWo3_0;
	wire w_dff_B_gHq1mxHV0_0;
	wire w_dff_B_JXVqcLXq8_0;
	wire w_dff_B_FJxIsRPF3_0;
	wire w_dff_B_mtzEfBpI2_0;
	wire w_dff_B_Ek0fZKhM6_0;
	wire w_dff_B_MFgqODb72_0;
	wire w_dff_B_E9BiMMfI4_0;
	wire w_dff_B_Z2B8rynr4_0;
	wire w_dff_B_qmjaMPIw1_0;
	wire w_dff_B_ECrHf2zC6_0;
	wire w_dff_B_N9Kjlmw54_0;
	wire w_dff_B_n9mxIqXi0_0;
	wire w_dff_B_EyMGRDZg7_0;
	wire w_dff_B_xU0f3KRl2_0;
	wire w_dff_B_3wEfpDUe2_0;
	wire w_dff_B_j2hspalA7_0;
	wire w_dff_B_8MbY1Ins3_0;
	wire w_dff_B_C58MuJw33_0;
	wire w_dff_B_it9OyEN43_0;
	wire w_dff_B_z1yQvdZP1_0;
	wire w_dff_B_2fj4AdYc9_0;
	wire w_dff_B_mZYvTbuO2_0;
	wire w_dff_B_hyCaKxBJ1_0;
	wire w_dff_B_yF0xLxvP5_0;
	wire w_dff_B_oSekbLOH3_0;
	wire w_dff_B_h5XniCCh9_0;
	wire w_dff_B_F36HbM4L5_0;
	wire w_dff_B_8jbe1RDh6_0;
	wire w_dff_B_MBsrpKVZ5_0;
	wire w_dff_B_No3w8VlE4_0;
	wire w_dff_B_iTvkgpvC3_0;
	wire w_dff_B_Q6i39hrm5_0;
	wire w_dff_B_jCPROOyD2_0;
	wire w_dff_B_Fb065wS42_0;
	wire w_dff_B_yX0WWuD12_0;
	wire w_dff_B_4OnC4kUA0_0;
	wire w_dff_B_NmIgjnUJ4_0;
	wire w_dff_B_9ffK5bGL2_0;
	wire w_dff_B_k6IMr95z9_0;
	wire w_dff_B_bJdwZxlZ6_0;
	wire w_dff_B_uIoZfzIv8_0;
	wire w_dff_B_aH30KB3z9_0;
	wire w_dff_B_lHzUY87g9_0;
	wire w_dff_B_KUCqu5vt6_0;
	wire w_dff_B_vd20wg4n1_0;
	wire w_dff_B_cNHPUzQw7_0;
	wire w_dff_B_EvEo9Pkn7_0;
	wire w_dff_B_HWib5OwB6_0;
	wire w_dff_B_lsQWPwDm6_0;
	wire w_dff_B_Fyj2NwWY0_0;
	wire w_dff_B_MaksMQu45_0;
	wire w_dff_B_tiLy5M3X9_0;
	wire w_dff_B_rEqIzkkt0_0;
	wire w_dff_B_UbiNwkFQ5_0;
	wire w_dff_B_fLIkzIlP5_0;
	wire w_dff_B_GKbXsgKF8_0;
	wire w_dff_B_Way09Ywm0_0;
	wire w_dff_B_KUii6ckP9_0;
	wire w_dff_B_646MqpjW3_0;
	wire w_dff_B_w3lR9CXB0_0;
	wire w_dff_B_fm8cLBpR6_0;
	wire w_dff_B_ju8l2vfT0_0;
	wire w_dff_B_JxWKhrsd3_0;
	wire w_dff_B_K8KR1v0h0_0;
	wire w_dff_B_UvqYw03W5_0;
	wire w_dff_B_h9uCuHdf8_0;
	wire w_dff_B_joHR6gXx1_0;
	wire w_dff_B_LJCweJus4_0;
	wire w_dff_B_6kHkPDp78_0;
	wire w_dff_B_yQxSAM1L6_0;
	wire w_dff_B_PhCI8RNz2_0;
	wire w_dff_B_SwtgvfxI4_0;
	wire w_dff_B_Ek657jhd9_0;
	wire w_dff_B_6vcnl2iQ6_0;
	wire w_dff_B_5SLe2eNO3_0;
	wire w_dff_B_CFDwVCYX8_0;
	wire w_dff_B_8XovsaSy3_0;
	wire w_dff_B_Lb1t9QhG6_0;
	wire w_dff_B_1bIKvqNO8_0;
	wire w_dff_B_HXQTeHnK9_0;
	wire w_dff_B_9xeGihgn1_0;
	wire w_dff_B_rqAiToFs3_0;
	wire w_dff_B_30v9Th3L5_0;
	wire w_dff_B_a1GkOzxU4_0;
	wire w_dff_B_sqLqSx5U8_0;
	wire w_dff_B_6AmJ106J1_0;
	wire w_dff_B_NwqyJ2OD2_0;
	wire w_dff_B_yEk5ecGq2_0;
	wire w_dff_B_AoKGARec0_0;
	wire w_dff_B_mrT4pSGv1_0;
	wire w_dff_B_b1mSl9DT0_0;
	wire w_dff_B_goXRnpUM6_0;
	wire w_dff_B_bVBNA7wK3_0;
	wire w_dff_B_R4Xup1eB1_0;
	wire w_dff_B_XdzVqCzX3_0;
	wire w_dff_B_HBiiIxZ67_0;
	wire w_dff_B_Kum9dh4r7_0;
	wire w_dff_B_u55DL7ub0_0;
	wire w_dff_B_GohZT36D3_0;
	wire w_dff_B_HvEYUVtu8_0;
	wire w_dff_B_zDTbwalz8_0;
	wire w_dff_B_DgA6ozJq1_0;
	wire w_dff_B_7b6bYiHg5_0;
	wire w_dff_B_zkA0H2TJ0_0;
	wire w_dff_B_7A5a7cYa4_0;
	wire w_dff_B_B0dLc4Kb9_0;
	wire w_dff_B_geok2ODD5_0;
	wire w_dff_B_TnBIMtmU7_0;
	wire w_dff_B_JktU5inu7_0;
	wire w_dff_B_Jv2UVd6g1_0;
	wire w_dff_B_VkFRakZ91_0;
	wire w_dff_B_xW0kb1In4_0;
	wire w_dff_B_TsWlvTGw2_0;
	wire w_dff_B_ghueHGkG3_0;
	wire w_dff_B_csVN0p779_0;
	wire w_dff_B_Fr2XhxCO7_0;
	wire w_dff_B_CY5I6Dgz8_0;
	wire w_dff_B_pmmZEC6D4_0;
	wire w_dff_B_WXt3uY0G0_0;
	wire w_dff_B_A0YB9WqP1_0;
	wire w_dff_B_IlM6eD5D1_0;
	wire w_dff_B_lIwnggMu4_0;
	wire w_dff_B_c7NH46Op4_0;
	wire w_dff_B_jrvJuDlt4_0;
	wire w_dff_B_Ah0VBcm17_0;
	wire w_dff_B_5orD6xrr6_0;
	wire w_dff_B_JMSRNqWX5_0;
	wire w_dff_B_1foiTy730_0;
	wire w_dff_B_VrOceuR77_0;
	wire w_dff_B_lsMFHzPE9_0;
	wire w_dff_B_pUFufnay7_0;
	wire w_dff_B_EUX6sfvJ6_0;
	wire w_dff_B_iG9NtK4K1_0;
	wire w_dff_B_pv3sBp5K2_0;
	wire w_dff_B_gjtWZT8u6_0;
	wire w_dff_B_U3Z9hAzM4_0;
	wire w_dff_B_BoShgiUc7_0;
	wire w_dff_B_c9yTcfM50_0;
	wire w_dff_B_hD1e3CLC0_0;
	wire w_dff_B_XBFHlLzf8_0;
	wire w_dff_B_bR8CSXxS3_0;
	wire w_dff_B_RYBOLw7n3_0;
	wire w_dff_B_0T3Nbega6_0;
	wire w_dff_B_VB5P8UTL5_0;
	wire w_dff_B_GePgwC936_0;
	wire w_dff_B_ukDCK8Vf6_0;
	wire w_dff_B_KAGeyIyS6_0;
	wire w_dff_B_QMxEWjXT3_0;
	wire w_dff_B_1DKQEo9i2_0;
	wire w_dff_B_GIOxWv5h3_0;
	wire w_dff_B_FUPMUI5t3_0;
	wire w_dff_B_lpcqvB2h3_0;
	wire w_dff_B_UUCqwFXR2_0;
	wire w_dff_B_PkJzX0Ml5_0;
	wire w_dff_B_CWeJCeTY4_0;
	wire w_dff_B_2A7qYmVr9_0;
	wire w_dff_B_Yx54bmGe0_0;
	wire w_dff_B_99vr0vfs6_0;
	wire w_dff_B_LWpVHPFi6_0;
	wire w_dff_B_LtqzSqf73_0;
	wire w_dff_B_nd50uFT93_0;
	wire w_dff_B_Sq60IGAl3_0;
	wire w_dff_B_WHj74Hgr6_0;
	wire w_dff_B_NKp9N87a6_0;
	wire w_dff_B_KqURzsvA4_0;
	wire w_dff_B_XHCHRC666_0;
	wire w_dff_B_luqQTiZz7_0;
	wire w_dff_B_aQrUFAWZ0_0;
	wire w_dff_B_vguzv9tU7_0;
	wire w_dff_B_USkauRet9_0;
	wire w_dff_B_Ugfr3I697_0;
	wire w_dff_B_8LO3tYGd8_0;
	wire w_dff_B_1Z9ckb7l5_0;
	wire w_dff_B_bc79WY4J3_0;
	wire w_dff_B_1Yuc01Af7_0;
	wire w_dff_B_zsrHNdGQ9_0;
	wire w_dff_B_63BceWwP8_0;
	wire w_dff_B_DyEX1x7T5_0;
	wire w_dff_B_oIFEkwfl4_0;
	wire w_dff_B_hK28HObY6_0;
	wire w_dff_B_73y1Gfaz3_0;
	wire w_dff_B_hqH6fwBA0_0;
	wire w_dff_B_CvrIixkZ0_0;
	wire w_dff_B_UWyGvAfr4_0;
	wire w_dff_B_becLxMS63_0;
	wire w_dff_B_vlsL3pMh2_0;
	wire w_dff_B_KApHAKxm1_0;
	wire w_dff_B_mmkX4I9b6_0;
	wire w_dff_B_EcdDGgM70_0;
	wire w_dff_B_y1qEE1vH6_0;
	wire w_dff_B_huZcUXJl1_0;
	wire w_dff_B_7ys95aUX5_0;
	wire w_dff_B_WOH18U781_0;
	wire w_dff_B_DwoezAJJ7_0;
	wire w_dff_B_gDS4yW2p0_0;
	wire w_dff_B_I0xZM2qy9_0;
	wire w_dff_B_LaiBGMm09_0;
	wire w_dff_B_p7xA06Kb4_0;
	wire w_dff_B_hwR3UXWw2_0;
	wire w_dff_B_tPJbIVE25_0;
	wire w_dff_B_98rxaBb90_0;
	wire w_dff_B_15IQasa12_0;
	wire w_dff_B_FdJzxjK20_0;
	wire w_dff_B_d3OJeoQD5_0;
	wire w_dff_B_mOyQaOUP6_0;
	wire w_dff_B_FMC2ALGB0_0;
	wire w_dff_B_J5hZN5sU2_0;
	wire w_dff_B_swrFznVd2_0;
	wire w_dff_B_V7Aqu1az5_0;
	wire w_dff_B_yyhY2Yw85_0;
	wire w_dff_B_Su83XJaR1_0;
	wire w_dff_B_CFUw9yfu4_0;
	wire w_dff_B_4pKocEiJ6_0;
	wire w_dff_B_FhqjgeKJ9_0;
	wire w_dff_B_Cz8B2XOQ2_0;
	wire w_dff_B_yZtfL8ho2_0;
	wire w_dff_B_AMRUMcIZ0_0;
	wire w_dff_B_0O8dBAK65_0;
	wire w_dff_B_eeSDeSIQ4_0;
	wire w_dff_B_AieIUgmS7_0;
	wire w_dff_B_L0WXBmqO4_0;
	wire w_dff_B_rKpeCilG4_0;
	wire w_dff_B_aoDqEjFW7_0;
	wire w_dff_B_BOz2XnWz8_0;
	wire w_dff_B_uLflUQtv0_0;
	wire w_dff_B_qpYuQQtv1_0;
	wire w_dff_B_sgXW8qAx8_0;
	wire w_dff_B_eSjjEMdr2_0;
	wire w_dff_B_OHrR9IVm0_0;
	wire w_dff_B_OfMJidXT3_0;
	wire w_dff_B_MOLD35Y74_0;
	wire w_dff_B_A7lgqtib8_0;
	wire w_dff_B_IgoGkVoq8_0;
	wire w_dff_B_5i4re2bm3_0;
	wire w_dff_B_VPrzomyO6_0;
	wire w_dff_B_p17P0aA03_0;
	wire w_dff_B_xsvbUtpc6_0;
	wire w_dff_B_em69dLqe0_0;
	wire w_dff_B_Gl0rW1Qn8_0;
	wire w_dff_B_PhuHTBhY4_0;
	wire w_dff_B_rP8ne3da3_0;
	wire w_dff_B_ERrrdDkU6_0;
	wire w_dff_B_qZ2VEzT82_0;
	wire w_dff_B_4HMDwuKd5_0;
	wire w_dff_B_S1Kc1tjD1_0;
	wire w_dff_B_P6SFdFZB3_0;
	wire w_dff_B_OMmmPeWO5_0;
	wire w_dff_B_bfp2AXte5_0;
	wire w_dff_B_ux7t2bqd3_0;
	wire w_dff_B_oJTqfavZ4_0;
	wire w_dff_B_sDKk6S8e7_0;
	wire w_dff_B_OfW4Jghg9_0;
	wire w_dff_B_2pB8xujb7_0;
	wire w_dff_B_pz7zkUlu3_0;
	wire w_dff_B_SROJpiDS2_0;
	wire w_dff_B_THjixmin7_0;
	wire w_dff_B_4af4m4Ov4_0;
	wire w_dff_B_6S96Z7S51_0;
	wire w_dff_B_i6YeeLqi1_0;
	wire w_dff_B_4PV1JVpJ3_0;
	wire w_dff_B_UGsB0gXX0_0;
	wire w_dff_B_g3aasNoc1_0;
	wire w_dff_B_4FAoKlbW9_0;
	wire w_dff_B_zkkXAhQn5_0;
	wire w_dff_B_OLxbQuH34_0;
	wire w_dff_B_KznebfxW6_0;
	wire w_dff_B_aRBAKbmy4_0;
	wire w_dff_B_bNmyuJte7_0;
	wire w_dff_B_wzlBs0G79_0;
	wire w_dff_B_7X1cEWH71_0;
	wire w_dff_B_Gi5pgYEa2_0;
	wire w_dff_B_uaSauKIB2_0;
	wire w_dff_B_EB2vTghp0_0;
	wire w_dff_B_3V14pkZT0_0;
	wire w_dff_B_SloTGfGm5_0;
	wire w_dff_B_YVnrL50z0_0;
	wire w_dff_B_2IlKruwx9_0;
	wire w_dff_B_kVoKSRtF3_0;
	wire w_dff_B_Zb3Aui4E2_0;
	wire w_dff_B_XIBVtP5T9_0;
	wire w_dff_B_hEIbsiQx7_0;
	wire w_dff_B_vVped8t61_0;
	wire w_dff_B_ZkDUw77u5_0;
	wire w_dff_B_MvzMNG2t9_0;
	wire w_dff_B_Ail5uBBE2_0;
	wire w_dff_B_qV1IbSDy5_0;
	wire w_dff_B_Or6PBY1k3_0;
	wire w_dff_B_gLQI5EyF4_0;
	wire w_dff_B_VUI7xP7N1_0;
	wire w_dff_B_ZrWmxTbZ5_0;
	wire w_dff_B_rKXDGhNW6_0;
	wire w_dff_B_CVSJZ2iq8_0;
	wire w_dff_B_rC8u444R3_0;
	wire w_dff_B_cL6aYRW21_0;
	wire w_dff_B_OGDHVhHV9_0;
	wire w_dff_B_btyvR2yp6_0;
	wire w_dff_B_X3Y9Qcy22_0;
	wire w_dff_B_JZJLzT7R1_0;
	wire w_dff_B_AJ7dbya17_0;
	wire w_dff_B_v3UYbTMW8_0;
	wire w_dff_B_DCkNC7O52_0;
	wire w_dff_B_ki1KXNyQ2_0;
	wire w_dff_B_G0kFSLcc6_0;
	wire w_dff_B_f8cyZzge4_0;
	wire w_dff_B_EzaRmUX02_0;
	wire w_dff_B_0f8mKj3l1_0;
	wire w_dff_B_kwHn0N3C3_0;
	wire w_dff_B_GH3kbN1A4_0;
	wire w_dff_B_Up5Zwngc3_0;
	wire w_dff_B_3M6pJRuC8_0;
	wire w_dff_B_1HnMSGBx7_0;
	wire w_dff_B_iTnGCJcI5_0;
	wire w_dff_B_J8qORiw16_0;
	wire w_dff_B_act0EzCl1_0;
	wire w_dff_B_MPgarCf60_0;
	wire w_dff_B_Zr5e05Kd9_0;
	wire w_dff_B_w7QyZyJX4_0;
	wire w_dff_B_VQl2595z1_0;
	wire w_dff_B_zGWPKchG6_0;
	wire w_dff_B_B4VkixQz7_0;
	wire w_dff_B_AZZAoUlg3_0;
	wire w_dff_B_fcLtakTq9_0;
	wire w_dff_B_GcsI27qI6_0;
	wire w_dff_B_79uVL9sZ7_0;
	wire w_dff_B_io6zSyI37_0;
	wire w_dff_B_ct3BczfG9_0;
	wire w_dff_B_NnkrXpG68_0;
	wire w_dff_B_82bDnHis2_0;
	wire w_dff_B_m7a7MgSH4_0;
	wire w_dff_B_eMbb14EB4_0;
	wire w_dff_B_AJnunAIe4_0;
	wire w_dff_B_mnp17btZ2_0;
	wire w_dff_B_Zd9dDlEE4_0;
	wire w_dff_B_24QlirJ28_0;
	wire w_dff_B_p5IueDTz1_0;
	wire w_dff_B_vbTSAZ3x6_0;
	wire w_dff_B_FmpoJySX5_0;
	wire w_dff_B_6clVDe9u5_0;
	wire w_dff_B_5TRClnVL4_0;
	wire w_dff_B_2MPg8mNX6_0;
	wire w_dff_B_ipLr3u053_0;
	wire w_dff_B_SP6w6syZ5_0;
	wire w_dff_B_yk90ZYBF7_0;
	wire w_dff_B_6WPlQnjn3_0;
	wire w_dff_B_3Psgfeor4_0;
	wire w_dff_B_GzQJe2hd3_0;
	wire w_dff_B_fFgdS6yr2_0;
	wire w_dff_B_wCqYeAoU5_0;
	wire w_dff_B_2QkoEW2i9_0;
	wire w_dff_B_NEl2t2WK5_0;
	wire w_dff_B_jkdSfD8o0_0;
	wire w_dff_B_d9YLOmDB7_0;
	wire w_dff_B_DhOwyyt05_0;
	wire w_dff_B_W0UFrXYB9_0;
	wire w_dff_B_J89MJakF3_0;
	wire w_dff_B_uENGzOBh2_0;
	wire w_dff_B_Ep7ZbnL90_0;
	wire w_dff_B_MsEOaw3U3_0;
	wire w_dff_B_Z1RMHlHD6_0;
	wire w_dff_B_BNmrJpzO8_0;
	wire w_dff_B_1mhdemTw3_0;
	wire w_dff_B_8DX3k4f20_0;
	wire w_dff_B_acAylcrc9_0;
	wire w_dff_B_setQDUl23_0;
	wire w_dff_B_TC9Jipj27_0;
	wire w_dff_B_9ufmnTMV7_0;
	wire w_dff_B_DMX1dXDT5_0;
	wire w_dff_B_1bnbnxWi5_0;
	wire w_dff_B_hYcRO49R2_0;
	wire w_dff_B_QoNs79Ag6_0;
	wire w_dff_B_7CXgmlU11_0;
	wire w_dff_B_O3LNg3lQ4_0;
	wire w_dff_B_zXATzSmg4_0;
	wire w_dff_B_DbHnkhoM2_0;
	wire w_dff_B_to6Tc7fS8_0;
	wire w_dff_B_r3egGGxX3_0;
	wire w_dff_B_ZHEFBFy70_0;
	wire w_dff_B_LGU3LcRJ3_0;
	wire w_dff_B_BCCiiD521_0;
	wire w_dff_B_BJ5MHOmb2_0;
	wire w_dff_B_EiHuVkh28_0;
	wire w_dff_B_9YBHhiIi4_0;
	wire w_dff_B_EzEAjWrM2_0;
	wire w_dff_B_Jt2KN0hA3_0;
	wire w_dff_B_W4sBaM5H5_0;
	wire w_dff_B_IIOII2UC9_0;
	wire w_dff_B_JCf1MSee8_0;
	wire w_dff_B_Xi9YM6Iy1_0;
	wire w_dff_B_Sg4YK8vp2_0;
	wire w_dff_B_0UMBkUdK0_0;
	wire w_dff_B_YX7CqXs84_0;
	wire w_dff_B_w9rZFh0P2_0;
	wire w_dff_B_nRU76yD61_0;
	wire w_dff_B_7QoyaaUP6_0;
	wire w_dff_B_xUbN0nya1_0;
	wire w_dff_B_2ioswjf45_0;
	wire w_dff_B_vKRXIBIi8_0;
	wire w_dff_B_0BiWx5La1_0;
	wire w_dff_B_429sELnG5_0;
	wire w_dff_B_B8sF3QoZ6_0;
	wire w_dff_B_VVKliftS9_0;
	wire w_dff_B_hC77Gjo20_0;
	wire w_dff_B_rdLexDQC7_0;
	wire w_dff_B_Kab0bn8L2_0;
	wire w_dff_B_yP51ITwX7_0;
	wire w_dff_B_73RWRYjg9_0;
	wire w_dff_B_D42ptgaw7_0;
	wire w_dff_B_l8pJKvwU4_0;
	wire w_dff_B_KbOYTM4W4_0;
	wire w_dff_B_udGSE7zz4_0;
	wire w_dff_B_eBtTxwtr5_0;
	wire w_dff_B_oJ7lkHKB1_0;
	wire w_dff_B_pYbb9aiH4_0;
	wire w_dff_B_tsHHG2pn2_0;
	wire w_dff_B_1GjYhWup4_0;
	wire w_dff_B_2va0z3ho3_0;
	wire w_dff_B_ZzbnFaOZ9_0;
	wire w_dff_B_Uoor99ov9_0;
	wire w_dff_B_mwaZx1Pw1_0;
	wire w_dff_B_KE9Wtkoq3_0;
	wire w_dff_B_neOY6BFx7_0;
	wire w_dff_B_LXqYXlFk4_0;
	wire w_dff_B_crEd0d0B0_0;
	wire w_dff_B_JVQanGuL2_0;
	wire w_dff_B_87ABA4220_0;
	wire w_dff_B_lWIE4kdJ0_0;
	wire w_dff_B_uUxQQKLa1_0;
	wire w_dff_B_djJxNpry8_0;
	wire w_dff_B_vM1UBh3N6_0;
	wire w_dff_B_bkQrWo0p1_0;
	wire w_dff_B_zLM4uuE45_0;
	wire w_dff_B_bOWF5lqG0_0;
	wire w_dff_B_LikD3aIF0_0;
	wire w_dff_B_zM8ZWNiA6_0;
	wire w_dff_B_bHdvkmT64_0;
	wire w_dff_B_vcWeeyN54_0;
	wire w_dff_B_4JebWuIn6_0;
	wire w_dff_B_FdzOElnO1_0;
	wire w_dff_B_oJrZnA5B5_0;
	wire w_dff_B_KuaKaXw61_0;
	wire w_dff_B_7QB61Y7k8_0;
	wire w_dff_B_6Zl32GTW5_0;
	wire w_dff_B_WiI8Ey2i9_0;
	wire w_dff_B_Bn0J8M762_0;
	wire w_dff_B_F93XNt5i5_0;
	wire w_dff_B_FXkoKMnn3_0;
	wire w_dff_B_7MmMkRQb7_0;
	wire w_dff_B_tmhoApgT1_0;
	wire w_dff_B_IaZj5f5E6_0;
	wire w_dff_B_MdaEq8cC1_0;
	wire w_dff_B_omNQpwgx2_0;
	wire w_dff_B_OMXlPSJV4_0;
	wire w_dff_B_DFUJyOSU3_0;
	wire w_dff_B_XhhwdUIa1_0;
	wire w_dff_B_wvHW04T62_0;
	wire w_dff_B_qWTm3oSy6_0;
	wire w_dff_B_fCIlhNPU1_0;
	wire w_dff_B_81eeMq5X9_0;
	wire w_dff_B_xnChlfi34_0;
	wire w_dff_B_Bjcvqyle8_0;
	wire w_dff_B_KAcvpLMI0_0;
	wire w_dff_B_c4IxKS9W8_0;
	wire w_dff_B_I6CjZlZ28_0;
	wire w_dff_B_D1jGAaK66_0;
	wire w_dff_B_zDv66KOB8_0;
	wire w_dff_B_GGYLst9G5_0;
	wire w_dff_B_bfxEIaek1_0;
	wire w_dff_B_8UT2cDNx0_0;
	wire w_dff_B_eA4AblRc4_0;
	wire w_dff_B_YXCUUzBE3_0;
	wire w_dff_B_RSXaTjSB4_0;
	wire w_dff_B_is0svj5R6_0;
	wire w_dff_B_HYzHSGIL5_0;
	wire w_dff_B_8axesWXT6_0;
	wire w_dff_B_4KtXTPat7_0;
	wire w_dff_B_qVdVgnM63_0;
	wire w_dff_B_mD6PHSB68_0;
	wire w_dff_B_kF0Imev28_0;
	wire w_dff_B_x7L4bWiu2_0;
	wire w_dff_B_DxTf15X22_0;
	wire w_dff_B_Spsqco3H4_0;
	wire w_dff_B_IgtOKXGT2_0;
	wire w_dff_B_qEgsXsUg9_0;
	wire w_dff_B_ov6Io3DL5_0;
	wire w_dff_B_iYpslwJ14_0;
	wire w_dff_B_BOwiWPIo6_0;
	wire w_dff_B_z94sYFJN8_0;
	wire w_dff_B_KfH6SYsc1_0;
	wire w_dff_B_IWC8jTjB4_0;
	wire w_dff_B_trIvCV9t3_0;
	wire w_dff_B_7X5463831_0;
	wire w_dff_B_snlhun002_0;
	wire w_dff_B_Fc8BozXS5_0;
	wire w_dff_B_znfAO9BJ3_0;
	wire w_dff_B_CcKhd9Sx9_0;
	wire w_dff_B_nprRhfRi8_0;
	wire w_dff_B_9AY16yQp7_0;
	wire w_dff_B_dHVmP7kB3_0;
	wire w_dff_B_uQCRUEsm3_0;
	wire w_dff_B_h1gGIhqh6_0;
	wire w_dff_B_iuEXXVGa8_0;
	wire w_dff_B_iwr7AWA66_0;
	wire w_dff_B_yAqiSVRh4_0;
	wire w_dff_B_uNf2OqZk3_0;
	wire w_dff_B_9HttA2JE1_0;
	wire w_dff_B_00ffjm2E0_0;
	wire w_dff_B_8bUDF9ix8_0;
	wire w_dff_B_KfswDMz35_0;
	wire w_dff_B_3ApTX3548_0;
	wire w_dff_B_y2TWio1J2_0;
	wire w_dff_B_xmyoRDTp1_0;
	wire w_dff_B_UijIED8f2_0;
	wire w_dff_B_KmQb0IHD9_0;
	wire w_dff_B_11gI7d5m0_0;
	wire w_dff_B_QsOjsc4Y2_0;
	wire w_dff_B_LTjmnrJO1_0;
	wire w_dff_B_zSrSj8Fp6_0;
	wire w_dff_B_DXl8iyb68_0;
	wire w_dff_B_53UoUw6A6_0;
	wire w_dff_B_9Q7JBnMj2_0;
	wire w_dff_B_MPkAfAVI9_0;
	wire w_dff_B_RjhTeT1N1_0;
	wire w_dff_B_rpzL0iEf5_0;
	wire w_dff_B_jtfNxXVo2_0;
	wire w_dff_B_epiKvRPA7_0;
	wire w_dff_B_NYAa6HbO8_0;
	wire w_dff_B_wrmKRBuO2_0;
	wire w_dff_B_epJUvQwS0_0;
	wire w_dff_B_UkRbA1kW0_0;
	wire w_dff_B_hUiR4VQm3_0;
	wire w_dff_B_eL98MWxO1_0;
	wire w_dff_B_Q4DkU52J5_0;
	wire w_dff_B_YV1gapoO4_0;
	wire w_dff_B_OalLZ1mB6_0;
	wire w_dff_B_7S2EpBCa6_0;
	wire w_dff_B_8DTpE4Zp1_0;
	wire w_dff_B_0Vln8Pqp2_0;
	wire w_dff_B_AdyZIk417_0;
	wire w_dff_B_iiHa9ajV1_0;
	wire w_dff_B_HHDt0loH9_0;
	wire w_dff_B_PCcJpXXW3_0;
	wire w_dff_B_8h4cd8Ej2_0;
	wire w_dff_B_vmtII7zd4_0;
	wire w_dff_B_5GZcVb409_0;
	wire w_dff_B_IuWpCWOI4_0;
	wire w_dff_B_vwhblVu44_0;
	wire w_dff_B_01JVspxS2_0;
	wire w_dff_B_fUUt94jj4_0;
	wire w_dff_B_AMBEo5So0_0;
	wire w_dff_B_GrQU66uW6_0;
	wire w_dff_B_dJ0ONYrp8_0;
	wire w_dff_B_mfVQhXaw7_0;
	wire w_dff_B_ztTZe4VO4_0;
	wire w_dff_B_UdbuoscS3_0;
	wire w_dff_B_qRYVwjpB6_0;
	wire w_dff_B_bI7CO9ur3_0;
	wire w_dff_B_tCIx70BC6_0;
	wire w_dff_B_4X4wSKmW6_0;
	wire w_dff_B_3gUUqtf63_0;
	wire w_dff_B_nUY4KDfq6_0;
	wire w_dff_B_POSGgnGY1_0;
	wire w_dff_B_a0I8Lziu0_0;
	wire w_dff_B_5Y0rdulh0_0;
	wire w_dff_B_VLP4Z1nt7_0;
	wire w_dff_B_5FA1RMFP5_0;
	wire w_dff_B_6SH55aU78_0;
	wire w_dff_B_FeHhwumd3_0;
	wire w_dff_B_As6YPZ1T8_0;
	wire w_dff_B_V85dXJTx9_0;
	wire w_dff_B_lD7eShyX9_0;
	wire w_dff_B_18Z8L0Bs1_0;
	wire w_dff_B_wBWQwLiz3_0;
	wire w_dff_B_XMZ24YTb2_0;
	wire w_dff_B_F7tJJUdp9_0;
	wire w_dff_B_pyH5qzWo2_0;
	wire w_dff_B_m6NqfXbK2_0;
	wire w_dff_B_71KChGh51_0;
	wire w_dff_B_8ADYl05n4_0;
	wire w_dff_B_pFbX0ArR1_0;
	wire w_dff_B_3xJwK9lW5_0;
	wire w_dff_B_F5vtCGLu7_0;
	wire w_dff_B_QF5uRPYv9_0;
	wire w_dff_B_Fxna4I119_0;
	wire w_dff_B_KiAsrvlZ4_0;
	wire w_dff_B_RHqzMPBN8_0;
	wire w_dff_B_C6RKWGWN4_0;
	wire w_dff_B_SGVKhsLi3_0;
	wire w_dff_B_rtGeXwMr4_0;
	wire w_dff_B_vHXhuWGI9_0;
	wire w_dff_B_kensvvsp9_0;
	wire w_dff_B_XKcXItV71_0;
	wire w_dff_B_7yEvBIrM2_0;
	wire w_dff_B_sJo82JNR4_0;
	wire w_dff_B_gAOLVwCc6_0;
	wire w_dff_B_pbsApzcG9_0;
	wire w_dff_B_O5VqGE7U3_0;
	wire w_dff_B_CBJcB2gf8_0;
	wire w_dff_B_NZ2hVoch4_0;
	wire w_dff_B_On6FOcow9_0;
	wire w_dff_B_9rn9yQoh0_0;
	wire w_dff_B_q8f9m24X0_0;
	wire w_dff_B_Sjsq87yN4_0;
	wire w_dff_B_L7HN03dK9_0;
	wire w_dff_B_C4wOqSqZ2_0;
	wire w_dff_B_mHLvCTdP8_0;
	wire w_dff_B_93BSnBvH2_0;
	wire w_dff_B_ty1O9y3B4_0;
	wire w_dff_B_bhcrfqRZ0_0;
	wire w_dff_B_oBStXrSG2_0;
	wire w_dff_B_KkurCbps6_0;
	wire w_dff_B_2Kk6QEAu6_0;
	wire w_dff_B_Jihq6Kvy5_0;
	wire w_dff_B_rn1yAsyk9_0;
	wire w_dff_B_sww4Gs9p2_0;
	wire w_dff_B_sQuyETEw9_0;
	wire w_dff_B_gfYolZw20_0;
	wire w_dff_B_tMeyRfLd1_0;
	wire w_dff_B_qgAHsxex2_0;
	wire w_dff_B_ccFyZxub5_0;
	wire w_dff_B_XpilEKo69_0;
	wire w_dff_B_UyXbQcRM5_0;
	wire w_dff_B_1c7ypbJ28_0;
	wire w_dff_B_quhpEhkV8_0;
	wire w_dff_B_ZPMSWbcO9_0;
	wire w_dff_B_FsO2KXY16_0;
	wire w_dff_B_fK7CgUWz2_0;
	wire w_dff_B_zmt3UkZY0_0;
	wire w_dff_B_jBxAI2UV6_0;
	wire w_dff_B_GgBdXz0U9_0;
	wire w_dff_B_03MzA0Kj3_0;
	wire w_dff_B_LdqzZI305_0;
	wire w_dff_B_o1V6vdcU0_0;
	wire w_dff_B_oo9mbzXF5_0;
	wire w_dff_B_UGdadZeY4_0;
	wire w_dff_B_7DLzRguY7_0;
	wire w_dff_B_yV9B1bcm9_0;
	wire w_dff_B_eqWLG71Y1_0;
	wire w_dff_B_QE3UhFth6_0;
	wire w_dff_B_h6mXwqX92_0;
	wire w_dff_B_HMGpbvyO1_0;
	wire w_dff_B_xBCyy7pN0_0;
	wire w_dff_B_W0K5zfFS9_0;
	wire w_dff_B_WlIzNb8K2_0;
	wire w_dff_B_rfckuJU06_0;
	wire w_dff_B_Eu8pChFF3_0;
	wire w_dff_B_S3pJhBGw0_0;
	wire w_dff_B_ZJUuqh130_0;
	wire w_dff_B_pIrIQHYH5_0;
	wire w_dff_B_ZluC5sUa1_0;
	wire w_dff_B_HWZ6xMrk3_0;
	wire w_dff_B_ZVI1toyV6_0;
	wire w_dff_B_e1ipzYgu1_0;
	wire w_dff_B_7P2MWAGJ5_0;
	wire w_dff_B_eXNMIxO55_0;
	wire w_dff_B_yypIunip2_0;
	wire w_dff_B_Sy7GwzC87_0;
	wire w_dff_B_tw0fiH2D9_0;
	wire w_dff_B_3EYGPgMO0_0;
	wire w_dff_B_9rEkfsRT6_0;
	wire w_dff_B_gKW1k3vP2_0;
	wire w_dff_B_WAKMJgJ61_0;
	wire w_dff_B_9Ci4xdAO5_0;
	wire w_dff_B_iA0KSU5s9_0;
	wire w_dff_B_tC36WRQz7_0;
	wire w_dff_B_oiCHdwmw3_0;
	wire w_dff_B_Yevv8j603_0;
	wire w_dff_B_rGjTU6yF8_0;
	wire w_dff_B_yl0RoV968_0;
	wire w_dff_B_1Z9pjIVe8_0;
	wire w_dff_B_dQiz3B5P5_0;
	wire w_dff_B_eiqSCjH55_0;
	wire w_dff_B_CVwiXj1l3_0;
	wire w_dff_B_06JyOsox7_0;
	wire w_dff_B_oq0Ad0me5_0;
	wire w_dff_B_jMoSSrJl9_0;
	wire w_dff_B_axok3U3t6_0;
	wire w_dff_B_ySucNKrO5_0;
	wire w_dff_B_4ThrRtdN4_0;
	wire w_dff_B_DUZzXQVu2_0;
	wire w_dff_B_okJl0APA3_0;
	wire w_dff_B_2lPoOPl03_0;
	wire w_dff_B_HaoU4eN69_0;
	wire w_dff_B_yj6azYvT2_0;
	wire w_dff_B_Eu2rFSWJ1_0;
	wire w_dff_B_PFeOYQaX8_0;
	wire w_dff_B_vMvenhfX3_0;
	wire w_dff_B_wZ3FJX3c1_0;
	wire w_dff_B_jFOUyfxY2_0;
	wire w_dff_B_MfeaioIt7_0;
	wire w_dff_B_9kRdCrj86_0;
	wire w_dff_B_pwd3PH0a4_0;
	wire w_dff_B_0Jx5mqXQ0_0;
	wire w_dff_B_VUuubfv55_0;
	wire w_dff_B_KFd18uWV7_0;
	wire w_dff_B_K8p4uDlq8_0;
	wire w_dff_B_MxdQpzyM1_0;
	wire w_dff_B_Uxw8tnbp2_0;
	wire w_dff_B_J8jYby6L9_0;
	wire w_dff_B_1hA3Zjco7_0;
	wire w_dff_B_KJK0PAH61_0;
	wire w_dff_B_dJuaSdJh4_0;
	wire w_dff_B_4U8x8mnJ7_0;
	wire w_dff_B_WPojmvGb3_0;
	wire w_dff_B_eX7TXg2U3_0;
	wire w_dff_B_oF2X9Cwx7_0;
	wire w_dff_B_Gy3LbCy64_0;
	wire w_dff_B_LHTXzUl40_0;
	wire w_dff_B_5PUROoBS0_0;
	wire w_dff_B_l7pV1nzR2_0;
	wire w_dff_B_hBR33tVC7_0;
	wire w_dff_B_rxxQYZmA9_0;
	wire w_dff_B_mDYmXbQU0_0;
	wire w_dff_B_mBpp0bFr9_0;
	wire w_dff_B_FjTeiGUe2_0;
	wire w_dff_B_q8d0M6PG0_0;
	wire w_dff_B_B5gUXouM3_0;
	wire w_dff_B_2yOO5nOM6_0;
	wire w_dff_B_sOUdE9qb5_0;
	wire w_dff_B_xcePaCNo1_0;
	wire w_dff_B_63vNJJiu5_0;
	wire w_dff_B_2PqNYrIe4_0;
	wire w_dff_B_8b1ag7og5_0;
	wire w_dff_B_gdeiR5LT7_0;
	wire w_dff_B_Da09Io531_0;
	wire w_dff_B_dVmv9vHg3_0;
	wire w_dff_B_eHQHT7xz2_0;
	wire w_dff_B_SWLTI55M8_0;
	wire w_dff_B_LYXJn9qz4_0;
	wire w_dff_B_KGVo2PeX0_0;
	wire w_dff_B_LAXjsAFB4_0;
	wire w_dff_B_rI9Nzwhg7_0;
	wire w_dff_B_ugvjlxaC5_0;
	wire w_dff_B_NANNXVAV9_0;
	wire w_dff_B_j73X8DON5_0;
	wire w_dff_B_nTtcdtcO5_0;
	wire w_dff_B_MXzxbtLz1_0;
	wire w_dff_B_3cPKHPvk6_0;
	wire w_dff_B_xD0LztTD2_0;
	wire w_dff_B_zkxrkWd16_0;
	wire w_dff_B_4dp5WdPe5_0;
	wire w_dff_B_kZo5hkEK7_0;
	wire w_dff_B_hKeteD9J5_0;
	wire w_dff_B_Qhoj792v0_0;
	wire w_dff_B_jzhPpdlh0_0;
	wire w_dff_B_i1rua6Vc3_0;
	wire w_dff_B_9tkhkb5q0_0;
	wire w_dff_B_ZJ1rabc32_0;
	wire w_dff_B_s5I3v4ig9_0;
	wire w_dff_B_LkQJ95b28_0;
	wire w_dff_B_sQSXIYc20_0;
	wire w_dff_B_rkanMmVt0_0;
	wire w_dff_B_QGHErctr7_0;
	wire w_dff_B_PT7i1Ttz8_0;
	wire w_dff_B_dBxtBld69_0;
	wire w_dff_B_r4VKMphT6_0;
	wire w_dff_B_31MmSSZo3_0;
	wire w_dff_B_5uiwG3cc4_0;
	wire w_dff_B_YJlMuXGB9_0;
	wire w_dff_B_IZ6uK1A32_0;
	wire w_dff_B_878j9qzM5_0;
	wire w_dff_B_BIiO9j742_0;
	wire w_dff_B_Vs9rDLX22_0;
	wire w_dff_B_jK6Lh1E11_0;
	wire w_dff_B_xHhRv1Kb7_0;
	wire w_dff_B_Sf1jbtGk8_0;
	wire w_dff_B_UhV715RX2_0;
	wire w_dff_B_5YX6nJMq1_0;
	wire w_dff_B_5OX6T6bd1_0;
	wire w_dff_B_d5wbN7sk9_0;
	wire w_dff_B_q7YBMCvj4_0;
	wire w_dff_B_lLGCBk5P2_0;
	wire w_dff_B_yHIi2Z015_0;
	wire w_dff_B_BbYLq30u9_0;
	wire w_dff_B_ySBxrBfl7_0;
	wire w_dff_B_9gUZrYLs3_0;
	wire w_dff_B_mHreAn3l5_0;
	wire w_dff_B_9LvwDiqm0_0;
	wire w_dff_B_pb9bVdYe1_0;
	wire w_dff_B_LzJaCswK7_0;
	wire w_dff_B_GVilGTTs0_0;
	wire w_dff_B_qTM2WJ6g7_0;
	wire w_dff_B_18PBxVR25_0;
	wire w_dff_B_HbKJ7URU3_0;
	wire w_dff_B_IEfb7JRR2_0;
	wire w_dff_B_h6f9s4XF0_0;
	wire w_dff_B_QYHw80FP7_0;
	wire w_dff_B_8Mtd3Naa9_0;
	wire w_dff_B_JFTcRt9D8_0;
	wire w_dff_B_wscGVvbY9_0;
	wire w_dff_B_mGCbnmdl5_0;
	wire w_dff_B_sQV7d8l79_0;
	wire w_dff_B_apYOr9S20_0;
	wire w_dff_B_qnnpzRAH0_0;
	wire w_dff_B_U0pY4BZE9_0;
	wire w_dff_B_BHea5s6y5_0;
	wire w_dff_B_tsVuorQg7_0;
	wire w_dff_B_3K9S219l0_0;
	wire w_dff_B_toQCYd3N5_0;
	wire w_dff_B_tHZmABeR8_0;
	wire w_dff_B_YGTEzjhz4_0;
	wire w_dff_B_CLYSVPik4_0;
	wire w_dff_B_DlDxpIud7_0;
	wire w_dff_B_wYSkosGg7_0;
	wire w_dff_B_jirmYym30_0;
	wire w_dff_B_w7WuqIQE6_0;
	wire w_dff_B_ZI38D2bb7_0;
	wire w_dff_B_MTN3bQAP2_0;
	wire w_dff_B_W9tLR0IX1_0;
	wire w_dff_B_iTYTaTfQ0_0;
	wire w_dff_B_kvU20JZV5_0;
	wire w_dff_B_E60WvHlZ6_0;
	wire w_dff_B_KlI0Ouxa1_0;
	wire w_dff_B_thqkTFDY1_0;
	wire w_dff_B_EGAh7bB19_0;
	wire w_dff_B_blrktEUo2_0;
	wire w_dff_B_DYUpT7FU2_0;
	wire w_dff_B_pJOCtfPc7_0;
	wire w_dff_B_kZscPfF05_0;
	wire w_dff_B_QcZZTuIQ3_0;
	wire w_dff_B_4Ib2ppjx9_0;
	wire w_dff_B_V3gwhS3V5_0;
	wire w_dff_B_IYFP5TKO1_0;
	wire w_dff_B_X7wuqdgo1_0;
	wire w_dff_B_VnuZ65KF6_0;
	wire w_dff_B_UdcxoF2j6_0;
	wire w_dff_B_fAYQjJsa9_0;
	wire w_dff_B_CA2U5DbZ0_0;
	wire w_dff_B_aEgfGQY88_0;
	wire w_dff_B_8cCJzAnO8_0;
	wire w_dff_B_n5UIEOHW0_0;
	wire w_dff_B_yA4ojZ635_0;
	wire w_dff_B_fo0qJLoY3_0;
	wire w_dff_B_BQtJWMuP1_0;
	wire w_dff_B_wdKNfiWz1_0;
	wire w_dff_B_mmNYz6hq6_0;
	wire w_dff_B_B7YPRWT83_0;
	wire w_dff_B_HQlYCfa04_0;
	wire w_dff_B_ZjO0DUm18_0;
	wire w_dff_B_xGL6q3Bd5_0;
	wire w_dff_B_GFMVAOmn4_0;
	wire w_dff_B_WN0PGnhN3_0;
	wire w_dff_B_Fe2F91ED4_0;
	wire w_dff_B_rOptkkxL5_0;
	wire w_dff_B_Aom7jxAB4_0;
	wire w_dff_B_FAEDgE524_0;
	wire w_dff_B_VyYYL8Qt5_0;
	wire w_dff_B_YlYKYX4Q4_0;
	wire w_dff_B_gSPGKa2r4_0;
	wire w_dff_B_p6f5tlaT1_0;
	wire w_dff_B_vC3vzaYd9_0;
	wire w_dff_B_X1RoAtF93_0;
	wire w_dff_B_vhYTa54k4_0;
	wire w_dff_B_Ak161OG79_0;
	wire w_dff_B_DrnpvY3C8_0;
	wire w_dff_B_QrDIbC9f0_0;
	wire w_dff_B_3Bo961OP5_0;
	wire w_dff_B_IshJWfsA0_0;
	wire w_dff_B_E3GkM9bh2_0;
	wire w_dff_B_AbrcW48E5_0;
	wire w_dff_B_BiVauN6W1_0;
	wire w_dff_B_Y8Oh2AcU8_0;
	wire w_dff_B_TFZwZyeR2_0;
	wire w_dff_B_ZiNsTG490_0;
	wire w_dff_B_bz2HqiGf4_0;
	wire w_dff_B_1XjZcdtT3_0;
	wire w_dff_B_VmNzdaB18_0;
	wire w_dff_B_O8iW6WIQ4_0;
	wire w_dff_B_dnKQIDC61_0;
	wire w_dff_B_N5uL4RCF3_0;
	wire w_dff_B_gccVeE6L6_0;
	wire w_dff_B_c6euSobx0_0;
	wire w_dff_B_bZIcHaS78_0;
	wire w_dff_B_vHG4tcom6_0;
	wire w_dff_B_jmbnj2jO3_0;
	wire w_dff_B_6hZiz89g1_0;
	wire w_dff_B_hemcgMxm7_0;
	wire w_dff_B_A09Z9Qnf5_0;
	wire w_dff_B_POhBay9D2_0;
	wire w_dff_B_Ixb1pRGX6_0;
	wire w_dff_B_wdvdLn5n6_0;
	wire w_dff_B_TDogG1D40_0;
	wire w_dff_B_1owVF1lH7_0;
	wire w_dff_B_ha0SSQzY4_0;
	wire w_dff_B_2tyf0Uhe8_0;
	wire w_dff_B_yzEFVarW7_0;
	wire w_dff_B_hNYMxaaS9_0;
	wire w_dff_B_dFPTtBWq1_0;
	wire w_dff_B_cxlppIV79_0;
	wire w_dff_B_YVnsYMzi1_0;
	wire w_dff_B_HRdAuiEo4_0;
	wire w_dff_B_dVvbJW963_0;
	wire w_dff_B_FCutw8t22_0;
	wire w_dff_B_QClhmHSt5_0;
	wire w_dff_B_zRyHnnjd2_0;
	wire w_dff_B_kMl9yicX5_0;
	wire w_dff_B_VyIGJ9183_0;
	wire w_dff_B_3OfqcGYA6_0;
	wire w_dff_B_SxCzBEj88_0;
	wire w_dff_B_pbwwiBwO7_0;
	wire w_dff_B_agrR3ZMU5_0;
	wire w_dff_B_lw8QH2W58_0;
	wire w_dff_B_Mnw9cP8y6_0;
	wire w_dff_B_Cnw9lZYv5_0;
	wire w_dff_B_ptAe97e99_0;
	wire w_dff_B_A0K3CV4S3_0;
	wire w_dff_B_mILDGCpi8_0;
	wire w_dff_B_3SwRcVo26_0;
	wire w_dff_B_3ImerPUB9_0;
	wire w_dff_B_iu3g6XT02_0;
	wire w_dff_B_tvgBNtyF3_0;
	wire w_dff_B_DrFDeCqs3_0;
	wire w_dff_B_Z7mhA6AK0_0;
	wire w_dff_B_a4r6e87p8_0;
	wire w_dff_B_DC1xpvVx2_0;
	wire w_dff_B_JqBnzML99_0;
	wire w_dff_B_N6Dlo1VF8_0;
	wire w_dff_B_ZNuhTeA95_0;
	wire w_dff_B_OcH0zM7x5_0;
	wire w_dff_B_56CMJVCQ0_0;
	wire w_dff_B_WsCZY6uQ7_0;
	wire w_dff_B_rZgtu4FG9_0;
	wire w_dff_B_HpNBxB2c7_0;
	wire w_dff_B_gEWsEq7B9_0;
	wire w_dff_B_fUB77CFx7_0;
	wire w_dff_B_xlEFsqaD2_0;
	wire w_dff_B_3TpX3y4U1_0;
	wire w_dff_B_Mh8Lk0sf7_0;
	wire w_dff_B_nINtHQCR5_0;
	wire w_dff_B_8RSEU8P33_0;
	wire w_dff_B_lmmmKN3Y3_0;
	wire w_dff_B_8rswPLN26_0;
	wire w_dff_B_C0bAdgVI9_0;
	wire w_dff_B_rVKRJUWc9_0;
	wire w_dff_B_YRYNKleJ7_0;
	wire w_dff_B_fOXKvkXw7_0;
	wire w_dff_B_sUKwU3dg7_0;
	wire w_dff_B_HePElIVO0_0;
	wire w_dff_B_PFUUA1jQ0_0;
	wire w_dff_B_NMYaTAso6_0;
	wire w_dff_B_n4a4ziBb1_0;
	wire w_dff_B_IwOBWZwc1_0;
	wire w_dff_B_lCjMimkk7_0;
	wire w_dff_B_6ns0qHdv5_0;
	wire w_dff_B_D1bVyfCg7_0;
	wire w_dff_B_2dn2Sa3d9_0;
	wire w_dff_B_P68jduJO0_0;
	wire w_dff_B_6IjaQztm7_0;
	wire w_dff_B_K1LDRKNf6_0;
	wire w_dff_B_GFKdPcj02_0;
	wire w_dff_B_nKk7wij81_0;
	wire w_dff_B_MalIJpMY9_0;
	wire w_dff_B_FVkGPY8A4_0;
	wire w_dff_B_v3TbuZbB4_0;
	wire w_dff_B_ltmXst6H8_0;
	wire w_dff_B_OV2vOiv01_0;
	wire w_dff_B_x9YPzonl1_0;
	wire w_dff_B_ROVXGLfr9_0;
	wire w_dff_B_VNtrsrO71_0;
	wire w_dff_B_BXxgX8dt2_0;
	wire w_dff_B_u7Hu8Xtq8_0;
	wire w_dff_B_scYSoCvN2_0;
	wire w_dff_B_Rx2TCi7i0_0;
	wire w_dff_B_YWeOlb322_0;
	wire w_dff_B_m1nicARd3_0;
	wire w_dff_B_K3vHac6Q0_0;
	wire w_dff_B_bpZWisHi2_0;
	wire w_dff_B_2WAT7UkG4_0;
	wire w_dff_B_AtxdfFTw1_0;
	wire w_dff_B_WJdnsCAZ5_0;
	wire w_dff_B_pbHjgkNb1_0;
	wire w_dff_B_jzXi2paf6_0;
	wire w_dff_B_iEMhaJPs0_0;
	wire w_dff_B_xri6LWbP8_0;
	wire w_dff_B_Zi36Nuu53_0;
	wire w_dff_B_kP1VHHiD0_0;
	wire w_dff_B_r4NWKp934_0;
	wire w_dff_B_cfr2EdJo8_0;
	wire w_dff_B_WXj5shUv8_0;
	wire w_dff_B_fHL9ewFY8_0;
	wire w_dff_B_pC36Z5Il9_0;
	wire w_dff_B_bMIFxpYM3_0;
	wire w_dff_B_rKsRR8B18_0;
	wire w_dff_B_vnNcVzFb2_0;
	wire w_dff_B_ypXc36Wq4_0;
	wire w_dff_B_LROI9fzx7_0;
	wire w_dff_B_0LUjabfV5_0;
	wire w_dff_B_dXjo6nTt4_0;
	wire w_dff_B_Jp0UzgZy1_0;
	wire w_dff_B_NPhRZJrd5_0;
	wire w_dff_B_1aR2wi9I6_0;
	wire w_dff_B_P9ww9zfi6_0;
	wire w_dff_B_iwGZ0xgm9_0;
	wire w_dff_B_WamPNYCx7_0;
	wire w_dff_B_0Dw2PQsd0_0;
	wire w_dff_B_uf1tXRsq0_0;
	wire w_dff_B_pwH8bMZx2_0;
	wire w_dff_B_p9vSNjcF4_0;
	wire w_dff_B_gMihCNna4_0;
	wire w_dff_B_AnQv7iFL8_0;
	wire w_dff_B_6RfPHC5O5_0;
	wire w_dff_B_CNbq6GG21_0;
	wire w_dff_B_cdO0cDLa8_0;
	wire w_dff_B_N8p7dnMX3_0;
	wire w_dff_B_wml7S8l84_0;
	wire w_dff_B_M3Xd1PhB9_0;
	wire w_dff_B_Gqd7YsOb9_0;
	wire w_dff_B_HE8KoRyj2_0;
	wire w_dff_B_e9oF98zB1_0;
	wire w_dff_B_4BEID9NH3_0;
	wire w_dff_B_Xcol17ju2_0;
	wire w_dff_B_9yfiXWsL3_0;
	wire w_dff_B_dtPwKSWL7_0;
	wire w_dff_B_26hbwKBH1_0;
	wire w_dff_B_2elusBl54_0;
	wire w_dff_B_hIGgbbcT3_0;
	wire w_dff_B_RbHYZcMO1_0;
	wire w_dff_B_ugTyCguP0_0;
	wire w_dff_B_Of2N23Ai3_0;
	wire w_dff_B_bs1bV4Vw5_0;
	wire w_dff_B_elqrmwr35_0;
	wire w_dff_B_0Yegmpe35_0;
	wire w_dff_B_HJwMHHa77_0;
	wire w_dff_B_XYONRpMX3_0;
	wire w_dff_B_5nRM0Uqo0_0;
	wire w_dff_B_csfMFrXb0_0;
	wire w_dff_B_gwaIQQGJ1_0;
	wire w_dff_B_IoPXxkKg5_0;
	wire w_dff_B_Y6tCexmv9_0;
	wire w_dff_B_TbGpQ9YR5_0;
	wire w_dff_B_V8nrYw8x2_0;
	wire w_dff_B_4AuacWxR4_0;
	wire w_dff_B_z6eD9FLQ9_0;
	wire w_dff_B_YtT6L74T6_0;
	wire w_dff_B_rQwbrXEg3_0;
	wire w_dff_B_MImpxCfY7_0;
	wire w_dff_B_RhWXRdSz7_0;
	wire w_dff_B_e3grjneL8_0;
	wire w_dff_B_z6SUyQQp6_0;
	wire w_dff_B_wvitVInD3_0;
	wire w_dff_B_EJHIp3Av6_0;
	wire w_dff_B_fJIXlK8j6_0;
	wire w_dff_B_Ws8gdIGU2_0;
	wire w_dff_B_rOlXoMoq9_0;
	wire w_dff_B_rZsyBN5D7_0;
	wire w_dff_B_zadZWYrj3_0;
	wire w_dff_B_dcTCKUgQ6_0;
	wire w_dff_B_Lw6x3nZ96_0;
	wire w_dff_B_PcOoyN266_0;
	wire w_dff_B_C55CvjRy9_0;
	wire w_dff_B_roifZn3K3_0;
	wire w_dff_B_pwWdYu5t7_0;
	wire w_dff_B_5ERMbAsv8_0;
	wire w_dff_B_9IDcgHzL3_0;
	wire w_dff_B_W05GYXOh1_0;
	wire w_dff_B_HeNdTa4F7_0;
	wire w_dff_B_Uz6RhHJw9_0;
	wire w_dff_B_gIlfMgXj1_0;
	wire w_dff_B_xT417Rx08_0;
	wire w_dff_B_OCjNPtMl5_0;
	wire w_dff_B_pagZ7sfW8_0;
	wire w_dff_B_fjVtRjPI3_0;
	wire w_dff_B_zS96C8NC1_0;
	wire w_dff_B_clO5nt7m5_0;
	wire w_dff_B_zUsR3Qhs2_0;
	wire w_dff_B_RbhAgwFf4_0;
	wire w_dff_B_gNa9njv67_0;
	wire w_dff_B_8M7dDNxy3_0;
	wire w_dff_B_q3ro8XNg6_0;
	wire w_dff_B_rkbdtrsH9_0;
	wire w_dff_B_r1GeerKW4_0;
	wire w_dff_B_HwS05xRY1_0;
	wire w_dff_B_npdJYG3I4_0;
	wire w_dff_B_koDB1nkq4_0;
	wire w_dff_B_Q6VX4Jaw0_0;
	wire w_dff_B_Qv1b7M2u7_0;
	wire w_dff_B_VWUtoWC62_0;
	wire w_dff_B_8WOLjRNy1_0;
	wire w_dff_B_0zJCpDAt8_0;
	wire w_dff_B_T6wLnEUA3_0;
	wire w_dff_B_e5rNi6qV1_0;
	wire w_dff_B_Zsje3hqI7_0;
	wire w_dff_B_88gHF54N1_0;
	wire w_dff_B_9lBvPZZl7_0;
	wire w_dff_B_QmEDQSCh9_0;
	wire w_dff_B_Fg25dwkf4_0;
	wire w_dff_B_49ZjzouG7_0;
	wire w_dff_B_4M59PWGc6_0;
	wire w_dff_B_wSdLjt7N9_0;
	wire w_dff_B_j11bFsza9_0;
	wire w_dff_B_OhATlEu27_0;
	wire w_dff_B_vRIIBHzo3_0;
	wire w_dff_B_X3atVQTg5_0;
	wire w_dff_B_JrwEpjyr2_0;
	wire w_dff_B_Y98Q8kZG6_0;
	wire w_dff_B_p54lXqII9_0;
	wire w_dff_B_NO92IF1B7_0;
	wire w_dff_B_jK6mh18C6_0;
	wire w_dff_B_96gAZREG5_0;
	wire w_dff_B_bwacqj0h4_0;
	wire w_dff_B_qOsBJCSs0_0;
	wire w_dff_B_ASwJeVNh8_0;
	wire w_dff_B_tu9n90Yi2_0;
	wire w_dff_B_cZXH2y5q2_0;
	wire w_dff_B_5fv9iXVj7_0;
	wire w_dff_B_HwpyzPsg3_0;
	wire w_dff_B_DWZvWsa45_0;
	wire w_dff_B_aIMOrtzc2_0;
	wire w_dff_B_qclTWQc92_0;
	wire w_dff_B_l9LFpjIh4_0;
	wire w_dff_B_mpEr5KH37_0;
	wire w_dff_B_52FqaxSt7_0;
	wire w_dff_B_hvLK5edJ2_0;
	wire w_dff_B_xdPZG6vH2_0;
	wire w_dff_B_ZtE1BT2l8_0;
	wire w_dff_B_fT6YRSrD8_0;
	wire w_dff_B_wcjQj3bN8_0;
	wire w_dff_B_bSi6h9OL1_0;
	wire w_dff_B_z2nodQ5C6_0;
	wire w_dff_B_n5fYwwXW8_0;
	wire w_dff_B_1ZNI3kEJ1_0;
	wire w_dff_B_LJZC9NRv6_0;
	wire w_dff_B_qjOYAvwg1_0;
	wire w_dff_B_U7aOzUv02_0;
	wire w_dff_B_X6D9I1ru0_0;
	wire w_dff_B_TnML09fW1_0;
	wire w_dff_B_WJrzA8LD4_0;
	wire w_dff_B_nAiRgwlH5_0;
	wire w_dff_B_i4A5QtzN0_0;
	wire w_dff_B_dXZMItQ46_0;
	wire w_dff_B_K8ukcugw7_0;
	wire w_dff_B_h61f6hzY5_0;
	wire w_dff_B_sVa8StLI5_0;
	wire w_dff_B_vCxsbMFU3_0;
	wire w_dff_B_9nQbLlzI0_0;
	wire w_dff_B_n1EMLMJy0_0;
	wire w_dff_B_EUPZZoSL6_0;
	wire w_dff_B_SSH81M866_0;
	wire w_dff_B_mM8auC6O1_0;
	wire w_dff_B_x3oRt3C52_0;
	wire w_dff_B_KrPqwPbq3_0;
	wire w_dff_B_DGGLKCV08_0;
	wire w_dff_B_Sl5uAGPc7_0;
	wire w_dff_B_5CJTdA2k2_0;
	wire w_dff_B_ku9hUzde0_0;
	wire w_dff_B_YBNOgsWi6_0;
	wire w_dff_B_4OTtZhrV7_0;
	wire w_dff_B_xRFEj3YO8_0;
	wire w_dff_B_tgwVYjIg3_0;
	wire w_dff_B_7fpLCNfK4_0;
	wire w_dff_B_F2e0qTWi8_0;
	wire w_dff_B_MxSY16zF0_0;
	wire w_dff_B_IrsYUVUH1_0;
	wire w_dff_B_MsxkzGhm3_0;
	wire w_dff_B_JFxKYQfw4_0;
	wire w_dff_B_SofAR1CR7_0;
	wire w_dff_B_z3DGAngw5_0;
	wire w_dff_B_hPdt6xMi3_0;
	wire w_dff_B_mFrJLiJ80_0;
	wire w_dff_B_bTwy420H5_0;
	wire w_dff_B_cLuCe9RC7_0;
	wire w_dff_B_jtPbMuU01_0;
	wire w_dff_B_k05MxG376_0;
	wire w_dff_B_BPzy3ys37_0;
	wire w_dff_B_VqP6rJBB0_0;
	wire w_dff_B_fOVkZ61s4_0;
	wire w_dff_B_DVNaRLwH1_0;
	wire w_dff_B_jmmV1UR48_0;
	wire w_dff_B_Kc2Vev8J5_0;
	wire w_dff_B_StlBTWAv5_0;
	wire w_dff_B_DTWPbApp7_0;
	wire w_dff_B_ImRRhKX16_0;
	wire w_dff_B_T7cuqgKe6_0;
	wire w_dff_B_26iXzTi24_0;
	wire w_dff_B_P5raa7iH5_0;
	wire w_dff_B_534qgITM8_0;
	wire w_dff_B_pjy9kEid4_0;
	wire w_dff_B_IrLGOxd82_0;
	wire w_dff_B_LfZuWKDf0_0;
	wire w_dff_B_oMjt1qKM8_0;
	wire w_dff_B_vO8bFBFu7_0;
	wire w_dff_B_RqF7z6ix8_0;
	wire w_dff_B_wboFmJWv1_0;
	wire w_dff_B_9oT9nGjG2_0;
	wire w_dff_B_zSCdU7MV5_0;
	wire w_dff_B_EV00l0fe4_0;
	wire w_dff_B_EcNQHBKi3_0;
	wire w_dff_B_ZRCvYCot5_0;
	wire w_dff_B_ptdetvH26_0;
	wire w_dff_B_kZfIIG5p1_0;
	wire w_dff_B_9E9LPpF47_0;
	wire w_dff_B_cHRf4jFS6_0;
	wire w_dff_B_GpbFh6gO8_0;
	wire w_dff_B_XhbPu0R95_0;
	wire w_dff_B_RZJPVBIw7_0;
	wire w_dff_B_e8Q3EY8E5_0;
	wire w_dff_B_wf6N3ee44_0;
	wire w_dff_B_2dPm7vnJ7_0;
	wire w_dff_B_4J1Mwn6u0_0;
	wire w_dff_B_Ih6mbkCq0_0;
	wire w_dff_B_tnW2TgI04_0;
	wire w_dff_B_dZv1TT1s8_0;
	wire w_dff_B_rNgmYX2U0_0;
	wire w_dff_B_ov8QcAIA5_0;
	wire w_dff_B_ONygDv806_0;
	wire w_dff_B_14ddiKh63_0;
	wire w_dff_B_Vqh54OtS2_0;
	wire w_dff_B_erkFpigz8_0;
	wire w_dff_B_qqggysAj0_0;
	wire w_dff_B_hsrFqxlp6_0;
	wire w_dff_B_DfPvFU655_0;
	wire w_dff_B_yB2s3Z0O7_0;
	wire w_dff_B_VEuNX9yI7_0;
	wire w_dff_B_8FKK6kC72_0;
	wire w_dff_B_ON72gYPy2_0;
	wire w_dff_B_uFgbbB2u8_0;
	wire w_dff_B_pj7MqDkE2_0;
	wire w_dff_B_FnWyRtqy7_0;
	wire w_dff_B_iLs3lp5Y6_0;
	wire w_dff_B_Q8vJVLDZ4_0;
	wire w_dff_B_aN0kJfLk4_0;
	wire w_dff_B_Cjr67EwA1_0;
	wire w_dff_B_RNMzg2Ln6_0;
	wire w_dff_B_PGCdp9MW6_0;
	wire w_dff_B_v6bMOoiR8_0;
	wire w_dff_B_a7LsIWB48_0;
	wire w_dff_B_rtATlEVn0_0;
	wire w_dff_B_kjdSeWsF1_0;
	wire w_dff_B_LOvX9Jjn0_0;
	wire w_dff_B_T27tXn7v0_0;
	wire w_dff_B_SvjAMgLx0_0;
	wire w_dff_B_ls4nVUQ24_0;
	wire w_dff_B_I7yf34Bu8_0;
	wire w_dff_B_EZvSDj9R9_0;
	wire w_dff_B_rBYNYFbH4_0;
	wire w_dff_B_RjY3VDr80_0;
	wire w_dff_B_44rcrMNH1_0;
	wire w_dff_B_dU7m9MNj5_0;
	wire w_dff_B_UmUYOyza3_0;
	wire w_dff_B_VKB6AZcp7_0;
	wire w_dff_B_Cx3jRaYD6_0;
	wire w_dff_B_1DdhqPrz2_0;
	wire w_dff_B_M6UwPZ8z2_0;
	wire w_dff_B_mOnru5Gv3_0;
	wire w_dff_B_CWkhzmp43_0;
	wire w_dff_B_Sdq46Lib7_0;
	wire w_dff_B_FGDPvwzl4_0;
	wire w_dff_B_9fRtXgjP7_0;
	wire w_dff_B_swH8lO7r2_0;
	wire w_dff_B_FbfisYWQ7_0;
	wire w_dff_B_VPGX3hye7_0;
	wire w_dff_B_3dQSkHhr5_0;
	wire w_dff_B_4749LPl88_0;
	wire w_dff_B_Kr3St3gd4_0;
	wire w_dff_B_HaJtJ9W44_0;
	wire w_dff_B_6KybQLdZ8_0;
	wire w_dff_B_1Nb0u8t70_0;
	wire w_dff_B_woAwXAuG2_0;
	wire w_dff_B_XIdjPbaG5_0;
	wire w_dff_B_KTNTSNLj0_0;
	wire w_dff_B_Y7OVtIdX1_0;
	wire w_dff_B_Kz2tAwq64_0;
	wire w_dff_B_84m8ypX36_0;
	wire w_dff_B_tWLcj1rx9_0;
	wire w_dff_B_rGPCty7D2_0;
	wire w_dff_B_D7fCJeVx6_0;
	wire w_dff_B_UwCUdrn85_0;
	wire w_dff_B_Bs5fgbR58_0;
	wire w_dff_B_6yx3Ua6u2_0;
	wire w_dff_B_Wu6WLvLu6_0;
	wire w_dff_B_EiWb5KYS5_0;
	wire w_dff_B_HcIa7fiQ1_0;
	wire w_dff_B_VjETb8KY5_0;
	wire w_dff_B_HsADwHgF2_0;
	wire w_dff_B_TM57K66V9_0;
	wire w_dff_B_vD6JUPlz0_0;
	wire w_dff_B_kAT3upPx2_0;
	wire w_dff_B_krlCTgMQ1_0;
	wire w_dff_B_FerMHviC0_0;
	wire w_dff_B_4ve86PSQ0_0;
	wire w_dff_B_aMV6Svoj8_0;
	wire w_dff_B_ejDlgELE4_0;
	wire w_dff_B_GN0qANP52_0;
	wire w_dff_B_c2Jq4dcx7_0;
	wire w_dff_B_1BWEqvbk0_0;
	wire w_dff_B_dWECNPgy9_0;
	wire w_dff_B_rm5EmWSX5_0;
	wire w_dff_B_x1BF1BUU3_0;
	wire w_dff_B_4D0e6DQI6_0;
	wire w_dff_B_PUUCstNx9_0;
	wire w_dff_B_XA1RQxyR7_0;
	wire w_dff_B_nAbfrSV09_0;
	wire w_dff_B_Ab3IT7Dh2_0;
	wire w_dff_B_o7WwTovS6_0;
	wire w_dff_B_nYsULZsA3_0;
	wire w_dff_B_I3nbp6qU3_0;
	wire w_dff_B_9biXOlce0_0;
	wire w_dff_B_jIivYryf8_0;
	wire w_dff_B_mwrykKhY9_0;
	wire w_dff_B_OgruAIXJ9_0;
	wire w_dff_B_YyVIEu8A4_0;
	wire w_dff_B_J4Tc4Nfx2_0;
	wire w_dff_B_puVG3F539_0;
	wire w_dff_B_0OjSc4mg1_0;
	wire w_dff_B_MUt2RQG45_0;
	wire w_dff_B_1JLdUdCP3_0;
	wire w_dff_B_o2WsywEg8_0;
	wire w_dff_B_qDb9SBpR7_0;
	wire w_dff_B_nRAWg75X2_0;
	wire w_dff_B_muX7q6CO0_0;
	wire w_dff_B_JhrC8uVe4_0;
	wire w_dff_B_QUTIphUX9_0;
	wire w_dff_B_JrjXALgH0_0;
	wire w_dff_B_5Ov3MkWU4_0;
	wire w_dff_B_WOL3ufiO1_0;
	wire w_dff_B_tWbNMCYe9_0;
	wire w_dff_B_RFIbUvxx2_0;
	wire w_dff_B_3fEKCzTR8_0;
	wire w_dff_B_pnxrMXfL6_0;
	wire w_dff_B_uUkfOFQn1_0;
	wire w_dff_B_QtSE2alq8_0;
	wire w_dff_B_a60LwpbU0_0;
	wire w_dff_B_1xKJMbsb7_0;
	wire w_dff_B_zyFmT5e05_0;
	wire w_dff_B_p5DSkSea4_0;
	wire w_dff_B_OMwW1Zbs2_0;
	wire w_dff_B_7ean7UXY0_0;
	wire w_dff_B_oitKwxnb4_0;
	wire w_dff_B_PeXnXtj88_0;
	wire w_dff_B_t2TBwC2m4_0;
	wire w_dff_B_xpfmd1fS5_0;
	wire w_dff_B_yiz34MsO2_0;
	wire w_dff_B_aZrBtuQV7_0;
	wire w_dff_B_hrLHjEyU9_0;
	wire w_dff_B_s3kqD9F70_0;
	wire w_dff_B_MRPGm56t9_0;
	wire w_dff_B_idYSafC78_0;
	wire w_dff_B_mzo147uB9_0;
	wire w_dff_B_wW80m5xJ7_0;
	wire w_dff_B_iX1elz686_0;
	wire w_dff_B_XWi7Zoti3_0;
	wire w_dff_B_9EyMk9Bx3_0;
	wire w_dff_B_jg09GqFo7_0;
	wire w_dff_B_cXvUOrSZ5_0;
	wire w_dff_B_IiXRSKqj0_0;
	wire w_dff_B_QaPpatWl3_0;
	wire w_dff_B_gmU7MplD8_0;
	wire w_dff_B_FKgzxNck2_0;
	wire w_dff_B_iuRBEMsL8_0;
	wire w_dff_B_zhWBGiw30_0;
	wire w_dff_B_c16mnQyi5_0;
	wire w_dff_B_kZoiANpD2_0;
	wire w_dff_B_Ue9aPG913_0;
	wire w_dff_B_GxxhsJjw6_0;
	wire w_dff_B_fviA1pj29_0;
	wire w_dff_B_0m1XsGUV5_0;
	wire w_dff_B_mFuzQE5A0_0;
	wire w_dff_B_yBF9yxPn5_0;
	wire w_dff_B_VOIcKW1j8_0;
	wire w_dff_B_SVgJJ2vo8_0;
	wire w_dff_B_OeJl0nhT7_0;
	wire w_dff_B_KBTawIzE0_0;
	wire w_dff_B_pb8aXKb90_0;
	wire w_dff_B_0fImpkSC8_0;
	wire w_dff_B_Sq1RSOax7_0;
	wire w_dff_B_iYF7zXYh2_0;
	wire w_dff_B_fl8zZlLZ3_0;
	wire w_dff_B_cbmYB3cD6_0;
	wire w_dff_B_JGvRZpqj5_0;
	wire w_dff_B_hrlz2aiW6_0;
	wire w_dff_B_h9Vbz6W55_0;
	wire w_dff_B_dmNLg6ON4_0;
	wire w_dff_B_DuZZPuLK1_0;
	wire w_dff_B_Cr0eBaQe4_0;
	wire w_dff_B_4FSo0TXl9_0;
	wire w_dff_B_3Vl08xmX6_0;
	wire w_dff_B_RGnPaSJw9_0;
	wire w_dff_B_7zZFrWzC0_0;
	wire w_dff_B_i0WlbGm57_0;
	wire w_dff_B_AKFeOXCo2_0;
	wire w_dff_B_rCV0ZODX8_0;
	wire w_dff_B_Y5tZFD296_0;
	wire w_dff_B_dYkw7LMd5_0;
	wire w_dff_B_79TJ03jF6_0;
	wire w_dff_B_KoJVSAfr6_0;
	wire w_dff_B_ninceOZA1_0;
	wire w_dff_B_ZLiEY06c5_0;
	wire w_dff_B_a0Wtax9k9_0;
	wire w_dff_B_KDAiu1qz2_0;
	wire w_dff_B_KvTUSNaz7_0;
	wire w_dff_B_x63XX1Ly6_0;
	wire w_dff_B_wbr0oOuf3_0;
	wire w_dff_B_87DRgOHA1_0;
	wire w_dff_B_k8hJc1TX5_0;
	wire w_dff_B_epM7xax95_0;
	wire w_dff_B_IiYF23UO4_0;
	wire w_dff_B_w13Ku9pw9_0;
	wire w_dff_B_nH9UmjbH6_0;
	wire w_dff_B_K5JydMTT7_0;
	wire w_dff_B_QcRFm2ko6_0;
	wire w_dff_B_OZsDaZDK5_0;
	wire w_dff_B_krgSRuj05_0;
	wire w_dff_B_VUY6y9pD5_0;
	wire w_dff_B_ifKdVjtU2_0;
	wire w_dff_B_YsAFealH2_0;
	wire w_dff_B_erm8ltah9_0;
	wire w_dff_B_ynh2rDWK5_0;
	wire w_dff_B_teUIUmXN2_0;
	wire w_dff_B_36Nr5e4v0_0;
	wire w_dff_B_evYzW6yN9_0;
	wire w_dff_B_A2EaiSLS2_0;
	wire w_dff_B_3WES9sEE4_0;
	wire w_dff_B_i8VZmfPt2_0;
	wire w_dff_B_VAXZtPOg8_0;
	wire w_dff_B_Q0AGl5hU8_0;
	wire w_dff_B_dckM39du9_0;
	wire w_dff_B_IzjaZ1XN1_0;
	wire w_dff_B_rJRZKPlQ9_0;
	wire w_dff_B_ZJ7IgyKt1_0;
	wire w_dff_B_GLeXHGI72_0;
	wire w_dff_B_8orOh9oT4_0;
	wire w_dff_B_DCVvUxlg7_0;
	wire w_dff_B_zfvIZB2u3_0;
	wire w_dff_B_alLn5dug9_0;
	wire w_dff_B_fNKQ5FxJ5_0;
	wire w_dff_B_zIFcmTRN6_0;
	wire w_dff_B_dIAPTpEE3_0;
	wire w_dff_B_SvocjBtu9_0;
	wire w_dff_B_5XM7lrJ18_0;
	wire w_dff_B_AvvWnsEE4_0;
	wire w_dff_B_LDPSWqN55_0;
	wire w_dff_B_Ne51fv8f4_0;
	wire w_dff_B_tiZ4KHiW2_0;
	wire w_dff_B_I2jlKbNp8_0;
	wire w_dff_B_cNBkCEVi1_0;
	wire w_dff_B_NQ03wBgH1_0;
	wire w_dff_B_Hlu0yAFh2_0;
	wire w_dff_B_9fjo0r898_0;
	wire w_dff_B_UJWMk3Z27_0;
	wire w_dff_B_euGD2qB86_0;
	wire w_dff_B_fjNKgvcU9_0;
	wire w_dff_B_4Vqi2sXR0_0;
	wire w_dff_B_EyBF3q6K5_0;
	wire w_dff_B_0JLHOIUQ5_0;
	wire w_dff_B_PA6TGe5t5_0;
	wire w_dff_B_LnVF8d2f1_0;
	wire w_dff_B_aPbt9GGI7_0;
	wire w_dff_B_7vk1Ogy88_0;
	wire w_dff_B_ZrbQErD96_0;
	wire w_dff_B_QlkWJsah4_0;
	wire w_dff_B_BZuEnWnu4_0;
	wire w_dff_B_QYwB1byA3_0;
	wire w_dff_B_6csUr0Hr4_0;
	wire w_dff_B_RA6pGNX62_0;
	wire w_dff_B_hdIg99Ys2_0;
	wire w_dff_B_l42FmOb26_0;
	wire w_dff_B_nE6sKC2a9_0;
	wire w_dff_B_cXEgdtn60_0;
	wire w_dff_B_xrPnkjAD4_0;
	wire w_dff_B_NyMCjCYC9_0;
	wire w_dff_B_FQKpehzb2_0;
	wire w_dff_B_0lyI64ZE3_0;
	wire w_dff_B_DVswJc5Z6_0;
	wire w_dff_B_BSKY3utX3_0;
	wire w_dff_B_K9SkFrZw4_0;
	wire w_dff_B_MCHK6wHv1_0;
	wire w_dff_B_PQbkRS7H2_0;
	wire w_dff_B_52sZSUvo4_0;
	wire w_dff_B_679TxmNw3_0;
	wire w_dff_B_h2KF3RLB3_0;
	wire w_dff_B_ILY51LBP4_0;
	wire w_dff_B_cs6IY91D8_0;
	wire w_dff_B_qFtykAGp8_0;
	wire w_dff_B_knLqfLUQ0_0;
	wire w_dff_B_lvEXTfsp2_0;
	wire w_dff_B_G4Gr10HC0_0;
	wire w_dff_B_vQpZ6Imv8_0;
	wire w_dff_B_zlbjkOeu8_0;
	wire w_dff_B_hAxxrdp33_0;
	wire w_dff_B_Xe44QXIQ1_0;
	wire w_dff_B_JthLW1dC9_0;
	wire w_dff_B_AfVvE9ms4_0;
	wire w_dff_B_yQndL1I96_0;
	wire w_dff_B_ZQpNBVcN9_0;
	wire w_dff_B_yhlUcBIH5_0;
	wire w_dff_B_CPhFAnYN7_0;
	wire w_dff_B_lbTHRrQO6_0;
	wire w_dff_B_Mx8h8HwG9_0;
	wire w_dff_B_yZr8mdDz5_0;
	wire w_dff_B_zsTH0Awc5_0;
	wire w_dff_B_miPfl8T48_0;
	wire w_dff_B_WoAWFxgM3_0;
	wire w_dff_B_sXDzow1e0_0;
	wire w_dff_B_Yo2B737v3_0;
	wire w_dff_B_HLQWv4eU2_0;
	wire w_dff_B_o6xCwdXu5_0;
	wire w_dff_B_tc3u8w468_0;
	wire w_dff_B_14EdoGIE1_0;
	wire w_dff_B_ykoox14D0_0;
	wire w_dff_B_V7sInmd47_0;
	wire w_dff_B_jNfKLFXS1_0;
	wire w_dff_B_mWjTHgVh6_0;
	wire w_dff_B_f7Ele7RO9_0;
	wire w_dff_B_piWs9FDx6_0;
	wire w_dff_B_XoVzFCJj4_0;
	wire w_dff_B_fLGqLtS47_0;
	wire w_dff_B_Hqg8jK0B1_0;
	wire w_dff_B_vqnhZzCs2_0;
	wire w_dff_B_E8l6wy0I3_0;
	wire w_dff_B_dvqeaSij1_0;
	wire w_dff_B_wl7LBGnw1_0;
	wire w_dff_B_GYR9jce80_0;
	wire w_dff_B_zuqBaa1S9_0;
	wire w_dff_B_FJzbmHpf0_0;
	wire w_dff_B_FvAWsfAE8_0;
	wire w_dff_B_tVs9R9vG9_0;
	wire w_dff_B_svSuWFHX8_0;
	wire w_dff_B_DDPQKyId7_0;
	wire w_dff_B_wwokALGe8_0;
	wire w_dff_B_yrfvQdy76_0;
	wire w_dff_B_pDVPPZn74_0;
	wire w_dff_B_LCgeEXT91_0;
	wire w_dff_B_mTHEaqJk3_0;
	wire w_dff_B_5tLVq2XS7_0;
	wire w_dff_B_Bb3m5DC66_0;
	wire w_dff_B_PKeVa7sH0_0;
	wire w_dff_B_zmvkgoz16_0;
	wire w_dff_B_xLHrsSlh6_0;
	wire w_dff_B_ZXpFUhLT6_0;
	wire w_dff_B_Ao1UVAxz4_0;
	wire w_dff_B_u3YMuD0w7_0;
	wire w_dff_B_TJU8CB1K9_0;
	wire w_dff_B_PJvjguEn8_0;
	wire w_dff_B_xopPfgnR5_0;
	wire w_dff_B_3fx4ymWY5_0;
	wire w_dff_B_ZbCqZhea4_0;
	wire w_dff_B_I8HSUCXM1_0;
	wire w_dff_B_vuPeDlkB9_0;
	wire w_dff_B_QIQQwm6M6_0;
	wire w_dff_B_3UBzza6x6_0;
	wire w_dff_B_RorxNhg46_0;
	wire w_dff_B_rr3m3kMy9_0;
	wire w_dff_B_u6N0CKnZ2_0;
	wire w_dff_B_I200MfGu1_0;
	wire w_dff_B_UnW3HPIw5_0;
	wire w_dff_B_7x7R4RIK4_0;
	wire w_dff_B_zj3vQalB8_0;
	wire w_dff_B_CaCXwbVA0_0;
	wire w_dff_B_KjEFd3Tr2_0;
	wire w_dff_B_eoRU2Dig8_0;
	wire w_dff_B_XF4TZrF18_0;
	wire w_dff_B_kFIBnhRV3_0;
	wire w_dff_B_bsb7w8Ld0_0;
	wire w_dff_B_BHGtaNg47_0;
	wire w_dff_B_ENYkbVwg8_0;
	wire w_dff_B_yippQWKC3_0;
	wire w_dff_B_vnYCDvKi3_0;
	wire w_dff_B_WxKeVE7v8_0;
	wire w_dff_B_0UN5UyyP6_0;
	wire w_dff_B_6h4QR3wu1_0;
	wire w_dff_B_mzldZlCK9_0;
	wire w_dff_B_CjJInOFP4_0;
	wire w_dff_B_tg9dYumo2_0;
	wire w_dff_B_atYxgtNA9_0;
	wire w_dff_B_ZBWtA7WT3_0;
	wire w_dff_B_llTlEFUM4_0;
	wire w_dff_B_JFgWisLP9_0;
	wire w_dff_B_WnrB3uOv4_0;
	wire w_dff_B_xl5GkG4S3_0;
	wire w_dff_B_evmwPmZp5_0;
	wire w_dff_B_9v14hgE90_0;
	wire w_dff_B_Vws8LjOK8_0;
	wire w_dff_B_5rb1BXV10_0;
	wire w_dff_B_nKYOxuLI3_0;
	wire w_dff_B_mecQYNlA7_0;
	wire w_dff_B_RCFoAGTf5_0;
	wire w_dff_B_hDJREAJx5_0;
	wire w_dff_B_ogBL6tSm1_0;
	wire w_dff_B_3Lz9qtbN5_0;
	wire w_dff_B_rtfxgeGM8_0;
	wire w_dff_B_0AH7p5RH7_0;
	wire w_dff_B_4x8jDMf12_0;
	wire w_dff_B_hUNL9Unj1_0;
	wire w_dff_B_jeAaxdpn6_0;
	wire w_dff_B_74tiN2Vz8_0;
	wire w_dff_B_krFHa4VO1_0;
	wire w_dff_B_l5MegGRP7_0;
	wire w_dff_B_SvCz5SVf1_0;
	wire w_dff_B_Ns6paOb38_0;
	wire w_dff_B_Mz12lt6A9_0;
	wire w_dff_B_RMoNROTT9_0;
	wire w_dff_B_v0WrVMHE7_0;
	wire w_dff_B_xb3SG3cp0_0;
	wire w_dff_B_YHXAcmMC2_0;
	wire w_dff_B_fVLAJgwU3_0;
	wire w_dff_B_bB01Exob1_0;
	wire w_dff_B_lOHYKota2_0;
	wire w_dff_B_9ql3TWyJ3_0;
	wire w_dff_B_1kldjOYI8_0;
	wire w_dff_B_oIgOlh7c4_0;
	wire w_dff_B_HyOB6jnY9_0;
	wire w_dff_B_jZviLZL95_0;
	wire w_dff_B_8MIPVDkK5_0;
	wire w_dff_B_gzTQnsKE7_0;
	wire w_dff_B_7gbW1flP8_0;
	wire w_dff_B_NsrK7wS07_0;
	wire w_dff_B_7x5hpzsk3_0;
	wire w_dff_B_7W05GFDH2_0;
	wire w_dff_B_yNH3dqqb9_0;
	wire w_dff_B_Jf7TFLmy3_0;
	wire w_dff_B_KyJ1suCw5_0;
	wire w_dff_B_RxOwBrzg8_0;
	wire w_dff_B_2KaLYNB77_0;
	wire w_dff_B_zAQfmmks4_0;
	wire w_dff_B_Coi5c6uW9_0;
	wire w_dff_B_xZpFUUVQ1_0;
	wire w_dff_B_VqPChw8q9_0;
	wire w_dff_B_8cFO0wxB1_0;
	wire w_dff_B_M2vePlTa1_0;
	wire w_dff_B_kfcsDZEe9_0;
	wire w_dff_B_4cvrNabJ5_0;
	wire w_dff_B_PeUrXRar1_0;
	wire w_dff_B_KwlAvEJO9_0;
	wire w_dff_B_M5Km0IC42_0;
	wire w_dff_B_WbF1jP9J5_0;
	wire w_dff_B_a3KQkaOj6_0;
	wire w_dff_B_YrVuElf97_0;
	wire w_dff_B_ZKgBPr5l0_0;
	wire w_dff_B_8dWM9WLj4_0;
	wire w_dff_B_OyaThRrB8_0;
	wire w_dff_B_BYGhXWV19_0;
	wire w_dff_B_KMMLpX870_0;
	wire w_dff_B_xE22n2gA2_0;
	wire w_dff_B_eek1d2Wg1_0;
	wire w_dff_B_6LtcpZ0P2_0;
	wire w_dff_B_PlLqyFs54_0;
	wire w_dff_B_2wn8wvNT5_0;
	wire w_dff_B_NJNmvW7d4_0;
	wire w_dff_B_HQtN0HWE1_0;
	wire w_dff_B_rsVJgZa16_0;
	wire w_dff_B_EWG3f3tx2_0;
	wire w_dff_B_cScT3Bku6_0;
	wire w_dff_B_2b5Edwz26_0;
	wire w_dff_B_m3vZCVYd5_0;
	wire w_dff_B_1WhLU8m30_0;
	wire w_dff_B_6amr7AjJ7_0;
	wire w_dff_B_HDFdf9d89_0;
	wire w_dff_B_v7kZVRhL5_0;
	wire w_dff_B_OleMdkzj5_0;
	wire w_dff_B_91Mn7IRd9_0;
	wire w_dff_B_IaacLBCk8_0;
	wire w_dff_B_HMJx3LXH4_0;
	wire w_dff_B_cYxv0T411_0;
	wire w_dff_B_8VYO2KIZ4_0;
	wire w_dff_B_Fv0xdtCj1_0;
	wire w_dff_B_ei42O0my7_0;
	wire w_dff_B_smcaRgdt0_0;
	wire w_dff_B_OmXcePvN4_0;
	wire w_dff_B_JwZqahIm8_0;
	wire w_dff_B_5gDMRACq6_0;
	wire w_dff_B_pgIX1swX2_0;
	wire w_dff_B_logAA0ks9_0;
	wire w_dff_B_BVXBqqUR5_0;
	wire w_dff_B_slySt0GR3_0;
	wire w_dff_B_zBnkBPnf2_0;
	wire w_dff_B_Noal6Ocm4_0;
	wire w_dff_B_2GmTQCri3_0;
	wire w_dff_B_vNriQ0Vb5_0;
	wire w_dff_B_dAe9zNSK3_0;
	wire w_dff_B_OC7rTDjS7_0;
	wire w_dff_B_kCm3iSPC2_0;
	wire w_dff_B_YgouYNVU9_0;
	wire w_dff_B_oBZLviGg4_0;
	wire w_dff_B_vgkiyEAh6_0;
	wire w_dff_B_fhcfjD9y4_0;
	wire w_dff_B_XPUb2IrR6_0;
	wire w_dff_B_Yi1rEeFd2_0;
	wire w_dff_B_HxQvK6lw6_0;
	wire w_dff_B_rNhTu0Fi9_0;
	wire w_dff_B_OcI7n4Lp2_0;
	wire w_dff_B_RsujpwAI8_0;
	wire w_dff_B_NrE4IRjb7_0;
	wire w_dff_B_Xfw0J6eh3_0;
	wire w_dff_B_UdcaEZAD4_0;
	wire w_dff_B_7pOuXS1g4_0;
	wire w_dff_B_QE1Q7emD3_0;
	wire w_dff_B_eA957Lio5_0;
	wire w_dff_B_9QEuLWPn3_0;
	wire w_dff_B_XVbpx3LL7_0;
	wire w_dff_B_IV28YlRB1_0;
	wire w_dff_B_YWPOyVwS0_0;
	wire w_dff_B_eNgZMEAZ9_0;
	wire w_dff_B_OA6rj82y0_0;
	wire w_dff_B_mjzcpdz86_0;
	wire w_dff_B_YHOhW1QB9_0;
	wire w_dff_B_Pdbx63Z19_0;
	wire w_dff_B_RNaotcwI3_0;
	wire w_dff_B_57BS15644_0;
	wire w_dff_B_55ZTfQup5_0;
	wire w_dff_B_HCgo7Hcf4_0;
	wire w_dff_B_OMyKHvgZ2_0;
	wire w_dff_B_x9ZWGzaE2_0;
	wire w_dff_B_IIiexAjM3_0;
	wire w_dff_B_mB6wE1yn1_0;
	wire w_dff_B_fL2y0fpg7_0;
	wire w_dff_B_0keNPwNm7_0;
	wire w_dff_B_0YU51EUf1_0;
	wire w_dff_B_1fRvMtBU8_0;
	wire w_dff_B_eNM5LHYZ1_0;
	wire w_dff_B_mmumLB8T4_0;
	wire w_dff_B_24OWo8On2_0;
	wire w_dff_B_Xnkv6wpE2_0;
	wire w_dff_B_ClGaX7et6_0;
	wire w_dff_B_ZkimcW9H4_0;
	wire w_dff_B_wuLaYuXU0_0;
	wire w_dff_B_6oRMzsHG0_0;
	wire w_dff_B_hcqYwIxD0_0;
	wire w_dff_B_GLy3QedQ0_0;
	wire w_dff_B_g7nyyOxt6_0;
	wire w_dff_B_Hj2cCQXp4_0;
	wire w_dff_B_7qQeG4ym9_0;
	wire w_dff_B_zj3Ax0SY9_0;
	wire w_dff_B_JVfwb49E3_0;
	wire w_dff_B_v0Ap766Z6_0;
	wire w_dff_B_OVzwgguU2_0;
	wire w_dff_B_enkNNa8E7_0;
	wire w_dff_B_5tjnvZyx1_0;
	wire w_dff_B_ldNbWkD46_0;
	wire w_dff_B_razZ34i70_0;
	wire w_dff_B_iA3bsgiS9_0;
	wire w_dff_B_WQN2CA9w4_0;
	wire w_dff_B_eqPSxxTU2_0;
	wire w_dff_B_hf3r0Hiu1_0;
	wire w_dff_B_hiOftxfl0_0;
	wire w_dff_B_30Lb7JtM3_0;
	wire w_dff_B_iU7lI2O91_0;
	wire w_dff_B_0cwLrV9z8_0;
	wire w_dff_B_tQitZD2H6_0;
	wire w_dff_B_mbBXjP7c9_0;
	wire w_dff_B_ctXXeX4L3_0;
	wire w_dff_B_aiRcMePC2_0;
	wire w_dff_B_sNHO2xgZ7_0;
	wire w_dff_B_ginmtGZ63_0;
	wire w_dff_B_K9pCFAio9_0;
	wire w_dff_B_K67xS4pS4_0;
	wire w_dff_B_hVqyHXBV9_0;
	wire w_dff_B_6z6HtBD57_0;
	wire w_dff_B_AUHRhyGt5_0;
	wire w_dff_B_TkgeNQY00_0;
	wire w_dff_B_zpwJvQ515_0;
	wire w_dff_B_WDjhrQKW0_0;
	wire w_dff_B_V270VAkB9_0;
	wire w_dff_B_ycw05gBQ0_0;
	wire w_dff_B_lcnAP0z92_0;
	wire w_dff_B_DfF5ngS37_0;
	wire w_dff_B_NXHrwrVd0_0;
	wire w_dff_B_AGThUvVk7_0;
	wire w_dff_B_RNRT9YyD6_0;
	wire w_dff_B_aBoh4ovx6_0;
	wire w_dff_B_JindIYki7_0;
	wire w_dff_B_c0dpcB5P3_0;
	wire w_dff_B_s7MyU8fC4_0;
	wire w_dff_B_MoIgWBGR4_0;
	wire w_dff_B_ub22zWvN3_0;
	wire w_dff_B_lJOSsY171_0;
	wire w_dff_B_L6XEqsQD2_0;
	wire w_dff_B_I4C07N0v0_0;
	wire w_dff_B_wXsBjVto8_0;
	wire w_dff_B_9vfeCqXL4_0;
	wire w_dff_B_cjd6mApc6_0;
	wire w_dff_B_ZuhHacUi8_0;
	wire w_dff_B_jqPInde50_0;
	wire w_dff_B_ItioxTAY9_0;
	wire w_dff_B_0QPZ31Wc8_0;
	wire w_dff_B_lpUMr7ja7_0;
	wire w_dff_B_MTK2mGuD8_0;
	wire w_dff_B_t0AoUYbB4_0;
	wire w_dff_B_LKPy1WfB0_0;
	wire w_dff_B_h8DSVQj50_0;
	wire w_dff_B_ikxjbfcP3_0;
	wire w_dff_B_SXAKrERt1_0;
	wire w_dff_B_57EwLenK7_0;
	wire w_dff_B_0bl1NVbR4_0;
	wire w_dff_B_cJmYllNu8_0;
	wire w_dff_B_S0eHrJej0_0;
	wire w_dff_B_pjfiUR7r9_0;
	wire w_dff_B_Twpr0dGv4_0;
	wire w_dff_B_eW4XODF99_0;
	wire w_dff_B_Jo1gIF7K4_0;
	wire w_dff_B_VnSgSmds6_0;
	wire w_dff_B_z06JAgyL8_0;
	wire w_dff_B_f9r7QJFW6_0;
	wire w_dff_B_BfgMa1Bj8_0;
	wire w_dff_B_i5lceecz9_0;
	wire w_dff_B_78vPS1tb1_0;
	wire w_dff_B_YgGHVgip6_0;
	wire w_dff_B_QBbMYkpT0_0;
	wire w_dff_B_V4yv1Dm83_0;
	wire w_dff_B_CPKzqgqd9_0;
	wire w_dff_B_0oeP7dUY2_0;
	wire w_dff_B_pumxgpUT7_0;
	wire w_dff_B_RlP2hxfb9_0;
	wire w_dff_B_H5RqFnkF4_0;
	wire w_dff_B_Vyawy5hR4_0;
	wire w_dff_B_TTvxEKge3_0;
	wire w_dff_B_lgsZtvDU5_0;
	wire w_dff_B_dXyKjo3Z3_0;
	wire w_dff_B_xqNNXwyF1_0;
	wire w_dff_B_e1hQjS0U0_0;
	wire w_dff_B_LyveZ1Xv9_0;
	wire w_dff_B_oQyy2W5V3_0;
	wire w_dff_B_l8okepPR3_0;
	wire w_dff_B_NgmasIYY3_0;
	wire w_dff_B_ValgLkKF1_0;
	wire w_dff_B_9g6oaCFv5_0;
	wire w_dff_B_CORAAWD78_0;
	wire w_dff_B_5MdrKi917_0;
	wire w_dff_B_qdA9zPt24_0;
	wire w_dff_B_HaUILZLG0_0;
	wire w_dff_B_0PzgsZbI1_0;
	wire w_dff_B_mpeAJpV75_0;
	wire w_dff_B_zrk2oeIB9_0;
	wire w_dff_B_ZSdTDVQk8_0;
	wire w_dff_B_sGHXupt62_0;
	wire w_dff_B_wDbBQEJO2_0;
	wire w_dff_B_ZbwhacVQ4_0;
	wire w_dff_B_IT05QkwA1_0;
	wire w_dff_B_6lP44hqT6_0;
	wire w_dff_B_tNCiAupb8_0;
	wire w_dff_B_DdJ72lJM3_0;
	wire w_dff_B_xj5rbALU6_0;
	wire w_dff_B_IeLeMarR4_0;
	wire w_dff_B_bI9VxqpI7_0;
	wire w_dff_B_CXeqhXDz3_0;
	wire w_dff_B_3yANIJ0n1_0;
	wire w_dff_B_SgKEG25y2_0;
	wire w_dff_B_rtLKtDF75_0;
	wire w_dff_B_tsJ7SVNS7_0;
	wire w_dff_B_cR2iWGNm2_0;
	wire w_dff_B_qXsr8YMz5_0;
	wire w_dff_B_1xXRNM1N8_0;
	wire w_dff_B_8vJgU9Pd0_0;
	wire w_dff_B_neOEgyy66_0;
	wire w_dff_B_g7yG9TCX9_0;
	wire w_dff_B_ObmE9enM5_0;
	wire w_dff_B_xG7ijfTh9_0;
	wire w_dff_B_r29RsP4F6_0;
	wire w_dff_B_GC0tytrT3_0;
	wire w_dff_B_maDeWo187_0;
	wire w_dff_B_99vLvXpZ7_0;
	wire w_dff_B_aOkopAdL7_0;
	wire w_dff_B_iENNeByh6_0;
	wire w_dff_B_lDGt7iS93_0;
	wire w_dff_B_ANGAEBR29_0;
	wire w_dff_B_EROz8aSS0_0;
	wire w_dff_B_HVTuliIy6_0;
	wire w_dff_B_pbghLIdh4_0;
	wire w_dff_B_OqqO1U7D9_0;
	wire w_dff_B_JiyGNTAj4_0;
	wire w_dff_B_XUnZMClu4_0;
	wire w_dff_B_DlU8PPoj8_0;
	wire w_dff_B_VxUgdIIL1_0;
	wire w_dff_B_mYBB8z7y8_0;
	wire w_dff_B_HjJ4US4Q1_0;
	wire w_dff_B_r3VVL3Wb7_0;
	wire w_dff_B_voI9mhzg2_0;
	wire w_dff_B_FqLqem4x5_0;
	wire w_dff_B_lShsHD8R7_0;
	wire w_dff_B_bkKN7mRm3_0;
	wire w_dff_B_c3wEEVfN9_0;
	wire w_dff_B_BQqbw3445_0;
	wire w_dff_B_lwQ1oD6S9_0;
	wire w_dff_B_y9Q5au4T4_0;
	wire w_dff_B_DxK7zWo11_0;
	wire w_dff_B_faQGBYKa9_0;
	wire w_dff_B_3I5pooTO7_0;
	wire w_dff_B_cfFB24pP0_0;
	wire w_dff_B_f9d0InF66_0;
	wire w_dff_B_YbfPydN56_0;
	wire w_dff_B_K80VNsHQ9_0;
	wire w_dff_B_eu2N1W3a8_0;
	wire w_dff_B_h2MQXie50_0;
	wire w_dff_B_ikzr0D3R1_0;
	wire w_dff_B_8PARjvWG7_0;
	wire w_dff_B_Svtva3j69_0;
	wire w_dff_B_Q6D2xxis9_0;
	wire w_dff_B_Wu2J385L5_0;
	wire w_dff_B_wGIDmibr0_0;
	wire w_dff_B_k2OEKT3Z2_0;
	wire w_dff_B_D44JhL0K2_0;
	wire w_dff_B_J0R6U13T8_0;
	wire w_dff_B_KaEd3tYK1_0;
	wire w_dff_B_ayg7Z1Jg7_0;
	wire w_dff_B_7wKYrfz42_0;
	wire w_dff_B_s1IFzW6e3_0;
	wire w_dff_B_KpSIdnJ37_0;
	wire w_dff_B_h7OzLhJK2_0;
	wire w_dff_B_i0PS1ePd4_0;
	wire w_dff_B_td55wW7w2_0;
	wire w_dff_B_7IFs5pdC3_0;
	wire w_dff_B_xwjNpZHV8_0;
	wire w_dff_B_7dkg0NBF5_0;
	wire w_dff_B_4Qpql1583_0;
	wire w_dff_B_G0Ooledi7_0;
	wire w_dff_B_mxh4ADsU8_0;
	wire w_dff_B_8gkTUaR25_0;
	wire w_dff_B_hSsav01T8_0;
	wire w_dff_B_ExAZPzVT2_0;
	wire w_dff_B_NTBAdT9P8_0;
	wire w_dff_B_mqYykUGY5_0;
	wire w_dff_B_NeAK7oRq0_0;
	wire w_dff_B_D8ClRm555_0;
	wire w_dff_B_xQhJdJjm4_0;
	wire w_dff_B_GxAMHFJ85_0;
	wire w_dff_B_qCQkSwOJ7_0;
	wire w_dff_B_U7lz97841_0;
	wire w_dff_B_bdOq4ceS9_0;
	wire w_dff_B_2tHVEpgi4_0;
	wire w_dff_B_tQoTk3u53_0;
	wire w_dff_B_k9QxEl460_0;
	wire w_dff_B_sEuHC5Mo6_0;
	wire w_dff_B_GinDUmHK9_0;
	wire w_dff_B_UZoZTpXC5_0;
	wire w_dff_B_cENIvTQT9_0;
	wire w_dff_B_f1xhoyIn4_0;
	wire w_dff_B_gKQuFc3l4_0;
	wire w_dff_B_IklnBEV54_0;
	wire w_dff_B_4WXZG6qv3_0;
	wire w_dff_B_2QXrUTUd8_0;
	wire w_dff_B_BaobjH3z8_0;
	wire w_dff_B_VbI1f1PP7_0;
	wire w_dff_B_r9Uzvsxa5_0;
	wire w_dff_B_yANSEPOJ6_0;
	wire w_dff_B_QK4P1QL93_0;
	wire w_dff_B_rtWKMnH03_0;
	wire w_dff_B_z2V96TGI1_0;
	wire w_dff_B_foUP6z4Q3_0;
	wire w_dff_B_htV8mfbF1_0;
	wire w_dff_B_ckD0w8RQ1_0;
	wire w_dff_B_34LSAjkY5_0;
	wire w_dff_B_I6ywWay94_0;
	wire w_dff_B_RYCCcu415_0;
	wire w_dff_B_5VobtnOs3_0;
	wire w_dff_B_mOQrCJ1g5_0;
	wire w_dff_B_hn22zHpw6_0;
	wire w_dff_B_OzpXqPiS3_0;
	wire w_dff_B_op4UQWkT3_0;
	wire w_dff_B_ropqRbhv4_0;
	wire w_dff_B_3oPLHGCN9_0;
	wire w_dff_B_NYqGAdoD6_0;
	wire w_dff_B_woMA8ku71_0;
	wire w_dff_B_q0pQxjt75_0;
	wire w_dff_B_naGqQuvO9_0;
	wire w_dff_B_I2oui9Xr6_0;
	wire w_dff_B_SwzWSLWO7_0;
	wire w_dff_B_EpZcCx541_0;
	wire w_dff_B_M9fh4NkT3_0;
	wire w_dff_B_mHcw9xNn8_0;
	wire w_dff_B_ysMQwcks0_0;
	wire w_dff_B_cIUo5hLy3_0;
	wire w_dff_B_vb3gKBLM7_0;
	wire w_dff_B_gYVT3xAL8_0;
	wire w_dff_B_JGeRqTgp0_0;
	wire w_dff_B_f9vcm3833_0;
	wire w_dff_B_GLGQKuXA2_0;
	wire w_dff_B_hJxcmQD65_0;
	wire w_dff_B_9KGl4FJm0_0;
	wire w_dff_B_lwNpq0MP0_0;
	wire w_dff_B_teryKs1E9_0;
	wire w_dff_B_ROpempxJ7_0;
	wire w_dff_B_atGRPXTu2_0;
	wire w_dff_B_b6Vmd6hu6_0;
	wire w_dff_B_xWQbYHu12_0;
	wire w_dff_B_MRurAhZu9_0;
	wire w_dff_B_KmfeMXeL1_0;
	wire w_dff_B_B0RNuat01_0;
	wire w_dff_B_xgkKze5a9_0;
	wire w_dff_B_LsEJxYeO3_0;
	wire w_dff_B_2xberylD4_0;
	wire w_dff_B_Wm3uww6j6_0;
	wire w_dff_B_RdooBz740_0;
	wire w_dff_B_rO48ehu66_0;
	wire w_dff_B_AzJFvXw91_0;
	wire w_dff_B_WrBPJO8w1_0;
	wire w_dff_B_jfiZURSu5_0;
	wire w_dff_B_dBqZMyST8_0;
	wire w_dff_B_SrYfIE7g4_0;
	wire w_dff_B_6IN9eImK6_0;
	wire w_dff_B_ScKd0CFw6_0;
	wire w_dff_B_jN7t1Vlh5_0;
	wire w_dff_B_9YeI7Kyf2_0;
	wire w_dff_B_v8tqkuBK2_0;
	wire w_dff_B_AaTuoEnF4_0;
	wire w_dff_B_wPQSnwg69_0;
	wire w_dff_B_1aNURhaJ6_0;
	wire w_dff_B_7rLlObMg7_0;
	wire w_dff_B_2RtrFZ1t1_0;
	wire w_dff_B_2WrZcO8O9_0;
	wire w_dff_B_3jRpLMvD3_0;
	wire w_dff_B_hiPsxWSI4_0;
	wire w_dff_B_S7PtYfzw0_0;
	wire w_dff_B_jxVEOjI58_0;
	wire w_dff_B_E1DGR5EH1_0;
	wire w_dff_B_pVqGtZit6_0;
	wire w_dff_B_Q5zWN9L96_0;
	wire w_dff_B_hLOJOK031_0;
	wire w_dff_B_OBw3k05s3_0;
	wire w_dff_B_mtmqLYXP7_0;
	wire w_dff_B_nbM3Jkn44_0;
	wire w_dff_B_EMQIW3ku3_0;
	wire w_dff_B_MO27MXk02_0;
	wire w_dff_B_pNgJRW8u2_0;
	wire w_dff_B_S7QUpJyY1_0;
	wire w_dff_B_PKjSGtUM3_0;
	wire w_dff_B_S4E3W6KN6_0;
	wire w_dff_B_1nhqSAKw3_0;
	wire w_dff_B_YCGHBEaW3_0;
	wire w_dff_B_VEAuRrIs0_0;
	wire w_dff_B_1etwaut50_0;
	wire w_dff_B_EEwoF9t74_0;
	wire w_dff_B_Cgg5vZzs0_0;
	wire w_dff_B_riVnUW115_0;
	wire w_dff_B_faeJll4c4_0;
	wire w_dff_B_kr0Y06bI5_0;
	wire w_dff_B_TGDg4Fxd3_0;
	wire w_dff_B_e7RI90VD9_0;
	wire w_dff_B_rxoS4dAY3_0;
	wire w_dff_B_i0tfqvMv1_0;
	wire w_dff_B_Z1AMaSaV8_0;
	wire w_dff_B_f6ZQH2494_0;
	wire w_dff_B_qbc8uBF02_0;
	wire w_dff_B_sykpQlV87_0;
	wire w_dff_B_1vaM9zZZ1_0;
	wire w_dff_B_szIUk8025_0;
	wire w_dff_B_xfmlBT012_0;
	wire w_dff_B_qjDb8Fo38_0;
	wire w_dff_B_fwgvE4TM6_0;
	wire w_dff_B_VpZyQ5rH6_0;
	wire w_dff_B_wOI1fQRM1_0;
	wire w_dff_B_fH6asaQR3_0;
	wire w_dff_B_1VBKnOCE2_0;
	wire w_dff_B_4k1t9D9Y9_0;
	wire w_dff_B_4MrxxEGB2_0;
	wire w_dff_B_q5yKBMhs4_0;
	wire w_dff_B_2BOfN6Q42_0;
	wire w_dff_B_VBPAzVx42_0;
	wire w_dff_B_ch7qP2NG1_0;
	wire w_dff_B_RKgqDM6U0_0;
	wire w_dff_B_zStsKIT92_0;
	wire w_dff_B_iQLqDQQa3_0;
	wire w_dff_B_jqAhKNPr6_0;
	wire w_dff_B_vXuMHGEW4_0;
	wire w_dff_B_p9tLmpFF4_0;
	wire w_dff_B_iEAyHtIg5_0;
	wire w_dff_B_aEReYzTB6_0;
	wire w_dff_B_QakGROrO1_0;
	wire w_dff_B_HQk9F0Lb4_0;
	wire w_dff_B_VWxzcZ9V8_0;
	wire w_dff_B_oyjkip7Q4_0;
	wire w_dff_B_HymvBPt40_0;
	wire w_dff_B_V683s9sJ4_0;
	wire w_dff_B_7p9o18fa3_0;
	wire w_dff_B_e7FJUkZD6_0;
	wire w_dff_B_1MKuaGmE3_0;
	wire w_dff_B_t93lsMUY1_0;
	wire w_dff_B_YoIkeLTo9_0;
	wire w_dff_B_m7xcYI0O7_0;
	wire w_dff_B_2ZJhUVNi1_0;
	wire w_dff_B_6UITKluf8_0;
	wire w_dff_B_jJ0IIAdr6_0;
	wire w_dff_B_e3sHNQI22_0;
	wire w_dff_B_rpCByu2K5_0;
	wire w_dff_B_UQJWJHC32_0;
	wire w_dff_B_9Ag1LGdL7_0;
	wire w_dff_B_DwXTjwsP2_0;
	wire w_dff_B_aoUktpXP3_0;
	wire w_dff_B_YxtDK2ns4_0;
	wire w_dff_B_KzlEm6Bm6_0;
	wire w_dff_B_ZpH52zS71_0;
	wire w_dff_B_sFUX0Vcj1_0;
	wire w_dff_B_lJORFGME9_0;
	wire w_dff_B_yxViGg4Z0_0;
	wire w_dff_B_SLWZZrER1_0;
	wire w_dff_B_n3tpDtvk4_0;
	wire w_dff_B_KFl4aPQk8_0;
	wire w_dff_B_vLRY4kvG6_0;
	wire w_dff_B_vrhL2Odi7_0;
	wire w_dff_B_NZ9iKc2M8_0;
	wire w_dff_B_DraEQZfK4_0;
	wire w_dff_B_x2KYQWpG7_0;
	wire w_dff_B_RlqI4oeM9_0;
	wire w_dff_B_bAGEFQEV4_0;
	wire w_dff_B_NIXTqOCw7_0;
	wire w_dff_B_5SrNQhXs1_0;
	wire w_dff_B_82bX7yMC9_0;
	wire w_dff_B_6WQrfXFa6_0;
	wire w_dff_B_0KcfeBgc0_0;
	wire w_dff_B_jXUP2hUX2_0;
	wire w_dff_B_G2shiP8a3_0;
	wire w_dff_B_gQgetMSG0_0;
	wire w_dff_B_vGY73Shj4_0;
	wire w_dff_B_x230VX6o2_0;
	wire w_dff_B_ITSwtqNg0_0;
	wire w_dff_B_wMKWB4GX3_0;
	wire w_dff_B_PPVQVJ4W0_0;
	wire w_dff_B_zW3vfONN5_0;
	wire w_dff_B_cQyTUBvz7_0;
	wire w_dff_B_e46jy3lO4_0;
	wire w_dff_B_Agii0MqL1_0;
	wire w_dff_B_KyY1UFWL3_0;
	wire w_dff_B_MRn3By8s7_0;
	wire w_dff_B_NzdugDE63_0;
	wire w_dff_B_ds7bxBFr3_0;
	wire w_dff_B_Z8d4rzGQ8_0;
	wire w_dff_B_x7i2vxLV7_0;
	wire w_dff_B_0D5LiEID7_0;
	wire w_dff_B_tv2RRyZy0_0;
	wire w_dff_B_vIJigdPa0_0;
	wire w_dff_B_N1hpe2jk4_0;
	wire w_dff_B_gzoHAuVw1_0;
	wire w_dff_B_IdfMHzSF1_0;
	wire w_dff_B_8EiCbJMz0_0;
	wire w_dff_B_UQGyPA3k6_0;
	wire w_dff_B_hgTGGOc43_0;
	wire w_dff_B_QpQdV85s5_0;
	wire w_dff_B_0Hoqw0ur1_0;
	wire w_dff_B_MwUmG7DW4_0;
	wire w_dff_B_2zi5FKpx8_0;
	wire w_dff_B_0f1eobwe8_0;
	wire w_dff_B_y052bCq92_0;
	wire w_dff_B_212jN4uS2_0;
	wire w_dff_B_SwnPAFRO8_0;
	wire w_dff_B_eHmUQnW99_0;
	wire w_dff_B_9nRjR8Ge1_0;
	wire w_dff_B_27INWU3O0_0;
	wire w_dff_B_xcDE6JbJ4_0;
	wire w_dff_B_35Zzwq683_0;
	wire w_dff_B_tZHTz3T80_0;
	wire w_dff_B_o3ojjpxb8_0;
	wire w_dff_B_K3RS2WYq3_0;
	wire w_dff_B_4DRHh5WT2_0;
	wire w_dff_B_mSflLm8e5_0;
	wire w_dff_B_DwvyECH30_0;
	wire w_dff_B_7cyNYUos6_0;
	wire w_dff_B_RVXe09fZ9_0;
	wire w_dff_B_ShfkVBKY4_0;
	wire w_dff_B_uOBXALGU9_0;
	wire w_dff_B_MGNhczvD5_0;
	wire w_dff_B_efcRf5aJ0_0;
	wire w_dff_B_404BsHmB4_0;
	wire w_dff_B_ZJdyszo40_0;
	wire w_dff_B_8zkucMzy0_0;
	wire w_dff_B_nrXNRODy9_0;
	wire w_dff_B_YTEajDhQ3_0;
	wire w_dff_B_iufXdTah5_0;
	wire w_dff_B_wLLIM7pj7_0;
	wire w_dff_B_N8mw2iaZ6_0;
	wire w_dff_B_I1xd5Q4t7_0;
	wire w_dff_B_OID3XpKU5_0;
	wire w_dff_B_zegGqo9K6_0;
	wire w_dff_B_BXAUWvT53_0;
	wire w_dff_B_OBBaTtj89_0;
	wire w_dff_B_mRCC0SPp1_0;
	wire w_dff_B_0BCVMXHX7_0;
	wire w_dff_B_VD3swhdo6_0;
	wire w_dff_B_aBjHiLyJ1_0;
	wire w_dff_B_ggOBYlC84_0;
	wire w_dff_B_cT2vDEWf8_0;
	wire w_dff_B_ut9FwjEy7_0;
	wire w_dff_B_cK8zPTj01_0;
	wire w_dff_B_RXPWPRzV5_0;
	wire w_dff_B_kPeAOuBD7_0;
	wire w_dff_B_jyeDho8c0_0;
	wire w_dff_B_uJdXKlai3_0;
	wire w_dff_B_xcaW26FH7_0;
	wire w_dff_B_T0Uq0v029_0;
	wire w_dff_B_34VbIJNH2_0;
	wire w_dff_B_0mp5ciba5_0;
	wire w_dff_B_wZxhmfKh1_0;
	wire w_dff_B_oqJu9l2M4_0;
	wire w_dff_B_Yf6Y7Qkm6_0;
	wire w_dff_B_VWqbhx1M7_0;
	wire w_dff_B_kHA0vOpM4_0;
	wire w_dff_B_nzF5mTP21_0;
	wire w_dff_B_mGRIYUKt8_0;
	wire w_dff_B_FWkg8djd8_0;
	wire w_dff_B_1OfimBcA7_0;
	wire w_dff_B_fx0rMpml0_0;
	wire w_dff_B_nJV9S1V85_0;
	wire w_dff_B_11Rp9fqm3_0;
	wire w_dff_B_8m9eHZXG5_0;
	wire w_dff_B_6UM1RTYG6_0;
	wire w_dff_B_9YbEg9pz2_0;
	wire w_dff_B_Q2i4jHJO6_0;
	wire w_dff_B_OznLmD8I1_0;
	wire w_dff_B_XKRgdknm6_0;
	wire w_dff_B_Ws4EjfI20_0;
	wire w_dff_B_9i1h24cq5_0;
	wire w_dff_B_DVy0fdLL7_0;
	wire w_dff_B_JlFHpbuF3_0;
	wire w_dff_B_puJfkekU4_0;
	wire w_dff_B_JYGiK5QG0_0;
	wire w_dff_B_8yzjh6dk0_0;
	wire w_dff_B_9LrSMCjv1_0;
	wire w_dff_B_SkSkI2WZ1_0;
	wire w_dff_B_uvsy7iJp5_0;
	wire w_dff_B_VwIXG8d25_0;
	wire w_dff_B_AkHjRKZN6_0;
	wire w_dff_B_IZTrinxD5_0;
	wire w_dff_B_XGyR95ZE2_0;
	wire w_dff_B_leeQw8rV5_0;
	wire w_dff_B_dbT628Vt1_0;
	wire w_dff_B_pwFhYqJa4_0;
	wire w_dff_B_99DJbLNY6_0;
	wire w_dff_B_BdhYscDh8_0;
	wire w_dff_B_fkXlF58S2_0;
	wire w_dff_B_fQiq6p2n4_0;
	wire w_dff_B_eCA2PY434_0;
	wire w_dff_B_ldcyIKZa3_0;
	wire w_dff_B_4rXeWAsx1_0;
	wire w_dff_B_Z3uASZtT0_0;
	wire w_dff_B_gf7kSrln3_0;
	wire w_dff_B_cgt4YXwf3_0;
	wire w_dff_B_kjUTgarz4_0;
	wire w_dff_B_DVUSMd3i4_0;
	wire w_dff_B_5Er3MTwe5_0;
	wire w_dff_B_vOhFNWy42_0;
	wire w_dff_B_5nUDXCC78_0;
	wire w_dff_B_7ldrUj3E3_0;
	wire w_dff_B_Q9tuIgl56_0;
	wire w_dff_B_70D0ZeN33_0;
	wire w_dff_B_IuMLLEF52_0;
	wire w_dff_B_rl0s45Hr5_0;
	wire w_dff_B_nBOkQzRW5_0;
	wire w_dff_B_IwDOjdtB9_0;
	wire w_dff_B_zePLxlzP2_0;
	wire w_dff_B_MrjC0Nsf0_0;
	wire w_dff_B_9BbWUDOQ9_0;
	wire w_dff_B_jkPyd1S97_0;
	wire w_dff_B_jvG7E53V9_0;
	wire w_dff_B_5Jo5qCoR7_0;
	wire w_dff_B_BYloEgoh5_0;
	wire w_dff_B_W53dzSHP3_0;
	wire w_dff_B_RzY5B0Ih6_0;
	wire w_dff_B_nXhlz6th7_0;
	wire w_dff_B_4ommtaw37_0;
	wire w_dff_B_5QIuwX2U4_0;
	wire w_dff_B_qZB9Bp031_0;
	wire w_dff_B_bofmnyac9_0;
	wire w_dff_B_N6cgR2tm7_0;
	wire w_dff_B_OE2ZdGDa7_0;
	wire w_dff_B_HgEHpkiR6_0;
	wire w_dff_B_bW5lx9K62_0;
	wire w_dff_B_wL4lbu5R9_0;
	wire w_dff_B_2HSkl1IC8_0;
	wire w_dff_B_36IAP31z6_0;
	wire w_dff_B_iK5aSvpx3_0;
	wire w_dff_B_Gejfezgl4_0;
	wire w_dff_B_dpREpI1S1_0;
	wire w_dff_B_xYMoj03v2_0;
	wire w_dff_B_x5s7SwfV5_0;
	wire w_dff_B_2fiKOFhJ7_0;
	wire w_dff_B_ozZFYezY5_0;
	wire w_dff_B_LGvLSvvD5_0;
	wire w_dff_B_bZi1lRHb1_0;
	wire w_dff_B_ff5GhsKM6_0;
	wire w_dff_B_ZdVKEATP0_0;
	wire w_dff_B_UZdRAZsF9_0;
	wire w_dff_B_GsetXVEG7_0;
	wire w_dff_B_38BnUpEY1_0;
	wire w_dff_B_vwLiHdnA7_0;
	wire w_dff_B_elyoLX7k0_0;
	wire w_dff_B_r45bNTik4_0;
	wire w_dff_B_wQU9GMd80_0;
	wire w_dff_B_9G1Awdc28_0;
	wire w_dff_B_yWAJKTy82_0;
	wire w_dff_B_x1qxu2m24_0;
	wire w_dff_B_sTDLdOkr7_0;
	wire w_dff_B_mMr1X3771_0;
	wire w_dff_B_VrrlWfUi7_0;
	wire w_dff_B_ZOYtTr2Y4_0;
	wire w_dff_B_iyWXhSBQ3_0;
	wire w_dff_B_D0Xw5fND1_0;
	wire w_dff_B_3jIFMp7Q2_0;
	wire w_dff_B_mcjqYnyk6_0;
	wire w_dff_B_9aVcTZ3Y9_0;
	wire w_dff_B_FpwJ6Q869_0;
	wire w_dff_B_w8O0C1gR8_0;
	wire w_dff_B_StbFnvXe7_0;
	wire w_dff_B_TEAACXXo2_0;
	wire w_dff_B_kw2VL7qC3_0;
	wire w_dff_B_bnlnVv9T9_0;
	wire w_dff_B_Odk6xkZY2_0;
	wire w_dff_B_wK6zk5NY4_0;
	wire w_dff_B_4eyLIK714_0;
	wire w_dff_B_enxBNapu3_0;
	wire w_dff_B_ARkgyqWn6_0;
	wire w_dff_B_aEspfCFZ7_0;
	wire w_dff_B_tADwWlsu9_0;
	wire w_dff_B_x73SyZpA3_0;
	wire w_dff_B_s8VjViHO6_0;
	wire w_dff_B_lggMrUCL2_0;
	wire w_dff_B_pN0pcOoO4_0;
	wire w_dff_B_zAf7mVbR5_0;
	wire w_dff_B_KZq9pLel7_0;
	wire w_dff_B_rzJcUxmw4_0;
	wire w_dff_B_fcTx2uAt0_0;
	wire w_dff_B_sqP8r64f5_0;
	wire w_dff_B_RGgWpfJX5_0;
	wire w_dff_B_FGsJKvD37_0;
	wire w_dff_B_AW3xLrzy1_0;
	wire w_dff_B_OI2C8o5U0_0;
	wire w_dff_B_RBkikNet9_0;
	wire w_dff_B_n9rM7yTo3_0;
	wire w_dff_B_Ku1mdLTr4_0;
	wire w_dff_B_wmDNkcw54_0;
	wire w_dff_B_ZOuSm1ZR2_0;
	wire w_dff_B_pmPJUOSx3_0;
	wire w_dff_B_OHhZ9ZR25_0;
	wire w_dff_B_PMhGhtTo9_0;
	wire w_dff_B_kVKoFsj77_0;
	wire w_dff_B_EGEXzWU93_0;
	wire w_dff_B_1OCYNory6_0;
	wire w_dff_B_nr5bGOBE5_0;
	wire w_dff_B_ELDzrqbW5_0;
	wire w_dff_B_TQAXlIAK4_0;
	wire w_dff_B_DhS8Ndcu3_0;
	wire w_dff_B_uh6izZ3S4_0;
	wire w_dff_B_AYDG4Pbd6_0;
	wire w_dff_B_fvzIQwTD7_0;
	wire w_dff_B_ulGJImFW4_0;
	wire w_dff_B_vwMgjcE08_0;
	wire w_dff_B_RUcxmNUm8_0;
	wire w_dff_B_uSh4msnA3_0;
	wire w_dff_B_jCAhsPsG8_0;
	wire w_dff_B_Q0DEtEDD9_0;
	wire w_dff_B_xGzCzgYc1_0;
	wire w_dff_B_47OiT29x9_0;
	wire w_dff_B_sjIkIasD6_0;
	wire w_dff_B_HL4vSb0i3_0;
	wire w_dff_B_GEubLeZ76_0;
	wire w_dff_B_eGuVSfhE3_0;
	wire w_dff_B_mWzpjlr73_0;
	wire w_dff_B_pPKBXpYt4_0;
	wire w_dff_B_ZKo11Bso6_0;
	wire w_dff_B_1xSGfU5p7_0;
	wire w_dff_B_oZEFHgBT9_0;
	wire w_dff_B_rizs14Rv1_0;
	wire w_dff_B_3Vr6j7Op8_0;
	wire w_dff_B_rCzTFrsx2_0;
	wire w_dff_B_SrrZ8mhG1_0;
	wire w_dff_B_mnuMK0k33_0;
	wire w_dff_B_w3hqzGoA0_0;
	wire w_dff_B_0TK6Qbt07_0;
	wire w_dff_B_pHykt49I6_0;
	wire w_dff_B_utkvrmZc7_0;
	wire w_dff_B_DkLiLsCZ5_0;
	wire w_dff_B_g23GuXx38_0;
	wire w_dff_B_hZb0JHan7_0;
	wire w_dff_B_Bx7CoowZ0_0;
	wire w_dff_B_X2L28eJj8_0;
	wire w_dff_B_eRGJXM1a2_0;
	wire w_dff_B_23mVQqz58_0;
	wire w_dff_B_xnHP6Dda9_0;
	wire w_dff_B_cf45dtR64_0;
	wire w_dff_B_lLthOjPU7_0;
	wire w_dff_B_80iKDJKN0_0;
	wire w_dff_B_vC3WVPAy4_0;
	wire w_dff_B_iUbw8r529_0;
	wire w_dff_B_qVWscI2K4_0;
	wire w_dff_B_UiUFMzzk8_0;
	wire w_dff_B_kNH1NCLK2_0;
	wire w_dff_B_NRWs1TjP5_0;
	wire w_dff_B_LOKC2fWL6_0;
	wire w_dff_B_8XA5MRG59_0;
	wire w_dff_B_5hP75AeK5_0;
	wire w_dff_B_CpvMz4mN2_0;
	wire w_dff_B_8TvSFsgr7_0;
	wire w_dff_B_skCZuw8K6_0;
	wire w_dff_B_yM04tRlt4_0;
	wire w_dff_B_R2yF4jim3_0;
	wire w_dff_B_6f3dN7QN8_0;
	wire w_dff_B_gDrtT0l58_0;
	wire w_dff_B_3MMhsFCd0_0;
	wire w_dff_B_kQ1dnboA2_0;
	wire w_dff_B_urpsbfi53_0;
	wire w_dff_B_MVOLU3ws7_0;
	wire w_dff_B_mvmwfVA57_0;
	wire w_dff_B_oDDBxuIg1_0;
	wire w_dff_B_fdSxHe9t4_0;
	wire w_dff_B_GFar60K43_0;
	wire w_dff_B_e4YMGjjT1_0;
	wire w_dff_B_WpG0zDRd4_0;
	wire w_dff_B_UtCXg2np6_0;
	wire w_dff_B_D3hAIm7G6_0;
	wire w_dff_B_L9ET4TqU5_0;
	wire w_dff_B_LTiPZO7K5_0;
	wire w_dff_B_LJ1iqzgF4_0;
	wire w_dff_B_yvo7MTYZ8_0;
	wire w_dff_B_UqTuvFWY4_0;
	wire w_dff_B_vUGz1A9w7_0;
	wire w_dff_B_hmjJ8dgr7_0;
	wire w_dff_B_RrUiokRv8_0;
	wire w_dff_B_jnL9yvYN9_0;
	wire w_dff_B_Ev7GUK5u2_0;
	wire w_dff_B_3tiwEpoL1_0;
	wire w_dff_B_VmvndDKD0_0;
	wire w_dff_B_WqPYqotT9_0;
	wire w_dff_B_meG3HzrP3_0;
	wire w_dff_B_GvEgjppo1_0;
	wire w_dff_B_24eN53Uy1_0;
	wire w_dff_B_x8EtnUJm3_0;
	wire w_dff_B_RBaqlklD2_0;
	wire w_dff_B_qIOzllUj9_0;
	wire w_dff_B_rF9TcJz53_0;
	wire w_dff_B_R4OJcZS96_0;
	wire w_dff_B_mWedHaVg3_0;
	wire w_dff_B_8cuSA7pD9_0;
	wire w_dff_B_O4Kzfig71_0;
	wire w_dff_B_UNVoVzip5_0;
	wire w_dff_B_CSnIVTiN1_0;
	wire w_dff_B_ybU4RxjG7_0;
	wire w_dff_B_HZggoPB68_0;
	wire w_dff_B_YQeXZEzV6_0;
	wire w_dff_B_DFALM1Vp0_0;
	wire w_dff_B_WRu66ThJ8_0;
	wire w_dff_B_SeIvU6JH0_0;
	wire w_dff_B_0c5FSzV43_0;
	wire w_dff_B_eft00hZo3_0;
	wire w_dff_B_M3z591OZ9_0;
	wire w_dff_B_DAlnCixT3_0;
	wire w_dff_B_480fpUpr1_0;
	wire w_dff_B_ygXPRUIH7_0;
	wire w_dff_B_H3ZEg4fS0_0;
	wire w_dff_B_OqYZB5g93_0;
	wire w_dff_B_LGS1kK4r4_0;
	wire w_dff_B_PihdAonI9_0;
	wire w_dff_B_q4GgwZBd6_0;
	wire w_dff_B_nkFkux7L2_0;
	wire w_dff_B_lrEKLnkW3_0;
	wire w_dff_B_gNWOrdoQ1_0;
	wire w_dff_B_Xv1sEiPb6_0;
	wire w_dff_B_WCh4pQGB0_0;
	wire w_dff_B_Ujz2OuiD1_0;
	wire w_dff_B_Hs7IZQoM5_0;
	wire w_dff_B_Dm54EjHG2_0;
	wire w_dff_B_87zPumQs9_0;
	wire w_dff_B_xfpY7DEM9_0;
	wire w_dff_B_GaJW3tMO1_0;
	wire w_dff_B_xcJtpljq5_0;
	wire w_dff_B_uOt7OzVK6_0;
	wire w_dff_B_7qeVJBD69_0;
	wire w_dff_B_yyuyMGT65_0;
	wire w_dff_B_zLZT0Tce6_0;
	wire w_dff_B_dS418c9I0_0;
	wire w_dff_B_VSsCDWao5_0;
	wire w_dff_B_RUBwzeCd5_0;
	wire w_dff_B_l0PYgtk60_0;
	wire w_dff_B_5ELIJgwc3_0;
	wire w_dff_B_Uz8gbmkX0_0;
	wire w_dff_B_brAe0uFP4_0;
	wire w_dff_B_OVIPcE9O7_0;
	wire w_dff_B_PupL3Jnj0_0;
	wire w_dff_B_Vx2dRgeS4_0;
	wire w_dff_B_RXjy7JkA5_0;
	wire w_dff_B_7OIIjJiv9_0;
	wire w_dff_B_tyhbdQX67_0;
	wire w_dff_B_sHGVczSf8_0;
	wire w_dff_B_vjNYtJUJ1_0;
	wire w_dff_B_jNUyLwVg0_0;
	wire w_dff_B_0hXimAm42_0;
	wire w_dff_B_g9lvzgj05_0;
	wire w_dff_B_nSFZB8ys0_0;
	wire w_dff_B_UNfF6J3U9_0;
	wire w_dff_B_RwnIKpvb8_0;
	wire w_dff_B_7RYfViia6_0;
	wire w_dff_B_guqjXXO03_0;
	wire w_dff_B_wxxFjGE56_0;
	wire w_dff_B_GPikOGZW1_0;
	wire w_dff_B_VdTOUKKa2_0;
	wire w_dff_B_m50nFDnK3_0;
	wire w_dff_B_oTXl1Gi04_0;
	wire w_dff_B_GNkyk62V2_0;
	wire w_dff_B_Nhts54gS1_0;
	wire w_dff_B_orZoKxgX9_0;
	wire w_dff_B_eYmwcwLz3_0;
	wire w_dff_B_vxh4chKb1_0;
	wire w_dff_B_O5XuocJf1_0;
	wire w_dff_B_qh0VNzGu2_0;
	wire w_dff_B_YlgCbFom8_0;
	wire w_dff_B_0JpBfqp46_0;
	wire w_dff_B_JyshFPPs6_0;
	wire w_dff_B_PPZZ7XJq1_0;
	wire w_dff_B_SbNY8Z5z6_0;
	wire w_dff_B_XuYarmnf2_0;
	wire w_dff_B_SgfYSBrd1_0;
	wire w_dff_B_jhOqBV6g7_0;
	wire w_dff_B_l5z5e8ni8_0;
	wire w_dff_B_mUrmYZRx9_0;
	wire w_dff_B_IJW5cSVS6_0;
	wire w_dff_B_aTXPPdsk3_0;
	wire w_dff_B_OwRqrd5q0_0;
	wire w_dff_B_MXU39VTA7_0;
	wire w_dff_B_zro1Avn13_0;
	wire w_dff_B_fJl1mHSm4_0;
	wire w_dff_B_AxD95VGg4_0;
	wire w_dff_B_vyxqTUgj3_0;
	wire w_dff_B_pofWpHeK6_0;
	wire w_dff_B_X7PrYFQ60_0;
	wire w_dff_B_DjC3kDmD0_0;
	wire w_dff_B_oXz1HTAS4_0;
	wire w_dff_B_wMNURBNE3_0;
	wire w_dff_B_6JZWmO0a8_0;
	wire w_dff_B_2ZXq0dxu8_0;
	wire w_dff_B_MxNAwhCS2_0;
	wire w_dff_B_bCxsUiei6_0;
	wire w_dff_B_9zTGPg8K3_0;
	wire w_dff_B_iARsXMcr3_0;
	wire w_dff_B_yT7kWIM38_0;
	wire w_dff_B_CRWWdflb4_0;
	wire w_dff_B_hZm8Mf0L9_0;
	wire w_dff_B_vz8V1pPd1_0;
	wire w_dff_B_GL4Grb4P3_0;
	wire w_dff_B_OBczsvOg4_0;
	wire w_dff_B_5KTdh6Ph9_0;
	wire w_dff_B_oeFDRw2b9_0;
	wire w_dff_B_7MhKQS0Y9_0;
	wire w_dff_B_7Or7W8OI3_0;
	wire w_dff_B_hGgjVT1m4_0;
	wire w_dff_B_cxQHbRrb4_0;
	wire w_dff_B_xdSkvs3I5_0;
	wire w_dff_B_rTwRzNAk7_0;
	wire w_dff_B_lf3cti9i9_0;
	wire w_dff_B_UfsG2AX90_0;
	wire w_dff_B_U6YoEVXG6_0;
	wire w_dff_B_W24lS6cO7_0;
	wire w_dff_B_yCVdShtp5_0;
	wire w_dff_B_a3YReHKm5_0;
	wire w_dff_B_H07vlX996_0;
	wire w_dff_B_p0WI3M5P7_0;
	wire w_dff_B_D8WtqPFi1_0;
	wire w_dff_B_XveV5cCh8_0;
	wire w_dff_B_tHAyiOmX3_0;
	wire w_dff_B_lm6QGgng2_0;
	wire w_dff_B_rJ30bGHP0_0;
	wire w_dff_B_93ISU1Se1_0;
	wire w_dff_B_QNtnG1XT5_0;
	wire w_dff_B_mbPHK5WD0_0;
	wire w_dff_B_U9DxhiUg5_0;
	wire w_dff_B_29c6tTxp3_0;
	wire w_dff_B_bGRpgUhq1_0;
	wire w_dff_B_vmCGCL2L4_0;
	wire w_dff_B_6uNI6KZv2_0;
	wire w_dff_B_9qI6ZFZn9_0;
	wire w_dff_B_9o382cXc3_0;
	wire w_dff_B_h3AaYqih9_0;
	wire w_dff_B_YaCtgqK82_0;
	wire w_dff_B_zanO9U3n3_0;
	wire w_dff_B_jBiVlFCR9_0;
	wire w_dff_B_kQXg7P1b7_0;
	wire w_dff_B_s5l04Gn46_0;
	wire w_dff_B_YZl2ArNk6_0;
	wire w_dff_B_dPN2vdxK9_0;
	wire w_dff_B_GOisHFjS3_0;
	wire w_dff_B_pg8VuWm85_0;
	wire w_dff_B_XFFpCov71_0;
	wire w_dff_B_4DmOdg1F0_0;
	wire w_dff_B_SztyR6N21_0;
	wire w_dff_B_cI1t0jWd4_0;
	wire w_dff_B_TYj3X4Pm0_0;
	wire w_dff_B_Ekk6QjLl5_0;
	wire w_dff_B_mUSciLFF7_0;
	wire w_dff_B_5TCqRFol3_0;
	wire w_dff_B_oQU9RbYs3_0;
	wire w_dff_B_j7ga9LeB6_0;
	wire w_dff_B_ltd9MiKv9_0;
	wire w_dff_B_bb7oX1hP5_0;
	wire w_dff_B_GzIPLYZ21_0;
	wire w_dff_B_Zl28QESE7_0;
	wire w_dff_B_uoX7Oait0_0;
	wire w_dff_B_UKPKORPl6_0;
	wire w_dff_B_YX7GABMR7_0;
	wire w_dff_B_U2ZnsQuv4_0;
	wire w_dff_B_JT82WYwF6_0;
	wire w_dff_B_apnq8xML3_0;
	wire w_dff_B_89uhpWyp0_0;
	wire w_dff_B_GIlVFjpc8_0;
	wire w_dff_B_muW3arSx4_0;
	wire w_dff_B_rlyya7Q45_0;
	wire w_dff_B_QZm4Rezf6_0;
	wire w_dff_B_1c7Ow9ex5_0;
	wire w_dff_B_1jNH5cUL4_0;
	wire w_dff_B_qbkdhUaH2_0;
	wire w_dff_B_VcCJnFgE2_0;
	wire w_dff_B_9tz9GHYq1_0;
	wire w_dff_B_ng2nA4ap7_0;
	wire w_dff_B_Q6yt5r8u4_0;
	wire w_dff_B_OGlxJj7O4_0;
	wire w_dff_B_xkBpH88v2_0;
	wire w_dff_B_nyNqJLOO5_0;
	wire w_dff_B_pj7yDpwE5_0;
	wire w_dff_B_Aq64c9ZN5_0;
	wire w_dff_B_XwKTvYa33_0;
	wire w_dff_B_P8lAmxvD7_0;
	wire w_dff_B_lmc9HCMD2_0;
	wire w_dff_B_eH62Bknl2_0;
	wire w_dff_B_m9vDMMVt4_0;
	wire w_dff_B_gfGgB88U4_0;
	wire w_dff_B_F95Yo3fz7_0;
	wire w_dff_B_C304g7ml1_0;
	wire w_dff_B_VNkkN1Qm1_0;
	wire w_dff_B_3k8weLLt7_0;
	wire w_dff_B_AyeCyypE6_0;
	wire w_dff_B_KrjLWKeI8_0;
	wire w_dff_B_MfQQ1Ux78_0;
	wire w_dff_B_3xIjYwtq8_0;
	wire w_dff_B_Pfm1yHMo5_0;
	wire w_dff_B_o7rBlzRd7_0;
	wire w_dff_B_aSXVF1Rs2_0;
	wire w_dff_B_bp9mHlMY2_0;
	wire w_dff_B_PFpFZXWe9_0;
	wire w_dff_B_djlnkOzk7_0;
	wire w_dff_B_h0WDq8K44_0;
	wire w_dff_B_63gHmbso9_0;
	wire w_dff_B_xtYKZpYA4_0;
	wire w_dff_B_I2OCK4JD0_0;
	wire w_dff_B_pvqwtDtB6_0;
	wire w_dff_B_7vugEMsJ2_0;
	wire w_dff_B_Rw2JWE0p7_0;
	wire w_dff_B_YpXZJu6A1_0;
	wire w_dff_B_NUMclR8m9_0;
	wire w_dff_B_Ohydm42G4_0;
	wire w_dff_B_lfNMoP7O0_0;
	wire w_dff_B_dh43NSpn4_0;
	wire w_dff_B_IAtPc13h2_0;
	wire w_dff_B_AX0gEQ749_0;
	wire w_dff_B_aGKJxMg95_0;
	wire w_dff_B_0DOMc9m97_0;
	wire w_dff_B_aNkRzRjd9_0;
	wire w_dff_B_FSOHVuNe4_0;
	wire w_dff_B_2fga3iRe5_0;
	wire w_dff_B_BVAOB23F3_0;
	wire w_dff_B_cQPiGk7P6_0;
	wire w_dff_B_cSBO8h2r9_0;
	wire w_dff_B_4O5uDLRc8_0;
	wire w_dff_B_mRhuBEzX7_0;
	wire w_dff_B_trsMTfJV7_0;
	wire w_dff_B_hs0bIqB05_0;
	wire w_dff_B_YuHPHLcZ5_0;
	wire w_dff_B_CKv0lEqe8_0;
	wire w_dff_B_0pCnJL7O1_0;
	wire w_dff_B_69MVTQxo8_0;
	wire w_dff_B_yX6tNH4N1_0;
	wire w_dff_B_YHoNSSNz7_0;
	wire w_dff_B_OrKrD8ZZ4_0;
	wire w_dff_B_kEuOdEsw4_0;
	wire w_dff_B_CKTaj6S72_0;
	wire w_dff_B_4mjVS48m6_0;
	wire w_dff_B_2HaBSoxF6_0;
	wire w_dff_B_OJZiK74L5_0;
	wire w_dff_B_iuslrgjc1_0;
	wire w_dff_B_R4X4vpoZ1_0;
	wire w_dff_B_6b6Ll4sr8_0;
	wire w_dff_B_0nen7ZoL0_0;
	wire w_dff_B_o5fE4GQ61_0;
	wire w_dff_B_pdB5P6nR6_0;
	wire w_dff_B_yrAlxNKZ0_0;
	wire w_dff_B_dO9dIBhX7_0;
	wire w_dff_B_PkSPLW072_0;
	wire w_dff_B_xiWc8TLK1_0;
	wire w_dff_B_lWhkR4ix3_0;
	wire w_dff_B_BU5Wzufg0_0;
	wire w_dff_B_J9WR5ZO72_0;
	wire w_dff_B_UosIINje5_0;
	wire w_dff_B_Ua7JFNbw0_0;
	wire w_dff_B_3oYeOmZE3_0;
	wire w_dff_B_cu7jrV3J3_0;
	wire w_dff_B_kpU3coUu6_0;
	wire w_dff_B_8L7DzqaR0_0;
	wire w_dff_B_esNMC7tL1_0;
	wire w_dff_B_yPwD44Iu3_0;
	wire w_dff_B_APOZFSFv5_0;
	wire w_dff_B_CWbYvsI17_0;
	wire w_dff_B_bdOlm3cp4_0;
	wire w_dff_B_bNXFubr90_0;
	wire w_dff_B_EEk01UaF8_0;
	wire w_dff_B_5EmVVvVd1_0;
	wire w_dff_B_oDm5FM826_0;
	wire w_dff_B_sMpz7B927_0;
	wire w_dff_B_i9iZlJfX8_0;
	wire w_dff_B_NFjNaAnv6_0;
	wire w_dff_B_wRkKeCvy3_0;
	wire w_dff_B_5tUusbz36_0;
	wire w_dff_B_PISKIqu05_0;
	wire w_dff_B_xHl8NOXM2_0;
	wire w_dff_B_lJWcNF2S1_0;
	wire w_dff_B_NjINS3uI3_0;
	wire w_dff_B_wlpGhfkl6_0;
	wire w_dff_B_v4RJQEfZ1_0;
	wire w_dff_B_OykUYMHQ7_0;
	wire w_dff_B_WPxIS6nV9_0;
	wire w_dff_B_y2gUNXh91_0;
	wire w_dff_B_qhYrMvwl3_0;
	wire w_dff_B_QibSu3MY0_0;
	wire w_dff_B_CrpXcl3L2_0;
	wire w_dff_B_XpzuIzld0_0;
	wire w_dff_B_dAExRaPu8_0;
	wire w_dff_B_CbTwYaLV0_0;
	wire w_dff_B_fv8mqUCh1_0;
	wire w_dff_B_89q5qkTY6_0;
	wire w_dff_B_Jn5J4HWP8_0;
	wire w_dff_B_tS5qMp922_0;
	wire w_dff_B_XYkhcZ5o5_0;
	wire w_dff_B_5oKoSGR99_0;
	wire w_dff_B_e0jBCEhW3_0;
	wire w_dff_B_4wpRwwEq3_0;
	wire w_dff_B_ymYVUOHL6_0;
	wire w_dff_B_Vw6llRE23_0;
	wire w_dff_B_PGzrBREj0_0;
	wire w_dff_B_pNTLlTIs9_0;
	wire w_dff_B_Hgrqy4jd9_0;
	wire w_dff_B_VvfcyPt59_0;
	wire w_dff_B_eeyNjUxG1_0;
	wire w_dff_B_u6K5nWz25_0;
	wire w_dff_B_pHriOpf62_0;
	wire w_dff_B_Ta2w5qNi1_0;
	wire w_dff_B_pZiIGT1H6_0;
	wire w_dff_B_hj2McUWr9_0;
	wire w_dff_B_K1KhT9JZ7_0;
	wire w_dff_B_YeW3yzi12_0;
	wire w_dff_B_FHk8Cm157_0;
	wire w_dff_B_3diL9t954_0;
	wire w_dff_B_CK8pLLj75_0;
	wire w_dff_B_OWI6VM5D4_0;
	wire w_dff_B_T0tTv2gd1_0;
	wire w_dff_B_GoTtdasZ9_0;
	wire w_dff_B_JZ0JOwL22_0;
	wire w_dff_B_ePoI6xiD8_0;
	wire w_dff_B_k6da1RbX4_0;
	wire w_dff_B_jaMlvBPg1_0;
	wire w_dff_B_fVVQV1n03_0;
	wire w_dff_B_j4anH7x76_0;
	wire w_dff_B_Wd8YoPrp2_0;
	wire w_dff_B_XunoqiqL6_0;
	wire w_dff_B_zt26dltR8_0;
	wire w_dff_B_MHc159FP6_0;
	wire w_dff_B_OlSTHSpf3_0;
	wire w_dff_B_4jV0ufxc0_0;
	wire w_dff_B_TG7EVUyF9_0;
	wire w_dff_B_gaWTXJfm1_0;
	wire w_dff_B_gQNYQKJR8_0;
	wire w_dff_B_FlbRwU2r1_0;
	wire w_dff_B_mX2v2CdV1_0;
	wire w_dff_B_OXjDVGjo3_0;
	wire w_dff_B_wKVifQ5f3_0;
	wire w_dff_B_1s8CBTXJ6_0;
	wire w_dff_B_PWFs6dZC6_0;
	wire w_dff_B_iCdOhtuk0_0;
	wire w_dff_B_EhGyXncz5_0;
	wire w_dff_B_xUKp0f8C8_0;
	wire w_dff_B_X80eaCwq1_0;
	wire w_dff_B_jiRS4z6o0_0;
	wire w_dff_B_tSNFly4b2_0;
	wire w_dff_B_VghliOnV8_0;
	wire w_dff_B_yEEv1zRe9_0;
	wire w_dff_B_F5HqIpao2_0;
	wire w_dff_B_c52XXpUA5_0;
	wire w_dff_B_0cXD8FQ38_0;
	wire w_dff_B_LNcVVJ9d0_0;
	wire w_dff_B_RU6yi0Qa3_0;
	wire w_dff_B_q09krvnU6_0;
	wire w_dff_B_0fo4sWsv3_0;
	wire w_dff_B_Lh9Y4DgO6_0;
	wire w_dff_B_fxLWi57l9_0;
	wire w_dff_B_y3sNygWR4_0;
	wire w_dff_B_EGbb2BET2_0;
	wire w_dff_B_49lUd3Sc1_0;
	wire w_dff_B_oXqwIjFO6_0;
	wire w_dff_B_2wnl7G8F9_0;
	wire w_dff_B_vPkjnst92_0;
	wire w_dff_B_tAmjocYI1_0;
	wire w_dff_B_j1i98p4f2_0;
	wire w_dff_B_ehXNnoXo2_0;
	wire w_dff_B_RcTolzv66_0;
	wire w_dff_B_oDb0BsKV0_0;
	wire w_dff_B_dcP9bSpQ5_0;
	wire w_dff_B_FAGp2f471_0;
	wire w_dff_B_eqmpm2GS2_0;
	wire w_dff_B_frSjzcuQ7_0;
	wire w_dff_B_vaFtvecJ7_0;
	wire w_dff_B_573kwaHL6_0;
	wire w_dff_B_KD4ObqjU1_0;
	wire w_dff_B_QA0shmqH6_0;
	wire w_dff_B_R1KPK5NJ0_0;
	wire w_dff_B_lQzeQN2u2_0;
	wire w_dff_B_XP6iymHU6_0;
	wire w_dff_B_frHC1SBb8_0;
	wire w_dff_B_31GTaWVV9_0;
	wire w_dff_B_W2uokUDX2_0;
	wire w_dff_B_XiXwICzV1_0;
	wire w_dff_B_0QqotNMq2_0;
	wire w_dff_B_zByqVL7c6_0;
	wire w_dff_B_eRYks9G98_0;
	wire w_dff_B_LdPmKlDJ3_0;
	wire w_dff_B_sfLimVBe8_0;
	wire w_dff_B_VIj0WmHF4_0;
	wire w_dff_B_QdNx6xj44_0;
	wire w_dff_B_wEb8Cs8S4_0;
	wire w_dff_B_MTgufgRd8_0;
	wire w_dff_B_hJv1keCv8_0;
	wire w_dff_B_MnU9pBJ17_0;
	wire w_dff_B_yJ8aqfJh2_0;
	wire w_dff_B_prLBWnEz1_0;
	wire w_dff_B_hjICNjmV5_0;
	wire w_dff_B_5ZnERbT50_0;
	wire w_dff_B_cVKHtW8N3_0;
	wire w_dff_B_UlkkA3XK1_0;
	wire w_dff_B_de56BOYi1_0;
	wire w_dff_B_1cD3vLbb4_0;
	wire w_dff_B_RYSkFlHW0_0;
	wire w_dff_B_epEwuMPm3_0;
	wire w_dff_B_LKugcwPw5_0;
	wire w_dff_B_A71mZpmU4_0;
	wire w_dff_B_z3akaDy54_0;
	wire w_dff_B_PKlVr9y60_0;
	wire w_dff_B_H1Ismx8S3_0;
	wire w_dff_B_ktnydPjl3_0;
	wire w_dff_B_W3Qac7z77_0;
	wire w_dff_B_R9mKPtUn2_0;
	wire w_dff_B_F2p7XeCT4_0;
	wire w_dff_B_m2GGTYQT1_0;
	wire w_dff_B_aQY9Vmue7_0;
	wire w_dff_B_xGN0Qqyt1_0;
	wire w_dff_B_fiuvY00G3_0;
	wire w_dff_B_aHO5VoQR0_0;
	wire w_dff_B_xQiSzY7V8_0;
	wire w_dff_B_iZFrfk9X7_0;
	wire w_dff_B_5OkbODOr5_0;
	wire w_dff_B_q7LqM9db3_0;
	wire w_dff_B_JYo2tjZt9_0;
	wire w_dff_B_BNeCqfF61_0;
	wire w_dff_B_lOIOhChm2_0;
	wire w_dff_B_QURScThB4_0;
	wire w_dff_B_ALmUfoUf8_0;
	wire w_dff_B_a5BqRznn5_0;
	wire w_dff_B_VE4kZJhC9_0;
	wire w_dff_B_j4MSl7Rl9_0;
	wire w_dff_B_C7b4GfIv0_0;
	wire w_dff_B_V6i0CRwj5_0;
	wire w_dff_B_1sZ7BzvQ7_0;
	wire w_dff_B_ZnChadNt0_0;
	wire w_dff_B_qQaYDmDp7_0;
	wire w_dff_B_G2hJzBq82_0;
	wire w_dff_B_Ycgvm1YK5_0;
	wire w_dff_B_C33CuETS7_0;
	wire w_dff_B_yPPObXP35_0;
	wire w_dff_B_tn4ZeCnK3_0;
	wire w_dff_B_pRYBAsFm7_0;
	wire w_dff_B_IrTON0Rr9_0;
	wire w_dff_B_2Y63atFT6_0;
	wire w_dff_B_rQNt04901_0;
	wire w_dff_B_JSfahvmV3_0;
	wire w_dff_B_IikKiVcf9_0;
	wire w_dff_B_ribwdkTf7_0;
	wire w_dff_B_pmANmI7m5_0;
	wire w_dff_B_37boURr84_0;
	wire w_dff_B_oNmT3o6l0_0;
	wire w_dff_B_Yt4gJOsA6_0;
	wire w_dff_B_96cPcaDV0_0;
	wire w_dff_B_JtbCCNnA0_0;
	wire w_dff_B_T0jVaiTr8_0;
	wire w_dff_B_AeZXTDz20_0;
	wire w_dff_B_LBHc8Nmn0_0;
	wire w_dff_B_NrqR9U6x4_0;
	wire w_dff_B_7D8Ni5ge8_0;
	wire w_dff_B_iV2cyu5Y3_0;
	wire w_dff_B_xaTPwzlo0_0;
	wire w_dff_B_1WGYhbD68_0;
	wire w_dff_B_l42Cru9g5_0;
	wire w_dff_B_LrX6lbra8_0;
	wire w_dff_B_bGSFoYhO9_0;
	wire w_dff_B_saKLDtS28_0;
	wire w_dff_B_6A7hocPr3_0;
	wire w_dff_B_yCU0xiTF1_0;
	wire w_dff_B_TtB7TcO89_0;
	wire w_dff_B_pIunSuZN1_0;
	wire w_dff_B_KhsCuYaB6_0;
	wire w_dff_B_OcbUrppn6_0;
	wire w_dff_B_PCXjid5C4_0;
	wire w_dff_B_y6Eorlus8_0;
	wire w_dff_B_owIG0yJ06_0;
	wire w_dff_B_Ln4sFxsX2_0;
	wire w_dff_B_eKwGPw7V8_0;
	wire w_dff_B_OlmF5qTe4_0;
	wire w_dff_B_5SYs1ChX1_0;
	wire w_dff_B_FOkIB6aE9_0;
	wire w_dff_B_2xMjHazF1_0;
	wire w_dff_B_ZrCyTODv6_0;
	wire w_dff_B_de0Eltu84_0;
	wire w_dff_B_dNu5LnJL2_0;
	wire w_dff_B_mAg1Ma4N2_0;
	wire w_dff_B_eUV9qe9P0_0;
	wire w_dff_B_u4s8MfAV2_0;
	wire w_dff_B_QI4t88Im4_0;
	wire w_dff_B_3Re7f7gr6_0;
	wire w_dff_B_LrvPmcfc6_0;
	wire w_dff_B_Jpyr0i3p5_0;
	wire w_dff_B_rgNpTVNe8_0;
	wire w_dff_B_hRgMZVDQ0_0;
	wire w_dff_B_8CMIGMki7_0;
	wire w_dff_B_8r5sT5Hj9_0;
	wire w_dff_B_agKJkgO88_0;
	wire w_dff_B_5tUUvYSs5_0;
	wire w_dff_B_SUUYl2Ql6_0;
	wire w_dff_B_2Kcfu0Ow9_0;
	wire w_dff_B_V3CPQKV23_0;
	wire w_dff_B_h8dfXeo67_0;
	wire w_dff_B_6fmHsrpf9_0;
	wire w_dff_B_vv05b3pP6_0;
	wire w_dff_B_iv0OTOHd3_0;
	wire w_dff_B_Lo11yvdl1_0;
	wire w_dff_B_pCR9Yfr53_0;
	wire w_dff_B_SPDzZlbu0_0;
	wire w_dff_B_XMqaOnrd7_0;
	wire w_dff_B_2FGhGH2k2_0;
	wire w_dff_B_k6gdoh4L9_0;
	wire w_dff_B_OEcg16PF4_0;
	wire w_dff_B_VuLpQPGO9_0;
	wire w_dff_B_FrmXP06D2_0;
	wire w_dff_B_geqgFR811_0;
	wire w_dff_B_20cXzEjq0_0;
	wire w_dff_B_moPeNJNd9_0;
	wire w_dff_B_N3qEAfNq3_0;
	wire w_dff_B_GtfoM1uq0_0;
	wire w_dff_B_pmoeat4U0_0;
	wire w_dff_B_E3ZUZcLs9_0;
	wire w_dff_B_ehJMKFQM6_0;
	wire w_dff_B_3XzqoR0D2_0;
	wire w_dff_B_ajXEGd817_0;
	wire w_dff_B_ZStMTwQe6_0;
	wire w_dff_B_q9ucs9dJ6_0;
	wire w_dff_B_22wiXwxE9_0;
	wire w_dff_B_Lk1S6Kbi7_0;
	wire w_dff_B_66sgbL4g3_0;
	wire w_dff_B_aTILEKEi7_0;
	wire w_dff_B_33JP8V1O5_0;
	wire w_dff_B_on5EDIln4_0;
	wire w_dff_B_MR96iNia7_0;
	wire w_dff_B_CDWAS9cZ7_0;
	wire w_dff_B_g9mHbIN76_0;
	wire w_dff_B_pXakBqg36_0;
	wire w_dff_B_1KvY9WdL1_0;
	wire w_dff_B_AqTpSvBg9_0;
	wire w_dff_B_ARkWtLDg2_0;
	wire w_dff_B_RVxQSl9z2_0;
	wire w_dff_B_MXapfCiO0_0;
	wire w_dff_B_NiJgqczZ6_0;
	wire w_dff_B_pJBJs51D7_0;
	wire w_dff_B_6VXoqg1k7_0;
	wire w_dff_B_a53JGxks9_0;
	wire w_dff_B_EvjNB68H3_0;
	wire w_dff_B_w96ba0o01_0;
	wire w_dff_B_jBxV5ZP92_0;
	wire w_dff_B_KBm0uTY37_0;
	wire w_dff_B_cu6Mvi1O3_0;
	wire w_dff_B_RHlAZacF5_0;
	wire w_dff_B_unqY8mlw0_0;
	wire w_dff_B_egQMpBlX8_0;
	wire w_dff_B_7EMz2fWV0_0;
	wire w_dff_B_frwXzutk5_0;
	wire w_dff_B_XoAPZ96H2_0;
	wire w_dff_B_VxpdCQyE4_0;
	wire w_dff_B_5nGgvKrc1_0;
	wire w_dff_B_EpWcbXQC9_0;
	wire w_dff_B_ikShCIX86_0;
	wire w_dff_B_MDGgDhvE2_0;
	wire w_dff_B_uO2yOCfx7_0;
	wire w_dff_B_AFpSPMYN9_0;
	wire w_dff_B_cTffIZWH2_0;
	wire w_dff_B_3ECHQIaU1_0;
	wire w_dff_B_F2Lyayif5_0;
	wire w_dff_B_6GcnVHFK3_0;
	wire w_dff_B_z70llqHZ0_0;
	wire w_dff_B_fuXnMRtv2_0;
	wire w_dff_B_UkzBpdJk3_0;
	wire w_dff_B_1KN2rOI35_0;
	wire w_dff_B_NDLYw4BX6_0;
	wire w_dff_B_4DQBQDm09_0;
	wire w_dff_B_0wTDjqhf0_0;
	wire w_dff_B_wblBllOt5_0;
	wire w_dff_B_ZlLBXL0q4_0;
	wire w_dff_B_IvDHNfVi3_0;
	wire w_dff_B_aGRkfmxy1_0;
	wire w_dff_B_tMWeQkwK3_0;
	wire w_dff_B_7mcESinR8_0;
	wire w_dff_B_w75cR5T45_0;
	wire w_dff_B_JgN08Anm3_0;
	wire w_dff_B_aFyF0oj45_0;
	wire w_dff_B_z4yGXYRC6_0;
	wire w_dff_B_NJX6h7iV3_0;
	wire w_dff_B_jkmHeVEt0_0;
	wire w_dff_B_M1OaGsg82_0;
	wire w_dff_B_n41gK4eS7_0;
	wire w_dff_B_UyrT6NAh6_0;
	wire w_dff_B_9rc0CAUg3_0;
	wire w_dff_B_pHlugRtT4_0;
	wire w_dff_B_1Nga2AzP5_0;
	wire w_dff_B_m0CZFsE05_0;
	wire w_dff_B_i6zH9xfd3_0;
	wire w_dff_B_cOdCS9p96_0;
	wire w_dff_B_bmx66jTE1_0;
	wire w_dff_B_5BYT7Hkh0_0;
	wire w_dff_B_iQ3YF5Pz9_0;
	wire w_dff_B_vC48mWBm1_0;
	wire w_dff_B_gwewANYg9_0;
	wire w_dff_B_y0CcsUWT2_0;
	wire w_dff_B_15W38iue0_0;
	wire w_dff_B_AlQcuCud8_0;
	wire w_dff_B_pNiayghy5_0;
	wire w_dff_B_0QBYYCfx6_0;
	wire w_dff_B_kSbs4dz32_0;
	wire w_dff_B_SYPE1Myu0_0;
	wire w_dff_B_gjU2VSrl5_0;
	wire w_dff_B_gIhryTrY2_0;
	wire w_dff_B_GGTpIqzJ3_0;
	wire w_dff_B_1sYlDTx17_0;
	wire w_dff_B_KHzhYfHX4_0;
	wire w_dff_B_sVLdLstf7_0;
	wire w_dff_B_aBDnNtof8_0;
	wire w_dff_B_rrcyax9y5_0;
	wire w_dff_B_iG7hTRaU5_0;
	wire w_dff_B_7FQBMSLZ2_0;
	wire w_dff_B_rrhZqAUJ7_0;
	wire w_dff_B_XAhX8icl7_0;
	wire w_dff_B_MHuBcaSt0_0;
	wire w_dff_B_WVMFfHbY1_0;
	wire w_dff_B_o7VqJYbT7_0;
	wire w_dff_B_SmeeZ4tL6_0;
	wire w_dff_B_73IF7KRg3_0;
	wire w_dff_B_BxbavUD39_0;
	wire w_dff_B_CHIrgCrR3_0;
	wire w_dff_B_LYTy6ISu5_0;
	wire w_dff_B_cquNgXv40_0;
	wire w_dff_B_HddT7aXK1_0;
	wire w_dff_B_9yP5DuKQ0_0;
	wire w_dff_B_PJMw2XNx9_0;
	wire w_dff_B_xYQ7Zcz49_0;
	wire w_dff_B_OCt7ZsUi7_0;
	wire w_dff_B_vtGN0D4r3_0;
	wire w_dff_B_YOwd49Y06_0;
	wire w_dff_B_XFNrNkxe1_0;
	wire w_dff_B_U4mECs0r7_0;
	wire w_dff_B_rXOMJpwB3_0;
	wire w_dff_B_NFllEoXk6_0;
	wire w_dff_B_0QsMHnpL9_0;
	wire w_dff_B_Twnfa97T6_0;
	wire w_dff_B_G6YcFTpg6_0;
	wire w_dff_B_vZZIn7do3_0;
	wire w_dff_B_9azuofPq2_0;
	wire w_dff_B_URUsk3MO0_0;
	wire w_dff_B_8wd0pn7A4_0;
	wire w_dff_B_8HpPVXXn4_0;
	wire w_dff_B_rGoXWfzz2_0;
	wire w_dff_B_1VWRbAFr3_0;
	wire w_dff_B_YsYCyOqW2_0;
	wire w_dff_B_QcCldeJf2_0;
	wire w_dff_B_REoL3ClF6_0;
	wire w_dff_B_rPfnGHDG2_0;
	wire w_dff_B_2fmDeasB9_0;
	wire w_dff_B_2I7LxLKF3_0;
	wire w_dff_B_baT2ARg28_0;
	wire w_dff_B_i2OGFSEI6_0;
	wire w_dff_B_670Xcgpe5_0;
	wire w_dff_B_QKAwfh3j5_0;
	wire w_dff_B_ZAFVuXJo2_0;
	wire w_dff_B_h9Owkg0i8_0;
	wire w_dff_B_jaV6vv2Y7_0;
	wire w_dff_B_SS39PbM01_0;
	wire w_dff_B_0mdxo3WL3_0;
	wire w_dff_B_Dsizarx17_0;
	wire w_dff_B_LEMRb8hz5_0;
	wire w_dff_B_8WRodDgi5_0;
	wire w_dff_B_2IYgpU4x5_0;
	wire w_dff_B_YfZSMbct1_0;
	wire w_dff_B_tJuO6fUj4_0;
	wire w_dff_B_4fDFzSel4_0;
	wire w_dff_B_OcSOR1jH6_0;
	wire w_dff_B_ybIv3Zc71_0;
	wire w_dff_B_1BAhsGEk5_0;
	wire w_dff_B_aO7mvjEi6_0;
	wire w_dff_B_buV9XsNC1_0;
	wire w_dff_B_KIVOnZwv2_0;
	wire w_dff_B_6yGBRLHY8_0;
	wire w_dff_B_j58iVanm4_0;
	wire w_dff_B_Pot2UTII2_0;
	wire w_dff_B_gbxrcPo36_0;
	wire w_dff_B_02TqhYHf2_0;
	wire w_dff_B_aqT3dCPg1_0;
	wire w_dff_B_8cWEkuD12_0;
	wire w_dff_B_71nkVB5p6_0;
	wire w_dff_B_KhVTjIfx9_0;
	wire w_dff_B_vHLCZ4pF0_0;
	wire w_dff_B_VBVqxeLI0_0;
	wire w_dff_B_F4s63S5p8_0;
	wire w_dff_B_CgB0dbMi4_0;
	wire w_dff_B_NzYinipm2_0;
	wire w_dff_B_nw5wdooD7_0;
	wire w_dff_B_Uqg6pbIw5_0;
	wire w_dff_B_MiHvLnEP0_0;
	wire w_dff_B_FUf4G8331_0;
	wire w_dff_B_iwmOFbya2_0;
	wire w_dff_B_EjbaOgTM5_0;
	wire w_dff_B_qasx58sI4_0;
	wire w_dff_B_PTt5yt1J9_0;
	wire w_dff_B_Na910Bfd1_0;
	wire w_dff_B_VfwFG6rv0_0;
	wire w_dff_B_araAvJEA9_0;
	wire w_dff_B_8SlINF8p7_0;
	wire w_dff_B_4u3RNrBc6_0;
	wire w_dff_B_Fn2T9zcL1_0;
	wire w_dff_B_HW9stFUS1_0;
	wire w_dff_B_a6v2rfvp2_0;
	wire w_dff_B_sJNIWidZ7_0;
	wire w_dff_B_yqVr2DNA1_0;
	wire w_dff_B_ckxNXAPc9_0;
	wire w_dff_B_GnCUwiQs6_0;
	wire w_dff_B_TDWLEqX25_0;
	wire w_dff_B_RMrYRhzl6_0;
	wire w_dff_B_IVWHdDRC6_0;
	wire w_dff_B_1cZnVxff6_0;
	wire w_dff_B_fQ0SBGcg6_0;
	wire w_dff_B_vtqh0Ppx6_0;
	wire w_dff_B_CNSv9hMK0_0;
	wire w_dff_B_e2ljy7uB0_0;
	wire w_dff_B_xwfdHKxM6_0;
	wire w_dff_B_YljmDFe52_0;
	wire w_dff_B_BqZk7xP18_0;
	wire w_dff_B_Ox9dIUWk2_0;
	wire w_dff_B_diLv3GE92_0;
	wire w_dff_B_jwYYhK3T4_0;
	wire w_dff_B_JOmqquYs5_0;
	wire w_dff_B_fTNL12B76_0;
	wire w_dff_B_YfaYofbG5_0;
	wire w_dff_B_iiL6A9U45_0;
	wire w_dff_B_6fqUfEJI2_0;
	wire w_dff_B_A1vohAOT1_0;
	wire w_dff_B_mX6zUOKX6_0;
	wire w_dff_B_h1C0nFZh6_0;
	wire w_dff_B_gBJF0tbC8_0;
	wire w_dff_B_1NOccfLd7_0;
	wire w_dff_B_tUimDyCa2_0;
	wire w_dff_B_OMh5HBhk3_0;
	wire w_dff_B_7ANrYdw48_0;
	wire w_dff_B_ZYkWAQb59_0;
	wire w_dff_B_ay4qsUHV1_0;
	wire w_dff_B_nGVVSN2v8_0;
	wire w_dff_B_YYwv4BJ15_0;
	wire w_dff_B_bO379u7c7_0;
	wire w_dff_B_Y7VsG9id8_0;
	wire w_dff_B_63KiuyzB9_0;
	wire w_dff_B_M3eWBkSk1_0;
	wire w_dff_B_qNnEAjzs4_0;
	wire w_dff_B_zT7O8DQ47_0;
	wire w_dff_B_6NlwGPmf9_0;
	wire w_dff_B_UYLTsiUC7_0;
	wire w_dff_B_kWONCJSn0_0;
	wire w_dff_B_MS6IPvQu3_0;
	wire w_dff_B_TTOrtpJ42_0;
	wire w_dff_B_epvi4E0Y5_0;
	wire w_dff_B_jHtEUOk53_0;
	wire w_dff_B_Z7NnmeeY3_0;
	wire w_dff_B_c3F1Tnwz8_0;
	wire w_dff_B_O2CgCM2y4_0;
	wire w_dff_B_YueCyedn2_0;
	wire w_dff_B_XIit2uNM3_0;
	wire w_dff_B_FIH0O3PE7_0;
	wire w_dff_B_9QwMtVZH7_0;
	wire w_dff_B_iGBc7U835_0;
	wire w_dff_B_zOBFKmIG1_0;
	wire w_dff_B_Gv7OQc6a9_0;
	wire w_dff_B_w0ObPVLr6_0;
	wire w_dff_B_wB3P3ZDn1_0;
	wire w_dff_B_QoK31wgl6_0;
	wire w_dff_B_hDGfCOUa7_0;
	wire w_dff_B_rbEKOed13_0;
	wire w_dff_B_9w62NqoI9_0;
	wire w_dff_B_lQ7h7CId1_0;
	wire w_dff_B_q7eixNu19_0;
	wire w_dff_B_aVtERWWg4_0;
	wire w_dff_B_BYV83VVI8_0;
	wire w_dff_B_NVMMmkC14_0;
	wire w_dff_B_42vFMTZd7_0;
	wire w_dff_B_oJnJh0Uw9_0;
	wire w_dff_B_9B4L9QN64_0;
	wire w_dff_B_8vhDov6l6_0;
	wire w_dff_B_eAj6qN8B3_0;
	wire w_dff_B_e84rrwvS3_0;
	wire w_dff_B_Q1KJMv9w1_0;
	wire w_dff_B_JfafIsUy1_0;
	wire w_dff_B_kevNxul21_0;
	wire w_dff_B_XYjokHdl6_0;
	wire w_dff_B_7U2tDgcl9_0;
	wire w_dff_B_ZKGdyJ900_0;
	wire w_dff_B_U6u55A9L6_0;
	wire w_dff_B_uaMqcePb5_0;
	wire w_dff_B_6UHE639p7_0;
	wire w_dff_B_HPdYf0aL0_0;
	wire w_dff_B_RSD11qq79_0;
	wire w_dff_B_H7RRcInR7_0;
	wire w_dff_B_PE1dnht06_0;
	wire w_dff_B_CZNzxYcS2_0;
	wire w_dff_B_Rdfaso0W9_0;
	wire w_dff_B_DLKGojIZ2_0;
	wire w_dff_B_jSkpze7G8_0;
	wire w_dff_B_oPKN4p3d5_0;
	wire w_dff_B_trvscKgr9_0;
	wire w_dff_B_TA6RxhDI3_0;
	wire w_dff_B_T0eBvAu56_0;
	wire w_dff_B_jQFfflpp8_0;
	wire w_dff_B_QLtcTgWz4_0;
	wire w_dff_B_SVOxw2tu7_0;
	wire w_dff_B_vvg8Ulfn5_0;
	wire w_dff_B_Gm9NC6fF6_0;
	wire w_dff_B_qpx5BBst8_0;
	wire w_dff_B_xQHFDjek1_0;
	wire w_dff_B_1VKNp4vS6_0;
	wire w_dff_B_6cTdRamm7_0;
	wire w_dff_B_Wjjk8S1x1_0;
	wire w_dff_B_9vcuXYfz0_0;
	wire w_dff_B_Z57goe1K3_0;
	wire w_dff_B_XBATHLZS6_0;
	wire w_dff_B_0IwsHbfy0_0;
	wire w_dff_B_udcVLTQG1_0;
	wire w_dff_B_67W1r02d3_0;
	wire w_dff_B_VjDlzsGQ4_0;
	wire w_dff_B_jVm8dfvb6_0;
	wire w_dff_B_On0BB9t34_0;
	wire w_dff_B_plYGxNwq3_0;
	wire w_dff_B_cDzvERom3_0;
	wire w_dff_B_gUGUsPZu9_0;
	wire w_dff_B_ztDlVhTp2_0;
	wire w_dff_B_tYqDB4EN6_0;
	wire w_dff_B_3Iw6unZh7_0;
	wire w_dff_B_HqxgmXPU3_0;
	wire w_dff_B_P7HVCpYw4_0;
	wire w_dff_B_JdbqUIM05_0;
	wire w_dff_B_uoTaioss2_0;
	wire w_dff_B_xDWWmLjZ9_0;
	wire w_dff_B_G5EJpep07_0;
	wire w_dff_B_T2YmP8GL7_0;
	wire w_dff_B_nklgWzpH4_0;
	wire w_dff_B_ZXZWAm6g6_0;
	wire w_dff_B_eoEoJo673_0;
	wire w_dff_B_h222w6BG3_0;
	wire w_dff_B_hdWqmTW64_0;
	wire w_dff_B_Ysh7bVVO8_0;
	wire w_dff_B_Y1clmQ7b1_0;
	wire w_dff_B_ZeTPjXIe8_0;
	wire w_dff_B_QZq85zmY8_0;
	wire w_dff_B_XGWhxQsZ8_0;
	wire w_dff_B_IuCCrDRT4_0;
	wire w_dff_B_0fR7u6Ys5_0;
	wire w_dff_B_Uwelh4V23_0;
	wire w_dff_B_VLEBRs3r6_0;
	wire w_dff_B_rQHQqHXQ8_0;
	wire w_dff_B_ODsOWPSp4_0;
	wire w_dff_B_3CI9vcSz1_0;
	wire w_dff_B_HvbPgBVb0_0;
	wire w_dff_B_DeuWbQdY2_0;
	wire w_dff_B_jpdZv3Q25_0;
	wire w_dff_B_8t2ohWji8_0;
	wire w_dff_B_w6YHkdCv7_0;
	wire w_dff_B_HtldMgdf0_0;
	wire w_dff_B_xpuZ1OLr7_0;
	wire w_dff_B_PrRvLsxZ6_0;
	wire w_dff_B_gySG7fem7_0;
	wire w_dff_B_IETOyFW67_0;
	wire w_dff_B_sEJhzPr62_0;
	wire w_dff_B_nOL90Hyt4_0;
	wire w_dff_B_2DN8uHtl7_0;
	wire w_dff_B_Pvyl37zS4_0;
	wire w_dff_B_jvhB9CbW7_0;
	wire w_dff_B_wSYc1CNi4_0;
	wire w_dff_B_Q3ek2Oyw4_0;
	wire w_dff_B_F4JkyPU58_0;
	wire w_dff_B_SieVe3Ol3_0;
	wire w_dff_B_PpvYVAPT6_0;
	wire w_dff_B_EIeNnAz38_0;
	wire w_dff_B_tmuq0qS35_0;
	wire w_dff_B_KdnVXJbt6_0;
	wire w_dff_B_Rv8hatbY5_0;
	wire w_dff_B_ZI6fjHmS7_0;
	wire w_dff_B_Ov2dgGlC1_0;
	wire w_dff_B_zleW9DY09_0;
	wire w_dff_B_o0Tnxdyx7_0;
	wire w_dff_B_qJtkcBIK4_0;
	wire w_dff_B_19YzJv9I1_0;
	wire w_dff_B_XiworvY53_0;
	wire w_dff_B_6MPsd7W32_0;
	wire w_dff_B_yaiIkwHR2_0;
	wire w_dff_B_2s1cPYZF4_0;
	wire w_dff_B_93uEfT1T0_0;
	wire w_dff_B_JZXIks4y6_0;
	wire w_dff_B_71haXrJZ1_0;
	wire w_dff_B_srYQ604o0_0;
	wire w_dff_B_tvxMLiiL9_0;
	wire w_dff_B_LSWn1x8e5_0;
	wire w_dff_B_hXgbemVz2_0;
	wire w_dff_B_bgpFdUFS2_0;
	wire w_dff_B_X4EZn1M13_0;
	wire w_dff_B_eyySQIqE6_0;
	wire w_dff_B_JWtMNE7Q6_0;
	wire w_dff_B_2pVWTnaL9_0;
	wire w_dff_B_0tIW24Sl2_0;
	wire w_dff_B_qmsSJ3yW5_0;
	wire w_dff_B_0wvE8l2H8_0;
	wire w_dff_B_QvXXgIOR5_0;
	wire w_dff_B_za769sNV7_0;
	wire w_dff_B_HpMsnEni5_0;
	wire w_dff_B_uWMn5IYn4_0;
	wire w_dff_B_DKyQyM5R7_0;
	wire w_dff_B_cl13aeGR4_0;
	wire w_dff_B_Y5qPERVi0_0;
	wire w_dff_B_AEjyVo2L5_0;
	wire w_dff_B_83bwYSdd1_0;
	wire w_dff_B_oGYS17yU6_0;
	wire w_dff_B_o7cLntBr9_0;
	wire w_dff_B_nzpOFU7Q8_0;
	wire w_dff_B_kd2ksk6b2_0;
	wire w_dff_B_4D1wTTfc6_0;
	wire w_dff_B_SfVIvRmZ1_0;
	wire w_dff_B_5voHPdDr7_0;
	wire w_dff_B_968wELXU8_0;
	wire w_dff_B_lBy4Ms0D5_0;
	wire w_dff_B_xZski9ev2_0;
	wire w_dff_B_bWWERdDD8_0;
	wire w_dff_B_3wGUs2am8_0;
	wire w_dff_B_g2ZISok74_0;
	wire w_dff_B_B7YvaD4A2_0;
	wire w_dff_B_2PViXef75_0;
	wire w_dff_B_mEc9Ho3k7_0;
	wire w_dff_B_wgUGMa0p2_0;
	wire w_dff_B_zAhRoE9u1_0;
	wire w_dff_B_zRVI6D4X9_0;
	wire w_dff_B_GYP6yAdF9_0;
	wire w_dff_B_ntjSw7dF6_0;
	wire w_dff_B_5Zwip4k81_0;
	wire w_dff_B_jmDuG3Jx0_0;
	wire w_dff_B_DJXJUhZN3_0;
	wire w_dff_B_GQHpvbFz1_0;
	wire w_dff_B_QHVEtMsV2_0;
	wire w_dff_B_ouP5JOAq0_0;
	wire w_dff_B_cqES8raJ6_0;
	wire w_dff_B_jOXGfaj73_0;
	wire w_dff_B_HoMEbkSw9_0;
	wire w_dff_B_bgcegKWU2_0;
	wire w_dff_B_dd0p0oAi6_0;
	wire w_dff_B_pusv550R7_0;
	wire w_dff_B_ZfxIdoRS3_0;
	wire w_dff_B_rZly37lq9_0;
	wire w_dff_B_1QrxlgIi3_0;
	wire w_dff_B_EZ3bjkOA6_0;
	wire w_dff_B_atZEI2L26_0;
	wire w_dff_B_zN2WAg558_0;
	wire w_dff_B_oqDDBQ8k8_0;
	wire w_dff_B_sPJWm7tm8_0;
	wire w_dff_B_cx7ciW4N5_0;
	wire w_dff_B_8jr8A6wf2_0;
	wire w_dff_B_fKPhdPw80_0;
	wire w_dff_B_ArPEip2A9_0;
	wire w_dff_B_w6Y4u58X5_0;
	wire w_dff_B_DyWZwweL9_0;
	wire w_dff_B_NTvxV2DC0_0;
	wire w_dff_B_Vyjyv6Y98_0;
	wire w_dff_B_hj3vrpnk2_0;
	wire w_dff_B_Yx31Y2yi2_0;
	wire w_dff_B_wzDVvkSD5_0;
	wire w_dff_B_NkXuCfbI5_0;
	wire w_dff_B_ApEmhpxu8_0;
	wire w_dff_B_iXWoM0wB9_0;
	wire w_dff_B_FDhDBvSa8_0;
	wire w_dff_B_U9FQO6r42_0;
	wire w_dff_B_AobR9bnN8_0;
	wire w_dff_B_DGFQE7b14_0;
	wire w_dff_B_z9SRrJur5_0;
	wire w_dff_B_VDGxEkFo7_0;
	wire w_dff_B_CVH01MXj6_0;
	wire w_dff_B_DGJOucNC7_0;
	wire w_dff_B_T0dICz7U5_0;
	wire w_dff_B_B1x4mKxj2_0;
	wire w_dff_B_oJ9BwWfd6_0;
	wire w_dff_B_9UTPLhqN1_0;
	wire w_dff_B_4OocKqtL1_0;
	wire w_dff_B_TA3qS7rS4_0;
	wire w_dff_B_lZUXb3am7_0;
	wire w_dff_B_1ztAo8ZS5_0;
	wire w_dff_B_SAc63fLB8_0;
	wire w_dff_B_anKfKQCv4_0;
	wire w_dff_B_P4nZcRXe7_0;
	wire w_dff_B_iddLDsQe1_0;
	wire w_dff_B_ac51NJ8M5_0;
	wire w_dff_B_YcwgTnpQ1_0;
	wire w_dff_B_o0JTq3177_0;
	wire w_dff_B_V8yniEIl3_0;
	wire w_dff_B_w0bV01dU2_0;
	wire w_dff_B_cHBo464i5_0;
	wire w_dff_B_kzpLcWcb2_0;
	wire w_dff_B_R52MuZJ14_0;
	wire w_dff_B_nQfUyDek2_0;
	wire w_dff_B_EM6Q6fXr3_0;
	wire w_dff_B_39990Mc98_0;
	wire w_dff_B_K8OexuYb9_0;
	wire w_dff_B_wiGiQNyH2_0;
	wire w_dff_B_reHKeMie8_0;
	wire w_dff_B_npM5Nl0O6_0;
	wire w_dff_B_2OoijRqk8_0;
	wire w_dff_B_mxRnyncP0_0;
	wire w_dff_B_u2obqZvQ8_0;
	wire w_dff_B_23XQ23Vq8_0;
	wire w_dff_B_HOoJjIW81_0;
	wire w_dff_B_8jGzfMY66_0;
	wire w_dff_B_Y5OzA62R8_0;
	wire w_dff_B_x052kdxA0_0;
	wire w_dff_B_WvdaZn920_0;
	wire w_dff_B_gjdPgoE86_0;
	wire w_dff_B_nzfeVEXt0_0;
	wire w_dff_B_JJ9rG2Gu2_0;
	wire w_dff_B_ajN1aV6p4_0;
	wire w_dff_B_4S2NTSbc2_0;
	wire w_dff_B_XyATiomv8_0;
	wire w_dff_B_CctImZ677_0;
	wire w_dff_B_yUO1rcyV8_0;
	wire w_dff_B_G1nS78DA1_0;
	wire w_dff_B_UWTf4VsK0_0;
	wire w_dff_B_Yks2LHNj7_0;
	wire w_dff_B_fAbiPnOI4_0;
	wire w_dff_B_Eg504Qtb6_0;
	wire w_dff_B_JDOlONTx1_0;
	wire w_dff_B_2tZ2TT418_0;
	wire w_dff_B_bQwu2pKW1_0;
	wire w_dff_B_a5tYb59C2_0;
	wire w_dff_B_ggmU1zId5_0;
	wire w_dff_B_NpqnGBF81_0;
	wire w_dff_B_txZuw9hH9_0;
	wire w_dff_B_LE2yWl298_0;
	wire w_dff_B_Cs0dg0j89_0;
	wire w_dff_B_HQ0WDu3E9_0;
	wire w_dff_B_COKo5FpP0_0;
	wire w_dff_B_nWq3XiFw8_0;
	wire w_dff_B_o12N0bDT3_0;
	wire w_dff_B_TY8mE9Li0_0;
	wire w_dff_B_Im30cn4y5_0;
	wire w_dff_B_KF5ZAWdU8_0;
	wire w_dff_B_t9e84WK16_0;
	wire w_dff_B_k6pbRaNT3_0;
	wire w_dff_B_MKvpkoCF0_0;
	wire w_dff_B_Yf7m6c1S4_0;
	wire w_dff_B_3rPiMYEK0_0;
	wire w_dff_B_MtbNuX5Z5_0;
	wire w_dff_B_8RA9EyCE0_0;
	wire w_dff_B_1yniShmk4_0;
	wire w_dff_B_3j4nDcev0_0;
	wire w_dff_B_rz3GLmFp6_0;
	wire w_dff_B_Ud3Dy1Eo2_0;
	wire w_dff_B_k9DFeDPe2_0;
	wire w_dff_B_lZUCSA9A3_0;
	wire w_dff_B_fDZ95RFP3_0;
	wire w_dff_B_3GgoQRQw0_0;
	wire w_dff_B_MXq7WG1f2_0;
	wire w_dff_B_I8btYOZ85_0;
	wire w_dff_B_nFWX1Tk75_0;
	wire w_dff_B_rLp89D2B8_0;
	wire w_dff_B_L7Kwj1N42_0;
	wire w_dff_B_b12LLiXT2_0;
	wire w_dff_B_mwOIfAEw8_0;
	wire w_dff_B_W8EQbhah2_0;
	wire w_dff_B_GDLg9PZ15_0;
	wire w_dff_B_QYj8j4lR1_0;
	wire w_dff_B_9L6RF8JV8_0;
	wire w_dff_B_uznJy0lY2_0;
	wire w_dff_B_ziTfRZrj3_0;
	wire w_dff_B_UwgeImGO4_0;
	wire w_dff_B_nF1qfK8k2_0;
	wire w_dff_B_7H5KW3lH4_0;
	wire w_dff_B_BvI3xdZn8_0;
	wire w_dff_B_OaUTPC2v7_0;
	wire w_dff_B_trzzL8lt6_0;
	wire w_dff_B_VHdkFBLW9_0;
	wire w_dff_B_ah5RcUrR1_0;
	wire w_dff_B_JPiWC0wi9_0;
	wire w_dff_B_L5Pucexw8_0;
	wire w_dff_B_docg3eac9_0;
	wire w_dff_B_EttfWhTC3_0;
	wire w_dff_B_nSUBjaxG9_0;
	wire w_dff_B_bdW7SarL9_0;
	wire w_dff_B_Jjdj1cZ71_0;
	wire w_dff_B_BdHYiJcT4_0;
	wire w_dff_B_3HtbydAD1_0;
	wire w_dff_B_g9GROpv34_0;
	wire w_dff_B_LrwqCsfY0_0;
	wire w_dff_B_Db0V13Qf3_0;
	wire w_dff_B_wAxo6ZkR6_0;
	wire w_dff_B_hcyqwcDR8_0;
	wire w_dff_B_ncfYkBw05_0;
	wire w_dff_B_NEcMygc96_0;
	wire w_dff_B_MnPQDsx59_0;
	wire w_dff_B_BfVf1e9F2_0;
	wire w_dff_B_Pw2BAIRZ8_0;
	wire w_dff_B_ciTHcdW91_0;
	wire w_dff_B_oMPmOW1m6_0;
	wire w_dff_B_0aip3RuV9_0;
	wire w_dff_B_WCUJ3gjy9_0;
	wire w_dff_B_Y5Tp0Aqu1_0;
	wire w_dff_B_ZSVpoMic1_0;
	wire w_dff_B_lUKJVG9c5_0;
	wire w_dff_B_53hN5EYA5_0;
	wire w_dff_B_BuFh8Hxo2_0;
	wire w_dff_B_4P6ybyWZ9_0;
	wire w_dff_B_oBP6ETy65_0;
	wire w_dff_B_POlv0clL2_0;
	wire w_dff_B_GQ59k3ax2_0;
	wire w_dff_B_q8D3XDFy9_0;
	wire w_dff_B_H4XpqHqe1_0;
	wire w_dff_B_OG2uWAfO8_0;
	wire w_dff_B_1ZXxUS0t8_0;
	wire w_dff_B_uSbo473H4_0;
	wire w_dff_B_G0PN0gDH2_0;
	wire w_dff_B_nVnr4XIg6_0;
	wire w_dff_B_w5tC6RVB7_0;
	wire w_dff_B_Cwao2zTs7_0;
	wire w_dff_B_IHOCXAD78_0;
	wire w_dff_B_WD6Z4xBB3_0;
	wire w_dff_B_m56xR5qt0_0;
	wire w_dff_B_ceT84vat9_0;
	wire w_dff_B_CdsB3iVe2_0;
	wire w_dff_B_G2vBjQl91_0;
	wire w_dff_B_FzuzKVaR2_0;
	wire w_dff_B_OXEH8LOc4_0;
	wire w_dff_B_phXZYXDE9_0;
	wire w_dff_B_tJjvCFaF8_0;
	wire w_dff_B_CG3qYiiH9_0;
	wire w_dff_B_LGaA90wP8_0;
	wire w_dff_B_8qh9t5cc0_0;
	wire w_dff_B_GP7jMlkS5_0;
	wire w_dff_B_QZNtyzr55_0;
	wire w_dff_B_QXBGWgRV9_0;
	wire w_dff_B_QjiUcXlb3_0;
	wire w_dff_B_eAL6qBVp8_0;
	wire w_dff_B_pPhVScum2_0;
	wire w_dff_B_Wn6DD4PA5_0;
	wire w_dff_B_o5K0aP9q2_0;
	wire w_dff_B_x1rHUAFq1_0;
	wire w_dff_B_uuZXmYkW8_0;
	wire w_dff_B_mzYG1aHG2_0;
	wire w_dff_B_9qakpVN09_0;
	wire w_dff_B_zUZPMoaj8_0;
	wire w_dff_B_28AEySVh9_0;
	wire w_dff_B_L4vt9y447_0;
	wire w_dff_B_cIYLqHl43_0;
	wire w_dff_B_jV6OSf7h7_0;
	wire w_dff_B_ifZD6cu69_0;
	wire w_dff_B_WQMoiER83_0;
	wire w_dff_B_pFexGzC92_0;
	wire w_dff_B_JqB01Iod7_0;
	wire w_dff_B_p3DsJkDf3_0;
	wire w_dff_B_utjsIphL0_0;
	wire w_dff_B_Fg3yS2qD6_0;
	wire w_dff_B_TATfofGL1_0;
	wire w_dff_B_mWTzbsI77_0;
	wire w_dff_B_o03zHjcG7_0;
	wire w_dff_B_YY7BsTrf3_0;
	wire w_dff_B_KgQKlFF93_0;
	wire w_dff_B_Ttqi03tx6_0;
	wire w_dff_B_H2Dnf3dc2_0;
	wire w_dff_B_CM7jz7L08_0;
	wire w_dff_B_PGqEwNli6_0;
	wire w_dff_B_jZykDcjk1_0;
	wire w_dff_B_BGJcRS4d6_0;
	wire w_dff_B_fTkniR4A9_0;
	wire w_dff_B_ma8ElqK70_0;
	wire w_dff_B_jo4cFnr11_0;
	wire w_dff_B_t9ovZgvW0_0;
	wire w_dff_B_meG5Ji8a6_0;
	wire w_dff_B_UpNu6R1R2_0;
	wire w_dff_B_ltHfzfbS9_0;
	wire w_dff_B_pW1NiX0c2_0;
	wire w_dff_B_5mzjNiO58_0;
	wire w_dff_B_QXSd3mEE7_0;
	wire w_dff_B_XQFCNxae4_0;
	wire w_dff_B_E5PzlMqY3_0;
	wire w_dff_B_qJ6D9iMz5_0;
	wire w_dff_B_Uo8qwJ6z1_0;
	wire w_dff_B_lf3JsRov0_0;
	wire w_dff_B_fykQMdf01_0;
	wire w_dff_B_neOMRHVV8_0;
	wire w_dff_B_KXmHRlCq2_0;
	wire w_dff_B_dI6UbY0n8_0;
	wire w_dff_B_xy4ZFNtu2_0;
	wire w_dff_B_mNkORTe84_0;
	wire w_dff_B_QvfpEdGf5_0;
	wire w_dff_B_pJs4pl4V2_0;
	wire w_dff_B_VPSKlS1d6_0;
	wire w_dff_B_PYd4ZtCy6_0;
	wire w_dff_B_iiWokwY60_0;
	wire w_dff_B_WP0JqA5K8_0;
	wire w_dff_B_0gnvdIXO5_0;
	wire w_dff_B_ZrazR2MC9_0;
	wire w_dff_B_Bbw3HlHC5_0;
	wire w_dff_B_WLcoUUuU8_0;
	wire w_dff_B_bkixuBlO8_0;
	wire w_dff_B_MbqnRTuo1_0;
	wire w_dff_B_expjBXjo4_0;
	wire w_dff_B_f3hIg0vi4_0;
	wire w_dff_B_J1HiIVl22_0;
	wire w_dff_B_ZUkjynjR4_0;
	wire w_dff_B_gDu2FW9f1_0;
	wire w_dff_B_Lz0r841V0_0;
	wire w_dff_B_O4JdixWM3_0;
	wire w_dff_B_XSzpCLky9_0;
	wire w_dff_B_cCy6XunU8_0;
	wire w_dff_B_esXN1fYe4_0;
	wire w_dff_B_4464nAZJ1_0;
	wire w_dff_B_hfxWRCUC1_0;
	wire w_dff_B_3xPxFbc54_0;
	wire w_dff_B_hefYU6vU4_0;
	wire w_dff_B_AnswcnUc9_0;
	wire w_dff_B_nywxU3Bl1_0;
	wire w_dff_B_t4sWVa0J3_0;
	wire w_dff_B_dC93gKEJ0_0;
	wire w_dff_B_GgBrDkta4_0;
	wire w_dff_B_ATHHpgLz9_0;
	wire w_dff_B_C7TWCQnK1_0;
	wire w_dff_B_RnCEMxAh9_0;
	wire w_dff_B_N56pYF8L2_0;
	wire w_dff_B_4t2jEr5f5_0;
	wire w_dff_B_8ausr4H82_0;
	wire w_dff_B_sLFdCexR5_0;
	wire w_dff_B_wbwvO3oo7_0;
	wire w_dff_B_wO1NqDRk2_0;
	wire w_dff_B_OG4wtSEy2_0;
	wire w_dff_B_CJvIfNUT8_0;
	wire w_dff_B_SuZOm4Q02_0;
	wire w_dff_B_z1ngT9Rg6_0;
	wire w_dff_B_gObonihq8_0;
	wire w_dff_B_v6wFi9fD8_0;
	wire w_dff_B_Y2LleHzL0_0;
	wire w_dff_B_7VoU9dqQ5_0;
	wire w_dff_B_0xq9NL2h4_0;
	wire w_dff_B_Q61pZNZz9_0;
	wire w_dff_B_OW9Ii3kI4_0;
	wire w_dff_B_s59uKsJl0_0;
	wire w_dff_B_6njFsaYT2_0;
	wire w_dff_B_vmD25BkI0_0;
	wire w_dff_B_zz2aymKs5_0;
	wire w_dff_B_4ibYHJsS0_0;
	wire w_dff_B_RNywH5tF7_0;
	wire w_dff_B_FvakI0Qn7_0;
	wire w_dff_B_REl8PntW2_0;
	wire w_dff_B_cUKjUDVY3_0;
	wire w_dff_B_wGFMoWCr4_0;
	wire w_dff_B_E6lARNtU6_0;
	wire w_dff_B_d8vXLIM54_0;
	wire w_dff_B_I4LX4cDH5_0;
	wire w_dff_B_zmexGCnF8_0;
	wire w_dff_B_lxFPLiYd2_0;
	wire w_dff_B_9l76CoSq6_0;
	wire w_dff_B_lcFptnhE4_0;
	wire w_dff_B_09iEg04s5_0;
	wire w_dff_B_xYXRn8HT4_0;
	wire w_dff_B_rJQqSIF11_0;
	wire w_dff_B_aSuPJBe29_0;
	wire w_dff_B_WIH07Xkj5_0;
	wire w_dff_B_PM8o8nAm7_0;
	wire w_dff_B_bWTiumqj8_0;
	wire w_dff_B_nXRDLqzk4_0;
	wire w_dff_B_qKmbI41y7_0;
	wire w_dff_B_zr09pa7n1_0;
	wire w_dff_B_E4Vg84Lj1_0;
	wire w_dff_B_ZK5CgouX2_0;
	wire w_dff_B_Kygmbtdm2_0;
	wire w_dff_B_zn43aFR24_0;
	wire w_dff_B_lW7n09O32_0;
	wire w_dff_B_mh8cKYwj2_0;
	wire w_dff_B_Yxb7eyNY0_0;
	wire w_dff_B_i03DsB0k9_0;
	wire w_dff_B_WyresKMq8_0;
	wire w_dff_B_JKNycuHs1_0;
	wire w_dff_B_To6n4iMm1_0;
	wire w_dff_B_9nB2Bezx5_0;
	wire w_dff_B_KcmTXtoY7_0;
	wire w_dff_B_ZaQbYrLH4_0;
	wire w_dff_B_T6otSM9I4_0;
	wire w_dff_B_dCkkux5u4_0;
	wire w_dff_B_nzw6BVd93_0;
	wire w_dff_B_AaXqchK28_0;
	wire w_dff_B_6cDGnhpg6_0;
	wire w_dff_B_bXGxEJQW8_0;
	wire w_dff_B_wdMnH8Ff5_0;
	wire w_dff_B_3iKPHi4K4_0;
	wire w_dff_B_FXQ3W1k68_0;
	wire w_dff_B_GZmZOvaj2_0;
	wire w_dff_B_RugSlYs21_0;
	wire w_dff_B_3vL4qTJL9_0;
	wire w_dff_B_N5UCnsYn8_0;
	wire w_dff_B_JS5nSguM2_0;
	wire w_dff_B_XReSzSqK2_0;
	wire w_dff_B_xrc0AWSP3_0;
	wire w_dff_B_EZTMbPfY5_0;
	wire w_dff_B_NfwtV7ar1_0;
	wire w_dff_B_U52sDTsA5_0;
	wire w_dff_B_papPhMdP6_0;
	wire w_dff_B_TdB2oZHS9_0;
	wire w_dff_B_jokVzOCq4_0;
	wire w_dff_B_rsrwPn7Q8_0;
	wire w_dff_B_f7OWNSBZ7_0;
	wire w_dff_B_qb1B3slN1_0;
	wire w_dff_B_mQ6sCzV03_0;
	wire w_dff_B_swq2P9Ax7_0;
	wire w_dff_B_ubxnuARn6_0;
	wire w_dff_B_bZTzS0SK2_0;
	wire w_dff_B_HQFZrY3k8_0;
	wire w_dff_B_amZiA1wi7_0;
	wire w_dff_B_Lhi9rStt0_0;
	wire w_dff_B_KvAc0izF4_0;
	wire w_dff_B_l114WAU63_0;
	wire w_dff_B_IrusQLRo6_0;
	wire w_dff_B_zEafl3z17_0;
	wire w_dff_B_Ef8Ppp8R5_0;
	wire w_dff_B_ltokuBCR5_0;
	wire w_dff_B_RXaRnNG89_0;
	wire w_dff_B_lmXu2mHI5_0;
	wire w_dff_B_fllAp6r39_0;
	wire w_dff_B_XhtHh4Cf7_0;
	wire w_dff_B_49LT0sZG0_0;
	wire w_dff_B_XpAbIZSD0_0;
	wire w_dff_B_Z8IhUQBi1_0;
	wire w_dff_B_B74k7I7U6_0;
	wire w_dff_B_hPdAM3bS5_0;
	wire w_dff_B_zmgDIyvg3_0;
	wire w_dff_B_xW1z9eYL7_0;
	wire w_dff_B_R6P5RagF3_0;
	wire w_dff_B_VGb6Ptq23_0;
	wire w_dff_B_47S8cGDP4_0;
	wire w_dff_B_eF1Y3tH79_0;
	wire w_dff_B_8Ib1lwHk3_0;
	wire w_dff_B_oWJ2uPW18_0;
	wire w_dff_B_WGZrHuMM2_0;
	wire w_dff_B_Gww81NxQ2_0;
	wire w_dff_B_z0UvKrVS2_0;
	wire w_dff_B_OhcBtwwL3_0;
	wire w_dff_B_mKRHJEaT7_0;
	wire w_dff_B_fLTydxC90_0;
	wire w_dff_B_SOymH8sV5_0;
	wire w_dff_B_MkJLb7yg8_0;
	wire w_dff_B_1uxv8di55_0;
	wire w_dff_B_lcCQC9FS8_0;
	wire w_dff_B_ZHC8vifY5_0;
	wire w_dff_B_3IkOFxUB6_0;
	wire w_dff_B_ncqogXVe4_0;
	wire w_dff_B_3LCKPhW87_0;
	wire w_dff_B_ldADEgEZ5_0;
	wire w_dff_B_Ti0fmlFP6_0;
	wire w_dff_B_1EDzcKgC8_0;
	wire w_dff_B_YkuWKzVy2_0;
	wire w_dff_B_Va3GCSV01_0;
	wire w_dff_B_idmhnMSV1_0;
	wire w_dff_B_z1JUa0KP3_0;
	wire w_dff_B_bm3uN25j4_0;
	wire w_dff_B_xgu7Fjgx7_0;
	wire w_dff_B_y8TBpVZY7_0;
	wire w_dff_B_5w3PXRDA6_0;
	wire w_dff_B_FKK7EtMa7_0;
	wire w_dff_B_tI9tqR8K8_0;
	wire w_dff_B_1A03e1BA0_0;
	wire w_dff_B_l0vnjnHH8_0;
	wire w_dff_B_o4NfDfSU4_0;
	wire w_dff_B_toxmDRH98_0;
	wire w_dff_B_8NjOG2gv0_0;
	wire w_dff_B_mw76b3jb4_0;
	wire w_dff_B_7EhcehT73_0;
	wire w_dff_B_IEqH6rZa1_0;
	wire w_dff_B_seimVXrJ4_0;
	wire w_dff_B_TYRcfwl23_0;
	wire w_dff_B_GNfOxe4K6_0;
	wire w_dff_B_ZfYPFTUU8_0;
	wire w_dff_B_fYLTMBXi1_0;
	wire w_dff_B_29YjHbro9_0;
	wire w_dff_B_JIb0ZRqE7_0;
	wire w_dff_B_LyjLC9yF7_0;
	wire w_dff_B_coRleIV87_0;
	wire w_dff_B_1vJFv3ZA9_0;
	wire w_dff_B_UoItZ67J8_0;
	wire w_dff_B_9eDKA3c71_0;
	wire w_dff_B_WU8fFmwC2_0;
	wire w_dff_B_hCzyrGpy3_0;
	wire w_dff_B_N2aM87v43_0;
	wire w_dff_B_pYnbF4kV5_0;
	wire w_dff_B_dSTR5RCM6_0;
	wire w_dff_B_FB6kOVCH1_0;
	wire w_dff_B_GR5pGJRg3_0;
	wire w_dff_B_Dd0LCtA33_0;
	wire w_dff_B_4CsqGgUw2_0;
	wire w_dff_B_RuXI1vk84_0;
	wire w_dff_B_R9eycxBg5_0;
	wire w_dff_B_iaVH9DLh4_0;
	wire w_dff_B_W98wexpC1_0;
	wire w_dff_B_7OmBOugY1_0;
	wire w_dff_B_AG6AZ9Nm4_0;
	wire w_dff_B_eMKqIWfC0_0;
	wire w_dff_B_0ymKUaxh0_0;
	wire w_dff_B_7ptmFTMB5_0;
	wire w_dff_B_5WLAdz2G9_0;
	wire w_dff_B_lH9PAfsY7_0;
	wire w_dff_B_iJ9OizwH7_0;
	wire w_dff_B_uHn64dBX9_0;
	wire w_dff_B_FYjWbd0t8_0;
	wire w_dff_B_fk039VRl4_0;
	wire w_dff_B_QN6PEh9G3_0;
	wire w_dff_B_NYGLRl3e2_0;
	wire w_dff_B_M6pBe7jj2_0;
	wire w_dff_B_WUa0vBEc0_0;
	wire w_dff_B_mBJ7qwKY5_0;
	wire w_dff_B_6DBQ2pi99_0;
	wire w_dff_B_8NEJDtKE8_0;
	wire w_dff_B_KnOqWmjK0_0;
	wire w_dff_B_6n7COUYF2_0;
	wire w_dff_B_FI0Lsdpt6_0;
	wire w_dff_B_QWLJXPU56_0;
	wire w_dff_B_vsx1C2pJ4_0;
	wire w_dff_B_8tXB6zb78_0;
	wire w_dff_B_T0nPAzhQ9_0;
	wire w_dff_B_B2i3kMnG5_0;
	wire w_dff_B_dJhWv3XA1_0;
	wire w_dff_B_KxI36ckE7_0;
	wire w_dff_B_s4iz3U4L5_0;
	wire w_dff_B_OZxBQ9Lg8_0;
	wire w_dff_B_sLqxUbDO1_0;
	wire w_dff_B_JZ1ZxhAg2_0;
	wire w_dff_B_OBtaPguL1_0;
	wire w_dff_B_jL7ZsxXN5_0;
	wire w_dff_B_6ig9KpOO3_0;
	wire w_dff_B_bNuv0OMU7_0;
	wire w_dff_B_WTB1Tm6Y4_0;
	wire w_dff_B_qEcBxoGU2_0;
	wire w_dff_B_uMtu1fbb4_0;
	wire w_dff_B_UbU53qU97_0;
	wire w_dff_B_b7uIGOd70_0;
	wire w_dff_B_fek6Kjkc8_0;
	wire w_dff_B_QwJVRI1J7_0;
	wire w_dff_B_OwB2scgS6_0;
	wire w_dff_B_JRmbTlP12_0;
	wire w_dff_B_DgPVVtDQ6_0;
	wire w_dff_B_Nog7bVeE8_0;
	wire w_dff_B_1L36KDnF5_0;
	wire w_dff_B_UpAFjjnA5_0;
	wire w_dff_B_Vn54Je6Y0_0;
	wire w_dff_B_AcNJ84GQ0_0;
	wire w_dff_B_cOzYuYH38_0;
	wire w_dff_B_FkT3Rce07_0;
	wire w_dff_B_09q1r8kV6_0;
	wire w_dff_B_sYCdQLvi8_0;
	wire w_dff_B_GIJFw0J56_0;
	wire w_dff_B_o5ByDST94_0;
	wire w_dff_B_VudLPSsx4_0;
	wire w_dff_B_Zi2pPeuQ7_0;
	wire w_dff_B_aVh0GrHE4_0;
	wire w_dff_B_nrDSOjCU1_0;
	wire w_dff_B_kxMPYsLc4_0;
	wire w_dff_B_u3QFuncY3_0;
	wire w_dff_B_MWhvCoPy3_0;
	wire w_dff_B_CF887ifs5_0;
	wire w_dff_B_3OLCiZsM8_0;
	wire w_dff_B_lu049csJ5_0;
	wire w_dff_B_PDdhCz2h6_0;
	wire w_dff_B_yvif2dZq0_0;
	wire w_dff_B_pZbcdhu90_0;
	wire w_dff_B_1bi4Tpbs2_0;
	wire w_dff_B_3UAlUXRr8_0;
	wire w_dff_B_lCsWWIAI8_0;
	wire w_dff_B_hSBtbjYK6_0;
	wire w_dff_B_CAx6TS4B1_0;
	wire w_dff_B_agazoS5v6_0;
	wire w_dff_B_dd8LGRTQ5_0;
	wire w_dff_B_9vgahaJ52_0;
	wire w_dff_B_TXxQZrVy5_0;
	wire w_dff_B_piQYU72g2_0;
	wire w_dff_B_PzGOo34e2_0;
	wire w_dff_B_qGzKW0d84_0;
	wire w_dff_B_PsTtP93w9_0;
	wire w_dff_B_wR1cEirQ8_0;
	wire w_dff_B_7pacKH3a8_0;
	wire w_dff_B_VY5VH9f41_0;
	wire w_dff_B_GFPnc5QO4_0;
	wire w_dff_B_0Q3FRUhx5_0;
	wire w_dff_B_tOzFoTvX9_0;
	wire w_dff_B_VfmXcYWC8_0;
	wire w_dff_B_UdsshWbY0_0;
	wire w_dff_B_wW5a0vz27_0;
	wire w_dff_B_tUgFNM0R2_0;
	wire w_dff_B_F50xyKXc6_0;
	wire w_dff_B_n9kt1zO44_0;
	wire w_dff_B_gZCxEFbs8_0;
	wire w_dff_B_qXkXsSem1_0;
	wire w_dff_B_AEFnbmRR7_0;
	wire w_dff_B_JMkSfCVw2_0;
	wire w_dff_B_iyPTWEUJ8_0;
	wire w_dff_B_xwHJtFQ73_0;
	wire w_dff_B_T6cy6adT3_0;
	wire w_dff_B_YCOrLBcA4_0;
	wire w_dff_B_8JBrw99v3_0;
	wire w_dff_B_azvmkemw2_0;
	wire w_dff_B_6qGfsBCE4_0;
	wire w_dff_B_k21MNWbT7_0;
	wire w_dff_B_vAXUboMo7_0;
	wire w_dff_B_yZCF1dRt3_0;
	wire w_dff_B_wBhNV9VT5_0;
	wire w_dff_B_Gq2Me05z8_0;
	wire w_dff_B_264E3Ppg9_0;
	wire w_dff_B_XtQtJtAB7_0;
	wire w_dff_B_QJcDwvRC7_0;
	wire w_dff_B_aFaLotrb9_0;
	wire w_dff_B_iKLFWyxf5_0;
	wire w_dff_B_CoH9D9UO9_0;
	wire w_dff_B_O4IoVMVJ8_0;
	wire w_dff_B_iYwXAFHP3_0;
	wire w_dff_B_DIIOGA3I4_0;
	wire w_dff_B_C6YddNUb1_0;
	wire w_dff_B_wDJANGWS5_0;
	wire w_dff_B_NG9S8L2O4_0;
	wire w_dff_B_K5VE6OX58_0;
	wire w_dff_B_uFWTbJsY4_0;
	wire w_dff_B_u5PZETdo0_0;
	wire w_dff_B_n62NxzBo2_0;
	wire w_dff_B_PQuwOxuc2_0;
	wire w_dff_B_aB2r7vXo0_0;
	wire w_dff_B_d9lEHOo34_0;
	wire w_dff_B_eWEJ0pE03_0;
	wire w_dff_B_SRTtuOkb1_0;
	wire w_dff_B_u6Kv1OwD1_0;
	wire w_dff_B_3eRuT4Cj6_0;
	wire w_dff_B_Q7H5VH3Y7_0;
	wire w_dff_B_C04OXU6R4_0;
	wire w_dff_B_aCBPNTXZ4_0;
	wire w_dff_B_syBLDzeQ2_0;
	wire w_dff_B_KdrNcJEW5_0;
	wire w_dff_B_YAiZB8iQ9_0;
	wire w_dff_B_DaitgYX06_0;
	wire w_dff_B_xsNgiLEd8_0;
	wire w_dff_B_qETm5rru0_0;
	wire w_dff_B_BGECBSbQ1_0;
	wire w_dff_B_NYC5UaPH9_0;
	wire w_dff_B_7Wv9h8JE6_0;
	wire w_dff_B_2avyXCgM7_0;
	wire w_dff_B_6TgpZSP71_0;
	wire w_dff_B_urBmP0Nt8_0;
	wire w_dff_B_KEEgq3Bz0_0;
	wire w_dff_B_Bi0EReY61_0;
	wire w_dff_B_juAbyvRb9_0;
	wire w_dff_B_d4AZS7cc9_0;
	wire w_dff_B_jsZ7rHLO3_0;
	wire w_dff_B_whb7k4OF9_0;
	wire w_dff_B_HsobfZOH9_0;
	wire w_dff_B_CxH25B2D8_0;
	wire w_dff_B_z7sBEGJ62_0;
	wire w_dff_B_hiOdseny2_0;
	wire w_dff_B_DZxoEhGy1_0;
	wire w_dff_B_3bixYwa48_0;
	wire w_dff_B_YOIBaXK64_0;
	wire w_dff_B_rSqV4Ts16_0;
	wire w_dff_B_3QdofVOX3_0;
	wire w_dff_B_Vm9xGCX25_0;
	wire w_dff_B_kuRuPFmE9_0;
	wire w_dff_B_k7ztCerr2_0;
	wire w_dff_B_mR9z6GsX2_0;
	wire w_dff_B_2MRfOOKE0_0;
	wire w_dff_B_DtUckFku0_0;
	wire w_dff_B_06xO03r36_0;
	wire w_dff_B_LDcoyRPN9_0;
	wire w_dff_B_ZsBkbrrA7_0;
	wire w_dff_B_6PSJnfqR9_0;
	wire w_dff_B_e1vuhETi1_0;
	wire w_dff_B_22inKnNB2_0;
	wire w_dff_B_1Zjtsvsj7_0;
	wire w_dff_B_2g7v0kq88_0;
	wire w_dff_B_dt23Tw214_0;
	wire w_dff_B_douDrV062_0;
	wire w_dff_B_bJA65jY69_0;
	wire w_dff_B_BocNrqby2_0;
	wire w_dff_B_4rdZMJyE1_0;
	wire w_dff_B_1MDfjnGS8_0;
	wire w_dff_B_19uc25ty4_0;
	wire w_dff_B_2sI8qR5D5_0;
	wire w_dff_B_iW29RgG02_0;
	wire w_dff_B_E0jSOTne1_0;
	wire w_dff_B_b2KFkNXt6_0;
	wire w_dff_B_3Gq8fW909_0;
	wire w_dff_B_3PMSX4V41_0;
	wire w_dff_B_dDmiZuzD1_0;
	wire w_dff_B_lKZf2caW0_0;
	wire w_dff_B_SDlL0hdy8_0;
	wire w_dff_B_e6Ujrzvl3_0;
	wire w_dff_B_FrcdP5mw2_0;
	wire w_dff_B_pDfIcIct4_0;
	wire w_dff_B_qvz13JqE2_0;
	wire w_dff_B_iBqUaBqm5_0;
	wire w_dff_B_DXCiLBRE0_0;
	wire w_dff_B_Iqv9HwlC3_0;
	wire w_dff_B_bD4khmYF5_0;
	wire w_dff_B_5XukiGgD6_0;
	wire w_dff_B_1acq1Ii29_0;
	wire w_dff_B_4xevaueD6_0;
	wire w_dff_B_Hx4PsOQz5_0;
	wire w_dff_B_mIiTho5V0_0;
	wire w_dff_B_P2vsFb309_0;
	wire w_dff_B_LXkLR1Fr3_0;
	wire w_dff_B_sW7lNcSW5_0;
	wire w_dff_B_xHzgBnZg4_0;
	wire w_dff_B_JpTlCLDr0_0;
	wire w_dff_B_9E4Kjc1o2_0;
	wire w_dff_B_qONrkGfY1_0;
	wire w_dff_B_I0TawrUE3_0;
	wire w_dff_B_vDHofyhm0_0;
	wire w_dff_B_c7yZhhEO9_0;
	wire w_dff_B_WuYUn96Y9_0;
	wire w_dff_B_Ol7JlfiZ4_0;
	wire w_dff_B_wSqtQmgq7_0;
	wire w_dff_B_bRCbm9Rl7_0;
	wire w_dff_B_R8zKQYmx3_0;
	wire w_dff_B_9bi76dWM7_0;
	wire w_dff_B_NhSMTdg49_0;
	wire w_dff_B_ETzjzWvT0_0;
	wire w_dff_B_wXohqQjK0_0;
	wire w_dff_B_fNxdkUYc6_0;
	wire w_dff_B_dplX0Cxl5_0;
	wire w_dff_B_TQvxEiMA4_0;
	wire w_dff_B_KL5N6nit9_0;
	wire w_dff_B_wh4smQiZ2_0;
	wire w_dff_B_tfZwkC5h7_0;
	wire w_dff_B_FDkpAuuP3_0;
	wire w_dff_B_CJRtQWYe7_0;
	wire w_dff_B_pDIF9pf89_0;
	wire w_dff_B_oxDHxBc66_0;
	wire w_dff_B_Gq7t7FSN6_0;
	wire w_dff_B_YiUz0Nwb5_0;
	wire w_dff_B_18Xtw7Oy7_0;
	wire w_dff_B_E9kwQgXP9_0;
	wire w_dff_B_RerU6hJo4_0;
	wire w_dff_B_rl6MY5LG7_0;
	wire w_dff_B_QEFc5zrY0_0;
	wire w_dff_B_JEUHMBWj4_0;
	wire w_dff_B_BsBwoum93_0;
	wire w_dff_B_lw6RVVWI9_0;
	wire w_dff_B_cHt50svL9_0;
	wire w_dff_B_1iwoqoe52_0;
	wire w_dff_B_77W1sNdN3_0;
	wire w_dff_B_VK2ZOAJp7_0;
	wire w_dff_B_GLVqlhWB9_0;
	wire w_dff_B_DCvC2j9c7_0;
	wire w_dff_B_bPIzqSKU1_0;
	wire w_dff_B_bkk4KhS27_0;
	wire w_dff_B_MHxfriwQ6_0;
	wire w_dff_B_hwvyEvxS0_0;
	wire w_dff_B_kyP5gtgY7_0;
	wire w_dff_B_HStEtvYq3_0;
	wire w_dff_B_Do2DXFxA7_0;
	wire w_dff_B_XfvIiYZg2_0;
	wire w_dff_B_0oGe2geI1_0;
	wire w_dff_B_qyJML38p0_0;
	wire w_dff_B_CPPLd22G2_0;
	wire w_dff_B_I7DcFExr6_0;
	wire w_dff_B_pQxhO0z48_0;
	wire w_dff_B_o7KTXB8A8_0;
	wire w_dff_B_QSbUKSIM0_0;
	wire w_dff_B_suCkceyA8_0;
	wire w_dff_B_m0wmeRoQ7_0;
	wire w_dff_B_eMtMOVyO5_0;
	wire w_dff_B_oWayQWxz7_0;
	wire w_dff_B_XuEhrRXj2_0;
	wire w_dff_B_P3abaly04_0;
	wire w_dff_B_4oLwDK1c6_0;
	wire w_dff_B_KRMzZgX74_0;
	wire w_dff_B_tKtF7Wnt0_0;
	wire w_dff_B_iaUguIy35_0;
	wire w_dff_B_5vyJka1y5_0;
	wire w_dff_B_SncPSBPK3_0;
	wire w_dff_B_JCIUJa659_0;
	wire w_dff_B_dW1k918b6_0;
	wire w_dff_B_ZCdyyF1Z7_0;
	wire w_dff_B_xUnVWRlw9_0;
	wire w_dff_B_ZmM808xo9_0;
	wire w_dff_B_4Se8GE2H7_0;
	wire w_dff_B_K4evWBVk3_0;
	wire w_dff_B_tGfKGrvW6_0;
	wire w_dff_B_xO6IeWhE7_0;
	wire w_dff_B_hMzYzdHY2_0;
	wire w_dff_B_9CZ7M2z41_0;
	wire w_dff_B_5PSKn6904_0;
	wire w_dff_B_yX6ftvJC7_0;
	wire w_dff_B_oasAignb1_0;
	wire w_dff_B_GJMisELy4_0;
	wire w_dff_B_LPmTurw50_0;
	wire w_dff_B_u6aglghB9_0;
	wire w_dff_B_VjkLqvdk3_0;
	wire w_dff_B_VlXGF5s78_0;
	wire w_dff_B_MHLMp1re6_0;
	wire w_dff_B_d4bCQ6kf9_0;
	wire w_dff_B_RVIQ57f00_0;
	wire w_dff_B_xFHBGtJE6_0;
	wire w_dff_B_JTUR309x7_0;
	wire w_dff_B_P52kOmzq7_0;
	wire w_dff_B_7oXEJaj02_0;
	wire w_dff_B_Dk9FjoTE4_0;
	wire w_dff_B_Et4U5xZw0_0;
	wire w_dff_B_C5dV5OGy2_0;
	wire w_dff_B_RTjt4pGP6_0;
	wire w_dff_B_46EfvZkW0_0;
	wire w_dff_B_BPGfvcvo7_0;
	wire w_dff_B_pIByHgSw4_0;
	wire w_dff_B_NeBzaGqv9_0;
	wire w_dff_B_RM4VGVsv5_0;
	wire w_dff_B_jWLrh7su1_0;
	wire w_dff_B_lo2pgxl81_0;
	wire w_dff_B_A495pgkA5_0;
	wire w_dff_B_VxyDIn9V8_0;
	wire w_dff_B_LU1BuPt49_0;
	wire w_dff_B_fSaz2gyY1_0;
	wire w_dff_B_rNCyxoNw2_0;
	wire w_dff_B_7k4Da50G6_0;
	wire w_dff_B_Xaq2Q8Nu8_0;
	wire w_dff_B_NKYKeJVu9_0;
	wire w_dff_B_hbroTsbw5_0;
	wire w_dff_B_lbstM2MV7_0;
	wire w_dff_B_2RgDHNzc0_0;
	wire w_dff_B_5DCwVdQC5_0;
	wire w_dff_B_mT5R6jG87_0;
	wire w_dff_B_mIhfyMt21_0;
	wire w_dff_B_QtSRwaCV7_0;
	wire w_dff_B_CZ2aD6hQ4_0;
	wire w_dff_B_GFrAB78X7_0;
	wire w_dff_B_lf7v4Nnh0_0;
	wire w_dff_B_tMnsVjYJ7_0;
	wire w_dff_B_p9OIkyt69_0;
	wire w_dff_B_rilLkg6K7_0;
	wire w_dff_B_qVUAyPpR9_0;
	wire w_dff_B_KSsHrZsN1_0;
	wire w_dff_B_k7tcXP4j7_0;
	wire w_dff_B_r9Mik5vs3_0;
	wire w_dff_B_NF5QXmlA3_0;
	wire w_dff_B_jNvoTVNr1_0;
	wire w_dff_B_i0mzmYiS7_0;
	wire w_dff_B_XFSAAHqQ4_0;
	wire w_dff_B_EhXTZVmp6_0;
	wire w_dff_B_eCEc1y8j3_0;
	wire w_dff_B_Gmku2spy9_0;
	wire w_dff_B_puhSnyon2_0;
	wire w_dff_B_zYqCHeFc9_0;
	wire w_dff_B_U8RzyLka3_0;
	wire w_dff_B_7q24LWYe6_0;
	wire w_dff_B_j10PvIAu6_0;
	wire w_dff_B_LycHESkq9_0;
	wire w_dff_B_J4jM6YNu7_0;
	wire w_dff_B_4BdIKe0Y2_0;
	wire w_dff_B_IT84bfga5_0;
	wire w_dff_B_zuwhgRWo6_0;
	wire w_dff_B_tqRdfYdx0_0;
	wire w_dff_B_SZrUMgEJ2_0;
	wire w_dff_B_kLHknRFj5_0;
	wire w_dff_B_04PfymOH4_0;
	wire w_dff_B_Qz3IzuF57_0;
	wire w_dff_B_rXGf7Xad9_0;
	wire w_dff_B_dVHsq43y5_0;
	wire w_dff_B_SA4ZvnlD5_0;
	wire w_dff_B_ZijGJxIu2_0;
	wire w_dff_B_aKc547s88_0;
	wire w_dff_B_yUzHJh7E5_0;
	wire w_dff_B_RTeMNHTZ5_0;
	wire w_dff_B_izNEmQzV3_0;
	wire w_dff_B_DsVZS0sS3_0;
	wire w_dff_B_ZN7c288f0_0;
	wire w_dff_B_SdSoa2yY1_0;
	wire w_dff_B_3uBwT7VQ4_0;
	wire w_dff_B_RCL9xhQg7_0;
	wire w_dff_B_8MrJ8lXq4_0;
	wire w_dff_B_vPkze0ct4_0;
	wire w_dff_B_usXJsdDZ1_0;
	wire w_dff_B_BIxuUcjS6_0;
	wire w_dff_B_3JNl8jYy3_0;
	wire w_dff_B_1pR10h4d4_0;
	wire w_dff_B_yH5iCWGi5_0;
	wire w_dff_B_MudU0od86_0;
	wire w_dff_B_8Tv1xEOP9_0;
	wire w_dff_B_Ic6ZXSpk0_0;
	wire w_dff_B_hXD6z7MN7_0;
	wire w_dff_B_xUfZZOJ30_0;
	wire w_dff_B_LKc93ApG2_0;
	wire w_dff_B_XuRZNCMp8_0;
	wire w_dff_B_vOnBnEEc6_0;
	wire w_dff_B_vBjaB1Kv5_0;
	wire w_dff_B_K8b7Wkp80_0;
	wire w_dff_B_4sGtHFz83_0;
	wire w_dff_B_D3wjCbNs9_0;
	wire w_dff_B_MIEFg4NP4_0;
	wire w_dff_B_VW2R976v3_0;
	wire w_dff_B_e1EDcwHP2_0;
	wire w_dff_B_0DL2AU736_0;
	wire w_dff_B_pGU1PONX9_0;
	wire w_dff_B_7vcrAh8U1_0;
	wire w_dff_B_QYa9mtG04_0;
	wire w_dff_B_0VzXXHas3_0;
	wire w_dff_B_heA6ovfd9_0;
	wire w_dff_B_WGCSYcQp2_0;
	wire w_dff_B_TepX1mJy4_0;
	wire w_dff_B_h8NG1vhQ1_0;
	wire w_dff_B_liZh6P9O6_0;
	wire w_dff_B_t7m5dmNK3_0;
	wire w_dff_B_jY8FVxd07_0;
	wire w_dff_B_ltuIUQgE2_0;
	wire w_dff_B_OijgP3js1_0;
	wire w_dff_B_J9gvKhVz0_0;
	wire w_dff_B_sA4odH6z4_0;
	wire w_dff_B_KKQcqHFT5_0;
	wire w_dff_B_iBJsnuCg0_0;
	wire w_dff_B_nRwV1o3D6_0;
	wire w_dff_B_NE8vMLC30_0;
	wire w_dff_B_jTuWiCzY7_0;
	wire w_dff_B_ruBSvo7p8_0;
	wire w_dff_B_5GLQo37P4_0;
	wire w_dff_B_G4SMXkX32_0;
	wire w_dff_B_Qus7NFco4_0;
	wire w_dff_B_6dujABMS3_0;
	wire w_dff_B_J6S3xhdH7_0;
	wire w_dff_B_Ld0uTr3D8_0;
	wire w_dff_B_8XdTk8ch5_0;
	wire w_dff_B_jfc1YHB47_0;
	wire w_dff_B_6vJjOm7R7_0;
	wire w_dff_B_kzx7Qa7Z2_0;
	wire w_dff_B_QvU9Dc3X3_0;
	wire w_dff_B_6yz624wj1_0;
	wire w_dff_B_zEJtToqs3_0;
	wire w_dff_B_p2OEjJJb5_0;
	wire w_dff_B_pPzyjyLF1_0;
	wire w_dff_B_dvlsUwcj9_0;
	wire w_dff_B_IBM8fJMC1_0;
	wire w_dff_B_irXSsmDw9_0;
	wire w_dff_B_y4jpDxnt1_0;
	wire w_dff_B_WrHyyegD7_0;
	wire w_dff_B_FAYirqBa0_0;
	wire w_dff_B_3eMcAsGG5_0;
	wire w_dff_B_t66iQooO7_0;
	wire w_dff_B_OgbsSv5y6_0;
	wire w_dff_B_bj17yU8k5_0;
	wire w_dff_B_DOU5GeaM0_0;
	wire w_dff_B_QJPgP2Ii8_0;
	wire w_dff_B_dvTrZ2uC7_0;
	wire w_dff_B_1J0CQA1T1_0;
	wire w_dff_B_O5pd8KNF2_0;
	wire w_dff_B_xKyJSnvx9_0;
	wire w_dff_B_xUxwdEOO4_0;
	wire w_dff_B_WvWxvWzg8_0;
	wire w_dff_B_4JurAnWO1_0;
	wire w_dff_B_1PywuMYM8_0;
	wire w_dff_B_qQK6xdmP0_0;
	wire w_dff_B_yHbwg9zI7_0;
	wire w_dff_B_e35l5UNQ1_0;
	wire w_dff_B_cdkBYG2h0_0;
	wire w_dff_B_IG7pST6V5_0;
	wire w_dff_B_EPH60IHt3_0;
	wire w_dff_B_l5qyYNxV1_0;
	wire w_dff_B_IAiQbhVG9_0;
	wire w_dff_B_fnq00r5f8_0;
	wire w_dff_B_hAq0AFvq7_0;
	wire w_dff_B_rwtN9Dwa0_0;
	wire w_dff_B_e8jJu26v3_0;
	wire w_dff_B_eHsvm46h3_0;
	wire w_dff_B_TtgmAGTn0_0;
	wire w_dff_B_4EMNny3E5_0;
	wire w_dff_B_u2LK2WNV2_0;
	wire w_dff_B_BfiVhUQz3_0;
	wire w_dff_B_7KHaRl9h8_0;
	wire w_dff_B_4ZgDo9038_0;
	wire w_dff_B_7vLfPSF12_0;
	wire w_dff_B_qwfiJ8jA7_0;
	wire w_dff_B_Gn6RKfnD8_0;
	wire w_dff_B_VoKB9te33_0;
	wire w_dff_B_i5Ln6cRk3_0;
	wire w_dff_B_dRIK55IK4_0;
	wire w_dff_B_yHwN6seX7_0;
	wire w_dff_B_1hYcPsh28_0;
	wire w_dff_B_iQdA0oYB7_0;
	wire w_dff_B_ONiY33U54_0;
	wire w_dff_B_SsvILKT16_0;
	wire w_dff_B_DPy1PlS17_0;
	wire w_dff_B_dQL4cCvp1_0;
	wire w_dff_B_zHY7OdU13_0;
	wire w_dff_B_EpjFEFeS6_0;
	wire w_dff_B_M9AbqevZ7_0;
	wire w_dff_B_N3uT70rS9_0;
	wire w_dff_B_Kzc4vf1Y8_0;
	wire w_dff_B_qeU1Jg9J3_0;
	wire w_dff_B_YxVz6JQl8_0;
	wire w_dff_B_FoBnzwng2_0;
	wire w_dff_B_ydFqt54R5_0;
	wire w_dff_B_0Yk60AUn4_0;
	wire w_dff_B_KWjZkP2Z7_0;
	wire w_dff_B_jaK0c1Xn0_0;
	wire w_dff_B_7EiIuLxG6_0;
	wire w_dff_B_yzxG5pAF8_0;
	wire w_dff_B_m2cDGtgO7_0;
	wire w_dff_B_KXAHi7d68_0;
	wire w_dff_B_OwyZ7XQu4_0;
	wire w_dff_B_8nhSkh2d0_0;
	wire w_dff_B_doTWgxu09_0;
	wire w_dff_B_DfJVRy199_0;
	wire w_dff_B_YryYg53B0_0;
	wire w_dff_B_tDNBPcBN1_0;
	wire w_dff_B_VYbjiQVo0_0;
	wire w_dff_B_SvvQIaor6_0;
	wire w_dff_B_Mbm0k7Ty0_0;
	wire w_dff_B_KNGBHHix8_0;
	wire w_dff_B_liyVAZm50_0;
	wire w_dff_B_tmovH3rI1_0;
	wire w_dff_B_vLltUVYY5_0;
	wire w_dff_B_AKb6EvBO0_0;
	wire w_dff_B_OCrwxUvx1_0;
	wire w_dff_B_w7pQ7NKj8_0;
	wire w_dff_B_k1aDtxx55_0;
	wire w_dff_B_NtITRMw89_0;
	wire w_dff_B_RvtWyrLH0_0;
	wire w_dff_B_9vinJAyS7_0;
	wire w_dff_B_hbD1bP0Y2_0;
	wire w_dff_B_KOeHJObt7_0;
	wire w_dff_B_ZlvCaaZo4_0;
	wire w_dff_B_aLUVpM9m6_0;
	wire w_dff_B_UwlWFzeN5_0;
	wire w_dff_B_UEFFLVhB1_0;
	wire w_dff_B_0LkHLgGP3_0;
	wire w_dff_B_G9OQg0hk8_0;
	wire w_dff_B_fZJ5prOr5_0;
	wire w_dff_B_MGTlem011_0;
	wire w_dff_B_P2bGgnOC2_0;
	wire w_dff_B_gKKZ7ijG5_0;
	wire w_dff_B_GZS0JPIc8_0;
	wire w_dff_B_BfDKFQb51_0;
	wire w_dff_B_TiIBP8De2_0;
	wire w_dff_B_ahi47YUR1_0;
	wire w_dff_B_2L9c7xNO9_0;
	wire w_dff_B_cirpKDKK6_0;
	wire w_dff_B_YTaqmtxP4_0;
	wire w_dff_B_pbCKghN20_0;
	wire w_dff_B_5ypTpoPi5_0;
	wire w_dff_B_z4G8Pj2d1_0;
	wire w_dff_B_jCrwUYlh1_0;
	wire w_dff_B_3jsugFd75_0;
	wire w_dff_B_h3kS9t0a5_0;
	wire w_dff_B_ZQaquU432_0;
	wire w_dff_B_LtIRXA7N4_0;
	wire w_dff_B_zsf56dpY7_0;
	wire w_dff_B_I6JZrKXq3_0;
	wire w_dff_B_euQRbziA8_0;
	wire w_dff_B_mGH4Jypu5_0;
	wire w_dff_B_4iPpF1Tk3_0;
	wire w_dff_B_mlscRo030_0;
	wire w_dff_B_ZTDC1JDE7_0;
	wire w_dff_B_TERbME9F8_0;
	wire w_dff_B_Y58xZaMx0_0;
	wire w_dff_B_U0SaqLbB5_0;
	wire w_dff_B_nlS8FHBj7_0;
	wire w_dff_B_6jrtoveD4_0;
	wire w_dff_B_nrJpjEzB0_0;
	wire w_dff_B_VCHSalno5_0;
	wire w_dff_B_sw1P9WON5_0;
	wire w_dff_B_mqJ7AQMa2_0;
	wire w_dff_B_0Eyj2soR8_0;
	wire w_dff_B_x8wOIjQS5_0;
	wire w_dff_B_T1tXy2XH0_0;
	wire w_dff_B_NQAJivaY7_0;
	wire w_dff_B_Hbnqvyz66_0;
	wire w_dff_B_wd0ZXQVw3_0;
	wire w_dff_B_yKICTire7_0;
	wire w_dff_B_YNYFKqvT1_0;
	wire w_dff_B_pzm6NvQh4_0;
	wire w_dff_B_yi97ZAmR0_0;
	wire w_dff_B_NysdbI4B7_0;
	wire w_dff_B_Z8oEXEOq5_0;
	wire w_dff_B_PrvvhIbo1_0;
	wire w_dff_B_0oklccaG4_0;
	wire w_dff_B_uiSXcZUB4_0;
	wire w_dff_B_mDeIGuJ43_0;
	wire w_dff_B_bPjvRbd34_0;
	wire w_dff_B_ENEpxAde1_0;
	wire w_dff_B_YYh6OEfL0_0;
	wire w_dff_B_m2uiIz561_0;
	wire w_dff_B_kNSsNfC44_0;
	wire w_dff_B_LiqLZPqr6_0;
	wire w_dff_B_17rldnQW9_0;
	wire w_dff_B_whrCssj15_0;
	wire w_dff_B_7HpG867R3_0;
	wire w_dff_B_3qU7Pgnd1_0;
	wire w_dff_B_VasuzH687_0;
	wire w_dff_B_jTSAjFIp4_0;
	wire w_dff_B_szxPUmwE9_0;
	wire w_dff_B_wILe7lwQ1_0;
	wire w_dff_B_jxkLKYS50_0;
	wire w_dff_B_FDORIHlv4_0;
	wire w_dff_B_aAOVCfFw2_0;
	wire w_dff_B_xzNnsrPZ7_0;
	wire w_dff_B_DvZpfQh54_0;
	wire w_dff_B_81zvE9Ef0_0;
	wire w_dff_B_bNJMmZSS0_0;
	wire w_dff_B_WEjQ75Xz2_0;
	wire w_dff_B_od168AOs0_0;
	wire w_dff_B_hkNZmOeF6_0;
	wire w_dff_B_0HABUdRj6_0;
	wire w_dff_B_1Ox4RIbi2_0;
	wire w_dff_B_urGQZy9D3_0;
	wire w_dff_B_Et0Ae4xm4_0;
	wire w_dff_B_eNc3Quge2_0;
	wire w_dff_B_nRcI7H9Q4_0;
	wire w_dff_B_kJjiz5uG4_0;
	wire w_dff_B_u2z4JjPk5_0;
	wire w_dff_B_aUXWCfaT5_0;
	wire w_dff_B_vSmmTJWj6_0;
	wire w_dff_B_4GQKI0Wq5_0;
	wire w_dff_B_l749LOFF5_0;
	wire w_dff_B_aRd4vaSr9_0;
	wire w_dff_B_vPSmcQff2_0;
	wire w_dff_B_kNchVSOD4_0;
	wire w_dff_B_qYjdLf3P0_0;
	wire w_dff_B_F0FQD6cg9_0;
	wire w_dff_B_hJIGDIrz4_0;
	wire w_dff_B_AR2FvIXN8_0;
	wire w_dff_B_d50zOTAp5_0;
	wire w_dff_B_k7v2pxiZ3_0;
	wire w_dff_B_lRwxMITQ8_0;
	wire w_dff_B_zex4fiO20_0;
	wire w_dff_B_97cjC2gG3_0;
	wire w_dff_B_ubt9NPi78_0;
	wire w_dff_B_Y2DU5Z5c3_0;
	wire w_dff_B_VULUXgp86_0;
	wire w_dff_B_Hg2syQxk9_0;
	wire w_dff_B_JB3M4uWh1_0;
	wire w_dff_B_aBle1NC62_0;
	wire w_dff_B_zM0TcW941_0;
	wire w_dff_B_n0oxOqpK1_0;
	wire w_dff_B_N8XFtalI6_0;
	wire w_dff_B_OaRocCCV1_0;
	wire w_dff_B_Bha0PZ8T5_0;
	wire w_dff_B_bdyIpRd64_0;
	wire w_dff_B_PayoqlsK8_0;
	wire w_dff_B_cJe2QCEx9_0;
	wire w_dff_B_OvBXG0gx8_0;
	wire w_dff_B_Dls3IOzT3_0;
	wire w_dff_B_gRUP5ac66_0;
	wire w_dff_B_JWa0fYzz7_0;
	wire w_dff_B_gfnlPPgT8_0;
	wire w_dff_B_X5fasANi6_0;
	wire w_dff_B_gELEVP791_0;
	wire w_dff_B_4FyXF39X4_0;
	wire w_dff_B_JzUETrMd5_0;
	wire w_dff_B_ZMSgl2eg8_0;
	wire w_dff_B_arvvqOuV6_0;
	wire w_dff_B_IJFnLUlT7_0;
	wire w_dff_B_OZzL7Krh5_0;
	wire w_dff_B_j68Ib33U5_0;
	wire w_dff_B_6zFH5uQN4_0;
	wire w_dff_B_hQxUX1WK5_0;
	wire w_dff_B_8itDHIDq3_0;
	wire w_dff_B_oIn76kGK6_0;
	wire w_dff_B_xRqNo4PA0_0;
	wire w_dff_B_UgChdVzk8_0;
	wire w_dff_B_enyuX2n99_0;
	wire w_dff_B_weeMWlHm2_0;
	wire w_dff_B_Cp0yVbP13_0;
	wire w_dff_B_SBebaV8n2_0;
	wire w_dff_B_oqHghBrO3_0;
	wire w_dff_B_F0e8169s2_0;
	wire w_dff_B_csu2yVde3_0;
	wire w_dff_B_Z7PCXxEK1_0;
	wire w_dff_B_XMyPOCWG6_0;
	wire w_dff_B_VlgJaTYI1_0;
	wire w_dff_B_rWJ1jfPs7_0;
	wire w_dff_B_M7vRvPIA2_0;
	wire w_dff_B_H52zktDU8_0;
	wire w_dff_B_jXczRxPA9_0;
	wire w_dff_B_qUOG4h1x1_0;
	wire w_dff_B_o2BsuHd70_0;
	wire w_dff_B_Uy391QM83_0;
	wire w_dff_B_yWsdAQQN4_0;
	wire w_dff_B_hSS5iuJ31_0;
	wire w_dff_B_QRoVHLTH5_0;
	wire w_dff_B_asFz572A4_0;
	wire w_dff_B_Q17GLZcN7_0;
	wire w_dff_B_enQSSbSI4_0;
	wire w_dff_B_7HO00lui4_0;
	wire w_dff_B_GRsMJyys5_0;
	wire w_dff_B_oYeez4Mp4_0;
	wire w_dff_B_OCCOYnUR6_0;
	wire w_dff_B_XykJq9xE8_0;
	wire w_dff_B_pSQIn4d31_0;
	wire w_dff_B_mrE4b4hj0_0;
	wire w_dff_B_FEC12HEQ4_0;
	wire w_dff_B_UkKKrox99_0;
	wire w_dff_B_rBIY3iHI6_0;
	wire w_dff_B_akrvIWaH5_0;
	wire w_dff_B_axc63lYQ5_0;
	wire w_dff_B_jgXX1eQ82_0;
	wire w_dff_B_PcGZrH3T8_0;
	wire w_dff_B_f3795ANB1_0;
	wire w_dff_B_FvBLlsaI2_0;
	wire w_dff_B_eAwVNVwG9_0;
	wire w_dff_B_ziZwOSYL3_0;
	wire w_dff_B_yPdosjHg9_0;
	wire w_dff_B_wymPk2af8_0;
	wire w_dff_B_R0WSs6Kl2_0;
	wire w_dff_B_pvkvl9fo4_0;
	wire w_dff_B_aitfsw0Y0_0;
	wire w_dff_B_7g7gUE3u9_0;
	wire w_dff_B_tPg7xZrw4_0;
	wire w_dff_B_iBS0wxeZ6_0;
	wire w_dff_B_jjVcmA4s4_0;
	wire w_dff_B_WQjdV6h15_0;
	wire w_dff_B_CZLR0oVD8_0;
	wire w_dff_B_OySqiWIz0_0;
	wire w_dff_B_LEjgoI5o0_0;
	wire w_dff_B_4WD5y66k1_0;
	wire w_dff_B_skvqbat10_0;
	wire w_dff_B_058xrlB73_0;
	wire w_dff_B_C1xAoHo36_0;
	wire w_dff_B_SP7zVPQj4_0;
	wire w_dff_B_eIXA1Ojg3_0;
	wire w_dff_B_VZFoyD096_0;
	wire w_dff_B_UXRrNooA3_0;
	wire w_dff_B_mx6QzdhE8_0;
	wire w_dff_B_lo3ftZGt8_0;
	wire w_dff_B_wJjz88Px4_0;
	wire w_dff_B_RcaFbYO23_0;
	wire w_dff_B_2dC1oWKF0_0;
	wire w_dff_B_9Syh3jcY8_0;
	wire w_dff_B_RGCJIKH71_0;
	wire w_dff_B_Ysl7iKtY3_0;
	wire w_dff_B_6dFmWfct1_0;
	wire w_dff_B_Ctcu9det7_0;
	wire w_dff_B_rdyuhxwe7_0;
	wire w_dff_B_o6lmB5kz9_0;
	wire w_dff_B_7igJX8uc5_0;
	wire w_dff_B_J1cj6hri7_0;
	wire w_dff_B_vqBhSY1U0_0;
	wire w_dff_B_2pDodbty5_0;
	wire w_dff_B_r6L3mB699_0;
	wire w_dff_B_hUioI3XI0_0;
	wire w_dff_B_h7a50YUe6_0;
	wire w_dff_B_R39OpCJ14_0;
	wire w_dff_B_R1MBCPqW0_0;
	wire w_dff_B_ayKbiZxB8_0;
	wire w_dff_B_mI9qiqLD3_0;
	wire w_dff_B_XQ5VNEIN0_0;
	wire w_dff_B_olB7Nf1l5_0;
	wire w_dff_B_Z8bPN8lA7_0;
	wire w_dff_B_a4ImkX0F1_0;
	wire w_dff_B_lDMaNvAY8_0;
	wire w_dff_B_PPVk8cTU1_0;
	wire w_dff_B_f06G2IVk1_0;
	wire w_dff_B_4G0r33FD6_0;
	wire w_dff_B_Uo9sTI2d6_0;
	wire w_dff_B_ceXLxFiL2_0;
	wire w_dff_B_3McNI1BL0_0;
	wire w_dff_B_zDAuNtQN3_0;
	wire w_dff_B_YzTcwtiy2_0;
	wire w_dff_B_JGsJ6wVA3_0;
	wire w_dff_B_8Y8lLYyy9_0;
	wire w_dff_B_D5b77H9w0_0;
	wire w_dff_B_1B8zarzA9_0;
	wire w_dff_B_TEwD6oFa2_0;
	wire w_dff_B_uBe9ALIw3_0;
	wire w_dff_B_g89ZXUxF9_0;
	wire w_dff_B_HQ3uB9VM1_0;
	wire w_dff_B_mtJwnctp2_0;
	wire w_dff_B_aCmArjJb1_0;
	wire w_dff_B_sQImK0oE6_0;
	wire w_dff_B_yvHaVn4I2_0;
	wire w_dff_B_2adiK2LN7_0;
	wire w_dff_B_pTGyYuFZ4_0;
	wire w_dff_B_7LYmdE161_0;
	wire w_dff_B_gH0gpuAR2_0;
	wire w_dff_B_5l3KvKCB6_0;
	wire w_dff_B_ONbJNmru1_0;
	wire w_dff_B_8YOxLtd12_0;
	wire w_dff_B_bda9rMd55_0;
	wire w_dff_B_zBiJ20cc7_0;
	wire w_dff_B_yw4Ht0p46_0;
	wire w_dff_B_QKXuQfY94_0;
	wire w_dff_B_xkcW9Ldj2_0;
	wire w_dff_B_YSC6YNxi9_0;
	wire w_dff_B_ht3ZNn0X2_0;
	wire w_dff_B_2y13gvOT4_0;
	wire w_dff_B_WHfWUouE0_0;
	wire w_dff_B_VaxtxZZ68_0;
	wire w_dff_B_8kTQRZpM2_0;
	wire w_dff_B_sLqCAoEz9_0;
	wire w_dff_B_f5k0RJ456_0;
	wire w_dff_B_uvwQYYe33_0;
	wire w_dff_B_PRHQDVjY9_0;
	wire w_dff_B_NfGs6jPv4_0;
	wire w_dff_B_br24ce4R8_0;
	wire w_dff_B_PfkViLOG8_0;
	wire w_dff_B_M3EDA1xX7_0;
	wire w_dff_B_Dv7mLFTF0_0;
	wire w_dff_B_lWCsIlXA3_0;
	wire w_dff_B_b6Ptx8On0_0;
	wire w_dff_B_JqoYJHNx4_0;
	wire w_dff_B_QUgVbbHD2_0;
	wire w_dff_B_tAlzt0PE9_0;
	wire w_dff_B_zFlF74da1_0;
	wire w_dff_B_KfmETYUc9_0;
	wire w_dff_B_h9TbfxFo9_0;
	wire w_dff_B_8yg7ndMK2_0;
	wire w_dff_B_3MpH5j2X5_0;
	wire w_dff_B_EWl41ZHf9_0;
	wire w_dff_B_XInmM5uu3_0;
	wire w_dff_B_dIrbEeRa3_0;
	wire w_dff_B_gBbA07bB9_0;
	wire w_dff_B_pghgJ4ba8_0;
	wire w_dff_B_Q37UsApI4_0;
	wire w_dff_B_yQhmpA628_0;
	wire w_dff_B_viVkT27L6_0;
	wire w_dff_B_XxWJ1Jxq1_0;
	wire w_dff_B_qJ6EI6jf5_0;
	wire w_dff_B_OrBgQSXt0_0;
	wire w_dff_B_949NfNXB3_0;
	wire w_dff_B_EZeSEKlo9_0;
	wire w_dff_B_RkqjMSOq9_0;
	wire w_dff_B_Mh3FBitm2_0;
	wire w_dff_B_Na2H7pV40_0;
	wire w_dff_B_YtrVJamn6_0;
	wire w_dff_B_YYP0CtYA1_0;
	wire w_dff_B_d6p7MoRg9_0;
	wire w_dff_B_8kAJQYO34_0;
	wire w_dff_B_qH5oY8uJ3_0;
	wire w_dff_B_D5Uc1jHX5_0;
	wire w_dff_B_oFWzUzBP3_0;
	wire w_dff_B_xqY3nI2K4_0;
	wire w_dff_B_OdI2Kmp07_0;
	wire w_dff_B_hjy5hvL31_0;
	wire w_dff_B_tO9ZQHds9_0;
	wire w_dff_B_XQ6nkice2_0;
	wire w_dff_B_255O0Gm10_0;
	wire w_dff_B_xkVcMmOa7_0;
	wire w_dff_B_3AGfhD7j7_0;
	wire w_dff_B_iAB8pE324_0;
	wire w_dff_B_0R0K3Tct8_0;
	wire w_dff_B_myEnWWZf3_0;
	wire w_dff_B_ALKRB9Qx1_0;
	wire w_dff_B_w5qCJn1V6_0;
	wire w_dff_B_4vYjZtvV4_0;
	wire w_dff_B_JW8XbCeJ8_0;
	wire w_dff_B_1NVcs1eF0_0;
	wire w_dff_B_XpuqO2R07_0;
	wire w_dff_B_9YuaLM9C6_0;
	wire w_dff_B_MXoq1Ttp7_0;
	wire w_dff_B_qGiSvxQb7_0;
	wire w_dff_B_ENTmt6wu3_0;
	wire w_dff_B_LEA0bSTb9_0;
	wire w_dff_B_hy3o6oGJ7_0;
	wire w_dff_B_bOmHALdH6_0;
	wire w_dff_B_lEZK15qY6_0;
	wire w_dff_B_qSxc1DSk1_0;
	wire w_dff_B_ctoUowCc3_0;
	wire w_dff_B_m3x6gj4X9_0;
	wire w_dff_B_Uo2YVoss8_0;
	wire w_dff_B_GjpHOfA39_0;
	wire w_dff_B_XejYHmwb3_0;
	wire w_dff_B_q3JTuYo19_0;
	wire w_dff_B_3NMrET7T2_0;
	wire w_dff_B_Q3ZifXet2_0;
	wire w_dff_B_zd7nAWJf9_0;
	wire w_dff_B_B7UsuSFP8_0;
	wire w_dff_B_xds5KlN45_0;
	wire w_dff_B_Xk0JZCvB8_0;
	wire w_dff_B_J7YFGtA00_0;
	wire w_dff_B_bv29g9Jy1_0;
	wire w_dff_B_lZGlEFem2_0;
	wire w_dff_B_FQSNxKtS7_0;
	wire w_dff_B_Hvq6Grez2_0;
	wire w_dff_B_TcFL9nsw1_0;
	wire w_dff_B_xRZ7eL2I9_0;
	wire w_dff_B_4uVeLXgT1_0;
	wire w_dff_B_S1hPxKk54_0;
	wire w_dff_B_pQEcvPJv2_0;
	wire w_dff_B_NHJIqKwT4_0;
	wire w_dff_B_64vqJbq99_0;
	wire w_dff_B_zcyh6tyj7_0;
	wire w_dff_B_OGYbucAE2_0;
	wire w_dff_B_5soQjnSu7_0;
	wire w_dff_B_Tfb2awxR8_0;
	wire w_dff_B_QW5uwTx62_0;
	wire w_dff_B_J79DAcIc8_0;
	wire w_dff_B_sYWKG7EC6_0;
	wire w_dff_B_VQvPcADU8_0;
	wire w_dff_B_AL82UpN57_0;
	wire w_dff_B_ZdleOjl17_0;
	wire w_dff_B_1R7ICl8B5_0;
	wire w_dff_B_6j3JQ2Ye1_0;
	wire w_dff_B_GwRlqcdt9_0;
	wire w_dff_B_aFU78AoU4_0;
	wire w_dff_B_k7Sv53oC8_0;
	wire w_dff_B_zNXCch063_0;
	wire w_dff_B_06188mbO7_0;
	wire w_dff_B_0T21YHHZ5_0;
	wire w_dff_B_4MTCsF4h5_0;
	wire w_dff_B_Z2ZYBYoe5_0;
	wire w_dff_B_9NJc5g0k8_0;
	wire w_dff_B_tsUyjEzS5_0;
	wire w_dff_B_dRJvOagH5_0;
	wire w_dff_B_X1ffWE3Q5_0;
	wire w_dff_B_rTAMs7736_0;
	wire w_dff_B_m05ehC0M4_0;
	wire w_dff_B_R0ah8XUb0_0;
	wire w_dff_B_R9A4UXxW7_0;
	wire w_dff_B_EPxWfQPV7_0;
	wire w_dff_B_Mf4bGIIs7_0;
	wire w_dff_B_QaQNlswz9_0;
	wire w_dff_B_EuzV3vtZ1_0;
	wire w_dff_B_QNasHvvk5_0;
	wire w_dff_B_y4hAOaeC8_0;
	wire w_dff_B_DW7Hd0zZ4_0;
	wire w_dff_B_pEIU1tti0_0;
	wire w_dff_B_ansSb8I39_0;
	wire w_dff_B_fAjzcvNj6_0;
	wire w_dff_B_QLIZezVG4_0;
	wire w_dff_B_Qg9q82gk7_0;
	wire w_dff_B_dRcAfLlT1_0;
	wire w_dff_B_03kc00be7_0;
	wire w_dff_B_tTmkozGb2_0;
	wire w_dff_B_mvqwZPIt5_0;
	wire w_dff_B_fsFWWfRn4_0;
	wire w_dff_B_ryLtxjvR4_0;
	wire w_dff_B_Zi7Kn8s95_0;
	wire w_dff_B_ewEgondB9_0;
	wire w_dff_B_s8fARmAD6_0;
	wire w_dff_B_eeDG3VW25_0;
	wire w_dff_B_DxlMODMl8_0;
	wire w_dff_B_ZaOHtoZ17_0;
	wire w_dff_B_f7st35aB7_0;
	wire w_dff_B_gX65ix2R6_0;
	wire w_dff_B_XaPkAPXA9_0;
	wire w_dff_B_YvAd3XN95_0;
	wire w_dff_B_If53B8Lr3_0;
	wire w_dff_B_3qhl4UMJ7_0;
	wire w_dff_B_FjrUDAfU4_0;
	wire w_dff_B_99w7Z6TT5_0;
	wire w_dff_B_gGSxsUmt7_0;
	wire w_dff_B_oHLn4Y4u5_0;
	wire w_dff_B_m1lKuX0E8_0;
	wire w_dff_B_FoVXwOim6_0;
	wire w_dff_B_Ci8weqxh9_0;
	wire w_dff_B_dvfqsnxx7_0;
	wire w_dff_B_uaufbcCs8_0;
	wire w_dff_B_VwnMBN5V0_0;
	wire w_dff_B_PAFSZUxB2_0;
	wire w_dff_B_fTJkyqac6_0;
	wire w_dff_B_Z5KanTJ08_0;
	wire w_dff_B_sumWS9Vf1_0;
	wire w_dff_B_Hs5hme0D4_0;
	wire w_dff_B_aUHOxU028_0;
	wire w_dff_B_bDPtbaLa9_0;
	wire w_dff_B_LWzBJ1wn8_0;
	wire w_dff_B_K9EmdHoN5_0;
	wire w_dff_B_VUr17GFe9_0;
	wire w_dff_B_Am7rY1bk0_0;
	wire w_dff_B_U4RWagem4_0;
	wire w_dff_B_xMv1cFCZ6_0;
	wire w_dff_B_iJ80qHxz8_0;
	wire w_dff_B_ZyQYSZ7M0_0;
	wire w_dff_B_vqi0rSWK0_0;
	wire w_dff_B_JNlauO5R2_0;
	wire w_dff_B_q8wKsiWr7_0;
	wire w_dff_B_BT95v4uZ1_0;
	wire w_dff_B_zUs7LGxC3_0;
	wire w_dff_B_dERnxNsj3_0;
	wire w_dff_B_5xRsFM2h0_0;
	wire w_dff_B_SVtCOT2J2_0;
	wire w_dff_B_HZqNBcJf9_0;
	wire w_dff_B_Pf0M2pUw5_0;
	wire w_dff_B_oft0TmF22_0;
	wire w_dff_B_MeInrIck5_0;
	wire w_dff_B_D7IZ15Xj8_0;
	wire w_dff_B_lex8LvAY0_0;
	wire w_dff_B_0EacPJrC4_0;
	wire w_dff_B_K6gDg8ps6_0;
	wire w_dff_B_R6jgogip4_0;
	wire w_dff_B_UxC2HckD4_0;
	wire w_dff_B_tTc713Uj8_0;
	wire w_dff_B_oRHtQbeD3_0;
	wire w_dff_B_9xMQN7mS8_0;
	wire w_dff_B_ywF9zxmX0_0;
	wire w_dff_B_b2mL7x6g3_0;
	wire w_dff_B_QA871eee6_0;
	wire w_dff_B_pyQmjL5f4_0;
	wire w_dff_B_Kz5OZ4SS3_0;
	wire w_dff_B_GX8upgfY9_0;
	wire w_dff_B_7KiseVrI1_0;
	wire w_dff_B_USkwMxb58_0;
	wire w_dff_B_1PbrWO2m0_0;
	wire w_dff_B_YL5KE44k3_0;
	wire w_dff_B_jr9TK7yz0_0;
	wire w_dff_B_YE7lnPud9_0;
	wire w_dff_B_6SYbh95w9_0;
	wire w_dff_B_BZZufOtI5_0;
	wire w_dff_B_yqvkyrSA5_0;
	wire w_dff_B_SsVTULxg1_0;
	wire w_dff_B_tWhdsU6j2_0;
	wire w_dff_B_ZMiI4tSI8_0;
	wire w_dff_B_28DVf9vj6_0;
	wire w_dff_B_WEwKMJx30_0;
	wire w_dff_B_EpwZydaA5_0;
	wire w_dff_B_eYXoIjyu2_0;
	wire w_dff_B_jrLI29pl5_0;
	wire w_dff_B_JG8DkIUd7_0;
	wire w_dff_B_OxKsOoDk2_0;
	wire w_dff_B_gSM54LjO2_0;
	wire w_dff_B_DW3JjsXk5_0;
	wire w_dff_B_bMYepiXd0_0;
	wire w_dff_B_RxDlKpGR1_0;
	wire w_dff_B_jgeBD7LJ0_0;
	wire w_dff_B_lSnu0hEj7_0;
	wire w_dff_B_voGnUNqX6_0;
	wire w_dff_B_RiP2rXi55_0;
	wire w_dff_B_Xj5IwNDZ3_0;
	wire w_dff_B_DreSfcaI6_0;
	wire w_dff_B_sKqGZVVb5_0;
	wire w_dff_B_c9qoYoWt5_0;
	wire w_dff_B_45FinX8J8_0;
	wire w_dff_B_QXacbdg74_0;
	wire w_dff_B_UhqzJBa99_0;
	wire w_dff_B_Ize3D40m1_0;
	wire w_dff_B_ddhj3QHk2_0;
	wire w_dff_B_8W09mOKq3_0;
	wire w_dff_B_em62HQD64_0;
	wire w_dff_B_qhYwhaxn2_0;
	wire w_dff_B_MI6HC4ki4_0;
	wire w_dff_B_hCdq7GtP3_0;
	wire w_dff_B_XsNGDlmV1_0;
	wire w_dff_B_yKkBc2z46_0;
	wire w_dff_B_snxZhQFr4_0;
	wire w_dff_B_8ObNGCI84_0;
	wire w_dff_B_HG9Vk3OM7_0;
	wire w_dff_B_r0rT2Is62_0;
	wire w_dff_B_5PrLCwF72_0;
	wire w_dff_B_lU5TZhx31_0;
	wire w_dff_B_gIvtSsaY3_0;
	wire w_dff_B_Io6IhENr2_0;
	wire w_dff_B_j2B6MhCB5_0;
	wire w_dff_B_1YfhAhGF9_0;
	wire w_dff_B_VGPns6hT5_0;
	wire w_dff_B_sW6nfMfl4_0;
	wire w_dff_B_dUGc9UGL1_0;
	wire w_dff_B_ssziijg54_0;
	wire w_dff_B_qBqDYGex6_0;
	wire w_dff_B_bvcHLzuZ9_0;
	wire w_dff_B_BdjdFfqJ5_0;
	wire w_dff_B_Lcy99c6n0_0;
	wire w_dff_B_8T58l3zu0_0;
	wire w_dff_B_MKoIYWEN1_0;
	wire w_dff_B_sFYOgUgD2_0;
	wire w_dff_B_iqj7Ez2z2_0;
	wire w_dff_B_1VTFtqw26_0;
	wire w_dff_B_QFCS8o9h9_0;
	wire w_dff_B_qCbSgFBQ9_0;
	wire w_dff_B_NCSjtdzZ5_0;
	wire w_dff_B_t0LAegjI5_0;
	wire w_dff_B_lGbTRTlI6_0;
	wire w_dff_B_2Mau76xd5_0;
	wire w_dff_B_ZYiFP1Iv4_0;
	wire w_dff_B_ESvanhO48_0;
	wire w_dff_B_mStUFvyr1_0;
	wire w_dff_B_qjSeEygS7_0;
	wire w_dff_B_NvsNP2829_0;
	wire w_dff_B_VDy8bCyP8_0;
	wire w_dff_B_o1pTnOrf9_0;
	wire w_dff_B_AOv7yzLK2_0;
	wire w_dff_B_UjFyqUbx8_0;
	wire w_dff_B_dZRukDxF5_0;
	wire w_dff_B_GfOiaw6Q0_0;
	wire w_dff_B_85W6pltF8_0;
	wire w_dff_B_c6d7m3HU2_0;
	wire w_dff_B_uZzhl7WP6_0;
	wire w_dff_B_NWbI1MMV8_0;
	wire w_dff_B_UEfEi3w39_0;
	wire w_dff_B_wiPKtVAr4_0;
	wire w_dff_B_DzQbWtaQ8_0;
	wire w_dff_B_U0D9RSqn3_0;
	wire w_dff_B_5Pb8sBBf1_0;
	wire w_dff_B_CovSE80Y8_0;
	wire w_dff_B_1Zq4LUxj6_0;
	wire w_dff_B_ISTrKf4C6_0;
	wire w_dff_B_JDhcM3W96_0;
	wire w_dff_B_sQoUExAW5_0;
	wire w_dff_B_ogw97NAZ1_0;
	wire w_dff_B_VQv6UVHk6_0;
	wire w_dff_B_QBMXYK116_0;
	wire w_dff_B_YHtLDvGi4_0;
	wire w_dff_B_DVQi1o885_0;
	wire w_dff_B_PP84ZHW99_0;
	wire w_dff_B_1SGkRLQA4_0;
	wire w_dff_B_qNjiej5C5_0;
	wire w_dff_B_ByIazu2g6_0;
	wire w_dff_B_zUO80eUi9_0;
	wire w_dff_B_5g0mg10I0_0;
	wire w_dff_B_xLNxPQP56_0;
	wire w_dff_B_BDrDtfkc8_0;
	wire w_dff_B_ZS5RtR481_0;
	wire w_dff_B_LEyHzAeA3_0;
	wire w_dff_B_zrSZD4I47_0;
	wire w_dff_B_gJ9PIjdI8_0;
	wire w_dff_B_HOTVZBKz6_0;
	wire w_dff_B_ka6z1FoH1_0;
	wire w_dff_B_8I44RRvp5_0;
	wire w_dff_B_atTc2hgQ9_0;
	wire w_dff_B_joWKk9zU8_0;
	wire w_dff_B_pzth4bdp0_0;
	wire w_dff_B_284155wq5_0;
	wire w_dff_B_1vZ8lB9m6_0;
	wire w_dff_B_0X0LIAop1_0;
	wire w_dff_B_XZ0A7KtN8_0;
	wire w_dff_B_mnnh0AzY7_0;
	wire w_dff_B_MKKp3jhp1_0;
	wire w_dff_B_RZoLLbOj0_0;
	wire w_dff_B_ENFkvwC06_0;
	wire w_dff_B_9mEdzbOZ5_0;
	wire w_dff_B_AgmQJTh00_0;
	wire w_dff_B_fToZhYKv6_0;
	wire w_dff_B_p9ed42J71_0;
	wire w_dff_B_GoAFN8DH7_0;
	wire w_dff_B_jQkod9A81_0;
	wire w_dff_B_Hgt3bEnx2_0;
	wire w_dff_B_C7skC0hb3_0;
	wire w_dff_B_V65TL54Q8_0;
	wire w_dff_B_IZRQj2473_0;
	wire w_dff_B_4eavRGSr6_0;
	wire w_dff_B_rZoTZyJt8_0;
	wire w_dff_B_3v5VLc1J9_0;
	wire w_dff_B_REMF3GuW0_0;
	wire w_dff_B_YL8zTHVl5_0;
	wire w_dff_B_9thUzuR96_0;
	wire w_dff_B_19GLMtJm4_0;
	wire w_dff_B_EbqXdmSo3_0;
	wire w_dff_B_6UmJmk6w2_0;
	wire w_dff_B_PPxofY7O6_0;
	wire w_dff_B_c4gdAp6b7_0;
	wire w_dff_B_vpmjKDyh7_0;
	wire w_dff_B_j2nwwKNV3_0;
	wire w_dff_B_rnPYDQLn4_0;
	wire w_dff_B_tcacvOZJ7_0;
	wire w_dff_B_w68Wzjw10_0;
	wire w_dff_B_8yU9wllU8_0;
	wire w_dff_B_FdVK2dLW7_0;
	wire w_dff_B_QI4Zre4z6_0;
	wire w_dff_B_0lZtMVcn2_0;
	wire w_dff_B_uFUJ54ht2_0;
	wire w_dff_B_sBZNRpfz4_0;
	wire w_dff_B_2QRWqBTN5_0;
	wire w_dff_B_smbicmKF2_0;
	wire w_dff_B_mdCtVYWR7_0;
	wire w_dff_B_HgspKiik1_0;
	wire w_dff_B_9Ky0V8JL3_0;
	wire w_dff_B_SeDHYRt34_0;
	wire w_dff_B_P7kR7Qdy5_0;
	wire w_dff_B_6G9lhlBa7_0;
	wire w_dff_B_pbLhd0ZI9_0;
	wire w_dff_B_m8tgTlRz8_0;
	wire w_dff_B_BKRcikdw8_0;
	wire w_dff_B_j67ywXjT4_0;
	wire w_dff_B_5Ra9CF982_0;
	wire w_dff_B_FiLo6R6S7_0;
	wire w_dff_B_5bEhIJ632_0;
	wire w_dff_B_jeXDElwt5_0;
	wire w_dff_B_bCG1tQmS9_0;
	wire w_dff_B_IjR9ApJg5_0;
	wire w_dff_B_7rPX4sM22_0;
	wire w_dff_B_sGrvLns29_0;
	wire w_dff_B_2OtMJ1Xt4_0;
	wire w_dff_B_68K6qTvt9_0;
	wire w_dff_B_eeev1QQd4_0;
	wire w_dff_B_hjcSyLNg5_0;
	wire w_dff_B_6M3CObuF1_0;
	wire w_dff_B_9eMXsrWy4_0;
	wire w_dff_B_Mh3FSkp80_0;
	wire w_dff_B_yWARzmpv9_0;
	wire w_dff_B_RxGkl3gm1_0;
	wire w_dff_B_qTLKcbfh6_0;
	wire w_dff_B_6KdzJKNr2_0;
	wire w_dff_B_Fbuael3j4_0;
	wire w_dff_B_QkoZ85Tr4_0;
	wire w_dff_B_1VDCeoYA1_0;
	wire w_dff_B_TxOxlGYx1_0;
	wire w_dff_B_g7IHH28r6_0;
	wire w_dff_B_OOLDaeKM9_0;
	wire w_dff_B_U5FsKTUb8_0;
	wire w_dff_B_bRcugeFv7_0;
	wire w_dff_B_oBKVmUkv2_0;
	wire w_dff_B_1uR9BjNH7_0;
	wire w_dff_B_3GpbkWYZ1_0;
	wire w_dff_B_yKw6r9jY3_0;
	wire w_dff_B_hHaX25Fb6_0;
	wire w_dff_B_qju38gGh4_0;
	wire w_dff_B_QE9vSeWv1_0;
	wire w_dff_B_jjYXaImP1_0;
	wire w_dff_B_javhpdaP0_0;
	wire w_dff_B_3cYRPfB37_0;
	wire w_dff_B_cfrql63o5_0;
	wire w_dff_B_JybZEV0g6_0;
	wire w_dff_B_3lg6fRCH6_0;
	wire w_dff_B_fMZ9bkJ64_0;
	wire w_dff_B_aMrycb0I8_0;
	wire w_dff_B_ErX8eh0w8_0;
	wire w_dff_B_fz9SrC2q4_0;
	wire w_dff_B_UOrXbJRB7_0;
	wire w_dff_B_FdPiqGdg7_0;
	wire w_dff_B_8Sw8H5AL9_0;
	wire w_dff_B_Kk8YkuMB3_0;
	wire w_dff_B_v4AOX7le2_0;
	wire w_dff_B_1OpR2KMz8_0;
	wire w_dff_B_b9FCcMva1_0;
	wire w_dff_B_TkMiZdKv2_0;
	wire w_dff_B_yXx7r8rJ8_0;
	wire w_dff_B_HDJXbPwf3_0;
	wire w_dff_B_NfgRmekj8_0;
	wire w_dff_B_8szD1fQj3_0;
	wire w_dff_B_XTu2tx6K5_0;
	wire w_dff_B_1Cp3Xlu70_0;
	wire w_dff_B_4i5xBvOj4_0;
	wire w_dff_B_sFCzxq8x1_0;
	wire w_dff_B_phmHkO1L6_0;
	wire w_dff_B_pUjW3O9p8_0;
	wire w_dff_B_anFKiTtd6_0;
	wire w_dff_B_H6faowjM1_0;
	wire w_dff_B_UMLMKIGX4_0;
	wire w_dff_B_3nIU2xaG7_0;
	wire w_dff_B_WuVoAzyj4_0;
	wire w_dff_B_B6fpBHaI4_0;
	wire w_dff_B_PCtYaWD78_0;
	wire w_dff_B_4nyGGiF76_0;
	wire w_dff_B_v7S6j6CY4_0;
	wire w_dff_B_9Q9O6KN22_0;
	wire w_dff_B_Ha3Ou0wu8_0;
	wire w_dff_B_1qy6kROB1_0;
	wire w_dff_B_kEvV7k6J1_0;
	wire w_dff_B_BziCGQdg9_0;
	wire w_dff_B_0mJkoMhS3_0;
	wire w_dff_B_IMvfyqJ12_0;
	wire w_dff_B_1yjF3upI3_0;
	wire w_dff_B_hU2xvfoD7_0;
	wire w_dff_B_jH1vbdlj8_0;
	wire w_dff_B_Q4Iyc5pC2_0;
	wire w_dff_B_GZusmrKV4_0;
	wire w_dff_B_kdLNS5yS3_0;
	wire w_dff_B_WHZpE7LF3_0;
	wire w_dff_B_3JNz2vpY1_0;
	wire w_dff_B_Gblky7394_0;
	wire w_dff_B_yf4HX0u41_0;
	wire w_dff_B_nvu97efN1_0;
	wire w_dff_B_qwVr1rC41_0;
	wire w_dff_B_2w3gAkD51_0;
	wire w_dff_B_GhXrqSip5_0;
	wire w_dff_B_Zt6Razf06_0;
	wire w_dff_B_sOUg29rq1_0;
	wire w_dff_B_iIcRMXxs5_0;
	wire w_dff_B_BUHZyAWR0_0;
	wire w_dff_B_FLyeW2pl1_0;
	wire w_dff_B_wWRlteQQ2_0;
	wire w_dff_B_PTeZlwlE6_0;
	wire w_dff_B_lHTRrGFV1_0;
	wire w_dff_B_ecVL8fmo2_0;
	wire w_dff_B_jVlAcpZ07_0;
	wire w_dff_B_KhIlBopL1_0;
	wire w_dff_B_eyergLvU9_0;
	wire w_dff_B_5meeMWcj3_0;
	wire w_dff_B_Xh6h7Du88_0;
	wire w_dff_B_bcVvLfRG8_0;
	wire w_dff_B_FSoIWlHL6_0;
	wire w_dff_B_xEbicrAq0_0;
	wire w_dff_B_A7qvzuar1_0;
	wire w_dff_B_aPcMadu43_0;
	wire w_dff_B_Oy2qUmD86_0;
	wire w_dff_B_DtXJgLC54_0;
	wire w_dff_B_3WtYBPXV5_0;
	wire w_dff_B_4eYAOaTo8_0;
	wire w_dff_B_T0S1fxii1_0;
	wire w_dff_B_b1Ymardl7_0;
	wire w_dff_B_pqJMNoT86_0;
	wire w_dff_B_NfLNTYs39_0;
	wire w_dff_B_KyDhcp9D5_0;
	wire w_dff_B_LCasklDP8_0;
	wire w_dff_B_MMDUX33q7_0;
	wire w_dff_B_An18KtIF3_0;
	wire w_dff_B_RAJSq0ts6_0;
	wire w_dff_B_HuWpDLE56_0;
	wire w_dff_B_NhwbHhev1_0;
	wire w_dff_B_YRI7OsJv7_0;
	wire w_dff_B_IL0XQ2Gf9_0;
	wire w_dff_B_ZSWQYgik1_0;
	wire w_dff_B_3UeKj0wI6_0;
	wire w_dff_B_td0aycKm9_0;
	wire w_dff_B_RtpiBDq05_0;
	wire w_dff_B_7OGDhqiW4_0;
	wire w_dff_B_eBH4Nj4a2_0;
	wire w_dff_B_bXyXzKVd9_0;
	wire w_dff_B_QDR0W5Gu0_0;
	wire w_dff_B_6u9PMJ075_0;
	wire w_dff_B_s74rdd5T0_0;
	wire w_dff_B_rLBFfNfn7_0;
	wire w_dff_B_ES4MEgR89_0;
	wire w_dff_B_T2zANDhP2_0;
	wire w_dff_B_2jSCno820_0;
	wire w_dff_B_vqvVnJq35_0;
	wire w_dff_B_jIGXsslq5_0;
	wire w_dff_B_KiDbaGfZ6_0;
	wire w_dff_B_fpRKzTs10_0;
	wire w_dff_B_sIING38w8_0;
	wire w_dff_B_ZsY46qQz4_0;
	wire w_dff_B_ErAW2XY51_0;
	wire w_dff_B_gEFk0bmc1_0;
	wire w_dff_B_3xKuW1hJ6_0;
	wire w_dff_B_HhkzoLIB2_0;
	wire w_dff_B_MuZniDyC9_0;
	wire w_dff_B_KuwhWxoR5_0;
	wire w_dff_B_fhhbusxU7_0;
	wire w_dff_B_hDHP5zhU4_0;
	wire w_dff_B_nzYEIVwr7_0;
	wire w_dff_B_46uvAGbh6_0;
	wire w_dff_B_AHKtGtyA9_0;
	wire w_dff_B_2ghRHon87_0;
	wire w_dff_B_bhSZisTk0_0;
	wire w_dff_B_p3naK36l8_0;
	wire w_dff_B_FVbAlllk6_0;
	wire w_dff_B_Dn0jecqQ2_0;
	wire w_dff_B_ohuDVRCW4_0;
	wire w_dff_B_2IA0E61U7_0;
	wire w_dff_B_Up3ANdop7_0;
	wire w_dff_B_yeLqkkRE2_0;
	wire w_dff_B_SVmc92bt7_0;
	wire w_dff_B_WJJ7y8Tu3_0;
	wire w_dff_B_C0Lb6Ahd1_0;
	wire w_dff_B_YuupTCKx4_0;
	wire w_dff_B_uDFyPzGp7_0;
	wire w_dff_B_ZhgGiEm79_0;
	wire w_dff_B_3WmfKVE20_0;
	wire w_dff_B_kz2WX4gh7_0;
	wire w_dff_B_n6Brr1eb3_0;
	wire w_dff_B_m9yS7dMG9_0;
	wire w_dff_B_LkM9bzTO1_0;
	wire w_dff_B_XA6Jgvc14_0;
	wire w_dff_B_ZvEhLFv78_0;
	wire w_dff_B_45o3fjhQ8_0;
	wire w_dff_B_EATydhzE5_0;
	wire w_dff_B_gVXHyWQB0_0;
	wire w_dff_B_DmkAllKZ6_0;
	wire w_dff_B_jn1ccoQw8_0;
	wire w_dff_B_G7wQ0CCE4_0;
	wire w_dff_B_HlSrfZPG6_0;
	wire w_dff_B_3yoVrpNn1_0;
	wire w_dff_B_6VPqM88X8_0;
	wire w_dff_B_ZmveveaH3_0;
	wire w_dff_B_FUMUhn2t4_0;
	wire w_dff_B_DRGqoQst1_0;
	wire w_dff_B_t56nAR5Z5_0;
	wire w_dff_B_bvUpw8fz1_0;
	wire w_dff_B_AGsYW8xa2_0;
	wire w_dff_B_rtt6Mkn48_0;
	wire w_dff_B_HLpB3qmL5_0;
	wire w_dff_B_9YJnsIyF7_0;
	wire w_dff_B_baHvFq3V2_0;
	wire w_dff_B_XFUunqJn0_0;
	wire w_dff_B_nlEza59P2_0;
	wire w_dff_B_5iTdFiWG2_0;
	wire w_dff_B_5ik7dOD48_0;
	wire w_dff_B_PaVAueOx8_0;
	wire w_dff_B_Y4t0NgXz6_0;
	wire w_dff_B_qsS8u5Pp1_0;
	wire w_dff_B_BRhErMvA7_0;
	wire w_dff_B_pHw6SCC42_0;
	wire w_dff_B_14qw1mBa3_0;
	wire w_dff_B_TE2W0Imk6_0;
	wire w_dff_B_MgAJtuB17_0;
	wire w_dff_B_XGT53Xsq2_0;
	wire w_dff_B_5TxQLPZP6_0;
	wire w_dff_B_YvLwp3Ut5_0;
	wire w_dff_B_ol8bmYDi8_0;
	wire w_dff_B_xKAiLwJm3_0;
	wire w_dff_B_bgj8K81M1_0;
	wire w_dff_B_uxuYl4C17_0;
	wire w_dff_B_qSlEKpkG6_0;
	wire w_dff_B_LsxtOyh74_0;
	wire w_dff_B_pa6Wo2BO4_0;
	wire w_dff_B_OfLeGgiB6_0;
	wire w_dff_B_zCGL2FI74_0;
	wire w_dff_B_AnGKKJt33_0;
	wire w_dff_B_w6bDZ4HN5_0;
	wire w_dff_B_Z5lumHrF3_0;
	wire w_dff_B_NqhsmJQc3_0;
	wire w_dff_B_2I9oic4J2_0;
	wire w_dff_B_jE3gGIn46_0;
	wire w_dff_B_QmriqQQA9_0;
	wire w_dff_B_E02EDSMt1_0;
	wire w_dff_B_P2qyRF8K4_0;
	wire w_dff_B_AnUBsgCg0_0;
	wire w_dff_B_ciRIYHl29_0;
	wire w_dff_B_bjaqF0ZD9_0;
	wire w_dff_B_7k9h5O3k6_0;
	wire w_dff_B_BNluhNy42_0;
	wire w_dff_B_QIT3SBBW6_0;
	wire w_dff_B_JQzpuMXS8_0;
	wire w_dff_B_bqCTjpcL9_0;
	wire w_dff_B_uX9IqRB81_0;
	wire w_dff_B_mzA3Cg8J6_0;
	wire w_dff_B_xO3KsHO66_0;
	wire w_dff_B_4SmdUwi71_0;
	wire w_dff_B_H8oqT6J93_0;
	wire w_dff_B_4XzJK8Gg6_0;
	wire w_dff_B_1XX0WgBP1_0;
	wire w_dff_B_R6YUz3z28_0;
	wire w_dff_B_8yFHfUiN2_0;
	wire w_dff_B_FeM8thi53_0;
	wire w_dff_B_F4p0snYn0_0;
	wire w_dff_B_AU3wcHUQ1_0;
	wire w_dff_B_3vKBcR4y2_0;
	wire w_dff_B_XevCGRFb7_0;
	wire w_dff_B_b9l9YqWJ8_0;
	wire w_dff_B_3JKDk23U9_0;
	wire w_dff_B_GdCBevGf7_0;
	wire w_dff_B_fjQdDwis8_0;
	wire w_dff_B_iOjoLuk30_0;
	wire w_dff_B_yVtB9mxq8_0;
	wire w_dff_B_y1DUNIKE2_0;
	wire w_dff_B_ktNdov5X8_0;
	wire w_dff_B_BKRWFx523_0;
	wire w_dff_B_EI038q2N7_0;
	wire w_dff_B_b1QayugI9_0;
	wire w_dff_B_gtdu5Yxn6_0;
	wire w_dff_B_7ZLA1AEU3_0;
	wire w_dff_B_kmfv2In99_0;
	wire w_dff_B_qYy2l2GS4_0;
	wire w_dff_B_4QyGyHa53_0;
	wire w_dff_B_z3YLYRms7_0;
	wire w_dff_B_uq6nkgFO0_0;
	wire w_dff_B_EVYUVjSW2_0;
	wire w_dff_B_Yyrez7Fi4_0;
	wire w_dff_B_bkkM4V7I5_0;
	wire w_dff_B_SSO2b7TT0_0;
	wire w_dff_B_4ybstWh80_0;
	wire w_dff_B_2xbCP0oy1_0;
	wire w_dff_B_6wLIYx6m8_0;
	wire w_dff_B_Dj6JnDZ11_0;
	wire w_dff_B_lHMxqmMG1_0;
	wire w_dff_B_Lu0eTXOt5_0;
	wire w_dff_B_M8n3SWsm2_0;
	wire w_dff_B_QFKVtpy08_0;
	wire w_dff_B_W9RkfTyR1_0;
	wire w_dff_B_WqYsR6aj0_0;
	wire w_dff_B_JG6RM1k87_0;
	wire w_dff_B_rtgGt7my7_0;
	wire w_dff_B_QlndlzQS4_0;
	wire w_dff_B_du85iw1C5_0;
	wire w_dff_B_s14OcBtD5_0;
	wire w_dff_B_tidPtZPJ4_0;
	wire w_dff_B_VZw7honL6_0;
	wire w_dff_B_TT45QkOS2_0;
	wire w_dff_B_bjiHRgdS3_0;
	wire w_dff_B_Ss7i2Bw90_0;
	wire w_dff_B_0zDidFUn2_0;
	wire w_dff_B_Qek5J5k80_0;
	wire w_dff_B_0QfYaqb86_0;
	wire w_dff_B_o9yTFobN5_0;
	wire w_dff_B_n0xpXh2y6_0;
	wire w_dff_B_Ajd5YtvK8_0;
	wire w_dff_B_FskJtOUr8_0;
	wire w_dff_B_b30rvFHq0_0;
	wire w_dff_B_pGdrETgs8_0;
	wire w_dff_B_7icUPGR23_0;
	wire w_dff_B_L2IWobFb8_0;
	wire w_dff_B_0t8LD5oz6_0;
	wire w_dff_B_YvoUw0471_0;
	wire w_dff_B_f7FrN3YU6_0;
	wire w_dff_B_Y1DsgdCH2_0;
	wire w_dff_B_aESggMQI6_0;
	wire w_dff_B_SsLNApqS7_0;
	wire w_dff_B_aBvX1duK8_0;
	wire w_dff_B_MuOTdBbz6_0;
	wire w_dff_B_sui8Kq456_0;
	wire w_dff_B_PcdbTwvc7_0;
	wire w_dff_B_aNnGcEt09_0;
	wire w_dff_B_PU1wLCQP7_0;
	wire w_dff_B_n7s0thyv7_0;
	wire w_dff_B_3QDAHMmj4_0;
	wire w_dff_B_QlbG0Nm58_0;
	wire w_dff_B_kdyOUyGn4_0;
	wire w_dff_B_RZbOA3Em1_0;
	wire w_dff_B_TSji5Tyv4_0;
	wire w_dff_B_DB401HXm8_0;
	wire w_dff_B_eFVXScsq6_0;
	wire w_dff_B_sEGwsu4a0_0;
	wire w_dff_B_AF3T9QpX6_0;
	wire w_dff_B_i4xc8eaS5_0;
	wire w_dff_B_YZX0D7ZM2_0;
	wire w_dff_B_07X3RyDd9_0;
	wire w_dff_B_Q8QjIA982_0;
	wire w_dff_B_0ji4sAsF1_0;
	wire w_dff_B_caf0nWoP4_0;
	wire w_dff_B_cEKkY6bt2_0;
	wire w_dff_B_hTmF8Qd97_0;
	wire w_dff_B_38UupXcB0_0;
	wire w_dff_B_rHs3VIWw9_0;
	wire w_dff_B_DsdfOOoK5_0;
	wire w_dff_B_LWTCzuch2_0;
	wire w_dff_B_wNh2ztIJ3_0;
	wire w_dff_B_d7f7UIjm7_0;
	wire w_dff_B_OQgYeVkg6_0;
	wire w_dff_B_GKypNqJd2_0;
	wire w_dff_B_qvwEj2Hf4_0;
	wire w_dff_B_YpJDZxaE6_0;
	wire w_dff_B_Ucig1agG3_0;
	wire w_dff_B_u9OY4RPb0_0;
	wire w_dff_B_uNC1l8Z80_0;
	wire w_dff_B_8U7G98lZ4_0;
	wire w_dff_B_YEsUQv1B3_0;
	wire w_dff_B_VxjKO3032_0;
	wire w_dff_B_KCv9h0wh2_0;
	wire w_dff_B_XuMixnZF9_0;
	wire w_dff_B_i84eCWYK5_0;
	wire w_dff_B_U6iwCUZI0_0;
	wire w_dff_B_a5doqkpu9_0;
	wire w_dff_B_57llpIob9_0;
	wire w_dff_B_7vRhbgR89_0;
	wire w_dff_B_oEK9mALP8_0;
	wire w_dff_B_vIkxOLPx8_0;
	wire w_dff_B_E6iKKrI60_0;
	wire w_dff_B_Uyuf2mfa0_0;
	wire w_dff_B_1Xzww8T78_0;
	wire w_dff_B_njK3vFMj2_0;
	wire w_dff_B_HhC6SGrG6_0;
	wire w_dff_B_TMD9qqX40_0;
	wire w_dff_B_sGe1J2sr6_0;
	wire w_dff_B_WgXCP8oB1_0;
	wire w_dff_B_WOjvGSCr8_0;
	wire w_dff_B_zakEMstQ7_0;
	wire w_dff_B_ss1rzqcX8_0;
	wire w_dff_B_6NJbhcMc8_0;
	wire w_dff_B_gEKVGIrr0_0;
	wire w_dff_B_TeeUhAJH4_0;
	wire w_dff_B_pwRMvVCF2_0;
	wire w_dff_B_0Btbh8ue2_0;
	wire w_dff_B_REEkhnWJ6_0;
	wire w_dff_B_osRhnc4L7_0;
	wire w_dff_B_urmRmVsn4_0;
	wire w_dff_B_DyS7xSXY7_0;
	wire w_dff_B_NRtyQ9LL2_0;
	wire w_dff_B_pSYE8h1n8_0;
	wire w_dff_B_CWAAsrHB5_0;
	wire w_dff_B_j4qLCyvR0_0;
	wire w_dff_B_AfDCJyYt4_0;
	wire w_dff_B_Rrv7Kelz8_0;
	wire w_dff_B_qX4CVjCr3_0;
	wire w_dff_B_CAupgnU25_0;
	wire w_dff_B_0a5auGct7_0;
	wire w_dff_B_OstfHIGV8_0;
	wire w_dff_B_JlgY5HaC6_0;
	wire w_dff_B_CArRZfBW6_0;
	wire w_dff_B_LhDuKVVU8_0;
	wire w_dff_B_5FrZBA1s4_0;
	wire w_dff_B_XQ9Rjv7h6_0;
	wire w_dff_B_a8gC8uVN9_0;
	wire w_dff_B_483hyO8g4_0;
	wire w_dff_B_qEAYffRl1_0;
	wire w_dff_B_kcLCUR772_0;
	wire w_dff_B_7szMmokO0_0;
	wire w_dff_B_KMCHcUBV0_0;
	wire w_dff_B_heNREE0Y6_0;
	wire w_dff_B_H6bPQElY1_0;
	wire w_dff_B_gz2OrYPI9_0;
	wire w_dff_B_nAxAlxz78_0;
	wire w_dff_B_5wyFce4n6_0;
	wire w_dff_B_quUKTcuk1_0;
	wire w_dff_B_oPL44UVW6_0;
	wire w_dff_B_iE6Jz1SW3_0;
	wire w_dff_B_DE3XsQ635_0;
	wire w_dff_B_jnOUUyph7_0;
	wire w_dff_B_nn041RUC8_0;
	wire w_dff_B_Ott5IRF98_0;
	wire w_dff_B_abhOlZYA7_0;
	wire w_dff_B_lQFKS9cz2_0;
	wire w_dff_B_M9azyQZp9_0;
	wire w_dff_B_0H2INgDW0_0;
	wire w_dff_B_ZiTnUagd1_0;
	wire w_dff_B_CbJ52ZMk7_0;
	wire w_dff_B_PQxVaC210_0;
	wire w_dff_B_OR5nETYs0_0;
	wire w_dff_B_T319vpfa4_0;
	wire w_dff_B_f8akAoUd3_0;
	wire w_dff_B_qyLKJi1A2_0;
	wire w_dff_B_aC6sKNmO2_0;
	wire w_dff_B_8d2RFYTT9_0;
	wire w_dff_B_i0l3dmF45_0;
	wire w_dff_B_byNuTY3P8_0;
	wire w_dff_B_XmlN3y7k5_0;
	wire w_dff_B_kTjdueIQ1_0;
	wire w_dff_B_1psdxSCW2_0;
	wire w_dff_B_WdQRaDsG6_0;
	wire w_dff_B_t91WNSGm1_0;
	wire w_dff_B_IEwWzTiz3_0;
	wire w_dff_B_mf48kb8J1_0;
	wire w_dff_B_AeV4wvcd9_0;
	wire w_dff_B_PJyJoXTf0_0;
	wire w_dff_B_t74qSl9a8_0;
	wire w_dff_B_IZc4wbgh8_0;
	wire w_dff_B_KbFwBhXd3_0;
	wire w_dff_B_oV4kSYUM3_0;
	wire w_dff_B_71zA2kTt4_0;
	wire w_dff_B_3ieDKJEX2_0;
	wire w_dff_B_goPzpxyf9_0;
	wire w_dff_B_8fhEuSZk1_0;
	wire w_dff_B_QdgWjF0B1_0;
	wire w_dff_B_9spmQcSQ7_0;
	wire w_dff_B_wvt8aCLK8_0;
	wire w_dff_B_LHvcpfcj5_0;
	wire w_dff_B_MkSo5soc6_0;
	wire w_dff_B_Z36m5uF72_0;
	wire w_dff_B_4RoGkf3r2_0;
	wire w_dff_B_hFDQBF8z9_0;
	wire w_dff_B_AeXMupvd9_0;
	wire w_dff_B_B3apuCFj8_0;
	wire w_dff_B_prjaBGQ89_0;
	wire w_dff_B_OMpeXpLq6_0;
	wire w_dff_B_g1TsJgxk4_0;
	wire w_dff_B_mUKxOZ513_0;
	wire w_dff_B_SeZRqgZB9_0;
	wire w_dff_B_wSkievnF8_0;
	wire w_dff_B_s2zO63RE6_0;
	wire w_dff_B_tyiABXnk7_0;
	wire w_dff_B_PkwEA4Rc9_0;
	wire w_dff_B_gVaUN1NU5_0;
	wire w_dff_B_9P7yv7Ye7_0;
	wire w_dff_B_Vr9tWKYM4_0;
	wire w_dff_B_yp9b0hnF4_0;
	wire w_dff_B_1D79UTZf5_0;
	wire w_dff_B_VAj705Ce6_0;
	wire w_dff_B_qTwxy58w0_0;
	wire w_dff_B_e8dfjaRZ9_0;
	wire w_dff_B_FJS06Muv8_0;
	wire w_dff_B_eMzPEEbX4_0;
	wire w_dff_B_gXpXSEfj8_0;
	wire w_dff_B_lewfv43k5_0;
	wire w_dff_B_xIRT4pZK3_0;
	wire w_dff_B_MT6YAPpC5_0;
	wire w_dff_B_3xJzgs0k4_0;
	wire w_dff_B_HjcxW1gs6_0;
	wire w_dff_B_EzdcUTXM9_0;
	wire w_dff_B_jx9QqAFk1_0;
	wire w_dff_B_pYIFf5wj1_0;
	wire w_dff_B_C8hsQ1t99_0;
	wire w_dff_B_um4WyG5E7_0;
	wire w_dff_B_Mh8g19Sk5_0;
	wire w_dff_B_eh7BWXtk3_0;
	wire w_dff_B_RRKtcs4q6_0;
	wire w_dff_B_MueYSLX36_0;
	wire w_dff_B_wooc5c0P3_0;
	wire w_dff_B_ziaGA0rp2_0;
	wire w_dff_B_WXptrmNp1_0;
	wire w_dff_B_3zbQGrC62_0;
	wire w_dff_B_y6XPv0xv4_0;
	wire w_dff_B_ci8m6xmH5_0;
	wire w_dff_B_DbwP4hdC4_0;
	wire w_dff_B_XE6q6rOO0_0;
	wire w_dff_B_5DMJKqlB4_0;
	wire w_dff_B_eCn7Nu3a1_0;
	wire w_dff_B_JolXBKwI8_0;
	wire w_dff_B_Bq8QRUuD3_0;
	wire w_dff_B_ck9hUul88_0;
	wire w_dff_B_WIJZ78gw8_0;
	wire w_dff_B_oZAz2n0E1_0;
	wire w_dff_B_3xVA9W6i1_0;
	wire w_dff_B_XQPE7p0h1_0;
	wire w_dff_B_cd2KeBby1_0;
	wire w_dff_B_1uRJoPpO1_0;
	wire w_dff_B_jTqEqb1H4_0;
	wire w_dff_B_hbt8k0ef1_0;
	wire w_dff_B_MYelRpm85_0;
	wire w_dff_B_pTlWKZ6x2_0;
	wire w_dff_B_d8VofKpQ0_0;
	wire w_dff_B_wbZG7QoE8_0;
	wire w_dff_B_phoMujdh2_0;
	wire w_dff_B_jVs3W3jJ7_0;
	wire w_dff_B_qI0VCpAH7_0;
	wire w_dff_B_GWSHrsgV9_0;
	wire w_dff_B_Qg6BnTtV9_0;
	wire w_dff_B_6hzz9GG38_0;
	wire w_dff_B_sbZw3v7L2_0;
	wire w_dff_B_BjYlc2CB4_0;
	wire w_dff_B_LXw0OWrp3_0;
	wire w_dff_B_UDcq6OOm5_0;
	wire w_dff_B_WuYhmjkv6_0;
	wire w_dff_B_oHjSdhyP1_0;
	wire w_dff_B_DvEsZjMl7_0;
	wire w_dff_B_AgOf2Dca6_0;
	wire w_dff_B_kaMqvGnX4_0;
	wire w_dff_B_LMcbZJOa8_0;
	wire w_dff_B_D4G1r1cU8_0;
	wire w_dff_B_6vOmPyiY1_0;
	wire w_dff_B_aeNsupF99_0;
	wire w_dff_B_T4j0H2KR2_0;
	wire w_dff_B_fphVRBL66_0;
	wire w_dff_B_2c6vUZbK5_0;
	wire w_dff_B_ZEmVIxwi4_0;
	wire w_dff_B_HnKcbF1T8_0;
	wire w_dff_B_9wjeYoBY6_0;
	wire w_dff_B_nWqcM3FS5_0;
	wire w_dff_B_7QFPOCrV6_0;
	wire w_dff_B_TgiI1lZR5_0;
	wire w_dff_B_ClKSzvHU7_0;
	wire w_dff_B_IfW2Sv7q7_0;
	wire w_dff_B_NeD4Nn9y8_0;
	wire w_dff_B_UPVdnHXy5_0;
	wire w_dff_B_6zU42Z0I9_0;
	wire w_dff_B_cAeYRSUq6_0;
	wire w_dff_B_rkqSrGhN4_0;
	wire w_dff_B_uw8WfP724_0;
	wire w_dff_B_SkhbmHSz9_0;
	wire w_dff_B_9rgiGrKw2_0;
	wire w_dff_B_DyeB2vL03_0;
	wire w_dff_B_mcwkPAkL2_0;
	wire w_dff_B_XuY9E4Ou4_0;
	wire w_dff_B_BppOGXt43_0;
	wire w_dff_B_pZ6P6bM07_0;
	wire w_dff_B_uuKE7prV9_0;
	wire w_dff_B_YFkhXDhi0_0;
	wire w_dff_B_ofaTlYyf5_0;
	wire w_dff_B_l1BQO1Bu9_0;
	wire w_dff_B_87RqLrR94_0;
	wire w_dff_B_BohxU8tM5_0;
	wire w_dff_B_FT6qOtrS4_0;
	wire w_dff_B_EuTOQkN66_0;
	wire w_dff_B_Kr4Saxpw5_0;
	wire w_dff_B_aN2YQPxw9_0;
	wire w_dff_B_lvOHKtlw4_0;
	wire w_dff_B_Bh5TkV9c9_0;
	wire w_dff_B_yBY6zIKE7_0;
	wire w_dff_B_OktgxKr12_0;
	wire w_dff_B_jXu0gceh6_0;
	wire w_dff_B_RdfHookR8_0;
	wire w_dff_B_H0luIVyz1_0;
	wire w_dff_B_zzFl00kT8_0;
	wire w_dff_B_Mpjw50Ap0_0;
	wire w_dff_B_IY2l35Pl2_0;
	wire w_dff_B_WO4CwQt12_0;
	wire w_dff_B_vTtcFnaX1_0;
	wire w_dff_B_Ov5Jfpqt1_0;
	wire w_dff_B_9CkXA9AG3_0;
	wire w_dff_B_gVkbTBwR4_0;
	wire w_dff_B_vlndYaxx5_0;
	wire w_dff_B_r3RtS4sf5_0;
	wire w_dff_B_20S2Q5oJ1_0;
	wire w_dff_B_ZaARAyP08_0;
	wire w_dff_B_aG5BVySM7_0;
	wire w_dff_B_vqfDjWX14_0;
	wire w_dff_B_lx4KyX9J6_0;
	wire w_dff_B_G6kldeH14_0;
	wire w_dff_B_v8aBzas02_0;
	wire w_dff_B_uVItd6s24_0;
	wire w_dff_B_ZLMwJtYI1_0;
	wire w_dff_B_1FVKKcoT6_0;
	wire w_dff_B_SRgO1VNq5_0;
	wire w_dff_B_TSH1xZyN5_0;
	wire w_dff_B_Vt8WOKXG1_0;
	wire w_dff_B_xOmJmBh08_0;
	wire w_dff_B_yMpw4ghJ6_0;
	wire w_dff_B_E0UEn0QU0_0;
	wire w_dff_B_lIfmeSyV2_0;
	wire w_dff_B_hcdQaGWh9_0;
	wire w_dff_B_GZvz9KB76_0;
	wire w_dff_B_Q2Hc1GQB1_0;
	wire w_dff_B_8Dm77OtX9_0;
	wire w_dff_B_atmx5RPm8_1;
	wire w_dff_B_RFADscL76_1;
	wire w_dff_B_rj31xIls3_1;
	wire w_dff_B_9RGDo8fL4_1;
	wire w_dff_B_oeDww5zt9_1;
	wire w_dff_B_RPTgCTBP0_1;
	wire w_dff_B_x6gtpROe7_1;
	wire w_dff_B_4EzZvJGs4_1;
	wire w_dff_B_AmluzxDU4_1;
	wire w_dff_B_tv8mwf8P2_1;
	wire w_dff_B_igS4eQLx5_1;
	wire w_dff_B_U48KMSgO0_1;
	wire w_dff_B_NczshOmV4_1;
	wire w_dff_B_THkn9HEh5_1;
	wire w_dff_B_9wMpNnnR9_1;
	wire w_dff_B_79Q61mpM9_1;
	wire w_dff_B_9PuQADfm2_1;
	wire w_dff_B_okaXoeu12_1;
	wire w_dff_B_JFAqEzkK9_1;
	wire w_dff_B_Z5PLn4Da1_1;
	wire w_dff_B_6CiEtYja6_1;
	wire w_dff_B_2vwo12f40_1;
	wire w_dff_B_rqpUrkEP4_1;
	wire w_dff_B_zt1VhDA51_1;
	wire w_dff_B_bd1VUPjf7_1;
	wire w_dff_B_HGpO0FUN8_1;
	wire w_dff_B_GsGj0xnB0_1;
	wire w_dff_B_WBxiJ5p85_1;
	wire w_dff_B_M7puSxrt0_1;
	wire w_dff_B_5OJSG2Qz4_1;
	wire w_dff_B_JJKXNAmW8_1;
	wire w_dff_B_XLWcYd4j3_1;
	wire w_dff_B_72ROqm773_1;
	wire w_dff_B_p25PetQz4_1;
	wire w_dff_B_67EOdVvO7_1;
	wire w_dff_B_AYhQO0aq8_1;
	wire w_dff_B_76oJad779_1;
	wire w_dff_B_rP15x5Rj0_1;
	wire w_dff_B_up7mT3Jm8_1;
	wire w_dff_B_KFzFLXDC0_1;
	wire w_dff_B_VY05avO17_1;
	wire w_dff_B_S5uGMGjZ9_1;
	wire w_dff_B_jCQhqh0Q3_1;
	wire w_dff_B_w0dy3pmO6_1;
	wire w_dff_B_T6It8k2d6_1;
	wire w_dff_B_rtoXt2Is2_1;
	wire w_dff_B_g2MJLP8o2_1;
	wire w_dff_B_whyfvX1e7_1;
	wire w_dff_B_HZYjyU0U5_1;
	wire w_dff_B_oQqu21dV9_1;
	wire w_dff_B_DRUxcFe53_1;
	wire w_dff_B_WzSQX1Jb5_1;
	wire w_dff_B_v9ivZ9ad6_1;
	wire w_dff_B_gYpFQRhC0_1;
	wire w_dff_B_6w1SuZ9p1_1;
	wire w_dff_B_3p7OZ9v27_1;
	wire w_dff_B_dMb07bMO2_1;
	wire w_dff_B_pItQfPMm5_1;
	wire w_dff_B_HX5bYkUY3_1;
	wire w_dff_B_1FMtGHUR4_1;
	wire w_dff_B_cYrW1LaP2_1;
	wire w_dff_B_XzpDLXSC2_1;
	wire w_dff_B_LfM2WKy50_1;
	wire w_dff_B_V5Hlthry0_1;
	wire w_dff_B_Y42FY6WM1_1;
	wire w_dff_B_4gytCVG11_1;
	wire w_dff_B_G4aqjBaa6_1;
	wire w_dff_B_Wnrjcml20_1;
	wire w_dff_B_94XqCZLk3_1;
	wire w_dff_B_PfKSA2qF1_1;
	wire w_dff_B_KgBkMctq7_1;
	wire w_dff_B_OjoujAV64_1;
	wire w_dff_B_HynhC1Us7_1;
	wire w_dff_B_NQC4b47e6_1;
	wire w_dff_B_1tKqnsoN1_1;
	wire w_dff_B_uGDjLqrh9_1;
	wire w_dff_B_Vl6FtdEh6_1;
	wire w_dff_B_C6bW0Lci0_1;
	wire w_dff_B_ZkHqpgI72_1;
	wire w_dff_B_G8a6zfWg1_1;
	wire w_dff_B_4LuSDWLC6_1;
	wire w_dff_B_9mDyfVzL3_1;
	wire w_dff_B_YPSKTM3S9_1;
	wire w_dff_B_PRKFr2OB3_1;
	wire w_dff_B_3jV6T0em6_1;
	wire w_dff_B_RFINkQKi6_1;
	wire w_dff_B_reVxmV880_1;
	wire w_dff_B_2zQ7FImu0_1;
	wire w_dff_B_dh03SZt34_1;
	wire w_dff_B_ldiTaqoA7_1;
	wire w_dff_B_C5rcPgpM8_1;
	wire w_dff_B_QPQLq1Oy9_1;
	wire w_dff_B_lvX0xXKI8_1;
	wire w_dff_B_rgz1z64h0_1;
	wire w_dff_B_PyqAeOa11_1;
	wire w_dff_B_wOfb5myz5_1;
	wire w_dff_B_xNcuImkN8_1;
	wire w_dff_B_t6eym27f6_1;
	wire w_dff_B_53l1Clmq1_1;
	wire w_dff_B_fCkwkyjV4_1;
	wire w_dff_B_DJ7IG5Eh6_1;
	wire w_dff_B_l3OTR7B54_1;
	wire w_dff_B_qMaKviYj5_1;
	wire w_dff_B_KaLZeSy47_1;
	wire w_dff_B_mv5YzRGw0_1;
	wire w_dff_B_e5DQr9QO4_1;
	wire w_dff_B_n6QN3WIB6_1;
	wire w_dff_B_x0BLhzmH2_1;
	wire w_dff_B_QdGEdET97_1;
	wire w_dff_B_4mX8BWrB6_1;
	wire w_dff_B_UigGvA6R5_1;
	wire w_dff_B_8QcYi2eM7_1;
	wire w_dff_B_QJqq90ea5_1;
	wire w_dff_B_9bOUD3e91_1;
	wire w_dff_B_LP806dpe2_1;
	wire w_dff_B_FTExwWGv4_1;
	wire w_dff_B_RCPZkv7G0_1;
	wire w_dff_B_NaKG4y3Z2_1;
	wire w_dff_B_HRz2cCEW6_1;
	wire w_dff_B_WC60V9Pu8_1;
	wire w_dff_B_gzY9tO7N6_1;
	wire w_dff_B_6uRnwMLP0_1;
	wire w_dff_B_5QD35np92_1;
	wire w_dff_B_d1nf5OLW0_1;
	wire w_dff_B_cokVGotX5_1;
	wire w_dff_B_tpBuigwr1_1;
	wire w_dff_B_66p7sXjF1_1;
	wire w_dff_B_ZhSybxxK6_0;
	wire w_dff_B_HR6ojHVk8_0;
	wire w_dff_B_7v69VILJ0_0;
	wire w_dff_B_pxZt5sZd2_0;
	wire w_dff_B_CTEC44q93_0;
	wire w_dff_B_tUSTaSsl3_0;
	wire w_dff_B_T9b8DQA04_0;
	wire w_dff_B_rGAOrHRK2_0;
	wire w_dff_B_fCOsxztJ2_0;
	wire w_dff_B_r98hkcrQ3_0;
	wire w_dff_B_Ah5Lmctq4_0;
	wire w_dff_B_JiODjbEz2_0;
	wire w_dff_B_U6Q9QYTM3_0;
	wire w_dff_B_ERbzeH3g0_0;
	wire w_dff_B_ia2eZ6ML2_0;
	wire w_dff_B_iVplwo8H9_0;
	wire w_dff_B_yUEcPzMJ8_0;
	wire w_dff_B_t1A2hG7x9_0;
	wire w_dff_B_QdtDZF1S8_0;
	wire w_dff_B_EVcLzrgm9_0;
	wire w_dff_B_slC5Nc3n2_0;
	wire w_dff_B_XXcTucB50_0;
	wire w_dff_B_2D1X5yUO2_0;
	wire w_dff_B_K180yQkN7_0;
	wire w_dff_B_qWhpoLDA6_0;
	wire w_dff_B_aT2LDygW3_0;
	wire w_dff_B_vXRpq0DC2_0;
	wire w_dff_B_V1JEaggK4_0;
	wire w_dff_B_izUq2Um46_0;
	wire w_dff_B_I0K9myuV1_0;
	wire w_dff_B_sTaUWHyB2_0;
	wire w_dff_B_fGAkXdOh0_0;
	wire w_dff_B_XO1po3HH2_0;
	wire w_dff_B_9tav4sVA3_0;
	wire w_dff_B_dFPmVX9Y9_0;
	wire w_dff_B_Wed9gell2_0;
	wire w_dff_B_Vwnu2Rxe2_0;
	wire w_dff_B_C9l0aCj93_0;
	wire w_dff_B_h369j09H8_0;
	wire w_dff_B_TAuZZkPz3_0;
	wire w_dff_B_HlRPPLr95_0;
	wire w_dff_B_QnUObPUF9_0;
	wire w_dff_B_Z1hgLreU2_0;
	wire w_dff_B_qv50o4BA2_0;
	wire w_dff_B_o0Xx4yWp2_0;
	wire w_dff_B_U0qfYNmh5_0;
	wire w_dff_B_ChDSmj630_0;
	wire w_dff_B_oFOHarpP0_0;
	wire w_dff_B_99EVfNFn0_0;
	wire w_dff_B_d3FmXBNv1_0;
	wire w_dff_B_P0Yr2uRG2_0;
	wire w_dff_B_1Va7SEkL2_0;
	wire w_dff_B_2fTAI0Us1_0;
	wire w_dff_B_6Eg9timZ0_0;
	wire w_dff_B_1pfZkSI01_0;
	wire w_dff_B_TibFc1XT8_0;
	wire w_dff_B_SR7b3DuN5_0;
	wire w_dff_B_Yj5jmHab9_0;
	wire w_dff_B_WOyGo2ic5_0;
	wire w_dff_B_ABWPYzyd1_0;
	wire w_dff_B_Clj5FDQq8_0;
	wire w_dff_B_DmpqHqSc8_0;
	wire w_dff_B_J1aLXGbI4_0;
	wire w_dff_B_N8wg7laN4_0;
	wire w_dff_B_GP5vLHyv2_0;
	wire w_dff_B_Be2Ysxib5_0;
	wire w_dff_B_gPsQtPnN3_0;
	wire w_dff_B_A36AN5835_0;
	wire w_dff_B_My5FkOem5_0;
	wire w_dff_B_AErbHNx32_0;
	wire w_dff_B_3lw6lXpq4_0;
	wire w_dff_B_e5kn9bDL4_0;
	wire w_dff_B_WOXC58xL9_0;
	wire w_dff_B_MBNxqEwQ0_0;
	wire w_dff_B_5wamTYmW5_0;
	wire w_dff_B_RdYtaUpK3_0;
	wire w_dff_B_nqSKNmyc3_0;
	wire w_dff_B_7h0FUDYy4_0;
	wire w_dff_B_QRFl5BpH5_0;
	wire w_dff_B_lHKGjeth2_0;
	wire w_dff_B_DzG9wZ8R8_0;
	wire w_dff_B_OetR8HtG3_0;
	wire w_dff_B_QD3eN4qy0_0;
	wire w_dff_B_xcOhM3897_0;
	wire w_dff_B_nsrOx64v5_0;
	wire w_dff_B_Lw4EMmik2_0;
	wire w_dff_B_vaPzb9Lh3_0;
	wire w_dff_B_twdsDPhj4_0;
	wire w_dff_B_2BgPyPxL1_0;
	wire w_dff_B_cdmP6FRm8_0;
	wire w_dff_B_3MLd8POT7_0;
	wire w_dff_B_Q6N4BjUs1_0;
	wire w_dff_B_ZwTS8L4J5_0;
	wire w_dff_B_5eT1uxPd5_0;
	wire w_dff_B_1znjDKfO1_0;
	wire w_dff_B_k7saA5fi9_0;
	wire w_dff_B_ScYLCaw14_0;
	wire w_dff_B_DGImIhA32_0;
	wire w_dff_B_XVsxPe4A7_0;
	wire w_dff_B_ZywCeo2z8_0;
	wire w_dff_B_lWlKqLvt3_0;
	wire w_dff_B_YtYriMyZ3_0;
	wire w_dff_B_IythJWoj7_0;
	wire w_dff_B_2877Msfg5_0;
	wire w_dff_B_JRRpibkr5_0;
	wire w_dff_B_q1Ka5dt06_0;
	wire w_dff_B_LbHYiKyu6_0;
	wire w_dff_B_8K7Rwd960_0;
	wire w_dff_B_UkkkbCyZ2_0;
	wire w_dff_B_V6CDGR0q8_0;
	wire w_dff_B_pTlsvhYO1_0;
	wire w_dff_B_QExLkNpv5_0;
	wire w_dff_B_XiOn47WN8_0;
	wire w_dff_B_l2bArXxB7_0;
	wire w_dff_B_Q93H77K29_0;
	wire w_dff_B_9qSwlpjO1_0;
	wire w_dff_B_x5VFf4df8_0;
	wire w_dff_B_htIWiGFV0_0;
	wire w_dff_B_rp9vt6i54_0;
	wire w_dff_B_qK05uAH65_0;
	wire w_dff_B_PLXBpS6r1_0;
	wire w_dff_B_lW1mhuSE7_0;
	wire w_dff_B_HMySgqvW9_0;
	wire w_dff_B_chQOsgIx4_0;
	wire w_dff_B_Ld72VMUp9_0;
	wire w_dff_B_LAftCvl50_0;
	wire w_dff_B_kagAjCL64_0;
	wire w_dff_B_qjFwTGxP1_1;
	wire w_dff_B_LtZsPGh25_1;
	wire w_dff_B_dW92EnaZ1_1;
	wire w_dff_B_rDobrcMO9_1;
	wire w_dff_B_TaIFXNXn5_1;
	wire w_dff_B_fTXL76RH1_1;
	wire w_dff_B_SWO1VNoZ6_1;
	wire w_dff_B_qtwiTqLc8_1;
	wire w_dff_B_MyLOtbVu5_1;
	wire w_dff_B_iTtCN6C14_1;
	wire w_dff_B_9xGNOBzr6_1;
	wire w_dff_B_TYMDtaDg2_1;
	wire w_dff_B_HpHI2JVg1_1;
	wire w_dff_B_yY55FNfD7_1;
	wire w_dff_B_IqeghPMR8_1;
	wire w_dff_B_keFfFJ6t8_1;
	wire w_dff_B_wsQ3WbNG3_1;
	wire w_dff_B_oboScFUG6_1;
	wire w_dff_B_xe0Kf96f6_1;
	wire w_dff_B_CGzX8wAP5_1;
	wire w_dff_B_ZSzkqT5D6_1;
	wire w_dff_B_LglLR6kE2_1;
	wire w_dff_B_QTPQCk5J0_1;
	wire w_dff_B_c8PZR3jf8_1;
	wire w_dff_B_K09zfacP0_1;
	wire w_dff_B_T5fnkjyI2_1;
	wire w_dff_B_v5OMq2pA1_1;
	wire w_dff_B_C0kMhk337_1;
	wire w_dff_B_7Mvjc0O61_1;
	wire w_dff_B_XM4TILbz7_1;
	wire w_dff_B_QpGGAeox1_1;
	wire w_dff_B_WeuonUrS6_1;
	wire w_dff_B_B7L9MCGb4_1;
	wire w_dff_B_ycXMBjR54_1;
	wire w_dff_B_KAGggqh48_1;
	wire w_dff_B_FoMRjuHa9_1;
	wire w_dff_B_TyMT8Oai1_1;
	wire w_dff_B_QThEvbVe3_1;
	wire w_dff_B_2qV6bWAY7_1;
	wire w_dff_B_QhCdLOFK5_1;
	wire w_dff_B_BlA5O6cd2_1;
	wire w_dff_B_KFzOiraL5_1;
	wire w_dff_B_7JGkfJtD3_1;
	wire w_dff_B_XV0pEo2l3_1;
	wire w_dff_B_LKNlVyBz8_1;
	wire w_dff_B_WNu5eXCK1_1;
	wire w_dff_B_gObKPTmG6_1;
	wire w_dff_B_cNENFW5t7_1;
	wire w_dff_B_0vsjRolz6_1;
	wire w_dff_B_Fxvm5vPZ1_1;
	wire w_dff_B_sFpfKT8X7_1;
	wire w_dff_B_pFdDnQGj7_1;
	wire w_dff_B_GNmagbj10_1;
	wire w_dff_B_VaZwxek65_1;
	wire w_dff_B_T70BR5b65_1;
	wire w_dff_B_nPV2hRap2_1;
	wire w_dff_B_BalEm5O52_1;
	wire w_dff_B_Rhqgx9ps7_1;
	wire w_dff_B_8yRd9DR00_1;
	wire w_dff_B_aiH2UxQ45_1;
	wire w_dff_B_0j3WZ4HX0_1;
	wire w_dff_B_DrP1uDhV9_1;
	wire w_dff_B_txnh3JSb9_1;
	wire w_dff_B_ACmiHmq19_1;
	wire w_dff_B_yiv7h9zv4_1;
	wire w_dff_B_5SoWRpiD4_1;
	wire w_dff_B_MpXvo99k6_1;
	wire w_dff_B_FUFG53Ln1_1;
	wire w_dff_B_cwwQTsWZ7_1;
	wire w_dff_B_UD1By94n0_1;
	wire w_dff_B_O3NfOOfO1_1;
	wire w_dff_B_5Oq74Rxk8_1;
	wire w_dff_B_XsxOnK867_1;
	wire w_dff_B_mN8OCDtM7_1;
	wire w_dff_B_nS57dSDL7_1;
	wire w_dff_B_BmHiU5VO6_1;
	wire w_dff_B_3VNwujLj4_1;
	wire w_dff_B_Q0alDEF74_1;
	wire w_dff_B_sa97GCRl4_1;
	wire w_dff_B_szP7HnQ50_1;
	wire w_dff_B_u3ipOcjU8_1;
	wire w_dff_B_kn1vR85C7_1;
	wire w_dff_B_G7DdSTmA4_1;
	wire w_dff_B_3nYI5KG06_1;
	wire w_dff_B_fBlOQnWp2_1;
	wire w_dff_B_94aJhMqB6_1;
	wire w_dff_B_KHP2p4OH7_1;
	wire w_dff_B_Ytc35zPu3_1;
	wire w_dff_B_JVQ57C7i9_1;
	wire w_dff_B_0s0dPjLj1_1;
	wire w_dff_B_t1GTVvN16_1;
	wire w_dff_B_0chOpwD94_1;
	wire w_dff_B_JawOBCjj5_1;
	wire w_dff_B_U16ejgIK9_1;
	wire w_dff_B_EGczAVq93_1;
	wire w_dff_B_uV8QYM7I5_1;
	wire w_dff_B_0KbJmfYC1_1;
	wire w_dff_B_OScwFDyr0_1;
	wire w_dff_B_j3dgmtwS6_1;
	wire w_dff_B_9LeGDpeM8_1;
	wire w_dff_B_Au9YUNtD6_1;
	wire w_dff_B_iTtZdKQ85_1;
	wire w_dff_B_3SuEsW770_1;
	wire w_dff_B_I7tw9qDa5_1;
	wire w_dff_B_LaZLcbmA8_1;
	wire w_dff_B_PXYmFUcf2_1;
	wire w_dff_B_vqCGRPoq9_1;
	wire w_dff_B_C5nm0R890_1;
	wire w_dff_B_jDEcKhfV6_1;
	wire w_dff_B_vbK5iP3S2_1;
	wire w_dff_B_fF9qNdta0_1;
	wire w_dff_B_fJF763LR9_1;
	wire w_dff_B_130cv7473_1;
	wire w_dff_B_JzjrsjBu9_1;
	wire w_dff_B_mJD14FKk0_1;
	wire w_dff_B_Qux1WfCy1_1;
	wire w_dff_B_YuEZvZoQ4_1;
	wire w_dff_B_N12tJPel7_1;
	wire w_dff_B_VtuFAYEw0_1;
	wire w_dff_B_es37bXV36_1;
	wire w_dff_B_VPzNwCch5_1;
	wire w_dff_B_QoliabzH9_1;
	wire w_dff_B_7vxyjbbi2_1;
	wire w_dff_B_xndqxWZN7_1;
	wire w_dff_B_DkDpKM995_1;
	wire w_dff_B_uZVHTY441_1;
	wire w_dff_B_UIfRMMo17_0;
	wire w_dff_B_sEYm1PnX8_0;
	wire w_dff_B_8KdiZ2Z47_0;
	wire w_dff_B_OIU4Vtun3_0;
	wire w_dff_B_vcMhgbVm8_0;
	wire w_dff_B_BDBknKSh5_0;
	wire w_dff_B_K4cpapNp1_0;
	wire w_dff_B_gh47d6QV4_0;
	wire w_dff_B_gYxJyOCt7_0;
	wire w_dff_B_nQcCXD8u0_0;
	wire w_dff_B_ehj63xts3_0;
	wire w_dff_B_7PaJGfIE5_0;
	wire w_dff_B_NWKKcmph6_0;
	wire w_dff_B_hJuN2ovf5_0;
	wire w_dff_B_SJH1WdSV3_0;
	wire w_dff_B_2OKllxAE7_0;
	wire w_dff_B_TAYlzFfb9_0;
	wire w_dff_B_wE5QgV1g8_0;
	wire w_dff_B_7KhKfUyC7_0;
	wire w_dff_B_HoSP0Or07_0;
	wire w_dff_B_Cn1zECOW4_0;
	wire w_dff_B_GfXPN2PZ0_0;
	wire w_dff_B_tTPtnnub5_0;
	wire w_dff_B_G10VaWMB6_0;
	wire w_dff_B_8T7Deinj5_0;
	wire w_dff_B_Wd5Ui0yN3_0;
	wire w_dff_B_0sixEjbQ6_0;
	wire w_dff_B_GDVSf4dv0_0;
	wire w_dff_B_mKPcTAxu1_0;
	wire w_dff_B_OlPObljC3_0;
	wire w_dff_B_oAcq70lk2_0;
	wire w_dff_B_XkINiefj9_0;
	wire w_dff_B_8bxpsKze5_0;
	wire w_dff_B_SF4PPvlF0_0;
	wire w_dff_B_CbEzOaUY6_0;
	wire w_dff_B_5EOOx0lr4_0;
	wire w_dff_B_A1tBblZP1_0;
	wire w_dff_B_Mat87lFi1_0;
	wire w_dff_B_mcHp6r683_0;
	wire w_dff_B_KU7I6zKP9_0;
	wire w_dff_B_QnzTMJqT8_0;
	wire w_dff_B_NMAoaklK0_0;
	wire w_dff_B_wdNxyA832_0;
	wire w_dff_B_3toypXCa5_0;
	wire w_dff_B_YKASeoiX4_0;
	wire w_dff_B_qAHBOJ486_0;
	wire w_dff_B_pzGJ38Re2_0;
	wire w_dff_B_2exID8Tl9_0;
	wire w_dff_B_Y6E4ZdBX8_0;
	wire w_dff_B_2s67h5uY5_0;
	wire w_dff_B_pbRwGNh50_0;
	wire w_dff_B_ReqN87sL7_0;
	wire w_dff_B_6FhJ5evS2_0;
	wire w_dff_B_3dqMHn1g2_0;
	wire w_dff_B_APLbVDTH9_0;
	wire w_dff_B_lMhO8JRY7_0;
	wire w_dff_B_2jCeuxHF1_0;
	wire w_dff_B_dXUYhB749_0;
	wire w_dff_B_W48yjts62_0;
	wire w_dff_B_p7p98mYh4_0;
	wire w_dff_B_j7c3tMRw0_0;
	wire w_dff_B_p5TH6L823_0;
	wire w_dff_B_6Xmhg7f57_0;
	wire w_dff_B_kT7l4loP3_0;
	wire w_dff_B_J1bnMWc63_0;
	wire w_dff_B_UAfeS6Mu0_0;
	wire w_dff_B_rdW3g0p80_0;
	wire w_dff_B_8m3f4Rrq7_0;
	wire w_dff_B_IOD82zOu5_0;
	wire w_dff_B_0uvycL3x0_0;
	wire w_dff_B_ZBjdw3w07_0;
	wire w_dff_B_oxf2Vwjv0_0;
	wire w_dff_B_DnBCThME5_0;
	wire w_dff_B_FdPlqoNF3_0;
	wire w_dff_B_NMFWkd9N5_0;
	wire w_dff_B_fTphxSUS6_0;
	wire w_dff_B_U7uYyPWd0_0;
	wire w_dff_B_FnDkmIOv6_0;
	wire w_dff_B_IzXv99gG7_0;
	wire w_dff_B_uW34HRL47_0;
	wire w_dff_B_pUcGSPB91_0;
	wire w_dff_B_PYBMFpUb9_0;
	wire w_dff_B_jm6gE8V13_0;
	wire w_dff_B_iF8OvDmU2_0;
	wire w_dff_B_TE85hIov6_0;
	wire w_dff_B_XETMNRd40_0;
	wire w_dff_B_YSZ4SavV4_0;
	wire w_dff_B_lji79BQR2_0;
	wire w_dff_B_gLPIv3Ty4_0;
	wire w_dff_B_ksQmPqfu1_0;
	wire w_dff_B_6x9ub2bx4_0;
	wire w_dff_B_Cl8mEKel8_0;
	wire w_dff_B_A4SJWYP19_0;
	wire w_dff_B_mTnZeH0p7_0;
	wire w_dff_B_fB6MDpEm1_0;
	wire w_dff_B_cqAod1e78_0;
	wire w_dff_B_W8rLN8me8_0;
	wire w_dff_B_PmHIsatk6_0;
	wire w_dff_B_8FhigV8A8_0;
	wire w_dff_B_3CUW0Tyv3_0;
	wire w_dff_B_agaIgjiY5_0;
	wire w_dff_B_5QoASS2s3_0;
	wire w_dff_B_F6829vpX1_0;
	wire w_dff_B_CTLNycMm9_0;
	wire w_dff_B_UkIALfw99_0;
	wire w_dff_B_DEayxWl14_0;
	wire w_dff_B_6i5RghSa5_0;
	wire w_dff_B_e2MUULoz3_0;
	wire w_dff_B_GUJnZhVb8_0;
	wire w_dff_B_qOClIXxQ1_0;
	wire w_dff_B_pllzwnu44_0;
	wire w_dff_B_7vzSVvY71_0;
	wire w_dff_B_RZx1FXN96_0;
	wire w_dff_B_K9G9WEws1_0;
	wire w_dff_B_dlKyWSjy4_0;
	wire w_dff_B_I3zJEqxf4_0;
	wire w_dff_B_bNbjF7No7_0;
	wire w_dff_B_yB78cJMU8_0;
	wire w_dff_B_05sQ1YAL9_0;
	wire w_dff_B_HurN6bGI8_0;
	wire w_dff_B_dXaR3gRJ0_0;
	wire w_dff_B_N9gTvttA7_0;
	wire w_dff_B_lrDVgVsa3_0;
	wire w_dff_B_t6WIj8CJ3_0;
	wire w_dff_B_3yjLCZJr2_0;
	wire w_dff_B_DNEnPLV67_0;
	wire w_dff_B_PeJMRXYm7_1;
	wire w_dff_B_Wiq7zt4W4_1;
	wire w_dff_B_2gazRcPi3_1;
	wire w_dff_B_sT1NyVZW5_1;
	wire w_dff_B_xeKHbRBE2_1;
	wire w_dff_B_MsoxdLTO7_1;
	wire w_dff_B_HA2m0Zgv2_1;
	wire w_dff_B_uZln1uGt9_1;
	wire w_dff_B_TfEDFa7M4_1;
	wire w_dff_B_VBNbnLRv9_1;
	wire w_dff_B_NMbhZqF13_1;
	wire w_dff_B_GRKZgOnA9_1;
	wire w_dff_B_fgWc8n1X0_1;
	wire w_dff_B_Y4Lnimlj8_1;
	wire w_dff_B_dW8iRuQT6_1;
	wire w_dff_B_3SXHIxi50_1;
	wire w_dff_B_tZaEXAva8_1;
	wire w_dff_B_ZYlAkPz61_1;
	wire w_dff_B_cLYFJyYG0_1;
	wire w_dff_B_y5VyVXjM1_1;
	wire w_dff_B_lZ3nBqQK4_1;
	wire w_dff_B_j5JC0dDh6_1;
	wire w_dff_B_dWwtbhsU4_1;
	wire w_dff_B_wQxpwdh25_1;
	wire w_dff_B_c6XBPG3H8_1;
	wire w_dff_B_YP6fwQ929_1;
	wire w_dff_B_ZTkp6LO53_1;
	wire w_dff_B_gXu6JrfR9_1;
	wire w_dff_B_9iLnkI9X5_1;
	wire w_dff_B_yBBxLciN0_1;
	wire w_dff_B_Gz5WVE5l6_1;
	wire w_dff_B_Ce3V9bNW4_1;
	wire w_dff_B_GnAuJlnv8_1;
	wire w_dff_B_ehn53vEQ9_1;
	wire w_dff_B_iiv3RP1D2_1;
	wire w_dff_B_FxNAlomB1_1;
	wire w_dff_B_u2AVdzzZ3_1;
	wire w_dff_B_3sFZ7W2j9_1;
	wire w_dff_B_EXsJSvgH9_1;
	wire w_dff_B_ntYIyMmg4_1;
	wire w_dff_B_Eskgs0l44_1;
	wire w_dff_B_fSiQxdSn4_1;
	wire w_dff_B_r5W895SF3_1;
	wire w_dff_B_B4JZwX4C6_1;
	wire w_dff_B_oI7yG2Ov5_1;
	wire w_dff_B_tw7DQOUz7_1;
	wire w_dff_B_vhFocqyv4_1;
	wire w_dff_B_NkncWFJK2_1;
	wire w_dff_B_rZ8NEeaP6_1;
	wire w_dff_B_OfHGrOCt1_1;
	wire w_dff_B_woq8m1pW8_1;
	wire w_dff_B_lCWMDEcX7_1;
	wire w_dff_B_mxIvtezJ4_1;
	wire w_dff_B_HLDupKPU2_1;
	wire w_dff_B_73FFJ3sa5_1;
	wire w_dff_B_CgV9igpK7_1;
	wire w_dff_B_Cj5fSiLs3_1;
	wire w_dff_B_9AuY64Sa9_1;
	wire w_dff_B_Q8xiu3zP2_1;
	wire w_dff_B_QZGKarUy1_1;
	wire w_dff_B_vClkgFhS3_1;
	wire w_dff_B_YT8xm2Iy4_1;
	wire w_dff_B_TO3BQIx44_1;
	wire w_dff_B_bz3EMpQq3_1;
	wire w_dff_B_moqXD66n7_1;
	wire w_dff_B_b5S2fOyC0_1;
	wire w_dff_B_ok1ZS0Ps8_1;
	wire w_dff_B_MrONCrF44_1;
	wire w_dff_B_kE4BFMRr0_1;
	wire w_dff_B_FgS4MFPD2_1;
	wire w_dff_B_q2OKyHLx5_1;
	wire w_dff_B_6KYO2uzd1_1;
	wire w_dff_B_GR044DAE2_1;
	wire w_dff_B_XcQe7W8l6_1;
	wire w_dff_B_OtRXcKN75_1;
	wire w_dff_B_vOTZvkpf8_1;
	wire w_dff_B_vKoWYKZv4_1;
	wire w_dff_B_djybVx9m5_1;
	wire w_dff_B_8fq1QfUs8_1;
	wire w_dff_B_cCfbTfJ69_1;
	wire w_dff_B_e1CJdju65_1;
	wire w_dff_B_q7oS9qaI6_1;
	wire w_dff_B_5fD5dJ1C8_1;
	wire w_dff_B_vlqhbnTp1_1;
	wire w_dff_B_1baSNXil2_1;
	wire w_dff_B_YyUQP1Yz7_1;
	wire w_dff_B_CgvCYpeL9_1;
	wire w_dff_B_KWmywiR21_1;
	wire w_dff_B_fA0kqpSB9_1;
	wire w_dff_B_jkzuCscJ6_1;
	wire w_dff_B_yP5rpBqu2_1;
	wire w_dff_B_iikdZxSv7_1;
	wire w_dff_B_W0jaPUOG6_1;
	wire w_dff_B_PXAohauM5_1;
	wire w_dff_B_j7qJ5wGm2_1;
	wire w_dff_B_TTGlPZDV5_1;
	wire w_dff_B_ZynYgw6A7_1;
	wire w_dff_B_bmzlTLMw4_1;
	wire w_dff_B_Uh1CetYi7_1;
	wire w_dff_B_LVp9OJPG9_1;
	wire w_dff_B_OTRMn5AT1_1;
	wire w_dff_B_XNx55mJc4_1;
	wire w_dff_B_WCVQQn2Z4_1;
	wire w_dff_B_8xeGuheq1_1;
	wire w_dff_B_8rWM0NSK2_1;
	wire w_dff_B_DpVfeCqn9_1;
	wire w_dff_B_FLooi0u00_1;
	wire w_dff_B_NxsP3JOE5_1;
	wire w_dff_B_xSyMuwPc9_1;
	wire w_dff_B_YPjSjgan5_1;
	wire w_dff_B_zHcoyCFp8_1;
	wire w_dff_B_GY0f20Nd8_1;
	wire w_dff_B_qZte3hRw7_1;
	wire w_dff_B_8PR18gDU6_1;
	wire w_dff_B_GtqqI2B20_1;
	wire w_dff_B_I3zmRXlp5_1;
	wire w_dff_B_qgE89aah3_1;
	wire w_dff_B_nj5brqWu0_1;
	wire w_dff_B_NmWQJAZR7_1;
	wire w_dff_B_yTS1F6IJ9_1;
	wire w_dff_B_ZVxn8VaI5_1;
	wire w_dff_B_zUudwbrL0_1;
	wire w_dff_B_19MZpVs95_1;
	wire w_dff_B_lUBrKJW10_1;
	wire w_dff_B_cdHtn6570_1;
	wire w_dff_B_IMnVun0Q4_0;
	wire w_dff_B_VAjhsi152_0;
	wire w_dff_B_Ixsoupfq3_0;
	wire w_dff_B_EQRSAtTk3_0;
	wire w_dff_B_TLcepq6k1_0;
	wire w_dff_B_fQZLxhSm3_0;
	wire w_dff_B_4uq5uk1e2_0;
	wire w_dff_B_ntVLpPRX3_0;
	wire w_dff_B_z1gylA3Q9_0;
	wire w_dff_B_OrwUJUdw2_0;
	wire w_dff_B_edf8jYCF8_0;
	wire w_dff_B_PnV34B7w1_0;
	wire w_dff_B_8DldS5Cp0_0;
	wire w_dff_B_oW1zYRmF0_0;
	wire w_dff_B_tgWlweE71_0;
	wire w_dff_B_J6Y7qPpE9_0;
	wire w_dff_B_qjzBuBzg3_0;
	wire w_dff_B_oqchZ6051_0;
	wire w_dff_B_V3QrYPJO2_0;
	wire w_dff_B_rjdoaBX81_0;
	wire w_dff_B_zAWkoLjI6_0;
	wire w_dff_B_JsKDRV3C8_0;
	wire w_dff_B_WhF391KJ4_0;
	wire w_dff_B_sB3hWUCX2_0;
	wire w_dff_B_66SgVw1a1_0;
	wire w_dff_B_kZMA0rtj5_0;
	wire w_dff_B_gdCCQYfR3_0;
	wire w_dff_B_4lD30sUO7_0;
	wire w_dff_B_wpCC2XWU0_0;
	wire w_dff_B_F6QzjSia3_0;
	wire w_dff_B_IEIK7X0Y5_0;
	wire w_dff_B_pG3rpEGJ8_0;
	wire w_dff_B_BGA3TmS48_0;
	wire w_dff_B_GU0xIJok8_0;
	wire w_dff_B_FDmijpER7_0;
	wire w_dff_B_7AEMpKiG2_0;
	wire w_dff_B_wJ749GZi2_0;
	wire w_dff_B_Rf01G3uW1_0;
	wire w_dff_B_WMy4NIXB7_0;
	wire w_dff_B_G4MNqFtJ3_0;
	wire w_dff_B_J9bsXzV72_0;
	wire w_dff_B_yX6gfEQc1_0;
	wire w_dff_B_lmlGSbUF3_0;
	wire w_dff_B_tT4OUdiy7_0;
	wire w_dff_B_MPcLLEvy5_0;
	wire w_dff_B_8sGAn65s6_0;
	wire w_dff_B_ZQuoN1vj4_0;
	wire w_dff_B_K7JEPbt00_0;
	wire w_dff_B_sO04ZVAK5_0;
	wire w_dff_B_9bIks27h4_0;
	wire w_dff_B_PGSfgcW68_0;
	wire w_dff_B_86JATPbA0_0;
	wire w_dff_B_QTuAey3s3_0;
	wire w_dff_B_UHWEwQSi7_0;
	wire w_dff_B_OcX2W1w95_0;
	wire w_dff_B_UAiq6hR03_0;
	wire w_dff_B_6ylJCuaV5_0;
	wire w_dff_B_MOSNjWBY3_0;
	wire w_dff_B_w3VS5xRg5_0;
	wire w_dff_B_1NVCE82i5_0;
	wire w_dff_B_8KX8VFWz4_0;
	wire w_dff_B_Cg23HPDG3_0;
	wire w_dff_B_mliKyHbN2_0;
	wire w_dff_B_V1byI0Ol4_0;
	wire w_dff_B_TMNy6PmX6_0;
	wire w_dff_B_Gew0W3Sr4_0;
	wire w_dff_B_a1U805450_0;
	wire w_dff_B_6f6WCIrx7_0;
	wire w_dff_B_vv5kaedV9_0;
	wire w_dff_B_n79wEXfz3_0;
	wire w_dff_B_6uJn5AC98_0;
	wire w_dff_B_o4nmDaC89_0;
	wire w_dff_B_OZuFnDnY0_0;
	wire w_dff_B_JXaLon864_0;
	wire w_dff_B_iOrtRVcg5_0;
	wire w_dff_B_ge1i3KHv5_0;
	wire w_dff_B_vcgDCCJj4_0;
	wire w_dff_B_LOUOG8p22_0;
	wire w_dff_B_MToH7Jdj3_0;
	wire w_dff_B_jHXk46My1_0;
	wire w_dff_B_pDBIaVaB3_0;
	wire w_dff_B_b9itHejq2_0;
	wire w_dff_B_sK6nx3kW4_0;
	wire w_dff_B_0NHkqqYB9_0;
	wire w_dff_B_Vw1HvXim9_0;
	wire w_dff_B_CEp2nxG80_0;
	wire w_dff_B_CQZJfCA03_0;
	wire w_dff_B_ciFCD8mz4_0;
	wire w_dff_B_vSHuAQsA7_0;
	wire w_dff_B_1PWnsKMM0_0;
	wire w_dff_B_VcH6Qt5e8_0;
	wire w_dff_B_ADb1uOCp2_0;
	wire w_dff_B_iVlYBZ2r1_0;
	wire w_dff_B_vjwpUNmO4_0;
	wire w_dff_B_LWLymFrt1_0;
	wire w_dff_B_G8sbiDlD9_0;
	wire w_dff_B_blWbO9755_0;
	wire w_dff_B_u6Rv9ZsP2_0;
	wire w_dff_B_n0eQyWeG0_0;
	wire w_dff_B_kwMRE6wA3_0;
	wire w_dff_B_FWLe1q7S2_0;
	wire w_dff_B_1ugbiaKb4_0;
	wire w_dff_B_cm9WZrdO1_0;
	wire w_dff_B_CbHCSJUA3_0;
	wire w_dff_B_DTokUmuG5_0;
	wire w_dff_B_0vreo1EL3_0;
	wire w_dff_B_cRzaImJV4_0;
	wire w_dff_B_A2ESqh3h9_0;
	wire w_dff_B_YrV7BLld1_0;
	wire w_dff_B_lJAXRhCf6_0;
	wire w_dff_B_OkhOkxN08_0;
	wire w_dff_B_DzyeuD2h9_0;
	wire w_dff_B_aMON1cWP4_0;
	wire w_dff_B_zdX2rrMt1_0;
	wire w_dff_B_JNK6Lsyf7_0;
	wire w_dff_B_Roaq9tY26_0;
	wire w_dff_B_pUvYqRzk6_0;
	wire w_dff_B_o4kFetsG5_0;
	wire w_dff_B_fTvzuKQH5_0;
	wire w_dff_B_bDPP2thR9_0;
	wire w_dff_B_s4dAHRDt0_0;
	wire w_dff_B_c2ue1IU29_0;
	wire w_dff_B_sfOAAu5Y1_0;
	wire w_dff_B_Q63QvkbE0_0;
	wire w_dff_B_B43o3NKK2_0;
	wire w_dff_B_oqYIPTeU4_1;
	wire w_dff_B_tczRxsH46_1;
	wire w_dff_B_94Gh0IAv1_1;
	wire w_dff_B_XvVnduTm9_1;
	wire w_dff_B_rNTs7xoz3_1;
	wire w_dff_B_6JR2JrYa2_1;
	wire w_dff_B_sQjGRBF71_1;
	wire w_dff_B_EDAuk2Xe2_1;
	wire w_dff_B_FgnK8xl14_1;
	wire w_dff_B_uBHNsLnf1_1;
	wire w_dff_B_INXEK2Sg7_1;
	wire w_dff_B_GmlP5Xla5_1;
	wire w_dff_B_MnxEDMVB5_1;
	wire w_dff_B_MTCX9mng9_1;
	wire w_dff_B_qYZaejB08_1;
	wire w_dff_B_cMZ91g1w8_1;
	wire w_dff_B_oMOrSPYN7_1;
	wire w_dff_B_BXYP1xeg3_1;
	wire w_dff_B_AHH63meh4_1;
	wire w_dff_B_d9kr3czF9_1;
	wire w_dff_B_UtVzCpwt7_1;
	wire w_dff_B_0WpDxjBa2_1;
	wire w_dff_B_ZcROiVMY9_1;
	wire w_dff_B_ufTqqo5U5_1;
	wire w_dff_B_CDvLvOWq8_1;
	wire w_dff_B_nvs7VNKf2_1;
	wire w_dff_B_FplUPSm90_1;
	wire w_dff_B_MahhnMRB5_1;
	wire w_dff_B_DFKLVSkq8_1;
	wire w_dff_B_txR1o5Zc9_1;
	wire w_dff_B_fyi9rg8v3_1;
	wire w_dff_B_LV0zw84p6_1;
	wire w_dff_B_FWEQGw1X9_1;
	wire w_dff_B_ZxzevGlQ1_1;
	wire w_dff_B_9ql3iZh97_1;
	wire w_dff_B_XVc5QF827_1;
	wire w_dff_B_fjNElSGi8_1;
	wire w_dff_B_vsWrkZtp1_1;
	wire w_dff_B_X9CsLi1a8_1;
	wire w_dff_B_hKtTLNWx7_1;
	wire w_dff_B_WPMBjTXD5_1;
	wire w_dff_B_ybwBwObn5_1;
	wire w_dff_B_dG6QAN7L1_1;
	wire w_dff_B_PUCooeSz0_1;
	wire w_dff_B_1jMSfx4V9_1;
	wire w_dff_B_j0u58wpI3_1;
	wire w_dff_B_w58al6FC3_1;
	wire w_dff_B_SmpS2Qz92_1;
	wire w_dff_B_ETZ2rAul2_1;
	wire w_dff_B_akscmYcW3_1;
	wire w_dff_B_b6lpjkdW7_1;
	wire w_dff_B_7jBWCWQc8_1;
	wire w_dff_B_1MyMxmme0_1;
	wire w_dff_B_A48oSovy9_1;
	wire w_dff_B_f3QWxPvS1_1;
	wire w_dff_B_FdaaEdc90_1;
	wire w_dff_B_WX9EqciO9_1;
	wire w_dff_B_JlDiXBcc5_1;
	wire w_dff_B_uJZLxMzu9_1;
	wire w_dff_B_ewjeKkt57_1;
	wire w_dff_B_zNb99BgK9_1;
	wire w_dff_B_yCb8gJMo4_1;
	wire w_dff_B_GwhiUGWz6_1;
	wire w_dff_B_PyafcMaX9_1;
	wire w_dff_B_1NTTxpba1_1;
	wire w_dff_B_TmiynQBN1_1;
	wire w_dff_B_ZCOOpv8o9_1;
	wire w_dff_B_W6zwAjlI8_1;
	wire w_dff_B_7T53m27X3_1;
	wire w_dff_B_JgzDgTE35_1;
	wire w_dff_B_voazf92t0_1;
	wire w_dff_B_tpLLy3Nz5_1;
	wire w_dff_B_yqCccnhz8_1;
	wire w_dff_B_dNhs6sjE3_1;
	wire w_dff_B_qs6ENmwM9_1;
	wire w_dff_B_FTFsp5691_1;
	wire w_dff_B_YgFGocW31_1;
	wire w_dff_B_alByZtzp2_1;
	wire w_dff_B_IRMbgUJC1_1;
	wire w_dff_B_v9XqOznu2_1;
	wire w_dff_B_0n6r3ASl7_1;
	wire w_dff_B_z25WlsvQ2_1;
	wire w_dff_B_pnGvleuN1_1;
	wire w_dff_B_diEdI7F51_1;
	wire w_dff_B_ZNS5qQJ09_1;
	wire w_dff_B_FIuPFV7o8_1;
	wire w_dff_B_nrVoCE1H5_1;
	wire w_dff_B_0DsO1CXd1_1;
	wire w_dff_B_YUEfFZ5L7_1;
	wire w_dff_B_v2mJS4Ls8_1;
	wire w_dff_B_wtPgOPWs2_1;
	wire w_dff_B_9ALlXqTx1_1;
	wire w_dff_B_G452Aqi41_1;
	wire w_dff_B_RMo9ksG02_1;
	wire w_dff_B_PvgHgzWU1_1;
	wire w_dff_B_p1QddroD8_1;
	wire w_dff_B_RS4PnBFr1_1;
	wire w_dff_B_33mC7kB02_1;
	wire w_dff_B_1NxulKpu3_1;
	wire w_dff_B_ONvdAm0F7_1;
	wire w_dff_B_LYWOGmNa2_1;
	wire w_dff_B_umajNF3R8_1;
	wire w_dff_B_VeU5RgRJ8_1;
	wire w_dff_B_s8eJBhyK0_1;
	wire w_dff_B_UWk2V1Pd2_1;
	wire w_dff_B_5evCLscw5_1;
	wire w_dff_B_T1nghpIG3_1;
	wire w_dff_B_e1tHOO0X9_1;
	wire w_dff_B_5bCn8Jlu3_1;
	wire w_dff_B_xE3dXEMe3_1;
	wire w_dff_B_peXNoHOm5_1;
	wire w_dff_B_9YhTGdo50_1;
	wire w_dff_B_ZJIp1DiE6_1;
	wire w_dff_B_Ro3hG1000_1;
	wire w_dff_B_IOCsQ4RV2_1;
	wire w_dff_B_604l9mpP4_1;
	wire w_dff_B_UO7xfXY45_1;
	wire w_dff_B_beTjcDsf8_1;
	wire w_dff_B_6TPkIcMj8_1;
	wire w_dff_B_dHP4styR0_1;
	wire w_dff_B_PKoAfIOJ3_1;
	wire w_dff_B_BiApeeNs4_1;
	wire w_dff_B_tBVIKrr45_1;
	wire w_dff_B_WOhTpZP77_1;
	wire w_dff_B_w2UCqheB3_0;
	wire w_dff_B_HpGTHQgg6_0;
	wire w_dff_B_CvmUCDRx5_0;
	wire w_dff_B_AujreAjX9_0;
	wire w_dff_B_R1Cc6msq6_0;
	wire w_dff_B_Xegf7MA70_0;
	wire w_dff_B_bxDlTe5U9_0;
	wire w_dff_B_ORPkQi6C5_0;
	wire w_dff_B_uufp58WE3_0;
	wire w_dff_B_DPYAbrse2_0;
	wire w_dff_B_jiF5o9EO0_0;
	wire w_dff_B_CgGeWtOV6_0;
	wire w_dff_B_u4tJx7aG3_0;
	wire w_dff_B_0GuDs4pM9_0;
	wire w_dff_B_UYsi4ikq6_0;
	wire w_dff_B_2MQqjAKP6_0;
	wire w_dff_B_Nwen2Gf48_0;
	wire w_dff_B_Oc2ksfoM5_0;
	wire w_dff_B_DEh6uNc78_0;
	wire w_dff_B_0bHlZmKc5_0;
	wire w_dff_B_i1XNPAwE8_0;
	wire w_dff_B_hasKDMsR0_0;
	wire w_dff_B_DEsPVo3N8_0;
	wire w_dff_B_HVt6udWA8_0;
	wire w_dff_B_NESNjduk9_0;
	wire w_dff_B_AMT9FJqQ7_0;
	wire w_dff_B_KnOO89J35_0;
	wire w_dff_B_2uodiFBb9_0;
	wire w_dff_B_GLG2pbkc1_0;
	wire w_dff_B_Bk5mbJEd8_0;
	wire w_dff_B_uioYmElR4_0;
	wire w_dff_B_gwao8SRb2_0;
	wire w_dff_B_NXEfhIWO4_0;
	wire w_dff_B_I6JWxblv6_0;
	wire w_dff_B_P1MrBnLi0_0;
	wire w_dff_B_rn3dF23u3_0;
	wire w_dff_B_fHEgJ9xt0_0;
	wire w_dff_B_WvEAAH396_0;
	wire w_dff_B_Or6unfsz9_0;
	wire w_dff_B_ZQ79dYv42_0;
	wire w_dff_B_VgMkRi0F4_0;
	wire w_dff_B_c1la2naF7_0;
	wire w_dff_B_8BlCHmGs9_0;
	wire w_dff_B_RTuFv2jB9_0;
	wire w_dff_B_NMI6u2Vm1_0;
	wire w_dff_B_bA1aj1Ja5_0;
	wire w_dff_B_mzhRBYUq3_0;
	wire w_dff_B_H5VpTsS30_0;
	wire w_dff_B_bxObI4uX7_0;
	wire w_dff_B_RK0TCsYA3_0;
	wire w_dff_B_eqjkK41L5_0;
	wire w_dff_B_n171pwKy9_0;
	wire w_dff_B_kYJw0nya1_0;
	wire w_dff_B_Vku1k3N08_0;
	wire w_dff_B_6k4dRwQa8_0;
	wire w_dff_B_I7H3BmAH6_0;
	wire w_dff_B_zsz0bKgE1_0;
	wire w_dff_B_4k8l3izr5_0;
	wire w_dff_B_5SfkRjzQ9_0;
	wire w_dff_B_aRzmjmHw2_0;
	wire w_dff_B_YBWHNTm40_0;
	wire w_dff_B_3YExAsal2_0;
	wire w_dff_B_cTy98Or30_0;
	wire w_dff_B_jXru8UAN5_0;
	wire w_dff_B_j4fPjshF6_0;
	wire w_dff_B_BcVUBeY14_0;
	wire w_dff_B_nodnidlk9_0;
	wire w_dff_B_Mo6z9htM5_0;
	wire w_dff_B_5lfFUUGb7_0;
	wire w_dff_B_HNKWwTdp5_0;
	wire w_dff_B_tgMHmLvg7_0;
	wire w_dff_B_yGx9XO0y1_0;
	wire w_dff_B_7wOukHDP7_0;
	wire w_dff_B_3mCMrSM53_0;
	wire w_dff_B_EjhPv0Ue1_0;
	wire w_dff_B_586AmrHn1_0;
	wire w_dff_B_sVeiOpTv3_0;
	wire w_dff_B_mHJk5P6P4_0;
	wire w_dff_B_SQy7amcp8_0;
	wire w_dff_B_JqvLh42k3_0;
	wire w_dff_B_kvx9Yotb4_0;
	wire w_dff_B_lvO8LczQ8_0;
	wire w_dff_B_iXWmVun97_0;
	wire w_dff_B_mQHMMDY13_0;
	wire w_dff_B_VeaFra8e0_0;
	wire w_dff_B_1oDJRiut2_0;
	wire w_dff_B_JOP3wQKt7_0;
	wire w_dff_B_QO7hosX06_0;
	wire w_dff_B_30HJfyvr3_0;
	wire w_dff_B_t5TBYdXg2_0;
	wire w_dff_B_hiulta0n9_0;
	wire w_dff_B_a0ANJVWH8_0;
	wire w_dff_B_eQDhJaQr8_0;
	wire w_dff_B_jblAHUSy8_0;
	wire w_dff_B_TeqD7gin4_0;
	wire w_dff_B_h49672xp6_0;
	wire w_dff_B_RPfYOhkB3_0;
	wire w_dff_B_NGWKogmw0_0;
	wire w_dff_B_Wk4KetGe0_0;
	wire w_dff_B_uTflJdG17_0;
	wire w_dff_B_UXItrIjW6_0;
	wire w_dff_B_EOLcdZNy0_0;
	wire w_dff_B_WiSVbLIf7_0;
	wire w_dff_B_YSwUJrZg9_0;
	wire w_dff_B_NDXc5CgD3_0;
	wire w_dff_B_oQb1CUJZ6_0;
	wire w_dff_B_yTiXYGqt9_0;
	wire w_dff_B_7QWeiGtI1_0;
	wire w_dff_B_zVUTpR733_0;
	wire w_dff_B_ErcSPY5p9_0;
	wire w_dff_B_Lso0hCi86_0;
	wire w_dff_B_oj9BPdGt0_0;
	wire w_dff_B_pETxBHAB6_0;
	wire w_dff_B_9oeEatje8_0;
	wire w_dff_B_CDVe9Lni1_0;
	wire w_dff_B_5AJeGuG53_0;
	wire w_dff_B_mD9JOMR65_0;
	wire w_dff_B_tAMSHKno7_0;
	wire w_dff_B_FE4voPy93_0;
	wire w_dff_B_3BlTFiyi6_0;
	wire w_dff_B_qlKuB7PC5_0;
	wire w_dff_B_w0Xu8MMm0_0;
	wire w_dff_B_yYEBiORo3_0;
	wire w_dff_B_niFMbCQe5_0;
	wire w_dff_B_xlvf58vQ1_1;
	wire w_dff_B_TTyx2DR68_1;
	wire w_dff_B_adBEQpWH4_1;
	wire w_dff_B_T9SsQlCm4_1;
	wire w_dff_B_YZTMGZrP2_1;
	wire w_dff_B_aqGz3X2U2_1;
	wire w_dff_B_1T0xIEXj0_1;
	wire w_dff_B_j4Qr55xX6_1;
	wire w_dff_B_X9ys2ipn3_1;
	wire w_dff_B_MZTRSDSN5_1;
	wire w_dff_B_wKjbdVkK8_1;
	wire w_dff_B_K65fyst61_1;
	wire w_dff_B_naMSC7bd7_1;
	wire w_dff_B_mFpoFg8w0_1;
	wire w_dff_B_ZNTO9vlu6_1;
	wire w_dff_B_JiBjjnmS5_1;
	wire w_dff_B_PGJdhn066_1;
	wire w_dff_B_g9jBuuxl1_1;
	wire w_dff_B_IORxOFa64_1;
	wire w_dff_B_EkBj8YK36_1;
	wire w_dff_B_JlYTub2w1_1;
	wire w_dff_B_tTXzqfwP3_1;
	wire w_dff_B_YCcPspPj9_1;
	wire w_dff_B_anQ1ieDQ0_1;
	wire w_dff_B_zHkaOqPY2_1;
	wire w_dff_B_xcwH6Zn87_1;
	wire w_dff_B_qRV4VmrB4_1;
	wire w_dff_B_7AeT5CL99_1;
	wire w_dff_B_wnJwFzY71_1;
	wire w_dff_B_Eli4ENS49_1;
	wire w_dff_B_8z4rXfXo1_1;
	wire w_dff_B_Q71ONbxz9_1;
	wire w_dff_B_so9NQCV50_1;
	wire w_dff_B_qF4M63Kt9_1;
	wire w_dff_B_WRQBdW015_1;
	wire w_dff_B_dpIq37uP5_1;
	wire w_dff_B_n7rxVgFO2_1;
	wire w_dff_B_EKVtwnh58_1;
	wire w_dff_B_RlNahTF76_1;
	wire w_dff_B_J8BvEfSI5_1;
	wire w_dff_B_MyWIFJO38_1;
	wire w_dff_B_nr4Ulwcs3_1;
	wire w_dff_B_CD4EsmfM2_1;
	wire w_dff_B_VZOseP6H2_1;
	wire w_dff_B_xH6WR0Bc1_1;
	wire w_dff_B_PXmMgz7r5_1;
	wire w_dff_B_B8ucmhgy9_1;
	wire w_dff_B_kSGBWEoK7_1;
	wire w_dff_B_8FwmaDCC8_1;
	wire w_dff_B_yHBsplJU6_1;
	wire w_dff_B_lEUKQ5Jh8_1;
	wire w_dff_B_GfxfQfyG5_1;
	wire w_dff_B_8nnEb4cf0_1;
	wire w_dff_B_0pJFpHVi2_1;
	wire w_dff_B_V243fT3F8_1;
	wire w_dff_B_H85nIkPZ7_1;
	wire w_dff_B_mBuljhDl0_1;
	wire w_dff_B_EPJKOdEc2_1;
	wire w_dff_B_25L9GQSA6_1;
	wire w_dff_B_35sVY74G7_1;
	wire w_dff_B_YzfdV7da7_1;
	wire w_dff_B_md59xA725_1;
	wire w_dff_B_U6lud0nQ2_1;
	wire w_dff_B_Q0IpHpA16_1;
	wire w_dff_B_hDsqDcpX3_1;
	wire w_dff_B_56ZfvXFK9_1;
	wire w_dff_B_cbNCLpXx7_1;
	wire w_dff_B_wiLcXbuD1_1;
	wire w_dff_B_wOYgkfWA2_1;
	wire w_dff_B_VenL9k034_1;
	wire w_dff_B_adRC1Spb7_1;
	wire w_dff_B_HWwsSvMW8_1;
	wire w_dff_B_yH7bPvti5_1;
	wire w_dff_B_teslDa011_1;
	wire w_dff_B_z5Xic96G8_1;
	wire w_dff_B_ZdRgUDh58_1;
	wire w_dff_B_YOC3YxSe5_1;
	wire w_dff_B_9Oysk1De1_1;
	wire w_dff_B_svYgorby7_1;
	wire w_dff_B_orUwcZHc5_1;
	wire w_dff_B_bZOTdtDJ1_1;
	wire w_dff_B_E0o0jsJD4_1;
	wire w_dff_B_7Xb5Yn1W7_1;
	wire w_dff_B_qfEGJUMP1_1;
	wire w_dff_B_uaPWsuno6_1;
	wire w_dff_B_PTdKFq1Z2_1;
	wire w_dff_B_sE6Z9dCs6_1;
	wire w_dff_B_vvcFx5Je0_1;
	wire w_dff_B_SLYAROsV1_1;
	wire w_dff_B_meIXkeyV2_1;
	wire w_dff_B_A7VceNDg4_1;
	wire w_dff_B_GzoORZZi1_1;
	wire w_dff_B_n6pIe9V38_1;
	wire w_dff_B_mlFwG6D14_1;
	wire w_dff_B_UVzWyeGm8_1;
	wire w_dff_B_i0Hw55dn2_1;
	wire w_dff_B_1K9eH9dv7_1;
	wire w_dff_B_XjxpKpjw4_1;
	wire w_dff_B_9QPXdl4i0_1;
	wire w_dff_B_NocTdLFw2_1;
	wire w_dff_B_tmehyRQF0_1;
	wire w_dff_B_jvRcFlPW4_1;
	wire w_dff_B_GpQlljSz4_1;
	wire w_dff_B_DJBJuvdo1_1;
	wire w_dff_B_RVAyDpQT0_1;
	wire w_dff_B_6tPjsgCX7_1;
	wire w_dff_B_F9qXrrgj8_1;
	wire w_dff_B_rjefnjaQ8_1;
	wire w_dff_B_gFjkcwoc6_1;
	wire w_dff_B_QTmH9Rgb2_1;
	wire w_dff_B_FNn87wEo1_1;
	wire w_dff_B_0wPVGqB70_1;
	wire w_dff_B_wyrOMR8X2_1;
	wire w_dff_B_0ShiLpUC5_1;
	wire w_dff_B_CPSFP8od5_1;
	wire w_dff_B_XFU1OhDk3_1;
	wire w_dff_B_7EmC7Be77_1;
	wire w_dff_B_5lYm1sbU4_1;
	wire w_dff_B_T057vtT76_1;
	wire w_dff_B_v0qgbIni3_1;
	wire w_dff_B_OXDQLYQM0_1;
	wire w_dff_B_R2r5urwW2_1;
	wire w_dff_B_LkmyUViD3_1;
	wire w_dff_B_ihlUGtXO8_0;
	wire w_dff_B_NkOGzgBJ9_0;
	wire w_dff_B_p09xVsVY1_0;
	wire w_dff_B_0x2a8bzk6_0;
	wire w_dff_B_2D9RksV12_0;
	wire w_dff_B_Jl3mnOkw2_0;
	wire w_dff_B_XjypEmla5_0;
	wire w_dff_B_tKy7lzpq7_0;
	wire w_dff_B_83FZHCaX8_0;
	wire w_dff_B_5bmOblIn6_0;
	wire w_dff_B_nYDAu46E0_0;
	wire w_dff_B_IoIH5eRg8_0;
	wire w_dff_B_sVYv0QnC7_0;
	wire w_dff_B_rLBMJeiD5_0;
	wire w_dff_B_FQUOScfA3_0;
	wire w_dff_B_s0pUiaCh4_0;
	wire w_dff_B_wUX6OwdT6_0;
	wire w_dff_B_mBlZF68n9_0;
	wire w_dff_B_xqzbBVX38_0;
	wire w_dff_B_0I10pM2n0_0;
	wire w_dff_B_mhdMjQlu8_0;
	wire w_dff_B_a4Wax3J05_0;
	wire w_dff_B_tTbJZN4b2_0;
	wire w_dff_B_5grlECEy6_0;
	wire w_dff_B_9ahz7QzT3_0;
	wire w_dff_B_qpkKpWaP2_0;
	wire w_dff_B_vEA4YN229_0;
	wire w_dff_B_SfiivDl58_0;
	wire w_dff_B_XhnCNJfe9_0;
	wire w_dff_B_Yae4X7aV0_0;
	wire w_dff_B_Lmsr50hD4_0;
	wire w_dff_B_o0rAgbcO7_0;
	wire w_dff_B_sMgtRZuH6_0;
	wire w_dff_B_BwpORKUs8_0;
	wire w_dff_B_1Ba3HmeU4_0;
	wire w_dff_B_Tqt3ylUe4_0;
	wire w_dff_B_O4Aey8852_0;
	wire w_dff_B_OaP1z9Xp8_0;
	wire w_dff_B_s9IXb4lF0_0;
	wire w_dff_B_Y4AE17Yg8_0;
	wire w_dff_B_zj0fm7Vz6_0;
	wire w_dff_B_TtMNznxo2_0;
	wire w_dff_B_LIHsrAjx8_0;
	wire w_dff_B_VzGHiERh0_0;
	wire w_dff_B_7h1ZVCIE7_0;
	wire w_dff_B_63WDjKph8_0;
	wire w_dff_B_OFGWtzhD9_0;
	wire w_dff_B_x9UyrlZa1_0;
	wire w_dff_B_MjH3lbxJ4_0;
	wire w_dff_B_k478VyFo3_0;
	wire w_dff_B_qz2r93Fu4_0;
	wire w_dff_B_69GanfH85_0;
	wire w_dff_B_lEHpw3uC9_0;
	wire w_dff_B_MBR4Bqag1_0;
	wire w_dff_B_uMesbX2l8_0;
	wire w_dff_B_lcmLEtLN4_0;
	wire w_dff_B_1cJYQPYZ4_0;
	wire w_dff_B_lbqFqpCt7_0;
	wire w_dff_B_voKNSnEL7_0;
	wire w_dff_B_MeW3wqjq1_0;
	wire w_dff_B_Zr6U3pSh6_0;
	wire w_dff_B_ZpdeBxHt9_0;
	wire w_dff_B_JNmQcTox4_0;
	wire w_dff_B_wccacKVF9_0;
	wire w_dff_B_kj4qZUcD2_0;
	wire w_dff_B_87nUqp621_0;
	wire w_dff_B_tg6XyGZ03_0;
	wire w_dff_B_SHyb2bd79_0;
	wire w_dff_B_Yt7Y0Cxy4_0;
	wire w_dff_B_rfBshHXY2_0;
	wire w_dff_B_Mr0V7Xre1_0;
	wire w_dff_B_NDj991vz6_0;
	wire w_dff_B_dGrQ0FDj8_0;
	wire w_dff_B_E5uY0JtH1_0;
	wire w_dff_B_ylzSd0Ly2_0;
	wire w_dff_B_PJUHQmdO7_0;
	wire w_dff_B_timsz4Qi5_0;
	wire w_dff_B_DHMhyWsv2_0;
	wire w_dff_B_MWCuFCjn1_0;
	wire w_dff_B_hqSiKuxP5_0;
	wire w_dff_B_ASvLsKR52_0;
	wire w_dff_B_4EYPuryV6_0;
	wire w_dff_B_bfXD3M9V8_0;
	wire w_dff_B_E8z8KThg7_0;
	wire w_dff_B_ARYa9xKC7_0;
	wire w_dff_B_XnBYhEer7_0;
	wire w_dff_B_39n8ryt86_0;
	wire w_dff_B_mFbzyEFd7_0;
	wire w_dff_B_mPsRocZH1_0;
	wire w_dff_B_H2ouOVSo6_0;
	wire w_dff_B_zqeayftb6_0;
	wire w_dff_B_1OcOLfLf1_0;
	wire w_dff_B_hLBaU4Vj8_0;
	wire w_dff_B_FSI0gpRE5_0;
	wire w_dff_B_QyQe0UJL1_0;
	wire w_dff_B_GPWikoaz1_0;
	wire w_dff_B_WA7ccQy34_0;
	wire w_dff_B_DiQtJIPr7_0;
	wire w_dff_B_wYuGZ2Ig5_0;
	wire w_dff_B_LEg1aN8I1_0;
	wire w_dff_B_OkPLZWAi8_0;
	wire w_dff_B_DufBxwSX9_0;
	wire w_dff_B_70nLApIG0_0;
	wire w_dff_B_TX9Xt2la9_0;
	wire w_dff_B_GapYUI1h5_0;
	wire w_dff_B_9svg7rmL1_0;
	wire w_dff_B_tWWdQgtJ4_0;
	wire w_dff_B_0CQMMybI4_0;
	wire w_dff_B_cYfT9H400_0;
	wire w_dff_B_aqla3uee8_0;
	wire w_dff_B_Idkb6SYB6_0;
	wire w_dff_B_se6qxCOK7_0;
	wire w_dff_B_a1OSw7zZ0_0;
	wire w_dff_B_O6ZXWT2t0_0;
	wire w_dff_B_4rJmYiWA4_0;
	wire w_dff_B_JXHIGKBh9_0;
	wire w_dff_B_zTMJ1CSA8_0;
	wire w_dff_B_r5wJPKfA1_0;
	wire w_dff_B_T0elTxmH8_0;
	wire w_dff_B_RHjZapdP3_0;
	wire w_dff_B_ziihU3C56_0;
	wire w_dff_B_kb0qb4o00_0;
	wire w_dff_B_oY8pBb783_0;
	wire w_dff_B_z01nDMwv4_1;
	wire w_dff_B_6EtclvnV9_1;
	wire w_dff_B_ZBcu8scr0_1;
	wire w_dff_B_LqkFspZw1_1;
	wire w_dff_B_tXP1X49f7_1;
	wire w_dff_B_eCcyG9jT8_1;
	wire w_dff_B_Uv9PxNtF9_1;
	wire w_dff_B_HpBrX3Se1_1;
	wire w_dff_B_MRgkquuw9_1;
	wire w_dff_B_HOA0lw9V2_1;
	wire w_dff_B_ONoDfZCu1_1;
	wire w_dff_B_MEYCNacy8_1;
	wire w_dff_B_WPOUJTJr9_1;
	wire w_dff_B_ppgNypcU2_1;
	wire w_dff_B_AVKslCmw2_1;
	wire w_dff_B_TgzzxENF2_1;
	wire w_dff_B_3PUyYZIX2_1;
	wire w_dff_B_DNpmCXYj4_1;
	wire w_dff_B_67KCkxOw9_1;
	wire w_dff_B_CUHpFrCa8_1;
	wire w_dff_B_zmYC0MD74_1;
	wire w_dff_B_gmcrlBtl9_1;
	wire w_dff_B_NesNbuze8_1;
	wire w_dff_B_cIPg8KD27_1;
	wire w_dff_B_2JZ92O8j0_1;
	wire w_dff_B_fVztKYZX7_1;
	wire w_dff_B_IzdbYgxG7_1;
	wire w_dff_B_1hjlMMYl6_1;
	wire w_dff_B_GLxaCAdr4_1;
	wire w_dff_B_MsmGbAwv0_1;
	wire w_dff_B_olb9qy8G0_1;
	wire w_dff_B_sBQ2Plh99_1;
	wire w_dff_B_sUg2zMX23_1;
	wire w_dff_B_M4JPRDYr3_1;
	wire w_dff_B_C4vEU0F57_1;
	wire w_dff_B_pBcnD1kN2_1;
	wire w_dff_B_YpoTIwnV5_1;
	wire w_dff_B_ecaywQ3W4_1;
	wire w_dff_B_SNpKsaVS6_1;
	wire w_dff_B_xDU3utD33_1;
	wire w_dff_B_IOoVO09q8_1;
	wire w_dff_B_r7OxnRq26_1;
	wire w_dff_B_ncp8gaxD0_1;
	wire w_dff_B_5AKjTN8n2_1;
	wire w_dff_B_KUJBXrMG0_1;
	wire w_dff_B_YREIpQpD8_1;
	wire w_dff_B_t3AX2Ue72_1;
	wire w_dff_B_la8TEb3D4_1;
	wire w_dff_B_xjVI8tzM6_1;
	wire w_dff_B_kkNod70o8_1;
	wire w_dff_B_bmzszsJ56_1;
	wire w_dff_B_o6lofO308_1;
	wire w_dff_B_kYVXWfTh4_1;
	wire w_dff_B_vLlqJdbV1_1;
	wire w_dff_B_K7P2meAE5_1;
	wire w_dff_B_XAzC2BvG2_1;
	wire w_dff_B_ip7Lp4sn8_1;
	wire w_dff_B_0OQMVJdH3_1;
	wire w_dff_B_anGpywdC9_1;
	wire w_dff_B_6oxiMOGB8_1;
	wire w_dff_B_NGvF5hsp6_1;
	wire w_dff_B_DHufxwt50_1;
	wire w_dff_B_rotnroWx9_1;
	wire w_dff_B_6vbS29bj1_1;
	wire w_dff_B_Jw6tLjP76_1;
	wire w_dff_B_oZMBEcqh6_1;
	wire w_dff_B_jTWHkSJH5_1;
	wire w_dff_B_6FxYUHsi9_1;
	wire w_dff_B_IlitXWrR5_1;
	wire w_dff_B_CKCoXO692_1;
	wire w_dff_B_SNgoNgaX4_1;
	wire w_dff_B_eriyZy030_1;
	wire w_dff_B_wNtVVCzX3_1;
	wire w_dff_B_KVFVZLHq7_1;
	wire w_dff_B_8KVgezxO5_1;
	wire w_dff_B_gFiwlnzb6_1;
	wire w_dff_B_sNmxpQxx6_1;
	wire w_dff_B_924ILho16_1;
	wire w_dff_B_9LdlSj4V6_1;
	wire w_dff_B_DFKto3wA5_1;
	wire w_dff_B_UWXbKLbW8_1;
	wire w_dff_B_trU4JIUl8_1;
	wire w_dff_B_Knj0R4De6_1;
	wire w_dff_B_yNA9Lu6y2_1;
	wire w_dff_B_4lLcYCez9_1;
	wire w_dff_B_HuepJOaS9_1;
	wire w_dff_B_2BHqe7X89_1;
	wire w_dff_B_itN1NFKy7_1;
	wire w_dff_B_oSek1iaI0_1;
	wire w_dff_B_YMziUT3Y2_1;
	wire w_dff_B_3rqvSSHv2_1;
	wire w_dff_B_ttCYVUMl4_1;
	wire w_dff_B_HD3rvZxt5_1;
	wire w_dff_B_zmpdtUQ97_1;
	wire w_dff_B_rManAGOy5_1;
	wire w_dff_B_UEUloay98_1;
	wire w_dff_B_SpQZ42fl5_1;
	wire w_dff_B_SeLCNm5T1_1;
	wire w_dff_B_jMmJiZJx6_1;
	wire w_dff_B_bNTJcCDt2_1;
	wire w_dff_B_6BHKAgrd5_1;
	wire w_dff_B_jxo5zOz77_1;
	wire w_dff_B_lbhvHxMg9_1;
	wire w_dff_B_xqOVZdHf7_1;
	wire w_dff_B_Jgzy3lKO9_1;
	wire w_dff_B_AJU9a7Vx9_1;
	wire w_dff_B_gS8sz9dN8_1;
	wire w_dff_B_uyZpVk0P3_1;
	wire w_dff_B_xGhH23sQ3_1;
	wire w_dff_B_nUbtSo662_1;
	wire w_dff_B_lx2Ms7HH6_1;
	wire w_dff_B_aTskClIk1_1;
	wire w_dff_B_q4H6WhDe7_1;
	wire w_dff_B_ac2BNYvd5_1;
	wire w_dff_B_P3pcQVXZ3_1;
	wire w_dff_B_qTfinytC8_1;
	wire w_dff_B_T4KtDsWT1_1;
	wire w_dff_B_Jt2yUwxU0_1;
	wire w_dff_B_72b234om0_1;
	wire w_dff_B_uyXBKvGh3_1;
	wire w_dff_B_QDVmiuHX6_1;
	wire w_dff_B_Dkr9JPcC7_1;
	wire w_dff_B_2QfVLIYH5_0;
	wire w_dff_B_Wes1Bi1r1_0;
	wire w_dff_B_UIsyTEMs9_0;
	wire w_dff_B_4BfkN1Pp6_0;
	wire w_dff_B_BrBkJX9S6_0;
	wire w_dff_B_XQSODnrH6_0;
	wire w_dff_B_95JaTi651_0;
	wire w_dff_B_0hjvQMEF6_0;
	wire w_dff_B_LI958ltJ2_0;
	wire w_dff_B_2Gtl6xCK7_0;
	wire w_dff_B_In46HT6Z1_0;
	wire w_dff_B_rxc7WBZp7_0;
	wire w_dff_B_5QllazsF0_0;
	wire w_dff_B_pd7me7DP9_0;
	wire w_dff_B_Ng3dVv7L3_0;
	wire w_dff_B_paORnNy44_0;
	wire w_dff_B_tYW6IXLz0_0;
	wire w_dff_B_PNkgAw1z0_0;
	wire w_dff_B_jFxQUTmn4_0;
	wire w_dff_B_KOUcbzYt3_0;
	wire w_dff_B_c4kYWWfy1_0;
	wire w_dff_B_E8XILlGk4_0;
	wire w_dff_B_uirCvuzF7_0;
	wire w_dff_B_qr4s4FB56_0;
	wire w_dff_B_X7dPO1SY9_0;
	wire w_dff_B_bLwAzQAS1_0;
	wire w_dff_B_NQR8LqCj4_0;
	wire w_dff_B_gx2VO75d9_0;
	wire w_dff_B_e80M7d9g1_0;
	wire w_dff_B_0dzIYKbP7_0;
	wire w_dff_B_kY197Etg9_0;
	wire w_dff_B_i7ozsX6s0_0;
	wire w_dff_B_9KdxYw2t2_0;
	wire w_dff_B_xoD3q1Lo0_0;
	wire w_dff_B_h0i9s6pm8_0;
	wire w_dff_B_gyFCuJcJ4_0;
	wire w_dff_B_dZZslLEA1_0;
	wire w_dff_B_zcoK2CbP8_0;
	wire w_dff_B_LtYDAigb7_0;
	wire w_dff_B_xC8rs0ZH0_0;
	wire w_dff_B_97RnY4z27_0;
	wire w_dff_B_wwrpkPNY5_0;
	wire w_dff_B_KPx9lQ8r3_0;
	wire w_dff_B_qHUuajeQ1_0;
	wire w_dff_B_Pm4eCqHe4_0;
	wire w_dff_B_wI1OGoCG9_0;
	wire w_dff_B_3RujAxvW8_0;
	wire w_dff_B_Uoqk2gai7_0;
	wire w_dff_B_lQMt7VwU9_0;
	wire w_dff_B_DlHCO0Au0_0;
	wire w_dff_B_qOQepiXU5_0;
	wire w_dff_B_MKtVx2j64_0;
	wire w_dff_B_1HUQQNxE1_0;
	wire w_dff_B_9n9MJrX61_0;
	wire w_dff_B_HoqXpdaz5_0;
	wire w_dff_B_t6nFwwmc3_0;
	wire w_dff_B_nKknmpYo9_0;
	wire w_dff_B_rKedzUXh7_0;
	wire w_dff_B_V7vZN6FK0_0;
	wire w_dff_B_lQpIsANE1_0;
	wire w_dff_B_7aoBpfmz5_0;
	wire w_dff_B_g49WO7MT8_0;
	wire w_dff_B_MMDdDQD77_0;
	wire w_dff_B_nmYTSN6j2_0;
	wire w_dff_B_d8TqjGOz3_0;
	wire w_dff_B_IcaMaKP03_0;
	wire w_dff_B_yGQm8Yee8_0;
	wire w_dff_B_QtqRXhAW0_0;
	wire w_dff_B_QeyUCVkz9_0;
	wire w_dff_B_ZqSRhkFK7_0;
	wire w_dff_B_luahPtJk9_0;
	wire w_dff_B_onDud58R2_0;
	wire w_dff_B_MLyS5MlY8_0;
	wire w_dff_B_BhJ4dnG18_0;
	wire w_dff_B_ldVdQmma7_0;
	wire w_dff_B_1aJlZVpr2_0;
	wire w_dff_B_upfcGmyu1_0;
	wire w_dff_B_xV9BH7HW1_0;
	wire w_dff_B_kVcx0yfU9_0;
	wire w_dff_B_T9G1J35g1_0;
	wire w_dff_B_EybFPoWC5_0;
	wire w_dff_B_1xv37al60_0;
	wire w_dff_B_YOXAaZZZ7_0;
	wire w_dff_B_Mg0wGt1V0_0;
	wire w_dff_B_POLVBjgc3_0;
	wire w_dff_B_ZQprZfvQ5_0;
	wire w_dff_B_DqUs78GW9_0;
	wire w_dff_B_BszbWXgZ0_0;
	wire w_dff_B_1umRlSl88_0;
	wire w_dff_B_rm6x90Wr2_0;
	wire w_dff_B_FeSijBGi5_0;
	wire w_dff_B_9B6tyNHQ4_0;
	wire w_dff_B_HpvtjtJC5_0;
	wire w_dff_B_uIwZqBG17_0;
	wire w_dff_B_QpDocHiI5_0;
	wire w_dff_B_9Wsz7g1n1_0;
	wire w_dff_B_QWohCsaE2_0;
	wire w_dff_B_DxydY4YS6_0;
	wire w_dff_B_HSoN7PQp5_0;
	wire w_dff_B_d291vfqe6_0;
	wire w_dff_B_jGs1Z1vX5_0;
	wire w_dff_B_MK4eVmub9_0;
	wire w_dff_B_TfcBQnjB7_0;
	wire w_dff_B_gjEZsume5_0;
	wire w_dff_B_aGv1906U0_0;
	wire w_dff_B_JIAURANF6_0;
	wire w_dff_B_0v4CG99s9_0;
	wire w_dff_B_zhjxi2Ld9_0;
	wire w_dff_B_RArV20Il7_0;
	wire w_dff_B_kHjcuUnU5_0;
	wire w_dff_B_tR6hnRcF9_0;
	wire w_dff_B_X4yn2Anp8_0;
	wire w_dff_B_wtkyyWPf7_0;
	wire w_dff_B_Sl9F6Et71_0;
	wire w_dff_B_jTE3N4Z76_0;
	wire w_dff_B_4rxem5xX4_0;
	wire w_dff_B_sqISUf5R2_0;
	wire w_dff_B_aHDWCnpi6_0;
	wire w_dff_B_r5P8x6jF2_0;
	wire w_dff_B_zb1bl7zN4_0;
	wire w_dff_B_cidGYdUa6_0;
	wire w_dff_B_SQmXewmR4_0;
	wire w_dff_B_f8qTgXte9_1;
	wire w_dff_B_wA3ayJKz9_1;
	wire w_dff_B_WyYKA7pW5_1;
	wire w_dff_B_DAvIUI0Y4_1;
	wire w_dff_B_NMD9kh3O2_1;
	wire w_dff_B_eqxDkH0O8_1;
	wire w_dff_B_QNlR3t9x8_1;
	wire w_dff_B_Pi83P7Jj1_1;
	wire w_dff_B_yLelrGJg4_1;
	wire w_dff_B_265rvvmm7_1;
	wire w_dff_B_VIpU8MEZ7_1;
	wire w_dff_B_IR4m8D4z1_1;
	wire w_dff_B_kR8xyHfm8_1;
	wire w_dff_B_xJsZXO0B1_1;
	wire w_dff_B_d532XBxq9_1;
	wire w_dff_B_lBPAWRUn6_1;
	wire w_dff_B_lAZCmoHB9_1;
	wire w_dff_B_s2oQhqpx5_1;
	wire w_dff_B_LwVyTjA67_1;
	wire w_dff_B_KxcTmLCk6_1;
	wire w_dff_B_ojx8xbw63_1;
	wire w_dff_B_pxnZdb897_1;
	wire w_dff_B_yrZG7lNJ0_1;
	wire w_dff_B_pXzA0Phq4_1;
	wire w_dff_B_FyDdRiCH4_1;
	wire w_dff_B_GsYgYjUL2_1;
	wire w_dff_B_Y6rFuYd22_1;
	wire w_dff_B_dcMSza5I3_1;
	wire w_dff_B_6kx3AJcv9_1;
	wire w_dff_B_b3YpRzjt5_1;
	wire w_dff_B_oUWhOode7_1;
	wire w_dff_B_wjF3NDpp9_1;
	wire w_dff_B_6gLk7Eoc2_1;
	wire w_dff_B_eFZlryEr7_1;
	wire w_dff_B_Wj3Se4Si7_1;
	wire w_dff_B_6C6wDDRI7_1;
	wire w_dff_B_ULOEeAsr5_1;
	wire w_dff_B_dhJpIDDa4_1;
	wire w_dff_B_z7DTt5rD6_1;
	wire w_dff_B_KlTVUsek4_1;
	wire w_dff_B_cBByDh8p3_1;
	wire w_dff_B_2z1bpdKs2_1;
	wire w_dff_B_z7AfpNzJ1_1;
	wire w_dff_B_Za6DAwDP4_1;
	wire w_dff_B_rLMbyeqU8_1;
	wire w_dff_B_fhjaWZTg6_1;
	wire w_dff_B_7jtK5JmY3_1;
	wire w_dff_B_omyDYBd36_1;
	wire w_dff_B_hnAAJgEf7_1;
	wire w_dff_B_QoQ55iHQ4_1;
	wire w_dff_B_E5bJ3CFB0_1;
	wire w_dff_B_mOjoM2Lg9_1;
	wire w_dff_B_DQsGlLso2_1;
	wire w_dff_B_Cdfil6tL6_1;
	wire w_dff_B_o8JT9GyU6_1;
	wire w_dff_B_6bKoZvuP1_1;
	wire w_dff_B_PxObT3Vs6_1;
	wire w_dff_B_3dBdoVri1_1;
	wire w_dff_B_vBOC7GO92_1;
	wire w_dff_B_IFAYAUit5_1;
	wire w_dff_B_yXVD7yRc9_1;
	wire w_dff_B_U7bVR98W5_1;
	wire w_dff_B_unEQqwuE6_1;
	wire w_dff_B_d8TCTVuy2_1;
	wire w_dff_B_ET6JeDMn7_1;
	wire w_dff_B_wDNmYvA14_1;
	wire w_dff_B_xt6JAc2B0_1;
	wire w_dff_B_60AoPMW41_1;
	wire w_dff_B_t8sMV8DN2_1;
	wire w_dff_B_R85AbA0R6_1;
	wire w_dff_B_HIYxCD2f2_1;
	wire w_dff_B_B2eYx8Q56_1;
	wire w_dff_B_uf7oa47w9_1;
	wire w_dff_B_YPJ9nDUz1_1;
	wire w_dff_B_nMc59K3H8_1;
	wire w_dff_B_bCwx0H6p0_1;
	wire w_dff_B_gu03SAMI3_1;
	wire w_dff_B_zt312RzB2_1;
	wire w_dff_B_UM1NDhb67_1;
	wire w_dff_B_hYu6J6jU6_1;
	wire w_dff_B_mhyCqDbY7_1;
	wire w_dff_B_FRFxtHCR1_1;
	wire w_dff_B_VuOuJlF88_1;
	wire w_dff_B_17FqGLs39_1;
	wire w_dff_B_OOADEoCA0_1;
	wire w_dff_B_x4DAf78o5_1;
	wire w_dff_B_ATNpuaLy3_1;
	wire w_dff_B_pCOqBZ5a6_1;
	wire w_dff_B_7JFpEUAY0_1;
	wire w_dff_B_oZIYArVl3_1;
	wire w_dff_B_D8FKC54r8_1;
	wire w_dff_B_5f3WTAVR3_1;
	wire w_dff_B_qkFObSEu1_1;
	wire w_dff_B_oGDOMs2B4_1;
	wire w_dff_B_QvyQniSd7_1;
	wire w_dff_B_yLWVVCBF6_1;
	wire w_dff_B_RJLZJt0h9_1;
	wire w_dff_B_N1hPepM65_1;
	wire w_dff_B_0OGwauoM3_1;
	wire w_dff_B_PnYoe6II7_1;
	wire w_dff_B_SCCLtmRc5_1;
	wire w_dff_B_zEYqtAP65_1;
	wire w_dff_B_AMsAyZTz4_1;
	wire w_dff_B_oi0tPcgv1_1;
	wire w_dff_B_IGwUYizm5_1;
	wire w_dff_B_vP1BvdZd9_1;
	wire w_dff_B_nSQTaVBp1_1;
	wire w_dff_B_yVI5i3fN6_1;
	wire w_dff_B_B88AtstK2_1;
	wire w_dff_B_Tc3infSS9_1;
	wire w_dff_B_BM859FES4_1;
	wire w_dff_B_3BFB0Ztv8_1;
	wire w_dff_B_SM8s8saF5_1;
	wire w_dff_B_sICl1CVE1_1;
	wire w_dff_B_DSAnUEkB6_1;
	wire w_dff_B_ComdkNfQ3_1;
	wire w_dff_B_XXu7XgUA8_1;
	wire w_dff_B_9RfZLfa71_1;
	wire w_dff_B_ksM03QlX8_1;
	wire w_dff_B_MPBIqVyH9_1;
	wire w_dff_B_OendyP6K5_1;
	wire w_dff_B_tM9vMwNR4_0;
	wire w_dff_B_uhfXwzUK0_0;
	wire w_dff_B_XHOQ2RTY8_0;
	wire w_dff_B_73KsFIbG8_0;
	wire w_dff_B_SxANcsW96_0;
	wire w_dff_B_ppFd768R0_0;
	wire w_dff_B_lpXl7YPL9_0;
	wire w_dff_B_J9MsiBFx0_0;
	wire w_dff_B_C60neQfg4_0;
	wire w_dff_B_NgVd2CZr6_0;
	wire w_dff_B_2JwzRc4A8_0;
	wire w_dff_B_w5pizpHP7_0;
	wire w_dff_B_EuSPMpIl3_0;
	wire w_dff_B_um4AIsXm5_0;
	wire w_dff_B_6MmOjB9R5_0;
	wire w_dff_B_9XSbfqsG5_0;
	wire w_dff_B_Bp5qn2KU0_0;
	wire w_dff_B_Kh6MxY7r6_0;
	wire w_dff_B_Sqbvxk8B1_0;
	wire w_dff_B_GhAuJcPK3_0;
	wire w_dff_B_BulXm3oD5_0;
	wire w_dff_B_UtNuC4Me2_0;
	wire w_dff_B_VvVgAdlR8_0;
	wire w_dff_B_xlFP8uDR4_0;
	wire w_dff_B_MwNB2qsV2_0;
	wire w_dff_B_J9oGn0sy9_0;
	wire w_dff_B_M22xxVJq7_0;
	wire w_dff_B_emQo0S9V2_0;
	wire w_dff_B_gj13ySDt2_0;
	wire w_dff_B_SdpwCDWy9_0;
	wire w_dff_B_PXt43aUE0_0;
	wire w_dff_B_PQZUbu0R6_0;
	wire w_dff_B_okE9LWUO4_0;
	wire w_dff_B_aFeTWQFj3_0;
	wire w_dff_B_lGd3crRN0_0;
	wire w_dff_B_03Ua75Cb7_0;
	wire w_dff_B_nL371TK89_0;
	wire w_dff_B_vMAzRO376_0;
	wire w_dff_B_Sfu57Pet3_0;
	wire w_dff_B_Vfxkiga97_0;
	wire w_dff_B_0Du4hO558_0;
	wire w_dff_B_FQwcILQr1_0;
	wire w_dff_B_7deU1YPm7_0;
	wire w_dff_B_U6WaxnyG7_0;
	wire w_dff_B_IE4XmMqO1_0;
	wire w_dff_B_XIDhGfYe4_0;
	wire w_dff_B_BbSW8EG01_0;
	wire w_dff_B_01j2suE16_0;
	wire w_dff_B_ZQNxCRW28_0;
	wire w_dff_B_qs0z4ASg3_0;
	wire w_dff_B_Hb5oaEBn9_0;
	wire w_dff_B_aIXkLAfO7_0;
	wire w_dff_B_hzIHzoj10_0;
	wire w_dff_B_S9no621i9_0;
	wire w_dff_B_zdSxhAjc0_0;
	wire w_dff_B_Ihpyj1898_0;
	wire w_dff_B_djmgujPx9_0;
	wire w_dff_B_HHXF1L2n9_0;
	wire w_dff_B_pfSse2or9_0;
	wire w_dff_B_yoLIBYJa9_0;
	wire w_dff_B_t3JcdQsG3_0;
	wire w_dff_B_s6VMMbPr3_0;
	wire w_dff_B_ZrFR8mMC6_0;
	wire w_dff_B_bd95D6VF7_0;
	wire w_dff_B_VOdgSkbG9_0;
	wire w_dff_B_ghxMdhcM0_0;
	wire w_dff_B_Oa236skM5_0;
	wire w_dff_B_VA5Wc4EH5_0;
	wire w_dff_B_LpvTUo541_0;
	wire w_dff_B_1BZtxsHt4_0;
	wire w_dff_B_4nt7qEs50_0;
	wire w_dff_B_0aC17Nfq2_0;
	wire w_dff_B_DiQQ739I5_0;
	wire w_dff_B_6ecbn7gn4_0;
	wire w_dff_B_lMrzd39c6_0;
	wire w_dff_B_1DV4jHEs3_0;
	wire w_dff_B_nBgWTI0J3_0;
	wire w_dff_B_OhnaNYWH1_0;
	wire w_dff_B_64tDrTxv7_0;
	wire w_dff_B_2LR4zyBv1_0;
	wire w_dff_B_K8ptnSmK4_0;
	wire w_dff_B_LwH556Dk7_0;
	wire w_dff_B_z0aXwVt17_0;
	wire w_dff_B_tDRux8yC0_0;
	wire w_dff_B_GM9gKOZD0_0;
	wire w_dff_B_ICeIw2zD9_0;
	wire w_dff_B_DvyPNxlV8_0;
	wire w_dff_B_4awwGqWm6_0;
	wire w_dff_B_wmcfKzZl8_0;
	wire w_dff_B_2TFoYEKO8_0;
	wire w_dff_B_PQZmsKa46_0;
	wire w_dff_B_n73NktSA9_0;
	wire w_dff_B_50ryWj8f7_0;
	wire w_dff_B_e8KebvRU4_0;
	wire w_dff_B_HoUCemaA0_0;
	wire w_dff_B_YrOPCbeR4_0;
	wire w_dff_B_WDW6ZdUQ4_0;
	wire w_dff_B_yjJ4ndBe6_0;
	wire w_dff_B_kPdv9fzy6_0;
	wire w_dff_B_ZQHcXbS85_0;
	wire w_dff_B_XgwZm5Cj9_0;
	wire w_dff_B_uClfECq68_0;
	wire w_dff_B_MTcd4K5W2_0;
	wire w_dff_B_RHYhS3Pp0_0;
	wire w_dff_B_l6aiJ5Rp7_0;
	wire w_dff_B_uRpD9wvm9_0;
	wire w_dff_B_189KW5Mw0_0;
	wire w_dff_B_1gXPrIcA9_0;
	wire w_dff_B_YJ3IFZiO7_0;
	wire w_dff_B_PEAcNf6L2_0;
	wire w_dff_B_brIu6GOx4_0;
	wire w_dff_B_Kxq0iqGR4_0;
	wire w_dff_B_rUdkOYQS7_0;
	wire w_dff_B_Qmh2opri7_0;
	wire w_dff_B_0yt44FnY0_0;
	wire w_dff_B_TVVClLn13_0;
	wire w_dff_B_dw3rFMsF8_0;
	wire w_dff_B_iNsE2v409_0;
	wire w_dff_B_QOuDUobD7_0;
	wire w_dff_B_6CFEKehx6_0;
	wire w_dff_B_nEpywF7H8_0;
	wire w_dff_B_hcPXkUGE1_1;
	wire w_dff_B_XavnPH2f0_1;
	wire w_dff_B_NiDlEVIN3_1;
	wire w_dff_B_tsdEwm0t4_1;
	wire w_dff_B_FCy9SeUg6_1;
	wire w_dff_B_0Exq71OG3_1;
	wire w_dff_B_NPApAPev3_1;
	wire w_dff_B_sBpTzv4r9_1;
	wire w_dff_B_G4lqCRRS9_1;
	wire w_dff_B_7IAmLvla7_1;
	wire w_dff_B_GPatByqn8_1;
	wire w_dff_B_ZKEP9MCn9_1;
	wire w_dff_B_D3tTMyic2_1;
	wire w_dff_B_IBo4gq5x8_1;
	wire w_dff_B_0icHqgb25_1;
	wire w_dff_B_n2e5uGBN9_1;
	wire w_dff_B_hRxZAZiG2_1;
	wire w_dff_B_Rd3qvTtt0_1;
	wire w_dff_B_Jep5mWU60_1;
	wire w_dff_B_hZbkHOKL3_1;
	wire w_dff_B_qszaWM906_1;
	wire w_dff_B_49zXDCoS0_1;
	wire w_dff_B_7ofKzIcq7_1;
	wire w_dff_B_8fFQuj1P1_1;
	wire w_dff_B_fAzq0rhf7_1;
	wire w_dff_B_ggWrBE816_1;
	wire w_dff_B_LfEh797H2_1;
	wire w_dff_B_veqfGzta2_1;
	wire w_dff_B_GbvyUG1R8_1;
	wire w_dff_B_8VBbc0aR6_1;
	wire w_dff_B_Zs2b4iHb1_1;
	wire w_dff_B_EZVwhznK9_1;
	wire w_dff_B_PoMe8pHi9_1;
	wire w_dff_B_LeNXRqvp5_1;
	wire w_dff_B_mZf2a6280_1;
	wire w_dff_B_WCvTiAP60_1;
	wire w_dff_B_sbOnY7HQ4_1;
	wire w_dff_B_ZKH5Vzcn5_1;
	wire w_dff_B_bntmMVLk9_1;
	wire w_dff_B_QJYQALB37_1;
	wire w_dff_B_meGUUGBf9_1;
	wire w_dff_B_000zO23n4_1;
	wire w_dff_B_TBAxneeS1_1;
	wire w_dff_B_73HDM3X21_1;
	wire w_dff_B_pknlHcXd7_1;
	wire w_dff_B_Znt4o8t94_1;
	wire w_dff_B_9EbzWdIs4_1;
	wire w_dff_B_ujnXSU5j3_1;
	wire w_dff_B_9v9Cnyda0_1;
	wire w_dff_B_yMQhW0og4_1;
	wire w_dff_B_A97W2rSp1_1;
	wire w_dff_B_NNlyL4r45_1;
	wire w_dff_B_jb6OiXs53_1;
	wire w_dff_B_bh6ScHfj7_1;
	wire w_dff_B_i73NuGwF8_1;
	wire w_dff_B_3oSRHMcu2_1;
	wire w_dff_B_MY1TNxua8_1;
	wire w_dff_B_Gpy4nZj66_1;
	wire w_dff_B_M8iJ3Vjo0_1;
	wire w_dff_B_9GKw9ZeA2_1;
	wire w_dff_B_C6w6ReHm6_1;
	wire w_dff_B_Gejv70dY2_1;
	wire w_dff_B_DMNb6yXX3_1;
	wire w_dff_B_iASjosPi7_1;
	wire w_dff_B_SqGZmNoZ8_1;
	wire w_dff_B_BxmfDQnp5_1;
	wire w_dff_B_aYsRzhlY7_1;
	wire w_dff_B_dPkQc1ws0_1;
	wire w_dff_B_6joKHa8G6_1;
	wire w_dff_B_Tmao4VgQ4_1;
	wire w_dff_B_aMb3kUaa9_1;
	wire w_dff_B_rLZvEJYF1_1;
	wire w_dff_B_6xpklti30_1;
	wire w_dff_B_2CwzFqti7_1;
	wire w_dff_B_OznFFY1o0_1;
	wire w_dff_B_EW07CUuS2_1;
	wire w_dff_B_6FfilXMI5_1;
	wire w_dff_B_94zh6EBI2_1;
	wire w_dff_B_mkwV1cs23_1;
	wire w_dff_B_TDFNha2V0_1;
	wire w_dff_B_kJuc7Mag6_1;
	wire w_dff_B_idxkDdah9_1;
	wire w_dff_B_EEKgkwFg3_1;
	wire w_dff_B_64Zi7aej0_1;
	wire w_dff_B_0JplkbLq1_1;
	wire w_dff_B_K6GtJeIq1_1;
	wire w_dff_B_YkZSwbtn1_1;
	wire w_dff_B_cj0DCRd02_1;
	wire w_dff_B_rbMxRyTo5_1;
	wire w_dff_B_5tzGr4sn5_1;
	wire w_dff_B_rHvzfJJ14_1;
	wire w_dff_B_i8VpmdVF1_1;
	wire w_dff_B_MAneHMCi1_1;
	wire w_dff_B_SpCXiGba5_1;
	wire w_dff_B_H16gR1LR8_1;
	wire w_dff_B_EtPlqHiY4_1;
	wire w_dff_B_mCInpfKO7_1;
	wire w_dff_B_3bP3hiG91_1;
	wire w_dff_B_X5cDXw4r7_1;
	wire w_dff_B_OJL8zPrG4_1;
	wire w_dff_B_hBHzNRVd9_1;
	wire w_dff_B_dwQb54sa4_1;
	wire w_dff_B_RJCOAlA64_1;
	wire w_dff_B_vwzyujkD1_1;
	wire w_dff_B_9l6upuw68_1;
	wire w_dff_B_7ltLWsBY1_1;
	wire w_dff_B_iQBBJXrU8_1;
	wire w_dff_B_VXYiMtsS7_1;
	wire w_dff_B_b0te6clD6_1;
	wire w_dff_B_dPftqRX89_1;
	wire w_dff_B_Zmadsj9k4_1;
	wire w_dff_B_Ix7BLOaU6_1;
	wire w_dff_B_VFrBBxDi6_1;
	wire w_dff_B_CozY5rtY7_1;
	wire w_dff_B_CK5ljyiq2_1;
	wire w_dff_B_wckZfDj72_1;
	wire w_dff_B_ElPFh7Of1_1;
	wire w_dff_B_cixnBFfE0_1;
	wire w_dff_B_sKL4thCY2_1;
	wire w_dff_B_1R6I2MTe0_1;
	wire w_dff_B_DmiS8B3L6_0;
	wire w_dff_B_xM345Y5V1_0;
	wire w_dff_B_oSVMpu7v5_0;
	wire w_dff_B_KouUV3Fd1_0;
	wire w_dff_B_Yy1fBsMj8_0;
	wire w_dff_B_nAvb8QQy7_0;
	wire w_dff_B_wkengbpg0_0;
	wire w_dff_B_dfED2d4k5_0;
	wire w_dff_B_dJHgZWeo9_0;
	wire w_dff_B_ljmptqht0_0;
	wire w_dff_B_Kyq8mKWQ1_0;
	wire w_dff_B_s1mHkyUz2_0;
	wire w_dff_B_0loYNIRv6_0;
	wire w_dff_B_jdQ8jHyh8_0;
	wire w_dff_B_E1V2KQSA9_0;
	wire w_dff_B_zMfk9k0r8_0;
	wire w_dff_B_3RRmFZWD3_0;
	wire w_dff_B_2c5LqGLI7_0;
	wire w_dff_B_lViASZIE5_0;
	wire w_dff_B_mPEnpJo82_0;
	wire w_dff_B_nNwMIVFG9_0;
	wire w_dff_B_7ktKAge17_0;
	wire w_dff_B_xsGop4tW1_0;
	wire w_dff_B_MPpvUto57_0;
	wire w_dff_B_W9XfOpxT6_0;
	wire w_dff_B_hZWpFjNb3_0;
	wire w_dff_B_x1rojjt17_0;
	wire w_dff_B_dNqLqrhV5_0;
	wire w_dff_B_T3qWaSKq3_0;
	wire w_dff_B_Xm1Erx5e7_0;
	wire w_dff_B_wHWGp6hT9_0;
	wire w_dff_B_bW9oJaLB3_0;
	wire w_dff_B_wu9PpQbf9_0;
	wire w_dff_B_iBx7VdQm5_0;
	wire w_dff_B_N72PAhuE2_0;
	wire w_dff_B_FFOjzuJe2_0;
	wire w_dff_B_slu5ZbCq0_0;
	wire w_dff_B_v9KEctaI6_0;
	wire w_dff_B_KBKTvPqe1_0;
	wire w_dff_B_mCLtrh4K2_0;
	wire w_dff_B_w7nRcUPN4_0;
	wire w_dff_B_m7SxjzDl7_0;
	wire w_dff_B_ZKKb9tCi2_0;
	wire w_dff_B_kR8FmrOM0_0;
	wire w_dff_B_tBfkhtXm6_0;
	wire w_dff_B_pLKwh8m85_0;
	wire w_dff_B_guDWjVXa2_0;
	wire w_dff_B_tw7DMU3u7_0;
	wire w_dff_B_AZ7Okffn0_0;
	wire w_dff_B_ppIKGOWx6_0;
	wire w_dff_B_uvX2sCY46_0;
	wire w_dff_B_obRL9Nk68_0;
	wire w_dff_B_qWD0E8fM5_0;
	wire w_dff_B_z0aR4dFB1_0;
	wire w_dff_B_0DOth7S28_0;
	wire w_dff_B_xeLSmYp20_0;
	wire w_dff_B_c2xrgluw2_0;
	wire w_dff_B_d6r4A8FF6_0;
	wire w_dff_B_JEvOvgSL6_0;
	wire w_dff_B_xYXnW7nk7_0;
	wire w_dff_B_SOqUhn952_0;
	wire w_dff_B_SAxdX41Y0_0;
	wire w_dff_B_Hcbg1YCr6_0;
	wire w_dff_B_PGV85OmQ9_0;
	wire w_dff_B_j54TmuRa9_0;
	wire w_dff_B_bztkgWoP0_0;
	wire w_dff_B_qjPM2jJE8_0;
	wire w_dff_B_okt0GNZc0_0;
	wire w_dff_B_25Fh1sIl3_0;
	wire w_dff_B_EKVjkUM46_0;
	wire w_dff_B_q9JfqPeX9_0;
	wire w_dff_B_uPnr1PXO2_0;
	wire w_dff_B_Ase3oQJF2_0;
	wire w_dff_B_ELk0EIzV2_0;
	wire w_dff_B_I3pdV6ZQ7_0;
	wire w_dff_B_VMtiRCuB4_0;
	wire w_dff_B_69LrehmD4_0;
	wire w_dff_B_FVWarx0c0_0;
	wire w_dff_B_WkrqLDnN7_0;
	wire w_dff_B_i0uWrgGi7_0;
	wire w_dff_B_YesU9k7I7_0;
	wire w_dff_B_e4Q0tUh28_0;
	wire w_dff_B_49iqi9vY3_0;
	wire w_dff_B_i0V7VUL25_0;
	wire w_dff_B_wU6ltCAi4_0;
	wire w_dff_B_mGSRjdud1_0;
	wire w_dff_B_iUAbyBWy9_0;
	wire w_dff_B_bZgMucZP1_0;
	wire w_dff_B_nRGCw61o8_0;
	wire w_dff_B_81XXrLxH6_0;
	wire w_dff_B_WFX7lA4x4_0;
	wire w_dff_B_ADdjmPg34_0;
	wire w_dff_B_xiMQvOmp7_0;
	wire w_dff_B_XHdonrsG8_0;
	wire w_dff_B_oQaVnIZW9_0;
	wire w_dff_B_wu6hGo3Y6_0;
	wire w_dff_B_wC10m9iq3_0;
	wire w_dff_B_5A8lEkG11_0;
	wire w_dff_B_ZQ3O21mD6_0;
	wire w_dff_B_oFzw8wIp7_0;
	wire w_dff_B_oVB96x231_0;
	wire w_dff_B_s6kolGIt8_0;
	wire w_dff_B_QmsGdkTE8_0;
	wire w_dff_B_IkOAgSwj0_0;
	wire w_dff_B_hRaer5xI2_0;
	wire w_dff_B_rwRBUbz36_0;
	wire w_dff_B_9ykGo8Rk9_0;
	wire w_dff_B_901ryyiL2_0;
	wire w_dff_B_kvAOLe5b5_0;
	wire w_dff_B_0gEsQm253_0;
	wire w_dff_B_gCBSyele0_0;
	wire w_dff_B_fToHlPGI9_0;
	wire w_dff_B_8veaDZvP9_0;
	wire w_dff_B_rYFOO46L8_0;
	wire w_dff_B_RXU664dX3_0;
	wire w_dff_B_GeyrJEWw2_0;
	wire w_dff_B_Xua6oPfC8_0;
	wire w_dff_B_f4y5YBEj1_0;
	wire w_dff_B_VUdKXJJA4_0;
	wire w_dff_B_urlYAJ559_0;
	wire w_dff_B_6ZJ2B90F4_1;
	wire w_dff_B_XgC1VJGa5_1;
	wire w_dff_B_WmFTPlty5_1;
	wire w_dff_B_8EtGIwQl3_1;
	wire w_dff_B_wkSUwda18_1;
	wire w_dff_B_VwBccq4w1_1;
	wire w_dff_B_M7KbPZg11_1;
	wire w_dff_B_C1gAATUa6_1;
	wire w_dff_B_qeGtAeP11_1;
	wire w_dff_B_20oawz8w8_1;
	wire w_dff_B_4brz1GLZ3_1;
	wire w_dff_B_zrub0edS1_1;
	wire w_dff_B_sM48ITAY0_1;
	wire w_dff_B_Xu8dHqAK3_1;
	wire w_dff_B_fL4r92p34_1;
	wire w_dff_B_WfLpBtFN7_1;
	wire w_dff_B_iz6GKrWj5_1;
	wire w_dff_B_wyixcF4B0_1;
	wire w_dff_B_AO8gYpzD9_1;
	wire w_dff_B_uOiJMq6z7_1;
	wire w_dff_B_WO3mDd509_1;
	wire w_dff_B_EDFrqSX08_1;
	wire w_dff_B_4SwMoBnw2_1;
	wire w_dff_B_YdzkRIGQ2_1;
	wire w_dff_B_e1ZjCM265_1;
	wire w_dff_B_LPgF5hbc9_1;
	wire w_dff_B_6dyapKtA8_1;
	wire w_dff_B_0QxXBDYG7_1;
	wire w_dff_B_98SYshbP6_1;
	wire w_dff_B_urFNhsEF8_1;
	wire w_dff_B_PIt4L3yH5_1;
	wire w_dff_B_EPL9IKN54_1;
	wire w_dff_B_Of9cqFmO5_1;
	wire w_dff_B_GISs8RJ51_1;
	wire w_dff_B_dYhzJzpb8_1;
	wire w_dff_B_8Ly5VTXd8_1;
	wire w_dff_B_DbFJDAab5_1;
	wire w_dff_B_ZG6E00pS5_1;
	wire w_dff_B_V9E5ZCbc0_1;
	wire w_dff_B_zPKZP7zU2_1;
	wire w_dff_B_BrVhiL6R4_1;
	wire w_dff_B_VutLSd6n2_1;
	wire w_dff_B_JFCPEFzO0_1;
	wire w_dff_B_30izPVSv6_1;
	wire w_dff_B_Wk0fSFGf1_1;
	wire w_dff_B_SXk16agu8_1;
	wire w_dff_B_PvVYcDLX3_1;
	wire w_dff_B_qoCEinwP9_1;
	wire w_dff_B_o1h7roaU7_1;
	wire w_dff_B_JB3fTzTe2_1;
	wire w_dff_B_jm7fkLfB0_1;
	wire w_dff_B_XNEXT1Yz7_1;
	wire w_dff_B_YRJHmesp2_1;
	wire w_dff_B_SqtNvor55_1;
	wire w_dff_B_iPznLBaZ5_1;
	wire w_dff_B_mMYuIlKN1_1;
	wire w_dff_B_2NAZTEHk9_1;
	wire w_dff_B_9Ww78L353_1;
	wire w_dff_B_kRLCanVC8_1;
	wire w_dff_B_HZqQIV0C5_1;
	wire w_dff_B_M1Si2zLj9_1;
	wire w_dff_B_2Y7KoNG93_1;
	wire w_dff_B_3cnDEG7O2_1;
	wire w_dff_B_NQ50Ym6f1_1;
	wire w_dff_B_PYA67cGF4_1;
	wire w_dff_B_nayPBG5B4_1;
	wire w_dff_B_4ulNaD3g2_1;
	wire w_dff_B_kDmaarHJ3_1;
	wire w_dff_B_Bnr84nrE0_1;
	wire w_dff_B_pq6LVOGV7_1;
	wire w_dff_B_drpfdpA27_1;
	wire w_dff_B_PJuHsV6V7_1;
	wire w_dff_B_fa5dLJkX3_1;
	wire w_dff_B_RTmzCHU50_1;
	wire w_dff_B_OLvzY3yV7_1;
	wire w_dff_B_n24jqsHS5_1;
	wire w_dff_B_PdbcKl9C7_1;
	wire w_dff_B_hsnAgIWa7_1;
	wire w_dff_B_ym7hkXN32_1;
	wire w_dff_B_7L1oB9EE3_1;
	wire w_dff_B_ApfBJJJa7_1;
	wire w_dff_B_q6X1lfWl7_1;
	wire w_dff_B_YTRcjFPY5_1;
	wire w_dff_B_Gcy5hbj28_1;
	wire w_dff_B_CZQncF1E6_1;
	wire w_dff_B_JBLnxQhL5_1;
	wire w_dff_B_VoUNmmqo6_1;
	wire w_dff_B_63FwWgcJ4_1;
	wire w_dff_B_pXt3VUrN4_1;
	wire w_dff_B_ybk2Lthi7_1;
	wire w_dff_B_sEFt6puM4_1;
	wire w_dff_B_InfOptXn7_1;
	wire w_dff_B_GJsT1EFX3_1;
	wire w_dff_B_KFZzT8EC1_1;
	wire w_dff_B_zeegFoI83_1;
	wire w_dff_B_oNZa8tcN5_1;
	wire w_dff_B_wEZ7oaDq3_1;
	wire w_dff_B_kdT267tF2_1;
	wire w_dff_B_ByNyOFpy6_1;
	wire w_dff_B_9P3BuhQo2_1;
	wire w_dff_B_vN3PQZCt4_1;
	wire w_dff_B_Gai0xEha7_1;
	wire w_dff_B_7UDU43za0_1;
	wire w_dff_B_2VUUf3kt9_1;
	wire w_dff_B_rZOacF6j8_1;
	wire w_dff_B_FPE0Tijx2_1;
	wire w_dff_B_ThiYQWt53_1;
	wire w_dff_B_VJrSGc3j8_1;
	wire w_dff_B_mddY9Gl86_1;
	wire w_dff_B_j3h3KUec4_1;
	wire w_dff_B_NSTQJrwo2_1;
	wire w_dff_B_o2gN1zCD0_1;
	wire w_dff_B_XTp20tg52_1;
	wire w_dff_B_Pv7emCxc2_1;
	wire w_dff_B_phve4e6S7_1;
	wire w_dff_B_2HboaWI04_1;
	wire w_dff_B_Gbt3fbkn3_1;
	wire w_dff_B_ClWslrlp8_1;
	wire w_dff_B_UxHmoAjS1_1;
	wire w_dff_B_OBvIyR2T2_0;
	wire w_dff_B_eWmltQAJ2_0;
	wire w_dff_B_Y72cGf7J8_0;
	wire w_dff_B_BC3x89br9_0;
	wire w_dff_B_MEM72NPB9_0;
	wire w_dff_B_Rxh12fnE0_0;
	wire w_dff_B_UoFrLTCG1_0;
	wire w_dff_B_3OINwGFg5_0;
	wire w_dff_B_mUYbJReH6_0;
	wire w_dff_B_TNRdxHUH4_0;
	wire w_dff_B_4YzXJCMG6_0;
	wire w_dff_B_1EZGvYVA3_0;
	wire w_dff_B_rVw9kkY29_0;
	wire w_dff_B_5xkRPJOT0_0;
	wire w_dff_B_euOwuYcp1_0;
	wire w_dff_B_3s9L8Xct4_0;
	wire w_dff_B_k7W7nsZ06_0;
	wire w_dff_B_7NcmlQOG5_0;
	wire w_dff_B_xTQDePxT7_0;
	wire w_dff_B_e5nEBnQ64_0;
	wire w_dff_B_Cf6qzudz3_0;
	wire w_dff_B_QXgl2pq38_0;
	wire w_dff_B_i3mZi5lB3_0;
	wire w_dff_B_8JW7Ni1S3_0;
	wire w_dff_B_LKO01fNs5_0;
	wire w_dff_B_eMsTXzsS2_0;
	wire w_dff_B_YuiZujfi8_0;
	wire w_dff_B_6eZnYLSU0_0;
	wire w_dff_B_dUlwXxJt7_0;
	wire w_dff_B_ymEwlZYF7_0;
	wire w_dff_B_3G7ikQ5o6_0;
	wire w_dff_B_pQvlhuLM9_0;
	wire w_dff_B_ufgw2k0D4_0;
	wire w_dff_B_SGEmeXaY1_0;
	wire w_dff_B_dClj0k4s2_0;
	wire w_dff_B_Jq6PPaxS6_0;
	wire w_dff_B_lRd8Bw9X9_0;
	wire w_dff_B_ZMqTcW402_0;
	wire w_dff_B_IZ6xCIZG4_0;
	wire w_dff_B_0GZFFMdT6_0;
	wire w_dff_B_6EBpYBOK9_0;
	wire w_dff_B_dUEPX3IQ8_0;
	wire w_dff_B_4EUFmaEt2_0;
	wire w_dff_B_EXZkEsnB0_0;
	wire w_dff_B_nNv8vYer8_0;
	wire w_dff_B_OtnZcrah8_0;
	wire w_dff_B_rLGjJ4bu1_0;
	wire w_dff_B_b07krKOj1_0;
	wire w_dff_B_0kuo0w8A7_0;
	wire w_dff_B_bzSXEorl7_0;
	wire w_dff_B_ujWic2xz4_0;
	wire w_dff_B_JqlrhBWN9_0;
	wire w_dff_B_edZwPy4H8_0;
	wire w_dff_B_fXIJTsZQ2_0;
	wire w_dff_B_atBFjTsy7_0;
	wire w_dff_B_sVCfwL192_0;
	wire w_dff_B_KZGo2XtR5_0;
	wire w_dff_B_uDWde4n81_0;
	wire w_dff_B_njBhggTg5_0;
	wire w_dff_B_P5Hzo2Zp1_0;
	wire w_dff_B_4BfguwV94_0;
	wire w_dff_B_HkBAUb3b0_0;
	wire w_dff_B_ngRyoD7x8_0;
	wire w_dff_B_oEZXVowk2_0;
	wire w_dff_B_8K6VsHfA3_0;
	wire w_dff_B_l6DYfbgB3_0;
	wire w_dff_B_mwtPgu9c0_0;
	wire w_dff_B_xFbV3PoU2_0;
	wire w_dff_B_AgqJIlai1_0;
	wire w_dff_B_1nPrVcnp2_0;
	wire w_dff_B_5zKXETA53_0;
	wire w_dff_B_8epVmzz87_0;
	wire w_dff_B_N5cJ9LNb5_0;
	wire w_dff_B_afPq0GAY8_0;
	wire w_dff_B_5XU8T3Mw8_0;
	wire w_dff_B_XQ2xL5tM2_0;
	wire w_dff_B_vzYWFa9T8_0;
	wire w_dff_B_nMCaWRfT6_0;
	wire w_dff_B_m2LfiuhB0_0;
	wire w_dff_B_RrwnGvqr5_0;
	wire w_dff_B_unXnc3AO8_0;
	wire w_dff_B_Hu2gvB395_0;
	wire w_dff_B_mWU2Bni57_0;
	wire w_dff_B_qxljZjVO0_0;
	wire w_dff_B_CNui0XvE3_0;
	wire w_dff_B_Eo4JERnf8_0;
	wire w_dff_B_d8B3KVR47_0;
	wire w_dff_B_P1cmW4xQ4_0;
	wire w_dff_B_LBXBeSez1_0;
	wire w_dff_B_8KmYPTae8_0;
	wire w_dff_B_14oMNk0D7_0;
	wire w_dff_B_Rnhj953L7_0;
	wire w_dff_B_ZvnWeP999_0;
	wire w_dff_B_3fAtqGT09_0;
	wire w_dff_B_aAhtehik0_0;
	wire w_dff_B_o6Rq3phW0_0;
	wire w_dff_B_cnh7sGxs4_0;
	wire w_dff_B_UhYaz45r0_0;
	wire w_dff_B_heSdbbWs5_0;
	wire w_dff_B_L3uyP2X62_0;
	wire w_dff_B_zIWosCQc7_0;
	wire w_dff_B_ZNc4ox7c3_0;
	wire w_dff_B_ZOLbvdtG2_0;
	wire w_dff_B_x1mt1XC68_0;
	wire w_dff_B_oIFa4bEX1_0;
	wire w_dff_B_iQmPgdEz3_0;
	wire w_dff_B_Ch1LW24n7_0;
	wire w_dff_B_rOyHgDks8_0;
	wire w_dff_B_kGDwxasu3_0;
	wire w_dff_B_wHLiDIXZ9_0;
	wire w_dff_B_j1x5kQTT0_0;
	wire w_dff_B_uAUjPAjr6_0;
	wire w_dff_B_rXf4j4Y44_0;
	wire w_dff_B_nEavyAKv3_0;
	wire w_dff_B_QcxVJFj87_0;
	wire w_dff_B_LrzuCVep6_0;
	wire w_dff_B_J9zqpGSM3_0;
	wire w_dff_B_mAq3ZGyQ2_0;
	wire w_dff_B_JSc81Qhc2_0;
	wire w_dff_B_sYq6oIB27_1;
	wire w_dff_B_Mc2PPan17_1;
	wire w_dff_B_4qKbGJTO6_1;
	wire w_dff_B_14xh7Ujc8_1;
	wire w_dff_B_xwiTDYel3_1;
	wire w_dff_B_rTuSd1994_1;
	wire w_dff_B_8cR0rBkV4_1;
	wire w_dff_B_5JI2EuHq8_1;
	wire w_dff_B_DZkDuAc95_1;
	wire w_dff_B_ATEK1pgC7_1;
	wire w_dff_B_U5pTLMyQ0_1;
	wire w_dff_B_S9U0rcYm5_1;
	wire w_dff_B_cfPrY5Fi9_1;
	wire w_dff_B_aXfLR1ZS2_1;
	wire w_dff_B_IKfIb25a1_1;
	wire w_dff_B_389xdMPT9_1;
	wire w_dff_B_3VHdWk4Q2_1;
	wire w_dff_B_5nYmQITp2_1;
	wire w_dff_B_oxm5N6Bn3_1;
	wire w_dff_B_qWa1F2rv8_1;
	wire w_dff_B_repZVBIo9_1;
	wire w_dff_B_TmJcs3DT1_1;
	wire w_dff_B_cyz57FfY7_1;
	wire w_dff_B_55ap0eZ79_1;
	wire w_dff_B_qv9xgGOe2_1;
	wire w_dff_B_GUSy8BVL6_1;
	wire w_dff_B_Tfg8qDL46_1;
	wire w_dff_B_QRI6PbSb5_1;
	wire w_dff_B_xAuy5jje1_1;
	wire w_dff_B_dmKlRpZe2_1;
	wire w_dff_B_64Fs2Iib3_1;
	wire w_dff_B_2K2x6IeT6_1;
	wire w_dff_B_SAKsbJUN6_1;
	wire w_dff_B_E07jwBMe0_1;
	wire w_dff_B_kMxHPedC1_1;
	wire w_dff_B_JYngolCI4_1;
	wire w_dff_B_ODzATTYR9_1;
	wire w_dff_B_GnLQI6qe3_1;
	wire w_dff_B_Z0zr7KT67_1;
	wire w_dff_B_ExfL3PUW8_1;
	wire w_dff_B_GNT1NYBN3_1;
	wire w_dff_B_uomdK2v57_1;
	wire w_dff_B_qRHjwwew8_1;
	wire w_dff_B_nB5crXne1_1;
	wire w_dff_B_kZAoHPhN5_1;
	wire w_dff_B_cxsi7iuI6_1;
	wire w_dff_B_pf5jKgF90_1;
	wire w_dff_B_VPlu4Mi47_1;
	wire w_dff_B_H3zG7Jxj5_1;
	wire w_dff_B_VEUU7NPZ3_1;
	wire w_dff_B_oIkXknC90_1;
	wire w_dff_B_6s7AcXor9_1;
	wire w_dff_B_SwbCaKMk0_1;
	wire w_dff_B_S9QDlWnx4_1;
	wire w_dff_B_pdKY1lxM4_1;
	wire w_dff_B_u3lptrnf8_1;
	wire w_dff_B_GbBouQ5h7_1;
	wire w_dff_B_EI245wFH6_1;
	wire w_dff_B_ETIGfcFn8_1;
	wire w_dff_B_2AMTPYFz5_1;
	wire w_dff_B_1HLApl003_1;
	wire w_dff_B_8JnTbCBE4_1;
	wire w_dff_B_N5jV3Jlw4_1;
	wire w_dff_B_34Yuk4Sg7_1;
	wire w_dff_B_E7KxLBXn5_1;
	wire w_dff_B_HAqv7guS4_1;
	wire w_dff_B_ZEdYL15L5_1;
	wire w_dff_B_z2K6vSV76_1;
	wire w_dff_B_EbPlB7874_1;
	wire w_dff_B_aene9t648_1;
	wire w_dff_B_8Henj0RT7_1;
	wire w_dff_B_lSUaYgkw1_1;
	wire w_dff_B_W1RGT3kX4_1;
	wire w_dff_B_L2Yyhw4X1_1;
	wire w_dff_B_OAK4GISu9_1;
	wire w_dff_B_n6MpM0oR2_1;
	wire w_dff_B_WgCHhUfe4_1;
	wire w_dff_B_V24btCTU1_1;
	wire w_dff_B_46iaAK8d8_1;
	wire w_dff_B_GRRWWKgJ3_1;
	wire w_dff_B_LSoTwvbM4_1;
	wire w_dff_B_5H1TghRK9_1;
	wire w_dff_B_nYUPnOY41_1;
	wire w_dff_B_WFoDYRVC3_1;
	wire w_dff_B_m5g4kFHf0_1;
	wire w_dff_B_uYMdIVgf0_1;
	wire w_dff_B_SVUFnekn2_1;
	wire w_dff_B_6OfZvN8s7_1;
	wire w_dff_B_ac5b9gd27_1;
	wire w_dff_B_9oCCIevO5_1;
	wire w_dff_B_6rRwW7Ws4_1;
	wire w_dff_B_tY1rLmmh2_1;
	wire w_dff_B_OCEhKZzF9_1;
	wire w_dff_B_Et1lDeqa9_1;
	wire w_dff_B_1VOxYzwg9_1;
	wire w_dff_B_64aPibxn5_1;
	wire w_dff_B_eKWjpM350_1;
	wire w_dff_B_V500e5aP3_1;
	wire w_dff_B_U74oms4w5_1;
	wire w_dff_B_p8i8DXbS3_1;
	wire w_dff_B_bSrTy1ev8_1;
	wire w_dff_B_aBlLHLBO6_1;
	wire w_dff_B_Bs4WsX2g9_1;
	wire w_dff_B_4JDGpC0g4_1;
	wire w_dff_B_p2Dyonl82_1;
	wire w_dff_B_BBY7MKTB9_1;
	wire w_dff_B_r2RFdo4Y5_1;
	wire w_dff_B_LIENfJEl4_1;
	wire w_dff_B_ZHJlxTIa7_1;
	wire w_dff_B_dGDIGRuM0_1;
	wire w_dff_B_TeLvXY2Y6_1;
	wire w_dff_B_Izmrb4xg5_1;
	wire w_dff_B_tuOP7eqL8_1;
	wire w_dff_B_dMzdyEiI6_1;
	wire w_dff_B_hB0Mxx1g3_1;
	wire w_dff_B_hhejUK2T5_1;
	wire w_dff_B_W6b68rBH3_1;
	wire w_dff_B_hW63y0Sx4_1;
	wire w_dff_B_syFTwmB93_0;
	wire w_dff_B_rGkd5r7P5_0;
	wire w_dff_B_OlmzySVc6_0;
	wire w_dff_B_Ut9vB0XY6_0;
	wire w_dff_B_EoLinNfp9_0;
	wire w_dff_B_6j2dYUEX7_0;
	wire w_dff_B_z2173c6s1_0;
	wire w_dff_B_On7zB16x4_0;
	wire w_dff_B_biyyJnSh6_0;
	wire w_dff_B_TezYp0Ra8_0;
	wire w_dff_B_braLNV6O5_0;
	wire w_dff_B_ZeUtcFsF7_0;
	wire w_dff_B_zC3DyTHw6_0;
	wire w_dff_B_SvOZJ9Gi3_0;
	wire w_dff_B_ky4sKzd06_0;
	wire w_dff_B_gE3zK0w63_0;
	wire w_dff_B_YAnSMdnK3_0;
	wire w_dff_B_9Q80FKWm6_0;
	wire w_dff_B_TR0D03kd1_0;
	wire w_dff_B_GRLNTJPk4_0;
	wire w_dff_B_22X2GU6B4_0;
	wire w_dff_B_b5lIMHw38_0;
	wire w_dff_B_K1i8waze1_0;
	wire w_dff_B_XFLWQoGc7_0;
	wire w_dff_B_GSByVAd25_0;
	wire w_dff_B_MtzmmXRR6_0;
	wire w_dff_B_cbNpikyc7_0;
	wire w_dff_B_YNm8l35B3_0;
	wire w_dff_B_7apRK40L8_0;
	wire w_dff_B_XIt328QY0_0;
	wire w_dff_B_7l6hmQ2M6_0;
	wire w_dff_B_pfmQUzfS4_0;
	wire w_dff_B_IPy17bNt9_0;
	wire w_dff_B_1Et8djZy2_0;
	wire w_dff_B_fCD8ZvnQ2_0;
	wire w_dff_B_l3TqqqL40_0;
	wire w_dff_B_5UKu6m229_0;
	wire w_dff_B_FHMUvI1i3_0;
	wire w_dff_B_tH7rGPYO5_0;
	wire w_dff_B_Lj3TNSSx7_0;
	wire w_dff_B_zviujcVA6_0;
	wire w_dff_B_rWTKYZYJ1_0;
	wire w_dff_B_6WqjrJA54_0;
	wire w_dff_B_ZHDe1QPz3_0;
	wire w_dff_B_Q4rko9hu3_0;
	wire w_dff_B_2O1AmU713_0;
	wire w_dff_B_NFRIOZh67_0;
	wire w_dff_B_lo9ZQOI16_0;
	wire w_dff_B_ofOAyfxh7_0;
	wire w_dff_B_fzgk1dLt9_0;
	wire w_dff_B_HS7BREav1_0;
	wire w_dff_B_uD5oK2bF2_0;
	wire w_dff_B_eOv37QLa0_0;
	wire w_dff_B_8bTL8iVs7_0;
	wire w_dff_B_Yn0zx3027_0;
	wire w_dff_B_z5vT4OBK5_0;
	wire w_dff_B_g87oetmx9_0;
	wire w_dff_B_gzj3X2n83_0;
	wire w_dff_B_xICX0ZDl7_0;
	wire w_dff_B_sBJqN9m51_0;
	wire w_dff_B_VH8U2p3E4_0;
	wire w_dff_B_SZttFc7V6_0;
	wire w_dff_B_JjBTIVlq7_0;
	wire w_dff_B_k8niOOyu4_0;
	wire w_dff_B_XnQzF0iA4_0;
	wire w_dff_B_RegjiEZj8_0;
	wire w_dff_B_NybTSBVG7_0;
	wire w_dff_B_3WTVIihh4_0;
	wire w_dff_B_T8lG7MNp5_0;
	wire w_dff_B_5ZteBW1k8_0;
	wire w_dff_B_TldflRhm2_0;
	wire w_dff_B_r1gEPlLE9_0;
	wire w_dff_B_yjFeG0Ie1_0;
	wire w_dff_B_pvQFLMEh1_0;
	wire w_dff_B_tN67ZL9p9_0;
	wire w_dff_B_2y2p9ZtR8_0;
	wire w_dff_B_oCxJMgs76_0;
	wire w_dff_B_QWiCdKsj9_0;
	wire w_dff_B_yaSwftAH4_0;
	wire w_dff_B_tpsQhyHM6_0;
	wire w_dff_B_TU5WsVp09_0;
	wire w_dff_B_VATC0ZSr1_0;
	wire w_dff_B_QbGTHADZ6_0;
	wire w_dff_B_sT7RScMQ8_0;
	wire w_dff_B_yKyhJFUi5_0;
	wire w_dff_B_fFXzhb695_0;
	wire w_dff_B_pYbeUMXS7_0;
	wire w_dff_B_P25KHeJ97_0;
	wire w_dff_B_4ghMgmNn1_0;
	wire w_dff_B_FaRzaNcD9_0;
	wire w_dff_B_v7bfzJ8b8_0;
	wire w_dff_B_ndlISqRV8_0;
	wire w_dff_B_wAapW3Cd0_0;
	wire w_dff_B_2a2fGktN2_0;
	wire w_dff_B_SUJAiTxQ9_0;
	wire w_dff_B_fvMxO81f6_0;
	wire w_dff_B_8XPyocbv2_0;
	wire w_dff_B_bnveSGRw9_0;
	wire w_dff_B_FmRSMsMy7_0;
	wire w_dff_B_ZkNNlGdm5_0;
	wire w_dff_B_vv73V3B65_0;
	wire w_dff_B_go8YdW1i5_0;
	wire w_dff_B_blbbGZV41_0;
	wire w_dff_B_0b0N0YCK5_0;
	wire w_dff_B_kQMGscL80_0;
	wire w_dff_B_xXGtxy0E0_0;
	wire w_dff_B_sSzFJBc48_0;
	wire w_dff_B_L0Gow7Jz5_0;
	wire w_dff_B_OSMMiefa9_0;
	wire w_dff_B_7v4lYdnc4_0;
	wire w_dff_B_XfwMWNn70_0;
	wire w_dff_B_wkxq2Bkn0_0;
	wire w_dff_B_59cngZlb0_0;
	wire w_dff_B_UHQtzWZl8_0;
	wire w_dff_B_vgJcCKrd6_0;
	wire w_dff_B_e0HN5Sku6_0;
	wire w_dff_B_xoZojuwa7_0;
	wire w_dff_B_PG2MTWyb5_0;
	wire w_dff_B_VHn9TJQs4_1;
	wire w_dff_B_weU0RXLM5_1;
	wire w_dff_B_mXLpm9LL5_1;
	wire w_dff_B_QQvrlayg6_1;
	wire w_dff_B_7yNumaUC6_1;
	wire w_dff_B_g2vZiXYP5_1;
	wire w_dff_B_8FnJnD3z7_1;
	wire w_dff_B_8d4CFpGF3_1;
	wire w_dff_B_FZaX2W3d6_1;
	wire w_dff_B_Ba1mraEJ8_1;
	wire w_dff_B_CvJGr1j23_1;
	wire w_dff_B_VrLSQstI7_1;
	wire w_dff_B_yp0kKRyi6_1;
	wire w_dff_B_alNwLkmM0_1;
	wire w_dff_B_M1rMyHoL3_1;
	wire w_dff_B_T6NVnOqK7_1;
	wire w_dff_B_TKF9hkmS6_1;
	wire w_dff_B_DfttxFvS3_1;
	wire w_dff_B_hz3xGkkH4_1;
	wire w_dff_B_mlrtrj4I8_1;
	wire w_dff_B_Z9uRKsnt5_1;
	wire w_dff_B_tbdN8ecb3_1;
	wire w_dff_B_8vwSmKNJ9_1;
	wire w_dff_B_IioFGClq1_1;
	wire w_dff_B_P91aLeGR0_1;
	wire w_dff_B_72K5SKWg9_1;
	wire w_dff_B_gMB6IRLs1_1;
	wire w_dff_B_Z6f4XFcB3_1;
	wire w_dff_B_hfhOpRUK7_1;
	wire w_dff_B_xOxumTwj5_1;
	wire w_dff_B_0GcyFVx43_1;
	wire w_dff_B_uzSnaecV0_1;
	wire w_dff_B_WSTVPVVF3_1;
	wire w_dff_B_QVr6NXvU1_1;
	wire w_dff_B_2X7izOS41_1;
	wire w_dff_B_rkbMdsOO8_1;
	wire w_dff_B_yph8wovY1_1;
	wire w_dff_B_tzqPMpLH0_1;
	wire w_dff_B_4iMasuAT4_1;
	wire w_dff_B_7BewOAbz1_1;
	wire w_dff_B_0wCuhX9P9_1;
	wire w_dff_B_HxRmiiOV9_1;
	wire w_dff_B_Legzqtl65_1;
	wire w_dff_B_9i2TSU313_1;
	wire w_dff_B_ORN53I3K0_1;
	wire w_dff_B_8DFnl29K3_1;
	wire w_dff_B_eQXs7xZY4_1;
	wire w_dff_B_QWKKtUMY4_1;
	wire w_dff_B_Pu7APPQZ1_1;
	wire w_dff_B_pUrO5l0j5_1;
	wire w_dff_B_zAqgsTp33_1;
	wire w_dff_B_NeOthQYI5_1;
	wire w_dff_B_OFPMgZrs6_1;
	wire w_dff_B_5qdPJeJF5_1;
	wire w_dff_B_9YZ0tzTb7_1;
	wire w_dff_B_dxokdYOo3_1;
	wire w_dff_B_BAh8xJSH5_1;
	wire w_dff_B_wUKF8ogW1_1;
	wire w_dff_B_3cFsxSls8_1;
	wire w_dff_B_MJ8qJrJc7_1;
	wire w_dff_B_YJ9BY6258_1;
	wire w_dff_B_IbaBSp9K6_1;
	wire w_dff_B_gphZL0c48_1;
	wire w_dff_B_zjBEs5kK9_1;
	wire w_dff_B_RCtKRZoy9_1;
	wire w_dff_B_CWTtPHLv0_1;
	wire w_dff_B_9vygHb7i0_1;
	wire w_dff_B_zrbP7GxY7_1;
	wire w_dff_B_vlgOJ9V45_1;
	wire w_dff_B_lQdenUxA3_1;
	wire w_dff_B_T9S4j88q1_1;
	wire w_dff_B_YMHPHOGC7_1;
	wire w_dff_B_e3vPg3aK4_1;
	wire w_dff_B_3haVZqPq3_1;
	wire w_dff_B_XWeteEXP6_1;
	wire w_dff_B_smQYrNTu9_1;
	wire w_dff_B_ubSYQkAp4_1;
	wire w_dff_B_S1mvOlBs1_1;
	wire w_dff_B_sVsR5Bib1_1;
	wire w_dff_B_THBBGuER1_1;
	wire w_dff_B_Fvn1pcjV7_1;
	wire w_dff_B_6kjFu5kD2_1;
	wire w_dff_B_QQqIqfzG1_1;
	wire w_dff_B_JUYeebX73_1;
	wire w_dff_B_ZcZAQ4h83_1;
	wire w_dff_B_KasNIBlK6_1;
	wire w_dff_B_PxF00urH7_1;
	wire w_dff_B_AhfhLbtx1_1;
	wire w_dff_B_6jqm9QDu1_1;
	wire w_dff_B_RAzeX9Ee3_1;
	wire w_dff_B_h5ZmYzif9_1;
	wire w_dff_B_Gq98wQqv7_1;
	wire w_dff_B_LJPx6NS17_1;
	wire w_dff_B_4wHqYd5m9_1;
	wire w_dff_B_TzECuIlT0_1;
	wire w_dff_B_CYelCk5L1_1;
	wire w_dff_B_MJQcLT6M0_1;
	wire w_dff_B_ES7KtxQN2_1;
	wire w_dff_B_BqWfWFbi0_1;
	wire w_dff_B_07dyed016_1;
	wire w_dff_B_F5vh5ikl9_1;
	wire w_dff_B_pqau9lx39_1;
	wire w_dff_B_71rkZhAP6_1;
	wire w_dff_B_GhOmgY1E2_1;
	wire w_dff_B_suawknRD1_1;
	wire w_dff_B_J6ckBTzW4_1;
	wire w_dff_B_GWvrKgw21_1;
	wire w_dff_B_20TtFKlF8_1;
	wire w_dff_B_dguU4IQa4_1;
	wire w_dff_B_0Xx7iimN3_1;
	wire w_dff_B_UiQkJDS42_1;
	wire w_dff_B_KQYMATR73_1;
	wire w_dff_B_Tm6JEVns6_1;
	wire w_dff_B_QmP3Pabd6_1;
	wire w_dff_B_I3kkLVVQ0_1;
	wire w_dff_B_rs3vVlKB5_1;
	wire w_dff_B_Pe1iiYr60_1;
	wire w_dff_B_M7EI9SW90_0;
	wire w_dff_B_5DlrnuB45_0;
	wire w_dff_B_4NvbCU4G1_0;
	wire w_dff_B_ifBdqo8a5_0;
	wire w_dff_B_oAaGdQqR9_0;
	wire w_dff_B_IeYAlWuO9_0;
	wire w_dff_B_JqH1fp9I9_0;
	wire w_dff_B_P673onFb5_0;
	wire w_dff_B_AgSz4TSZ3_0;
	wire w_dff_B_OZ0h0jjA9_0;
	wire w_dff_B_xxaRuZgU2_0;
	wire w_dff_B_bPA1eVCN6_0;
	wire w_dff_B_QiiZuJe62_0;
	wire w_dff_B_rSHWIbpy0_0;
	wire w_dff_B_5nrxxgvh5_0;
	wire w_dff_B_ytaZtXJp0_0;
	wire w_dff_B_5RqGnWwl9_0;
	wire w_dff_B_PYHhmXPH4_0;
	wire w_dff_B_4eOcVJVv8_0;
	wire w_dff_B_wSv5OMIn7_0;
	wire w_dff_B_rCGn6ZpC6_0;
	wire w_dff_B_FDrzNFow4_0;
	wire w_dff_B_nM0r0Jkc4_0;
	wire w_dff_B_JZkn5b0e9_0;
	wire w_dff_B_n0IIdDsi3_0;
	wire w_dff_B_JYv0oRdD6_0;
	wire w_dff_B_tMe3Qlhx6_0;
	wire w_dff_B_YAvOovI92_0;
	wire w_dff_B_mhDkDj2e1_0;
	wire w_dff_B_iPZzOWWJ1_0;
	wire w_dff_B_oWM6jmUt7_0;
	wire w_dff_B_cN3zvUzP9_0;
	wire w_dff_B_Jd1DXDNY2_0;
	wire w_dff_B_ReW7hyrU9_0;
	wire w_dff_B_kPvfq4EU7_0;
	wire w_dff_B_eNJRRZPe3_0;
	wire w_dff_B_0JaJ4R4P9_0;
	wire w_dff_B_yQhDGsuU4_0;
	wire w_dff_B_whvYdmgG3_0;
	wire w_dff_B_sJQDvEHQ2_0;
	wire w_dff_B_hLcmAr003_0;
	wire w_dff_B_N5ZZWG9P9_0;
	wire w_dff_B_E9XpuREw2_0;
	wire w_dff_B_tHJtXSo34_0;
	wire w_dff_B_pvKd1m2w5_0;
	wire w_dff_B_unjXOp8p0_0;
	wire w_dff_B_ZI0RRKRl2_0;
	wire w_dff_B_CnP0slgD6_0;
	wire w_dff_B_Pu8KmmXN5_0;
	wire w_dff_B_IzNaHN1V0_0;
	wire w_dff_B_8ejwgIiy8_0;
	wire w_dff_B_maSwbOzT1_0;
	wire w_dff_B_HiyVQhUE9_0;
	wire w_dff_B_OreHujBm1_0;
	wire w_dff_B_snYMKc227_0;
	wire w_dff_B_hv0woxsA1_0;
	wire w_dff_B_mC0dDsO84_0;
	wire w_dff_B_gFIsGDk84_0;
	wire w_dff_B_A5aTERoy1_0;
	wire w_dff_B_2gLOA8Ld4_0;
	wire w_dff_B_IT5vkL4H7_0;
	wire w_dff_B_qO9ITuGd6_0;
	wire w_dff_B_1nPCrTZm5_0;
	wire w_dff_B_6iS57Xmq5_0;
	wire w_dff_B_YHJplSgl9_0;
	wire w_dff_B_12qGtThZ1_0;
	wire w_dff_B_NxXlxi6j0_0;
	wire w_dff_B_iVAxyb5X0_0;
	wire w_dff_B_kZAyKJ1V6_0;
	wire w_dff_B_CPMIU3Et0_0;
	wire w_dff_B_yKLMkLdr5_0;
	wire w_dff_B_t9ulnEnL3_0;
	wire w_dff_B_ZYEy1BOh6_0;
	wire w_dff_B_1eWsj6Xp4_0;
	wire w_dff_B_PNx1tVtz4_0;
	wire w_dff_B_25zsk5Pn9_0;
	wire w_dff_B_Kqqn8YoK4_0;
	wire w_dff_B_H6KRydry6_0;
	wire w_dff_B_Zbe0OBqx2_0;
	wire w_dff_B_h6ThyQlb0_0;
	wire w_dff_B_LDP8luwg1_0;
	wire w_dff_B_Rfes5znt0_0;
	wire w_dff_B_h0BAPlbY7_0;
	wire w_dff_B_2pwfBrSc6_0;
	wire w_dff_B_zIGcAts16_0;
	wire w_dff_B_WwPZX7ES5_0;
	wire w_dff_B_v3N7St3I6_0;
	wire w_dff_B_lpQCQZH77_0;
	wire w_dff_B_Zoxst3704_0;
	wire w_dff_B_T8aQEHVr2_0;
	wire w_dff_B_qxcsQPKH3_0;
	wire w_dff_B_WFv9DYoH8_0;
	wire w_dff_B_tWf3XB4i8_0;
	wire w_dff_B_iJS4LuBa1_0;
	wire w_dff_B_P2oTfjLT0_0;
	wire w_dff_B_V9TZ42Uf4_0;
	wire w_dff_B_JKBWP2Ai8_0;
	wire w_dff_B_UjaNzp175_0;
	wire w_dff_B_m9DS1XgK6_0;
	wire w_dff_B_CaNEwa7s6_0;
	wire w_dff_B_huh2ku8H8_0;
	wire w_dff_B_Z6mUNCq97_0;
	wire w_dff_B_znD4ty7R5_0;
	wire w_dff_B_TnCyVnkM8_0;
	wire w_dff_B_kNPdqaCW7_0;
	wire w_dff_B_nRrdxhvB4_0;
	wire w_dff_B_u4rFfE759_0;
	wire w_dff_B_jRJlZfOd8_0;
	wire w_dff_B_7SiybSqA8_0;
	wire w_dff_B_0oAT4Rev5_0;
	wire w_dff_B_s2gsltDL7_0;
	wire w_dff_B_Va5VyfBr5_0;
	wire w_dff_B_YEIBzdqU3_0;
	wire w_dff_B_1330L5tP0_0;
	wire w_dff_B_7DRwlRO77_0;
	wire w_dff_B_kLMAFHjd5_0;
	wire w_dff_B_YHtR4fi00_0;
	wire w_dff_B_Mva6TcQC3_1;
	wire w_dff_B_kokxEdVW1_1;
	wire w_dff_B_DuHvCeXp9_1;
	wire w_dff_B_8HTLUvlt4_1;
	wire w_dff_B_IVq4IGff9_1;
	wire w_dff_B_X4mKLp5N4_1;
	wire w_dff_B_KmwrLEB03_1;
	wire w_dff_B_0esGfP8z2_1;
	wire w_dff_B_f7vGlDzW6_1;
	wire w_dff_B_DasWWJJw4_1;
	wire w_dff_B_mWMed6LW1_1;
	wire w_dff_B_fOpm9S0e6_1;
	wire w_dff_B_QMMBpxF42_1;
	wire w_dff_B_rRAhMiLx1_1;
	wire w_dff_B_Iogz5Cyt4_1;
	wire w_dff_B_eMcL5tkk0_1;
	wire w_dff_B_5UlNxpAs9_1;
	wire w_dff_B_2jjWzCxk8_1;
	wire w_dff_B_9SLRow335_1;
	wire w_dff_B_7LXNU9WD0_1;
	wire w_dff_B_YPTKF3bv0_1;
	wire w_dff_B_8YfUqkGs4_1;
	wire w_dff_B_RvV3B9Lk6_1;
	wire w_dff_B_16YwknhO5_1;
	wire w_dff_B_pCxzE4MB2_1;
	wire w_dff_B_80BoNJFi1_1;
	wire w_dff_B_pm0YsuEi7_1;
	wire w_dff_B_jh7lPzj90_1;
	wire w_dff_B_XJpTwJ1N0_1;
	wire w_dff_B_TgmkPTjJ5_1;
	wire w_dff_B_MlefUiER5_1;
	wire w_dff_B_BQFQkRKn1_1;
	wire w_dff_B_uKilCTj05_1;
	wire w_dff_B_rfi7v14r4_1;
	wire w_dff_B_wOr8EqwB9_1;
	wire w_dff_B_Y5ha6kkK4_1;
	wire w_dff_B_agJMqJbA9_1;
	wire w_dff_B_7cWnK8Ja1_1;
	wire w_dff_B_lJyKqemu5_1;
	wire w_dff_B_gFAVYVfM6_1;
	wire w_dff_B_wpEhMsoK1_1;
	wire w_dff_B_pMpQUgLF2_1;
	wire w_dff_B_R5Emixij0_1;
	wire w_dff_B_gAskS9d85_1;
	wire w_dff_B_SO7QG9tp3_1;
	wire w_dff_B_0LAQqcji3_1;
	wire w_dff_B_wjK4LdHO2_1;
	wire w_dff_B_m3Z1pYuz1_1;
	wire w_dff_B_40pTdnTV4_1;
	wire w_dff_B_9cYSHblH7_1;
	wire w_dff_B_R0KXtrdP2_1;
	wire w_dff_B_haSwwdUt8_1;
	wire w_dff_B_vwQnEUg09_1;
	wire w_dff_B_IzzOXkwY4_1;
	wire w_dff_B_OxkcOqHu1_1;
	wire w_dff_B_oGgbXCnT8_1;
	wire w_dff_B_7AuRGt5N5_1;
	wire w_dff_B_5r4wPzZq0_1;
	wire w_dff_B_yJ5n5j3l9_1;
	wire w_dff_B_nFZjQded9_1;
	wire w_dff_B_dUut2OlH6_1;
	wire w_dff_B_oAvWXRvp2_1;
	wire w_dff_B_9eImSTrN9_1;
	wire w_dff_B_j3wGZEew6_1;
	wire w_dff_B_S52isB6i7_1;
	wire w_dff_B_5RxK6jmr7_1;
	wire w_dff_B_SGuEypJX3_1;
	wire w_dff_B_6HNUGjpl2_1;
	wire w_dff_B_X2BqJM3K4_1;
	wire w_dff_B_2LKZDNeI3_1;
	wire w_dff_B_QhYOYsAE4_1;
	wire w_dff_B_zuJZW8bC6_1;
	wire w_dff_B_idOx3eYX8_1;
	wire w_dff_B_7Tzfi5aE0_1;
	wire w_dff_B_Nee9REeW2_1;
	wire w_dff_B_a6PbQl1x4_1;
	wire w_dff_B_kpwezgEs1_1;
	wire w_dff_B_WKnQEFf81_1;
	wire w_dff_B_tN7muEOo9_1;
	wire w_dff_B_pj5Q2XNi2_1;
	wire w_dff_B_glfGUBZ16_1;
	wire w_dff_B_nXjSbwsS7_1;
	wire w_dff_B_Gz2BeENo0_1;
	wire w_dff_B_8nUXdlyh2_1;
	wire w_dff_B_ECD4Emfb9_1;
	wire w_dff_B_1XgQn9YC1_1;
	wire w_dff_B_lUQjkxGn7_1;
	wire w_dff_B_qUO7qdcq1_1;
	wire w_dff_B_ZwrzRpIa0_1;
	wire w_dff_B_r2zxWOiQ3_1;
	wire w_dff_B_wjrD4Gba7_1;
	wire w_dff_B_omgaa8xX0_1;
	wire w_dff_B_vpfARLRc8_1;
	wire w_dff_B_fFrIurs99_1;
	wire w_dff_B_oO9qGIbb9_1;
	wire w_dff_B_kq1FULtz0_1;
	wire w_dff_B_vzduoSy73_1;
	wire w_dff_B_CSU5Exqh4_1;
	wire w_dff_B_eGVwxzAz7_1;
	wire w_dff_B_NhGUpUZd7_1;
	wire w_dff_B_Ymc7dSyE2_1;
	wire w_dff_B_3aAy86DJ0_1;
	wire w_dff_B_HLeWyBgG7_1;
	wire w_dff_B_k9kLOO4a2_1;
	wire w_dff_B_qEvwrYGp8_1;
	wire w_dff_B_P4oizCHC4_1;
	wire w_dff_B_MvLDE62y9_1;
	wire w_dff_B_c8t4eMk40_1;
	wire w_dff_B_ST0q4Qjd2_1;
	wire w_dff_B_XxBlAudr6_1;
	wire w_dff_B_YGBlSZ3u7_1;
	wire w_dff_B_7Z2MS1fk0_1;
	wire w_dff_B_drTDZiCu1_1;
	wire w_dff_B_3iG0t9it0_1;
	wire w_dff_B_y9BNTbnt8_1;
	wire w_dff_B_0nN0BSNX5_1;
	wire w_dff_B_CEcVRHjZ2_0;
	wire w_dff_B_rtlwDItD9_0;
	wire w_dff_B_of6DTMrQ5_0;
	wire w_dff_B_aGCFd8mm2_0;
	wire w_dff_B_yZyw2owQ2_0;
	wire w_dff_B_Dlo29GBj3_0;
	wire w_dff_B_zbDTd6015_0;
	wire w_dff_B_eR62aRzx5_0;
	wire w_dff_B_PZtNmySa7_0;
	wire w_dff_B_Rfo3o5cV2_0;
	wire w_dff_B_uSCRDwjQ9_0;
	wire w_dff_B_ctbF1Ulq7_0;
	wire w_dff_B_D07dR8wm2_0;
	wire w_dff_B_XaUGYvOY0_0;
	wire w_dff_B_rVRna2Hg5_0;
	wire w_dff_B_xJHVUlZX9_0;
	wire w_dff_B_G8boljKA9_0;
	wire w_dff_B_d1IG8QGg3_0;
	wire w_dff_B_sr4Fp0DC8_0;
	wire w_dff_B_AQh94kD40_0;
	wire w_dff_B_Lp8ee4nw7_0;
	wire w_dff_B_HYqQiyx82_0;
	wire w_dff_B_aQcdx7hr4_0;
	wire w_dff_B_S2Wl7Q1L0_0;
	wire w_dff_B_nWgaLhR66_0;
	wire w_dff_B_aXF9oQJA9_0;
	wire w_dff_B_24trkB455_0;
	wire w_dff_B_I1UaNswh3_0;
	wire w_dff_B_kBbz9s5V5_0;
	wire w_dff_B_OaRGEu4p4_0;
	wire w_dff_B_3jpsfhIq4_0;
	wire w_dff_B_hb446n6I6_0;
	wire w_dff_B_vD5iaqfe1_0;
	wire w_dff_B_dbx7uHRZ9_0;
	wire w_dff_B_2hUrxHKo4_0;
	wire w_dff_B_hGpOnTPN3_0;
	wire w_dff_B_O15gnHGa9_0;
	wire w_dff_B_dKN9ee4Y3_0;
	wire w_dff_B_yTcj7qUT3_0;
	wire w_dff_B_ib5h5OsW0_0;
	wire w_dff_B_ddup17tU2_0;
	wire w_dff_B_2UOiuz2B8_0;
	wire w_dff_B_LUjfoTF04_0;
	wire w_dff_B_GtbWfExF2_0;
	wire w_dff_B_HBYounN53_0;
	wire w_dff_B_mzyMEDLv4_0;
	wire w_dff_B_MbtIKZL59_0;
	wire w_dff_B_Pj03Arrf8_0;
	wire w_dff_B_IyBTYlXi1_0;
	wire w_dff_B_8FEiPlDW9_0;
	wire w_dff_B_pqfQ7txp5_0;
	wire w_dff_B_dtxSjQuc6_0;
	wire w_dff_B_wifl28q81_0;
	wire w_dff_B_SHW4TUzh0_0;
	wire w_dff_B_selpxYZT2_0;
	wire w_dff_B_VBGAhItr7_0;
	wire w_dff_B_HW5IhkaJ7_0;
	wire w_dff_B_iQMTKuhs4_0;
	wire w_dff_B_TqCDsnul8_0;
	wire w_dff_B_GBPh6MQS4_0;
	wire w_dff_B_QI3oEd8p6_0;
	wire w_dff_B_LfXWihqg3_0;
	wire w_dff_B_iM4xOC2P8_0;
	wire w_dff_B_q8o5KloS6_0;
	wire w_dff_B_Xtx4G3vh9_0;
	wire w_dff_B_OlsHckU21_0;
	wire w_dff_B_fiU3edQc3_0;
	wire w_dff_B_TfRCJYOG4_0;
	wire w_dff_B_im0ifTAi2_0;
	wire w_dff_B_G0vFep251_0;
	wire w_dff_B_RGRYrxUn1_0;
	wire w_dff_B_hC79WNhS4_0;
	wire w_dff_B_dZ5dLyHX5_0;
	wire w_dff_B_52nLrKKd8_0;
	wire w_dff_B_4bzjMXpP9_0;
	wire w_dff_B_U0vtRxJ48_0;
	wire w_dff_B_TJG1b6v82_0;
	wire w_dff_B_AQV777Rz8_0;
	wire w_dff_B_20FlKqlq1_0;
	wire w_dff_B_pAha6tjz5_0;
	wire w_dff_B_PvD6pQJi1_0;
	wire w_dff_B_hN9yoSho4_0;
	wire w_dff_B_yKt2x2n35_0;
	wire w_dff_B_fzOSd82d7_0;
	wire w_dff_B_nxMiRQsR4_0;
	wire w_dff_B_jWjuFFjz3_0;
	wire w_dff_B_QUhzDHYV7_0;
	wire w_dff_B_UhNmhSVy5_0;
	wire w_dff_B_FWBfXhrK8_0;
	wire w_dff_B_8b2KP5PT2_0;
	wire w_dff_B_WnWnmiv69_0;
	wire w_dff_B_QJWQ2UHw3_0;
	wire w_dff_B_RhzAqGUo2_0;
	wire w_dff_B_objedPYf6_0;
	wire w_dff_B_6keo17Jm9_0;
	wire w_dff_B_e7wX5awP2_0;
	wire w_dff_B_3m9OCgPF3_0;
	wire w_dff_B_4N8ppNo25_0;
	wire w_dff_B_FTJBg4vB8_0;
	wire w_dff_B_5vL8vtHN2_0;
	wire w_dff_B_jTacgAvb5_0;
	wire w_dff_B_KxjvUQzK3_0;
	wire w_dff_B_mtt3OAM07_0;
	wire w_dff_B_JNEE5kdi4_0;
	wire w_dff_B_qZNb5GWQ4_0;
	wire w_dff_B_w9DRzh0n4_0;
	wire w_dff_B_YHspHjoT1_0;
	wire w_dff_B_2BPQpjbO1_0;
	wire w_dff_B_kA9YYPZO5_0;
	wire w_dff_B_vtBo1Mg96_0;
	wire w_dff_B_6X3X32i51_0;
	wire w_dff_B_mMX3SkrN1_0;
	wire w_dff_B_ImCUCeM42_0;
	wire w_dff_B_GTZSpFw73_0;
	wire w_dff_B_QRImenJk5_0;
	wire w_dff_B_k7K9XKQ61_0;
	wire w_dff_B_J6E6OeuB3_1;
	wire w_dff_B_ekydRNRm6_1;
	wire w_dff_B_suaHM4gB9_1;
	wire w_dff_B_5EltmYY89_1;
	wire w_dff_B_lD71pSi28_1;
	wire w_dff_B_u8T8jq7S0_1;
	wire w_dff_B_NE17rn8J7_1;
	wire w_dff_B_yBgVfDsw0_1;
	wire w_dff_B_AATsKAgO0_1;
	wire w_dff_B_GiCsjwu04_1;
	wire w_dff_B_qlHzmWSj8_1;
	wire w_dff_B_Gx5ECXYr8_1;
	wire w_dff_B_poKQ7djP9_1;
	wire w_dff_B_vTuWXpzW1_1;
	wire w_dff_B_aims8asC2_1;
	wire w_dff_B_ET657AIj5_1;
	wire w_dff_B_ahSjjnQt0_1;
	wire w_dff_B_5Nle80dz1_1;
	wire w_dff_B_tPvJuUk45_1;
	wire w_dff_B_BVn2FPyB8_1;
	wire w_dff_B_HlVO66GQ5_1;
	wire w_dff_B_u0lvtJJE5_1;
	wire w_dff_B_RVNTHlCb6_1;
	wire w_dff_B_SuN8QHy73_1;
	wire w_dff_B_TUfV9tun7_1;
	wire w_dff_B_E6WB9u2o6_1;
	wire w_dff_B_KUEmSiAk1_1;
	wire w_dff_B_BQQkszUf4_1;
	wire w_dff_B_BtVFA8sJ2_1;
	wire w_dff_B_crFtoYkU7_1;
	wire w_dff_B_DN9HcD6v8_1;
	wire w_dff_B_oXzvce9N8_1;
	wire w_dff_B_sQSF0xzh9_1;
	wire w_dff_B_CXs5HuYa5_1;
	wire w_dff_B_vbxfDsLv8_1;
	wire w_dff_B_NBisfOiF6_1;
	wire w_dff_B_SjS2hqwN4_1;
	wire w_dff_B_pCJ7e4FS0_1;
	wire w_dff_B_zTB39jfD1_1;
	wire w_dff_B_c9y4j0191_1;
	wire w_dff_B_VQULySjX2_1;
	wire w_dff_B_2RLTwiEG8_1;
	wire w_dff_B_xP8l1tt87_1;
	wire w_dff_B_qId6cRTo7_1;
	wire w_dff_B_2STgaVi67_1;
	wire w_dff_B_KDy1Bz6A2_1;
	wire w_dff_B_IpbddDJP9_1;
	wire w_dff_B_P0XRYMY91_1;
	wire w_dff_B_RHvkn7l22_1;
	wire w_dff_B_08w6AZx02_1;
	wire w_dff_B_5pmxiRyR9_1;
	wire w_dff_B_L6DvscGH8_1;
	wire w_dff_B_pupEmGhs4_1;
	wire w_dff_B_DeJ34ZzK6_1;
	wire w_dff_B_GIgX8GWm1_1;
	wire w_dff_B_xCUqtNJg5_1;
	wire w_dff_B_Jcg7lNh85_1;
	wire w_dff_B_EqrXVh3y8_1;
	wire w_dff_B_LbTHXGcd5_1;
	wire w_dff_B_FjYwjX1l2_1;
	wire w_dff_B_Wtk5BMNj5_1;
	wire w_dff_B_5yVe6hZN7_1;
	wire w_dff_B_56GWUrSm9_1;
	wire w_dff_B_8R9OaSo16_1;
	wire w_dff_B_81DG4xZv0_1;
	wire w_dff_B_hvsfi7SJ6_1;
	wire w_dff_B_HLXjHnPc8_1;
	wire w_dff_B_xDhUz0eA5_1;
	wire w_dff_B_23oKKmbI4_1;
	wire w_dff_B_2emqIVQY5_1;
	wire w_dff_B_JKcatsSO6_1;
	wire w_dff_B_LghcBRfS2_1;
	wire w_dff_B_JpVDBtyl4_1;
	wire w_dff_B_pA2MZHhR0_1;
	wire w_dff_B_JtLkvqGU5_1;
	wire w_dff_B_fzcsPpco2_1;
	wire w_dff_B_aEjRS6Me4_1;
	wire w_dff_B_SXLNZ0VT1_1;
	wire w_dff_B_AMj6Dc9L6_1;
	wire w_dff_B_pLuib1cd8_1;
	wire w_dff_B_1JDqF20i7_1;
	wire w_dff_B_kGF785tx7_1;
	wire w_dff_B_i3F51tK17_1;
	wire w_dff_B_EoSNBCoy9_1;
	wire w_dff_B_L6UfDWSe7_1;
	wire w_dff_B_iePPLRq35_1;
	wire w_dff_B_qD8wQudE5_1;
	wire w_dff_B_MxFvXjqI2_1;
	wire w_dff_B_ghFUSEBb1_1;
	wire w_dff_B_nsOANQZh1_1;
	wire w_dff_B_DE0PeJcg4_1;
	wire w_dff_B_i4sfX0Pi6_1;
	wire w_dff_B_S3nrAXFr5_1;
	wire w_dff_B_u6tmZq4Y7_1;
	wire w_dff_B_pyCIjXkf4_1;
	wire w_dff_B_QnA1DRYy5_1;
	wire w_dff_B_9MMvWxuV1_1;
	wire w_dff_B_sxf07jmx3_1;
	wire w_dff_B_I6aAMcYr7_1;
	wire w_dff_B_TOH2blfR3_1;
	wire w_dff_B_sJRHqjKW8_1;
	wire w_dff_B_DMXGwRS08_1;
	wire w_dff_B_3ppe9bG11_1;
	wire w_dff_B_GVRlRWhZ4_1;
	wire w_dff_B_SEb04kH37_1;
	wire w_dff_B_V6SJyvHn0_1;
	wire w_dff_B_brRxbKFR7_1;
	wire w_dff_B_ME5l3UJt3_1;
	wire w_dff_B_mvUyxB3H1_1;
	wire w_dff_B_Wa3rStW03_1;
	wire w_dff_B_P9Er4em07_1;
	wire w_dff_B_TUvV9uPf5_1;
	wire w_dff_B_XqHKqY9F6_1;
	wire w_dff_B_Calt62xu3_1;
	wire w_dff_B_DmeXqhOy3_1;
	wire w_dff_B_pfbTqXXG1_0;
	wire w_dff_B_Uw8Pseyl7_0;
	wire w_dff_B_7fLCgk2S3_0;
	wire w_dff_B_MmQqyFOf1_0;
	wire w_dff_B_itpXekh08_0;
	wire w_dff_B_h23wqXfC7_0;
	wire w_dff_B_DOUJuvoL0_0;
	wire w_dff_B_2j34fPCF0_0;
	wire w_dff_B_QHYXr5C66_0;
	wire w_dff_B_ABtQpvYU0_0;
	wire w_dff_B_nL1OYnUx2_0;
	wire w_dff_B_XzTRCcCo3_0;
	wire w_dff_B_b9FQ16xm8_0;
	wire w_dff_B_4vLICp688_0;
	wire w_dff_B_Yv3JoQzG6_0;
	wire w_dff_B_QQNqunm91_0;
	wire w_dff_B_pZb2KrV00_0;
	wire w_dff_B_Q4ztJBHL6_0;
	wire w_dff_B_SmBl1Bcb9_0;
	wire w_dff_B_hFgz3um19_0;
	wire w_dff_B_tOH1vVKL3_0;
	wire w_dff_B_5Ws8UyBA0_0;
	wire w_dff_B_HszMZe0m8_0;
	wire w_dff_B_MVLtSCjV3_0;
	wire w_dff_B_bOnyNOFe7_0;
	wire w_dff_B_fkoJ5Jjw0_0;
	wire w_dff_B_Q90IWg9Q2_0;
	wire w_dff_B_KN1fh3TJ9_0;
	wire w_dff_B_rqRohDcD8_0;
	wire w_dff_B_aH8b8GyH8_0;
	wire w_dff_B_qrJMhkEn0_0;
	wire w_dff_B_gpbDAU8f9_0;
	wire w_dff_B_rPBKxsxN2_0;
	wire w_dff_B_MjESDd3Q7_0;
	wire w_dff_B_RycHrpEV1_0;
	wire w_dff_B_nhS8BPsd1_0;
	wire w_dff_B_ZIVdhz7i0_0;
	wire w_dff_B_vjqSo6t65_0;
	wire w_dff_B_v4lwbTeb6_0;
	wire w_dff_B_xXxxeBEB6_0;
	wire w_dff_B_xX9ZufBE2_0;
	wire w_dff_B_WYln5OOG2_0;
	wire w_dff_B_TQay20PG3_0;
	wire w_dff_B_9EfsfU6D7_0;
	wire w_dff_B_bEE8t4SK3_0;
	wire w_dff_B_vWmN97LW1_0;
	wire w_dff_B_m5khuecM8_0;
	wire w_dff_B_shrIfdo19_0;
	wire w_dff_B_Q7YSl3iw1_0;
	wire w_dff_B_m0afCjyx2_0;
	wire w_dff_B_s8DUX3p31_0;
	wire w_dff_B_eVwcYOHQ0_0;
	wire w_dff_B_sfgFyjIt5_0;
	wire w_dff_B_LhS3JG1z7_0;
	wire w_dff_B_bSNws27A1_0;
	wire w_dff_B_11pDVKuv4_0;
	wire w_dff_B_wV4uZ5Sm8_0;
	wire w_dff_B_oV9dxKqX1_0;
	wire w_dff_B_VBE0HBhG1_0;
	wire w_dff_B_6fngLBZU7_0;
	wire w_dff_B_VQwpoh080_0;
	wire w_dff_B_YEKvAFMu1_0;
	wire w_dff_B_cbIx5wA74_0;
	wire w_dff_B_t0Hsi3QP9_0;
	wire w_dff_B_eJSab3Vq4_0;
	wire w_dff_B_rie5fYW03_0;
	wire w_dff_B_vmrkeYnu7_0;
	wire w_dff_B_2oe3zhVW3_0;
	wire w_dff_B_DLgEEcHe4_0;
	wire w_dff_B_Wgfequ1T0_0;
	wire w_dff_B_gtK7CO3B1_0;
	wire w_dff_B_freIDPdd8_0;
	wire w_dff_B_bKzCqqpN1_0;
	wire w_dff_B_MAeA0RML4_0;
	wire w_dff_B_YQAMhp5n0_0;
	wire w_dff_B_wapMKsOJ8_0;
	wire w_dff_B_Lo3ItOgO2_0;
	wire w_dff_B_pXkKd7Kz1_0;
	wire w_dff_B_b5IQTnp33_0;
	wire w_dff_B_D9rd5KXP6_0;
	wire w_dff_B_lkMRwUoy4_0;
	wire w_dff_B_UOZ77J6s6_0;
	wire w_dff_B_4dmaQakO5_0;
	wire w_dff_B_HfHV0p9z3_0;
	wire w_dff_B_2h1MaLiM2_0;
	wire w_dff_B_RU2aNEET8_0;
	wire w_dff_B_l5c4V3iN3_0;
	wire w_dff_B_w1tZACVk8_0;
	wire w_dff_B_Fl7D7wAm4_0;
	wire w_dff_B_pshJjRMi3_0;
	wire w_dff_B_aQv0bGNk7_0;
	wire w_dff_B_ae7OEHZp0_0;
	wire w_dff_B_kvtzmL0r4_0;
	wire w_dff_B_oDI3aSF29_0;
	wire w_dff_B_mqkx78xk3_0;
	wire w_dff_B_0seXyGFE9_0;
	wire w_dff_B_lR7n1kre2_0;
	wire w_dff_B_q9sw8fpB1_0;
	wire w_dff_B_pDiftYiS6_0;
	wire w_dff_B_4Mik9kMM2_0;
	wire w_dff_B_2Gw5om041_0;
	wire w_dff_B_0xMzr56d5_0;
	wire w_dff_B_Bc3aEgHa3_0;
	wire w_dff_B_Jr5rAzQK1_0;
	wire w_dff_B_Z0Qj2PC29_0;
	wire w_dff_B_5Iw6WGuZ5_0;
	wire w_dff_B_M4XffYyu2_0;
	wire w_dff_B_sOSJEZFe8_0;
	wire w_dff_B_Fiym9kQc9_0;
	wire w_dff_B_4gkEbQSM5_0;
	wire w_dff_B_ekHpHopO6_0;
	wire w_dff_B_t9WZNTWu4_0;
	wire w_dff_B_tAY2Yj6h5_0;
	wire w_dff_B_EYJkHRuW1_0;
	wire w_dff_B_ihbYCldo3_0;
	wire w_dff_B_MCq281UY6_1;
	wire w_dff_B_1ADqnZNQ4_1;
	wire w_dff_B_7t9HJ7sx2_1;
	wire w_dff_B_tkwL7lN16_1;
	wire w_dff_B_LS2fiSKH2_1;
	wire w_dff_B_TcM1PmAn2_1;
	wire w_dff_B_4uTXGvEq7_1;
	wire w_dff_B_dWw8OsXj0_1;
	wire w_dff_B_JbviCirz7_1;
	wire w_dff_B_aYarJ7CU1_1;
	wire w_dff_B_FSEIA4MW4_1;
	wire w_dff_B_aoJppHH29_1;
	wire w_dff_B_QLFHExor6_1;
	wire w_dff_B_zFQXqWL58_1;
	wire w_dff_B_7QDYzYvG2_1;
	wire w_dff_B_Mp43LeOg9_1;
	wire w_dff_B_F1SHhpCQ7_1;
	wire w_dff_B_VQv64JSq9_1;
	wire w_dff_B_3wJaWl3d6_1;
	wire w_dff_B_B1q10AOM0_1;
	wire w_dff_B_clg6xez41_1;
	wire w_dff_B_xDt5lsgj7_1;
	wire w_dff_B_8pKmFt6G3_1;
	wire w_dff_B_kmhcdLiB8_1;
	wire w_dff_B_PyKYIiaX0_1;
	wire w_dff_B_d0BVUFZ00_1;
	wire w_dff_B_JZeDEizN3_1;
	wire w_dff_B_6V9OAOSy1_1;
	wire w_dff_B_AOGEX5kr0_1;
	wire w_dff_B_cl58WqLZ2_1;
	wire w_dff_B_bzBy4IcZ8_1;
	wire w_dff_B_D3X6rZeS0_1;
	wire w_dff_B_cAPbxwEv0_1;
	wire w_dff_B_rhVk8whC4_1;
	wire w_dff_B_mhBkypJF1_1;
	wire w_dff_B_rTK8PBFd5_1;
	wire w_dff_B_8YIYuS5L0_1;
	wire w_dff_B_d7sc9C9q5_1;
	wire w_dff_B_AEfYuPVR1_1;
	wire w_dff_B_1mAkaiIM9_1;
	wire w_dff_B_1dwby9fs1_1;
	wire w_dff_B_6zeCK66Z0_1;
	wire w_dff_B_ScERKzgl5_1;
	wire w_dff_B_vIYE3bUe5_1;
	wire w_dff_B_kIQ57ik54_1;
	wire w_dff_B_hVvEonaG5_1;
	wire w_dff_B_PcC3HCUZ7_1;
	wire w_dff_B_uAN9qSbH8_1;
	wire w_dff_B_v2YTIsda9_1;
	wire w_dff_B_iAVuv22D1_1;
	wire w_dff_B_d1gWu6fs3_1;
	wire w_dff_B_vpO54gNf1_1;
	wire w_dff_B_2e7ZQvDb0_1;
	wire w_dff_B_mx0LxQZu7_1;
	wire w_dff_B_0Ugtxr3R0_1;
	wire w_dff_B_1WfTxDNM8_1;
	wire w_dff_B_5HYuIW3Y0_1;
	wire w_dff_B_l6t5TALj6_1;
	wire w_dff_B_GzfykcJo7_1;
	wire w_dff_B_JGt70JuB2_1;
	wire w_dff_B_AdA6CQ5C8_1;
	wire w_dff_B_ykauX71l3_1;
	wire w_dff_B_A1KMzE375_1;
	wire w_dff_B_C60JWqCY9_1;
	wire w_dff_B_guAiUpl23_1;
	wire w_dff_B_Qgnwv9a00_1;
	wire w_dff_B_wp7I8PDh1_1;
	wire w_dff_B_PGq0nBXZ0_1;
	wire w_dff_B_Jt5JYBMu5_1;
	wire w_dff_B_aVZHfeaP9_1;
	wire w_dff_B_uT9UZBIX0_1;
	wire w_dff_B_L5Bx4XHE3_1;
	wire w_dff_B_T9MpUjrF1_1;
	wire w_dff_B_btAq2qi01_1;
	wire w_dff_B_nyAcjzIt9_1;
	wire w_dff_B_EBQj51um8_1;
	wire w_dff_B_eoCRFH6e6_1;
	wire w_dff_B_QM9cp9qm2_1;
	wire w_dff_B_MSkuuZ4p9_1;
	wire w_dff_B_crHZNiH82_1;
	wire w_dff_B_Y3HQ5Wur3_1;
	wire w_dff_B_0SguyIlg0_1;
	wire w_dff_B_06qyFdKf7_1;
	wire w_dff_B_6xfsC01k5_1;
	wire w_dff_B_VBOUQcis4_1;
	wire w_dff_B_crKgyBc98_1;
	wire w_dff_B_mCFwTzhf3_1;
	wire w_dff_B_XuCysnJ71_1;
	wire w_dff_B_iLbXeH9p5_1;
	wire w_dff_B_FwauJUrI0_1;
	wire w_dff_B_iB5XbIjn2_1;
	wire w_dff_B_lSJMyNrK1_1;
	wire w_dff_B_WsG7DlL11_1;
	wire w_dff_B_VUxvO5sy1_1;
	wire w_dff_B_Eypraqwc0_1;
	wire w_dff_B_66VSaaGL4_1;
	wire w_dff_B_cAtCcmj90_1;
	wire w_dff_B_Lh9aLFRP8_1;
	wire w_dff_B_Hh59ncTe1_1;
	wire w_dff_B_5KD1EUHe7_1;
	wire w_dff_B_yRZwIymy7_1;
	wire w_dff_B_Gpc3FdUr1_1;
	wire w_dff_B_ZdtaE59g7_1;
	wire w_dff_B_uJ1qSNMa2_1;
	wire w_dff_B_Ipw2d4wE4_1;
	wire w_dff_B_1SY2ypEI3_1;
	wire w_dff_B_nUFQeGhJ8_1;
	wire w_dff_B_HllRApmp6_1;
	wire w_dff_B_Th2DnWdp4_1;
	wire w_dff_B_ZsBjt1bw8_1;
	wire w_dff_B_vDC3FAL36_1;
	wire w_dff_B_dBiYiSsG8_1;
	wire w_dff_B_N3sp0qOL9_1;
	wire w_dff_B_SjyTVPLT6_1;
	wire w_dff_B_rg3QJQk22_0;
	wire w_dff_B_Nx6dgmj31_0;
	wire w_dff_B_KysPl3gz9_0;
	wire w_dff_B_SeUWHHwM7_0;
	wire w_dff_B_eGxZdXiI3_0;
	wire w_dff_B_Ep13Dq9T0_0;
	wire w_dff_B_ceXWccHN8_0;
	wire w_dff_B_zj6XrN4j8_0;
	wire w_dff_B_gMo14vJs2_0;
	wire w_dff_B_PDxzq8wM0_0;
	wire w_dff_B_K4PqtKp17_0;
	wire w_dff_B_B7TEkhld6_0;
	wire w_dff_B_jcJlavc00_0;
	wire w_dff_B_NnIjIV0h6_0;
	wire w_dff_B_6Fdzq0SK4_0;
	wire w_dff_B_l1raEnt12_0;
	wire w_dff_B_aDh62mhu6_0;
	wire w_dff_B_7Ee6opFT4_0;
	wire w_dff_B_siN5GXkT0_0;
	wire w_dff_B_b6AujLj70_0;
	wire w_dff_B_kXQa8VgV0_0;
	wire w_dff_B_z3JHWaLb1_0;
	wire w_dff_B_k3kLrxQj5_0;
	wire w_dff_B_Bwpn8EZg4_0;
	wire w_dff_B_c0DkvoDH8_0;
	wire w_dff_B_lflksyiR1_0;
	wire w_dff_B_U5P7Atke3_0;
	wire w_dff_B_NjVlTxqN8_0;
	wire w_dff_B_LtIpXpqa0_0;
	wire w_dff_B_JeA7Omf62_0;
	wire w_dff_B_hkxHifVD3_0;
	wire w_dff_B_1InYddIc5_0;
	wire w_dff_B_YbkFbB3G2_0;
	wire w_dff_B_bWMHe5lm3_0;
	wire w_dff_B_brMV1ppe7_0;
	wire w_dff_B_168MpKru2_0;
	wire w_dff_B_7HhTAQmD7_0;
	wire w_dff_B_aMaKUyGa1_0;
	wire w_dff_B_KYvt7k1M0_0;
	wire w_dff_B_eDN03dgm5_0;
	wire w_dff_B_5IxD8TV83_0;
	wire w_dff_B_dcqs8CCV5_0;
	wire w_dff_B_oDmOby2X9_0;
	wire w_dff_B_c6WqCTZd7_0;
	wire w_dff_B_acMX1Wc62_0;
	wire w_dff_B_6PQFdLeR0_0;
	wire w_dff_B_uhdn1nIl4_0;
	wire w_dff_B_8LyOA8hz0_0;
	wire w_dff_B_uNcXXOMv4_0;
	wire w_dff_B_3J9Fc0WC8_0;
	wire w_dff_B_3zEPpAuD4_0;
	wire w_dff_B_1k8uGg8o9_0;
	wire w_dff_B_JmP4pRMn8_0;
	wire w_dff_B_ue8z7mek9_0;
	wire w_dff_B_ObduV78a6_0;
	wire w_dff_B_13KbV9xF6_0;
	wire w_dff_B_Kx3hxUf32_0;
	wire w_dff_B_ZLSlyOH09_0;
	wire w_dff_B_M2jtz1wW7_0;
	wire w_dff_B_0Ko6pMOz6_0;
	wire w_dff_B_hkrtPrUb0_0;
	wire w_dff_B_kL9ZBm5j1_0;
	wire w_dff_B_mMhx6LXN6_0;
	wire w_dff_B_4bl9Za4H4_0;
	wire w_dff_B_3sapSiPS0_0;
	wire w_dff_B_KhuvoFix5_0;
	wire w_dff_B_lMUXr4I70_0;
	wire w_dff_B_f6r8Q5kc6_0;
	wire w_dff_B_oLrwJps75_0;
	wire w_dff_B_t9Iu0MLT7_0;
	wire w_dff_B_sez2YKZZ9_0;
	wire w_dff_B_NamGkoJa6_0;
	wire w_dff_B_xBEy1UkH8_0;
	wire w_dff_B_FkU27wbF6_0;
	wire w_dff_B_pBSIRIN01_0;
	wire w_dff_B_9nAlsUlr3_0;
	wire w_dff_B_u4rYNDtK3_0;
	wire w_dff_B_PSnlgtFe9_0;
	wire w_dff_B_kkT2CKVd4_0;
	wire w_dff_B_GPuOuC477_0;
	wire w_dff_B_QVnjppW31_0;
	wire w_dff_B_KVxzluwI4_0;
	wire w_dff_B_4luu63Vb9_0;
	wire w_dff_B_TiySji0B7_0;
	wire w_dff_B_Px9S1YhM1_0;
	wire w_dff_B_rAMLmSKL9_0;
	wire w_dff_B_tY4ONek58_0;
	wire w_dff_B_8PiApWfS9_0;
	wire w_dff_B_N3vIpLre2_0;
	wire w_dff_B_Cr822LdL2_0;
	wire w_dff_B_6oH8S5ZE0_0;
	wire w_dff_B_f1r3VukZ1_0;
	wire w_dff_B_10cwXiW89_0;
	wire w_dff_B_5xQYjxiu8_0;
	wire w_dff_B_QUlRPTPT1_0;
	wire w_dff_B_umu8oH3l7_0;
	wire w_dff_B_xDl0uCko9_0;
	wire w_dff_B_wldbdp9X1_0;
	wire w_dff_B_DEzZXAY44_0;
	wire w_dff_B_fgFgXz0K2_0;
	wire w_dff_B_TJfmdXyR9_0;
	wire w_dff_B_jITTrzJr3_0;
	wire w_dff_B_dfkGlCKW3_0;
	wire w_dff_B_2HsMWCV05_0;
	wire w_dff_B_IGnLiNoR8_0;
	wire w_dff_B_Ee0N77Yf4_0;
	wire w_dff_B_2yz6TJGX7_0;
	wire w_dff_B_B35LWGEU2_0;
	wire w_dff_B_CQUcic3R1_0;
	wire w_dff_B_T7Gd17DH7_0;
	wire w_dff_B_ujDnUcL90_0;
	wire w_dff_B_MNUzXlcS1_0;
	wire w_dff_B_niRhq5lk6_0;
	wire w_dff_B_ImrDGPBo9_0;
	wire w_dff_B_3YQA7GhO9_1;
	wire w_dff_B_7EGcvmRq3_1;
	wire w_dff_B_pUnIl0Xh3_1;
	wire w_dff_B_5gwzeTxg7_1;
	wire w_dff_B_6jaL3z8x1_1;
	wire w_dff_B_NvKWCXoq0_1;
	wire w_dff_B_znCzwP0g0_1;
	wire w_dff_B_cbogA8Uf5_1;
	wire w_dff_B_s9dFUFog4_1;
	wire w_dff_B_B9SRpaRN6_1;
	wire w_dff_B_nCnhwQNR3_1;
	wire w_dff_B_FOYIMpm94_1;
	wire w_dff_B_M6mVhZ1P9_1;
	wire w_dff_B_KdElwcez9_1;
	wire w_dff_B_yQ7FiiUG3_1;
	wire w_dff_B_vq1MESMN7_1;
	wire w_dff_B_uRYvc69a5_1;
	wire w_dff_B_FurXDm5T5_1;
	wire w_dff_B_YZp21Yuy0_1;
	wire w_dff_B_d6l3VUG36_1;
	wire w_dff_B_fcZjSejq7_1;
	wire w_dff_B_NNZYOxKS1_1;
	wire w_dff_B_spvH7CPH3_1;
	wire w_dff_B_I2keuj8g4_1;
	wire w_dff_B_hdTPNeFH5_1;
	wire w_dff_B_3uxEPy1t5_1;
	wire w_dff_B_hdaFrKyw2_1;
	wire w_dff_B_7CmvGMNf7_1;
	wire w_dff_B_IQOONsFh7_1;
	wire w_dff_B_VtDU580u3_1;
	wire w_dff_B_FSdbyO547_1;
	wire w_dff_B_AVrF9Nqd9_1;
	wire w_dff_B_ETEiR65W2_1;
	wire w_dff_B_j3AUtkRy7_1;
	wire w_dff_B_aOgU4ELB6_1;
	wire w_dff_B_jBp8iQ3Q9_1;
	wire w_dff_B_g0i2eiEM2_1;
	wire w_dff_B_naq7KaiY9_1;
	wire w_dff_B_m4BD1M7t1_1;
	wire w_dff_B_qFC3XSkr0_1;
	wire w_dff_B_2H7MoZBm6_1;
	wire w_dff_B_4ffmlxfy8_1;
	wire w_dff_B_qkn14MKe0_1;
	wire w_dff_B_GV0mab0N4_1;
	wire w_dff_B_fzBtasrw2_1;
	wire w_dff_B_5dTKk3Gk5_1;
	wire w_dff_B_5rHczfM12_1;
	wire w_dff_B_BARQITdw4_1;
	wire w_dff_B_S6Xp7R9T7_1;
	wire w_dff_B_CJy5Xudd4_1;
	wire w_dff_B_UYfj7fOI1_1;
	wire w_dff_B_yS4atw2d4_1;
	wire w_dff_B_NswG0Ans4_1;
	wire w_dff_B_un6YYT3w5_1;
	wire w_dff_B_cd3W0sKe7_1;
	wire w_dff_B_PxnsfXQZ8_1;
	wire w_dff_B_s8ZLoxsW1_1;
	wire w_dff_B_68u018ga6_1;
	wire w_dff_B_FqSwABMJ7_1;
	wire w_dff_B_DQBQpGpU6_1;
	wire w_dff_B_c6elk3rw8_1;
	wire w_dff_B_2LS1FMrT4_1;
	wire w_dff_B_J0Fw0MuX7_1;
	wire w_dff_B_TjlvXwnq4_1;
	wire w_dff_B_svhjiGLW0_1;
	wire w_dff_B_y1tLFf3b4_1;
	wire w_dff_B_dXwZTh0u6_1;
	wire w_dff_B_2MiLxxwT9_1;
	wire w_dff_B_5h9EYBja3_1;
	wire w_dff_B_uuDfBczC4_1;
	wire w_dff_B_bodVyx9Q6_1;
	wire w_dff_B_0YEbGJsP3_1;
	wire w_dff_B_mKcGy4RO9_1;
	wire w_dff_B_Zofr1Qmk2_1;
	wire w_dff_B_UCeFjkBI3_1;
	wire w_dff_B_Bi5E5g4R2_1;
	wire w_dff_B_HWGdJFXr9_1;
	wire w_dff_B_Y3aalqrp4_1;
	wire w_dff_B_694Nfgxd3_1;
	wire w_dff_B_5nkSaVSg7_1;
	wire w_dff_B_3ae3CVYA4_1;
	wire w_dff_B_qwKXXEMs6_1;
	wire w_dff_B_vwIKYOXo0_1;
	wire w_dff_B_EkvemZGx2_1;
	wire w_dff_B_GWiituuR1_1;
	wire w_dff_B_cAicZc2D5_1;
	wire w_dff_B_EJZE4J9r1_1;
	wire w_dff_B_h1oZradx8_1;
	wire w_dff_B_1yxZmgRd1_1;
	wire w_dff_B_uDLlYtDu1_1;
	wire w_dff_B_leKrtHrF3_1;
	wire w_dff_B_oAT0uDd04_1;
	wire w_dff_B_LBcou8w18_1;
	wire w_dff_B_edF1hDSZ5_1;
	wire w_dff_B_trYikcLE6_1;
	wire w_dff_B_2ijSUluq4_1;
	wire w_dff_B_cK3bqB2z0_1;
	wire w_dff_B_X3eQIbMu3_1;
	wire w_dff_B_1wTGGqE21_1;
	wire w_dff_B_RChdCOTh8_1;
	wire w_dff_B_wh6kJdJV9_1;
	wire w_dff_B_YNnywHuL3_1;
	wire w_dff_B_V2jjIySG7_1;
	wire w_dff_B_JXQfFvYb1_1;
	wire w_dff_B_ktrX3pFw7_1;
	wire w_dff_B_g5pGDcfh4_1;
	wire w_dff_B_ls9plk3d3_1;
	wire w_dff_B_Wtb0mdY08_1;
	wire w_dff_B_TtFRaT1f7_1;
	wire w_dff_B_bcnFMOvs1_1;
	wire w_dff_B_kx5kWE2b9_1;
	wire w_dff_B_VQf37a1h2_1;
	wire w_dff_B_XYc0K6132_1;
	wire w_dff_B_EzaJodqS8_0;
	wire w_dff_B_zP9IFLva5_0;
	wire w_dff_B_Tbfqh9zA3_0;
	wire w_dff_B_Cwt730ap3_0;
	wire w_dff_B_cy1KuHkc1_0;
	wire w_dff_B_CSikebnx7_0;
	wire w_dff_B_t9C8YF5G1_0;
	wire w_dff_B_s8yVXaTS5_0;
	wire w_dff_B_aJeEXzM93_0;
	wire w_dff_B_QdFdyFSq2_0;
	wire w_dff_B_jdvTHacl8_0;
	wire w_dff_B_wDvCAyRX8_0;
	wire w_dff_B_RMSbwqqE2_0;
	wire w_dff_B_xDL61mur8_0;
	wire w_dff_B_ZO8MFldP8_0;
	wire w_dff_B_X0KhYbQ66_0;
	wire w_dff_B_dVn7ltZl7_0;
	wire w_dff_B_vxWHWu4e2_0;
	wire w_dff_B_W9yqDw8o0_0;
	wire w_dff_B_CjTMqDBl6_0;
	wire w_dff_B_hInJTAAg2_0;
	wire w_dff_B_HXswUPXO0_0;
	wire w_dff_B_1Rl8B2Dz8_0;
	wire w_dff_B_v0oqxoB94_0;
	wire w_dff_B_MIFTPmTL7_0;
	wire w_dff_B_bBDwxaEU5_0;
	wire w_dff_B_WXLUjImo9_0;
	wire w_dff_B_NK50IKiS3_0;
	wire w_dff_B_2YiMrnQS0_0;
	wire w_dff_B_tVBaLwx42_0;
	wire w_dff_B_fLtHDs0x3_0;
	wire w_dff_B_Xjiu6Mnu7_0;
	wire w_dff_B_XFhThrOF0_0;
	wire w_dff_B_FA6HpplW5_0;
	wire w_dff_B_ojhXwi681_0;
	wire w_dff_B_9NYK3v9Z0_0;
	wire w_dff_B_MCt5C8fh3_0;
	wire w_dff_B_bCCKn63x3_0;
	wire w_dff_B_q0ybYMd12_0;
	wire w_dff_B_euud8xNN7_0;
	wire w_dff_B_Y2Vo3erM5_0;
	wire w_dff_B_qhJxRSJ44_0;
	wire w_dff_B_EBNT5MeV9_0;
	wire w_dff_B_YnX8SGd08_0;
	wire w_dff_B_2kQGa55j6_0;
	wire w_dff_B_obwXsIGL8_0;
	wire w_dff_B_gdTSAvy01_0;
	wire w_dff_B_mHLn9DCy3_0;
	wire w_dff_B_A1Djr5mL5_0;
	wire w_dff_B_Vp1hRAYR3_0;
	wire w_dff_B_YtUm7cWw3_0;
	wire w_dff_B_snbSRhzY7_0;
	wire w_dff_B_7mOYbSHb8_0;
	wire w_dff_B_RxgRsp3S6_0;
	wire w_dff_B_TTEbFWa84_0;
	wire w_dff_B_pJYDz0MA3_0;
	wire w_dff_B_W5BfMJYa0_0;
	wire w_dff_B_Zd3kwPHU1_0;
	wire w_dff_B_SFBUncDH0_0;
	wire w_dff_B_Dp1BL3Ip1_0;
	wire w_dff_B_KlGlmZea4_0;
	wire w_dff_B_8bIsnR6f2_0;
	wire w_dff_B_VwcpeNwQ2_0;
	wire w_dff_B_zjprAQc92_0;
	wire w_dff_B_zlkwCEOt7_0;
	wire w_dff_B_jGVr0YIp3_0;
	wire w_dff_B_IlVMj93h0_0;
	wire w_dff_B_rWdFK9hF0_0;
	wire w_dff_B_ViOOoSv25_0;
	wire w_dff_B_8nK4QXOd6_0;
	wire w_dff_B_gxbzngQU7_0;
	wire w_dff_B_NSLytmao5_0;
	wire w_dff_B_7hn2KMY03_0;
	wire w_dff_B_avi2Sthf6_0;
	wire w_dff_B_Z6X1g8iq5_0;
	wire w_dff_B_i4Og4My66_0;
	wire w_dff_B_mdAtJWfp1_0;
	wire w_dff_B_v8vyGl5N8_0;
	wire w_dff_B_0QReq4ua6_0;
	wire w_dff_B_W21oVGa69_0;
	wire w_dff_B_AI11iYyS8_0;
	wire w_dff_B_1cVDvt215_0;
	wire w_dff_B_5L1xQX1p4_0;
	wire w_dff_B_TlSqn3Pj0_0;
	wire w_dff_B_swBtowFI2_0;
	wire w_dff_B_T8dJDN1p1_0;
	wire w_dff_B_8Z3eKigZ2_0;
	wire w_dff_B_fihr9Zdv1_0;
	wire w_dff_B_rSXCiBYb8_0;
	wire w_dff_B_Cb0KbrkC5_0;
	wire w_dff_B_c9NF1VNd0_0;
	wire w_dff_B_hg4UEku54_0;
	wire w_dff_B_ZAsXg52V5_0;
	wire w_dff_B_L3vW8Ise2_0;
	wire w_dff_B_ODlMj3Lr1_0;
	wire w_dff_B_LYbrjwl59_0;
	wire w_dff_B_Eipc1ETl2_0;
	wire w_dff_B_Xt1ZESqP2_0;
	wire w_dff_B_NKXseSeN5_0;
	wire w_dff_B_05y7fX6B6_0;
	wire w_dff_B_aRt1Bn6g6_0;
	wire w_dff_B_opvjvs1u1_0;
	wire w_dff_B_kAHZOL9x7_0;
	wire w_dff_B_sAfaT4qB9_0;
	wire w_dff_B_INXXsf2p8_0;
	wire w_dff_B_mv8K2Y7q9_0;
	wire w_dff_B_F9qpmOda1_0;
	wire w_dff_B_yF8jyCHj7_0;
	wire w_dff_B_cCpjDktR2_0;
	wire w_dff_B_SjSOfdQk3_0;
	wire w_dff_B_RljpaGqd9_0;
	wire w_dff_B_9stgRsss9_0;
	wire w_dff_B_mK9qdiWp4_0;
	wire w_dff_B_6gTBK1EM9_1;
	wire w_dff_B_uO3UTTnK8_1;
	wire w_dff_B_5EwD6ijE8_1;
	wire w_dff_B_SS19RUqy0_1;
	wire w_dff_B_3Auiu3ZY0_1;
	wire w_dff_B_PyWlXHIR0_1;
	wire w_dff_B_8YIlveUk2_1;
	wire w_dff_B_1irRMUgK8_1;
	wire w_dff_B_KABtyeGH4_1;
	wire w_dff_B_OuEdJBBJ2_1;
	wire w_dff_B_s25cA4pm4_1;
	wire w_dff_B_On2QhlCc3_1;
	wire w_dff_B_WgDPmVKq6_1;
	wire w_dff_B_oespMl3E3_1;
	wire w_dff_B_JtFFY2kH1_1;
	wire w_dff_B_Ywq9y5Pz7_1;
	wire w_dff_B_ShCw1KZ54_1;
	wire w_dff_B_I1gBqC4w6_1;
	wire w_dff_B_M9LTqsTF1_1;
	wire w_dff_B_rTrhKZFH4_1;
	wire w_dff_B_3C1foqNi2_1;
	wire w_dff_B_6gFS1gOo3_1;
	wire w_dff_B_shiMa7fG2_1;
	wire w_dff_B_rVLoYAcl3_1;
	wire w_dff_B_no7Scwuv7_1;
	wire w_dff_B_EiUnT0Xk6_1;
	wire w_dff_B_gMfcn3ey0_1;
	wire w_dff_B_ZJad3ImK8_1;
	wire w_dff_B_Zx9Qqb762_1;
	wire w_dff_B_aFJm5bRw2_1;
	wire w_dff_B_OPZyebUE7_1;
	wire w_dff_B_1dzxiVp58_1;
	wire w_dff_B_xz3eF4Kt5_1;
	wire w_dff_B_1ISlxlMM6_1;
	wire w_dff_B_fUyMmErb8_1;
	wire w_dff_B_IqkULnpB5_1;
	wire w_dff_B_UvgY0M8H1_1;
	wire w_dff_B_21IILwOy6_1;
	wire w_dff_B_JpGOYLhV7_1;
	wire w_dff_B_kNQKgbCZ1_1;
	wire w_dff_B_x22SxgCY9_1;
	wire w_dff_B_qnhqOrjf0_1;
	wire w_dff_B_nW3xrQnc4_1;
	wire w_dff_B_yil0NI7m4_1;
	wire w_dff_B_ViHlSzoC8_1;
	wire w_dff_B_SHNQ3Gih2_1;
	wire w_dff_B_WBZVi2Sp6_1;
	wire w_dff_B_fhZXCH4n9_1;
	wire w_dff_B_OxdEpg1X7_1;
	wire w_dff_B_rTh80AY43_1;
	wire w_dff_B_KCrW0SRh0_1;
	wire w_dff_B_4SdYkNW89_1;
	wire w_dff_B_rQo4x9RC5_1;
	wire w_dff_B_4Y1khT4L6_1;
	wire w_dff_B_uvutIR678_1;
	wire w_dff_B_igaI8JiZ5_1;
	wire w_dff_B_SOzl5xTF5_1;
	wire w_dff_B_IxxP0Bnh6_1;
	wire w_dff_B_kXPR3RWX8_1;
	wire w_dff_B_pF9ZeJ1X1_1;
	wire w_dff_B_Q7o9wOw31_1;
	wire w_dff_B_zUheRpOz1_1;
	wire w_dff_B_tlrv0vL40_1;
	wire w_dff_B_3vKfztKj3_1;
	wire w_dff_B_lNyLmvjt8_1;
	wire w_dff_B_EFXnHh7B1_1;
	wire w_dff_B_hJto8FeZ3_1;
	wire w_dff_B_YJbujVQj7_1;
	wire w_dff_B_wcygeEKr6_1;
	wire w_dff_B_EmmdnPCY9_1;
	wire w_dff_B_5W2tTDgZ9_1;
	wire w_dff_B_iAO25kjD1_1;
	wire w_dff_B_mK9JxwEz8_1;
	wire w_dff_B_bLpnqNvP2_1;
	wire w_dff_B_yDw2jqZu1_1;
	wire w_dff_B_zNwX4zva2_1;
	wire w_dff_B_jd7v22GO3_1;
	wire w_dff_B_GAORwh6C2_1;
	wire w_dff_B_EFQ4ScXG5_1;
	wire w_dff_B_b6GgD02e2_1;
	wire w_dff_B_MManmxoV8_1;
	wire w_dff_B_iqZtTlaH8_1;
	wire w_dff_B_8WEQ1V9L1_1;
	wire w_dff_B_srh5O0R77_1;
	wire w_dff_B_iMUG4Dhp3_1;
	wire w_dff_B_8u58h2Jp6_1;
	wire w_dff_B_KPr0hUaE8_1;
	wire w_dff_B_nbLOdoHx7_1;
	wire w_dff_B_vyLBmnSz8_1;
	wire w_dff_B_BKCZKVgF8_1;
	wire w_dff_B_K6ApCmot7_1;
	wire w_dff_B_CIxcN1lw0_1;
	wire w_dff_B_XCbllKuC4_1;
	wire w_dff_B_iMNuduJf2_1;
	wire w_dff_B_h9sZE2aB1_1;
	wire w_dff_B_u3sIVnAp9_1;
	wire w_dff_B_0GqivLDO1_1;
	wire w_dff_B_JSLl1Kq75_1;
	wire w_dff_B_Po7J7QsB6_1;
	wire w_dff_B_JLVVm7ep3_1;
	wire w_dff_B_AsiLObze4_1;
	wire w_dff_B_SIE3tkeY9_1;
	wire w_dff_B_1PvzNOCJ8_1;
	wire w_dff_B_JAPcQGai3_1;
	wire w_dff_B_r2QWZnGR7_1;
	wire w_dff_B_5GQWkxxL9_1;
	wire w_dff_B_Q1JYRqwz0_1;
	wire w_dff_B_Yc7NSR7p0_1;
	wire w_dff_B_hK4Xk5986_1;
	wire w_dff_B_mcQ4cN8r2_1;
	wire w_dff_B_cCB9zJ452_1;
	wire w_dff_B_3fsHmRIV7_1;
	wire w_dff_B_lXcbVTn96_0;
	wire w_dff_B_EuJsqeSg3_0;
	wire w_dff_B_MJDckVra5_0;
	wire w_dff_B_fisQWwGe5_0;
	wire w_dff_B_BQ24fjm62_0;
	wire w_dff_B_lu8MqvrR3_0;
	wire w_dff_B_jB1zSSsy8_0;
	wire w_dff_B_UjEPFYd52_0;
	wire w_dff_B_HOV4m2ek6_0;
	wire w_dff_B_6CVtGBpH5_0;
	wire w_dff_B_4aEeEHUi2_0;
	wire w_dff_B_JU99LIya2_0;
	wire w_dff_B_zrv6oWNC5_0;
	wire w_dff_B_6Gb5miR04_0;
	wire w_dff_B_5847u9wZ4_0;
	wire w_dff_B_1unM9Mx92_0;
	wire w_dff_B_iOepQaZo4_0;
	wire w_dff_B_rEz9W7s84_0;
	wire w_dff_B_uN2cxeDa8_0;
	wire w_dff_B_sctwvjzm9_0;
	wire w_dff_B_adZ2zJHA6_0;
	wire w_dff_B_OqUCJmYU8_0;
	wire w_dff_B_BX3hv6YD1_0;
	wire w_dff_B_m449Yf9y4_0;
	wire w_dff_B_8EmH85VL8_0;
	wire w_dff_B_3uZFVLjP4_0;
	wire w_dff_B_k3wenEl10_0;
	wire w_dff_B_v0QZ1dRM0_0;
	wire w_dff_B_U6EboWYB7_0;
	wire w_dff_B_XJ4iQiS00_0;
	wire w_dff_B_TkPSQJkp3_0;
	wire w_dff_B_jtbekEci6_0;
	wire w_dff_B_i71EgrhA0_0;
	wire w_dff_B_C9pjuqWt5_0;
	wire w_dff_B_dbes4qhe8_0;
	wire w_dff_B_aMUB5w0v3_0;
	wire w_dff_B_oWn261va5_0;
	wire w_dff_B_sgTcgaU81_0;
	wire w_dff_B_77tqyWvs1_0;
	wire w_dff_B_6APz98kU2_0;
	wire w_dff_B_TNhIk7Ih1_0;
	wire w_dff_B_cU0C33If0_0;
	wire w_dff_B_yJYmNmdh6_0;
	wire w_dff_B_iBtXgot99_0;
	wire w_dff_B_u5Mo357n1_0;
	wire w_dff_B_4DzhqyBu8_0;
	wire w_dff_B_WVUnn1F30_0;
	wire w_dff_B_lprqYsYz7_0;
	wire w_dff_B_hl4FJUbS7_0;
	wire w_dff_B_9A3Ssd8G5_0;
	wire w_dff_B_G9RerJcH4_0;
	wire w_dff_B_pLT6T9RD8_0;
	wire w_dff_B_PYAqlhWT4_0;
	wire w_dff_B_QemTcCs89_0;
	wire w_dff_B_3rWWJz0e4_0;
	wire w_dff_B_sVnjoQA17_0;
	wire w_dff_B_Ofwh46kp5_0;
	wire w_dff_B_hXscZl9E6_0;
	wire w_dff_B_jWCIsWrH5_0;
	wire w_dff_B_YoOEgNyD2_0;
	wire w_dff_B_56Jk0nau2_0;
	wire w_dff_B_i0LZErHj4_0;
	wire w_dff_B_PFUkBZh20_0;
	wire w_dff_B_WEzCsKLz3_0;
	wire w_dff_B_QvVvh4vt2_0;
	wire w_dff_B_dRo1ao7J4_0;
	wire w_dff_B_3x7bGVQX6_0;
	wire w_dff_B_GN6mD94b7_0;
	wire w_dff_B_JrVCeRGC2_0;
	wire w_dff_B_s3qJXBc55_0;
	wire w_dff_B_jjGFx3J51_0;
	wire w_dff_B_D5UzCQQy8_0;
	wire w_dff_B_tCqMjmsc2_0;
	wire w_dff_B_WKO7QTfx5_0;
	wire w_dff_B_p2rxYZOF2_0;
	wire w_dff_B_dHDv6ACA9_0;
	wire w_dff_B_rXzd1AYa1_0;
	wire w_dff_B_OkYKvnMa5_0;
	wire w_dff_B_6dTMppZA8_0;
	wire w_dff_B_AOGUaZLi2_0;
	wire w_dff_B_ApRG4ieU7_0;
	wire w_dff_B_Phgmjnkl1_0;
	wire w_dff_B_OL8cJkMh9_0;
	wire w_dff_B_z2bLtqbT5_0;
	wire w_dff_B_ALr5Fe5X0_0;
	wire w_dff_B_ClUh65WD4_0;
	wire w_dff_B_M2iqKTpG7_0;
	wire w_dff_B_UpJ9WE8l1_0;
	wire w_dff_B_lnFB99Bj8_0;
	wire w_dff_B_VAiZdZvZ6_0;
	wire w_dff_B_KgQSo1s25_0;
	wire w_dff_B_kJ8if1Rz8_0;
	wire w_dff_B_aevcQyYO9_0;
	wire w_dff_B_HkGrW22G5_0;
	wire w_dff_B_cPtHhfw96_0;
	wire w_dff_B_xMjn9can3_0;
	wire w_dff_B_qT5hyHnX6_0;
	wire w_dff_B_1ivdly6U4_0;
	wire w_dff_B_MlZiuXDQ4_0;
	wire w_dff_B_waMMDDVc1_0;
	wire w_dff_B_2CHPNr9c3_0;
	wire w_dff_B_KuGm4Giw7_0;
	wire w_dff_B_7eOg1sdf3_0;
	wire w_dff_B_1e0svXtD7_0;
	wire w_dff_B_zqxBeI1X0_0;
	wire w_dff_B_fcgveMbB5_0;
	wire w_dff_B_vHQ6kjWz2_0;
	wire w_dff_B_phBEkl3m2_0;
	wire w_dff_B_8wUH5XTf9_0;
	wire w_dff_B_aUAVFcQw1_0;
	wire w_dff_B_ncmA4MoC6_0;
	wire w_dff_B_9kk8s8Kj0_0;
	wire w_dff_B_f5fJqnrM7_1;
	wire w_dff_B_SCRBDtFc7_1;
	wire w_dff_B_kFZcFra90_1;
	wire w_dff_B_z9Ief7Ks5_1;
	wire w_dff_B_3ahmI1Xs7_1;
	wire w_dff_B_5AiS494R3_1;
	wire w_dff_B_3WgcX6Ds9_1;
	wire w_dff_B_0NYHveAO2_1;
	wire w_dff_B_MNNzQLw34_1;
	wire w_dff_B_wuIGaYfu8_1;
	wire w_dff_B_ZP15QZ0T1_1;
	wire w_dff_B_WTNqxCAK8_1;
	wire w_dff_B_x243EKgh1_1;
	wire w_dff_B_HbOt34VG0_1;
	wire w_dff_B_Yn3RuMFN6_1;
	wire w_dff_B_87KBbj4Y4_1;
	wire w_dff_B_4GRhYBde0_1;
	wire w_dff_B_iw1OlsIB4_1;
	wire w_dff_B_p8x0bEBn2_1;
	wire w_dff_B_O8akJU065_1;
	wire w_dff_B_xIEFSa847_1;
	wire w_dff_B_pXrq6MKO9_1;
	wire w_dff_B_xzS58Tau8_1;
	wire w_dff_B_BCZ9PQjd4_1;
	wire w_dff_B_booaxSNR1_1;
	wire w_dff_B_D1ghgW416_1;
	wire w_dff_B_I0RR89VS4_1;
	wire w_dff_B_Syn8FOEL2_1;
	wire w_dff_B_tQKZaWqY5_1;
	wire w_dff_B_KRNn8g490_1;
	wire w_dff_B_n4Cih7Cs0_1;
	wire w_dff_B_V8is0NG60_1;
	wire w_dff_B_uCXvTn7W7_1;
	wire w_dff_B_DfgfrNC04_1;
	wire w_dff_B_PoDMF17E9_1;
	wire w_dff_B_GvWs4D6b5_1;
	wire w_dff_B_jt6GZ1SQ9_1;
	wire w_dff_B_VEjB5MWe7_1;
	wire w_dff_B_JNWa2Hc12_1;
	wire w_dff_B_YedQTxBc1_1;
	wire w_dff_B_MWVEk7Yy2_1;
	wire w_dff_B_SGVrIX835_1;
	wire w_dff_B_iViIFdnS5_1;
	wire w_dff_B_s0cNhQew7_1;
	wire w_dff_B_c9Bs7ZZT3_1;
	wire w_dff_B_wbRhDBm88_1;
	wire w_dff_B_9iNe9YHu5_1;
	wire w_dff_B_AjXH0r3u6_1;
	wire w_dff_B_thVnRWrT7_1;
	wire w_dff_B_0PTJ0m2x9_1;
	wire w_dff_B_x67HYtzZ6_1;
	wire w_dff_B_Wyg9oLko4_1;
	wire w_dff_B_m7XQnY6f9_1;
	wire w_dff_B_86GG1ANT4_1;
	wire w_dff_B_fn7ngN5V4_1;
	wire w_dff_B_0NQxYXRW8_1;
	wire w_dff_B_dJdFIWHo0_1;
	wire w_dff_B_z9XltW5J7_1;
	wire w_dff_B_3mqeqZlv1_1;
	wire w_dff_B_0ZoUOAI12_1;
	wire w_dff_B_VsP0cSah0_1;
	wire w_dff_B_JcEcZDWL8_1;
	wire w_dff_B_krdChQNe4_1;
	wire w_dff_B_MZqqAY5K4_1;
	wire w_dff_B_iOZ3gROo8_1;
	wire w_dff_B_92w27m5X0_1;
	wire w_dff_B_ZglMHgYd9_1;
	wire w_dff_B_PbFPI6Fe5_1;
	wire w_dff_B_jchvVAJs1_1;
	wire w_dff_B_1DlG3P9Z6_1;
	wire w_dff_B_dNz23Tyv9_1;
	wire w_dff_B_E7DbAjSu7_1;
	wire w_dff_B_eHpZEKlY6_1;
	wire w_dff_B_Qj8FgEmd8_1;
	wire w_dff_B_XnaP1RXz3_1;
	wire w_dff_B_Jucbebss1_1;
	wire w_dff_B_EYBMdIFj3_1;
	wire w_dff_B_gwICwd4J7_1;
	wire w_dff_B_hEZ8aKD22_1;
	wire w_dff_B_68lFFIXZ4_1;
	wire w_dff_B_w4VXy8Sb4_1;
	wire w_dff_B_ny3alXd71_1;
	wire w_dff_B_MSi1KQ8d1_1;
	wire w_dff_B_HIsATejX5_1;
	wire w_dff_B_EFcE9LzN3_1;
	wire w_dff_B_r09dneTc2_1;
	wire w_dff_B_oOjE5vBU7_1;
	wire w_dff_B_SVsaNuYL0_1;
	wire w_dff_B_QUH1PpSS8_1;
	wire w_dff_B_bMwO5Ksz5_1;
	wire w_dff_B_FatS89pc5_1;
	wire w_dff_B_GbeDqxmI8_1;
	wire w_dff_B_NOPoR7ZS0_1;
	wire w_dff_B_rgwx18Bc2_1;
	wire w_dff_B_mEZrt6z78_1;
	wire w_dff_B_PgCb1xBM1_1;
	wire w_dff_B_gGE28DBO2_1;
	wire w_dff_B_9xckHE418_1;
	wire w_dff_B_LHB3u8c70_1;
	wire w_dff_B_DZ6NZwNS8_1;
	wire w_dff_B_PMS6C3Ib7_1;
	wire w_dff_B_Y81h77nn0_1;
	wire w_dff_B_YKDPraiS0_1;
	wire w_dff_B_dI7R08Xx1_1;
	wire w_dff_B_TNs070wt2_1;
	wire w_dff_B_9kifPkEd3_1;
	wire w_dff_B_Ss2Uaxdz6_1;
	wire w_dff_B_vm75blfX0_1;
	wire w_dff_B_2X6D9LyI9_1;
	wire w_dff_B_3ncbrnNb2_1;
	wire w_dff_B_7nEsIUQP7_1;
	wire w_dff_B_vh99L45W1_0;
	wire w_dff_B_WpPMkpzG4_0;
	wire w_dff_B_Q6ZTjjX75_0;
	wire w_dff_B_xKamv6vY8_0;
	wire w_dff_B_VCua7QkI4_0;
	wire w_dff_B_oxsb2J787_0;
	wire w_dff_B_9u38LOqB5_0;
	wire w_dff_B_loVxnU1V7_0;
	wire w_dff_B_scLkIwhk8_0;
	wire w_dff_B_18gcbKV37_0;
	wire w_dff_B_jBeGjqSL4_0;
	wire w_dff_B_LucZaYKp2_0;
	wire w_dff_B_f1DNbYTn6_0;
	wire w_dff_B_DjVneDZu7_0;
	wire w_dff_B_HRpiISse9_0;
	wire w_dff_B_DsmGcOrD9_0;
	wire w_dff_B_gnlDjTcb3_0;
	wire w_dff_B_Ns3pgPzD7_0;
	wire w_dff_B_oMCrHf1M1_0;
	wire w_dff_B_WaEEoS817_0;
	wire w_dff_B_JJ8F5yyf2_0;
	wire w_dff_B_8pAQ3Lj87_0;
	wire w_dff_B_atqK1YFV5_0;
	wire w_dff_B_jzaHvS473_0;
	wire w_dff_B_Mr5QEqgj0_0;
	wire w_dff_B_fR3Luis86_0;
	wire w_dff_B_XbWQcGBV3_0;
	wire w_dff_B_hfM7cqph0_0;
	wire w_dff_B_303QQDhd6_0;
	wire w_dff_B_RCfuaQTD0_0;
	wire w_dff_B_Kt9M91KE3_0;
	wire w_dff_B_KbOef6La6_0;
	wire w_dff_B_hLPLZt4l5_0;
	wire w_dff_B_AhxYsQDU0_0;
	wire w_dff_B_Gg644Uby4_0;
	wire w_dff_B_3Bnn5R344_0;
	wire w_dff_B_CqDmdEoC8_0;
	wire w_dff_B_QFhFRcxg6_0;
	wire w_dff_B_AC1xFoOV4_0;
	wire w_dff_B_o8P8HGCg4_0;
	wire w_dff_B_tCCy3xBw1_0;
	wire w_dff_B_2uK9qrsP1_0;
	wire w_dff_B_Zu7Qzsol6_0;
	wire w_dff_B_LuA8ccpT0_0;
	wire w_dff_B_LXIS0KMU6_0;
	wire w_dff_B_nudrdhfk0_0;
	wire w_dff_B_qaIlPDop6_0;
	wire w_dff_B_hzPq7EEo2_0;
	wire w_dff_B_61XcsiEZ2_0;
	wire w_dff_B_hWMclC1a1_0;
	wire w_dff_B_dPHn03oe7_0;
	wire w_dff_B_aTFnL8Uf6_0;
	wire w_dff_B_l0d8bZ0v1_0;
	wire w_dff_B_HufA5ZQ70_0;
	wire w_dff_B_KVVOJQLQ0_0;
	wire w_dff_B_bgNzMwST0_0;
	wire w_dff_B_SlPhwksZ4_0;
	wire w_dff_B_tQrdhgjC0_0;
	wire w_dff_B_kynfNtjN7_0;
	wire w_dff_B_Y2yw4CJS2_0;
	wire w_dff_B_DlBbqP5E9_0;
	wire w_dff_B_Twf2Fwju5_0;
	wire w_dff_B_aQaGiu9v3_0;
	wire w_dff_B_LyVO3kP23_0;
	wire w_dff_B_3fAnSOOd2_0;
	wire w_dff_B_i9OJ2SyL0_0;
	wire w_dff_B_eMBNXdNB4_0;
	wire w_dff_B_HtrNzdA12_0;
	wire w_dff_B_8k0y6odc7_0;
	wire w_dff_B_zzKyXlL40_0;
	wire w_dff_B_FqdQTw0W7_0;
	wire w_dff_B_WpwrAOeV6_0;
	wire w_dff_B_51kRVBih6_0;
	wire w_dff_B_cVlwItkV7_0;
	wire w_dff_B_p7WDw7xv5_0;
	wire w_dff_B_Zjihcsk99_0;
	wire w_dff_B_6C0fUjTS9_0;
	wire w_dff_B_PZt9ZuhX2_0;
	wire w_dff_B_l9IeCJRH7_0;
	wire w_dff_B_LO9LHHVb9_0;
	wire w_dff_B_LDV9GZol4_0;
	wire w_dff_B_5NpUfDCB0_0;
	wire w_dff_B_VmNsO4Go8_0;
	wire w_dff_B_MYjzijZW4_0;
	wire w_dff_B_SMQciwVq1_0;
	wire w_dff_B_ix9eixGn3_0;
	wire w_dff_B_JY5qLTsg5_0;
	wire w_dff_B_kGbyK0P85_0;
	wire w_dff_B_VSIalSkS8_0;
	wire w_dff_B_zzr6kFSZ2_0;
	wire w_dff_B_iwC1qx737_0;
	wire w_dff_B_LGOGR9YC7_0;
	wire w_dff_B_YpLf8Nod4_0;
	wire w_dff_B_au9UPdnR0_0;
	wire w_dff_B_g94g8swf6_0;
	wire w_dff_B_D1UWS14P5_0;
	wire w_dff_B_XmXDk5Sm5_0;
	wire w_dff_B_oXxfIAPA4_0;
	wire w_dff_B_zEaB8Ke58_0;
	wire w_dff_B_oDifmN1a4_0;
	wire w_dff_B_DvpOnxyT4_0;
	wire w_dff_B_2Q35UFnP7_0;
	wire w_dff_B_MODqHYDS0_0;
	wire w_dff_B_aGYC2kHH9_0;
	wire w_dff_B_eNX3bVES5_0;
	wire w_dff_B_t3PLhM7D0_0;
	wire w_dff_B_6luBvCat5_0;
	wire w_dff_B_iK4jWOFR2_0;
	wire w_dff_B_uw84qvIf3_0;
	wire w_dff_B_vOcnNdYY1_0;
	wire w_dff_B_JR5SiCzG0_0;
	wire w_dff_B_TNJgKzWo1_1;
	wire w_dff_B_lBCSnp2r7_1;
	wire w_dff_B_AVtLB6jr6_1;
	wire w_dff_B_24zzqBRI7_1;
	wire w_dff_B_x00mff6S6_1;
	wire w_dff_B_CDoGWpv02_1;
	wire w_dff_B_VGwfrrk02_1;
	wire w_dff_B_R7azb7Nd0_1;
	wire w_dff_B_v3RRxXsr0_1;
	wire w_dff_B_sFTrb7JH8_1;
	wire w_dff_B_JXW2zXQv5_1;
	wire w_dff_B_qLZvhUXn6_1;
	wire w_dff_B_Zs7x17fS0_1;
	wire w_dff_B_htye1RPi7_1;
	wire w_dff_B_uveo5U1G9_1;
	wire w_dff_B_FC3OSfkT6_1;
	wire w_dff_B_URjIChGw1_1;
	wire w_dff_B_cilZ3TtY0_1;
	wire w_dff_B_P8JUk6yn2_1;
	wire w_dff_B_sY810B3m1_1;
	wire w_dff_B_yfXeADdj6_1;
	wire w_dff_B_AUyAgJEw7_1;
	wire w_dff_B_oYwKGmbN0_1;
	wire w_dff_B_WNN78y1p2_1;
	wire w_dff_B_BmZiL57t3_1;
	wire w_dff_B_l01DRcmO0_1;
	wire w_dff_B_IIxIsKNe0_1;
	wire w_dff_B_0EvjvlxC6_1;
	wire w_dff_B_d0vS4m3V9_1;
	wire w_dff_B_ZUldIZr71_1;
	wire w_dff_B_cV71bmen7_1;
	wire w_dff_B_zWCE6COk1_1;
	wire w_dff_B_YgtXdsHb7_1;
	wire w_dff_B_iRSEWnqw4_1;
	wire w_dff_B_e1hi6Rn85_1;
	wire w_dff_B_3NjjINVj8_1;
	wire w_dff_B_RAtNW0Gg1_1;
	wire w_dff_B_AqJAn9bb1_1;
	wire w_dff_B_gZsuQJOZ9_1;
	wire w_dff_B_7qyUS5Wd2_1;
	wire w_dff_B_ACuUdNia4_1;
	wire w_dff_B_X5gl6zrp8_1;
	wire w_dff_B_9o42I44L6_1;
	wire w_dff_B_5mx11BE19_1;
	wire w_dff_B_iMrH0NZ31_1;
	wire w_dff_B_78QfnOWx4_1;
	wire w_dff_B_iJowQtKq0_1;
	wire w_dff_B_cf3m5jsR2_1;
	wire w_dff_B_uSgMIlFd1_1;
	wire w_dff_B_czIanC4b1_1;
	wire w_dff_B_0SsKP0wG1_1;
	wire w_dff_B_kMOcvVJd2_1;
	wire w_dff_B_AryzQLz15_1;
	wire w_dff_B_DQxIC9Z15_1;
	wire w_dff_B_bOKXOzTI4_1;
	wire w_dff_B_PJynUqyP3_1;
	wire w_dff_B_BXe3PbWw8_1;
	wire w_dff_B_gIFHpA6r4_1;
	wire w_dff_B_l9MmpgVJ6_1;
	wire w_dff_B_BSPTMW9T6_1;
	wire w_dff_B_z6XbKa2O2_1;
	wire w_dff_B_zMf20qIv4_1;
	wire w_dff_B_lESTFKZ39_1;
	wire w_dff_B_a72zZHwv7_1;
	wire w_dff_B_fvfuyOux9_1;
	wire w_dff_B_laBtyieW9_1;
	wire w_dff_B_tfNxG1O59_1;
	wire w_dff_B_xSu9ZqGL9_1;
	wire w_dff_B_byiIojBQ1_1;
	wire w_dff_B_TcMM18NK4_1;
	wire w_dff_B_iYUPolPE7_1;
	wire w_dff_B_gYVM8Glb9_1;
	wire w_dff_B_Sfr4aSJK3_1;
	wire w_dff_B_VCcD85Xm0_1;
	wire w_dff_B_dsvKWkqG3_1;
	wire w_dff_B_LKHs9SzN2_1;
	wire w_dff_B_EHMgFfpX0_1;
	wire w_dff_B_NN6hkRKp7_1;
	wire w_dff_B_8Z3PMryr0_1;
	wire w_dff_B_MWsgv9wk2_1;
	wire w_dff_B_6XyXBagH2_1;
	wire w_dff_B_9IMyFUuV7_1;
	wire w_dff_B_Ybge9p9p6_1;
	wire w_dff_B_BZ0kkJPv2_1;
	wire w_dff_B_3aSt7qKB5_1;
	wire w_dff_B_8D7NpUrs5_1;
	wire w_dff_B_1U6ocUSr9_1;
	wire w_dff_B_MZcbJ2FL9_1;
	wire w_dff_B_ZbzCUrij7_1;
	wire w_dff_B_Iy6YBLzm9_1;
	wire w_dff_B_zo0eN7VF1_1;
	wire w_dff_B_LetsnoQ83_1;
	wire w_dff_B_QMtwEum80_1;
	wire w_dff_B_XOHB2wXJ3_1;
	wire w_dff_B_M33UaZg95_1;
	wire w_dff_B_8nKa2SG72_1;
	wire w_dff_B_6ys3D0sJ8_1;
	wire w_dff_B_o0TBXR9R3_1;
	wire w_dff_B_p2oBQjh34_1;
	wire w_dff_B_9abC3eYk2_1;
	wire w_dff_B_DV8yiukN4_1;
	wire w_dff_B_vUmolh8w9_1;
	wire w_dff_B_7DHWEMMT2_1;
	wire w_dff_B_FMeYhrLy9_1;
	wire w_dff_B_V0ivtjd62_1;
	wire w_dff_B_H8tSLsLj6_1;
	wire w_dff_B_Vf5hwBZA4_1;
	wire w_dff_B_ZTG1a3co6_1;
	wire w_dff_B_3DnFUkNN0_1;
	wire w_dff_B_sX8cRBX78_1;
	wire w_dff_B_eijfc5pg6_0;
	wire w_dff_B_Kki71dkq6_0;
	wire w_dff_B_8tQuyefM2_0;
	wire w_dff_B_FaedtkvH6_0;
	wire w_dff_B_kpbLbBbY0_0;
	wire w_dff_B_wPp5KZpI7_0;
	wire w_dff_B_1bxbF8on2_0;
	wire w_dff_B_vSXwfNEF7_0;
	wire w_dff_B_eijOniyI3_0;
	wire w_dff_B_nV3SEymu4_0;
	wire w_dff_B_8kv3raGy9_0;
	wire w_dff_B_eV68pfbm2_0;
	wire w_dff_B_100189Eh1_0;
	wire w_dff_B_OX60F6sO5_0;
	wire w_dff_B_2ZhW6l159_0;
	wire w_dff_B_ZxPYZXRq7_0;
	wire w_dff_B_2hpBib9f8_0;
	wire w_dff_B_wh6eX9fk6_0;
	wire w_dff_B_rKbtq0A12_0;
	wire w_dff_B_uYH3qtOg1_0;
	wire w_dff_B_2yYLkmNq7_0;
	wire w_dff_B_31P7kpkf3_0;
	wire w_dff_B_KnAeTAsA9_0;
	wire w_dff_B_rrOkmwmw6_0;
	wire w_dff_B_1mOsWA3e8_0;
	wire w_dff_B_vNc2k22x5_0;
	wire w_dff_B_H9jodjJU9_0;
	wire w_dff_B_MuNVOHU85_0;
	wire w_dff_B_bS1gtJIQ2_0;
	wire w_dff_B_Fy5hxjQG2_0;
	wire w_dff_B_ESI79r7D6_0;
	wire w_dff_B_pN7FLYz65_0;
	wire w_dff_B_aRPsBVvL0_0;
	wire w_dff_B_x117IfYm2_0;
	wire w_dff_B_ayDpPYeB9_0;
	wire w_dff_B_8c211PYI1_0;
	wire w_dff_B_JurUsh7g3_0;
	wire w_dff_B_Ny1UPnCN7_0;
	wire w_dff_B_jb4Whx431_0;
	wire w_dff_B_JdekCFq97_0;
	wire w_dff_B_bCh4qLeT5_0;
	wire w_dff_B_larob4IN7_0;
	wire w_dff_B_59UCg4tp4_0;
	wire w_dff_B_zWSRUSon2_0;
	wire w_dff_B_VmeH1jGz6_0;
	wire w_dff_B_0U550N7F1_0;
	wire w_dff_B_ukIxxz0y6_0;
	wire w_dff_B_0t9lsczO6_0;
	wire w_dff_B_hrQNrluM5_0;
	wire w_dff_B_Uai1f90i2_0;
	wire w_dff_B_STa2ezN83_0;
	wire w_dff_B_Ldlh7Pm86_0;
	wire w_dff_B_ERu4tLOb4_0;
	wire w_dff_B_RiBaRBtP4_0;
	wire w_dff_B_GW4R7AIJ5_0;
	wire w_dff_B_uPnO5vJ01_0;
	wire w_dff_B_TzLWDAsc6_0;
	wire w_dff_B_3H9T2crH9_0;
	wire w_dff_B_IBPXt5Ow0_0;
	wire w_dff_B_4hqYCYAG7_0;
	wire w_dff_B_BH0Ge5NT6_0;
	wire w_dff_B_2daF8TP68_0;
	wire w_dff_B_o39NmiNr7_0;
	wire w_dff_B_sF22bwQT7_0;
	wire w_dff_B_Ph1O0jJO8_0;
	wire w_dff_B_mis7YoWy3_0;
	wire w_dff_B_SMG1l1Rg5_0;
	wire w_dff_B_BFBtnrUY2_0;
	wire w_dff_B_T2qhl3b43_0;
	wire w_dff_B_819bPhog1_0;
	wire w_dff_B_CyGo6Nfs8_0;
	wire w_dff_B_JIafjria0_0;
	wire w_dff_B_YHutGRmb3_0;
	wire w_dff_B_OInsV6VW0_0;
	wire w_dff_B_WjXlSdFp5_0;
	wire w_dff_B_hCeTkbMk3_0;
	wire w_dff_B_WNUB00xy9_0;
	wire w_dff_B_SZ4VXvos9_0;
	wire w_dff_B_yzzc5q2Q3_0;
	wire w_dff_B_pkRr9Hfb7_0;
	wire w_dff_B_O7jpM7Rg7_0;
	wire w_dff_B_vL7lzYGD0_0;
	wire w_dff_B_YkZUb3pQ5_0;
	wire w_dff_B_2qwDEWHw7_0;
	wire w_dff_B_7WIssvmJ4_0;
	wire w_dff_B_Mal5DAro1_0;
	wire w_dff_B_qycH0BtL6_0;
	wire w_dff_B_RKNvS5rk7_0;
	wire w_dff_B_dtoruauM9_0;
	wire w_dff_B_UqsaClGw3_0;
	wire w_dff_B_j79nUqGF6_0;
	wire w_dff_B_RMfEebmb3_0;
	wire w_dff_B_y1FZ4rqb3_0;
	wire w_dff_B_CVQQtmVk9_0;
	wire w_dff_B_l6CIO8uO6_0;
	wire w_dff_B_a8iR5bg72_0;
	wire w_dff_B_smNCzs7c0_0;
	wire w_dff_B_IBJgy6V73_0;
	wire w_dff_B_N68b2DFq4_0;
	wire w_dff_B_euMyhzMj6_0;
	wire w_dff_B_0jmMO6n58_0;
	wire w_dff_B_WF6q6UMt6_0;
	wire w_dff_B_L9nTN4eZ4_0;
	wire w_dff_B_IrRSRxVR0_0;
	wire w_dff_B_GpeT42fu3_0;
	wire w_dff_B_wmA091ne9_0;
	wire w_dff_B_fs04zcVl2_0;
	wire w_dff_B_3duPMmKT4_0;
	wire w_dff_B_0ST06S6Z7_0;
	wire w_dff_B_gYw3T9cY7_0;
	wire w_dff_B_GdXnogvr7_1;
	wire w_dff_B_XQwIbR8p4_1;
	wire w_dff_B_XRW2itrt9_1;
	wire w_dff_B_W5fOSvQ24_1;
	wire w_dff_B_cIPUVuF94_1;
	wire w_dff_B_7XdPC3LR4_1;
	wire w_dff_B_5T81fUaD8_1;
	wire w_dff_B_8bQZlJOO0_1;
	wire w_dff_B_XqgXzWwt8_1;
	wire w_dff_B_oftdZZa24_1;
	wire w_dff_B_tT9aN8G51_1;
	wire w_dff_B_40NbgsGD4_1;
	wire w_dff_B_rvr7EOT11_1;
	wire w_dff_B_aKGcBlSp4_1;
	wire w_dff_B_vcQiqavX5_1;
	wire w_dff_B_mDKkOzfl8_1;
	wire w_dff_B_qaB5zHrA2_1;
	wire w_dff_B_Jya1gP1o4_1;
	wire w_dff_B_OlbHQIYo5_1;
	wire w_dff_B_DvvFtIW32_1;
	wire w_dff_B_WGVbmZp47_1;
	wire w_dff_B_Fpv9YHTV0_1;
	wire w_dff_B_6d2eINSq6_1;
	wire w_dff_B_aKp1oa0J7_1;
	wire w_dff_B_0tMQlvNh4_1;
	wire w_dff_B_Ac7jinqw7_1;
	wire w_dff_B_VmsNyaTt1_1;
	wire w_dff_B_HGFYq3Nj1_1;
	wire w_dff_B_LUdSKeJ88_1;
	wire w_dff_B_7L2Keg130_1;
	wire w_dff_B_kLnz6kAV0_1;
	wire w_dff_B_yOOvbO6P0_1;
	wire w_dff_B_PbUxpgOp0_1;
	wire w_dff_B_VBS6iIeL7_1;
	wire w_dff_B_U0YrBBnK6_1;
	wire w_dff_B_nE5ZQDb68_1;
	wire w_dff_B_9gi2erYH8_1;
	wire w_dff_B_70vy9pFs4_1;
	wire w_dff_B_YLQZl8bD2_1;
	wire w_dff_B_DrxjVXPS8_1;
	wire w_dff_B_gicHjYTq4_1;
	wire w_dff_B_IC5KiwpU8_1;
	wire w_dff_B_LCAQhOok8_1;
	wire w_dff_B_Lcdse3FY4_1;
	wire w_dff_B_BEtKi7yH2_1;
	wire w_dff_B_20XgnWZD6_1;
	wire w_dff_B_7tWUc2sC8_1;
	wire w_dff_B_MbLVCZ504_1;
	wire w_dff_B_sj3oHv8P8_1;
	wire w_dff_B_1SWLi7Mg2_1;
	wire w_dff_B_BynzUjIH6_1;
	wire w_dff_B_lWhhEMYP5_1;
	wire w_dff_B_RebZUSRG0_1;
	wire w_dff_B_dEw66dmo6_1;
	wire w_dff_B_08QWJ17r5_1;
	wire w_dff_B_e10YDfn47_1;
	wire w_dff_B_WWg7wf7O1_1;
	wire w_dff_B_7u2dcfEg9_1;
	wire w_dff_B_5lpFBKTS5_1;
	wire w_dff_B_YdZFmXL88_1;
	wire w_dff_B_JfFWg1iW5_1;
	wire w_dff_B_Uk3Po1dr8_1;
	wire w_dff_B_8Mb32oqK2_1;
	wire w_dff_B_0Wk9LVZs3_1;
	wire w_dff_B_wuCGhu0J9_1;
	wire w_dff_B_QHXnIcX82_1;
	wire w_dff_B_z7rfscAq7_1;
	wire w_dff_B_Uq6s8GXI7_1;
	wire w_dff_B_gbo5BqUI5_1;
	wire w_dff_B_ecgcdOhE0_1;
	wire w_dff_B_ijMlERTJ4_1;
	wire w_dff_B_ipn2A3FN3_1;
	wire w_dff_B_Wb3hR7mj1_1;
	wire w_dff_B_LnGiy3TB1_1;
	wire w_dff_B_eLaz2e8v5_1;
	wire w_dff_B_WCavkgzK5_1;
	wire w_dff_B_PvztYaNT4_1;
	wire w_dff_B_0jZGnh2v2_1;
	wire w_dff_B_EGczUprh7_1;
	wire w_dff_B_6Lyd6ATI7_1;
	wire w_dff_B_MQg2O00O6_1;
	wire w_dff_B_vQT0tWoq5_1;
	wire w_dff_B_l3qwcyBC1_1;
	wire w_dff_B_CRG8t1ah8_1;
	wire w_dff_B_LNlJZs1C4_1;
	wire w_dff_B_IWux2oHZ9_1;
	wire w_dff_B_hxw07n0o8_1;
	wire w_dff_B_Jx6ohcKw2_1;
	wire w_dff_B_pldm7iwc9_1;
	wire w_dff_B_Ey1Bv6j82_1;
	wire w_dff_B_V78sD6Ie7_1;
	wire w_dff_B_rj64pd9j9_1;
	wire w_dff_B_amElfdG16_1;
	wire w_dff_B_lH6RBAX57_1;
	wire w_dff_B_cxCprxkp4_1;
	wire w_dff_B_eBYFtK4C2_1;
	wire w_dff_B_oq2MWXEb3_1;
	wire w_dff_B_ievQsVz30_1;
	wire w_dff_B_EMh02utm5_1;
	wire w_dff_B_1N4e48Hr0_1;
	wire w_dff_B_2rj0tbAx3_1;
	wire w_dff_B_3cLY4mMu9_1;
	wire w_dff_B_lPQkhTh67_1;
	wire w_dff_B_vzwRcvaQ5_1;
	wire w_dff_B_47jZaQhx6_1;
	wire w_dff_B_KQtw1Zjg3_1;
	wire w_dff_B_ji1m2Zy14_1;
	wire w_dff_B_Zeu5QyPt7_1;
	wire w_dff_B_mscM20U91_1;
	wire w_dff_B_OjgH8gAT8_0;
	wire w_dff_B_TQ78zH5j3_0;
	wire w_dff_B_K24HpLYV1_0;
	wire w_dff_B_R63ClVW62_0;
	wire w_dff_B_ELKXiSbI5_0;
	wire w_dff_B_GTop6alx5_0;
	wire w_dff_B_isnod7H93_0;
	wire w_dff_B_hYN94gql4_0;
	wire w_dff_B_TYDkehFz3_0;
	wire w_dff_B_1R1iEFKn7_0;
	wire w_dff_B_hc0wCGcQ3_0;
	wire w_dff_B_0kox4D0f8_0;
	wire w_dff_B_fSunZdvb8_0;
	wire w_dff_B_br6IXRvj1_0;
	wire w_dff_B_s0DMGbSC6_0;
	wire w_dff_B_9lKQl8VW9_0;
	wire w_dff_B_yke4QKy12_0;
	wire w_dff_B_aah6ulmI7_0;
	wire w_dff_B_04M2D68W8_0;
	wire w_dff_B_rZvBXlim7_0;
	wire w_dff_B_zD41bNiG7_0;
	wire w_dff_B_lkQPnXny1_0;
	wire w_dff_B_AMlU3bff0_0;
	wire w_dff_B_ih9AxHTJ2_0;
	wire w_dff_B_xvhPIzqt6_0;
	wire w_dff_B_Uchh0Bas0_0;
	wire w_dff_B_PEgbaQ6E7_0;
	wire w_dff_B_K10P0fQr3_0;
	wire w_dff_B_P15aDoTu2_0;
	wire w_dff_B_SCaMJe4u7_0;
	wire w_dff_B_Nd7Fues73_0;
	wire w_dff_B_Z1ueymbs7_0;
	wire w_dff_B_nuJkUSOm2_0;
	wire w_dff_B_XaRpYCAd6_0;
	wire w_dff_B_6Df0zqfJ4_0;
	wire w_dff_B_dtFngcJS1_0;
	wire w_dff_B_dCvPrrXy3_0;
	wire w_dff_B_ihgSkygg2_0;
	wire w_dff_B_DwdcsoqK5_0;
	wire w_dff_B_vZ2dBD3F2_0;
	wire w_dff_B_ALJcwdXU8_0;
	wire w_dff_B_h4lfzINb3_0;
	wire w_dff_B_uVu2H0jH1_0;
	wire w_dff_B_oK6EAMFd5_0;
	wire w_dff_B_szAD2Rne6_0;
	wire w_dff_B_V8BeWNtC3_0;
	wire w_dff_B_pgydElYJ8_0;
	wire w_dff_B_LDp9m6jh6_0;
	wire w_dff_B_253hTXaZ8_0;
	wire w_dff_B_shgoIpAe2_0;
	wire w_dff_B_JjU0kbAT0_0;
	wire w_dff_B_Nyf1tyS72_0;
	wire w_dff_B_EVOVZtAd7_0;
	wire w_dff_B_lSezfx319_0;
	wire w_dff_B_EeTvjZ833_0;
	wire w_dff_B_E1nOEVE68_0;
	wire w_dff_B_1mmysII87_0;
	wire w_dff_B_Z1nAeDqs7_0;
	wire w_dff_B_jiqGkYTx0_0;
	wire w_dff_B_QXsj9D0E1_0;
	wire w_dff_B_NLb17XNZ9_0;
	wire w_dff_B_6IIpGqTX5_0;
	wire w_dff_B_0vwFyDdw3_0;
	wire w_dff_B_NkBj7BcQ2_0;
	wire w_dff_B_DZerjOCU2_0;
	wire w_dff_B_uKsc8miY8_0;
	wire w_dff_B_jZYYgkKq1_0;
	wire w_dff_B_H8ickXxF7_0;
	wire w_dff_B_A8pRry767_0;
	wire w_dff_B_GWmOgk2V0_0;
	wire w_dff_B_rnm3cO2Q2_0;
	wire w_dff_B_0eO1sDOQ9_0;
	wire w_dff_B_Arb0ROCA4_0;
	wire w_dff_B_hETQgg9q5_0;
	wire w_dff_B_bbwbSTyP8_0;
	wire w_dff_B_X6Gir7cf1_0;
	wire w_dff_B_L7CtLO6o6_0;
	wire w_dff_B_K2JIZ6ZI1_0;
	wire w_dff_B_uMd8AryD2_0;
	wire w_dff_B_GrNRIarL1_0;
	wire w_dff_B_5Rpe5MKA3_0;
	wire w_dff_B_25jn3B9A7_0;
	wire w_dff_B_P9VzfJ9J9_0;
	wire w_dff_B_KN53MaCM1_0;
	wire w_dff_B_2XawnBzw4_0;
	wire w_dff_B_k9FJG9Do2_0;
	wire w_dff_B_TArSJXeg5_0;
	wire w_dff_B_qY3vTnCq5_0;
	wire w_dff_B_toHFjzK43_0;
	wire w_dff_B_UtQbRfGY3_0;
	wire w_dff_B_qnPVfik00_0;
	wire w_dff_B_ZGFz7tMl6_0;
	wire w_dff_B_Ml1jO7Ic0_0;
	wire w_dff_B_QRC27lcQ5_0;
	wire w_dff_B_FJ4WNLA39_0;
	wire w_dff_B_Lbc52OQP8_0;
	wire w_dff_B_Y5afw0ZB8_0;
	wire w_dff_B_LpU5trMT0_0;
	wire w_dff_B_eRQIpvKz8_0;
	wire w_dff_B_0Z7hCwz47_0;
	wire w_dff_B_o4Svj9Vj3_0;
	wire w_dff_B_HIERyfhj0_0;
	wire w_dff_B_s6bl0pUF6_0;
	wire w_dff_B_BbZnq9aI1_0;
	wire w_dff_B_AVz3ik2a7_0;
	wire w_dff_B_6W81Yg0D1_0;
	wire w_dff_B_LJocUySI0_0;
	wire w_dff_B_CZKMbq7t9_0;
	wire w_dff_B_C9QaqcpL4_0;
	wire w_dff_B_bFVN0Qed9_1;
	wire w_dff_B_HSBDnd5v7_1;
	wire w_dff_B_gWDft5LV8_1;
	wire w_dff_B_KN7UEH1d6_1;
	wire w_dff_B_IoYVsFeU4_1;
	wire w_dff_B_Ko52s5Hi0_1;
	wire w_dff_B_wXNFg8NA9_1;
	wire w_dff_B_cAPzcAbI6_1;
	wire w_dff_B_HyxNk1rF9_1;
	wire w_dff_B_leZFrgEh6_1;
	wire w_dff_B_DN4pplCX5_1;
	wire w_dff_B_xXPd4XLS3_1;
	wire w_dff_B_pY5DrhnD9_1;
	wire w_dff_B_ntVByL6G6_1;
	wire w_dff_B_3RDIIUFW3_1;
	wire w_dff_B_jtTKa6VD9_1;
	wire w_dff_B_nhs8tYnY3_1;
	wire w_dff_B_vZ7nAznE0_1;
	wire w_dff_B_kY1zTx6Z7_1;
	wire w_dff_B_jWKVX2Bb9_1;
	wire w_dff_B_Pm851Ymt1_1;
	wire w_dff_B_k3WSiMb69_1;
	wire w_dff_B_z7az5cOA5_1;
	wire w_dff_B_9jCkwasi9_1;
	wire w_dff_B_8SKuRgD08_1;
	wire w_dff_B_WQO8gDls8_1;
	wire w_dff_B_LGoYdaZg6_1;
	wire w_dff_B_AbSDOs336_1;
	wire w_dff_B_osv36UEq6_1;
	wire w_dff_B_4SZA163P8_1;
	wire w_dff_B_UesKWUS14_1;
	wire w_dff_B_gNPo2dzH8_1;
	wire w_dff_B_ODqNautq3_1;
	wire w_dff_B_jgcXi6pZ7_1;
	wire w_dff_B_IXx4TcSe3_1;
	wire w_dff_B_Ur0U9lGf8_1;
	wire w_dff_B_L0XYUffd4_1;
	wire w_dff_B_Tlk9GDzm3_1;
	wire w_dff_B_cJvfzVON1_1;
	wire w_dff_B_k4Z7XCDJ6_1;
	wire w_dff_B_vv4ZDUyh9_1;
	wire w_dff_B_8iqiTTzx3_1;
	wire w_dff_B_QP7WfLZS6_1;
	wire w_dff_B_3IwECteJ0_1;
	wire w_dff_B_ZxEmBrr27_1;
	wire w_dff_B_YaaUE8zO1_1;
	wire w_dff_B_hYH7VbdA0_1;
	wire w_dff_B_5x7Mp2Lx7_1;
	wire w_dff_B_H83HnVeM9_1;
	wire w_dff_B_VDg9BtRN8_1;
	wire w_dff_B_5D26V9wt3_1;
	wire w_dff_B_r9KLOEtj1_1;
	wire w_dff_B_94rmknWS0_1;
	wire w_dff_B_LF4wsQji1_1;
	wire w_dff_B_5IofoIbI0_1;
	wire w_dff_B_wwyyc6zB6_1;
	wire w_dff_B_5sj9XZwc7_1;
	wire w_dff_B_yOAEe7IH2_1;
	wire w_dff_B_IHkCUzU34_1;
	wire w_dff_B_XaAe5UmA1_1;
	wire w_dff_B_cBESAYhG1_1;
	wire w_dff_B_JceMSJ8I2_1;
	wire w_dff_B_1zQC9HOu0_1;
	wire w_dff_B_gv1fmmBW4_1;
	wire w_dff_B_5IyfkmIV0_1;
	wire w_dff_B_hDpjD3FY8_1;
	wire w_dff_B_taonE3Hk0_1;
	wire w_dff_B_P747L8WS5_1;
	wire w_dff_B_LciAk2zr4_1;
	wire w_dff_B_tMB6SiXu4_1;
	wire w_dff_B_Qf773v530_1;
	wire w_dff_B_HtvzNgK15_1;
	wire w_dff_B_uIqRUHnO5_1;
	wire w_dff_B_uTzEIOu43_1;
	wire w_dff_B_zpmvfynv2_1;
	wire w_dff_B_QSY34u1X5_1;
	wire w_dff_B_JGl9DQes3_1;
	wire w_dff_B_uQaNhLDe6_1;
	wire w_dff_B_YISJmDUl2_1;
	wire w_dff_B_qZMmcBxe9_1;
	wire w_dff_B_xgwmgfx24_1;
	wire w_dff_B_ymgcPYnU6_1;
	wire w_dff_B_Ne01avRW2_1;
	wire w_dff_B_oH1sQqBu3_1;
	wire w_dff_B_ImXwsVgn7_1;
	wire w_dff_B_5QWsOaar3_1;
	wire w_dff_B_8zszqGh32_1;
	wire w_dff_B_d0QARxKa6_1;
	wire w_dff_B_ZOjvBBCA8_1;
	wire w_dff_B_tAY6tdAr0_1;
	wire w_dff_B_ss4fYgPG1_1;
	wire w_dff_B_PJbZVXZ39_1;
	wire w_dff_B_UaA2q3QW0_1;
	wire w_dff_B_zXuXbAg94_1;
	wire w_dff_B_kg0aVgPW1_1;
	wire w_dff_B_qXDo8E5j9_1;
	wire w_dff_B_FvOkDus66_1;
	wire w_dff_B_ORaioyxN3_1;
	wire w_dff_B_ENSVAwRI7_1;
	wire w_dff_B_ZjnuHFbu0_1;
	wire w_dff_B_2rSl9HV12_1;
	wire w_dff_B_yqZitFZj4_1;
	wire w_dff_B_ANVA01PR5_1;
	wire w_dff_B_gvgNoTLP7_1;
	wire w_dff_B_nwX3XGbn2_1;
	wire w_dff_B_JdwvomK95_1;
	wire w_dff_B_D1eNItdK8_1;
	wire w_dff_B_BMacVM8n4_1;
	wire w_dff_B_8deQ3RaC2_0;
	wire w_dff_B_LZL8vLaM7_0;
	wire w_dff_B_zCoLkU1W2_0;
	wire w_dff_B_Sjo7tciE3_0;
	wire w_dff_B_1TG6dtgk4_0;
	wire w_dff_B_sDs86Ikx2_0;
	wire w_dff_B_z6PUWR8z2_0;
	wire w_dff_B_slbc8sEX2_0;
	wire w_dff_B_0abywTc20_0;
	wire w_dff_B_Nxc9yxPb6_0;
	wire w_dff_B_Tt9BHrTK8_0;
	wire w_dff_B_3UweyeU27_0;
	wire w_dff_B_oA47j4YF9_0;
	wire w_dff_B_xvD4s9IZ5_0;
	wire w_dff_B_GtepwspG4_0;
	wire w_dff_B_wtsmixzP9_0;
	wire w_dff_B_xqHyY5m65_0;
	wire w_dff_B_CHnjgpIv6_0;
	wire w_dff_B_h0Bglps86_0;
	wire w_dff_B_DSK2wJdV5_0;
	wire w_dff_B_4DyduRFv9_0;
	wire w_dff_B_5ZiI9uBl4_0;
	wire w_dff_B_2QQkHLUC3_0;
	wire w_dff_B_kVDEMbO49_0;
	wire w_dff_B_pNVNweeH6_0;
	wire w_dff_B_crShAWPu0_0;
	wire w_dff_B_AFVvm6CW1_0;
	wire w_dff_B_NuyCH00F5_0;
	wire w_dff_B_Aj2o48NQ3_0;
	wire w_dff_B_16tKTqVr7_0;
	wire w_dff_B_oB0TbDs02_0;
	wire w_dff_B_PlGcQ7vB6_0;
	wire w_dff_B_aNbozymt3_0;
	wire w_dff_B_vPiBtOGQ3_0;
	wire w_dff_B_kLl3hZl09_0;
	wire w_dff_B_3mgr8RtU0_0;
	wire w_dff_B_iva8plW76_0;
	wire w_dff_B_KC5tcFuK8_0;
	wire w_dff_B_7jJfqrHH6_0;
	wire w_dff_B_fHA6wVgn7_0;
	wire w_dff_B_yj70ytnF2_0;
	wire w_dff_B_rVhPHQmC7_0;
	wire w_dff_B_Kh6NGusd7_0;
	wire w_dff_B_7kj2tfp01_0;
	wire w_dff_B_AyE07pT04_0;
	wire w_dff_B_dvzjfVSt7_0;
	wire w_dff_B_CDxmYxKr7_0;
	wire w_dff_B_XS4DU9tw4_0;
	wire w_dff_B_2bF4EF9Z5_0;
	wire w_dff_B_a5K1c3Bo8_0;
	wire w_dff_B_53qxiWqd2_0;
	wire w_dff_B_U8Cra25v2_0;
	wire w_dff_B_goAZPxvf2_0;
	wire w_dff_B_9jiy1SYX1_0;
	wire w_dff_B_HkdNSkfs4_0;
	wire w_dff_B_HZ9we5PL3_0;
	wire w_dff_B_fRQ8TtFq2_0;
	wire w_dff_B_CSKFWIas1_0;
	wire w_dff_B_hbmTbEWi8_0;
	wire w_dff_B_XeCv7cN38_0;
	wire w_dff_B_O85L9Tk05_0;
	wire w_dff_B_PUUBZXtq3_0;
	wire w_dff_B_Z6CSjm9I1_0;
	wire w_dff_B_KpPV1p3s6_0;
	wire w_dff_B_0XYGvi6T6_0;
	wire w_dff_B_zecfbCZG9_0;
	wire w_dff_B_MSyEWdwW9_0;
	wire w_dff_B_zFxI68wS8_0;
	wire w_dff_B_xayqS21i1_0;
	wire w_dff_B_vtoGmsN28_0;
	wire w_dff_B_g513HMU55_0;
	wire w_dff_B_3ZnT0QOE9_0;
	wire w_dff_B_e61vckDh0_0;
	wire w_dff_B_aiVXdiAC4_0;
	wire w_dff_B_7hFEtFMA2_0;
	wire w_dff_B_Ym1v7XJ56_0;
	wire w_dff_B_wySjj1zN5_0;
	wire w_dff_B_Hdu3tnUH8_0;
	wire w_dff_B_H3Xc0WrE1_0;
	wire w_dff_B_KLDaTWHJ2_0;
	wire w_dff_B_YEwlDs3x4_0;
	wire w_dff_B_nmLBtDhF4_0;
	wire w_dff_B_M91nXk6g2_0;
	wire w_dff_B_QiLGjchY4_0;
	wire w_dff_B_c15dFlmW2_0;
	wire w_dff_B_Re2vektU1_0;
	wire w_dff_B_taHjV3hZ3_0;
	wire w_dff_B_ZjJR6ow80_0;
	wire w_dff_B_wkcVbRyr8_0;
	wire w_dff_B_cIvUoP7m0_0;
	wire w_dff_B_w7N7Xmkr3_0;
	wire w_dff_B_NlewqK2G4_0;
	wire w_dff_B_0bBG0e9p3_0;
	wire w_dff_B_FgaDW4t81_0;
	wire w_dff_B_spk9uJHE8_0;
	wire w_dff_B_hxXzLpOP1_0;
	wire w_dff_B_cIoKiF850_0;
	wire w_dff_B_l2or20CR9_0;
	wire w_dff_B_zvXq4FAs6_0;
	wire w_dff_B_v6DhjobE1_0;
	wire w_dff_B_6QK2jsIT8_0;
	wire w_dff_B_Tt7TPj6N2_0;
	wire w_dff_B_a35uhzbZ9_0;
	wire w_dff_B_4c2yPfRT6_0;
	wire w_dff_B_G9smq10s2_0;
	wire w_dff_B_cJVNtqKO5_0;
	wire w_dff_B_bJrEKCoO4_0;
	wire w_dff_B_ISqqPwDn9_0;
	wire w_dff_B_sNp6ShSz7_1;
	wire w_dff_B_kJFprg0r5_1;
	wire w_dff_B_dINkKPxx1_1;
	wire w_dff_B_W2v9cfAu0_1;
	wire w_dff_B_DUGQt5qn9_1;
	wire w_dff_B_73CLID8z0_1;
	wire w_dff_B_oRCSPhpP4_1;
	wire w_dff_B_ZlMj3kR61_1;
	wire w_dff_B_KX2LgwsS9_1;
	wire w_dff_B_vuUqtOWm6_1;
	wire w_dff_B_Auwu0XXj6_1;
	wire w_dff_B_KB4ZfdLj2_1;
	wire w_dff_B_HngxO0Uj0_1;
	wire w_dff_B_2rAo27ek3_1;
	wire w_dff_B_1yuMyIff2_1;
	wire w_dff_B_bwOPwuYv2_1;
	wire w_dff_B_MTk4h14h7_1;
	wire w_dff_B_d7WeVBrS5_1;
	wire w_dff_B_FrWhF4Cz9_1;
	wire w_dff_B_hJUC7WUN2_1;
	wire w_dff_B_CxKcba1o0_1;
	wire w_dff_B_6vUiK6130_1;
	wire w_dff_B_mjDMx4ul9_1;
	wire w_dff_B_tYKbNTyW2_1;
	wire w_dff_B_A3wnPson6_1;
	wire w_dff_B_j9Jg9zDH3_1;
	wire w_dff_B_QYaEuE2X5_1;
	wire w_dff_B_tJoPPfBW7_1;
	wire w_dff_B_BcfQLpAq2_1;
	wire w_dff_B_fGdEvZyL9_1;
	wire w_dff_B_lt2uSuFn2_1;
	wire w_dff_B_eOwKKlvL6_1;
	wire w_dff_B_Kb5eZCR04_1;
	wire w_dff_B_HmmRyGwv2_1;
	wire w_dff_B_9gwTku3U3_1;
	wire w_dff_B_Ob6jiuSn0_1;
	wire w_dff_B_8HEUaogz5_1;
	wire w_dff_B_Ii1lU8fb6_1;
	wire w_dff_B_DtZdYFLU3_1;
	wire w_dff_B_AFAxx7y61_1;
	wire w_dff_B_6sH0kz1P9_1;
	wire w_dff_B_ljYpIwnb2_1;
	wire w_dff_B_AFjh8EhR3_1;
	wire w_dff_B_OMRA4bCC0_1;
	wire w_dff_B_GVnabYUt7_1;
	wire w_dff_B_Xl68Rniz2_1;
	wire w_dff_B_3zNbge5I6_1;
	wire w_dff_B_5mWCnpXf3_1;
	wire w_dff_B_80a8rMpB4_1;
	wire w_dff_B_LcBIPVk52_1;
	wire w_dff_B_wkt9KDvl9_1;
	wire w_dff_B_eXYZBust9_1;
	wire w_dff_B_UtRC0vIv2_1;
	wire w_dff_B_eSV6K7Yu5_1;
	wire w_dff_B_XHpJ1g3i7_1;
	wire w_dff_B_tMf2eBS41_1;
	wire w_dff_B_sRPbSVa98_1;
	wire w_dff_B_Cv2hXfG22_1;
	wire w_dff_B_0jGqNUTS9_1;
	wire w_dff_B_XmiSzfrw1_1;
	wire w_dff_B_jDHWSs2W6_1;
	wire w_dff_B_1GmN4tGU8_1;
	wire w_dff_B_Dc44K48P5_1;
	wire w_dff_B_LCACFbPS9_1;
	wire w_dff_B_r6Eb3GYB8_1;
	wire w_dff_B_exURoR631_1;
	wire w_dff_B_6sERNQHn1_1;
	wire w_dff_B_DwNa9UBF4_1;
	wire w_dff_B_Fv0wd9zd4_1;
	wire w_dff_B_frV9Zoog4_1;
	wire w_dff_B_mUuqq02s2_1;
	wire w_dff_B_2Kp7A3SX6_1;
	wire w_dff_B_p73HMTjL8_1;
	wire w_dff_B_2AFVpd2l3_1;
	wire w_dff_B_KJa3pqMR3_1;
	wire w_dff_B_T5YsAIWP2_1;
	wire w_dff_B_jzbrsWDm2_1;
	wire w_dff_B_GMzh451l4_1;
	wire w_dff_B_ycIpniEc3_1;
	wire w_dff_B_cZ3tMkVU1_1;
	wire w_dff_B_0W3BNHKB2_1;
	wire w_dff_B_D9zm9QL63_1;
	wire w_dff_B_RjxutSIJ3_1;
	wire w_dff_B_LehWGyme1_1;
	wire w_dff_B_IzGGpkGF4_1;
	wire w_dff_B_hG9jjS9b1_1;
	wire w_dff_B_Rb3hY0CN6_1;
	wire w_dff_B_c9CPLuWJ3_1;
	wire w_dff_B_PHTDjAR21_1;
	wire w_dff_B_OK4Cbq2N3_1;
	wire w_dff_B_SCKtyKSI8_1;
	wire w_dff_B_XJeY6c0D5_1;
	wire w_dff_B_SHLLeqqr4_1;
	wire w_dff_B_uP8GFxyD6_1;
	wire w_dff_B_iijEBp3U2_1;
	wire w_dff_B_sTOnEMhS8_1;
	wire w_dff_B_GblG97w47_1;
	wire w_dff_B_A36wNVHx6_1;
	wire w_dff_B_USqdnUqB5_1;
	wire w_dff_B_KEVR8POg8_1;
	wire w_dff_B_JxTT3yEo9_1;
	wire w_dff_B_MaMNWOS70_1;
	wire w_dff_B_JELEf7Sw8_1;
	wire w_dff_B_tHHHLE2j9_1;
	wire w_dff_B_VSuAiR5z5_1;
	wire w_dff_B_vJde0YQf8_1;
	wire w_dff_B_XTpaCHU28_1;
	wire w_dff_B_pomrhoKX3_0;
	wire w_dff_B_baCcp0oq8_0;
	wire w_dff_B_XOUVEuQM9_0;
	wire w_dff_B_iIRRvqXo2_0;
	wire w_dff_B_4ZDaoUx90_0;
	wire w_dff_B_uZ8VJFde1_0;
	wire w_dff_B_fFfeAyoS5_0;
	wire w_dff_B_vrRmLZtB7_0;
	wire w_dff_B_34i4JCfy4_0;
	wire w_dff_B_e0H4W5wI5_0;
	wire w_dff_B_MxyzzHXk8_0;
	wire w_dff_B_ID4vhbKP0_0;
	wire w_dff_B_lCi4MSn69_0;
	wire w_dff_B_qJifAUfl6_0;
	wire w_dff_B_z8m25sLp9_0;
	wire w_dff_B_gxbjblo96_0;
	wire w_dff_B_3yvVl3l50_0;
	wire w_dff_B_QABOeMfz6_0;
	wire w_dff_B_YZSuemMn5_0;
	wire w_dff_B_omGWFeWB4_0;
	wire w_dff_B_CRL12axe7_0;
	wire w_dff_B_SiufHU2S1_0;
	wire w_dff_B_FKrAPskI5_0;
	wire w_dff_B_ee2L7aO76_0;
	wire w_dff_B_1hrnuihP5_0;
	wire w_dff_B_0iKcyB6a0_0;
	wire w_dff_B_Me5b1PGq4_0;
	wire w_dff_B_oyEvkl4H7_0;
	wire w_dff_B_gDCeEwbQ4_0;
	wire w_dff_B_3iU4jI8b5_0;
	wire w_dff_B_gLWVFxL25_0;
	wire w_dff_B_xZNckrrA1_0;
	wire w_dff_B_0BLRsOe23_0;
	wire w_dff_B_KcUXHiAH5_0;
	wire w_dff_B_nKmcGCwL3_0;
	wire w_dff_B_hR41QYdD6_0;
	wire w_dff_B_D48VAFVc8_0;
	wire w_dff_B_J36eJ6qG6_0;
	wire w_dff_B_DpDdnZDY4_0;
	wire w_dff_B_xoxvbiiT5_0;
	wire w_dff_B_jXZa1wDf4_0;
	wire w_dff_B_SKy6bEDi4_0;
	wire w_dff_B_i2msDnMm6_0;
	wire w_dff_B_QlPHvjD14_0;
	wire w_dff_B_WWffVfOq9_0;
	wire w_dff_B_gByYrllJ4_0;
	wire w_dff_B_SoARTfZF5_0;
	wire w_dff_B_CTyDAvbT0_0;
	wire w_dff_B_pAICIYvP2_0;
	wire w_dff_B_QDJNz9Tm3_0;
	wire w_dff_B_ztoT0opx6_0;
	wire w_dff_B_JxICGcUt9_0;
	wire w_dff_B_myoXOUum0_0;
	wire w_dff_B_E5W8l5If0_0;
	wire w_dff_B_Ft7QBMg95_0;
	wire w_dff_B_qiBKn6Kg7_0;
	wire w_dff_B_sTK66WS13_0;
	wire w_dff_B_mV9AOvXr2_0;
	wire w_dff_B_btB1mEKx3_0;
	wire w_dff_B_0wtbn10a4_0;
	wire w_dff_B_nxcFl2bI5_0;
	wire w_dff_B_JVtan3Qz4_0;
	wire w_dff_B_IKBhzfGn2_0;
	wire w_dff_B_xBRBwFRm5_0;
	wire w_dff_B_xxfuCkD96_0;
	wire w_dff_B_BNuSu2Ox9_0;
	wire w_dff_B_BUFmk3Cl2_0;
	wire w_dff_B_3RqGMbzc2_0;
	wire w_dff_B_KF1K7Qfd5_0;
	wire w_dff_B_PoVtOAqm5_0;
	wire w_dff_B_5AHgWFZh4_0;
	wire w_dff_B_Mlpajz0y5_0;
	wire w_dff_B_sOaWQa9i1_0;
	wire w_dff_B_P5NahKIs3_0;
	wire w_dff_B_jpCQUsBu6_0;
	wire w_dff_B_cOIt78Ng7_0;
	wire w_dff_B_cvbQq8QU1_0;
	wire w_dff_B_rdF4XIZ41_0;
	wire w_dff_B_qrvbyXEo2_0;
	wire w_dff_B_6qNdAErD0_0;
	wire w_dff_B_RjWmkJTb4_0;
	wire w_dff_B_zFAUXzQW6_0;
	wire w_dff_B_YAx3gkgB4_0;
	wire w_dff_B_VbXmrZlD6_0;
	wire w_dff_B_gO0JsDvz1_0;
	wire w_dff_B_ONFmeABu9_0;
	wire w_dff_B_LKNqEdxf1_0;
	wire w_dff_B_aJ5CKMW35_0;
	wire w_dff_B_McxDPGt43_0;
	wire w_dff_B_wZAa0PfI2_0;
	wire w_dff_B_iuIi85S93_0;
	wire w_dff_B_xHnBmQFG1_0;
	wire w_dff_B_TWSyTdm77_0;
	wire w_dff_B_sZjpofVw6_0;
	wire w_dff_B_NsxZKiOO6_0;
	wire w_dff_B_oHPeoiAT6_0;
	wire w_dff_B_KT71PfDa5_0;
	wire w_dff_B_AKO3xROQ2_0;
	wire w_dff_B_Ew6PCfXS9_0;
	wire w_dff_B_cdTRIFdt5_0;
	wire w_dff_B_jEqqGPwr8_0;
	wire w_dff_B_DmEpAyja3_0;
	wire w_dff_B_upEAL2tH7_0;
	wire w_dff_B_pZy9ywM63_0;
	wire w_dff_B_RSVqasus7_0;
	wire w_dff_B_UcLcfnEH4_0;
	wire w_dff_B_rQs1ywwY3_0;
	wire w_dff_B_ziLTM7Mv0_1;
	wire w_dff_B_JppgMvTB2_1;
	wire w_dff_B_5zp088EI0_1;
	wire w_dff_B_unK8V57A2_1;
	wire w_dff_B_JXqkLCk36_1;
	wire w_dff_B_zkiwK9dx7_1;
	wire w_dff_B_bVzakFPN1_1;
	wire w_dff_B_rV34xDOI2_1;
	wire w_dff_B_HaBCZKri7_1;
	wire w_dff_B_uvp4uylE9_1;
	wire w_dff_B_uUagZVog8_1;
	wire w_dff_B_pdrJnaYb7_1;
	wire w_dff_B_W7msf6WW5_1;
	wire w_dff_B_wm3x5N3G3_1;
	wire w_dff_B_DYvucooa8_1;
	wire w_dff_B_71pfdEjU0_1;
	wire w_dff_B_j5GrO96V5_1;
	wire w_dff_B_Q8RSgHzH0_1;
	wire w_dff_B_qFIK46ND6_1;
	wire w_dff_B_i1GCqMrP5_1;
	wire w_dff_B_quhWUEMl4_1;
	wire w_dff_B_9QliUMWL2_1;
	wire w_dff_B_nWU6iosP7_1;
	wire w_dff_B_3munYuCa3_1;
	wire w_dff_B_QMnnd6x60_1;
	wire w_dff_B_n5KH8bNc1_1;
	wire w_dff_B_2Fa5s8bH3_1;
	wire w_dff_B_X9InJHaX0_1;
	wire w_dff_B_0mtu47He4_1;
	wire w_dff_B_sdshQXGJ1_1;
	wire w_dff_B_kc1a2mbG4_1;
	wire w_dff_B_krp0yNrd0_1;
	wire w_dff_B_SuZoj0JQ9_1;
	wire w_dff_B_jF7oMYoN4_1;
	wire w_dff_B_84jn34NM7_1;
	wire w_dff_B_GEe2zmwU5_1;
	wire w_dff_B_o7y7ePYZ2_1;
	wire w_dff_B_DmdVwadQ2_1;
	wire w_dff_B_s0Zdac2D0_1;
	wire w_dff_B_d6Jw8NPt8_1;
	wire w_dff_B_VJ2ycxkd5_1;
	wire w_dff_B_yBKYa5tC2_1;
	wire w_dff_B_WwlNXJEA9_1;
	wire w_dff_B_VNuqwP7b9_1;
	wire w_dff_B_MDKUS8Pu5_1;
	wire w_dff_B_O0H5SKCC9_1;
	wire w_dff_B_XPoRxyEJ4_1;
	wire w_dff_B_iIYXcv9I7_1;
	wire w_dff_B_cGpMQEVd7_1;
	wire w_dff_B_A8motzwi4_1;
	wire w_dff_B_XSAuaGPJ8_1;
	wire w_dff_B_jVEmj9RX3_1;
	wire w_dff_B_pBRve9tm9_1;
	wire w_dff_B_RW1RUIVr6_1;
	wire w_dff_B_clRH3NjO5_1;
	wire w_dff_B_3al7Lryt9_1;
	wire w_dff_B_qM4pHBPP0_1;
	wire w_dff_B_3VREC1Y76_1;
	wire w_dff_B_oaf5EENS7_1;
	wire w_dff_B_frKGwZtW4_1;
	wire w_dff_B_WKOv21Kw1_1;
	wire w_dff_B_Mn5eYnsu7_1;
	wire w_dff_B_rExBtcga4_1;
	wire w_dff_B_8J85daFQ8_1;
	wire w_dff_B_ygfmDo1b7_1;
	wire w_dff_B_KvnvNw4R9_1;
	wire w_dff_B_7QLk3Ih44_1;
	wire w_dff_B_FZMpEpWQ3_1;
	wire w_dff_B_DSFliSsu4_1;
	wire w_dff_B_878ETSX64_1;
	wire w_dff_B_J93ErqUJ7_1;
	wire w_dff_B_NC08NBCG9_1;
	wire w_dff_B_uGapLXyd4_1;
	wire w_dff_B_dVujtNXs2_1;
	wire w_dff_B_1MsgKfBg1_1;
	wire w_dff_B_LFvfSxTj5_1;
	wire w_dff_B_0IluKIdd7_1;
	wire w_dff_B_U1BsWREF0_1;
	wire w_dff_B_0fLTMB6u3_1;
	wire w_dff_B_DbXPuAl33_1;
	wire w_dff_B_cXuSid1T2_1;
	wire w_dff_B_OvgwmrmJ3_1;
	wire w_dff_B_aRnlNRVT0_1;
	wire w_dff_B_dhbKDunM6_1;
	wire w_dff_B_IuWdFmHJ7_1;
	wire w_dff_B_AlI43VYf3_1;
	wire w_dff_B_fQDL9vth7_1;
	wire w_dff_B_TDh6r4uK3_1;
	wire w_dff_B_ANVQHhKt8_1;
	wire w_dff_B_lodUgsRh3_1;
	wire w_dff_B_1ynOt1R01_1;
	wire w_dff_B_RF6UXE7p6_1;
	wire w_dff_B_h0Ac4r5T2_1;
	wire w_dff_B_YJVK6OyD2_1;
	wire w_dff_B_ib1jukmZ7_1;
	wire w_dff_B_p1guUylt9_1;
	wire w_dff_B_yREBVfuC2_1;
	wire w_dff_B_bE3hAoWJ1_1;
	wire w_dff_B_fMz32HQt4_1;
	wire w_dff_B_DhLmN5zo3_1;
	wire w_dff_B_2F0z03f70_1;
	wire w_dff_B_JP2X0w3b5_1;
	wire w_dff_B_X4nabGQI4_1;
	wire w_dff_B_9FOoyu9q4_1;
	wire w_dff_B_r6CCakIW7_1;
	wire w_dff_B_P8u9UvcR2_1;
	wire w_dff_B_29wQ6VC00_0;
	wire w_dff_B_95cyNm3X7_0;
	wire w_dff_B_0pkdsav03_0;
	wire w_dff_B_VpEujyx84_0;
	wire w_dff_B_DcU3epRh2_0;
	wire w_dff_B_3psZYbWh2_0;
	wire w_dff_B_mekTVtDp1_0;
	wire w_dff_B_AFdrrYpY1_0;
	wire w_dff_B_YlpETyDe2_0;
	wire w_dff_B_LtoigXS11_0;
	wire w_dff_B_lnAMYQyf8_0;
	wire w_dff_B_gOMiQl1u6_0;
	wire w_dff_B_LS5sbzif0_0;
	wire w_dff_B_i6BHeBTb2_0;
	wire w_dff_B_mIN3d78w1_0;
	wire w_dff_B_Ye3TTZcF1_0;
	wire w_dff_B_UHk4d3Nb3_0;
	wire w_dff_B_ipLikkw02_0;
	wire w_dff_B_2WoFnMBh7_0;
	wire w_dff_B_QGd9Swlp7_0;
	wire w_dff_B_Wu4FZKd05_0;
	wire w_dff_B_Vmrp97804_0;
	wire w_dff_B_s9xnr6Pe2_0;
	wire w_dff_B_dyBrehPs0_0;
	wire w_dff_B_yR7n3T0A8_0;
	wire w_dff_B_zdOnvQdf9_0;
	wire w_dff_B_HJGwPcYa6_0;
	wire w_dff_B_aWjKBzaV0_0;
	wire w_dff_B_N3vJtnMD5_0;
	wire w_dff_B_jXdoLGA43_0;
	wire w_dff_B_rTapqOOZ4_0;
	wire w_dff_B_IearAhPt4_0;
	wire w_dff_B_ac09Q1978_0;
	wire w_dff_B_SbLJRpJj8_0;
	wire w_dff_B_aTemLyWC2_0;
	wire w_dff_B_dm1uwraT0_0;
	wire w_dff_B_a33z0QD25_0;
	wire w_dff_B_cmh8g24U9_0;
	wire w_dff_B_378AIIW14_0;
	wire w_dff_B_qo1I6EWH6_0;
	wire w_dff_B_pmlBNUhK6_0;
	wire w_dff_B_DKcVkPuE7_0;
	wire w_dff_B_EFQSQSk04_0;
	wire w_dff_B_J6XpONsp2_0;
	wire w_dff_B_ucZBbHJ59_0;
	wire w_dff_B_HnAuSiv57_0;
	wire w_dff_B_8QqAeA4W4_0;
	wire w_dff_B_zDbyTkJw2_0;
	wire w_dff_B_HXOPrIN76_0;
	wire w_dff_B_bblFn69R8_0;
	wire w_dff_B_wpTdDqGr0_0;
	wire w_dff_B_GxbX4Cab4_0;
	wire w_dff_B_VTwEPMHl6_0;
	wire w_dff_B_gctUakBU0_0;
	wire w_dff_B_AgrqmcjW6_0;
	wire w_dff_B_tyPWyxTl2_0;
	wire w_dff_B_syhUo1cF2_0;
	wire w_dff_B_HPMSueB41_0;
	wire w_dff_B_eNs7Ry896_0;
	wire w_dff_B_j4lf7bYQ0_0;
	wire w_dff_B_ycY1IlSU3_0;
	wire w_dff_B_FS5rStR61_0;
	wire w_dff_B_hBpdjPmG0_0;
	wire w_dff_B_hrLVEVHK7_0;
	wire w_dff_B_nSITv95n9_0;
	wire w_dff_B_8CZYt4qo7_0;
	wire w_dff_B_at2HwvLi3_0;
	wire w_dff_B_9ygDQVEG6_0;
	wire w_dff_B_fZS1BtOV9_0;
	wire w_dff_B_xELxgy789_0;
	wire w_dff_B_U09uoXR96_0;
	wire w_dff_B_ccBwl2gZ4_0;
	wire w_dff_B_ayx3pwgB2_0;
	wire w_dff_B_YzWvd2OB0_0;
	wire w_dff_B_9famPQo49_0;
	wire w_dff_B_5lZb1mgG9_0;
	wire w_dff_B_stvrphk09_0;
	wire w_dff_B_17cXq4X46_0;
	wire w_dff_B_7vIoF1Qc0_0;
	wire w_dff_B_PknXh2HB1_0;
	wire w_dff_B_mVbVs9gG9_0;
	wire w_dff_B_05A0b1yf0_0;
	wire w_dff_B_GW1rbx2z6_0;
	wire w_dff_B_fAmRyzbQ8_0;
	wire w_dff_B_OWtdytaD9_0;
	wire w_dff_B_FuTTeeuX1_0;
	wire w_dff_B_JFml0BBk6_0;
	wire w_dff_B_Q8dQkKOd8_0;
	wire w_dff_B_OKNTs6kD0_0;
	wire w_dff_B_frAbasL66_0;
	wire w_dff_B_cX2qw0Z04_0;
	wire w_dff_B_tlsd6gJ52_0;
	wire w_dff_B_9jvOhias7_0;
	wire w_dff_B_CDenmHyS5_0;
	wire w_dff_B_wNaBnSyQ9_0;
	wire w_dff_B_Dw3ibZ2E1_0;
	wire w_dff_B_ztDSc3fz3_0;
	wire w_dff_B_GNKytxFO3_0;
	wire w_dff_B_AUYca1hl2_0;
	wire w_dff_B_WifhNf3n2_0;
	wire w_dff_B_8t38Yj9U5_0;
	wire w_dff_B_whkEqGju9_0;
	wire w_dff_B_1m4hZpYQ7_0;
	wire w_dff_B_r0fBw0CL6_0;
	wire w_dff_B_dFlcaupd5_0;
	wire w_dff_B_OmEewm5z6_0;
	wire w_dff_B_JUUjm9XO7_1;
	wire w_dff_B_ugGZOQGc4_1;
	wire w_dff_B_aaS0NVKT3_1;
	wire w_dff_B_Mag5RAyv4_1;
	wire w_dff_B_nvlWEInm8_1;
	wire w_dff_B_PyDChZAP3_1;
	wire w_dff_B_bTtMVvBi8_1;
	wire w_dff_B_6ipDwSkz7_1;
	wire w_dff_B_fvOamn8j9_1;
	wire w_dff_B_W2BfAWBI3_1;
	wire w_dff_B_ZDPbW5Ud3_1;
	wire w_dff_B_66A2Y7jx4_1;
	wire w_dff_B_rv9Pg3UY2_1;
	wire w_dff_B_9EsukJjn0_1;
	wire w_dff_B_4NZxd1G13_1;
	wire w_dff_B_9ILGoqVG4_1;
	wire w_dff_B_mKx1xcwS8_1;
	wire w_dff_B_XG1AWsmw1_1;
	wire w_dff_B_AXlW9Mng1_1;
	wire w_dff_B_0DBCNyFy1_1;
	wire w_dff_B_pbbm2fMz0_1;
	wire w_dff_B_5WUfzSRl8_1;
	wire w_dff_B_Ajc4k1FC6_1;
	wire w_dff_B_NMq6UkGZ4_1;
	wire w_dff_B_ruVKIaDw4_1;
	wire w_dff_B_tmlXTsKA8_1;
	wire w_dff_B_zEGyTuKT3_1;
	wire w_dff_B_k3xLNKhO6_1;
	wire w_dff_B_5zoKq7im8_1;
	wire w_dff_B_K0pL3mhG2_1;
	wire w_dff_B_1Hy5iJpa9_1;
	wire w_dff_B_rf3tRyeL7_1;
	wire w_dff_B_JJx3DrRV3_1;
	wire w_dff_B_hFXxEyka4_1;
	wire w_dff_B_qLlHQfSq7_1;
	wire w_dff_B_BLywJjcP4_1;
	wire w_dff_B_g31FVAto9_1;
	wire w_dff_B_KKO4CKx77_1;
	wire w_dff_B_n9wBg8Et9_1;
	wire w_dff_B_SIJUhVml3_1;
	wire w_dff_B_YjRPGwob9_1;
	wire w_dff_B_tdYXr8Ue5_1;
	wire w_dff_B_2z6Xm6jk5_1;
	wire w_dff_B_g8eVitQw0_1;
	wire w_dff_B_vTYPfvl81_1;
	wire w_dff_B_UhU2nAds0_1;
	wire w_dff_B_zUPJRTCT3_1;
	wire w_dff_B_jBODE7sf7_1;
	wire w_dff_B_mvsYVhxU3_1;
	wire w_dff_B_VewwZZgh6_1;
	wire w_dff_B_tdA69xAC3_1;
	wire w_dff_B_TLG4aLnL8_1;
	wire w_dff_B_kdqW6lY40_1;
	wire w_dff_B_tqVtFNve8_1;
	wire w_dff_B_Rw87Cy3u6_1;
	wire w_dff_B_xRC3sDTn0_1;
	wire w_dff_B_SqEdrAAx5_1;
	wire w_dff_B_m3C534ZW5_1;
	wire w_dff_B_ewtK5mJ97_1;
	wire w_dff_B_2GYbysjL2_1;
	wire w_dff_B_uJXetQbI6_1;
	wire w_dff_B_5p2Uwr378_1;
	wire w_dff_B_hSYqCOIf6_1;
	wire w_dff_B_pdGh6DDR5_1;
	wire w_dff_B_FU5WNjug3_1;
	wire w_dff_B_KeLjHwOo0_1;
	wire w_dff_B_E7WElCnm2_1;
	wire w_dff_B_iG6VsE8q8_1;
	wire w_dff_B_ttvzSkoR7_1;
	wire w_dff_B_yIVzYWdx2_1;
	wire w_dff_B_iX6WM2vv0_1;
	wire w_dff_B_k2zSO25V4_1;
	wire w_dff_B_kQ2MLCEU3_1;
	wire w_dff_B_vaP66fZx3_1;
	wire w_dff_B_rXWxyiOV1_1;
	wire w_dff_B_UcXmYYVp5_1;
	wire w_dff_B_fRNd6gK80_1;
	wire w_dff_B_knJcnDia6_1;
	wire w_dff_B_cBgUkfGc0_1;
	wire w_dff_B_GlqGkDHz4_1;
	wire w_dff_B_3Kd18oPV1_1;
	wire w_dff_B_cJyLxk779_1;
	wire w_dff_B_8IXRVP938_1;
	wire w_dff_B_83sdgtFi5_1;
	wire w_dff_B_2mSg8kJD8_1;
	wire w_dff_B_ItvNy3gS8_1;
	wire w_dff_B_zLaIRpRP6_1;
	wire w_dff_B_RZjEuioS1_1;
	wire w_dff_B_58PEEVGP1_1;
	wire w_dff_B_cVjkXz2t7_1;
	wire w_dff_B_dyNkmlfy8_1;
	wire w_dff_B_3oPKDMJ41_1;
	wire w_dff_B_cj7yehJr8_1;
	wire w_dff_B_NHEvEhQa4_1;
	wire w_dff_B_72IqebV26_1;
	wire w_dff_B_ETzYWIxJ7_1;
	wire w_dff_B_BErVn2rC2_1;
	wire w_dff_B_LQNZ0gjG7_1;
	wire w_dff_B_bLOwMUpj1_1;
	wire w_dff_B_c7EIYxgT3_1;
	wire w_dff_B_R7FpmBCw1_1;
	wire w_dff_B_3dT33HA32_1;
	wire w_dff_B_w0HbWKII0_1;
	wire w_dff_B_r6KoXOnJ3_1;
	wire w_dff_B_opUbMGB49_1;
	wire w_dff_B_sopoYNE76_0;
	wire w_dff_B_0eGGHMlu3_0;
	wire w_dff_B_ZR57yI1Z8_0;
	wire w_dff_B_gm6BWLov8_0;
	wire w_dff_B_4pl9aWMf4_0;
	wire w_dff_B_leq9d4qL3_0;
	wire w_dff_B_duTWINYO1_0;
	wire w_dff_B_vB43oCBE1_0;
	wire w_dff_B_MatlSzIi3_0;
	wire w_dff_B_iclNGsXo1_0;
	wire w_dff_B_aomv0Fqh8_0;
	wire w_dff_B_fRw8MDn73_0;
	wire w_dff_B_wsODJM8E6_0;
	wire w_dff_B_zcawso2S7_0;
	wire w_dff_B_nNxa7va32_0;
	wire w_dff_B_JXSP59g56_0;
	wire w_dff_B_zr89SJry3_0;
	wire w_dff_B_anzB9ocb7_0;
	wire w_dff_B_0Ha5SysI8_0;
	wire w_dff_B_lai9bFW44_0;
	wire w_dff_B_Bcn4AlFl6_0;
	wire w_dff_B_qFwM2U1V6_0;
	wire w_dff_B_1KrcOf3k7_0;
	wire w_dff_B_ubAMaq8Q2_0;
	wire w_dff_B_QmfOAmNk3_0;
	wire w_dff_B_LdaOF7WW8_0;
	wire w_dff_B_nGiKIEOw8_0;
	wire w_dff_B_NjEYtfRS3_0;
	wire w_dff_B_s7NG6gVf6_0;
	wire w_dff_B_joyQhANH8_0;
	wire w_dff_B_MlBXG8Bf0_0;
	wire w_dff_B_sALFBYPA4_0;
	wire w_dff_B_4l5xCi2h6_0;
	wire w_dff_B_E4ajtg692_0;
	wire w_dff_B_Mv7yniZq2_0;
	wire w_dff_B_4hxiN5Og8_0;
	wire w_dff_B_Odmd7uzu3_0;
	wire w_dff_B_YLWAYSjY3_0;
	wire w_dff_B_sRipMn8T2_0;
	wire w_dff_B_vg4Gf6lg3_0;
	wire w_dff_B_k3pfXuHF7_0;
	wire w_dff_B_eXGVUCuG5_0;
	wire w_dff_B_33YCekoC2_0;
	wire w_dff_B_87DN9wnS0_0;
	wire w_dff_B_0baUcS5p7_0;
	wire w_dff_B_0nZm7Sdy8_0;
	wire w_dff_B_mk7sEWke6_0;
	wire w_dff_B_fIYAB21S1_0;
	wire w_dff_B_nD5jHmAZ0_0;
	wire w_dff_B_u3xd9PFr8_0;
	wire w_dff_B_lH8XCHC72_0;
	wire w_dff_B_DbuqCntg1_0;
	wire w_dff_B_3OlBQqIe5_0;
	wire w_dff_B_QjbMqjXH9_0;
	wire w_dff_B_WMDwby1R5_0;
	wire w_dff_B_Mfct0s1v0_0;
	wire w_dff_B_6DT5gzTT1_0;
	wire w_dff_B_L4UskE3C7_0;
	wire w_dff_B_bp8t7ZE46_0;
	wire w_dff_B_17eGOwd79_0;
	wire w_dff_B_Kmw9BlMH2_0;
	wire w_dff_B_aLWfetc56_0;
	wire w_dff_B_A0xtEKIQ1_0;
	wire w_dff_B_b5VN4p2H0_0;
	wire w_dff_B_B2RodtiT9_0;
	wire w_dff_B_l0O7bCit6_0;
	wire w_dff_B_fzHBgx1X3_0;
	wire w_dff_B_u8OwdW1U7_0;
	wire w_dff_B_l6H5NuBV9_0;
	wire w_dff_B_bJFMvIC76_0;
	wire w_dff_B_4r81DgCj2_0;
	wire w_dff_B_eZdSR4q52_0;
	wire w_dff_B_6Js46pfn6_0;
	wire w_dff_B_QVqjuezl8_0;
	wire w_dff_B_2qPGzj4G6_0;
	wire w_dff_B_8yTE7N012_0;
	wire w_dff_B_n41vpbyU5_0;
	wire w_dff_B_jKZdXvcN2_0;
	wire w_dff_B_us1IIPa28_0;
	wire w_dff_B_HgbC4rMv0_0;
	wire w_dff_B_y5QRl9T57_0;
	wire w_dff_B_xWkFxl7Y9_0;
	wire w_dff_B_J3Ebs7Pn4_0;
	wire w_dff_B_ZW4dlhnT8_0;
	wire w_dff_B_jR8AcVOh7_0;
	wire w_dff_B_sKchNxYA3_0;
	wire w_dff_B_RpgGaSTt0_0;
	wire w_dff_B_Xd3u2lNs0_0;
	wire w_dff_B_Ix4QkzFX5_0;
	wire w_dff_B_YRvKzS0T1_0;
	wire w_dff_B_CtZzvZcf9_0;
	wire w_dff_B_IOd6Jlkx8_0;
	wire w_dff_B_z8sCIKSH0_0;
	wire w_dff_B_Dp7MEQVe0_0;
	wire w_dff_B_hf9tfxjv8_0;
	wire w_dff_B_VwSvjwLC5_0;
	wire w_dff_B_A13X0RKi1_0;
	wire w_dff_B_69jdkr2X4_0;
	wire w_dff_B_rOPpMwfn2_0;
	wire w_dff_B_m3eUTp5i8_0;
	wire w_dff_B_KHpBvGl34_0;
	wire w_dff_B_fE6COzPy2_0;
	wire w_dff_B_BsF4gmAC7_0;
	wire w_dff_B_NEKHiB8j6_0;
	wire w_dff_B_IzQy6DU01_0;
	wire w_dff_B_HJ6lVrTb0_1;
	wire w_dff_B_HkwNynPJ9_1;
	wire w_dff_B_a6fYzwqM7_1;
	wire w_dff_B_W8m1CUOh6_1;
	wire w_dff_B_ZcbKwOBE0_1;
	wire w_dff_B_xkLvKH0P2_1;
	wire w_dff_B_5uwaqEZk0_1;
	wire w_dff_B_GrGmLSE58_1;
	wire w_dff_B_JYWOJZGU1_1;
	wire w_dff_B_gLcofKyE3_1;
	wire w_dff_B_Eim1cGsx4_1;
	wire w_dff_B_Y5O0ij5F6_1;
	wire w_dff_B_ofxVtgf67_1;
	wire w_dff_B_7diVCkaV2_1;
	wire w_dff_B_pMh7tMWD6_1;
	wire w_dff_B_fmQNbMFh3_1;
	wire w_dff_B_2q9IsWxb7_1;
	wire w_dff_B_RACxajck2_1;
	wire w_dff_B_aA4nJKB04_1;
	wire w_dff_B_HFsZEE1F0_1;
	wire w_dff_B_GXQsBL7t1_1;
	wire w_dff_B_UHuE8k1I4_1;
	wire w_dff_B_THM0uF6f7_1;
	wire w_dff_B_PGzZk2nL0_1;
	wire w_dff_B_0PKHyQ317_1;
	wire w_dff_B_KR5q2HIy6_1;
	wire w_dff_B_RydqBP1p9_1;
	wire w_dff_B_Y22SUoGK6_1;
	wire w_dff_B_yHwmgnXE8_1;
	wire w_dff_B_G2gFgPUO7_1;
	wire w_dff_B_8dit25wa2_1;
	wire w_dff_B_90FidDOm4_1;
	wire w_dff_B_NUURd4pn0_1;
	wire w_dff_B_u5sGMKrC3_1;
	wire w_dff_B_kdSgblys0_1;
	wire w_dff_B_08D9uipu3_1;
	wire w_dff_B_N8AFf5hJ8_1;
	wire w_dff_B_pvAnsIew8_1;
	wire w_dff_B_iZzPuJhS9_1;
	wire w_dff_B_SKauuycG8_1;
	wire w_dff_B_0rekuKli1_1;
	wire w_dff_B_OTPE3UwP1_1;
	wire w_dff_B_BwG9m3In4_1;
	wire w_dff_B_DTH32o8H2_1;
	wire w_dff_B_SKS1RfRB5_1;
	wire w_dff_B_rtdb7BK05_1;
	wire w_dff_B_YTvAxG3Q3_1;
	wire w_dff_B_J7rm1AFB5_1;
	wire w_dff_B_f6BytXrQ8_1;
	wire w_dff_B_y0Lqhrfb8_1;
	wire w_dff_B_djeOODWI7_1;
	wire w_dff_B_uliD3X7z1_1;
	wire w_dff_B_vbnuL4pR8_1;
	wire w_dff_B_atxwU3iB6_1;
	wire w_dff_B_v2jjmF4A6_1;
	wire w_dff_B_wDE1PLUR8_1;
	wire w_dff_B_3H8ZsqCZ7_1;
	wire w_dff_B_YXFcmwWs9_1;
	wire w_dff_B_LHKzxVsH5_1;
	wire w_dff_B_9sC2MBoT7_1;
	wire w_dff_B_jt4JEY7O0_1;
	wire w_dff_B_Rr9mJgn85_1;
	wire w_dff_B_MJ99dW0b5_1;
	wire w_dff_B_CeGqMrfq0_1;
	wire w_dff_B_gU7WsBuK3_1;
	wire w_dff_B_J15nntqZ7_1;
	wire w_dff_B_WM8n7qpW1_1;
	wire w_dff_B_3e0YboH48_1;
	wire w_dff_B_ocQ8UxSp3_1;
	wire w_dff_B_BfuFaR1d6_1;
	wire w_dff_B_07ZFZeeX9_1;
	wire w_dff_B_qvImErpT1_1;
	wire w_dff_B_Q3Hnkmqj8_1;
	wire w_dff_B_dBKNN4PM7_1;
	wire w_dff_B_SsCfeRrd7_1;
	wire w_dff_B_beMOGVr14_1;
	wire w_dff_B_yAAegxo65_1;
	wire w_dff_B_Wq0Zzxw80_1;
	wire w_dff_B_O2Ynz6V51_1;
	wire w_dff_B_IfGIIln55_1;
	wire w_dff_B_jOvVRSwm4_1;
	wire w_dff_B_uSbS7F3I1_1;
	wire w_dff_B_fWQu58r08_1;
	wire w_dff_B_5UACoK6j5_1;
	wire w_dff_B_8GVe9j025_1;
	wire w_dff_B_ngKcFJy79_1;
	wire w_dff_B_jZBtkeVy6_1;
	wire w_dff_B_at6GQTXv8_1;
	wire w_dff_B_dHtBVGU23_1;
	wire w_dff_B_KT2elHrl6_1;
	wire w_dff_B_t8xirMW40_1;
	wire w_dff_B_8urqMdUE3_1;
	wire w_dff_B_U53R5WUf2_1;
	wire w_dff_B_8l0aIOKA3_1;
	wire w_dff_B_zTD1JsW25_1;
	wire w_dff_B_kN8FSfJV4_1;
	wire w_dff_B_dO9uMtjr9_1;
	wire w_dff_B_E1yN1Em58_1;
	wire w_dff_B_joxinVQu3_1;
	wire w_dff_B_mvlqfd8N7_1;
	wire w_dff_B_OBSvF7gD7_1;
	wire w_dff_B_GAkGCBbr8_1;
	wire w_dff_B_LVI8cSBi3_1;
	wire w_dff_B_8BuCOaXp1_1;
	wire w_dff_B_LI1muG7X8_0;
	wire w_dff_B_egmYcb4j8_0;
	wire w_dff_B_HfoUMNU27_0;
	wire w_dff_B_leG3NFcU0_0;
	wire w_dff_B_eoOSUF5U2_0;
	wire w_dff_B_qCOw17NJ7_0;
	wire w_dff_B_8qF4oLp59_0;
	wire w_dff_B_sxL51aso2_0;
	wire w_dff_B_7JLICGiQ1_0;
	wire w_dff_B_ZkmMBWjr2_0;
	wire w_dff_B_b77E3YUu2_0;
	wire w_dff_B_Dhb34zyI0_0;
	wire w_dff_B_Hjcx7EUi8_0;
	wire w_dff_B_8N8u9eN09_0;
	wire w_dff_B_sI6GdHPP9_0;
	wire w_dff_B_ZnyUfvvH2_0;
	wire w_dff_B_AFG806F59_0;
	wire w_dff_B_XEjjwvcA2_0;
	wire w_dff_B_iWd2cdY69_0;
	wire w_dff_B_HWk4etxo7_0;
	wire w_dff_B_fghiXM9g4_0;
	wire w_dff_B_D4NjwCDp5_0;
	wire w_dff_B_muBPgzAl6_0;
	wire w_dff_B_n9eQtlS83_0;
	wire w_dff_B_3OjDPwgO6_0;
	wire w_dff_B_EjSBSspc0_0;
	wire w_dff_B_4mltlmjF4_0;
	wire w_dff_B_IWj7SB838_0;
	wire w_dff_B_r5X8XCsD4_0;
	wire w_dff_B_q9kbxnmm7_0;
	wire w_dff_B_DefmhDpX7_0;
	wire w_dff_B_eVJhgeTY2_0;
	wire w_dff_B_fsDrF0vM9_0;
	wire w_dff_B_0tQLHKNs6_0;
	wire w_dff_B_63DrpowM4_0;
	wire w_dff_B_YF2Zahn03_0;
	wire w_dff_B_Ey5PKPlS0_0;
	wire w_dff_B_3oz5WrYv2_0;
	wire w_dff_B_op98yKlS5_0;
	wire w_dff_B_mcsgzguU6_0;
	wire w_dff_B_tLYShEHZ0_0;
	wire w_dff_B_6S6tvjRH1_0;
	wire w_dff_B_jplVcPNJ0_0;
	wire w_dff_B_Qhxplqxv4_0;
	wire w_dff_B_9RVKo98I3_0;
	wire w_dff_B_IpDIJSNC8_0;
	wire w_dff_B_fNMQA6Vj7_0;
	wire w_dff_B_7S6qvp1Z9_0;
	wire w_dff_B_3IngINET2_0;
	wire w_dff_B_qecdS1VE6_0;
	wire w_dff_B_pXJIDVD74_0;
	wire w_dff_B_LeWZ4lhu7_0;
	wire w_dff_B_Rr7I6YOX2_0;
	wire w_dff_B_dIapvW9Q9_0;
	wire w_dff_B_UBSKpJyw0_0;
	wire w_dff_B_nZt4nX8L4_0;
	wire w_dff_B_K5UkPmBo3_0;
	wire w_dff_B_11k69KHb6_0;
	wire w_dff_B_YWR2y9KU3_0;
	wire w_dff_B_3gak01wb9_0;
	wire w_dff_B_m7ehzTDk3_0;
	wire w_dff_B_NEgDjvWA6_0;
	wire w_dff_B_ffiE4x1C0_0;
	wire w_dff_B_r4Lt7h438_0;
	wire w_dff_B_ycii6xhC3_0;
	wire w_dff_B_m9B9t76Q1_0;
	wire w_dff_B_EhxT2tTV8_0;
	wire w_dff_B_oXh7r5bD6_0;
	wire w_dff_B_QNMF3iAj8_0;
	wire w_dff_B_xzEZGPjV0_0;
	wire w_dff_B_VeDMNrz93_0;
	wire w_dff_B_N9e2qZxf6_0;
	wire w_dff_B_UJ4GEoou0_0;
	wire w_dff_B_EwpETrgg3_0;
	wire w_dff_B_X3WEBxMB5_0;
	wire w_dff_B_zZOEJAJj1_0;
	wire w_dff_B_cTcYrSu97_0;
	wire w_dff_B_S9bhGfzF2_0;
	wire w_dff_B_aYcVxeT15_0;
	wire w_dff_B_ap8LFJF55_0;
	wire w_dff_B_LgZlzfhn2_0;
	wire w_dff_B_1CkPniOb4_0;
	wire w_dff_B_EE51UNaF4_0;
	wire w_dff_B_NdNDA36K1_0;
	wire w_dff_B_pwtiHkDR5_0;
	wire w_dff_B_A0JEfiZv9_0;
	wire w_dff_B_cTLRItGK3_0;
	wire w_dff_B_Z75AlfVW4_0;
	wire w_dff_B_SRJLofgB3_0;
	wire w_dff_B_aW6HM6pg6_0;
	wire w_dff_B_l5e3fs230_0;
	wire w_dff_B_WK19l0Xf4_0;
	wire w_dff_B_SdlSwMMp4_0;
	wire w_dff_B_zHS1dsAy1_0;
	wire w_dff_B_ODRF0p9l2_0;
	wire w_dff_B_dDPTvBqu6_0;
	wire w_dff_B_ZhfzBMLk8_0;
	wire w_dff_B_NwPrT38H6_0;
	wire w_dff_B_s6THB9RY5_0;
	wire w_dff_B_uYhXifJN1_0;
	wire w_dff_B_Rd53p9bN8_0;
	wire w_dff_B_GpMM8Ys45_0;
	wire w_dff_B_GLfXb2JO5_0;
	wire w_dff_B_lEwdgnFZ1_0;
	wire w_dff_B_fMaqATnV1_1;
	wire w_dff_B_LczZ2fgD9_1;
	wire w_dff_B_gLfPJs2k8_1;
	wire w_dff_B_z5jm6e2X4_1;
	wire w_dff_B_wLqXc8Eh1_1;
	wire w_dff_B_SIIPbB0c8_1;
	wire w_dff_B_4AM10sF09_1;
	wire w_dff_B_pd3vKY0h6_1;
	wire w_dff_B_0zMj7xj78_1;
	wire w_dff_B_GMOIlGUD1_1;
	wire w_dff_B_Ywh1KOHj5_1;
	wire w_dff_B_b8Wb6kc55_1;
	wire w_dff_B_Xr7aWDK08_1;
	wire w_dff_B_7DXUnPAy7_1;
	wire w_dff_B_LGzYi79Y5_1;
	wire w_dff_B_WM1q6cKc9_1;
	wire w_dff_B_FLPkBcsF3_1;
	wire w_dff_B_i6NWirmn7_1;
	wire w_dff_B_Iw7HvS4c2_1;
	wire w_dff_B_RCjBSv8K1_1;
	wire w_dff_B_OD2pNKbW2_1;
	wire w_dff_B_5TNBViO54_1;
	wire w_dff_B_QWOOMs9C9_1;
	wire w_dff_B_ztaprmkK6_1;
	wire w_dff_B_SEkV0cOO8_1;
	wire w_dff_B_LabkkwI49_1;
	wire w_dff_B_swE72mfm0_1;
	wire w_dff_B_N2aQWDGN4_1;
	wire w_dff_B_IRWKwa7E2_1;
	wire w_dff_B_Bl3593RG5_1;
	wire w_dff_B_ExjWkram7_1;
	wire w_dff_B_da6W8suy0_1;
	wire w_dff_B_337b6h9I7_1;
	wire w_dff_B_YlBZKN7q4_1;
	wire w_dff_B_r02HyutI4_1;
	wire w_dff_B_0wmaVvbr9_1;
	wire w_dff_B_J2tPZ8I21_1;
	wire w_dff_B_RvfKmCGE5_1;
	wire w_dff_B_iT8shnqG8_1;
	wire w_dff_B_elOvhyhE2_1;
	wire w_dff_B_0OAcjmcj5_1;
	wire w_dff_B_DB2vbbvL0_1;
	wire w_dff_B_crSU5yex0_1;
	wire w_dff_B_BNfHpmXF5_1;
	wire w_dff_B_SAf1DYnP0_1;
	wire w_dff_B_PdDpRUEt9_1;
	wire w_dff_B_PzdBbhbu4_1;
	wire w_dff_B_23cEm7iu6_1;
	wire w_dff_B_dfyFE99p5_1;
	wire w_dff_B_wnOzjbsO2_1;
	wire w_dff_B_x64VKMPF9_1;
	wire w_dff_B_WGIs6CrK3_1;
	wire w_dff_B_NDHVr71m4_1;
	wire w_dff_B_jU6j1S9I3_1;
	wire w_dff_B_bBW133xo7_1;
	wire w_dff_B_j1gTpmQG3_1;
	wire w_dff_B_nu4wcaFe2_1;
	wire w_dff_B_d5ww5trd6_1;
	wire w_dff_B_vxSjOymS8_1;
	wire w_dff_B_BLHDNoIe6_1;
	wire w_dff_B_JjtDlUbO9_1;
	wire w_dff_B_caypdeIr4_1;
	wire w_dff_B_UcCUvmwO2_1;
	wire w_dff_B_VjqQEqSk0_1;
	wire w_dff_B_Z0I00MCQ1_1;
	wire w_dff_B_CINVDIGM1_1;
	wire w_dff_B_caZpxfEV1_1;
	wire w_dff_B_xhE3hfVr6_1;
	wire w_dff_B_DdifxwCM3_1;
	wire w_dff_B_FI4q1Rkk4_1;
	wire w_dff_B_hkOWJ4OF2_1;
	wire w_dff_B_vLWd5O6c7_1;
	wire w_dff_B_NZd7Lg3u7_1;
	wire w_dff_B_0Jq5KK763_1;
	wire w_dff_B_CSNzOrFa7_1;
	wire w_dff_B_aOAiC69s0_1;
	wire w_dff_B_8cz2WsSi6_1;
	wire w_dff_B_vNNqIT0k0_1;
	wire w_dff_B_am6QIwSN5_1;
	wire w_dff_B_D7UeQCsY6_1;
	wire w_dff_B_WcqaJ2jn3_1;
	wire w_dff_B_it3M0FVM2_1;
	wire w_dff_B_SsrF3jtx4_1;
	wire w_dff_B_5rekw1lX6_1;
	wire w_dff_B_enA95C2F9_1;
	wire w_dff_B_0LDZx56T0_1;
	wire w_dff_B_LYGoZoG09_1;
	wire w_dff_B_2PWh1po04_1;
	wire w_dff_B_3VfNJbtd4_1;
	wire w_dff_B_U3MKcYr33_1;
	wire w_dff_B_JZl7bUXj2_1;
	wire w_dff_B_EtMzor9e5_1;
	wire w_dff_B_09753Men2_1;
	wire w_dff_B_SRo4UDe63_1;
	wire w_dff_B_TdRn8OID0_1;
	wire w_dff_B_9r3EyRnt9_1;
	wire w_dff_B_RV449SGC0_1;
	wire w_dff_B_TrlzIL7K6_1;
	wire w_dff_B_Rv29iDqX4_1;
	wire w_dff_B_EY4FzuFX5_1;
	wire w_dff_B_TtaQ10hk0_1;
	wire w_dff_B_ndlMbPLS5_1;
	wire w_dff_B_GI8cjqgr1_1;
	wire w_dff_B_e6lz4nSd7_0;
	wire w_dff_B_QP1HIkg01_0;
	wire w_dff_B_ej58O5Cg7_0;
	wire w_dff_B_c1OS9FIc1_0;
	wire w_dff_B_UxUQjaGq6_0;
	wire w_dff_B_3IGJFiRl8_0;
	wire w_dff_B_BYw3f24c1_0;
	wire w_dff_B_GCMdQVue7_0;
	wire w_dff_B_joe4ZUSL2_0;
	wire w_dff_B_WhWE3lOn2_0;
	wire w_dff_B_XHUCO0FG0_0;
	wire w_dff_B_QN1rs2GM8_0;
	wire w_dff_B_6zu9grEN8_0;
	wire w_dff_B_A8dbrEFY8_0;
	wire w_dff_B_75cvf8bH4_0;
	wire w_dff_B_cKKOVBjd7_0;
	wire w_dff_B_qtYDwSyy0_0;
	wire w_dff_B_YVmHd4Qa5_0;
	wire w_dff_B_uzPZcTdB4_0;
	wire w_dff_B_LrDCyk2e9_0;
	wire w_dff_B_22TBqFiZ7_0;
	wire w_dff_B_uOgljo4N5_0;
	wire w_dff_B_YmNN57yQ9_0;
	wire w_dff_B_Q2Omy1N32_0;
	wire w_dff_B_p3PFj3k72_0;
	wire w_dff_B_xnokRXv86_0;
	wire w_dff_B_Vo3ZFT8P1_0;
	wire w_dff_B_XSpMbBMq5_0;
	wire w_dff_B_eSd5pEHh6_0;
	wire w_dff_B_qiRjCs3g2_0;
	wire w_dff_B_M9DkvZxp0_0;
	wire w_dff_B_W4DMuDQH8_0;
	wire w_dff_B_2bo03jgs9_0;
	wire w_dff_B_WLNjEQDx7_0;
	wire w_dff_B_I4SY4MPK0_0;
	wire w_dff_B_fJliKFbw1_0;
	wire w_dff_B_MisHAYvD7_0;
	wire w_dff_B_Pa2q46Wb6_0;
	wire w_dff_B_OMLl9mby1_0;
	wire w_dff_B_ezRSevQT2_0;
	wire w_dff_B_iJCBvH4N1_0;
	wire w_dff_B_hzOjO8wT3_0;
	wire w_dff_B_vZED4JAN8_0;
	wire w_dff_B_BpALgirx8_0;
	wire w_dff_B_eKWoX3Js4_0;
	wire w_dff_B_oxXNSdov8_0;
	wire w_dff_B_L5epyQPQ9_0;
	wire w_dff_B_QOkAJBUi8_0;
	wire w_dff_B_VmPocXDV2_0;
	wire w_dff_B_CSBB6bv62_0;
	wire w_dff_B_1yL7wUaL1_0;
	wire w_dff_B_v3NoQaqj4_0;
	wire w_dff_B_YZYvtNtZ8_0;
	wire w_dff_B_ePVZN5wl8_0;
	wire w_dff_B_kLgxzR3X1_0;
	wire w_dff_B_xGpjraOR2_0;
	wire w_dff_B_iXyjUXoo0_0;
	wire w_dff_B_fmJptW6U6_0;
	wire w_dff_B_e2nzqi1Y5_0;
	wire w_dff_B_TakbssWp7_0;
	wire w_dff_B_zW8bEz0W9_0;
	wire w_dff_B_vOcimzpI5_0;
	wire w_dff_B_ra5hyIxk1_0;
	wire w_dff_B_j9rX7nar7_0;
	wire w_dff_B_ii5VuVHj2_0;
	wire w_dff_B_KvW3IjMc5_0;
	wire w_dff_B_ILjjkCgc1_0;
	wire w_dff_B_OSjB8WzJ2_0;
	wire w_dff_B_FSfjnVL29_0;
	wire w_dff_B_EkDOfp9y1_0;
	wire w_dff_B_Iiumm3eR9_0;
	wire w_dff_B_z4Gd4soa7_0;
	wire w_dff_B_BKECVXw49_0;
	wire w_dff_B_6I1gYRnV6_0;
	wire w_dff_B_yhQaCsgT9_0;
	wire w_dff_B_T3heKXXc3_0;
	wire w_dff_B_VAsiJoMd5_0;
	wire w_dff_B_18tnDX7V4_0;
	wire w_dff_B_MtOzHtfH3_0;
	wire w_dff_B_QprVbgpW7_0;
	wire w_dff_B_P2XHdSjZ6_0;
	wire w_dff_B_kRXfaSXs7_0;
	wire w_dff_B_eAO4Gal12_0;
	wire w_dff_B_ZsIhPlMI7_0;
	wire w_dff_B_Pj30zCB80_0;
	wire w_dff_B_AZ6NrpXW4_0;
	wire w_dff_B_6Lf2J6yg9_0;
	wire w_dff_B_DcjTsauK2_0;
	wire w_dff_B_rjautiqH2_0;
	wire w_dff_B_jnCsBWIj1_0;
	wire w_dff_B_aGNge5uQ5_0;
	wire w_dff_B_RDjbSkuj4_0;
	wire w_dff_B_MpVggaHh6_0;
	wire w_dff_B_4Ys50if07_0;
	wire w_dff_B_i1o0bDT82_0;
	wire w_dff_B_YniSy8aB5_0;
	wire w_dff_B_lck7UEvD2_0;
	wire w_dff_B_VU70DES38_0;
	wire w_dff_B_X0285ssm4_0;
	wire w_dff_B_ms0rmQyj3_0;
	wire w_dff_B_CyFTqv8S8_0;
	wire w_dff_B_ap8PWfKR3_0;
	wire w_dff_B_ISBRX9kG4_0;
	wire w_dff_B_Uc08YVKY5_1;
	wire w_dff_B_JNr4uM3S9_1;
	wire w_dff_B_9h76yTlC5_1;
	wire w_dff_B_Y0ZwGY1U7_1;
	wire w_dff_B_Jlfr7Qml8_1;
	wire w_dff_B_gM9vXp6G5_1;
	wire w_dff_B_kRwJcoUK7_1;
	wire w_dff_B_u1EZgqHf5_1;
	wire w_dff_B_ushofyMb6_1;
	wire w_dff_B_rpfBrktU3_1;
	wire w_dff_B_w8AP4Hsl0_1;
	wire w_dff_B_Ktjdo2Ns7_1;
	wire w_dff_B_9Pr1Z7lQ3_1;
	wire w_dff_B_KnE6zQED7_1;
	wire w_dff_B_3waKnxTt1_1;
	wire w_dff_B_DA1DP4Xd1_1;
	wire w_dff_B_MWTz8cpq3_1;
	wire w_dff_B_eiujRRXT5_1;
	wire w_dff_B_nhnZyIlb3_1;
	wire w_dff_B_PKKnjG4f4_1;
	wire w_dff_B_QIQrqbdL7_1;
	wire w_dff_B_F0X5ybIW2_1;
	wire w_dff_B_nVXWQ8082_1;
	wire w_dff_B_I7uVEbnw8_1;
	wire w_dff_B_ER6QXdeH7_1;
	wire w_dff_B_SqcqtdqA5_1;
	wire w_dff_B_iaPnzZ829_1;
	wire w_dff_B_J5R3M07j5_1;
	wire w_dff_B_8n1HrsKJ1_1;
	wire w_dff_B_AtOdfwoZ3_1;
	wire w_dff_B_mVlI4WCx0_1;
	wire w_dff_B_GvCzs7de9_1;
	wire w_dff_B_xpU7rWtj2_1;
	wire w_dff_B_7ZeUikwx8_1;
	wire w_dff_B_HlQd3npy0_1;
	wire w_dff_B_timINsCF3_1;
	wire w_dff_B_DXrU1c7V2_1;
	wire w_dff_B_GeIx1So29_1;
	wire w_dff_B_hdMRwFTk8_1;
	wire w_dff_B_3fpwr5H99_1;
	wire w_dff_B_V8LVNEXd4_1;
	wire w_dff_B_nsx127bK8_1;
	wire w_dff_B_uJq1wClp0_1;
	wire w_dff_B_z0YzCurh0_1;
	wire w_dff_B_qGAIjcRr7_1;
	wire w_dff_B_xPHGV7GV4_1;
	wire w_dff_B_DUlgI1nE0_1;
	wire w_dff_B_wa9rmqy67_1;
	wire w_dff_B_DqfPtgYI7_1;
	wire w_dff_B_YK0ZpN1t9_1;
	wire w_dff_B_w6EAt5FU2_1;
	wire w_dff_B_QzbbztSb7_1;
	wire w_dff_B_AT81xLg10_1;
	wire w_dff_B_9MNWekpF7_1;
	wire w_dff_B_FS5iXezl4_1;
	wire w_dff_B_k6rbrxsV2_1;
	wire w_dff_B_YFAysJ3K5_1;
	wire w_dff_B_YHznMhmx8_1;
	wire w_dff_B_E5LZrr773_1;
	wire w_dff_B_8XugjQEe6_1;
	wire w_dff_B_YGeeYzEU1_1;
	wire w_dff_B_f02OrG1J2_1;
	wire w_dff_B_hr9zR0DI5_1;
	wire w_dff_B_O2uIn6pg7_1;
	wire w_dff_B_Sl5BtnIU1_1;
	wire w_dff_B_ntE6AoX12_1;
	wire w_dff_B_anVdO9Di7_1;
	wire w_dff_B_KtpZAMZl6_1;
	wire w_dff_B_PQoiDZgy6_1;
	wire w_dff_B_2hYxQ0tg1_1;
	wire w_dff_B_31yiIhMV2_1;
	wire w_dff_B_c0EmdxH57_1;
	wire w_dff_B_vptXheoI2_1;
	wire w_dff_B_nXwVgPLW3_1;
	wire w_dff_B_JuDNfIgZ0_1;
	wire w_dff_B_ozJvyKhd1_1;
	wire w_dff_B_nqLzc8YF2_1;
	wire w_dff_B_VftNLq0q5_1;
	wire w_dff_B_4wMeMZnu6_1;
	wire w_dff_B_KKWyLyDV6_1;
	wire w_dff_B_R8iTdVWC7_1;
	wire w_dff_B_S0zR8KcJ7_1;
	wire w_dff_B_UBVTSTPL7_1;
	wire w_dff_B_8YY9fMqH0_1;
	wire w_dff_B_0oEdJGk36_1;
	wire w_dff_B_o4qTf8jB5_1;
	wire w_dff_B_MPDSEuom9_1;
	wire w_dff_B_c8ylioBm9_1;
	wire w_dff_B_nWFNcPuy9_1;
	wire w_dff_B_0SwTFmC67_1;
	wire w_dff_B_CeOU4EFo6_1;
	wire w_dff_B_UY8LQKXX4_1;
	wire w_dff_B_fno0KeT45_1;
	wire w_dff_B_JlRKt4Hh9_1;
	wire w_dff_B_v3VyVP3u6_1;
	wire w_dff_B_0VnddscN1_1;
	wire w_dff_B_YQVrJRo68_1;
	wire w_dff_B_MQ8eRaQ16_1;
	wire w_dff_B_Q2hFncA24_1;
	wire w_dff_B_90HziY8o0_1;
	wire w_dff_B_R7LC8kK87_1;
	wire w_dff_B_CTOAbFb57_1;
	wire w_dff_B_2DMqRswL7_0;
	wire w_dff_B_xBuCHRR42_0;
	wire w_dff_B_XKbh560A8_0;
	wire w_dff_B_lKBUYmLM9_0;
	wire w_dff_B_ScFiBwxj0_0;
	wire w_dff_B_YcTdU1gp2_0;
	wire w_dff_B_GJAjsNRd6_0;
	wire w_dff_B_MfxeiVbI4_0;
	wire w_dff_B_QcEt8eNG0_0;
	wire w_dff_B_7x8H3DV25_0;
	wire w_dff_B_aekMSfWk4_0;
	wire w_dff_B_KXjnSbXn0_0;
	wire w_dff_B_J1nJZVwh3_0;
	wire w_dff_B_qHR0xegx2_0;
	wire w_dff_B_bOy7XOuS1_0;
	wire w_dff_B_ypOF11ny7_0;
	wire w_dff_B_mxDxIay68_0;
	wire w_dff_B_OOC2jVv87_0;
	wire w_dff_B_Cy9UViWe1_0;
	wire w_dff_B_MrbGNQYL7_0;
	wire w_dff_B_BWYUbXs32_0;
	wire w_dff_B_cGcQ3dir2_0;
	wire w_dff_B_IjwtMq1Q2_0;
	wire w_dff_B_YrkQIZLi8_0;
	wire w_dff_B_83JO0qDw7_0;
	wire w_dff_B_u4zdLjIr7_0;
	wire w_dff_B_OvoTV3iT5_0;
	wire w_dff_B_AKxmYToU0_0;
	wire w_dff_B_rB8X50qJ6_0;
	wire w_dff_B_Xxzgxo4c9_0;
	wire w_dff_B_SxquOrW65_0;
	wire w_dff_B_KZGxgImK6_0;
	wire w_dff_B_PJp2lxaC5_0;
	wire w_dff_B_ChAtkDs68_0;
	wire w_dff_B_nZxjo0XW2_0;
	wire w_dff_B_5nBc7xwK0_0;
	wire w_dff_B_Xv7jY3EZ5_0;
	wire w_dff_B_THzs32C03_0;
	wire w_dff_B_I7MFPJDM5_0;
	wire w_dff_B_2Cn5U2F45_0;
	wire w_dff_B_lLJQocVo0_0;
	wire w_dff_B_H3HluzHI1_0;
	wire w_dff_B_Oe8ll1Ws8_0;
	wire w_dff_B_FnJBjWar1_0;
	wire w_dff_B_G0qZVe1L0_0;
	wire w_dff_B_bZvfMu5U8_0;
	wire w_dff_B_VFHLz0Y14_0;
	wire w_dff_B_cMimULRD4_0;
	wire w_dff_B_jtKpkOcZ6_0;
	wire w_dff_B_IztNoIMf2_0;
	wire w_dff_B_K3mqoUfs1_0;
	wire w_dff_B_fsw5iKBs5_0;
	wire w_dff_B_MZQyXlyG3_0;
	wire w_dff_B_NlwdAv251_0;
	wire w_dff_B_4qZsYSHs0_0;
	wire w_dff_B_lhi9bC4H7_0;
	wire w_dff_B_VD3Wc7S56_0;
	wire w_dff_B_JVLbNvhS5_0;
	wire w_dff_B_I1RSLtRl2_0;
	wire w_dff_B_jiebWjNd1_0;
	wire w_dff_B_ZjkdADfx0_0;
	wire w_dff_B_FfLSB3rV3_0;
	wire w_dff_B_JUguTPI86_0;
	wire w_dff_B_PcIGDrxO4_0;
	wire w_dff_B_BDNe8ZEZ7_0;
	wire w_dff_B_KH5FZZGx9_0;
	wire w_dff_B_5DURdh370_0;
	wire w_dff_B_q4K6CRfJ5_0;
	wire w_dff_B_vXlbygkA6_0;
	wire w_dff_B_VGTIDXsV5_0;
	wire w_dff_B_XXOZJK8q0_0;
	wire w_dff_B_aaQvUOy22_0;
	wire w_dff_B_WpE5i4M96_0;
	wire w_dff_B_8qzNuaiB0_0;
	wire w_dff_B_zJ6k3pij6_0;
	wire w_dff_B_tNMA2gKW9_0;
	wire w_dff_B_UcgRjmm15_0;
	wire w_dff_B_FdCSyEd02_0;
	wire w_dff_B_AXYDZMNB2_0;
	wire w_dff_B_z1wmerGy6_0;
	wire w_dff_B_MdDCbMdU2_0;
	wire w_dff_B_qpSaXMca4_0;
	wire w_dff_B_FIpSm2XP9_0;
	wire w_dff_B_BAYi9v7u5_0;
	wire w_dff_B_Uz99iBGr7_0;
	wire w_dff_B_SaRDTlUT9_0;
	wire w_dff_B_aKphVdIy6_0;
	wire w_dff_B_VGjpTU1u9_0;
	wire w_dff_B_E2S8nRC23_0;
	wire w_dff_B_x0fgemQS2_0;
	wire w_dff_B_fi93cS7e7_0;
	wire w_dff_B_X6rYgYGA1_0;
	wire w_dff_B_LFeU1zzp4_0;
	wire w_dff_B_diSNUr6c2_0;
	wire w_dff_B_k0Svme9a1_0;
	wire w_dff_B_Gzgy1Qhg2_0;
	wire w_dff_B_G7Zm8O1g3_0;
	wire w_dff_B_iFZ3HDaO6_0;
	wire w_dff_B_pkVu7UHh8_0;
	wire w_dff_B_gJWoYztq2_0;
	wire w_dff_B_QphMgtJX7_0;
	wire w_dff_B_MNe3cJhP9_0;
	wire w_dff_B_Kj5AR5fJ7_1;
	wire w_dff_B_oovlYFa64_1;
	wire w_dff_B_Oq3sHPJg2_1;
	wire w_dff_B_xjPrILrz4_1;
	wire w_dff_B_F4lLoHk67_1;
	wire w_dff_B_7PrOpdYl8_1;
	wire w_dff_B_wHjuVeUC1_1;
	wire w_dff_B_bRPaR6oL3_1;
	wire w_dff_B_CdFqOPkU0_1;
	wire w_dff_B_Q6drcGUE6_1;
	wire w_dff_B_JWBxPnSI7_1;
	wire w_dff_B_s9wLR4hg0_1;
	wire w_dff_B_CTnX0Qhc5_1;
	wire w_dff_B_8iFRSUQ14_1;
	wire w_dff_B_0gBtGdap6_1;
	wire w_dff_B_15GUVvqO8_1;
	wire w_dff_B_zPMx39Ge7_1;
	wire w_dff_B_yC50Oo7z4_1;
	wire w_dff_B_i2gZfiC96_1;
	wire w_dff_B_W1GlwIdV2_1;
	wire w_dff_B_GqDpNLGt6_1;
	wire w_dff_B_6jh7DCiL5_1;
	wire w_dff_B_oX0dvEqh0_1;
	wire w_dff_B_Ox9u8pFD1_1;
	wire w_dff_B_0XUaaG3w6_1;
	wire w_dff_B_QbeXYslI5_1;
	wire w_dff_B_hdejZx0q3_1;
	wire w_dff_B_NsNeJRRP7_1;
	wire w_dff_B_rCFS9CA73_1;
	wire w_dff_B_UG2dEszc7_1;
	wire w_dff_B_4ekLntUr4_1;
	wire w_dff_B_KSbivQYk5_1;
	wire w_dff_B_jwm2cIUf8_1;
	wire w_dff_B_wDMddMnV5_1;
	wire w_dff_B_cTG46KWu8_1;
	wire w_dff_B_2B57DeYB5_1;
	wire w_dff_B_LpvxXFYX9_1;
	wire w_dff_B_w4YPEJlc9_1;
	wire w_dff_B_gKUC1bO50_1;
	wire w_dff_B_7nXJ67Dt8_1;
	wire w_dff_B_lfdK1lJW1_1;
	wire w_dff_B_7L3Oi4Vy0_1;
	wire w_dff_B_PBi1OoMT8_1;
	wire w_dff_B_9auMD5uR7_1;
	wire w_dff_B_eqS0iseN6_1;
	wire w_dff_B_Cet8uBUu6_1;
	wire w_dff_B_k0F8m3NB9_1;
	wire w_dff_B_SZQUkxMM3_1;
	wire w_dff_B_v36G6yS04_1;
	wire w_dff_B_BkwC78Od6_1;
	wire w_dff_B_uwb9k4xF1_1;
	wire w_dff_B_nmsBbPLB4_1;
	wire w_dff_B_K8EOOJ1M7_1;
	wire w_dff_B_5mIDOJEl0_1;
	wire w_dff_B_ynEJA2Cc8_1;
	wire w_dff_B_fERPU5X67_1;
	wire w_dff_B_25EwPB4s3_1;
	wire w_dff_B_9AC2eQed8_1;
	wire w_dff_B_wMCjXOI78_1;
	wire w_dff_B_M7JlE5Aj8_1;
	wire w_dff_B_vms5oa6r8_1;
	wire w_dff_B_xNZqeWOU9_1;
	wire w_dff_B_TBbIDfG28_1;
	wire w_dff_B_nSaVU8LB8_1;
	wire w_dff_B_Li1VsOmH7_1;
	wire w_dff_B_zfahlay29_1;
	wire w_dff_B_dUFONw517_1;
	wire w_dff_B_xF30TW5R7_1;
	wire w_dff_B_XTErd2bd2_1;
	wire w_dff_B_SKDCRRov5_1;
	wire w_dff_B_EufDlfqr8_1;
	wire w_dff_B_yc8vxl173_1;
	wire w_dff_B_S2LNM6L52_1;
	wire w_dff_B_TXNrvu3H2_1;
	wire w_dff_B_wVkADsaW7_1;
	wire w_dff_B_7pjHbMAI4_1;
	wire w_dff_B_CZyv6MJn5_1;
	wire w_dff_B_RjzaxENB5_1;
	wire w_dff_B_ws037e9S8_1;
	wire w_dff_B_1RiDqpM92_1;
	wire w_dff_B_7iulf4eM9_1;
	wire w_dff_B_AmMmxHSs5_1;
	wire w_dff_B_L4mSRr4i5_1;
	wire w_dff_B_GDBqg1AN6_1;
	wire w_dff_B_R12BfaXI8_1;
	wire w_dff_B_IuPAEgwk6_1;
	wire w_dff_B_fcZduaqd0_1;
	wire w_dff_B_VoNjxuvq5_1;
	wire w_dff_B_wktnuJFL4_1;
	wire w_dff_B_12byotXl6_1;
	wire w_dff_B_aaVNcO7N2_1;
	wire w_dff_B_aZasClLY4_1;
	wire w_dff_B_qn2brB9g5_1;
	wire w_dff_B_SiLJdpvG4_1;
	wire w_dff_B_4VtBdByz4_1;
	wire w_dff_B_hUe7bFZi0_1;
	wire w_dff_B_Iw8yfBaD8_1;
	wire w_dff_B_D9pND7lJ6_1;
	wire w_dff_B_RfhM5a1Q5_1;
	wire w_dff_B_b3qpPrCX5_1;
	wire w_dff_B_eOrMuw528_1;
	wire w_dff_B_PQRirv0m1_0;
	wire w_dff_B_D9gpv3kI4_0;
	wire w_dff_B_4K39FXIG9_0;
	wire w_dff_B_8PdTeILF8_0;
	wire w_dff_B_2T2924mg3_0;
	wire w_dff_B_v4SQFyul6_0;
	wire w_dff_B_ri0HYp239_0;
	wire w_dff_B_1ypkeiBu2_0;
	wire w_dff_B_y9nRsGxj9_0;
	wire w_dff_B_TTfgeIOM0_0;
	wire w_dff_B_aHfEl3WP9_0;
	wire w_dff_B_BYKjJXzo3_0;
	wire w_dff_B_gCklSXy41_0;
	wire w_dff_B_7IFKvv5m7_0;
	wire w_dff_B_i8Xq67pF2_0;
	wire w_dff_B_FfZUezRD1_0;
	wire w_dff_B_ecgCzsY40_0;
	wire w_dff_B_rTBFtG2P6_0;
	wire w_dff_B_XDrDrEvz3_0;
	wire w_dff_B_ewOkrIJn8_0;
	wire w_dff_B_nn3scauF5_0;
	wire w_dff_B_dcrNNsXE3_0;
	wire w_dff_B_xVkHm4c43_0;
	wire w_dff_B_m4vONICa3_0;
	wire w_dff_B_lnc1Snmr9_0;
	wire w_dff_B_cw030unO2_0;
	wire w_dff_B_TEO5YD8Z8_0;
	wire w_dff_B_LQrZYVFJ6_0;
	wire w_dff_B_DYhN7bMT4_0;
	wire w_dff_B_DoVj4msS1_0;
	wire w_dff_B_AN4TmMtZ1_0;
	wire w_dff_B_r1HvdoVy1_0;
	wire w_dff_B_v8ivtiXS6_0;
	wire w_dff_B_Ng9qgkXr5_0;
	wire w_dff_B_mCWpCiQC9_0;
	wire w_dff_B_TVLkAODu4_0;
	wire w_dff_B_gssSvAKg1_0;
	wire w_dff_B_Nt8AkM2W0_0;
	wire w_dff_B_uW15OETl6_0;
	wire w_dff_B_OSrkWgmF6_0;
	wire w_dff_B_5WZOjuU90_0;
	wire w_dff_B_zRNUK3wv8_0;
	wire w_dff_B_rx6J8DIR6_0;
	wire w_dff_B_T5e4P5jh1_0;
	wire w_dff_B_Tw7YyZQy8_0;
	wire w_dff_B_qzOjTNJG6_0;
	wire w_dff_B_cIeubwr68_0;
	wire w_dff_B_dOMyglfL4_0;
	wire w_dff_B_r2oqDg6g1_0;
	wire w_dff_B_DP5UyGLi3_0;
	wire w_dff_B_GOXbqGGt6_0;
	wire w_dff_B_qUf7scos5_0;
	wire w_dff_B_hXwger6Q0_0;
	wire w_dff_B_qaG96RCx0_0;
	wire w_dff_B_jR6pJF6b9_0;
	wire w_dff_B_hGWJW1Oi3_0;
	wire w_dff_B_m69YFwVh8_0;
	wire w_dff_B_XP178ACT1_0;
	wire w_dff_B_Tyz7FRDj5_0;
	wire w_dff_B_Kvp7cwzZ7_0;
	wire w_dff_B_WmtFT1UX8_0;
	wire w_dff_B_WaZiaEi05_0;
	wire w_dff_B_YcrveNHU9_0;
	wire w_dff_B_XzUjWw8I8_0;
	wire w_dff_B_ro1gLVvR6_0;
	wire w_dff_B_4x0fcnX07_0;
	wire w_dff_B_ALyepbeq7_0;
	wire w_dff_B_f6iUujuk5_0;
	wire w_dff_B_IB6jH9PE8_0;
	wire w_dff_B_g88kN3uI6_0;
	wire w_dff_B_D4X58SKJ5_0;
	wire w_dff_B_4nhufPn46_0;
	wire w_dff_B_ELMaxXhd1_0;
	wire w_dff_B_5GHwduaf2_0;
	wire w_dff_B_hycexgJs7_0;
	wire w_dff_B_9D3h1bEM0_0;
	wire w_dff_B_2w9i8F3i2_0;
	wire w_dff_B_eqgPPYbX5_0;
	wire w_dff_B_G5rtZoew6_0;
	wire w_dff_B_v9otEqz79_0;
	wire w_dff_B_Fe5Cztr34_0;
	wire w_dff_B_HluWOPtu2_0;
	wire w_dff_B_4llKQOpS1_0;
	wire w_dff_B_Aog8pcXj5_0;
	wire w_dff_B_hSYLk0sV3_0;
	wire w_dff_B_yRRRiyKJ6_0;
	wire w_dff_B_95jaZ1ps3_0;
	wire w_dff_B_vU336DFM7_0;
	wire w_dff_B_HyPNRr7b0_0;
	wire w_dff_B_aK28yDJq0_0;
	wire w_dff_B_RNu8fyVC8_0;
	wire w_dff_B_wzn4mPF53_0;
	wire w_dff_B_bFsrc20v8_0;
	wire w_dff_B_7jmY5U6d3_0;
	wire w_dff_B_w04qloms2_0;
	wire w_dff_B_Hdq9eNO36_0;
	wire w_dff_B_4tDfSGdR2_0;
	wire w_dff_B_SX4kGZlS9_0;
	wire w_dff_B_wm6uFC186_0;
	wire w_dff_B_jse6aP2y1_0;
	wire w_dff_B_WKYHnQ064_0;
	wire w_dff_B_dW3bOQsl4_1;
	wire w_dff_B_EAtwghzA5_1;
	wire w_dff_B_bZUiXPwS2_1;
	wire w_dff_B_tqVeCLjJ6_1;
	wire w_dff_B_TZVevdMK9_1;
	wire w_dff_B_JSUQAoxZ4_1;
	wire w_dff_B_vzk5YVgY7_1;
	wire w_dff_B_ahVDdP2N6_1;
	wire w_dff_B_ZxNxXE353_1;
	wire w_dff_B_cd5oMpdK5_1;
	wire w_dff_B_eVM8NMRf2_1;
	wire w_dff_B_ZhpnEFfF8_1;
	wire w_dff_B_Ft4cEAzk5_1;
	wire w_dff_B_dHnhehqL8_1;
	wire w_dff_B_0hhvlaJU9_1;
	wire w_dff_B_Z2f1xnDL8_1;
	wire w_dff_B_ACiDnWhG9_1;
	wire w_dff_B_H9atbfUk1_1;
	wire w_dff_B_z6reGHio0_1;
	wire w_dff_B_8prjGHfW0_1;
	wire w_dff_B_6PZ9zAgl7_1;
	wire w_dff_B_404R34Wx4_1;
	wire w_dff_B_QFVLQk999_1;
	wire w_dff_B_ZdvJztze0_1;
	wire w_dff_B_jtUU8lLt4_1;
	wire w_dff_B_ErfJELrv8_1;
	wire w_dff_B_SfgdcvMN5_1;
	wire w_dff_B_y6mhtZWH9_1;
	wire w_dff_B_SxZQYWiU0_1;
	wire w_dff_B_Ym66mhjs3_1;
	wire w_dff_B_zk0lrBTR9_1;
	wire w_dff_B_sBKj8tvH3_1;
	wire w_dff_B_9RGFGaUs8_1;
	wire w_dff_B_b8F8wylu8_1;
	wire w_dff_B_FoGxaiXO7_1;
	wire w_dff_B_htFtFf5k4_1;
	wire w_dff_B_efNeOYOv9_1;
	wire w_dff_B_nb21rX101_1;
	wire w_dff_B_cyE9GT2i1_1;
	wire w_dff_B_H3vbTa5N0_1;
	wire w_dff_B_0K4W2rfU6_1;
	wire w_dff_B_fU3HWTrg4_1;
	wire w_dff_B_CEJbSzhb7_1;
	wire w_dff_B_Ha899IwM9_1;
	wire w_dff_B_q3iHuL7x8_1;
	wire w_dff_B_rWaVp7W00_1;
	wire w_dff_B_V6nJ2JND0_1;
	wire w_dff_B_tKpXAavf9_1;
	wire w_dff_B_W9iXaONO1_1;
	wire w_dff_B_dhxVqzlD7_1;
	wire w_dff_B_U7TsXFN70_1;
	wire w_dff_B_41vyKhgg0_1;
	wire w_dff_B_CGViD9Ra2_1;
	wire w_dff_B_VlY5E9vk3_1;
	wire w_dff_B_PfXaZAgN8_1;
	wire w_dff_B_RHPfq9Ac8_1;
	wire w_dff_B_PM0i3fPu5_1;
	wire w_dff_B_qwWAUPHb8_1;
	wire w_dff_B_6ndAXiJ42_1;
	wire w_dff_B_P4W8IZrJ2_1;
	wire w_dff_B_rtr0nblm8_1;
	wire w_dff_B_48IR0VUc0_1;
	wire w_dff_B_Cl5xRC565_1;
	wire w_dff_B_tm8WBy4I7_1;
	wire w_dff_B_yFhqCxz27_1;
	wire w_dff_B_Tlc9wAFJ4_1;
	wire w_dff_B_Sc1HFL605_1;
	wire w_dff_B_QzYujono6_1;
	wire w_dff_B_ST20qWtV2_1;
	wire w_dff_B_IMsnHKjp4_1;
	wire w_dff_B_eEqRptMH7_1;
	wire w_dff_B_tEtvD5pC8_1;
	wire w_dff_B_PkbUtv1R1_1;
	wire w_dff_B_XQiqryRZ3_1;
	wire w_dff_B_u1hQWf5a5_1;
	wire w_dff_B_QPZUVCc46_1;
	wire w_dff_B_VcIic6js6_1;
	wire w_dff_B_ZVojjKw26_1;
	wire w_dff_B_ZM3RHWZj3_1;
	wire w_dff_B_nMZBmZ6Y5_1;
	wire w_dff_B_KxGC3tHv5_1;
	wire w_dff_B_46pT0eQ89_1;
	wire w_dff_B_PQ9oIgaA7_1;
	wire w_dff_B_Z0StsYyh3_1;
	wire w_dff_B_iZeFzGdY0_1;
	wire w_dff_B_eEUI45IG3_1;
	wire w_dff_B_j1mj19K26_1;
	wire w_dff_B_NIH6EfS74_1;
	wire w_dff_B_iwPjKlG56_1;
	wire w_dff_B_8mtLIjRB2_1;
	wire w_dff_B_aWVqOKkb0_1;
	wire w_dff_B_U5fTCsZj0_1;
	wire w_dff_B_1CDbxVMk3_1;
	wire w_dff_B_OhiKHpSY6_1;
	wire w_dff_B_pPjbgOal2_1;
	wire w_dff_B_9L9tzgWz6_1;
	wire w_dff_B_bHi0BR043_1;
	wire w_dff_B_5Nk4raz90_1;
	wire w_dff_B_JYPc6Jnl2_1;
	wire w_dff_B_ihOKXM3G5_1;
	wire w_dff_B_eEkl9s2m0_0;
	wire w_dff_B_D8KUBLF05_0;
	wire w_dff_B_qf2xbpia8_0;
	wire w_dff_B_cF2Sw4nS1_0;
	wire w_dff_B_F8K1U4a32_0;
	wire w_dff_B_gzVC7ztD2_0;
	wire w_dff_B_kfUrLfsQ6_0;
	wire w_dff_B_dK0S79aT7_0;
	wire w_dff_B_x0nMv34b8_0;
	wire w_dff_B_eyLtVXlI7_0;
	wire w_dff_B_X5hgcZze5_0;
	wire w_dff_B_Pz5HTgqD6_0;
	wire w_dff_B_y4rYCSiz6_0;
	wire w_dff_B_6ThmlYtL4_0;
	wire w_dff_B_Qt5IzyyR1_0;
	wire w_dff_B_ObpYJLW88_0;
	wire w_dff_B_bHDtyw2h2_0;
	wire w_dff_B_Rq0JrPuX7_0;
	wire w_dff_B_F34YsqpI4_0;
	wire w_dff_B_eDZTykKZ1_0;
	wire w_dff_B_x5VNB92I5_0;
	wire w_dff_B_aI8VEOIL6_0;
	wire w_dff_B_etFAJqn31_0;
	wire w_dff_B_MHIml8f18_0;
	wire w_dff_B_1atySNUl8_0;
	wire w_dff_B_FdquoYvk6_0;
	wire w_dff_B_CFKLh3J16_0;
	wire w_dff_B_yENi3WCZ7_0;
	wire w_dff_B_279KTDcr6_0;
	wire w_dff_B_ovzb43mE2_0;
	wire w_dff_B_KWKTiTHN0_0;
	wire w_dff_B_9z2B29rq6_0;
	wire w_dff_B_evTDnltg1_0;
	wire w_dff_B_rTLjHJzu6_0;
	wire w_dff_B_zlJc4Iql7_0;
	wire w_dff_B_BRXTv2Ar3_0;
	wire w_dff_B_8ew50BET9_0;
	wire w_dff_B_Jvy36XlD1_0;
	wire w_dff_B_Gzfj7Rtr1_0;
	wire w_dff_B_L9JCj7Nh2_0;
	wire w_dff_B_DHosqy593_0;
	wire w_dff_B_4Vx0avMy9_0;
	wire w_dff_B_9JBOmamy5_0;
	wire w_dff_B_94Vg3t2Y5_0;
	wire w_dff_B_N0GTgjBi0_0;
	wire w_dff_B_NAw1NFwm6_0;
	wire w_dff_B_SV7uZX0U3_0;
	wire w_dff_B_l3YsVBH02_0;
	wire w_dff_B_r5fRi3ip8_0;
	wire w_dff_B_ntCgpe8A0_0;
	wire w_dff_B_35GHKOE14_0;
	wire w_dff_B_FQSkhLyP4_0;
	wire w_dff_B_IvlD4qZH5_0;
	wire w_dff_B_SL43gV0Q9_0;
	wire w_dff_B_afRyoNGk8_0;
	wire w_dff_B_88uefvSS1_0;
	wire w_dff_B_kUwJ55Pl8_0;
	wire w_dff_B_jyvSWpbW0_0;
	wire w_dff_B_MHLF0uRC8_0;
	wire w_dff_B_mVgsqD6c4_0;
	wire w_dff_B_SClotsqa5_0;
	wire w_dff_B_LfPBmi6M8_0;
	wire w_dff_B_SJrdyF1v3_0;
	wire w_dff_B_X9qmn73p7_0;
	wire w_dff_B_9jzDUsxY1_0;
	wire w_dff_B_GRKnsCBI3_0;
	wire w_dff_B_caQ1HtKN7_0;
	wire w_dff_B_sWDZ9yAP0_0;
	wire w_dff_B_FxuBYA3C1_0;
	wire w_dff_B_AMLNUDZa6_0;
	wire w_dff_B_gL9ovFQ70_0;
	wire w_dff_B_v3OMlvve5_0;
	wire w_dff_B_HTPqckhM9_0;
	wire w_dff_B_9mpvb3V42_0;
	wire w_dff_B_uhuyayo28_0;
	wire w_dff_B_prU3UkQf5_0;
	wire w_dff_B_fkAOM1JZ7_0;
	wire w_dff_B_n9KTjp973_0;
	wire w_dff_B_s6T8f5YH9_0;
	wire w_dff_B_j09wXN7a2_0;
	wire w_dff_B_vJFA0Str3_0;
	wire w_dff_B_MNoNaIff9_0;
	wire w_dff_B_sdvHJx4Z4_0;
	wire w_dff_B_DIOzZIet3_0;
	wire w_dff_B_Ly8V1W0a0_0;
	wire w_dff_B_K1JjLZHY3_0;
	wire w_dff_B_z2W0T16R9_0;
	wire w_dff_B_rAvTOp0k3_0;
	wire w_dff_B_kHJmpJSC1_0;
	wire w_dff_B_tdDJgPSW1_0;
	wire w_dff_B_VVqaybmK0_0;
	wire w_dff_B_hHQUy4MR1_0;
	wire w_dff_B_5SgonsWr9_0;
	wire w_dff_B_ut7QM3Hu0_0;
	wire w_dff_B_VHq0bp8e0_0;
	wire w_dff_B_ACyBYY7T7_0;
	wire w_dff_B_YtryxROZ1_0;
	wire w_dff_B_1a6uerT96_0;
	wire w_dff_B_dYjiT6bc3_0;
	wire w_dff_B_ZBeU3nCK4_0;
	wire w_dff_B_n82feeXJ6_1;
	wire w_dff_B_WkAQ7u6W2_1;
	wire w_dff_B_Gy6kPcyJ2_1;
	wire w_dff_B_0wgGlcsX2_1;
	wire w_dff_B_agtoXMUa0_1;
	wire w_dff_B_7l8pwWSl6_1;
	wire w_dff_B_tVJkpn0z3_1;
	wire w_dff_B_MfLCiWjv1_1;
	wire w_dff_B_6B6ifIgf0_1;
	wire w_dff_B_6Vvsb01V8_1;
	wire w_dff_B_JFGj1o086_1;
	wire w_dff_B_4kEhO6654_1;
	wire w_dff_B_gaFn8EE36_1;
	wire w_dff_B_js56byEH9_1;
	wire w_dff_B_7FPHmqli1_1;
	wire w_dff_B_bNkFueRe3_1;
	wire w_dff_B_7tcyyuyz4_1;
	wire w_dff_B_F14aY1DM8_1;
	wire w_dff_B_vNrMpOOE0_1;
	wire w_dff_B_U6VQecYl7_1;
	wire w_dff_B_kVVFQFnb7_1;
	wire w_dff_B_TfQjYiCO0_1;
	wire w_dff_B_FipZUJmv2_1;
	wire w_dff_B_Ut6LkS6c3_1;
	wire w_dff_B_UiYvUax80_1;
	wire w_dff_B_K0Lk56Wa1_1;
	wire w_dff_B_Vqz7au1b1_1;
	wire w_dff_B_C6rk0dxg7_1;
	wire w_dff_B_t9OXnGY12_1;
	wire w_dff_B_0efPE6rr3_1;
	wire w_dff_B_HAJIT6Na0_1;
	wire w_dff_B_jcnzE5Jb5_1;
	wire w_dff_B_h02VGJpv7_1;
	wire w_dff_B_rMtvu2vC1_1;
	wire w_dff_B_t1jv47dd1_1;
	wire w_dff_B_X7HolBmJ8_1;
	wire w_dff_B_DQgBa13G7_1;
	wire w_dff_B_g5DcuphP8_1;
	wire w_dff_B_cwx6rjzh1_1;
	wire w_dff_B_sAG6e7xv6_1;
	wire w_dff_B_n8VY4oYC7_1;
	wire w_dff_B_JnI5wO649_1;
	wire w_dff_B_97GSGcyp0_1;
	wire w_dff_B_VH4azXFr3_1;
	wire w_dff_B_zasPMfwE5_1;
	wire w_dff_B_6Y1kiCmQ0_1;
	wire w_dff_B_Uyk3Gpn20_1;
	wire w_dff_B_DyElRSxN3_1;
	wire w_dff_B_2yGZeXi54_1;
	wire w_dff_B_615Gw5Dn4_1;
	wire w_dff_B_YY4UgXBP1_1;
	wire w_dff_B_geC9abhG8_1;
	wire w_dff_B_wJW0CYU81_1;
	wire w_dff_B_Hdfepvd84_1;
	wire w_dff_B_pRnUMcW69_1;
	wire w_dff_B_NzppTr7Z4_1;
	wire w_dff_B_6LFlVRea8_1;
	wire w_dff_B_eBTKs3XB0_1;
	wire w_dff_B_oGBfP9N66_1;
	wire w_dff_B_O5hCadVz8_1;
	wire w_dff_B_2Kb5B5Pe9_1;
	wire w_dff_B_vbs6i2S92_1;
	wire w_dff_B_Ci4Wnzv17_1;
	wire w_dff_B_Yxo4r10Z5_1;
	wire w_dff_B_F5hhH1ky1_1;
	wire w_dff_B_ZrPO1EYw8_1;
	wire w_dff_B_NHXs0VmM5_1;
	wire w_dff_B_pJnEtqX11_1;
	wire w_dff_B_JAiFItIv1_1;
	wire w_dff_B_aWURpxMI8_1;
	wire w_dff_B_RD3jpQJC6_1;
	wire w_dff_B_fjmJSJfd4_1;
	wire w_dff_B_WSqCwYOX8_1;
	wire w_dff_B_3IJIS5TI0_1;
	wire w_dff_B_KkQQOTJO7_1;
	wire w_dff_B_yRMPGGna3_1;
	wire w_dff_B_1b4SG3UD4_1;
	wire w_dff_B_rjPrTpep2_1;
	wire w_dff_B_v8vo6aph6_1;
	wire w_dff_B_GPP20TpI9_1;
	wire w_dff_B_DxnqTG731_1;
	wire w_dff_B_f4A6OvnA9_1;
	wire w_dff_B_sXFj5RV76_1;
	wire w_dff_B_t6n5teLA0_1;
	wire w_dff_B_eGtIiAFY6_1;
	wire w_dff_B_N1GsdJ2a5_1;
	wire w_dff_B_pkTK782F8_1;
	wire w_dff_B_HmTlhb8b1_1;
	wire w_dff_B_gfNzXfd36_1;
	wire w_dff_B_ykuba2Ed6_1;
	wire w_dff_B_83jJYclD3_1;
	wire w_dff_B_R4vn3LvQ9_1;
	wire w_dff_B_KK540xpY0_1;
	wire w_dff_B_IlqIn0Sw2_1;
	wire w_dff_B_q4NvRVS12_1;
	wire w_dff_B_24Tvryrg2_1;
	wire w_dff_B_6VIr25WK5_1;
	wire w_dff_B_VbfHAiNn1_1;
	wire w_dff_B_miF1RlLv4_1;
	wire w_dff_B_3nrQhyw92_0;
	wire w_dff_B_CbbIn7De4_0;
	wire w_dff_B_TNhXpKTA8_0;
	wire w_dff_B_XBKPienL3_0;
	wire w_dff_B_J4QZxdaB8_0;
	wire w_dff_B_VZKRyolt2_0;
	wire w_dff_B_Gq4cEV8O4_0;
	wire w_dff_B_z5bhuvm83_0;
	wire w_dff_B_Cfaw5fL02_0;
	wire w_dff_B_lLSfw8h66_0;
	wire w_dff_B_ZPjS357q8_0;
	wire w_dff_B_6cCCoO4T4_0;
	wire w_dff_B_51NaMtTy6_0;
	wire w_dff_B_nBtYDfgE3_0;
	wire w_dff_B_lrnpdaoP4_0;
	wire w_dff_B_PsZmjjBa3_0;
	wire w_dff_B_YjOEHnX96_0;
	wire w_dff_B_zjCVIRYL7_0;
	wire w_dff_B_LBY4wlAw6_0;
	wire w_dff_B_Zh5f54wP8_0;
	wire w_dff_B_evLOa2o75_0;
	wire w_dff_B_UJHFRTpn2_0;
	wire w_dff_B_DEjALPo85_0;
	wire w_dff_B_P4sEBclQ3_0;
	wire w_dff_B_LBIBHDpo6_0;
	wire w_dff_B_Z8GiTpec7_0;
	wire w_dff_B_4vyCtkBr9_0;
	wire w_dff_B_RVhu7ODk2_0;
	wire w_dff_B_NxIVddl43_0;
	wire w_dff_B_7d8uokgC2_0;
	wire w_dff_B_13CNFcAF2_0;
	wire w_dff_B_PK67j5m66_0;
	wire w_dff_B_vXvQQ8JZ8_0;
	wire w_dff_B_fEHuOur00_0;
	wire w_dff_B_pYGG8UsA7_0;
	wire w_dff_B_lJW7bXCv6_0;
	wire w_dff_B_AMZD781e0_0;
	wire w_dff_B_AzafLKOk8_0;
	wire w_dff_B_XiEVUsl41_0;
	wire w_dff_B_eKyToK7j1_0;
	wire w_dff_B_VgmczsXf0_0;
	wire w_dff_B_fgcGeT7F4_0;
	wire w_dff_B_yGCbEa8h2_0;
	wire w_dff_B_VGknEvuL7_0;
	wire w_dff_B_wHcIpB151_0;
	wire w_dff_B_BciolMIY8_0;
	wire w_dff_B_MmtSn4mq0_0;
	wire w_dff_B_dPdT549G8_0;
	wire w_dff_B_GxU8k5yj6_0;
	wire w_dff_B_aAA4G1Hu8_0;
	wire w_dff_B_z08MuNHr2_0;
	wire w_dff_B_VrgYqoUE8_0;
	wire w_dff_B_PppM4nIV6_0;
	wire w_dff_B_bWRkCA5q7_0;
	wire w_dff_B_Cdr4sT0g5_0;
	wire w_dff_B_Pktez2lp6_0;
	wire w_dff_B_8blY9eG88_0;
	wire w_dff_B_eXlQ8K6D0_0;
	wire w_dff_B_NaI5Py8a7_0;
	wire w_dff_B_AoIHz6HU1_0;
	wire w_dff_B_7e28TEzI6_0;
	wire w_dff_B_6pzLgnTy5_0;
	wire w_dff_B_RWrg3STi4_0;
	wire w_dff_B_yFNyU4lr3_0;
	wire w_dff_B_G57TeDAz0_0;
	wire w_dff_B_zmQ0upcc8_0;
	wire w_dff_B_2OW9FTIb4_0;
	wire w_dff_B_F8qd2xgs0_0;
	wire w_dff_B_7EkivCwc2_0;
	wire w_dff_B_mI2TrU6G2_0;
	wire w_dff_B_UgSyorgU1_0;
	wire w_dff_B_Ib6ErwfP1_0;
	wire w_dff_B_t8JDe3iy9_0;
	wire w_dff_B_SwrFF9Aw4_0;
	wire w_dff_B_Vzfxnqkl2_0;
	wire w_dff_B_MyO7Scdb6_0;
	wire w_dff_B_RSFQF9bE8_0;
	wire w_dff_B_WTJABp3A8_0;
	wire w_dff_B_ZRJ9Tv5i7_0;
	wire w_dff_B_FzWP0Bfa9_0;
	wire w_dff_B_xsN5xeiE2_0;
	wire w_dff_B_UBkYUe9l1_0;
	wire w_dff_B_cWja660D3_0;
	wire w_dff_B_T6L9ubBb7_0;
	wire w_dff_B_yY9hNZMB2_0;
	wire w_dff_B_KWycYczW1_0;
	wire w_dff_B_IHMLO9jW2_0;
	wire w_dff_B_rI0sIsJW4_0;
	wire w_dff_B_2dm7WGKX0_0;
	wire w_dff_B_1toynP512_0;
	wire w_dff_B_COeXabQJ7_0;
	wire w_dff_B_SfJJgq0q0_0;
	wire w_dff_B_PmwnDScI5_0;
	wire w_dff_B_f6wAjAeX6_0;
	wire w_dff_B_o5qM1l3d5_0;
	wire w_dff_B_HMy8kcEr3_0;
	wire w_dff_B_ZXdUhwdU2_0;
	wire w_dff_B_qEjfMrsJ3_0;
	wire w_dff_B_wOyfHYTt8_0;
	wire w_dff_B_Z5B1ifAp1_1;
	wire w_dff_B_smI5au8k5_1;
	wire w_dff_B_6BILCbsP8_1;
	wire w_dff_B_dKxRMyPF3_1;
	wire w_dff_B_Bfm9nvDd8_1;
	wire w_dff_B_JFlUgZlJ2_1;
	wire w_dff_B_VGVnmGfa2_1;
	wire w_dff_B_mHTX2EBj4_1;
	wire w_dff_B_2kMjsHUf0_1;
	wire w_dff_B_klBU5ysp5_1;
	wire w_dff_B_NyVsTaYp6_1;
	wire w_dff_B_UJoFoob13_1;
	wire w_dff_B_mA1B7HbN8_1;
	wire w_dff_B_Rlwfmm4F2_1;
	wire w_dff_B_UIxNoNV49_1;
	wire w_dff_B_fwXK3dgO4_1;
	wire w_dff_B_X8d1YTXT0_1;
	wire w_dff_B_y4DbhuP14_1;
	wire w_dff_B_7ZzlPaq74_1;
	wire w_dff_B_JUCpOFes5_1;
	wire w_dff_B_sRnnoN4f1_1;
	wire w_dff_B_UQ6ky9QJ5_1;
	wire w_dff_B_Hc39as0V8_1;
	wire w_dff_B_kkQSVCxI2_1;
	wire w_dff_B_tjrJW4Jp7_1;
	wire w_dff_B_6iEMUaG30_1;
	wire w_dff_B_Dicl31VT7_1;
	wire w_dff_B_o9uwlSEE9_1;
	wire w_dff_B_fBunnmMH4_1;
	wire w_dff_B_vSdZt5K19_1;
	wire w_dff_B_oEcHW4UD8_1;
	wire w_dff_B_hBQGymFB7_1;
	wire w_dff_B_YFRf7nCJ4_1;
	wire w_dff_B_UjkGPIGk1_1;
	wire w_dff_B_0L0OPBlx1_1;
	wire w_dff_B_dDq2mjJ57_1;
	wire w_dff_B_a33gikOx4_1;
	wire w_dff_B_cfv2yNw21_1;
	wire w_dff_B_mbMDqcV79_1;
	wire w_dff_B_rsbBSUQk8_1;
	wire w_dff_B_ArvOWERt6_1;
	wire w_dff_B_GKY25DZB1_1;
	wire w_dff_B_P2HXyoyy1_1;
	wire w_dff_B_rFmaUZyg2_1;
	wire w_dff_B_OfaP09Nb3_1;
	wire w_dff_B_5EIl57YG4_1;
	wire w_dff_B_lW5Lng6G3_1;
	wire w_dff_B_nJrWBbhn9_1;
	wire w_dff_B_OlKgHFTO7_1;
	wire w_dff_B_LHGOzpwD8_1;
	wire w_dff_B_6r7IHxOB7_1;
	wire w_dff_B_vyPhRNvO9_1;
	wire w_dff_B_nNk2b9Pr5_1;
	wire w_dff_B_eZ1gYnSV0_1;
	wire w_dff_B_UcLdKzOT7_1;
	wire w_dff_B_PfQFCLM56_1;
	wire w_dff_B_3X21uRNw3_1;
	wire w_dff_B_i7oZEuPT7_1;
	wire w_dff_B_jnun1KzD2_1;
	wire w_dff_B_QDCFAuB92_1;
	wire w_dff_B_R5voHkfq6_1;
	wire w_dff_B_7dJi9ygn3_1;
	wire w_dff_B_XV6BtSFk7_1;
	wire w_dff_B_tCpZB0Im2_1;
	wire w_dff_B_iVbImZAW4_1;
	wire w_dff_B_MyOzqX2M7_1;
	wire w_dff_B_hv7jnx4o7_1;
	wire w_dff_B_btcU6MIV7_1;
	wire w_dff_B_d6zJbC1Z1_1;
	wire w_dff_B_P7aMs2qJ9_1;
	wire w_dff_B_Bd1rbLsN2_1;
	wire w_dff_B_0vveAfYR4_1;
	wire w_dff_B_wQrgJvMG9_1;
	wire w_dff_B_jMEt6kbz1_1;
	wire w_dff_B_7DcZmRHA5_1;
	wire w_dff_B_FyB1FXnj4_1;
	wire w_dff_B_TxpvTaAI6_1;
	wire w_dff_B_EtMdV7Et3_1;
	wire w_dff_B_ddOF38Ih3_1;
	wire w_dff_B_yGYLIp2W9_1;
	wire w_dff_B_TjlEfZXk4_1;
	wire w_dff_B_l8Ja5oxY8_1;
	wire w_dff_B_U2AwKyTz1_1;
	wire w_dff_B_ApzrNSSa7_1;
	wire w_dff_B_kMolEM8f1_1;
	wire w_dff_B_RiZp2iRJ1_1;
	wire w_dff_B_CqAEFC1Z7_1;
	wire w_dff_B_pYDoLRgG2_1;
	wire w_dff_B_YezcYCFo5_1;
	wire w_dff_B_fOm82p1F7_1;
	wire w_dff_B_Wse4aiTd1_1;
	wire w_dff_B_yqELsMRu5_1;
	wire w_dff_B_thnOzZPD3_1;
	wire w_dff_B_0hf5fLIH0_1;
	wire w_dff_B_grgCfZ3C4_1;
	wire w_dff_B_TUo8Ckd70_1;
	wire w_dff_B_8mMDisi62_1;
	wire w_dff_B_sukvz7S18_1;
	wire w_dff_B_rUqvxiH18_0;
	wire w_dff_B_Xldh1oT70_0;
	wire w_dff_B_o2HIcIT42_0;
	wire w_dff_B_6wcPQrus1_0;
	wire w_dff_B_VeBO6M3b3_0;
	wire w_dff_B_H9JAqf418_0;
	wire w_dff_B_Xac74v3o8_0;
	wire w_dff_B_i61dsSQq3_0;
	wire w_dff_B_5g92NNFy2_0;
	wire w_dff_B_HtbQ3uBa8_0;
	wire w_dff_B_P8OExxy25_0;
	wire w_dff_B_fHPKsPlV9_0;
	wire w_dff_B_WeKWfWe80_0;
	wire w_dff_B_LW4ghJrl4_0;
	wire w_dff_B_LhLFQMKr0_0;
	wire w_dff_B_SJQK9jwT8_0;
	wire w_dff_B_M158QfaG4_0;
	wire w_dff_B_pcL1Gjfy1_0;
	wire w_dff_B_kI75E0aa1_0;
	wire w_dff_B_LpKS0x3B7_0;
	wire w_dff_B_uPgbB2Bz0_0;
	wire w_dff_B_Fo9bFWL57_0;
	wire w_dff_B_tvfTDtLb4_0;
	wire w_dff_B_nnFWtXnt4_0;
	wire w_dff_B_HMgYkUtU6_0;
	wire w_dff_B_y9doERtt2_0;
	wire w_dff_B_FAGuU0yQ9_0;
	wire w_dff_B_H5aKfxvI6_0;
	wire w_dff_B_Fvu5ov6C6_0;
	wire w_dff_B_UcH42UBV5_0;
	wire w_dff_B_LB0ACfsO5_0;
	wire w_dff_B_VzTEqsHa6_0;
	wire w_dff_B_Zg4NCMYi9_0;
	wire w_dff_B_AnzSAkka4_0;
	wire w_dff_B_7GdqVjWD1_0;
	wire w_dff_B_sPuPpmIu0_0;
	wire w_dff_B_pXV3OwQB5_0;
	wire w_dff_B_GGwFsP557_0;
	wire w_dff_B_CBJ2Dphc7_0;
	wire w_dff_B_8pPbuVo30_0;
	wire w_dff_B_qNXc3wRs9_0;
	wire w_dff_B_lvk3HfUk8_0;
	wire w_dff_B_uq5ctBI36_0;
	wire w_dff_B_1Zi5DzAv1_0;
	wire w_dff_B_Qd6rnflo3_0;
	wire w_dff_B_itOgf6c80_0;
	wire w_dff_B_l33AUiP30_0;
	wire w_dff_B_FGTJPmTo6_0;
	wire w_dff_B_pTSbL3mH8_0;
	wire w_dff_B_CCqJujbK5_0;
	wire w_dff_B_l6N3iB2r2_0;
	wire w_dff_B_AKznrzuT1_0;
	wire w_dff_B_FhE4lZ2I0_0;
	wire w_dff_B_spDVAovP0_0;
	wire w_dff_B_AUuyQZPs7_0;
	wire w_dff_B_BjrK1yoO2_0;
	wire w_dff_B_oJApgSLa1_0;
	wire w_dff_B_wYkdhPUN9_0;
	wire w_dff_B_HUBeeWJM7_0;
	wire w_dff_B_M9d0kA6r8_0;
	wire w_dff_B_IKCL7hOb2_0;
	wire w_dff_B_yCSblpJ54_0;
	wire w_dff_B_KiYAU9YB4_0;
	wire w_dff_B_DtAXHXqJ7_0;
	wire w_dff_B_WeGVkTtR1_0;
	wire w_dff_B_GR4eUGU35_0;
	wire w_dff_B_9jjULUl33_0;
	wire w_dff_B_LL6Z1eYE5_0;
	wire w_dff_B_pRfGqLQ09_0;
	wire w_dff_B_n1N6rYyn8_0;
	wire w_dff_B_VtPbto6B5_0;
	wire w_dff_B_Kd1WDuCv8_0;
	wire w_dff_B_hWNAZ5To5_0;
	wire w_dff_B_kq8Swrjc6_0;
	wire w_dff_B_ezraewP35_0;
	wire w_dff_B_wOHk7AAH8_0;
	wire w_dff_B_U8kJ5bLc9_0;
	wire w_dff_B_kxCeRf143_0;
	wire w_dff_B_0cRfT15D3_0;
	wire w_dff_B_sBhSsg0t4_0;
	wire w_dff_B_1Fyhinto4_0;
	wire w_dff_B_O72zvYXv9_0;
	wire w_dff_B_nbRar6NA3_0;
	wire w_dff_B_F1EQOuCM8_0;
	wire w_dff_B_oLhzaB2K7_0;
	wire w_dff_B_UzQxTQzl6_0;
	wire w_dff_B_Q4uhzlvz5_0;
	wire w_dff_B_4ghgTtho9_0;
	wire w_dff_B_bPed92S03_0;
	wire w_dff_B_QEs5bxR17_0;
	wire w_dff_B_ClyVqHKy8_0;
	wire w_dff_B_UkR6PPJC2_0;
	wire w_dff_B_AWx6xZS86_0;
	wire w_dff_B_ekSGesoT8_0;
	wire w_dff_B_p6MYarz92_0;
	wire w_dff_B_lsj58b6A4_0;
	wire w_dff_B_MJq8zZki6_0;
	wire w_dff_B_CzElqIeo4_0;
	wire w_dff_B_Dbr4hHKB7_1;
	wire w_dff_B_M1V8pSCe2_1;
	wire w_dff_B_jt412CnA5_1;
	wire w_dff_B_tYMQQef54_1;
	wire w_dff_B_oTXRj5Ij4_1;
	wire w_dff_B_J52uqJQr5_1;
	wire w_dff_B_AdCRbKfF8_1;
	wire w_dff_B_Fh2SNVTx3_1;
	wire w_dff_B_AfDDOqbi3_1;
	wire w_dff_B_KumwjENN5_1;
	wire w_dff_B_ullppxKj1_1;
	wire w_dff_B_AXN01XtF4_1;
	wire w_dff_B_NX2ttHWO1_1;
	wire w_dff_B_06IpgZUI4_1;
	wire w_dff_B_zQ5EMnhY8_1;
	wire w_dff_B_iQFTAae45_1;
	wire w_dff_B_XUbB55pQ4_1;
	wire w_dff_B_fejEvfLA7_1;
	wire w_dff_B_HxlJQza61_1;
	wire w_dff_B_I30PErWL7_1;
	wire w_dff_B_s2I7wNWS1_1;
	wire w_dff_B_2GqcAZlD1_1;
	wire w_dff_B_PPIq027W4_1;
	wire w_dff_B_yHUIvbsh8_1;
	wire w_dff_B_HHagNUqw6_1;
	wire w_dff_B_E88OA8zG6_1;
	wire w_dff_B_0MySkf4y8_1;
	wire w_dff_B_4DcEFcyJ8_1;
	wire w_dff_B_3nZ7x0qX0_1;
	wire w_dff_B_RGNbmbDh7_1;
	wire w_dff_B_ead1Dbqk2_1;
	wire w_dff_B_dtfXQUXA3_1;
	wire w_dff_B_YcKNjoIO3_1;
	wire w_dff_B_k6ckExfr4_1;
	wire w_dff_B_b02joubA6_1;
	wire w_dff_B_lFo2OMaH8_1;
	wire w_dff_B_UcOtnxf13_1;
	wire w_dff_B_6tBjxt1n6_1;
	wire w_dff_B_25EGAsJT6_1;
	wire w_dff_B_NNt2IY2d5_1;
	wire w_dff_B_P5Ut0wK42_1;
	wire w_dff_B_eXW653uy9_1;
	wire w_dff_B_mmHEHHQ00_1;
	wire w_dff_B_X2SMlDZf2_1;
	wire w_dff_B_Gp9j5lie5_1;
	wire w_dff_B_1xe2xa2b7_1;
	wire w_dff_B_xl4ky81B8_1;
	wire w_dff_B_Nf1JW0Sy8_1;
	wire w_dff_B_N3H7juG44_1;
	wire w_dff_B_RVBQFYe26_1;
	wire w_dff_B_SehHSgxe9_1;
	wire w_dff_B_q9NQ572J1_1;
	wire w_dff_B_WygCBZrl0_1;
	wire w_dff_B_iCdOZC8v7_1;
	wire w_dff_B_u78A3r9W2_1;
	wire w_dff_B_WRVShjn52_1;
	wire w_dff_B_oO46UanB4_1;
	wire w_dff_B_2ET4CGcy3_1;
	wire w_dff_B_3WVvWm4U8_1;
	wire w_dff_B_elvslTpM4_1;
	wire w_dff_B_0M3DidwV5_1;
	wire w_dff_B_OtgaCh0k0_1;
	wire w_dff_B_yzn87wbr0_1;
	wire w_dff_B_EtQioman0_1;
	wire w_dff_B_X4TrKgAK2_1;
	wire w_dff_B_12GyJk4w6_1;
	wire w_dff_B_1iR8VOcz6_1;
	wire w_dff_B_YDgGnJyk4_1;
	wire w_dff_B_TnMoPJkA0_1;
	wire w_dff_B_RrvzXPOb5_1;
	wire w_dff_B_KdMpr6kL5_1;
	wire w_dff_B_o6atlUfx5_1;
	wire w_dff_B_vA0AJS1L9_1;
	wire w_dff_B_G6sJ2W8p0_1;
	wire w_dff_B_mPQaqsW65_1;
	wire w_dff_B_0QETm1X44_1;
	wire w_dff_B_nOrAbU4z0_1;
	wire w_dff_B_JgYCvPNL1_1;
	wire w_dff_B_Sb8o7SrZ3_1;
	wire w_dff_B_Fx8y1IPI6_1;
	wire w_dff_B_BLTTxahc2_1;
	wire w_dff_B_eBj6S86y0_1;
	wire w_dff_B_7W2V7Ewn4_1;
	wire w_dff_B_jZPdK1kZ9_1;
	wire w_dff_B_NvPygvMp7_1;
	wire w_dff_B_Vor6ZZVU5_1;
	wire w_dff_B_vZsSDmqN4_1;
	wire w_dff_B_dtYczj4u5_1;
	wire w_dff_B_OcRBzI3e0_1;
	wire w_dff_B_6uWEU51u0_1;
	wire w_dff_B_CPLyEXKS6_1;
	wire w_dff_B_Arn7DGHt6_1;
	wire w_dff_B_ZbMRvaeY4_1;
	wire w_dff_B_Gg0qI4IW3_1;
	wire w_dff_B_KdYG81lr0_1;
	wire w_dff_B_DvnUCB5e3_1;
	wire w_dff_B_WB80gDUQ3_1;
	wire w_dff_B_GjGh3WJu0_0;
	wire w_dff_B_87AHIjf61_0;
	wire w_dff_B_vha20V114_0;
	wire w_dff_B_IIWhL9Oy6_0;
	wire w_dff_B_0xPVz5iZ6_0;
	wire w_dff_B_c73mP7TR4_0;
	wire w_dff_B_KMt2Vp601_0;
	wire w_dff_B_56mdr7yb8_0;
	wire w_dff_B_INlpUnzy1_0;
	wire w_dff_B_5iQ9aL7I9_0;
	wire w_dff_B_K2iAn8p76_0;
	wire w_dff_B_EHRxyDpz5_0;
	wire w_dff_B_tkwPMeTL4_0;
	wire w_dff_B_k2dibsWK2_0;
	wire w_dff_B_Z9ofRIyT9_0;
	wire w_dff_B_QMMpuiUz2_0;
	wire w_dff_B_kkRvZaQa9_0;
	wire w_dff_B_RrEFziYm2_0;
	wire w_dff_B_UkeEDUmI1_0;
	wire w_dff_B_thld9spP1_0;
	wire w_dff_B_5vfUe3Zu0_0;
	wire w_dff_B_YNbHDSyk2_0;
	wire w_dff_B_XPehuPkM0_0;
	wire w_dff_B_ZdPUWvF32_0;
	wire w_dff_B_xelrXhYO3_0;
	wire w_dff_B_4mo0fLKN6_0;
	wire w_dff_B_JNHaoWyZ1_0;
	wire w_dff_B_bZujMI7a4_0;
	wire w_dff_B_axWWilLA8_0;
	wire w_dff_B_nyEmfRx03_0;
	wire w_dff_B_xxQqm72r2_0;
	wire w_dff_B_sJLemPYT6_0;
	wire w_dff_B_7sprYiKU5_0;
	wire w_dff_B_e76x8MDY9_0;
	wire w_dff_B_KrEvJ6Em0_0;
	wire w_dff_B_9VOd76IC5_0;
	wire w_dff_B_kdcXW1Dn7_0;
	wire w_dff_B_a3CTIul14_0;
	wire w_dff_B_GtMlnX143_0;
	wire w_dff_B_kF67EOkP8_0;
	wire w_dff_B_dvgxW1fE9_0;
	wire w_dff_B_fqpPdD304_0;
	wire w_dff_B_CAJyC8AI6_0;
	wire w_dff_B_NsncFfJi6_0;
	wire w_dff_B_1Sn1fci71_0;
	wire w_dff_B_cartHQiF5_0;
	wire w_dff_B_K7ajf5zH2_0;
	wire w_dff_B_9T7E4BJm4_0;
	wire w_dff_B_cBsNe0Kj1_0;
	wire w_dff_B_EhJ4eNRk3_0;
	wire w_dff_B_JzYWfGWg9_0;
	wire w_dff_B_6VMSdjb25_0;
	wire w_dff_B_3pd9mDXE9_0;
	wire w_dff_B_Ti5ZiTDw4_0;
	wire w_dff_B_Y8s4ZyLT4_0;
	wire w_dff_B_rQT0WRwO0_0;
	wire w_dff_B_QNrAjY2s8_0;
	wire w_dff_B_THshr7nV5_0;
	wire w_dff_B_q2b5Mr069_0;
	wire w_dff_B_QcFVbgt62_0;
	wire w_dff_B_npoZexg99_0;
	wire w_dff_B_eyeMZbHu8_0;
	wire w_dff_B_gpj5eUpe6_0;
	wire w_dff_B_RTy8gz0z3_0;
	wire w_dff_B_NN3NZ2ah9_0;
	wire w_dff_B_hhjmCZRY8_0;
	wire w_dff_B_dAOVQXDY8_0;
	wire w_dff_B_fsAZWSZI7_0;
	wire w_dff_B_M5DZCPvj6_0;
	wire w_dff_B_pdNiP3hC7_0;
	wire w_dff_B_W2REQXXw7_0;
	wire w_dff_B_r47RgOHP5_0;
	wire w_dff_B_V7Vyc3sJ1_0;
	wire w_dff_B_S4OLg2yr2_0;
	wire w_dff_B_ar8XvTH63_0;
	wire w_dff_B_pJ7az45L4_0;
	wire w_dff_B_ag80TtA29_0;
	wire w_dff_B_udxludNu2_0;
	wire w_dff_B_c4uWKt9O0_0;
	wire w_dff_B_d8k9JwJL6_0;
	wire w_dff_B_KQa96zfY2_0;
	wire w_dff_B_HMMi7YPO4_0;
	wire w_dff_B_VMDwLyZ19_0;
	wire w_dff_B_x1VH9U9f5_0;
	wire w_dff_B_e5ZhdMUD9_0;
	wire w_dff_B_c32iPo0W0_0;
	wire w_dff_B_NvmzhQFe8_0;
	wire w_dff_B_QJlmnVcJ9_0;
	wire w_dff_B_OwnieKJd8_0;
	wire w_dff_B_fdbEgXEg2_0;
	wire w_dff_B_FiNcMpAP6_0;
	wire w_dff_B_X7BNpBXy1_0;
	wire w_dff_B_DfkeKuht3_0;
	wire w_dff_B_0kwJxems0_0;
	wire w_dff_B_rO5HQhB26_0;
	wire w_dff_B_mULJ6y7Q6_0;
	wire w_dff_B_XE2iBHU27_0;
	wire w_dff_B_X6k1QGWv0_1;
	wire w_dff_B_OhruMBzk6_1;
	wire w_dff_B_gsAuGk6a3_1;
	wire w_dff_B_qDbiWVZy8_1;
	wire w_dff_B_mdI0Fwlk3_1;
	wire w_dff_B_v0aIkXA33_1;
	wire w_dff_B_eoAtNEcx1_1;
	wire w_dff_B_tYpqItOU8_1;
	wire w_dff_B_PgdDTKDx1_1;
	wire w_dff_B_3mETEtpF9_1;
	wire w_dff_B_fTJalLeC5_1;
	wire w_dff_B_1HEa7eRm2_1;
	wire w_dff_B_hlHz8Q0g6_1;
	wire w_dff_B_tEVcGN6p7_1;
	wire w_dff_B_ECeAd9Bq2_1;
	wire w_dff_B_JMLzCD4R4_1;
	wire w_dff_B_UdIWccTE0_1;
	wire w_dff_B_BpAHrHRS0_1;
	wire w_dff_B_BBfgyF8V9_1;
	wire w_dff_B_tHrlVO5A4_1;
	wire w_dff_B_bdKhbPu02_1;
	wire w_dff_B_ndFRSCRI2_1;
	wire w_dff_B_8jsUJxoz9_1;
	wire w_dff_B_LN3jD4Wz5_1;
	wire w_dff_B_IiLloUit1_1;
	wire w_dff_B_gaRITIlM0_1;
	wire w_dff_B_Eyru6rLW5_1;
	wire w_dff_B_prMpyePJ0_1;
	wire w_dff_B_M0QL4oJg0_1;
	wire w_dff_B_mW5VNVn62_1;
	wire w_dff_B_IYu9f9W17_1;
	wire w_dff_B_8aiJyBES7_1;
	wire w_dff_B_OvqpOZDC8_1;
	wire w_dff_B_iVESutl40_1;
	wire w_dff_B_j1Bhpc6S4_1;
	wire w_dff_B_sR7Zp4OF8_1;
	wire w_dff_B_CQ8Y6tTp1_1;
	wire w_dff_B_MFws36604_1;
	wire w_dff_B_XtPZyC9D8_1;
	wire w_dff_B_Tmu3Mwki4_1;
	wire w_dff_B_GC8IoMHt4_1;
	wire w_dff_B_voBOfHj30_1;
	wire w_dff_B_01dYlaXF0_1;
	wire w_dff_B_5k79iCEF9_1;
	wire w_dff_B_z15N4nXr3_1;
	wire w_dff_B_cmbJVVmN0_1;
	wire w_dff_B_uVjcN9o64_1;
	wire w_dff_B_C5TPksbH6_1;
	wire w_dff_B_itlApGNA6_1;
	wire w_dff_B_Kv4cd13c7_1;
	wire w_dff_B_fEarABeZ6_1;
	wire w_dff_B_kVYTvMoH9_1;
	wire w_dff_B_c9ljnnf46_1;
	wire w_dff_B_bIXfaSag4_1;
	wire w_dff_B_gUG2cZ7F5_1;
	wire w_dff_B_edydH8W29_1;
	wire w_dff_B_a3cgnRV14_1;
	wire w_dff_B_WA2kttRh7_1;
	wire w_dff_B_gSjKMQhC3_1;
	wire w_dff_B_uorQ4rQZ4_1;
	wire w_dff_B_8UMElZlA7_1;
	wire w_dff_B_JT2icPdU2_1;
	wire w_dff_B_jFKnzbEl5_1;
	wire w_dff_B_ODhwVTrS3_1;
	wire w_dff_B_48nzjYbs5_1;
	wire w_dff_B_Rsc1aUEr9_1;
	wire w_dff_B_Z7YP2Vpt9_1;
	wire w_dff_B_9sDBfI0c8_1;
	wire w_dff_B_hiEntRbO6_1;
	wire w_dff_B_1gglhluY3_1;
	wire w_dff_B_dStCm4rp2_1;
	wire w_dff_B_aiL9QGwt6_1;
	wire w_dff_B_1Mm6isHR0_1;
	wire w_dff_B_N1y6wS8K6_1;
	wire w_dff_B_HyXTneoF4_1;
	wire w_dff_B_ezmF7k1U0_1;
	wire w_dff_B_t0svJczu1_1;
	wire w_dff_B_NGAQV2UX8_1;
	wire w_dff_B_etEj1QAX0_1;
	wire w_dff_B_JXLDJJ4g0_1;
	wire w_dff_B_17ZWHBFQ0_1;
	wire w_dff_B_91IWJTxR5_1;
	wire w_dff_B_xfwwyH7Y4_1;
	wire w_dff_B_0LZhZyG82_1;
	wire w_dff_B_Tm3iqxpu1_1;
	wire w_dff_B_gNXKhCuS8_1;
	wire w_dff_B_Ju22jkuY5_1;
	wire w_dff_B_nMUlxsrx1_1;
	wire w_dff_B_SUXm0i3Q9_1;
	wire w_dff_B_7YGRiLKz7_1;
	wire w_dff_B_wS9Y9S1n7_1;
	wire w_dff_B_o6dyVh8f7_1;
	wire w_dff_B_mGVgvzrS8_1;
	wire w_dff_B_zk07ZSL38_1;
	wire w_dff_B_66FJgh837_1;
	wire w_dff_B_i16ixeFE0_1;
	wire w_dff_B_pB9ohBpz5_0;
	wire w_dff_B_qN5gVHgU3_0;
	wire w_dff_B_4t1mlIvC3_0;
	wire w_dff_B_FURDTsYV5_0;
	wire w_dff_B_MBdieqMe0_0;
	wire w_dff_B_BfFCQTJe0_0;
	wire w_dff_B_EFUNuYVk1_0;
	wire w_dff_B_yMFnqjzX7_0;
	wire w_dff_B_4T15hbcn8_0;
	wire w_dff_B_AvT02vpZ9_0;
	wire w_dff_B_1xIKDRRx5_0;
	wire w_dff_B_QTM9pWrH4_0;
	wire w_dff_B_IM8AeYQh7_0;
	wire w_dff_B_5owa66a82_0;
	wire w_dff_B_m2vHSqeq3_0;
	wire w_dff_B_UNtdUWQm7_0;
	wire w_dff_B_lIOBYjns0_0;
	wire w_dff_B_2faxuY1F8_0;
	wire w_dff_B_PM3aSWS50_0;
	wire w_dff_B_Is3GgUso7_0;
	wire w_dff_B_4UZQvBcp9_0;
	wire w_dff_B_hvYMu4RO9_0;
	wire w_dff_B_jx8JTva21_0;
	wire w_dff_B_h27Zusum7_0;
	wire w_dff_B_m1Zy5TGV2_0;
	wire w_dff_B_ZtObcjWI4_0;
	wire w_dff_B_5LIHS1Z84_0;
	wire w_dff_B_avFI0M5V7_0;
	wire w_dff_B_9TosqZQv6_0;
	wire w_dff_B_dKLAarJG8_0;
	wire w_dff_B_IF2GADLm1_0;
	wire w_dff_B_7izdc4V76_0;
	wire w_dff_B_RGkywMA92_0;
	wire w_dff_B_xjN6BYGZ6_0;
	wire w_dff_B_RsrFWTXq7_0;
	wire w_dff_B_zNMF2o3f1_0;
	wire w_dff_B_UbMj15YF7_0;
	wire w_dff_B_cZ5BOPwq0_0;
	wire w_dff_B_qUsKM4NW5_0;
	wire w_dff_B_uEIeSmiW0_0;
	wire w_dff_B_mXB4ko7Q7_0;
	wire w_dff_B_Y5CH93RO1_0;
	wire w_dff_B_rJlmCpRD9_0;
	wire w_dff_B_BDrkrepj7_0;
	wire w_dff_B_A92dBLID0_0;
	wire w_dff_B_Zzoca1WP0_0;
	wire w_dff_B_J7xGRWWQ8_0;
	wire w_dff_B_jfthEalt2_0;
	wire w_dff_B_UaJJ4Jr95_0;
	wire w_dff_B_K5ygOkS13_0;
	wire w_dff_B_PN1cuHp77_0;
	wire w_dff_B_GejEV5Eg6_0;
	wire w_dff_B_pY928UbG4_0;
	wire w_dff_B_vJdTy1Ut0_0;
	wire w_dff_B_Yi05wNmp9_0;
	wire w_dff_B_CJr9sUpv0_0;
	wire w_dff_B_1olkKZCp9_0;
	wire w_dff_B_Yh6q8TR29_0;
	wire w_dff_B_iXekFgxa6_0;
	wire w_dff_B_crnV6jVU5_0;
	wire w_dff_B_KzHaswyh6_0;
	wire w_dff_B_knf8fCeI9_0;
	wire w_dff_B_NaGBnOLk0_0;
	wire w_dff_B_jL9UKd2c2_0;
	wire w_dff_B_W3sTHeaQ4_0;
	wire w_dff_B_smls63i15_0;
	wire w_dff_B_rbMoLEQl6_0;
	wire w_dff_B_C6MyzLOf9_0;
	wire w_dff_B_YttT4K8E7_0;
	wire w_dff_B_A8X96XcQ6_0;
	wire w_dff_B_0X58FGYH0_0;
	wire w_dff_B_CQz7a8gO4_0;
	wire w_dff_B_zhWzqRpU0_0;
	wire w_dff_B_5sh32TL86_0;
	wire w_dff_B_34Xqphlm5_0;
	wire w_dff_B_SHxPIKwg2_0;
	wire w_dff_B_78ZLS5812_0;
	wire w_dff_B_MksQTyno0_0;
	wire w_dff_B_zdOcxGy39_0;
	wire w_dff_B_wsW4U1dB3_0;
	wire w_dff_B_w98e7xUS0_0;
	wire w_dff_B_pdbfvMqH3_0;
	wire w_dff_B_5cks2KkI7_0;
	wire w_dff_B_7sd8C4268_0;
	wire w_dff_B_sfEETGGb8_0;
	wire w_dff_B_pVwxEO8f4_0;
	wire w_dff_B_Ob5xSnvX8_0;
	wire w_dff_B_9a0vFLUn0_0;
	wire w_dff_B_S9GyfjEX9_0;
	wire w_dff_B_qiQhmBhK7_0;
	wire w_dff_B_zfZaybuE0_0;
	wire w_dff_B_R8gm21p73_0;
	wire w_dff_B_X1oxPpZf6_0;
	wire w_dff_B_lxbb6iv81_0;
	wire w_dff_B_5r1rrR6p3_0;
	wire w_dff_B_3XsPByS46_0;
	wire w_dff_B_5h5pEzoJ1_1;
	wire w_dff_B_TW22cvRH5_1;
	wire w_dff_B_34SK0ARe2_1;
	wire w_dff_B_J7p5oi1M9_1;
	wire w_dff_B_GHZwEY2s1_1;
	wire w_dff_B_g2jdiwii1_1;
	wire w_dff_B_svz0r1ll2_1;
	wire w_dff_B_s4S94kZ96_1;
	wire w_dff_B_f7AWNVNL8_1;
	wire w_dff_B_tfsKzCkX8_1;
	wire w_dff_B_1EsPREt61_1;
	wire w_dff_B_sEmo0SZx6_1;
	wire w_dff_B_fZEKeNit1_1;
	wire w_dff_B_1xevbUJr4_1;
	wire w_dff_B_k0KJEXRo3_1;
	wire w_dff_B_KGEILHza1_1;
	wire w_dff_B_FfVwj9YX7_1;
	wire w_dff_B_3ASk24GQ2_1;
	wire w_dff_B_NlwZVyxn1_1;
	wire w_dff_B_7pbXjwHD1_1;
	wire w_dff_B_Gg6UT4Z16_1;
	wire w_dff_B_aa0nRbpH3_1;
	wire w_dff_B_0InrlveO2_1;
	wire w_dff_B_1WjlFOcE2_1;
	wire w_dff_B_S8jNN0zf1_1;
	wire w_dff_B_SuZBlx139_1;
	wire w_dff_B_3AMKNiPJ1_1;
	wire w_dff_B_jUzV742W3_1;
	wire w_dff_B_FNbz4A4v3_1;
	wire w_dff_B_ec8KbeNC6_1;
	wire w_dff_B_LUTxwJ8h0_1;
	wire w_dff_B_CahfPJlh5_1;
	wire w_dff_B_lx8D4W2E5_1;
	wire w_dff_B_qbMiveIy7_1;
	wire w_dff_B_dwX66ODU5_1;
	wire w_dff_B_hb4NwXxJ8_1;
	wire w_dff_B_pLZg3z3p0_1;
	wire w_dff_B_GF7WkCUh3_1;
	wire w_dff_B_lBmk3FQv6_1;
	wire w_dff_B_rJkdbwcB7_1;
	wire w_dff_B_pjohpkrt4_1;
	wire w_dff_B_iwgyciuB1_1;
	wire w_dff_B_GO4a9lSi5_1;
	wire w_dff_B_WSA9MvCL1_1;
	wire w_dff_B_kL7HkD6D4_1;
	wire w_dff_B_EioNTpVY9_1;
	wire w_dff_B_LNBmf1Xn8_1;
	wire w_dff_B_d9FZL5962_1;
	wire w_dff_B_RWQrh6mq0_1;
	wire w_dff_B_9XaHFRwg9_1;
	wire w_dff_B_xxKQ4Ia91_1;
	wire w_dff_B_qCh9Ijb56_1;
	wire w_dff_B_m1QcDzfL5_1;
	wire w_dff_B_UvLUOwdL7_1;
	wire w_dff_B_af2ln9mi4_1;
	wire w_dff_B_2l1X0JWa3_1;
	wire w_dff_B_azVg8IOu7_1;
	wire w_dff_B_h6ukKkiD4_1;
	wire w_dff_B_c1aLeOMc0_1;
	wire w_dff_B_Z2zhRQzZ5_1;
	wire w_dff_B_Z2l5jexn7_1;
	wire w_dff_B_PQjUwcbL3_1;
	wire w_dff_B_K8NNNrRb2_1;
	wire w_dff_B_R3hbC0lI4_1;
	wire w_dff_B_kBZLhqis3_1;
	wire w_dff_B_pBhMXUKh1_1;
	wire w_dff_B_vodXbVJ26_1;
	wire w_dff_B_EDTYywnX5_1;
	wire w_dff_B_Ci0YArzd4_1;
	wire w_dff_B_4j9UoHSZ4_1;
	wire w_dff_B_l9QuPTnE5_1;
	wire w_dff_B_IdMkGcYU3_1;
	wire w_dff_B_oaAdyzia2_1;
	wire w_dff_B_AKnU10zy5_1;
	wire w_dff_B_hK7GLm3G0_1;
	wire w_dff_B_4EnP114U3_1;
	wire w_dff_B_htkj9dM24_1;
	wire w_dff_B_VuImE7Zp1_1;
	wire w_dff_B_V79VZpFO3_1;
	wire w_dff_B_O1HARNWQ3_1;
	wire w_dff_B_Z2mbYRCK4_1;
	wire w_dff_B_aKjDdA3e7_1;
	wire w_dff_B_e8ZoBi5d2_1;
	wire w_dff_B_mRoO8x6R9_1;
	wire w_dff_B_fIOfh2wh3_1;
	wire w_dff_B_kR8LnsSr2_1;
	wire w_dff_B_W13wPvvM4_1;
	wire w_dff_B_HNZ5Rhd77_1;
	wire w_dff_B_AeohlU5a3_1;
	wire w_dff_B_Rugfoc3L6_1;
	wire w_dff_B_FndFkS8U0_1;
	wire w_dff_B_6tvLxXyI9_1;
	wire w_dff_B_l2Y8TxU44_1;
	wire w_dff_B_fqdrpVbN6_1;
	wire w_dff_B_Jf6mJkjd5_1;
	wire w_dff_B_i8hjuhlu9_0;
	wire w_dff_B_76ubyzjk6_0;
	wire w_dff_B_2JUcnE6Z6_0;
	wire w_dff_B_5kkV5XQC7_0;
	wire w_dff_B_aSytXVeC2_0;
	wire w_dff_B_QJPEGd597_0;
	wire w_dff_B_5vittjnS2_0;
	wire w_dff_B_PR9goVpm3_0;
	wire w_dff_B_RP3oI6Nd4_0;
	wire w_dff_B_VLf54wtn9_0;
	wire w_dff_B_pzfAHvHI0_0;
	wire w_dff_B_ceaM2JMS6_0;
	wire w_dff_B_hXAQVowD9_0;
	wire w_dff_B_qEQVx2xH9_0;
	wire w_dff_B_MuLgi9Fk0_0;
	wire w_dff_B_xbaeqHf26_0;
	wire w_dff_B_WvpMQQrw0_0;
	wire w_dff_B_NaE259Mg0_0;
	wire w_dff_B_GA25x1Px6_0;
	wire w_dff_B_71eXY0lQ7_0;
	wire w_dff_B_JbEUF7ot4_0;
	wire w_dff_B_Umb7swJJ7_0;
	wire w_dff_B_FnUuINN84_0;
	wire w_dff_B_Uu3FwLVp4_0;
	wire w_dff_B_AHExV0Qf9_0;
	wire w_dff_B_7VMRMB8y0_0;
	wire w_dff_B_CDaOiJ8J3_0;
	wire w_dff_B_iXaF2lDd6_0;
	wire w_dff_B_qtMibAbp3_0;
	wire w_dff_B_xAxUj8Os9_0;
	wire w_dff_B_VFQ2YYTI0_0;
	wire w_dff_B_B1jgPaIN5_0;
	wire w_dff_B_L5f7ZURS5_0;
	wire w_dff_B_DaGiZrT46_0;
	wire w_dff_B_nJ4Ku9xO9_0;
	wire w_dff_B_w0F39Ppm7_0;
	wire w_dff_B_yu8tBKAE9_0;
	wire w_dff_B_CjkOfixa4_0;
	wire w_dff_B_S90VgQyU2_0;
	wire w_dff_B_eDsKeAmE1_0;
	wire w_dff_B_haItXVPK8_0;
	wire w_dff_B_VgwNIEZi6_0;
	wire w_dff_B_ezp1duFy8_0;
	wire w_dff_B_1zbwQ8W52_0;
	wire w_dff_B_FWRkZ8sw0_0;
	wire w_dff_B_6UqfWH3R3_0;
	wire w_dff_B_6V0miGFq3_0;
	wire w_dff_B_6r4CoxRh4_0;
	wire w_dff_B_GwnGBeS01_0;
	wire w_dff_B_lemZ41vD2_0;
	wire w_dff_B_SM5vYIv53_0;
	wire w_dff_B_iYKu0jZI7_0;
	wire w_dff_B_xWCNrAXh6_0;
	wire w_dff_B_THDKSGDB9_0;
	wire w_dff_B_zJsyjVAl8_0;
	wire w_dff_B_UoGT25TO7_0;
	wire w_dff_B_3BTz2QOv8_0;
	wire w_dff_B_d8DVl0Zv9_0;
	wire w_dff_B_ghMBkZe21_0;
	wire w_dff_B_irOuD0Bm1_0;
	wire w_dff_B_lgET5Av46_0;
	wire w_dff_B_aK22A6Ah9_0;
	wire w_dff_B_xhbP446k1_0;
	wire w_dff_B_b8voxjEf1_0;
	wire w_dff_B_WYhARzM81_0;
	wire w_dff_B_kFiFUhd77_0;
	wire w_dff_B_im71HWpd0_0;
	wire w_dff_B_g2Gqysx42_0;
	wire w_dff_B_cgxSuDDf5_0;
	wire w_dff_B_MlQT6Hfu7_0;
	wire w_dff_B_HjqrmXjg3_0;
	wire w_dff_B_sGzGMXpn6_0;
	wire w_dff_B_wRIOv2bx6_0;
	wire w_dff_B_DaHKbmqu1_0;
	wire w_dff_B_x1fxOtZK0_0;
	wire w_dff_B_65OhVyop0_0;
	wire w_dff_B_aYKMZH9H4_0;
	wire w_dff_B_sW0rXPWk3_0;
	wire w_dff_B_lZ9HvCBD6_0;
	wire w_dff_B_vkmjfrXb3_0;
	wire w_dff_B_2xHZtOgN5_0;
	wire w_dff_B_qluoOv0f5_0;
	wire w_dff_B_bQ5oZYPx1_0;
	wire w_dff_B_CSdErt2L5_0;
	wire w_dff_B_w4uv4KX34_0;
	wire w_dff_B_DrNNixjE3_0;
	wire w_dff_B_GsquZjmj7_0;
	wire w_dff_B_JLDbsI091_0;
	wire w_dff_B_laECUqgj7_0;
	wire w_dff_B_h80dNyXL3_0;
	wire w_dff_B_vfu81PqA8_0;
	wire w_dff_B_JqtnApUX2_0;
	wire w_dff_B_7QfGz7AH0_0;
	wire w_dff_B_l5iuMxeB6_0;
	wire w_dff_B_gF4cW8n67_0;
	wire w_dff_B_V4Id4OKl3_1;
	wire w_dff_B_FUwoILhq4_1;
	wire w_dff_B_gOmB6Gj76_1;
	wire w_dff_B_jqRGrULa6_1;
	wire w_dff_B_W8txnoBr5_1;
	wire w_dff_B_ak6byy5r4_1;
	wire w_dff_B_PXvfUu7z8_1;
	wire w_dff_B_JM3H6XI40_1;
	wire w_dff_B_VVtGThzh2_1;
	wire w_dff_B_QDX8E3WK0_1;
	wire w_dff_B_PyLaqtzv6_1;
	wire w_dff_B_D4rFeW5n7_1;
	wire w_dff_B_vtFGlBHl9_1;
	wire w_dff_B_YL9ZDojH2_1;
	wire w_dff_B_vww5tgWF5_1;
	wire w_dff_B_uR5b9UZr9_1;
	wire w_dff_B_nUOTufvf3_1;
	wire w_dff_B_KcqX1aL82_1;
	wire w_dff_B_efyeNG8K8_1;
	wire w_dff_B_1njcdvY62_1;
	wire w_dff_B_7eyUq7aC7_1;
	wire w_dff_B_ev5jeRdp2_1;
	wire w_dff_B_nOTZb0mq6_1;
	wire w_dff_B_g5AosEdZ8_1;
	wire w_dff_B_axowICWa3_1;
	wire w_dff_B_sNAt40SC3_1;
	wire w_dff_B_K9tW33W14_1;
	wire w_dff_B_JByQrClz1_1;
	wire w_dff_B_qxZzGxFs4_1;
	wire w_dff_B_dTiwJBqc5_1;
	wire w_dff_B_TYG1D1pQ0_1;
	wire w_dff_B_Ob6aHVnN7_1;
	wire w_dff_B_jwyhO8Vs8_1;
	wire w_dff_B_7AnpxpV43_1;
	wire w_dff_B_OkSfpMsf8_1;
	wire w_dff_B_WCrdtPIC6_1;
	wire w_dff_B_ElMsHhza8_1;
	wire w_dff_B_RHRuAJWm6_1;
	wire w_dff_B_PyBmSSVk2_1;
	wire w_dff_B_B7CZDynS5_1;
	wire w_dff_B_50wj6ssY4_1;
	wire w_dff_B_lOZSlXPt3_1;
	wire w_dff_B_ODOVFQ8H0_1;
	wire w_dff_B_JGTGbXnm5_1;
	wire w_dff_B_DMB2Lh6Q1_1;
	wire w_dff_B_dhqkdMmc0_1;
	wire w_dff_B_5fkAPVop7_1;
	wire w_dff_B_CfX0MTeq8_1;
	wire w_dff_B_f3zwWfhV4_1;
	wire w_dff_B_3WLiYBPk8_1;
	wire w_dff_B_xGimSENv5_1;
	wire w_dff_B_CKn9l4Kr1_1;
	wire w_dff_B_9ocvr2sP9_1;
	wire w_dff_B_O20G46hs7_1;
	wire w_dff_B_PoK5GwyZ2_1;
	wire w_dff_B_Cv7ae5305_1;
	wire w_dff_B_mGo7EScm5_1;
	wire w_dff_B_lWeG9KZw3_1;
	wire w_dff_B_LX5pjq8p0_1;
	wire w_dff_B_O7S507ih5_1;
	wire w_dff_B_YfIyJNHL8_1;
	wire w_dff_B_zJTwdKRq9_1;
	wire w_dff_B_m8jD3M1a0_1;
	wire w_dff_B_igDalDOA5_1;
	wire w_dff_B_73dKzfCz6_1;
	wire w_dff_B_RTDxXUBi6_1;
	wire w_dff_B_Gzeak3hw2_1;
	wire w_dff_B_ndxTx1pN5_1;
	wire w_dff_B_5dI8zPV48_1;
	wire w_dff_B_OtzK438z1_1;
	wire w_dff_B_UN7YaIu62_1;
	wire w_dff_B_RwGBgBiC1_1;
	wire w_dff_B_sfZVOxTI8_1;
	wire w_dff_B_q7asw41e8_1;
	wire w_dff_B_lrD7kicI6_1;
	wire w_dff_B_7dA3H1dG9_1;
	wire w_dff_B_MBBr2bSI5_1;
	wire w_dff_B_taRdgtTr3_1;
	wire w_dff_B_SDLOufBX6_1;
	wire w_dff_B_TIWcSlAI4_1;
	wire w_dff_B_dEodIcwZ0_1;
	wire w_dff_B_yGIVbhBp8_1;
	wire w_dff_B_pW7hpMga7_1;
	wire w_dff_B_07A6QlD61_1;
	wire w_dff_B_1SKjaigN2_1;
	wire w_dff_B_vpwAAi2W0_1;
	wire w_dff_B_Vdv0FRq96_1;
	wire w_dff_B_I9OgCQ9m8_1;
	wire w_dff_B_nSgMasaR8_1;
	wire w_dff_B_jablWl1A6_1;
	wire w_dff_B_x0zFPHjr0_1;
	wire w_dff_B_HY9tid950_1;
	wire w_dff_B_prkOEvLy1_1;
	wire w_dff_B_gjoULGb32_1;
	wire w_dff_B_zIDCfSlT4_0;
	wire w_dff_B_MRH0kbpu9_0;
	wire w_dff_B_7ZV0rU0I7_0;
	wire w_dff_B_Y1Z3YWoP0_0;
	wire w_dff_B_vP4xMjMZ2_0;
	wire w_dff_B_wgVcbYj93_0;
	wire w_dff_B_RedyTcYe6_0;
	wire w_dff_B_mqeMtM671_0;
	wire w_dff_B_J1cb6B2A0_0;
	wire w_dff_B_91c1GROD5_0;
	wire w_dff_B_vVVEWpUC4_0;
	wire w_dff_B_d3JOicTv0_0;
	wire w_dff_B_fQw0xfZT9_0;
	wire w_dff_B_ztxYsfqY5_0;
	wire w_dff_B_5vK0gKNH0_0;
	wire w_dff_B_a46F5i661_0;
	wire w_dff_B_VO89RzTc6_0;
	wire w_dff_B_TOZpVuYs8_0;
	wire w_dff_B_tcfODsTj9_0;
	wire w_dff_B_Ddb5UEzH3_0;
	wire w_dff_B_rbOTEwN20_0;
	wire w_dff_B_JuoW0pJP8_0;
	wire w_dff_B_DXGRnf9x0_0;
	wire w_dff_B_QkUpHHBg5_0;
	wire w_dff_B_Ny9nz9O93_0;
	wire w_dff_B_hGEzkZkF7_0;
	wire w_dff_B_8b7OOEIj0_0;
	wire w_dff_B_Db4PHfoP2_0;
	wire w_dff_B_f6hIX16U3_0;
	wire w_dff_B_WngVcNBa7_0;
	wire w_dff_B_It7XBfVE7_0;
	wire w_dff_B_vf99utdR5_0;
	wire w_dff_B_CJ835o1m4_0;
	wire w_dff_B_kU7BB5eZ1_0;
	wire w_dff_B_Mt64mcxQ1_0;
	wire w_dff_B_9tpLwi0n1_0;
	wire w_dff_B_X769e3gl8_0;
	wire w_dff_B_wCynEx8b6_0;
	wire w_dff_B_nPENxYqD9_0;
	wire w_dff_B_8LAVOjQi0_0;
	wire w_dff_B_C4fUTGvb4_0;
	wire w_dff_B_mQJFSKgO3_0;
	wire w_dff_B_mxi2saeZ8_0;
	wire w_dff_B_dhazEBQh2_0;
	wire w_dff_B_narvYCok5_0;
	wire w_dff_B_HZYWSKlb8_0;
	wire w_dff_B_qxmaXVaL1_0;
	wire w_dff_B_exqnjkt53_0;
	wire w_dff_B_GMIO81oT5_0;
	wire w_dff_B_8oGHIq6R9_0;
	wire w_dff_B_JL310I535_0;
	wire w_dff_B_WNY353GA7_0;
	wire w_dff_B_Z8jo0LFH6_0;
	wire w_dff_B_iLpQhrys9_0;
	wire w_dff_B_grDKkQ9S1_0;
	wire w_dff_B_YMInR4TI5_0;
	wire w_dff_B_YpBGOVyZ3_0;
	wire w_dff_B_xOTPnXLV3_0;
	wire w_dff_B_kfb600uh7_0;
	wire w_dff_B_MbfewOqH4_0;
	wire w_dff_B_EeUGYaSy1_0;
	wire w_dff_B_sbNHupP22_0;
	wire w_dff_B_U6z1YcMv7_0;
	wire w_dff_B_TFRxEf5t4_0;
	wire w_dff_B_AV1Y5qNW1_0;
	wire w_dff_B_rZ5LQRvG9_0;
	wire w_dff_B_W6Urze7c0_0;
	wire w_dff_B_2QpAcxgm7_0;
	wire w_dff_B_ic3lSNup9_0;
	wire w_dff_B_oLoM5QvQ7_0;
	wire w_dff_B_UPe20AvG6_0;
	wire w_dff_B_ifnVewRr5_0;
	wire w_dff_B_NPkroi0A1_0;
	wire w_dff_B_irbehqs29_0;
	wire w_dff_B_vZDPM6ka0_0;
	wire w_dff_B_711Y4oqI9_0;
	wire w_dff_B_j5S9OtfC6_0;
	wire w_dff_B_VGSlfaPw1_0;
	wire w_dff_B_ZCImlmkd5_0;
	wire w_dff_B_eJoBJKN96_0;
	wire w_dff_B_jbulfgBo7_0;
	wire w_dff_B_TFUZBVYt3_0;
	wire w_dff_B_cbkSIbUg6_0;
	wire w_dff_B_N8TKDq7N2_0;
	wire w_dff_B_5R023Dvz3_0;
	wire w_dff_B_Z81DTIDr7_0;
	wire w_dff_B_EF3hGMje8_0;
	wire w_dff_B_CuIHmZcq4_0;
	wire w_dff_B_Qd2FPUwi0_0;
	wire w_dff_B_q3n5TzjL9_0;
	wire w_dff_B_YuvgbGU55_0;
	wire w_dff_B_bzPWadtA9_0;
	wire w_dff_B_G4FiTUOn2_0;
	wire w_dff_B_Tlk8jcgs4_0;
	wire w_dff_B_NIPgnmvE5_1;
	wire w_dff_B_GNazyr6z7_1;
	wire w_dff_B_SRafIkTg8_1;
	wire w_dff_B_jfyKVKxb6_1;
	wire w_dff_B_Gqoq2WRY9_1;
	wire w_dff_B_hOjwb8ou8_1;
	wire w_dff_B_nmnt5xcc6_1;
	wire w_dff_B_qfNir07L8_1;
	wire w_dff_B_tjXsTbGM0_1;
	wire w_dff_B_yThbUDN74_1;
	wire w_dff_B_i8uCCkZj0_1;
	wire w_dff_B_jc9rBImC3_1;
	wire w_dff_B_sQd0kZYn2_1;
	wire w_dff_B_qfWNX0J09_1;
	wire w_dff_B_GWYui08G5_1;
	wire w_dff_B_8HrnCfnF9_1;
	wire w_dff_B_9Psa5Rir3_1;
	wire w_dff_B_0pvI4qSP4_1;
	wire w_dff_B_8NRA4ImH2_1;
	wire w_dff_B_K3liEBnP7_1;
	wire w_dff_B_CaDbtZGg6_1;
	wire w_dff_B_LWQCpjxd2_1;
	wire w_dff_B_ZP2U6ziC1_1;
	wire w_dff_B_6dO1q6LA8_1;
	wire w_dff_B_3UhEkn1c9_1;
	wire w_dff_B_aqhEYIpX5_1;
	wire w_dff_B_TUtVtCGX2_1;
	wire w_dff_B_8f0LtSgp4_1;
	wire w_dff_B_aSMH59jL4_1;
	wire w_dff_B_ihorJH7F9_1;
	wire w_dff_B_uJabjRPI5_1;
	wire w_dff_B_prlyCjJM6_1;
	wire w_dff_B_xqfmdQEK4_1;
	wire w_dff_B_UTUw33b70_1;
	wire w_dff_B_YuVuYVtA3_1;
	wire w_dff_B_y3eYixxI9_1;
	wire w_dff_B_4Z6DRA540_1;
	wire w_dff_B_4bmZvCzy4_1;
	wire w_dff_B_4hvkd2lt9_1;
	wire w_dff_B_Agmltuqy7_1;
	wire w_dff_B_02laE88z8_1;
	wire w_dff_B_VZAiEAtY7_1;
	wire w_dff_B_U9UiiICj9_1;
	wire w_dff_B_mhImDYsm1_1;
	wire w_dff_B_vkZSsfgU6_1;
	wire w_dff_B_UzAKZNwJ9_1;
	wire w_dff_B_M0O8gISK1_1;
	wire w_dff_B_URlhlWey0_1;
	wire w_dff_B_uUawEShs2_1;
	wire w_dff_B_lRsGibNx9_1;
	wire w_dff_B_EVhfsF6W8_1;
	wire w_dff_B_aE2G8XQ32_1;
	wire w_dff_B_QTu7zUnH1_1;
	wire w_dff_B_evK6g61U2_1;
	wire w_dff_B_F1YmhZjp0_1;
	wire w_dff_B_BJPIFfZJ7_1;
	wire w_dff_B_v4m9yThQ1_1;
	wire w_dff_B_1Rcas2YK4_1;
	wire w_dff_B_hU198oK02_1;
	wire w_dff_B_YRXOFSQW0_1;
	wire w_dff_B_OsRxHc9o2_1;
	wire w_dff_B_HyBK42dg7_1;
	wire w_dff_B_RfcIotNc5_1;
	wire w_dff_B_11nXivdv5_1;
	wire w_dff_B_p8GAccRn6_1;
	wire w_dff_B_NKa6mCVm3_1;
	wire w_dff_B_qKm0c2PR6_1;
	wire w_dff_B_QqTC3GqG1_1;
	wire w_dff_B_d67I1yEw2_1;
	wire w_dff_B_Yvz8a1Zj4_1;
	wire w_dff_B_DTmqrhI77_1;
	wire w_dff_B_YTMw8jbj6_1;
	wire w_dff_B_ntFNMbjf3_1;
	wire w_dff_B_G2p7C0LJ4_1;
	wire w_dff_B_kkYTFtPX6_1;
	wire w_dff_B_nyE2hOSS6_1;
	wire w_dff_B_fFWDEjXN2_1;
	wire w_dff_B_H7D2VEHU0_1;
	wire w_dff_B_zyLsYVRs4_1;
	wire w_dff_B_ZPxGnCnY7_1;
	wire w_dff_B_W0U7m01G1_1;
	wire w_dff_B_PUzwXvxc8_1;
	wire w_dff_B_6PVqFGWO6_1;
	wire w_dff_B_DIuDIFah8_1;
	wire w_dff_B_f3Wh9rEy8_1;
	wire w_dff_B_ouW4klhi7_1;
	wire w_dff_B_5JJMuoK85_1;
	wire w_dff_B_5xbvey3D3_1;
	wire w_dff_B_DqZ3krW32_1;
	wire w_dff_B_uLIT2wYr9_1;
	wire w_dff_B_CdufCjmh8_1;
	wire w_dff_B_MLhHLfZ69_1;
	wire w_dff_B_qRRscppg1_1;
	wire w_dff_B_lu0jKwhg7_0;
	wire w_dff_B_LMG6sXCp5_0;
	wire w_dff_B_jQimGCcU4_0;
	wire w_dff_B_UGbJwrK80_0;
	wire w_dff_B_JbfWrsew3_0;
	wire w_dff_B_vvLnYKPt0_0;
	wire w_dff_B_SX9cjsYO7_0;
	wire w_dff_B_a7zfLXLZ1_0;
	wire w_dff_B_0RKhL6QD0_0;
	wire w_dff_B_PYQyE1yt0_0;
	wire w_dff_B_TjxINM5T6_0;
	wire w_dff_B_LaGT85EI4_0;
	wire w_dff_B_98401wJs5_0;
	wire w_dff_B_7H3l43WF2_0;
	wire w_dff_B_KkNAJwhW1_0;
	wire w_dff_B_kMbZVk0N2_0;
	wire w_dff_B_uhlipbo12_0;
	wire w_dff_B_eU1ZMQl38_0;
	wire w_dff_B_FYgBgGkM1_0;
	wire w_dff_B_tdaCUUCh3_0;
	wire w_dff_B_zjaA3UCz9_0;
	wire w_dff_B_j9zhAkxk0_0;
	wire w_dff_B_bjGQrSQw3_0;
	wire w_dff_B_zKR3BpMY3_0;
	wire w_dff_B_Fsv1XcOM9_0;
	wire w_dff_B_eP80DWHN1_0;
	wire w_dff_B_uMTO6AbD9_0;
	wire w_dff_B_LqzZ19jE2_0;
	wire w_dff_B_FoXkDSWr9_0;
	wire w_dff_B_ewDUfnrO5_0;
	wire w_dff_B_bYYMEXXA5_0;
	wire w_dff_B_swqyUwyx9_0;
	wire w_dff_B_4L96TeJJ7_0;
	wire w_dff_B_XowcDu7J3_0;
	wire w_dff_B_ZdD6P1kc7_0;
	wire w_dff_B_n4T3GGwq1_0;
	wire w_dff_B_Q1ZtM9W36_0;
	wire w_dff_B_yD4ZP8Ky7_0;
	wire w_dff_B_JFMKQI0n4_0;
	wire w_dff_B_BXXTbmW67_0;
	wire w_dff_B_9OzdXUnA5_0;
	wire w_dff_B_6ClUdtnQ0_0;
	wire w_dff_B_8AQy0azS0_0;
	wire w_dff_B_yYGzIpmp6_0;
	wire w_dff_B_eIOcBpCL5_0;
	wire w_dff_B_soHxIGkn1_0;
	wire w_dff_B_Zj7Agyuo8_0;
	wire w_dff_B_GUERlje50_0;
	wire w_dff_B_bLc4jksm0_0;
	wire w_dff_B_DHPiFWKz8_0;
	wire w_dff_B_V8YMXhhG4_0;
	wire w_dff_B_0tOAmo6v5_0;
	wire w_dff_B_mXHFyDR38_0;
	wire w_dff_B_3DUEDxSV2_0;
	wire w_dff_B_CFDZZqPX4_0;
	wire w_dff_B_iUZnEXYf3_0;
	wire w_dff_B_6XQagl4x4_0;
	wire w_dff_B_045SAdZ08_0;
	wire w_dff_B_6iOHQxq56_0;
	wire w_dff_B_ZlnGgaU10_0;
	wire w_dff_B_7SNsgknd4_0;
	wire w_dff_B_UkjGFXeC6_0;
	wire w_dff_B_ZM99NR263_0;
	wire w_dff_B_giyBhSGG8_0;
	wire w_dff_B_bC88Rmr72_0;
	wire w_dff_B_BFiisW189_0;
	wire w_dff_B_6e7R4Sh14_0;
	wire w_dff_B_WbJF2mNq0_0;
	wire w_dff_B_Pd1XC5Qu7_0;
	wire w_dff_B_eyJLCFYt9_0;
	wire w_dff_B_FKDsgxv23_0;
	wire w_dff_B_n4YjFBQ69_0;
	wire w_dff_B_qbF6fOU16_0;
	wire w_dff_B_tcBIdS1F9_0;
	wire w_dff_B_5yv60ErV3_0;
	wire w_dff_B_PV6UTCN74_0;
	wire w_dff_B_DN0IvlKQ2_0;
	wire w_dff_B_4JQHIIHQ9_0;
	wire w_dff_B_VlFtOg230_0;
	wire w_dff_B_iRaeLmCR6_0;
	wire w_dff_B_pS5Sx5fS8_0;
	wire w_dff_B_LHsiC0Jf1_0;
	wire w_dff_B_5madsnMo3_0;
	wire w_dff_B_208MumJ28_0;
	wire w_dff_B_XvplUUQN7_0;
	wire w_dff_B_d2zxyvRn8_0;
	wire w_dff_B_Vs4X5a7l1_0;
	wire w_dff_B_dEEZRkyX6_0;
	wire w_dff_B_5OC06DAu9_0;
	wire w_dff_B_RAmAeZvY4_0;
	wire w_dff_B_gBxUcg4g0_0;
	wire w_dff_B_ikZRNFc48_0;
	wire w_dff_B_Z53VFgFh4_0;
	wire w_dff_B_gJdq2iFW4_1;
	wire w_dff_B_kxp8UXUu7_1;
	wire w_dff_B_Y8AS3hzT7_1;
	wire w_dff_B_rYUKApbL1_1;
	wire w_dff_B_1D6fcqmm4_1;
	wire w_dff_B_XTDzDp7s6_1;
	wire w_dff_B_o8HThdOc9_1;
	wire w_dff_B_BVLnBUKQ7_1;
	wire w_dff_B_Q72bFlLb5_1;
	wire w_dff_B_7w8HJnUw1_1;
	wire w_dff_B_Earm1Lbh5_1;
	wire w_dff_B_AQCtyrYs0_1;
	wire w_dff_B_XLPQlUWJ3_1;
	wire w_dff_B_a40VwrMN9_1;
	wire w_dff_B_OXHbIwbY8_1;
	wire w_dff_B_nClTPOUA0_1;
	wire w_dff_B_x0WGYBFI3_1;
	wire w_dff_B_l0Mk3j9i2_1;
	wire w_dff_B_oTfozGIW0_1;
	wire w_dff_B_WWOZ8LHr2_1;
	wire w_dff_B_z7ZTOhm55_1;
	wire w_dff_B_yQOybGYQ3_1;
	wire w_dff_B_AkQFHqJJ2_1;
	wire w_dff_B_nN68PjVC6_1;
	wire w_dff_B_2kpzQNDz3_1;
	wire w_dff_B_Juay2Nov4_1;
	wire w_dff_B_FXvrNmQ59_1;
	wire w_dff_B_VBUE0oDI6_1;
	wire w_dff_B_fqREJ3yI4_1;
	wire w_dff_B_p4o6w6TL1_1;
	wire w_dff_B_umbdZvZk2_1;
	wire w_dff_B_T0G0K86w9_1;
	wire w_dff_B_gjYt8e504_1;
	wire w_dff_B_WxshiquB5_1;
	wire w_dff_B_pvL3FjqO3_1;
	wire w_dff_B_Oo9lCkc38_1;
	wire w_dff_B_LqZkMe9J7_1;
	wire w_dff_B_bdmcPQ3E0_1;
	wire w_dff_B_UKYfU18j8_1;
	wire w_dff_B_xgvNeYYX7_1;
	wire w_dff_B_pf5bLrZd2_1;
	wire w_dff_B_2qVzltxa0_1;
	wire w_dff_B_iXjBJbqQ0_1;
	wire w_dff_B_GQOHcUtf8_1;
	wire w_dff_B_G6aCvdQ98_1;
	wire w_dff_B_VQFU9dlP5_1;
	wire w_dff_B_HGr7RPbD3_1;
	wire w_dff_B_dDCKUA7p7_1;
	wire w_dff_B_Q4Trv6Kx3_1;
	wire w_dff_B_Ky9FZmxw7_1;
	wire w_dff_B_kp9m1rdh1_1;
	wire w_dff_B_dNsFh5629_1;
	wire w_dff_B_CMXQOyfh5_1;
	wire w_dff_B_g0dV1RIx1_1;
	wire w_dff_B_SLZO7cTh8_1;
	wire w_dff_B_v30Q16nc3_1;
	wire w_dff_B_sFRDUQyu4_1;
	wire w_dff_B_c3qqaAIE7_1;
	wire w_dff_B_1Z84bdlj8_1;
	wire w_dff_B_HeBMupr65_1;
	wire w_dff_B_ZtZW9Vkp9_1;
	wire w_dff_B_bTWyxHBG4_1;
	wire w_dff_B_JSjapsW71_1;
	wire w_dff_B_modIlHbJ9_1;
	wire w_dff_B_ju0FS38I7_1;
	wire w_dff_B_SR7yMiT46_1;
	wire w_dff_B_qPlGZ4Op4_1;
	wire w_dff_B_zgHESNBO2_1;
	wire w_dff_B_6MyFkASg8_1;
	wire w_dff_B_1jpzhTsR7_1;
	wire w_dff_B_f17KTT2q2_1;
	wire w_dff_B_thw9dMyV7_1;
	wire w_dff_B_7tDgPT6H2_1;
	wire w_dff_B_XM37YRli8_1;
	wire w_dff_B_AL8Jhazv9_1;
	wire w_dff_B_aHVoLH9V4_1;
	wire w_dff_B_PCRJhqxl5_1;
	wire w_dff_B_6Zi3mZRg6_1;
	wire w_dff_B_5p6VndcG9_1;
	wire w_dff_B_hK8IBF6Z7_1;
	wire w_dff_B_xBgQUeLM5_1;
	wire w_dff_B_pUYlLAwu1_1;
	wire w_dff_B_riFVKxaT3_1;
	wire w_dff_B_CAxX5keN2_1;
	wire w_dff_B_hT9uO1Sj6_1;
	wire w_dff_B_2XG7dEL79_1;
	wire w_dff_B_aRJdYECd0_1;
	wire w_dff_B_Q8vzqKRK2_1;
	wire w_dff_B_NJXi8wR85_1;
	wire w_dff_B_HmwWwxAw6_1;
	wire w_dff_B_ATTpfHUD2_1;
	wire w_dff_B_Vnmk2IHa8_1;
	wire w_dff_B_lM2dOOfg6_0;
	wire w_dff_B_UVBbWmA94_0;
	wire w_dff_B_O5EZFslc0_0;
	wire w_dff_B_wpQvMyOr8_0;
	wire w_dff_B_ffZKLTDW9_0;
	wire w_dff_B_AtwWn1ak4_0;
	wire w_dff_B_JFXGJ8Q57_0;
	wire w_dff_B_cM0XTWPi0_0;
	wire w_dff_B_gBbmHKQx9_0;
	wire w_dff_B_8wkIgPVT6_0;
	wire w_dff_B_7IbJrvUK8_0;
	wire w_dff_B_ZFjcT3Mm6_0;
	wire w_dff_B_vyqccrap3_0;
	wire w_dff_B_wBEh1cYs8_0;
	wire w_dff_B_LEvP48ZI4_0;
	wire w_dff_B_O7o0v4391_0;
	wire w_dff_B_Vu0dGa9d7_0;
	wire w_dff_B_ScmTPTjs2_0;
	wire w_dff_B_CSPiqqkT7_0;
	wire w_dff_B_DAvgV9gY4_0;
	wire w_dff_B_dbwZnmVb1_0;
	wire w_dff_B_b4oSywtt6_0;
	wire w_dff_B_heADqEni1_0;
	wire w_dff_B_jaJEzduF5_0;
	wire w_dff_B_ZI4LEGYH2_0;
	wire w_dff_B_yYDFQRsZ7_0;
	wire w_dff_B_goIIgDJs7_0;
	wire w_dff_B_wydOFzRy6_0;
	wire w_dff_B_eWJ5OrwX9_0;
	wire w_dff_B_dg6eiWIh2_0;
	wire w_dff_B_WOH5FebT2_0;
	wire w_dff_B_SuOwa5ZY2_0;
	wire w_dff_B_ztuftAGP7_0;
	wire w_dff_B_jWwmd1iH4_0;
	wire w_dff_B_qrkXPVzr1_0;
	wire w_dff_B_NeygJGxY4_0;
	wire w_dff_B_5mlTtPy62_0;
	wire w_dff_B_SgFXI4tH1_0;
	wire w_dff_B_9xBA2FgC8_0;
	wire w_dff_B_Pn8DZBJI7_0;
	wire w_dff_B_6BNrlVVG6_0;
	wire w_dff_B_mSbK4Cra5_0;
	wire w_dff_B_DTSA04BY1_0;
	wire w_dff_B_BB6gZxnl4_0;
	wire w_dff_B_mU06QV8i2_0;
	wire w_dff_B_ZZPsf6WI2_0;
	wire w_dff_B_e1xU3K620_0;
	wire w_dff_B_vsYwFBOP4_0;
	wire w_dff_B_AQzJivG39_0;
	wire w_dff_B_B26oeoLo6_0;
	wire w_dff_B_TLcpQ3IQ1_0;
	wire w_dff_B_MGPMoaRv0_0;
	wire w_dff_B_wuhFgHP11_0;
	wire w_dff_B_vYUpdkdO0_0;
	wire w_dff_B_sbK29lDI3_0;
	wire w_dff_B_GH1p1qcc2_0;
	wire w_dff_B_SNATx7hZ5_0;
	wire w_dff_B_Sx5BBdHK2_0;
	wire w_dff_B_uKMBZZ7b1_0;
	wire w_dff_B_B2AAVMVs9_0;
	wire w_dff_B_T3LNFtu92_0;
	wire w_dff_B_x2ILHnnz5_0;
	wire w_dff_B_x9qszdhL8_0;
	wire w_dff_B_UftfQlIV1_0;
	wire w_dff_B_vz3zVUZd8_0;
	wire w_dff_B_fmk6QcDA9_0;
	wire w_dff_B_cJOc17Dj2_0;
	wire w_dff_B_lzFljsCR2_0;
	wire w_dff_B_PtfeqFIx3_0;
	wire w_dff_B_yep4vL4G0_0;
	wire w_dff_B_NheNfkYk8_0;
	wire w_dff_B_UebbZUQr0_0;
	wire w_dff_B_br2B6fth1_0;
	wire w_dff_B_syA4iOfo1_0;
	wire w_dff_B_QJiujBaq8_0;
	wire w_dff_B_2FUlOjPf6_0;
	wire w_dff_B_VBqk8ThL3_0;
	wire w_dff_B_TncV616K6_0;
	wire w_dff_B_c5JrsnKV6_0;
	wire w_dff_B_RbbPDLYO1_0;
	wire w_dff_B_kOGm8zEs9_0;
	wire w_dff_B_KBgZBmGc5_0;
	wire w_dff_B_ZtxR5PI36_0;
	wire w_dff_B_l6ocIsuX2_0;
	wire w_dff_B_eMlvmWyc5_0;
	wire w_dff_B_waAhaXlM4_0;
	wire w_dff_B_yIo0sQNo8_0;
	wire w_dff_B_Tjg5JjoQ5_0;
	wire w_dff_B_c3Num61Z6_0;
	wire w_dff_B_RiUHyLMr8_0;
	wire w_dff_B_t57R8BJk5_0;
	wire w_dff_B_2tpIruTy5_0;
	wire w_dff_B_ZQKKpnKS0_1;
	wire w_dff_B_hyvVoXDq5_1;
	wire w_dff_B_2rlWrmKE8_1;
	wire w_dff_B_b77XAnMR0_1;
	wire w_dff_B_XTx48BFZ6_1;
	wire w_dff_B_qdXgJKKH5_1;
	wire w_dff_B_OeO1Wmeq0_1;
	wire w_dff_B_TZxNTdXT0_1;
	wire w_dff_B_i6woalFV3_1;
	wire w_dff_B_WQiHXRey7_1;
	wire w_dff_B_eKpshZld5_1;
	wire w_dff_B_rBhIkbGK4_1;
	wire w_dff_B_5AcocSIw2_1;
	wire w_dff_B_upL5tNg77_1;
	wire w_dff_B_hAwyS8Ed9_1;
	wire w_dff_B_hMCqLxTx9_1;
	wire w_dff_B_ABREldef9_1;
	wire w_dff_B_Za16KxHz1_1;
	wire w_dff_B_g9BEGyV38_1;
	wire w_dff_B_q2dsZIkH5_1;
	wire w_dff_B_HCkqZFVx7_1;
	wire w_dff_B_wuh39z5h0_1;
	wire w_dff_B_KZVJ1Uil1_1;
	wire w_dff_B_BWpVNCCC2_1;
	wire w_dff_B_DKdYYBA96_1;
	wire w_dff_B_qwEHv9v82_1;
	wire w_dff_B_kTqFJaj26_1;
	wire w_dff_B_NOLA7Ut27_1;
	wire w_dff_B_fsJEECv94_1;
	wire w_dff_B_LuYGpeAY1_1;
	wire w_dff_B_le184tYM0_1;
	wire w_dff_B_T9eTpHAR9_1;
	wire w_dff_B_uH14Dbid2_1;
	wire w_dff_B_2Lkym8bN9_1;
	wire w_dff_B_a9kFii4x0_1;
	wire w_dff_B_lmmnAsfP6_1;
	wire w_dff_B_EnxXsfQC6_1;
	wire w_dff_B_RVIrtoho8_1;
	wire w_dff_B_V8mjDS7W3_1;
	wire w_dff_B_jnQNt3aD2_1;
	wire w_dff_B_7gg0bx6b0_1;
	wire w_dff_B_JY0KhHLO8_1;
	wire w_dff_B_iLXZ0D6q2_1;
	wire w_dff_B_FsLwiPBW3_1;
	wire w_dff_B_loGaXOrq4_1;
	wire w_dff_B_5aBw9nLi5_1;
	wire w_dff_B_mZpK3axG0_1;
	wire w_dff_B_XyRs4s4z3_1;
	wire w_dff_B_ACmCXSDy4_1;
	wire w_dff_B_GJh7p58r5_1;
	wire w_dff_B_2frT5aZ90_1;
	wire w_dff_B_KzN9yxYq6_1;
	wire w_dff_B_AJZCYnvk9_1;
	wire w_dff_B_DbsOHvFM7_1;
	wire w_dff_B_BP6jGezL7_1;
	wire w_dff_B_VamXzUl30_1;
	wire w_dff_B_AWRB28MV2_1;
	wire w_dff_B_5AjSqHfD8_1;
	wire w_dff_B_9dV47HvI6_1;
	wire w_dff_B_bOBWRJGc1_1;
	wire w_dff_B_Mvp7oTsm1_1;
	wire w_dff_B_bZJSGiR79_1;
	wire w_dff_B_Pfl3HMCX3_1;
	wire w_dff_B_UiKAMvgk0_1;
	wire w_dff_B_dIa7nWvw1_1;
	wire w_dff_B_IG3ckOWe8_1;
	wire w_dff_B_8nE5qFnE0_1;
	wire w_dff_B_HL2xPlH74_1;
	wire w_dff_B_mcEoyKTN6_1;
	wire w_dff_B_oXFS6tjS9_1;
	wire w_dff_B_3Mi9Gsdu5_1;
	wire w_dff_B_ELejFTVp7_1;
	wire w_dff_B_sn5Wp6Fr4_1;
	wire w_dff_B_j8SCVz7e6_1;
	wire w_dff_B_VUiFq6jH9_1;
	wire w_dff_B_IxpQ1gpW4_1;
	wire w_dff_B_MP9moO1H6_1;
	wire w_dff_B_CMYRLp6X7_1;
	wire w_dff_B_uNurphcp6_1;
	wire w_dff_B_XktcUBUX7_1;
	wire w_dff_B_iN8WgXyO6_1;
	wire w_dff_B_3XjSxaxE6_1;
	wire w_dff_B_MlD79jp26_1;
	wire w_dff_B_bA6E01ro1_1;
	wire w_dff_B_J5bPjCEh8_1;
	wire w_dff_B_PKpGVWci4_1;
	wire w_dff_B_b4Yyg7Wb8_1;
	wire w_dff_B_y35aUNqV9_1;
	wire w_dff_B_8Kymw5863_1;
	wire w_dff_B_YvcDHCUq5_1;
	wire w_dff_B_eoY4eUdu5_1;
	wire w_dff_B_r6oiuFx05_0;
	wire w_dff_B_2bawyn1r8_0;
	wire w_dff_B_ziqfpptT1_0;
	wire w_dff_B_37JprzNU9_0;
	wire w_dff_B_akUv6lz74_0;
	wire w_dff_B_OGMDRS3F7_0;
	wire w_dff_B_UnjYyCk78_0;
	wire w_dff_B_nhdnsPRK0_0;
	wire w_dff_B_HQE5uNHq0_0;
	wire w_dff_B_HHmdn0UE9_0;
	wire w_dff_B_V6tFQHXl8_0;
	wire w_dff_B_nXVvsL5x3_0;
	wire w_dff_B_1wvDl6qs8_0;
	wire w_dff_B_ravbEzCR9_0;
	wire w_dff_B_8KhRWNQ71_0;
	wire w_dff_B_cyzAh48f6_0;
	wire w_dff_B_s5e8FSEN1_0;
	wire w_dff_B_mK1nylq38_0;
	wire w_dff_B_Um5pdJSm4_0;
	wire w_dff_B_oZzS8cBA7_0;
	wire w_dff_B_Rsw4HFE22_0;
	wire w_dff_B_FUtx1SPN0_0;
	wire w_dff_B_FJrcUHrM5_0;
	wire w_dff_B_qVH48R986_0;
	wire w_dff_B_VKbE30s90_0;
	wire w_dff_B_otbRIaFe2_0;
	wire w_dff_B_oSXLY6E07_0;
	wire w_dff_B_XEENkSAO6_0;
	wire w_dff_B_9avH78Dr5_0;
	wire w_dff_B_SwwZKrUg8_0;
	wire w_dff_B_Dzixfz0g7_0;
	wire w_dff_B_jYBkZqFp1_0;
	wire w_dff_B_DHIPo0I45_0;
	wire w_dff_B_wx8zFKNI8_0;
	wire w_dff_B_PmlhirSB8_0;
	wire w_dff_B_6RWenhc93_0;
	wire w_dff_B_mzqpiX8W6_0;
	wire w_dff_B_PjwitYUW4_0;
	wire w_dff_B_nYfbVR5P4_0;
	wire w_dff_B_ud0NlXKT4_0;
	wire w_dff_B_hR6qfRFe9_0;
	wire w_dff_B_ojaHAo0n5_0;
	wire w_dff_B_iIXUgi9K5_0;
	wire w_dff_B_RQfKjI439_0;
	wire w_dff_B_a8ZPmP1q9_0;
	wire w_dff_B_7zFFgnua2_0;
	wire w_dff_B_7gxoReoM7_0;
	wire w_dff_B_8cXdFcyZ5_0;
	wire w_dff_B_oaQ0FsZ10_0;
	wire w_dff_B_oZvnS2510_0;
	wire w_dff_B_EXC8SVu56_0;
	wire w_dff_B_2PcolzLq4_0;
	wire w_dff_B_LDhGuWmx4_0;
	wire w_dff_B_M4qapaot3_0;
	wire w_dff_B_pCRKaWQa6_0;
	wire w_dff_B_QD9euuLG9_0;
	wire w_dff_B_a88WwJJP7_0;
	wire w_dff_B_9iyKrfid3_0;
	wire w_dff_B_4HyRwzR37_0;
	wire w_dff_B_EaD88TUA8_0;
	wire w_dff_B_r4dh04yK0_0;
	wire w_dff_B_wqR3NJMA7_0;
	wire w_dff_B_Qnjbbc5T4_0;
	wire w_dff_B_C0f42nzF8_0;
	wire w_dff_B_lo9QwvLM4_0;
	wire w_dff_B_vTH0mWKG9_0;
	wire w_dff_B_Kt6wot8k7_0;
	wire w_dff_B_epyffjIx6_0;
	wire w_dff_B_wm3QBzfu2_0;
	wire w_dff_B_umGt7O0q9_0;
	wire w_dff_B_UngqZoyv3_0;
	wire w_dff_B_l87SoIcI6_0;
	wire w_dff_B_oVjMHjQe7_0;
	wire w_dff_B_63sWTRei1_0;
	wire w_dff_B_SkGqrsQ32_0;
	wire w_dff_B_1f1zlaui2_0;
	wire w_dff_B_VhcQO4xz5_0;
	wire w_dff_B_XpQCptHj0_0;
	wire w_dff_B_UCouXUMV6_0;
	wire w_dff_B_dpDwdH1y6_0;
	wire w_dff_B_nOwIypRd1_0;
	wire w_dff_B_2ACqmBer0_0;
	wire w_dff_B_sLkbvnto5_0;
	wire w_dff_B_0fb6EK129_0;
	wire w_dff_B_LJfbNuao1_0;
	wire w_dff_B_QaEH5rye9_0;
	wire w_dff_B_aldOUR2M3_0;
	wire w_dff_B_E5Shiag94_0;
	wire w_dff_B_iHxN2qeg1_0;
	wire w_dff_B_uiXlNlYP1_0;
	wire w_dff_B_yQ9eGirj0_0;
	wire w_dff_B_se6uw62Z3_1;
	wire w_dff_B_YDFTS4SQ8_1;
	wire w_dff_B_cpUYpy5L2_1;
	wire w_dff_B_At484BH01_1;
	wire w_dff_B_TwSipUUb6_1;
	wire w_dff_B_442PVjyk4_1;
	wire w_dff_B_VeLr0Mw59_1;
	wire w_dff_B_LxYosw3b0_1;
	wire w_dff_B_fiyfH08J3_1;
	wire w_dff_B_pg9ajxEX1_1;
	wire w_dff_B_BHOL2XNv4_1;
	wire w_dff_B_Dnw9AESR8_1;
	wire w_dff_B_vuaxBBiN0_1;
	wire w_dff_B_fm1ljZqU0_1;
	wire w_dff_B_Pi1MUNvl8_1;
	wire w_dff_B_xiWacX7r8_1;
	wire w_dff_B_ZmshhO0M4_1;
	wire w_dff_B_2RM2zhVA6_1;
	wire w_dff_B_aadhiS0u7_1;
	wire w_dff_B_ODs7ZHdc9_1;
	wire w_dff_B_uuTht2yX7_1;
	wire w_dff_B_8PNwltkp0_1;
	wire w_dff_B_UagfwMXB8_1;
	wire w_dff_B_N9UWKVbL3_1;
	wire w_dff_B_UenmgPv27_1;
	wire w_dff_B_l8eCAZ7q8_1;
	wire w_dff_B_e4SZfojh6_1;
	wire w_dff_B_MahyBmm61_1;
	wire w_dff_B_poG3bfMf7_1;
	wire w_dff_B_hXyV80Eh8_1;
	wire w_dff_B_96Y8Y0Xn7_1;
	wire w_dff_B_u8LgfXdD4_1;
	wire w_dff_B_YZrnAZso7_1;
	wire w_dff_B_6q36HsiP7_1;
	wire w_dff_B_gfBpOPU05_1;
	wire w_dff_B_ayQVFRgc6_1;
	wire w_dff_B_D7Bq0hXG9_1;
	wire w_dff_B_RAqRx4YC3_1;
	wire w_dff_B_rrTAiO973_1;
	wire w_dff_B_PdmRQyhx4_1;
	wire w_dff_B_jlTdkK9s5_1;
	wire w_dff_B_q6r7xMLt3_1;
	wire w_dff_B_v7cnN4s29_1;
	wire w_dff_B_SX529mAj1_1;
	wire w_dff_B_girElLVg7_1;
	wire w_dff_B_4016CAJ11_1;
	wire w_dff_B_cMLBt9kp1_1;
	wire w_dff_B_uLTtgTGu2_1;
	wire w_dff_B_zF8Wz0fX8_1;
	wire w_dff_B_DzR02vbf7_1;
	wire w_dff_B_EsGhCumm9_1;
	wire w_dff_B_tyTJrobg6_1;
	wire w_dff_B_xZ1dsy4Y4_1;
	wire w_dff_B_0rzug1X50_1;
	wire w_dff_B_9yUdXD7Q0_1;
	wire w_dff_B_P6ZBZUna8_1;
	wire w_dff_B_ehxFBoAy6_1;
	wire w_dff_B_O6uoHPkp0_1;
	wire w_dff_B_KXCWaXlA1_1;
	wire w_dff_B_h5SArAYA8_1;
	wire w_dff_B_67xymoO71_1;
	wire w_dff_B_fhEPmXiH3_1;
	wire w_dff_B_dTsEZXC33_1;
	wire w_dff_B_yogbt60R8_1;
	wire w_dff_B_9EkWQFFq8_1;
	wire w_dff_B_gAaNQ4jQ3_1;
	wire w_dff_B_Ab1nIuMG4_1;
	wire w_dff_B_xfIxl0zk7_1;
	wire w_dff_B_T7EngNF43_1;
	wire w_dff_B_Z4x5vGIF6_1;
	wire w_dff_B_mSYnoF7c0_1;
	wire w_dff_B_eMqWX1mv4_1;
	wire w_dff_B_2j8yGB2t7_1;
	wire w_dff_B_oBGuM9CJ9_1;
	wire w_dff_B_xjNVOoN11_1;
	wire w_dff_B_V0t9D08C8_1;
	wire w_dff_B_u67vymPe9_1;
	wire w_dff_B_uEGT0HKF9_1;
	wire w_dff_B_bwbXM5zf9_1;
	wire w_dff_B_vPk5cKqa5_1;
	wire w_dff_B_ENDknJRO4_1;
	wire w_dff_B_AoiiewfB8_1;
	wire w_dff_B_aXE0BQV53_1;
	wire w_dff_B_rhDmmGVz7_1;
	wire w_dff_B_9Ny2l7y05_1;
	wire w_dff_B_MR3g1Rmd9_1;
	wire w_dff_B_GJxbffZN1_1;
	wire w_dff_B_VrVeXKav6_1;
	wire w_dff_B_QhDgwt0p3_1;
	wire w_dff_B_8T9xx6qV1_1;
	wire w_dff_B_9TIwEGfL8_0;
	wire w_dff_B_sIteoKyL8_0;
	wire w_dff_B_00Epb6yB9_0;
	wire w_dff_B_tk6ZurhK2_0;
	wire w_dff_B_TDPGJW6W9_0;
	wire w_dff_B_r0bZlsZ27_0;
	wire w_dff_B_P55q99eh7_0;
	wire w_dff_B_qOMxUOQB0_0;
	wire w_dff_B_GA7N7gGi1_0;
	wire w_dff_B_KM0OfOSB7_0;
	wire w_dff_B_63mw0JeE4_0;
	wire w_dff_B_CeIS1ebV3_0;
	wire w_dff_B_ZuLkiFml4_0;
	wire w_dff_B_CUCnWHdZ8_0;
	wire w_dff_B_UImQlz6O0_0;
	wire w_dff_B_RnKs8BBT4_0;
	wire w_dff_B_XrGY9wZF1_0;
	wire w_dff_B_D7Gg0IyA5_0;
	wire w_dff_B_RyOQ2TAX1_0;
	wire w_dff_B_Ud0Mwmln4_0;
	wire w_dff_B_Qi56saku0_0;
	wire w_dff_B_dM2qqaU35_0;
	wire w_dff_B_cW5EmClX9_0;
	wire w_dff_B_jn3TTuLa2_0;
	wire w_dff_B_ME6W3FR53_0;
	wire w_dff_B_fGtxDOeT3_0;
	wire w_dff_B_Yl4aPK3S6_0;
	wire w_dff_B_LQGJATPE7_0;
	wire w_dff_B_zgYswCqo8_0;
	wire w_dff_B_qJVr2lAM9_0;
	wire w_dff_B_iKbkbYNq5_0;
	wire w_dff_B_wbbMIOMZ0_0;
	wire w_dff_B_qK2JSXFx0_0;
	wire w_dff_B_0ENvKeQX2_0;
	wire w_dff_B_2nv5Y9tz5_0;
	wire w_dff_B_NwWtRiby8_0;
	wire w_dff_B_8f9lUmVY2_0;
	wire w_dff_B_MOJaemYw3_0;
	wire w_dff_B_ubiPk2dv7_0;
	wire w_dff_B_4Ah5fmIz1_0;
	wire w_dff_B_eo5i8lER0_0;
	wire w_dff_B_fSBLeV4Y6_0;
	wire w_dff_B_8FG9T9k87_0;
	wire w_dff_B_RLiXS2969_0;
	wire w_dff_B_MnNLDbuF8_0;
	wire w_dff_B_oKEFgqO73_0;
	wire w_dff_B_cbwPiUJS3_0;
	wire w_dff_B_1eid7WdF0_0;
	wire w_dff_B_CytOpRm93_0;
	wire w_dff_B_A5aCXa3M9_0;
	wire w_dff_B_Sr9ARhcy1_0;
	wire w_dff_B_O2MXcG8D1_0;
	wire w_dff_B_fw0AaPIr8_0;
	wire w_dff_B_8DxRkOeI1_0;
	wire w_dff_B_ChaCEjcx6_0;
	wire w_dff_B_LE7h1kVx6_0;
	wire w_dff_B_SR7lmSk17_0;
	wire w_dff_B_upYOXlrG2_0;
	wire w_dff_B_ETyYKwbI8_0;
	wire w_dff_B_A3JkxCNg8_0;
	wire w_dff_B_3sgCRIyf1_0;
	wire w_dff_B_SjXgULOd1_0;
	wire w_dff_B_Mqk47ZQl3_0;
	wire w_dff_B_39aR6EaX5_0;
	wire w_dff_B_ZNXax4Ux1_0;
	wire w_dff_B_lL0rgrqc6_0;
	wire w_dff_B_zWHxyE0u6_0;
	wire w_dff_B_azEX5QrN2_0;
	wire w_dff_B_39Hqd9fk9_0;
	wire w_dff_B_cYGe8lOB3_0;
	wire w_dff_B_XzuFU1fd3_0;
	wire w_dff_B_GVEkaWq78_0;
	wire w_dff_B_SPYaZBIt9_0;
	wire w_dff_B_IKK8GyuH4_0;
	wire w_dff_B_WPAHE3mh3_0;
	wire w_dff_B_nIdPCuCc6_0;
	wire w_dff_B_LyL1bnj37_0;
	wire w_dff_B_r3MtVTUV4_0;
	wire w_dff_B_49A45O3U7_0;
	wire w_dff_B_SPYIYyVM1_0;
	wire w_dff_B_3ITYnHvH3_0;
	wire w_dff_B_JIjQ7XFx8_0;
	wire w_dff_B_xJ5r5Fbi2_0;
	wire w_dff_B_uVjbqEq83_0;
	wire w_dff_B_tDjI2Xgg9_0;
	wire w_dff_B_PDwlWK5J4_0;
	wire w_dff_B_jxrQ0aod0_0;
	wire w_dff_B_zzWVvkcD6_0;
	wire w_dff_B_dh0e9h5F0_0;
	wire w_dff_B_wsbERzgk2_0;
	wire w_dff_B_rKDKmjhn1_1;
	wire w_dff_B_er6DPLDV9_1;
	wire w_dff_B_ODFTmzQx6_1;
	wire w_dff_B_cdw8X4H16_1;
	wire w_dff_B_mD0hgiOU4_1;
	wire w_dff_B_XLPWQ5T59_1;
	wire w_dff_B_mHQpz9YE1_1;
	wire w_dff_B_KyEJI5Bt8_1;
	wire w_dff_B_wq03rv2k6_1;
	wire w_dff_B_aiNAYzaR4_1;
	wire w_dff_B_bx2HPkwq1_1;
	wire w_dff_B_6zDt640a2_1;
	wire w_dff_B_XxjHxdxX5_1;
	wire w_dff_B_XxhCUhdQ1_1;
	wire w_dff_B_Zc7zOHuv6_1;
	wire w_dff_B_o8Akz7Mt5_1;
	wire w_dff_B_QEHvMTz34_1;
	wire w_dff_B_JsxK5gxm1_1;
	wire w_dff_B_CQRFALly7_1;
	wire w_dff_B_Uf6KxqXy3_1;
	wire w_dff_B_nl9xqzwR2_1;
	wire w_dff_B_jPPhEZsJ2_1;
	wire w_dff_B_FiU7s8qO1_1;
	wire w_dff_B_kNypXD1Q4_1;
	wire w_dff_B_0RkdU8Dk8_1;
	wire w_dff_B_EZSTBJhw7_1;
	wire w_dff_B_tsV3vvCx4_1;
	wire w_dff_B_zL04EztH8_1;
	wire w_dff_B_bnYS9BIZ0_1;
	wire w_dff_B_0HmWMjm60_1;
	wire w_dff_B_7cLCiQrE9_1;
	wire w_dff_B_a43D8jlE0_1;
	wire w_dff_B_ClCzBaz86_1;
	wire w_dff_B_H59AaPml8_1;
	wire w_dff_B_zGXCVR4D2_1;
	wire w_dff_B_yowb84Xb8_1;
	wire w_dff_B_bkDWcV3o3_1;
	wire w_dff_B_VLrIIkL24_1;
	wire w_dff_B_HuOV8PjD9_1;
	wire w_dff_B_8dftSuwz0_1;
	wire w_dff_B_SSKgH0KB3_1;
	wire w_dff_B_JMRYtb9y7_1;
	wire w_dff_B_NEnxLnDV7_1;
	wire w_dff_B_amkxZG7q1_1;
	wire w_dff_B_3HSDIFXS2_1;
	wire w_dff_B_9wVIedni4_1;
	wire w_dff_B_ZSRuF6jb7_1;
	wire w_dff_B_US6vRUHY0_1;
	wire w_dff_B_RzfUZ08N9_1;
	wire w_dff_B_S7D9ZjUa7_1;
	wire w_dff_B_V1bKtOVA2_1;
	wire w_dff_B_ltlyL98u1_1;
	wire w_dff_B_GiMVxJ3q9_1;
	wire w_dff_B_fKLzQruU2_1;
	wire w_dff_B_IMDbmNky4_1;
	wire w_dff_B_2YRG67FH6_1;
	wire w_dff_B_YM06LLsm5_1;
	wire w_dff_B_3e0Nst5O6_1;
	wire w_dff_B_MBWRp3Ey3_1;
	wire w_dff_B_PLdqrGPO2_1;
	wire w_dff_B_BLqyRjBX1_1;
	wire w_dff_B_DKc8bUBK8_1;
	wire w_dff_B_GAlLQwWb0_1;
	wire w_dff_B_pwXVKTPS2_1;
	wire w_dff_B_2YBe1GuN5_1;
	wire w_dff_B_ieOnnjQB6_1;
	wire w_dff_B_ScSKBDkm6_1;
	wire w_dff_B_tr7FRnQa7_1;
	wire w_dff_B_bWrAbkGA7_1;
	wire w_dff_B_gohdcBDQ3_1;
	wire w_dff_B_Dql4hhBu7_1;
	wire w_dff_B_WVh3pUMT9_1;
	wire w_dff_B_WKXVA4Ld0_1;
	wire w_dff_B_k2AYrc4j4_1;
	wire w_dff_B_AdKJ3Hcc8_1;
	wire w_dff_B_jcSfwrUx9_1;
	wire w_dff_B_csSKlNFX4_1;
	wire w_dff_B_ar2mZ5eW9_1;
	wire w_dff_B_6iVhIGeW4_1;
	wire w_dff_B_404uCMXz1_1;
	wire w_dff_B_kYuYXyIp6_1;
	wire w_dff_B_k7t0G1JG8_1;
	wire w_dff_B_qxFNxcRM7_1;
	wire w_dff_B_FpTQl5Wl9_1;
	wire w_dff_B_flJCG5ug4_1;
	wire w_dff_B_aOkUFpOL7_1;
	wire w_dff_B_OLNO1eLj9_1;
	wire w_dff_B_AVhDbNiO2_1;
	wire w_dff_B_fXOzDmTA4_1;
	wire w_dff_B_CWY8rxXl1_0;
	wire w_dff_B_Ny70iVOY9_0;
	wire w_dff_B_Q9H4HAL91_0;
	wire w_dff_B_30UWpCw58_0;
	wire w_dff_B_omDmp2vB0_0;
	wire w_dff_B_LGRf6koU9_0;
	wire w_dff_B_vwZCHmW48_0;
	wire w_dff_B_af6AY2XI5_0;
	wire w_dff_B_zDJTeMAT6_0;
	wire w_dff_B_oifYlsDu9_0;
	wire w_dff_B_zSKEdXgu0_0;
	wire w_dff_B_FLTnRCvU1_0;
	wire w_dff_B_EWjKqhVF3_0;
	wire w_dff_B_uEblP9m40_0;
	wire w_dff_B_vLSkXsNv3_0;
	wire w_dff_B_0WWw44gL1_0;
	wire w_dff_B_cT684YBL8_0;
	wire w_dff_B_2iu8I3dq9_0;
	wire w_dff_B_n8Z6Ey0N6_0;
	wire w_dff_B_8kuPXEBp8_0;
	wire w_dff_B_n25xiboc3_0;
	wire w_dff_B_DM63jPwM4_0;
	wire w_dff_B_q4Bj0sIl0_0;
	wire w_dff_B_I0hi6NFe2_0;
	wire w_dff_B_EtL3VBlb5_0;
	wire w_dff_B_FSx0JAlp5_0;
	wire w_dff_B_x1PaXvSn0_0;
	wire w_dff_B_rMpptube3_0;
	wire w_dff_B_4LXFm2cM8_0;
	wire w_dff_B_MEdwn9WO6_0;
	wire w_dff_B_YZA7a6bx2_0;
	wire w_dff_B_pGg2c7GD7_0;
	wire w_dff_B_eCMr5V4a0_0;
	wire w_dff_B_3PDhePEA7_0;
	wire w_dff_B_YjJH8gE13_0;
	wire w_dff_B_DtD70DHb6_0;
	wire w_dff_B_JPIFBaPW5_0;
	wire w_dff_B_fC8vDLJp1_0;
	wire w_dff_B_R3uBh1WE3_0;
	wire w_dff_B_xX63uc1T8_0;
	wire w_dff_B_IBGy8Mal3_0;
	wire w_dff_B_CRlFtMDL1_0;
	wire w_dff_B_fhayUEiM1_0;
	wire w_dff_B_CTT2RzvP6_0;
	wire w_dff_B_GNpGWrch2_0;
	wire w_dff_B_79o3CK3J5_0;
	wire w_dff_B_wJccEvqV2_0;
	wire w_dff_B_qZc6Kva81_0;
	wire w_dff_B_58n5S6Og6_0;
	wire w_dff_B_gbbwywZx9_0;
	wire w_dff_B_DBQAm4B07_0;
	wire w_dff_B_M1BI0gGk2_0;
	wire w_dff_B_2qmu4oG88_0;
	wire w_dff_B_FT5BDjny3_0;
	wire w_dff_B_Q9hu3h5h6_0;
	wire w_dff_B_MVyVtx7U7_0;
	wire w_dff_B_ksW94IBm2_0;
	wire w_dff_B_edURTfez4_0;
	wire w_dff_B_moy20kW28_0;
	wire w_dff_B_AES7Vx9z9_0;
	wire w_dff_B_wTLA7ySI6_0;
	wire w_dff_B_KKmk6h587_0;
	wire w_dff_B_mUBHhjhV0_0;
	wire w_dff_B_6t2YTT5n9_0;
	wire w_dff_B_iyju2Npd6_0;
	wire w_dff_B_MbGZNfAM5_0;
	wire w_dff_B_n0UEG5tt1_0;
	wire w_dff_B_gf76WM7O6_0;
	wire w_dff_B_BUsnqW3l9_0;
	wire w_dff_B_O49HHtdK9_0;
	wire w_dff_B_U0LAbCxi3_0;
	wire w_dff_B_tmd08aPY9_0;
	wire w_dff_B_gLwQOAJk1_0;
	wire w_dff_B_ouLHRigy8_0;
	wire w_dff_B_tPkjOYBy4_0;
	wire w_dff_B_vILfiHHU9_0;
	wire w_dff_B_R2PnrNGY4_0;
	wire w_dff_B_FqO1L7OJ6_0;
	wire w_dff_B_wyKOe8zS5_0;
	wire w_dff_B_ufcbxOSq4_0;
	wire w_dff_B_D7GKjPWf6_0;
	wire w_dff_B_sD6exW0m0_0;
	wire w_dff_B_MoMNsD464_0;
	wire w_dff_B_a01Bcux69_0;
	wire w_dff_B_HWHgsry20_0;
	wire w_dff_B_QsNjBccf5_0;
	wire w_dff_B_TgKETz5Q9_0;
	wire w_dff_B_JZOXfO6O4_0;
	wire w_dff_B_AOA64WTK7_0;
	wire w_dff_B_UPtvfWU60_1;
	wire w_dff_B_UuOGWOQp9_1;
	wire w_dff_B_yMt3zrPz8_1;
	wire w_dff_B_8P3Gnk313_1;
	wire w_dff_B_LYUouN115_1;
	wire w_dff_B_h0DfzFCB3_1;
	wire w_dff_B_knu0rVNO2_1;
	wire w_dff_B_CZDWk2PV0_1;
	wire w_dff_B_EA5nR9F51_1;
	wire w_dff_B_duyFeznp0_1;
	wire w_dff_B_TcBiiXrJ3_1;
	wire w_dff_B_uLSGMLcW8_1;
	wire w_dff_B_v0TSw7JI3_1;
	wire w_dff_B_4t17URdi6_1;
	wire w_dff_B_vE3UuXuF7_1;
	wire w_dff_B_R5k7A6RI9_1;
	wire w_dff_B_WlfhKH3U5_1;
	wire w_dff_B_cI3IDdS14_1;
	wire w_dff_B_aeAVzOg09_1;
	wire w_dff_B_cFj5Rkyd6_1;
	wire w_dff_B_qTb8J63n7_1;
	wire w_dff_B_uOx7elwQ2_1;
	wire w_dff_B_JSZ2VZWM4_1;
	wire w_dff_B_F7FYp8q85_1;
	wire w_dff_B_V1ZQmTS75_1;
	wire w_dff_B_g8Zm9LJX0_1;
	wire w_dff_B_iufyHvuQ4_1;
	wire w_dff_B_Wa2XdwjX7_1;
	wire w_dff_B_K6xUvzdL9_1;
	wire w_dff_B_OgvBeiFM7_1;
	wire w_dff_B_sLV6BVkR5_1;
	wire w_dff_B_Ej2EvRIy2_1;
	wire w_dff_B_HGsJMk7P0_1;
	wire w_dff_B_gjfCaYEd9_1;
	wire w_dff_B_urQqdP6W4_1;
	wire w_dff_B_rd9rnUmv2_1;
	wire w_dff_B_7zEgOf3D5_1;
	wire w_dff_B_R4kYRWuP0_1;
	wire w_dff_B_7yUVFmDn0_1;
	wire w_dff_B_WUXOmaGF5_1;
	wire w_dff_B_AyXoPT2q4_1;
	wire w_dff_B_yoITZG6x9_1;
	wire w_dff_B_j8H2qCDz2_1;
	wire w_dff_B_cxJ5m42a9_1;
	wire w_dff_B_3kJ06I5f3_1;
	wire w_dff_B_7G3xDoNL0_1;
	wire w_dff_B_kdItoFeT0_1;
	wire w_dff_B_qPjCYXlb9_1;
	wire w_dff_B_KjKFHHGJ3_1;
	wire w_dff_B_4H8rZfp22_1;
	wire w_dff_B_I6ZHTxQ72_1;
	wire w_dff_B_mAIZ0iRx5_1;
	wire w_dff_B_N671BKDk2_1;
	wire w_dff_B_zoxs8NpC1_1;
	wire w_dff_B_Q8WXGUNJ9_1;
	wire w_dff_B_Eq45sx0L3_1;
	wire w_dff_B_pYASwdi28_1;
	wire w_dff_B_tMOh0O4u2_1;
	wire w_dff_B_0roOkXH24_1;
	wire w_dff_B_MH69ShYO8_1;
	wire w_dff_B_vSiNR5eF4_1;
	wire w_dff_B_YPeD6d7k1_1;
	wire w_dff_B_fHsyco9E6_1;
	wire w_dff_B_CnWOAJ7q1_1;
	wire w_dff_B_Mxv6c0mD9_1;
	wire w_dff_B_yAllGcT59_1;
	wire w_dff_B_qWiGnwCm2_1;
	wire w_dff_B_iZqOtCPt9_1;
	wire w_dff_B_BBhfh24u9_1;
	wire w_dff_B_rI29TUNV0_1;
	wire w_dff_B_4zmlxP5B9_1;
	wire w_dff_B_9BlZBOlK0_1;
	wire w_dff_B_dGbXgqSD7_1;
	wire w_dff_B_vfag6Alh2_1;
	wire w_dff_B_viRKEOL81_1;
	wire w_dff_B_GwWNSl3K4_1;
	wire w_dff_B_mmGaHJCF4_1;
	wire w_dff_B_EuDKPksJ8_1;
	wire w_dff_B_vJdIGQTd9_1;
	wire w_dff_B_6Q20xzzj1_1;
	wire w_dff_B_z6lZE8jM0_1;
	wire w_dff_B_JzzNGpKQ4_1;
	wire w_dff_B_EoiDjHmx8_1;
	wire w_dff_B_aYMo1f8Q1_1;
	wire w_dff_B_9wosPKm44_1;
	wire w_dff_B_cAUCsaW39_1;
	wire w_dff_B_TPpqxXKK1_1;
	wire w_dff_B_brSNaHyt4_1;
	wire w_dff_B_gj9BSaQ32_0;
	wire w_dff_B_zScffpru6_0;
	wire w_dff_B_eRTzEZpJ6_0;
	wire w_dff_B_01rWgdmJ3_0;
	wire w_dff_B_QuU0yevI8_0;
	wire w_dff_B_WuP55TXA7_0;
	wire w_dff_B_zn9j9xCW5_0;
	wire w_dff_B_wqVOPVUm3_0;
	wire w_dff_B_dN4gfwnQ8_0;
	wire w_dff_B_RenkfMsc9_0;
	wire w_dff_B_cqGmaX3E7_0;
	wire w_dff_B_PtwmYSdd5_0;
	wire w_dff_B_WuZw9MOB7_0;
	wire w_dff_B_IXVE1zvs5_0;
	wire w_dff_B_fimdODgY4_0;
	wire w_dff_B_O4nudeKV7_0;
	wire w_dff_B_HjBxPVmu6_0;
	wire w_dff_B_QNx5d1kF9_0;
	wire w_dff_B_u8AICUb41_0;
	wire w_dff_B_Nw9h7WSn4_0;
	wire w_dff_B_WFLAkxCm6_0;
	wire w_dff_B_dIO8Od0q6_0;
	wire w_dff_B_OnURPUhk5_0;
	wire w_dff_B_1fbtBmKS0_0;
	wire w_dff_B_wX4S2dqZ2_0;
	wire w_dff_B_weSLLnbF3_0;
	wire w_dff_B_hEbhc98o2_0;
	wire w_dff_B_O5FKdVO75_0;
	wire w_dff_B_lwZGOtEz8_0;
	wire w_dff_B_j8v2niyu4_0;
	wire w_dff_B_Cgw5QtpC0_0;
	wire w_dff_B_2b8Jtanv8_0;
	wire w_dff_B_kBRfDvoP4_0;
	wire w_dff_B_Nw7jXWAZ9_0;
	wire w_dff_B_Mf0LqrWX5_0;
	wire w_dff_B_qyZixoqC9_0;
	wire w_dff_B_aiZLZEq63_0;
	wire w_dff_B_1AaDvqDm1_0;
	wire w_dff_B_gH7gHrNK6_0;
	wire w_dff_B_EIVlY7Gq6_0;
	wire w_dff_B_hAg9ZTMY9_0;
	wire w_dff_B_fiBGJqbq1_0;
	wire w_dff_B_ZGRaC1kQ2_0;
	wire w_dff_B_eNxLlYtU5_0;
	wire w_dff_B_oNVlvjEm9_0;
	wire w_dff_B_ypipYVnK0_0;
	wire w_dff_B_G3wt2Ihy5_0;
	wire w_dff_B_LbuN2S981_0;
	wire w_dff_B_TW3FMs1W4_0;
	wire w_dff_B_qKGSCiFM8_0;
	wire w_dff_B_0Sd2KXnC8_0;
	wire w_dff_B_QNWKoSPe6_0;
	wire w_dff_B_xLmYmdXH5_0;
	wire w_dff_B_hYBJVPYE0_0;
	wire w_dff_B_XMqHatDK8_0;
	wire w_dff_B_f5WRGiSU7_0;
	wire w_dff_B_YBjguptx0_0;
	wire w_dff_B_cFs0iOoL4_0;
	wire w_dff_B_kzJ4k9HD4_0;
	wire w_dff_B_vHReqyac4_0;
	wire w_dff_B_lXj30V6V2_0;
	wire w_dff_B_Yr3uBJhz8_0;
	wire w_dff_B_P8fyoIaN1_0;
	wire w_dff_B_ooeeHe1Z9_0;
	wire w_dff_B_1qN8zhd62_0;
	wire w_dff_B_q8WGGNTC8_0;
	wire w_dff_B_Ofpdrk672_0;
	wire w_dff_B_dmE7wIib9_0;
	wire w_dff_B_WCARSoGH8_0;
	wire w_dff_B_RMTzlVVX2_0;
	wire w_dff_B_gPiENw7M9_0;
	wire w_dff_B_cx2KtWNM1_0;
	wire w_dff_B_jgNPEzhL6_0;
	wire w_dff_B_vyv3QZRw0_0;
	wire w_dff_B_ATufaRAT8_0;
	wire w_dff_B_RMFUD2fO6_0;
	wire w_dff_B_IGVwytqN2_0;
	wire w_dff_B_VkCKYLEW6_0;
	wire w_dff_B_p465ngL27_0;
	wire w_dff_B_44xOJOdM7_0;
	wire w_dff_B_UGl0cc1T6_0;
	wire w_dff_B_fBiDhWsS6_0;
	wire w_dff_B_w8lFOCaz9_0;
	wire w_dff_B_fKUl863m0_0;
	wire w_dff_B_UYLDZLJM4_0;
	wire w_dff_B_WTuT0sRw7_0;
	wire w_dff_B_D1pBStHq0_0;
	wire w_dff_B_N7vmbMkQ0_0;
	wire w_dff_B_3nxITtqi1_1;
	wire w_dff_B_OY2rNriK2_1;
	wire w_dff_B_KxDJtCsC5_1;
	wire w_dff_B_MRznJZ2V8_1;
	wire w_dff_B_6hJao4te2_1;
	wire w_dff_B_aNDxRmSo2_1;
	wire w_dff_B_9mDzCuTh4_1;
	wire w_dff_B_TkGFrCbe0_1;
	wire w_dff_B_MvI5NZum1_1;
	wire w_dff_B_OvDfYURa0_1;
	wire w_dff_B_seEix5eN4_1;
	wire w_dff_B_YGK7MZPn7_1;
	wire w_dff_B_YMcqpjlG1_1;
	wire w_dff_B_oR5AoGfk2_1;
	wire w_dff_B_M2eZ4DfO4_1;
	wire w_dff_B_UJmA2lav7_1;
	wire w_dff_B_hfkTVK7o6_1;
	wire w_dff_B_EIInKr7E9_1;
	wire w_dff_B_b9XhOSpz8_1;
	wire w_dff_B_i8DE75Ze0_1;
	wire w_dff_B_etvdKZ7e5_1;
	wire w_dff_B_xT6XSek77_1;
	wire w_dff_B_N8ze5nwB4_1;
	wire w_dff_B_2fPf9uIc4_1;
	wire w_dff_B_pWiraKkQ6_1;
	wire w_dff_B_hxGFuNEE1_1;
	wire w_dff_B_9uXZVZ7o6_1;
	wire w_dff_B_2n8yYbkH4_1;
	wire w_dff_B_qGvwWjX74_1;
	wire w_dff_B_570ADOlS3_1;
	wire w_dff_B_fGGrn6YP6_1;
	wire w_dff_B_JhhTo1ZE2_1;
	wire w_dff_B_g5NZvvAt8_1;
	wire w_dff_B_LaGgbmqZ2_1;
	wire w_dff_B_PAlhKosg6_1;
	wire w_dff_B_gyA1OFlq0_1;
	wire w_dff_B_ovgXJbXd2_1;
	wire w_dff_B_A5e2ravW8_1;
	wire w_dff_B_6Q0caIYh0_1;
	wire w_dff_B_TJLpKMo57_1;
	wire w_dff_B_Iwu02DDs8_1;
	wire w_dff_B_sskXV6pq5_1;
	wire w_dff_B_RixVdW8j2_1;
	wire w_dff_B_CDB3Pimm3_1;
	wire w_dff_B_TsnxBlJj6_1;
	wire w_dff_B_gnt9diSQ7_1;
	wire w_dff_B_ahDyzhe43_1;
	wire w_dff_B_fl9kYm1H7_1;
	wire w_dff_B_KySJAlVy8_1;
	wire w_dff_B_kGAcvuc99_1;
	wire w_dff_B_IBE3bsOk7_1;
	wire w_dff_B_U3epGkXT2_1;
	wire w_dff_B_K1CLJtb48_1;
	wire w_dff_B_Rqg5JfTZ5_1;
	wire w_dff_B_1hafOUpw8_1;
	wire w_dff_B_kc0k9wSE7_1;
	wire w_dff_B_vtFiJc4h0_1;
	wire w_dff_B_tEBBFEtC9_1;
	wire w_dff_B_0nZBMp6Y4_1;
	wire w_dff_B_zJ7KyBYy5_1;
	wire w_dff_B_gsENW5VE5_1;
	wire w_dff_B_z2nQMeJU1_1;
	wire w_dff_B_ccxG0Q207_1;
	wire w_dff_B_o24hhAGX8_1;
	wire w_dff_B_NYlA2kK67_1;
	wire w_dff_B_z2U4Prsj6_1;
	wire w_dff_B_y6G2xfc01_1;
	wire w_dff_B_CAzTvFjT7_1;
	wire w_dff_B_HZtwRYYs1_1;
	wire w_dff_B_2wOj47B74_1;
	wire w_dff_B_3Sqezcf91_1;
	wire w_dff_B_4jvZRNPu1_1;
	wire w_dff_B_zNbb8qII5_1;
	wire w_dff_B_6ySqU7NU6_1;
	wire w_dff_B_4sa4L1va5_1;
	wire w_dff_B_bVK9UKFi6_1;
	wire w_dff_B_mLXAfc796_1;
	wire w_dff_B_TRjy6evf4_1;
	wire w_dff_B_QDBbrq6c2_1;
	wire w_dff_B_fvWpofjd2_1;
	wire w_dff_B_pM9LgozB4_1;
	wire w_dff_B_LswJxzVi3_1;
	wire w_dff_B_KBOyUbQG1_1;
	wire w_dff_B_axP6W0ux6_1;
	wire w_dff_B_1eQjlJ7B5_1;
	wire w_dff_B_LPntHGIh3_1;
	wire w_dff_B_utDSKdr27_1;
	wire w_dff_B_9OfuBhph8_0;
	wire w_dff_B_fSvMGx083_0;
	wire w_dff_B_PbQQjmcP1_0;
	wire w_dff_B_UmIzH0ra0_0;
	wire w_dff_B_2EOuS1kW7_0;
	wire w_dff_B_HJjDZQ491_0;
	wire w_dff_B_FsIxBUry9_0;
	wire w_dff_B_QdOryrZ81_0;
	wire w_dff_B_qDO5vPBl7_0;
	wire w_dff_B_tszjXaEA4_0;
	wire w_dff_B_wlJRwORz2_0;
	wire w_dff_B_SK5LwVko8_0;
	wire w_dff_B_YeYxrDAV9_0;
	wire w_dff_B_5Qp7hdX02_0;
	wire w_dff_B_8ICqi3Ox9_0;
	wire w_dff_B_vyJ9grxt2_0;
	wire w_dff_B_bfs9zKE79_0;
	wire w_dff_B_bxdeaFXv6_0;
	wire w_dff_B_QsY6qUnX4_0;
	wire w_dff_B_j59beE0U8_0;
	wire w_dff_B_z0hlPxAr6_0;
	wire w_dff_B_4tL7UEOV2_0;
	wire w_dff_B_1dkoGQx85_0;
	wire w_dff_B_lm0gTiO35_0;
	wire w_dff_B_srwZ13vA8_0;
	wire w_dff_B_T9q9rx4k3_0;
	wire w_dff_B_S07tiac19_0;
	wire w_dff_B_xUgD5UNb5_0;
	wire w_dff_B_A6fW8pRB0_0;
	wire w_dff_B_crgzXCqM1_0;
	wire w_dff_B_aIqpclKv9_0;
	wire w_dff_B_rYpOO1Mu6_0;
	wire w_dff_B_vm8WZ0yM2_0;
	wire w_dff_B_L3hDfd8S0_0;
	wire w_dff_B_wMRyWpiD0_0;
	wire w_dff_B_Vf80f1Lw3_0;
	wire w_dff_B_zraub0fj5_0;
	wire w_dff_B_uY4V9vDI4_0;
	wire w_dff_B_hPLKAhbe9_0;
	wire w_dff_B_XeI2PEdj6_0;
	wire w_dff_B_byRcTbez4_0;
	wire w_dff_B_aUxFGFSR6_0;
	wire w_dff_B_GONssTcG3_0;
	wire w_dff_B_hZS5ek4N0_0;
	wire w_dff_B_mYEE4hLh4_0;
	wire w_dff_B_utaoV4oG5_0;
	wire w_dff_B_l9AqLoT11_0;
	wire w_dff_B_uexlpWaD7_0;
	wire w_dff_B_3UwJZ2Us6_0;
	wire w_dff_B_ph05CXZ16_0;
	wire w_dff_B_CW0eQWU43_0;
	wire w_dff_B_SmHGQilD7_0;
	wire w_dff_B_Rzn23w105_0;
	wire w_dff_B_QnCJ3FFM2_0;
	wire w_dff_B_egwZnSYa0_0;
	wire w_dff_B_0yDvGr9g3_0;
	wire w_dff_B_0598e1ao2_0;
	wire w_dff_B_QSoSxXWZ6_0;
	wire w_dff_B_VdjDn69y3_0;
	wire w_dff_B_fTT29wPF9_0;
	wire w_dff_B_zxfVbPlO8_0;
	wire w_dff_B_TA34UdTz7_0;
	wire w_dff_B_MoN52Izk1_0;
	wire w_dff_B_Sor7zlqY9_0;
	wire w_dff_B_ZANXWw0N6_0;
	wire w_dff_B_qkDf3kKX9_0;
	wire w_dff_B_b1Qaza8E9_0;
	wire w_dff_B_cpmt8CvA4_0;
	wire w_dff_B_SHVva91F4_0;
	wire w_dff_B_r6PKqLfI1_0;
	wire w_dff_B_AAvzp0KW5_0;
	wire w_dff_B_p3uAXoKr8_0;
	wire w_dff_B_WmF1feBH6_0;
	wire w_dff_B_gIrCgn8u6_0;
	wire w_dff_B_SwLUpiyP0_0;
	wire w_dff_B_XHHSkZBs7_0;
	wire w_dff_B_ZmfgwsEv4_0;
	wire w_dff_B_fJU91JOB5_0;
	wire w_dff_B_SK2pSLPr2_0;
	wire w_dff_B_KSDyklnh5_0;
	wire w_dff_B_AfyInHg87_0;
	wire w_dff_B_bIh4yIkm9_0;
	wire w_dff_B_bD2ZHqTj2_0;
	wire w_dff_B_hc8SK1Fi3_0;
	wire w_dff_B_PPPR0yO03_0;
	wire w_dff_B_NxxGUlsv8_0;
	wire w_dff_B_dfcAYDfk0_0;
	wire w_dff_B_qcSVTYBt6_1;
	wire w_dff_B_kCUZfYTp3_1;
	wire w_dff_B_l9JmYZuV0_1;
	wire w_dff_B_MUTLEILN0_1;
	wire w_dff_B_t1DlIuwm4_1;
	wire w_dff_B_MDmwKUKd8_1;
	wire w_dff_B_ggdNpTeq7_1;
	wire w_dff_B_Sl6ehuhW1_1;
	wire w_dff_B_L2g6XaFm5_1;
	wire w_dff_B_IX9sPtvr1_1;
	wire w_dff_B_faNiQ44i5_1;
	wire w_dff_B_5teCjQA89_1;
	wire w_dff_B_pHMIlqKv2_1;
	wire w_dff_B_0WXk4iqa7_1;
	wire w_dff_B_BU8p5kxc3_1;
	wire w_dff_B_KwNJ0nR89_1;
	wire w_dff_B_HD1v7Uex0_1;
	wire w_dff_B_1XKQHulc3_1;
	wire w_dff_B_uYRl3mGy6_1;
	wire w_dff_B_O7LXoTaD2_1;
	wire w_dff_B_H1ESkHXW7_1;
	wire w_dff_B_NN6KyhtX9_1;
	wire w_dff_B_Pd2Ycupa4_1;
	wire w_dff_B_03GxbXdr8_1;
	wire w_dff_B_MaSD429G4_1;
	wire w_dff_B_DRNPArfw6_1;
	wire w_dff_B_wVgaMNmO0_1;
	wire w_dff_B_CNG9TtUj2_1;
	wire w_dff_B_fDJqvT1B2_1;
	wire w_dff_B_0UytVQ538_1;
	wire w_dff_B_1Zi6cly41_1;
	wire w_dff_B_ZfrVhfV95_1;
	wire w_dff_B_FKubNhMB5_1;
	wire w_dff_B_il7oxq9A9_1;
	wire w_dff_B_r4gNjLID6_1;
	wire w_dff_B_gBvwLckV9_1;
	wire w_dff_B_KAgHEonp2_1;
	wire w_dff_B_NWOYjdxL1_1;
	wire w_dff_B_w5kPSTO77_1;
	wire w_dff_B_mBurp2Wg1_1;
	wire w_dff_B_8ikH037v5_1;
	wire w_dff_B_Jc5yxD6j4_1;
	wire w_dff_B_RIpNZff03_1;
	wire w_dff_B_D6Qr4FjS6_1;
	wire w_dff_B_hatumkC54_1;
	wire w_dff_B_xvc7aVNj9_1;
	wire w_dff_B_dJmtbbsb4_1;
	wire w_dff_B_fH8U0KNH8_1;
	wire w_dff_B_DVfUTmGv6_1;
	wire w_dff_B_wkFIHAjd8_1;
	wire w_dff_B_eQUQcj2A8_1;
	wire w_dff_B_5mEazVqq0_1;
	wire w_dff_B_z8quFIX49_1;
	wire w_dff_B_5ehHha4I4_1;
	wire w_dff_B_B7sZWNWV2_1;
	wire w_dff_B_1R8BjQso5_1;
	wire w_dff_B_4aMiubAG9_1;
	wire w_dff_B_El0fXTge8_1;
	wire w_dff_B_RtkevHbs4_1;
	wire w_dff_B_eagTtNFW7_1;
	wire w_dff_B_HnY2EmTT9_1;
	wire w_dff_B_yibIVmkH0_1;
	wire w_dff_B_DMfWNayZ1_1;
	wire w_dff_B_AdMQCjDj7_1;
	wire w_dff_B_VE2qHRlP4_1;
	wire w_dff_B_5PgKb5Di1_1;
	wire w_dff_B_kJwU9FMJ3_1;
	wire w_dff_B_WCDyewqD5_1;
	wire w_dff_B_Rsfv1YQS6_1;
	wire w_dff_B_20oLA5Fu7_1;
	wire w_dff_B_NEh4Ars43_1;
	wire w_dff_B_MuZtmzvI0_1;
	wire w_dff_B_VqP7gHLh7_1;
	wire w_dff_B_EXarQuNl8_1;
	wire w_dff_B_SYtHEa4P5_1;
	wire w_dff_B_fmhA17n98_1;
	wire w_dff_B_yhtsF8Sz7_1;
	wire w_dff_B_Cn2hHtih0_1;
	wire w_dff_B_8xIVSn6b0_1;
	wire w_dff_B_toIxr72N6_1;
	wire w_dff_B_BFLvQCNi1_1;
	wire w_dff_B_zlMrmKcm4_1;
	wire w_dff_B_cO5bJQqp0_1;
	wire w_dff_B_phmxwEJS6_1;
	wire w_dff_B_cCTExRmf2_1;
	wire w_dff_B_epsTtTK93_1;
	wire w_dff_B_lJKhvoH82_0;
	wire w_dff_B_tYJqsr5I9_0;
	wire w_dff_B_Z3Z7ZH8q4_0;
	wire w_dff_B_RGMB55Qg6_0;
	wire w_dff_B_DpLshpnH9_0;
	wire w_dff_B_UT2eOLfP0_0;
	wire w_dff_B_rhzop9Wj6_0;
	wire w_dff_B_8Lx8gHrN0_0;
	wire w_dff_B_3cAwkOm45_0;
	wire w_dff_B_HNHTCCXO0_0;
	wire w_dff_B_F8LxUllA6_0;
	wire w_dff_B_rX82UoT69_0;
	wire w_dff_B_Ak7edaud8_0;
	wire w_dff_B_RCebTlL39_0;
	wire w_dff_B_59V0tLYw0_0;
	wire w_dff_B_D3UdOmYb1_0;
	wire w_dff_B_xxoqTyml6_0;
	wire w_dff_B_BMkInMR34_0;
	wire w_dff_B_xc42WZ2K7_0;
	wire w_dff_B_3u70UCbM7_0;
	wire w_dff_B_qcnVjCEA7_0;
	wire w_dff_B_3t1jWBqX8_0;
	wire w_dff_B_3sEaB4hb2_0;
	wire w_dff_B_bOJPNF9p3_0;
	wire w_dff_B_LSbV7o3T6_0;
	wire w_dff_B_0gVHR0mp2_0;
	wire w_dff_B_CcVqdpX83_0;
	wire w_dff_B_HhYHRB5A6_0;
	wire w_dff_B_xdK0AGMy6_0;
	wire w_dff_B_mNqA4OR71_0;
	wire w_dff_B_DuajkWtH8_0;
	wire w_dff_B_yiRRm0pg0_0;
	wire w_dff_B_dquNXKj92_0;
	wire w_dff_B_MY61xwSR8_0;
	wire w_dff_B_OqlVEJAF1_0;
	wire w_dff_B_Z3LdAn8U1_0;
	wire w_dff_B_4WiDP0Jz6_0;
	wire w_dff_B_zNVdezlO2_0;
	wire w_dff_B_6G5koO6k8_0;
	wire w_dff_B_qnyw3YUh8_0;
	wire w_dff_B_hVQt8W721_0;
	wire w_dff_B_h6j9IioH2_0;
	wire w_dff_B_qpQOSbSI1_0;
	wire w_dff_B_dtO7tGe90_0;
	wire w_dff_B_XtxS4THl4_0;
	wire w_dff_B_LyroC0pO7_0;
	wire w_dff_B_se7GK7f21_0;
	wire w_dff_B_DlLxr2Yu4_0;
	wire w_dff_B_HD8vbn4S1_0;
	wire w_dff_B_oDuOkmWK7_0;
	wire w_dff_B_9TE1E8X39_0;
	wire w_dff_B_noti4kox8_0;
	wire w_dff_B_tdplmZdU6_0;
	wire w_dff_B_7EeOCSTE5_0;
	wire w_dff_B_BzLW0QeY4_0;
	wire w_dff_B_TfodfJ7I6_0;
	wire w_dff_B_TeAOA5997_0;
	wire w_dff_B_O2GFG1zm8_0;
	wire w_dff_B_mFtGdxyv1_0;
	wire w_dff_B_wuYptM569_0;
	wire w_dff_B_sIjMrqwr4_0;
	wire w_dff_B_2PfwSk4k2_0;
	wire w_dff_B_Lgz7XXpd8_0;
	wire w_dff_B_mvmbzmkD9_0;
	wire w_dff_B_RMiPg7n25_0;
	wire w_dff_B_hE5szb6K7_0;
	wire w_dff_B_Qvfx0zTR0_0;
	wire w_dff_B_3ElEBm7Y3_0;
	wire w_dff_B_sSJRl0zJ3_0;
	wire w_dff_B_nkWTR3151_0;
	wire w_dff_B_9XRJmcUB6_0;
	wire w_dff_B_J2wQ01T72_0;
	wire w_dff_B_weR9CNAu3_0;
	wire w_dff_B_81W8Bcd78_0;
	wire w_dff_B_WEX9TPsK2_0;
	wire w_dff_B_CxjRKDCx8_0;
	wire w_dff_B_sKnetmQq7_0;
	wire w_dff_B_oA16ioMu6_0;
	wire w_dff_B_TLmonIpi5_0;
	wire w_dff_B_HqjuU3ck9_0;
	wire w_dff_B_jG98F9on0_0;
	wire w_dff_B_GwOesIIM8_0;
	wire w_dff_B_ni1zVnKN5_0;
	wire w_dff_B_xJLu7Dhv0_0;
	wire w_dff_B_BTdgaiJE3_0;
	wire w_dff_B_f56FFK1t6_0;
	wire w_dff_B_zbQvJ6C20_1;
	wire w_dff_B_qkZKEyZM5_1;
	wire w_dff_B_j4xkmDK01_1;
	wire w_dff_B_zatxTxgJ2_1;
	wire w_dff_B_z23GvKJy1_1;
	wire w_dff_B_FU5uW0LL5_1;
	wire w_dff_B_0JOslABT7_1;
	wire w_dff_B_zfaeMbhO7_1;
	wire w_dff_B_By6RENUn8_1;
	wire w_dff_B_Cm0JmzQM0_1;
	wire w_dff_B_MRWRJWiv5_1;
	wire w_dff_B_bKcHDVgq7_1;
	wire w_dff_B_agEp6D0J7_1;
	wire w_dff_B_yXzGxSnQ9_1;
	wire w_dff_B_27yZqm3R3_1;
	wire w_dff_B_jOX0Y95X4_1;
	wire w_dff_B_JG3sCRf83_1;
	wire w_dff_B_ofZCAthg4_1;
	wire w_dff_B_Wlj5ZjIk6_1;
	wire w_dff_B_Ct3kltv05_1;
	wire w_dff_B_lp7XH4td4_1;
	wire w_dff_B_t8nnAsFa4_1;
	wire w_dff_B_iIHAmn9P9_1;
	wire w_dff_B_9QUtU3ri9_1;
	wire w_dff_B_JJZDMfo27_1;
	wire w_dff_B_hdB5Vu0Y0_1;
	wire w_dff_B_GCPQZIcq3_1;
	wire w_dff_B_aLlYiWik5_1;
	wire w_dff_B_grzNRwks5_1;
	wire w_dff_B_XYADlfYb7_1;
	wire w_dff_B_MiP3P8gZ6_1;
	wire w_dff_B_L2NoJ0596_1;
	wire w_dff_B_8RkYEkTS8_1;
	wire w_dff_B_k2IuLtRU2_1;
	wire w_dff_B_05SpV9JD0_1;
	wire w_dff_B_vRPA8CpO5_1;
	wire w_dff_B_Iss29SFq5_1;
	wire w_dff_B_MkWsVnk81_1;
	wire w_dff_B_SnWspLte0_1;
	wire w_dff_B_v7h1jybE7_1;
	wire w_dff_B_tWfbd1wB9_1;
	wire w_dff_B_uiYCYSo46_1;
	wire w_dff_B_hef6HTNh4_1;
	wire w_dff_B_KsnqZkag3_1;
	wire w_dff_B_zoYKeZuQ2_1;
	wire w_dff_B_lqUlsJr93_1;
	wire w_dff_B_2qg6iKSM7_1;
	wire w_dff_B_caYLUQbm4_1;
	wire w_dff_B_0rqwwXhM5_1;
	wire w_dff_B_xfgpOJRk4_1;
	wire w_dff_B_QrJq7BVy9_1;
	wire w_dff_B_r62YTe5a1_1;
	wire w_dff_B_wXIeoSUK9_1;
	wire w_dff_B_FtB8rJSI9_1;
	wire w_dff_B_889gqyHm2_1;
	wire w_dff_B_yRAVixMX4_1;
	wire w_dff_B_Kv6Gql8K6_1;
	wire w_dff_B_9ongw8eY6_1;
	wire w_dff_B_VFdd7dNM6_1;
	wire w_dff_B_johDkqTX1_1;
	wire w_dff_B_xG0IAOyf5_1;
	wire w_dff_B_ontINZd45_1;
	wire w_dff_B_mponBiiv1_1;
	wire w_dff_B_7oyNpD7Y9_1;
	wire w_dff_B_MHFPgTmc5_1;
	wire w_dff_B_Un8VFwHd3_1;
	wire w_dff_B_AZY4aIGL8_1;
	wire w_dff_B_hWbl4can7_1;
	wire w_dff_B_zTtvZ0Ge9_1;
	wire w_dff_B_HgqGc6jD2_1;
	wire w_dff_B_kbJGJARV1_1;
	wire w_dff_B_3TvpvZzv1_1;
	wire w_dff_B_q0e6NACN2_1;
	wire w_dff_B_Pb5dlJDf5_1;
	wire w_dff_B_rZYql6Ih7_1;
	wire w_dff_B_RPzSUgBZ5_1;
	wire w_dff_B_ugtsLmQ65_1;
	wire w_dff_B_U3ER6DbH1_1;
	wire w_dff_B_BMdQNpqJ9_1;
	wire w_dff_B_BClkdMQc4_1;
	wire w_dff_B_gBg1UEpp0_1;
	wire w_dff_B_qFVlKnSy1_1;
	wire w_dff_B_TBbi45624_1;
	wire w_dff_B_nZFY3ZaV0_1;
	wire w_dff_B_8UlPWcMp1_1;
	wire w_dff_B_3msDc8HK9_0;
	wire w_dff_B_dmrV2Ji61_0;
	wire w_dff_B_FdG9gOQB6_0;
	wire w_dff_B_0n35iexP7_0;
	wire w_dff_B_QWhhxulS7_0;
	wire w_dff_B_EVumF80J0_0;
	wire w_dff_B_PTML7Nqq4_0;
	wire w_dff_B_4esAWS705_0;
	wire w_dff_B_lMgLuAUV7_0;
	wire w_dff_B_UVXGxXoK5_0;
	wire w_dff_B_iBUuvlbL8_0;
	wire w_dff_B_g7anM3Pd5_0;
	wire w_dff_B_MFxd858v7_0;
	wire w_dff_B_k18YaPRN6_0;
	wire w_dff_B_yFmWwlCQ8_0;
	wire w_dff_B_aRYMJqhW1_0;
	wire w_dff_B_VZTQcXus1_0;
	wire w_dff_B_QdAZzkMb6_0;
	wire w_dff_B_SoPw7wRM5_0;
	wire w_dff_B_5BTjZDLb8_0;
	wire w_dff_B_FHSyB3Yj9_0;
	wire w_dff_B_aX53TefW5_0;
	wire w_dff_B_QIUiqdd55_0;
	wire w_dff_B_qLMAomy10_0;
	wire w_dff_B_dzJuL4r81_0;
	wire w_dff_B_qExanZTJ3_0;
	wire w_dff_B_DMVlJJIf6_0;
	wire w_dff_B_b6kgwMDK7_0;
	wire w_dff_B_BC2WxAwk3_0;
	wire w_dff_B_z3GeC4HW3_0;
	wire w_dff_B_ihpTs5eF0_0;
	wire w_dff_B_sETUEPwu2_0;
	wire w_dff_B_4U1pC6Ie1_0;
	wire w_dff_B_RtEXnXBG7_0;
	wire w_dff_B_udzItZ6C4_0;
	wire w_dff_B_weMw1psK9_0;
	wire w_dff_B_C2G07WEF1_0;
	wire w_dff_B_8TRDEEBO4_0;
	wire w_dff_B_QB1IXyew8_0;
	wire w_dff_B_qp26auB63_0;
	wire w_dff_B_kI2dXGRk5_0;
	wire w_dff_B_XqOtYwS99_0;
	wire w_dff_B_YFmMzJDX4_0;
	wire w_dff_B_puvZOHJr3_0;
	wire w_dff_B_MnVza0pd2_0;
	wire w_dff_B_GIMAJzJL7_0;
	wire w_dff_B_4exDOfFQ0_0;
	wire w_dff_B_UnNaBk9q7_0;
	wire w_dff_B_6jzhcUbu5_0;
	wire w_dff_B_eM0hB67C3_0;
	wire w_dff_B_s4pMU2ic3_0;
	wire w_dff_B_WV0Zihy29_0;
	wire w_dff_B_A4ytXW2y6_0;
	wire w_dff_B_3mDjKqEZ6_0;
	wire w_dff_B_bf2FZPon1_0;
	wire w_dff_B_xJBqJB2M5_0;
	wire w_dff_B_ZZU372l87_0;
	wire w_dff_B_F0kdrYZa2_0;
	wire w_dff_B_UiJ1EqSr9_0;
	wire w_dff_B_uWwRSsrZ1_0;
	wire w_dff_B_haQDWQAZ6_0;
	wire w_dff_B_SwhZn6SF5_0;
	wire w_dff_B_wezeHtDL5_0;
	wire w_dff_B_RBTvXJq86_0;
	wire w_dff_B_mSny4DcO2_0;
	wire w_dff_B_KtRvRu983_0;
	wire w_dff_B_TFZFbgvc4_0;
	wire w_dff_B_H4O1GOiU3_0;
	wire w_dff_B_VSQ0QRtf2_0;
	wire w_dff_B_TuVIazGH6_0;
	wire w_dff_B_nB4Z9b8r8_0;
	wire w_dff_B_qTBND50X4_0;
	wire w_dff_B_DoYeaq9e6_0;
	wire w_dff_B_ijtOPvtT0_0;
	wire w_dff_B_YUpIWiZ31_0;
	wire w_dff_B_s266H8zw3_0;
	wire w_dff_B_D3oVOrNU8_0;
	wire w_dff_B_7aN59Uv71_0;
	wire w_dff_B_uSN6thyP8_0;
	wire w_dff_B_ldrRvn527_0;
	wire w_dff_B_eHTTBcll6_0;
	wire w_dff_B_vdCbUMJ06_0;
	wire w_dff_B_HvHUCB9z8_0;
	wire w_dff_B_Sx2NmIou8_0;
	wire w_dff_B_LbDxoEnS2_0;
	wire w_dff_B_GKtRYPrW2_1;
	wire w_dff_B_3F1aMPwX3_1;
	wire w_dff_B_7ipyUibD1_1;
	wire w_dff_B_3Z4uc6Es6_1;
	wire w_dff_B_RprIe1Dt1_1;
	wire w_dff_B_rjLJBud54_1;
	wire w_dff_B_8fv1Bf5S2_1;
	wire w_dff_B_ZrPlNy286_1;
	wire w_dff_B_9W4sielV8_1;
	wire w_dff_B_Kt2JAZpY6_1;
	wire w_dff_B_HCpcGmzM1_1;
	wire w_dff_B_cx7bQocO7_1;
	wire w_dff_B_EhfcKy846_1;
	wire w_dff_B_tphxZSMk1_1;
	wire w_dff_B_Ndad2jbe8_1;
	wire w_dff_B_hS1wXzlv5_1;
	wire w_dff_B_jtawZMZS5_1;
	wire w_dff_B_rqfDRn3X2_1;
	wire w_dff_B_r6g8H71W1_1;
	wire w_dff_B_sqEqgQik3_1;
	wire w_dff_B_Ws5szzQx2_1;
	wire w_dff_B_sjsLXqOQ3_1;
	wire w_dff_B_GmlnaTke8_1;
	wire w_dff_B_B5BYmlYS1_1;
	wire w_dff_B_QKoKqY614_1;
	wire w_dff_B_7Chx3MfP0_1;
	wire w_dff_B_LGkYfDpn3_1;
	wire w_dff_B_gudizypC1_1;
	wire w_dff_B_jHkHUqva5_1;
	wire w_dff_B_dQCzMzMy0_1;
	wire w_dff_B_OF3ywdzv0_1;
	wire w_dff_B_E3TqWAjh0_1;
	wire w_dff_B_HBSvAhJa4_1;
	wire w_dff_B_itaB3R5g2_1;
	wire w_dff_B_SD4QNh4g1_1;
	wire w_dff_B_XvZXIE296_1;
	wire w_dff_B_K87zYtj92_1;
	wire w_dff_B_2qWdqTH73_1;
	wire w_dff_B_4odDBRJw6_1;
	wire w_dff_B_BBh2S4Na3_1;
	wire w_dff_B_cnhIEryX7_1;
	wire w_dff_B_ztrWRd7J8_1;
	wire w_dff_B_j39FyQzb7_1;
	wire w_dff_B_eBM8205w1_1;
	wire w_dff_B_CURzSjlm4_1;
	wire w_dff_B_Q4VwXRyH6_1;
	wire w_dff_B_8xYdzrIY1_1;
	wire w_dff_B_4yV7nJBP4_1;
	wire w_dff_B_l6Ltd7GT5_1;
	wire w_dff_B_qMEhjrSU0_1;
	wire w_dff_B_tnyo2G0o6_1;
	wire w_dff_B_u3kneydC3_1;
	wire w_dff_B_nj8hUOoP3_1;
	wire w_dff_B_S1fm64og5_1;
	wire w_dff_B_8e04RCjO4_1;
	wire w_dff_B_JIUf7FBz2_1;
	wire w_dff_B_5pIGDXSh9_1;
	wire w_dff_B_bu60NKrG4_1;
	wire w_dff_B_97A3pkXr7_1;
	wire w_dff_B_tuagi6Ba0_1;
	wire w_dff_B_u5SYOHUA9_1;
	wire w_dff_B_Kd09eGeT9_1;
	wire w_dff_B_UWURkiLl8_1;
	wire w_dff_B_bHHS2Dnx6_1;
	wire w_dff_B_CYcAG6bC2_1;
	wire w_dff_B_ZQ5XIhPt2_1;
	wire w_dff_B_9DhvbhLG9_1;
	wire w_dff_B_mwg3qWgc6_1;
	wire w_dff_B_Od2dIDMp2_1;
	wire w_dff_B_PY1v2Rwt9_1;
	wire w_dff_B_vSuWtJfl2_1;
	wire w_dff_B_MukH1qL56_1;
	wire w_dff_B_oC8QApYL6_1;
	wire w_dff_B_2AeYhtpO0_1;
	wire w_dff_B_nyqwvJoK4_1;
	wire w_dff_B_ysxui0172_1;
	wire w_dff_B_LVVtV4Qm1_1;
	wire w_dff_B_FMVPXCWy1_1;
	wire w_dff_B_COstpe8X7_1;
	wire w_dff_B_CBkZ6ETZ4_1;
	wire w_dff_B_Vbuzfyop4_1;
	wire w_dff_B_FjY0zC7k0_1;
	wire w_dff_B_n0qrL1M48_1;
	wire w_dff_B_etx97ig43_1;
	wire w_dff_B_IS9gqbo12_0;
	wire w_dff_B_9Vj3Nt8X5_0;
	wire w_dff_B_SXu1pMQS5_0;
	wire w_dff_B_n3WVT6mU1_0;
	wire w_dff_B_raRSMuC74_0;
	wire w_dff_B_fPUHfe4T1_0;
	wire w_dff_B_5vzL2BVh1_0;
	wire w_dff_B_2OmAh31x7_0;
	wire w_dff_B_zJ4FtWxm1_0;
	wire w_dff_B_JsgkxfMI9_0;
	wire w_dff_B_blQQ2uMx4_0;
	wire w_dff_B_gepnvB4j8_0;
	wire w_dff_B_oX5E9BmF8_0;
	wire w_dff_B_HVeHePan1_0;
	wire w_dff_B_zHp0ZRjP8_0;
	wire w_dff_B_vXtK9Mlt5_0;
	wire w_dff_B_h7tdAW7D8_0;
	wire w_dff_B_Zlikh2j86_0;
	wire w_dff_B_VPTpC2H45_0;
	wire w_dff_B_VvMr97nE3_0;
	wire w_dff_B_NahAC0Eo9_0;
	wire w_dff_B_280qH7kL6_0;
	wire w_dff_B_MlKTwdTh4_0;
	wire w_dff_B_aGjj0Nh93_0;
	wire w_dff_B_LAOfmeim3_0;
	wire w_dff_B_h0ZQAsrA1_0;
	wire w_dff_B_Rbgkyd2G8_0;
	wire w_dff_B_RUOWKRLc3_0;
	wire w_dff_B_Zqy47IMD9_0;
	wire w_dff_B_Xck9EUzY8_0;
	wire w_dff_B_ypyvD6Bz4_0;
	wire w_dff_B_HpUYi8oQ3_0;
	wire w_dff_B_cRZ5Imnm4_0;
	wire w_dff_B_mDCQl1v25_0;
	wire w_dff_B_mIiKfnyG8_0;
	wire w_dff_B_lgZJCgZP1_0;
	wire w_dff_B_7ndmbS6K9_0;
	wire w_dff_B_rTCVd5N99_0;
	wire w_dff_B_7E3pJjH17_0;
	wire w_dff_B_g6nplmB82_0;
	wire w_dff_B_h9cRijoQ3_0;
	wire w_dff_B_fFVisHlT2_0;
	wire w_dff_B_FIWK01KE2_0;
	wire w_dff_B_gs5iODbn6_0;
	wire w_dff_B_DMyofCCZ7_0;
	wire w_dff_B_bhVr24TV4_0;
	wire w_dff_B_tI6gCD1J8_0;
	wire w_dff_B_Q3fAfedx4_0;
	wire w_dff_B_2hHLb52J6_0;
	wire w_dff_B_UXHygEj31_0;
	wire w_dff_B_MPWVDqaN0_0;
	wire w_dff_B_dwHbIRQV6_0;
	wire w_dff_B_kFtrtvSs1_0;
	wire w_dff_B_Ys4FiAHx0_0;
	wire w_dff_B_9YrrfuX94_0;
	wire w_dff_B_5AGYM25N5_0;
	wire w_dff_B_qHUkpTyI3_0;
	wire w_dff_B_fOUDaivR3_0;
	wire w_dff_B_alYZk9ks1_0;
	wire w_dff_B_IO2CtH3y3_0;
	wire w_dff_B_KtHIdWub0_0;
	wire w_dff_B_XP0zdyAC9_0;
	wire w_dff_B_zU4AQxrN6_0;
	wire w_dff_B_UcJWm4uf0_0;
	wire w_dff_B_uiSNVyjp4_0;
	wire w_dff_B_QZiYkCeo5_0;
	wire w_dff_B_V9sIaIe34_0;
	wire w_dff_B_mRo9FUhG9_0;
	wire w_dff_B_32yQTYIV2_0;
	wire w_dff_B_50EwaRSy4_0;
	wire w_dff_B_ekMlRWdn7_0;
	wire w_dff_B_Em4aZHXi9_0;
	wire w_dff_B_kEpVFEnH7_0;
	wire w_dff_B_YZgb51P05_0;
	wire w_dff_B_WxaoF8hO3_0;
	wire w_dff_B_44JFbs0e0_0;
	wire w_dff_B_bWFses4t8_0;
	wire w_dff_B_EVWYhNQk7_0;
	wire w_dff_B_fEoxjw221_0;
	wire w_dff_B_SJ3NDSfr7_0;
	wire w_dff_B_xf81cLkS2_0;
	wire w_dff_B_NfmeXSyA9_0;
	wire w_dff_B_ihb62fBO1_0;
	wire w_dff_B_mRYvO6bw1_0;
	wire w_dff_B_Mq8qISei8_1;
	wire w_dff_B_zVwl7onX2_1;
	wire w_dff_B_jkhEDHER3_1;
	wire w_dff_B_sjCYmBud1_1;
	wire w_dff_B_jovfwT9y8_1;
	wire w_dff_B_dByslP4G1_1;
	wire w_dff_B_TqaYnsJW8_1;
	wire w_dff_B_2N9Enggv5_1;
	wire w_dff_B_M2l7D4P54_1;
	wire w_dff_B_CUaXZ9OF8_1;
	wire w_dff_B_ajq5lKV57_1;
	wire w_dff_B_0Oeh6Ivd1_1;
	wire w_dff_B_ALDAxfQp4_1;
	wire w_dff_B_XujCND2b7_1;
	wire w_dff_B_YZ3L0UOX4_1;
	wire w_dff_B_wLzp8yy96_1;
	wire w_dff_B_1W53RdhW9_1;
	wire w_dff_B_8sVhLcJ53_1;
	wire w_dff_B_VneuQfHg2_1;
	wire w_dff_B_d9oWTCcI3_1;
	wire w_dff_B_Ib90Bc2V6_1;
	wire w_dff_B_ZO7bX5aP4_1;
	wire w_dff_B_fy2DG2792_1;
	wire w_dff_B_x9u41iBL8_1;
	wire w_dff_B_qBqDGxo13_1;
	wire w_dff_B_HZUFPXbX1_1;
	wire w_dff_B_piUxztbY6_1;
	wire w_dff_B_KTdvDgsl7_1;
	wire w_dff_B_0ejnl01W7_1;
	wire w_dff_B_gmtA3fTG3_1;
	wire w_dff_B_ZeE6vPmm5_1;
	wire w_dff_B_pkTlWEEt6_1;
	wire w_dff_B_K0xiAILb1_1;
	wire w_dff_B_Fa6nHqKX9_1;
	wire w_dff_B_iP1Y05CH9_1;
	wire w_dff_B_hSyM2ESL0_1;
	wire w_dff_B_SUJ9gpXS1_1;
	wire w_dff_B_Gj7GG32j2_1;
	wire w_dff_B_o68rxA8H6_1;
	wire w_dff_B_Rr9TWc367_1;
	wire w_dff_B_NDxObvPn9_1;
	wire w_dff_B_dPqgRTiZ7_1;
	wire w_dff_B_6vK1fI4O5_1;
	wire w_dff_B_IYn3bxHz2_1;
	wire w_dff_B_qVwDrg6t2_1;
	wire w_dff_B_ia5XpHfb1_1;
	wire w_dff_B_Q9RYIJyk5_1;
	wire w_dff_B_zoX5ATlX5_1;
	wire w_dff_B_wbM3uAG80_1;
	wire w_dff_B_7Xdc5KDA2_1;
	wire w_dff_B_eMjTXNVt2_1;
	wire w_dff_B_OyvQbfIX6_1;
	wire w_dff_B_LkLd7c4S5_1;
	wire w_dff_B_D1JzKo7d1_1;
	wire w_dff_B_8eNJeAIF6_1;
	wire w_dff_B_VMsSEPD41_1;
	wire w_dff_B_3V3AGUMO8_1;
	wire w_dff_B_n5zI5kEv0_1;
	wire w_dff_B_cOFKFadO3_1;
	wire w_dff_B_PwtDI52T9_1;
	wire w_dff_B_09g35pyA2_1;
	wire w_dff_B_FeR02UvE6_1;
	wire w_dff_B_5kcb8wRv6_1;
	wire w_dff_B_XLby0v3k4_1;
	wire w_dff_B_YIcD3ovG5_1;
	wire w_dff_B_lJ7GpQk82_1;
	wire w_dff_B_CbZ06e4w7_1;
	wire w_dff_B_g0qywdFH7_1;
	wire w_dff_B_R7UTxnki4_1;
	wire w_dff_B_wri3YED41_1;
	wire w_dff_B_O8bczUst3_1;
	wire w_dff_B_38fwY4Ln6_1;
	wire w_dff_B_faHhFQx39_1;
	wire w_dff_B_rAkmUrHa2_1;
	wire w_dff_B_8IY2qjMo0_1;
	wire w_dff_B_DVsHxG738_1;
	wire w_dff_B_Dz1BOvfe3_1;
	wire w_dff_B_2OLArSu79_1;
	wire w_dff_B_uvEgy2uw2_1;
	wire w_dff_B_gFNdgW0F4_1;
	wire w_dff_B_9iZ9wvN55_1;
	wire w_dff_B_R04kQDea7_1;
	wire w_dff_B_pqpOHVfn2_1;
	wire w_dff_B_lbx0bJ3I1_0;
	wire w_dff_B_UgaUlG2h9_0;
	wire w_dff_B_bgm9I2RO3_0;
	wire w_dff_B_YQcMCGIS2_0;
	wire w_dff_B_w58wDCjv1_0;
	wire w_dff_B_kywKR1cJ6_0;
	wire w_dff_B_ulUMzjEr8_0;
	wire w_dff_B_4ZxSj76o7_0;
	wire w_dff_B_eMYbxtrk4_0;
	wire w_dff_B_fSm2hHlu7_0;
	wire w_dff_B_yXjcUZOK0_0;
	wire w_dff_B_1zLrhq7K1_0;
	wire w_dff_B_5wjrOJs38_0;
	wire w_dff_B_XMzR0ZiJ0_0;
	wire w_dff_B_gPfC5QxC4_0;
	wire w_dff_B_syhuGrkJ1_0;
	wire w_dff_B_xMp1MZqg5_0;
	wire w_dff_B_5RpfC5KX3_0;
	wire w_dff_B_8mrylY1Q0_0;
	wire w_dff_B_ovHkF9IV0_0;
	wire w_dff_B_rvcFtqMG9_0;
	wire w_dff_B_2sfw3t971_0;
	wire w_dff_B_rlgkM11P5_0;
	wire w_dff_B_N7gOJYOh8_0;
	wire w_dff_B_Ipbu9Ot25_0;
	wire w_dff_B_wYqg17or3_0;
	wire w_dff_B_52rEqSmP5_0;
	wire w_dff_B_Y4dLJha30_0;
	wire w_dff_B_1dsZkoae8_0;
	wire w_dff_B_TAyn4PGm2_0;
	wire w_dff_B_zR8DzHqz5_0;
	wire w_dff_B_JPxwGHbe9_0;
	wire w_dff_B_F1bEbhZw3_0;
	wire w_dff_B_Ovtj5Uu34_0;
	wire w_dff_B_mlE9rzgM9_0;
	wire w_dff_B_F2dJ8WjC6_0;
	wire w_dff_B_LQ3kaRtF8_0;
	wire w_dff_B_Qb5hRfiD2_0;
	wire w_dff_B_luqFBp6l0_0;
	wire w_dff_B_JSXjiCEQ0_0;
	wire w_dff_B_nyu6l83o3_0;
	wire w_dff_B_DUPsTurq4_0;
	wire w_dff_B_3J4ZgUEC1_0;
	wire w_dff_B_1IBbH39q0_0;
	wire w_dff_B_pn6a7Tt96_0;
	wire w_dff_B_Bbq4SO8H0_0;
	wire w_dff_B_ujHpbwvQ9_0;
	wire w_dff_B_TNQBdK2p8_0;
	wire w_dff_B_UoMHYi4T2_0;
	wire w_dff_B_ZVSmNbLf7_0;
	wire w_dff_B_49oXdpNJ2_0;
	wire w_dff_B_nTfSG4iy3_0;
	wire w_dff_B_Oy80N22j5_0;
	wire w_dff_B_CHQb8XLy8_0;
	wire w_dff_B_YJkhyArE6_0;
	wire w_dff_B_QAH5LVWN5_0;
	wire w_dff_B_mh4uii889_0;
	wire w_dff_B_zfdsILgT3_0;
	wire w_dff_B_SzkvICuc8_0;
	wire w_dff_B_uqsLirJX5_0;
	wire w_dff_B_uskQaVMn5_0;
	wire w_dff_B_BHZ6k7Y53_0;
	wire w_dff_B_XH8yS9iD4_0;
	wire w_dff_B_R5zlN7zy5_0;
	wire w_dff_B_V8anR2zM2_0;
	wire w_dff_B_ETi7pgUl8_0;
	wire w_dff_B_lVz8UHwx9_0;
	wire w_dff_B_KvRRpVXS0_0;
	wire w_dff_B_wPXMR1n72_0;
	wire w_dff_B_RgdBGlg80_0;
	wire w_dff_B_dCaPC60s2_0;
	wire w_dff_B_zftcPdEp8_0;
	wire w_dff_B_3UL5uNh81_0;
	wire w_dff_B_XBqXH6D92_0;
	wire w_dff_B_QmfgcSuP6_0;
	wire w_dff_B_tNRYvELa2_0;
	wire w_dff_B_QGUwBrrA3_0;
	wire w_dff_B_vOhWD8ma3_0;
	wire w_dff_B_fNLVoglA7_0;
	wire w_dff_B_oeLcs5Fp4_0;
	wire w_dff_B_v73dFm1n7_0;
	wire w_dff_B_AtsoBtob9_0;
	wire w_dff_B_XuAALr0W2_0;
	wire w_dff_B_Xd3qesh12_1;
	wire w_dff_B_Eokc923Z1_1;
	wire w_dff_B_oAHzyOSn4_1;
	wire w_dff_B_ICP5pvP52_1;
	wire w_dff_B_QXMlNoS57_1;
	wire w_dff_B_HhcMAKUO9_1;
	wire w_dff_B_z2dU9mrH0_1;
	wire w_dff_B_DTG1yr730_1;
	wire w_dff_B_kPYFWJQU5_1;
	wire w_dff_B_eldJobIu1_1;
	wire w_dff_B_seIxoZZz2_1;
	wire w_dff_B_L1ssJrKX0_1;
	wire w_dff_B_zjULwgap5_1;
	wire w_dff_B_1gm5Ydf39_1;
	wire w_dff_B_8eSX5zWY4_1;
	wire w_dff_B_DFHIWMFM8_1;
	wire w_dff_B_oXXmaJfU7_1;
	wire w_dff_B_E88Fkyhd9_1;
	wire w_dff_B_sGUqVLio2_1;
	wire w_dff_B_9uUW4FKq6_1;
	wire w_dff_B_cApTODzx3_1;
	wire w_dff_B_u9Y1Kk1M2_1;
	wire w_dff_B_yzvPv0Gf2_1;
	wire w_dff_B_e277gc5k7_1;
	wire w_dff_B_5yP6dijU2_1;
	wire w_dff_B_syBHCo5S8_1;
	wire w_dff_B_s6tREeMO8_1;
	wire w_dff_B_RnLjzHSX0_1;
	wire w_dff_B_eCalJcio6_1;
	wire w_dff_B_ksb7gZyq3_1;
	wire w_dff_B_9qaNjVeX6_1;
	wire w_dff_B_O8bgULBf5_1;
	wire w_dff_B_qY474FcQ6_1;
	wire w_dff_B_CFFeTcxm3_1;
	wire w_dff_B_399lFJV69_1;
	wire w_dff_B_53UHsDp51_1;
	wire w_dff_B_tYs46H4D0_1;
	wire w_dff_B_rt75IlMh2_1;
	wire w_dff_B_2O0ggyf76_1;
	wire w_dff_B_0o1vNFXX9_1;
	wire w_dff_B_5rKo3sG89_1;
	wire w_dff_B_YRGyUjuk0_1;
	wire w_dff_B_doE5mHOh9_1;
	wire w_dff_B_fmMw772B1_1;
	wire w_dff_B_KvZawl2d8_1;
	wire w_dff_B_u9Yjhk0a5_1;
	wire w_dff_B_kgyJzPCJ1_1;
	wire w_dff_B_O1FazG0M5_1;
	wire w_dff_B_w4H1VIdU4_1;
	wire w_dff_B_774dSw5z2_1;
	wire w_dff_B_lMaWDzSI2_1;
	wire w_dff_B_y6CplWrf0_1;
	wire w_dff_B_bnYHiXBW9_1;
	wire w_dff_B_3kQGj0Cf9_1;
	wire w_dff_B_2WtXukM07_1;
	wire w_dff_B_sSUNASYl8_1;
	wire w_dff_B_zveSQgSV5_1;
	wire w_dff_B_b3HkcRC63_1;
	wire w_dff_B_DCuFrT1Q1_1;
	wire w_dff_B_FqulapPz9_1;
	wire w_dff_B_jACIDB1M8_1;
	wire w_dff_B_PqOy7b1u8_1;
	wire w_dff_B_ef8zidSD8_1;
	wire w_dff_B_ly868IGg7_1;
	wire w_dff_B_48xh1Xbv7_1;
	wire w_dff_B_ENuE0Vz92_1;
	wire w_dff_B_POWywMl40_1;
	wire w_dff_B_vImdWakB7_1;
	wire w_dff_B_hx1EwlHH6_1;
	wire w_dff_B_rdN34DIu8_1;
	wire w_dff_B_AyvGowR26_1;
	wire w_dff_B_z7cI5L9c8_1;
	wire w_dff_B_25t8uufX2_1;
	wire w_dff_B_x7ePNm8y5_1;
	wire w_dff_B_aUdLdDXa1_1;
	wire w_dff_B_IjxD3l1I6_1;
	wire w_dff_B_gisVeJyT4_1;
	wire w_dff_B_9oyZfYz89_1;
	wire w_dff_B_PTXz50yE3_1;
	wire w_dff_B_PkGbuQfZ3_1;
	wire w_dff_B_RuSpPh4Y8_1;
	wire w_dff_B_GzgJUVn93_1;
	wire w_dff_B_XcvAxMVt9_0;
	wire w_dff_B_RpVKE8vT4_0;
	wire w_dff_B_9vBSIjVw6_0;
	wire w_dff_B_NRtPG4HM1_0;
	wire w_dff_B_iTFCQodU7_0;
	wire w_dff_B_eNZRrUkz9_0;
	wire w_dff_B_FNGg0k8D4_0;
	wire w_dff_B_a50DlNCi9_0;
	wire w_dff_B_bTonFqOW3_0;
	wire w_dff_B_b73D48xU6_0;
	wire w_dff_B_wiavP2YL6_0;
	wire w_dff_B_xDx47EjO1_0;
	wire w_dff_B_t4SJtfgz5_0;
	wire w_dff_B_m8rltR9S8_0;
	wire w_dff_B_FUZynIAS5_0;
	wire w_dff_B_SNJC5Cqh2_0;
	wire w_dff_B_PuTqYIrU5_0;
	wire w_dff_B_bswICrJG7_0;
	wire w_dff_B_jr1mpQMw5_0;
	wire w_dff_B_IpenWHNU5_0;
	wire w_dff_B_T7qsEW3G4_0;
	wire w_dff_B_bVuI5yqA8_0;
	wire w_dff_B_xJ3iZ2ii1_0;
	wire w_dff_B_rusifKPM8_0;
	wire w_dff_B_32aZPd3X6_0;
	wire w_dff_B_L8Cgwdgs0_0;
	wire w_dff_B_6rAVLAmc7_0;
	wire w_dff_B_yg4SBqH26_0;
	wire w_dff_B_6wzUchkh8_0;
	wire w_dff_B_XAEVdv4h6_0;
	wire w_dff_B_sseBOyvc7_0;
	wire w_dff_B_GlzUnj512_0;
	wire w_dff_B_f2oUjk3w3_0;
	wire w_dff_B_2zzWnXtA3_0;
	wire w_dff_B_T2vaAMqJ2_0;
	wire w_dff_B_dYNyFugB3_0;
	wire w_dff_B_XxUQXtJi6_0;
	wire w_dff_B_ptd5B7Z85_0;
	wire w_dff_B_49ppE5Yu2_0;
	wire w_dff_B_EIqH16tS9_0;
	wire w_dff_B_s72BTiyB5_0;
	wire w_dff_B_IULCqqVL5_0;
	wire w_dff_B_OPCZ2pQK8_0;
	wire w_dff_B_ttK48AQt5_0;
	wire w_dff_B_yUjJGqob2_0;
	wire w_dff_B_a3fZ0Rio8_0;
	wire w_dff_B_3GhrjSsy0_0;
	wire w_dff_B_3i1rE0Li9_0;
	wire w_dff_B_iz6Tp54D5_0;
	wire w_dff_B_eDt15EWn3_0;
	wire w_dff_B_QNakKLW77_0;
	wire w_dff_B_HDVIR3J11_0;
	wire w_dff_B_UCeS1BTq5_0;
	wire w_dff_B_1GCpW4xq1_0;
	wire w_dff_B_SCkx9vpA6_0;
	wire w_dff_B_sUS44pZR7_0;
	wire w_dff_B_Jz3Hz0aB0_0;
	wire w_dff_B_HPb3SAhM2_0;
	wire w_dff_B_GCwkzC5l9_0;
	wire w_dff_B_SSiLXWJO5_0;
	wire w_dff_B_GSc3vhSl1_0;
	wire w_dff_B_SzGCLdj83_0;
	wire w_dff_B_ny6XWGds6_0;
	wire w_dff_B_cQbPTwoj5_0;
	wire w_dff_B_tKxglLIJ7_0;
	wire w_dff_B_wDB7Jm120_0;
	wire w_dff_B_JpQ9tElH8_0;
	wire w_dff_B_FSeBSD4l2_0;
	wire w_dff_B_m2PCLPWI8_0;
	wire w_dff_B_foavRE1o9_0;
	wire w_dff_B_3iAyf6st6_0;
	wire w_dff_B_x7wKRM273_0;
	wire w_dff_B_FYwZKf7J8_0;
	wire w_dff_B_VgtKyPMi1_0;
	wire w_dff_B_AL7UwVBw4_0;
	wire w_dff_B_7KeJblEc5_0;
	wire w_dff_B_DPn3BabI4_0;
	wire w_dff_B_JmnLm2Ir4_0;
	wire w_dff_B_OZ0Y5C9I6_0;
	wire w_dff_B_urhxRM5H3_0;
	wire w_dff_B_HnA7n8nv2_0;
	wire w_dff_B_kq0cFdQ24_0;
	wire w_dff_B_HGLUILcM4_1;
	wire w_dff_B_FAQyOcLZ7_1;
	wire w_dff_B_ecvuUYPK7_1;
	wire w_dff_B_rHN2QkmK2_1;
	wire w_dff_B_oSpA3vca2_1;
	wire w_dff_B_5ogCHQop0_1;
	wire w_dff_B_LLEgP7sp0_1;
	wire w_dff_B_WtEFNwD22_1;
	wire w_dff_B_SdvpqJ9I0_1;
	wire w_dff_B_kmjw1zPo7_1;
	wire w_dff_B_9tJZEBie7_1;
	wire w_dff_B_ZL2b8DO29_1;
	wire w_dff_B_Oytvunn13_1;
	wire w_dff_B_bqTIOM818_1;
	wire w_dff_B_zvgoz3Or6_1;
	wire w_dff_B_DjlqhmOH2_1;
	wire w_dff_B_HRPm5ceE0_1;
	wire w_dff_B_y0e9V7Le4_1;
	wire w_dff_B_D3sBofnd3_1;
	wire w_dff_B_bIqpzd0J6_1;
	wire w_dff_B_w46QEcus9_1;
	wire w_dff_B_VnurZ78S7_1;
	wire w_dff_B_rvsf82Hy9_1;
	wire w_dff_B_KCY6jKxL8_1;
	wire w_dff_B_neuIDJ094_1;
	wire w_dff_B_LLlnUf0X8_1;
	wire w_dff_B_XnIRbzHe1_1;
	wire w_dff_B_GlfsU0pY0_1;
	wire w_dff_B_HkvM7tUT2_1;
	wire w_dff_B_Jc0uU5PP2_1;
	wire w_dff_B_t8S2V3MC4_1;
	wire w_dff_B_aaEYDhan0_1;
	wire w_dff_B_pPZqv6HN4_1;
	wire w_dff_B_6Q9PEvRh8_1;
	wire w_dff_B_zwpm3GUc5_1;
	wire w_dff_B_uJWYmW7H4_1;
	wire w_dff_B_NZk7PCDX8_1;
	wire w_dff_B_7EzHJnX21_1;
	wire w_dff_B_cqLup7jz7_1;
	wire w_dff_B_P6j9Uit05_1;
	wire w_dff_B_yjodbsVS4_1;
	wire w_dff_B_HJUaiY828_1;
	wire w_dff_B_qzyPgkD27_1;
	wire w_dff_B_X0uR2JGV6_1;
	wire w_dff_B_ER3U3fqg6_1;
	wire w_dff_B_OKF48mbL2_1;
	wire w_dff_B_VthZKeJx5_1;
	wire w_dff_B_BZMoRq1H3_1;
	wire w_dff_B_1556L6KT5_1;
	wire w_dff_B_rg0cl9838_1;
	wire w_dff_B_Dvmvkiei3_1;
	wire w_dff_B_dS5eIGWr2_1;
	wire w_dff_B_G9zIIImv0_1;
	wire w_dff_B_7ka1G4sx6_1;
	wire w_dff_B_KWT6pzHw7_1;
	wire w_dff_B_VpeHMeY28_1;
	wire w_dff_B_IXZHpsWX0_1;
	wire w_dff_B_XMZThkG69_1;
	wire w_dff_B_OJU6tlcr3_1;
	wire w_dff_B_2FY1RBD26_1;
	wire w_dff_B_XUKOerNr6_1;
	wire w_dff_B_cSjM4ZjR3_1;
	wire w_dff_B_xiwPHwZO0_1;
	wire w_dff_B_rmy2HHye7_1;
	wire w_dff_B_4A1CkX5B4_1;
	wire w_dff_B_vbbWAHtj0_1;
	wire w_dff_B_smF1nojO0_1;
	wire w_dff_B_57FFLbto4_1;
	wire w_dff_B_C2Y1m1Yv7_1;
	wire w_dff_B_wtrTuE9s1_1;
	wire w_dff_B_7V0Zc7gS5_1;
	wire w_dff_B_fRWjVBnI8_1;
	wire w_dff_B_svFv9JXO5_1;
	wire w_dff_B_UIKRhfJj1_1;
	wire w_dff_B_lfWYUkE89_1;
	wire w_dff_B_jz0eAxfA5_1;
	wire w_dff_B_p5Y4LAwZ6_1;
	wire w_dff_B_4ZXn5FRc7_1;
	wire w_dff_B_fNWVTgnR3_1;
	wire w_dff_B_yXHeBq5g7_1;
	wire w_dff_B_tvjawTBP1_1;
	wire w_dff_B_G5qkCL0X7_0;
	wire w_dff_B_W0Qjtbz47_0;
	wire w_dff_B_FrTXzQKt6_0;
	wire w_dff_B_85UZipWH4_0;
	wire w_dff_B_Qwhn3Ko87_0;
	wire w_dff_B_cKlewMrP2_0;
	wire w_dff_B_LjzyfdRH7_0;
	wire w_dff_B_ZXyzgNCw8_0;
	wire w_dff_B_6uLSzrLn5_0;
	wire w_dff_B_Sr54sdTA5_0;
	wire w_dff_B_AyMcy5ei3_0;
	wire w_dff_B_JLvX7JJU4_0;
	wire w_dff_B_bBz64bGA2_0;
	wire w_dff_B_pKhh7Bse3_0;
	wire w_dff_B_QMFevvUf8_0;
	wire w_dff_B_ixUx4s6R0_0;
	wire w_dff_B_e4ioJ66S3_0;
	wire w_dff_B_mcwjGYuR6_0;
	wire w_dff_B_W2uRE0Cp8_0;
	wire w_dff_B_e3df2hCj1_0;
	wire w_dff_B_WWMhl39V7_0;
	wire w_dff_B_KuPQB4Se4_0;
	wire w_dff_B_cCXIpIxk5_0;
	wire w_dff_B_j3AMZp8F3_0;
	wire w_dff_B_Qy23gWSG3_0;
	wire w_dff_B_8ZKhRNLZ9_0;
	wire w_dff_B_2IFjmLoA3_0;
	wire w_dff_B_HWP9ru513_0;
	wire w_dff_B_0CdQbKA81_0;
	wire w_dff_B_tHPKEO575_0;
	wire w_dff_B_snBOq5kJ0_0;
	wire w_dff_B_oTZTnS232_0;
	wire w_dff_B_lAezKzTq6_0;
	wire w_dff_B_pQvZFp9X9_0;
	wire w_dff_B_yqLXZtf07_0;
	wire w_dff_B_fhzR3x2f4_0;
	wire w_dff_B_PZZ92WMf6_0;
	wire w_dff_B_xV5VhJBE8_0;
	wire w_dff_B_udSN2HBo6_0;
	wire w_dff_B_UznRq11J3_0;
	wire w_dff_B_UwRvC1K20_0;
	wire w_dff_B_E6zqEYfG2_0;
	wire w_dff_B_vAcTpdOW4_0;
	wire w_dff_B_pdYnTYPI3_0;
	wire w_dff_B_4NhGbutW7_0;
	wire w_dff_B_xKT1u53Y9_0;
	wire w_dff_B_bgmYoS3D8_0;
	wire w_dff_B_K9nWt2Yx3_0;
	wire w_dff_B_zzyP0Zp78_0;
	wire w_dff_B_Izliwfpz0_0;
	wire w_dff_B_s2TekWhD5_0;
	wire w_dff_B_zucnam1y8_0;
	wire w_dff_B_7zs0lD3d3_0;
	wire w_dff_B_fU7zMoX06_0;
	wire w_dff_B_ql6LDvXf6_0;
	wire w_dff_B_G3bu3MRX2_0;
	wire w_dff_B_VCVnfmzm3_0;
	wire w_dff_B_TPK0c9xf2_0;
	wire w_dff_B_nlsQP6292_0;
	wire w_dff_B_WAmrd0AY3_0;
	wire w_dff_B_vVMEnPU32_0;
	wire w_dff_B_xQkZ1Kwc9_0;
	wire w_dff_B_CnnuCVmE3_0;
	wire w_dff_B_bCsX3cDJ5_0;
	wire w_dff_B_41grjv8w0_0;
	wire w_dff_B_cudNGoO26_0;
	wire w_dff_B_chimribU5_0;
	wire w_dff_B_UHzd7LdG8_0;
	wire w_dff_B_3wWRXdiY2_0;
	wire w_dff_B_xbj2Qh1V4_0;
	wire w_dff_B_UnoDeeOr7_0;
	wire w_dff_B_tCwpCsJa9_0;
	wire w_dff_B_pCwSTHxS9_0;
	wire w_dff_B_Tfa6iLBB6_0;
	wire w_dff_B_JCmdtD7q6_0;
	wire w_dff_B_FIzmcAae6_0;
	wire w_dff_B_WYMQiob36_0;
	wire w_dff_B_anDCubS42_0;
	wire w_dff_B_PygIc9OI4_0;
	wire w_dff_B_nSy1uQnu2_0;
	wire w_dff_B_JvDs4JAs1_0;
	wire w_dff_B_1fNWwNfy0_1;
	wire w_dff_B_0hMFpWJF4_1;
	wire w_dff_B_ohVW7VIx3_1;
	wire w_dff_B_bojFVHxi6_1;
	wire w_dff_B_U1RRFvWX4_1;
	wire w_dff_B_k6RWaLjO8_1;
	wire w_dff_B_kwOVKXfA7_1;
	wire w_dff_B_5UzRbjzr2_1;
	wire w_dff_B_FODG8SnM9_1;
	wire w_dff_B_e6TUD5kF7_1;
	wire w_dff_B_3ahSLU0f5_1;
	wire w_dff_B_GIKKA03y8_1;
	wire w_dff_B_SS6WDjzM5_1;
	wire w_dff_B_cWw19qAf3_1;
	wire w_dff_B_BFNjEJig8_1;
	wire w_dff_B_Kjp1X3wj4_1;
	wire w_dff_B_yxCjC1Eo5_1;
	wire w_dff_B_SeajZeG01_1;
	wire w_dff_B_1brRFTAQ7_1;
	wire w_dff_B_jVBvabbt5_1;
	wire w_dff_B_1ZYustJz1_1;
	wire w_dff_B_YVdG32KG6_1;
	wire w_dff_B_P6WDcFKN9_1;
	wire w_dff_B_IGqHtOAZ5_1;
	wire w_dff_B_oCAn17SR0_1;
	wire w_dff_B_KXbAAbK76_1;
	wire w_dff_B_pwEezPyR0_1;
	wire w_dff_B_A5znvr275_1;
	wire w_dff_B_VXehlGKy3_1;
	wire w_dff_B_EdIecont7_1;
	wire w_dff_B_tx1DN6rz5_1;
	wire w_dff_B_fnIfyBF51_1;
	wire w_dff_B_bAT882n93_1;
	wire w_dff_B_OhRJB9ro3_1;
	wire w_dff_B_cZfPFW8I5_1;
	wire w_dff_B_DQG9O0KZ1_1;
	wire w_dff_B_pRpKWNyO9_1;
	wire w_dff_B_aWFkOS0o6_1;
	wire w_dff_B_dRiK9Ukz0_1;
	wire w_dff_B_cduITGCM4_1;
	wire w_dff_B_gqbX7jdF0_1;
	wire w_dff_B_hFQT1YAU5_1;
	wire w_dff_B_hkJ3ShXI0_1;
	wire w_dff_B_5vb6oOpc8_1;
	wire w_dff_B_nZg0GdcQ2_1;
	wire w_dff_B_EFlFV7KA5_1;
	wire w_dff_B_FSmo0P7R4_1;
	wire w_dff_B_3J7wgZMo8_1;
	wire w_dff_B_sYvKG95B8_1;
	wire w_dff_B_YJaQeKRC6_1;
	wire w_dff_B_ZxSgdjvF3_1;
	wire w_dff_B_eLDVdvK05_1;
	wire w_dff_B_leSJa8mv3_1;
	wire w_dff_B_emB1c9tb6_1;
	wire w_dff_B_ovrDLKBA1_1;
	wire w_dff_B_CSf3cnQF3_1;
	wire w_dff_B_qWbXoKNO7_1;
	wire w_dff_B_ODxQMLDb6_1;
	wire w_dff_B_ZwTNwGA55_1;
	wire w_dff_B_R3xUGviu9_1;
	wire w_dff_B_EN1NQcku8_1;
	wire w_dff_B_1LGb7X9i6_1;
	wire w_dff_B_y4Vxv6FO7_1;
	wire w_dff_B_csX0uRYy5_1;
	wire w_dff_B_mFe7Unt29_1;
	wire w_dff_B_WAZikE3v7_1;
	wire w_dff_B_8tIQy2SM3_1;
	wire w_dff_B_1S442Ar52_1;
	wire w_dff_B_aj23fqra7_1;
	wire w_dff_B_8SQNheKS0_1;
	wire w_dff_B_nviS5O506_1;
	wire w_dff_B_eIl5V82O6_1;
	wire w_dff_B_3pOx5mzZ5_1;
	wire w_dff_B_w3vnM6zc0_1;
	wire w_dff_B_5SuKWVLd3_1;
	wire w_dff_B_PDF1HE6X2_1;
	wire w_dff_B_xD6nLRAA9_1;
	wire w_dff_B_5Zwwjfqu1_1;
	wire w_dff_B_nRpberWk8_1;
	wire w_dff_B_e84DdMJl5_1;
	wire w_dff_B_LA8nUIhW1_0;
	wire w_dff_B_UlwaVDyo4_0;
	wire w_dff_B_WsGbYJHm5_0;
	wire w_dff_B_joZJAjTz7_0;
	wire w_dff_B_bGHwirTb0_0;
	wire w_dff_B_sjPjaM7I3_0;
	wire w_dff_B_uA4c2xIE5_0;
	wire w_dff_B_5EoqFvgV4_0;
	wire w_dff_B_ohalHl3I7_0;
	wire w_dff_B_VuRCtj7r9_0;
	wire w_dff_B_93txWX9V4_0;
	wire w_dff_B_fjicCr5Z6_0;
	wire w_dff_B_mGafTpnt9_0;
	wire w_dff_B_hOdSlX2K2_0;
	wire w_dff_B_BusYKFN71_0;
	wire w_dff_B_yJ07B1S13_0;
	wire w_dff_B_07V96llp4_0;
	wire w_dff_B_hjFWNCWA7_0;
	wire w_dff_B_SOpCPN7r2_0;
	wire w_dff_B_FTtsVcvj6_0;
	wire w_dff_B_EtWZMNfG2_0;
	wire w_dff_B_L677Jlfv4_0;
	wire w_dff_B_sZfXbixm5_0;
	wire w_dff_B_IPzOYziY9_0;
	wire w_dff_B_1XvA1Jmo0_0;
	wire w_dff_B_9gBZcg8H3_0;
	wire w_dff_B_12hH4dGZ5_0;
	wire w_dff_B_7LbisSyT2_0;
	wire w_dff_B_mtPh5xJ10_0;
	wire w_dff_B_FPDXdtsm1_0;
	wire w_dff_B_07N54mPD2_0;
	wire w_dff_B_gJ0yOhSL0_0;
	wire w_dff_B_R6xK6GA07_0;
	wire w_dff_B_Nz9McD6Q8_0;
	wire w_dff_B_tsPwY25c3_0;
	wire w_dff_B_Sa3VBwqB5_0;
	wire w_dff_B_QPv0mvlg0_0;
	wire w_dff_B_eO1IIRFA4_0;
	wire w_dff_B_S1UjzQh42_0;
	wire w_dff_B_N5ROz9rz6_0;
	wire w_dff_B_eFnN80HK4_0;
	wire w_dff_B_O5e8Amcy6_0;
	wire w_dff_B_VD38JG0M7_0;
	wire w_dff_B_mEcvTa2v6_0;
	wire w_dff_B_MvVy2GtC7_0;
	wire w_dff_B_BMZ9kfZd3_0;
	wire w_dff_B_EISWj2oM1_0;
	wire w_dff_B_BzdIBGA48_0;
	wire w_dff_B_iSM6W20w8_0;
	wire w_dff_B_sogyuxOg0_0;
	wire w_dff_B_VE8BkZXE0_0;
	wire w_dff_B_cpt6ZdiB9_0;
	wire w_dff_B_8Ywpla247_0;
	wire w_dff_B_CHNqhXo22_0;
	wire w_dff_B_DsBOklLR6_0;
	wire w_dff_B_fVhNd03m0_0;
	wire w_dff_B_inBtQ2Fh1_0;
	wire w_dff_B_LvRMYlsV7_0;
	wire w_dff_B_mWZPlMUn1_0;
	wire w_dff_B_FG0yEm768_0;
	wire w_dff_B_Wgklik3i7_0;
	wire w_dff_B_e4ZRLmT65_0;
	wire w_dff_B_uc4EemAt8_0;
	wire w_dff_B_v62cHd8i6_0;
	wire w_dff_B_8bZh3vep5_0;
	wire w_dff_B_IN6Z1lU39_0;
	wire w_dff_B_xO2ENmm82_0;
	wire w_dff_B_bc4YtK6Z7_0;
	wire w_dff_B_YhHx2WQc0_0;
	wire w_dff_B_JSwaYugR5_0;
	wire w_dff_B_XRyY7pT98_0;
	wire w_dff_B_sKB8gmvT8_0;
	wire w_dff_B_VaegOeAt7_0;
	wire w_dff_B_gXkYNe7n9_0;
	wire w_dff_B_pW8kc4Be2_0;
	wire w_dff_B_tnRPek717_0;
	wire w_dff_B_ysmONgPT3_0;
	wire w_dff_B_o5w7wT8k3_0;
	wire w_dff_B_HgzYxPhY9_0;
	wire w_dff_B_MhnprG8l9_0;
	wire w_dff_B_qceRoBmQ1_1;
	wire w_dff_B_nuicdX2j0_1;
	wire w_dff_B_KhD2OBuk3_1;
	wire w_dff_B_4JJj7Ghw4_1;
	wire w_dff_B_QHMVQmaQ1_1;
	wire w_dff_B_706k3QG64_1;
	wire w_dff_B_i0ZmiZkZ5_1;
	wire w_dff_B_RWCUxv5t6_1;
	wire w_dff_B_7B9YVItL2_1;
	wire w_dff_B_oO4vhS9F3_1;
	wire w_dff_B_uEi0WiuB0_1;
	wire w_dff_B_abEnW9Zc4_1;
	wire w_dff_B_UzQodXDE8_1;
	wire w_dff_B_zPdKUbsG2_1;
	wire w_dff_B_CYJARK1g6_1;
	wire w_dff_B_Oii4CUX08_1;
	wire w_dff_B_hF4uKHVr3_1;
	wire w_dff_B_lOMYp8Kt3_1;
	wire w_dff_B_2ahuWX887_1;
	wire w_dff_B_JMGiE6G57_1;
	wire w_dff_B_TDtMm0XF1_1;
	wire w_dff_B_UWnr3xXR6_1;
	wire w_dff_B_lFTYaQDp8_1;
	wire w_dff_B_L7kOx4Gv5_1;
	wire w_dff_B_sAWqPKB59_1;
	wire w_dff_B_VzLpQoOw6_1;
	wire w_dff_B_rhEZciPG6_1;
	wire w_dff_B_fVOMApE95_1;
	wire w_dff_B_jgMf64ZO3_1;
	wire w_dff_B_FjREz1Ko1_1;
	wire w_dff_B_RWsC1hqg3_1;
	wire w_dff_B_YcC5qUWt7_1;
	wire w_dff_B_OjJcsPVX5_1;
	wire w_dff_B_rddN5v7d1_1;
	wire w_dff_B_0VDSB8Kz6_1;
	wire w_dff_B_n7bb6j482_1;
	wire w_dff_B_27vDazFn0_1;
	wire w_dff_B_cgp6ZmvE8_1;
	wire w_dff_B_PcwTg4Nf8_1;
	wire w_dff_B_q5rNOSs75_1;
	wire w_dff_B_yFqsHu4m0_1;
	wire w_dff_B_QYl9RcJo7_1;
	wire w_dff_B_zwRJYAip8_1;
	wire w_dff_B_cB6U3jUe6_1;
	wire w_dff_B_CWf4T7Q14_1;
	wire w_dff_B_YXNjCd5l2_1;
	wire w_dff_B_I7mOOrUk8_1;
	wire w_dff_B_xWYdAhSV0_1;
	wire w_dff_B_LWVgbbQf8_1;
	wire w_dff_B_ro2YST8v1_1;
	wire w_dff_B_LYP36CjP9_1;
	wire w_dff_B_FWGwVdIL3_1;
	wire w_dff_B_SZmvxS565_1;
	wire w_dff_B_osRZc0eC4_1;
	wire w_dff_B_UIZFMvfW9_1;
	wire w_dff_B_YcXqJC6S0_1;
	wire w_dff_B_w7HSpxz76_1;
	wire w_dff_B_a33IaeeV4_1;
	wire w_dff_B_kVzCrytA1_1;
	wire w_dff_B_8PC2PrYQ7_1;
	wire w_dff_B_hA6Esfvs9_1;
	wire w_dff_B_tUvVXCne1_1;
	wire w_dff_B_n8NVf91s7_1;
	wire w_dff_B_7dc5sPpq5_1;
	wire w_dff_B_ELIHhym96_1;
	wire w_dff_B_VFbNHcqM6_1;
	wire w_dff_B_xIwOwtEl0_1;
	wire w_dff_B_KFRsv0e36_1;
	wire w_dff_B_WErrMpK48_1;
	wire w_dff_B_IY6u5P0P2_1;
	wire w_dff_B_T8tVNFsk9_1;
	wire w_dff_B_HGObvQ0B4_1;
	wire w_dff_B_WmVuxury4_1;
	wire w_dff_B_rrrI6D1L4_1;
	wire w_dff_B_kWY03dVN0_1;
	wire w_dff_B_qABRW3tr6_1;
	wire w_dff_B_RYu0Dyl48_1;
	wire w_dff_B_HNvMBpKf9_1;
	wire w_dff_B_sIPXzDkp4_1;
	wire w_dff_B_C0HHHzh75_0;
	wire w_dff_B_0unVWWyq5_0;
	wire w_dff_B_DYKWDjoX2_0;
	wire w_dff_B_IYubbnKR7_0;
	wire w_dff_B_QQk97jog6_0;
	wire w_dff_B_01JquW444_0;
	wire w_dff_B_bJg4TdHi2_0;
	wire w_dff_B_qIRSSsbt1_0;
	wire w_dff_B_ahFmu9QF6_0;
	wire w_dff_B_ldvR4YwX7_0;
	wire w_dff_B_tn0WhfQ49_0;
	wire w_dff_B_aIbwPofl7_0;
	wire w_dff_B_gDq3y9cm1_0;
	wire w_dff_B_jh7p3t3W0_0;
	wire w_dff_B_Azk00dkJ0_0;
	wire w_dff_B_GkE1YKNl1_0;
	wire w_dff_B_DRBOY5cU8_0;
	wire w_dff_B_YyZ3OxUL0_0;
	wire w_dff_B_qSezP5MA4_0;
	wire w_dff_B_EwXafume2_0;
	wire w_dff_B_SidiTEaW2_0;
	wire w_dff_B_WI4iuNYk9_0;
	wire w_dff_B_gC1FqZfa3_0;
	wire w_dff_B_5dywQ92U5_0;
	wire w_dff_B_Y9gyQyNF6_0;
	wire w_dff_B_RBi06g3M8_0;
	wire w_dff_B_xYbX8bbr1_0;
	wire w_dff_B_WImmKUQa0_0;
	wire w_dff_B_i13Vv1PM3_0;
	wire w_dff_B_k4qQKCLj6_0;
	wire w_dff_B_Yd0LhWEN2_0;
	wire w_dff_B_Eej5KYxV4_0;
	wire w_dff_B_wgeHFxXT0_0;
	wire w_dff_B_LKW7eHky4_0;
	wire w_dff_B_lLoufkls1_0;
	wire w_dff_B_4rSgmUun2_0;
	wire w_dff_B_cfoVcOpw7_0;
	wire w_dff_B_2xrE3NSH1_0;
	wire w_dff_B_CcYX6sPK8_0;
	wire w_dff_B_Jwr9ud9u8_0;
	wire w_dff_B_Y05VgRx63_0;
	wire w_dff_B_tv9e17wr1_0;
	wire w_dff_B_yjmp301p1_0;
	wire w_dff_B_WFn3IAxy3_0;
	wire w_dff_B_fuOQSH5C1_0;
	wire w_dff_B_5ITfGVaQ2_0;
	wire w_dff_B_0VD5m62i0_0;
	wire w_dff_B_not8cW135_0;
	wire w_dff_B_9jvl69mj8_0;
	wire w_dff_B_4TrvZjcd5_0;
	wire w_dff_B_FSKLiabn8_0;
	wire w_dff_B_qb8zBmN64_0;
	wire w_dff_B_isw0vxTt7_0;
	wire w_dff_B_4AHxuAkV4_0;
	wire w_dff_B_SH38UfqO5_0;
	wire w_dff_B_ezIRKy3t8_0;
	wire w_dff_B_OCQCRQcb0_0;
	wire w_dff_B_05Kch9JF6_0;
	wire w_dff_B_XO7Wi3Gt8_0;
	wire w_dff_B_dOPWldWu1_0;
	wire w_dff_B_u0CkkhaS3_0;
	wire w_dff_B_SWGrBkMc8_0;
	wire w_dff_B_Y4tj5F2l3_0;
	wire w_dff_B_AVhl6SGa2_0;
	wire w_dff_B_k68Mwf0C2_0;
	wire w_dff_B_gUV6Cqb07_0;
	wire w_dff_B_uJ8bQSmx0_0;
	wire w_dff_B_EnIhzMOw3_0;
	wire w_dff_B_qNCpt48b4_0;
	wire w_dff_B_YQu8q8eu7_0;
	wire w_dff_B_QQoj9x9n2_0;
	wire w_dff_B_hccerYTj0_0;
	wire w_dff_B_cAvIqjhH2_0;
	wire w_dff_B_lvBtN87r4_0;
	wire w_dff_B_N9aWi0P60_0;
	wire w_dff_B_srqhhSHi4_0;
	wire w_dff_B_nqBuXuO03_0;
	wire w_dff_B_8VOKdXdQ9_0;
	wire w_dff_B_OkjULAnL9_0;
	wire w_dff_B_9NJgM24b5_1;
	wire w_dff_B_Ee89ZGrN4_1;
	wire w_dff_B_ZF42x9ts0_1;
	wire w_dff_B_QjswzR6b7_1;
	wire w_dff_B_Louy74bJ1_1;
	wire w_dff_B_KSXvOQt49_1;
	wire w_dff_B_vWIbbuSJ2_1;
	wire w_dff_B_FenRkLh27_1;
	wire w_dff_B_26b3Zlqq7_1;
	wire w_dff_B_Muweay6I7_1;
	wire w_dff_B_CMWFYgjn0_1;
	wire w_dff_B_j8KqCyKQ6_1;
	wire w_dff_B_sT0Hmm989_1;
	wire w_dff_B_tozgOeZS8_1;
	wire w_dff_B_Y7x8ms9G3_1;
	wire w_dff_B_bsT20mAX8_1;
	wire w_dff_B_tINAJHrN2_1;
	wire w_dff_B_zjO5cdOm8_1;
	wire w_dff_B_4DUWaUx61_1;
	wire w_dff_B_Ol3ZBT5B5_1;
	wire w_dff_B_A1uC9sbx9_1;
	wire w_dff_B_pwMQRzIi0_1;
	wire w_dff_B_mjZS1bgC8_1;
	wire w_dff_B_ysFgUrBC8_1;
	wire w_dff_B_co0ctbka3_1;
	wire w_dff_B_iS99qmpY0_1;
	wire w_dff_B_9VmRnF7I2_1;
	wire w_dff_B_t4eQxJZH6_1;
	wire w_dff_B_XwUgOE3E5_1;
	wire w_dff_B_Nm5IPIl41_1;
	wire w_dff_B_JaKKb2p29_1;
	wire w_dff_B_ICBZ6n092_1;
	wire w_dff_B_oo2OxxsJ1_1;
	wire w_dff_B_tTj9umva9_1;
	wire w_dff_B_Wy7hGWI61_1;
	wire w_dff_B_IQJhi7uQ9_1;
	wire w_dff_B_qhye2kpX3_1;
	wire w_dff_B_cVDBCvHa0_1;
	wire w_dff_B_hcdN6NNH1_1;
	wire w_dff_B_52ms6wAm9_1;
	wire w_dff_B_e8cBAJ450_1;
	wire w_dff_B_BFddvJTE7_1;
	wire w_dff_B_FsUz8bED2_1;
	wire w_dff_B_F7zOgjsA2_1;
	wire w_dff_B_ed99a9fb5_1;
	wire w_dff_B_901DdbOZ7_1;
	wire w_dff_B_NcAKWOW76_1;
	wire w_dff_B_45zR5xGK2_1;
	wire w_dff_B_O7c4UxYo3_1;
	wire w_dff_B_v0LDFqJ10_1;
	wire w_dff_B_VHa9mYIA3_1;
	wire w_dff_B_ktlZVb6b6_1;
	wire w_dff_B_CGC6woTF7_1;
	wire w_dff_B_40M3lrbG9_1;
	wire w_dff_B_EJ4RaDyY2_1;
	wire w_dff_B_PRIf5Z2A2_1;
	wire w_dff_B_qCgnp5tw7_1;
	wire w_dff_B_2WZarVJq6_1;
	wire w_dff_B_Lg6v5lBM4_1;
	wire w_dff_B_s43XP0Le3_1;
	wire w_dff_B_wfRhvxgL3_1;
	wire w_dff_B_TndS5KXC9_1;
	wire w_dff_B_r8PlXZlq0_1;
	wire w_dff_B_UuuzylPH3_1;
	wire w_dff_B_zftX87tM0_1;
	wire w_dff_B_bbA0ckeX8_1;
	wire w_dff_B_HlBBpU5P9_1;
	wire w_dff_B_jfFDA3w71_1;
	wire w_dff_B_15P4j7GD1_1;
	wire w_dff_B_u8RZ4i7D2_1;
	wire w_dff_B_jtXBEZHH1_1;
	wire w_dff_B_rg7QbqaU7_1;
	wire w_dff_B_kAeLitOl4_1;
	wire w_dff_B_TejR0zQI9_1;
	wire w_dff_B_xdTQ0fQL4_1;
	wire w_dff_B_CQwcGSaj4_1;
	wire w_dff_B_Amfob1qH1_1;
	wire w_dff_B_PPpQ5mdn1_1;
	wire w_dff_B_AKYzejYo5_0;
	wire w_dff_B_7IDtgNJk7_0;
	wire w_dff_B_8HrLto0e2_0;
	wire w_dff_B_JpX2n4bg1_0;
	wire w_dff_B_IaEbr7209_0;
	wire w_dff_B_nSyI0P9w4_0;
	wire w_dff_B_vrUairEN8_0;
	wire w_dff_B_wcO3udsH0_0;
	wire w_dff_B_QMIJgd9Z3_0;
	wire w_dff_B_olCUdMbx8_0;
	wire w_dff_B_vOpYVEes8_0;
	wire w_dff_B_Mj2dEgYd3_0;
	wire w_dff_B_ZdScPvL71_0;
	wire w_dff_B_mtYlnKgr1_0;
	wire w_dff_B_eMSlw0Pt4_0;
	wire w_dff_B_MaRdwAHT1_0;
	wire w_dff_B_ZmpmK7St6_0;
	wire w_dff_B_VaDQCl2Y8_0;
	wire w_dff_B_KvghZkei9_0;
	wire w_dff_B_gi1vx5sq4_0;
	wire w_dff_B_7EnuHvxh9_0;
	wire w_dff_B_qwhUHJDk8_0;
	wire w_dff_B_xpLm7AOd1_0;
	wire w_dff_B_37slPqMN9_0;
	wire w_dff_B_gtWRKnly7_0;
	wire w_dff_B_gECJYpll1_0;
	wire w_dff_B_I4muCoFR5_0;
	wire w_dff_B_3Vo90gVp6_0;
	wire w_dff_B_J97ykhr25_0;
	wire w_dff_B_lhCECIPs9_0;
	wire w_dff_B_Af5AdqYE5_0;
	wire w_dff_B_p88eS73Q0_0;
	wire w_dff_B_H7hjs9Kc4_0;
	wire w_dff_B_gkb9CDrm3_0;
	wire w_dff_B_aIyQQONY1_0;
	wire w_dff_B_HrQm4c5a8_0;
	wire w_dff_B_wvS1Pqwl2_0;
	wire w_dff_B_oYJAh0cj9_0;
	wire w_dff_B_gDE3kUwP1_0;
	wire w_dff_B_IpocvKzj5_0;
	wire w_dff_B_hMYQshit6_0;
	wire w_dff_B_vvfUGRbh0_0;
	wire w_dff_B_stdu2BJX2_0;
	wire w_dff_B_4rpeBBVQ0_0;
	wire w_dff_B_hEZrfaVQ7_0;
	wire w_dff_B_dk8Gjgog4_0;
	wire w_dff_B_i2eCqOGc5_0;
	wire w_dff_B_BolPvYss6_0;
	wire w_dff_B_uoqHmwnq3_0;
	wire w_dff_B_iMLRkoUN5_0;
	wire w_dff_B_QIBLQZZa0_0;
	wire w_dff_B_bFJKcIP87_0;
	wire w_dff_B_lhZFRcmq9_0;
	wire w_dff_B_z6rvqgCH2_0;
	wire w_dff_B_oQcsgDTN6_0;
	wire w_dff_B_qPjFxPqP6_0;
	wire w_dff_B_cfFdhhoE2_0;
	wire w_dff_B_18yjfYTz5_0;
	wire w_dff_B_jsRJJOYz8_0;
	wire w_dff_B_5xgLIorn9_0;
	wire w_dff_B_mmH7ljqM2_0;
	wire w_dff_B_qA1OOnNy6_0;
	wire w_dff_B_QcxskTGc8_0;
	wire w_dff_B_MPlmTR1w1_0;
	wire w_dff_B_seD2LrPD7_0;
	wire w_dff_B_2s0OEdS27_0;
	wire w_dff_B_4OOlJfPb9_0;
	wire w_dff_B_sE3eZfIE4_0;
	wire w_dff_B_whJyrNNb9_0;
	wire w_dff_B_fgDz39rj3_0;
	wire w_dff_B_c5MKNbQr9_0;
	wire w_dff_B_1dUNJKul3_0;
	wire w_dff_B_vSJ6okrh6_0;
	wire w_dff_B_7HOhPr9F3_0;
	wire w_dff_B_eDTMfV4R7_0;
	wire w_dff_B_7OfKxHUE9_0;
	wire w_dff_B_OAi2xSZU9_0;
	wire w_dff_B_nx8MnoHd2_0;
	wire w_dff_B_lCknWwrj8_1;
	wire w_dff_B_xZsUVpB96_1;
	wire w_dff_B_OdyCepR85_1;
	wire w_dff_B_TdQA974I2_1;
	wire w_dff_B_1OLK7WvQ2_1;
	wire w_dff_B_QRCLJIzF2_1;
	wire w_dff_B_zgky6dEv8_1;
	wire w_dff_B_FGEnxrmt2_1;
	wire w_dff_B_iHU1lMPN3_1;
	wire w_dff_B_JdgEoIGi3_1;
	wire w_dff_B_vbCn5soC4_1;
	wire w_dff_B_pwwNt5c28_1;
	wire w_dff_B_ROq1uc8L7_1;
	wire w_dff_B_MurowAlE7_1;
	wire w_dff_B_6XfR9vIt1_1;
	wire w_dff_B_WXvnlxJT5_1;
	wire w_dff_B_yaRblRQ46_1;
	wire w_dff_B_DIohpfQV5_1;
	wire w_dff_B_YvKgTTZQ7_1;
	wire w_dff_B_kG1QNLdi9_1;
	wire w_dff_B_sXuXqJmA8_1;
	wire w_dff_B_iNq0GzVs2_1;
	wire w_dff_B_fXK9lR2Q4_1;
	wire w_dff_B_LvndWEaJ3_1;
	wire w_dff_B_H74PVpH53_1;
	wire w_dff_B_8qyhmj779_1;
	wire w_dff_B_LlZHsgZg7_1;
	wire w_dff_B_vnR7Vhd15_1;
	wire w_dff_B_hJS2rmOb2_1;
	wire w_dff_B_lPCprq4y1_1;
	wire w_dff_B_JwWZkULi6_1;
	wire w_dff_B_T1QzJsnp7_1;
	wire w_dff_B_yuMrqQsK6_1;
	wire w_dff_B_hFX3SBAr1_1;
	wire w_dff_B_VvxhphEV2_1;
	wire w_dff_B_KP6iEftl2_1;
	wire w_dff_B_wHB3vvVW5_1;
	wire w_dff_B_bQ9tjdIx0_1;
	wire w_dff_B_rXxfZgr74_1;
	wire w_dff_B_0l0nvwRK1_1;
	wire w_dff_B_knOUVsni5_1;
	wire w_dff_B_ANDRZreF6_1;
	wire w_dff_B_it1pg5m83_1;
	wire w_dff_B_T6y7wXMy3_1;
	wire w_dff_B_eUYgLd0Z4_1;
	wire w_dff_B_Q01jJjEK7_1;
	wire w_dff_B_jI1RE9so4_1;
	wire w_dff_B_uQNoylBf7_1;
	wire w_dff_B_i6FkjAbK9_1;
	wire w_dff_B_jKzmRNqQ0_1;
	wire w_dff_B_4FQAICTw7_1;
	wire w_dff_B_nYL3Nx2S9_1;
	wire w_dff_B_WENE3vIV8_1;
	wire w_dff_B_qxrqIai26_1;
	wire w_dff_B_EffnkreD7_1;
	wire w_dff_B_QNB56xWq6_1;
	wire w_dff_B_r5AYdCqd9_1;
	wire w_dff_B_2YAzXdR91_1;
	wire w_dff_B_cMVQaYHH7_1;
	wire w_dff_B_Qyq5nCpg1_1;
	wire w_dff_B_3sp0g04m1_1;
	wire w_dff_B_tpDNhVmN3_1;
	wire w_dff_B_WYLn8ZGZ6_1;
	wire w_dff_B_GYHJmo1p7_1;
	wire w_dff_B_BDprvJWN4_1;
	wire w_dff_B_o8C8aFx62_1;
	wire w_dff_B_gYgMndHP4_1;
	wire w_dff_B_2iKCVqqj6_1;
	wire w_dff_B_IDPg7c2D3_1;
	wire w_dff_B_UrHN7OS58_1;
	wire w_dff_B_tKxokccA5_1;
	wire w_dff_B_9jxuSUNa7_1;
	wire w_dff_B_GCQ35GD83_1;
	wire w_dff_B_EBMD30yN5_1;
	wire w_dff_B_oI973qly7_1;
	wire w_dff_B_jqQA2aqk2_1;
	wire w_dff_B_HA2BJTtt9_1;
	wire w_dff_B_8pR5AibF7_0;
	wire w_dff_B_PTgSigU62_0;
	wire w_dff_B_XbVtRYNq9_0;
	wire w_dff_B_Rt1ZJNqG2_0;
	wire w_dff_B_vbS1gE4f5_0;
	wire w_dff_B_ezEXvfl51_0;
	wire w_dff_B_d37Hi4Od5_0;
	wire w_dff_B_IO1WzdKW2_0;
	wire w_dff_B_SEyXEGbi5_0;
	wire w_dff_B_888l08rT3_0;
	wire w_dff_B_1irBXwd25_0;
	wire w_dff_B_Lvej4ssC6_0;
	wire w_dff_B_j8jljDa79_0;
	wire w_dff_B_3RhFFOSC6_0;
	wire w_dff_B_4JDAeqte3_0;
	wire w_dff_B_iWkEtxVz3_0;
	wire w_dff_B_yaX44PMA7_0;
	wire w_dff_B_k3pIdAEr1_0;
	wire w_dff_B_LD2sgsV22_0;
	wire w_dff_B_ufiDitnS4_0;
	wire w_dff_B_OhJ9YZ951_0;
	wire w_dff_B_74CaXz5Z5_0;
	wire w_dff_B_DOQQAgLu4_0;
	wire w_dff_B_dsp8lnif5_0;
	wire w_dff_B_aAp71gpb7_0;
	wire w_dff_B_T0LA9Nw03_0;
	wire w_dff_B_10nzDHj67_0;
	wire w_dff_B_DahEASI98_0;
	wire w_dff_B_C5OsTMEn8_0;
	wire w_dff_B_bLvUkQ5E1_0;
	wire w_dff_B_afsvWgQ33_0;
	wire w_dff_B_KXhgsZnd3_0;
	wire w_dff_B_x37VCLaJ0_0;
	wire w_dff_B_fjmfZY1A0_0;
	wire w_dff_B_In4uh2SE9_0;
	wire w_dff_B_fH5HQvAi4_0;
	wire w_dff_B_dVSyXFwA2_0;
	wire w_dff_B_F18WAuQ17_0;
	wire w_dff_B_RxYBCtvV6_0;
	wire w_dff_B_DeLRJMnl2_0;
	wire w_dff_B_BaBZuiMe0_0;
	wire w_dff_B_zFfxEav43_0;
	wire w_dff_B_cKbfnsVF5_0;
	wire w_dff_B_QoErXhUF6_0;
	wire w_dff_B_ab9VWgkK0_0;
	wire w_dff_B_3NTnxzKy3_0;
	wire w_dff_B_lMaiTyyr7_0;
	wire w_dff_B_tRYKaLhl0_0;
	wire w_dff_B_XIlI9xkP5_0;
	wire w_dff_B_RSF77Hhi8_0;
	wire w_dff_B_jqJrSM7f2_0;
	wire w_dff_B_MRsiVjKc1_0;
	wire w_dff_B_ZXbgPzE16_0;
	wire w_dff_B_odyB82xQ8_0;
	wire w_dff_B_Jm9rZfzg2_0;
	wire w_dff_B_E3fYC9Lc7_0;
	wire w_dff_B_OZmjox1e6_0;
	wire w_dff_B_0DRsR5bf0_0;
	wire w_dff_B_ktgXCOXu0_0;
	wire w_dff_B_IbSg46bX1_0;
	wire w_dff_B_QBBQkVIG8_0;
	wire w_dff_B_J6L1RD5k0_0;
	wire w_dff_B_uzcBvMxk0_0;
	wire w_dff_B_JKpHx7LD2_0;
	wire w_dff_B_ma2r9Cls1_0;
	wire w_dff_B_kgpuzd063_0;
	wire w_dff_B_h483iYpH0_0;
	wire w_dff_B_LDmWxb6H9_0;
	wire w_dff_B_sZwG3PZS6_0;
	wire w_dff_B_K19q3U5j0_0;
	wire w_dff_B_SfYFSYlY8_0;
	wire w_dff_B_0At1ML9x5_0;
	wire w_dff_B_4vR1Fg8b0_0;
	wire w_dff_B_y4cCk3QS7_0;
	wire w_dff_B_kjQazQ2J0_0;
	wire w_dff_B_tFfMyx684_0;
	wire w_dff_B_tkkHea3i0_0;
	wire w_dff_B_vWkwsoob5_1;
	wire w_dff_B_kHKmM3Us2_1;
	wire w_dff_B_QuhYpKCW9_1;
	wire w_dff_B_LALH7kbx2_1;
	wire w_dff_B_M6b94v5q0_1;
	wire w_dff_B_dIFwdDTK5_1;
	wire w_dff_B_cyp5PYob1_1;
	wire w_dff_B_AC1l9Bnu7_1;
	wire w_dff_B_UNxvzmta7_1;
	wire w_dff_B_dwMsz9xw0_1;
	wire w_dff_B_pX2UXhnk6_1;
	wire w_dff_B_pzGV0cx13_1;
	wire w_dff_B_Tr32mQqt8_1;
	wire w_dff_B_Qzrdw8Sa6_1;
	wire w_dff_B_PdTKADZr3_1;
	wire w_dff_B_gM71vmhI7_1;
	wire w_dff_B_Rhwm3rHQ4_1;
	wire w_dff_B_OWsBmfZN5_1;
	wire w_dff_B_iD3D3xJB5_1;
	wire w_dff_B_ThbPfWDJ1_1;
	wire w_dff_B_UKXhGR6F1_1;
	wire w_dff_B_5kQ52v5b1_1;
	wire w_dff_B_PenMa5rR3_1;
	wire w_dff_B_t7zXDa3p1_1;
	wire w_dff_B_u732Smtf0_1;
	wire w_dff_B_td6gkA3P9_1;
	wire w_dff_B_URAlXzOj5_1;
	wire w_dff_B_wLs0cD850_1;
	wire w_dff_B_EcA06yZa4_1;
	wire w_dff_B_Dsiq8tRm8_1;
	wire w_dff_B_5RzThljG4_1;
	wire w_dff_B_iD28wjrw3_1;
	wire w_dff_B_nt5ccctD4_1;
	wire w_dff_B_bWOW1rZQ6_1;
	wire w_dff_B_9Vz53FNo6_1;
	wire w_dff_B_TFANf9cN6_1;
	wire w_dff_B_74ruwPTI7_1;
	wire w_dff_B_8UFPFhdU6_1;
	wire w_dff_B_qVFtB9gW4_1;
	wire w_dff_B_E8ov80fE0_1;
	wire w_dff_B_saiEfAmf8_1;
	wire w_dff_B_yVTKt6Cz2_1;
	wire w_dff_B_YLArECpI4_1;
	wire w_dff_B_dmi9TOxo7_1;
	wire w_dff_B_W2j8eTxx6_1;
	wire w_dff_B_XB4D5V0k0_1;
	wire w_dff_B_1ir5ZE9B3_1;
	wire w_dff_B_8fEKguUf5_1;
	wire w_dff_B_Q2SbXHbd3_1;
	wire w_dff_B_jMQM2M6y5_1;
	wire w_dff_B_nzRnGZpe3_1;
	wire w_dff_B_ReEGW0oi9_1;
	wire w_dff_B_K5gh1g9W8_1;
	wire w_dff_B_vgk24bdc8_1;
	wire w_dff_B_i4rzaCrW7_1;
	wire w_dff_B_NdjYAE8v1_1;
	wire w_dff_B_hqtRGZx85_1;
	wire w_dff_B_jpfjsvFt6_1;
	wire w_dff_B_aypb6kBz2_1;
	wire w_dff_B_PkxuWRtq7_1;
	wire w_dff_B_c8JM0jut5_1;
	wire w_dff_B_PBpMSWtP2_1;
	wire w_dff_B_AmIYtOuT1_1;
	wire w_dff_B_dI38pliI1_1;
	wire w_dff_B_EayRjbrE3_1;
	wire w_dff_B_RWW4oKsi1_1;
	wire w_dff_B_cDBqrpOP5_1;
	wire w_dff_B_D8ukmdFy4_1;
	wire w_dff_B_W8Vmw1lW3_1;
	wire w_dff_B_JlLdtDBr9_1;
	wire w_dff_B_GyjGYEKW3_1;
	wire w_dff_B_SSsgMMn53_1;
	wire w_dff_B_1BfijTHY6_1;
	wire w_dff_B_B2QvJI0J3_1;
	wire w_dff_B_7CxKjaeA3_1;
	wire w_dff_B_NwsfVLEn3_1;
	wire w_dff_B_xhrH6Nm59_0;
	wire w_dff_B_IIVCRSfT9_0;
	wire w_dff_B_Vz75Hc9N1_0;
	wire w_dff_B_ryUncve94_0;
	wire w_dff_B_fzwsv5Ng7_0;
	wire w_dff_B_02ur9dbA6_0;
	wire w_dff_B_Ukbytt5a0_0;
	wire w_dff_B_upfwbd9v5_0;
	wire w_dff_B_jVU0m9z81_0;
	wire w_dff_B_m6jinLyX8_0;
	wire w_dff_B_q3f2w4hW9_0;
	wire w_dff_B_EelgDfDz9_0;
	wire w_dff_B_YWDRUUir3_0;
	wire w_dff_B_2jGsQFbT9_0;
	wire w_dff_B_FFxz1r686_0;
	wire w_dff_B_LjfOJKfn9_0;
	wire w_dff_B_bhF2X3nJ8_0;
	wire w_dff_B_q78C42SI4_0;
	wire w_dff_B_ZTfgykT46_0;
	wire w_dff_B_MFr8crzT2_0;
	wire w_dff_B_C5Pddw0X6_0;
	wire w_dff_B_Qw0Yx3lN7_0;
	wire w_dff_B_yZ4UumJW5_0;
	wire w_dff_B_t9XNvqfh7_0;
	wire w_dff_B_Naen5Ig93_0;
	wire w_dff_B_iJ5WC9Jq0_0;
	wire w_dff_B_SLGAKHsB9_0;
	wire w_dff_B_6Ays6BV72_0;
	wire w_dff_B_h98fre8B9_0;
	wire w_dff_B_M0PymkID7_0;
	wire w_dff_B_8VV1FZOi7_0;
	wire w_dff_B_npTNlMOa8_0;
	wire w_dff_B_cUMyGulG0_0;
	wire w_dff_B_o8G2JyCb5_0;
	wire w_dff_B_myRu39ur8_0;
	wire w_dff_B_xZA5tJ8K2_0;
	wire w_dff_B_61J9Poug7_0;
	wire w_dff_B_2baMkR5X5_0;
	wire w_dff_B_SshvMVj89_0;
	wire w_dff_B_X2z7ayJJ8_0;
	wire w_dff_B_Yg0dPY2j1_0;
	wire w_dff_B_2G52tnv12_0;
	wire w_dff_B_0hAfMPkm1_0;
	wire w_dff_B_rD9euaHI7_0;
	wire w_dff_B_hEsduBhp0_0;
	wire w_dff_B_V7sCtpSY6_0;
	wire w_dff_B_qOv9yfU77_0;
	wire w_dff_B_PoNosoNN3_0;
	wire w_dff_B_lIBmC1Rw9_0;
	wire w_dff_B_t16Darf14_0;
	wire w_dff_B_0han21e32_0;
	wire w_dff_B_q0Txbzls2_0;
	wire w_dff_B_bd2CmCoH1_0;
	wire w_dff_B_DFh0NfmB0_0;
	wire w_dff_B_0ACsdpkW0_0;
	wire w_dff_B_OSkzEPVq1_0;
	wire w_dff_B_IGcDcHAI4_0;
	wire w_dff_B_IhMaCvDh6_0;
	wire w_dff_B_dySYdNLk3_0;
	wire w_dff_B_q5toYGPF8_0;
	wire w_dff_B_gaqWYEvY9_0;
	wire w_dff_B_WE0qIHoN2_0;
	wire w_dff_B_X4w4jAka2_0;
	wire w_dff_B_0r5nbhGq5_0;
	wire w_dff_B_en0bcXGN9_0;
	wire w_dff_B_F4xZ3c6h7_0;
	wire w_dff_B_ViVPGS8l2_0;
	wire w_dff_B_l0Yf07rA0_0;
	wire w_dff_B_B5LtcFVG6_0;
	wire w_dff_B_vRbftr4M2_0;
	wire w_dff_B_pC7rqyHu3_0;
	wire w_dff_B_hlndAAMl5_0;
	wire w_dff_B_qozOIvyD4_0;
	wire w_dff_B_XAE10I893_0;
	wire w_dff_B_SeDS6H6O2_0;
	wire w_dff_B_ogHkkQPV9_0;
	wire w_dff_B_fHBzS1Qj2_1;
	wire w_dff_B_GRopQDNe2_1;
	wire w_dff_B_mHqdaL8S5_1;
	wire w_dff_B_NkKEE4hf8_1;
	wire w_dff_B_5HJd2Ywu1_1;
	wire w_dff_B_0V7iFQOI8_1;
	wire w_dff_B_yzYSvzCT6_1;
	wire w_dff_B_J5V2NcVn0_1;
	wire w_dff_B_iG1sVmlX9_1;
	wire w_dff_B_aaq4mC4U7_1;
	wire w_dff_B_Pz9yoNB81_1;
	wire w_dff_B_5htoz7wO1_1;
	wire w_dff_B_IMRkCq3l5_1;
	wire w_dff_B_jfHSZsx56_1;
	wire w_dff_B_SqclJWp48_1;
	wire w_dff_B_keN5G0ag7_1;
	wire w_dff_B_pEHqStHt6_1;
	wire w_dff_B_Fpis1flx9_1;
	wire w_dff_B_ENUDrgFV6_1;
	wire w_dff_B_QiucTPP74_1;
	wire w_dff_B_0bzNuzCC6_1;
	wire w_dff_B_WKWUERgi6_1;
	wire w_dff_B_CE07WeNE8_1;
	wire w_dff_B_6Gxr33yF0_1;
	wire w_dff_B_smrgTVRZ0_1;
	wire w_dff_B_HKmPsPlD7_1;
	wire w_dff_B_w4gle9Fi8_1;
	wire w_dff_B_0l6Fwr7h9_1;
	wire w_dff_B_yX8FJu2R6_1;
	wire w_dff_B_rfFExPzG2_1;
	wire w_dff_B_mVKGQXKT0_1;
	wire w_dff_B_wRfypqQU9_1;
	wire w_dff_B_FFaY4lUK9_1;
	wire w_dff_B_iTYtuHjh7_1;
	wire w_dff_B_A6BE0GtO2_1;
	wire w_dff_B_cJyNYkpL9_1;
	wire w_dff_B_vTdJpKuB7_1;
	wire w_dff_B_SBVp6tmq7_1;
	wire w_dff_B_XIgoaezm7_1;
	wire w_dff_B_fgqZTn0Y2_1;
	wire w_dff_B_dBGCToTY4_1;
	wire w_dff_B_f1na4EFN5_1;
	wire w_dff_B_5RN1rz7j2_1;
	wire w_dff_B_KL748LSw3_1;
	wire w_dff_B_LVEgZ2y84_1;
	wire w_dff_B_Pz0C8YGX5_1;
	wire w_dff_B_fIIhbOo01_1;
	wire w_dff_B_AgVwI4mG7_1;
	wire w_dff_B_gb5X35pF6_1;
	wire w_dff_B_lTF4DvuM2_1;
	wire w_dff_B_fpQBtV6F4_1;
	wire w_dff_B_cXx7hrRE8_1;
	wire w_dff_B_yU8IOQd13_1;
	wire w_dff_B_EBuIYaZv1_1;
	wire w_dff_B_NhG75iV78_1;
	wire w_dff_B_P1xugy5g5_1;
	wire w_dff_B_qJKTQRMG5_1;
	wire w_dff_B_HSAtnPCm9_1;
	wire w_dff_B_2OI6n3n12_1;
	wire w_dff_B_HNtekZpL1_1;
	wire w_dff_B_reYtGFKb0_1;
	wire w_dff_B_RlHvAOD07_1;
	wire w_dff_B_sPPHuCiZ6_1;
	wire w_dff_B_FazavZOt9_1;
	wire w_dff_B_JtloA87w9_1;
	wire w_dff_B_XMzLTVwp1_1;
	wire w_dff_B_e0QxKCJC7_1;
	wire w_dff_B_fYxI2bvJ1_1;
	wire w_dff_B_29qVH3sF3_1;
	wire w_dff_B_yDHr625w2_1;
	wire w_dff_B_2nt6yQUH0_1;
	wire w_dff_B_BMA8R8kp0_1;
	wire w_dff_B_CWvGASmY1_1;
	wire w_dff_B_zXeAHdLL5_1;
	wire w_dff_B_iCcYTe8i1_1;
	wire w_dff_B_KKQakevS5_0;
	wire w_dff_B_IhDGF9wD5_0;
	wire w_dff_B_4RNSSUwD7_0;
	wire w_dff_B_pJYJVPvG1_0;
	wire w_dff_B_MeZqI1Vs8_0;
	wire w_dff_B_NUmgf4hR3_0;
	wire w_dff_B_NaEsykuF6_0;
	wire w_dff_B_djV25LEY0_0;
	wire w_dff_B_5Ye4GQGV8_0;
	wire w_dff_B_S1Ux8Jpl1_0;
	wire w_dff_B_BuJDb4Zd8_0;
	wire w_dff_B_vyYoU76S7_0;
	wire w_dff_B_j4eDO0iq0_0;
	wire w_dff_B_vzYntVQH4_0;
	wire w_dff_B_DhLw4Sf48_0;
	wire w_dff_B_kRnq9FQR5_0;
	wire w_dff_B_Clh0ZgdA4_0;
	wire w_dff_B_s7LPLWVc3_0;
	wire w_dff_B_HUEhu5CO6_0;
	wire w_dff_B_4ABZhlbX6_0;
	wire w_dff_B_t4q3b0OU9_0;
	wire w_dff_B_l9eIGpDQ4_0;
	wire w_dff_B_I20CSoCB9_0;
	wire w_dff_B_w5YhRXmd8_0;
	wire w_dff_B_en541yeg8_0;
	wire w_dff_B_wdo74DPK9_0;
	wire w_dff_B_KQ7vyMZB6_0;
	wire w_dff_B_QqJtAtlP6_0;
	wire w_dff_B_HpDSNcJq8_0;
	wire w_dff_B_nhUFAeSf1_0;
	wire w_dff_B_Lrerls4A4_0;
	wire w_dff_B_yL4zEJyM6_0;
	wire w_dff_B_YUfHx6So4_0;
	wire w_dff_B_co16vS2v1_0;
	wire w_dff_B_eJ5ImPck9_0;
	wire w_dff_B_GvsBcK7a3_0;
	wire w_dff_B_DDvavwnA4_0;
	wire w_dff_B_XG1tvJuA4_0;
	wire w_dff_B_i4gwd2VF1_0;
	wire w_dff_B_OOAWPb6Z3_0;
	wire w_dff_B_Df0fWIFc7_0;
	wire w_dff_B_hHnVT1au1_0;
	wire w_dff_B_gGPz1dSO0_0;
	wire w_dff_B_kQFMvZhe5_0;
	wire w_dff_B_bUueOIPZ0_0;
	wire w_dff_B_PfqZblfI4_0;
	wire w_dff_B_J0s7zKTJ6_0;
	wire w_dff_B_lmfqUDMB1_0;
	wire w_dff_B_LVKqfL9B0_0;
	wire w_dff_B_q7Ocs7Ei2_0;
	wire w_dff_B_kW0hc2Fd0_0;
	wire w_dff_B_kOk8aa1D3_0;
	wire w_dff_B_4Mppnres1_0;
	wire w_dff_B_u23GWRg08_0;
	wire w_dff_B_JQaMCbOl3_0;
	wire w_dff_B_tzwRobKE2_0;
	wire w_dff_B_6GPTC3jI3_0;
	wire w_dff_B_0A23CzIg8_0;
	wire w_dff_B_1gHyfTLa9_0;
	wire w_dff_B_VBw2aKEP2_0;
	wire w_dff_B_DttoBILE6_0;
	wire w_dff_B_Qop7ZEK13_0;
	wire w_dff_B_Sd9TXsMA3_0;
	wire w_dff_B_nXZZwd4K5_0;
	wire w_dff_B_NmUpZhn23_0;
	wire w_dff_B_YO3I10x21_0;
	wire w_dff_B_uLZagXrY4_0;
	wire w_dff_B_0adFijnY2_0;
	wire w_dff_B_OPUjSWhz6_0;
	wire w_dff_B_vBjknD2k1_0;
	wire w_dff_B_Ze6FlNRD1_0;
	wire w_dff_B_ZGHgKduP7_0;
	wire w_dff_B_6xRazE0Z0_0;
	wire w_dff_B_1LX0OJy92_0;
	wire w_dff_B_eQj5PWyb8_0;
	wire w_dff_B_fzcQWGjQ1_1;
	wire w_dff_B_iWqqy8Ef0_1;
	wire w_dff_B_9Av6yP9T3_1;
	wire w_dff_B_YXx2SfdY1_1;
	wire w_dff_B_oIYmjxts5_1;
	wire w_dff_B_p8yNM6qJ2_1;
	wire w_dff_B_FCCUOyOc5_1;
	wire w_dff_B_QT1NzXQi2_1;
	wire w_dff_B_U8HTmwp55_1;
	wire w_dff_B_FUmWtdDH4_1;
	wire w_dff_B_MEOVQKAS1_1;
	wire w_dff_B_UdPpq5NB9_1;
	wire w_dff_B_Mhc9hgNk9_1;
	wire w_dff_B_Qapas9H97_1;
	wire w_dff_B_eLBOgaF59_1;
	wire w_dff_B_MoASXsnZ0_1;
	wire w_dff_B_5jhs2Gql9_1;
	wire w_dff_B_rHroq8Um7_1;
	wire w_dff_B_hM0BHclV2_1;
	wire w_dff_B_XIoaE5mR7_1;
	wire w_dff_B_5orr76Oy5_1;
	wire w_dff_B_MBvwhF022_1;
	wire w_dff_B_1ZAhBf8L2_1;
	wire w_dff_B_on9oBKIb0_1;
	wire w_dff_B_nuwwpKgZ5_1;
	wire w_dff_B_Ce1x3yho2_1;
	wire w_dff_B_DhjtPnGr8_1;
	wire w_dff_B_2oCfYTSA5_1;
	wire w_dff_B_Xm2qg5Nn8_1;
	wire w_dff_B_CAmA70hQ5_1;
	wire w_dff_B_Ql0RvhiW8_1;
	wire w_dff_B_UD7L9CII8_1;
	wire w_dff_B_CpsaaURa7_1;
	wire w_dff_B_VSOnUax70_1;
	wire w_dff_B_bTZjxV3X9_1;
	wire w_dff_B_m9XojbnU1_1;
	wire w_dff_B_ec05QcVN4_1;
	wire w_dff_B_UWWylQYY9_1;
	wire w_dff_B_UBv1pgTI6_1;
	wire w_dff_B_93kHH1z81_1;
	wire w_dff_B_vh4YDzLy3_1;
	wire w_dff_B_ngm6uAAi4_1;
	wire w_dff_B_0H8Cm9Ip6_1;
	wire w_dff_B_li0ODhpa9_1;
	wire w_dff_B_ICpyKWgS1_1;
	wire w_dff_B_POTFi3md5_1;
	wire w_dff_B_pXRCJx5B8_1;
	wire w_dff_B_g56UXDze6_1;
	wire w_dff_B_0Gx8e77j0_1;
	wire w_dff_B_JWiXsLj33_1;
	wire w_dff_B_HdJm9LvW7_1;
	wire w_dff_B_WiI54ckC1_1;
	wire w_dff_B_WTtqsecn6_1;
	wire w_dff_B_idsXCX3d9_1;
	wire w_dff_B_y2F4RiEV4_1;
	wire w_dff_B_11Vt3sBK0_1;
	wire w_dff_B_wM9oTRtT9_1;
	wire w_dff_B_aaiF4Yzg2_1;
	wire w_dff_B_WJdfKBfg4_1;
	wire w_dff_B_cwwrwLCm6_1;
	wire w_dff_B_Y6qNhR5p3_1;
	wire w_dff_B_sUdhBr9E5_1;
	wire w_dff_B_cA5cZ6907_1;
	wire w_dff_B_b9BLn1h61_1;
	wire w_dff_B_hnEdSN8A2_1;
	wire w_dff_B_W7FVO3aG1_1;
	wire w_dff_B_9cvDDs469_1;
	wire w_dff_B_2K7tkW5v1_1;
	wire w_dff_B_pbgoh5Qd8_1;
	wire w_dff_B_rBwhVI587_1;
	wire w_dff_B_cVeA81v10_1;
	wire w_dff_B_c4AgP0Gh0_1;
	wire w_dff_B_h5ChKpm86_1;
	wire w_dff_B_yknhl01q3_1;
	wire w_dff_B_NXdUOz5k1_0;
	wire w_dff_B_rvLNVcuE6_0;
	wire w_dff_B_gHuqydpu1_0;
	wire w_dff_B_Womz66i84_0;
	wire w_dff_B_AyNzqpIh4_0;
	wire w_dff_B_AXGHcgiM1_0;
	wire w_dff_B_OLgFLNcu7_0;
	wire w_dff_B_fGmBEd840_0;
	wire w_dff_B_LAE4i4Nd7_0;
	wire w_dff_B_5nYvM20E9_0;
	wire w_dff_B_FLISnqZ31_0;
	wire w_dff_B_kgskhX5U8_0;
	wire w_dff_B_pseM8KBi5_0;
	wire w_dff_B_NCZ3iCjn1_0;
	wire w_dff_B_yfd8K9kw0_0;
	wire w_dff_B_soHwuBmQ0_0;
	wire w_dff_B_ttlUcDMf3_0;
	wire w_dff_B_wDJ7CNjL7_0;
	wire w_dff_B_DBH5LdSb4_0;
	wire w_dff_B_aSbcZRhu5_0;
	wire w_dff_B_BU8ADFap7_0;
	wire w_dff_B_2QBwY8623_0;
	wire w_dff_B_NMCoNdre5_0;
	wire w_dff_B_4JlLuIGm7_0;
	wire w_dff_B_7k2r6Ht79_0;
	wire w_dff_B_kuLBzDew0_0;
	wire w_dff_B_VbRP7utx1_0;
	wire w_dff_B_BgjkTimB9_0;
	wire w_dff_B_pOWyAVL76_0;
	wire w_dff_B_txbNW4CK3_0;
	wire w_dff_B_8YcG4hoe3_0;
	wire w_dff_B_VHsc707M3_0;
	wire w_dff_B_FoqpMuCn2_0;
	wire w_dff_B_MOUfJ2bf1_0;
	wire w_dff_B_zKYMz6YK5_0;
	wire w_dff_B_W1CSDG8t9_0;
	wire w_dff_B_lkMNodfX8_0;
	wire w_dff_B_DeuUb19m8_0;
	wire w_dff_B_2T2l4kmR7_0;
	wire w_dff_B_vildeu6e0_0;
	wire w_dff_B_CG00E0vw7_0;
	wire w_dff_B_ApCQjulg9_0;
	wire w_dff_B_74o4HdjE8_0;
	wire w_dff_B_zDCkAEWQ3_0;
	wire w_dff_B_fK4nLh8r9_0;
	wire w_dff_B_3fBo5HpL0_0;
	wire w_dff_B_FKZmoGFT1_0;
	wire w_dff_B_UShcwkED6_0;
	wire w_dff_B_4PUDOwNs3_0;
	wire w_dff_B_9Fa55XcT1_0;
	wire w_dff_B_sLTfuto52_0;
	wire w_dff_B_etjT0UeA0_0;
	wire w_dff_B_nr2Yngns4_0;
	wire w_dff_B_ttamoL4V1_0;
	wire w_dff_B_40zbkknR9_0;
	wire w_dff_B_0WwOXIgK8_0;
	wire w_dff_B_VKAWpe2X1_0;
	wire w_dff_B_uSx5Ur0E4_0;
	wire w_dff_B_JDqwaRfV9_0;
	wire w_dff_B_mo9r74Aw1_0;
	wire w_dff_B_J9W8VrJi2_0;
	wire w_dff_B_w1JhITiY6_0;
	wire w_dff_B_3YhGHSeV9_0;
	wire w_dff_B_T9IyBr3I4_0;
	wire w_dff_B_DRhjfae82_0;
	wire w_dff_B_G75xdA971_0;
	wire w_dff_B_ZcdO2RPK4_0;
	wire w_dff_B_E2sDRwcC4_0;
	wire w_dff_B_vnDJJop06_0;
	wire w_dff_B_6K4WLKcr8_0;
	wire w_dff_B_3n7DBwv68_0;
	wire w_dff_B_7Ak4wJe99_0;
	wire w_dff_B_PLV9oANz4_0;
	wire w_dff_B_zTdSogfq8_0;
	wire w_dff_B_P1a241067_1;
	wire w_dff_B_WBtJ2fqY2_1;
	wire w_dff_B_9jD9mowu5_1;
	wire w_dff_B_0fmoSMOy1_1;
	wire w_dff_B_VTyKecC02_1;
	wire w_dff_B_4C4bnUWE3_1;
	wire w_dff_B_SKBPGTCL9_1;
	wire w_dff_B_OvVv21AE5_1;
	wire w_dff_B_k11z6bDt0_1;
	wire w_dff_B_OQ1vd6TP3_1;
	wire w_dff_B_9Uxuewrh6_1;
	wire w_dff_B_UQpsdQPT1_1;
	wire w_dff_B_3NH9F9hi3_1;
	wire w_dff_B_XDXpJEb01_1;
	wire w_dff_B_G1DgOKdE8_1;
	wire w_dff_B_pwewoXo13_1;
	wire w_dff_B_pAjrQGmh3_1;
	wire w_dff_B_Aw8S6JcH2_1;
	wire w_dff_B_CKKMrjSH4_1;
	wire w_dff_B_OiZm2VEm8_1;
	wire w_dff_B_A3iCMKUs1_1;
	wire w_dff_B_10It760G9_1;
	wire w_dff_B_DX4UyAc42_1;
	wire w_dff_B_lU8vVODj6_1;
	wire w_dff_B_H2pjsWzT9_1;
	wire w_dff_B_AcJPtQK80_1;
	wire w_dff_B_bNtDkg091_1;
	wire w_dff_B_YpFb5RHt5_1;
	wire w_dff_B_MwbFFXpn5_1;
	wire w_dff_B_MGixn9EF7_1;
	wire w_dff_B_CrK3a6ka5_1;
	wire w_dff_B_fADA8nPu2_1;
	wire w_dff_B_iDDLOMSv5_1;
	wire w_dff_B_bupoSeDY8_1;
	wire w_dff_B_E9pOElhA6_1;
	wire w_dff_B_VPlwSNKi2_1;
	wire w_dff_B_9UZzjdqH8_1;
	wire w_dff_B_N1eUPrLV7_1;
	wire w_dff_B_fXdK2AGn0_1;
	wire w_dff_B_mErZx3rd6_1;
	wire w_dff_B_pe0G3Tzl6_1;
	wire w_dff_B_80W7Q4dK1_1;
	wire w_dff_B_kE4D6ikc6_1;
	wire w_dff_B_NZR66vAv1_1;
	wire w_dff_B_i7grhFx50_1;
	wire w_dff_B_41zHWW3w6_1;
	wire w_dff_B_7bi29k8c5_1;
	wire w_dff_B_LpPMhu5y7_1;
	wire w_dff_B_0zcTE1Bs3_1;
	wire w_dff_B_0qLLWQmH0_1;
	wire w_dff_B_kSOBHOgB4_1;
	wire w_dff_B_GejgVfJ74_1;
	wire w_dff_B_Jl2NPXL00_1;
	wire w_dff_B_2lcY77pa2_1;
	wire w_dff_B_8L5gM2XY0_1;
	wire w_dff_B_3ktVkiK66_1;
	wire w_dff_B_a3npL29q4_1;
	wire w_dff_B_IWrQNUuz6_1;
	wire w_dff_B_aZkSvajn3_1;
	wire w_dff_B_l8u35DY66_1;
	wire w_dff_B_8igXaLMG6_1;
	wire w_dff_B_JrGG7lIa6_1;
	wire w_dff_B_JnJbw1BE6_1;
	wire w_dff_B_ZOZbBxey3_1;
	wire w_dff_B_jXTzPP9m4_1;
	wire w_dff_B_NoabEJFQ3_1;
	wire w_dff_B_LoQRTAu85_1;
	wire w_dff_B_btPsXjUD0_1;
	wire w_dff_B_NQmElksK9_1;
	wire w_dff_B_Gv8tLM9X0_1;
	wire w_dff_B_3omyXlQ26_1;
	wire w_dff_B_LnUCF9vy8_1;
	wire w_dff_B_yBmv7bjw0_1;
	wire w_dff_B_RAHituV56_0;
	wire w_dff_B_aA9MMUZg1_0;
	wire w_dff_B_MiQYWdBZ7_0;
	wire w_dff_B_ZEsAe6eD3_0;
	wire w_dff_B_i6VhmQwu4_0;
	wire w_dff_B_L3ynKQpL0_0;
	wire w_dff_B_S3mZmyAG0_0;
	wire w_dff_B_ZYTmjL1Y3_0;
	wire w_dff_B_VOoMSUSD9_0;
	wire w_dff_B_zFqCZzvi4_0;
	wire w_dff_B_uSlPX1qB3_0;
	wire w_dff_B_VlSZki5Q5_0;
	wire w_dff_B_6IxXXMo99_0;
	wire w_dff_B_tS0SPITA0_0;
	wire w_dff_B_dLKL2beP3_0;
	wire w_dff_B_0GqKqaxd3_0;
	wire w_dff_B_x9E4GK9J7_0;
	wire w_dff_B_H8rbAbgZ0_0;
	wire w_dff_B_eAxQyGb48_0;
	wire w_dff_B_DOSvCxMA8_0;
	wire w_dff_B_nZ7TMs2t3_0;
	wire w_dff_B_Q4jb6NL63_0;
	wire w_dff_B_Rrqr1Uj90_0;
	wire w_dff_B_mfjnUpzA1_0;
	wire w_dff_B_jRAkfUvh2_0;
	wire w_dff_B_OZJFt1Jz9_0;
	wire w_dff_B_oYk5U38s2_0;
	wire w_dff_B_HWRZgDLW4_0;
	wire w_dff_B_MlqYv43V0_0;
	wire w_dff_B_5ej493qt9_0;
	wire w_dff_B_NqJiMSj51_0;
	wire w_dff_B_87PaAeXd0_0;
	wire w_dff_B_pruRAMB99_0;
	wire w_dff_B_1MNEhZdI5_0;
	wire w_dff_B_IpnBBlcW6_0;
	wire w_dff_B_hiA6z7NU1_0;
	wire w_dff_B_QzJp9Tl70_0;
	wire w_dff_B_7O96u6dz3_0;
	wire w_dff_B_6dwmHMj61_0;
	wire w_dff_B_lsEPhBgi2_0;
	wire w_dff_B_0qBd94Ap8_0;
	wire w_dff_B_fEVehGMh4_0;
	wire w_dff_B_DSndmckA4_0;
	wire w_dff_B_2ogHnr3U7_0;
	wire w_dff_B_qrPuhFOX2_0;
	wire w_dff_B_su8gd8sq2_0;
	wire w_dff_B_KbhraIE22_0;
	wire w_dff_B_iKk4QUEi2_0;
	wire w_dff_B_zyjU2V6i8_0;
	wire w_dff_B_dlmvgXlg2_0;
	wire w_dff_B_VNb5ncHS1_0;
	wire w_dff_B_KfjkTy7X0_0;
	wire w_dff_B_Bb9Mwo246_0;
	wire w_dff_B_YnB2EQJc4_0;
	wire w_dff_B_qpnWWWUU5_0;
	wire w_dff_B_FgWrSpTH5_0;
	wire w_dff_B_BYDiHvZm4_0;
	wire w_dff_B_Do5MkOoQ6_0;
	wire w_dff_B_yrz9v0t61_0;
	wire w_dff_B_5z3U7XQD0_0;
	wire w_dff_B_3XnMhdo41_0;
	wire w_dff_B_eBPAsBAR6_0;
	wire w_dff_B_IZUlk9BH6_0;
	wire w_dff_B_dxMJb1gP3_0;
	wire w_dff_B_vPvwatj83_0;
	wire w_dff_B_wRo5T9ko6_0;
	wire w_dff_B_Zc2pNYTa5_0;
	wire w_dff_B_lpghyYVv7_0;
	wire w_dff_B_2Hi23M2r2_0;
	wire w_dff_B_PZz4M9hI3_0;
	wire w_dff_B_Y9Cdh24Z6_0;
	wire w_dff_B_BODBuvVB6_0;
	wire w_dff_B_rKut0M2W1_0;
	wire w_dff_B_b4HSidhS9_1;
	wire w_dff_B_GrqHro6J9_1;
	wire w_dff_B_QwqtT17P6_1;
	wire w_dff_B_SvqzD8iR4_1;
	wire w_dff_B_5N730P6n1_1;
	wire w_dff_B_PN4JjQXV6_1;
	wire w_dff_B_xvcyzseX9_1;
	wire w_dff_B_SmHblLy75_1;
	wire w_dff_B_T5smbZTS3_1;
	wire w_dff_B_GACa4STw2_1;
	wire w_dff_B_M4lhjITy5_1;
	wire w_dff_B_PRzfMe5g1_1;
	wire w_dff_B_5OcTVZmz6_1;
	wire w_dff_B_1g5NA4Bn0_1;
	wire w_dff_B_AtgLpfYf0_1;
	wire w_dff_B_pl2Jfj7l2_1;
	wire w_dff_B_l2TMvDHP2_1;
	wire w_dff_B_6MYnmPOk8_1;
	wire w_dff_B_7up5ZRKX0_1;
	wire w_dff_B_WkErKG0L6_1;
	wire w_dff_B_mun8BVp62_1;
	wire w_dff_B_epqHRWpi1_1;
	wire w_dff_B_Oy2Vne6r4_1;
	wire w_dff_B_2Y9W4CfV7_1;
	wire w_dff_B_NNLff3Lt3_1;
	wire w_dff_B_K686eWDB7_1;
	wire w_dff_B_r7aCH8wM3_1;
	wire w_dff_B_zSS8ZzN40_1;
	wire w_dff_B_9LHZBG0E0_1;
	wire w_dff_B_xk1N7SbQ3_1;
	wire w_dff_B_tcFwzUeZ0_1;
	wire w_dff_B_cJsWbnMT9_1;
	wire w_dff_B_cpxgLhzs4_1;
	wire w_dff_B_PNSolVS35_1;
	wire w_dff_B_KTV7JitT7_1;
	wire w_dff_B_S5kF8oyp1_1;
	wire w_dff_B_4eOrq1hD2_1;
	wire w_dff_B_jYEZptSz4_1;
	wire w_dff_B_84AFV4wZ4_1;
	wire w_dff_B_SbOqHVtP9_1;
	wire w_dff_B_PihnK1wM7_1;
	wire w_dff_B_pC7Qi3dg8_1;
	wire w_dff_B_kFReKYZS6_1;
	wire w_dff_B_HgL6vTZ53_1;
	wire w_dff_B_M6R53h0c2_1;
	wire w_dff_B_jVlFUBsW6_1;
	wire w_dff_B_o9X0LLj41_1;
	wire w_dff_B_ydGaxygF9_1;
	wire w_dff_B_pvG1Bkes5_1;
	wire w_dff_B_zJdmmRxx5_1;
	wire w_dff_B_hZMGqjXs4_1;
	wire w_dff_B_pM2AWCf15_1;
	wire w_dff_B_BWm5S38Q9_1;
	wire w_dff_B_pJmzltft3_1;
	wire w_dff_B_aH3rfv8h8_1;
	wire w_dff_B_TK7dTSFu2_1;
	wire w_dff_B_apqCesxp5_1;
	wire w_dff_B_fTtlmO4F2_1;
	wire w_dff_B_9JdUVkl86_1;
	wire w_dff_B_gfWeo0Ef7_1;
	wire w_dff_B_B2rUbfEZ7_1;
	wire w_dff_B_A6hKXfm65_1;
	wire w_dff_B_rgd4q4JO6_1;
	wire w_dff_B_qTTQQUpr0_1;
	wire w_dff_B_ATxwmUt31_1;
	wire w_dff_B_HaKLKpFt1_1;
	wire w_dff_B_GYiACixA2_1;
	wire w_dff_B_O8vQytY30_1;
	wire w_dff_B_qARWhyZh9_1;
	wire w_dff_B_XT4w1tQi0_1;
	wire w_dff_B_nAL383XY7_1;
	wire w_dff_B_CmLHlizM1_1;
	wire w_dff_B_GFyTLlSL7_0;
	wire w_dff_B_PxTmtekB1_0;
	wire w_dff_B_QHM1ATau8_0;
	wire w_dff_B_dRDueS452_0;
	wire w_dff_B_AH6aannt7_0;
	wire w_dff_B_3rV3KiuU9_0;
	wire w_dff_B_9YAuWKnM3_0;
	wire w_dff_B_ssRh6omy8_0;
	wire w_dff_B_B8JeIfJd8_0;
	wire w_dff_B_cjHgWY2H3_0;
	wire w_dff_B_ywvVU7Mf4_0;
	wire w_dff_B_BwVmR7SR8_0;
	wire w_dff_B_nfUXkAuU9_0;
	wire w_dff_B_NQ3hdSku8_0;
	wire w_dff_B_DBcCHZp04_0;
	wire w_dff_B_n4cvWEd38_0;
	wire w_dff_B_b02EVVu31_0;
	wire w_dff_B_tmeqqpIg0_0;
	wire w_dff_B_aaBQF0Cn8_0;
	wire w_dff_B_Fk1cmqpc9_0;
	wire w_dff_B_jAcp4NRB0_0;
	wire w_dff_B_z424nFrH6_0;
	wire w_dff_B_5gWowZOH2_0;
	wire w_dff_B_5n6abP317_0;
	wire w_dff_B_4AL1rcrm0_0;
	wire w_dff_B_NxJ7c8hl3_0;
	wire w_dff_B_YUV4qxrB6_0;
	wire w_dff_B_WBcw1FaZ6_0;
	wire w_dff_B_Y40OrlF30_0;
	wire w_dff_B_n08nwpdU0_0;
	wire w_dff_B_zVLiVMKA8_0;
	wire w_dff_B_ddsPfdrH4_0;
	wire w_dff_B_nK1cSWgf8_0;
	wire w_dff_B_zhO5B4ZN8_0;
	wire w_dff_B_GLenQ7nM6_0;
	wire w_dff_B_rURqX3Tj8_0;
	wire w_dff_B_DvVKpehl2_0;
	wire w_dff_B_WVedm75X3_0;
	wire w_dff_B_zkc0RCJ48_0;
	wire w_dff_B_etj6C3jq1_0;
	wire w_dff_B_pow9Xqhp8_0;
	wire w_dff_B_IM238BUL5_0;
	wire w_dff_B_BvDFv2aE3_0;
	wire w_dff_B_goKe2PLj9_0;
	wire w_dff_B_GtVZ4Owg1_0;
	wire w_dff_B_bB84obzN0_0;
	wire w_dff_B_TVpGm1bL0_0;
	wire w_dff_B_iGMFxjY16_0;
	wire w_dff_B_HftuvI6x5_0;
	wire w_dff_B_6KgP9fnU4_0;
	wire w_dff_B_n1c7whd10_0;
	wire w_dff_B_utgJJrcv4_0;
	wire w_dff_B_pSIxGsn99_0;
	wire w_dff_B_ZbWtIy7L5_0;
	wire w_dff_B_Z3Qc2kDf4_0;
	wire w_dff_B_L1VMpWZE9_0;
	wire w_dff_B_sTh5CHzI9_0;
	wire w_dff_B_cf2HexZ64_0;
	wire w_dff_B_qgPPnmKV3_0;
	wire w_dff_B_JKcuVPDt2_0;
	wire w_dff_B_k51KdTd10_0;
	wire w_dff_B_mdfpRZoz6_0;
	wire w_dff_B_hwjwXKxG5_0;
	wire w_dff_B_duZOeWpI5_0;
	wire w_dff_B_HAoUd2zw6_0;
	wire w_dff_B_chVpCn8l2_0;
	wire w_dff_B_KZNYSLRT7_0;
	wire w_dff_B_vLichBWZ1_0;
	wire w_dff_B_xgV7aKI32_0;
	wire w_dff_B_ukBXUbxV1_0;
	wire w_dff_B_XnXEUs236_0;
	wire w_dff_B_FLEVHsvk5_0;
	wire w_dff_B_Fn07mpj66_1;
	wire w_dff_B_CPMG4O5U9_1;
	wire w_dff_B_SZoP2WA16_1;
	wire w_dff_B_21kpJTjy4_1;
	wire w_dff_B_sREIaAun7_1;
	wire w_dff_B_rHsmr3kF0_1;
	wire w_dff_B_iJqtsLo26_1;
	wire w_dff_B_ofuibS3N9_1;
	wire w_dff_B_dWbTqyrF3_1;
	wire w_dff_B_5ycJ3PHi8_1;
	wire w_dff_B_23mOysOv2_1;
	wire w_dff_B_wt0vfdau2_1;
	wire w_dff_B_5Gfz4Cbu7_1;
	wire w_dff_B_0z0OIQZK0_1;
	wire w_dff_B_Qucn0uoQ0_1;
	wire w_dff_B_u2B7voVP8_1;
	wire w_dff_B_OsrTxzBq6_1;
	wire w_dff_B_D08ZMa047_1;
	wire w_dff_B_evWj6xiq4_1;
	wire w_dff_B_J40iZ6Ho9_1;
	wire w_dff_B_nWKsqVu08_1;
	wire w_dff_B_viNll7tx8_1;
	wire w_dff_B_qGJVV4M45_1;
	wire w_dff_B_HkIhst496_1;
	wire w_dff_B_VZq9cFdL7_1;
	wire w_dff_B_ounaAOLQ4_1;
	wire w_dff_B_2duDj88d2_1;
	wire w_dff_B_XGy4m2J89_1;
	wire w_dff_B_s29Eg6PN9_1;
	wire w_dff_B_NmxiH5lS5_1;
	wire w_dff_B_nBGMMrt79_1;
	wire w_dff_B_NjWXLlhu1_1;
	wire w_dff_B_QJaX1yLt5_1;
	wire w_dff_B_1nZXS5tk2_1;
	wire w_dff_B_HgjxWLeM9_1;
	wire w_dff_B_QzBSIu435_1;
	wire w_dff_B_NBZzaYUS9_1;
	wire w_dff_B_GqbdVfgC8_1;
	wire w_dff_B_erHLbXQL4_1;
	wire w_dff_B_eUUKJn3q6_1;
	wire w_dff_B_H1ytEKT36_1;
	wire w_dff_B_GGB3ALZY0_1;
	wire w_dff_B_JAfcG5719_1;
	wire w_dff_B_Mxvq50P53_1;
	wire w_dff_B_lVh7q02f0_1;
	wire w_dff_B_yJxWgjrK7_1;
	wire w_dff_B_7bj5zypn6_1;
	wire w_dff_B_bWnn7mRa7_1;
	wire w_dff_B_YFgZ2xtI1_1;
	wire w_dff_B_2q3ifhJd6_1;
	wire w_dff_B_br2dRU665_1;
	wire w_dff_B_jcF9v2hz5_1;
	wire w_dff_B_mNc6PFXQ0_1;
	wire w_dff_B_nFYobDWW9_1;
	wire w_dff_B_AmehRiI93_1;
	wire w_dff_B_YCHQ6EdZ0_1;
	wire w_dff_B_n1SoDHzL9_1;
	wire w_dff_B_DLIX49hN9_1;
	wire w_dff_B_k8xOooFM4_1;
	wire w_dff_B_XwnUYPgR2_1;
	wire w_dff_B_3UQkUfI68_1;
	wire w_dff_B_POirTfb49_1;
	wire w_dff_B_Jm5xqbpj7_1;
	wire w_dff_B_sgnaPnVx9_1;
	wire w_dff_B_zxY0mHzY3_1;
	wire w_dff_B_iWu0Xn025_1;
	wire w_dff_B_VGUWiZmZ8_1;
	wire w_dff_B_w3E6nsfT5_1;
	wire w_dff_B_5nh3WXtJ0_1;
	wire w_dff_B_VkNunJB06_1;
	wire w_dff_B_2xeLz8H77_1;
	wire w_dff_B_nvl1DsuF6_0;
	wire w_dff_B_UxUSEnrq9_0;
	wire w_dff_B_qk7OKlME8_0;
	wire w_dff_B_ljzoi7Gx0_0;
	wire w_dff_B_GyxbHnTi1_0;
	wire w_dff_B_RF2xT56F1_0;
	wire w_dff_B_qtiZPLq51_0;
	wire w_dff_B_poDzi82x6_0;
	wire w_dff_B_F7jtAGL09_0;
	wire w_dff_B_u5nVXoww7_0;
	wire w_dff_B_TT9lRUQV8_0;
	wire w_dff_B_xUbNhu9M1_0;
	wire w_dff_B_TjgeKRwY9_0;
	wire w_dff_B_k8kRByqR6_0;
	wire w_dff_B_tnZDjq6y5_0;
	wire w_dff_B_rCJs1lad9_0;
	wire w_dff_B_PoxsRFmk6_0;
	wire w_dff_B_dd5hwphR4_0;
	wire w_dff_B_CNylEeYP7_0;
	wire w_dff_B_At2ilMbM0_0;
	wire w_dff_B_Jd4F5Olk6_0;
	wire w_dff_B_4QhqIe667_0;
	wire w_dff_B_i9pUHtxJ6_0;
	wire w_dff_B_uRen2yrE3_0;
	wire w_dff_B_vafBg3Vk3_0;
	wire w_dff_B_xuIisjlp4_0;
	wire w_dff_B_eWLD32ma0_0;
	wire w_dff_B_SNQz7Q316_0;
	wire w_dff_B_GsUAQ68U8_0;
	wire w_dff_B_RSaTXRfz7_0;
	wire w_dff_B_USp6mICs2_0;
	wire w_dff_B_4ExvazqS9_0;
	wire w_dff_B_Jd1gpXR12_0;
	wire w_dff_B_5M7EyEsQ4_0;
	wire w_dff_B_IcM4Ep1U6_0;
	wire w_dff_B_I4kbpMhW8_0;
	wire w_dff_B_S3z89LHJ1_0;
	wire w_dff_B_XLnaXlOQ9_0;
	wire w_dff_B_h5fbgJQb2_0;
	wire w_dff_B_4HukJdoK4_0;
	wire w_dff_B_5IG5ManI3_0;
	wire w_dff_B_rkLa2H1l3_0;
	wire w_dff_B_ZEcAbrYv0_0;
	wire w_dff_B_2E1Auvo42_0;
	wire w_dff_B_3isJtvCp9_0;
	wire w_dff_B_rW8HDDwB0_0;
	wire w_dff_B_rM39nGdq6_0;
	wire w_dff_B_0wB66zH80_0;
	wire w_dff_B_oFUvSo5u3_0;
	wire w_dff_B_NOZCM0cf2_0;
	wire w_dff_B_x0K9wlQz2_0;
	wire w_dff_B_NhC7MEUy1_0;
	wire w_dff_B_vRFCuuG98_0;
	wire w_dff_B_UzQOeXxz6_0;
	wire w_dff_B_uuGrenYI4_0;
	wire w_dff_B_HfD8uDU70_0;
	wire w_dff_B_hfjeN3Wx6_0;
	wire w_dff_B_ECUwhUDy0_0;
	wire w_dff_B_fU2RXRtI8_0;
	wire w_dff_B_CbEXAH8a8_0;
	wire w_dff_B_iR9EAUy26_0;
	wire w_dff_B_Le0kiDce0_0;
	wire w_dff_B_7QGzODXK6_0;
	wire w_dff_B_fRDxdxij7_0;
	wire w_dff_B_c4Pa7EKc0_0;
	wire w_dff_B_nQwA0zln9_0;
	wire w_dff_B_LmJdCNY68_0;
	wire w_dff_B_hgg32NFA5_0;
	wire w_dff_B_m9LK9m683_0;
	wire w_dff_B_FuCsEnzB2_0;
	wire w_dff_B_opoKmvzR0_0;
	wire w_dff_B_fPtnV4ne1_1;
	wire w_dff_B_u5KB2iBC0_1;
	wire w_dff_B_jdWkOwwN7_1;
	wire w_dff_B_uwYk1ykc6_1;
	wire w_dff_B_SiluVxBi9_1;
	wire w_dff_B_VAACcGSx5_1;
	wire w_dff_B_h3w4uTr13_1;
	wire w_dff_B_39zBnsb43_1;
	wire w_dff_B_aZtWOlo36_1;
	wire w_dff_B_A1Dsif1O2_1;
	wire w_dff_B_UNfAREHO0_1;
	wire w_dff_B_Sgz1soDP7_1;
	wire w_dff_B_2JK0dxAD0_1;
	wire w_dff_B_iFw6OVHl8_1;
	wire w_dff_B_RjclR5278_1;
	wire w_dff_B_6uAudWPB3_1;
	wire w_dff_B_plIOSQUf0_1;
	wire w_dff_B_jKEPCnNX6_1;
	wire w_dff_B_YVaQyCet2_1;
	wire w_dff_B_iz4QeOnO6_1;
	wire w_dff_B_rFPliHwR7_1;
	wire w_dff_B_awJCPDGO5_1;
	wire w_dff_B_2C25k7Jb7_1;
	wire w_dff_B_rVS7Kz5u7_1;
	wire w_dff_B_trc6snZY1_1;
	wire w_dff_B_eQjwPyqC5_1;
	wire w_dff_B_jP9xQUtG5_1;
	wire w_dff_B_jqdsOLBy4_1;
	wire w_dff_B_9wvJyR1H1_1;
	wire w_dff_B_5tdoIqmD1_1;
	wire w_dff_B_1McRnk3w4_1;
	wire w_dff_B_NuFG2oGH1_1;
	wire w_dff_B_0NdLb2sr3_1;
	wire w_dff_B_EdpR58VJ4_1;
	wire w_dff_B_vCoVINpe7_1;
	wire w_dff_B_q3H8vo2M7_1;
	wire w_dff_B_gU6I6iIH9_1;
	wire w_dff_B_X8rZibmw1_1;
	wire w_dff_B_8BSjqyq00_1;
	wire w_dff_B_MZKGPgIk0_1;
	wire w_dff_B_vfoBeLG48_1;
	wire w_dff_B_pxtXzr5M9_1;
	wire w_dff_B_akxC9Onn9_1;
	wire w_dff_B_kAmT2Wwo3_1;
	wire w_dff_B_x9OiuhUO1_1;
	wire w_dff_B_sDbcG5VX0_1;
	wire w_dff_B_ohXgzFRg6_1;
	wire w_dff_B_tuFLE2z73_1;
	wire w_dff_B_a8Wm1DCm6_1;
	wire w_dff_B_nTMYM4Ce6_1;
	wire w_dff_B_1Zj5aoxT5_1;
	wire w_dff_B_khpJAC276_1;
	wire w_dff_B_5h2KiXqU1_1;
	wire w_dff_B_3OZt11gE3_1;
	wire w_dff_B_Z14jyo114_1;
	wire w_dff_B_vIyHb3Mq2_1;
	wire w_dff_B_aCtDj9Ow4_1;
	wire w_dff_B_mR77MZ8I0_1;
	wire w_dff_B_DBZVxHnp3_1;
	wire w_dff_B_AhsGIHbx2_1;
	wire w_dff_B_yhVf4j9i5_1;
	wire w_dff_B_u2csuEJ05_1;
	wire w_dff_B_qgLzhbVe3_1;
	wire w_dff_B_QWLTNVuz7_1;
	wire w_dff_B_Nn3e0hev5_1;
	wire w_dff_B_aCH4LLod8_1;
	wire w_dff_B_shoRslMY0_1;
	wire w_dff_B_uXXOUjCv2_1;
	wire w_dff_B_9VcyI3r83_1;
	wire w_dff_B_pVF4M0wG0_1;
	wire w_dff_B_5Ni2CrgP5_0;
	wire w_dff_B_FSDDnmCR6_0;
	wire w_dff_B_UM8lSR7m2_0;
	wire w_dff_B_D21i3gug7_0;
	wire w_dff_B_9ObiCvZv1_0;
	wire w_dff_B_Lm0XaGbR3_0;
	wire w_dff_B_2YMpziwZ3_0;
	wire w_dff_B_C44ROdL24_0;
	wire w_dff_B_TabcxDqg2_0;
	wire w_dff_B_h2KZ6CGk5_0;
	wire w_dff_B_sAvbZ5hM3_0;
	wire w_dff_B_quVmLe8D7_0;
	wire w_dff_B_vdaOlCqG6_0;
	wire w_dff_B_yQqVSCO33_0;
	wire w_dff_B_eH7kOKHS9_0;
	wire w_dff_B_FLRfAfIX1_0;
	wire w_dff_B_kGFRuOZH4_0;
	wire w_dff_B_eXcRlOOD7_0;
	wire w_dff_B_TaQKXIL92_0;
	wire w_dff_B_7sHwa8Mc9_0;
	wire w_dff_B_zO5Y0dJj3_0;
	wire w_dff_B_FUHHROpm6_0;
	wire w_dff_B_hg6yJ2KZ4_0;
	wire w_dff_B_3U56scaO3_0;
	wire w_dff_B_0IdauRGb0_0;
	wire w_dff_B_6E5XANT57_0;
	wire w_dff_B_0LwHkpT39_0;
	wire w_dff_B_W5LqX5Ho0_0;
	wire w_dff_B_GB0jboq45_0;
	wire w_dff_B_RfGtvzon1_0;
	wire w_dff_B_vA3eJbty0_0;
	wire w_dff_B_fMkP9Uic2_0;
	wire w_dff_B_hyPuF6Ow8_0;
	wire w_dff_B_RIhNgZz05_0;
	wire w_dff_B_EKHbUWMj5_0;
	wire w_dff_B_geDmSBno5_0;
	wire w_dff_B_OriJUwel6_0;
	wire w_dff_B_xgMQCIlB4_0;
	wire w_dff_B_zsbImneq4_0;
	wire w_dff_B_sk0oR1Kf4_0;
	wire w_dff_B_q3RSenw00_0;
	wire w_dff_B_Tx9pgges0_0;
	wire w_dff_B_1PuhqfBk1_0;
	wire w_dff_B_S3oheR1K1_0;
	wire w_dff_B_lxh7nCk79_0;
	wire w_dff_B_T7cWo3xx4_0;
	wire w_dff_B_7GSxoU2g5_0;
	wire w_dff_B_zHi0uYkY5_0;
	wire w_dff_B_eGWX7n3w8_0;
	wire w_dff_B_h0nfvhi62_0;
	wire w_dff_B_vFEo9h5K5_0;
	wire w_dff_B_0SoYbOul9_0;
	wire w_dff_B_mpidmNvA2_0;
	wire w_dff_B_1MmgSsZ66_0;
	wire w_dff_B_3azS8yEz2_0;
	wire w_dff_B_dYF03m3J8_0;
	wire w_dff_B_7wkog4mP8_0;
	wire w_dff_B_mOWiLkdh4_0;
	wire w_dff_B_6AcOMnso4_0;
	wire w_dff_B_OTTj2QL28_0;
	wire w_dff_B_VYksLNI65_0;
	wire w_dff_B_Z8NxScdf1_0;
	wire w_dff_B_3ldWa6gA5_0;
	wire w_dff_B_C0O7QFSI4_0;
	wire w_dff_B_wSLYOuqJ4_0;
	wire w_dff_B_JrId8InE1_0;
	wire w_dff_B_7K3aF9Vz9_0;
	wire w_dff_B_5f4GkgB66_0;
	wire w_dff_B_1ntz2iTa3_0;
	wire w_dff_B_ok8xe67Q0_0;
	wire w_dff_B_ptW8XoVC7_1;
	wire w_dff_B_3pJQMJoW5_1;
	wire w_dff_B_cekGFxVL7_1;
	wire w_dff_B_ixlxO9H45_1;
	wire w_dff_B_dA0IOJR33_1;
	wire w_dff_B_FlMMIyM59_1;
	wire w_dff_B_Jxka773Z0_1;
	wire w_dff_B_rdR2pFcl4_1;
	wire w_dff_B_DTbs7MKm6_1;
	wire w_dff_B_XPvgE4Qs9_1;
	wire w_dff_B_jz8Re5ZI2_1;
	wire w_dff_B_zJlMaynd1_1;
	wire w_dff_B_KqMN3XV17_1;
	wire w_dff_B_h1jjEvu12_1;
	wire w_dff_B_nmVmKBVL3_1;
	wire w_dff_B_QTPcrAO08_1;
	wire w_dff_B_KuOuFnyX7_1;
	wire w_dff_B_MFUfr5Qa6_1;
	wire w_dff_B_8qzSMwtE9_1;
	wire w_dff_B_mxmjQZhX3_1;
	wire w_dff_B_nOE1QFe26_1;
	wire w_dff_B_0YsZnwW28_1;
	wire w_dff_B_gfXIpjCS2_1;
	wire w_dff_B_6Yu3s5tv7_1;
	wire w_dff_B_8DQWRRrg3_1;
	wire w_dff_B_D82Loipc7_1;
	wire w_dff_B_8r3015HU7_1;
	wire w_dff_B_JtQLUTeL5_1;
	wire w_dff_B_8Cr0TDEK8_1;
	wire w_dff_B_delF4Zas1_1;
	wire w_dff_B_tbdtF29X5_1;
	wire w_dff_B_shH6qQGn7_1;
	wire w_dff_B_RpVWgE2a6_1;
	wire w_dff_B_hZ079ath5_1;
	wire w_dff_B_6VVkpMPZ1_1;
	wire w_dff_B_hFiHPxHv8_1;
	wire w_dff_B_faYWkUvB7_1;
	wire w_dff_B_ncU3zyj54_1;
	wire w_dff_B_b47Ey68k6_1;
	wire w_dff_B_04oEdqq83_1;
	wire w_dff_B_sYoD3wKb8_1;
	wire w_dff_B_U3ijMOQ21_1;
	wire w_dff_B_xuERZg8e0_1;
	wire w_dff_B_C0aIYlpK2_1;
	wire w_dff_B_AUKxi8sQ2_1;
	wire w_dff_B_MkIcXSec5_1;
	wire w_dff_B_hLk0iwCI2_1;
	wire w_dff_B_kAZSBhwF8_1;
	wire w_dff_B_car6Iadq0_1;
	wire w_dff_B_JQLYd7Gz9_1;
	wire w_dff_B_6TxBxlq59_1;
	wire w_dff_B_8j8EdYPm6_1;
	wire w_dff_B_eTmHU9F74_1;
	wire w_dff_B_vdi7sNWe8_1;
	wire w_dff_B_UVST5Psl6_1;
	wire w_dff_B_sV5OFSWG8_1;
	wire w_dff_B_TnQ11QdE6_1;
	wire w_dff_B_r7INjLgL2_1;
	wire w_dff_B_Vf8B4GpP1_1;
	wire w_dff_B_hvlMPTQU4_1;
	wire w_dff_B_o8Q9QmFf8_1;
	wire w_dff_B_VyhL9ZbR7_1;
	wire w_dff_B_Vx6SkBpy5_1;
	wire w_dff_B_V3roUK6J2_1;
	wire w_dff_B_j0hqHtfN0_1;
	wire w_dff_B_79PLedoF0_1;
	wire w_dff_B_IYp0UUHq6_1;
	wire w_dff_B_kANsNCpt4_1;
	wire w_dff_B_7PPvMfFA7_1;
	wire w_dff_B_I6WIoN6h9_0;
	wire w_dff_B_v20YfTkz6_0;
	wire w_dff_B_PfraoEG97_0;
	wire w_dff_B_imbyAO0c0_0;
	wire w_dff_B_W1o7TQaN3_0;
	wire w_dff_B_okqyDaim1_0;
	wire w_dff_B_OfCh70Dx4_0;
	wire w_dff_B_u4IfrlRY8_0;
	wire w_dff_B_tu2SQGoP4_0;
	wire w_dff_B_V96De1zx0_0;
	wire w_dff_B_6rRrfUwT2_0;
	wire w_dff_B_gleQx6wI2_0;
	wire w_dff_B_qf9QqL4M3_0;
	wire w_dff_B_mmjojyzO8_0;
	wire w_dff_B_PUgkccG65_0;
	wire w_dff_B_bzzPzEFh1_0;
	wire w_dff_B_LY3rvpL17_0;
	wire w_dff_B_zQxkMZYt4_0;
	wire w_dff_B_vtTpJuU04_0;
	wire w_dff_B_AcgPGI5J9_0;
	wire w_dff_B_3ISiST9S4_0;
	wire w_dff_B_Hny5F13O7_0;
	wire w_dff_B_KoMGABHe1_0;
	wire w_dff_B_AYmvd9PC9_0;
	wire w_dff_B_VTqx7xA56_0;
	wire w_dff_B_jFSt2hhA9_0;
	wire w_dff_B_2ElLLR002_0;
	wire w_dff_B_VBmHLkhk4_0;
	wire w_dff_B_uu8e0X9u2_0;
	wire w_dff_B_rxm1CEDV3_0;
	wire w_dff_B_POCj02fA0_0;
	wire w_dff_B_QZmL1ut17_0;
	wire w_dff_B_is1RNg5Z7_0;
	wire w_dff_B_F448UmfK5_0;
	wire w_dff_B_dYvtZ8Df4_0;
	wire w_dff_B_Jlo8iZXm1_0;
	wire w_dff_B_1lD11DCz5_0;
	wire w_dff_B_X7lFK10V4_0;
	wire w_dff_B_ByIfzr0X7_0;
	wire w_dff_B_IM7RNfKI9_0;
	wire w_dff_B_l25djXMi1_0;
	wire w_dff_B_NtXcXJe15_0;
	wire w_dff_B_7tdbdGb58_0;
	wire w_dff_B_b3nx18Dx2_0;
	wire w_dff_B_wSys2fMt6_0;
	wire w_dff_B_RQiFxszD5_0;
	wire w_dff_B_TJy3hCGi0_0;
	wire w_dff_B_QAVTeGs81_0;
	wire w_dff_B_SHZTPkSY3_0;
	wire w_dff_B_BVceaEl17_0;
	wire w_dff_B_oEZnnk893_0;
	wire w_dff_B_g2qzq5Uk0_0;
	wire w_dff_B_pZ0wTiXF3_0;
	wire w_dff_B_pRlFmw680_0;
	wire w_dff_B_PrE4Y01E3_0;
	wire w_dff_B_UPycdJTr5_0;
	wire w_dff_B_REgZMpD55_0;
	wire w_dff_B_kvaykdB33_0;
	wire w_dff_B_l5TD8cJi8_0;
	wire w_dff_B_bKY8m1741_0;
	wire w_dff_B_He72oM2c0_0;
	wire w_dff_B_1Nni3J8A7_0;
	wire w_dff_B_FQYrsurh4_0;
	wire w_dff_B_IKOjdOM87_0;
	wire w_dff_B_paRCc5t83_0;
	wire w_dff_B_RQgA9OTF1_0;
	wire w_dff_B_LscnLPzu1_0;
	wire w_dff_B_ZVOHQZK42_0;
	wire w_dff_B_iAHi3cHM6_0;
	wire w_dff_B_ccPsAbWf9_1;
	wire w_dff_B_dmbCAVom9_1;
	wire w_dff_B_MgeQSUbk5_1;
	wire w_dff_B_0DkQeKzB3_1;
	wire w_dff_B_24do6nwZ7_1;
	wire w_dff_B_5CsvRKcR9_1;
	wire w_dff_B_BwLXSL496_1;
	wire w_dff_B_X5SdyCPi4_1;
	wire w_dff_B_pBcaSdze7_1;
	wire w_dff_B_oF7TpXhf2_1;
	wire w_dff_B_0Jb9fXQB2_1;
	wire w_dff_B_uMDf2A0X9_1;
	wire w_dff_B_TgXIkbVz9_1;
	wire w_dff_B_bn0PNVvC9_1;
	wire w_dff_B_Rs4oPUVF0_1;
	wire w_dff_B_FgAafpcG0_1;
	wire w_dff_B_UwaFiXc28_1;
	wire w_dff_B_gm5GmJDo1_1;
	wire w_dff_B_bF6joxCt6_1;
	wire w_dff_B_P5K6vhlN1_1;
	wire w_dff_B_7ry2rKjK0_1;
	wire w_dff_B_lMzls0By5_1;
	wire w_dff_B_qtCAoueu8_1;
	wire w_dff_B_nyelgwX72_1;
	wire w_dff_B_RU54vTfO6_1;
	wire w_dff_B_dhGlGXz38_1;
	wire w_dff_B_TJvcmoAJ6_1;
	wire w_dff_B_VGuaFH3C4_1;
	wire w_dff_B_bCdNpNb82_1;
	wire w_dff_B_cd4ZdLXE0_1;
	wire w_dff_B_gCWmVbHO2_1;
	wire w_dff_B_uIH1LtwR0_1;
	wire w_dff_B_aBLe5VPw2_1;
	wire w_dff_B_Mew2iMBG1_1;
	wire w_dff_B_B1HOIyvz8_1;
	wire w_dff_B_x7a7HDjW2_1;
	wire w_dff_B_MVEgX4ZT6_1;
	wire w_dff_B_X6gl0TC57_1;
	wire w_dff_B_RnXb8XwF7_1;
	wire w_dff_B_WdejpLEj2_1;
	wire w_dff_B_tGg6C0Gf2_1;
	wire w_dff_B_bYaLPosM8_1;
	wire w_dff_B_96qtvItC4_1;
	wire w_dff_B_1DzZ794W0_1;
	wire w_dff_B_V0YdEzAl6_1;
	wire w_dff_B_u9Iyaxzs1_1;
	wire w_dff_B_10iTyhZc8_1;
	wire w_dff_B_jQCpIzdn1_1;
	wire w_dff_B_Y7qClh7w5_1;
	wire w_dff_B_Jl6hGn6p0_1;
	wire w_dff_B_rXbfx66U8_1;
	wire w_dff_B_pnOqBFsZ5_1;
	wire w_dff_B_PfcHVto03_1;
	wire w_dff_B_R5prVtWR3_1;
	wire w_dff_B_g0FnvyOO0_1;
	wire w_dff_B_X5WDxEki9_1;
	wire w_dff_B_6rFnZItM8_1;
	wire w_dff_B_rVcEjktx8_1;
	wire w_dff_B_bZcmDoP90_1;
	wire w_dff_B_9yJEvkvp4_1;
	wire w_dff_B_kbGi0tiY5_1;
	wire w_dff_B_qIt9bu6a7_1;
	wire w_dff_B_W5g0AisX0_1;
	wire w_dff_B_uccJS0r33_1;
	wire w_dff_B_zZI2lwkB3_1;
	wire w_dff_B_Q2rwYFRl1_1;
	wire w_dff_B_uEErvOl90_1;
	wire w_dff_B_qVRyJbno5_1;
	wire w_dff_B_Z7Sirpij6_0;
	wire w_dff_B_Xt0IZgU98_0;
	wire w_dff_B_SscclUei3_0;
	wire w_dff_B_06Ha8EZo0_0;
	wire w_dff_B_rW9Os9Be3_0;
	wire w_dff_B_aLTFwZJy5_0;
	wire w_dff_B_tNkFvcdR8_0;
	wire w_dff_B_tcxaZwbW0_0;
	wire w_dff_B_Q4pd3c0U9_0;
	wire w_dff_B_aEOuJAQW1_0;
	wire w_dff_B_sXlyN3LW9_0;
	wire w_dff_B_ysnb1nD20_0;
	wire w_dff_B_ZDo2W9112_0;
	wire w_dff_B_pH8Al40V3_0;
	wire w_dff_B_h3AyDBmA5_0;
	wire w_dff_B_BTcpYFCC2_0;
	wire w_dff_B_2TLyYWgn4_0;
	wire w_dff_B_1PXVEvfi7_0;
	wire w_dff_B_j9uYYPGg2_0;
	wire w_dff_B_FMkCthkR8_0;
	wire w_dff_B_OzMDdI7f5_0;
	wire w_dff_B_B3Qfqtdn6_0;
	wire w_dff_B_azkTL9Ge3_0;
	wire w_dff_B_167uqdjx2_0;
	wire w_dff_B_pbofjOQ73_0;
	wire w_dff_B_WBFFFfyu5_0;
	wire w_dff_B_lSLEwKtG5_0;
	wire w_dff_B_in8KpmEK3_0;
	wire w_dff_B_lpWVG82G3_0;
	wire w_dff_B_196kHsNn6_0;
	wire w_dff_B_DaWn44x37_0;
	wire w_dff_B_ixTnrwlj0_0;
	wire w_dff_B_TZ6t1DcZ9_0;
	wire w_dff_B_73Eyf9sN5_0;
	wire w_dff_B_JUgVaWZe5_0;
	wire w_dff_B_HQt7KFSI4_0;
	wire w_dff_B_nljmBTFz4_0;
	wire w_dff_B_XUqcbzYd3_0;
	wire w_dff_B_qEBXuOTc1_0;
	wire w_dff_B_0IUP9tQc4_0;
	wire w_dff_B_1N6TIWUA9_0;
	wire w_dff_B_NqEojNv73_0;
	wire w_dff_B_dZXrFEHE3_0;
	wire w_dff_B_fquEqgDn0_0;
	wire w_dff_B_NipIEUO12_0;
	wire w_dff_B_H2nginmZ3_0;
	wire w_dff_B_zNukDOmz4_0;
	wire w_dff_B_OcdQusVV4_0;
	wire w_dff_B_Z3I96UfL8_0;
	wire w_dff_B_GR16x9f84_0;
	wire w_dff_B_YWVEAJNb3_0;
	wire w_dff_B_DTwAlIz35_0;
	wire w_dff_B_pESVZrL72_0;
	wire w_dff_B_oIGVC5e15_0;
	wire w_dff_B_z9VmCxm43_0;
	wire w_dff_B_nAAcQ5dS9_0;
	wire w_dff_B_qBEN5rIH6_0;
	wire w_dff_B_LdGie02W9_0;
	wire w_dff_B_q6hamDKF4_0;
	wire w_dff_B_EWIV7aT86_0;
	wire w_dff_B_XgdVLFX05_0;
	wire w_dff_B_da93tegn2_0;
	wire w_dff_B_oTCFVaiB9_0;
	wire w_dff_B_yN0uHUf27_0;
	wire w_dff_B_Ql5QI0JW4_0;
	wire w_dff_B_4WKBwRrS5_0;
	wire w_dff_B_jLpXYLo19_0;
	wire w_dff_B_2OXQnYqp2_0;
	wire w_dff_B_GYLbdOCX1_1;
	wire w_dff_B_XTMiRIhg6_1;
	wire w_dff_B_fca62qz78_1;
	wire w_dff_B_CA96vvcK6_1;
	wire w_dff_B_AxC8Bn919_1;
	wire w_dff_B_VnGEQUVf8_1;
	wire w_dff_B_gz805dBu9_1;
	wire w_dff_B_OYSgM1FI7_1;
	wire w_dff_B_kVgENUOB3_1;
	wire w_dff_B_a5FLGmfM2_1;
	wire w_dff_B_pudAD3l09_1;
	wire w_dff_B_Ry7mGxoA4_1;
	wire w_dff_B_ayRfBUuD5_1;
	wire w_dff_B_8TdiQmeR0_1;
	wire w_dff_B_15tzuv726_1;
	wire w_dff_B_a4rhMODF8_1;
	wire w_dff_B_h5kncKbx2_1;
	wire w_dff_B_c7UWHLAU3_1;
	wire w_dff_B_vK6RYFCF5_1;
	wire w_dff_B_dV7qbMGB7_1;
	wire w_dff_B_nIhwms0s2_1;
	wire w_dff_B_5xgyrkik8_1;
	wire w_dff_B_kXpfZHYh6_1;
	wire w_dff_B_P4D5bdzx3_1;
	wire w_dff_B_nbDHKJqV7_1;
	wire w_dff_B_VBapY2Xc5_1;
	wire w_dff_B_m3ahZ0hv3_1;
	wire w_dff_B_npLZaldD7_1;
	wire w_dff_B_rY1AjtU16_1;
	wire w_dff_B_OB3r4e8T6_1;
	wire w_dff_B_3EkqwtWF6_1;
	wire w_dff_B_FlCYy9XC2_1;
	wire w_dff_B_7WQkiWTC5_1;
	wire w_dff_B_ekxYldbM2_1;
	wire w_dff_B_4nrSJw3b6_1;
	wire w_dff_B_eSczoEVk3_1;
	wire w_dff_B_VfiN7Kqr7_1;
	wire w_dff_B_yDWaDszt7_1;
	wire w_dff_B_KV7PT3no8_1;
	wire w_dff_B_Mamc8fYB6_1;
	wire w_dff_B_R7fWHnxx9_1;
	wire w_dff_B_ebdebRnl0_1;
	wire w_dff_B_IMkukUns7_1;
	wire w_dff_B_BHFm5u7A9_1;
	wire w_dff_B_Fh8EvCGF5_1;
	wire w_dff_B_aSirw5ni6_1;
	wire w_dff_B_MckXILbF5_1;
	wire w_dff_B_7b54I00q0_1;
	wire w_dff_B_ew2uIHn05_1;
	wire w_dff_B_E9YuMPL53_1;
	wire w_dff_B_JlnpJguO9_1;
	wire w_dff_B_t6xqW9AH7_1;
	wire w_dff_B_GUvPEhZy4_1;
	wire w_dff_B_fKPjesXu7_1;
	wire w_dff_B_QqPNInrF5_1;
	wire w_dff_B_9BafUZ3m2_1;
	wire w_dff_B_r4FeSYkW5_1;
	wire w_dff_B_qqW4rb7h8_1;
	wire w_dff_B_bd0Chshm7_1;
	wire w_dff_B_YNTY3V7G0_1;
	wire w_dff_B_bFmVn5FG1_1;
	wire w_dff_B_mfpjVyzb5_1;
	wire w_dff_B_Hqpq0lHO1_1;
	wire w_dff_B_q8PTZoPo1_1;
	wire w_dff_B_webqAdQe2_1;
	wire w_dff_B_xE1QwoiX4_1;
	wire w_dff_B_cSmyQJfw1_1;
	wire w_dff_B_2kuov4Ma5_0;
	wire w_dff_B_hgcS7yAr1_0;
	wire w_dff_B_VFTWXQwn3_0;
	wire w_dff_B_IyIOkS585_0;
	wire w_dff_B_J5TPWZ5A2_0;
	wire w_dff_B_xpa1SDpE3_0;
	wire w_dff_B_MEZD3l295_0;
	wire w_dff_B_pMjUpsoh0_0;
	wire w_dff_B_eCCIluiV0_0;
	wire w_dff_B_JcJcVjnT0_0;
	wire w_dff_B_Y3F6E1Cv9_0;
	wire w_dff_B_aUYGUOPZ0_0;
	wire w_dff_B_tmivuLWk9_0;
	wire w_dff_B_JHQmj32y2_0;
	wire w_dff_B_x6STL4N87_0;
	wire w_dff_B_f79Gd9jy3_0;
	wire w_dff_B_nT9Ppg2E5_0;
	wire w_dff_B_g4wSRRW03_0;
	wire w_dff_B_vcQEEfC96_0;
	wire w_dff_B_X1PT3bfU4_0;
	wire w_dff_B_zOmvvbsf7_0;
	wire w_dff_B_pa1ivYoB2_0;
	wire w_dff_B_gNrW1Hqd8_0;
	wire w_dff_B_VCz6KMAP0_0;
	wire w_dff_B_LIMABhSd5_0;
	wire w_dff_B_vzyPKbW73_0;
	wire w_dff_B_imAPqwS29_0;
	wire w_dff_B_bNVQeznS5_0;
	wire w_dff_B_LXjMrRfl1_0;
	wire w_dff_B_4GDqU3Y27_0;
	wire w_dff_B_L6Md8L6y4_0;
	wire w_dff_B_1JB8yVNP5_0;
	wire w_dff_B_gj84PKrv2_0;
	wire w_dff_B_WTAsiURZ6_0;
	wire w_dff_B_GqDHW8ku9_0;
	wire w_dff_B_arDvEw2o7_0;
	wire w_dff_B_9O6ALU7A7_0;
	wire w_dff_B_AyMsjAM11_0;
	wire w_dff_B_kSiyrEyt6_0;
	wire w_dff_B_nYpzzvIZ5_0;
	wire w_dff_B_BTwfQMWg4_0;
	wire w_dff_B_HcS9eDNk2_0;
	wire w_dff_B_bfB4mSgk7_0;
	wire w_dff_B_zqzTntQx4_0;
	wire w_dff_B_BPyDJHz75_0;
	wire w_dff_B_Zy20p5QQ9_0;
	wire w_dff_B_78wEVBwe5_0;
	wire w_dff_B_olI84OtP1_0;
	wire w_dff_B_mAjfHW8s2_0;
	wire w_dff_B_IJube8Tl3_0;
	wire w_dff_B_bLRExcag1_0;
	wire w_dff_B_otck3mYW7_0;
	wire w_dff_B_OW0lfqG68_0;
	wire w_dff_B_KLDZkxPv9_0;
	wire w_dff_B_0ioHCZkX2_0;
	wire w_dff_B_8wWhhm1t0_0;
	wire w_dff_B_Ye7Ynpi14_0;
	wire w_dff_B_4OiEwAw81_0;
	wire w_dff_B_tCwxgcz61_0;
	wire w_dff_B_n8ypLifR2_0;
	wire w_dff_B_9f3vnqCZ2_0;
	wire w_dff_B_q22xhbRt6_0;
	wire w_dff_B_8bx1wEvl6_0;
	wire w_dff_B_Ok9Fv8JV6_0;
	wire w_dff_B_SAdbhHjd5_0;
	wire w_dff_B_K3XBmhG19_0;
	wire w_dff_B_bDbh5nUT3_0;
	wire w_dff_B_56bX8R0X1_1;
	wire w_dff_B_J1VBtjpb7_1;
	wire w_dff_B_kT8blCOC1_1;
	wire w_dff_B_TSzDlOlD2_1;
	wire w_dff_B_mONv6dmT2_1;
	wire w_dff_B_zpmgjFJA0_1;
	wire w_dff_B_tOzNchBf7_1;
	wire w_dff_B_McKFDm483_1;
	wire w_dff_B_kN4zv8fZ9_1;
	wire w_dff_B_lkp6yAJk8_1;
	wire w_dff_B_Kx9gPkVX2_1;
	wire w_dff_B_knTFINpX0_1;
	wire w_dff_B_BdKWTzfq3_1;
	wire w_dff_B_ue7wsvFG8_1;
	wire w_dff_B_9ZMM5I1P3_1;
	wire w_dff_B_Btqj4csN3_1;
	wire w_dff_B_FuXT22V75_1;
	wire w_dff_B_9XYUF4Y51_1;
	wire w_dff_B_7fcbPlL34_1;
	wire w_dff_B_KbrJpvMN9_1;
	wire w_dff_B_wHeGzfyO0_1;
	wire w_dff_B_rbCrlYIc2_1;
	wire w_dff_B_XlYlYdku0_1;
	wire w_dff_B_LU0eBLHF4_1;
	wire w_dff_B_9KSkMU2o8_1;
	wire w_dff_B_wt0LdzhI8_1;
	wire w_dff_B_G8hwBcFe3_1;
	wire w_dff_B_Berkjg9t1_1;
	wire w_dff_B_7Rl9qeDe3_1;
	wire w_dff_B_EuE4d9l20_1;
	wire w_dff_B_NYdYAMfg2_1;
	wire w_dff_B_SJoVikYW5_1;
	wire w_dff_B_q6GBacby4_1;
	wire w_dff_B_JrXM8Gur7_1;
	wire w_dff_B_srMCdosz4_1;
	wire w_dff_B_4hKse7bY4_1;
	wire w_dff_B_TFs6LkqF2_1;
	wire w_dff_B_go67H1jV6_1;
	wire w_dff_B_c3DWREm90_1;
	wire w_dff_B_wcaO8rLs8_1;
	wire w_dff_B_Goglo8i51_1;
	wire w_dff_B_gxgFigMS6_1;
	wire w_dff_B_1MknRRtB0_1;
	wire w_dff_B_FYp2ifzv6_1;
	wire w_dff_B_tBEhIhY80_1;
	wire w_dff_B_URwioq5W9_1;
	wire w_dff_B_rH3K16z08_1;
	wire w_dff_B_Z4XxR2Vj7_1;
	wire w_dff_B_POg0RIHh7_1;
	wire w_dff_B_pB6jNztE3_1;
	wire w_dff_B_gAWATq4q7_1;
	wire w_dff_B_zmDSTPOg8_1;
	wire w_dff_B_7HZk2J4Z2_1;
	wire w_dff_B_x19aOJ4G4_1;
	wire w_dff_B_7YOlw7Rq5_1;
	wire w_dff_B_rADkxrbZ0_1;
	wire w_dff_B_xvXgV9UQ2_1;
	wire w_dff_B_CrMqGhrX5_1;
	wire w_dff_B_tazpeA5A9_1;
	wire w_dff_B_3mG95Zq31_1;
	wire w_dff_B_VeAwDMtq4_1;
	wire w_dff_B_qzF6vHka3_1;
	wire w_dff_B_CX5qG5KJ2_1;
	wire w_dff_B_jT6bcSwr0_1;
	wire w_dff_B_0jkwT1wb5_1;
	wire w_dff_B_SvQrjUup5_1;
	wire w_dff_B_lC8L2YxA4_0;
	wire w_dff_B_UPgIhrhr4_0;
	wire w_dff_B_51ulyRTI6_0;
	wire w_dff_B_IQ0VR6wP1_0;
	wire w_dff_B_ZjGJvPSI4_0;
	wire w_dff_B_tvqjYEwZ2_0;
	wire w_dff_B_Le8Canjh3_0;
	wire w_dff_B_lhdOWkJI7_0;
	wire w_dff_B_sfWgnykp5_0;
	wire w_dff_B_nQjRrXT37_0;
	wire w_dff_B_9dfk2v6l8_0;
	wire w_dff_B_4Sk6MFFu2_0;
	wire w_dff_B_0sNlxbt18_0;
	wire w_dff_B_0F3aU7Xk2_0;
	wire w_dff_B_IETck1EM7_0;
	wire w_dff_B_iDnLCt3V6_0;
	wire w_dff_B_oT6Q1veI4_0;
	wire w_dff_B_Qddfi4658_0;
	wire w_dff_B_asck50dK0_0;
	wire w_dff_B_xc1yyz7X4_0;
	wire w_dff_B_4WbD3Ruu4_0;
	wire w_dff_B_ygJPhuTH1_0;
	wire w_dff_B_t4ihs8jP1_0;
	wire w_dff_B_OOmlmDZy0_0;
	wire w_dff_B_q3sb1ZZ37_0;
	wire w_dff_B_fDvSImvh6_0;
	wire w_dff_B_eAv5gTy56_0;
	wire w_dff_B_tu1W32LA1_0;
	wire w_dff_B_4fpJw69N2_0;
	wire w_dff_B_j8top92t0_0;
	wire w_dff_B_giU7u6ow1_0;
	wire w_dff_B_ybnAhAMc9_0;
	wire w_dff_B_pEIs1MsE1_0;
	wire w_dff_B_Iv4h4NTC2_0;
	wire w_dff_B_uixhFbrS8_0;
	wire w_dff_B_VdGqVnLr0_0;
	wire w_dff_B_zQLbocjZ8_0;
	wire w_dff_B_7zcYi1To6_0;
	wire w_dff_B_v4lHygoC3_0;
	wire w_dff_B_proeNED82_0;
	wire w_dff_B_Ud0vc5AS6_0;
	wire w_dff_B_JAvHcDPl3_0;
	wire w_dff_B_x19qJt542_0;
	wire w_dff_B_Xo2I9Atg9_0;
	wire w_dff_B_dVLQmnYY3_0;
	wire w_dff_B_AlsrzvHm5_0;
	wire w_dff_B_zVmuojRz8_0;
	wire w_dff_B_gr65bRSH8_0;
	wire w_dff_B_Vih6pky98_0;
	wire w_dff_B_DREh6Ggg1_0;
	wire w_dff_B_kVLy3ipX6_0;
	wire w_dff_B_Di5LgRRX3_0;
	wire w_dff_B_kvlNU53N1_0;
	wire w_dff_B_0aMKTrjg4_0;
	wire w_dff_B_yFJWLOEU1_0;
	wire w_dff_B_6ZjTiqxA7_0;
	wire w_dff_B_JA9I5uAh1_0;
	wire w_dff_B_Vr1dtRmG6_0;
	wire w_dff_B_nFCXKPYZ1_0;
	wire w_dff_B_1TqtO5gz9_0;
	wire w_dff_B_vwtDePh67_0;
	wire w_dff_B_efUGQzXU9_0;
	wire w_dff_B_c2gXUocZ1_0;
	wire w_dff_B_a7wPIu1f1_0;
	wire w_dff_B_8SgZofGF7_0;
	wire w_dff_B_Mcr16eGs4_0;
	wire w_dff_B_7RUTZ4zU2_1;
	wire w_dff_B_zh4yBwlC6_1;
	wire w_dff_B_6kluDntq0_1;
	wire w_dff_B_69QmJAUD5_1;
	wire w_dff_B_eUsldsk62_1;
	wire w_dff_B_eDqPIPgc3_1;
	wire w_dff_B_CKXEPosv7_1;
	wire w_dff_B_g71M3N2a3_1;
	wire w_dff_B_ROXgn1xk4_1;
	wire w_dff_B_UBk1rUiz5_1;
	wire w_dff_B_grIg65Bo8_1;
	wire w_dff_B_3su8UvJ92_1;
	wire w_dff_B_y2O6myBI6_1;
	wire w_dff_B_JMfa18Nx5_1;
	wire w_dff_B_d1WlfRUu6_1;
	wire w_dff_B_Bgc7zlAf7_1;
	wire w_dff_B_tLE6cLRp7_1;
	wire w_dff_B_CiVge8Qz6_1;
	wire w_dff_B_hjHbACXu9_1;
	wire w_dff_B_iUWCiWiG5_1;
	wire w_dff_B_ym415l320_1;
	wire w_dff_B_RR2qjc2W0_1;
	wire w_dff_B_G7vkg4dJ7_1;
	wire w_dff_B_kfw8nkjS4_1;
	wire w_dff_B_L2I1VkNL2_1;
	wire w_dff_B_pCmAb4DC9_1;
	wire w_dff_B_CkGmlYcr0_1;
	wire w_dff_B_02oPRZOV9_1;
	wire w_dff_B_saTYnvjd4_1;
	wire w_dff_B_xSds98j35_1;
	wire w_dff_B_8G5Feubv2_1;
	wire w_dff_B_il0oKbyf7_1;
	wire w_dff_B_gKyPP9wD0_1;
	wire w_dff_B_2tFGeIHX4_1;
	wire w_dff_B_6IZBCQvH0_1;
	wire w_dff_B_3bwl2I039_1;
	wire w_dff_B_0bTe5xoN7_1;
	wire w_dff_B_gho2VcCs6_1;
	wire w_dff_B_3gaMNsXM6_1;
	wire w_dff_B_BbFk8HaN1_1;
	wire w_dff_B_ffg2xW9O3_1;
	wire w_dff_B_IeNIno6q0_1;
	wire w_dff_B_XBQnb87s0_1;
	wire w_dff_B_wgL2iy9s2_1;
	wire w_dff_B_ulxkTynz5_1;
	wire w_dff_B_iSyD2i7a9_1;
	wire w_dff_B_zVhLE4EG2_1;
	wire w_dff_B_mFwyxYtW1_1;
	wire w_dff_B_KqXYvtun4_1;
	wire w_dff_B_0zHvMaRL8_1;
	wire w_dff_B_FTiAOK5M1_1;
	wire w_dff_B_k13IfzzH0_1;
	wire w_dff_B_x5Xq9cFG9_1;
	wire w_dff_B_6yQkGmP23_1;
	wire w_dff_B_qzzrmTg50_1;
	wire w_dff_B_xMjyzten7_1;
	wire w_dff_B_uaBMf0Ov5_1;
	wire w_dff_B_rrrKqrcF5_1;
	wire w_dff_B_JsQwJtSs2_1;
	wire w_dff_B_O21dVdx15_1;
	wire w_dff_B_ZideBjrU7_1;
	wire w_dff_B_Gjyh2fKb3_1;
	wire w_dff_B_1rSLPhl06_1;
	wire w_dff_B_hKx3fuL67_1;
	wire w_dff_B_NsY7JH502_1;
	wire w_dff_B_GEUzZB1m6_0;
	wire w_dff_B_EgxhAFsZ9_0;
	wire w_dff_B_lmHDZMkk9_0;
	wire w_dff_B_NtrhFY9P1_0;
	wire w_dff_B_Era2yddZ9_0;
	wire w_dff_B_u1dbi5Aj6_0;
	wire w_dff_B_wfLV2Djz7_0;
	wire w_dff_B_p6vknCGc5_0;
	wire w_dff_B_rk60TxdO8_0;
	wire w_dff_B_wOTquhKX1_0;
	wire w_dff_B_cabrGrRQ6_0;
	wire w_dff_B_172tfGOf4_0;
	wire w_dff_B_AA3vfSq39_0;
	wire w_dff_B_ZVdcox9C2_0;
	wire w_dff_B_cspLt6N93_0;
	wire w_dff_B_EDBypqyU3_0;
	wire w_dff_B_4HkFUDsW2_0;
	wire w_dff_B_RKuAUXUZ9_0;
	wire w_dff_B_1USPPnLV9_0;
	wire w_dff_B_66L2saSR9_0;
	wire w_dff_B_WFUGenHp2_0;
	wire w_dff_B_uOZQLOrV2_0;
	wire w_dff_B_uW1X7DZu7_0;
	wire w_dff_B_hoaUnRl34_0;
	wire w_dff_B_hkM24vPM3_0;
	wire w_dff_B_l2EG3j3S2_0;
	wire w_dff_B_CfEy3taW2_0;
	wire w_dff_B_Skt9gxQk7_0;
	wire w_dff_B_y8oJOJv10_0;
	wire w_dff_B_Zp8rVhpO8_0;
	wire w_dff_B_sdxLvkqM2_0;
	wire w_dff_B_dz5ojoSk0_0;
	wire w_dff_B_D09QsuvI5_0;
	wire w_dff_B_vYWBSVrn3_0;
	wire w_dff_B_EQZcIIy48_0;
	wire w_dff_B_fPOg4O0G3_0;
	wire w_dff_B_ze07Q5ma2_0;
	wire w_dff_B_0xlaqssf2_0;
	wire w_dff_B_N9PkOXHb4_0;
	wire w_dff_B_M94hMR660_0;
	wire w_dff_B_W8njf6Rr0_0;
	wire w_dff_B_VHMMMsFQ0_0;
	wire w_dff_B_wViNcPEe6_0;
	wire w_dff_B_dmqzSnUX6_0;
	wire w_dff_B_do8guoy77_0;
	wire w_dff_B_IR1vPNZS1_0;
	wire w_dff_B_X2HsWHIV2_0;
	wire w_dff_B_uOFHBJ8Q2_0;
	wire w_dff_B_G6aAfiPF9_0;
	wire w_dff_B_m4LbWDCE6_0;
	wire w_dff_B_wGnGLw7v7_0;
	wire w_dff_B_JEVXnVFX1_0;
	wire w_dff_B_eD2NTRBl2_0;
	wire w_dff_B_m5t01a8u0_0;
	wire w_dff_B_FKoGc5pu2_0;
	wire w_dff_B_cLQrrrTq9_0;
	wire w_dff_B_8OAmP6dJ4_0;
	wire w_dff_B_JupuSsmG5_0;
	wire w_dff_B_ZYq0H2iY3_0;
	wire w_dff_B_blAMKkR16_0;
	wire w_dff_B_q2LgQ0Gs2_0;
	wire w_dff_B_SEkSkBZV6_0;
	wire w_dff_B_GAvcsof61_0;
	wire w_dff_B_m8F3KBwR0_0;
	wire w_dff_B_CuQ7QQJA6_0;
	wire w_dff_B_nS8rjJeB5_1;
	wire w_dff_B_VTPBg5wx6_1;
	wire w_dff_B_eBidpytV4_1;
	wire w_dff_B_Jj6e9lh24_1;
	wire w_dff_B_A7suurIY2_1;
	wire w_dff_B_hsOgVLe48_1;
	wire w_dff_B_yjjAjc7x8_1;
	wire w_dff_B_QpFQWZ810_1;
	wire w_dff_B_nQ7HpCc60_1;
	wire w_dff_B_AHIsHExp9_1;
	wire w_dff_B_I3MQ57Gs4_1;
	wire w_dff_B_FH0zwPGi3_1;
	wire w_dff_B_d78C6Lkt9_1;
	wire w_dff_B_Hz39arMe4_1;
	wire w_dff_B_2toyf6gO0_1;
	wire w_dff_B_S4z1YssN2_1;
	wire w_dff_B_w668kYAL8_1;
	wire w_dff_B_7Odta9Xs7_1;
	wire w_dff_B_FK8CKacm3_1;
	wire w_dff_B_A6gyFyOH3_1;
	wire w_dff_B_laPivbMg4_1;
	wire w_dff_B_vyb1i9MF2_1;
	wire w_dff_B_3KTwAvUB4_1;
	wire w_dff_B_zs3MaSr95_1;
	wire w_dff_B_7OdJvSyP8_1;
	wire w_dff_B_4jD6a6Bo2_1;
	wire w_dff_B_iNB1kBqi3_1;
	wire w_dff_B_IoUT6ftK3_1;
	wire w_dff_B_9TmBcy0q4_1;
	wire w_dff_B_NwqlbZuE0_1;
	wire w_dff_B_7PxXoN4N0_1;
	wire w_dff_B_spE9vrh28_1;
	wire w_dff_B_S176hAA30_1;
	wire w_dff_B_8AQbBgk44_1;
	wire w_dff_B_kqP8Zlwi1_1;
	wire w_dff_B_63wyduLu5_1;
	wire w_dff_B_tIK3KKXj6_1;
	wire w_dff_B_UJK6vTrf5_1;
	wire w_dff_B_2NviqDDV3_1;
	wire w_dff_B_AYUOc8Gs5_1;
	wire w_dff_B_j15IcKmA1_1;
	wire w_dff_B_OhtQOzVD0_1;
	wire w_dff_B_KLCzHLKu7_1;
	wire w_dff_B_MdeiuEh41_1;
	wire w_dff_B_5EvCmtn50_1;
	wire w_dff_B_SZYbdwEX3_1;
	wire w_dff_B_6oy73FDB8_1;
	wire w_dff_B_REoTtRit1_1;
	wire w_dff_B_9avp0UTU2_1;
	wire w_dff_B_hWNOZcnz8_1;
	wire w_dff_B_HEGWyX2r6_1;
	wire w_dff_B_nfwDGdAw9_1;
	wire w_dff_B_d6AQp35w2_1;
	wire w_dff_B_4jLjwKaP1_1;
	wire w_dff_B_H4M4vGHf9_1;
	wire w_dff_B_waGw9LyA0_1;
	wire w_dff_B_2Qva7Bku8_1;
	wire w_dff_B_j2zzwqhC0_1;
	wire w_dff_B_JUIiLmhv4_1;
	wire w_dff_B_dhkiUpHi9_1;
	wire w_dff_B_vuJXoeI63_1;
	wire w_dff_B_JYX8rV1H7_1;
	wire w_dff_B_8Wtnif2L2_1;
	wire w_dff_B_7KmGZ0V04_1;
	wire w_dff_B_8jvt49m20_0;
	wire w_dff_B_y8kKgoeP1_0;
	wire w_dff_B_0dx886Ab3_0;
	wire w_dff_B_sUlcGnsL9_0;
	wire w_dff_B_Wa7HuQ6Q1_0;
	wire w_dff_B_ZNWjGReA2_0;
	wire w_dff_B_PAZl7fDR1_0;
	wire w_dff_B_32Fn1vWW5_0;
	wire w_dff_B_uc1vmQNc3_0;
	wire w_dff_B_AQwrQfHK9_0;
	wire w_dff_B_bC5jBocF6_0;
	wire w_dff_B_ci4c5CF33_0;
	wire w_dff_B_nuzmbeWP1_0;
	wire w_dff_B_B7Hw1spn0_0;
	wire w_dff_B_mlnM6kO62_0;
	wire w_dff_B_EuUOriNB7_0;
	wire w_dff_B_gV2aYLZu5_0;
	wire w_dff_B_SzQKEmyD2_0;
	wire w_dff_B_CTKMIZTy8_0;
	wire w_dff_B_3gdFVuvg4_0;
	wire w_dff_B_cewDTCxe9_0;
	wire w_dff_B_XcDV76281_0;
	wire w_dff_B_zInW8uel6_0;
	wire w_dff_B_180jp84y5_0;
	wire w_dff_B_i6YDqOyM0_0;
	wire w_dff_B_pSF9T5Pf2_0;
	wire w_dff_B_bVFiigHL8_0;
	wire w_dff_B_lHP5kb4g2_0;
	wire w_dff_B_dYhXjvMW5_0;
	wire w_dff_B_zV3Bh9KR9_0;
	wire w_dff_B_p2uARIOa3_0;
	wire w_dff_B_PYTZ8VtL4_0;
	wire w_dff_B_EGkNCrWW0_0;
	wire w_dff_B_SV1DUznb6_0;
	wire w_dff_B_OOSxOqMm7_0;
	wire w_dff_B_0TrsDzSo0_0;
	wire w_dff_B_sOPMhTBd5_0;
	wire w_dff_B_qRRGCDx71_0;
	wire w_dff_B_kU4aM4Ij4_0;
	wire w_dff_B_isPekpHg1_0;
	wire w_dff_B_sUxngRBc5_0;
	wire w_dff_B_mO4k8g2u9_0;
	wire w_dff_B_zaxnlJSa6_0;
	wire w_dff_B_xBDjz1107_0;
	wire w_dff_B_WGiSRHLC9_0;
	wire w_dff_B_SiXnnu6K5_0;
	wire w_dff_B_aXmc2KFr1_0;
	wire w_dff_B_XQ8nriLS7_0;
	wire w_dff_B_zELcjJ1u1_0;
	wire w_dff_B_F516xxhK4_0;
	wire w_dff_B_LN8GzzQ85_0;
	wire w_dff_B_SDd9pG3g6_0;
	wire w_dff_B_n2BpADnQ6_0;
	wire w_dff_B_hYq1GgVC3_0;
	wire w_dff_B_le5p1kjZ9_0;
	wire w_dff_B_JcQE2Eb47_0;
	wire w_dff_B_G0PReR3J0_0;
	wire w_dff_B_9PGRykE52_0;
	wire w_dff_B_UEunsgaB1_0;
	wire w_dff_B_hx8YtgrH1_0;
	wire w_dff_B_KuEIbo5y0_0;
	wire w_dff_B_kits9ir32_0;
	wire w_dff_B_4e2hgKf74_0;
	wire w_dff_B_Xj7EsTj23_0;
	wire w_dff_B_7cu7BDBS8_1;
	wire w_dff_B_uDqwjLj17_1;
	wire w_dff_B_4Yb516S16_1;
	wire w_dff_B_2YcgcUE42_1;
	wire w_dff_B_odBgWBtx6_1;
	wire w_dff_B_cbCgOXKC4_1;
	wire w_dff_B_vhwz3dOr6_1;
	wire w_dff_B_PsA58lrt6_1;
	wire w_dff_B_imCIvpUZ8_1;
	wire w_dff_B_IdW1OJU97_1;
	wire w_dff_B_OsfbAIuW6_1;
	wire w_dff_B_z2fJUlJw0_1;
	wire w_dff_B_XCUHLsZ74_1;
	wire w_dff_B_j9NGT5YK2_1;
	wire w_dff_B_IGRL3lqn4_1;
	wire w_dff_B_vXANSm6S1_1;
	wire w_dff_B_gcJo1ROv2_1;
	wire w_dff_B_CjMoUz0g9_1;
	wire w_dff_B_aZ8nqmGT8_1;
	wire w_dff_B_A7PZ9GsO1_1;
	wire w_dff_B_iT5MW0qn5_1;
	wire w_dff_B_n9Ig3jhR8_1;
	wire w_dff_B_Cu5mas7q6_1;
	wire w_dff_B_I65WPdcW8_1;
	wire w_dff_B_kFN790u39_1;
	wire w_dff_B_S5lGZ8J95_1;
	wire w_dff_B_uIpOpjSU2_1;
	wire w_dff_B_2Isikgdt0_1;
	wire w_dff_B_1uaBUYjd8_1;
	wire w_dff_B_6BWM4xHe6_1;
	wire w_dff_B_D2t2dySb7_1;
	wire w_dff_B_z6WYQSXk4_1;
	wire w_dff_B_JWFXxkoL4_1;
	wire w_dff_B_FDYeKO5A5_1;
	wire w_dff_B_c8TtplOB7_1;
	wire w_dff_B_c0MzHVnU4_1;
	wire w_dff_B_TPpuQTEn7_1;
	wire w_dff_B_BVr4Ymur2_1;
	wire w_dff_B_Cx89FCXi5_1;
	wire w_dff_B_2hlkU6Dy2_1;
	wire w_dff_B_zwqOC2Hw2_1;
	wire w_dff_B_wuoZo4Q99_1;
	wire w_dff_B_m0kHz9zy9_1;
	wire w_dff_B_oZnF0VNm8_1;
	wire w_dff_B_vaqKKXb76_1;
	wire w_dff_B_n1oRl45p3_1;
	wire w_dff_B_VMz29ONC9_1;
	wire w_dff_B_bx9muena6_1;
	wire w_dff_B_0UuwdQhS5_1;
	wire w_dff_B_1imDCN9U1_1;
	wire w_dff_B_l6Oug9xJ1_1;
	wire w_dff_B_4fQmefUB9_1;
	wire w_dff_B_dKIuqhRF8_1;
	wire w_dff_B_saMclL7J2_1;
	wire w_dff_B_M5nzTvhP9_1;
	wire w_dff_B_bvtfSewb1_1;
	wire w_dff_B_15G1G7e40_1;
	wire w_dff_B_XMoTTNRF2_1;
	wire w_dff_B_QcjToezX0_1;
	wire w_dff_B_mXyo8GpD5_1;
	wire w_dff_B_oyx70XJx7_1;
	wire w_dff_B_4g3ciLln4_1;
	wire w_dff_B_HRhAL3Ck5_1;
	wire w_dff_B_Iq5SIEBg6_0;
	wire w_dff_B_bmrF8RiS9_0;
	wire w_dff_B_r7MNbbqV7_0;
	wire w_dff_B_gQHgiSjD3_0;
	wire w_dff_B_qnPmHTNX8_0;
	wire w_dff_B_TAEV7iu27_0;
	wire w_dff_B_SZ66MXMF7_0;
	wire w_dff_B_YHjvIQoi4_0;
	wire w_dff_B_xoksyxlb4_0;
	wire w_dff_B_KvxheGpT2_0;
	wire w_dff_B_Ea58jBqh6_0;
	wire w_dff_B_4Y4zcUxE3_0;
	wire w_dff_B_2kjiat809_0;
	wire w_dff_B_I780kHOK0_0;
	wire w_dff_B_7Xq193pV4_0;
	wire w_dff_B_zNDcUXjD9_0;
	wire w_dff_B_ZoZt7Vke9_0;
	wire w_dff_B_yAXdDuId3_0;
	wire w_dff_B_FNPm2xdt1_0;
	wire w_dff_B_MSY8yK4a2_0;
	wire w_dff_B_UllGlyU07_0;
	wire w_dff_B_yHPFuprz2_0;
	wire w_dff_B_uT4LyiFS9_0;
	wire w_dff_B_i90G6ENc0_0;
	wire w_dff_B_2VnWw6Lw7_0;
	wire w_dff_B_dgSVkDSR7_0;
	wire w_dff_B_yw9Aq1s27_0;
	wire w_dff_B_xiVuwzzH4_0;
	wire w_dff_B_ZOEY9g4g0_0;
	wire w_dff_B_8yuHZmbB1_0;
	wire w_dff_B_D11GE3nS0_0;
	wire w_dff_B_6Di2tpgr8_0;
	wire w_dff_B_gfZQfCSD6_0;
	wire w_dff_B_n1wrFb1w8_0;
	wire w_dff_B_cVAJMW9Z7_0;
	wire w_dff_B_5E48SLub1_0;
	wire w_dff_B_qsyeCCur8_0;
	wire w_dff_B_8rvzTbZY2_0;
	wire w_dff_B_gGh3ub9W9_0;
	wire w_dff_B_JtWItMy44_0;
	wire w_dff_B_CuhD3rm99_0;
	wire w_dff_B_tpLSu2OR1_0;
	wire w_dff_B_QSQ8UDAV1_0;
	wire w_dff_B_GrGS9iFN1_0;
	wire w_dff_B_MU7OR6QM1_0;
	wire w_dff_B_fflddMHi4_0;
	wire w_dff_B_1gjHNwWc6_0;
	wire w_dff_B_50W7jHId4_0;
	wire w_dff_B_D1TrHkD97_0;
	wire w_dff_B_RqaAzPuO6_0;
	wire w_dff_B_1FnkpiRx8_0;
	wire w_dff_B_TvPafgFc4_0;
	wire w_dff_B_oRv6gGLj3_0;
	wire w_dff_B_FZhMXYUO1_0;
	wire w_dff_B_AvlaCdJf9_0;
	wire w_dff_B_IGcHJelU4_0;
	wire w_dff_B_C1ixfA4R2_0;
	wire w_dff_B_dnzUGiSt8_0;
	wire w_dff_B_6qouszEI7_0;
	wire w_dff_B_ouioeusH9_0;
	wire w_dff_B_er01xbRt3_0;
	wire w_dff_B_pzmkeITL1_0;
	wire w_dff_B_J5sqkVLr6_0;
	wire w_dff_B_pCM6Lm6q5_1;
	wire w_dff_B_6g0XpZPS6_1;
	wire w_dff_B_HIcw1Ujt6_1;
	wire w_dff_B_JSWdv6P78_1;
	wire w_dff_B_q0KVr8gt5_1;
	wire w_dff_B_FAsyEvzp0_1;
	wire w_dff_B_FJCFVEKQ8_1;
	wire w_dff_B_4OO3EZD56_1;
	wire w_dff_B_RyX0zQpk7_1;
	wire w_dff_B_zeC7bnIP2_1;
	wire w_dff_B_TnpxSOum1_1;
	wire w_dff_B_M3WoWmAY6_1;
	wire w_dff_B_4MO54Gg99_1;
	wire w_dff_B_kJHuamjg4_1;
	wire w_dff_B_AZrgnmcb3_1;
	wire w_dff_B_WsjUi3Z02_1;
	wire w_dff_B_wnGOngvr1_1;
	wire w_dff_B_4o4fRPLS7_1;
	wire w_dff_B_GffUK5y29_1;
	wire w_dff_B_r3xQzSi28_1;
	wire w_dff_B_G4vRyjta4_1;
	wire w_dff_B_SoEiGnIc9_1;
	wire w_dff_B_cSy2rZTF5_1;
	wire w_dff_B_jcpNYGoa8_1;
	wire w_dff_B_V7x0HHom5_1;
	wire w_dff_B_YhIb3nKD3_1;
	wire w_dff_B_BSNDtTVs0_1;
	wire w_dff_B_8fXS1JJJ3_1;
	wire w_dff_B_bgE0axYw4_1;
	wire w_dff_B_5wZkBvJB4_1;
	wire w_dff_B_TSyG6yGQ7_1;
	wire w_dff_B_GnSoo2yZ0_1;
	wire w_dff_B_ApU1RraW2_1;
	wire w_dff_B_dXxRocCG3_1;
	wire w_dff_B_NyCSVVwW0_1;
	wire w_dff_B_SkTkYTez9_1;
	wire w_dff_B_ThLrF0L50_1;
	wire w_dff_B_EGNoTHZr6_1;
	wire w_dff_B_iAAgjrVY4_1;
	wire w_dff_B_Ch9Js3uL3_1;
	wire w_dff_B_BJJQJOLT0_1;
	wire w_dff_B_COHzw3Zv6_1;
	wire w_dff_B_QireFWjw0_1;
	wire w_dff_B_iDWWtNtt6_1;
	wire w_dff_B_NwnT28Ys4_1;
	wire w_dff_B_8w4rU8iO1_1;
	wire w_dff_B_Nnsn6uhN7_1;
	wire w_dff_B_sTCo5yyV6_1;
	wire w_dff_B_JfrxKUFD2_1;
	wire w_dff_B_hFcX7sdE2_1;
	wire w_dff_B_0Eg3HpmP6_1;
	wire w_dff_B_XiZ30F528_1;
	wire w_dff_B_SkJKHoaU3_1;
	wire w_dff_B_vkt6hixL8_1;
	wire w_dff_B_8C6yja3S5_1;
	wire w_dff_B_L2a0jLLv7_1;
	wire w_dff_B_3DIWUwOC8_1;
	wire w_dff_B_dsiL7QO31_1;
	wire w_dff_B_bZkssdEr2_1;
	wire w_dff_B_AoekRums7_1;
	wire w_dff_B_uPtNt3TD0_1;
	wire w_dff_B_cMTGAhWx0_1;
	wire w_dff_B_Gb948lxH1_0;
	wire w_dff_B_xCgC25rv5_0;
	wire w_dff_B_0T5yJljr6_0;
	wire w_dff_B_Cx6GdO1b6_0;
	wire w_dff_B_9FA9bqwa3_0;
	wire w_dff_B_omhxUjMQ2_0;
	wire w_dff_B_RWbulGMU8_0;
	wire w_dff_B_biOsRHvH5_0;
	wire w_dff_B_AajU3Poq2_0;
	wire w_dff_B_9k83aELm8_0;
	wire w_dff_B_twXb4y336_0;
	wire w_dff_B_nwoVfyvi7_0;
	wire w_dff_B_oTNcbAP31_0;
	wire w_dff_B_Mluztiq98_0;
	wire w_dff_B_NkpLAXM08_0;
	wire w_dff_B_2Oxc3Bb70_0;
	wire w_dff_B_fcvkr44d8_0;
	wire w_dff_B_GZpZuG998_0;
	wire w_dff_B_7bd4c1KM4_0;
	wire w_dff_B_g3XloexJ9_0;
	wire w_dff_B_zHKfXbTo6_0;
	wire w_dff_B_L79zxG8M9_0;
	wire w_dff_B_H7AFWyFd4_0;
	wire w_dff_B_MI2VsTuJ0_0;
	wire w_dff_B_R5A55xmn6_0;
	wire w_dff_B_bocE3cjN9_0;
	wire w_dff_B_3iMJ1vi79_0;
	wire w_dff_B_XH7l6pFw1_0;
	wire w_dff_B_xkz7X7su9_0;
	wire w_dff_B_P7Ttqsm60_0;
	wire w_dff_B_r78hXM8n4_0;
	wire w_dff_B_QnUHT7aa9_0;
	wire w_dff_B_Aaj1fTkD9_0;
	wire w_dff_B_NiN5AGtF5_0;
	wire w_dff_B_wlC7SorM1_0;
	wire w_dff_B_eSmT3Kxy0_0;
	wire w_dff_B_En9mGDM56_0;
	wire w_dff_B_JU8Pvl128_0;
	wire w_dff_B_qUFc0Ed45_0;
	wire w_dff_B_JPN8PLhI2_0;
	wire w_dff_B_IMtlwL1c8_0;
	wire w_dff_B_U9HNst065_0;
	wire w_dff_B_W0AM2YSI3_0;
	wire w_dff_B_NiNbrwPS6_0;
	wire w_dff_B_qPNot8fL7_0;
	wire w_dff_B_bTkhISM76_0;
	wire w_dff_B_3zXwjCk84_0;
	wire w_dff_B_qSeJNasX3_0;
	wire w_dff_B_VsC3ZK6P6_0;
	wire w_dff_B_mbanrVUj6_0;
	wire w_dff_B_mKZRQVP83_0;
	wire w_dff_B_ukn8lQJC0_0;
	wire w_dff_B_07t8K00Q6_0;
	wire w_dff_B_ln577FH27_0;
	wire w_dff_B_wAbb5i1f6_0;
	wire w_dff_B_PggIU1MR3_0;
	wire w_dff_B_csLlCdeo0_0;
	wire w_dff_B_1wKRBaic4_0;
	wire w_dff_B_A5xpSkoS7_0;
	wire w_dff_B_D316AO3t0_0;
	wire w_dff_B_M4MGvFqE3_0;
	wire w_dff_B_fIXrmCN75_0;
	wire w_dff_B_cJXCeA0y1_1;
	wire w_dff_B_59HshVZs5_1;
	wire w_dff_B_7TbwzYyW6_1;
	wire w_dff_B_VYJOMNCg2_1;
	wire w_dff_B_zyAYYDJ41_1;
	wire w_dff_B_KEu0eFlD6_1;
	wire w_dff_B_z3BTkWCm6_1;
	wire w_dff_B_IEYnuEbp6_1;
	wire w_dff_B_WocVIAZP4_1;
	wire w_dff_B_16KqC2lq3_1;
	wire w_dff_B_f52Galrs2_1;
	wire w_dff_B_79iSBHbn9_1;
	wire w_dff_B_MREGjirp4_1;
	wire w_dff_B_lcyCrvdg1_1;
	wire w_dff_B_cjHB07l78_1;
	wire w_dff_B_cQVTuwlt3_1;
	wire w_dff_B_NFXRdkBp2_1;
	wire w_dff_B_bw4tAdz56_1;
	wire w_dff_B_MmC0O3Jy9_1;
	wire w_dff_B_2m4yg1en4_1;
	wire w_dff_B_b9Pjx3a21_1;
	wire w_dff_B_MCwlDmhL0_1;
	wire w_dff_B_HkRpkuox2_1;
	wire w_dff_B_3EPNxRK11_1;
	wire w_dff_B_kMm4iLo02_1;
	wire w_dff_B_mwm4f3jj5_1;
	wire w_dff_B_2Z2DBqI25_1;
	wire w_dff_B_AMwvfgvg0_1;
	wire w_dff_B_Lm7HFJFP8_1;
	wire w_dff_B_CocpBhrM1_1;
	wire w_dff_B_bTMeguTl4_1;
	wire w_dff_B_dbV42ggt3_1;
	wire w_dff_B_X5Nj5lhu8_1;
	wire w_dff_B_3TZnnSnD0_1;
	wire w_dff_B_7qc1KcHe9_1;
	wire w_dff_B_gnWiF34h1_1;
	wire w_dff_B_6GIRifoM8_1;
	wire w_dff_B_HhwQyiw53_1;
	wire w_dff_B_3txzdJ769_1;
	wire w_dff_B_Vz5VF6nz6_1;
	wire w_dff_B_KLbxjjcm3_1;
	wire w_dff_B_phGo1tTR9_1;
	wire w_dff_B_yTcGv9Tp8_1;
	wire w_dff_B_SShyMNgN8_1;
	wire w_dff_B_yKFOmL6P5_1;
	wire w_dff_B_RkEsnCnM8_1;
	wire w_dff_B_m9lvf0eN6_1;
	wire w_dff_B_qc9FyenM2_1;
	wire w_dff_B_LNX9EyJ24_1;
	wire w_dff_B_wyWpdCvO3_1;
	wire w_dff_B_jmD3nOY58_1;
	wire w_dff_B_bi72tpfm5_1;
	wire w_dff_B_bVL4ArLi6_1;
	wire w_dff_B_OLHl6SlF6_1;
	wire w_dff_B_cC1TbIde8_1;
	wire w_dff_B_npTdC99a0_1;
	wire w_dff_B_BCnOsJAV2_1;
	wire w_dff_B_B2GyJLRl2_1;
	wire w_dff_B_zTg9Asyt2_1;
	wire w_dff_B_6HxPxKS97_1;
	wire w_dff_B_uGDXx6qa1_1;
	wire w_dff_B_iCIplsYd1_0;
	wire w_dff_B_R032ZZRg9_0;
	wire w_dff_B_lIV4UJEk4_0;
	wire w_dff_B_xTqWbW790_0;
	wire w_dff_B_ixbL4vuu8_0;
	wire w_dff_B_s5uNid6B0_0;
	wire w_dff_B_Gx1wuIWB0_0;
	wire w_dff_B_QLhEGMfl8_0;
	wire w_dff_B_GyKup3Yz8_0;
	wire w_dff_B_pG0Tfhxu4_0;
	wire w_dff_B_Y0MESBHd9_0;
	wire w_dff_B_0GCi309a2_0;
	wire w_dff_B_qr15E9pm1_0;
	wire w_dff_B_SviJMRe40_0;
	wire w_dff_B_98L6txer0_0;
	wire w_dff_B_pQ67VDW02_0;
	wire w_dff_B_Riw8sEhq4_0;
	wire w_dff_B_8d5uUr404_0;
	wire w_dff_B_2BDAb8Ld1_0;
	wire w_dff_B_gaPI7QpK9_0;
	wire w_dff_B_bckyv8fy8_0;
	wire w_dff_B_z2CUQsrk8_0;
	wire w_dff_B_UFE4WZqR9_0;
	wire w_dff_B_kc1zoTdG8_0;
	wire w_dff_B_Umk802Ry1_0;
	wire w_dff_B_zpBsNDiN3_0;
	wire w_dff_B_0jKSU1ix0_0;
	wire w_dff_B_koYusXgY5_0;
	wire w_dff_B_BoSNCSfl0_0;
	wire w_dff_B_NxkGtQvq7_0;
	wire w_dff_B_6Q9rhIwi3_0;
	wire w_dff_B_Md306bRj5_0;
	wire w_dff_B_Qbf0zgD62_0;
	wire w_dff_B_zvgZVG6U5_0;
	wire w_dff_B_7M3zvLsv9_0;
	wire w_dff_B_iGEiv4fl9_0;
	wire w_dff_B_bXOGno0P0_0;
	wire w_dff_B_mE0JMGW64_0;
	wire w_dff_B_LpsdSPht5_0;
	wire w_dff_B_4PbJHVNJ1_0;
	wire w_dff_B_KBNebchZ7_0;
	wire w_dff_B_ymRIN3jK2_0;
	wire w_dff_B_nsGtLrzT6_0;
	wire w_dff_B_eXgiMATL4_0;
	wire w_dff_B_eDqZ8lPw9_0;
	wire w_dff_B_otWcS33k2_0;
	wire w_dff_B_5NocYk2f2_0;
	wire w_dff_B_BHGDl4sJ3_0;
	wire w_dff_B_0ot5iYN30_0;
	wire w_dff_B_aB7eZaWZ9_0;
	wire w_dff_B_8uCdyeHM3_0;
	wire w_dff_B_yg1H9zqC3_0;
	wire w_dff_B_jUvToiwx6_0;
	wire w_dff_B_JAIq4SKV0_0;
	wire w_dff_B_CIQ32VdY8_0;
	wire w_dff_B_JYr9aXgA9_0;
	wire w_dff_B_PWDjvkGs6_0;
	wire w_dff_B_POJGLbQe0_0;
	wire w_dff_B_VobqMd4O4_0;
	wire w_dff_B_SLEJI2E67_0;
	wire w_dff_B_nUECFkPE3_0;
	wire w_dff_B_4r2a8qYn0_1;
	wire w_dff_B_Sly2Rx7X7_1;
	wire w_dff_B_hlydHVMl8_1;
	wire w_dff_B_yzeIPWWA1_1;
	wire w_dff_B_wPodME3e2_1;
	wire w_dff_B_7GjLbvzm7_1;
	wire w_dff_B_juRmGHoY0_1;
	wire w_dff_B_nDTvbOWK6_1;
	wire w_dff_B_p0CKGQ2U5_1;
	wire w_dff_B_lvVXzTXP7_1;
	wire w_dff_B_ojAQA5Aw1_1;
	wire w_dff_B_gDSCbj817_1;
	wire w_dff_B_mbs9phc69_1;
	wire w_dff_B_I94G633r6_1;
	wire w_dff_B_dnST0awd2_1;
	wire w_dff_B_IZg8B82I0_1;
	wire w_dff_B_gtrt0q9Z4_1;
	wire w_dff_B_jKTcvnDw0_1;
	wire w_dff_B_HT2QJnO22_1;
	wire w_dff_B_Ewicx5MI8_1;
	wire w_dff_B_7Uusi3WG0_1;
	wire w_dff_B_Pj6balu61_1;
	wire w_dff_B_Su5dXGqT0_1;
	wire w_dff_B_1CGdUx5Y7_1;
	wire w_dff_B_tDR81CLx2_1;
	wire w_dff_B_bs1PMIkH7_1;
	wire w_dff_B_Y7OhseaZ9_1;
	wire w_dff_B_BOeVL6ve7_1;
	wire w_dff_B_g0tsrqBD1_1;
	wire w_dff_B_h5QnmR809_1;
	wire w_dff_B_xRkDJq5h9_1;
	wire w_dff_B_WWKSD8Cq4_1;
	wire w_dff_B_Ig8YdTV84_1;
	wire w_dff_B_pXHdOA077_1;
	wire w_dff_B_t2l5o3Ta6_1;
	wire w_dff_B_boxmnPnb1_1;
	wire w_dff_B_HoysxmWq2_1;
	wire w_dff_B_cEPoh1h64_1;
	wire w_dff_B_u9DOPFVB9_1;
	wire w_dff_B_JmMp7Cdw4_1;
	wire w_dff_B_JQVCBCXc7_1;
	wire w_dff_B_pZzBcMIm0_1;
	wire w_dff_B_l9WmSUtg4_1;
	wire w_dff_B_WgfPajVu1_1;
	wire w_dff_B_mzaSY1Zu9_1;
	wire w_dff_B_OfoRcyLI7_1;
	wire w_dff_B_9ZXlClCf9_1;
	wire w_dff_B_M4UGntXx5_1;
	wire w_dff_B_LDXOTzf36_1;
	wire w_dff_B_yIbndY3H6_1;
	wire w_dff_B_A9D3q4lP5_1;
	wire w_dff_B_n5TTfjRT9_1;
	wire w_dff_B_LzQpxSza9_1;
	wire w_dff_B_NN0hhJfy2_1;
	wire w_dff_B_AZxMxgX31_1;
	wire w_dff_B_f9dMONXb3_1;
	wire w_dff_B_0HXGUKem9_1;
	wire w_dff_B_IBvWu3Eh6_1;
	wire w_dff_B_ma7LURTy0_1;
	wire w_dff_B_gZ9xFATs7_1;
	wire w_dff_B_bK7ToB561_0;
	wire w_dff_B_vrl6EvLN9_0;
	wire w_dff_B_iyGeSKHv5_0;
	wire w_dff_B_wKyKD5oY3_0;
	wire w_dff_B_xh3lNg544_0;
	wire w_dff_B_33RCGcIN7_0;
	wire w_dff_B_yAEvh6ME1_0;
	wire w_dff_B_TqNbQJRH0_0;
	wire w_dff_B_C7RB8ZTe4_0;
	wire w_dff_B_etSwmNbZ3_0;
	wire w_dff_B_uZAVrlBY3_0;
	wire w_dff_B_xe8Wi7jE8_0;
	wire w_dff_B_VOWqZwoz5_0;
	wire w_dff_B_zESnTcPO2_0;
	wire w_dff_B_OxueMZJc8_0;
	wire w_dff_B_pGG8WJUa9_0;
	wire w_dff_B_Oq0fkz0l7_0;
	wire w_dff_B_3RUhCgWm2_0;
	wire w_dff_B_iKVZ2m0e4_0;
	wire w_dff_B_HzNFQLS72_0;
	wire w_dff_B_6I4EmERV8_0;
	wire w_dff_B_EYevRhXP5_0;
	wire w_dff_B_CUAjfqae4_0;
	wire w_dff_B_OY5QezOA2_0;
	wire w_dff_B_xrVkakDe4_0;
	wire w_dff_B_o9dmVp507_0;
	wire w_dff_B_bwGMiDeP9_0;
	wire w_dff_B_jvm9tsOV5_0;
	wire w_dff_B_AVi0ttD09_0;
	wire w_dff_B_xTLU9toU0_0;
	wire w_dff_B_BUuWtqCV3_0;
	wire w_dff_B_VO0v5epf5_0;
	wire w_dff_B_oOuD9jeo5_0;
	wire w_dff_B_EXleF4Sd9_0;
	wire w_dff_B_kKqLcXHM0_0;
	wire w_dff_B_zbY4bD9a6_0;
	wire w_dff_B_zQyWVxrd6_0;
	wire w_dff_B_nmKAHa1f6_0;
	wire w_dff_B_3aWDFIBf9_0;
	wire w_dff_B_IEBmjdSg9_0;
	wire w_dff_B_Bjty1Tt67_0;
	wire w_dff_B_53aklnda2_0;
	wire w_dff_B_Bu79q6876_0;
	wire w_dff_B_1yWYUlkS8_0;
	wire w_dff_B_0XKY71Rh7_0;
	wire w_dff_B_0XRA4b5v2_0;
	wire w_dff_B_rpPTQowr0_0;
	wire w_dff_B_5TswgD3O8_0;
	wire w_dff_B_ckk5nHEA2_0;
	wire w_dff_B_lQqTLJ0Q0_0;
	wire w_dff_B_yXlWp8g34_0;
	wire w_dff_B_4J8UpfmA3_0;
	wire w_dff_B_xnoGFQho2_0;
	wire w_dff_B_83aPIXcz7_0;
	wire w_dff_B_UAS5stHz9_0;
	wire w_dff_B_TP3oONU42_0;
	wire w_dff_B_iPaydoqZ6_0;
	wire w_dff_B_Ryv6wlV94_0;
	wire w_dff_B_i64hvzJ48_0;
	wire w_dff_B_LsprbBuG0_0;
	wire w_dff_B_1Cx2caxz2_1;
	wire w_dff_B_vbRcEPTh3_1;
	wire w_dff_B_LvCxr4V80_1;
	wire w_dff_B_z3WnlphU0_1;
	wire w_dff_B_mn7LwfYp9_1;
	wire w_dff_B_KzmADoTA4_1;
	wire w_dff_B_QODcd1RD4_1;
	wire w_dff_B_5L3Io06b1_1;
	wire w_dff_B_K7cmhTgc0_1;
	wire w_dff_B_IoDvpxl32_1;
	wire w_dff_B_fv4E2Fld4_1;
	wire w_dff_B_sjdERbEs4_1;
	wire w_dff_B_zfoIswA72_1;
	wire w_dff_B_5l7hGFXW0_1;
	wire w_dff_B_bRSljdGJ7_1;
	wire w_dff_B_ZgQK24zP8_1;
	wire w_dff_B_naXpGiBI6_1;
	wire w_dff_B_JMiN8GXZ6_1;
	wire w_dff_B_HUg9T4C80_1;
	wire w_dff_B_eq6ugiHg7_1;
	wire w_dff_B_aPGmollr7_1;
	wire w_dff_B_mB9Nlvsz9_1;
	wire w_dff_B_ViyzJoYs0_1;
	wire w_dff_B_AtqpOaXn3_1;
	wire w_dff_B_FpYOZrTm9_1;
	wire w_dff_B_BHwGjug68_1;
	wire w_dff_B_DDfvJhH70_1;
	wire w_dff_B_y389G3vK0_1;
	wire w_dff_B_5FgpWpnl6_1;
	wire w_dff_B_U3JRfg9Z1_1;
	wire w_dff_B_ClW58C9k4_1;
	wire w_dff_B_FK5tsFwb2_1;
	wire w_dff_B_IYCZTfX03_1;
	wire w_dff_B_PCAzmfHq9_1;
	wire w_dff_B_wODzMxyA4_1;
	wire w_dff_B_1gQkhwGp9_1;
	wire w_dff_B_8Ue2Hj8O5_1;
	wire w_dff_B_90SkqCke5_1;
	wire w_dff_B_LaURsvA52_1;
	wire w_dff_B_K1nORJFn0_1;
	wire w_dff_B_3LbkweKt7_1;
	wire w_dff_B_J0NPgAzB3_1;
	wire w_dff_B_Datb44zb4_1;
	wire w_dff_B_0trhLKQ41_1;
	wire w_dff_B_JhjYVBbm1_1;
	wire w_dff_B_WU9ViVsG2_1;
	wire w_dff_B_sT70E6fh1_1;
	wire w_dff_B_g8JdIeNz5_1;
	wire w_dff_B_C8dI7RKM9_1;
	wire w_dff_B_dogrt0bY4_1;
	wire w_dff_B_VAGySKC93_1;
	wire w_dff_B_U7uE6QrZ9_1;
	wire w_dff_B_9aBkHysO8_1;
	wire w_dff_B_DWyBmJIV0_1;
	wire w_dff_B_ozCyyVsh4_1;
	wire w_dff_B_cI4GD7xH9_1;
	wire w_dff_B_0U4Zp4el5_1;
	wire w_dff_B_6BCzzzIk1_1;
	wire w_dff_B_NtYVoxbX5_1;
	wire w_dff_B_xMJ8Ciao7_0;
	wire w_dff_B_vSFhHKni3_0;
	wire w_dff_B_w1imK7my9_0;
	wire w_dff_B_pjCs8IJ28_0;
	wire w_dff_B_aNzkU1O32_0;
	wire w_dff_B_vYZOsSVd9_0;
	wire w_dff_B_DZYx8Q680_0;
	wire w_dff_B_0oRIfecE9_0;
	wire w_dff_B_JzWFCzIV0_0;
	wire w_dff_B_mltLMu050_0;
	wire w_dff_B_ZjHoYKYX7_0;
	wire w_dff_B_7xxrVNAZ8_0;
	wire w_dff_B_f6YrUZjQ6_0;
	wire w_dff_B_zrv7936S3_0;
	wire w_dff_B_GnqGi2xD8_0;
	wire w_dff_B_ubtHYmWE4_0;
	wire w_dff_B_AdTpG3142_0;
	wire w_dff_B_VNBffzMG2_0;
	wire w_dff_B_NIWY21Si3_0;
	wire w_dff_B_tu8JMW301_0;
	wire w_dff_B_qwIKNpJb1_0;
	wire w_dff_B_b68fVYw63_0;
	wire w_dff_B_MYI5QRP06_0;
	wire w_dff_B_mpMpEfFL5_0;
	wire w_dff_B_msFyOpjd9_0;
	wire w_dff_B_kUPQ2jMn5_0;
	wire w_dff_B_bTjTUVwT6_0;
	wire w_dff_B_WxdEABRo7_0;
	wire w_dff_B_lGW2T8n41_0;
	wire w_dff_B_1X46zTKq0_0;
	wire w_dff_B_QwWCDhRA2_0;
	wire w_dff_B_CdquVX552_0;
	wire w_dff_B_wkifLEgs5_0;
	wire w_dff_B_J60MzZXP7_0;
	wire w_dff_B_GzHbQOhD1_0;
	wire w_dff_B_tUntfrAW0_0;
	wire w_dff_B_Ey4vlT174_0;
	wire w_dff_B_YxR7vpTH6_0;
	wire w_dff_B_dpcinvtm0_0;
	wire w_dff_B_K9nMNI3k6_0;
	wire w_dff_B_6Pgs1x7T0_0;
	wire w_dff_B_0b8BnNLT3_0;
	wire w_dff_B_wqsYkcVq0_0;
	wire w_dff_B_SEL0GGUA1_0;
	wire w_dff_B_tjrxL4aE1_0;
	wire w_dff_B_UKmlommC3_0;
	wire w_dff_B_wVFqXuWr5_0;
	wire w_dff_B_UdpaqKrt7_0;
	wire w_dff_B_4gwA4mz83_0;
	wire w_dff_B_vkPQatIp2_0;
	wire w_dff_B_LvLXhLf50_0;
	wire w_dff_B_9yAIr1Ce7_0;
	wire w_dff_B_iH32c2aR6_0;
	wire w_dff_B_8aJjRu5i1_0;
	wire w_dff_B_FnTFnsir7_0;
	wire w_dff_B_JKwARmW67_0;
	wire w_dff_B_hxxUxdVp6_0;
	wire w_dff_B_LgOqTvTR3_0;
	wire w_dff_B_pQOVSYfd7_0;
	wire w_dff_B_QtN5qD899_1;
	wire w_dff_B_BhK3uIPd2_1;
	wire w_dff_B_nVyzy8dO1_1;
	wire w_dff_B_M2GbGVRc7_1;
	wire w_dff_B_rON9mXIN5_1;
	wire w_dff_B_ZbMvnJ8n7_1;
	wire w_dff_B_Ww93OQfn0_1;
	wire w_dff_B_Q8dcIBKq6_1;
	wire w_dff_B_2tNelLJL8_1;
	wire w_dff_B_9oDwAZwX2_1;
	wire w_dff_B_qytbBNr40_1;
	wire w_dff_B_DQzX6z0F2_1;
	wire w_dff_B_qsKPAzlQ3_1;
	wire w_dff_B_XaqLyrZn8_1;
	wire w_dff_B_gumfe9L20_1;
	wire w_dff_B_6pAGLQS84_1;
	wire w_dff_B_jyyO2smQ6_1;
	wire w_dff_B_QMgJQDr59_1;
	wire w_dff_B_UkEvQpEm5_1;
	wire w_dff_B_rxigErof6_1;
	wire w_dff_B_xBO1dK357_1;
	wire w_dff_B_rHaX9fF95_1;
	wire w_dff_B_GAd2QaDS8_1;
	wire w_dff_B_GclAZwzu5_1;
	wire w_dff_B_7vnjpK433_1;
	wire w_dff_B_qul3X06P7_1;
	wire w_dff_B_RwsYYg4w0_1;
	wire w_dff_B_PqEnw8Th4_1;
	wire w_dff_B_4hwD080H1_1;
	wire w_dff_B_GWk0qToj9_1;
	wire w_dff_B_tV5ewyNb8_1;
	wire w_dff_B_OFBrhHVk2_1;
	wire w_dff_B_ZPdKca7b7_1;
	wire w_dff_B_WMiaqdY48_1;
	wire w_dff_B_50aNQJna7_1;
	wire w_dff_B_YTBJ8uZ56_1;
	wire w_dff_B_ZEWd1Usu6_1;
	wire w_dff_B_Ro5PxidI0_1;
	wire w_dff_B_fxRK22Ws0_1;
	wire w_dff_B_ebgIrvys7_1;
	wire w_dff_B_BCWSgJn99_1;
	wire w_dff_B_vv69iHma1_1;
	wire w_dff_B_SpovpCDb4_1;
	wire w_dff_B_01gwM5td1_1;
	wire w_dff_B_3ydsrsbU9_1;
	wire w_dff_B_19EKRhkE9_1;
	wire w_dff_B_GPuZbTUg8_1;
	wire w_dff_B_KcXhrDlg6_1;
	wire w_dff_B_s7jEAdkM2_1;
	wire w_dff_B_m3mI4AfZ0_1;
	wire w_dff_B_LhlkRvhW5_1;
	wire w_dff_B_t3UiMecJ2_1;
	wire w_dff_B_c2MWpj7p1_1;
	wire w_dff_B_MmIq7VXG8_1;
	wire w_dff_B_92kAfPWp0_1;
	wire w_dff_B_PMoP7dQt5_1;
	wire w_dff_B_vdKdPBZQ8_1;
	wire w_dff_B_WezfSukm9_1;
	wire w_dff_B_3EbZKUZW6_0;
	wire w_dff_B_m5xhbG9y8_0;
	wire w_dff_B_xVRGVVqd6_0;
	wire w_dff_B_OLecySnw0_0;
	wire w_dff_B_RdAXibh13_0;
	wire w_dff_B_A5rMYJBz8_0;
	wire w_dff_B_qobfzLXL2_0;
	wire w_dff_B_Nyf5Y3g61_0;
	wire w_dff_B_Hkf1kb616_0;
	wire w_dff_B_kF2fPO3l1_0;
	wire w_dff_B_EvNMMVMc0_0;
	wire w_dff_B_EHP7Ju2R1_0;
	wire w_dff_B_nov3DkHn6_0;
	wire w_dff_B_skjKwW3f6_0;
	wire w_dff_B_rcR9tqwC3_0;
	wire w_dff_B_O1mV4QtD9_0;
	wire w_dff_B_mTyNPoAB0_0;
	wire w_dff_B_rv76iRzu1_0;
	wire w_dff_B_9BhQMxDU9_0;
	wire w_dff_B_E03CVzQb8_0;
	wire w_dff_B_3YGaRqIu4_0;
	wire w_dff_B_qOrN67cM1_0;
	wire w_dff_B_ZlhKjNc12_0;
	wire w_dff_B_dOn35z4Y0_0;
	wire w_dff_B_58atLflz6_0;
	wire w_dff_B_njGhdoid9_0;
	wire w_dff_B_58U6EFxH0_0;
	wire w_dff_B_GKoaAw8s3_0;
	wire w_dff_B_bAz2h1C45_0;
	wire w_dff_B_UO4rzyae3_0;
	wire w_dff_B_095kRksM1_0;
	wire w_dff_B_lcov63Po0_0;
	wire w_dff_B_V6tpfWNY7_0;
	wire w_dff_B_0pDBbWT35_0;
	wire w_dff_B_Lm5xfr8P1_0;
	wire w_dff_B_W3tYjjy10_0;
	wire w_dff_B_6as0KEqd5_0;
	wire w_dff_B_6CVVIedW9_0;
	wire w_dff_B_cgymDpta2_0;
	wire w_dff_B_OxTSltq28_0;
	wire w_dff_B_NYBhYppf2_0;
	wire w_dff_B_oMx0QT8S6_0;
	wire w_dff_B_84DNG2JZ9_0;
	wire w_dff_B_EWryNmyW9_0;
	wire w_dff_B_arYWH0Ma9_0;
	wire w_dff_B_ug4mcUrf6_0;
	wire w_dff_B_pPom2blk5_0;
	wire w_dff_B_8LByvSlY7_0;
	wire w_dff_B_vxmWHeNr3_0;
	wire w_dff_B_C0ENE8n84_0;
	wire w_dff_B_HRkudgNT9_0;
	wire w_dff_B_Gcz3vLz62_0;
	wire w_dff_B_EhHOQVgi4_0;
	wire w_dff_B_zJxe281o8_0;
	wire w_dff_B_vMQXSUN57_0;
	wire w_dff_B_Z2LiN9iz2_0;
	wire w_dff_B_nQBMPS0x9_0;
	wire w_dff_B_jX94jsrp1_0;
	wire w_dff_B_2Fh0fFQ36_1;
	wire w_dff_B_cna6aabl3_1;
	wire w_dff_B_8pNKKJkC4_1;
	wire w_dff_B_IEwzXTD45_1;
	wire w_dff_B_Lvyjbjhr6_1;
	wire w_dff_B_BvQqoA6l3_1;
	wire w_dff_B_wqk3qosK7_1;
	wire w_dff_B_4wpnnK5J2_1;
	wire w_dff_B_3Jf4ZWm04_1;
	wire w_dff_B_YwLuvEKI6_1;
	wire w_dff_B_4YHJtBmE0_1;
	wire w_dff_B_Vr3CkPg10_1;
	wire w_dff_B_eUPKISmw4_1;
	wire w_dff_B_jioS5rU41_1;
	wire w_dff_B_k4Cw3Myd1_1;
	wire w_dff_B_DZv0marw9_1;
	wire w_dff_B_AdoR8d0i0_1;
	wire w_dff_B_zUmhhjUJ0_1;
	wire w_dff_B_g0wot8bn0_1;
	wire w_dff_B_863NnPMp2_1;
	wire w_dff_B_bwXv3Nma9_1;
	wire w_dff_B_POVRJj548_1;
	wire w_dff_B_0V30eLpk9_1;
	wire w_dff_B_5gds8XUZ4_1;
	wire w_dff_B_lPqfSb8b0_1;
	wire w_dff_B_fipJqsSe8_1;
	wire w_dff_B_dLIrZH2K6_1;
	wire w_dff_B_4Rz9h9rD4_1;
	wire w_dff_B_S4w2GT5n6_1;
	wire w_dff_B_eQ1qDrA86_1;
	wire w_dff_B_eiYeq4ox4_1;
	wire w_dff_B_ou0RgOdy9_1;
	wire w_dff_B_gDyc3p8b0_1;
	wire w_dff_B_Hb4m2qnY3_1;
	wire w_dff_B_1K76nVgS4_1;
	wire w_dff_B_eoP3Yex09_1;
	wire w_dff_B_2Uj1LSKp3_1;
	wire w_dff_B_ghSR0Zmw4_1;
	wire w_dff_B_5RaPRw7l4_1;
	wire w_dff_B_27uAV64G6_1;
	wire w_dff_B_JgpuGL5Q5_1;
	wire w_dff_B_7N4MKayX3_1;
	wire w_dff_B_GhL8ah425_1;
	wire w_dff_B_IGujUGsJ2_1;
	wire w_dff_B_gesBFxlK8_1;
	wire w_dff_B_5Mzt9yVe4_1;
	wire w_dff_B_3672zwHl0_1;
	wire w_dff_B_OsJ4Xwr37_1;
	wire w_dff_B_MjGSkulR6_1;
	wire w_dff_B_TmOPLkar1_1;
	wire w_dff_B_T9xEWAhQ2_1;
	wire w_dff_B_c8fB6bqp0_1;
	wire w_dff_B_cjFPaJhc7_1;
	wire w_dff_B_do1dJ43T8_1;
	wire w_dff_B_lG5DkX6d0_1;
	wire w_dff_B_Tf7WMqGk9_1;
	wire w_dff_B_oG1alkJt9_1;
	wire w_dff_B_dBdjK4Go2_0;
	wire w_dff_B_wyPIm1UZ3_0;
	wire w_dff_B_BjFyTSEJ1_0;
	wire w_dff_B_jXLLyTQO5_0;
	wire w_dff_B_OMiCFaPv5_0;
	wire w_dff_B_OP7PK68l7_0;
	wire w_dff_B_FpX1ZdTa1_0;
	wire w_dff_B_8DMekzTk8_0;
	wire w_dff_B_G4sePo7S0_0;
	wire w_dff_B_t8rmk72t4_0;
	wire w_dff_B_LlxRW8C52_0;
	wire w_dff_B_Ky9pUCVw5_0;
	wire w_dff_B_Oy0NuylO8_0;
	wire w_dff_B_2noy2oTJ2_0;
	wire w_dff_B_dLBVVI7u3_0;
	wire w_dff_B_NRbQ4r6x2_0;
	wire w_dff_B_NBvesLd92_0;
	wire w_dff_B_K3H4kZND4_0;
	wire w_dff_B_MjByZoJH9_0;
	wire w_dff_B_56sHsrca8_0;
	wire w_dff_B_cwC5cs5I1_0;
	wire w_dff_B_g9qqL6A16_0;
	wire w_dff_B_TuWm4ZfD5_0;
	wire w_dff_B_4xiv5mHj9_0;
	wire w_dff_B_YRzchkIR9_0;
	wire w_dff_B_K74nRoLS3_0;
	wire w_dff_B_cLWezrlL6_0;
	wire w_dff_B_qcSg3F8k4_0;
	wire w_dff_B_3aZscX4A1_0;
	wire w_dff_B_s7nhyX6k9_0;
	wire w_dff_B_rTPn8nXI6_0;
	wire w_dff_B_kGnHDunW8_0;
	wire w_dff_B_dQRXvK4c9_0;
	wire w_dff_B_LPBJXOcQ8_0;
	wire w_dff_B_b5AQC59K3_0;
	wire w_dff_B_dhivIDxT2_0;
	wire w_dff_B_6vd3IVKb2_0;
	wire w_dff_B_P0g11IjR1_0;
	wire w_dff_B_DGjguLL43_0;
	wire w_dff_B_dTFCTEre2_0;
	wire w_dff_B_ciAR4HWn8_0;
	wire w_dff_B_IbE5Bi4l7_0;
	wire w_dff_B_Q59msCFu4_0;
	wire w_dff_B_jXcU14ww5_0;
	wire w_dff_B_eWohGabJ7_0;
	wire w_dff_B_T7F6FABL1_0;
	wire w_dff_B_2JdPZ1OT5_0;
	wire w_dff_B_4NRa4jZy9_0;
	wire w_dff_B_q8M4SDgg7_0;
	wire w_dff_B_NMOeFRYK4_0;
	wire w_dff_B_Ju8OmXTI0_0;
	wire w_dff_B_Iwn6LkHQ1_0;
	wire w_dff_B_pvhokLI60_0;
	wire w_dff_B_YdQR1MtD3_0;
	wire w_dff_B_MuFHsWWb0_0;
	wire w_dff_B_DJknTa6t8_0;
	wire w_dff_B_y4LeRC6T7_0;
	wire w_dff_B_GpWeFU1s5_1;
	wire w_dff_B_FgTKZoKY3_1;
	wire w_dff_B_aiiSi7yj2_1;
	wire w_dff_B_k9uGIfOT2_1;
	wire w_dff_B_VsnQUbqM6_1;
	wire w_dff_B_H86GVT4Y9_1;
	wire w_dff_B_noW4LybY3_1;
	wire w_dff_B_v5JRCwk38_1;
	wire w_dff_B_WZSkCvgY7_1;
	wire w_dff_B_zhg9jDwQ9_1;
	wire w_dff_B_dI8eMT2e2_1;
	wire w_dff_B_OOl40zg64_1;
	wire w_dff_B_a2jHVhPZ4_1;
	wire w_dff_B_2ew70LjY4_1;
	wire w_dff_B_2QNNBvTf6_1;
	wire w_dff_B_sFOQtUNk8_1;
	wire w_dff_B_87nCt9bA0_1;
	wire w_dff_B_buDyeB7T7_1;
	wire w_dff_B_6KmE9TuB0_1;
	wire w_dff_B_eVO0fgWg6_1;
	wire w_dff_B_NQZZxeGt0_1;
	wire w_dff_B_daK270jr9_1;
	wire w_dff_B_Ehbjd6Ch0_1;
	wire w_dff_B_MniuClbY7_1;
	wire w_dff_B_3uFndIfq4_1;
	wire w_dff_B_NGaQbojq4_1;
	wire w_dff_B_IiwrG0eu4_1;
	wire w_dff_B_v5Inhmz92_1;
	wire w_dff_B_3x5CRNck3_1;
	wire w_dff_B_dPvXVYw16_1;
	wire w_dff_B_x6ouehoS0_1;
	wire w_dff_B_Py0FRrTG8_1;
	wire w_dff_B_vZXReVgw5_1;
	wire w_dff_B_T7n84AaM3_1;
	wire w_dff_B_vYEUeJoc9_1;
	wire w_dff_B_2T110TmO9_1;
	wire w_dff_B_GCyTDkA14_1;
	wire w_dff_B_sNmnjWOY1_1;
	wire w_dff_B_YEnXssFw8_1;
	wire w_dff_B_0iwNGo6Z5_1;
	wire w_dff_B_9V7Hm9qW8_1;
	wire w_dff_B_pKtxPdUH5_1;
	wire w_dff_B_U05Knw5y5_1;
	wire w_dff_B_pzI1WzRe5_1;
	wire w_dff_B_98pEpBOP1_1;
	wire w_dff_B_3VVTgbij2_1;
	wire w_dff_B_dsFFpdN42_1;
	wire w_dff_B_QdYTwScb1_1;
	wire w_dff_B_IAurgHSJ4_1;
	wire w_dff_B_BgMUHX8R5_1;
	wire w_dff_B_yCjwOozj4_1;
	wire w_dff_B_OQj0EPzU8_1;
	wire w_dff_B_OUMAHm6x3_1;
	wire w_dff_B_CW9Chxyz6_1;
	wire w_dff_B_PhaSoyuf9_1;
	wire w_dff_B_7hG8iOrA5_1;
	wire w_dff_B_lCwjjydv0_0;
	wire w_dff_B_ucmcO5Ml9_0;
	wire w_dff_B_0mLqRJyn2_0;
	wire w_dff_B_7nWxuOlI8_0;
	wire w_dff_B_qAiuHkW09_0;
	wire w_dff_B_XoioK0yV9_0;
	wire w_dff_B_9GQ1TgWU3_0;
	wire w_dff_B_59gJDSWg4_0;
	wire w_dff_B_Fqri8rU17_0;
	wire w_dff_B_fusZp0wO4_0;
	wire w_dff_B_qfiPzsTJ0_0;
	wire w_dff_B_1IHRjypV6_0;
	wire w_dff_B_Mt73eZIK8_0;
	wire w_dff_B_L8tAwmN70_0;
	wire w_dff_B_Rg5dGiZJ9_0;
	wire w_dff_B_U09o2vKe9_0;
	wire w_dff_B_UBub5VMl4_0;
	wire w_dff_B_Y5Hjnyb33_0;
	wire w_dff_B_izX1EhWs3_0;
	wire w_dff_B_GFojTKFQ4_0;
	wire w_dff_B_HgByJuwt0_0;
	wire w_dff_B_AAhMz0cT7_0;
	wire w_dff_B_IVtehnJB2_0;
	wire w_dff_B_ppAay2wQ0_0;
	wire w_dff_B_fvd8OPgU6_0;
	wire w_dff_B_ud6T4sad7_0;
	wire w_dff_B_R2RMJGAo2_0;
	wire w_dff_B_Udu3LCzL3_0;
	wire w_dff_B_cPRnuFfU0_0;
	wire w_dff_B_VfYi89cV3_0;
	wire w_dff_B_crlkUjKD0_0;
	wire w_dff_B_lnwW7c1Z6_0;
	wire w_dff_B_MjnPmnjI0_0;
	wire w_dff_B_5rPxPaU28_0;
	wire w_dff_B_TAYMsVAj8_0;
	wire w_dff_B_m0gHZEVP0_0;
	wire w_dff_B_CHvgD6cr3_0;
	wire w_dff_B_Swy415Fb5_0;
	wire w_dff_B_rS4why0S1_0;
	wire w_dff_B_FAS5VmN86_0;
	wire w_dff_B_8bMGc5ws7_0;
	wire w_dff_B_TamJ9C3q4_0;
	wire w_dff_B_EDiQGhZA2_0;
	wire w_dff_B_tG9RCre11_0;
	wire w_dff_B_9HgKTcxd6_0;
	wire w_dff_B_jE0d3Y2q4_0;
	wire w_dff_B_IewIwsfG9_0;
	wire w_dff_B_u20dojIx1_0;
	wire w_dff_B_4pg06WGH8_0;
	wire w_dff_B_3KJRWdtl7_0;
	wire w_dff_B_EFceaqyR5_0;
	wire w_dff_B_J9OGBn7A9_0;
	wire w_dff_B_nN040jiK9_0;
	wire w_dff_B_tVW8F4P63_0;
	wire w_dff_B_qRjaLalN4_0;
	wire w_dff_B_3PM2Wo7i4_0;
	wire w_dff_B_u3TmHQQg3_1;
	wire w_dff_B_WyI1cjee2_1;
	wire w_dff_B_QwI2VE026_1;
	wire w_dff_B_f3OOC1vX5_1;
	wire w_dff_B_kObOhMPQ6_1;
	wire w_dff_B_UXXiYhTZ7_1;
	wire w_dff_B_vSzIN6NW1_1;
	wire w_dff_B_zx7wZkaR9_1;
	wire w_dff_B_qjQmHTsH3_1;
	wire w_dff_B_gxCBoZzF0_1;
	wire w_dff_B_T1Nxxa6N3_1;
	wire w_dff_B_aItBSbms7_1;
	wire w_dff_B_m9z39zzQ9_1;
	wire w_dff_B_wLFJeXXi6_1;
	wire w_dff_B_98y3Vefh8_1;
	wire w_dff_B_TOqFGqCT9_1;
	wire w_dff_B_WWse1KpF5_1;
	wire w_dff_B_QNEaobnf7_1;
	wire w_dff_B_mSkhTW764_1;
	wire w_dff_B_xMWIwYl62_1;
	wire w_dff_B_x02PzPzH6_1;
	wire w_dff_B_VLUkPEy28_1;
	wire w_dff_B_8sX3xPsl3_1;
	wire w_dff_B_GBVOD50H0_1;
	wire w_dff_B_jNtNys3P5_1;
	wire w_dff_B_OubD3WKZ2_1;
	wire w_dff_B_pcaQ4YbL7_1;
	wire w_dff_B_7Ni4p2F14_1;
	wire w_dff_B_URUERMh85_1;
	wire w_dff_B_KsDpCKZB3_1;
	wire w_dff_B_xx3DzdvC8_1;
	wire w_dff_B_3vi7eenL8_1;
	wire w_dff_B_xm2P1eNU0_1;
	wire w_dff_B_1hSD98Bj1_1;
	wire w_dff_B_31MJ7sCG5_1;
	wire w_dff_B_qFsfFMl80_1;
	wire w_dff_B_MVByffY11_1;
	wire w_dff_B_rlPV8eVZ9_1;
	wire w_dff_B_iVd6ZCv73_1;
	wire w_dff_B_XQftyCr26_1;
	wire w_dff_B_bCEJJ1tn6_1;
	wire w_dff_B_N7h1wGxT8_1;
	wire w_dff_B_YXV3KCnD0_1;
	wire w_dff_B_W7Dg6nDB7_1;
	wire w_dff_B_jdkH2UOj7_1;
	wire w_dff_B_Ra4Icv467_1;
	wire w_dff_B_oBUgjbJu4_1;
	wire w_dff_B_5LUFVdB82_1;
	wire w_dff_B_x8gIbswR4_1;
	wire w_dff_B_83yftHTo3_1;
	wire w_dff_B_5pXggwZi5_1;
	wire w_dff_B_S4ZFBNfZ5_1;
	wire w_dff_B_Eq02vrvz2_1;
	wire w_dff_B_ObDGcnQU8_1;
	wire w_dff_B_2n0kw3zB1_1;
	wire w_dff_B_EsGJzq0m3_0;
	wire w_dff_B_sU19rznP3_0;
	wire w_dff_B_IPWvB2Wl9_0;
	wire w_dff_B_6bizC6M54_0;
	wire w_dff_B_sCD3mHk49_0;
	wire w_dff_B_fhRiEnQz3_0;
	wire w_dff_B_bmpbmBlk3_0;
	wire w_dff_B_9umcwsmN4_0;
	wire w_dff_B_0IDKInX46_0;
	wire w_dff_B_LA6dKFUh9_0;
	wire w_dff_B_uAfYTa8O8_0;
	wire w_dff_B_g6jccsU59_0;
	wire w_dff_B_1iButynI2_0;
	wire w_dff_B_sQowIlt83_0;
	wire w_dff_B_PAiQ2VbV8_0;
	wire w_dff_B_jVnUIAVA9_0;
	wire w_dff_B_cINYgPb58_0;
	wire w_dff_B_rDEHEZWj5_0;
	wire w_dff_B_6KIz9v888_0;
	wire w_dff_B_JOgEGpBe8_0;
	wire w_dff_B_cUoiqd011_0;
	wire w_dff_B_n5qNuo1S7_0;
	wire w_dff_B_RmDJbPsU9_0;
	wire w_dff_B_sa9SjKqv1_0;
	wire w_dff_B_PBFYuqlC4_0;
	wire w_dff_B_hkSqgQ6W2_0;
	wire w_dff_B_TwtWAeLD6_0;
	wire w_dff_B_5YaTVtET9_0;
	wire w_dff_B_VftSinlm9_0;
	wire w_dff_B_bhnbH8kj1_0;
	wire w_dff_B_UxywJgzz8_0;
	wire w_dff_B_OtYc43D56_0;
	wire w_dff_B_LC9d0Ljk9_0;
	wire w_dff_B_gku3dSbK8_0;
	wire w_dff_B_Rbpqcn241_0;
	wire w_dff_B_FDtEjWJY3_0;
	wire w_dff_B_QUl09qph3_0;
	wire w_dff_B_AaQaOd5P7_0;
	wire w_dff_B_ovWruR753_0;
	wire w_dff_B_cgX8LBHo8_0;
	wire w_dff_B_rjylf6od7_0;
	wire w_dff_B_Bt632EuU5_0;
	wire w_dff_B_WMWMEPWe4_0;
	wire w_dff_B_3BR8YzSM9_0;
	wire w_dff_B_dk3ZerKI6_0;
	wire w_dff_B_i6kUDe318_0;
	wire w_dff_B_33Nb1gZU4_0;
	wire w_dff_B_EA8KARRM1_0;
	wire w_dff_B_vWQAAiWQ6_0;
	wire w_dff_B_WM0tBsn91_0;
	wire w_dff_B_z8rNMEFI7_0;
	wire w_dff_B_W4LRAtjG4_0;
	wire w_dff_B_n2SzxAAr1_0;
	wire w_dff_B_m5ibI5Kj7_0;
	wire w_dff_B_krSKQ8iz1_0;
	wire w_dff_B_b5cRaWfO3_1;
	wire w_dff_B_xlaGHZpv9_1;
	wire w_dff_B_gFzSFs251_1;
	wire w_dff_B_RAkB4lKs8_1;
	wire w_dff_B_J0A4sMAg3_1;
	wire w_dff_B_qITCs0Z54_1;
	wire w_dff_B_z81S9qzx5_1;
	wire w_dff_B_9O7j9BaX8_1;
	wire w_dff_B_eBqnDMTA3_1;
	wire w_dff_B_ZS581Y7Y7_1;
	wire w_dff_B_RNOrmn2G3_1;
	wire w_dff_B_GWmmUahR8_1;
	wire w_dff_B_5dtNx9NK9_1;
	wire w_dff_B_pHCAYkUu6_1;
	wire w_dff_B_6ooHb8145_1;
	wire w_dff_B_6z6YJeSJ8_1;
	wire w_dff_B_ZDPkAR0O8_1;
	wire w_dff_B_yV5BnaNt6_1;
	wire w_dff_B_aZkUgmSp5_1;
	wire w_dff_B_iNNRgKN24_1;
	wire w_dff_B_qvEcccPS0_1;
	wire w_dff_B_ogrzD7CN0_1;
	wire w_dff_B_V7mgggxv6_1;
	wire w_dff_B_0qy9Xb9k3_1;
	wire w_dff_B_hV2arTAE2_1;
	wire w_dff_B_0gg7424s5_1;
	wire w_dff_B_cN3qZ7nT9_1;
	wire w_dff_B_QmAHih4Q6_1;
	wire w_dff_B_lNAl2PBD8_1;
	wire w_dff_B_FEOjUxHq4_1;
	wire w_dff_B_GqgF33Vm5_1;
	wire w_dff_B_dpeDIHqQ1_1;
	wire w_dff_B_3GytPG7M5_1;
	wire w_dff_B_eYVPShpD2_1;
	wire w_dff_B_czpvQJoN5_1;
	wire w_dff_B_OwoURhs59_1;
	wire w_dff_B_BtgBJ39c3_1;
	wire w_dff_B_uwsbOTxx4_1;
	wire w_dff_B_Vnojznox4_1;
	wire w_dff_B_ZeRwnd7x6_1;
	wire w_dff_B_dtjxjMSz0_1;
	wire w_dff_B_jTDhGBs07_1;
	wire w_dff_B_PTcwSUUh3_1;
	wire w_dff_B_QnUnaBCc7_1;
	wire w_dff_B_GBGM6Wqj1_1;
	wire w_dff_B_ycVE9GKq1_1;
	wire w_dff_B_UM3geSuB2_1;
	wire w_dff_B_in75Yttl2_1;
	wire w_dff_B_sYnq7Z1t6_1;
	wire w_dff_B_G1EGA7eb7_1;
	wire w_dff_B_9TEw2b3a3_1;
	wire w_dff_B_7gPiBWga2_1;
	wire w_dff_B_Y1BbdXkY5_1;
	wire w_dff_B_o4QB8nIG6_1;
	wire w_dff_B_qgluD6W81_0;
	wire w_dff_B_P3tZvSFY8_0;
	wire w_dff_B_cjmn3daQ8_0;
	wire w_dff_B_lkP51Fe28_0;
	wire w_dff_B_RX372wIP1_0;
	wire w_dff_B_LODRxVuP3_0;
	wire w_dff_B_CMvbWlZI9_0;
	wire w_dff_B_Qw4zpn3i3_0;
	wire w_dff_B_XSkCxKzz4_0;
	wire w_dff_B_kdriNoI87_0;
	wire w_dff_B_U6JGT3CN0_0;
	wire w_dff_B_AYF1fGEB5_0;
	wire w_dff_B_NsXxB5lA3_0;
	wire w_dff_B_5EflqxPj3_0;
	wire w_dff_B_ltqeW4Ki0_0;
	wire w_dff_B_ktfDYClP5_0;
	wire w_dff_B_lt1VzINv0_0;
	wire w_dff_B_cc3jXEfG1_0;
	wire w_dff_B_bzOPL8I80_0;
	wire w_dff_B_qWehV0hB2_0;
	wire w_dff_B_xlDhjvz07_0;
	wire w_dff_B_pUaOUwjp9_0;
	wire w_dff_B_UIwajwPo0_0;
	wire w_dff_B_d0BF7Ojp6_0;
	wire w_dff_B_izH7tfVv4_0;
	wire w_dff_B_LfQudMwg9_0;
	wire w_dff_B_hhFLWRJV0_0;
	wire w_dff_B_OXUtnckG6_0;
	wire w_dff_B_eOyAxgCh7_0;
	wire w_dff_B_XVCZhUN09_0;
	wire w_dff_B_0v9ArSCW1_0;
	wire w_dff_B_Yw3riKHO0_0;
	wire w_dff_B_OtOLNGDa9_0;
	wire w_dff_B_yYSI4l345_0;
	wire w_dff_B_Ax22BgcJ8_0;
	wire w_dff_B_M1iRof4g1_0;
	wire w_dff_B_HqLo0pTa7_0;
	wire w_dff_B_ios72luL7_0;
	wire w_dff_B_S4FK22xX7_0;
	wire w_dff_B_KfRSqJR12_0;
	wire w_dff_B_4UyExW7n7_0;
	wire w_dff_B_eQU5zz4z1_0;
	wire w_dff_B_4oDxjTBS4_0;
	wire w_dff_B_Xo416V730_0;
	wire w_dff_B_Vqvyy7Tn2_0;
	wire w_dff_B_4xJChCV04_0;
	wire w_dff_B_Oi3s39gH7_0;
	wire w_dff_B_pIXfFVxd7_0;
	wire w_dff_B_ie4FZ6xV3_0;
	wire w_dff_B_LJi9gYe52_0;
	wire w_dff_B_UPmU200N5_0;
	wire w_dff_B_5KI7Y7LT5_0;
	wire w_dff_B_f3oqTQmX3_0;
	wire w_dff_B_PGiiN9Zt6_0;
	wire w_dff_B_3NitMkSn5_1;
	wire w_dff_B_TD2Z713j1_1;
	wire w_dff_B_fP6arkUA1_1;
	wire w_dff_B_5hibjoB12_1;
	wire w_dff_B_SBj1vHub8_1;
	wire w_dff_B_zbKmpZxD4_1;
	wire w_dff_B_lqY1FCXF4_1;
	wire w_dff_B_dM9s1a8J8_1;
	wire w_dff_B_LM3SgKNk9_1;
	wire w_dff_B_SDopu2EN1_1;
	wire w_dff_B_N4MNZalv6_1;
	wire w_dff_B_YiirUJhj9_1;
	wire w_dff_B_OwSdZTxt6_1;
	wire w_dff_B_2VqZHS2R7_1;
	wire w_dff_B_XHsRDCG96_1;
	wire w_dff_B_6q7Z3Cw30_1;
	wire w_dff_B_EkEgcoTD9_1;
	wire w_dff_B_hXtkLu3D3_1;
	wire w_dff_B_ZcVTmXbd9_1;
	wire w_dff_B_A1XMNnPh8_1;
	wire w_dff_B_WI4lMTSO2_1;
	wire w_dff_B_tREcRG0L5_1;
	wire w_dff_B_U0HNQjfI9_1;
	wire w_dff_B_mG0IVshm0_1;
	wire w_dff_B_t6azt6QS3_1;
	wire w_dff_B_dRas7cl43_1;
	wire w_dff_B_J8Lii8eP9_1;
	wire w_dff_B_Lvmat3IV1_1;
	wire w_dff_B_cIoF13n37_1;
	wire w_dff_B_WXyncf266_1;
	wire w_dff_B_SbnysYY39_1;
	wire w_dff_B_mB3fUMUv3_1;
	wire w_dff_B_NFX3FAcm5_1;
	wire w_dff_B_34KXOmbo1_1;
	wire w_dff_B_gntJ5zFW8_1;
	wire w_dff_B_Fd5aVKKW5_1;
	wire w_dff_B_V1Fzn0Hz3_1;
	wire w_dff_B_SHzVeHZz1_1;
	wire w_dff_B_ABl7DXHU3_1;
	wire w_dff_B_Oa0XLna62_1;
	wire w_dff_B_NSKaInd08_1;
	wire w_dff_B_jrGGJek59_1;
	wire w_dff_B_mD9wOaOj6_1;
	wire w_dff_B_XdEyA1PA6_1;
	wire w_dff_B_GUKttWlt3_1;
	wire w_dff_B_7TkwSu6j1_1;
	wire w_dff_B_MC81BYoT1_1;
	wire w_dff_B_pOxdbK7F9_1;
	wire w_dff_B_SGlrsFHN7_1;
	wire w_dff_B_BwevHhOt9_1;
	wire w_dff_B_aeNYWdBC5_1;
	wire w_dff_B_ASGowOXa9_1;
	wire w_dff_B_NmBOBsht4_1;
	wire w_dff_B_LZiz5Mk84_0;
	wire w_dff_B_Cg7oUIvo6_0;
	wire w_dff_B_qmpjg2xX3_0;
	wire w_dff_B_8MeaT4Re8_0;
	wire w_dff_B_rU1WovaH5_0;
	wire w_dff_B_cCDqW4AS3_0;
	wire w_dff_B_bSODKpen8_0;
	wire w_dff_B_59KfPeM54_0;
	wire w_dff_B_CQIrmEjv0_0;
	wire w_dff_B_M5z9CxST4_0;
	wire w_dff_B_uOUHpAvM3_0;
	wire w_dff_B_tFlWG7Wd3_0;
	wire w_dff_B_s4OlzC849_0;
	wire w_dff_B_jogyRlTu0_0;
	wire w_dff_B_8KxzbwZY6_0;
	wire w_dff_B_KZvx0bmv9_0;
	wire w_dff_B_ENkhQy1m6_0;
	wire w_dff_B_Q8vIP5FK5_0;
	wire w_dff_B_wvrTyQXF7_0;
	wire w_dff_B_qIg12tJV1_0;
	wire w_dff_B_4R10EknX2_0;
	wire w_dff_B_x6m6PfM41_0;
	wire w_dff_B_IuGJVSDc4_0;
	wire w_dff_B_EaB2OiFS9_0;
	wire w_dff_B_7tLK8jSy8_0;
	wire w_dff_B_abJ5S8bA8_0;
	wire w_dff_B_wyHXDwFz2_0;
	wire w_dff_B_nqfoKhld4_0;
	wire w_dff_B_UeIP226U6_0;
	wire w_dff_B_hMQyWIQ96_0;
	wire w_dff_B_rY8jcPou3_0;
	wire w_dff_B_77ox5Eyr9_0;
	wire w_dff_B_ARztImsF2_0;
	wire w_dff_B_9Ieo69JZ3_0;
	wire w_dff_B_yaH6cuNL9_0;
	wire w_dff_B_P9wUUOL93_0;
	wire w_dff_B_cDXCglxj5_0;
	wire w_dff_B_OiBhCLLK5_0;
	wire w_dff_B_PmXYMJ4Q5_0;
	wire w_dff_B_J8TpZcJc0_0;
	wire w_dff_B_cA507CoC5_0;
	wire w_dff_B_XjlxePQq2_0;
	wire w_dff_B_KdPouap28_0;
	wire w_dff_B_caKrQ1o24_0;
	wire w_dff_B_fiSm5DT83_0;
	wire w_dff_B_uocp1eZa9_0;
	wire w_dff_B_tlaMApI32_0;
	wire w_dff_B_yFCLzRZ81_0;
	wire w_dff_B_hNPlTbA14_0;
	wire w_dff_B_fy7XqznP4_0;
	wire w_dff_B_OOSx4D8S7_0;
	wire w_dff_B_YAYWLjIP7_0;
	wire w_dff_B_PKOhVjuX2_0;
	wire w_dff_B_UaRV9XiG9_1;
	wire w_dff_B_ai6QQYtD2_1;
	wire w_dff_B_6ulGzJuO0_1;
	wire w_dff_B_Yh8x01by5_1;
	wire w_dff_B_cZz7PcrI2_1;
	wire w_dff_B_HXraKzYR1_1;
	wire w_dff_B_hDoW6Imj0_1;
	wire w_dff_B_9BhmjCQ98_1;
	wire w_dff_B_z1A0BqMQ0_1;
	wire w_dff_B_cQw5Ygzh8_1;
	wire w_dff_B_geHnPb5o1_1;
	wire w_dff_B_rL0o6L9n1_1;
	wire w_dff_B_fGXVZiE07_1;
	wire w_dff_B_r5eIxA1C1_1;
	wire w_dff_B_5Zr7A37h7_1;
	wire w_dff_B_8YGySTQb1_1;
	wire w_dff_B_qkQiWXg85_1;
	wire w_dff_B_Lnf1Vxmy8_1;
	wire w_dff_B_gNg2Bj4n7_1;
	wire w_dff_B_F5BkbjlA0_1;
	wire w_dff_B_nSSjuBxj0_1;
	wire w_dff_B_jRNSO7Ad9_1;
	wire w_dff_B_CfZtREaj7_1;
	wire w_dff_B_pcNBA27f6_1;
	wire w_dff_B_YjQIUFxD7_1;
	wire w_dff_B_elgCwbZ71_1;
	wire w_dff_B_nOIukjqm0_1;
	wire w_dff_B_vSQHOlay9_1;
	wire w_dff_B_HagQRFEJ2_1;
	wire w_dff_B_moWyMS6c6_1;
	wire w_dff_B_FgbhDgid5_1;
	wire w_dff_B_YnndI7fC7_1;
	wire w_dff_B_8AjHEswg3_1;
	wire w_dff_B_omF8WcBY1_1;
	wire w_dff_B_4cQ0tuWt0_1;
	wire w_dff_B_y9xgnwPd1_1;
	wire w_dff_B_Ssa1m4iN3_1;
	wire w_dff_B_JRrVcOLQ0_1;
	wire w_dff_B_ym9V9iZV0_1;
	wire w_dff_B_vQyt8eDB7_1;
	wire w_dff_B_CWijj2xq6_1;
	wire w_dff_B_sYfMa7sh8_1;
	wire w_dff_B_zYeuVKsX5_1;
	wire w_dff_B_0qKHwpwa0_1;
	wire w_dff_B_LrrV8GhS1_1;
	wire w_dff_B_YxQft1Qn7_1;
	wire w_dff_B_GUSPqldz7_1;
	wire w_dff_B_tHHP3yKU1_1;
	wire w_dff_B_hlgryvHg4_1;
	wire w_dff_B_4o7gxzqN8_1;
	wire w_dff_B_cluyeuU07_1;
	wire w_dff_B_79nILaoK7_1;
	wire w_dff_B_pGUbVjsV3_0;
	wire w_dff_B_d3rqFy5D5_0;
	wire w_dff_B_BNdNpxkY9_0;
	wire w_dff_B_Jeo6SBNY1_0;
	wire w_dff_B_kOYnA20F5_0;
	wire w_dff_B_rGvnW9783_0;
	wire w_dff_B_kOfgVrCm8_0;
	wire w_dff_B_4vEHYa0W6_0;
	wire w_dff_B_1OLEl31J2_0;
	wire w_dff_B_bnqNQYyD9_0;
	wire w_dff_B_yI2g0aOB6_0;
	wire w_dff_B_8q1AVIyY0_0;
	wire w_dff_B_9uoMbIDX1_0;
	wire w_dff_B_90ENeEdu6_0;
	wire w_dff_B_wTcAe09v7_0;
	wire w_dff_B_PxMenEEx5_0;
	wire w_dff_B_KAVa2u9w1_0;
	wire w_dff_B_NZpfTpyH8_0;
	wire w_dff_B_1e1mwxTc2_0;
	wire w_dff_B_LBSYbJPY9_0;
	wire w_dff_B_FL3l4UmT4_0;
	wire w_dff_B_egqqIj7F9_0;
	wire w_dff_B_uGfySTqf5_0;
	wire w_dff_B_FBFGkjD36_0;
	wire w_dff_B_9bywbQDE0_0;
	wire w_dff_B_p0RUlMGR9_0;
	wire w_dff_B_NvXMLp5e8_0;
	wire w_dff_B_cIy6U2Dg3_0;
	wire w_dff_B_RpSPZDMK5_0;
	wire w_dff_B_cpjiHNqP9_0;
	wire w_dff_B_bo1EpKJ08_0;
	wire w_dff_B_0Jjtd9Ny6_0;
	wire w_dff_B_NRRVuZBu9_0;
	wire w_dff_B_9inLRKhL5_0;
	wire w_dff_B_10rHqYex3_0;
	wire w_dff_B_oQ31CafH6_0;
	wire w_dff_B_psv2ZGRp5_0;
	wire w_dff_B_S5DVYHzT2_0;
	wire w_dff_B_nHiGZgZ04_0;
	wire w_dff_B_XF69njg37_0;
	wire w_dff_B_vnNfoRqy5_0;
	wire w_dff_B_6job68c48_0;
	wire w_dff_B_ZvxRwRnz6_0;
	wire w_dff_B_ODhguznM4_0;
	wire w_dff_B_il1gIN9f0_0;
	wire w_dff_B_BD0PLByC2_0;
	wire w_dff_B_NjlY0O9g5_0;
	wire w_dff_B_VEx44Apl7_0;
	wire w_dff_B_DeHnzkIw8_0;
	wire w_dff_B_OJQ39A6f8_0;
	wire w_dff_B_YTJNs6OE9_0;
	wire w_dff_B_YyW5ipZv0_0;
	wire w_dff_B_bQJvc0Ve4_1;
	wire w_dff_B_zpqlmqQV7_1;
	wire w_dff_B_rXaYLGdB1_1;
	wire w_dff_B_tDQKSBf49_1;
	wire w_dff_B_ZgIzSM0g2_1;
	wire w_dff_B_EzlASfqV0_1;
	wire w_dff_B_zOtsgs4y5_1;
	wire w_dff_B_3HiJEepv8_1;
	wire w_dff_B_mH5nxX8w0_1;
	wire w_dff_B_yXRxkrjl3_1;
	wire w_dff_B_EsEpf7x14_1;
	wire w_dff_B_ePEQmxLZ0_1;
	wire w_dff_B_cwlunOWY5_1;
	wire w_dff_B_2raQsTBN5_1;
	wire w_dff_B_VtKk39hK5_1;
	wire w_dff_B_GDcWeBkl4_1;
	wire w_dff_B_0nDkNwCJ9_1;
	wire w_dff_B_xQaQhewD5_1;
	wire w_dff_B_NwSl4ljJ9_1;
	wire w_dff_B_fzFNLoXH8_1;
	wire w_dff_B_THQVFNnC3_1;
	wire w_dff_B_BVvyncLx5_1;
	wire w_dff_B_oBdoHUk20_1;
	wire w_dff_B_77BlTrmI7_1;
	wire w_dff_B_Akj4xQoO2_1;
	wire w_dff_B_F63teBN88_1;
	wire w_dff_B_I2cJFXtg8_1;
	wire w_dff_B_1cEWMqRE4_1;
	wire w_dff_B_okmk8ej78_1;
	wire w_dff_B_kkLOaFPG5_1;
	wire w_dff_B_EjC2iTcd4_1;
	wire w_dff_B_vHvRE9FN1_1;
	wire w_dff_B_BI742HCc7_1;
	wire w_dff_B_MqfxA0Lp3_1;
	wire w_dff_B_Nn016g5K1_1;
	wire w_dff_B_nfwkgyr70_1;
	wire w_dff_B_HYC4HdS17_1;
	wire w_dff_B_4Y4qqm3i7_1;
	wire w_dff_B_CozIy5H87_1;
	wire w_dff_B_06amHgLg0_1;
	wire w_dff_B_dlS9G38y9_1;
	wire w_dff_B_eCym5FEC1_1;
	wire w_dff_B_rmWpV3nV5_1;
	wire w_dff_B_fTEJk2RJ7_1;
	wire w_dff_B_YmAS7Fvg3_1;
	wire w_dff_B_ypTX0I4J3_1;
	wire w_dff_B_VLimmRyo2_1;
	wire w_dff_B_OmDnhRHM5_1;
	wire w_dff_B_ALskcCGj8_1;
	wire w_dff_B_qfGrphfe9_1;
	wire w_dff_B_YvJN65Kw3_1;
	wire w_dff_B_M2Z2Zpi32_0;
	wire w_dff_B_9BNZtYOb1_0;
	wire w_dff_B_urkHJcp67_0;
	wire w_dff_B_HYUQAbQz0_0;
	wire w_dff_B_6dR6rfDE6_0;
	wire w_dff_B_NdN26ESU3_0;
	wire w_dff_B_bcAtTlFa1_0;
	wire w_dff_B_cjyUP6Kr0_0;
	wire w_dff_B_3AjLE3qU1_0;
	wire w_dff_B_QfEyjW9I7_0;
	wire w_dff_B_I8jMhcO03_0;
	wire w_dff_B_k7RHcAAU8_0;
	wire w_dff_B_FAE4LRK28_0;
	wire w_dff_B_Tsy8CsY51_0;
	wire w_dff_B_qzVPgNDZ8_0;
	wire w_dff_B_Gezd239A1_0;
	wire w_dff_B_nyhxF0bx7_0;
	wire w_dff_B_d24qscAP0_0;
	wire w_dff_B_DDGoja6p3_0;
	wire w_dff_B_HLsuJNa15_0;
	wire w_dff_B_sTveYXAB5_0;
	wire w_dff_B_HidMJlhl6_0;
	wire w_dff_B_ls5QBqFE3_0;
	wire w_dff_B_RJOXyWdE1_0;
	wire w_dff_B_GPTPpF4S8_0;
	wire w_dff_B_jnx3XdYU8_0;
	wire w_dff_B_pD6aRnsO7_0;
	wire w_dff_B_U3E4HFq46_0;
	wire w_dff_B_lyp4tZrL0_0;
	wire w_dff_B_9hDLQRiJ7_0;
	wire w_dff_B_HoUpFYSE5_0;
	wire w_dff_B_TvI30jHQ4_0;
	wire w_dff_B_5V8MuIts4_0;
	wire w_dff_B_G1HHMFcq3_0;
	wire w_dff_B_KGGzbHOG1_0;
	wire w_dff_B_3F0HRwKR7_0;
	wire w_dff_B_UfRH370V6_0;
	wire w_dff_B_p0lZTIYI2_0;
	wire w_dff_B_6Sp6LpxQ3_0;
	wire w_dff_B_mYyvAyXV9_0;
	wire w_dff_B_qPvW9PJ80_0;
	wire w_dff_B_a5RrtU5Q3_0;
	wire w_dff_B_Tcb12aoD3_0;
	wire w_dff_B_JIoB9FaU8_0;
	wire w_dff_B_6YMK5mcd7_0;
	wire w_dff_B_K2CBbsIh3_0;
	wire w_dff_B_nDNyBPl96_0;
	wire w_dff_B_K3fYR1rs1_0;
	wire w_dff_B_4RgPXNwX4_0;
	wire w_dff_B_zD5kcOtr8_0;
	wire w_dff_B_pJXXJjmH2_0;
	wire w_dff_B_Bn0ayf4l4_1;
	wire w_dff_B_OPBHspa78_1;
	wire w_dff_B_bUr2KpR36_1;
	wire w_dff_B_wcblMY8k6_1;
	wire w_dff_B_icjOWe594_1;
	wire w_dff_B_gZfppW2h5_1;
	wire w_dff_B_si1WYAmm3_1;
	wire w_dff_B_zm2c9Z7N0_1;
	wire w_dff_B_72KwYpSV6_1;
	wire w_dff_B_8NxQKTM29_1;
	wire w_dff_B_d5auuZ082_1;
	wire w_dff_B_zUOcucZ45_1;
	wire w_dff_B_9Doe7fob0_1;
	wire w_dff_B_IItQNjhK6_1;
	wire w_dff_B_JjFlQL1Y5_1;
	wire w_dff_B_CNa3mE9S8_1;
	wire w_dff_B_CTxuITsz9_1;
	wire w_dff_B_AiRXKI9w3_1;
	wire w_dff_B_5UzYnNcM5_1;
	wire w_dff_B_UKfwHjPq0_1;
	wire w_dff_B_me5Mvwh82_1;
	wire w_dff_B_C7YKzlWL4_1;
	wire w_dff_B_SiCu6AZd6_1;
	wire w_dff_B_1f6dY7SB4_1;
	wire w_dff_B_cBkaatC65_1;
	wire w_dff_B_Py9Fyv2e4_1;
	wire w_dff_B_XR1rBt5N7_1;
	wire w_dff_B_TUCQCzOL1_1;
	wire w_dff_B_b9Fa4T0N5_1;
	wire w_dff_B_dLhp6r1k5_1;
	wire w_dff_B_KesjSdmP3_1;
	wire w_dff_B_y5dEn2zu7_1;
	wire w_dff_B_U8JxLU4j7_1;
	wire w_dff_B_rDJUI1sC4_1;
	wire w_dff_B_Xk4bNTa88_1;
	wire w_dff_B_n4Po8Bdw4_1;
	wire w_dff_B_srHselSA2_1;
	wire w_dff_B_OdB1l3Ip0_1;
	wire w_dff_B_wF9PpH6P0_1;
	wire w_dff_B_923Ba2Vi2_1;
	wire w_dff_B_t9LnWkL38_1;
	wire w_dff_B_R1frhqzv4_1;
	wire w_dff_B_XTZGcLFe9_1;
	wire w_dff_B_2bzqm8vX8_1;
	wire w_dff_B_giOac33U5_1;
	wire w_dff_B_juqi6SO07_1;
	wire w_dff_B_bkVmEFIp3_1;
	wire w_dff_B_NpUfs0ua2_1;
	wire w_dff_B_j6Xz2bdg7_1;
	wire w_dff_B_YfcGYVQq4_1;
	wire w_dff_B_o8lKl7m83_0;
	wire w_dff_B_m9OuHavv5_0;
	wire w_dff_B_gNsFavlC5_0;
	wire w_dff_B_GNFIWxiW6_0;
	wire w_dff_B_yztwk1Wg8_0;
	wire w_dff_B_J5gNqZO42_0;
	wire w_dff_B_jecSgOEO2_0;
	wire w_dff_B_nAMmXpDe1_0;
	wire w_dff_B_2CGPr0jL7_0;
	wire w_dff_B_C8aTMibt1_0;
	wire w_dff_B_oEasvFXR1_0;
	wire w_dff_B_jX7N9V0l2_0;
	wire w_dff_B_nhHmOG3l9_0;
	wire w_dff_B_2zfAyqfA1_0;
	wire w_dff_B_79j2RWhB7_0;
	wire w_dff_B_Mipow4lI7_0;
	wire w_dff_B_tgjkLOLF0_0;
	wire w_dff_B_M8j2y6Gb9_0;
	wire w_dff_B_GcV2SYhj9_0;
	wire w_dff_B_3wIQeuvn5_0;
	wire w_dff_B_6PdG8ZXr7_0;
	wire w_dff_B_nSRU9s8V7_0;
	wire w_dff_B_XQuVQhQs3_0;
	wire w_dff_B_0ZJBcOC74_0;
	wire w_dff_B_lTAhuV0P1_0;
	wire w_dff_B_iZTbxxbL3_0;
	wire w_dff_B_xNYiCHiy4_0;
	wire w_dff_B_ZdkeEZqT4_0;
	wire w_dff_B_6wYHZRJa3_0;
	wire w_dff_B_nLpqIPr92_0;
	wire w_dff_B_rypsM0rh5_0;
	wire w_dff_B_oJrbA7549_0;
	wire w_dff_B_2MgsdNv10_0;
	wire w_dff_B_nvUQFevb7_0;
	wire w_dff_B_Qz2Aludt3_0;
	wire w_dff_B_aFt5mB8r1_0;
	wire w_dff_B_nCJQ1OO02_0;
	wire w_dff_B_GOrBIJIZ5_0;
	wire w_dff_B_HWXM8W3R5_0;
	wire w_dff_B_0HvLrBnk7_0;
	wire w_dff_B_wMph96Ty8_0;
	wire w_dff_B_Bf7cOeaZ6_0;
	wire w_dff_B_tVxHdxMC3_0;
	wire w_dff_B_cCv8HaBD0_0;
	wire w_dff_B_0Tpg07rk5_0;
	wire w_dff_B_bKzotIXb8_0;
	wire w_dff_B_QTJk9WmN1_0;
	wire w_dff_B_XUO0cnc56_0;
	wire w_dff_B_zAV1WpsN2_0;
	wire w_dff_B_puRmXWhG3_0;
	wire w_dff_B_5kNCBtc74_1;
	wire w_dff_B_uoXHR67E5_1;
	wire w_dff_B_1ZwEeslb3_1;
	wire w_dff_B_Vu1XErOu6_1;
	wire w_dff_B_S0oXXYtW8_1;
	wire w_dff_B_8hiwjcQm3_1;
	wire w_dff_B_VaCA9vCu2_1;
	wire w_dff_B_NEOb3VVp4_1;
	wire w_dff_B_uxmPXaA96_1;
	wire w_dff_B_SeGm6zRR2_1;
	wire w_dff_B_plgHfCGH5_1;
	wire w_dff_B_C5jDYmwz1_1;
	wire w_dff_B_VwM0htNJ5_1;
	wire w_dff_B_0JdZOWma5_1;
	wire w_dff_B_wK7wchF66_1;
	wire w_dff_B_tDKb11eW6_1;
	wire w_dff_B_xLCAc80U8_1;
	wire w_dff_B_snmgibni4_1;
	wire w_dff_B_P3rbp7P50_1;
	wire w_dff_B_D5Y9nkM24_1;
	wire w_dff_B_7esFzaJc1_1;
	wire w_dff_B_Vj0rlalk2_1;
	wire w_dff_B_6YqNFGIg7_1;
	wire w_dff_B_v0ep1tLh9_1;
	wire w_dff_B_dkWHpMiA5_1;
	wire w_dff_B_N6bZIXBS3_1;
	wire w_dff_B_Vw5v93c62_1;
	wire w_dff_B_Y7f2ZDFI3_1;
	wire w_dff_B_nw43XgZG2_1;
	wire w_dff_B_2BrZbtDu9_1;
	wire w_dff_B_tokFQjsw5_1;
	wire w_dff_B_nulaadlk4_1;
	wire w_dff_B_wUKrFFBA3_1;
	wire w_dff_B_V4imVhSE2_1;
	wire w_dff_B_ifZ4tcSX1_1;
	wire w_dff_B_5B80bnKd4_1;
	wire w_dff_B_wtpp65Ik2_1;
	wire w_dff_B_zkt4Jsye9_1;
	wire w_dff_B_QTuSFALZ7_1;
	wire w_dff_B_Fflv2MGN1_1;
	wire w_dff_B_gSOESurT3_1;
	wire w_dff_B_zLpnZT2N8_1;
	wire w_dff_B_MS6rJ1o08_1;
	wire w_dff_B_1bb3jT2z7_1;
	wire w_dff_B_UxfLqzNf8_1;
	wire w_dff_B_rvgwMEOG7_1;
	wire w_dff_B_ftd9imrv6_1;
	wire w_dff_B_ITNKsc4Y9_1;
	wire w_dff_B_GecnHXzy9_1;
	wire w_dff_B_RYLpmxO94_0;
	wire w_dff_B_G13H5dCi3_0;
	wire w_dff_B_ezjcyRii5_0;
	wire w_dff_B_XVFFCW5k8_0;
	wire w_dff_B_1X2vffpK4_0;
	wire w_dff_B_5quM9VZJ2_0;
	wire w_dff_B_xqYvSQZX6_0;
	wire w_dff_B_OynyNYX33_0;
	wire w_dff_B_wmDOAMH98_0;
	wire w_dff_B_ymvk5kmL8_0;
	wire w_dff_B_jyUaxdDZ9_0;
	wire w_dff_B_TwIaURru0_0;
	wire w_dff_B_lVYmrqF10_0;
	wire w_dff_B_jQ2558Mk1_0;
	wire w_dff_B_96muY35c1_0;
	wire w_dff_B_zC14Kwyq9_0;
	wire w_dff_B_QnUjg5pl5_0;
	wire w_dff_B_Wn9SE4811_0;
	wire w_dff_B_arigDJuU6_0;
	wire w_dff_B_hHmelqxt8_0;
	wire w_dff_B_wDalVPYk4_0;
	wire w_dff_B_XgFvN2AZ3_0;
	wire w_dff_B_Idhox2Iw6_0;
	wire w_dff_B_5cvJRhJw0_0;
	wire w_dff_B_TYDBNPwG1_0;
	wire w_dff_B_46eipWmF1_0;
	wire w_dff_B_VQPO9YMH9_0;
	wire w_dff_B_nCrUplG55_0;
	wire w_dff_B_mise7VtT4_0;
	wire w_dff_B_9nz9xISJ3_0;
	wire w_dff_B_XEwqnxQC9_0;
	wire w_dff_B_9Y7rA5TP6_0;
	wire w_dff_B_50PypCeG2_0;
	wire w_dff_B_rqJwqihk6_0;
	wire w_dff_B_fhUqZg6j4_0;
	wire w_dff_B_3HJqArCw7_0;
	wire w_dff_B_uEFjUHwe5_0;
	wire w_dff_B_kYsVhlIg9_0;
	wire w_dff_B_gzPfgmdf1_0;
	wire w_dff_B_eQqM7EEQ8_0;
	wire w_dff_B_zKUvKSTu6_0;
	wire w_dff_B_H8PZzNAC0_0;
	wire w_dff_B_Rb4ms70y4_0;
	wire w_dff_B_uaqzDU7K0_0;
	wire w_dff_B_yvUUtoGq8_0;
	wire w_dff_B_6PmNXT3k8_0;
	wire w_dff_B_9D24XVkK7_0;
	wire w_dff_B_5p3UXoCp3_0;
	wire w_dff_B_CtINLd6Q5_0;
	wire w_dff_B_6sCSTLSj4_1;
	wire w_dff_B_GvGqxZ3V3_1;
	wire w_dff_B_hWFjEYmV3_1;
	wire w_dff_B_6crFkfLe6_1;
	wire w_dff_B_DjMlEltp7_1;
	wire w_dff_B_Gry2k59O3_1;
	wire w_dff_B_VYsM1v2D8_1;
	wire w_dff_B_VmyNWgjk3_1;
	wire w_dff_B_JDJFjqGW1_1;
	wire w_dff_B_DkBYT4ie2_1;
	wire w_dff_B_PwBl56if5_1;
	wire w_dff_B_yLKumY2s4_1;
	wire w_dff_B_KLAVQKdh3_1;
	wire w_dff_B_t4pfyRXO9_1;
	wire w_dff_B_Rqu0kexE4_1;
	wire w_dff_B_NIkRan838_1;
	wire w_dff_B_31ln5hJh9_1;
	wire w_dff_B_99R7wNjY7_1;
	wire w_dff_B_Rj55s4yc2_1;
	wire w_dff_B_FWEtqpvL3_1;
	wire w_dff_B_W78dtbey3_1;
	wire w_dff_B_pqhKhvzM5_1;
	wire w_dff_B_EEOq5RlS0_1;
	wire w_dff_B_WUkmjuyB8_1;
	wire w_dff_B_ExzLkwKL5_1;
	wire w_dff_B_wxpM6EWG3_1;
	wire w_dff_B_BePO5IXJ4_1;
	wire w_dff_B_5nJkuluL7_1;
	wire w_dff_B_LOqAfdhc0_1;
	wire w_dff_B_mc8q4U0a2_1;
	wire w_dff_B_oPu8Kb6S7_1;
	wire w_dff_B_7C3ASDbp1_1;
	wire w_dff_B_Yk31x2LH0_1;
	wire w_dff_B_k65tflB37_1;
	wire w_dff_B_ufgvtTPv4_1;
	wire w_dff_B_cifzNKpT5_1;
	wire w_dff_B_xojATAs66_1;
	wire w_dff_B_2s4vnN7u1_1;
	wire w_dff_B_3u3MEhQz3_1;
	wire w_dff_B_CrhhMABa3_1;
	wire w_dff_B_6zXPqvjK6_1;
	wire w_dff_B_ZvnD84cz9_1;
	wire w_dff_B_hFt9XGbI9_1;
	wire w_dff_B_I5dzgASW8_1;
	wire w_dff_B_ap2KaO5W2_1;
	wire w_dff_B_CWsNdAS21_1;
	wire w_dff_B_w8Vn2nOt6_1;
	wire w_dff_B_jwcKYoSU1_1;
	wire w_dff_B_40axs05m0_0;
	wire w_dff_B_OffUMx7R8_0;
	wire w_dff_B_Q8B2xwor8_0;
	wire w_dff_B_sGD3YZEY0_0;
	wire w_dff_B_kZ11lPUx2_0;
	wire w_dff_B_ISezBBuN8_0;
	wire w_dff_B_taLFUeXC6_0;
	wire w_dff_B_IgyaCaAn1_0;
	wire w_dff_B_XgiNsoNh7_0;
	wire w_dff_B_z3zWNLWx9_0;
	wire w_dff_B_CuBVRx4n9_0;
	wire w_dff_B_7Hc6tHMn0_0;
	wire w_dff_B_IYDyJz1m5_0;
	wire w_dff_B_fr9wnS0u6_0;
	wire w_dff_B_soMDuZBG4_0;
	wire w_dff_B_h8BXpw9J3_0;
	wire w_dff_B_RONKxCzt3_0;
	wire w_dff_B_xpjWN0uD0_0;
	wire w_dff_B_k0chVUju2_0;
	wire w_dff_B_aD44xSYH9_0;
	wire w_dff_B_7hruGXbF7_0;
	wire w_dff_B_QZPvQEjj7_0;
	wire w_dff_B_AGfo1Rsu2_0;
	wire w_dff_B_d1aLTJp94_0;
	wire w_dff_B_fxd2ASEM6_0;
	wire w_dff_B_8EJ4AQyt2_0;
	wire w_dff_B_QVV9mnIC8_0;
	wire w_dff_B_Buunm74Z4_0;
	wire w_dff_B_CZLvVthy3_0;
	wire w_dff_B_uAu4QFrV7_0;
	wire w_dff_B_36JBPEQP6_0;
	wire w_dff_B_gpGrFkiB2_0;
	wire w_dff_B_JE3xncqI2_0;
	wire w_dff_B_lA9ksrmU5_0;
	wire w_dff_B_rgWBQvSp3_0;
	wire w_dff_B_cH9MFqUT0_0;
	wire w_dff_B_ERfPkje79_0;
	wire w_dff_B_SzbEFIL33_0;
	wire w_dff_B_z8ogwEuY9_0;
	wire w_dff_B_xHe58wJT7_0;
	wire w_dff_B_35IDh1Zl0_0;
	wire w_dff_B_h8D3TgeQ2_0;
	wire w_dff_B_i1O2QFby3_0;
	wire w_dff_B_dM1kPNpR2_0;
	wire w_dff_B_uDBbSCPA7_0;
	wire w_dff_B_ms9K776m3_0;
	wire w_dff_B_VLbvT5nE1_0;
	wire w_dff_B_YAxWtq8t8_0;
	wire w_dff_B_vvWIz1QP5_1;
	wire w_dff_B_x6ed2YVm7_1;
	wire w_dff_B_vhBEouJ16_1;
	wire w_dff_B_JOnOab7Y5_1;
	wire w_dff_B_H8TNWflg5_1;
	wire w_dff_B_rYuSiGpX3_1;
	wire w_dff_B_PjNOFRsW3_1;
	wire w_dff_B_yzUMUqn91_1;
	wire w_dff_B_MPCpsYqI3_1;
	wire w_dff_B_NU2sOvR51_1;
	wire w_dff_B_CKTlIbPr3_1;
	wire w_dff_B_2Cj7x41M4_1;
	wire w_dff_B_FG7SWVwj6_1;
	wire w_dff_B_rR0cphWL9_1;
	wire w_dff_B_1h989HLm3_1;
	wire w_dff_B_QuJVjKsV6_1;
	wire w_dff_B_IKAiJwAl0_1;
	wire w_dff_B_WtPJZocd1_1;
	wire w_dff_B_QAdpB0jX0_1;
	wire w_dff_B_1Px8bGZx0_1;
	wire w_dff_B_vRPiREMc6_1;
	wire w_dff_B_kBMyCMHf2_1;
	wire w_dff_B_8Ezv7QT95_1;
	wire w_dff_B_sBBygfT39_1;
	wire w_dff_B_GW2KJw0R7_1;
	wire w_dff_B_jGursqEB5_1;
	wire w_dff_B_PQpomRoH7_1;
	wire w_dff_B_Ge2ue2aj0_1;
	wire w_dff_B_p1WsVsb60_1;
	wire w_dff_B_ZNo9H01j1_1;
	wire w_dff_B_Ty8hcaE66_1;
	wire w_dff_B_FZGIMHUy7_1;
	wire w_dff_B_qA0QAqjM5_1;
	wire w_dff_B_FHvAcDl31_1;
	wire w_dff_B_0gOv2HX11_1;
	wire w_dff_B_l8qcYsiU9_1;
	wire w_dff_B_WIxcTGWV3_1;
	wire w_dff_B_SKbqsVY74_1;
	wire w_dff_B_GCQuWFux6_1;
	wire w_dff_B_x5IXtwpv7_1;
	wire w_dff_B_2yyDiDP56_1;
	wire w_dff_B_GsfZAp0v5_1;
	wire w_dff_B_8Ynj0uPy0_1;
	wire w_dff_B_2FLoPUoD0_1;
	wire w_dff_B_RieSgn2L4_1;
	wire w_dff_B_jyOn7VFb8_1;
	wire w_dff_B_HGuNeMUK0_1;
	wire w_dff_B_X5L2oJc08_0;
	wire w_dff_B_hsMdZii72_0;
	wire w_dff_B_sFIILIqp7_0;
	wire w_dff_B_KqsKhx3Y1_0;
	wire w_dff_B_uJogh1Xe0_0;
	wire w_dff_B_wS9chUuM1_0;
	wire w_dff_B_rPv7w3865_0;
	wire w_dff_B_8KAfykP25_0;
	wire w_dff_B_NOPEF98n0_0;
	wire w_dff_B_sH6WML8f9_0;
	wire w_dff_B_wWCohYwY7_0;
	wire w_dff_B_4KyL94eA2_0;
	wire w_dff_B_ayAxIPLi7_0;
	wire w_dff_B_S1d0e5Lm2_0;
	wire w_dff_B_SxZayiWL5_0;
	wire w_dff_B_cC3Lp0en3_0;
	wire w_dff_B_YIIPcC1A9_0;
	wire w_dff_B_A4xCihqY4_0;
	wire w_dff_B_3xONO7RM1_0;
	wire w_dff_B_Xepa6ujA6_0;
	wire w_dff_B_LkWWh7pG9_0;
	wire w_dff_B_hr4JckW02_0;
	wire w_dff_B_yxJkppAV7_0;
	wire w_dff_B_t4NlzVy80_0;
	wire w_dff_B_XRwplYNf4_0;
	wire w_dff_B_7mztHKZu6_0;
	wire w_dff_B_5AhiBGHR0_0;
	wire w_dff_B_9G4rxd8p1_0;
	wire w_dff_B_sVtwLxFP0_0;
	wire w_dff_B_6uOiN1TZ0_0;
	wire w_dff_B_23IPDeYb4_0;
	wire w_dff_B_8O8qpHJS1_0;
	wire w_dff_B_GM8Q3bDK6_0;
	wire w_dff_B_0RpHrqHE3_0;
	wire w_dff_B_V7TIGBT59_0;
	wire w_dff_B_2D6U3nw51_0;
	wire w_dff_B_Xp7snU9d4_0;
	wire w_dff_B_so8Tqb4r7_0;
	wire w_dff_B_Maa3dE9Q0_0;
	wire w_dff_B_u8uo5R6K2_0;
	wire w_dff_B_RApRDQZK1_0;
	wire w_dff_B_Kn0gZBDs8_0;
	wire w_dff_B_kizdjsid5_0;
	wire w_dff_B_IgXKponO7_0;
	wire w_dff_B_YoVBKepe5_0;
	wire w_dff_B_7FHPGv6J7_0;
	wire w_dff_B_dL6uwy6j5_0;
	wire w_dff_B_RareMZ3a0_1;
	wire w_dff_B_yF59gkoW3_1;
	wire w_dff_B_tBiJ8S9k1_1;
	wire w_dff_B_jLAeV3cH0_1;
	wire w_dff_B_3wzp0HUu3_1;
	wire w_dff_B_CrgpEJ4p0_1;
	wire w_dff_B_6Ja2co3F4_1;
	wire w_dff_B_59DVj8Js9_1;
	wire w_dff_B_bJyV7eUw5_1;
	wire w_dff_B_3OZ1ouUr1_1;
	wire w_dff_B_bYOqyUOC4_1;
	wire w_dff_B_BNbpJa2r6_1;
	wire w_dff_B_gHbPwMYe9_1;
	wire w_dff_B_6gQnOMtJ9_1;
	wire w_dff_B_HEfMyAge5_1;
	wire w_dff_B_gbJFsDfJ5_1;
	wire w_dff_B_40aohpb96_1;
	wire w_dff_B_IZQeTgDk9_1;
	wire w_dff_B_FBiPRHqU8_1;
	wire w_dff_B_diTHVDpi4_1;
	wire w_dff_B_vKbaXYpi3_1;
	wire w_dff_B_cg8SRKwx1_1;
	wire w_dff_B_VRL8Nveg9_1;
	wire w_dff_B_SUNP9bmW7_1;
	wire w_dff_B_UCtUPBnI0_1;
	wire w_dff_B_UfQaruGv7_1;
	wire w_dff_B_LkXJbTM55_1;
	wire w_dff_B_JFCnja7Y7_1;
	wire w_dff_B_WeVK8C5h8_1;
	wire w_dff_B_lAsJRaTI5_1;
	wire w_dff_B_12mobeAb1_1;
	wire w_dff_B_zbkT3Di76_1;
	wire w_dff_B_CRcalJ793_1;
	wire w_dff_B_7eNX7ec42_1;
	wire w_dff_B_lIez84FE3_1;
	wire w_dff_B_P4nF0UWT6_1;
	wire w_dff_B_W62ryUpn4_1;
	wire w_dff_B_mHjw1S9M1_1;
	wire w_dff_B_oMqc1zsx4_1;
	wire w_dff_B_0Nh5DdFJ8_1;
	wire w_dff_B_aIL6VXuh6_1;
	wire w_dff_B_lmVL6hjy9_1;
	wire w_dff_B_gSQlFaGW5_1;
	wire w_dff_B_2fXr4ntQ1_1;
	wire w_dff_B_dT5YuAQX7_1;
	wire w_dff_B_ka8N4w5F3_1;
	wire w_dff_B_aBsTRinM6_0;
	wire w_dff_B_4EqVSWda4_0;
	wire w_dff_B_yOsaRBXF0_0;
	wire w_dff_B_Xj56PTnV0_0;
	wire w_dff_B_PXMx5Mmx9_0;
	wire w_dff_B_xNgy5rF84_0;
	wire w_dff_B_8Ci4NS0g4_0;
	wire w_dff_B_9YgRv75p1_0;
	wire w_dff_B_OACoJPxt3_0;
	wire w_dff_B_TRn10SlH3_0;
	wire w_dff_B_icnd60Cb2_0;
	wire w_dff_B_0FwPjB7W8_0;
	wire w_dff_B_vryRiryW3_0;
	wire w_dff_B_ZK0JBD3a4_0;
	wire w_dff_B_e7eddv003_0;
	wire w_dff_B_FjTq0QQM7_0;
	wire w_dff_B_IdUpPekU8_0;
	wire w_dff_B_dOBM42Mt6_0;
	wire w_dff_B_XjpTKGfm1_0;
	wire w_dff_B_yfMw7pnX1_0;
	wire w_dff_B_O6QePwCH2_0;
	wire w_dff_B_zrIknAPE4_0;
	wire w_dff_B_kHdafHAP4_0;
	wire w_dff_B_8zBUV71a6_0;
	wire w_dff_B_wfWOYZJ37_0;
	wire w_dff_B_KNhaQbf18_0;
	wire w_dff_B_O3YF9qtD9_0;
	wire w_dff_B_oP3PMArx1_0;
	wire w_dff_B_ycfeH6QV9_0;
	wire w_dff_B_zdHLg6hv5_0;
	wire w_dff_B_UmV4s7tZ3_0;
	wire w_dff_B_1HiDBbvd4_0;
	wire w_dff_B_JZZIy4KT8_0;
	wire w_dff_B_fjntXGqZ9_0;
	wire w_dff_B_vBqpgiy78_0;
	wire w_dff_B_dW4CplXG6_0;
	wire w_dff_B_VASnbmaW8_0;
	wire w_dff_B_FGMHauze8_0;
	wire w_dff_B_48aUyuVU1_0;
	wire w_dff_B_JyRHmNJl6_0;
	wire w_dff_B_60oyD4mx1_0;
	wire w_dff_B_UcLgOXrH5_0;
	wire w_dff_B_SxEj46qu5_0;
	wire w_dff_B_6cpYQZsk3_0;
	wire w_dff_B_8LNWvVGh4_0;
	wire w_dff_B_ZUFZvbyO9_0;
	wire w_dff_B_BfJV4Ur19_1;
	wire w_dff_B_xjnpz65V7_1;
	wire w_dff_B_4u32G6LM7_1;
	wire w_dff_B_PhsnOrBz1_1;
	wire w_dff_B_n3k8eKwb9_1;
	wire w_dff_B_Bhppne3H4_1;
	wire w_dff_B_BHZXVDlh5_1;
	wire w_dff_B_3DZdZwSO7_1;
	wire w_dff_B_qgjwp6H59_1;
	wire w_dff_B_FjISFoFn0_1;
	wire w_dff_B_eVP6afzg4_1;
	wire w_dff_B_dGAnLv7S1_1;
	wire w_dff_B_wrltKf9t8_1;
	wire w_dff_B_E6wfKDYf8_1;
	wire w_dff_B_zstLw8Pf6_1;
	wire w_dff_B_iJZwrhS32_1;
	wire w_dff_B_zW7vuYN68_1;
	wire w_dff_B_8qToVnRD6_1;
	wire w_dff_B_c3uE6Jvq8_1;
	wire w_dff_B_aFajiWuF4_1;
	wire w_dff_B_9SPTMo1L0_1;
	wire w_dff_B_UkSdvZEm2_1;
	wire w_dff_B_KuA1hRWS2_1;
	wire w_dff_B_mQKcb8SE7_1;
	wire w_dff_B_tLUqMK891_1;
	wire w_dff_B_qsRDDkov8_1;
	wire w_dff_B_g8KZL2Hr0_1;
	wire w_dff_B_qeGANq7a7_1;
	wire w_dff_B_MxjdNVv43_1;
	wire w_dff_B_dZSiIDYK9_1;
	wire w_dff_B_5aDJs0GN8_1;
	wire w_dff_B_6T6hcWBO8_1;
	wire w_dff_B_bTpRRFzg5_1;
	wire w_dff_B_YGtQo8gn1_1;
	wire w_dff_B_zrDe780f4_1;
	wire w_dff_B_rxgdsmxm4_1;
	wire w_dff_B_oKnqqtqY3_1;
	wire w_dff_B_GvHDDkT62_1;
	wire w_dff_B_UlL2W78Z6_1;
	wire w_dff_B_V41fX9643_1;
	wire w_dff_B_6bVTpYNH6_1;
	wire w_dff_B_yOlqlKDM7_1;
	wire w_dff_B_QdvKYQ2L9_1;
	wire w_dff_B_06brwXGZ0_1;
	wire w_dff_B_Fx8sXFkn9_1;
	wire w_dff_B_FbtI6Of34_0;
	wire w_dff_B_XDIlVbMV0_0;
	wire w_dff_B_eCaRibv90_0;
	wire w_dff_B_kW2IixvL6_0;
	wire w_dff_B_LfgYQ0ge5_0;
	wire w_dff_B_E23eIArt9_0;
	wire w_dff_B_uMppIBr96_0;
	wire w_dff_B_XoByUtor9_0;
	wire w_dff_B_N2Xmux2n4_0;
	wire w_dff_B_y7iCFvdQ0_0;
	wire w_dff_B_ZZ2qEJM67_0;
	wire w_dff_B_WhCYHgX61_0;
	wire w_dff_B_fRebIAFe5_0;
	wire w_dff_B_GHVhWHSr4_0;
	wire w_dff_B_Bxujhhbu5_0;
	wire w_dff_B_7Hpz5qb68_0;
	wire w_dff_B_Ccp5HXRm9_0;
	wire w_dff_B_s72c2n8R6_0;
	wire w_dff_B_2DLnntdb6_0;
	wire w_dff_B_QDRaTnnQ7_0;
	wire w_dff_B_WFGXknLw9_0;
	wire w_dff_B_AUaRfcRm1_0;
	wire w_dff_B_rXCzInwj3_0;
	wire w_dff_B_yaLJiO3n9_0;
	wire w_dff_B_5DQoXppv8_0;
	wire w_dff_B_5s19uiwV6_0;
	wire w_dff_B_xuj8m10v6_0;
	wire w_dff_B_rlN7NpqB4_0;
	wire w_dff_B_46Uwhuwb6_0;
	wire w_dff_B_z4UHXo5W6_0;
	wire w_dff_B_6dwXgyjx3_0;
	wire w_dff_B_YmFpfVVW8_0;
	wire w_dff_B_TU7GA8Qi2_0;
	wire w_dff_B_W9Xb6OZx8_0;
	wire w_dff_B_2UNFf4Ty5_0;
	wire w_dff_B_IDcAj2xk5_0;
	wire w_dff_B_IIK19u7o6_0;
	wire w_dff_B_cgSfWJbn2_0;
	wire w_dff_B_5uh1eMy41_0;
	wire w_dff_B_ltZQHJzB0_0;
	wire w_dff_B_picAWtcF3_0;
	wire w_dff_B_yOnKICW88_0;
	wire w_dff_B_AaGCz7o39_0;
	wire w_dff_B_Tc3H8Sc58_0;
	wire w_dff_B_ru1ByfvL1_0;
	wire w_dff_B_ZbhWhr9i0_1;
	wire w_dff_B_pwsoJJEN3_1;
	wire w_dff_B_wq6ka6iV3_1;
	wire w_dff_B_uAgzUDyg8_1;
	wire w_dff_B_AeRvJUhx5_1;
	wire w_dff_B_2CW2rMrE2_1;
	wire w_dff_B_5beuRPkf9_1;
	wire w_dff_B_U3TaZbq12_1;
	wire w_dff_B_7XCG2brg3_1;
	wire w_dff_B_2IDYKDSB4_1;
	wire w_dff_B_qv8EtgK93_1;
	wire w_dff_B_OInE0V554_1;
	wire w_dff_B_I4qmYqrl8_1;
	wire w_dff_B_FJ1p4NKB9_1;
	wire w_dff_B_yTzjFn1Z3_1;
	wire w_dff_B_SRSGRlyT9_1;
	wire w_dff_B_DSZxKQR17_1;
	wire w_dff_B_cErlBgLi0_1;
	wire w_dff_B_iAiTcOsN1_1;
	wire w_dff_B_UvuNRS5J0_1;
	wire w_dff_B_3Ojifvup9_1;
	wire w_dff_B_IN6YxyS01_1;
	wire w_dff_B_riZB7D8v0_1;
	wire w_dff_B_zSBr4CkT5_1;
	wire w_dff_B_w9foHQ6s1_1;
	wire w_dff_B_4LRWFXGT3_1;
	wire w_dff_B_O0b8v42C3_1;
	wire w_dff_B_bYfmDYht4_1;
	wire w_dff_B_5qgNxNOJ5_1;
	wire w_dff_B_L9jk8hv28_1;
	wire w_dff_B_bf80tCGe1_1;
	wire w_dff_B_CICJpYsg8_1;
	wire w_dff_B_aSlR0yiB8_1;
	wire w_dff_B_Ipg9G7pv1_1;
	wire w_dff_B_OkRAWWVb1_1;
	wire w_dff_B_WeMiE7JE1_1;
	wire w_dff_B_5BgT35oh5_1;
	wire w_dff_B_Oyu48oAj2_1;
	wire w_dff_B_uaEDwFjn2_1;
	wire w_dff_B_2RX2wqtp4_1;
	wire w_dff_B_DiaR3j2k7_1;
	wire w_dff_B_Yf4r0V2C1_1;
	wire w_dff_B_OdLRh7Za6_1;
	wire w_dff_B_y5N9hr4K5_1;
	wire w_dff_B_rkFLpgaS2_0;
	wire w_dff_B_S3LOZWvw8_0;
	wire w_dff_B_LoTvtAJc4_0;
	wire w_dff_B_d0CprS0L3_0;
	wire w_dff_B_buPdR9c42_0;
	wire w_dff_B_wDac1SNJ8_0;
	wire w_dff_B_JrZRhLJN3_0;
	wire w_dff_B_93tL2AYf2_0;
	wire w_dff_B_YhpaIu4D4_0;
	wire w_dff_B_q1a5rF7N6_0;
	wire w_dff_B_crQsYrUo4_0;
	wire w_dff_B_4VnZWyum0_0;
	wire w_dff_B_vlxWcSOz7_0;
	wire w_dff_B_sQ58d6Wc9_0;
	wire w_dff_B_KCxSDtfF1_0;
	wire w_dff_B_GkdOq5lE8_0;
	wire w_dff_B_N9cRcq5A6_0;
	wire w_dff_B_ivW5Zqpi7_0;
	wire w_dff_B_Mmm72eLt8_0;
	wire w_dff_B_cqGSFRGD7_0;
	wire w_dff_B_DT1w3ZyN0_0;
	wire w_dff_B_1UFxYQH18_0;
	wire w_dff_B_CuM2w5TT6_0;
	wire w_dff_B_nIyt3SmD3_0;
	wire w_dff_B_vq6JB6IU9_0;
	wire w_dff_B_Lbvj6yNV7_0;
	wire w_dff_B_dLcS5xX39_0;
	wire w_dff_B_I3EZLtz33_0;
	wire w_dff_B_69D6oSmW9_0;
	wire w_dff_B_9mL590f38_0;
	wire w_dff_B_oRwYY0Nh0_0;
	wire w_dff_B_Bn0kH5WL1_0;
	wire w_dff_B_hgQsWDyx3_0;
	wire w_dff_B_ReiD0qrT1_0;
	wire w_dff_B_al2HzM9O1_0;
	wire w_dff_B_SlrMrmXS7_0;
	wire w_dff_B_DCBYSJg66_0;
	wire w_dff_B_lUAmwcSL1_0;
	wire w_dff_B_Aug3b18x0_0;
	wire w_dff_B_Tny9fVpg8_0;
	wire w_dff_B_5AZs62he7_0;
	wire w_dff_B_ZzddWN548_0;
	wire w_dff_B_hy209J786_0;
	wire w_dff_B_XJ6b8ERc3_0;
	wire w_dff_B_hmXEDbDG4_1;
	wire w_dff_B_tAKMLcDx5_1;
	wire w_dff_B_qcy2NM5A9_1;
	wire w_dff_B_nvNvYJlT6_1;
	wire w_dff_B_OldzLEIo1_1;
	wire w_dff_B_rYqClixL7_1;
	wire w_dff_B_VwjJ68u28_1;
	wire w_dff_B_4kQ3BXYM6_1;
	wire w_dff_B_qZprjZLy9_1;
	wire w_dff_B_ZvKlv1NG2_1;
	wire w_dff_B_uPgYOZAa7_1;
	wire w_dff_B_PWeIYkio6_1;
	wire w_dff_B_evfM2W0p2_1;
	wire w_dff_B_XfqALNc12_1;
	wire w_dff_B_zomaaGNg7_1;
	wire w_dff_B_rwxtLz4s9_1;
	wire w_dff_B_5TDEQuhY7_1;
	wire w_dff_B_kZhyqGCq0_1;
	wire w_dff_B_hvCzCf3a9_1;
	wire w_dff_B_TKJIU4lu4_1;
	wire w_dff_B_DW4uxPVp3_1;
	wire w_dff_B_sc1hreCE8_1;
	wire w_dff_B_4Uyq7GMV3_1;
	wire w_dff_B_iAIZ3eEk3_1;
	wire w_dff_B_jpco5LcG1_1;
	wire w_dff_B_JLALGLXw4_1;
	wire w_dff_B_sNirE9If7_1;
	wire w_dff_B_45hiEaMW8_1;
	wire w_dff_B_OOFHBLuB8_1;
	wire w_dff_B_BBfyzCDk5_1;
	wire w_dff_B_EfMLlRon4_1;
	wire w_dff_B_GQ9mPjde4_1;
	wire w_dff_B_ncShczgI2_1;
	wire w_dff_B_eqgTEXam7_1;
	wire w_dff_B_ltCw1BIv3_1;
	wire w_dff_B_zl72ZCTT2_1;
	wire w_dff_B_vI4GBiwP8_1;
	wire w_dff_B_lqeuXDbv6_1;
	wire w_dff_B_QDNHosOz1_1;
	wire w_dff_B_94wIuLld1_1;
	wire w_dff_B_RY0SM2dq1_1;
	wire w_dff_B_INBVpObJ2_1;
	wire w_dff_B_OGZRqfWA9_1;
	wire w_dff_B_VVBVUF222_0;
	wire w_dff_B_dJiUKVNg4_0;
	wire w_dff_B_sxj8NmoB9_0;
	wire w_dff_B_4CuSmZZ12_0;
	wire w_dff_B_4eXe4Rzb2_0;
	wire w_dff_B_9qxlf1dl6_0;
	wire w_dff_B_qZOEJsS60_0;
	wire w_dff_B_7iZNVHLr6_0;
	wire w_dff_B_8HD9x4128_0;
	wire w_dff_B_e47r6vrl8_0;
	wire w_dff_B_uNUhQLKP7_0;
	wire w_dff_B_GqCWByrM3_0;
	wire w_dff_B_3mZkS0QV7_0;
	wire w_dff_B_rH3stAxW8_0;
	wire w_dff_B_eNzgpg0A5_0;
	wire w_dff_B_j8Sjl2VU8_0;
	wire w_dff_B_squWjeIf5_0;
	wire w_dff_B_Un8OMywj5_0;
	wire w_dff_B_nSBg6gC83_0;
	wire w_dff_B_HW9QDRPy6_0;
	wire w_dff_B_KW0rY31m7_0;
	wire w_dff_B_7xpzeyZY0_0;
	wire w_dff_B_5fY9Roe13_0;
	wire w_dff_B_EjbYz7756_0;
	wire w_dff_B_fA27xfmz5_0;
	wire w_dff_B_AFUcymdh8_0;
	wire w_dff_B_IyRtfTsA2_0;
	wire w_dff_B_zciLAZl70_0;
	wire w_dff_B_UTBQFDlX6_0;
	wire w_dff_B_YXvOjyel5_0;
	wire w_dff_B_Fcp0nyhg4_0;
	wire w_dff_B_i7pyVAgt8_0;
	wire w_dff_B_K2PKQ5uq7_0;
	wire w_dff_B_FoR2v05a5_0;
	wire w_dff_B_9SxyD6vQ9_0;
	wire w_dff_B_XafsW9UQ1_0;
	wire w_dff_B_BTAE8Es11_0;
	wire w_dff_B_yT7dIv8Q0_0;
	wire w_dff_B_OKsCZfTR4_0;
	wire w_dff_B_y7gRlNEB5_0;
	wire w_dff_B_5T8yzaqJ1_0;
	wire w_dff_B_ntLbGJVc0_0;
	wire w_dff_B_O1mNMYi88_0;
	wire w_dff_B_I7LqbT2f6_1;
	wire w_dff_B_wVR5WhD46_1;
	wire w_dff_B_D7PpRXsQ3_1;
	wire w_dff_B_KagA3vx81_1;
	wire w_dff_B_WS2gRnrE3_1;
	wire w_dff_B_diIbVVjn3_1;
	wire w_dff_B_vBFGn19E8_1;
	wire w_dff_B_s9J8fvom2_1;
	wire w_dff_B_GdFp3fIg8_1;
	wire w_dff_B_CLfn7nv39_1;
	wire w_dff_B_9LbufJdN7_1;
	wire w_dff_B_HXBPWuK24_1;
	wire w_dff_B_Y0L3hPQ42_1;
	wire w_dff_B_QwcrBjxJ0_1;
	wire w_dff_B_AYkb6pPK8_1;
	wire w_dff_B_UvpjWccQ2_1;
	wire w_dff_B_zfncn8f53_1;
	wire w_dff_B_EjYAWdsV3_1;
	wire w_dff_B_bNEs9cej4_1;
	wire w_dff_B_woE3QMSV8_1;
	wire w_dff_B_vGS18eus3_1;
	wire w_dff_B_BGuh95xX6_1;
	wire w_dff_B_SKbrTr5H8_1;
	wire w_dff_B_1dRHI08r1_1;
	wire w_dff_B_W4yY2TYG2_1;
	wire w_dff_B_2FBvsjGC4_1;
	wire w_dff_B_0eAzUOTC7_1;
	wire w_dff_B_mLwQ88MO4_1;
	wire w_dff_B_WeXoqRHL7_1;
	wire w_dff_B_5Ok4u67t8_1;
	wire w_dff_B_fd6fsVzN1_1;
	wire w_dff_B_ff2Mmcw55_1;
	wire w_dff_B_WHqckdFZ1_1;
	wire w_dff_B_A2aximwh1_1;
	wire w_dff_B_Y6BkQyQw2_1;
	wire w_dff_B_hFmPcJDa1_1;
	wire w_dff_B_Ii4Oanhf1_1;
	wire w_dff_B_CpGhp91t1_1;
	wire w_dff_B_2twUHnhx1_1;
	wire w_dff_B_zIWJSRtM2_1;
	wire w_dff_B_AkqcSZze2_1;
	wire w_dff_B_JMCouiXX8_1;
	wire w_dff_B_AcSz1DMq5_0;
	wire w_dff_B_PJePDGCS2_0;
	wire w_dff_B_NqHLJzGF9_0;
	wire w_dff_B_il8JkgqN6_0;
	wire w_dff_B_zQJPEKn48_0;
	wire w_dff_B_crfEaEZ47_0;
	wire w_dff_B_7zA5mFRp7_0;
	wire w_dff_B_n6y0sVy43_0;
	wire w_dff_B_KpbAV0gT4_0;
	wire w_dff_B_pkI9WEZY4_0;
	wire w_dff_B_0fdd2xVV6_0;
	wire w_dff_B_5LduqPRo9_0;
	wire w_dff_B_yPThiWtg6_0;
	wire w_dff_B_42s6Ek1s7_0;
	wire w_dff_B_jINLYooY0_0;
	wire w_dff_B_H9n2s8wP1_0;
	wire w_dff_B_zlMEz8vm0_0;
	wire w_dff_B_OcQJchxO8_0;
	wire w_dff_B_lXsVs8a26_0;
	wire w_dff_B_ufQptKRw5_0;
	wire w_dff_B_lfl0aAXB5_0;
	wire w_dff_B_O1QkvmHl2_0;
	wire w_dff_B_mFnNs4YD8_0;
	wire w_dff_B_A8Lo3swX6_0;
	wire w_dff_B_LE03pELK4_0;
	wire w_dff_B_Lb21lxX88_0;
	wire w_dff_B_1eUFobsA4_0;
	wire w_dff_B_5WtdonBp8_0;
	wire w_dff_B_vuYe2YEX1_0;
	wire w_dff_B_Io1QzfOL0_0;
	wire w_dff_B_Q32EF3Z83_0;
	wire w_dff_B_sS1Du8u40_0;
	wire w_dff_B_Ow6NRkMo4_0;
	wire w_dff_B_ew8IcJrQ3_0;
	wire w_dff_B_vgmPifxO3_0;
	wire w_dff_B_Cn1Ozxvh4_0;
	wire w_dff_B_lzsM3vLa5_0;
	wire w_dff_B_mWy09Jvh2_0;
	wire w_dff_B_e3BiTXmW2_0;
	wire w_dff_B_v9og7iuP2_0;
	wire w_dff_B_r5gEe0757_0;
	wire w_dff_B_Fe0B8YFI0_0;
	wire w_dff_B_LfvVBueY0_1;
	wire w_dff_B_NcKvCmdt5_1;
	wire w_dff_B_DJ6o65Lq3_1;
	wire w_dff_B_q0Psu5Uy0_1;
	wire w_dff_B_Je1FYDtC3_1;
	wire w_dff_B_iFxXbCNx8_1;
	wire w_dff_B_oC44ZmXv2_1;
	wire w_dff_B_uinjqs4z6_1;
	wire w_dff_B_pDoJZss74_1;
	wire w_dff_B_5SihKAo75_1;
	wire w_dff_B_JRksUubY9_1;
	wire w_dff_B_nJegQheD2_1;
	wire w_dff_B_h87hwmAm7_1;
	wire w_dff_B_DB7syB5h6_1;
	wire w_dff_B_QQxYH7d35_1;
	wire w_dff_B_gWGgSwGM6_1;
	wire w_dff_B_X5apSPjd9_1;
	wire w_dff_B_8gCECxur4_1;
	wire w_dff_B_6z21e0oO0_1;
	wire w_dff_B_jdSjGdEz7_1;
	wire w_dff_B_437FKpI84_1;
	wire w_dff_B_wA7ZMEcc7_1;
	wire w_dff_B_H7zLB2vL5_1;
	wire w_dff_B_ykok26La2_1;
	wire w_dff_B_EsPOWioc0_1;
	wire w_dff_B_Kq9F65Lt1_1;
	wire w_dff_B_MkO2miZq2_1;
	wire w_dff_B_TElzeroM0_1;
	wire w_dff_B_oQrqWhYX1_1;
	wire w_dff_B_iXFk4EJZ2_1;
	wire w_dff_B_O8NN1KSx5_1;
	wire w_dff_B_DM7PYOeZ4_1;
	wire w_dff_B_9jHn0Qrs3_1;
	wire w_dff_B_xh44CqbF7_1;
	wire w_dff_B_4ChyFnB71_1;
	wire w_dff_B_lqlvHr5s5_1;
	wire w_dff_B_aKvZTimR6_1;
	wire w_dff_B_UfLN8bv23_1;
	wire w_dff_B_rNYfaluK9_1;
	wire w_dff_B_daPY71Er5_1;
	wire w_dff_B_AyOrLbF03_1;
	wire w_dff_B_8QmPIgxg7_0;
	wire w_dff_B_gdpXlBXN8_0;
	wire w_dff_B_AugFBj339_0;
	wire w_dff_B_JC1E4JBT7_0;
	wire w_dff_B_ymUm0FtD5_0;
	wire w_dff_B_57KJpRgz0_0;
	wire w_dff_B_wtk4BUCI5_0;
	wire w_dff_B_UpULRIn27_0;
	wire w_dff_B_AmpsyZsk8_0;
	wire w_dff_B_tmnkAl681_0;
	wire w_dff_B_JoB70bx69_0;
	wire w_dff_B_hMab1QwY0_0;
	wire w_dff_B_4eDjRmk35_0;
	wire w_dff_B_iWtDPUc90_0;
	wire w_dff_B_qaMoqtoE5_0;
	wire w_dff_B_RaTFKHR32_0;
	wire w_dff_B_30aKGob80_0;
	wire w_dff_B_fErKBY4y9_0;
	wire w_dff_B_YzZSBsJV3_0;
	wire w_dff_B_m6Ympzvr4_0;
	wire w_dff_B_2oURZFRQ9_0;
	wire w_dff_B_RtKZtlBg9_0;
	wire w_dff_B_mj71ook10_0;
	wire w_dff_B_2mmi0acZ2_0;
	wire w_dff_B_bbiEC2Of8_0;
	wire w_dff_B_COsaEQCG9_0;
	wire w_dff_B_yFeoltQO1_0;
	wire w_dff_B_TCUhTIcm8_0;
	wire w_dff_B_o364N6ic5_0;
	wire w_dff_B_KWOueVoT5_0;
	wire w_dff_B_I8390tJR1_0;
	wire w_dff_B_kJwWrDQw3_0;
	wire w_dff_B_RHzLpNHa0_0;
	wire w_dff_B_bDxRWC8G9_0;
	wire w_dff_B_DvLBN5eN1_0;
	wire w_dff_B_D78bRx178_0;
	wire w_dff_B_6zdCY1st4_0;
	wire w_dff_B_jrGRcu648_0;
	wire w_dff_B_OjIGXFHP6_0;
	wire w_dff_B_LpJVmWzl0_0;
	wire w_dff_B_Vysb7cc73_0;
	wire w_dff_B_JtBXUdKo9_1;
	wire w_dff_B_tnuR8YWP5_1;
	wire w_dff_B_ylFQdDCL4_1;
	wire w_dff_B_FEWVQ50k5_1;
	wire w_dff_B_l6SyDGht7_1;
	wire w_dff_B_NJVX5EQd2_1;
	wire w_dff_B_Snv4rtsR1_1;
	wire w_dff_B_XGof5jkU7_1;
	wire w_dff_B_lX3DDY6P2_1;
	wire w_dff_B_xrqOj9PN6_1;
	wire w_dff_B_6ijP604D0_1;
	wire w_dff_B_DsvsmWQi6_1;
	wire w_dff_B_MNC9zpYz2_1;
	wire w_dff_B_Bny0fsYb5_1;
	wire w_dff_B_9e1uVB6s3_1;
	wire w_dff_B_loMNqfOv9_1;
	wire w_dff_B_Y1r64aQ38_1;
	wire w_dff_B_9qjEfqHL5_1;
	wire w_dff_B_1mpgSUft4_1;
	wire w_dff_B_eZTibyd20_1;
	wire w_dff_B_vnDv5Lrd5_1;
	wire w_dff_B_XJpXZniX4_1;
	wire w_dff_B_j8My0uqp8_1;
	wire w_dff_B_CKDDbEDM3_1;
	wire w_dff_B_YZortXJx0_1;
	wire w_dff_B_PZV5GHdW1_1;
	wire w_dff_B_J6hPIZzi6_1;
	wire w_dff_B_QuZ4fmUX1_1;
	wire w_dff_B_nbjg4KOP4_1;
	wire w_dff_B_LH6xMYq93_1;
	wire w_dff_B_7kXgOwiy2_1;
	wire w_dff_B_gocHhJhU6_1;
	wire w_dff_B_4RytfaR86_1;
	wire w_dff_B_wRNdkMcH9_1;
	wire w_dff_B_0GN34qzU1_1;
	wire w_dff_B_LaLGX4Cn7_1;
	wire w_dff_B_Ihdgu3SC3_1;
	wire w_dff_B_NcT0vIXU4_1;
	wire w_dff_B_2FaxzmXI9_1;
	wire w_dff_B_snRizMBV3_1;
	wire w_dff_B_o8mfxGyU6_0;
	wire w_dff_B_PUPElYb84_0;
	wire w_dff_B_dLpcJHua6_0;
	wire w_dff_B_TkbtOCnL5_0;
	wire w_dff_B_fDi3aK9J6_0;
	wire w_dff_B_Ul0Z20f02_0;
	wire w_dff_B_1sqn5kY48_0;
	wire w_dff_B_zTtg9Q927_0;
	wire w_dff_B_AqwG4Rta1_0;
	wire w_dff_B_poKcUpzJ3_0;
	wire w_dff_B_X6h0VplD7_0;
	wire w_dff_B_RNKjgaXI1_0;
	wire w_dff_B_oQRgSYB33_0;
	wire w_dff_B_rm1TJM0X5_0;
	wire w_dff_B_wKmXwpRf0_0;
	wire w_dff_B_iXGhHx0F6_0;
	wire w_dff_B_I4H8JLQ83_0;
	wire w_dff_B_xdM7t0hJ0_0;
	wire w_dff_B_G7AG8Hem0_0;
	wire w_dff_B_RWt0LnXB7_0;
	wire w_dff_B_U1BaAeiV1_0;
	wire w_dff_B_TAUiwysf0_0;
	wire w_dff_B_m61JRhu45_0;
	wire w_dff_B_D0X3Pn096_0;
	wire w_dff_B_QdgAXuHb7_0;
	wire w_dff_B_TMJA1A3w8_0;
	wire w_dff_B_XhNtbCfn9_0;
	wire w_dff_B_4zRtAuoH9_0;
	wire w_dff_B_dAH1Q7QK9_0;
	wire w_dff_B_19RreQQs1_0;
	wire w_dff_B_94366zT98_0;
	wire w_dff_B_juOMJ1AY3_0;
	wire w_dff_B_aA85Jycj4_0;
	wire w_dff_B_5fCnl3QD9_0;
	wire w_dff_B_qXgoHIwS3_0;
	wire w_dff_B_nBYX7AaE3_0;
	wire w_dff_B_7BmlLgs43_0;
	wire w_dff_B_pBBtc8UM7_0;
	wire w_dff_B_6O2Govit3_0;
	wire w_dff_B_v6JmAK7j4_0;
	wire w_dff_B_xzNs3A4M6_1;
	wire w_dff_B_s01y1Wtc1_1;
	wire w_dff_B_wCtWxCcz4_1;
	wire w_dff_B_8yP6upqU5_1;
	wire w_dff_B_C5GJfc6h0_1;
	wire w_dff_B_8tpjvD302_1;
	wire w_dff_B_qaTYaa3Z7_1;
	wire w_dff_B_6DXjRWWV4_1;
	wire w_dff_B_7yuGZxwu6_1;
	wire w_dff_B_irM2ab3R0_1;
	wire w_dff_B_psde5juB8_1;
	wire w_dff_B_O2O1igCC1_1;
	wire w_dff_B_HJPnBiZm2_1;
	wire w_dff_B_LQo44HpF2_1;
	wire w_dff_B_n7IBoHt73_1;
	wire w_dff_B_Nb6mRhav0_1;
	wire w_dff_B_iVfYt3Xp8_1;
	wire w_dff_B_x1f5z0VI7_1;
	wire w_dff_B_51nqEt9r5_1;
	wire w_dff_B_HChZ5S6X1_1;
	wire w_dff_B_KKocAJDS9_1;
	wire w_dff_B_xANEwfpg5_1;
	wire w_dff_B_N9aBp7x86_1;
	wire w_dff_B_rjpQ0Vrr7_1;
	wire w_dff_B_eVLvNr9U2_1;
	wire w_dff_B_wzZLjjXc3_1;
	wire w_dff_B_LCB8nkvn4_1;
	wire w_dff_B_IaVkYITB1_1;
	wire w_dff_B_TJtf2OrS3_1;
	wire w_dff_B_4shiWAZO0_1;
	wire w_dff_B_TX61vdvN2_1;
	wire w_dff_B_NEYiPyj59_1;
	wire w_dff_B_wCBlSHfj3_1;
	wire w_dff_B_gp754SI74_1;
	wire w_dff_B_5KZNcjZo2_1;
	wire w_dff_B_ojL8Y5TK5_1;
	wire w_dff_B_URhAnzRc0_1;
	wire w_dff_B_84Hiap2m8_1;
	wire w_dff_B_1cZChDiV8_1;
	wire w_dff_B_i5VTpo2H0_0;
	wire w_dff_B_RQmDHBCp0_0;
	wire w_dff_B_rvxlBOtD2_0;
	wire w_dff_B_yqNj9LDA3_0;
	wire w_dff_B_RIATV5hH1_0;
	wire w_dff_B_jMsOL3vp7_0;
	wire w_dff_B_r9zowARR0_0;
	wire w_dff_B_Zg4iFbBX0_0;
	wire w_dff_B_lCXmiMOp9_0;
	wire w_dff_B_g4UFrxPP1_0;
	wire w_dff_B_jFPiEOD57_0;
	wire w_dff_B_QMMJIS8c6_0;
	wire w_dff_B_4lmsmhQq7_0;
	wire w_dff_B_bCrYGWew7_0;
	wire w_dff_B_GK3lBu273_0;
	wire w_dff_B_Bgr8ryv43_0;
	wire w_dff_B_0ltDi3rS8_0;
	wire w_dff_B_bedNWeIh6_0;
	wire w_dff_B_CZhY63wi9_0;
	wire w_dff_B_6AxVyPtV2_0;
	wire w_dff_B_o4vlHLg51_0;
	wire w_dff_B_ejQ3axLP1_0;
	wire w_dff_B_pj9IPYEV4_0;
	wire w_dff_B_YC3DZGqd5_0;
	wire w_dff_B_p7v87gs65_0;
	wire w_dff_B_Q1FbSoin3_0;
	wire w_dff_B_Isxlw9op1_0;
	wire w_dff_B_GEdcbSpu6_0;
	wire w_dff_B_9UGnkm8S6_0;
	wire w_dff_B_ul4Emnel7_0;
	wire w_dff_B_mReWuBRi7_0;
	wire w_dff_B_80BJIkHo9_0;
	wire w_dff_B_qhgaY1TM3_0;
	wire w_dff_B_h0ypPEU98_0;
	wire w_dff_B_4waKMxF29_0;
	wire w_dff_B_TAYMfE5T9_0;
	wire w_dff_B_CwvfHwiR1_0;
	wire w_dff_B_l4zQADy20_0;
	wire w_dff_B_GoygnPeZ7_0;
	wire w_dff_B_iOAW5AkF8_1;
	wire w_dff_B_9L0ukpX21_1;
	wire w_dff_B_bwvSSOEo8_1;
	wire w_dff_B_ROFAGxLi7_1;
	wire w_dff_B_jT6Ym0JL5_1;
	wire w_dff_B_SqxwqfOG2_1;
	wire w_dff_B_cLvbRdyC2_1;
	wire w_dff_B_7bK7jhrl1_1;
	wire w_dff_B_ckTpkfs12_1;
	wire w_dff_B_Pb7DM3cE3_1;
	wire w_dff_B_3g2H9eTP3_1;
	wire w_dff_B_coVYVmSq1_1;
	wire w_dff_B_6odMHASB8_1;
	wire w_dff_B_VFhPuvlR3_1;
	wire w_dff_B_u2oY7gAH2_1;
	wire w_dff_B_eNekqtlL6_1;
	wire w_dff_B_0vTuaUAb2_1;
	wire w_dff_B_bC4I7ru02_1;
	wire w_dff_B_5uaozvxf7_1;
	wire w_dff_B_cZmWyixe1_1;
	wire w_dff_B_2Mq98epl1_1;
	wire w_dff_B_DVyKpPt54_1;
	wire w_dff_B_Ug8Xamma4_1;
	wire w_dff_B_zWjkUzMy5_1;
	wire w_dff_B_LTJcstDk5_1;
	wire w_dff_B_3tjs6x592_1;
	wire w_dff_B_ONjHRyg59_1;
	wire w_dff_B_9PreDRWH4_1;
	wire w_dff_B_xPSeyFCx0_1;
	wire w_dff_B_xdN6Hr634_1;
	wire w_dff_B_wNfL7A9v3_1;
	wire w_dff_B_l18RPvVU6_1;
	wire w_dff_B_TO7PzIaj3_1;
	wire w_dff_B_bipiOQLK9_1;
	wire w_dff_B_3s3EH4Fk3_1;
	wire w_dff_B_cycLBPrn5_1;
	wire w_dff_B_NHJKcyqZ4_1;
	wire w_dff_B_u1eB0U854_1;
	wire w_dff_B_Z8jCkfZY6_0;
	wire w_dff_B_Bt7Owyjw5_0;
	wire w_dff_B_TlvrmO933_0;
	wire w_dff_B_LgIM5swc7_0;
	wire w_dff_B_Cqf05TVk4_0;
	wire w_dff_B_hD6wqKc17_0;
	wire w_dff_B_aRhaC4cG6_0;
	wire w_dff_B_3nAD1CKi8_0;
	wire w_dff_B_QOAJRXMM4_0;
	wire w_dff_B_76qjEiyE8_0;
	wire w_dff_B_HRdRkrcI1_0;
	wire w_dff_B_yhZHwnXK9_0;
	wire w_dff_B_B8um4RKu0_0;
	wire w_dff_B_MBAOr4b09_0;
	wire w_dff_B_et7e8b3V1_0;
	wire w_dff_B_L0nYeOLq4_0;
	wire w_dff_B_IqrIqAQr5_0;
	wire w_dff_B_UV6KRfwW4_0;
	wire w_dff_B_tFgU9Iza0_0;
	wire w_dff_B_L3DnhOEG3_0;
	wire w_dff_B_UsxwXYhk4_0;
	wire w_dff_B_zCxnUZ4G7_0;
	wire w_dff_B_l5QxuTNN1_0;
	wire w_dff_B_j8HtY50C2_0;
	wire w_dff_B_A1hVmr8q2_0;
	wire w_dff_B_b3bUlmRR2_0;
	wire w_dff_B_G1iaj4CP7_0;
	wire w_dff_B_8KVtQ9Jx0_0;
	wire w_dff_B_zVaeqir66_0;
	wire w_dff_B_X2EG9XJK3_0;
	wire w_dff_B_LD9DlGyG4_0;
	wire w_dff_B_wRbo9ZCb1_0;
	wire w_dff_B_I2GqYFZV5_0;
	wire w_dff_B_20nn7j327_0;
	wire w_dff_B_m4ydpTvG5_0;
	wire w_dff_B_4f0BJZaz9_0;
	wire w_dff_B_ccXyxJ5S1_0;
	wire w_dff_B_wdau1vMx1_0;
	wire w_dff_B_f4hct7133_1;
	wire w_dff_B_UXIyiguw6_1;
	wire w_dff_B_ozl04Lbd5_1;
	wire w_dff_B_JJnQpDCe3_1;
	wire w_dff_B_20Iin53p2_1;
	wire w_dff_B_CPAQ9Htg8_1;
	wire w_dff_B_bXOSEEV56_1;
	wire w_dff_B_mH2SAvxU1_1;
	wire w_dff_B_MixDna5N6_1;
	wire w_dff_B_t8szfHZc6_1;
	wire w_dff_B_lDBahBDa5_1;
	wire w_dff_B_Qc5i2W7l6_1;
	wire w_dff_B_jlMKZlRA4_1;
	wire w_dff_B_HsOv0bM55_1;
	wire w_dff_B_hcChzzT21_1;
	wire w_dff_B_jOZWmHiB3_1;
	wire w_dff_B_6W51sSxp6_1;
	wire w_dff_B_yVQvIEVZ7_1;
	wire w_dff_B_ctGeb99d9_1;
	wire w_dff_B_eUTnZ67z0_1;
	wire w_dff_B_EEHIYTbk5_1;
	wire w_dff_B_jLjqArVF7_1;
	wire w_dff_B_ycN4tM0G0_1;
	wire w_dff_B_65HPNs7T0_1;
	wire w_dff_B_2jEWg2ys7_1;
	wire w_dff_B_ljjvTOLC3_1;
	wire w_dff_B_v3B2YGPr4_1;
	wire w_dff_B_IQ7KbHQ30_1;
	wire w_dff_B_ihQOhxU36_1;
	wire w_dff_B_U1veCSAc6_1;
	wire w_dff_B_X53RkT039_1;
	wire w_dff_B_MRkHPJkR3_1;
	wire w_dff_B_uxWcVFyM7_1;
	wire w_dff_B_pskpqPuo7_1;
	wire w_dff_B_R3I60Yzp2_1;
	wire w_dff_B_5fIXPGLI4_1;
	wire w_dff_B_S6RAvCjq6_1;
	wire w_dff_B_DmHFh1vJ1_0;
	wire w_dff_B_VqROpL253_0;
	wire w_dff_B_jIHgcl5h1_0;
	wire w_dff_B_Sgdhq7o45_0;
	wire w_dff_B_ilIt7LCa6_0;
	wire w_dff_B_R0DJgRiQ3_0;
	wire w_dff_B_5R8mmLHp8_0;
	wire w_dff_B_CguuiksR8_0;
	wire w_dff_B_FGXbcDCf4_0;
	wire w_dff_B_OqgE3CEy2_0;
	wire w_dff_B_ns4710rp3_0;
	wire w_dff_B_dyeMjlIy7_0;
	wire w_dff_B_CFUDoG6Z3_0;
	wire w_dff_B_B0sOZkZM6_0;
	wire w_dff_B_5gcYsIoH5_0;
	wire w_dff_B_xiOR2scU6_0;
	wire w_dff_B_BzsR9TK23_0;
	wire w_dff_B_bhrvY4bm6_0;
	wire w_dff_B_REKnead37_0;
	wire w_dff_B_1mNAH0Ly8_0;
	wire w_dff_B_Auq973zI4_0;
	wire w_dff_B_h3Z9Bh2Q6_0;
	wire w_dff_B_ilqOOL8z3_0;
	wire w_dff_B_J1VZ0xkc1_0;
	wire w_dff_B_9DyUJqlf7_0;
	wire w_dff_B_Otk4fYEB1_0;
	wire w_dff_B_dr9GPM9O7_0;
	wire w_dff_B_gskPMh415_0;
	wire w_dff_B_BzhcQmsX5_0;
	wire w_dff_B_tT4ya5nE6_0;
	wire w_dff_B_5Vz0mAoU0_0;
	wire w_dff_B_BGDhAFpM9_0;
	wire w_dff_B_YfzPuViz1_0;
	wire w_dff_B_ZEuUTuhN9_0;
	wire w_dff_B_xR5NWHE36_0;
	wire w_dff_B_LviJle7c6_0;
	wire w_dff_B_vt7Bt9w49_0;
	wire w_dff_B_h5xdW6Ka7_1;
	wire w_dff_B_sMzxXgdl5_1;
	wire w_dff_B_icuzylNk4_1;
	wire w_dff_B_52MpWRoQ2_1;
	wire w_dff_B_tt2ib7Qh9_1;
	wire w_dff_B_UPDmu91F1_1;
	wire w_dff_B_HcO25vxE5_1;
	wire w_dff_B_jpD1P5a48_1;
	wire w_dff_B_qfrnzzyn2_1;
	wire w_dff_B_MxZOwriT5_1;
	wire w_dff_B_Hu6DelX76_1;
	wire w_dff_B_hQHzplWL8_1;
	wire w_dff_B_D4IoxlfC7_1;
	wire w_dff_B_gFuvVzQ31_1;
	wire w_dff_B_7X2EEtLC2_1;
	wire w_dff_B_0cN8V0ev7_1;
	wire w_dff_B_kNX0wAeJ9_1;
	wire w_dff_B_sWp3WGKN7_1;
	wire w_dff_B_kKOGdNK46_1;
	wire w_dff_B_KYBZSZZK0_1;
	wire w_dff_B_VtTivnjq1_1;
	wire w_dff_B_caDg5JJH9_1;
	wire w_dff_B_el37d9oH3_1;
	wire w_dff_B_94qDdOOI4_1;
	wire w_dff_B_bxI4QB295_1;
	wire w_dff_B_lMWKw1qL3_1;
	wire w_dff_B_lpHH3xJE8_1;
	wire w_dff_B_xcIt5GSE5_1;
	wire w_dff_B_juPcgAlV9_1;
	wire w_dff_B_p3GPETM53_1;
	wire w_dff_B_z0YRF4gu7_1;
	wire w_dff_B_GX55SWVr3_1;
	wire w_dff_B_pIXeCOyP1_1;
	wire w_dff_B_ltcYCDCy1_1;
	wire w_dff_B_t23r44QK3_1;
	wire w_dff_B_ntOAyf159_1;
	wire w_dff_B_BA3uUTcD5_0;
	wire w_dff_B_IY37tbG36_0;
	wire w_dff_B_rX8QeA4w1_0;
	wire w_dff_B_UunReUbN6_0;
	wire w_dff_B_GO1xSD9R9_0;
	wire w_dff_B_QdCBvY8M0_0;
	wire w_dff_B_WYNtXSG78_0;
	wire w_dff_B_vw1qRB0Y3_0;
	wire w_dff_B_21VJfEaJ9_0;
	wire w_dff_B_cMFwrMor9_0;
	wire w_dff_B_HypVbknO8_0;
	wire w_dff_B_U6v6e7Ma9_0;
	wire w_dff_B_7JABikK63_0;
	wire w_dff_B_Wcy97j6v0_0;
	wire w_dff_B_wAZV1ICG5_0;
	wire w_dff_B_RnExXpTC8_0;
	wire w_dff_B_M6EWYHAY4_0;
	wire w_dff_B_ztlmdiCI5_0;
	wire w_dff_B_gOvI0Pqc2_0;
	wire w_dff_B_BedvMGyv6_0;
	wire w_dff_B_12UjqWxY1_0;
	wire w_dff_B_Hr36akQr9_0;
	wire w_dff_B_9E4UyoDN3_0;
	wire w_dff_B_KU25avqa7_0;
	wire w_dff_B_BvqJYc5o9_0;
	wire w_dff_B_g3pE7bqQ3_0;
	wire w_dff_B_bjj7b4G76_0;
	wire w_dff_B_ts6zT4X01_0;
	wire w_dff_B_1WI8exoW7_0;
	wire w_dff_B_dQzew06Y4_0;
	wire w_dff_B_s5s1FNvm2_0;
	wire w_dff_B_LTklb7IV9_0;
	wire w_dff_B_3OBW9knB7_0;
	wire w_dff_B_ksPxZ7WT3_0;
	wire w_dff_B_T2Fc7qLA3_0;
	wire w_dff_B_Giv88Gjw1_0;
	wire w_dff_B_RFleY3cT7_1;
	wire w_dff_B_o0SdHfrv0_1;
	wire w_dff_B_PKCgycnV4_1;
	wire w_dff_B_n7CGMQ451_1;
	wire w_dff_B_aaMGmXGc4_1;
	wire w_dff_B_n3t1iiLE1_1;
	wire w_dff_B_zoIudX5I5_1;
	wire w_dff_B_0uGNVUpk4_1;
	wire w_dff_B_N5OF68FT9_1;
	wire w_dff_B_oxLipQWa5_1;
	wire w_dff_B_d3Tt3NNn6_1;
	wire w_dff_B_gLIVBpqf8_1;
	wire w_dff_B_gLSRRrlu8_1;
	wire w_dff_B_DCCReXPn7_1;
	wire w_dff_B_RhH8y4yo4_1;
	wire w_dff_B_5kKUMZGE4_1;
	wire w_dff_B_Vy6giZbs8_1;
	wire w_dff_B_4HeTjNQa2_1;
	wire w_dff_B_jHqlPfIE7_1;
	wire w_dff_B_m88H5LkI7_1;
	wire w_dff_B_NxU417Uu9_1;
	wire w_dff_B_K7fU8ITe9_1;
	wire w_dff_B_QG2BfaTf6_1;
	wire w_dff_B_5V6RjaT84_1;
	wire w_dff_B_wI1eJqcb0_1;
	wire w_dff_B_ZPIO6g0O6_1;
	wire w_dff_B_6hHLCboa5_1;
	wire w_dff_B_8UPRRRSB7_1;
	wire w_dff_B_QkHjKDoB8_1;
	wire w_dff_B_4kZcQGWj4_1;
	wire w_dff_B_s8fbOKAE3_1;
	wire w_dff_B_TtdLCU858_1;
	wire w_dff_B_VY1D2qEV5_1;
	wire w_dff_B_9XkkEIKa9_1;
	wire w_dff_B_PbcuSyj41_1;
	wire w_dff_B_Rqvx2lkt1_0;
	wire w_dff_B_MUXDV8y82_0;
	wire w_dff_B_Hib5v7zF8_0;
	wire w_dff_B_36deffBk1_0;
	wire w_dff_B_Z4trfWgg6_0;
	wire w_dff_B_w1i2sHnu1_0;
	wire w_dff_B_xJyfTY1R9_0;
	wire w_dff_B_nkW5Mc1L2_0;
	wire w_dff_B_hr540QWz5_0;
	wire w_dff_B_s5CVi2OT9_0;
	wire w_dff_B_Zrlwuc2h1_0;
	wire w_dff_B_lk1kZ6Oj4_0;
	wire w_dff_B_IoEansJ12_0;
	wire w_dff_B_vKcd36FX3_0;
	wire w_dff_B_yPl8uL8o9_0;
	wire w_dff_B_dxNMwbHM4_0;
	wire w_dff_B_1Bp3UrTf9_0;
	wire w_dff_B_bdrTM9D63_0;
	wire w_dff_B_S2GLdNs63_0;
	wire w_dff_B_UogI0Y4z9_0;
	wire w_dff_B_ZGwpUHiZ3_0;
	wire w_dff_B_AW74jYXA5_0;
	wire w_dff_B_G1gWiONj5_0;
	wire w_dff_B_otHs145F4_0;
	wire w_dff_B_J6HEMNNZ1_0;
	wire w_dff_B_nzuQA4Fm8_0;
	wire w_dff_B_qK5Sdcws0_0;
	wire w_dff_B_3OTtlZsH6_0;
	wire w_dff_B_U8xbl7qB7_0;
	wire w_dff_B_rwAlfQEC1_0;
	wire w_dff_B_WD8zd9KI8_0;
	wire w_dff_B_tgrF5Hzc9_0;
	wire w_dff_B_NBNeCR8Y4_0;
	wire w_dff_B_UgeCLmEn2_0;
	wire w_dff_B_N2n8UqAM7_0;
	wire w_dff_B_02b2xEfn2_1;
	wire w_dff_B_gkzTkmCx1_1;
	wire w_dff_B_jRWgKmn68_1;
	wire w_dff_B_plYVua4g6_1;
	wire w_dff_B_tjH0DXuC6_1;
	wire w_dff_B_Ipjlbscu2_1;
	wire w_dff_B_50Lqqz3j7_1;
	wire w_dff_B_oeLEYTe21_1;
	wire w_dff_B_oomihasE2_1;
	wire w_dff_B_Una2FvI36_1;
	wire w_dff_B_xASc30645_1;
	wire w_dff_B_ZSFXmSrz0_1;
	wire w_dff_B_Klg170KV7_1;
	wire w_dff_B_926dC0rJ0_1;
	wire w_dff_B_FjgoKXaQ8_1;
	wire w_dff_B_FIntbdhJ6_1;
	wire w_dff_B_RjS4d5lB5_1;
	wire w_dff_B_1Ct1ObmX7_1;
	wire w_dff_B_RnbTfalx4_1;
	wire w_dff_B_BbDgaJkA2_1;
	wire w_dff_B_A4O1rxU15_1;
	wire w_dff_B_yYNvWGU08_1;
	wire w_dff_B_KuIDJd9f3_1;
	wire w_dff_B_TdjAzBHD0_1;
	wire w_dff_B_CoN9U1CR8_1;
	wire w_dff_B_R2j7WGDG4_1;
	wire w_dff_B_A74IMyT57_1;
	wire w_dff_B_Ky1Ma0gz9_1;
	wire w_dff_B_IUzz9bHI1_1;
	wire w_dff_B_LLMWUEpr8_1;
	wire w_dff_B_bWlS1lQp9_1;
	wire w_dff_B_faX2aisv2_1;
	wire w_dff_B_RvlOhSxn9_1;
	wire w_dff_B_xBRXkssz2_1;
	wire w_dff_B_jPjE4w566_0;
	wire w_dff_B_Ri33JLN58_0;
	wire w_dff_B_qzVPKuyH0_0;
	wire w_dff_B_Z9Wml6E79_0;
	wire w_dff_B_DpwaP6ej4_0;
	wire w_dff_B_FO1BGuR42_0;
	wire w_dff_B_CGZ7jiuy1_0;
	wire w_dff_B_Zzm804cc2_0;
	wire w_dff_B_PQ69IjpM0_0;
	wire w_dff_B_DNhqEuWv9_0;
	wire w_dff_B_ZLY8E1Ar3_0;
	wire w_dff_B_AbBPNhSW3_0;
	wire w_dff_B_g4mkXwWN6_0;
	wire w_dff_B_aAQAtjIZ1_0;
	wire w_dff_B_lAOr0Neg3_0;
	wire w_dff_B_PxYGi3lK2_0;
	wire w_dff_B_m9edO10P9_0;
	wire w_dff_B_8m53RdS99_0;
	wire w_dff_B_OqzuyDLw2_0;
	wire w_dff_B_87Cmlgxq5_0;
	wire w_dff_B_KwyDwHQw0_0;
	wire w_dff_B_Advn2Nhl0_0;
	wire w_dff_B_r1lyi1PS9_0;
	wire w_dff_B_sTmFQkDr7_0;
	wire w_dff_B_r2VTro4A7_0;
	wire w_dff_B_YavBotb38_0;
	wire w_dff_B_J4vcTPkf5_0;
	wire w_dff_B_CiejrLnL6_0;
	wire w_dff_B_s0ABvs464_0;
	wire w_dff_B_IXBbbxc29_0;
	wire w_dff_B_aHx5w51h0_0;
	wire w_dff_B_mEZxTeOo9_0;
	wire w_dff_B_iI1rlTwq7_0;
	wire w_dff_B_NuWicBqk2_0;
	wire w_dff_B_02Ap5I3I2_1;
	wire w_dff_B_KMkF11mo1_1;
	wire w_dff_B_wFI2wHrj4_1;
	wire w_dff_B_l9DDrO862_1;
	wire w_dff_B_80uY3sSQ4_1;
	wire w_dff_B_zWWTpkUM0_1;
	wire w_dff_B_4hoZaLfJ4_1;
	wire w_dff_B_64h7T9QD7_1;
	wire w_dff_B_6ZBuhXOA6_1;
	wire w_dff_B_M2iBSq8J2_1;
	wire w_dff_B_Eujl7wjc8_1;
	wire w_dff_B_i60bOPkj2_1;
	wire w_dff_B_F6HgQXgX6_1;
	wire w_dff_B_wFnbaeXT9_1;
	wire w_dff_B_QfdSnFPW9_1;
	wire w_dff_B_UdEM3CIt5_1;
	wire w_dff_B_N8lCJAP71_1;
	wire w_dff_B_9KpUejbz4_1;
	wire w_dff_B_u6uv26L64_1;
	wire w_dff_B_gwihwOcj1_1;
	wire w_dff_B_12ndL5kl2_1;
	wire w_dff_B_w7LtAWwv4_1;
	wire w_dff_B_8DU8tLtq3_1;
	wire w_dff_B_ZQQIIxgW6_1;
	wire w_dff_B_rHDfCPm65_1;
	wire w_dff_B_BLOZd5o33_1;
	wire w_dff_B_ybr6fgZm2_1;
	wire w_dff_B_JfQCiZAS3_1;
	wire w_dff_B_vD1Xj51c1_1;
	wire w_dff_B_zqSHb1R55_1;
	wire w_dff_B_zlZ0WpMP4_1;
	wire w_dff_B_anBghBRu9_1;
	wire w_dff_B_D2kiPHXL3_1;
	wire w_dff_B_7RJiBTay1_0;
	wire w_dff_B_VpafdGyq6_0;
	wire w_dff_B_LOxNFQMu9_0;
	wire w_dff_B_xdQIF0Ce8_0;
	wire w_dff_B_JhyBeqdV9_0;
	wire w_dff_B_ypxhoOHo6_0;
	wire w_dff_B_RtYdGEuc6_0;
	wire w_dff_B_kCbcZnUt0_0;
	wire w_dff_B_JmmLgQQy9_0;
	wire w_dff_B_bud2Cav66_0;
	wire w_dff_B_Qacz87Np6_0;
	wire w_dff_B_roIrZ3r95_0;
	wire w_dff_B_INQJCmsq4_0;
	wire w_dff_B_S2YUjpry2_0;
	wire w_dff_B_hQvhKyRF0_0;
	wire w_dff_B_gBAv87676_0;
	wire w_dff_B_eMJv1uhA0_0;
	wire w_dff_B_pbKGzT0D2_0;
	wire w_dff_B_xy3halQ76_0;
	wire w_dff_B_R019oiuF3_0;
	wire w_dff_B_Esw8TCrc8_0;
	wire w_dff_B_wU4KaYnM5_0;
	wire w_dff_B_Gmqk0wQw5_0;
	wire w_dff_B_38OZjszQ5_0;
	wire w_dff_B_QLzSVlP16_0;
	wire w_dff_B_YnqMNmTs9_0;
	wire w_dff_B_rJLGgzlb4_0;
	wire w_dff_B_SmFLyRQE5_0;
	wire w_dff_B_Lqoqfaep2_0;
	wire w_dff_B_Nqo52NhK6_0;
	wire w_dff_B_4FBdH4nN3_0;
	wire w_dff_B_HZFIiVPS6_0;
	wire w_dff_B_76wrGEuj0_0;
	wire w_dff_B_tcHJDcFR1_1;
	wire w_dff_B_9WZlktg52_1;
	wire w_dff_B_70J7M71a6_1;
	wire w_dff_B_0bNe4Y0s1_1;
	wire w_dff_B_nL0y6gwC7_1;
	wire w_dff_B_oLYZUBoU8_1;
	wire w_dff_B_8e33wE607_1;
	wire w_dff_B_cwZcdbUu5_1;
	wire w_dff_B_AZBe0AUB8_1;
	wire w_dff_B_Q8rdd7TP9_1;
	wire w_dff_B_ihvEdK217_1;
	wire w_dff_B_HKvyjCvR1_1;
	wire w_dff_B_AHs9aKfS6_1;
	wire w_dff_B_cL4iQgTA6_1;
	wire w_dff_B_bBfx54BQ6_1;
	wire w_dff_B_K7JRSSOa8_1;
	wire w_dff_B_Y4PA8f7k0_1;
	wire w_dff_B_UrbgIzAO2_1;
	wire w_dff_B_z7F38Wm55_1;
	wire w_dff_B_M7kYfyXx9_1;
	wire w_dff_B_3tsAD5WQ5_1;
	wire w_dff_B_vt5r96si8_1;
	wire w_dff_B_vo4VCx545_1;
	wire w_dff_B_6boj367I4_1;
	wire w_dff_B_9lkMKfrF3_1;
	wire w_dff_B_qCwmP2Bx2_1;
	wire w_dff_B_SnPkuC3J6_1;
	wire w_dff_B_nJDSxQzd6_1;
	wire w_dff_B_M8fpqb9M1_1;
	wire w_dff_B_r7PLsI4y8_1;
	wire w_dff_B_ObSE17NU7_1;
	wire w_dff_B_vpzfAeXc3_1;
	wire w_dff_B_LTNSCy3T5_0;
	wire w_dff_B_Kq8KMKH56_0;
	wire w_dff_B_j5jfyqWt5_0;
	wire w_dff_B_oZlHD0Yl6_0;
	wire w_dff_B_HepHhI2P1_0;
	wire w_dff_B_8Efjhcm60_0;
	wire w_dff_B_ONwbUvE51_0;
	wire w_dff_B_VPLQHarR4_0;
	wire w_dff_B_lYpDM30S8_0;
	wire w_dff_B_gkWjX6SZ2_0;
	wire w_dff_B_xHe8vVaJ7_0;
	wire w_dff_B_yMdjtUHY0_0;
	wire w_dff_B_NJJYcFd94_0;
	wire w_dff_B_JYBt8lY52_0;
	wire w_dff_B_rjhanWVQ0_0;
	wire w_dff_B_N8FOrpxZ3_0;
	wire w_dff_B_1qRgo3sm0_0;
	wire w_dff_B_ZehycAL99_0;
	wire w_dff_B_F8h5tk9C4_0;
	wire w_dff_B_xxiTipoX3_0;
	wire w_dff_B_Z51J2Y152_0;
	wire w_dff_B_FSbsuUJ49_0;
	wire w_dff_B_c2Ni1VaX3_0;
	wire w_dff_B_hJYS97bM5_0;
	wire w_dff_B_uZPAnIg84_0;
	wire w_dff_B_rxbIYFOS9_0;
	wire w_dff_B_pjsjn3Lx1_0;
	wire w_dff_B_AXIT0TSo2_0;
	wire w_dff_B_MJXNOGvL3_0;
	wire w_dff_B_LtvlIL626_0;
	wire w_dff_B_SOMmHbp60_0;
	wire w_dff_B_cOSHsCTW4_0;
	wire w_dff_B_samYFRy26_1;
	wire w_dff_B_v8zPcZTW1_1;
	wire w_dff_B_ckoCJW2f2_1;
	wire w_dff_B_UGRsZrVB2_1;
	wire w_dff_B_Z7KUzV076_1;
	wire w_dff_B_7ie9hnnY2_1;
	wire w_dff_B_aCNE0rnf2_1;
	wire w_dff_B_zi007nmq0_1;
	wire w_dff_B_zHr8XPjf7_1;
	wire w_dff_B_QVu79ELB2_1;
	wire w_dff_B_rpOfhEHv6_1;
	wire w_dff_B_kW7Ee0re6_1;
	wire w_dff_B_O1W0Lwt47_1;
	wire w_dff_B_5P8jtjQX2_1;
	wire w_dff_B_WIAfGV192_1;
	wire w_dff_B_PX7GPVOA0_1;
	wire w_dff_B_0idppEZJ3_1;
	wire w_dff_B_XoIYF6co2_1;
	wire w_dff_B_c93rijkr7_1;
	wire w_dff_B_2xgoZpIf0_1;
	wire w_dff_B_WyJIYZMM9_1;
	wire w_dff_B_9aIXKL2h6_1;
	wire w_dff_B_ArO8sxJ99_1;
	wire w_dff_B_B6nLJOJA8_1;
	wire w_dff_B_dlr1o53y1_1;
	wire w_dff_B_s88bDLvV1_1;
	wire w_dff_B_jhR3FbZ11_1;
	wire w_dff_B_Hu4pUPJp1_1;
	wire w_dff_B_bEJ5Q8kn7_1;
	wire w_dff_B_6b8ZfWk11_1;
	wire w_dff_B_MqGZ9eEe7_1;
	wire w_dff_B_9Ggorrgr6_0;
	wire w_dff_B_ug1THLAA8_0;
	wire w_dff_B_p2njF8Wy0_0;
	wire w_dff_B_7BqpENEe4_0;
	wire w_dff_B_VQ8RXdVW7_0;
	wire w_dff_B_m0Aee3JC2_0;
	wire w_dff_B_5rh7trX38_0;
	wire w_dff_B_yGaqTppP6_0;
	wire w_dff_B_eg2ny05c4_0;
	wire w_dff_B_0VrRwCMq1_0;
	wire w_dff_B_s2sZnpMk3_0;
	wire w_dff_B_214eGyoe3_0;
	wire w_dff_B_YmbertBM1_0;
	wire w_dff_B_iNuIMc615_0;
	wire w_dff_B_UgRoswJS6_0;
	wire w_dff_B_ol2PWX3g7_0;
	wire w_dff_B_QqvKBaoG2_0;
	wire w_dff_B_1R9OOYbQ0_0;
	wire w_dff_B_s3RzwFa12_0;
	wire w_dff_B_3BVcZBgW8_0;
	wire w_dff_B_2G1Aa0kZ9_0;
	wire w_dff_B_45XYBINy1_0;
	wire w_dff_B_ynroTsRQ3_0;
	wire w_dff_B_EN9YDQum1_0;
	wire w_dff_B_NkzF3NyE6_0;
	wire w_dff_B_jhDoapJP3_0;
	wire w_dff_B_ip3MrRlz8_0;
	wire w_dff_B_1F86GwH13_0;
	wire w_dff_B_7JgE58Gx7_0;
	wire w_dff_B_ppIkGrU39_0;
	wire w_dff_B_znPY8YBC7_0;
	wire w_dff_B_Cz4WtRxM5_1;
	wire w_dff_B_hX4DDc072_1;
	wire w_dff_B_vO4oC1wC1_1;
	wire w_dff_B_N4QkzRah0_1;
	wire w_dff_B_noq5BmFc8_1;
	wire w_dff_B_wot6X4XY2_1;
	wire w_dff_B_SoZ8p6EM4_1;
	wire w_dff_B_AzSalxIW5_1;
	wire w_dff_B_8lhDmClm5_1;
	wire w_dff_B_upPOgiH16_1;
	wire w_dff_B_vdn2loSW0_1;
	wire w_dff_B_ovjpKjld3_1;
	wire w_dff_B_iF3FEifp1_1;
	wire w_dff_B_bCE7ygWT0_1;
	wire w_dff_B_2WFUWllr6_1;
	wire w_dff_B_Hn1ui6Rj0_1;
	wire w_dff_B_6Ko2H74B0_1;
	wire w_dff_B_kOy0lbw30_1;
	wire w_dff_B_v1EP3kgw5_1;
	wire w_dff_B_9zav3DDa1_1;
	wire w_dff_B_orFt2uhv8_1;
	wire w_dff_B_lOUweBA10_1;
	wire w_dff_B_pAQzK9x95_1;
	wire w_dff_B_4FvCS16N8_1;
	wire w_dff_B_KXpwsZS63_1;
	wire w_dff_B_kd2gB3L62_1;
	wire w_dff_B_QVdUCIrd3_1;
	wire w_dff_B_Q3XMAHfH4_1;
	wire w_dff_B_LTDwHoxl1_1;
	wire w_dff_B_fYp7rwhu5_1;
	wire w_dff_B_KVAaujiM8_0;
	wire w_dff_B_qau2pyoL4_0;
	wire w_dff_B_cERkMASt4_0;
	wire w_dff_B_CL07I3La5_0;
	wire w_dff_B_VekVdwrf9_0;
	wire w_dff_B_gw8GjGg32_0;
	wire w_dff_B_dIFaRqJ38_0;
	wire w_dff_B_s0SY6L6P3_0;
	wire w_dff_B_xZqCvfWm9_0;
	wire w_dff_B_rR833kho1_0;
	wire w_dff_B_f4Hjsnyc5_0;
	wire w_dff_B_HIFK3fD29_0;
	wire w_dff_B_7GAWPKnJ8_0;
	wire w_dff_B_pMq7HHim5_0;
	wire w_dff_B_Hpll6Zaz4_0;
	wire w_dff_B_3bOyimU30_0;
	wire w_dff_B_0r66Rra19_0;
	wire w_dff_B_sc2CgKKH6_0;
	wire w_dff_B_bhTrfgfj9_0;
	wire w_dff_B_zBU8oC3W8_0;
	wire w_dff_B_Wp6clGhC6_0;
	wire w_dff_B_gyKCnTy02_0;
	wire w_dff_B_mue6Cm2y2_0;
	wire w_dff_B_sBWbgYsk6_0;
	wire w_dff_B_DobI48jM4_0;
	wire w_dff_B_Iae9FgpR7_0;
	wire w_dff_B_SW8NICzc1_0;
	wire w_dff_B_jrdi6QfX3_0;
	wire w_dff_B_FuBS1k7T9_0;
	wire w_dff_B_norHvl765_0;
	wire w_dff_B_M14cBlRa3_1;
	wire w_dff_B_5uJWKH683_1;
	wire w_dff_B_ORDz8jHr0_1;
	wire w_dff_B_Y9B4bwQp3_1;
	wire w_dff_B_SXpLQFZD3_1;
	wire w_dff_B_HVIgRfMF6_1;
	wire w_dff_B_9zRL7yZl3_1;
	wire w_dff_B_5P3N4tZX5_1;
	wire w_dff_B_1UtBCH3i9_1;
	wire w_dff_B_6qhYjcvS4_1;
	wire w_dff_B_yBwEhq9Y5_1;
	wire w_dff_B_vKMEa47W2_1;
	wire w_dff_B_tSIC5Z2N9_1;
	wire w_dff_B_R4LvJLUz9_1;
	wire w_dff_B_f4LXkT1g6_1;
	wire w_dff_B_k0qWQIyd3_1;
	wire w_dff_B_I3VXEj6g5_1;
	wire w_dff_B_nHVGy9fB0_1;
	wire w_dff_B_JLI54C3i4_1;
	wire w_dff_B_6GlsA9Pl1_1;
	wire w_dff_B_baVt6ZSl9_1;
	wire w_dff_B_3xuXNVe27_1;
	wire w_dff_B_DytvXwob2_1;
	wire w_dff_B_ddtiVxdK6_1;
	wire w_dff_B_bTFY9pP37_1;
	wire w_dff_B_Z8zTQmtf6_1;
	wire w_dff_B_vlazR5UV4_1;
	wire w_dff_B_ycAvA3bo6_1;
	wire w_dff_B_8BjQK9zd0_1;
	wire w_dff_B_K955MgLd2_0;
	wire w_dff_B_0bFrWliJ3_0;
	wire w_dff_B_u3xurdFd9_0;
	wire w_dff_B_qEPqL1lz8_0;
	wire w_dff_B_FRy9Sbe00_0;
	wire w_dff_B_usV5zQIJ5_0;
	wire w_dff_B_ZCAcNYzC6_0;
	wire w_dff_B_mfWO26go4_0;
	wire w_dff_B_7j8eGKHU3_0;
	wire w_dff_B_CReshun12_0;
	wire w_dff_B_6TAgUcO31_0;
	wire w_dff_B_GjDh4VHQ9_0;
	wire w_dff_B_6hsWPD6h3_0;
	wire w_dff_B_2SC8oVLH8_0;
	wire w_dff_B_ZpiByu876_0;
	wire w_dff_B_FzaFPmnd4_0;
	wire w_dff_B_EkXR9rup5_0;
	wire w_dff_B_9EgvbX9c9_0;
	wire w_dff_B_qGVosCTG1_0;
	wire w_dff_B_1DYf3zti2_0;
	wire w_dff_B_k3atWQ127_0;
	wire w_dff_B_KqOdcc988_0;
	wire w_dff_B_0ldvzPUH2_0;
	wire w_dff_B_VRpTGNTt2_0;
	wire w_dff_B_XRq1WP6W0_0;
	wire w_dff_B_STiWvv1c6_0;
	wire w_dff_B_5GKmYqIk5_0;
	wire w_dff_B_dxJBpCHf6_0;
	wire w_dff_B_qICniHxc5_0;
	wire w_dff_B_WwGsn7LM4_1;
	wire w_dff_B_f5ScmcyJ6_1;
	wire w_dff_B_aCLgWyNj8_1;
	wire w_dff_B_NSG7h4PV7_1;
	wire w_dff_B_Nm7SQCST1_1;
	wire w_dff_B_jHSFzABG5_1;
	wire w_dff_B_pdZ06Urv9_1;
	wire w_dff_B_nG97F2Ex8_1;
	wire w_dff_B_c7ZVKITz0_1;
	wire w_dff_B_Gt7NUnjt0_1;
	wire w_dff_B_VbnvtDzw0_1;
	wire w_dff_B_sCBkMioo1_1;
	wire w_dff_B_mlholDQR6_1;
	wire w_dff_B_ASDanwoZ2_1;
	wire w_dff_B_NmEhouA63_1;
	wire w_dff_B_puvOBG1g8_1;
	wire w_dff_B_3ALvuP1T5_1;
	wire w_dff_B_rA6yFVJI6_1;
	wire w_dff_B_4CQIpvhh0_1;
	wire w_dff_B_9rjun1La0_1;
	wire w_dff_B_OxW1yAXT0_1;
	wire w_dff_B_cKJveguF8_1;
	wire w_dff_B_tHXTKG4t0_1;
	wire w_dff_B_dQwJwBfQ7_1;
	wire w_dff_B_OgDtmjCn6_1;
	wire w_dff_B_ET19mGkv9_1;
	wire w_dff_B_dbGglKDe6_1;
	wire w_dff_B_2YMJeXnr4_1;
	wire w_dff_B_jB9dqKE43_0;
	wire w_dff_B_Xa6ExE5U8_0;
	wire w_dff_B_Xe2eAvbj2_0;
	wire w_dff_B_utP8Au306_0;
	wire w_dff_B_pJQs1Bcx6_0;
	wire w_dff_B_7Z1s3hJ50_0;
	wire w_dff_B_2yVGrjXx0_0;
	wire w_dff_B_PshY9lv55_0;
	wire w_dff_B_CkzlWNUu7_0;
	wire w_dff_B_XrQqis6x0_0;
	wire w_dff_B_zd0ukQpz7_0;
	wire w_dff_B_qB9AiSgF4_0;
	wire w_dff_B_6lqgn5wN8_0;
	wire w_dff_B_UurPIyiQ3_0;
	wire w_dff_B_AZTO00TC7_0;
	wire w_dff_B_1zuWxfB68_0;
	wire w_dff_B_yVylfGHH5_0;
	wire w_dff_B_2pixfssf7_0;
	wire w_dff_B_bqLpzn4O5_0;
	wire w_dff_B_cLRNaMk04_0;
	wire w_dff_B_dWHjnBLA2_0;
	wire w_dff_B_Sp28x1Ar4_0;
	wire w_dff_B_STtDZsFd2_0;
	wire w_dff_B_k6gMftkm4_0;
	wire w_dff_B_v4YSt8vz1_0;
	wire w_dff_B_mQg6QTo99_0;
	wire w_dff_B_rAcpl1I21_0;
	wire w_dff_B_X8LY3C7p1_0;
	wire w_dff_B_jEbGC2eA4_1;
	wire w_dff_B_N1xf8Rcn6_1;
	wire w_dff_B_Muv2PFjB5_1;
	wire w_dff_B_xw8Q4aK42_1;
	wire w_dff_B_p7z4SON57_1;
	wire w_dff_B_7jxHsP4f2_1;
	wire w_dff_B_ViqrtEds8_1;
	wire w_dff_B_hPARAbyN5_1;
	wire w_dff_B_QjBjnzj84_1;
	wire w_dff_B_Yyp7tIBm2_1;
	wire w_dff_B_x3H8XNX06_1;
	wire w_dff_B_8EszFODT5_1;
	wire w_dff_B_81DWx3yH1_1;
	wire w_dff_B_DvNlnxOf2_1;
	wire w_dff_B_pJ6Gmn2H1_1;
	wire w_dff_B_giWiqLOj7_1;
	wire w_dff_B_UY4LD7Fn5_1;
	wire w_dff_B_Vp0VVceo5_1;
	wire w_dff_B_0GsAUBrv1_1;
	wire w_dff_B_2QT99DA90_1;
	wire w_dff_B_6PQDSOM19_1;
	wire w_dff_B_SKkqFQD85_1;
	wire w_dff_B_PZ5OFXo40_1;
	wire w_dff_B_mcYUlvgW4_1;
	wire w_dff_B_W1aVsd749_1;
	wire w_dff_B_zPLs8g880_1;
	wire w_dff_B_UIEJM1lk8_1;
	wire w_dff_B_AWw7MNe60_0;
	wire w_dff_B_kF1uaxWH8_0;
	wire w_dff_B_a28HfzOT6_0;
	wire w_dff_B_bUKqhQLd8_0;
	wire w_dff_B_UAXnDc7f5_0;
	wire w_dff_B_EI4oPBKI2_0;
	wire w_dff_B_K9sMFS0A1_0;
	wire w_dff_B_Sg9hxv1q9_0;
	wire w_dff_B_CMnCBKYk6_0;
	wire w_dff_B_BbvIvvKF4_0;
	wire w_dff_B_4VpBNvBM1_0;
	wire w_dff_B_XYAcKEcw3_0;
	wire w_dff_B_K1Tmd6IG7_0;
	wire w_dff_B_wAtzXDS95_0;
	wire w_dff_B_TNLldSDC0_0;
	wire w_dff_B_RWGFRdYC9_0;
	wire w_dff_B_RAAQqzSZ3_0;
	wire w_dff_B_DISV63gQ0_0;
	wire w_dff_B_DhzvxISg0_0;
	wire w_dff_B_sSsDZT0G4_0;
	wire w_dff_B_QUxvVfjt7_0;
	wire w_dff_B_lDnu2xxq9_0;
	wire w_dff_B_CV1cKdzL0_0;
	wire w_dff_B_qhHkb7Ch0_0;
	wire w_dff_B_euxuPu5B7_0;
	wire w_dff_B_9Xff2Fa12_0;
	wire w_dff_B_d3Bc1Lmg9_0;
	wire w_dff_B_m47kjmmf6_1;
	wire w_dff_B_zEKrbGf94_1;
	wire w_dff_B_H1UwU8lb9_1;
	wire w_dff_B_cJefzE431_1;
	wire w_dff_B_upxIZDjY4_1;
	wire w_dff_B_p0hMUHHl6_1;
	wire w_dff_B_SD1wIlEX0_1;
	wire w_dff_B_UXLwP4lR4_1;
	wire w_dff_B_MsRu5ljh5_1;
	wire w_dff_B_aSlCRTCN1_1;
	wire w_dff_B_Yjl4ESYk8_1;
	wire w_dff_B_jq0aeaTg8_1;
	wire w_dff_B_mSQQUG2e5_1;
	wire w_dff_B_vmZPRSBL5_1;
	wire w_dff_B_W3oA2bFZ1_1;
	wire w_dff_B_qhDGW6su6_1;
	wire w_dff_B_XrYy7vtE8_1;
	wire w_dff_B_gTMcphaj8_1;
	wire w_dff_B_LuUPDFaz9_1;
	wire w_dff_B_eVAlL21p9_1;
	wire w_dff_B_gGkGFiGi3_1;
	wire w_dff_B_sYS25J7f9_1;
	wire w_dff_B_YYnhOVjW6_1;
	wire w_dff_B_qpi6SN8X2_1;
	wire w_dff_B_LQskBW503_1;
	wire w_dff_B_YvVPAofT6_1;
	wire w_dff_B_6LkOjHvA7_0;
	wire w_dff_B_4XYmqwGw4_0;
	wire w_dff_B_iolOQF2d8_0;
	wire w_dff_B_RnfMtriw1_0;
	wire w_dff_B_sUsicH7W0_0;
	wire w_dff_B_QJnco1Dq8_0;
	wire w_dff_B_Hh5ikDDx5_0;
	wire w_dff_B_IR9jkgZl4_0;
	wire w_dff_B_scrGlXOA1_0;
	wire w_dff_B_V1Yi3vbE7_0;
	wire w_dff_B_UobApmHn1_0;
	wire w_dff_B_bePznbIU0_0;
	wire w_dff_B_wPzL3Mn84_0;
	wire w_dff_B_5s9X372m0_0;
	wire w_dff_B_g9XD0cEj8_0;
	wire w_dff_B_DRy4QOlE3_0;
	wire w_dff_B_p395qPK33_0;
	wire w_dff_B_H9PsgRw26_0;
	wire w_dff_B_pXTfVs3i5_0;
	wire w_dff_B_H3VVbSMP6_0;
	wire w_dff_B_FvACIz0R3_0;
	wire w_dff_B_3u3wk3C94_0;
	wire w_dff_B_g8Cm3rJN0_0;
	wire w_dff_B_HIycXObK2_0;
	wire w_dff_B_CT7QS0sv9_0;
	wire w_dff_B_bFwFmeEw7_0;
	wire w_dff_B_Wb0mxUq91_1;
	wire w_dff_B_WiO3QQhK2_1;
	wire w_dff_B_GYWvVFsF0_1;
	wire w_dff_B_qhkzfFXX1_1;
	wire w_dff_B_nylJwnYH2_1;
	wire w_dff_B_pdQynfY53_1;
	wire w_dff_B_FbVuU11Y5_1;
	wire w_dff_B_uEDEhPiX2_1;
	wire w_dff_B_VGYtJ86v7_1;
	wire w_dff_B_2QwbOco99_1;
	wire w_dff_B_B9VzruyW8_1;
	wire w_dff_B_5l5KD6jS0_1;
	wire w_dff_B_uhAMMFSz4_1;
	wire w_dff_B_WJ0QK7hy6_1;
	wire w_dff_B_1URQWq077_1;
	wire w_dff_B_GTxav8wm7_1;
	wire w_dff_B_WDFwtscJ7_1;
	wire w_dff_B_8qsrFrGL2_1;
	wire w_dff_B_Zm5x2N2B7_1;
	wire w_dff_B_0pT00Q9e4_1;
	wire w_dff_B_RzrTjCVQ8_1;
	wire w_dff_B_QElwnxde8_1;
	wire w_dff_B_fdLvrelX7_1;
	wire w_dff_B_Gzqg4BA45_1;
	wire w_dff_B_nk8Q4hzv5_1;
	wire w_dff_B_db5T3eSR1_0;
	wire w_dff_B_AYPQc4Vq2_0;
	wire w_dff_B_jHtMmMs17_0;
	wire w_dff_B_UHjYbtox8_0;
	wire w_dff_B_sYdTR8HW9_0;
	wire w_dff_B_QPRMV83g6_0;
	wire w_dff_B_TY2eUKX81_0;
	wire w_dff_B_duOTAfbj6_0;
	wire w_dff_B_0LrOqCnH6_0;
	wire w_dff_B_G6daYLZo1_0;
	wire w_dff_B_WT7QBB8j8_0;
	wire w_dff_B_UXiN6msR9_0;
	wire w_dff_B_z0k8JdLs2_0;
	wire w_dff_B_tvfgLy9T5_0;
	wire w_dff_B_YBtL3Jbo1_0;
	wire w_dff_B_xjmg3mpv1_0;
	wire w_dff_B_vDtxa8cd9_0;
	wire w_dff_B_4e90aYLG8_0;
	wire w_dff_B_i3Jja0yv6_0;
	wire w_dff_B_HQalQ15v3_0;
	wire w_dff_B_Q8dyLceV7_0;
	wire w_dff_B_rBGac74U7_0;
	wire w_dff_B_f359shWt5_0;
	wire w_dff_B_VuXxQXSH5_0;
	wire w_dff_B_kc8HMq882_0;
	wire w_dff_B_AnRFY6P59_1;
	wire w_dff_B_1ilWoncE7_1;
	wire w_dff_B_TtVvSwnO9_1;
	wire w_dff_B_2e2GW7yY0_1;
	wire w_dff_B_XfbvT7Nc6_1;
	wire w_dff_B_ahL5U5e97_1;
	wire w_dff_B_8pAs6gXb9_1;
	wire w_dff_B_pzbWGiv33_1;
	wire w_dff_B_zmTmNv9A8_1;
	wire w_dff_B_SFd7vEGX0_1;
	wire w_dff_B_mPM0y6mF0_1;
	wire w_dff_B_Fg9q1f5W4_1;
	wire w_dff_B_hby8E9yb4_1;
	wire w_dff_B_KO7H60of7_1;
	wire w_dff_B_esIAVLEp6_1;
	wire w_dff_B_NmX60Cay4_1;
	wire w_dff_B_VSgvxO1I9_1;
	wire w_dff_B_XhQg9Mxx1_1;
	wire w_dff_B_qHdW0Lby3_1;
	wire w_dff_B_0rJbQZPN9_1;
	wire w_dff_B_UqtMZYYs4_1;
	wire w_dff_B_2STSG4oh5_1;
	wire w_dff_B_FXFRtHln0_1;
	wire w_dff_B_mAYLtnxH0_1;
	wire w_dff_B_ORB5OVYO5_0;
	wire w_dff_B_dsD3knkv5_0;
	wire w_dff_B_rBiIlAy80_0;
	wire w_dff_B_0wGjaba27_0;
	wire w_dff_B_RgCIjfmT8_0;
	wire w_dff_B_BQDcfmLy4_0;
	wire w_dff_B_xUWZgGL89_0;
	wire w_dff_B_hsB7URDw7_0;
	wire w_dff_B_phT04UDP8_0;
	wire w_dff_B_FQMjJqiN4_0;
	wire w_dff_B_C64ubjqN9_0;
	wire w_dff_B_EUN409DQ7_0;
	wire w_dff_B_2dXi4wSe8_0;
	wire w_dff_B_JCRcWhEw7_0;
	wire w_dff_B_3HENdVeT2_0;
	wire w_dff_B_lutsWKzk8_0;
	wire w_dff_B_iXN2t8V27_0;
	wire w_dff_B_uft6ISGb8_0;
	wire w_dff_B_qNlsMg7G1_0;
	wire w_dff_B_2PO0njAe1_0;
	wire w_dff_B_PsqNBR7s9_0;
	wire w_dff_B_7Ptke34g1_0;
	wire w_dff_B_duuzWikO5_0;
	wire w_dff_B_WEHr8swc1_0;
	wire w_dff_B_7edgnBR81_1;
	wire w_dff_B_0MAQMHq53_1;
	wire w_dff_B_QQdnpqgp6_1;
	wire w_dff_B_piijkjuC6_1;
	wire w_dff_B_EqSLs5iI7_1;
	wire w_dff_B_3AwOmlqM8_1;
	wire w_dff_B_AGCKqSXE6_1;
	wire w_dff_B_flH8TDKj3_1;
	wire w_dff_B_HR7UytV38_1;
	wire w_dff_B_39c2frOG5_1;
	wire w_dff_B_CiMxmFWS0_1;
	wire w_dff_B_Duad9wHL9_1;
	wire w_dff_B_mUQ0sMOW8_1;
	wire w_dff_B_xH0H4AfA9_1;
	wire w_dff_B_MBpaSc8S3_1;
	wire w_dff_B_9VgXWMOX3_1;
	wire w_dff_B_rMCj5kZg9_1;
	wire w_dff_B_LEkqTHx12_1;
	wire w_dff_B_8gaKvIj29_1;
	wire w_dff_B_IPopdG0o3_1;
	wire w_dff_B_CdY3vwIN9_1;
	wire w_dff_B_QYAa0j5h3_1;
	wire w_dff_B_fxvTyWRy8_1;
	wire w_dff_B_VxcVUf7H5_0;
	wire w_dff_B_BJxiAccS9_0;
	wire w_dff_B_vh1CGSU90_0;
	wire w_dff_B_qhTbMA485_0;
	wire w_dff_B_gH3C0luF2_0;
	wire w_dff_B_O6BkGu1Z7_0;
	wire w_dff_B_ubtcXv1d0_0;
	wire w_dff_B_huwtojip9_0;
	wire w_dff_B_wNLgOwHR6_0;
	wire w_dff_B_yboVqc1q9_0;
	wire w_dff_B_UTxHv5kQ9_0;
	wire w_dff_B_WGzj0TcJ3_0;
	wire w_dff_B_Io800KAz5_0;
	wire w_dff_B_cjg6KSmO8_0;
	wire w_dff_B_nH0wW2JQ2_0;
	wire w_dff_B_CGyoJYNY3_0;
	wire w_dff_B_CjT98AnT2_0;
	wire w_dff_B_NFjf6lvI5_0;
	wire w_dff_B_mKaBape88_0;
	wire w_dff_B_IG5BdfI66_0;
	wire w_dff_B_iCQC6N7R7_0;
	wire w_dff_B_YCCdy70h4_0;
	wire w_dff_B_vffmUHZP1_0;
	wire w_dff_B_DXhPNNpz1_1;
	wire w_dff_B_mTtX9v0t9_1;
	wire w_dff_B_Y2ANFewa3_1;
	wire w_dff_B_jgzopvEA0_1;
	wire w_dff_B_Aq5Ikao38_1;
	wire w_dff_B_UhfBFeYt6_1;
	wire w_dff_B_fHb0j4ew5_1;
	wire w_dff_B_hEoaFcUm6_1;
	wire w_dff_B_6JB7cQ9z3_1;
	wire w_dff_B_jpBio3oi6_1;
	wire w_dff_B_cS71ko3Z0_1;
	wire w_dff_B_tP12ks5X0_1;
	wire w_dff_B_P0wl6mZ51_1;
	wire w_dff_B_BeJoeIXj7_1;
	wire w_dff_B_79b0qMv45_1;
	wire w_dff_B_vnx7SaAd2_1;
	wire w_dff_B_Lk6oOYTe4_1;
	wire w_dff_B_mL0PLyNd4_1;
	wire w_dff_B_wFhZGdBy9_1;
	wire w_dff_B_O0Gb9j260_1;
	wire w_dff_B_BMUS3aHp6_1;
	wire w_dff_B_tOY8ECp76_1;
	wire w_dff_B_GwfYFLQG5_0;
	wire w_dff_B_CS57lDA07_0;
	wire w_dff_B_By5F7GgY5_0;
	wire w_dff_B_RtcdwQQd6_0;
	wire w_dff_B_7Do5rFZp5_0;
	wire w_dff_B_WOqwXhkh7_0;
	wire w_dff_B_IxbFk8cI6_0;
	wire w_dff_B_0bOUT9uw7_0;
	wire w_dff_B_kwMH0CsE1_0;
	wire w_dff_B_jOj3r1vQ2_0;
	wire w_dff_B_sfI0GuZh1_0;
	wire w_dff_B_haoZ0fGm4_0;
	wire w_dff_B_QDtWVFUm6_0;
	wire w_dff_B_VSll0QuP2_0;
	wire w_dff_B_s0KFDVXq0_0;
	wire w_dff_B_lPBRUhZt3_0;
	wire w_dff_B_T52oUi9m8_0;
	wire w_dff_B_QIfhqqZY6_0;
	wire w_dff_B_h1TRqlBE7_0;
	wire w_dff_B_xxmYYP6a8_0;
	wire w_dff_B_y6CzhVen1_0;
	wire w_dff_B_nKZIowO61_0;
	wire w_dff_B_cnQQSUWE9_1;
	wire w_dff_B_oUTwsU4C2_1;
	wire w_dff_B_zlOAONAj5_1;
	wire w_dff_B_IFtzdkkf5_1;
	wire w_dff_B_Nu8LDJL90_1;
	wire w_dff_B_FvjXZquD1_1;
	wire w_dff_B_FK3KUyQ09_1;
	wire w_dff_B_ogbSYZp63_1;
	wire w_dff_B_lR3wgXjs6_1;
	wire w_dff_B_rnEWP2BY7_1;
	wire w_dff_B_nl7gEe5Z0_1;
	wire w_dff_B_syBgmKT68_1;
	wire w_dff_B_pvIK8Qgf1_1;
	wire w_dff_B_ZPySYxyv9_1;
	wire w_dff_B_1b9OPo4x8_1;
	wire w_dff_B_qAcmV4t20_1;
	wire w_dff_B_8r8vNDIX4_1;
	wire w_dff_B_zECH9nE16_1;
	wire w_dff_B_cXOIeajH7_1;
	wire w_dff_B_GNMk3aiO0_1;
	wire w_dff_B_k8b5cujs9_1;
	wire w_dff_B_LhQmirqn3_0;
	wire w_dff_B_3m5Josyl8_0;
	wire w_dff_B_MPMk29jj0_0;
	wire w_dff_B_Orp2IKKa9_0;
	wire w_dff_B_hxwCphf05_0;
	wire w_dff_B_fXmjm7Bw7_0;
	wire w_dff_B_Fg94zmG79_0;
	wire w_dff_B_Yarf2wHy0_0;
	wire w_dff_B_xgEYqYuX6_0;
	wire w_dff_B_n4gDINIR7_0;
	wire w_dff_B_IqiUbNfT0_0;
	wire w_dff_B_n6VTFJq68_0;
	wire w_dff_B_ieku2ZGi2_0;
	wire w_dff_B_3GFJHEF15_0;
	wire w_dff_B_FXOG0ofc5_0;
	wire w_dff_B_kxgwOpN27_0;
	wire w_dff_B_U8RnmLws4_0;
	wire w_dff_B_sCjKKZX31_0;
	wire w_dff_B_ZJUtsRPy0_0;
	wire w_dff_B_mO2p0KBo5_0;
	wire w_dff_B_TpJykMPA5_0;
	wire w_dff_B_xa5x4JPM2_1;
	wire w_dff_B_av4abSpH4_1;
	wire w_dff_B_7RVwqZRE9_1;
	wire w_dff_B_EpxKxves7_1;
	wire w_dff_B_dahhMMJK4_1;
	wire w_dff_B_bTUnJ4mk9_1;
	wire w_dff_B_FtDA7Hzj1_1;
	wire w_dff_B_jVOJ518L1_1;
	wire w_dff_B_YrimiXEq6_1;
	wire w_dff_B_fwlunybC8_1;
	wire w_dff_B_SRurwE5R8_1;
	wire w_dff_B_pcsLQWjT7_1;
	wire w_dff_B_I4OBEttl2_1;
	wire w_dff_B_d9HUysRq7_1;
	wire w_dff_B_z3ugAY2a0_1;
	wire w_dff_B_1lZkDcvQ6_1;
	wire w_dff_B_3ZXPQKqH3_1;
	wire w_dff_B_k3RquIqD7_1;
	wire w_dff_B_LlQSbhOp9_1;
	wire w_dff_B_wFlt2aWE8_1;
	wire w_dff_B_H3SsZrFy0_0;
	wire w_dff_B_H5otAfpI1_0;
	wire w_dff_B_9b3gyfzp3_0;
	wire w_dff_B_cVUdhSle8_0;
	wire w_dff_B_E2LqWjd31_0;
	wire w_dff_B_iANMbePJ3_0;
	wire w_dff_B_204ll75a2_0;
	wire w_dff_B_Qpz3pLeL0_0;
	wire w_dff_B_RdFzMQdt7_0;
	wire w_dff_B_nun3bSB21_0;
	wire w_dff_B_2oQtiWqH0_0;
	wire w_dff_B_D7yUlmOE0_0;
	wire w_dff_B_HjwDF7Qh8_0;
	wire w_dff_B_lxJyeo6e9_0;
	wire w_dff_B_Rptzv1ER2_0;
	wire w_dff_B_P6S8frr96_0;
	wire w_dff_B_sgXZrIhN5_0;
	wire w_dff_B_JPDt3g8i0_0;
	wire w_dff_B_RpyLTre07_0;
	wire w_dff_B_srqfiaFR0_0;
	wire w_dff_B_7xK6EmhU6_1;
	wire w_dff_B_SPsZqQtm8_1;
	wire w_dff_B_imSWdBGf4_1;
	wire w_dff_B_VGJaJ7kk0_1;
	wire w_dff_B_SGCN2dbh9_1;
	wire w_dff_B_ZCKVZTnK8_1;
	wire w_dff_B_jDUYEp0T5_1;
	wire w_dff_B_Z3LhNeMH3_1;
	wire w_dff_B_TqNQSCfI3_1;
	wire w_dff_B_vBA2cLxo4_1;
	wire w_dff_B_fEmIoLXP6_1;
	wire w_dff_B_CysGEYLx3_1;
	wire w_dff_B_ukjc9Gao2_1;
	wire w_dff_B_sGVK40HI1_1;
	wire w_dff_B_cdALOMMl5_1;
	wire w_dff_B_duGQQq2r0_1;
	wire w_dff_B_LwqrRRbV9_1;
	wire w_dff_B_o61DiKme9_1;
	wire w_dff_B_eyYJitxH0_1;
	wire w_dff_B_8w5aLc5T3_0;
	wire w_dff_B_gJywaFgx6_0;
	wire w_dff_B_aBDAsdZZ9_0;
	wire w_dff_B_Q5n57uH98_0;
	wire w_dff_B_JCX5X2EQ6_0;
	wire w_dff_B_YMf9Wzeq2_0;
	wire w_dff_B_xxDpY2CJ6_0;
	wire w_dff_B_iWetE3sI0_0;
	wire w_dff_B_OFNgbhx92_0;
	wire w_dff_B_gMdIllk53_0;
	wire w_dff_B_7jKOpOTx5_0;
	wire w_dff_B_SZvlTEXt2_0;
	wire w_dff_B_yW0M5Jdg2_0;
	wire w_dff_B_glbPXlE80_0;
	wire w_dff_B_iCpyig4C6_0;
	wire w_dff_B_VkNIvHyH4_0;
	wire w_dff_B_5aHwBBEa3_0;
	wire w_dff_B_TNHDgILC3_0;
	wire w_dff_B_CcU9AiUi0_0;
	wire w_dff_B_DsqcDONC2_1;
	wire w_dff_B_qEY7xbD11_1;
	wire w_dff_B_AZSKonBw8_1;
	wire w_dff_B_T86nmV2p3_1;
	wire w_dff_B_1fBNeVli2_1;
	wire w_dff_B_82Rxo4n26_1;
	wire w_dff_B_99fEhW9B9_1;
	wire w_dff_B_M1gUdRdO6_1;
	wire w_dff_B_idh8pFW65_1;
	wire w_dff_B_Ew5zMVam9_1;
	wire w_dff_B_hMLPG4LO5_1;
	wire w_dff_B_EEc5s4PX5_1;
	wire w_dff_B_qdyNlzfl1_1;
	wire w_dff_B_AW4wJHbW8_1;
	wire w_dff_B_lLRNHaXk1_1;
	wire w_dff_B_nUz2s5yt4_1;
	wire w_dff_B_pP5A4g558_1;
	wire w_dff_B_EWKSzcRm1_1;
	wire w_dff_B_qPGFOp2M9_0;
	wire w_dff_B_Q6xMljOf6_0;
	wire w_dff_B_TzODdsoK2_0;
	wire w_dff_B_1HHyb4Xq0_0;
	wire w_dff_B_aGWFNs8B4_0;
	wire w_dff_B_atTLjLDJ8_0;
	wire w_dff_B_akv8Vddd3_0;
	wire w_dff_B_QOhnN9BP5_0;
	wire w_dff_B_ak1MbCZO2_0;
	wire w_dff_B_eubY1vOU3_0;
	wire w_dff_B_OeRke0uK6_0;
	wire w_dff_B_JX7VGQvK9_0;
	wire w_dff_B_mOpQjRKP9_0;
	wire w_dff_B_upekkd5I8_0;
	wire w_dff_B_Vql2Za4h8_0;
	wire w_dff_B_QMvYmRMk4_0;
	wire w_dff_B_IGdmWZAf5_0;
	wire w_dff_B_bS2zNEr15_0;
	wire w_dff_B_DtGIA1Qr8_1;
	wire w_dff_B_TClm6Gwg8_1;
	wire w_dff_B_cQPMdY607_1;
	wire w_dff_B_OWOQHXBv3_1;
	wire w_dff_B_zJjkWGXe6_1;
	wire w_dff_B_3jo62fHS0_1;
	wire w_dff_B_hSUjpPmh8_1;
	wire w_dff_B_Ub5VEuQF6_1;
	wire w_dff_B_peaUIY4i2_1;
	wire w_dff_B_SW51JjHT7_1;
	wire w_dff_B_Lla3yk331_1;
	wire w_dff_B_1PU1J8NF4_1;
	wire w_dff_B_RGGE4mWw1_1;
	wire w_dff_B_CQkr8GgQ9_1;
	wire w_dff_B_ejvwjjJS3_1;
	wire w_dff_B_aIm1Iwxd0_1;
	wire w_dff_B_LxQ84mjb0_1;
	wire w_dff_B_4cj0w4qp2_0;
	wire w_dff_B_ttfr3fBJ7_0;
	wire w_dff_B_IjsRDjAf5_0;
	wire w_dff_B_Q4n4QISs2_0;
	wire w_dff_B_UzWE0xuc0_0;
	wire w_dff_B_G8UOLQmu2_0;
	wire w_dff_B_SRkte2WQ7_0;
	wire w_dff_B_y7IBRBiF8_0;
	wire w_dff_B_XVFsoCZ73_0;
	wire w_dff_B_5geMDvRG6_0;
	wire w_dff_B_StHB7Yd60_0;
	wire w_dff_B_AL3LKkyJ7_0;
	wire w_dff_B_lNiXWzoT9_0;
	wire w_dff_B_I0pcZiVS8_0;
	wire w_dff_B_ylFPqo4h2_0;
	wire w_dff_B_UXzqSjqs2_0;
	wire w_dff_B_M2JhGCeu4_0;
	wire w_dff_B_5S7dBTMF2_1;
	wire w_dff_B_H66g06Jv7_1;
	wire w_dff_B_eqgmM5eX7_1;
	wire w_dff_B_nrlqClN77_1;
	wire w_dff_B_zDiHmWge8_1;
	wire w_dff_B_3T24PzSq4_1;
	wire w_dff_B_6v6jhMIb4_1;
	wire w_dff_B_9YuYCD3O9_1;
	wire w_dff_B_bUSViud42_1;
	wire w_dff_B_egv2g8IU9_1;
	wire w_dff_B_Cvh92W7r2_1;
	wire w_dff_B_mowFca6I7_1;
	wire w_dff_B_hZppC5Ry8_1;
	wire w_dff_B_buqsmvbG4_1;
	wire w_dff_B_rZuwkguI5_1;
	wire w_dff_B_ghzowI0M3_1;
	wire w_dff_B_Gs3icwdR1_0;
	wire w_dff_B_2m4GT23m8_0;
	wire w_dff_B_6fJxv6bY6_0;
	wire w_dff_B_sBPeg4QF7_0;
	wire w_dff_B_DrHk8ME58_0;
	wire w_dff_B_ge20eKXn4_0;
	wire w_dff_B_YzzD5oRv5_0;
	wire w_dff_B_m4ChRGeD3_0;
	wire w_dff_B_tBNOCMDy4_0;
	wire w_dff_B_TKgZ6uI55_0;
	wire w_dff_B_Wq8VXjwJ4_0;
	wire w_dff_B_cyAFaND39_0;
	wire w_dff_B_cSwYfqwq8_0;
	wire w_dff_B_aBR3e6eT0_0;
	wire w_dff_B_w2W4jLg07_0;
	wire w_dff_B_Ps1HkcOR8_0;
	wire w_dff_B_CUOXvnUc5_1;
	wire w_dff_B_HPfjBPEr9_1;
	wire w_dff_B_PGPELzGd7_1;
	wire w_dff_B_Kb2hf6kc5_1;
	wire w_dff_B_sjwpyMU29_1;
	wire w_dff_B_tspZSzwa7_1;
	wire w_dff_B_NVQoXH6E9_1;
	wire w_dff_B_YUo1Ygd56_1;
	wire w_dff_B_6Rm8qGhB8_1;
	wire w_dff_B_lvZN4CVJ2_1;
	wire w_dff_B_gxtRfNv60_1;
	wire w_dff_B_ikB8jArh1_1;
	wire w_dff_B_odm2xBLw5_1;
	wire w_dff_B_m9q3uzCY6_1;
	wire w_dff_B_ORoqjfaO4_1;
	wire w_dff_B_sXbzJ5Q78_0;
	wire w_dff_B_rQsG1VQ11_0;
	wire w_dff_B_gHa8KuJC1_0;
	wire w_dff_B_UTQABHOg7_0;
	wire w_dff_B_AbJRHRrv1_0;
	wire w_dff_B_46AXX8fY8_0;
	wire w_dff_B_3z2JPzpZ4_0;
	wire w_dff_B_JTqh1Zvp5_0;
	wire w_dff_B_pi3yEozm0_0;
	wire w_dff_B_HQGS0GVA7_0;
	wire w_dff_B_lO38nP6x1_0;
	wire w_dff_B_sknHGjTq1_0;
	wire w_dff_B_phSHpzuI8_0;
	wire w_dff_B_YlwRzazy5_0;
	wire w_dff_B_Azuoeek25_0;
	wire w_dff_B_hyJeNg6b4_1;
	wire w_dff_B_eiqVd13B5_1;
	wire w_dff_B_zyDhBBD60_1;
	wire w_dff_B_Mi3poAXu6_1;
	wire w_dff_B_gE4KwiDc3_1;
	wire w_dff_B_Ev1G5wgk2_1;
	wire w_dff_B_fNerFjHe8_1;
	wire w_dff_B_Qe6Tvfbg1_1;
	wire w_dff_B_vcXp2qKs8_1;
	wire w_dff_B_zpcHU6sG8_1;
	wire w_dff_B_XDopxJbJ5_1;
	wire w_dff_B_vbZvn9X06_1;
	wire w_dff_B_WgGQvFyk8_1;
	wire w_dff_B_LgXnSLIA1_1;
	wire w_dff_B_fEYIY6q44_0;
	wire w_dff_B_kXVhlyVg4_0;
	wire w_dff_B_kpZkyfY87_0;
	wire w_dff_B_uy1hztZS6_0;
	wire w_dff_B_69c0OADM1_0;
	wire w_dff_B_QJzL0RRy6_0;
	wire w_dff_B_ibk2HsTc8_0;
	wire w_dff_B_86zqUp2N9_0;
	wire w_dff_B_OW9IdvrP2_0;
	wire w_dff_B_2h6rtg9U0_0;
	wire w_dff_B_TDMm0ipE7_0;
	wire w_dff_B_FxCCraqz2_0;
	wire w_dff_B_b858IeTD0_0;
	wire w_dff_B_bY5KWRW79_0;
	wire w_dff_B_EVgls9Hj2_1;
	wire w_dff_B_wKsM1TJx2_1;
	wire w_dff_B_llvWFGdo3_1;
	wire w_dff_B_hNfCcbQL1_1;
	wire w_dff_B_36yABsft3_1;
	wire w_dff_B_FMp0B9V20_1;
	wire w_dff_B_p7VG3Aqa4_1;
	wire w_dff_B_YlZbSA8n2_1;
	wire w_dff_B_GTIBmeFe0_1;
	wire w_dff_B_BjNPsRSJ7_1;
	wire w_dff_B_4bEbYv7J7_1;
	wire w_dff_B_lUDUU1OZ7_1;
	wire w_dff_B_EbOdpOXS9_1;
	wire w_dff_B_5CeuyEaX6_0;
	wire w_dff_B_a5tanuw44_0;
	wire w_dff_B_p1SXfKS10_0;
	wire w_dff_B_yHilQjpp3_0;
	wire w_dff_B_RTwv84eT1_0;
	wire w_dff_B_sI2dhu6C0_0;
	wire w_dff_B_s6pp4PGW1_0;
	wire w_dff_B_NlD4pJqc0_0;
	wire w_dff_B_1AX1uVCb8_0;
	wire w_dff_B_VugXbhlk9_0;
	wire w_dff_B_q5dE9HBj3_0;
	wire w_dff_B_RKWmxwpd3_0;
	wire w_dff_B_hz8fGERr9_0;
	wire w_dff_B_xgqsNOXB1_1;
	wire w_dff_B_NWHntx2t2_1;
	wire w_dff_B_AlPmFwRW4_1;
	wire w_dff_B_2a8lfKA75_1;
	wire w_dff_B_XxLjBnFw8_1;
	wire w_dff_B_NBWtTwgR2_1;
	wire w_dff_B_Okr54iu12_1;
	wire w_dff_B_6Jsg1KBg1_1;
	wire w_dff_B_g5zSm0bu7_1;
	wire w_dff_B_FPt83beR7_1;
	wire w_dff_B_8JMvHWgE6_1;
	wire w_dff_B_Uziv0Vnv8_1;
	wire w_dff_B_9AR7u68N2_0;
	wire w_dff_B_TbnkcOLG4_0;
	wire w_dff_B_RR9bi7VC1_0;
	wire w_dff_B_oT1a1THS1_0;
	wire w_dff_B_uZLVjhAF8_0;
	wire w_dff_B_DHQwpGTR8_0;
	wire w_dff_B_u02w9fFj6_0;
	wire w_dff_B_sfoT66hB2_0;
	wire w_dff_B_dmAlHyGz0_0;
	wire w_dff_B_8Ts70Iic0_0;
	wire w_dff_B_M0RIAs7T5_0;
	wire w_dff_B_PT2aeLqK8_0;
	wire w_dff_B_iK8IYRs33_1;
	wire w_dff_B_RvBrkqoy3_1;
	wire w_dff_B_b93Wd1dM7_1;
	wire w_dff_B_cL4TKsTY2_1;
	wire w_dff_B_8KTSPmul4_1;
	wire w_dff_B_qcBfZHT42_1;
	wire w_dff_B_WgmbwlWN9_1;
	wire w_dff_B_hl8ngWvW5_1;
	wire w_dff_B_gP2Ricw43_1;
	wire w_dff_B_FeH8ThDA8_1;
	wire w_dff_B_27LeE5x30_1;
	wire w_dff_B_WzittY0J2_0;
	wire w_dff_B_digy4ypN5_0;
	wire w_dff_B_IyXXLOIo4_0;
	wire w_dff_B_4SFULI4g1_0;
	wire w_dff_B_NHHorC111_0;
	wire w_dff_B_Qu85MC6D7_0;
	wire w_dff_B_CWlIy23N7_0;
	wire w_dff_B_FXDHyn1B9_0;
	wire w_dff_B_2pvDVzF08_0;
	wire w_dff_B_kd5CM0fw2_0;
	wire w_dff_B_nKJsQ9ti3_0;
	wire w_dff_B_u8Aqn7YY6_1;
	wire w_dff_B_2fzYDzLE3_1;
	wire w_dff_B_61jnnUxf9_1;
	wire w_dff_B_XVXDV8qX3_1;
	wire w_dff_B_a7TVaVEo9_1;
	wire w_dff_B_Dp5bon0S1_1;
	wire w_dff_B_ME01Jysm8_1;
	wire w_dff_B_hYK1Ehqo1_1;
	wire w_dff_B_C6X7E3jq9_1;
	wire w_dff_B_o5sfoxtN0_1;
	wire w_dff_B_2CqZQwGP3_0;
	wire w_dff_B_Xidoqr8P2_0;
	wire w_dff_B_PbfwgGb02_0;
	wire w_dff_B_HzSKeLUp3_0;
	wire w_dff_B_t7oo0FTl8_0;
	wire w_dff_B_k5jTnxDk4_0;
	wire w_dff_B_0NEvZZis7_0;
	wire w_dff_B_1UqxfKPV0_0;
	wire w_dff_B_2VgunHW36_0;
	wire w_dff_B_njqcx4ts3_0;
	wire w_dff_B_WZxvvIYD2_1;
	wire w_dff_B_TSlxqhxh6_1;
	wire w_dff_B_G7hfJw6t8_1;
	wire w_dff_B_KFMw82Hu5_1;
	wire w_dff_B_mfGu0USy7_1;
	wire w_dff_B_Ds146Ekz3_1;
	wire w_dff_B_42Jk9NQm2_1;
	wire w_dff_B_EbeYix8q6_1;
	wire w_dff_B_uSgQnbDf2_1;
	wire w_dff_B_vUH7yW4f1_0;
	wire w_dff_B_YJXgnpGf7_0;
	wire w_dff_B_iBuwANGT9_0;
	wire w_dff_B_UhDLPyJA2_0;
	wire w_dff_B_A5abHHqR5_0;
	wire w_dff_B_7S0Ebel80_0;
	wire w_dff_B_cIvKwSkV4_0;
	wire w_dff_B_hpnBngai8_0;
	wire w_dff_B_oTv1F9FH9_0;
	wire w_dff_B_2kSTW6Sd7_1;
	wire w_dff_B_HihNYsOz6_1;
	wire w_dff_B_rwmtQSBt7_1;
	wire w_dff_B_zGrYmkmI8_1;
	wire w_dff_B_C55HPewp1_1;
	wire w_dff_B_ydCb9c8S3_1;
	wire w_dff_B_fZ9qS8y43_1;
	wire w_dff_B_N7wdEcYt6_1;
	wire w_dff_B_vKddPc6J4_0;
	wire w_dff_B_SFgyGw4V0_0;
	wire w_dff_B_A2G2QvTk2_0;
	wire w_dff_B_9Td78AnT3_0;
	wire w_dff_B_RaHIRqRo3_0;
	wire w_dff_B_kXvKi1aH9_0;
	wire w_dff_B_Jh6s40yZ9_0;
	wire w_dff_B_mJs1Nkki5_0;
	wire w_dff_B_OB2obTJX4_1;
	wire w_dff_B_zaoNu5t89_1;
	wire w_dff_B_vrBd0hBk1_1;
	wire w_dff_B_yJ2vPBkx1_1;
	wire w_dff_B_qcTM0oYr3_1;
	wire w_dff_B_hRNmHLjc4_1;
	wire w_dff_B_hLXcHmzy9_1;
	wire w_dff_B_pxoEL8Ao6_0;
	wire w_dff_B_u7GZB3fE3_0;
	wire w_dff_B_VAKcFD7K6_0;
	wire w_dff_B_2mjUAZxI7_0;
	wire w_dff_B_1STAXDoW0_0;
	wire w_dff_B_dTc5u5NJ3_0;
	wire w_dff_B_ct1c3ZgN9_0;
	wire w_dff_B_CHUBRtFA7_1;
	wire w_dff_B_n0X03tB08_1;
	wire w_dff_B_ASNfjgOR3_1;
	wire w_dff_B_GHlrtJBt5_1;
	wire w_dff_B_6Ozoswgv6_1;
	wire w_dff_B_7AXejlE29_1;
	wire w_dff_B_OW2MPfgS2_0;
	wire w_dff_B_8V7YNLIH4_0;
	wire w_dff_B_xLIWOsd62_0;
	wire w_dff_B_pLV3pkIm4_0;
	wire w_dff_B_BxtlValQ7_0;
	wire w_dff_B_jwfquIHg2_0;
	wire w_dff_B_HuqhDjQS5_1;
	wire w_dff_B_IE6E3WZZ4_1;
	wire w_dff_B_sMlnHecV2_1;
	wire w_dff_B_3RzBsZo46_1;
	wire w_dff_B_IAJMsY3O3_1;
	wire w_dff_B_1XUtnL036_0;
	wire w_dff_B_dumKUOU95_0;
	wire w_dff_B_IhzeJ2iA2_0;
	wire w_dff_B_6HLLPz0U0_0;
	wire w_dff_B_D2KL4nNr1_0;
	wire w_dff_B_91yUkRCn4_1;
	wire w_dff_B_fO5HpThl3_1;
	wire w_dff_B_nHghsEwQ6_1;
	wire w_dff_B_9DVgFh9T1_1;
	wire w_dff_B_DBi1JzBL5_0;
	wire w_dff_B_OSgiaOyx3_0;
	wire w_dff_B_jpsm4AHP2_0;
	wire w_dff_B_NsJlHOhQ0_0;
	wire w_dff_B_rrHAuH711_1;
	wire w_dff_B_AAX4DMaO0_1;
	wire w_dff_B_RYyduIeI2_1;
	wire w_dff_B_U5MNQmS86_0;
	wire w_dff_B_6rt9170L4_0;
	wire w_dff_B_tOSk0HiB9_0;
	wire w_dff_B_q4293DRu4_1;
	wire w_dff_B_XC6XIR9e5_1;
	wire w_dff_B_yaQER63f8_0;
	wire w_dff_B_MevlBocM3_0;
	wire w_dff_B_bq66TJJL2_1;
	wire w_dff_B_7v1bBDjM8_0;
	wire w_dff_A_i0Y4neCV3_2;
	wire w_dff_A_j9T031q05_0;
	wire w_dff_A_vOiNMKYP3_0;
	wire w_dff_A_g7jlr3ng4_0;
	wire w_dff_A_7xO2jXg01_0;
	wire w_dff_A_iMKXw20r6_0;
	wire w_dff_A_MsCrJjMJ8_0;
	wire w_dff_A_4vHSuZu70_0;
	wire w_dff_A_WjGq4SrP5_0;
	wire w_dff_A_UD7Fx71E9_0;
	wire w_dff_A_BlG5FfJJ3_0;
	wire w_dff_A_u78ECBzG5_0;
	wire w_dff_A_IjlLUlhH9_0;
	wire w_dff_A_DeVWj5dN4_0;
	wire w_dff_A_NGHM5wy50_0;
	wire w_dff_A_fmaRaMD69_0;
	wire w_dff_A_1QE0PPCo6_0;
	wire w_dff_A_MtM8rSW48_0;
	wire w_dff_A_FVQJGeqJ3_0;
	wire w_dff_A_qyRq3uJQ5_0;
	wire w_dff_A_3jDPCLoI8_0;
	wire w_dff_A_1hGM26PS8_0;
	wire w_dff_A_BsNAX5yA1_0;
	wire w_dff_A_BbLFrTpV2_0;
	wire w_dff_A_Br5jEmCl2_0;
	wire w_dff_A_5cjTzbmW6_0;
	wire w_dff_A_Q4HY9n4w0_0;
	wire w_dff_A_KSDQi7Sr8_0;
	wire w_dff_A_9Esn0sSu7_0;
	wire w_dff_A_NYjX1kI69_0;
	wire w_dff_A_PAv4FYSN4_0;
	wire w_dff_A_fZbm0Pb18_0;
	wire w_dff_A_CpTsBUrx7_0;
	wire w_dff_A_wpibraiv9_0;
	wire w_dff_A_YECaqBxJ3_0;
	wire w_dff_A_YvPcmbAA1_0;
	wire w_dff_A_h1bwGIX91_0;
	wire w_dff_A_mytFLC8s0_0;
	wire w_dff_A_ChQHW2bi6_0;
	wire w_dff_A_Bfpumz2I0_0;
	wire w_dff_A_AQlr7wG59_0;
	wire w_dff_A_p3fLkJ6r9_0;
	wire w_dff_A_FfFHmd7v3_0;
	wire w_dff_A_a5Oc9kr70_0;
	wire w_dff_A_Ra95uvKl2_0;
	wire w_dff_A_wQ78edMl3_0;
	wire w_dff_A_lNWXIFlC6_0;
	wire w_dff_A_EQajtwzB7_0;
	wire w_dff_A_nS0N2j9E4_0;
	wire w_dff_A_F7vrl6TH5_0;
	wire w_dff_A_F82sm3Qg5_0;
	wire w_dff_A_DWlzNtNs3_0;
	wire w_dff_A_lzKWaH0E2_0;
	wire w_dff_A_MdGhRnUY2_0;
	wire w_dff_A_QwkWUQC88_0;
	wire w_dff_A_s16Kjcf04_0;
	wire w_dff_A_8C1R7pBF0_0;
	wire w_dff_A_A698ntck9_0;
	wire w_dff_A_XMpNqoHx8_0;
	wire w_dff_A_mbphToWb7_0;
	wire w_dff_A_h8kgWcfH2_0;
	wire w_dff_A_wdiR9ZbH8_0;
	wire w_dff_A_9aXA21gj8_0;
	wire w_dff_A_dllhdTsZ5_0;
	wire w_dff_A_hkntw2iQ3_0;
	wire w_dff_A_F2R2oWU87_0;
	wire w_dff_A_Yz94n4vv2_0;
	wire w_dff_A_mW3QoIE34_0;
	wire w_dff_A_p0NmxDOf5_0;
	wire w_dff_A_hAjsqHFs7_0;
	wire w_dff_A_XSuWdF6A5_0;
	wire w_dff_A_oU0ETh9J1_0;
	wire w_dff_A_b8zCdsUw4_0;
	wire w_dff_A_tNUiQJeN7_0;
	wire w_dff_A_sBerItzw4_0;
	wire w_dff_A_Ck24AXEd6_0;
	wire w_dff_A_zLwlimAo0_0;
	wire w_dff_A_q7N8tmnv2_0;
	wire w_dff_A_s07mlbpA8_0;
	wire w_dff_A_xN753xVm5_0;
	wire w_dff_A_ltBC9pjb9_0;
	wire w_dff_A_rsthNRDN8_0;
	wire w_dff_A_6VmHlJVB6_0;
	wire w_dff_A_Rd7ZK2f16_0;
	wire w_dff_A_MhIDTrRH2_0;
	wire w_dff_A_2084AwKm7_0;
	wire w_dff_A_dyLYxj1m9_0;
	wire w_dff_A_r76cTSru5_0;
	wire w_dff_A_9upUtRfy7_0;
	wire w_dff_A_R3GFswzi0_0;
	wire w_dff_A_qDpZEltD3_0;
	wire w_dff_A_tQ21VjHR8_0;
	wire w_dff_A_APJkiJjk3_0;
	wire w_dff_A_f0jsEngB0_0;
	wire w_dff_A_bj5kxm8C9_0;
	wire w_dff_A_892gOQmY8_0;
	wire w_dff_A_CXFTnmf38_0;
	wire w_dff_A_n5VIXJVX0_0;
	wire w_dff_A_OvUzNb0a9_0;
	wire w_dff_A_3T7R4z2L7_0;
	wire w_dff_A_6hVGcGjn7_0;
	wire w_dff_A_1bs2MkNT3_0;
	wire w_dff_A_hq1hQlX82_0;
	wire w_dff_A_K6RhxdqK9_0;
	wire w_dff_A_lB4foRKx4_0;
	wire w_dff_A_SyYyACrh3_0;
	wire w_dff_A_vrg7IbP29_0;
	wire w_dff_A_hw9WaR1E0_0;
	wire w_dff_A_FnaEgvJL6_0;
	wire w_dff_A_L5GZFCwL1_0;
	wire w_dff_A_7Ge97Kqv7_0;
	wire w_dff_A_5dlhIaId4_0;
	wire w_dff_A_kAsFlyjP4_0;
	wire w_dff_A_TzGzpJ4C3_0;
	wire w_dff_A_a3hY8lG88_0;
	wire w_dff_A_TtW8gwUa3_0;
	wire w_dff_A_jJJCywzm0_0;
	wire w_dff_A_3anXx5NG1_0;
	wire w_dff_A_LsjfsP1Y6_0;
	wire w_dff_A_crqbojAo4_0;
	wire w_dff_A_jC9vxI7n8_0;
	wire w_dff_A_xxv6f08e9_0;
	wire w_dff_A_IVoLt4XJ3_0;
	wire w_dff_A_vf1lBtKz5_0;
	wire w_dff_A_jWt7kMj01_0;
	wire w_dff_A_LsCziHwc8_0;
	wire w_dff_A_dYHDCUxr5_0;
	wire w_dff_A_0HyOVMXh8_2;
	wire w_dff_A_3G23CtSw0_0;
	wire w_dff_A_0nIw1xIb5_0;
	wire w_dff_A_QYm95bez2_0;
	wire w_dff_A_own2PeE63_0;
	wire w_dff_A_PnCakQKp7_0;
	wire w_dff_A_95eyG7NE0_0;
	wire w_dff_A_j6fh7tBp4_0;
	wire w_dff_A_dCXANpXg1_0;
	wire w_dff_A_6RytlC7I6_0;
	wire w_dff_A_Ai7zWDjI4_0;
	wire w_dff_A_dssNx9xZ2_0;
	wire w_dff_A_X5qBjmyC9_0;
	wire w_dff_A_dXWKlv5p2_0;
	wire w_dff_A_caK9uQfT4_0;
	wire w_dff_A_WgiQCrIh1_0;
	wire w_dff_A_H2n7MluO8_0;
	wire w_dff_A_lzT9a55J2_0;
	wire w_dff_A_ru8uTTJN4_0;
	wire w_dff_A_8iTMwZxx2_0;
	wire w_dff_A_vclqBMNU4_0;
	wire w_dff_A_u65A8I2k2_0;
	wire w_dff_A_40WVdttX2_0;
	wire w_dff_A_vX7CEtcz9_0;
	wire w_dff_A_Sz6NsqZl6_0;
	wire w_dff_A_JBr9KMOI3_0;
	wire w_dff_A_O0W1wJmi4_0;
	wire w_dff_A_chSHBBma5_0;
	wire w_dff_A_tNvW27wX0_0;
	wire w_dff_A_vL2PBhjs8_0;
	wire w_dff_A_Li7ZzbTp0_0;
	wire w_dff_A_CRD7aBrp1_0;
	wire w_dff_A_85BVUYDg4_0;
	wire w_dff_A_Ur617CXp1_0;
	wire w_dff_A_xR42W3dx1_0;
	wire w_dff_A_MUBBZAyu8_0;
	wire w_dff_A_0IqHmckP5_0;
	wire w_dff_A_mtVZU8B56_0;
	wire w_dff_A_yHrDEpg68_0;
	wire w_dff_A_1ED0imto9_0;
	wire w_dff_A_nNi07eYW2_0;
	wire w_dff_A_4Nomh9bM3_0;
	wire w_dff_A_SQNXA9Wl9_0;
	wire w_dff_A_irmpFzn86_0;
	wire w_dff_A_WcITGojs6_0;
	wire w_dff_A_5CVuS75m4_0;
	wire w_dff_A_xgR6y6b96_0;
	wire w_dff_A_UMmVYahG3_0;
	wire w_dff_A_t58Ms7ZG9_0;
	wire w_dff_A_9JTQdnKu9_0;
	wire w_dff_A_noVY6HwB7_0;
	wire w_dff_A_v1rMq7UA9_0;
	wire w_dff_A_WExnmypd3_0;
	wire w_dff_A_RcP08nNg3_0;
	wire w_dff_A_Z179FsCr8_0;
	wire w_dff_A_VOwnRV5i0_0;
	wire w_dff_A_MGRIkIPv5_0;
	wire w_dff_A_B68fX2v50_0;
	wire w_dff_A_KqVPuXUG4_0;
	wire w_dff_A_9whzdQBg6_0;
	wire w_dff_A_Cq0ZoSVK5_0;
	wire w_dff_A_4ihd7n8u0_0;
	wire w_dff_A_uX8FinwS8_0;
	wire w_dff_A_tbCkAZXf3_0;
	wire w_dff_A_L9QagEZF0_0;
	wire w_dff_A_Bd0HKDFY7_0;
	wire w_dff_A_LcE5VPro2_0;
	wire w_dff_A_BCS6BT2t9_0;
	wire w_dff_A_O5mNMmaB9_0;
	wire w_dff_A_aqz37mCq3_0;
	wire w_dff_A_g7eRWlGo3_0;
	wire w_dff_A_Xqb01NrL2_0;
	wire w_dff_A_CLSGyjeC9_0;
	wire w_dff_A_S1Yusywy5_0;
	wire w_dff_A_Sr2E2Dy67_0;
	wire w_dff_A_Juu2DPc14_0;
	wire w_dff_A_sFEwPaDj8_0;
	wire w_dff_A_VzD49Oyz8_0;
	wire w_dff_A_ubPW59ec6_0;
	wire w_dff_A_5rY6TR0a9_0;
	wire w_dff_A_TRIlYsW30_0;
	wire w_dff_A_6KJfzSC90_0;
	wire w_dff_A_dBw8ThP34_0;
	wire w_dff_A_r5IGKeUn0_0;
	wire w_dff_A_Hy53EKJI8_0;
	wire w_dff_A_tpdXvOML4_0;
	wire w_dff_A_va51BmCQ9_0;
	wire w_dff_A_YN7tNNay4_0;
	wire w_dff_A_imQL9fn46_0;
	wire w_dff_A_396hJunk3_0;
	wire w_dff_A_IVgNkzZM8_0;
	wire w_dff_A_QCtLnjdX3_0;
	wire w_dff_A_1m1hyP6z8_0;
	wire w_dff_A_R7HV63Vw0_0;
	wire w_dff_A_TgzLISqZ2_0;
	wire w_dff_A_0NBdKgS54_0;
	wire w_dff_A_19S5qRxr3_0;
	wire w_dff_A_PnlfMz8I5_0;
	wire w_dff_A_EyVPaNEH4_0;
	wire w_dff_A_JLEnT9bs8_0;
	wire w_dff_A_EMfMitW65_0;
	wire w_dff_A_yZ71UeeG4_0;
	wire w_dff_A_bV8uCmZ90_0;
	wire w_dff_A_L75unZ0w2_0;
	wire w_dff_A_V2N1sjSX9_0;
	wire w_dff_A_QEKkZaOf6_0;
	wire w_dff_A_fbbg29LL4_0;
	wire w_dff_A_tmdxY3We9_0;
	wire w_dff_A_Z5AYQiKM9_0;
	wire w_dff_A_RwuSfQ1A3_0;
	wire w_dff_A_xU7Yr7KA6_0;
	wire w_dff_A_GQwdU88m4_0;
	wire w_dff_A_SSoRjrpe6_0;
	wire w_dff_A_Lqcg1Ngn9_0;
	wire w_dff_A_SGLJI8Q25_0;
	wire w_dff_A_WhjorSEl2_0;
	wire w_dff_A_ajTaRkWl7_0;
	wire w_dff_A_GPrw2l8F5_0;
	wire w_dff_A_6f4VSBjy6_0;
	wire w_dff_A_98OqeYdm1_0;
	wire w_dff_A_pFjwNU4X6_0;
	wire w_dff_A_KP3JqESX0_0;
	wire w_dff_A_7m0DZKCr2_0;
	wire w_dff_A_QFuhrs5q5_0;
	wire w_dff_A_V6W5MPpX4_0;
	wire w_dff_A_BhZgMGEA0_0;
	wire w_dff_A_BvD62S921_2;
	wire w_dff_A_gMz6Lb5D8_0;
	wire w_dff_A_yLtN7iw95_0;
	wire w_dff_A_IA3oxORP5_0;
	wire w_dff_A_AUiNijlD2_0;
	wire w_dff_A_zMekuf8x1_0;
	wire w_dff_A_C5IQIOJW6_0;
	wire w_dff_A_j6WANsVL1_0;
	wire w_dff_A_JUMS4rlL9_0;
	wire w_dff_A_b7MWDKxD3_0;
	wire w_dff_A_L0p1xxS55_0;
	wire w_dff_A_QPb7BxDj1_0;
	wire w_dff_A_zQBw3Rtn4_0;
	wire w_dff_A_La4d9nsL1_0;
	wire w_dff_A_FhHZAgEC8_0;
	wire w_dff_A_m1qLRZr12_0;
	wire w_dff_A_AOAbQvcI2_0;
	wire w_dff_A_0frBFz460_0;
	wire w_dff_A_FZdDIpnV1_0;
	wire w_dff_A_pcJmtdQc1_0;
	wire w_dff_A_hi8IlDSj0_0;
	wire w_dff_A_6eUrlbcC0_0;
	wire w_dff_A_CiCKQe8J9_0;
	wire w_dff_A_uwkglmLH0_0;
	wire w_dff_A_Fxxmc7iO8_0;
	wire w_dff_A_F57YYRhM2_0;
	wire w_dff_A_ChVRGd0L0_0;
	wire w_dff_A_7IDO9qf89_0;
	wire w_dff_A_34iojwkP1_0;
	wire w_dff_A_DUHIAmDv9_0;
	wire w_dff_A_sDpan7jS9_0;
	wire w_dff_A_WVVgc9Sf9_0;
	wire w_dff_A_53N0H0zX5_0;
	wire w_dff_A_6MXTdlQ91_0;
	wire w_dff_A_C97PlHyO2_0;
	wire w_dff_A_tLb5D9S65_0;
	wire w_dff_A_t7G32yOC5_0;
	wire w_dff_A_H54wYtCl3_0;
	wire w_dff_A_XfdL9HlW6_0;
	wire w_dff_A_pIdsk8F65_0;
	wire w_dff_A_ZMs4jKWp8_0;
	wire w_dff_A_nkNIQKSY4_0;
	wire w_dff_A_0Fk5wTtC2_0;
	wire w_dff_A_o4DQiZVa7_0;
	wire w_dff_A_h1Jt0UWn1_0;
	wire w_dff_A_GCnye3ZX9_0;
	wire w_dff_A_7NPpwmKi3_0;
	wire w_dff_A_cfpTaVgI3_0;
	wire w_dff_A_ZAB4PPed8_0;
	wire w_dff_A_EJeNXIFi1_0;
	wire w_dff_A_X1nkO6wo0_0;
	wire w_dff_A_1RnWr8J29_0;
	wire w_dff_A_nDsazNLQ9_0;
	wire w_dff_A_3nqhLmj45_0;
	wire w_dff_A_bN1SHJC38_0;
	wire w_dff_A_zME2Tpf04_0;
	wire w_dff_A_7k56kaHd7_0;
	wire w_dff_A_1hCIaHIB3_0;
	wire w_dff_A_yngkKjXy7_0;
	wire w_dff_A_xMFeIU907_0;
	wire w_dff_A_HcXcIV3N6_0;
	wire w_dff_A_fR0Ob4G44_0;
	wire w_dff_A_2ykFKu2t5_0;
	wire w_dff_A_jm9LYl8C6_0;
	wire w_dff_A_tUp7NdTr2_0;
	wire w_dff_A_bwTsA3Q15_0;
	wire w_dff_A_eXAvG3xU4_0;
	wire w_dff_A_KDyacK611_0;
	wire w_dff_A_jPiwoq8Q8_0;
	wire w_dff_A_fGDojP762_0;
	wire w_dff_A_VyoFmQkw5_0;
	wire w_dff_A_T8khXwxt6_0;
	wire w_dff_A_K73VURR94_0;
	wire w_dff_A_EUMWAIkn3_0;
	wire w_dff_A_WEXHHw9z4_0;
	wire w_dff_A_eazaBLVO4_0;
	wire w_dff_A_rjirzV5f0_0;
	wire w_dff_A_Czdqyu6Y0_0;
	wire w_dff_A_Z1Laxp9i4_0;
	wire w_dff_A_15Gtg2h36_0;
	wire w_dff_A_QpFTH8B80_0;
	wire w_dff_A_V9QrQztm9_0;
	wire w_dff_A_qRYXWz9X8_0;
	wire w_dff_A_xFtAuA2J5_0;
	wire w_dff_A_fmsyS0um0_0;
	wire w_dff_A_m9HoNS8u7_0;
	wire w_dff_A_YY7pLLwB6_0;
	wire w_dff_A_pkQtA9eJ2_0;
	wire w_dff_A_PCclndeQ9_0;
	wire w_dff_A_4kthRXsq7_0;
	wire w_dff_A_kNM1InUm8_0;
	wire w_dff_A_5LvdS70S0_0;
	wire w_dff_A_pK93onTu3_0;
	wire w_dff_A_YX6yAdRf8_0;
	wire w_dff_A_rckmqZmE9_0;
	wire w_dff_A_dZJDu4xZ9_0;
	wire w_dff_A_0jpG0GS89_0;
	wire w_dff_A_93fubIHx8_0;
	wire w_dff_A_IuzcCOiA7_0;
	wire w_dff_A_ISeyzKuN8_0;
	wire w_dff_A_grOGOaF14_0;
	wire w_dff_A_ZzJuS0Wi2_0;
	wire w_dff_A_bPAKUw0p5_0;
	wire w_dff_A_VNSZvRpl0_0;
	wire w_dff_A_ab6HyjvL7_0;
	wire w_dff_A_95N8oCST4_0;
	wire w_dff_A_kDxktsP28_0;
	wire w_dff_A_k9lIUXm30_0;
	wire w_dff_A_jpGpTGH53_0;
	wire w_dff_A_57lRtJJu5_0;
	wire w_dff_A_ozZC3i9t3_0;
	wire w_dff_A_FL5FHqTE2_0;
	wire w_dff_A_ou4I5wYa1_0;
	wire w_dff_A_4lFlDF7p6_0;
	wire w_dff_A_bxIXJpTJ0_0;
	wire w_dff_A_gTy9ccLO5_0;
	wire w_dff_A_xDWTr75G7_0;
	wire w_dff_A_MV3cRGsb8_0;
	wire w_dff_A_plKD2YaN9_0;
	wire w_dff_A_5a8Is8P98_0;
	wire w_dff_A_ZQfeTGbs4_0;
	wire w_dff_A_xLY0Q4XN2_0;
	wire w_dff_A_25MA11i46_0;
	wire w_dff_A_P1xX5SoN3_0;
	wire w_dff_A_qRlywRaA1_0;
	wire w_dff_A_lRUw1Ruu2_2;
	wire w_dff_A_La1LKto64_0;
	wire w_dff_A_bdp3MxDE8_0;
	wire w_dff_A_WqgofUlT6_0;
	wire w_dff_A_HURVWnDK0_0;
	wire w_dff_A_tE3EP4Gv0_0;
	wire w_dff_A_aq0xns4Z7_0;
	wire w_dff_A_3nR77eZh3_0;
	wire w_dff_A_Ah14sbfU8_0;
	wire w_dff_A_1WcRL1Tj4_0;
	wire w_dff_A_ONCu3cv30_0;
	wire w_dff_A_KDg5tI2k3_0;
	wire w_dff_A_235zJRRa7_0;
	wire w_dff_A_aOiZ6Bzx1_0;
	wire w_dff_A_FChoMAaX2_0;
	wire w_dff_A_pCtOXO764_0;
	wire w_dff_A_0h8zISNG9_0;
	wire w_dff_A_fF46Ozse3_0;
	wire w_dff_A_gi1fmzJE6_0;
	wire w_dff_A_gaqTL2bo9_0;
	wire w_dff_A_Ax5bWosD2_0;
	wire w_dff_A_ctSG34BC7_0;
	wire w_dff_A_IaQmkzvh0_0;
	wire w_dff_A_rgU0Bqgn6_0;
	wire w_dff_A_hqA5agcV1_0;
	wire w_dff_A_h3XBLhf63_0;
	wire w_dff_A_G2k3SXBg8_0;
	wire w_dff_A_3GpCjouF8_0;
	wire w_dff_A_yHuxXgw80_0;
	wire w_dff_A_RRLV3ErP9_0;
	wire w_dff_A_zj0CkmKh7_0;
	wire w_dff_A_lem8Aolv3_0;
	wire w_dff_A_6Vmug3QF6_0;
	wire w_dff_A_fDNILKEJ8_0;
	wire w_dff_A_9lTlUCnX7_0;
	wire w_dff_A_24lpbOJf9_0;
	wire w_dff_A_kbYCQ5jM7_0;
	wire w_dff_A_Utn0vbNx7_0;
	wire w_dff_A_ik0m86LA5_0;
	wire w_dff_A_0bcUWQKt5_0;
	wire w_dff_A_MiWzcOCo6_0;
	wire w_dff_A_o6g47jgN2_0;
	wire w_dff_A_Ojr2sefc3_0;
	wire w_dff_A_fpXtYxcH7_0;
	wire w_dff_A_tzuzDKzW6_0;
	wire w_dff_A_REThOIV03_0;
	wire w_dff_A_nssv3Qjd3_0;
	wire w_dff_A_9zVim3YN2_0;
	wire w_dff_A_NzYZyxNE7_0;
	wire w_dff_A_zwYNBsE24_0;
	wire w_dff_A_hAQEzWNP0_0;
	wire w_dff_A_8fjYSDN06_0;
	wire w_dff_A_8nW0GRpX9_0;
	wire w_dff_A_BMshOraN6_0;
	wire w_dff_A_0N8IAiOv9_0;
	wire w_dff_A_hahuCbq42_0;
	wire w_dff_A_6ykzNZKe3_0;
	wire w_dff_A_INdv5qFp5_0;
	wire w_dff_A_duTSnfOO7_0;
	wire w_dff_A_nwTJnMl86_0;
	wire w_dff_A_V6AQytRS5_0;
	wire w_dff_A_Hl27t9hM6_0;
	wire w_dff_A_dRyg1Mam4_0;
	wire w_dff_A_6FlbFwlC6_0;
	wire w_dff_A_v13qb5nq7_0;
	wire w_dff_A_c6hh5IUo6_0;
	wire w_dff_A_hbFtzmBo3_0;
	wire w_dff_A_kxGQXqtr9_0;
	wire w_dff_A_JDnZjqQp7_0;
	wire w_dff_A_fKgz4nob1_0;
	wire w_dff_A_KkpAdIZ04_0;
	wire w_dff_A_b6SKdcWb7_0;
	wire w_dff_A_i3payFii8_0;
	wire w_dff_A_R6ME8LkR2_0;
	wire w_dff_A_vHWmL4bY5_0;
	wire w_dff_A_fxuGvgar1_0;
	wire w_dff_A_monQdnWv6_0;
	wire w_dff_A_vYhJ3o3P3_0;
	wire w_dff_A_qOYDpDCm0_0;
	wire w_dff_A_PcI56gSH0_0;
	wire w_dff_A_L7RLkWpq5_0;
	wire w_dff_A_APOk7nlo8_0;
	wire w_dff_A_V8oT1Aak0_0;
	wire w_dff_A_6Wo7BBeT1_0;
	wire w_dff_A_AVszMIfw3_0;
	wire w_dff_A_ndAAfpjO1_0;
	wire w_dff_A_MycMRMU68_0;
	wire w_dff_A_o6KCc00R9_0;
	wire w_dff_A_ElfwmsAm5_0;
	wire w_dff_A_QncfXZiP9_0;
	wire w_dff_A_cFHV3YQ45_0;
	wire w_dff_A_OTrGdUVH8_0;
	wire w_dff_A_N2ERbr8I4_0;
	wire w_dff_A_ZIs4rbFq8_0;
	wire w_dff_A_AZUEEfxO7_0;
	wire w_dff_A_iLufhf6o8_0;
	wire w_dff_A_MyMyPt571_0;
	wire w_dff_A_tRzYee8n4_0;
	wire w_dff_A_iYOAAS3t5_0;
	wire w_dff_A_B8MDTUpb8_0;
	wire w_dff_A_IfozyU0f6_0;
	wire w_dff_A_TeAQgpvl3_0;
	wire w_dff_A_N8imk39S0_0;
	wire w_dff_A_SFT6a6JL3_0;
	wire w_dff_A_z2m4hU9P3_0;
	wire w_dff_A_zfpi0cDF6_0;
	wire w_dff_A_vG7Wtfqb2_0;
	wire w_dff_A_Q6MQmU7a3_0;
	wire w_dff_A_kqxinkmM3_0;
	wire w_dff_A_27Y7HHIo6_0;
	wire w_dff_A_GxAGMbpU9_0;
	wire w_dff_A_6mZaMQ2u8_0;
	wire w_dff_A_OPV7AuyA9_0;
	wire w_dff_A_Mvev92x47_0;
	wire w_dff_A_FSH3reNl4_0;
	wire w_dff_A_LxDiXIh96_0;
	wire w_dff_A_mRkKIUyw0_0;
	wire w_dff_A_4heoCdeK5_0;
	wire w_dff_A_NrVXIPUz6_0;
	wire w_dff_A_yDjtFI9Y3_0;
	wire w_dff_A_1Bt2Y9695_0;
	wire w_dff_A_U3ZrDMSm2_0;
	wire w_dff_A_9yc2b15b4_0;
	wire w_dff_A_6mwv8tLa6_0;
	wire w_dff_A_1VQG7qnR4_2;
	wire w_dff_A_5Fa9cNUP9_0;
	wire w_dff_A_XszYuBZn6_0;
	wire w_dff_A_rYDI6ieU0_0;
	wire w_dff_A_Mb7TeTvB7_0;
	wire w_dff_A_7oPnku5t2_0;
	wire w_dff_A_zXBJKvOz5_0;
	wire w_dff_A_L0Frk5Ii6_0;
	wire w_dff_A_uumZ1lpo8_0;
	wire w_dff_A_7xBWhwoN9_0;
	wire w_dff_A_ZkF2pzgP4_0;
	wire w_dff_A_iNMcl5751_0;
	wire w_dff_A_25m6uuBK2_0;
	wire w_dff_A_jH9p5tME8_0;
	wire w_dff_A_FoMYKH7m5_0;
	wire w_dff_A_QMiARZyX8_0;
	wire w_dff_A_5a6wVnjT2_0;
	wire w_dff_A_HjFceiDg1_0;
	wire w_dff_A_77u0j4Uq4_0;
	wire w_dff_A_sICGys189_0;
	wire w_dff_A_8WD7kccW5_0;
	wire w_dff_A_XPVG3QX59_0;
	wire w_dff_A_5xDpoGie3_0;
	wire w_dff_A_fDdvouAS8_0;
	wire w_dff_A_CX8XH9k80_0;
	wire w_dff_A_wWsff6kH7_0;
	wire w_dff_A_tyOQC1gb4_0;
	wire w_dff_A_JOM0hDP27_0;
	wire w_dff_A_VxOcX4fM4_0;
	wire w_dff_A_9XJ5I31a5_0;
	wire w_dff_A_vNiNP8Ud7_0;
	wire w_dff_A_iFD7q3yd1_0;
	wire w_dff_A_9lFpBAUQ4_0;
	wire w_dff_A_j4kMoJ2N8_0;
	wire w_dff_A_koYqHtAr5_0;
	wire w_dff_A_j6EMyffI1_0;
	wire w_dff_A_deUhHxrn3_0;
	wire w_dff_A_iYXB5tPh6_0;
	wire w_dff_A_jRDIlC7w5_0;
	wire w_dff_A_X1yj2HMP6_0;
	wire w_dff_A_J0VsU88V9_0;
	wire w_dff_A_UJPKrkUT0_0;
	wire w_dff_A_l0OsOiUk9_0;
	wire w_dff_A_Y7gaWkRM9_0;
	wire w_dff_A_XgrdThwL7_0;
	wire w_dff_A_zukOVIFp0_0;
	wire w_dff_A_aMkd7sWD0_0;
	wire w_dff_A_ynriJyoJ2_0;
	wire w_dff_A_JselGAOv0_0;
	wire w_dff_A_dhQ5W5hO5_0;
	wire w_dff_A_3fFDjsAL8_0;
	wire w_dff_A_2KmSNbko8_0;
	wire w_dff_A_2ubffZrC5_0;
	wire w_dff_A_b2XEM6J21_0;
	wire w_dff_A_lqauPCNQ4_0;
	wire w_dff_A_RLWv6Flx1_0;
	wire w_dff_A_ZUVhd7L38_0;
	wire w_dff_A_IejkbUIe2_0;
	wire w_dff_A_wIRfZAe26_0;
	wire w_dff_A_IzkQeg2s2_0;
	wire w_dff_A_N9cHApKK5_0;
	wire w_dff_A_IhvCVoOx3_0;
	wire w_dff_A_rWO4psWV7_0;
	wire w_dff_A_mgZclAPZ3_0;
	wire w_dff_A_y43MHAER3_0;
	wire w_dff_A_cnBx4Qn79_0;
	wire w_dff_A_6upFUy2T4_0;
	wire w_dff_A_ab4oi3PL5_0;
	wire w_dff_A_No1HjYZc6_0;
	wire w_dff_A_BrZnQq3L7_0;
	wire w_dff_A_NyZpidZa7_0;
	wire w_dff_A_PZvrJR4n4_0;
	wire w_dff_A_TzN4dReA4_0;
	wire w_dff_A_HFSgiQ2O8_0;
	wire w_dff_A_Rk5annqX2_0;
	wire w_dff_A_MThSq39d1_0;
	wire w_dff_A_loObXrDX8_0;
	wire w_dff_A_Re12mYPe0_0;
	wire w_dff_A_sbmHq4qd3_0;
	wire w_dff_A_GacHLWK03_0;
	wire w_dff_A_Rqd5EoRH3_0;
	wire w_dff_A_VRTcxhZo9_0;
	wire w_dff_A_mXfj60WY4_0;
	wire w_dff_A_AGYcJ9yt6_0;
	wire w_dff_A_g5sCEzc00_0;
	wire w_dff_A_662Q5HJj8_0;
	wire w_dff_A_wMkIaqNk1_0;
	wire w_dff_A_pYKCuL1D1_0;
	wire w_dff_A_OtkchGOg2_0;
	wire w_dff_A_GteGHVar9_0;
	wire w_dff_A_ewLSiq3B8_0;
	wire w_dff_A_DBsiDWtA6_0;
	wire w_dff_A_x2X0pvH39_0;
	wire w_dff_A_y1iJf8Sb3_0;
	wire w_dff_A_J9sa2Ghz4_0;
	wire w_dff_A_SVoKgd9P2_0;
	wire w_dff_A_h3Bnk4hO7_0;
	wire w_dff_A_mBo9V4g62_0;
	wire w_dff_A_eEd3ROE53_0;
	wire w_dff_A_yZK3LxT81_0;
	wire w_dff_A_JXfeZ7db4_0;
	wire w_dff_A_Xb6kUgQI5_0;
	wire w_dff_A_WL7gqoW80_0;
	wire w_dff_A_e8WV26aU0_0;
	wire w_dff_A_00jNVlvt5_0;
	wire w_dff_A_GUGBYtzZ5_0;
	wire w_dff_A_i41Ga4qU9_0;
	wire w_dff_A_XBBCXx695_0;
	wire w_dff_A_Qe5cWNkw4_0;
	wire w_dff_A_6Flh009Z9_0;
	wire w_dff_A_E4APkXAG5_0;
	wire w_dff_A_asgeTDbE9_0;
	wire w_dff_A_UxgsX2GP6_0;
	wire w_dff_A_ZT6miqI60_0;
	wire w_dff_A_aSIs1bdk3_0;
	wire w_dff_A_MV6fgJqE2_0;
	wire w_dff_A_0JsU6p5D3_0;
	wire w_dff_A_t2Ktl2Mx2_0;
	wire w_dff_A_MM7DwEUX2_0;
	wire w_dff_A_THFzVDnS6_0;
	wire w_dff_A_3Qz4fLsn5_0;
	wire w_dff_A_Q0j0c46J3_0;
	wire w_dff_A_IuqKgyK03_0;
	wire w_dff_A_IdkFl4Xp4_2;
	wire w_dff_A_7WOSKiuK6_0;
	wire w_dff_A_whqaaO4I3_0;
	wire w_dff_A_dWZmbI9c4_0;
	wire w_dff_A_cLSxEBWv5_0;
	wire w_dff_A_js64y1LC4_0;
	wire w_dff_A_LmWZIKY74_0;
	wire w_dff_A_0lvHdkUq6_0;
	wire w_dff_A_k1VAt9Tt4_0;
	wire w_dff_A_68DsUUIw2_0;
	wire w_dff_A_ZZVkgg8w2_0;
	wire w_dff_A_FYyBu26T7_0;
	wire w_dff_A_6ZGFAdw08_0;
	wire w_dff_A_FYqQvUoA1_0;
	wire w_dff_A_NI6BFi2u9_0;
	wire w_dff_A_M1XSP2in8_0;
	wire w_dff_A_CkbEmAKk1_0;
	wire w_dff_A_Wtm3Bdwb3_0;
	wire w_dff_A_4RlHqDPm5_0;
	wire w_dff_A_WCIIhXIK5_0;
	wire w_dff_A_mzThEMH35_0;
	wire w_dff_A_RdHcBSkH5_0;
	wire w_dff_A_dCB1WaR64_0;
	wire w_dff_A_KuwRXycy1_0;
	wire w_dff_A_ydza07DE2_0;
	wire w_dff_A_imZOv0kF7_0;
	wire w_dff_A_2j8Kcy691_0;
	wire w_dff_A_FaqfAlgy0_0;
	wire w_dff_A_YggbqMBl2_0;
	wire w_dff_A_8kmZQxlg9_0;
	wire w_dff_A_AmeYctPz0_0;
	wire w_dff_A_BCkLTDGX2_0;
	wire w_dff_A_wn8ICb4d3_0;
	wire w_dff_A_0DNGrGX60_0;
	wire w_dff_A_KkoH3SFT0_0;
	wire w_dff_A_K0V2sZl95_0;
	wire w_dff_A_b64RPAkx2_0;
	wire w_dff_A_i8Bw4ziX8_0;
	wire w_dff_A_LynwnBL54_0;
	wire w_dff_A_pbUMnuaJ6_0;
	wire w_dff_A_eenawJlp6_0;
	wire w_dff_A_h68K7PFM5_0;
	wire w_dff_A_MM1znDoQ2_0;
	wire w_dff_A_wQnt1osF4_0;
	wire w_dff_A_jBqP9Rno1_0;
	wire w_dff_A_6SPblfPN8_0;
	wire w_dff_A_Q4FfvqYs8_0;
	wire w_dff_A_MdaOHuhM2_0;
	wire w_dff_A_yT3Zyqar2_0;
	wire w_dff_A_JBeftkVZ9_0;
	wire w_dff_A_80DNT7ja4_0;
	wire w_dff_A_aYGx0Sx09_0;
	wire w_dff_A_Za84DtOn4_0;
	wire w_dff_A_CAfnn6Ln6_0;
	wire w_dff_A_iX3mfOFH4_0;
	wire w_dff_A_GIAv927z8_0;
	wire w_dff_A_GJeHbi3J5_0;
	wire w_dff_A_AVEVBteC2_0;
	wire w_dff_A_3owZC4ri1_0;
	wire w_dff_A_fsC9gKLw2_0;
	wire w_dff_A_EWpfq3hw8_0;
	wire w_dff_A_qk84iQld3_0;
	wire w_dff_A_Wu21gRUj5_0;
	wire w_dff_A_0GjjQOdK3_0;
	wire w_dff_A_ug4j69FI0_0;
	wire w_dff_A_fCZfGh1d4_0;
	wire w_dff_A_NWCLG5AO6_0;
	wire w_dff_A_2ktIlevG8_0;
	wire w_dff_A_ueVTdPtx1_0;
	wire w_dff_A_LSNEDSnm8_0;
	wire w_dff_A_5xGXelTX6_0;
	wire w_dff_A_bghyKuUI2_0;
	wire w_dff_A_E2i1ybhL0_0;
	wire w_dff_A_EK1Gfz8W8_0;
	wire w_dff_A_uLktFuWB3_0;
	wire w_dff_A_MAndBeXK5_0;
	wire w_dff_A_yYgzJu3u3_0;
	wire w_dff_A_wqBpYfAS3_0;
	wire w_dff_A_Yj1onD7G7_0;
	wire w_dff_A_jkjdi0Vl0_0;
	wire w_dff_A_KIVEmHgf9_0;
	wire w_dff_A_386dJLEL3_0;
	wire w_dff_A_sHLcL5qa6_0;
	wire w_dff_A_24Glr9AA7_0;
	wire w_dff_A_v1VNd8VQ7_0;
	wire w_dff_A_nvOXj3F57_0;
	wire w_dff_A_NTJ7VvsC7_0;
	wire w_dff_A_CQN2ArvX2_0;
	wire w_dff_A_U0yJrItQ5_0;
	wire w_dff_A_rBEuEehq5_0;
	wire w_dff_A_fn0Ukzzx7_0;
	wire w_dff_A_NUOEiGJw3_0;
	wire w_dff_A_vNswGoVS3_0;
	wire w_dff_A_Cg96wRru5_0;
	wire w_dff_A_36QFqgDz7_0;
	wire w_dff_A_RGa31G8G5_0;
	wire w_dff_A_YCPseZMm8_0;
	wire w_dff_A_UvlBsSF25_0;
	wire w_dff_A_kpiZTyzw1_0;
	wire w_dff_A_ayqQ7A1i2_0;
	wire w_dff_A_NjUHC57B1_0;
	wire w_dff_A_r2mKJ7wF9_0;
	wire w_dff_A_57AD0IWV2_0;
	wire w_dff_A_6P8UH6uW9_0;
	wire w_dff_A_60bRszFd5_0;
	wire w_dff_A_8sKKRmnR2_0;
	wire w_dff_A_xV2v85oK2_0;
	wire w_dff_A_DvCj09hQ3_0;
	wire w_dff_A_I1weYQuB4_0;
	wire w_dff_A_q27U2D9o8_0;
	wire w_dff_A_yPvM6QNu6_0;
	wire w_dff_A_lvQAJwyq8_0;
	wire w_dff_A_uIAXNmT81_0;
	wire w_dff_A_oHDaYBC27_0;
	wire w_dff_A_4WTwgyoU7_0;
	wire w_dff_A_dz8QVQCV4_0;
	wire w_dff_A_Id0BBLu50_0;
	wire w_dff_A_Yi8Wyf0m3_0;
	wire w_dff_A_ZDKNtDlh6_0;
	wire w_dff_A_F2IbXNIW0_0;
	wire w_dff_A_u8FpD4uR5_0;
	wire w_dff_A_9oP0trCv0_0;
	wire w_dff_A_IFRtoXuS7_2;
	wire w_dff_A_dNM5ioeY8_0;
	wire w_dff_A_0ygzNt811_0;
	wire w_dff_A_EedsJ0zS4_0;
	wire w_dff_A_nR94jSnj8_0;
	wire w_dff_A_eXjQiPQt7_0;
	wire w_dff_A_OfoPCtRU5_0;
	wire w_dff_A_1HGnTNNH6_0;
	wire w_dff_A_H0D9fyRI8_0;
	wire w_dff_A_O8ywRI6V9_0;
	wire w_dff_A_2puUNEVy8_0;
	wire w_dff_A_e63m2zQL1_0;
	wire w_dff_A_x7oyIXNW4_0;
	wire w_dff_A_8k4OgaXM9_0;
	wire w_dff_A_GQZndfBN9_0;
	wire w_dff_A_78akKty68_0;
	wire w_dff_A_jDohhRzZ7_0;
	wire w_dff_A_sigLi1SZ7_0;
	wire w_dff_A_KyI08DTP9_0;
	wire w_dff_A_ay1uCFuY0_0;
	wire w_dff_A_PTBc4VHW4_0;
	wire w_dff_A_UhzCJEAI6_0;
	wire w_dff_A_wZntfqmn0_0;
	wire w_dff_A_QiAw9Cso6_0;
	wire w_dff_A_I2m3H2mn7_0;
	wire w_dff_A_qb9nrwjr8_0;
	wire w_dff_A_vxNMFwka9_0;
	wire w_dff_A_lv50pEPm8_0;
	wire w_dff_A_QNnuq1g22_0;
	wire w_dff_A_Qdj1UiX54_0;
	wire w_dff_A_iUDjuwIf4_0;
	wire w_dff_A_sRzHDofR2_0;
	wire w_dff_A_lXIBZskz4_0;
	wire w_dff_A_ieKkynYu2_0;
	wire w_dff_A_GqLd6dGd4_0;
	wire w_dff_A_yNASuVxS7_0;
	wire w_dff_A_mpq0EkWt2_0;
	wire w_dff_A_PzDfoN9w7_0;
	wire w_dff_A_79FKcPhC3_0;
	wire w_dff_A_aAE1O8N46_0;
	wire w_dff_A_mL4QLLKf1_0;
	wire w_dff_A_8nu04Mvj3_0;
	wire w_dff_A_dKUoN67J0_0;
	wire w_dff_A_PWoB4sES5_0;
	wire w_dff_A_SSWeRzZ21_0;
	wire w_dff_A_jUfcUwEM8_0;
	wire w_dff_A_dIno3LGr7_0;
	wire w_dff_A_lLTkimK53_0;
	wire w_dff_A_nDAF2WLG0_0;
	wire w_dff_A_H1RYwhUX7_0;
	wire w_dff_A_zREFLy8k6_0;
	wire w_dff_A_KFr37E3a6_0;
	wire w_dff_A_UUGkqhtd8_0;
	wire w_dff_A_bKg73B4J5_0;
	wire w_dff_A_cT9CC3GP3_0;
	wire w_dff_A_w2BcjzP62_0;
	wire w_dff_A_uSPJcw9i8_0;
	wire w_dff_A_UmoshPVG6_0;
	wire w_dff_A_SjfTFShX6_0;
	wire w_dff_A_PtLRR8HG1_0;
	wire w_dff_A_sJrkBDuJ7_0;
	wire w_dff_A_6ggOcCn26_0;
	wire w_dff_A_AENC41aY6_0;
	wire w_dff_A_4UL4ueNJ7_0;
	wire w_dff_A_dk8ZWBl44_0;
	wire w_dff_A_7wjnj2BV3_0;
	wire w_dff_A_phvBqXQN8_0;
	wire w_dff_A_xgz9OHjq8_0;
	wire w_dff_A_3npU9qCm6_0;
	wire w_dff_A_8MquYxoq7_0;
	wire w_dff_A_pRYTgd5Y3_0;
	wire w_dff_A_QSxdLCdb2_0;
	wire w_dff_A_0JuxbPDB7_0;
	wire w_dff_A_lZSBKMYh7_0;
	wire w_dff_A_UvC2xjUo2_0;
	wire w_dff_A_xceiiTia7_0;
	wire w_dff_A_cto6lBMf8_0;
	wire w_dff_A_hzLgh0216_0;
	wire w_dff_A_pQLE9Es92_0;
	wire w_dff_A_8xlRWhvp6_0;
	wire w_dff_A_3V3HZntB9_0;
	wire w_dff_A_F5KFFyef7_0;
	wire w_dff_A_go6OBVaW8_0;
	wire w_dff_A_RX5tRT9m0_0;
	wire w_dff_A_Be4yMm239_0;
	wire w_dff_A_uOdvJjvm4_0;
	wire w_dff_A_42nriZNs1_0;
	wire w_dff_A_ppgYe0Kr6_0;
	wire w_dff_A_otdmyLKD7_0;
	wire w_dff_A_rWF4A0gh4_0;
	wire w_dff_A_UwWgvn8a0_0;
	wire w_dff_A_w2czANKh2_0;
	wire w_dff_A_CJ26oO9q6_0;
	wire w_dff_A_jpbqLsyl6_0;
	wire w_dff_A_bHTNkRPH6_0;
	wire w_dff_A_tnzXvyKY8_0;
	wire w_dff_A_TSwnZtYR1_0;
	wire w_dff_A_q8ytKrrd2_0;
	wire w_dff_A_Ue1GZ5cq5_0;
	wire w_dff_A_Ywq21yhK5_0;
	wire w_dff_A_xG9KR7KU8_0;
	wire w_dff_A_lVxRtu1v4_0;
	wire w_dff_A_TZjE7A617_0;
	wire w_dff_A_hPOK1ZsB9_0;
	wire w_dff_A_4j3yS4H37_0;
	wire w_dff_A_TluW0DJW4_0;
	wire w_dff_A_GnHab2jC0_0;
	wire w_dff_A_RfhKmTB59_0;
	wire w_dff_A_UJYzzDkr1_0;
	wire w_dff_A_925rrjgO8_0;
	wire w_dff_A_a1tI1IAw9_0;
	wire w_dff_A_EWxKoSIP0_0;
	wire w_dff_A_t1uDvSzH4_0;
	wire w_dff_A_yyWyHS926_0;
	wire w_dff_A_Wdkx0ujD7_0;
	wire w_dff_A_TYoTy2uZ8_0;
	wire w_dff_A_ZmqUekGv8_0;
	wire w_dff_A_PCLwuSUy5_0;
	wire w_dff_A_iGyCGKtU5_0;
	wire w_dff_A_hnlozL1W4_0;
	wire w_dff_A_yaVjxPvn7_0;
	wire w_dff_A_sGoHlvcX8_2;
	wire w_dff_A_4W6QZxc78_0;
	wire w_dff_A_egHFEAyw0_0;
	wire w_dff_A_xQncDKc42_0;
	wire w_dff_A_g4eQNZOc3_0;
	wire w_dff_A_hOLSdc635_0;
	wire w_dff_A_fqYRsZHI8_0;
	wire w_dff_A_Jb19i3wQ9_0;
	wire w_dff_A_kYfU3JQz5_0;
	wire w_dff_A_8gRy1Co38_0;
	wire w_dff_A_lVyFbCZS6_0;
	wire w_dff_A_KQxBJq8i3_0;
	wire w_dff_A_dj9Kq0th5_0;
	wire w_dff_A_kCgK3GXG1_0;
	wire w_dff_A_U1RU7iWf1_0;
	wire w_dff_A_Q8udJ7bo7_0;
	wire w_dff_A_nkJA41tR4_0;
	wire w_dff_A_8HcvDrca6_0;
	wire w_dff_A_ydAZef970_0;
	wire w_dff_A_P6LCG2DZ0_0;
	wire w_dff_A_nLTMRlbh1_0;
	wire w_dff_A_n3ZpOXDP8_0;
	wire w_dff_A_VdA4E3q73_0;
	wire w_dff_A_eBOsIbtN9_0;
	wire w_dff_A_sRNozZAn6_0;
	wire w_dff_A_SHwXN1RT1_0;
	wire w_dff_A_cFyh7PrA6_0;
	wire w_dff_A_VskicEZp3_0;
	wire w_dff_A_IfunqZdA5_0;
	wire w_dff_A_2RpfZK663_0;
	wire w_dff_A_ZbZntsYK3_0;
	wire w_dff_A_v5ncrlI21_0;
	wire w_dff_A_4eNYktAA3_0;
	wire w_dff_A_un74S38m7_0;
	wire w_dff_A_zM36sHxC7_0;
	wire w_dff_A_nCJAiT6V4_0;
	wire w_dff_A_1mMAkSBq5_0;
	wire w_dff_A_qkvT121X8_0;
	wire w_dff_A_JMf8sMHM2_0;
	wire w_dff_A_93Ktuyfd4_0;
	wire w_dff_A_r1GFEXQe4_0;
	wire w_dff_A_6yJ42Ukp5_0;
	wire w_dff_A_iNarG90M1_0;
	wire w_dff_A_N3XvRgar4_0;
	wire w_dff_A_XsHZS8VK4_0;
	wire w_dff_A_0Cz0pDGs1_0;
	wire w_dff_A_1Wr2h8cN8_0;
	wire w_dff_A_xRp3GTiY1_0;
	wire w_dff_A_eHpDtK417_0;
	wire w_dff_A_ZVNAuxVq1_0;
	wire w_dff_A_UO38ASv10_0;
	wire w_dff_A_bB9O1liK7_0;
	wire w_dff_A_lXbVM0Hc0_0;
	wire w_dff_A_AFab10RQ2_0;
	wire w_dff_A_ZwNktAb33_0;
	wire w_dff_A_sczRJfeQ8_0;
	wire w_dff_A_ljBd9yWV3_0;
	wire w_dff_A_6EPYn6hh2_0;
	wire w_dff_A_sEQHXFxK6_0;
	wire w_dff_A_9BSO4exH9_0;
	wire w_dff_A_g06sEK4S9_0;
	wire w_dff_A_YTQR9xzP1_0;
	wire w_dff_A_zwNUoZ8I6_0;
	wire w_dff_A_OwqRkI7r5_0;
	wire w_dff_A_Xi4fSevg6_0;
	wire w_dff_A_SEvnLM3O7_0;
	wire w_dff_A_Af7rwO4Z3_0;
	wire w_dff_A_cPeZ6SD53_0;
	wire w_dff_A_5hx7B5lh3_0;
	wire w_dff_A_Q6Nl3oap9_0;
	wire w_dff_A_zRuQDe172_0;
	wire w_dff_A_grXBwiRm9_0;
	wire w_dff_A_Sr2siA583_0;
	wire w_dff_A_ESw6a8MQ7_0;
	wire w_dff_A_4BjnqR7I0_0;
	wire w_dff_A_cRTrEahq9_0;
	wire w_dff_A_qmuqNwqD7_0;
	wire w_dff_A_YLFiNG3B4_0;
	wire w_dff_A_J1xrbLhx1_0;
	wire w_dff_A_OGLOL5e16_0;
	wire w_dff_A_NZ6qgRVI9_0;
	wire w_dff_A_yDktkIvR3_0;
	wire w_dff_A_6izQlhzq8_0;
	wire w_dff_A_7YKBEPnx5_0;
	wire w_dff_A_IoSZqDpj8_0;
	wire w_dff_A_5EeVt9Zi0_0;
	wire w_dff_A_XhSkDvQV1_0;
	wire w_dff_A_TVkwsmJZ4_0;
	wire w_dff_A_GNGWReUy8_0;
	wire w_dff_A_hsVe60Ms8_0;
	wire w_dff_A_7KETfTpp2_0;
	wire w_dff_A_QhwUvnqZ9_0;
	wire w_dff_A_FRo5TK4e1_0;
	wire w_dff_A_t2taBbP39_0;
	wire w_dff_A_rheuBGEr4_0;
	wire w_dff_A_rKnPW2378_0;
	wire w_dff_A_DFP2rKdu3_0;
	wire w_dff_A_xuXzxhla2_0;
	wire w_dff_A_sFJmA4jD6_0;
	wire w_dff_A_oVxZavgL9_0;
	wire w_dff_A_awQuYCXd9_0;
	wire w_dff_A_J4a8nY809_0;
	wire w_dff_A_2FgvZGJk8_0;
	wire w_dff_A_KmD7Mh4p8_0;
	wire w_dff_A_IjoCFhh39_0;
	wire w_dff_A_1RoD7IHH2_0;
	wire w_dff_A_qfEw5MSI1_0;
	wire w_dff_A_bJGkmqbU5_0;
	wire w_dff_A_jXJoTtAM3_0;
	wire w_dff_A_Vg6NI2J61_0;
	wire w_dff_A_qDULmxVk6_0;
	wire w_dff_A_LFMid0cB6_0;
	wire w_dff_A_2VakWFqR1_0;
	wire w_dff_A_7EZaGmYx2_0;
	wire w_dff_A_R4ues0R64_0;
	wire w_dff_A_YG7bvOdM3_0;
	wire w_dff_A_MgyK0MRL9_0;
	wire w_dff_A_R7FH4fbX2_0;
	wire w_dff_A_58MSGd9a7_0;
	wire w_dff_A_ZLwKLtJq3_0;
	wire w_dff_A_hqBdsfmR3_2;
	wire w_dff_A_sWOG7FHo8_0;
	wire w_dff_A_k077Uut50_0;
	wire w_dff_A_bADamjWn4_0;
	wire w_dff_A_Q60y1mUk9_0;
	wire w_dff_A_1mVcQcAE2_0;
	wire w_dff_A_fe1zIwkf6_0;
	wire w_dff_A_0VUjgbwC6_0;
	wire w_dff_A_As6ONpT40_0;
	wire w_dff_A_xnxkpoyT4_0;
	wire w_dff_A_HMsgNolo4_0;
	wire w_dff_A_gtfnUHQE7_0;
	wire w_dff_A_A3i2bFjX6_0;
	wire w_dff_A_UbUe2Kf17_0;
	wire w_dff_A_U1S8mGzU5_0;
	wire w_dff_A_Z6zYKh7O3_0;
	wire w_dff_A_ewdPHNFY3_0;
	wire w_dff_A_yuhBwgqv6_0;
	wire w_dff_A_wl9MechG2_0;
	wire w_dff_A_yCspxLdO2_0;
	wire w_dff_A_yaYyfitw1_0;
	wire w_dff_A_Xty69Cur9_0;
	wire w_dff_A_grMN48ne6_0;
	wire w_dff_A_LROwg5h05_0;
	wire w_dff_A_Uhaay64q2_0;
	wire w_dff_A_wmNJ4NLZ6_0;
	wire w_dff_A_bpGILDte4_0;
	wire w_dff_A_yiPhruxa3_0;
	wire w_dff_A_aC4K7Shp1_0;
	wire w_dff_A_KB6IMC2P3_0;
	wire w_dff_A_HZmqnJB74_0;
	wire w_dff_A_oyuTAxmT1_0;
	wire w_dff_A_IflzbrZW3_0;
	wire w_dff_A_xbGI44Ak3_0;
	wire w_dff_A_fSU4pXCM5_0;
	wire w_dff_A_QQ0lJoft1_0;
	wire w_dff_A_JqtMtWun6_0;
	wire w_dff_A_kv7h2Yzn8_0;
	wire w_dff_A_tKN3LHxy9_0;
	wire w_dff_A_DsBILMrL1_0;
	wire w_dff_A_33D6SsAU4_0;
	wire w_dff_A_hcMwm2DF9_0;
	wire w_dff_A_bLdxEBzI7_0;
	wire w_dff_A_feBtEQQh4_0;
	wire w_dff_A_6pYcdlUK1_0;
	wire w_dff_A_YB4C5e1F9_0;
	wire w_dff_A_8OiCmwzk0_0;
	wire w_dff_A_rDGj7Q1i0_0;
	wire w_dff_A_FxwGHjLl7_0;
	wire w_dff_A_8mrxMDRD8_0;
	wire w_dff_A_w5XAm7Bf9_0;
	wire w_dff_A_uhtTf1z16_0;
	wire w_dff_A_Hi1W0WRm2_0;
	wire w_dff_A_SZ4ePauA4_0;
	wire w_dff_A_cYOgFdTT7_0;
	wire w_dff_A_zFO9lnkS7_0;
	wire w_dff_A_QnOwsA0K0_0;
	wire w_dff_A_yUI10Bf42_0;
	wire w_dff_A_SbCVwLaa2_0;
	wire w_dff_A_lK38vy6x5_0;
	wire w_dff_A_435CGDln8_0;
	wire w_dff_A_mnr3JpNV6_0;
	wire w_dff_A_IMd2R1Fa5_0;
	wire w_dff_A_KrUrWVju1_0;
	wire w_dff_A_vWNn7eQH1_0;
	wire w_dff_A_vP6t7DhO5_0;
	wire w_dff_A_muhXB0j46_0;
	wire w_dff_A_w15OVzbB4_0;
	wire w_dff_A_bQyoU5vk1_0;
	wire w_dff_A_tsgWoKuc9_0;
	wire w_dff_A_mMoeQG1x2_0;
	wire w_dff_A_GZeM7Lgj3_0;
	wire w_dff_A_Tcs5UMHB1_0;
	wire w_dff_A_mVINKIeB2_0;
	wire w_dff_A_4yW2qVps5_0;
	wire w_dff_A_ioWvvnrU1_0;
	wire w_dff_A_QVFiNPEC8_0;
	wire w_dff_A_Koe9jSw08_0;
	wire w_dff_A_RCzhCTvV3_0;
	wire w_dff_A_y0RdezRs4_0;
	wire w_dff_A_IKfcsEwg4_0;
	wire w_dff_A_MHankf090_0;
	wire w_dff_A_uvgGtS777_0;
	wire w_dff_A_jYvkSs9A3_0;
	wire w_dff_A_VSOwTyg44_0;
	wire w_dff_A_ZpoxRcY69_0;
	wire w_dff_A_k9ra6rwE2_0;
	wire w_dff_A_prvXHNpo0_0;
	wire w_dff_A_dgwlu9WA5_0;
	wire w_dff_A_uxnVYdDa8_0;
	wire w_dff_A_6LswrDbN6_0;
	wire w_dff_A_GfsIvQtw0_0;
	wire w_dff_A_KSLFMHLk7_0;
	wire w_dff_A_sQckYULF7_0;
	wire w_dff_A_OmyVFBLf8_0;
	wire w_dff_A_3Lb1IWRL3_0;
	wire w_dff_A_NSTjunAr1_0;
	wire w_dff_A_BkhXo2AL4_0;
	wire w_dff_A_xaEYEOJW9_0;
	wire w_dff_A_D4qYnBMC2_0;
	wire w_dff_A_w0dYMDYg0_0;
	wire w_dff_A_getjz7V28_0;
	wire w_dff_A_7LpYKxFt5_0;
	wire w_dff_A_28W5aH2K6_0;
	wire w_dff_A_U5RnASk11_0;
	wire w_dff_A_r0GVk2Pe7_0;
	wire w_dff_A_TBVMeCGo8_0;
	wire w_dff_A_ErTjsSXk7_0;
	wire w_dff_A_2OZLHZDr4_0;
	wire w_dff_A_2ZqmUP6w1_0;
	wire w_dff_A_1riIuvg58_0;
	wire w_dff_A_CBWZWl9S5_0;
	wire w_dff_A_sx9ATPQC2_0;
	wire w_dff_A_6OrMUFPu2_0;
	wire w_dff_A_kf5oJuF46_0;
	wire w_dff_A_PFaQGYxK9_0;
	wire w_dff_A_pPuynFWl5_0;
	wire w_dff_A_XfMAWmc97_0;
	wire w_dff_A_gQEtfDcs9_0;
	wire w_dff_A_TPd6RMHY6_2;
	wire w_dff_A_5qhc1AdK0_0;
	wire w_dff_A_oKwebBb92_0;
	wire w_dff_A_ELgAvyqV1_0;
	wire w_dff_A_Fo1cNxNA2_0;
	wire w_dff_A_C4diHBCU1_0;
	wire w_dff_A_uG1H5xEk7_0;
	wire w_dff_A_VjwGpPpD4_0;
	wire w_dff_A_oFbnVh4y7_0;
	wire w_dff_A_BGYlffrk1_0;
	wire w_dff_A_Rvpn2TQb6_0;
	wire w_dff_A_TuUKr8CC7_0;
	wire w_dff_A_Kr0BLb9U2_0;
	wire w_dff_A_C8WuXlrQ4_0;
	wire w_dff_A_fJE7ZlUa4_0;
	wire w_dff_A_ng8tJ7AN0_0;
	wire w_dff_A_gTG3JZtX0_0;
	wire w_dff_A_pdKGmA085_0;
	wire w_dff_A_9jyAnHEI8_0;
	wire w_dff_A_soDGOWyV4_0;
	wire w_dff_A_J540FnmE3_0;
	wire w_dff_A_oapD8LyZ5_0;
	wire w_dff_A_ekk7WLap6_0;
	wire w_dff_A_odu7KFF12_0;
	wire w_dff_A_5O5Xh0b56_0;
	wire w_dff_A_0dyfs50F7_0;
	wire w_dff_A_8MJ5XxQ18_0;
	wire w_dff_A_YfwHMbUa5_0;
	wire w_dff_A_4rG5yjCy7_0;
	wire w_dff_A_Xw86b9FC6_0;
	wire w_dff_A_Qs1lpwUU0_0;
	wire w_dff_A_JiPUreyM7_0;
	wire w_dff_A_jvkWY0FK8_0;
	wire w_dff_A_zUZYuJGC7_0;
	wire w_dff_A_wWAf9Xjw7_0;
	wire w_dff_A_81tWg6aq9_0;
	wire w_dff_A_P0IYBxEW8_0;
	wire w_dff_A_mrvY481p7_0;
	wire w_dff_A_vHQRbkbV7_0;
	wire w_dff_A_F0mOwgfQ5_0;
	wire w_dff_A_yWa4bRM23_0;
	wire w_dff_A_yI9ITnt29_0;
	wire w_dff_A_nkufeQnA9_0;
	wire w_dff_A_nTY9AT0U0_0;
	wire w_dff_A_S4GDwsci3_0;
	wire w_dff_A_ZhhuA6U36_0;
	wire w_dff_A_okZIWMFN2_0;
	wire w_dff_A_MJUYoofZ8_0;
	wire w_dff_A_bnwczqnS6_0;
	wire w_dff_A_XhCA6d1Z8_0;
	wire w_dff_A_lYO78a6M6_0;
	wire w_dff_A_TEOSqEFu7_0;
	wire w_dff_A_1vOBBOuH5_0;
	wire w_dff_A_RHaFhZBA5_0;
	wire w_dff_A_cAjkRbEU0_0;
	wire w_dff_A_a2hoNyqg4_0;
	wire w_dff_A_uIWdLd6w0_0;
	wire w_dff_A_bGLF6RKs0_0;
	wire w_dff_A_UOjJV8NZ0_0;
	wire w_dff_A_gE4pJxjk0_0;
	wire w_dff_A_ZvmtSwUG1_0;
	wire w_dff_A_MXobBHJP2_0;
	wire w_dff_A_hebXh9ER7_0;
	wire w_dff_A_SRDDYPek9_0;
	wire w_dff_A_evICsUMv8_0;
	wire w_dff_A_f3h2CkNv2_0;
	wire w_dff_A_iQBt9nmS5_0;
	wire w_dff_A_SziMIP2j1_0;
	wire w_dff_A_UJJV25nb3_0;
	wire w_dff_A_uYoSwYDn7_0;
	wire w_dff_A_ts7zJ5Tb7_0;
	wire w_dff_A_F6w6UlAx6_0;
	wire w_dff_A_sYp8UMwn9_0;
	wire w_dff_A_EJo59HU06_0;
	wire w_dff_A_pbbhVIpa0_0;
	wire w_dff_A_AFHu6rDq3_0;
	wire w_dff_A_sN6r5Psz8_0;
	wire w_dff_A_9zncHu7w2_0;
	wire w_dff_A_Ixb7AvpI6_0;
	wire w_dff_A_d2qge45n1_0;
	wire w_dff_A_gploWS1K6_0;
	wire w_dff_A_a1G9LEd90_0;
	wire w_dff_A_VKvFcBOQ3_0;
	wire w_dff_A_kPzPb2ib5_0;
	wire w_dff_A_KT5Pzb5p2_0;
	wire w_dff_A_2UifLQiR5_0;
	wire w_dff_A_WOZEytYC2_0;
	wire w_dff_A_VKkH7hu57_0;
	wire w_dff_A_8ovRG4gm6_0;
	wire w_dff_A_coIA58xT9_0;
	wire w_dff_A_5lQMfcsz7_0;
	wire w_dff_A_HydVFWFi0_0;
	wire w_dff_A_cbBspt3o2_0;
	wire w_dff_A_Cug2ntA18_0;
	wire w_dff_A_JItWcIBc7_0;
	wire w_dff_A_YfheOsXd8_0;
	wire w_dff_A_bXFhU7yJ8_0;
	wire w_dff_A_fqp1ss0R2_0;
	wire w_dff_A_aW1GduXA8_0;
	wire w_dff_A_qgbVWWsa7_0;
	wire w_dff_A_2dzkjre17_0;
	wire w_dff_A_ti3AE9Nx9_0;
	wire w_dff_A_3PPjiAZw2_0;
	wire w_dff_A_GblVuIFG4_0;
	wire w_dff_A_orpG6eH67_0;
	wire w_dff_A_AoYMz5245_0;
	wire w_dff_A_jP4YGIUT1_0;
	wire w_dff_A_B3R1hoNp8_0;
	wire w_dff_A_g0A8uaiE3_0;
	wire w_dff_A_Qqr0eMQf2_0;
	wire w_dff_A_gk7QQ19M1_0;
	wire w_dff_A_cICvejxt9_0;
	wire w_dff_A_g7qhwGua2_0;
	wire w_dff_A_0YxtZ9R23_0;
	wire w_dff_A_lmO3bB5r4_0;
	wire w_dff_A_Vn8QyEAP3_0;
	wire w_dff_A_CCCqz7dS7_0;
	wire w_dff_A_GSewm7ZW8_0;
	wire w_dff_A_K99ijCAz4_2;
	wire w_dff_A_jjVoD3AR3_0;
	wire w_dff_A_760m2NFX7_0;
	wire w_dff_A_iu1oGKb55_0;
	wire w_dff_A_Pb5Ssgcu6_0;
	wire w_dff_A_Czh0R1hf9_0;
	wire w_dff_A_uMob2VTh3_0;
	wire w_dff_A_4mW44HZk6_0;
	wire w_dff_A_awGgXWEf0_0;
	wire w_dff_A_Efs3Kc2K5_0;
	wire w_dff_A_KNXOpXvx0_0;
	wire w_dff_A_XOKGgzQL0_0;
	wire w_dff_A_MvhTjEBJ9_0;
	wire w_dff_A_aAZ6A1kX5_0;
	wire w_dff_A_IGLhGCm57_0;
	wire w_dff_A_B0VJY4VC9_0;
	wire w_dff_A_UsEBKtdf5_0;
	wire w_dff_A_zHZPFIvM2_0;
	wire w_dff_A_vDSd9rkY7_0;
	wire w_dff_A_WYATVSAs8_0;
	wire w_dff_A_jIQYJQWf5_0;
	wire w_dff_A_SDmt4iOz2_0;
	wire w_dff_A_iKBXCCy35_0;
	wire w_dff_A_8oz9Wyhx9_0;
	wire w_dff_A_5fPehC8h2_0;
	wire w_dff_A_q02Z14UO1_0;
	wire w_dff_A_k0u9xkPa3_0;
	wire w_dff_A_A4EBHP5a6_0;
	wire w_dff_A_JXLuhsgi7_0;
	wire w_dff_A_fT2p0KIq1_0;
	wire w_dff_A_Y6hv9qId6_0;
	wire w_dff_A_mMrFIkb33_0;
	wire w_dff_A_OkStu4Nd7_0;
	wire w_dff_A_SRX7Yj785_0;
	wire w_dff_A_diBiWOwM1_0;
	wire w_dff_A_joy2avoE4_0;
	wire w_dff_A_6qUWlzKo3_0;
	wire w_dff_A_Nw2b6nGT1_0;
	wire w_dff_A_pGLygNaG3_0;
	wire w_dff_A_h9KHelO10_0;
	wire w_dff_A_1zDzRekS7_0;
	wire w_dff_A_2y0DEzx67_0;
	wire w_dff_A_QShYQLxL0_0;
	wire w_dff_A_1pWeIyes3_0;
	wire w_dff_A_wBuutEON8_0;
	wire w_dff_A_LHfcZzWz7_0;
	wire w_dff_A_GMAWCa3R2_0;
	wire w_dff_A_ktH5KyYO5_0;
	wire w_dff_A_yws4mdaT6_0;
	wire w_dff_A_PulnezTO5_0;
	wire w_dff_A_m9ajVUs85_0;
	wire w_dff_A_ic4iOkUk1_0;
	wire w_dff_A_L0Gnt5tY2_0;
	wire w_dff_A_Vt3B8Vjt5_0;
	wire w_dff_A_NE52HxQy2_0;
	wire w_dff_A_0CpsxfaY4_0;
	wire w_dff_A_7QVX24J51_0;
	wire w_dff_A_zgn1OfDh1_0;
	wire w_dff_A_KGSIwgul8_0;
	wire w_dff_A_p7PSgJBZ2_0;
	wire w_dff_A_yv9LbyyV0_0;
	wire w_dff_A_1VLkec4L8_0;
	wire w_dff_A_ZhHCxTWs3_0;
	wire w_dff_A_hmLEYL4z4_0;
	wire w_dff_A_ZfWKkrDK8_0;
	wire w_dff_A_r3SQdPc77_0;
	wire w_dff_A_ORuSLANz5_0;
	wire w_dff_A_rFJeUEJU0_0;
	wire w_dff_A_nGz2vt9n0_0;
	wire w_dff_A_zbZiWfSE7_0;
	wire w_dff_A_8ux4ot8R9_0;
	wire w_dff_A_xU0AWXYE5_0;
	wire w_dff_A_WCdDihVX1_0;
	wire w_dff_A_XDqWUvbp7_0;
	wire w_dff_A_4iZsL2TP3_0;
	wire w_dff_A_GGLarvz40_0;
	wire w_dff_A_ycCWEksQ1_0;
	wire w_dff_A_Pe75E43a6_0;
	wire w_dff_A_SNd5FNiI3_0;
	wire w_dff_A_fiMYGD467_0;
	wire w_dff_A_ZpZkZq6D0_0;
	wire w_dff_A_Zdi3dTfX2_0;
	wire w_dff_A_mGmPoZMn2_0;
	wire w_dff_A_hpHhMutO5_0;
	wire w_dff_A_rZsGNHMR6_0;
	wire w_dff_A_wHLYRihD5_0;
	wire w_dff_A_fQ9m1BRv2_0;
	wire w_dff_A_582nucf89_0;
	wire w_dff_A_8lCQdlDI3_0;
	wire w_dff_A_tAdABm3I0_0;
	wire w_dff_A_L9hMv4S83_0;
	wire w_dff_A_XL0RG6jC6_0;
	wire w_dff_A_YoNPNwg12_0;
	wire w_dff_A_QswfTllp6_0;
	wire w_dff_A_QBQbdsmn7_0;
	wire w_dff_A_XSgTPFmZ9_0;
	wire w_dff_A_oTrKD4mT9_0;
	wire w_dff_A_6ntrtNGS0_0;
	wire w_dff_A_Bt5YQ6nr5_0;
	wire w_dff_A_5UkpyXkc2_0;
	wire w_dff_A_kRMDWBnH1_0;
	wire w_dff_A_TWfXQ2Sl3_0;
	wire w_dff_A_TfOavHbc7_0;
	wire w_dff_A_UPVyrwD12_0;
	wire w_dff_A_bSkYozi36_0;
	wire w_dff_A_Jh2bbCCl4_0;
	wire w_dff_A_LOhNhGVW7_0;
	wire w_dff_A_ySUfGGmy5_0;
	wire w_dff_A_qqT8UNDI9_0;
	wire w_dff_A_6cVKGCjB0_0;
	wire w_dff_A_LvN6XhM73_0;
	wire w_dff_A_jQgHP0PG2_0;
	wire w_dff_A_qQcI16md6_0;
	wire w_dff_A_3ZXZ8AV16_0;
	wire w_dff_A_ZOzEY6Re4_0;
	wire w_dff_A_LUoCgbM72_0;
	wire w_dff_A_HvvODXkS3_0;
	wire w_dff_A_ZrWr9ERl4_2;
	wire w_dff_A_15HcQg9U7_0;
	wire w_dff_A_UgVoAuRx9_0;
	wire w_dff_A_6bKLCRhg7_0;
	wire w_dff_A_HnbtIPTM7_0;
	wire w_dff_A_bNSqxWpw3_0;
	wire w_dff_A_yZdg2bYG1_0;
	wire w_dff_A_C7rHcHnE5_0;
	wire w_dff_A_aBedArzx6_0;
	wire w_dff_A_ihv0gZ9z8_0;
	wire w_dff_A_7UajP3OS9_0;
	wire w_dff_A_ql6x8v0S3_0;
	wire w_dff_A_4NZ6UZoi0_0;
	wire w_dff_A_TFI8iHyh5_0;
	wire w_dff_A_pXWqM8PU1_0;
	wire w_dff_A_MP4QBkco0_0;
	wire w_dff_A_2hcH2NAN2_0;
	wire w_dff_A_Zbo3kZsU8_0;
	wire w_dff_A_8iylWzLJ3_0;
	wire w_dff_A_qiiQj4bI9_0;
	wire w_dff_A_4F24Tn4b3_0;
	wire w_dff_A_02mVP7GQ0_0;
	wire w_dff_A_rTUjMI7x2_0;
	wire w_dff_A_EyhoHLkS2_0;
	wire w_dff_A_bpx99x1V6_0;
	wire w_dff_A_7leawFfC3_0;
	wire w_dff_A_VJA0fGUk6_0;
	wire w_dff_A_qJeP7gsc4_0;
	wire w_dff_A_9JithcuB7_0;
	wire w_dff_A_Xprvgxjm3_0;
	wire w_dff_A_YiEK16rm4_0;
	wire w_dff_A_fYv0izgo3_0;
	wire w_dff_A_3dcNZQKF6_0;
	wire w_dff_A_yEf3t1Fx3_0;
	wire w_dff_A_hOFFA0jj0_0;
	wire w_dff_A_fBuzkhkP4_0;
	wire w_dff_A_5iiAkiTO5_0;
	wire w_dff_A_W9OkXWNG4_0;
	wire w_dff_A_kHYDAXqZ8_0;
	wire w_dff_A_gbD6eOfb5_0;
	wire w_dff_A_YOzaICmi4_0;
	wire w_dff_A_vpE0DHAH5_0;
	wire w_dff_A_wS7BklKo3_0;
	wire w_dff_A_jzKdHl3s1_0;
	wire w_dff_A_epCTTsWm8_0;
	wire w_dff_A_9HpT1eWw8_0;
	wire w_dff_A_nCzWPstu1_0;
	wire w_dff_A_SUSXpkHA8_0;
	wire w_dff_A_0VmBQBJr8_0;
	wire w_dff_A_bFYvkhAP3_0;
	wire w_dff_A_IxllTX1D4_0;
	wire w_dff_A_ePPRqBus1_0;
	wire w_dff_A_fb60NbWI2_0;
	wire w_dff_A_pSZQOTxJ4_0;
	wire w_dff_A_dC2NcBKJ1_0;
	wire w_dff_A_JrCTLoXY6_0;
	wire w_dff_A_SkJD0Apt5_0;
	wire w_dff_A_yIkeT2ln9_0;
	wire w_dff_A_S6bOPlNl4_0;
	wire w_dff_A_axCSck3S7_0;
	wire w_dff_A_cK4FlwEo1_0;
	wire w_dff_A_wUOK7QKQ4_0;
	wire w_dff_A_10TaH3VO1_0;
	wire w_dff_A_J2CPWDlv9_0;
	wire w_dff_A_hpt6nDx61_0;
	wire w_dff_A_unztLCtB1_0;
	wire w_dff_A_1zCq4sQO2_0;
	wire w_dff_A_dFoNTzyt0_0;
	wire w_dff_A_1bn6RTcI0_0;
	wire w_dff_A_fE1ekTHR0_0;
	wire w_dff_A_6wjvUxBG5_0;
	wire w_dff_A_tsagRu9B4_0;
	wire w_dff_A_nbLw0WLj6_0;
	wire w_dff_A_qVOIaLGz1_0;
	wire w_dff_A_pQj4XA6F6_0;
	wire w_dff_A_lenHzLJi4_0;
	wire w_dff_A_eEBgcmwB1_0;
	wire w_dff_A_dNFtxpV62_0;
	wire w_dff_A_EZCKI5Vp6_0;
	wire w_dff_A_TlBzjPzF9_0;
	wire w_dff_A_DZcnUb4g1_0;
	wire w_dff_A_5T5pFwlh1_0;
	wire w_dff_A_pNhYQ22y8_0;
	wire w_dff_A_rr4vJImw4_0;
	wire w_dff_A_rfMzGpFH8_0;
	wire w_dff_A_RblJ08sR7_0;
	wire w_dff_A_eRWA5Weh2_0;
	wire w_dff_A_bUCnsmSF5_0;
	wire w_dff_A_3G2OhcFT1_0;
	wire w_dff_A_ZbdzZVdS4_0;
	wire w_dff_A_k3DCA6SB9_0;
	wire w_dff_A_ET9lZcgD0_0;
	wire w_dff_A_OQNcGgK65_0;
	wire w_dff_A_QG532PEa1_0;
	wire w_dff_A_XNzX6bgo5_0;
	wire w_dff_A_7ZavvGFy8_0;
	wire w_dff_A_jltbk1ix3_0;
	wire w_dff_A_o3bY3S3Y3_0;
	wire w_dff_A_H0hyyIro3_0;
	wire w_dff_A_uoAR7BSt3_0;
	wire w_dff_A_ZIn0HoNO2_0;
	wire w_dff_A_B9WWfpk30_0;
	wire w_dff_A_FO6D9ciQ6_0;
	wire w_dff_A_b3l3KliC4_0;
	wire w_dff_A_UYf7O8Tk2_0;
	wire w_dff_A_7aOcJt900_0;
	wire w_dff_A_6bqglOVK8_0;
	wire w_dff_A_AHXZk2rw1_0;
	wire w_dff_A_dKkO9qPk8_0;
	wire w_dff_A_ZQNDci8i0_0;
	wire w_dff_A_oN8lrO2u9_0;
	wire w_dff_A_B0zb1x6Q7_0;
	wire w_dff_A_PivgCzWd9_0;
	wire w_dff_A_QE7SKFjN1_0;
	wire w_dff_A_ZFs8B1zb2_0;
	wire w_dff_A_5DUOrROx7_0;
	wire w_dff_A_fR6FTcm21_2;
	wire w_dff_A_y7WhSNYQ7_0;
	wire w_dff_A_6z1nnNHl4_0;
	wire w_dff_A_XaOXOBOL0_0;
	wire w_dff_A_fodcdQKs6_0;
	wire w_dff_A_7BXV6UXY4_0;
	wire w_dff_A_tm0QLkmT1_0;
	wire w_dff_A_fZ3G0fIF0_0;
	wire w_dff_A_sihbW0vt7_0;
	wire w_dff_A_SVDLCNvx2_0;
	wire w_dff_A_6wDwT20S0_0;
	wire w_dff_A_bmPmeZCt2_0;
	wire w_dff_A_7RF50jCU8_0;
	wire w_dff_A_zAJRgU9d4_0;
	wire w_dff_A_3ToLIOZR1_0;
	wire w_dff_A_ikKcsmME0_0;
	wire w_dff_A_I3KAtPI58_0;
	wire w_dff_A_LCDkvxGM6_0;
	wire w_dff_A_WzzIVol07_0;
	wire w_dff_A_IaCWVXSM4_0;
	wire w_dff_A_nP8h33mC4_0;
	wire w_dff_A_trIiBRfK7_0;
	wire w_dff_A_FbYro3jv7_0;
	wire w_dff_A_TS5kjr0u8_0;
	wire w_dff_A_2jmUOqW10_0;
	wire w_dff_A_IYyeKXR31_0;
	wire w_dff_A_lqPIHeOr2_0;
	wire w_dff_A_AwcBvLbG3_0;
	wire w_dff_A_5w7Gfoom7_0;
	wire w_dff_A_GZnb6yT07_0;
	wire w_dff_A_U3YbTNFS4_0;
	wire w_dff_A_8j1E2ceg7_0;
	wire w_dff_A_SbMbh9sX0_0;
	wire w_dff_A_dnfJeEbh7_0;
	wire w_dff_A_dvvq5irm7_0;
	wire w_dff_A_iGp2IYsb1_0;
	wire w_dff_A_584jK6gU6_0;
	wire w_dff_A_iaokvyBS5_0;
	wire w_dff_A_B2cji4F71_0;
	wire w_dff_A_IHyt1oMD4_0;
	wire w_dff_A_kllMZS7q3_0;
	wire w_dff_A_NJSNWmYt1_0;
	wire w_dff_A_9n9jj4344_0;
	wire w_dff_A_FoO0ayB03_0;
	wire w_dff_A_j6Ts3P5a0_0;
	wire w_dff_A_P99ZzB4Y7_0;
	wire w_dff_A_75W9U8704_0;
	wire w_dff_A_c1z5pt989_0;
	wire w_dff_A_PPjWTK8L3_0;
	wire w_dff_A_6SzfAzzR1_0;
	wire w_dff_A_sWS2HhKH6_0;
	wire w_dff_A_tRTxfeMJ1_0;
	wire w_dff_A_BxW6PY2o8_0;
	wire w_dff_A_EHoXfIBY4_0;
	wire w_dff_A_1J4FoOdO4_0;
	wire w_dff_A_gAqIS2lD5_0;
	wire w_dff_A_xCvvQE6d4_0;
	wire w_dff_A_R8kdQ0IK5_0;
	wire w_dff_A_lTAphZi96_0;
	wire w_dff_A_5Swu2wGt3_0;
	wire w_dff_A_OlcjcwmA3_0;
	wire w_dff_A_LNM75Euf6_0;
	wire w_dff_A_cPrvOmTY3_0;
	wire w_dff_A_058Cf25e8_0;
	wire w_dff_A_KDS1bbSl9_0;
	wire w_dff_A_YNJYXBCF9_0;
	wire w_dff_A_xleCjhWi7_0;
	wire w_dff_A_rq4jptBu8_0;
	wire w_dff_A_UaFuHvic3_0;
	wire w_dff_A_9QAQU2qe9_0;
	wire w_dff_A_Y4dGORsR3_0;
	wire w_dff_A_aY0ry2Gg2_0;
	wire w_dff_A_ldrmDmAz6_0;
	wire w_dff_A_4ql2nkjp8_0;
	wire w_dff_A_Iht7PWfw9_0;
	wire w_dff_A_5LtbLBHI5_0;
	wire w_dff_A_UUERqg471_0;
	wire w_dff_A_iKFmuGJR0_0;
	wire w_dff_A_GdrE35gt8_0;
	wire w_dff_A_pJSrhPX42_0;
	wire w_dff_A_3h1DO1Y98_0;
	wire w_dff_A_kB1qCdO48_0;
	wire w_dff_A_tciRGW9O9_0;
	wire w_dff_A_1IZjxcza9_0;
	wire w_dff_A_EelNvNHN2_0;
	wire w_dff_A_tRxX3MST2_0;
	wire w_dff_A_NjMjIRqf6_0;
	wire w_dff_A_MSuLK1OP9_0;
	wire w_dff_A_7MM59aGF9_0;
	wire w_dff_A_X3Qqwu5C6_0;
	wire w_dff_A_epdSzUUA3_0;
	wire w_dff_A_UKxYtE504_0;
	wire w_dff_A_G6vb3wgD2_0;
	wire w_dff_A_jvt5CBJk3_0;
	wire w_dff_A_cqwQ3lgT8_0;
	wire w_dff_A_PWeN0vfI1_0;
	wire w_dff_A_30WlPK1O7_0;
	wire w_dff_A_KjMxXW2Z7_0;
	wire w_dff_A_rWHmgSme1_0;
	wire w_dff_A_GKLPcDGC0_0;
	wire w_dff_A_I863mCVa7_0;
	wire w_dff_A_na5gntbZ1_0;
	wire w_dff_A_yD6dehP53_0;
	wire w_dff_A_HNdbQz9a0_0;
	wire w_dff_A_JgLAJzPS0_0;
	wire w_dff_A_HT3oSSMJ1_0;
	wire w_dff_A_HT34WWlX5_0;
	wire w_dff_A_cBHBIEwD0_0;
	wire w_dff_A_hZAJBVeo9_0;
	wire w_dff_A_9HjBetnd0_0;
	wire w_dff_A_oATdPfMO9_0;
	wire w_dff_A_VuFtPo5K3_0;
	wire w_dff_A_dGceOg5Q2_0;
	wire w_dff_A_rI8AILxN3_0;
	wire w_dff_A_LMG2NbA00_0;
	wire w_dff_A_4btOcuhR0_2;
	wire w_dff_A_hXttFBOs2_0;
	wire w_dff_A_NvtMBi6u3_0;
	wire w_dff_A_03ZgzymL3_0;
	wire w_dff_A_y94CJZe51_0;
	wire w_dff_A_oYuZa7Dx0_0;
	wire w_dff_A_hoG73kf65_0;
	wire w_dff_A_cuhbW1WL3_0;
	wire w_dff_A_m8zZi9If8_0;
	wire w_dff_A_PD4rlpDZ4_0;
	wire w_dff_A_UZk2ijKF5_0;
	wire w_dff_A_m7OtoNr67_0;
	wire w_dff_A_mcqoY2Nm9_0;
	wire w_dff_A_Yx0d6Ig68_0;
	wire w_dff_A_4GUKwdtm9_0;
	wire w_dff_A_Js0auYev8_0;
	wire w_dff_A_jH6ElGOA3_0;
	wire w_dff_A_iINnE84N6_0;
	wire w_dff_A_oXY8KzHG9_0;
	wire w_dff_A_wSsS3qDZ9_0;
	wire w_dff_A_Tk2tLxqK3_0;
	wire w_dff_A_YHSGDYhC2_0;
	wire w_dff_A_nxc5s4eE8_0;
	wire w_dff_A_C9PjyOXE4_0;
	wire w_dff_A_shMjUDjF5_0;
	wire w_dff_A_WLnTsOxJ1_0;
	wire w_dff_A_Ke7AJq487_0;
	wire w_dff_A_IK6Sb2gW9_0;
	wire w_dff_A_CROxuNKx5_0;
	wire w_dff_A_6pD50PzY3_0;
	wire w_dff_A_DZ94IGi22_0;
	wire w_dff_A_Q5TRQSnK2_0;
	wire w_dff_A_qySVJRl90_0;
	wire w_dff_A_oTrtil7C2_0;
	wire w_dff_A_awa57HLB7_0;
	wire w_dff_A_ZWbfvXf69_0;
	wire w_dff_A_hX1HJ0Sl6_0;
	wire w_dff_A_paQmIG9L8_0;
	wire w_dff_A_wkUkTNpX6_0;
	wire w_dff_A_959lsYZv3_0;
	wire w_dff_A_dkQiuSUf5_0;
	wire w_dff_A_KtPPWwrf5_0;
	wire w_dff_A_MN2bDWSH3_0;
	wire w_dff_A_CTxRTJUc4_0;
	wire w_dff_A_ppYLMWDX7_0;
	wire w_dff_A_gOKEH9Mi3_0;
	wire w_dff_A_lwFhZSV63_0;
	wire w_dff_A_lFXtpmMq2_0;
	wire w_dff_A_5IykvP8q6_0;
	wire w_dff_A_D9s2Wfyp0_0;
	wire w_dff_A_903UcYyy5_0;
	wire w_dff_A_MADuVCyn5_0;
	wire w_dff_A_WJgNyte32_0;
	wire w_dff_A_9PASpTxr3_0;
	wire w_dff_A_ZgXvYBUH0_0;
	wire w_dff_A_dnv5g5VS8_0;
	wire w_dff_A_vr9q5a4S4_0;
	wire w_dff_A_7q12eyA13_0;
	wire w_dff_A_OjjTLHzT5_0;
	wire w_dff_A_BaVuN3mm1_0;
	wire w_dff_A_9VScVT5G7_0;
	wire w_dff_A_yCVnoLKQ1_0;
	wire w_dff_A_iSAmVDXf0_0;
	wire w_dff_A_09faWQrZ7_0;
	wire w_dff_A_Z3QjOCNN7_0;
	wire w_dff_A_iQgFg42F6_0;
	wire w_dff_A_WMZk7W2y7_0;
	wire w_dff_A_oVGfMUpW3_0;
	wire w_dff_A_gmPSRknr4_0;
	wire w_dff_A_FbCGl2cr6_0;
	wire w_dff_A_O8zju9cV9_0;
	wire w_dff_A_3wkPSCpg4_0;
	wire w_dff_A_u5nLHFer9_0;
	wire w_dff_A_mGWophlX7_0;
	wire w_dff_A_D8zotPIB7_0;
	wire w_dff_A_ZOKX4UXf0_0;
	wire w_dff_A_EMskCxFE2_0;
	wire w_dff_A_SSE4Bm1T4_0;
	wire w_dff_A_Whknq80S8_0;
	wire w_dff_A_kf3sdHL45_0;
	wire w_dff_A_sqeAyzXR3_0;
	wire w_dff_A_hNqkMtzr7_0;
	wire w_dff_A_ZDeP8kxK7_0;
	wire w_dff_A_ZE0cJZ223_0;
	wire w_dff_A_iXdsnQH82_0;
	wire w_dff_A_Rgooxdmk6_0;
	wire w_dff_A_FRqZLU7g3_0;
	wire w_dff_A_WkppzNmy0_0;
	wire w_dff_A_OLWEjz9g8_0;
	wire w_dff_A_q8xt3tDc8_0;
	wire w_dff_A_WLIDP5Zz4_0;
	wire w_dff_A_GNTGMBKc9_0;
	wire w_dff_A_sHjPr8Sp6_0;
	wire w_dff_A_wMIC8CQo7_0;
	wire w_dff_A_HYOM6pDn3_0;
	wire w_dff_A_DcSnrUzy5_0;
	wire w_dff_A_d8TqntnM0_0;
	wire w_dff_A_9KmiWiT92_0;
	wire w_dff_A_CT2Q01WD5_0;
	wire w_dff_A_AN1R04cO2_0;
	wire w_dff_A_V85UJkYn6_0;
	wire w_dff_A_bP85bTp89_0;
	wire w_dff_A_JyAypsUK6_0;
	wire w_dff_A_T9KwLQ7H4_0;
	wire w_dff_A_1GdOwlCq2_0;
	wire w_dff_A_7Vw4aZnR7_0;
	wire w_dff_A_WU4B3Z2E4_0;
	wire w_dff_A_Nde80F1o6_0;
	wire w_dff_A_E2eAmiMl8_0;
	wire w_dff_A_911xVSQE4_0;
	wire w_dff_A_SYbQqYQ70_0;
	wire w_dff_A_AUQl2ueY1_0;
	wire w_dff_A_PkaHEOyh8_0;
	wire w_dff_A_I02I6plj8_0;
	wire w_dff_A_KPqmqRhW5_2;
	wire w_dff_A_SgEdjVGx2_0;
	wire w_dff_A_HetkYEha4_0;
	wire w_dff_A_FH4ChRH80_0;
	wire w_dff_A_3cukWHsP5_0;
	wire w_dff_A_hm9tdfo84_0;
	wire w_dff_A_abnwBoSd5_0;
	wire w_dff_A_KyhkWLMK4_0;
	wire w_dff_A_mB5zRLED2_0;
	wire w_dff_A_MtOVPXtJ6_0;
	wire w_dff_A_vx89dJhg2_0;
	wire w_dff_A_mApcxBhK0_0;
	wire w_dff_A_1Bw9t0Vv9_0;
	wire w_dff_A_WUYuQ3Ax1_0;
	wire w_dff_A_tE06Q4IP3_0;
	wire w_dff_A_t6Yvze558_0;
	wire w_dff_A_vnJpdQZV7_0;
	wire w_dff_A_kw3bRMWl0_0;
	wire w_dff_A_3SqsgBYE9_0;
	wire w_dff_A_OtfD1YTa1_0;
	wire w_dff_A_vrtYWndX5_0;
	wire w_dff_A_czRBBvUL5_0;
	wire w_dff_A_vRp4RSR39_0;
	wire w_dff_A_IGtA3qJy1_0;
	wire w_dff_A_jKrfyg6H5_0;
	wire w_dff_A_0muZVTpA4_0;
	wire w_dff_A_lPGHCTwF3_0;
	wire w_dff_A_PK428G8O8_0;
	wire w_dff_A_CTONW30k7_0;
	wire w_dff_A_qEYXtEOp1_0;
	wire w_dff_A_EdgR7YUl9_0;
	wire w_dff_A_aqlmcIsW4_0;
	wire w_dff_A_5TzlW5AR2_0;
	wire w_dff_A_D39lk0xg3_0;
	wire w_dff_A_UM0DZMHy4_0;
	wire w_dff_A_2JFILxsC6_0;
	wire w_dff_A_NEVK5IJE1_0;
	wire w_dff_A_zyzHFxkr2_0;
	wire w_dff_A_xlZHsfPf5_0;
	wire w_dff_A_vEICNVV24_0;
	wire w_dff_A_iuatYexV2_0;
	wire w_dff_A_rKCpqKrG3_0;
	wire w_dff_A_CqEKkPbK0_0;
	wire w_dff_A_TQXV4JQl7_0;
	wire w_dff_A_UabOpz156_0;
	wire w_dff_A_5HSLAxjs0_0;
	wire w_dff_A_74n0dB3u6_0;
	wire w_dff_A_yFPpCaQx4_0;
	wire w_dff_A_c4edFJCv7_0;
	wire w_dff_A_lDQQ5RYS4_0;
	wire w_dff_A_XnkbO31U1_0;
	wire w_dff_A_DzICmh9B7_0;
	wire w_dff_A_dcAgGSrA6_0;
	wire w_dff_A_K2pbJSQb0_0;
	wire w_dff_A_GQwykDTQ5_0;
	wire w_dff_A_EXnHnrBS4_0;
	wire w_dff_A_v9AW4DIs7_0;
	wire w_dff_A_HNUIv0sg7_0;
	wire w_dff_A_dfeB26CL8_0;
	wire w_dff_A_SqOiAhrx1_0;
	wire w_dff_A_s8GkfFRS9_0;
	wire w_dff_A_UNxOZJac6_0;
	wire w_dff_A_NjGcVTVh4_0;
	wire w_dff_A_Xi0GEigo5_0;
	wire w_dff_A_hCSux4bt4_0;
	wire w_dff_A_Q0QoWgoU9_0;
	wire w_dff_A_6Ey0CQTk8_0;
	wire w_dff_A_DezHMF1g1_0;
	wire w_dff_A_tzD4vyM12_0;
	wire w_dff_A_H186WLXv5_0;
	wire w_dff_A_nmNhH4aX5_0;
	wire w_dff_A_CGWHNEyM2_0;
	wire w_dff_A_pSnjdBT06_0;
	wire w_dff_A_YukesCli4_0;
	wire w_dff_A_f9DTe8DA1_0;
	wire w_dff_A_F5QjwUTG0_0;
	wire w_dff_A_SxUiaafq4_0;
	wire w_dff_A_D5JkIpho2_0;
	wire w_dff_A_f53AXXp54_0;
	wire w_dff_A_8hkLduPJ5_0;
	wire w_dff_A_TbkNVXXF9_0;
	wire w_dff_A_9B3bhSv31_0;
	wire w_dff_A_0NWDLrLV9_0;
	wire w_dff_A_CdA1pW6V7_0;
	wire w_dff_A_dP6BUQ6o9_0;
	wire w_dff_A_zwJ9pYKE7_0;
	wire w_dff_A_pHlrahvY2_0;
	wire w_dff_A_4BsRjjQK7_0;
	wire w_dff_A_5RTGDfZC7_0;
	wire w_dff_A_BkQHaBjS7_0;
	wire w_dff_A_c8tUtC9C0_0;
	wire w_dff_A_b9qcIKjf4_0;
	wire w_dff_A_ijFYYkgr2_0;
	wire w_dff_A_VW6FtWRb6_0;
	wire w_dff_A_jpkbdgbo6_0;
	wire w_dff_A_fHGKWQYF2_0;
	wire w_dff_A_WmNQ3cQ84_0;
	wire w_dff_A_efv7ck776_0;
	wire w_dff_A_Trn2HCBl7_0;
	wire w_dff_A_iPbWYITl4_0;
	wire w_dff_A_p483Fs4E8_0;
	wire w_dff_A_3xps0bi00_0;
	wire w_dff_A_96dI2mB01_0;
	wire w_dff_A_9BsK8oIj7_0;
	wire w_dff_A_mcXaiTRj5_0;
	wire w_dff_A_oRANdWsb5_0;
	wire w_dff_A_UFtg8Tvl1_0;
	wire w_dff_A_Ge4dLXhI6_0;
	wire w_dff_A_yucONrb61_0;
	wire w_dff_A_16ubPdRp1_0;
	wire w_dff_A_6Y58dUmr3_0;
	wire w_dff_A_IB8T7nYI1_0;
	wire w_dff_A_QpC3Hlss6_0;
	wire w_dff_A_3a83FO075_2;
	wire w_dff_A_R5ZzPwYw2_0;
	wire w_dff_A_unp3g2o18_0;
	wire w_dff_A_eYMK1qX39_0;
	wire w_dff_A_EaUr1SQN4_0;
	wire w_dff_A_NuzNO3OM4_0;
	wire w_dff_A_sfNFdMeh4_0;
	wire w_dff_A_3j91GzBb3_0;
	wire w_dff_A_N2MMRaGm8_0;
	wire w_dff_A_DZP6L6OB8_0;
	wire w_dff_A_pk7boYRo2_0;
	wire w_dff_A_3qZArAa61_0;
	wire w_dff_A_tDox3vvh5_0;
	wire w_dff_A_cNGGygDf1_0;
	wire w_dff_A_IGh0fp031_0;
	wire w_dff_A_WdwOJxi03_0;
	wire w_dff_A_NL3YWKon8_0;
	wire w_dff_A_gjwROSFG1_0;
	wire w_dff_A_4JmmDfE36_0;
	wire w_dff_A_WeoA5Rhf4_0;
	wire w_dff_A_loOnmAaY9_0;
	wire w_dff_A_YSxOoQvQ5_0;
	wire w_dff_A_lHSMrh6f6_0;
	wire w_dff_A_M8U3bskl4_0;
	wire w_dff_A_87QjXuSx7_0;
	wire w_dff_A_59sXhw6V9_0;
	wire w_dff_A_jpEupxkm3_0;
	wire w_dff_A_4PHBpZHu2_0;
	wire w_dff_A_VTL1HRAQ7_0;
	wire w_dff_A_t9adHGTj8_0;
	wire w_dff_A_i9JuflxC9_0;
	wire w_dff_A_PE6HJHdD0_0;
	wire w_dff_A_K49rF0yR2_0;
	wire w_dff_A_d0fHLS2q5_0;
	wire w_dff_A_MDIZ812e6_0;
	wire w_dff_A_sG4CTWPm4_0;
	wire w_dff_A_7xy2MAdt6_0;
	wire w_dff_A_e3Ng8x4E9_0;
	wire w_dff_A_edfSKao57_0;
	wire w_dff_A_83GvkYMm0_0;
	wire w_dff_A_f7suxt9F0_0;
	wire w_dff_A_owo9Ua9h9_0;
	wire w_dff_A_RwQSpl3F0_0;
	wire w_dff_A_sveZIsL14_0;
	wire w_dff_A_vwk37Yfm0_0;
	wire w_dff_A_7bz1RmbR8_0;
	wire w_dff_A_GIx2hT7U5_0;
	wire w_dff_A_1bKXmKbl0_0;
	wire w_dff_A_a9df2deA1_0;
	wire w_dff_A_4DD8ByeP8_0;
	wire w_dff_A_HvTO4E3w0_0;
	wire w_dff_A_i6CM3pXk4_0;
	wire w_dff_A_Zwph8O7S6_0;
	wire w_dff_A_4KREGJ5L7_0;
	wire w_dff_A_nFH0Xs6i1_0;
	wire w_dff_A_CrnPe1sW4_0;
	wire w_dff_A_ABcuLraL3_0;
	wire w_dff_A_msE5VSQQ4_0;
	wire w_dff_A_tjiL7swM1_0;
	wire w_dff_A_Urgu16Ef1_0;
	wire w_dff_A_RceBeY541_0;
	wire w_dff_A_IvFCHQvF9_0;
	wire w_dff_A_k891ORud8_0;
	wire w_dff_A_kz74VQLS6_0;
	wire w_dff_A_fqgSZzc77_0;
	wire w_dff_A_fafwZQnB2_0;
	wire w_dff_A_tiMs8Q3l6_0;
	wire w_dff_A_ogkJcjLT2_0;
	wire w_dff_A_C4X5lUbO2_0;
	wire w_dff_A_rNeKw7dI1_0;
	wire w_dff_A_8UcDCQ3i0_0;
	wire w_dff_A_E8tb1b9J8_0;
	wire w_dff_A_xndHYYXf6_0;
	wire w_dff_A_gUB4rCDK7_0;
	wire w_dff_A_tptklpjh5_0;
	wire w_dff_A_Jn8tbMwm5_0;
	wire w_dff_A_w2Ir4HAT0_0;
	wire w_dff_A_wGQeSFoD1_0;
	wire w_dff_A_wxSmVvdS0_0;
	wire w_dff_A_b6tAiDf00_0;
	wire w_dff_A_CHbzrRqv8_0;
	wire w_dff_A_fvvU2Bu84_0;
	wire w_dff_A_toWNEzfK3_0;
	wire w_dff_A_fPSmFcHY0_0;
	wire w_dff_A_7BnloomA7_0;
	wire w_dff_A_eUc7EgCD2_0;
	wire w_dff_A_pNNbcazj4_0;
	wire w_dff_A_YkKEgnKf8_0;
	wire w_dff_A_dKuJHMS67_0;
	wire w_dff_A_zCf0S6xz3_0;
	wire w_dff_A_5IgKgJGL1_0;
	wire w_dff_A_AOmInIwT4_0;
	wire w_dff_A_BX8cZWal2_0;
	wire w_dff_A_8zXJQ6Xx0_0;
	wire w_dff_A_iKuApldO0_0;
	wire w_dff_A_VBo9wto11_0;
	wire w_dff_A_rLAOYLtl7_0;
	wire w_dff_A_vnaebWSB6_0;
	wire w_dff_A_PQ6lY9By3_0;
	wire w_dff_A_IbySE8iU2_0;
	wire w_dff_A_DjASBRg76_0;
	wire w_dff_A_a6Yv4szI3_0;
	wire w_dff_A_Z7QZXcGI3_0;
	wire w_dff_A_ijbCtb7n5_0;
	wire w_dff_A_vGTkiiCQ3_0;
	wire w_dff_A_Fh9HDm058_0;
	wire w_dff_A_b9HBXwYE4_0;
	wire w_dff_A_pR7WgH8F8_0;
	wire w_dff_A_HWlffA8n1_0;
	wire w_dff_A_V2ySCPy10_0;
	wire w_dff_A_d1KRSa3g7_0;
	wire w_dff_A_V3pZY9iN1_0;
	wire w_dff_A_LnRVlKwa4_2;
	wire w_dff_A_GK17Zi180_0;
	wire w_dff_A_lW9ue4Dn2_0;
	wire w_dff_A_BE9RXxIO3_0;
	wire w_dff_A_ixFFjpir3_0;
	wire w_dff_A_AJc7r0aX4_0;
	wire w_dff_A_uEnheoL41_0;
	wire w_dff_A_daE6IegH4_0;
	wire w_dff_A_vpGSQ5t40_0;
	wire w_dff_A_06lDjxKk2_0;
	wire w_dff_A_QeflJm1n3_0;
	wire w_dff_A_Jz3tUiPJ3_0;
	wire w_dff_A_vVpFV9RF8_0;
	wire w_dff_A_iUb9M4Mt3_0;
	wire w_dff_A_UpoWBSax6_0;
	wire w_dff_A_NAlYSviQ2_0;
	wire w_dff_A_DxhC7mnd2_0;
	wire w_dff_A_cUSAUAH70_0;
	wire w_dff_A_Q9WX1Wb54_0;
	wire w_dff_A_GfLPjbmh9_0;
	wire w_dff_A_gSi30ZFL0_0;
	wire w_dff_A_BqiiYC0T5_0;
	wire w_dff_A_YzG78xio8_0;
	wire w_dff_A_VLOdgHGE5_0;
	wire w_dff_A_dCxFqYyP6_0;
	wire w_dff_A_BMzsJ6o49_0;
	wire w_dff_A_gIkgkHOE3_0;
	wire w_dff_A_38zmTKvG5_0;
	wire w_dff_A_AQbHBeld3_0;
	wire w_dff_A_utVQxiDS8_0;
	wire w_dff_A_8GKWIRTR2_0;
	wire w_dff_A_JccYcWe10_0;
	wire w_dff_A_JFnIfDDo6_0;
	wire w_dff_A_0npYbGSR7_0;
	wire w_dff_A_E3ewEzc74_0;
	wire w_dff_A_z2wogqZx3_0;
	wire w_dff_A_zefGtloA3_0;
	wire w_dff_A_jxbUBYPm1_0;
	wire w_dff_A_qSkxmWZR6_0;
	wire w_dff_A_RijoFnLp3_0;
	wire w_dff_A_XFr3uI0x3_0;
	wire w_dff_A_crkcGPVa3_0;
	wire w_dff_A_wmX7xsHM9_0;
	wire w_dff_A_6NvJomrV2_0;
	wire w_dff_A_VGtyecpn9_0;
	wire w_dff_A_MC0aPK002_0;
	wire w_dff_A_QsANbYHm3_0;
	wire w_dff_A_FvPki2c32_0;
	wire w_dff_A_i3SnkOgy5_0;
	wire w_dff_A_MUwsc3Zd2_0;
	wire w_dff_A_aQ2v3rbt2_0;
	wire w_dff_A_azkOg4LF7_0;
	wire w_dff_A_dS4JQigv7_0;
	wire w_dff_A_bRfeQZ0Q2_0;
	wire w_dff_A_3AuhCwAT9_0;
	wire w_dff_A_2KtKK2LF4_0;
	wire w_dff_A_mFvcxgRC2_0;
	wire w_dff_A_Xub2dLhQ8_0;
	wire w_dff_A_S9fstQr57_0;
	wire w_dff_A_EbOiH5BD5_0;
	wire w_dff_A_DViXWFGQ6_0;
	wire w_dff_A_N9AWNA2D5_0;
	wire w_dff_A_xi5hklZm5_0;
	wire w_dff_A_jZbA6zbg0_0;
	wire w_dff_A_sPo61Znb1_0;
	wire w_dff_A_IZ3BHVys4_0;
	wire w_dff_A_fshhcu145_0;
	wire w_dff_A_o8F1Q50S3_0;
	wire w_dff_A_azSwqbDW3_0;
	wire w_dff_A_jXDBjFuD2_0;
	wire w_dff_A_9EwgyWNC7_0;
	wire w_dff_A_gNkFYLLe6_0;
	wire w_dff_A_Dkc77BML4_0;
	wire w_dff_A_zVH8nU5U0_0;
	wire w_dff_A_MeA5eeRx0_0;
	wire w_dff_A_TcuLzh6s8_0;
	wire w_dff_A_nkMtUgND0_0;
	wire w_dff_A_oMBxkO476_0;
	wire w_dff_A_TYV4Z4B59_0;
	wire w_dff_A_M8y88Keo2_0;
	wire w_dff_A_wfUlKs3q1_0;
	wire w_dff_A_Z1NBHCMx2_0;
	wire w_dff_A_CBSOZ4se8_0;
	wire w_dff_A_CJCdGsZp1_0;
	wire w_dff_A_yfK9XDiI3_0;
	wire w_dff_A_xsbLQR2Z2_0;
	wire w_dff_A_afvFzpEu6_0;
	wire w_dff_A_8gKV97629_0;
	wire w_dff_A_4B0Q3ecX3_0;
	wire w_dff_A_McgJoamV3_0;
	wire w_dff_A_nWNxZivz4_0;
	wire w_dff_A_pjIBkap30_0;
	wire w_dff_A_Tv38rjXd5_0;
	wire w_dff_A_BbUfIVL53_0;
	wire w_dff_A_Dpw7lItZ4_0;
	wire w_dff_A_LvQWLnqK0_0;
	wire w_dff_A_pe22L4Xn7_0;
	wire w_dff_A_cfbyEwWr9_0;
	wire w_dff_A_VDMuFJSj8_0;
	wire w_dff_A_pOvi5AFl4_0;
	wire w_dff_A_aenLQ3jJ3_0;
	wire w_dff_A_E53xgmrV7_0;
	wire w_dff_A_H3iOXkfp6_0;
	wire w_dff_A_gN7IGKPd0_0;
	wire w_dff_A_Jt9BIdY34_0;
	wire w_dff_A_eVtOGUf78_0;
	wire w_dff_A_8bU3y6LR7_0;
	wire w_dff_A_WdVxd6TF5_0;
	wire w_dff_A_TlbkNLvE8_0;
	wire w_dff_A_XhSVAIJU8_0;
	wire w_dff_A_bMqwp1pC8_0;
	wire w_dff_A_xWMjmKJE2_2;
	wire w_dff_A_DkJMFBsl0_0;
	wire w_dff_A_eRpe2XwF9_0;
	wire w_dff_A_xYvshyNj1_0;
	wire w_dff_A_7L2wVWA19_0;
	wire w_dff_A_ntlnEkbs6_0;
	wire w_dff_A_YhBG0bmk5_0;
	wire w_dff_A_L9buB5Kh1_0;
	wire w_dff_A_m7YZYDBO0_0;
	wire w_dff_A_mdTfVhnM0_0;
	wire w_dff_A_dGB1DOfZ8_0;
	wire w_dff_A_j7Jxdgcg1_0;
	wire w_dff_A_VsohchKp2_0;
	wire w_dff_A_nm58TXz85_0;
	wire w_dff_A_6V0Sn0jg2_0;
	wire w_dff_A_yTKuAOOy3_0;
	wire w_dff_A_YuarT5dq3_0;
	wire w_dff_A_ypgxAohj8_0;
	wire w_dff_A_Cj4NbuNv3_0;
	wire w_dff_A_obf4KN2F3_0;
	wire w_dff_A_DepMQ3AP1_0;
	wire w_dff_A_54Ip8c1M8_0;
	wire w_dff_A_VafUtmqL6_0;
	wire w_dff_A_EwmlLQ6J8_0;
	wire w_dff_A_OMJ54ela6_0;
	wire w_dff_A_dmZJhJio1_0;
	wire w_dff_A_MTfHFV5n7_0;
	wire w_dff_A_HYYEK37L1_0;
	wire w_dff_A_vQ5WQZWB1_0;
	wire w_dff_A_rerBWFOs2_0;
	wire w_dff_A_JTqmsg9W8_0;
	wire w_dff_A_olKsJiUt0_0;
	wire w_dff_A_zhWekP025_0;
	wire w_dff_A_Xo1T2vJN0_0;
	wire w_dff_A_IUeXKzG53_0;
	wire w_dff_A_bWo59w982_0;
	wire w_dff_A_V6IQTE7s5_0;
	wire w_dff_A_d29VOzQS2_0;
	wire w_dff_A_g0NGThwQ6_0;
	wire w_dff_A_5IJPJmME5_0;
	wire w_dff_A_n3zITi9s8_0;
	wire w_dff_A_NG8jV5401_0;
	wire w_dff_A_bm2zZj0w4_0;
	wire w_dff_A_sbe9cv5T4_0;
	wire w_dff_A_WuyrlZ9q5_0;
	wire w_dff_A_NnwocXyi6_0;
	wire w_dff_A_U5PCJfn73_0;
	wire w_dff_A_YM0Hm7P92_0;
	wire w_dff_A_pzdTgPyN8_0;
	wire w_dff_A_5p6oRS8A0_0;
	wire w_dff_A_ozu1WvW45_0;
	wire w_dff_A_DvLvGVYE7_0;
	wire w_dff_A_kw1oR4ST3_0;
	wire w_dff_A_0NnmIXzU9_0;
	wire w_dff_A_oVjXKx4p9_0;
	wire w_dff_A_X3R2WtyE0_0;
	wire w_dff_A_Ir5YRAR96_0;
	wire w_dff_A_02kA5U2F1_0;
	wire w_dff_A_Z5HPi5Ou3_0;
	wire w_dff_A_FDiGOMEP9_0;
	wire w_dff_A_ElnAZ9DI8_0;
	wire w_dff_A_By2I0aJz1_0;
	wire w_dff_A_PASuZudb7_0;
	wire w_dff_A_E3JSNpSC3_0;
	wire w_dff_A_5bCIY7b58_0;
	wire w_dff_A_ZoejADoS4_0;
	wire w_dff_A_8DNFPTKt0_0;
	wire w_dff_A_jnB6bsRC0_0;
	wire w_dff_A_sbXDQhRO6_0;
	wire w_dff_A_oFQ072T27_0;
	wire w_dff_A_bLN9Z6Uf8_0;
	wire w_dff_A_zjLxCi0u5_0;
	wire w_dff_A_r9vIrRWV2_0;
	wire w_dff_A_zPvoC2co9_0;
	wire w_dff_A_lVeMbgJN4_0;
	wire w_dff_A_XvciFmFD8_0;
	wire w_dff_A_lPrlWIuJ9_0;
	wire w_dff_A_IasE0Rks4_0;
	wire w_dff_A_VWjgA6Ef2_0;
	wire w_dff_A_DbaijFgF9_0;
	wire w_dff_A_H6dru41O1_0;
	wire w_dff_A_3GNLmASH0_0;
	wire w_dff_A_Q2SslOAA9_0;
	wire w_dff_A_vKmCJMEw4_0;
	wire w_dff_A_q8dPJcMt0_0;
	wire w_dff_A_OvWTKkgz4_0;
	wire w_dff_A_WTyIX9jb5_0;
	wire w_dff_A_OADpagla0_0;
	wire w_dff_A_FUwEQ77B5_0;
	wire w_dff_A_pX6Q9gKC1_0;
	wire w_dff_A_Gjdp805S9_0;
	wire w_dff_A_LniBg7fT7_0;
	wire w_dff_A_JaJrjXgB0_0;
	wire w_dff_A_qF9wrIKC8_0;
	wire w_dff_A_kEawaRxa6_0;
	wire w_dff_A_XZr9GQfw1_0;
	wire w_dff_A_jpdcxZII7_0;
	wire w_dff_A_rqyXRseC1_0;
	wire w_dff_A_EVc1WssU0_0;
	wire w_dff_A_PmvkQFem2_0;
	wire w_dff_A_9qVp0lul8_0;
	wire w_dff_A_WgOfwrNZ0_0;
	wire w_dff_A_EhHxeAZK8_0;
	wire w_dff_A_25Va3Ja75_0;
	wire w_dff_A_Awe5Cts26_0;
	wire w_dff_A_uNrlZAZy5_0;
	wire w_dff_A_qWAggIwb1_0;
	wire w_dff_A_UxmRffia0_0;
	wire w_dff_A_v0QMzmHJ8_0;
	wire w_dff_A_1VMuFBuy4_0;
	wire w_dff_A_0NVR8Dal9_2;
	wire w_dff_A_TOmvvoze0_0;
	wire w_dff_A_TJfhYb0O1_0;
	wire w_dff_A_40TqYhct7_0;
	wire w_dff_A_Skvnf2ON2_0;
	wire w_dff_A_nO7DapF13_0;
	wire w_dff_A_8SgC1x9o9_0;
	wire w_dff_A_XFjIpT4g5_0;
	wire w_dff_A_CHOiVaJH3_0;
	wire w_dff_A_EQ8jbN8w5_0;
	wire w_dff_A_P37psMpY6_0;
	wire w_dff_A_753iWZkq8_0;
	wire w_dff_A_Ary1l48t2_0;
	wire w_dff_A_feVFlSEw9_0;
	wire w_dff_A_ISOWXJsA6_0;
	wire w_dff_A_GHdujyMQ9_0;
	wire w_dff_A_96SLxyII2_0;
	wire w_dff_A_GjciuaJ36_0;
	wire w_dff_A_3l9Pyy6i2_0;
	wire w_dff_A_hyth8iQW3_0;
	wire w_dff_A_5oR0vOOk1_0;
	wire w_dff_A_nV2GqiOP5_0;
	wire w_dff_A_hzttibKQ1_0;
	wire w_dff_A_imLKk0GV8_0;
	wire w_dff_A_VVAacT5S3_0;
	wire w_dff_A_vhxvB4Ou2_0;
	wire w_dff_A_sDNlSzfV3_0;
	wire w_dff_A_elwENFas5_0;
	wire w_dff_A_NPrINVDs1_0;
	wire w_dff_A_pmABDIji3_0;
	wire w_dff_A_liuXLDjP6_0;
	wire w_dff_A_BdY8vhzM2_0;
	wire w_dff_A_PyFFHFsP3_0;
	wire w_dff_A_7fXEossO1_0;
	wire w_dff_A_pIAhj8wx5_0;
	wire w_dff_A_RlDydzZl0_0;
	wire w_dff_A_KS40lmps3_0;
	wire w_dff_A_lCu3HYrF7_0;
	wire w_dff_A_RboOhAq06_0;
	wire w_dff_A_lJOf4rp12_0;
	wire w_dff_A_ay8oj7dI7_0;
	wire w_dff_A_1lKNpT6U8_0;
	wire w_dff_A_Zgo8m8nF6_0;
	wire w_dff_A_WlivYmsQ1_0;
	wire w_dff_A_rWIXssFJ6_0;
	wire w_dff_A_O5Joij324_0;
	wire w_dff_A_joFGlk3w6_0;
	wire w_dff_A_D4Z40p0y1_0;
	wire w_dff_A_bVLZghZy9_0;
	wire w_dff_A_NNAFmcZQ7_0;
	wire w_dff_A_orrABZaF8_0;
	wire w_dff_A_Z6bh4OCV3_0;
	wire w_dff_A_rMCwQX3i9_0;
	wire w_dff_A_W8z0B9583_0;
	wire w_dff_A_6jgMqxPI5_0;
	wire w_dff_A_if9xx1hj8_0;
	wire w_dff_A_u5eysuuu2_0;
	wire w_dff_A_o4m5kJR06_0;
	wire w_dff_A_2UwW5H9A9_0;
	wire w_dff_A_V5watVz60_0;
	wire w_dff_A_VZO3lMIw3_0;
	wire w_dff_A_ItVFv0Rj3_0;
	wire w_dff_A_3yisev2b6_0;
	wire w_dff_A_KBTOBMpK8_0;
	wire w_dff_A_c9kv7l3X8_0;
	wire w_dff_A_ubitWyl53_0;
	wire w_dff_A_O8refhWl5_0;
	wire w_dff_A_EIX1avql9_0;
	wire w_dff_A_xfh00RZ62_0;
	wire w_dff_A_oK5ygvzo9_0;
	wire w_dff_A_7v9Wf43s3_0;
	wire w_dff_A_zAzllwME4_0;
	wire w_dff_A_Z4izq7vp3_0;
	wire w_dff_A_zQu47Bh95_0;
	wire w_dff_A_SdGxpUpS2_0;
	wire w_dff_A_QumTBtFd0_0;
	wire w_dff_A_Y61zjZ820_0;
	wire w_dff_A_TWfwnIWv2_0;
	wire w_dff_A_HMKdSwET0_0;
	wire w_dff_A_vx4Y2RsJ8_0;
	wire w_dff_A_AQ955nqT1_0;
	wire w_dff_A_srhVHj253_0;
	wire w_dff_A_hbHulm8i7_0;
	wire w_dff_A_c55O5gyO6_0;
	wire w_dff_A_Cg7tF7AY1_0;
	wire w_dff_A_KgTGfBXg1_0;
	wire w_dff_A_5orPkeyk6_0;
	wire w_dff_A_AReFv5yH3_0;
	wire w_dff_A_UD8aM2XE4_0;
	wire w_dff_A_4jtmBBXC2_0;
	wire w_dff_A_oXPoMipA6_0;
	wire w_dff_A_Axfa65bU2_0;
	wire w_dff_A_WsrByzpk8_0;
	wire w_dff_A_uDueegk10_0;
	wire w_dff_A_lpwNtV4M6_0;
	wire w_dff_A_aK4I4rg72_0;
	wire w_dff_A_ujGyJ2Zj2_0;
	wire w_dff_A_r8ob65RH6_0;
	wire w_dff_A_TlFtjFoC9_0;
	wire w_dff_A_LxbOVs2i8_0;
	wire w_dff_A_2JmFVYJO4_0;
	wire w_dff_A_WcGcB9Zg8_0;
	wire w_dff_A_yMd3x3Gg2_0;
	wire w_dff_A_N5rLyz2h2_0;
	wire w_dff_A_b718xl0k7_0;
	wire w_dff_A_yBtdBJDA7_0;
	wire w_dff_A_BUXDYlMr2_0;
	wire w_dff_A_EKQCWszx3_0;
	wire w_dff_A_1sh2seEG3_0;
	wire w_dff_A_Bp4ITOiF1_2;
	wire w_dff_A_jvMhEy0w4_0;
	wire w_dff_A_puiqbAQJ0_0;
	wire w_dff_A_7OyJ08e32_0;
	wire w_dff_A_K9STGv5v8_0;
	wire w_dff_A_hc21YYuw8_0;
	wire w_dff_A_cK8QsWnQ6_0;
	wire w_dff_A_pqJQEVZj6_0;
	wire w_dff_A_Ve5qVmpp5_0;
	wire w_dff_A_m1YTylw03_0;
	wire w_dff_A_G9UEDFcj5_0;
	wire w_dff_A_hNduPF7j8_0;
	wire w_dff_A_Pcauvq6G2_0;
	wire w_dff_A_SeaAQBJf7_0;
	wire w_dff_A_rC2d8dQ85_0;
	wire w_dff_A_m8Ls7nyl0_0;
	wire w_dff_A_nqunztJd7_0;
	wire w_dff_A_m6k4tKll4_0;
	wire w_dff_A_yZxNEeS50_0;
	wire w_dff_A_DiBA0nA22_0;
	wire w_dff_A_XRJDC3bM5_0;
	wire w_dff_A_6CoknTaN6_0;
	wire w_dff_A_qTtQNH2l9_0;
	wire w_dff_A_30UqPXbZ2_0;
	wire w_dff_A_yzdiOauz1_0;
	wire w_dff_A_EGFE87tl0_0;
	wire w_dff_A_9GPV57NR4_0;
	wire w_dff_A_DCyGSsyH7_0;
	wire w_dff_A_J7K5a11g6_0;
	wire w_dff_A_JMdkWgCK1_0;
	wire w_dff_A_uQewDmo25_0;
	wire w_dff_A_ryzdhsBi2_0;
	wire w_dff_A_8sXp3TtB0_0;
	wire w_dff_A_iR67T7ca6_0;
	wire w_dff_A_5xm66XVX3_0;
	wire w_dff_A_L2ZpyEHo1_0;
	wire w_dff_A_J5C6ccrW5_0;
	wire w_dff_A_5OHCCJXW4_0;
	wire w_dff_A_7jfb9PZq1_0;
	wire w_dff_A_6IHFroO32_0;
	wire w_dff_A_4KQsbQom0_0;
	wire w_dff_A_6u5Tfjln1_0;
	wire w_dff_A_el4kXqXE6_0;
	wire w_dff_A_cTMl91cR1_0;
	wire w_dff_A_cdypmyVO9_0;
	wire w_dff_A_pg18zwdY9_0;
	wire w_dff_A_1RWiZGir1_0;
	wire w_dff_A_Yqaqp5Sk0_0;
	wire w_dff_A_1NlbArOp3_0;
	wire w_dff_A_VrEsTOyr9_0;
	wire w_dff_A_ij3597uh2_0;
	wire w_dff_A_LJrcCYPh6_0;
	wire w_dff_A_DUX6RMZG2_0;
	wire w_dff_A_ojpIOoXX6_0;
	wire w_dff_A_vCU6N5y40_0;
	wire w_dff_A_RgvLKoKM6_0;
	wire w_dff_A_g8Oi2kgh1_0;
	wire w_dff_A_nq8tb7K39_0;
	wire w_dff_A_ymovtUPC6_0;
	wire w_dff_A_gs5PXvFi5_0;
	wire w_dff_A_jouTIX5H4_0;
	wire w_dff_A_x00fOAnh5_0;
	wire w_dff_A_qwQib3Cc3_0;
	wire w_dff_A_3qVRkpfc8_0;
	wire w_dff_A_Djd8YOcl7_0;
	wire w_dff_A_7VSZ3mKu9_0;
	wire w_dff_A_0dP8F4lu6_0;
	wire w_dff_A_91S9c9Zg9_0;
	wire w_dff_A_scFQk9JK8_0;
	wire w_dff_A_38WyhstZ1_0;
	wire w_dff_A_EBnWxIgM4_0;
	wire w_dff_A_ZWMmg8BO0_0;
	wire w_dff_A_htbS2hd94_0;
	wire w_dff_A_B99DhVL18_0;
	wire w_dff_A_tq71fueL5_0;
	wire w_dff_A_BvJn82Ka8_0;
	wire w_dff_A_dEFFalXI5_0;
	wire w_dff_A_HC7qwXAW2_0;
	wire w_dff_A_GoYp4wky2_0;
	wire w_dff_A_LkpETppz5_0;
	wire w_dff_A_im0SIaHK6_0;
	wire w_dff_A_JnZ8YA4g9_0;
	wire w_dff_A_x7cJdx304_0;
	wire w_dff_A_weVeiff28_0;
	wire w_dff_A_v3kfMOSZ9_0;
	wire w_dff_A_VnI56l6h0_0;
	wire w_dff_A_TeswHEfx1_0;
	wire w_dff_A_3AM0Dykc1_0;
	wire w_dff_A_s8HIqjjZ9_0;
	wire w_dff_A_POiu1HVf9_0;
	wire w_dff_A_iD2LdKTY9_0;
	wire w_dff_A_7twhiEC58_0;
	wire w_dff_A_LfWqBv3s9_0;
	wire w_dff_A_NXIQYlJs4_0;
	wire w_dff_A_a7MwbyCF7_0;
	wire w_dff_A_qDSEG6sJ3_0;
	wire w_dff_A_R2IheBoY1_0;
	wire w_dff_A_qQ7bp2U02_0;
	wire w_dff_A_O8aSecI10_0;
	wire w_dff_A_2IWgLiww5_0;
	wire w_dff_A_1J7GUhos8_0;
	wire w_dff_A_Vbg1HtEm6_0;
	wire w_dff_A_8nBXHZve6_0;
	wire w_dff_A_IU0ZPoAs6_0;
	wire w_dff_A_45yVBPQW0_0;
	wire w_dff_A_VpiuJnI57_0;
	wire w_dff_A_pUbe4B8Y8_0;
	wire w_dff_A_vNKOVZgK2_0;
	wire w_dff_A_UvvGn9rX2_2;
	wire w_dff_A_8qGKI0RE0_0;
	wire w_dff_A_wZEg82Zz8_0;
	wire w_dff_A_mncMAK0q7_0;
	wire w_dff_A_lGkx8MuB8_0;
	wire w_dff_A_UIzdue6V0_0;
	wire w_dff_A_gLD5VCrV3_0;
	wire w_dff_A_gi3QU3QK9_0;
	wire w_dff_A_uLKcvOBz3_0;
	wire w_dff_A_4FTt6KVL3_0;
	wire w_dff_A_cVuFZiSb1_0;
	wire w_dff_A_IUTnGK8V2_0;
	wire w_dff_A_C3rhQdvh8_0;
	wire w_dff_A_8Zpd6bTi0_0;
	wire w_dff_A_h4tYWMGz7_0;
	wire w_dff_A_zubNrUp77_0;
	wire w_dff_A_FTlVkIkD3_0;
	wire w_dff_A_G5w5MOZf8_0;
	wire w_dff_A_iTK3nIE62_0;
	wire w_dff_A_w0SUd0hn6_0;
	wire w_dff_A_rr4a6nIK1_0;
	wire w_dff_A_JKnHVHzs3_0;
	wire w_dff_A_wT7ix1Px7_0;
	wire w_dff_A_QWACnWA75_0;
	wire w_dff_A_4elQGf0A5_0;
	wire w_dff_A_3EDvDyQh8_0;
	wire w_dff_A_4H2rBl3T7_0;
	wire w_dff_A_xaEvi8XX3_0;
	wire w_dff_A_AFE4a6kQ6_0;
	wire w_dff_A_4LrasE4A6_0;
	wire w_dff_A_AbuQaFpq7_0;
	wire w_dff_A_n6VYAloR6_0;
	wire w_dff_A_8C69epkn0_0;
	wire w_dff_A_6sCTv7YC9_0;
	wire w_dff_A_fvWKkfVd2_0;
	wire w_dff_A_Ps6BVgVk1_0;
	wire w_dff_A_EgPX5KQE0_0;
	wire w_dff_A_E7idzcbD4_0;
	wire w_dff_A_YZ4GsjPS8_0;
	wire w_dff_A_oH7Srzv53_0;
	wire w_dff_A_oxZpepLt2_0;
	wire w_dff_A_AmMRAFFv3_0;
	wire w_dff_A_mrpUq6Z82_0;
	wire w_dff_A_nRjCnJhy4_0;
	wire w_dff_A_n3nWSkU31_0;
	wire w_dff_A_rUNMMlhJ6_0;
	wire w_dff_A_SKnDkxxv6_0;
	wire w_dff_A_kAlCYB6y2_0;
	wire w_dff_A_Iqo0yklh8_0;
	wire w_dff_A_zMWDgjx27_0;
	wire w_dff_A_A0xLaTrl7_0;
	wire w_dff_A_HfKHwlDi5_0;
	wire w_dff_A_iDy24gsk4_0;
	wire w_dff_A_KfmWXslX6_0;
	wire w_dff_A_psXl9lrP8_0;
	wire w_dff_A_zvymgTgE2_0;
	wire w_dff_A_vm4ecouK0_0;
	wire w_dff_A_iFKsiyEU8_0;
	wire w_dff_A_tYvWPRNK3_0;
	wire w_dff_A_JahjJTGg0_0;
	wire w_dff_A_KwwizCYN5_0;
	wire w_dff_A_VOgAkZLq2_0;
	wire w_dff_A_ReRfwaqf9_0;
	wire w_dff_A_8lXzZFzS5_0;
	wire w_dff_A_kV1xeooL7_0;
	wire w_dff_A_Ug59nff18_0;
	wire w_dff_A_dljAIf8o1_0;
	wire w_dff_A_90qzFw8Z0_0;
	wire w_dff_A_cwBFOqul1_0;
	wire w_dff_A_qzhBt72e5_0;
	wire w_dff_A_jZLHhsEk4_0;
	wire w_dff_A_blQi8cHc4_0;
	wire w_dff_A_jR5xStDa0_0;
	wire w_dff_A_7dgUCgTw7_0;
	wire w_dff_A_CUVlYVML3_0;
	wire w_dff_A_g6xHjmhg3_0;
	wire w_dff_A_9wBVthNS5_0;
	wire w_dff_A_HWuUvGrz7_0;
	wire w_dff_A_KgwQzC4l7_0;
	wire w_dff_A_MHZkWSvw5_0;
	wire w_dff_A_UGOO3Pty4_0;
	wire w_dff_A_d8Av83NJ8_0;
	wire w_dff_A_rFsdYm2n6_0;
	wire w_dff_A_q1h92xXi7_0;
	wire w_dff_A_PqUmnpAS6_0;
	wire w_dff_A_gfZByBoH1_0;
	wire w_dff_A_Ze3Tq36k7_0;
	wire w_dff_A_Y9kY4jDj7_0;
	wire w_dff_A_Ta9DDjfu9_0;
	wire w_dff_A_FVsT9Xjy5_0;
	wire w_dff_A_B3dhimzS7_0;
	wire w_dff_A_k6yMc0VY5_0;
	wire w_dff_A_MRHDy74K5_0;
	wire w_dff_A_Jb5HEV1x5_0;
	wire w_dff_A_s3YVPPW46_0;
	wire w_dff_A_c6QvyV1A1_0;
	wire w_dff_A_atiBqafO7_0;
	wire w_dff_A_HFVpFWCU2_0;
	wire w_dff_A_viN9fqdh0_0;
	wire w_dff_A_4vPXxwVj5_0;
	wire w_dff_A_89L2DePF6_0;
	wire w_dff_A_WBX00K669_0;
	wire w_dff_A_FesiCaIL4_0;
	wire w_dff_A_nAGDZfi66_0;
	wire w_dff_A_KE3h50LS1_0;
	wire w_dff_A_bgW4cfhb5_0;
	wire w_dff_A_gT40v9Uv7_0;
	wire w_dff_A_lCHLbsXY9_2;
	wire w_dff_A_5pd3pxCd0_0;
	wire w_dff_A_izdYvg859_0;
	wire w_dff_A_Rnq3BGaR9_0;
	wire w_dff_A_xLXJHLSE6_0;
	wire w_dff_A_hmZBM0wt7_0;
	wire w_dff_A_csFKwb7y5_0;
	wire w_dff_A_b3HbDjZj1_0;
	wire w_dff_A_mtH9pT4D9_0;
	wire w_dff_A_DAeIv3Tt1_0;
	wire w_dff_A_1X6Bji5v1_0;
	wire w_dff_A_da7VZ5i46_0;
	wire w_dff_A_Efcg6eXY2_0;
	wire w_dff_A_igECOkQg8_0;
	wire w_dff_A_xT9E5Qgl6_0;
	wire w_dff_A_sWHgN6M18_0;
	wire w_dff_A_6x1RHjpr7_0;
	wire w_dff_A_u4KgYuln5_0;
	wire w_dff_A_txc1f1B08_0;
	wire w_dff_A_J1rU6GpA4_0;
	wire w_dff_A_PGt4U0254_0;
	wire w_dff_A_eRyfysyt0_0;
	wire w_dff_A_PMs9oPPU5_0;
	wire w_dff_A_S2133bGj5_0;
	wire w_dff_A_UXqeLZWi2_0;
	wire w_dff_A_OevOKfvM9_0;
	wire w_dff_A_WM6lGyIs4_0;
	wire w_dff_A_2ldw2KTm9_0;
	wire w_dff_A_3R25R7Af4_0;
	wire w_dff_A_J0OSiSBk0_0;
	wire w_dff_A_RyVAaV5H7_0;
	wire w_dff_A_KdelyN9K4_0;
	wire w_dff_A_KmxVKamR8_0;
	wire w_dff_A_u6FvbWQy9_0;
	wire w_dff_A_ejHZVtyW7_0;
	wire w_dff_A_Q2r438ol0_0;
	wire w_dff_A_RFrBKZ1D2_0;
	wire w_dff_A_3kqEJFzN1_0;
	wire w_dff_A_U2hHdySL3_0;
	wire w_dff_A_B185ummz5_0;
	wire w_dff_A_Vt4CpBhV9_0;
	wire w_dff_A_IWSCJtX40_0;
	wire w_dff_A_gk2j205J0_0;
	wire w_dff_A_a0GYr0En4_0;
	wire w_dff_A_v1KTRN0H7_0;
	wire w_dff_A_C0WmJupj1_0;
	wire w_dff_A_m1omsexu0_0;
	wire w_dff_A_UhxrpWp47_0;
	wire w_dff_A_42kPPQaw7_0;
	wire w_dff_A_IfHcsQ6I8_0;
	wire w_dff_A_hIWv5xfW4_0;
	wire w_dff_A_SDFz8boM9_0;
	wire w_dff_A_gjvaAsRC3_0;
	wire w_dff_A_RSnX1Ozu6_0;
	wire w_dff_A_FJ2goiww9_0;
	wire w_dff_A_kAO5oVl70_0;
	wire w_dff_A_VyA3rdJQ5_0;
	wire w_dff_A_RWsENUmU9_0;
	wire w_dff_A_1iGcRfvK9_0;
	wire w_dff_A_ewafylVO7_0;
	wire w_dff_A_bu0qEqds3_0;
	wire w_dff_A_83a87D6G6_0;
	wire w_dff_A_9jMDtlyG7_0;
	wire w_dff_A_j0h2hltR9_0;
	wire w_dff_A_dPTtqRAw3_0;
	wire w_dff_A_vTbSlqOB8_0;
	wire w_dff_A_tsBUC5qc9_0;
	wire w_dff_A_WbpGKj4t4_0;
	wire w_dff_A_ArDe8fKK7_0;
	wire w_dff_A_UNmXbe9h8_0;
	wire w_dff_A_9uWF6XgJ1_0;
	wire w_dff_A_ABs5pq959_0;
	wire w_dff_A_WGMF3nzx0_0;
	wire w_dff_A_IHkl6Zr74_0;
	wire w_dff_A_DN5ZxBeK5_0;
	wire w_dff_A_KhAGHMYt3_0;
	wire w_dff_A_FhHNseIR4_0;
	wire w_dff_A_vjBGIUKh4_0;
	wire w_dff_A_QHQv3pTk9_0;
	wire w_dff_A_ix0FDSO22_0;
	wire w_dff_A_QPBq49vp8_0;
	wire w_dff_A_Ok8pvOZ99_0;
	wire w_dff_A_RRr3kmrq1_0;
	wire w_dff_A_RCd0t5l57_0;
	wire w_dff_A_UfZNiuRo8_0;
	wire w_dff_A_ULDYjV6J5_0;
	wire w_dff_A_qO7GpZOl8_0;
	wire w_dff_A_fUmXCxD37_0;
	wire w_dff_A_8b28aMpw2_0;
	wire w_dff_A_hfGCvspW4_0;
	wire w_dff_A_8gZjpzUU4_0;
	wire w_dff_A_gKELwUX22_0;
	wire w_dff_A_PyKsbI6B2_0;
	wire w_dff_A_woH1tcJQ1_0;
	wire w_dff_A_7mvaKFp77_0;
	wire w_dff_A_eECTUFPl2_0;
	wire w_dff_A_HZ4hGMrp8_0;
	wire w_dff_A_XqSGPLTf6_0;
	wire w_dff_A_g7joznxS5_0;
	wire w_dff_A_kCotj0PF2_0;
	wire w_dff_A_oGC5CTXB7_0;
	wire w_dff_A_vuLBUkkB2_0;
	wire w_dff_A_galTre5O3_0;
	wire w_dff_A_tOPjkisW3_0;
	wire w_dff_A_d1ZSvvVt7_0;
	wire w_dff_A_ArwO2Kdi0_0;
	wire w_dff_A_bwlIPVrT6_2;
	wire w_dff_A_8FzXY3168_0;
	wire w_dff_A_A6vbtUuC7_0;
	wire w_dff_A_HM2WTPae1_0;
	wire w_dff_A_tyIBQehs4_0;
	wire w_dff_A_WlOGOG2d7_0;
	wire w_dff_A_hWB6KHfc7_0;
	wire w_dff_A_FAqR5UKH3_0;
	wire w_dff_A_vmz8Sacf3_0;
	wire w_dff_A_5DryWorU4_0;
	wire w_dff_A_kdmAfC7Z2_0;
	wire w_dff_A_PDTG4Lyu3_0;
	wire w_dff_A_GVbLDY1S5_0;
	wire w_dff_A_8KN4RRSD1_0;
	wire w_dff_A_f4brMCd86_0;
	wire w_dff_A_DEthHJvO7_0;
	wire w_dff_A_OhHAtnqY5_0;
	wire w_dff_A_cS62FSNa3_0;
	wire w_dff_A_479AbONi3_0;
	wire w_dff_A_pJXoKSvf1_0;
	wire w_dff_A_PTaAt3HY8_0;
	wire w_dff_A_C9sVdWhH5_0;
	wire w_dff_A_n8rPqkCb9_0;
	wire w_dff_A_qiCgNgwo3_0;
	wire w_dff_A_5TEwIZ6n8_0;
	wire w_dff_A_0LSKHq6e7_0;
	wire w_dff_A_fWBXEgeT7_0;
	wire w_dff_A_OAO0GRfY1_0;
	wire w_dff_A_uHDcmhm02_0;
	wire w_dff_A_2E8jZQuZ7_0;
	wire w_dff_A_2rVGI5XN3_0;
	wire w_dff_A_iu0JGMa19_0;
	wire w_dff_A_Fjw2Ypi53_0;
	wire w_dff_A_SLd5HLax5_0;
	wire w_dff_A_kQ2WuSwu9_0;
	wire w_dff_A_RgpQF4Kq8_0;
	wire w_dff_A_zETwFmI94_0;
	wire w_dff_A_0D30lWH01_0;
	wire w_dff_A_IfvT1kZq6_0;
	wire w_dff_A_pqMGsv5r8_0;
	wire w_dff_A_lkIyvNq03_0;
	wire w_dff_A_4Fxy4zKq1_0;
	wire w_dff_A_TE1MwDsW3_0;
	wire w_dff_A_okusVvoe8_0;
	wire w_dff_A_O0H93BUF7_0;
	wire w_dff_A_9FL475L33_0;
	wire w_dff_A_giBoKNlS9_0;
	wire w_dff_A_M5zGQe7H2_0;
	wire w_dff_A_C8dMslQp0_0;
	wire w_dff_A_SSgz4MOR5_0;
	wire w_dff_A_BXKlKgrx6_0;
	wire w_dff_A_P9FQj71Z8_0;
	wire w_dff_A_Yw7D2DO90_0;
	wire w_dff_A_Ooc3W83r8_0;
	wire w_dff_A_YKupuHdO1_0;
	wire w_dff_A_O4BJ1L9Y0_0;
	wire w_dff_A_IAQ9ylwU0_0;
	wire w_dff_A_g58qylQv7_0;
	wire w_dff_A_cmqRq9ll9_0;
	wire w_dff_A_fJqLOD2P9_0;
	wire w_dff_A_biog2G9A6_0;
	wire w_dff_A_6sZx2PC66_0;
	wire w_dff_A_x1WcYlPQ0_0;
	wire w_dff_A_O4guebVd9_0;
	wire w_dff_A_9DOVMoJo9_0;
	wire w_dff_A_NFWUJqb86_0;
	wire w_dff_A_wHv1RlhK1_0;
	wire w_dff_A_ZIxYcDhK3_0;
	wire w_dff_A_LCoKL0Ld5_0;
	wire w_dff_A_kXkge0Qz3_0;
	wire w_dff_A_ZFNKyjxw1_0;
	wire w_dff_A_r4XED1Wz4_0;
	wire w_dff_A_QdUAVXYu7_0;
	wire w_dff_A_KtnQqaVm6_0;
	wire w_dff_A_m6aHDcbn9_0;
	wire w_dff_A_De8Moz1T5_0;
	wire w_dff_A_PanXAJOA6_0;
	wire w_dff_A_y90BUh0h2_0;
	wire w_dff_A_hF4kyPRr1_0;
	wire w_dff_A_4MD2y8Ik0_0;
	wire w_dff_A_EjK1JFvn1_0;
	wire w_dff_A_GDqZ6AHT0_0;
	wire w_dff_A_rA8UT6oB1_0;
	wire w_dff_A_GHux770v4_0;
	wire w_dff_A_fUOA2d2I4_0;
	wire w_dff_A_3rFeyepe7_0;
	wire w_dff_A_QxMgPICO1_0;
	wire w_dff_A_1L4XGj2E6_0;
	wire w_dff_A_lzFKR7sV0_0;
	wire w_dff_A_I3oSY4fj2_0;
	wire w_dff_A_JQcrzHkQ3_0;
	wire w_dff_A_pUp2hiZi9_0;
	wire w_dff_A_hEbO0vre1_0;
	wire w_dff_A_xUjPFYO97_0;
	wire w_dff_A_9N7vfbIU5_0;
	wire w_dff_A_1BnerdXf2_0;
	wire w_dff_A_pgrUrioX3_0;
	wire w_dff_A_Xjqc7oiz3_0;
	wire w_dff_A_RzMdwBna3_0;
	wire w_dff_A_d0zoPeGb8_0;
	wire w_dff_A_kPT4fht42_0;
	wire w_dff_A_a2phIt3T8_0;
	wire w_dff_A_g3gFHxxZ7_0;
	wire w_dff_A_gR2LLfUO8_0;
	wire w_dff_A_akm2I8wf7_0;
	wire w_dff_A_SzoSoT3h7_2;
	wire w_dff_A_LXu8MeCK4_0;
	wire w_dff_A_PVWHarOq6_0;
	wire w_dff_A_vifkcGun8_0;
	wire w_dff_A_MdeSnA3n3_0;
	wire w_dff_A_vqkNSrdK9_0;
	wire w_dff_A_mF9lCjQ08_0;
	wire w_dff_A_Iyd8w0tZ1_0;
	wire w_dff_A_TeFjgyX76_0;
	wire w_dff_A_YHZd3Amb7_0;
	wire w_dff_A_GIadcR8T8_0;
	wire w_dff_A_dtlDCxQZ1_0;
	wire w_dff_A_xpG3ulbz0_0;
	wire w_dff_A_imuh9k5R6_0;
	wire w_dff_A_IfgThEwV6_0;
	wire w_dff_A_IRrpS1iv1_0;
	wire w_dff_A_jD2jZJ493_0;
	wire w_dff_A_p1HjCQLw3_0;
	wire w_dff_A_jCV2xufZ5_0;
	wire w_dff_A_qykpVwGV0_0;
	wire w_dff_A_qB5FPRrW5_0;
	wire w_dff_A_owfNYa9D9_0;
	wire w_dff_A_mIU6Bse73_0;
	wire w_dff_A_2DbPMeuB7_0;
	wire w_dff_A_bW4x1qXE8_0;
	wire w_dff_A_bY11Q5mg8_0;
	wire w_dff_A_BAEbRGrc1_0;
	wire w_dff_A_ASg1x7au3_0;
	wire w_dff_A_gDgu3THB4_0;
	wire w_dff_A_BDvUB8TI5_0;
	wire w_dff_A_jYfVz6oW2_0;
	wire w_dff_A_a8l5C6Ap1_0;
	wire w_dff_A_8R47zttB4_0;
	wire w_dff_A_G4aae9Zw2_0;
	wire w_dff_A_sW7Q7Knw0_0;
	wire w_dff_A_2JXXtMpv3_0;
	wire w_dff_A_kJ7juJXl2_0;
	wire w_dff_A_wxOnMeeI0_0;
	wire w_dff_A_ODt5AzzS7_0;
	wire w_dff_A_KcJqTdHP8_0;
	wire w_dff_A_kWPWQpGd3_0;
	wire w_dff_A_3TjJOnOC7_0;
	wire w_dff_A_sgXkth8x3_0;
	wire w_dff_A_7eD9rVRi0_0;
	wire w_dff_A_4cms8jLp0_0;
	wire w_dff_A_KWhctdji3_0;
	wire w_dff_A_QBDjBpOu8_0;
	wire w_dff_A_TgFxIp3s3_0;
	wire w_dff_A_6iBUmoJf0_0;
	wire w_dff_A_aejISBg08_0;
	wire w_dff_A_uOcqpVc64_0;
	wire w_dff_A_ArBlX3jn0_0;
	wire w_dff_A_klpiuytj8_0;
	wire w_dff_A_o56JiOSW0_0;
	wire w_dff_A_gyPJsgey1_0;
	wire w_dff_A_kWZIIHBJ2_0;
	wire w_dff_A_IpEj3raU0_0;
	wire w_dff_A_YmNhCS0B9_0;
	wire w_dff_A_CCATSn5H4_0;
	wire w_dff_A_CGOYnW5O9_0;
	wire w_dff_A_7LiUCqHo5_0;
	wire w_dff_A_9sODmkT92_0;
	wire w_dff_A_7KUhGUFr0_0;
	wire w_dff_A_oi1zJ8CS5_0;
	wire w_dff_A_eKZGL1246_0;
	wire w_dff_A_FsmKzGuw4_0;
	wire w_dff_A_AFrjmDBM4_0;
	wire w_dff_A_Gw0mfJZS8_0;
	wire w_dff_A_6tpPbB2I3_0;
	wire w_dff_A_0lWJ2Xti3_0;
	wire w_dff_A_t4W4Gd1K1_0;
	wire w_dff_A_iyPVEQDl4_0;
	wire w_dff_A_QZ18hAHR0_0;
	wire w_dff_A_2DG7GwYF4_0;
	wire w_dff_A_VoWJFzLW5_0;
	wire w_dff_A_zkdlMpUx4_0;
	wire w_dff_A_3OQZIldj0_0;
	wire w_dff_A_4z0tI5rq0_0;
	wire w_dff_A_vPiJCUxB6_0;
	wire w_dff_A_funNv0lY2_0;
	wire w_dff_A_6M6BaDUw3_0;
	wire w_dff_A_CoDM5QjP2_0;
	wire w_dff_A_EYDQ1SN71_0;
	wire w_dff_A_ekhQo3kf1_0;
	wire w_dff_A_RynvRZny4_0;
	wire w_dff_A_TKbnUnwF1_0;
	wire w_dff_A_WTAQeAF97_0;
	wire w_dff_A_mnZVhNVH6_0;
	wire w_dff_A_QQcMw8Fl8_0;
	wire w_dff_A_HTZAA6WZ7_0;
	wire w_dff_A_1OmNtLNt8_0;
	wire w_dff_A_8xAFlvmf0_0;
	wire w_dff_A_xWTpfVgj4_0;
	wire w_dff_A_GLwGk8Zm5_0;
	wire w_dff_A_UjABIs6o9_0;
	wire w_dff_A_jhWgGv0K1_0;
	wire w_dff_A_DWIOOwgf4_0;
	wire w_dff_A_wAvlJOGm1_0;
	wire w_dff_A_3DiWJpNI4_0;
	wire w_dff_A_Si5NIZHx2_0;
	wire w_dff_A_HHgAH7bn6_0;
	wire w_dff_A_fKfOJnKl3_0;
	wire w_dff_A_Aun1bA194_0;
	wire w_dff_A_VMJTXdB51_0;
	wire w_dff_A_ejqy7DXE0_2;
	wire w_dff_A_W9qGWd5L5_0;
	wire w_dff_A_ggFuGkP97_0;
	wire w_dff_A_BVcr5RcT9_0;
	wire w_dff_A_PNMtgzvZ3_0;
	wire w_dff_A_9EZohE6J0_0;
	wire w_dff_A_Y7RBP92s3_0;
	wire w_dff_A_lWHrxWO81_0;
	wire w_dff_A_1sFEfer31_0;
	wire w_dff_A_ViTw3MGF1_0;
	wire w_dff_A_kymaJul48_0;
	wire w_dff_A_fUzRDZZ14_0;
	wire w_dff_A_QK7TvgVu8_0;
	wire w_dff_A_KOdloJ791_0;
	wire w_dff_A_L7sNwnTe5_0;
	wire w_dff_A_MuG62oUz0_0;
	wire w_dff_A_dRlNogGM5_0;
	wire w_dff_A_X46SUInS2_0;
	wire w_dff_A_xZYRmbfw9_0;
	wire w_dff_A_LYTxWNRW4_0;
	wire w_dff_A_bf0aTqXI7_0;
	wire w_dff_A_aCxSvOX66_0;
	wire w_dff_A_cIsj3QxJ3_0;
	wire w_dff_A_J9hs0yzB5_0;
	wire w_dff_A_vQAFlWTx8_0;
	wire w_dff_A_m3L4hsq31_0;
	wire w_dff_A_KtCpX6E49_0;
	wire w_dff_A_Fx8sSX2J7_0;
	wire w_dff_A_0aKUwqfo4_0;
	wire w_dff_A_rUdDsgZT2_0;
	wire w_dff_A_ZzRGaad17_0;
	wire w_dff_A_hyzJehtM7_0;
	wire w_dff_A_FVIX3Ia43_0;
	wire w_dff_A_bI80vFUL4_0;
	wire w_dff_A_WwcYynn03_0;
	wire w_dff_A_3SeYvBSO4_0;
	wire w_dff_A_dvq20nJy5_0;
	wire w_dff_A_V0TiymFn5_0;
	wire w_dff_A_InSpKmGW0_0;
	wire w_dff_A_vKNoR8dw6_0;
	wire w_dff_A_bgz3aLVs5_0;
	wire w_dff_A_33If5CeM2_0;
	wire w_dff_A_Yl1H3zSP4_0;
	wire w_dff_A_YSGDg2aq6_0;
	wire w_dff_A_yRgScSfz9_0;
	wire w_dff_A_emNbOSB58_0;
	wire w_dff_A_0joguT0n8_0;
	wire w_dff_A_e95w1D3H2_0;
	wire w_dff_A_7oxaZ6G89_0;
	wire w_dff_A_PsMZRVYY6_0;
	wire w_dff_A_3jfRZvRo2_0;
	wire w_dff_A_L1gTztii4_0;
	wire w_dff_A_mZvLRIe05_0;
	wire w_dff_A_2zqT3RIj3_0;
	wire w_dff_A_bwyy7mFv5_0;
	wire w_dff_A_QiJKv5Qp0_0;
	wire w_dff_A_bc5x8CLy1_0;
	wire w_dff_A_CYhoSLiY4_0;
	wire w_dff_A_H1dQJ4ez0_0;
	wire w_dff_A_IFsKeohE3_0;
	wire w_dff_A_ouXkB9Sb2_0;
	wire w_dff_A_V0XTjOvB4_0;
	wire w_dff_A_k1r1iZuP7_0;
	wire w_dff_A_7RQ14DhJ7_0;
	wire w_dff_A_8iuAEy5I8_0;
	wire w_dff_A_RHyheddQ1_0;
	wire w_dff_A_e8wzgcAC0_0;
	wire w_dff_A_vkPOIoEu2_0;
	wire w_dff_A_LnAJKT816_0;
	wire w_dff_A_ZaC6eVBr4_0;
	wire w_dff_A_EWZwgFVi5_0;
	wire w_dff_A_DhLQcXRh7_0;
	wire w_dff_A_2V8rt1eX1_0;
	wire w_dff_A_98aflCDi5_0;
	wire w_dff_A_qf0SAwA50_0;
	wire w_dff_A_vtUIdmVH0_0;
	wire w_dff_A_4KwMGY9a7_0;
	wire w_dff_A_aBb5MOyb7_0;
	wire w_dff_A_DD5cBLyN5_0;
	wire w_dff_A_Lg4EKZAv1_0;
	wire w_dff_A_NkcCgnAP7_0;
	wire w_dff_A_uQb8QUWy7_0;
	wire w_dff_A_S4Zgh2Bs1_0;
	wire w_dff_A_K7UdTQ9A0_0;
	wire w_dff_A_HirujnNS7_0;
	wire w_dff_A_ZVRApH6F5_0;
	wire w_dff_A_UqiPodn99_0;
	wire w_dff_A_Isp1yFap2_0;
	wire w_dff_A_n6pbBf6Z1_0;
	wire w_dff_A_EH6GaQiO8_0;
	wire w_dff_A_B6MKY3l67_0;
	wire w_dff_A_Rxo852FK5_0;
	wire w_dff_A_2k5F1CB89_0;
	wire w_dff_A_tJBO9hAc8_0;
	wire w_dff_A_oNekGLhW2_0;
	wire w_dff_A_Ao97cxID1_0;
	wire w_dff_A_I8fmg2eM1_0;
	wire w_dff_A_Byqdnubd4_0;
	wire w_dff_A_jRUa5FoK4_0;
	wire w_dff_A_ymB7fdEt0_0;
	wire w_dff_A_uKaxxzL60_0;
	wire w_dff_A_yQiRHdtT6_0;
	wire w_dff_A_lRdahrlG0_0;
	wire w_dff_A_0nEZ1YGf2_2;
	wire w_dff_A_XpUQpVdN7_0;
	wire w_dff_A_5thKmnai7_0;
	wire w_dff_A_n8SdQJkF4_0;
	wire w_dff_A_z2uBN0HD1_0;
	wire w_dff_A_uZ0XBi0R4_0;
	wire w_dff_A_Piisp0vd7_0;
	wire w_dff_A_t59uKDX81_0;
	wire w_dff_A_cvH13HmV0_0;
	wire w_dff_A_G2JPCfLJ4_0;
	wire w_dff_A_LDlLZ7Ya8_0;
	wire w_dff_A_CZNR46Kc9_0;
	wire w_dff_A_JycQkhvU5_0;
	wire w_dff_A_ESgeG3L03_0;
	wire w_dff_A_lgBszO8L4_0;
	wire w_dff_A_qyI2Er4q2_0;
	wire w_dff_A_HTx9f88E5_0;
	wire w_dff_A_siduIdft4_0;
	wire w_dff_A_LcJTspSp3_0;
	wire w_dff_A_C3kAR2FE0_0;
	wire w_dff_A_Zz4CQQak3_0;
	wire w_dff_A_iuF9XDjk1_0;
	wire w_dff_A_AruhJiPA3_0;
	wire w_dff_A_9sxbnDaN2_0;
	wire w_dff_A_OyjrpZtk1_0;
	wire w_dff_A_QbxKWqba6_0;
	wire w_dff_A_Q9vYBh663_0;
	wire w_dff_A_2Hs9V9YX4_0;
	wire w_dff_A_K1c8lOqV3_0;
	wire w_dff_A_XQrGES744_0;
	wire w_dff_A_mOFz25wK9_0;
	wire w_dff_A_LiVm21O92_0;
	wire w_dff_A_E6f6xOtF7_0;
	wire w_dff_A_tS6CCnjV3_0;
	wire w_dff_A_XNF6ZSNS0_0;
	wire w_dff_A_fiiYCJKr0_0;
	wire w_dff_A_9eUdAo6S2_0;
	wire w_dff_A_0JQKAZh02_0;
	wire w_dff_A_8ToBNj5J8_0;
	wire w_dff_A_BVLiAXXL2_0;
	wire w_dff_A_CYUuieAQ3_0;
	wire w_dff_A_TqA6t0059_0;
	wire w_dff_A_sQrLNdjJ9_0;
	wire w_dff_A_ZaJ6jopY8_0;
	wire w_dff_A_VuPzxNaY5_0;
	wire w_dff_A_ciMS16dp8_0;
	wire w_dff_A_Az1NZDsQ0_0;
	wire w_dff_A_SNYxVHDd6_0;
	wire w_dff_A_fOppy9ci6_0;
	wire w_dff_A_PM4uTAe31_0;
	wire w_dff_A_KAdNvwF04_0;
	wire w_dff_A_pYFBSyyQ3_0;
	wire w_dff_A_gE1KLIn52_0;
	wire w_dff_A_j15LUhPb0_0;
	wire w_dff_A_IzFGJGlB4_0;
	wire w_dff_A_9ih4B6lu8_0;
	wire w_dff_A_4pfPp2v81_0;
	wire w_dff_A_4UTkAK6z4_0;
	wire w_dff_A_ac8uZy296_0;
	wire w_dff_A_lxtRVMAD0_0;
	wire w_dff_A_Sf8lL5I23_0;
	wire w_dff_A_kwuv0SpU5_0;
	wire w_dff_A_joiyyHKD8_0;
	wire w_dff_A_2KleqGgU8_0;
	wire w_dff_A_poGmEZQK4_0;
	wire w_dff_A_6QcNXvES6_0;
	wire w_dff_A_IxqDbUPP0_0;
	wire w_dff_A_ElvEYsr06_0;
	wire w_dff_A_b953PdWO9_0;
	wire w_dff_A_AfY7WRZe5_0;
	wire w_dff_A_4dCduNFl5_0;
	wire w_dff_A_r11WoBd07_0;
	wire w_dff_A_IcebyBVR6_0;
	wire w_dff_A_cw0ijJ1f5_0;
	wire w_dff_A_Wkt1B6bc8_0;
	wire w_dff_A_l7zRAedK6_0;
	wire w_dff_A_cRCBYTGX2_0;
	wire w_dff_A_6fQmR3Kw0_0;
	wire w_dff_A_pTfgEiJ99_0;
	wire w_dff_A_JkVtL0DQ6_0;
	wire w_dff_A_uJ4KZjgh4_0;
	wire w_dff_A_QrqrotYQ9_0;
	wire w_dff_A_i14hUG3K5_0;
	wire w_dff_A_TEveETai2_0;
	wire w_dff_A_k1wJ2nx67_0;
	wire w_dff_A_0HSHNax31_0;
	wire w_dff_A_dJYTji9n6_0;
	wire w_dff_A_ZCqFWlPC1_0;
	wire w_dff_A_g7sfD5oQ3_0;
	wire w_dff_A_N2RzlP2m1_0;
	wire w_dff_A_aEDIY8A09_0;
	wire w_dff_A_symwYzaY6_0;
	wire w_dff_A_Nlm5jXQU7_0;
	wire w_dff_A_bRV5paq16_0;
	wire w_dff_A_GvoORiBG0_0;
	wire w_dff_A_LZe8Cn5W9_0;
	wire w_dff_A_s4pctpVC2_0;
	wire w_dff_A_yyPkTCU93_0;
	wire w_dff_A_SesGA1bx1_0;
	wire w_dff_A_uEVqlit24_0;
	wire w_dff_A_W90yQBs47_0;
	wire w_dff_A_x3X9er1E3_0;
	wire w_dff_A_M4eemYt31_2;
	wire w_dff_A_AwhbLbvS6_0;
	wire w_dff_A_rSr6SRMx2_0;
	wire w_dff_A_SmA2fzwJ5_0;
	wire w_dff_A_5rHiVLHD0_0;
	wire w_dff_A_bmCnJbg39_0;
	wire w_dff_A_mPkeNnAl7_0;
	wire w_dff_A_ow920u5m8_0;
	wire w_dff_A_EIR3NQ3l0_0;
	wire w_dff_A_47tVZ46P3_0;
	wire w_dff_A_8DzQKIKq7_0;
	wire w_dff_A_IJqun7Xu4_0;
	wire w_dff_A_0bdPYpd87_0;
	wire w_dff_A_4iyrtd2z5_0;
	wire w_dff_A_aX7UIuPX4_0;
	wire w_dff_A_1gQezk1d7_0;
	wire w_dff_A_CbxhIpxn5_0;
	wire w_dff_A_wfJAe4av2_0;
	wire w_dff_A_UMDqXr348_0;
	wire w_dff_A_pr0ZCi2E3_0;
	wire w_dff_A_W0E2eudA5_0;
	wire w_dff_A_jvXVb8bu4_0;
	wire w_dff_A_A4t18bvA2_0;
	wire w_dff_A_NPMz15Gh0_0;
	wire w_dff_A_j3DzRLm82_0;
	wire w_dff_A_CRZMfwm49_0;
	wire w_dff_A_Jtu5BTpk1_0;
	wire w_dff_A_gBldQUzH8_0;
	wire w_dff_A_v7uE4mJ59_0;
	wire w_dff_A_Ep5WBgiY6_0;
	wire w_dff_A_IXnFGN1c5_0;
	wire w_dff_A_gkPPHvL01_0;
	wire w_dff_A_5IEqqgjo9_0;
	wire w_dff_A_qpDgwJBG4_0;
	wire w_dff_A_3Gxms4ll2_0;
	wire w_dff_A_jEq3sh0o6_0;
	wire w_dff_A_6DiZT4nb9_0;
	wire w_dff_A_lnjxgXyp8_0;
	wire w_dff_A_uIFJt6je6_0;
	wire w_dff_A_72ADBfXj2_0;
	wire w_dff_A_FsRRNwpR8_0;
	wire w_dff_A_lvE2aJxj2_0;
	wire w_dff_A_xxvSkDpq0_0;
	wire w_dff_A_BQ0CF9jx4_0;
	wire w_dff_A_VO8oeS5O6_0;
	wire w_dff_A_qYblETKR2_0;
	wire w_dff_A_h5e7WUCW0_0;
	wire w_dff_A_0YyHPbH77_0;
	wire w_dff_A_do74JSrz6_0;
	wire w_dff_A_H4O3llyJ9_0;
	wire w_dff_A_hjpWyEbc5_0;
	wire w_dff_A_qoroFDrB1_0;
	wire w_dff_A_teEdXXph2_0;
	wire w_dff_A_adhHJpla8_0;
	wire w_dff_A_68o9WCJt7_0;
	wire w_dff_A_5TlTkyEc5_0;
	wire w_dff_A_VMd8OwCf6_0;
	wire w_dff_A_cDe528kn5_0;
	wire w_dff_A_OA3KMFzw5_0;
	wire w_dff_A_ORsblvhe9_0;
	wire w_dff_A_QlqjVhUC7_0;
	wire w_dff_A_OcZ2RIcp8_0;
	wire w_dff_A_YWlqxvnI8_0;
	wire w_dff_A_tSju8ERv6_0;
	wire w_dff_A_l3p1HFJs9_0;
	wire w_dff_A_LCy2irS62_0;
	wire w_dff_A_S2HXu8WE8_0;
	wire w_dff_A_lGd6oMyr3_0;
	wire w_dff_A_nZMV21yo1_0;
	wire w_dff_A_2dDEbAuI8_0;
	wire w_dff_A_mvSkrnOo8_0;
	wire w_dff_A_JDqeIWOB3_0;
	wire w_dff_A_zLa4xw4d8_0;
	wire w_dff_A_NHTmnWzZ6_0;
	wire w_dff_A_kBywAWeH1_0;
	wire w_dff_A_s41c1RUy2_0;
	wire w_dff_A_Pow3qPc02_0;
	wire w_dff_A_YZtryBzI5_0;
	wire w_dff_A_ThqVqPIM1_0;
	wire w_dff_A_N18mvCOA7_0;
	wire w_dff_A_dCrDcmGc0_0;
	wire w_dff_A_NFr1gWhT7_0;
	wire w_dff_A_jSzvHIwD2_0;
	wire w_dff_A_bZEafMQb4_0;
	wire w_dff_A_CrFqYhE37_0;
	wire w_dff_A_uz0G5zVt6_0;
	wire w_dff_A_5YEyLRgp1_0;
	wire w_dff_A_une5EDtn3_0;
	wire w_dff_A_HHmjhqcT3_0;
	wire w_dff_A_ABjHjKIJ1_0;
	wire w_dff_A_L3Vo3gBg8_0;
	wire w_dff_A_AWlYYlg03_0;
	wire w_dff_A_JPX9N0WJ6_0;
	wire w_dff_A_19a4yM0v1_0;
	wire w_dff_A_eVPz5MYC9_0;
	wire w_dff_A_GGaeYQ9t8_0;
	wire w_dff_A_JgsCMeoa0_0;
	wire w_dff_A_kAXY9dL53_0;
	wire w_dff_A_2Ly2Dkto3_0;
	wire w_dff_A_flgrYN4N1_0;
	wire w_dff_A_DGVT5jvk5_0;
	wire w_dff_A_JIss0YJB5_2;
	wire w_dff_A_dFCI4bb25_0;
	wire w_dff_A_GFVnMEX32_0;
	wire w_dff_A_PdhYMYTa6_0;
	wire w_dff_A_uwY7OENu0_0;
	wire w_dff_A_DwBmud3r9_0;
	wire w_dff_A_QcemS1tT2_0;
	wire w_dff_A_dF2stYhj8_0;
	wire w_dff_A_QEWyKXxR0_0;
	wire w_dff_A_BP5s2Fs15_0;
	wire w_dff_A_sCdy9pmJ7_0;
	wire w_dff_A_BAY9jtZM7_0;
	wire w_dff_A_3DrsgkwA4_0;
	wire w_dff_A_O7FILHmv1_0;
	wire w_dff_A_dCCpwe6g4_0;
	wire w_dff_A_ccFSYTPt6_0;
	wire w_dff_A_z7sxxBzn0_0;
	wire w_dff_A_WiuD2U8K2_0;
	wire w_dff_A_NDPKldIP0_0;
	wire w_dff_A_uv4kS5KF2_0;
	wire w_dff_A_EInzX4nG2_0;
	wire w_dff_A_SXRDNqca6_0;
	wire w_dff_A_UeQg360x7_0;
	wire w_dff_A_nmm01ZeL2_0;
	wire w_dff_A_T7UI2LqQ6_0;
	wire w_dff_A_lFapPDyx4_0;
	wire w_dff_A_UKtNuHeG7_0;
	wire w_dff_A_mz5OpgzS5_0;
	wire w_dff_A_djjwCMzg8_0;
	wire w_dff_A_0jpo4vPB3_0;
	wire w_dff_A_V90F3OSd8_0;
	wire w_dff_A_renxw8Dy1_0;
	wire w_dff_A_yJ4zkDVc7_0;
	wire w_dff_A_vaM0UJ282_0;
	wire w_dff_A_O8PSyLRJ1_0;
	wire w_dff_A_Y7eQ8eLF1_0;
	wire w_dff_A_58NvqY4K1_0;
	wire w_dff_A_fa3M0Vwx4_0;
	wire w_dff_A_L4fIWzaq4_0;
	wire w_dff_A_4hDSqpYX9_0;
	wire w_dff_A_69heILq08_0;
	wire w_dff_A_lDrRWOtQ4_0;
	wire w_dff_A_iUBY8FeP4_0;
	wire w_dff_A_TIR4IRzl3_0;
	wire w_dff_A_JDijeVCl4_0;
	wire w_dff_A_vKPhDFbO0_0;
	wire w_dff_A_6ns2hWIN5_0;
	wire w_dff_A_Na6CQS4z7_0;
	wire w_dff_A_tXYMzNL66_0;
	wire w_dff_A_E54WVSOc3_0;
	wire w_dff_A_BSKt0ocr1_0;
	wire w_dff_A_dHs4lF3q7_0;
	wire w_dff_A_0fw8tlyi2_0;
	wire w_dff_A_Ilb9BIp96_0;
	wire w_dff_A_IAU5FW1b1_0;
	wire w_dff_A_idXBsFgP0_0;
	wire w_dff_A_EcQN55hq3_0;
	wire w_dff_A_LHHL1ujd8_0;
	wire w_dff_A_piItm0YG7_0;
	wire w_dff_A_uzv6tZZ44_0;
	wire w_dff_A_07i9yxNv3_0;
	wire w_dff_A_mX6H77rn3_0;
	wire w_dff_A_p7gXbnKb1_0;
	wire w_dff_A_b46PmH9S7_0;
	wire w_dff_A_DwpVE6mL5_0;
	wire w_dff_A_915szK9h8_0;
	wire w_dff_A_lQtbeT7y7_0;
	wire w_dff_A_MJ0uYOoe6_0;
	wire w_dff_A_FNQX1sKs5_0;
	wire w_dff_A_jnRz40jd9_0;
	wire w_dff_A_OnAJmf9o9_0;
	wire w_dff_A_knavpqI26_0;
	wire w_dff_A_kQK27dXJ2_0;
	wire w_dff_A_l7Fvddct6_0;
	wire w_dff_A_le0X9G589_0;
	wire w_dff_A_jphLi6kC3_0;
	wire w_dff_A_ZygH8nJ06_0;
	wire w_dff_A_SYgmEh182_0;
	wire w_dff_A_1jPWKSFF8_0;
	wire w_dff_A_O9VFiXuI4_0;
	wire w_dff_A_KvTgUuRd4_0;
	wire w_dff_A_TbFnflIP9_0;
	wire w_dff_A_shMaAjZz3_0;
	wire w_dff_A_yDHJuRpm3_0;
	wire w_dff_A_4V0cJoRk8_0;
	wire w_dff_A_UNa3qPhz6_0;
	wire w_dff_A_fv0KZ2QH1_0;
	wire w_dff_A_DBhMB6uc9_0;
	wire w_dff_A_tZewAjMR5_0;
	wire w_dff_A_DYovrw3X8_0;
	wire w_dff_A_Mek4U3ad6_0;
	wire w_dff_A_VQLu4bnW8_0;
	wire w_dff_A_b5cjhAkL5_0;
	wire w_dff_A_JArkOiN17_0;
	wire w_dff_A_7MLLdLaI6_0;
	wire w_dff_A_MNkbdDQn4_0;
	wire w_dff_A_wzovpAgm6_0;
	wire w_dff_A_U7lON1Fz3_0;
	wire w_dff_A_biKLaRG36_0;
	wire w_dff_A_8lnx8x7n9_0;
	wire w_dff_A_7BbhU6Rh4_2;
	wire w_dff_A_LfqjixaV1_0;
	wire w_dff_A_CzG9471b4_0;
	wire w_dff_A_r9azPEcN4_0;
	wire w_dff_A_Pdgj5oec8_0;
	wire w_dff_A_Q2gWDUY78_0;
	wire w_dff_A_ptNq7EdW8_0;
	wire w_dff_A_UdO4ShWI5_0;
	wire w_dff_A_ubKkkyBH8_0;
	wire w_dff_A_tP9rBEk95_0;
	wire w_dff_A_JUBlxMuu0_0;
	wire w_dff_A_rTagaEW07_0;
	wire w_dff_A_Gwi2Ek4F6_0;
	wire w_dff_A_mWuA76ee5_0;
	wire w_dff_A_hRvtBTWC3_0;
	wire w_dff_A_9NKhObai5_0;
	wire w_dff_A_ms7K6n391_0;
	wire w_dff_A_2pCs6kaU2_0;
	wire w_dff_A_VcXGayQJ3_0;
	wire w_dff_A_Xomayz0X0_0;
	wire w_dff_A_4zi2NolQ5_0;
	wire w_dff_A_EDA33RRY5_0;
	wire w_dff_A_EOLFbbpO6_0;
	wire w_dff_A_wRLglZug3_0;
	wire w_dff_A_mAvKB8PR2_0;
	wire w_dff_A_6siqoi348_0;
	wire w_dff_A_aXlJ4mY71_0;
	wire w_dff_A_pjUxnIH16_0;
	wire w_dff_A_GLfpGtGX4_0;
	wire w_dff_A_c4LuTLzM0_0;
	wire w_dff_A_BAqqw0lj6_0;
	wire w_dff_A_g8teRVBZ3_0;
	wire w_dff_A_vxhYtxqg9_0;
	wire w_dff_A_b8AYPQMS8_0;
	wire w_dff_A_SSDggxQG5_0;
	wire w_dff_A_WPudK0A88_0;
	wire w_dff_A_KCBKK5vs7_0;
	wire w_dff_A_7oTS1dvG8_0;
	wire w_dff_A_LJMblzin1_0;
	wire w_dff_A_YqGI9qVV9_0;
	wire w_dff_A_96B7wQuc6_0;
	wire w_dff_A_lxNJOSC74_0;
	wire w_dff_A_QVdlgMqI3_0;
	wire w_dff_A_X3plMJtd9_0;
	wire w_dff_A_Jk0J2XwE4_0;
	wire w_dff_A_OdOqU9Bt2_0;
	wire w_dff_A_rIEtuhjR9_0;
	wire w_dff_A_p3Obv0Sw7_0;
	wire w_dff_A_T2tSucid8_0;
	wire w_dff_A_RU3Ti26G0_0;
	wire w_dff_A_kHFJTMML4_0;
	wire w_dff_A_SHxhsyGG1_0;
	wire w_dff_A_g72auxyq1_0;
	wire w_dff_A_j3Hgo9yH8_0;
	wire w_dff_A_3iuzaVec6_0;
	wire w_dff_A_an3tkXxa8_0;
	wire w_dff_A_6PciCPRA1_0;
	wire w_dff_A_T998yKGk5_0;
	wire w_dff_A_iBNgGZqc7_0;
	wire w_dff_A_Wx6HAjrJ9_0;
	wire w_dff_A_AmtJ0Lvy4_0;
	wire w_dff_A_iLT03WhG6_0;
	wire w_dff_A_cCFA310V2_0;
	wire w_dff_A_3BkecCwr9_0;
	wire w_dff_A_TD3hJ0WH6_0;
	wire w_dff_A_La7zAyyV0_0;
	wire w_dff_A_WkkvUzwc0_0;
	wire w_dff_A_MgnvXWx85_0;
	wire w_dff_A_gahUMigD7_0;
	wire w_dff_A_xLjB74ZW7_0;
	wire w_dff_A_FOiBFNYk7_0;
	wire w_dff_A_fIS3s7qB9_0;
	wire w_dff_A_1BufGXZm1_0;
	wire w_dff_A_B1CbZCMp7_0;
	wire w_dff_A_scuF2Pnb9_0;
	wire w_dff_A_W4kKV87n5_0;
	wire w_dff_A_0qtbZQjT4_0;
	wire w_dff_A_0wX0dJp43_0;
	wire w_dff_A_N6EuIn5d5_0;
	wire w_dff_A_mBWVEsDc6_0;
	wire w_dff_A_wyw8CGco8_0;
	wire w_dff_A_XIoD1hcd4_0;
	wire w_dff_A_0L0o0DIo3_0;
	wire w_dff_A_7zhPa08u0_0;
	wire w_dff_A_GDXXn1gl2_0;
	wire w_dff_A_bYiZELNT2_0;
	wire w_dff_A_tJV84ufY1_0;
	wire w_dff_A_Nd6E7wDl2_0;
	wire w_dff_A_gUiLEGFE7_0;
	wire w_dff_A_W0ruTNHa6_0;
	wire w_dff_A_GbwNOgds9_0;
	wire w_dff_A_Yx9e2PyO5_0;
	wire w_dff_A_SW6Hhg3R3_0;
	wire w_dff_A_OMKRgBxR8_0;
	wire w_dff_A_QOgItMQH7_0;
	wire w_dff_A_cqMWJ4D96_0;
	wire w_dff_A_kNwMTneU3_0;
	wire w_dff_A_pQd90E2v8_0;
	wire w_dff_A_RaNHooAH3_0;
	wire w_dff_A_MfypuXxv4_2;
	wire w_dff_A_zdOlqrlj4_0;
	wire w_dff_A_42fAdlNi0_0;
	wire w_dff_A_p9M1fOqB7_0;
	wire w_dff_A_aundsJR19_0;
	wire w_dff_A_jlRrOq8l8_0;
	wire w_dff_A_57Jc3TMY4_0;
	wire w_dff_A_fBVi7L3t4_0;
	wire w_dff_A_TQQ8eY0j7_0;
	wire w_dff_A_cQ2JmozW7_0;
	wire w_dff_A_3jynR71t7_0;
	wire w_dff_A_QEwdM94c7_0;
	wire w_dff_A_a2MCaISr1_0;
	wire w_dff_A_malu6XMK8_0;
	wire w_dff_A_IEqFLfRv0_0;
	wire w_dff_A_RBHYtUxk6_0;
	wire w_dff_A_iRyGJHqH5_0;
	wire w_dff_A_ZZbYLUlh6_0;
	wire w_dff_A_QDjTkkt51_0;
	wire w_dff_A_I3djsEor7_0;
	wire w_dff_A_wFNrXV636_0;
	wire w_dff_A_QzkpQ2G45_0;
	wire w_dff_A_lXLczKgJ3_0;
	wire w_dff_A_j4EINsUi7_0;
	wire w_dff_A_h5xR87ZD9_0;
	wire w_dff_A_E7yf5PqQ5_0;
	wire w_dff_A_bpHb6z6x1_0;
	wire w_dff_A_9ijk4KA32_0;
	wire w_dff_A_i49vIbw44_0;
	wire w_dff_A_N45sGNyX9_0;
	wire w_dff_A_qX3iKmqT5_0;
	wire w_dff_A_0mLib3Ic1_0;
	wire w_dff_A_3zze6v4u0_0;
	wire w_dff_A_0noVYfVc3_0;
	wire w_dff_A_JsOfsVKn6_0;
	wire w_dff_A_keJyqdro0_0;
	wire w_dff_A_Rl8vP1is3_0;
	wire w_dff_A_KR1HlduH4_0;
	wire w_dff_A_yt6d0OFb4_0;
	wire w_dff_A_JCZDrZux9_0;
	wire w_dff_A_qk3nEWK17_0;
	wire w_dff_A_Z9KNJgDX7_0;
	wire w_dff_A_drbAPcoA8_0;
	wire w_dff_A_Qh0Fs5Pk3_0;
	wire w_dff_A_XeMNdYYl4_0;
	wire w_dff_A_7kClTru31_0;
	wire w_dff_A_3DXMF5qy5_0;
	wire w_dff_A_aV71sszD9_0;
	wire w_dff_A_LzAA1TkY3_0;
	wire w_dff_A_Fdw45Z5A7_0;
	wire w_dff_A_cn5LbfD82_0;
	wire w_dff_A_s8eDJzvw0_0;
	wire w_dff_A_fF8YfCvq9_0;
	wire w_dff_A_mVi9qIpC7_0;
	wire w_dff_A_UOAuhCY19_0;
	wire w_dff_A_ixGzX1ZG5_0;
	wire w_dff_A_xjvzFRTM7_0;
	wire w_dff_A_3TgUbAwo5_0;
	wire w_dff_A_IOBOnBpN0_0;
	wire w_dff_A_aZHK1LBo3_0;
	wire w_dff_A_UlPb7xGx1_0;
	wire w_dff_A_3iSZb6iK8_0;
	wire w_dff_A_wIa54FeD1_0;
	wire w_dff_A_NcGd930p7_0;
	wire w_dff_A_Kf3VFY2b2_0;
	wire w_dff_A_N3bVx1ge8_0;
	wire w_dff_A_B8Vtbp0b0_0;
	wire w_dff_A_duyq20ZB4_0;
	wire w_dff_A_Kl1xbcvj7_0;
	wire w_dff_A_ZpfVUx930_0;
	wire w_dff_A_p8UVQvug3_0;
	wire w_dff_A_C4bcxwWo5_0;
	wire w_dff_A_XulejHAB3_0;
	wire w_dff_A_VsEKWqlu7_0;
	wire w_dff_A_eVRwYDbN9_0;
	wire w_dff_A_mWXkjwms5_0;
	wire w_dff_A_v5ozceBS8_0;
	wire w_dff_A_0f6rSJEj0_0;
	wire w_dff_A_g9mNr2lb5_0;
	wire w_dff_A_amNppAe01_0;
	wire w_dff_A_fHmNsu873_0;
	wire w_dff_A_u8klzVdW5_0;
	wire w_dff_A_MXTUzSFv4_0;
	wire w_dff_A_RWccJ74E2_0;
	wire w_dff_A_lEp38xPX1_0;
	wire w_dff_A_UgxBCfoA6_0;
	wire w_dff_A_EGnWsPIg8_0;
	wire w_dff_A_iQZxSYWs6_0;
	wire w_dff_A_y9gAim2U1_0;
	wire w_dff_A_St7HXQh97_0;
	wire w_dff_A_RXPWyulM1_0;
	wire w_dff_A_9vfmBxph2_0;
	wire w_dff_A_lX9CmjXJ9_0;
	wire w_dff_A_rWTbbxb21_0;
	wire w_dff_A_a3s3Pj7Q9_0;
	wire w_dff_A_Q5uI4hct1_0;
	wire w_dff_A_Qwv4GP0i3_0;
	wire w_dff_A_P9WI9vn16_0;
	wire w_dff_A_m45eyEAd4_2;
	wire w_dff_A_Wx2kalZ99_0;
	wire w_dff_A_EvLJEHTp5_0;
	wire w_dff_A_XlS8aBvx3_0;
	wire w_dff_A_v0r4CZtO2_0;
	wire w_dff_A_Penvwuy62_0;
	wire w_dff_A_RT75uAev7_0;
	wire w_dff_A_1P7i1joJ7_0;
	wire w_dff_A_PoWmjduH7_0;
	wire w_dff_A_QoIRXqco0_0;
	wire w_dff_A_ziKmwNuf6_0;
	wire w_dff_A_Iito4yRU6_0;
	wire w_dff_A_vJsyDuPA2_0;
	wire w_dff_A_CpnoYG6B6_0;
	wire w_dff_A_1jpseo286_0;
	wire w_dff_A_nLWBu4Cq4_0;
	wire w_dff_A_bAqmkQ7I7_0;
	wire w_dff_A_uluriX6K5_0;
	wire w_dff_A_RstTxIl16_0;
	wire w_dff_A_9f3Ev0xc5_0;
	wire w_dff_A_MNhZlhs06_0;
	wire w_dff_A_5FB3KJOx8_0;
	wire w_dff_A_JVTUOxxr4_0;
	wire w_dff_A_V1OTSyzX4_0;
	wire w_dff_A_4OoHZF5N3_0;
	wire w_dff_A_vXNH0Y9J2_0;
	wire w_dff_A_hvv1rbL06_0;
	wire w_dff_A_dvYP2lsa1_0;
	wire w_dff_A_ARgXA8Kr9_0;
	wire w_dff_A_Us18klBO3_0;
	wire w_dff_A_Bz56m29g8_0;
	wire w_dff_A_buRIKoaZ1_0;
	wire w_dff_A_VAWnMiBM9_0;
	wire w_dff_A_cv5Zs6vR2_0;
	wire w_dff_A_757iSOvs6_0;
	wire w_dff_A_vs1lzyKN0_0;
	wire w_dff_A_snFj8Xpl5_0;
	wire w_dff_A_rtq30XW18_0;
	wire w_dff_A_x0DbNDtM6_0;
	wire w_dff_A_346KtL4V2_0;
	wire w_dff_A_xWrAODEW4_0;
	wire w_dff_A_NsReiRRY4_0;
	wire w_dff_A_HnZohz3y1_0;
	wire w_dff_A_BT3erJOD0_0;
	wire w_dff_A_TboxvwgO8_0;
	wire w_dff_A_NO6JhiHs4_0;
	wire w_dff_A_sdL7SRKG8_0;
	wire w_dff_A_AHAq9gor6_0;
	wire w_dff_A_iBGnvnJm3_0;
	wire w_dff_A_SPMYRRwN1_0;
	wire w_dff_A_UET1ivrO7_0;
	wire w_dff_A_oBLNfSXw3_0;
	wire w_dff_A_wHq79Frn5_0;
	wire w_dff_A_ADugQLl23_0;
	wire w_dff_A_SmTcV4mc6_0;
	wire w_dff_A_IXIcvFv44_0;
	wire w_dff_A_o8PPN4bL5_0;
	wire w_dff_A_heM0Ijud4_0;
	wire w_dff_A_wO4uCGDJ5_0;
	wire w_dff_A_1MrudNvZ3_0;
	wire w_dff_A_t7LQzEWn2_0;
	wire w_dff_A_ILTVRGTn0_0;
	wire w_dff_A_JNX0A4MM6_0;
	wire w_dff_A_PAEzTRqn5_0;
	wire w_dff_A_ybZFxMBl2_0;
	wire w_dff_A_jrz5Vp8X8_0;
	wire w_dff_A_9BSXmlwp0_0;
	wire w_dff_A_b3eRhrYR7_0;
	wire w_dff_A_A2gXLhvE6_0;
	wire w_dff_A_9ko22dCP5_0;
	wire w_dff_A_Mc04vk5y2_0;
	wire w_dff_A_D4EhNa4Z4_0;
	wire w_dff_A_I8X08HfC5_0;
	wire w_dff_A_CUzDiWlv2_0;
	wire w_dff_A_mP6rND1o0_0;
	wire w_dff_A_0EGG93Ll7_0;
	wire w_dff_A_tg31B4vn7_0;
	wire w_dff_A_ADCqHYX24_0;
	wire w_dff_A_hUd96aIE0_0;
	wire w_dff_A_d6y7TEOy1_0;
	wire w_dff_A_PIVki6Pr5_0;
	wire w_dff_A_sSpUrxNE5_0;
	wire w_dff_A_sqMkZJiv2_0;
	wire w_dff_A_BJ6vWbrU0_0;
	wire w_dff_A_LogdoRNP9_0;
	wire w_dff_A_LFxHf0T66_0;
	wire w_dff_A_8im5i1fx1_0;
	wire w_dff_A_wb0OGDCr6_0;
	wire w_dff_A_a9tlW0gb4_0;
	wire w_dff_A_gXPX3UOS7_0;
	wire w_dff_A_qjwJ2l7P5_0;
	wire w_dff_A_KQr5rPeX5_0;
	wire w_dff_A_q30YGg2D0_0;
	wire w_dff_A_ypL7O0d37_0;
	wire w_dff_A_PvH6dXMl1_0;
	wire w_dff_A_L37lSGjN8_0;
	wire w_dff_A_2iosBtlP0_0;
	wire w_dff_A_HDJk7IDG5_2;
	wire w_dff_A_1KMSk5ni1_0;
	wire w_dff_A_LBQ3UZQS9_0;
	wire w_dff_A_iIf5jTlO5_0;
	wire w_dff_A_tkt2TCsn4_0;
	wire w_dff_A_QQpFWzS42_0;
	wire w_dff_A_PSWnTCZk3_0;
	wire w_dff_A_F4svAYcv1_0;
	wire w_dff_A_Xv5YH3f47_0;
	wire w_dff_A_v5s7pVLT7_0;
	wire w_dff_A_ZL25zWmZ5_0;
	wire w_dff_A_52hs2BNB6_0;
	wire w_dff_A_Va2DCOu51_0;
	wire w_dff_A_6LX25aEP9_0;
	wire w_dff_A_hRtGsuXF9_0;
	wire w_dff_A_RWPh9Knb3_0;
	wire w_dff_A_zyqUGTLi3_0;
	wire w_dff_A_Jgwcf05p3_0;
	wire w_dff_A_hwqlJh622_0;
	wire w_dff_A_jdzatfsk0_0;
	wire w_dff_A_A9VfYmQc4_0;
	wire w_dff_A_8LbLg9rS0_0;
	wire w_dff_A_Oz9q12bm0_0;
	wire w_dff_A_C8PnyTQS7_0;
	wire w_dff_A_Ku3Iad2r5_0;
	wire w_dff_A_DqvvcaWd6_0;
	wire w_dff_A_LN1mXno33_0;
	wire w_dff_A_xdNAfvfx0_0;
	wire w_dff_A_VLLhdAlN0_0;
	wire w_dff_A_8tA0gMe51_0;
	wire w_dff_A_XKr94d6V6_0;
	wire w_dff_A_yQpU0N8V2_0;
	wire w_dff_A_I2tGDJvr7_0;
	wire w_dff_A_4CUjPcWF2_0;
	wire w_dff_A_7vczdNd62_0;
	wire w_dff_A_Tfn1NlVW9_0;
	wire w_dff_A_IcjXBsl08_0;
	wire w_dff_A_sf6HM8qM6_0;
	wire w_dff_A_ANAj00bb7_0;
	wire w_dff_A_Vu4xvi6C5_0;
	wire w_dff_A_P3IcNp4f3_0;
	wire w_dff_A_RooPtbgS0_0;
	wire w_dff_A_H6FfmfWI9_0;
	wire w_dff_A_1yy10Jbe9_0;
	wire w_dff_A_lsjMGliR7_0;
	wire w_dff_A_rgfsf5Yy5_0;
	wire w_dff_A_jr8yS74M4_0;
	wire w_dff_A_HVcr2GXv0_0;
	wire w_dff_A_tdYKs75q0_0;
	wire w_dff_A_QVztt8No4_0;
	wire w_dff_A_9fYhtoq06_0;
	wire w_dff_A_x0KInFsh7_0;
	wire w_dff_A_BCufJ05V9_0;
	wire w_dff_A_bdueen1P7_0;
	wire w_dff_A_tUX7ATe30_0;
	wire w_dff_A_C9jqr3F16_0;
	wire w_dff_A_Lft4Y8zd6_0;
	wire w_dff_A_h6lxUglG7_0;
	wire w_dff_A_DOeJSmlX8_0;
	wire w_dff_A_DaUJHaia9_0;
	wire w_dff_A_1pd9r7Lz1_0;
	wire w_dff_A_Zt2DUzCI9_0;
	wire w_dff_A_yAguPVvr3_0;
	wire w_dff_A_HD5dY2QX6_0;
	wire w_dff_A_C8Vla8lD6_0;
	wire w_dff_A_aTsiJJrv4_0;
	wire w_dff_A_9mqD6HUG9_0;
	wire w_dff_A_Iw5anqG08_0;
	wire w_dff_A_X4pmaQtB5_0;
	wire w_dff_A_IPFAysBJ2_0;
	wire w_dff_A_KmQYMo2f8_0;
	wire w_dff_A_kSpLcaRg0_0;
	wire w_dff_A_gwo3cl2g1_0;
	wire w_dff_A_RNmscOtN0_0;
	wire w_dff_A_e21daD3A5_0;
	wire w_dff_A_FL5nlnuk2_0;
	wire w_dff_A_mF38GD9n2_0;
	wire w_dff_A_MCCRLRZ42_0;
	wire w_dff_A_Q6wfGJAf8_0;
	wire w_dff_A_SDIwXHON3_0;
	wire w_dff_A_xzUct8pV1_0;
	wire w_dff_A_ZVXFcrWg6_0;
	wire w_dff_A_NjyRr0XE5_0;
	wire w_dff_A_qi0spAow0_0;
	wire w_dff_A_IKJdRuNe5_0;
	wire w_dff_A_tyFnN7DZ0_0;
	wire w_dff_A_qmyFeJwd2_0;
	wire w_dff_A_pqhGVZIS8_0;
	wire w_dff_A_040MvXAb1_0;
	wire w_dff_A_DIwhYRBt6_0;
	wire w_dff_A_LtSWvQew5_0;
	wire w_dff_A_4zHkLZ1s7_0;
	wire w_dff_A_urxoGnKd6_0;
	wire w_dff_A_f51uoYlA1_0;
	wire w_dff_A_gf7ecoOt2_0;
	wire w_dff_A_hY9hUxCJ7_0;
	wire w_dff_A_Vbwd5rP60_2;
	wire w_dff_A_acguHRy91_0;
	wire w_dff_A_eWBgmLM32_0;
	wire w_dff_A_JSH2BpPH9_0;
	wire w_dff_A_HMEXUphm2_0;
	wire w_dff_A_bcVfDLXc9_0;
	wire w_dff_A_5WXv0ir40_0;
	wire w_dff_A_qFOHSeqv5_0;
	wire w_dff_A_ghqATLCH7_0;
	wire w_dff_A_jtc57SmF2_0;
	wire w_dff_A_TxwVwgWQ2_0;
	wire w_dff_A_YJb9zqtS3_0;
	wire w_dff_A_clURgq829_0;
	wire w_dff_A_B9nmkbPJ4_0;
	wire w_dff_A_2k5Gk8BW7_0;
	wire w_dff_A_xhVLUZNi0_0;
	wire w_dff_A_Eq0bb39p0_0;
	wire w_dff_A_lZWxKl9K6_0;
	wire w_dff_A_Bkm471TL8_0;
	wire w_dff_A_mbXB2Dlq7_0;
	wire w_dff_A_8cDSucz92_0;
	wire w_dff_A_zH2D31n48_0;
	wire w_dff_A_IllvKo8r0_0;
	wire w_dff_A_F20VDSIx8_0;
	wire w_dff_A_Gy8blDOL3_0;
	wire w_dff_A_R4YmRgQh0_0;
	wire w_dff_A_ZdZ8LIVF8_0;
	wire w_dff_A_lYwOT3XD6_0;
	wire w_dff_A_8NbSjTYQ0_0;
	wire w_dff_A_8zrlZBVF5_0;
	wire w_dff_A_f4lrLZTC3_0;
	wire w_dff_A_gDeO2G2C8_0;
	wire w_dff_A_FYGNwlxr1_0;
	wire w_dff_A_pfDFAsdz6_0;
	wire w_dff_A_zhWHKqVw6_0;
	wire w_dff_A_nxdqapsb6_0;
	wire w_dff_A_9Ifi4L7F7_0;
	wire w_dff_A_e6CBJ4h21_0;
	wire w_dff_A_PyiqqjOK3_0;
	wire w_dff_A_0aj8yugc3_0;
	wire w_dff_A_Kbk3X0P69_0;
	wire w_dff_A_ZFyWwRUf5_0;
	wire w_dff_A_LjKvTvfa8_0;
	wire w_dff_A_pKhsl2lB8_0;
	wire w_dff_A_mg62jM3S4_0;
	wire w_dff_A_AAqXqg4v1_0;
	wire w_dff_A_7y4CXdXA3_0;
	wire w_dff_A_VeG9PlFa4_0;
	wire w_dff_A_VHCXykxR6_0;
	wire w_dff_A_r2eJsA1e5_0;
	wire w_dff_A_lyLOCxks8_0;
	wire w_dff_A_NKwRdkeW2_0;
	wire w_dff_A_pb51qD7V7_0;
	wire w_dff_A_Dh9H56nq3_0;
	wire w_dff_A_e3fK55SL2_0;
	wire w_dff_A_aSqW5MCq7_0;
	wire w_dff_A_FIlD0ynx6_0;
	wire w_dff_A_1jOcEIC86_0;
	wire w_dff_A_ErHwsI9U1_0;
	wire w_dff_A_E0UGvoOz7_0;
	wire w_dff_A_b4I4O6NT4_0;
	wire w_dff_A_Qvjglidr8_0;
	wire w_dff_A_7hICxZOP3_0;
	wire w_dff_A_b3ZCy4If2_0;
	wire w_dff_A_iNXygzty4_0;
	wire w_dff_A_I6CWKPnt2_0;
	wire w_dff_A_Ij6AZunJ7_0;
	wire w_dff_A_J8aEbPPM5_0;
	wire w_dff_A_8LEMS8j92_0;
	wire w_dff_A_zuTy6rDg4_0;
	wire w_dff_A_lMoM9Gie5_0;
	wire w_dff_A_63TjIIhN6_0;
	wire w_dff_A_9U3JIBlW5_0;
	wire w_dff_A_dOXYVYLk3_0;
	wire w_dff_A_iQkxLnZO6_0;
	wire w_dff_A_e9uXjCFR8_0;
	wire w_dff_A_D1x8SWGG8_0;
	wire w_dff_A_EN0b0VM04_0;
	wire w_dff_A_hOUe51KZ0_0;
	wire w_dff_A_RASIn91O7_0;
	wire w_dff_A_C5xiiUX07_0;
	wire w_dff_A_5ocXhG7j9_0;
	wire w_dff_A_lrIdjV6O5_0;
	wire w_dff_A_v27JInPy5_0;
	wire w_dff_A_JwrjPW391_0;
	wire w_dff_A_b3eubL1g9_0;
	wire w_dff_A_SVuujN5B0_0;
	wire w_dff_A_clOeg2UJ0_0;
	wire w_dff_A_IQkFWOGN0_0;
	wire w_dff_A_VZcJ0Hsj1_0;
	wire w_dff_A_371ihWaD5_0;
	wire w_dff_A_l6xAvpDk0_0;
	wire w_dff_A_YGN7U03v6_0;
	wire w_dff_A_PR52G4kM5_0;
	wire w_dff_A_xGcvzYlW6_0;
	wire w_dff_A_AA7idxgZ2_2;
	wire w_dff_A_IXmzJoD52_0;
	wire w_dff_A_SUiDWMsI0_0;
	wire w_dff_A_8ttcsU1w2_0;
	wire w_dff_A_BtjTE1X13_0;
	wire w_dff_A_iIJyQgKl8_0;
	wire w_dff_A_4BgOiuQ80_0;
	wire w_dff_A_ar2v2KAu2_0;
	wire w_dff_A_OI9oBg3b5_0;
	wire w_dff_A_Fvd5Iqva9_0;
	wire w_dff_A_e4DhpLi45_0;
	wire w_dff_A_AdpjdJE36_0;
	wire w_dff_A_uAxjzFmT5_0;
	wire w_dff_A_oiCFDegG8_0;
	wire w_dff_A_LZFLbM197_0;
	wire w_dff_A_DDdq2hdP1_0;
	wire w_dff_A_4swA2f0R9_0;
	wire w_dff_A_pD2JoyfP9_0;
	wire w_dff_A_JkLgDBAh7_0;
	wire w_dff_A_6atLCMun9_0;
	wire w_dff_A_FzUfkCb47_0;
	wire w_dff_A_s28azhb96_0;
	wire w_dff_A_BKabnSNy7_0;
	wire w_dff_A_abzSJv9j8_0;
	wire w_dff_A_moYeier78_0;
	wire w_dff_A_3rJjjKxc2_0;
	wire w_dff_A_nXxWogiK6_0;
	wire w_dff_A_pYxWmkhq9_0;
	wire w_dff_A_9I0NvBXT3_0;
	wire w_dff_A_BSRWfDZO2_0;
	wire w_dff_A_Rqpj8eeM9_0;
	wire w_dff_A_D1MWBfai8_0;
	wire w_dff_A_ylUcUOKr0_0;
	wire w_dff_A_7HtJzcqB7_0;
	wire w_dff_A_RGHXKlFs4_0;
	wire w_dff_A_h7P5aI7x7_0;
	wire w_dff_A_smmsHfTa6_0;
	wire w_dff_A_EyUiVyjx5_0;
	wire w_dff_A_e4bPu2DX3_0;
	wire w_dff_A_3sr77xXo2_0;
	wire w_dff_A_DDofauw05_0;
	wire w_dff_A_uB5FBS4F3_0;
	wire w_dff_A_IiNkcaVJ4_0;
	wire w_dff_A_BjqJnB1N6_0;
	wire w_dff_A_RHqTVs6M4_0;
	wire w_dff_A_ziibFKak8_0;
	wire w_dff_A_obMBmyXc1_0;
	wire w_dff_A_WxsrymzD2_0;
	wire w_dff_A_H1viYh4t5_0;
	wire w_dff_A_OfYT7qSR0_0;
	wire w_dff_A_0DiFCaFh0_0;
	wire w_dff_A_f98SiEhU9_0;
	wire w_dff_A_iomll8mg2_0;
	wire w_dff_A_pd95cPaR6_0;
	wire w_dff_A_NAWgwRXy1_0;
	wire w_dff_A_zS2cQVBn4_0;
	wire w_dff_A_8LnUQHd07_0;
	wire w_dff_A_J6dmwfBt1_0;
	wire w_dff_A_f5mH1I341_0;
	wire w_dff_A_SnITCqxm0_0;
	wire w_dff_A_1wiy9psF6_0;
	wire w_dff_A_b7nmvzCl5_0;
	wire w_dff_A_B24VU6qr8_0;
	wire w_dff_A_BKMY13M98_0;
	wire w_dff_A_bGXrTSQm1_0;
	wire w_dff_A_0gfJ2qsd5_0;
	wire w_dff_A_qwMrHx5C7_0;
	wire w_dff_A_X7FPCX4q5_0;
	wire w_dff_A_o07PCTzF8_0;
	wire w_dff_A_Yk0FZKU76_0;
	wire w_dff_A_FlwsofEx2_0;
	wire w_dff_A_OnR1Doqj1_0;
	wire w_dff_A_2he1DkqY1_0;
	wire w_dff_A_F0QLvxFp8_0;
	wire w_dff_A_doVAtjvv4_0;
	wire w_dff_A_YNwZFz0b5_0;
	wire w_dff_A_iiS1uhtG2_0;
	wire w_dff_A_mSnl7QXm0_0;
	wire w_dff_A_qtMP3eTI2_0;
	wire w_dff_A_8gSwC1OM6_0;
	wire w_dff_A_4vJTNDWE6_0;
	wire w_dff_A_BXTRr1C68_0;
	wire w_dff_A_byH2M9Em8_0;
	wire w_dff_A_DCC8dUoA2_0;
	wire w_dff_A_mW4mUuKi0_0;
	wire w_dff_A_RG18yxmP6_0;
	wire w_dff_A_YrIiJjdx1_0;
	wire w_dff_A_7RQJdfYD5_0;
	wire w_dff_A_rELg6bc66_0;
	wire w_dff_A_GRm0XSQP3_0;
	wire w_dff_A_ecCi7hRr4_0;
	wire w_dff_A_LXFfsDD52_0;
	wire w_dff_A_VcVhUY0c1_0;
	wire w_dff_A_rOMkywIm4_0;
	wire w_dff_A_RzzGmYzn3_2;
	wire w_dff_A_dBfSA6ub2_0;
	wire w_dff_A_XVUpZ1zt4_0;
	wire w_dff_A_ujn4DM6Y2_0;
	wire w_dff_A_l1mlQqA58_0;
	wire w_dff_A_muVwVuO97_0;
	wire w_dff_A_3CqjXeza9_0;
	wire w_dff_A_qSonBavG7_0;
	wire w_dff_A_jMbSoduW0_0;
	wire w_dff_A_TqndA2fP0_0;
	wire w_dff_A_5wxTBUxl4_0;
	wire w_dff_A_S6H1fwlD7_0;
	wire w_dff_A_K6qO0xqR0_0;
	wire w_dff_A_im83zL383_0;
	wire w_dff_A_9DOqdkgc0_0;
	wire w_dff_A_WJCw94Aj0_0;
	wire w_dff_A_KWN1dpvq2_0;
	wire w_dff_A_kxCmcfCc4_0;
	wire w_dff_A_lHHp85zP6_0;
	wire w_dff_A_BYrGi2QE3_0;
	wire w_dff_A_zk1BHnw74_0;
	wire w_dff_A_64r3MPyM1_0;
	wire w_dff_A_m3JAd3kv5_0;
	wire w_dff_A_0coZ5S9K5_0;
	wire w_dff_A_QB0Ew6V78_0;
	wire w_dff_A_5iNSLTx45_0;
	wire w_dff_A_bYHfNVbu0_0;
	wire w_dff_A_iJkKEHDC9_0;
	wire w_dff_A_pCb7MVQY4_0;
	wire w_dff_A_0A1tRegP0_0;
	wire w_dff_A_7IqpVO0B0_0;
	wire w_dff_A_AW8ITODf7_0;
	wire w_dff_A_fqASo0au1_0;
	wire w_dff_A_me17I2Uh7_0;
	wire w_dff_A_SHmfCT5H6_0;
	wire w_dff_A_XnnE3lZb4_0;
	wire w_dff_A_CAYP4COO3_0;
	wire w_dff_A_vT7dtpOs6_0;
	wire w_dff_A_0CCWzmD37_0;
	wire w_dff_A_rtpnFsbC4_0;
	wire w_dff_A_CNta6gfV7_0;
	wire w_dff_A_h1jEWET94_0;
	wire w_dff_A_PRPja86B6_0;
	wire w_dff_A_XmzsLt3A5_0;
	wire w_dff_A_4s28Zs3r3_0;
	wire w_dff_A_6DZhO1yC4_0;
	wire w_dff_A_J8SHmDK24_0;
	wire w_dff_A_Kfi0iQGv1_0;
	wire w_dff_A_lRlRaB3M2_0;
	wire w_dff_A_Duc2nt1T2_0;
	wire w_dff_A_tQeUDxrn0_0;
	wire w_dff_A_uXAl6YYf0_0;
	wire w_dff_A_F9UTqTjf7_0;
	wire w_dff_A_ktsnwwmm6_0;
	wire w_dff_A_yTS93qct5_0;
	wire w_dff_A_EkQB7zjQ9_0;
	wire w_dff_A_tQ0JowUq0_0;
	wire w_dff_A_PVT7U1Ql3_0;
	wire w_dff_A_sSql4X0H4_0;
	wire w_dff_A_Umyqc3P18_0;
	wire w_dff_A_cbI1DzSd1_0;
	wire w_dff_A_caKcpMok2_0;
	wire w_dff_A_LUG9mbHN3_0;
	wire w_dff_A_TxDL49bF2_0;
	wire w_dff_A_ArgMUspD6_0;
	wire w_dff_A_d8aAiL6X2_0;
	wire w_dff_A_PSF79s9m0_0;
	wire w_dff_A_jPrwRqPh1_0;
	wire w_dff_A_yJ53mRLy5_0;
	wire w_dff_A_14G7cpxf1_0;
	wire w_dff_A_SD4vpAb10_0;
	wire w_dff_A_PfqZXFCM0_0;
	wire w_dff_A_aIEP0Nlq5_0;
	wire w_dff_A_Jyw4jyqW7_0;
	wire w_dff_A_SCuselYG2_0;
	wire w_dff_A_7Z92uT2d2_0;
	wire w_dff_A_2j4uVMqg2_0;
	wire w_dff_A_0fuoSUpE0_0;
	wire w_dff_A_PLux0Fem7_0;
	wire w_dff_A_sZAgWQbQ5_0;
	wire w_dff_A_ST7RWL082_0;
	wire w_dff_A_miTjf7vK9_0;
	wire w_dff_A_QJTWqxwc1_0;
	wire w_dff_A_yI6rIQoi0_0;
	wire w_dff_A_naKFjRhr9_0;
	wire w_dff_A_g43cBc1v4_0;
	wire w_dff_A_hpfzuxVx6_0;
	wire w_dff_A_JDOqkfEf8_0;
	wire w_dff_A_gU9MVpxj7_0;
	wire w_dff_A_egeb3Qdl9_0;
	wire w_dff_A_BiyTWZcm5_0;
	wire w_dff_A_X1eUhFJm8_0;
	wire w_dff_A_Ilp4LSRo3_0;
	wire w_dff_A_tKTU1hRn7_2;
	wire w_dff_A_Ch2Oc2vb5_0;
	wire w_dff_A_nEGB37bK5_0;
	wire w_dff_A_ZiGXwpii3_0;
	wire w_dff_A_Q8VRtOFn1_0;
	wire w_dff_A_VHdbFjJo8_0;
	wire w_dff_A_hObWfp1Q2_0;
	wire w_dff_A_tpi6swYx9_0;
	wire w_dff_A_wlGiXxif3_0;
	wire w_dff_A_ujbI0SNB8_0;
	wire w_dff_A_DliQZfyC6_0;
	wire w_dff_A_fOcyHfS14_0;
	wire w_dff_A_NFEmeulP6_0;
	wire w_dff_A_RO69BTiY7_0;
	wire w_dff_A_URj2PuUt2_0;
	wire w_dff_A_7Jdxw4nk7_0;
	wire w_dff_A_TzpHA0bX3_0;
	wire w_dff_A_bzazDJTk5_0;
	wire w_dff_A_eE9Ur35R2_0;
	wire w_dff_A_LJpxmHmg6_0;
	wire w_dff_A_aS182kDO4_0;
	wire w_dff_A_0iGgeNPM6_0;
	wire w_dff_A_btKxdY4I0_0;
	wire w_dff_A_0z5DsSvY5_0;
	wire w_dff_A_TIZn6i9V6_0;
	wire w_dff_A_bIGOQxb50_0;
	wire w_dff_A_rsTvC55X9_0;
	wire w_dff_A_fAX1yO723_0;
	wire w_dff_A_AWg4IurG0_0;
	wire w_dff_A_vZOxgZKa5_0;
	wire w_dff_A_SHEgAk5h7_0;
	wire w_dff_A_sf0PebLT0_0;
	wire w_dff_A_kQl7OQ3c1_0;
	wire w_dff_A_ADZ85spc2_0;
	wire w_dff_A_LorQSN5d3_0;
	wire w_dff_A_rEbafI8f1_0;
	wire w_dff_A_JpdLi8XN8_0;
	wire w_dff_A_EH7Uq0tc1_0;
	wire w_dff_A_hYcRuqmh7_0;
	wire w_dff_A_GrHDx2OA1_0;
	wire w_dff_A_Ua3RxwqY9_0;
	wire w_dff_A_5nrNoENL2_0;
	wire w_dff_A_u4BwEYyt4_0;
	wire w_dff_A_rr7t9NPn8_0;
	wire w_dff_A_M0ZSeS8F3_0;
	wire w_dff_A_hNN00mLk6_0;
	wire w_dff_A_LFaK89Zb7_0;
	wire w_dff_A_TPKgoR8J2_0;
	wire w_dff_A_g8p3WKfb4_0;
	wire w_dff_A_cuh9UZAW3_0;
	wire w_dff_A_EJB30njP4_0;
	wire w_dff_A_Bf6PewtZ0_0;
	wire w_dff_A_kF9UhB5E9_0;
	wire w_dff_A_tAcKHAuS4_0;
	wire w_dff_A_vioj2Pha6_0;
	wire w_dff_A_CStbZH4x4_0;
	wire w_dff_A_3rH5S1gQ1_0;
	wire w_dff_A_a63eicb86_0;
	wire w_dff_A_6fDPp9Ko2_0;
	wire w_dff_A_xXjgOvOx6_0;
	wire w_dff_A_qsEblaWp6_0;
	wire w_dff_A_VE8F3smc3_0;
	wire w_dff_A_7dyisAIS6_0;
	wire w_dff_A_BlMmpKU17_0;
	wire w_dff_A_UmSf4Fxd1_0;
	wire w_dff_A_m9VmeOCU6_0;
	wire w_dff_A_JDSlJP507_0;
	wire w_dff_A_kwUMshQW9_0;
	wire w_dff_A_H1DIgAo81_0;
	wire w_dff_A_cDG6dHMF3_0;
	wire w_dff_A_wTl97SuH3_0;
	wire w_dff_A_fOBCRBWX0_0;
	wire w_dff_A_UW2g8f6K7_0;
	wire w_dff_A_Jzq2nXK18_0;
	wire w_dff_A_qML8P6q92_0;
	wire w_dff_A_rNbqGuBL8_0;
	wire w_dff_A_IJbS29KA6_0;
	wire w_dff_A_VpMBkWWc6_0;
	wire w_dff_A_VXEiqVYQ0_0;
	wire w_dff_A_J3s55izY0_0;
	wire w_dff_A_lBsBNlMg3_0;
	wire w_dff_A_KGShAaPC6_0;
	wire w_dff_A_iYupWikI9_0;
	wire w_dff_A_Ky1TfkKH7_0;
	wire w_dff_A_yg6YV2HR6_0;
	wire w_dff_A_daVDB4VH8_0;
	wire w_dff_A_tW5EWCgl4_0;
	wire w_dff_A_0Yg2Inx50_0;
	wire w_dff_A_araptS9w7_0;
	wire w_dff_A_qtWGmOkL9_0;
	wire w_dff_A_MsxhfmAU1_0;
	wire w_dff_A_WB1oNc4C1_0;
	wire w_dff_A_F7Oq80ij2_2;
	wire w_dff_A_bvG6h68p8_0;
	wire w_dff_A_kKbT802A6_0;
	wire w_dff_A_TicpFAni1_0;
	wire w_dff_A_e1ZMROkg9_0;
	wire w_dff_A_xtQuLvzQ0_0;
	wire w_dff_A_FyNeBQTy3_0;
	wire w_dff_A_ajSyLEgZ9_0;
	wire w_dff_A_UuGRcLn26_0;
	wire w_dff_A_0GLxM1s98_0;
	wire w_dff_A_uyO9Rpkf1_0;
	wire w_dff_A_EeGEq80i9_0;
	wire w_dff_A_5Pbfy8tK5_0;
	wire w_dff_A_GlZW5Kgo0_0;
	wire w_dff_A_wrqmMmbC5_0;
	wire w_dff_A_L6InOzRZ7_0;
	wire w_dff_A_h48qxO9F9_0;
	wire w_dff_A_SEgcmIzs9_0;
	wire w_dff_A_PVqVZHZZ2_0;
	wire w_dff_A_Dt7Yzrww5_0;
	wire w_dff_A_0fVxvMb70_0;
	wire w_dff_A_pMf4uDEF6_0;
	wire w_dff_A_knFVBxyb9_0;
	wire w_dff_A_BypINXjO1_0;
	wire w_dff_A_w2M4RpAV5_0;
	wire w_dff_A_w4BLgTFP6_0;
	wire w_dff_A_hkIpvIyN3_0;
	wire w_dff_A_by0cmANi0_0;
	wire w_dff_A_gKUxMeCj6_0;
	wire w_dff_A_yIdPt0dq0_0;
	wire w_dff_A_k6mVzKPC9_0;
	wire w_dff_A_OGdVz8h07_0;
	wire w_dff_A_JR1LEqV33_0;
	wire w_dff_A_oA4uXYQI7_0;
	wire w_dff_A_YeIbYm5q5_0;
	wire w_dff_A_Fad9lO6K7_0;
	wire w_dff_A_fP4VwOhA7_0;
	wire w_dff_A_wPGXAP1T8_0;
	wire w_dff_A_X5uy6Ul89_0;
	wire w_dff_A_5MU8qTkR3_0;
	wire w_dff_A_mta8aeIC9_0;
	wire w_dff_A_lCezDUmS6_0;
	wire w_dff_A_GE9EpR9Y7_0;
	wire w_dff_A_gbC5Q28i4_0;
	wire w_dff_A_oOrZQhdc6_0;
	wire w_dff_A_MshdEHUA3_0;
	wire w_dff_A_GTVZegty5_0;
	wire w_dff_A_upm7cW246_0;
	wire w_dff_A_sFSjVZGK3_0;
	wire w_dff_A_Hs4VEL4d4_0;
	wire w_dff_A_sOsttbQ18_0;
	wire w_dff_A_YYe81kyk5_0;
	wire w_dff_A_9BGgxj7j8_0;
	wire w_dff_A_vhGKTBuB6_0;
	wire w_dff_A_GNCaruMB7_0;
	wire w_dff_A_xye2GpFu8_0;
	wire w_dff_A_q4ossp9T8_0;
	wire w_dff_A_gQtgonkD1_0;
	wire w_dff_A_AbmdYSKy3_0;
	wire w_dff_A_NB4PiZFN3_0;
	wire w_dff_A_qTodR5Bt9_0;
	wire w_dff_A_Wt4m43OV1_0;
	wire w_dff_A_tRnFLsr66_0;
	wire w_dff_A_QTLzNcJ88_0;
	wire w_dff_A_wMLmqWG17_0;
	wire w_dff_A_eZVlgkM91_0;
	wire w_dff_A_CQOseGOU6_0;
	wire w_dff_A_7TdwLPkn1_0;
	wire w_dff_A_NCc31cjr8_0;
	wire w_dff_A_KRXCyJt87_0;
	wire w_dff_A_GkQWWBe95_0;
	wire w_dff_A_mkdNoieO8_0;
	wire w_dff_A_qGr3qz6b0_0;
	wire w_dff_A_9hMEaNkN1_0;
	wire w_dff_A_L6ecBm7o4_0;
	wire w_dff_A_TivH4GlN0_0;
	wire w_dff_A_vdxWXSlF0_0;
	wire w_dff_A_MelRwXzO6_0;
	wire w_dff_A_BR0LuR3Q9_0;
	wire w_dff_A_N1YXJyvb9_0;
	wire w_dff_A_gnlIbS416_0;
	wire w_dff_A_lkE8GRpU2_0;
	wire w_dff_A_XOL0iivq7_0;
	wire w_dff_A_5Gv1WFMd0_0;
	wire w_dff_A_nv1F8qll0_0;
	wire w_dff_A_t7giiDop1_0;
	wire w_dff_A_Io4Iw7zF1_0;
	wire w_dff_A_I3u4EcEE3_0;
	wire w_dff_A_DdJUbF8B1_0;
	wire w_dff_A_IJBDKL7L4_0;
	wire w_dff_A_FK59F2FA3_0;
	wire w_dff_A_nym5NQ194_2;
	wire w_dff_A_z8rrjKwU6_0;
	wire w_dff_A_I4QKR9tw3_0;
	wire w_dff_A_Qkr7HnZx3_0;
	wire w_dff_A_3eRx8es30_0;
	wire w_dff_A_qreLIVrI2_0;
	wire w_dff_A_DMbCWc4Y4_0;
	wire w_dff_A_wG63FlUr6_0;
	wire w_dff_A_qL5P0RMW8_0;
	wire w_dff_A_2bR3qjOS5_0;
	wire w_dff_A_LFSaiEVS3_0;
	wire w_dff_A_HlvMhO3J8_0;
	wire w_dff_A_RMJfd49g2_0;
	wire w_dff_A_CYTDBucW7_0;
	wire w_dff_A_SodQK0h88_0;
	wire w_dff_A_S8cMXxxy9_0;
	wire w_dff_A_K5EtG5RS6_0;
	wire w_dff_A_artkEDXD3_0;
	wire w_dff_A_Vly9DdtO7_0;
	wire w_dff_A_1kFvQbYh5_0;
	wire w_dff_A_XEVR1Y7w9_0;
	wire w_dff_A_ZPbTvxwl7_0;
	wire w_dff_A_BOSLCrtr8_0;
	wire w_dff_A_DHHMuR2n9_0;
	wire w_dff_A_qj7VCTNE5_0;
	wire w_dff_A_n0SqvMtf9_0;
	wire w_dff_A_gA2cuz2X1_0;
	wire w_dff_A_bYe5LaRl5_0;
	wire w_dff_A_LTMo0VBu4_0;
	wire w_dff_A_3KheANi86_0;
	wire w_dff_A_JdqDOIb96_0;
	wire w_dff_A_V9D0exUG8_0;
	wire w_dff_A_43DpmDBQ5_0;
	wire w_dff_A_8g3R5jU41_0;
	wire w_dff_A_medKfdVW2_0;
	wire w_dff_A_tMBVcawi7_0;
	wire w_dff_A_Qb1M4P9u9_0;
	wire w_dff_A_d2p1vxxE4_0;
	wire w_dff_A_yOyycVXV7_0;
	wire w_dff_A_nyf4qYJ29_0;
	wire w_dff_A_ODP5KXIC3_0;
	wire w_dff_A_8nOVQr7W5_0;
	wire w_dff_A_pfXDxnML3_0;
	wire w_dff_A_qP8o6VDr9_0;
	wire w_dff_A_LkUz6N6u9_0;
	wire w_dff_A_nlAmtiG30_0;
	wire w_dff_A_MaaPbLPz7_0;
	wire w_dff_A_7mtMJiAr6_0;
	wire w_dff_A_M5zgZ8059_0;
	wire w_dff_A_H2KMaoOE6_0;
	wire w_dff_A_GMgvfOpi1_0;
	wire w_dff_A_ggWpBlY67_0;
	wire w_dff_A_nKF4HeOX3_0;
	wire w_dff_A_hr0nIN654_0;
	wire w_dff_A_E8388oFY9_0;
	wire w_dff_A_IMqEEpQW4_0;
	wire w_dff_A_54XMmjVF9_0;
	wire w_dff_A_3MGLJkYM7_0;
	wire w_dff_A_l27ASzcF2_0;
	wire w_dff_A_IXlO26rX6_0;
	wire w_dff_A_jiV4oIti1_0;
	wire w_dff_A_IthNF00f4_0;
	wire w_dff_A_A0HzUWp40_0;
	wire w_dff_A_I4rSGf2Q4_0;
	wire w_dff_A_EMnpFW7I4_0;
	wire w_dff_A_SPFTZNXB6_0;
	wire w_dff_A_YHKBeXrG2_0;
	wire w_dff_A_xoIaY69s6_0;
	wire w_dff_A_GTIU1wQ27_0;
	wire w_dff_A_2cuCh8Y87_0;
	wire w_dff_A_vo8qKwrs9_0;
	wire w_dff_A_PfDLiwR91_0;
	wire w_dff_A_aQ8ttUdW6_0;
	wire w_dff_A_Y00BZPE67_0;
	wire w_dff_A_FVU385FV6_0;
	wire w_dff_A_28daTBMc4_0;
	wire w_dff_A_azsgFpCz9_0;
	wire w_dff_A_MQptl2Hn9_0;
	wire w_dff_A_BHMXI4SY3_0;
	wire w_dff_A_Cj3jlpbe7_0;
	wire w_dff_A_wvFR0Uve3_0;
	wire w_dff_A_JgJPasJh5_0;
	wire w_dff_A_N6lR6jMC6_0;
	wire w_dff_A_hhYbkQx20_0;
	wire w_dff_A_wKjpYrWy5_0;
	wire w_dff_A_ZeZ8qDSk1_0;
	wire w_dff_A_J2mufkAo7_0;
	wire w_dff_A_dB4bUQiS8_0;
	wire w_dff_A_JnsKETaU9_0;
	wire w_dff_A_PXMtGslz3_0;
	wire w_dff_A_4Rn8acWn9_2;
	wire w_dff_A_9ym0hURn8_0;
	wire w_dff_A_yvKFYDyW6_0;
	wire w_dff_A_rB3bBYAo8_0;
	wire w_dff_A_oPNcd0GF2_0;
	wire w_dff_A_NGB2M9Hx0_0;
	wire w_dff_A_WbLPtOR91_0;
	wire w_dff_A_Tan51rf57_0;
	wire w_dff_A_9LDDF9eD7_0;
	wire w_dff_A_oZC6NZOM0_0;
	wire w_dff_A_K9CinZsf7_0;
	wire w_dff_A_DSjOBXel1_0;
	wire w_dff_A_ycxBJLah5_0;
	wire w_dff_A_wxiRA0pH7_0;
	wire w_dff_A_mrlzsnng6_0;
	wire w_dff_A_eTtNNSoP9_0;
	wire w_dff_A_XsOaRDLz0_0;
	wire w_dff_A_vJWiNudq2_0;
	wire w_dff_A_LS9J4qHz0_0;
	wire w_dff_A_kakepyhG6_0;
	wire w_dff_A_gO8O1W7W3_0;
	wire w_dff_A_gVSjW9hB3_0;
	wire w_dff_A_tLv7LdDn5_0;
	wire w_dff_A_kDbAWkJD9_0;
	wire w_dff_A_VVQFFhE27_0;
	wire w_dff_A_Q6keX4yH6_0;
	wire w_dff_A_QxCZyVeY1_0;
	wire w_dff_A_pYp2jd4T7_0;
	wire w_dff_A_gefk1dwu5_0;
	wire w_dff_A_mDn3iTYk4_0;
	wire w_dff_A_vqwfpaBb5_0;
	wire w_dff_A_Y56fIn5Q0_0;
	wire w_dff_A_2T2wMx4o9_0;
	wire w_dff_A_X156pY411_0;
	wire w_dff_A_dgAWoQu22_0;
	wire w_dff_A_n9Uuorpr4_0;
	wire w_dff_A_JKTKpB1N1_0;
	wire w_dff_A_K3aRhSSR0_0;
	wire w_dff_A_NoKsbhUR5_0;
	wire w_dff_A_xenreQ6W3_0;
	wire w_dff_A_vQwwAsJD1_0;
	wire w_dff_A_SU4m2x337_0;
	wire w_dff_A_1PygVFLS0_0;
	wire w_dff_A_pF3xXOZR0_0;
	wire w_dff_A_EiAoH38c6_0;
	wire w_dff_A_IiF9nW1Z6_0;
	wire w_dff_A_jWIFUvVH0_0;
	wire w_dff_A_JrEEMHtX9_0;
	wire w_dff_A_0H0kz2tT0_0;
	wire w_dff_A_6FBUCSAl3_0;
	wire w_dff_A_r3JLqB512_0;
	wire w_dff_A_l4bRaizl6_0;
	wire w_dff_A_zJMehraY4_0;
	wire w_dff_A_SRFL3jk26_0;
	wire w_dff_A_quz5vkU68_0;
	wire w_dff_A_j5hplv7a5_0;
	wire w_dff_A_dLDI33Zv4_0;
	wire w_dff_A_YOUNvOLs8_0;
	wire w_dff_A_sjtAweMc6_0;
	wire w_dff_A_M2WtbFEk0_0;
	wire w_dff_A_uMYP7TBh0_0;
	wire w_dff_A_75g1qZ7J7_0;
	wire w_dff_A_weRWmR114_0;
	wire w_dff_A_tLhWpRaf3_0;
	wire w_dff_A_CpyKdXUj2_0;
	wire w_dff_A_3n6zaMjq7_0;
	wire w_dff_A_OeMeC6hR8_0;
	wire w_dff_A_VVtjRuJU5_0;
	wire w_dff_A_jt50o2VL2_0;
	wire w_dff_A_arD3n7N57_0;
	wire w_dff_A_KkJXCeBg6_0;
	wire w_dff_A_CwQrxJiv6_0;
	wire w_dff_A_m6Z1D3HT6_0;
	wire w_dff_A_KPaFgBGL2_0;
	wire w_dff_A_jpVJqQs63_0;
	wire w_dff_A_gLpbDhbH4_0;
	wire w_dff_A_x7EIawcx8_0;
	wire w_dff_A_RHxXTx2I8_0;
	wire w_dff_A_0nPt8unl8_0;
	wire w_dff_A_pH3EjJnN6_0;
	wire w_dff_A_459ve60a5_0;
	wire w_dff_A_UGa98vKo1_0;
	wire w_dff_A_mbKVm1rI9_0;
	wire w_dff_A_I10fOUxm7_0;
	wire w_dff_A_zmyJ6ohw2_0;
	wire w_dff_A_ulqR7j5G3_0;
	wire w_dff_A_5NYrJ0xk2_0;
	wire w_dff_A_7qSoFryb6_0;
	wire w_dff_A_fi0uRMCN2_0;
	wire w_dff_A_f746W3Pr1_2;
	wire w_dff_A_E1Mfhl4N4_0;
	wire w_dff_A_nAJmMpoC7_0;
	wire w_dff_A_2IQuxUlC9_0;
	wire w_dff_A_GFnFqxHF0_0;
	wire w_dff_A_HZzxVe5R7_0;
	wire w_dff_A_xIPXtjfh6_0;
	wire w_dff_A_RXBPeT6X3_0;
	wire w_dff_A_FspnMCwp2_0;
	wire w_dff_A_Gxfb6Dm70_0;
	wire w_dff_A_PyzkpODJ4_0;
	wire w_dff_A_zMxAzMzW4_0;
	wire w_dff_A_N89C6uF51_0;
	wire w_dff_A_U2YbtVln0_0;
	wire w_dff_A_LTjzwddC6_0;
	wire w_dff_A_s7wbO6Lb9_0;
	wire w_dff_A_RsstR8tj8_0;
	wire w_dff_A_H2ew9FRo0_0;
	wire w_dff_A_5lX0hUKw1_0;
	wire w_dff_A_cyLsIclr2_0;
	wire w_dff_A_JhO5zw7r0_0;
	wire w_dff_A_Uy8oZC2A1_0;
	wire w_dff_A_kgBQQ83n1_0;
	wire w_dff_A_r8NL11tE5_0;
	wire w_dff_A_8dAtUHwX9_0;
	wire w_dff_A_p51L4Dw08_0;
	wire w_dff_A_cH12S2Tx8_0;
	wire w_dff_A_Y3Kn1imC6_0;
	wire w_dff_A_3RkeztCx5_0;
	wire w_dff_A_wdQkdX3V4_0;
	wire w_dff_A_Jnch4fUi1_0;
	wire w_dff_A_z6PWRfF86_0;
	wire w_dff_A_EwKBplcw3_0;
	wire w_dff_A_l9ADmwb05_0;
	wire w_dff_A_AFILsLV16_0;
	wire w_dff_A_fqef3RN83_0;
	wire w_dff_A_0NBBSGke1_0;
	wire w_dff_A_epF3FsQ92_0;
	wire w_dff_A_RoRATiEh5_0;
	wire w_dff_A_1VL2fA4n8_0;
	wire w_dff_A_pkrC71cH4_0;
	wire w_dff_A_rl4ed3tV0_0;
	wire w_dff_A_nzrpFkXX7_0;
	wire w_dff_A_1h4k5g802_0;
	wire w_dff_A_hPVc5LxE5_0;
	wire w_dff_A_CxjkIRIS8_0;
	wire w_dff_A_yC9zI7aD6_0;
	wire w_dff_A_Z8kFUtuq4_0;
	wire w_dff_A_c8DXcmZi7_0;
	wire w_dff_A_wdUWkAd01_0;
	wire w_dff_A_0sYeAFDC2_0;
	wire w_dff_A_ckcRrgRj0_0;
	wire w_dff_A_t9wIPvBX3_0;
	wire w_dff_A_Kabk8kkV2_0;
	wire w_dff_A_gpdwEzTC9_0;
	wire w_dff_A_D4QrJoqY0_0;
	wire w_dff_A_w2rtCkcZ5_0;
	wire w_dff_A_NnX9lT930_0;
	wire w_dff_A_S1DvLhHm1_0;
	wire w_dff_A_iEoEVDmH4_0;
	wire w_dff_A_7gGC4gM24_0;
	wire w_dff_A_kqH80jDy3_0;
	wire w_dff_A_UPhesf4B9_0;
	wire w_dff_A_oppNHXX38_0;
	wire w_dff_A_aWjCQfwP4_0;
	wire w_dff_A_bsVY1f6c5_0;
	wire w_dff_A_qOnrAXDp1_0;
	wire w_dff_A_591tFOw36_0;
	wire w_dff_A_9sf7j4QP6_0;
	wire w_dff_A_sjwMV4JZ0_0;
	wire w_dff_A_NK0Uaf4n7_0;
	wire w_dff_A_OGGO79F78_0;
	wire w_dff_A_8pWyg9LJ3_0;
	wire w_dff_A_1BWoCeRx2_0;
	wire w_dff_A_ZSsTMc9r7_0;
	wire w_dff_A_1acBxVBM3_0;
	wire w_dff_A_aFoE6i4s8_0;
	wire w_dff_A_k9hEVnLb9_0;
	wire w_dff_A_p1Bx8YHV3_0;
	wire w_dff_A_mWnRbqn53_0;
	wire w_dff_A_HeGKQYiV1_0;
	wire w_dff_A_jJQY80bG2_0;
	wire w_dff_A_2VATXkln2_0;
	wire w_dff_A_V24kuI7C0_0;
	wire w_dff_A_ZAAuTILi3_0;
	wire w_dff_A_mpexeJvC7_0;
	wire w_dff_A_XgAcfQmd8_0;
	wire w_dff_A_if8icmPh1_0;
	wire w_dff_A_m6wDD8ja6_2;
	wire w_dff_A_BHl71OzP6_0;
	wire w_dff_A_S4GDVtfe7_0;
	wire w_dff_A_cRmTUQN44_0;
	wire w_dff_A_uWQhdzul9_0;
	wire w_dff_A_a5vYoFVz5_0;
	wire w_dff_A_rnPYtGdE9_0;
	wire w_dff_A_NLeXx2aM6_0;
	wire w_dff_A_MB8CsnD64_0;
	wire w_dff_A_o9waanZ98_0;
	wire w_dff_A_83Q7eVzm6_0;
	wire w_dff_A_MhHoKnEJ1_0;
	wire w_dff_A_qZx5AP5s3_0;
	wire w_dff_A_6gVuoz968_0;
	wire w_dff_A_clfWsd9i5_0;
	wire w_dff_A_4IrE0puv3_0;
	wire w_dff_A_7yK4No5Y2_0;
	wire w_dff_A_NNZst9LK6_0;
	wire w_dff_A_fS440rFR4_0;
	wire w_dff_A_2n9xBBUw3_0;
	wire w_dff_A_DgkeoheS6_0;
	wire w_dff_A_ZONus89Q2_0;
	wire w_dff_A_RXs2uRQk6_0;
	wire w_dff_A_iMfpHmTI1_0;
	wire w_dff_A_NGEBiC2z9_0;
	wire w_dff_A_XofUm5kU4_0;
	wire w_dff_A_EQsX8gc47_0;
	wire w_dff_A_bX8uZ8OQ0_0;
	wire w_dff_A_XthixKrH0_0;
	wire w_dff_A_mg4tjIf27_0;
	wire w_dff_A_7CHxDIrY9_0;
	wire w_dff_A_YJUfiYMX4_0;
	wire w_dff_A_MDdt7uyp0_0;
	wire w_dff_A_NoRviJwv3_0;
	wire w_dff_A_bcLj5S4W0_0;
	wire w_dff_A_iE0weS3a2_0;
	wire w_dff_A_OPQnamKv6_0;
	wire w_dff_A_AAQLtQEV3_0;
	wire w_dff_A_zoQbiNIp2_0;
	wire w_dff_A_QY7m5XD97_0;
	wire w_dff_A_IltStdH92_0;
	wire w_dff_A_ZmXyIiqy5_0;
	wire w_dff_A_qZMfuUDk2_0;
	wire w_dff_A_GsGgvVHS6_0;
	wire w_dff_A_wLewi5y66_0;
	wire w_dff_A_4PdaJDLe5_0;
	wire w_dff_A_CxMkWETV2_0;
	wire w_dff_A_MNSEKAZY8_0;
	wire w_dff_A_CIxn2oFn2_0;
	wire w_dff_A_sXMgN7PZ6_0;
	wire w_dff_A_KwnQ1ZhS6_0;
	wire w_dff_A_1MX8UB0b3_0;
	wire w_dff_A_PFFVTUPD0_0;
	wire w_dff_A_Rl1XKOgL6_0;
	wire w_dff_A_G2ptjs5y9_0;
	wire w_dff_A_m7hKvn1g7_0;
	wire w_dff_A_mKaa2Wjo9_0;
	wire w_dff_A_iAXsZpMl6_0;
	wire w_dff_A_oNiRWPRy6_0;
	wire w_dff_A_XiOtLwJA8_0;
	wire w_dff_A_w8IQmPQa7_0;
	wire w_dff_A_DoDLtp033_0;
	wire w_dff_A_ErMBmMqg0_0;
	wire w_dff_A_VtrilmPI6_0;
	wire w_dff_A_nes9wCju9_0;
	wire w_dff_A_aSF9Ppk55_0;
	wire w_dff_A_RfruNhaw6_0;
	wire w_dff_A_9wL3LaY63_0;
	wire w_dff_A_ZIXCrHd76_0;
	wire w_dff_A_5CPZt2DX2_0;
	wire w_dff_A_JjvqSUFo5_0;
	wire w_dff_A_ki65u2I14_0;
	wire w_dff_A_fMg8iQoO7_0;
	wire w_dff_A_Z7rjPR5j1_0;
	wire w_dff_A_fUzznTMX5_0;
	wire w_dff_A_DKGdcBaW3_0;
	wire w_dff_A_jEmefuQ65_0;
	wire w_dff_A_DfENg6Lk5_0;
	wire w_dff_A_GrHit8J09_0;
	wire w_dff_A_C22bGiM54_0;
	wire w_dff_A_wn6vPOZK6_0;
	wire w_dff_A_hioXIX2W7_0;
	wire w_dff_A_TtlENguc7_0;
	wire w_dff_A_S0rUy7ha6_0;
	wire w_dff_A_MARckjvl6_0;
	wire w_dff_A_Uie4O28Q1_0;
	wire w_dff_A_0pMDkLN33_0;
	wire w_dff_A_6JBK2nPW1_2;
	wire w_dff_A_Ig44NJbk9_0;
	wire w_dff_A_LRmVccAH5_0;
	wire w_dff_A_Am39zBpf9_0;
	wire w_dff_A_q6bkMG3r5_0;
	wire w_dff_A_ofzib6Ux9_0;
	wire w_dff_A_7zVHYnFG1_0;
	wire w_dff_A_9GPFFWsn2_0;
	wire w_dff_A_RwRYpOlV1_0;
	wire w_dff_A_eUeSG9P08_0;
	wire w_dff_A_XahTCvEH2_0;
	wire w_dff_A_eElY7Vk07_0;
	wire w_dff_A_CFuzPRoq3_0;
	wire w_dff_A_HCXVOM8T0_0;
	wire w_dff_A_dmlUJlRM8_0;
	wire w_dff_A_0BVAuxGp3_0;
	wire w_dff_A_9SlYBCUY1_0;
	wire w_dff_A_6E7u8WM83_0;
	wire w_dff_A_GGuJuZlR5_0;
	wire w_dff_A_MTP2Fc0D0_0;
	wire w_dff_A_TzeoYon48_0;
	wire w_dff_A_wVUOj4Hb5_0;
	wire w_dff_A_bxlmQx078_0;
	wire w_dff_A_0yjJIeKB8_0;
	wire w_dff_A_pIANq9rP9_0;
	wire w_dff_A_vniFLQhn9_0;
	wire w_dff_A_HLNnf8aX0_0;
	wire w_dff_A_SUcwoulU3_0;
	wire w_dff_A_bzGrdG5L8_0;
	wire w_dff_A_3trIzNcl2_0;
	wire w_dff_A_6wlYvITz1_0;
	wire w_dff_A_RFj2KSND7_0;
	wire w_dff_A_aYNYGUpa4_0;
	wire w_dff_A_9VJhQXUh0_0;
	wire w_dff_A_xvgY8m9d7_0;
	wire w_dff_A_ernyu3e28_0;
	wire w_dff_A_4uFfwBbG9_0;
	wire w_dff_A_mckkwymu8_0;
	wire w_dff_A_weLrtYMy0_0;
	wire w_dff_A_vRFb8hrF5_0;
	wire w_dff_A_GP5KH0aN7_0;
	wire w_dff_A_0YryPYix4_0;
	wire w_dff_A_Idl9YaUA0_0;
	wire w_dff_A_YuSX56it9_0;
	wire w_dff_A_RNJFjpIk6_0;
	wire w_dff_A_p0UhPUEZ0_0;
	wire w_dff_A_HNCAy7Cb2_0;
	wire w_dff_A_SqR5GScA3_0;
	wire w_dff_A_zCCKVcRW1_0;
	wire w_dff_A_Qevygbzi0_0;
	wire w_dff_A_pGSbur8B1_0;
	wire w_dff_A_JXc14ZzH6_0;
	wire w_dff_A_Xa9PaJDy1_0;
	wire w_dff_A_JodmWguB4_0;
	wire w_dff_A_1VCMknYK8_0;
	wire w_dff_A_xPOqCAD35_0;
	wire w_dff_A_JGEFaSEz3_0;
	wire w_dff_A_bTiUZa0d0_0;
	wire w_dff_A_bFtFCiV93_0;
	wire w_dff_A_JDnTg7Wy2_0;
	wire w_dff_A_0xGYnvYT9_0;
	wire w_dff_A_Rx2AkfOZ7_0;
	wire w_dff_A_Id7s039g1_0;
	wire w_dff_A_FeHNKsXG8_0;
	wire w_dff_A_373RZLtH2_0;
	wire w_dff_A_cy6TiKAY7_0;
	wire w_dff_A_zqHffu1C6_0;
	wire w_dff_A_yBIXVU8B0_0;
	wire w_dff_A_hohG6Ava7_0;
	wire w_dff_A_YrozW7jp0_0;
	wire w_dff_A_ozpiGovK3_0;
	wire w_dff_A_dqAuvGf84_0;
	wire w_dff_A_MjaYf2H42_0;
	wire w_dff_A_fh10UvDM3_0;
	wire w_dff_A_GftTKNNO5_0;
	wire w_dff_A_LOkLnOjh0_0;
	wire w_dff_A_vKPllyVC5_0;
	wire w_dff_A_d0RxXPR64_0;
	wire w_dff_A_QvVkHKpg3_0;
	wire w_dff_A_GaRmSQ3Z4_0;
	wire w_dff_A_MLa1aEM94_0;
	wire w_dff_A_npUhE63i2_0;
	wire w_dff_A_h3uBRfXY5_0;
	wire w_dff_A_UrcCR59f5_0;
	wire w_dff_A_wWJe65Pb1_0;
	wire w_dff_A_j2CmVjSk5_0;
	wire w_dff_A_09ujqjlu8_2;
	wire w_dff_A_be74fz819_0;
	wire w_dff_A_I8xteb4F9_0;
	wire w_dff_A_VGF7z3iy1_0;
	wire w_dff_A_sDZi5Mfg2_0;
	wire w_dff_A_tbda1U0P4_0;
	wire w_dff_A_MufNjFSd8_0;
	wire w_dff_A_DlmJ5lzi0_0;
	wire w_dff_A_WVLj8wRy6_0;
	wire w_dff_A_xtE0Ueya9_0;
	wire w_dff_A_bjSse2pa1_0;
	wire w_dff_A_hoWIJ4us4_0;
	wire w_dff_A_upKxRkym8_0;
	wire w_dff_A_RJCqsJvr3_0;
	wire w_dff_A_nzmIOttB8_0;
	wire w_dff_A_UeRAWBye8_0;
	wire w_dff_A_kiyyZw0H3_0;
	wire w_dff_A_JCNxAO7s4_0;
	wire w_dff_A_SEjjlhd79_0;
	wire w_dff_A_dPGrPTZq1_0;
	wire w_dff_A_pXA8IV9V3_0;
	wire w_dff_A_CKqMEaNF6_0;
	wire w_dff_A_aQhVcq0b3_0;
	wire w_dff_A_hRhEXDo67_0;
	wire w_dff_A_LrdEYM1a5_0;
	wire w_dff_A_AjIxpUJS5_0;
	wire w_dff_A_BnDQLnGE7_0;
	wire w_dff_A_Jnzh4Z970_0;
	wire w_dff_A_LIVMCQeI7_0;
	wire w_dff_A_9bO3gilc0_0;
	wire w_dff_A_91CtK90a0_0;
	wire w_dff_A_0V7efWrM5_0;
	wire w_dff_A_KO6zhEyl8_0;
	wire w_dff_A_zgXRiywV5_0;
	wire w_dff_A_zGfviu9u3_0;
	wire w_dff_A_66rZtyR85_0;
	wire w_dff_A_CLw6JZE77_0;
	wire w_dff_A_tO3ncZsQ3_0;
	wire w_dff_A_zhxgy1SI9_0;
	wire w_dff_A_F02IGJHi6_0;
	wire w_dff_A_vlgSZwsw9_0;
	wire w_dff_A_QvmUDdwW1_0;
	wire w_dff_A_qs5sUFd54_0;
	wire w_dff_A_tvvEPsvj5_0;
	wire w_dff_A_m2rz8ZOa0_0;
	wire w_dff_A_7b5xt8Jb6_0;
	wire w_dff_A_RMLMDYql2_0;
	wire w_dff_A_RxVrpxhD1_0;
	wire w_dff_A_KsCP3sLU8_0;
	wire w_dff_A_CgPlzuhz8_0;
	wire w_dff_A_cNLxJw9X6_0;
	wire w_dff_A_fniQDc2H5_0;
	wire w_dff_A_9xlETZAD4_0;
	wire w_dff_A_JL50S49p1_0;
	wire w_dff_A_MlwASfw96_0;
	wire w_dff_A_dygkZ9gN4_0;
	wire w_dff_A_7NS9T6Ij1_0;
	wire w_dff_A_ArA2uCLg4_0;
	wire w_dff_A_jCK4P6Gw0_0;
	wire w_dff_A_V7HGuMDS9_0;
	wire w_dff_A_LCFq9c2U4_0;
	wire w_dff_A_RhWuPDMP0_0;
	wire w_dff_A_UrqmSOGO9_0;
	wire w_dff_A_B6kVDOoH6_0;
	wire w_dff_A_u49tUYXQ0_0;
	wire w_dff_A_VSIPmh6y8_0;
	wire w_dff_A_OAqUtPXc4_0;
	wire w_dff_A_OFsA9OWJ8_0;
	wire w_dff_A_ic1PIJyN5_0;
	wire w_dff_A_zckYKGVP9_0;
	wire w_dff_A_vdsyRhqH3_0;
	wire w_dff_A_zp7XrHna3_0;
	wire w_dff_A_CvWdVhc81_0;
	wire w_dff_A_30dp7QUw0_0;
	wire w_dff_A_JYfTop5S5_0;
	wire w_dff_A_CTAMHKIb9_0;
	wire w_dff_A_3NHchMO86_0;
	wire w_dff_A_YhkumKvG9_0;
	wire w_dff_A_8gLtMPJH2_0;
	wire w_dff_A_1KkeRVA44_0;
	wire w_dff_A_E6sukExO1_0;
	wire w_dff_A_muRFRCui3_0;
	wire w_dff_A_ouyj3V846_0;
	wire w_dff_A_pwOQZeRs9_0;
	wire w_dff_A_mr6hoPYX7_0;
	wire w_dff_A_I2YmvXsD7_2;
	wire w_dff_A_iwwCAYjP4_0;
	wire w_dff_A_9p7EbxrT3_0;
	wire w_dff_A_mBoupQAV6_0;
	wire w_dff_A_dazKTbJF6_0;
	wire w_dff_A_YV3D9fTu4_0;
	wire w_dff_A_5ICCUItY9_0;
	wire w_dff_A_KAtL8Svj9_0;
	wire w_dff_A_o0tbN3Rf5_0;
	wire w_dff_A_3aglvj2B9_0;
	wire w_dff_A_0QZOk1Tt1_0;
	wire w_dff_A_RlsEu0s89_0;
	wire w_dff_A_mrf5lEzd8_0;
	wire w_dff_A_K7n24jrx6_0;
	wire w_dff_A_KhX8Zs792_0;
	wire w_dff_A_8XcG8xDf8_0;
	wire w_dff_A_fRkOhPgT2_0;
	wire w_dff_A_1Aflo9lq5_0;
	wire w_dff_A_Z1ZPN1hd9_0;
	wire w_dff_A_Aj3mC7Yq8_0;
	wire w_dff_A_ctIBh6Wp8_0;
	wire w_dff_A_zuvrfReM5_0;
	wire w_dff_A_xOdwzxux1_0;
	wire w_dff_A_IVGsGoaU6_0;
	wire w_dff_A_0WhriuVL4_0;
	wire w_dff_A_CQDIP57e0_0;
	wire w_dff_A_jTXsJJre9_0;
	wire w_dff_A_ivmbgxt15_0;
	wire w_dff_A_oF0LvA588_0;
	wire w_dff_A_YaiEmU210_0;
	wire w_dff_A_ePXmgAeT0_0;
	wire w_dff_A_CrFaqAzs6_0;
	wire w_dff_A_sd9WIwLu6_0;
	wire w_dff_A_cyhdTi2s7_0;
	wire w_dff_A_Ebrbe4Ro5_0;
	wire w_dff_A_oUJM2Xul3_0;
	wire w_dff_A_BbnissWg5_0;
	wire w_dff_A_EG7x2Eyy4_0;
	wire w_dff_A_wV8ZhxCo5_0;
	wire w_dff_A_47GtF05j5_0;
	wire w_dff_A_loQ3y2CI1_0;
	wire w_dff_A_8PssS20B1_0;
	wire w_dff_A_dxvju1Yp4_0;
	wire w_dff_A_5GFDt7Em0_0;
	wire w_dff_A_vf1L7Tlg0_0;
	wire w_dff_A_jMxMaCax5_0;
	wire w_dff_A_y0aBSAA14_0;
	wire w_dff_A_UcENqhBs2_0;
	wire w_dff_A_8i7DLpwY8_0;
	wire w_dff_A_lLY9jVsG9_0;
	wire w_dff_A_KVDN2Mls1_0;
	wire w_dff_A_68UTzHBK5_0;
	wire w_dff_A_4qDqqGwG1_0;
	wire w_dff_A_kHXU97Lc7_0;
	wire w_dff_A_XpPYjHLw5_0;
	wire w_dff_A_flJKFsXs7_0;
	wire w_dff_A_D7MGyajg3_0;
	wire w_dff_A_phhfLAtf2_0;
	wire w_dff_A_lEEZB3fQ8_0;
	wire w_dff_A_KDeHjTUE0_0;
	wire w_dff_A_Bbf8bry06_0;
	wire w_dff_A_bohYFnGH5_0;
	wire w_dff_A_EicDp3dW2_0;
	wire w_dff_A_gRCiM6iH3_0;
	wire w_dff_A_P87bsD3U0_0;
	wire w_dff_A_58f8sd3p0_0;
	wire w_dff_A_YhN4a1Q65_0;
	wire w_dff_A_egnquzXW2_0;
	wire w_dff_A_dXhZkiuG8_0;
	wire w_dff_A_JHVMi7LS0_0;
	wire w_dff_A_QzZnwF7e5_0;
	wire w_dff_A_6HgVXsN02_0;
	wire w_dff_A_hbakRN0M2_0;
	wire w_dff_A_QAEXknsg6_0;
	wire w_dff_A_QnYlALgD3_0;
	wire w_dff_A_J769Eo012_0;
	wire w_dff_A_dIiHWuHW0_0;
	wire w_dff_A_awPYj27s3_0;
	wire w_dff_A_6RgqpFib8_0;
	wire w_dff_A_FgVjMgpT8_0;
	wire w_dff_A_Fhux8ibn9_0;
	wire w_dff_A_ExWud07P6_0;
	wire w_dff_A_yDKO6jnY6_0;
	wire w_dff_A_i9TXfYjA3_0;
	wire w_dff_A_QwZFXhVA9_2;
	wire w_dff_A_nvkloFpO9_0;
	wire w_dff_A_LbIgM0Sr3_0;
	wire w_dff_A_H0iNvINO7_0;
	wire w_dff_A_RundX8An2_0;
	wire w_dff_A_9rxmYfdH1_0;
	wire w_dff_A_xFel332I6_0;
	wire w_dff_A_af9wKAWX3_0;
	wire w_dff_A_YsM1BgCH8_0;
	wire w_dff_A_GadyavqL7_0;
	wire w_dff_A_xEiZUlON1_0;
	wire w_dff_A_mUMsLDWr3_0;
	wire w_dff_A_ZVXD2CPn3_0;
	wire w_dff_A_JSxkZfCp4_0;
	wire w_dff_A_AmTlAO325_0;
	wire w_dff_A_Pvxw8xvc6_0;
	wire w_dff_A_81QK1hPd9_0;
	wire w_dff_A_GOB7TVp82_0;
	wire w_dff_A_Yli3KqZy3_0;
	wire w_dff_A_yfOL9Q0B2_0;
	wire w_dff_A_vLarxcGg2_0;
	wire w_dff_A_xe0yl61c4_0;
	wire w_dff_A_uTizlrAL6_0;
	wire w_dff_A_ku1iD0Y45_0;
	wire w_dff_A_EGR2RRYy4_0;
	wire w_dff_A_Zcrx2RQa9_0;
	wire w_dff_A_s9LAINHP7_0;
	wire w_dff_A_2z9xenZG0_0;
	wire w_dff_A_NoDevIiG5_0;
	wire w_dff_A_KuJ735h86_0;
	wire w_dff_A_aQ3KPV1F1_0;
	wire w_dff_A_B6ElxsZl8_0;
	wire w_dff_A_b7mtH4VV7_0;
	wire w_dff_A_q3qkhjU29_0;
	wire w_dff_A_4u9iplea2_0;
	wire w_dff_A_9EGFBIGa0_0;
	wire w_dff_A_K4YooPV45_0;
	wire w_dff_A_l7cCkc5d2_0;
	wire w_dff_A_sOC4NZV84_0;
	wire w_dff_A_PuxORUE67_0;
	wire w_dff_A_CDTko9DL1_0;
	wire w_dff_A_WFz45bpl7_0;
	wire w_dff_A_boFmAM0m4_0;
	wire w_dff_A_acxQhCmO9_0;
	wire w_dff_A_blJxPUGY0_0;
	wire w_dff_A_Aig1CN4X5_0;
	wire w_dff_A_VbChy4NS9_0;
	wire w_dff_A_hDHVBNZY4_0;
	wire w_dff_A_iOHFtmFf5_0;
	wire w_dff_A_2MTiY6nB1_0;
	wire w_dff_A_1n4N6PNy0_0;
	wire w_dff_A_BctyuwEo3_0;
	wire w_dff_A_TNhBJMbf5_0;
	wire w_dff_A_xUUKkhNU0_0;
	wire w_dff_A_6orM6LHi7_0;
	wire w_dff_A_MwbP0iqd2_0;
	wire w_dff_A_CljpVI755_0;
	wire w_dff_A_XZcBWpOe8_0;
	wire w_dff_A_N6QmLFWO4_0;
	wire w_dff_A_9XtA2kaC0_0;
	wire w_dff_A_jhlepn2y3_0;
	wire w_dff_A_hjDgVkUM7_0;
	wire w_dff_A_m1JHBSk70_0;
	wire w_dff_A_IunuhWCv9_0;
	wire w_dff_A_y8jHW5686_0;
	wire w_dff_A_aWhpgFXZ8_0;
	wire w_dff_A_Ze0Tjzul6_0;
	wire w_dff_A_Tvg1wBCr4_0;
	wire w_dff_A_GvUqMuMM9_0;
	wire w_dff_A_PgcqJA811_0;
	wire w_dff_A_51nk0jiv9_0;
	wire w_dff_A_QLhtEXxF2_0;
	wire w_dff_A_EQqmmGRC4_0;
	wire w_dff_A_PNHhgyPK1_0;
	wire w_dff_A_NAGUwB5e0_0;
	wire w_dff_A_AkjmE9m44_0;
	wire w_dff_A_PJpTeiGq5_0;
	wire w_dff_A_pss17xV59_0;
	wire w_dff_A_Q9GGttvB4_0;
	wire w_dff_A_wP2gzpTS6_0;
	wire w_dff_A_sDTcExYP1_0;
	wire w_dff_A_spfe5KAf1_0;
	wire w_dff_A_liL365568_0;
	wire w_dff_A_VA8FezrL8_2;
	wire w_dff_A_b226qRnN3_0;
	wire w_dff_A_pZPQjE2g3_0;
	wire w_dff_A_8iIdkfKF8_0;
	wire w_dff_A_o1GZ0zij0_0;
	wire w_dff_A_if8Baa843_0;
	wire w_dff_A_UAz8SeHi6_0;
	wire w_dff_A_sg4Csuqz8_0;
	wire w_dff_A_4o1VsA5K8_0;
	wire w_dff_A_iCI7vs3b9_0;
	wire w_dff_A_UMYRLIK44_0;
	wire w_dff_A_oYqbKALq1_0;
	wire w_dff_A_y2unAVqf9_0;
	wire w_dff_A_gI3iWxhH5_0;
	wire w_dff_A_wMP0kDfA4_0;
	wire w_dff_A_aYdScR2t7_0;
	wire w_dff_A_XCCaEhXv4_0;
	wire w_dff_A_1uG86Qwl6_0;
	wire w_dff_A_xRbjSe2j1_0;
	wire w_dff_A_SmxzjB9o1_0;
	wire w_dff_A_OPR2Dgfc7_0;
	wire w_dff_A_2g2TVycB8_0;
	wire w_dff_A_vIvx6jIH3_0;
	wire w_dff_A_eRmnPQA45_0;
	wire w_dff_A_zz7xbobE6_0;
	wire w_dff_A_GNkl9cSO1_0;
	wire w_dff_A_dLlbPJj91_0;
	wire w_dff_A_HsZ4XLDi9_0;
	wire w_dff_A_lnF6INVy1_0;
	wire w_dff_A_PtH2FU308_0;
	wire w_dff_A_bLRHLw6I0_0;
	wire w_dff_A_qTs8cf0U2_0;
	wire w_dff_A_4AX9puio9_0;
	wire w_dff_A_gJHyPL2e9_0;
	wire w_dff_A_WisRR6O13_0;
	wire w_dff_A_19Do98xE4_0;
	wire w_dff_A_kczk54597_0;
	wire w_dff_A_myTyPijs6_0;
	wire w_dff_A_4kvYeWPA1_0;
	wire w_dff_A_S9e7LfMG8_0;
	wire w_dff_A_XgxjNJ0K7_0;
	wire w_dff_A_FKlQSajr2_0;
	wire w_dff_A_xedhvIKq8_0;
	wire w_dff_A_LvhQ5N1D1_0;
	wire w_dff_A_LtTvRMsL8_0;
	wire w_dff_A_w4u5U6lP8_0;
	wire w_dff_A_4SoVkHw83_0;
	wire w_dff_A_uI1Xt1Ht0_0;
	wire w_dff_A_2xt2lJfA0_0;
	wire w_dff_A_VJFz8Uom7_0;
	wire w_dff_A_4mVtzz5I9_0;
	wire w_dff_A_Jh0Pbxth0_0;
	wire w_dff_A_ep2o8L4k1_0;
	wire w_dff_A_ZfGnjXiW7_0;
	wire w_dff_A_pWPCIsz71_0;
	wire w_dff_A_catsBTZK1_0;
	wire w_dff_A_mlRZ4bO28_0;
	wire w_dff_A_CTOicfeF0_0;
	wire w_dff_A_TJ5n8bcQ7_0;
	wire w_dff_A_laPYLZzS2_0;
	wire w_dff_A_4FOur9j23_0;
	wire w_dff_A_Sf8DfBWg5_0;
	wire w_dff_A_zbu4IAnq0_0;
	wire w_dff_A_58knblez0_0;
	wire w_dff_A_1rYtvV0Z8_0;
	wire w_dff_A_F8kjRSmg6_0;
	wire w_dff_A_lPw9gapI9_0;
	wire w_dff_A_dfkK1r7m6_0;
	wire w_dff_A_SeZGPuyv4_0;
	wire w_dff_A_HZStFoNn9_0;
	wire w_dff_A_KIP5wquy5_0;
	wire w_dff_A_HXrZOhLr9_0;
	wire w_dff_A_Znn79pgt7_0;
	wire w_dff_A_3sEmRykW0_0;
	wire w_dff_A_Qlwi5kWE7_0;
	wire w_dff_A_6t05PBfO9_0;
	wire w_dff_A_hNUpVLeR7_0;
	wire w_dff_A_9yqlOFht4_0;
	wire w_dff_A_pskIfvvL5_0;
	wire w_dff_A_6FTNQ2Kh1_0;
	wire w_dff_A_uhHD4lyL4_0;
	wire w_dff_A_aDYoSPHZ4_0;
	wire w_dff_A_HG05Fu3s6_2;
	wire w_dff_A_1Y3ZXEOD9_0;
	wire w_dff_A_rsaC8EOD4_0;
	wire w_dff_A_yJa8GiY56_0;
	wire w_dff_A_d2U2JZ351_0;
	wire w_dff_A_eiabcs987_0;
	wire w_dff_A_oT8JnhJB9_0;
	wire w_dff_A_4O6DHlfK5_0;
	wire w_dff_A_Axp9Kb249_0;
	wire w_dff_A_JtWxbxBH8_0;
	wire w_dff_A_BNiSuHog3_0;
	wire w_dff_A_Itc1YIAW7_0;
	wire w_dff_A_YKCK1I1K7_0;
	wire w_dff_A_JjPsMhjR4_0;
	wire w_dff_A_vSPqQAyF0_0;
	wire w_dff_A_m9NmUZsP0_0;
	wire w_dff_A_WCnoFlRp1_0;
	wire w_dff_A_q1nV2qLW9_0;
	wire w_dff_A_QYTzw6fn8_0;
	wire w_dff_A_3b2N48St1_0;
	wire w_dff_A_QvS2scxK0_0;
	wire w_dff_A_cj63GRbJ6_0;
	wire w_dff_A_qGrn4L5R4_0;
	wire w_dff_A_nTSRAmSa6_0;
	wire w_dff_A_BOoo0Xz64_0;
	wire w_dff_A_7q1MmhDE7_0;
	wire w_dff_A_pbsXAUVu7_0;
	wire w_dff_A_NNkfLj2L5_0;
	wire w_dff_A_JSNZxt6X2_0;
	wire w_dff_A_UjzPN8SU4_0;
	wire w_dff_A_qEJrqRI55_0;
	wire w_dff_A_38cUQZwu9_0;
	wire w_dff_A_cfAXH0Q49_0;
	wire w_dff_A_ezuQ3fGf2_0;
	wire w_dff_A_7hofpAoX7_0;
	wire w_dff_A_44GbYigZ9_0;
	wire w_dff_A_17OAx2DH4_0;
	wire w_dff_A_8TO0W6bo3_0;
	wire w_dff_A_fczQbtFl7_0;
	wire w_dff_A_NdHswp9u8_0;
	wire w_dff_A_yEneimwF9_0;
	wire w_dff_A_4owuKtWK4_0;
	wire w_dff_A_RwptPYlL4_0;
	wire w_dff_A_LDHXtFyS9_0;
	wire w_dff_A_7dAVMnmv3_0;
	wire w_dff_A_orhT70XV3_0;
	wire w_dff_A_GHWlDHQF7_0;
	wire w_dff_A_F0gPMduf0_0;
	wire w_dff_A_Kh7bOlBZ0_0;
	wire w_dff_A_4SMjnric5_0;
	wire w_dff_A_HEtPXXun2_0;
	wire w_dff_A_hU4xo7TJ9_0;
	wire w_dff_A_cNq82MEO3_0;
	wire w_dff_A_v9ERO0Hi2_0;
	wire w_dff_A_p6fawIhc5_0;
	wire w_dff_A_xjzdKE530_0;
	wire w_dff_A_72mGvg8Z2_0;
	wire w_dff_A_aZYbpUCt3_0;
	wire w_dff_A_ISOq6j5g6_0;
	wire w_dff_A_wHy9NTg48_0;
	wire w_dff_A_ko4ok0sf2_0;
	wire w_dff_A_U4Jpn1HQ1_0;
	wire w_dff_A_ymMe0Kz95_0;
	wire w_dff_A_4g7pn8cp7_0;
	wire w_dff_A_h9ctqVME7_0;
	wire w_dff_A_AIfM2gNc4_0;
	wire w_dff_A_Q59DK8NO1_0;
	wire w_dff_A_KdUAUdq19_0;
	wire w_dff_A_FX5IWUoc2_0;
	wire w_dff_A_q7cZZz3O8_0;
	wire w_dff_A_3On6WqYB1_0;
	wire w_dff_A_63tcd6cp9_0;
	wire w_dff_A_7iAXgQrL4_0;
	wire w_dff_A_2JdxGfgq4_0;
	wire w_dff_A_LycyT0BB9_0;
	wire w_dff_A_B1YASNI46_0;
	wire w_dff_A_lQ5xWwDV2_0;
	wire w_dff_A_UQL8PhEg0_0;
	wire w_dff_A_dqLrMj3M3_0;
	wire w_dff_A_cSsadq7C0_0;
	wire w_dff_A_WLW2og5L4_0;
	wire w_dff_A_AIhCfEsq4_2;
	wire w_dff_A_Mcd8r44t0_0;
	wire w_dff_A_Qz76Zm9s4_0;
	wire w_dff_A_2G23Zo3b2_0;
	wire w_dff_A_pwAFPXiY0_0;
	wire w_dff_A_VJQ4SxBm8_0;
	wire w_dff_A_LBYLBaZf6_0;
	wire w_dff_A_npyf1nAS8_0;
	wire w_dff_A_x4ZsDeE40_0;
	wire w_dff_A_pb2gld0l1_0;
	wire w_dff_A_m0P8Dk0L5_0;
	wire w_dff_A_LKxYA0WB2_0;
	wire w_dff_A_MJpTqKJE0_0;
	wire w_dff_A_k1udsWbK9_0;
	wire w_dff_A_oWtbHikt8_0;
	wire w_dff_A_QUJegnHs2_0;
	wire w_dff_A_BPIXwtwp8_0;
	wire w_dff_A_11srEgQN9_0;
	wire w_dff_A_DbDtTKK26_0;
	wire w_dff_A_uztct3wy2_0;
	wire w_dff_A_IsPJJbj62_0;
	wire w_dff_A_ulaPoL4U6_0;
	wire w_dff_A_JEDaHwzL6_0;
	wire w_dff_A_XgUakTwu2_0;
	wire w_dff_A_yVBiuFpG4_0;
	wire w_dff_A_Zkot34Qt5_0;
	wire w_dff_A_GuYhh4d83_0;
	wire w_dff_A_pzCSfwi07_0;
	wire w_dff_A_AqDyW98h9_0;
	wire w_dff_A_aXjtoTK27_0;
	wire w_dff_A_CyR4yuNj0_0;
	wire w_dff_A_JnkblOjK9_0;
	wire w_dff_A_CY9bIOQj4_0;
	wire w_dff_A_eKWNEgVB3_0;
	wire w_dff_A_axhDMKbh6_0;
	wire w_dff_A_Fz6TVdNW7_0;
	wire w_dff_A_Dr6sawMl5_0;
	wire w_dff_A_I2VRxduo4_0;
	wire w_dff_A_Go1GYNxA0_0;
	wire w_dff_A_y8QegFjn5_0;
	wire w_dff_A_TLN9vnk87_0;
	wire w_dff_A_Uq4FoVBv9_0;
	wire w_dff_A_W2W9dNqC7_0;
	wire w_dff_A_x2objUkJ2_0;
	wire w_dff_A_H9VUiw3e3_0;
	wire w_dff_A_ZoFSIXa75_0;
	wire w_dff_A_396Ek8fd9_0;
	wire w_dff_A_uqgLOtsS9_0;
	wire w_dff_A_QeEHURnA2_0;
	wire w_dff_A_BYUnO9Sh1_0;
	wire w_dff_A_3HYrIsu11_0;
	wire w_dff_A_1Cox9EfY1_0;
	wire w_dff_A_vHYudDBo5_0;
	wire w_dff_A_YqHoSDXs5_0;
	wire w_dff_A_9790vaaC0_0;
	wire w_dff_A_gvXChzq40_0;
	wire w_dff_A_T56Os9rB3_0;
	wire w_dff_A_7x7hpyfc0_0;
	wire w_dff_A_4VmKR2rn3_0;
	wire w_dff_A_6pZ9RTP72_0;
	wire w_dff_A_qXLvXRzj6_0;
	wire w_dff_A_o8iW57Rc1_0;
	wire w_dff_A_4cUt3PnS1_0;
	wire w_dff_A_oa0VrNQq6_0;
	wire w_dff_A_be0FEAY46_0;
	wire w_dff_A_uTgQXcrR3_0;
	wire w_dff_A_0xZV8J2l9_0;
	wire w_dff_A_o13xOGmh6_0;
	wire w_dff_A_GgOvRwNH3_0;
	wire w_dff_A_n1h1dw9K3_0;
	wire w_dff_A_lVS80qA86_0;
	wire w_dff_A_fk6lzoKa2_0;
	wire w_dff_A_BEdpB4C30_0;
	wire w_dff_A_b1dLA96G0_0;
	wire w_dff_A_QR4EX62S0_0;
	wire w_dff_A_MFAyzbx46_0;
	wire w_dff_A_GVp1UVPk7_0;
	wire w_dff_A_PM5ZtlQD7_0;
	wire w_dff_A_2ycVZnh81_0;
	wire w_dff_A_tQit25iN5_0;
	wire w_dff_A_aJxExRy15_2;
	wire w_dff_A_NJQV6SZi2_0;
	wire w_dff_A_MhBca7KV1_0;
	wire w_dff_A_9OlWWsqQ2_0;
	wire w_dff_A_Zqv09oBS6_0;
	wire w_dff_A_VVASM3SG2_0;
	wire w_dff_A_YVPc6j3h6_0;
	wire w_dff_A_0z8fme2q7_0;
	wire w_dff_A_nGHTJf3E0_0;
	wire w_dff_A_JdMdHrXo9_0;
	wire w_dff_A_CjQsWB2y3_0;
	wire w_dff_A_61ToQZPn3_0;
	wire w_dff_A_7HDDk0Ny2_0;
	wire w_dff_A_CA81cROY1_0;
	wire w_dff_A_jDJVLSTG9_0;
	wire w_dff_A_Dukm22Qj1_0;
	wire w_dff_A_5wF390iD5_0;
	wire w_dff_A_XGe4BT3r3_0;
	wire w_dff_A_RedMbgfE6_0;
	wire w_dff_A_yORgae439_0;
	wire w_dff_A_2c5OQJUM8_0;
	wire w_dff_A_uumfmRZn3_0;
	wire w_dff_A_aAakDUJN0_0;
	wire w_dff_A_fl4wvd8T3_0;
	wire w_dff_A_kQ5Oqr6u0_0;
	wire w_dff_A_lrb8EH9h7_0;
	wire w_dff_A_SBhgyTjs2_0;
	wire w_dff_A_zq4e2W0W9_0;
	wire w_dff_A_6gFVf2vb0_0;
	wire w_dff_A_VAGS6w1e8_0;
	wire w_dff_A_p8DQ8MmW0_0;
	wire w_dff_A_SaFZpYw31_0;
	wire w_dff_A_2schEaM23_0;
	wire w_dff_A_WVuOI4ok0_0;
	wire w_dff_A_ZAWf4ALq5_0;
	wire w_dff_A_toFNROMF5_0;
	wire w_dff_A_OL7lrtJo9_0;
	wire w_dff_A_FJXgFxuv3_0;
	wire w_dff_A_hnOh2mkZ4_0;
	wire w_dff_A_fsZYiXue4_0;
	wire w_dff_A_i19eDR6q7_0;
	wire w_dff_A_f8MnNG2o7_0;
	wire w_dff_A_Rc2w68Zs3_0;
	wire w_dff_A_Ng4GBPnK8_0;
	wire w_dff_A_SZzkyurj3_0;
	wire w_dff_A_sTSzT9z68_0;
	wire w_dff_A_i1cHP5Pz3_0;
	wire w_dff_A_ZOeMV3mx5_0;
	wire w_dff_A_BVmgYYX16_0;
	wire w_dff_A_Dcy9FYHD4_0;
	wire w_dff_A_53TW0JYo5_0;
	wire w_dff_A_kD4t3t1u3_0;
	wire w_dff_A_MjW4Y4X77_0;
	wire w_dff_A_jset7Hrp4_0;
	wire w_dff_A_bo5hM1YX6_0;
	wire w_dff_A_OeEAXBqx7_0;
	wire w_dff_A_gvOndYL90_0;
	wire w_dff_A_Sv6v8ZMG7_0;
	wire w_dff_A_SgPoUcIc4_0;
	wire w_dff_A_t5CxSU6p2_0;
	wire w_dff_A_2sxTJBzf2_0;
	wire w_dff_A_SCp9anKm5_0;
	wire w_dff_A_SilJIt3L9_0;
	wire w_dff_A_jdVbzgzD8_0;
	wire w_dff_A_Z2UORUHY9_0;
	wire w_dff_A_HV3OpqiV2_0;
	wire w_dff_A_sTbfWvpH0_0;
	wire w_dff_A_WIHKVHEv6_0;
	wire w_dff_A_vYxh0iqH1_0;
	wire w_dff_A_CKoeG2LA3_0;
	wire w_dff_A_Ajoa1CTr4_0;
	wire w_dff_A_0E6OY1vP3_0;
	wire w_dff_A_BSzPQ1cr8_0;
	wire w_dff_A_GODjdHIs6_0;
	wire w_dff_A_vsh7Yx6j7_0;
	wire w_dff_A_iLtnmXgW9_0;
	wire w_dff_A_tQSgV8Ht4_0;
	wire w_dff_A_aDglIXsz2_0;
	wire w_dff_A_tpByKxB19_0;
	wire w_dff_A_3mKSz1HS2_2;
	wire w_dff_A_Ayv7Ppx06_0;
	wire w_dff_A_VRZQs1TI6_0;
	wire w_dff_A_qsKJ5qbk2_0;
	wire w_dff_A_1HZKPwpJ8_0;
	wire w_dff_A_dYhEOeAy8_0;
	wire w_dff_A_RSd7YNyE2_0;
	wire w_dff_A_A9abrbx92_0;
	wire w_dff_A_Rf4Lq1LW1_0;
	wire w_dff_A_hjLywgXr8_0;
	wire w_dff_A_ww7T9sFt0_0;
	wire w_dff_A_rSdSHtaX5_0;
	wire w_dff_A_I55otHc79_0;
	wire w_dff_A_m6HZRIDq8_0;
	wire w_dff_A_0GsZJ3Mb8_0;
	wire w_dff_A_0pK4sGkm1_0;
	wire w_dff_A_hyf7lwvX0_0;
	wire w_dff_A_HvcpWl597_0;
	wire w_dff_A_rJki5nAi1_0;
	wire w_dff_A_9VJqhq2B5_0;
	wire w_dff_A_BdMtPa6c2_0;
	wire w_dff_A_NZQ6XDaE5_0;
	wire w_dff_A_JptcqQKJ8_0;
	wire w_dff_A_LqMDoJNm5_0;
	wire w_dff_A_q90xRDts9_0;
	wire w_dff_A_TpJpQaKf0_0;
	wire w_dff_A_orumTqvT2_0;
	wire w_dff_A_7xJ4e79C4_0;
	wire w_dff_A_5B6tToZH1_0;
	wire w_dff_A_qYJIAWMz3_0;
	wire w_dff_A_xHpIpZJQ9_0;
	wire w_dff_A_4qI47ELd3_0;
	wire w_dff_A_aEUSdggI8_0;
	wire w_dff_A_9MjpSZ2L5_0;
	wire w_dff_A_mJdFMrsI5_0;
	wire w_dff_A_GVM2uqUo8_0;
	wire w_dff_A_FCk9xpC88_0;
	wire w_dff_A_yVTWZZlE3_0;
	wire w_dff_A_BwnN4wyZ6_0;
	wire w_dff_A_zsLCgcyH6_0;
	wire w_dff_A_QJ9RmIWD8_0;
	wire w_dff_A_CnvvP1RT2_0;
	wire w_dff_A_lloiz32N1_0;
	wire w_dff_A_pmP8KUow4_0;
	wire w_dff_A_FPm68tqi3_0;
	wire w_dff_A_PuULeQOX4_0;
	wire w_dff_A_oVV6jfYC5_0;
	wire w_dff_A_F38qtnoU0_0;
	wire w_dff_A_QboQC8Am2_0;
	wire w_dff_A_nG0DJOaO2_0;
	wire w_dff_A_J4pwPtEZ7_0;
	wire w_dff_A_L3RBCFh35_0;
	wire w_dff_A_hIz7n9vM4_0;
	wire w_dff_A_AbiGTZzy0_0;
	wire w_dff_A_Qbl7wfZu4_0;
	wire w_dff_A_r6IAGJNV0_0;
	wire w_dff_A_5tez9fPY8_0;
	wire w_dff_A_4Rk2jIV46_0;
	wire w_dff_A_WKEXg25Z4_0;
	wire w_dff_A_VU38RyNS6_0;
	wire w_dff_A_EiwL64n56_0;
	wire w_dff_A_uhc33KPv8_0;
	wire w_dff_A_JwDn17xS7_0;
	wire w_dff_A_2U74uBbJ9_0;
	wire w_dff_A_rpX69VDC6_0;
	wire w_dff_A_E4GIdYLV5_0;
	wire w_dff_A_6WTvRgv09_0;
	wire w_dff_A_4Yw9ASMd9_0;
	wire w_dff_A_gzOCrBSk3_0;
	wire w_dff_A_6EzLwRpF3_0;
	wire w_dff_A_Jaj8X0jw9_0;
	wire w_dff_A_rwzbeZNn0_0;
	wire w_dff_A_b67luegq1_0;
	wire w_dff_A_MC6t3PqP5_0;
	wire w_dff_A_NqoWYY8r9_0;
	wire w_dff_A_MIjE16wO4_0;
	wire w_dff_A_P2YgcVvb8_0;
	wire w_dff_A_Tr8mwIHU2_0;
	wire w_dff_A_s2adAl7P4_2;
	wire w_dff_A_p9e74CQN8_0;
	wire w_dff_A_nPiZY0MH4_0;
	wire w_dff_A_dzEbedML5_0;
	wire w_dff_A_NOpDgdU14_0;
	wire w_dff_A_lXzMcDau3_0;
	wire w_dff_A_VYRVjvVu5_0;
	wire w_dff_A_xGtHPyAS5_0;
	wire w_dff_A_w1U5qlyc9_0;
	wire w_dff_A_E43w3Iwf1_0;
	wire w_dff_A_OqgKUni50_0;
	wire w_dff_A_aIvvBTVq1_0;
	wire w_dff_A_lodkKEjr8_0;
	wire w_dff_A_1oWgng8M0_0;
	wire w_dff_A_Mt25iuGA4_0;
	wire w_dff_A_uamHzhzN6_0;
	wire w_dff_A_3t3oRcwu8_0;
	wire w_dff_A_P9yYoLt63_0;
	wire w_dff_A_iuz09znQ0_0;
	wire w_dff_A_eMwdA4SH8_0;
	wire w_dff_A_axXOLZgR8_0;
	wire w_dff_A_9X9chWfX8_0;
	wire w_dff_A_DYOmGE027_0;
	wire w_dff_A_J8qY0DHt8_0;
	wire w_dff_A_3Lz4mhlJ9_0;
	wire w_dff_A_UMUx6kGP8_0;
	wire w_dff_A_mNB4LWA62_0;
	wire w_dff_A_0cpTtEaZ6_0;
	wire w_dff_A_VLKZEIgi1_0;
	wire w_dff_A_ftD70KiW2_0;
	wire w_dff_A_76xFgNlE8_0;
	wire w_dff_A_7okjH4Kb2_0;
	wire w_dff_A_fxSkxYUh1_0;
	wire w_dff_A_wST5657d5_0;
	wire w_dff_A_nBRekPHZ8_0;
	wire w_dff_A_mb2ngAR64_0;
	wire w_dff_A_5KIViX3l8_0;
	wire w_dff_A_AGWHZpDO6_0;
	wire w_dff_A_zMLwvWqH8_0;
	wire w_dff_A_qd6bs8PP5_0;
	wire w_dff_A_P2Ro2ra41_0;
	wire w_dff_A_2xv3eXLA9_0;
	wire w_dff_A_Mnry7XKU8_0;
	wire w_dff_A_Nxp6sLEB9_0;
	wire w_dff_A_2Ad0xBuh4_0;
	wire w_dff_A_PlYmFzEy7_0;
	wire w_dff_A_xgwGsZFZ7_0;
	wire w_dff_A_3yhwGmLo8_0;
	wire w_dff_A_Vz30GvIZ3_0;
	wire w_dff_A_7DQC3X7E3_0;
	wire w_dff_A_zb6EAGno7_0;
	wire w_dff_A_RPUJQJwf1_0;
	wire w_dff_A_Wfq44m7z6_0;
	wire w_dff_A_2P7uytly9_0;
	wire w_dff_A_XfE6Rlyr3_0;
	wire w_dff_A_xDalQPYM0_0;
	wire w_dff_A_OtFyS5E27_0;
	wire w_dff_A_pIqfvuvg1_0;
	wire w_dff_A_aTfSc5CN2_0;
	wire w_dff_A_unE3wgMZ3_0;
	wire w_dff_A_vs8e6brq8_0;
	wire w_dff_A_IoCGsAx39_0;
	wire w_dff_A_TPugt1ud5_0;
	wire w_dff_A_RoiPUm8A4_0;
	wire w_dff_A_wBzyuGAx4_0;
	wire w_dff_A_ZzMkZ7tJ5_0;
	wire w_dff_A_gi9R00dn4_0;
	wire w_dff_A_jT6H4wEd8_0;
	wire w_dff_A_c5sFRDUV9_0;
	wire w_dff_A_4QgCc8kE3_0;
	wire w_dff_A_maY7meEX3_0;
	wire w_dff_A_SmiJYLCg8_0;
	wire w_dff_A_WAI2As8U6_0;
	wire w_dff_A_cg1LW6JN5_0;
	wire w_dff_A_fLyeR8lw5_0;
	wire w_dff_A_msZXrXJB8_0;
	wire w_dff_A_1EaWz1YO0_0;
	wire w_dff_A_FVUuRbF61_2;
	wire w_dff_A_za6uKTJo8_0;
	wire w_dff_A_C1vBaGHQ0_0;
	wire w_dff_A_yy1oYe0Q9_0;
	wire w_dff_A_Ka45KprM5_0;
	wire w_dff_A_1v5LnPC65_0;
	wire w_dff_A_99xxFQsX7_0;
	wire w_dff_A_0V0sCq0t5_0;
	wire w_dff_A_xRnN0fqv0_0;
	wire w_dff_A_3w4Bxij31_0;
	wire w_dff_A_y8L2Rgy94_0;
	wire w_dff_A_bHjadYxX0_0;
	wire w_dff_A_vwBaucBK1_0;
	wire w_dff_A_hRggI1r32_0;
	wire w_dff_A_SpUHXYxh5_0;
	wire w_dff_A_OZDyMNbJ0_0;
	wire w_dff_A_hscaPDxD1_0;
	wire w_dff_A_oIPBw6n24_0;
	wire w_dff_A_ZrTDPSko0_0;
	wire w_dff_A_jISupvsL9_0;
	wire w_dff_A_Z6Wte2wt5_0;
	wire w_dff_A_DMbG3TAN0_0;
	wire w_dff_A_ty99He0M5_0;
	wire w_dff_A_FpQrcYFN9_0;
	wire w_dff_A_eTyRV7Uv1_0;
	wire w_dff_A_9tQgvxoD1_0;
	wire w_dff_A_uKFy8WHt6_0;
	wire w_dff_A_FaUFIllK8_0;
	wire w_dff_A_r3Jz7kyX5_0;
	wire w_dff_A_DPpqnHGu3_0;
	wire w_dff_A_sJ8FYyXE7_0;
	wire w_dff_A_fkBJLsLl2_0;
	wire w_dff_A_uInRUfya7_0;
	wire w_dff_A_AZHjDvnt3_0;
	wire w_dff_A_LFFSWndL4_0;
	wire w_dff_A_uwP9rW7q0_0;
	wire w_dff_A_iTMrYELx1_0;
	wire w_dff_A_dKru4FVS3_0;
	wire w_dff_A_gc6PomZM1_0;
	wire w_dff_A_wgS1mZES9_0;
	wire w_dff_A_A7ogKbe88_0;
	wire w_dff_A_GGEAhZFD1_0;
	wire w_dff_A_EMU3bqyG5_0;
	wire w_dff_A_sZdgB3DU9_0;
	wire w_dff_A_qh8CFvTP9_0;
	wire w_dff_A_Oa0Eoz0O7_0;
	wire w_dff_A_F4vtuYJg5_0;
	wire w_dff_A_C1QnvXea3_0;
	wire w_dff_A_Z0XmoKy22_0;
	wire w_dff_A_mLieapSf5_0;
	wire w_dff_A_wki21UKd6_0;
	wire w_dff_A_V2QxSvUa3_0;
	wire w_dff_A_3SMUQ99Y2_0;
	wire w_dff_A_NTZvkYIE1_0;
	wire w_dff_A_v6gqwMek3_0;
	wire w_dff_A_P5UemhMJ4_0;
	wire w_dff_A_rAzB2KhL6_0;
	wire w_dff_A_BXZ6q2DB4_0;
	wire w_dff_A_iMMJWG2L5_0;
	wire w_dff_A_zhj8ihkX4_0;
	wire w_dff_A_kZ7tR5Vs6_0;
	wire w_dff_A_J25sRFb05_0;
	wire w_dff_A_qTXuH1Rl1_0;
	wire w_dff_A_wJzBZD5p8_0;
	wire w_dff_A_o6BtxZ6k7_0;
	wire w_dff_A_DGm31C3J9_0;
	wire w_dff_A_XvQxqeEL5_0;
	wire w_dff_A_tyEDMw7H2_0;
	wire w_dff_A_lS2OuWMh8_0;
	wire w_dff_A_AiLT5bqw0_0;
	wire w_dff_A_oZeBMBU93_0;
	wire w_dff_A_RCoLPb1E4_0;
	wire w_dff_A_8aHZwmOH9_0;
	wire w_dff_A_6p1zyRIY9_0;
	wire w_dff_A_gEO0PD3S4_0;
	wire w_dff_A_t0EGDvpx4_0;
	wire w_dff_A_G7GNSuM17_2;
	wire w_dff_A_l1Vh7YgW6_0;
	wire w_dff_A_YRgofBZ27_0;
	wire w_dff_A_t781VRLc6_0;
	wire w_dff_A_OpGV8T1d9_0;
	wire w_dff_A_ZZI8jzxH0_0;
	wire w_dff_A_BTmzGfix2_0;
	wire w_dff_A_iMOunIXD4_0;
	wire w_dff_A_uZkFKS1K2_0;
	wire w_dff_A_7qGuwbAV7_0;
	wire w_dff_A_dVrQ63pj9_0;
	wire w_dff_A_EiR4OOmW4_0;
	wire w_dff_A_2wySulYn7_0;
	wire w_dff_A_FyJTiNBa6_0;
	wire w_dff_A_POP8tHOu1_0;
	wire w_dff_A_09a3uzDm5_0;
	wire w_dff_A_86xese044_0;
	wire w_dff_A_wvbbBwei4_0;
	wire w_dff_A_QaWOJcub3_0;
	wire w_dff_A_G7bYDsnd0_0;
	wire w_dff_A_ge6JoBjL4_0;
	wire w_dff_A_iXzRamAH7_0;
	wire w_dff_A_YWdabcHF9_0;
	wire w_dff_A_kZ4PPs6C3_0;
	wire w_dff_A_hjCbWuiG0_0;
	wire w_dff_A_zIAZchVZ0_0;
	wire w_dff_A_6k73NZF09_0;
	wire w_dff_A_u39syC7A8_0;
	wire w_dff_A_DLjQm3Yl1_0;
	wire w_dff_A_cghGQbgO7_0;
	wire w_dff_A_BSLORxXU8_0;
	wire w_dff_A_t89g5p5Z7_0;
	wire w_dff_A_jwDQdgv20_0;
	wire w_dff_A_SSNR797D2_0;
	wire w_dff_A_OdDu2nXl1_0;
	wire w_dff_A_xp0xzVgW6_0;
	wire w_dff_A_3UVpfIHH2_0;
	wire w_dff_A_eWAChmSl3_0;
	wire w_dff_A_B2x0OPTf8_0;
	wire w_dff_A_svCp7Kuf3_0;
	wire w_dff_A_3Y9U3X1j0_0;
	wire w_dff_A_BlOuYw4O7_0;
	wire w_dff_A_UiZeewtW8_0;
	wire w_dff_A_G9vZRCnT1_0;
	wire w_dff_A_pdE64WSt8_0;
	wire w_dff_A_a8wci0QL2_0;
	wire w_dff_A_HVtc20pM6_0;
	wire w_dff_A_HoqDBzTy0_0;
	wire w_dff_A_rvGeCKCp4_0;
	wire w_dff_A_5lX71WQ05_0;
	wire w_dff_A_lRr46IbB3_0;
	wire w_dff_A_D2B9kVQh6_0;
	wire w_dff_A_Ng1EtVUH7_0;
	wire w_dff_A_6TU938Al0_0;
	wire w_dff_A_cjivnYUC6_0;
	wire w_dff_A_ph7VmcbG0_0;
	wire w_dff_A_psBOdpLB2_0;
	wire w_dff_A_5wUvn2Aa6_0;
	wire w_dff_A_o5aCjrWi9_0;
	wire w_dff_A_yX64Na0j3_0;
	wire w_dff_A_ybwSwN4q5_0;
	wire w_dff_A_eqIXxdOv3_0;
	wire w_dff_A_EMdEozSn7_0;
	wire w_dff_A_EqCpjty86_0;
	wire w_dff_A_qJzw7aX38_0;
	wire w_dff_A_Ih6dXHZ23_0;
	wire w_dff_A_dWAEoDRf8_0;
	wire w_dff_A_ExzG3lhp8_0;
	wire w_dff_A_gmVidBMn2_0;
	wire w_dff_A_ge5HwoRn0_0;
	wire w_dff_A_2zNkM9dH8_0;
	wire w_dff_A_YJ1UD6012_0;
	wire w_dff_A_xg3ILKV69_0;
	wire w_dff_A_hekdlsy96_0;
	wire w_dff_A_ZkGIJPPY3_0;
	wire w_dff_A_J9A7hwTx6_2;
	wire w_dff_A_OT3GK1AG8_0;
	wire w_dff_A_z88WRpUP4_0;
	wire w_dff_A_6aCdpau06_0;
	wire w_dff_A_Z2SxVOMq0_0;
	wire w_dff_A_t9pJlqlj0_0;
	wire w_dff_A_mBrLKQAS5_0;
	wire w_dff_A_pPYqN8QY9_0;
	wire w_dff_A_nDxfWVzy4_0;
	wire w_dff_A_aKs1sSID5_0;
	wire w_dff_A_SaDtsbVW5_0;
	wire w_dff_A_rskkAhRw5_0;
	wire w_dff_A_d16tCrGm7_0;
	wire w_dff_A_RrPLuR4w6_0;
	wire w_dff_A_JPkdiDbF3_0;
	wire w_dff_A_CIZG3EZr5_0;
	wire w_dff_A_HrWvwZoa3_0;
	wire w_dff_A_T6keuIcK0_0;
	wire w_dff_A_byhhlgXr4_0;
	wire w_dff_A_HQtRgNkz1_0;
	wire w_dff_A_REKRK8Lc4_0;
	wire w_dff_A_mHslQZmo1_0;
	wire w_dff_A_LPYnCjel0_0;
	wire w_dff_A_aiC8ujeM9_0;
	wire w_dff_A_npbiUpmV7_0;
	wire w_dff_A_WLuGQe8X5_0;
	wire w_dff_A_ARD4GBYd6_0;
	wire w_dff_A_6vOwHz3W0_0;
	wire w_dff_A_1mVz9cx33_0;
	wire w_dff_A_CezH1A4P9_0;
	wire w_dff_A_WkD4XFm68_0;
	wire w_dff_A_egb0vbE24_0;
	wire w_dff_A_mUUSMgpW1_0;
	wire w_dff_A_tplcAAZk3_0;
	wire w_dff_A_cugwLUWM2_0;
	wire w_dff_A_gCBjj5To0_0;
	wire w_dff_A_jS5ZeMDw7_0;
	wire w_dff_A_Kc14vn7P7_0;
	wire w_dff_A_ieTvplCn3_0;
	wire w_dff_A_prZETgUx6_0;
	wire w_dff_A_CfTi23LL4_0;
	wire w_dff_A_W5YcOg6s9_0;
	wire w_dff_A_Y1xhP8IX0_0;
	wire w_dff_A_i1ZkUOO01_0;
	wire w_dff_A_ZpMOjCMn8_0;
	wire w_dff_A_pdcznA3U1_0;
	wire w_dff_A_90PSYUac0_0;
	wire w_dff_A_vYZoLNUU9_0;
	wire w_dff_A_clk9LFOM3_0;
	wire w_dff_A_SiZXybuQ0_0;
	wire w_dff_A_zX62wHPB0_0;
	wire w_dff_A_LDuhTvzO4_0;
	wire w_dff_A_utt3HlAP6_0;
	wire w_dff_A_0kol8nHv1_0;
	wire w_dff_A_1dTZoTcV6_0;
	wire w_dff_A_prsExu7H8_0;
	wire w_dff_A_qpW5m0wq7_0;
	wire w_dff_A_oLgD2FYp6_0;
	wire w_dff_A_tFvLmla28_0;
	wire w_dff_A_astKMbRC9_0;
	wire w_dff_A_DR0N3oYZ3_0;
	wire w_dff_A_6ervdhKj7_0;
	wire w_dff_A_YDBDD9XM0_0;
	wire w_dff_A_szJk4oae9_0;
	wire w_dff_A_dzOdhbct6_0;
	wire w_dff_A_Z9iGPVmW6_0;
	wire w_dff_A_WReiHmMH0_0;
	wire w_dff_A_1PpJj5r82_0;
	wire w_dff_A_H7MVETaQ9_0;
	wire w_dff_A_bfht0aHI1_0;
	wire w_dff_A_yDaHJsnz9_0;
	wire w_dff_A_pn6SeXyP7_0;
	wire w_dff_A_9SIcFGXG8_0;
	wire w_dff_A_PdGDE0w11_0;
	wire w_dff_A_VAnnSBRN8_2;
	wire w_dff_A_9dclbZFg8_0;
	wire w_dff_A_H1Vz3KZD4_0;
	wire w_dff_A_714oKhDN7_0;
	wire w_dff_A_Dbo2qgqC8_0;
	wire w_dff_A_knKqIHwR8_0;
	wire w_dff_A_HLs8llKn5_0;
	wire w_dff_A_wjyhKIaP9_0;
	wire w_dff_A_dlGzekG65_0;
	wire w_dff_A_44mmG9RV8_0;
	wire w_dff_A_4KtgLMUH1_0;
	wire w_dff_A_5Y1m7mUl0_0;
	wire w_dff_A_TrnfOlBA5_0;
	wire w_dff_A_9Q3mkgmn8_0;
	wire w_dff_A_TWfIS3Y48_0;
	wire w_dff_A_3OYjzytK3_0;
	wire w_dff_A_b28BH3sI6_0;
	wire w_dff_A_dfu5OI8d7_0;
	wire w_dff_A_FLLW9SZi4_0;
	wire w_dff_A_eurZLrOl5_0;
	wire w_dff_A_J4lRUlM41_0;
	wire w_dff_A_FH8Jbixz1_0;
	wire w_dff_A_AU04OJJb4_0;
	wire w_dff_A_z1Ip7aOA5_0;
	wire w_dff_A_3rq6zMSZ4_0;
	wire w_dff_A_1FgSU8u30_0;
	wire w_dff_A_nU5DdzsQ8_0;
	wire w_dff_A_jHgPgV3P6_0;
	wire w_dff_A_f78FGPY04_0;
	wire w_dff_A_xxjc11Jw2_0;
	wire w_dff_A_pHY3wEVz0_0;
	wire w_dff_A_woeJLyyP5_0;
	wire w_dff_A_shKRasrK3_0;
	wire w_dff_A_e4VjbQK76_0;
	wire w_dff_A_laEcLmxb5_0;
	wire w_dff_A_VnS7i1n47_0;
	wire w_dff_A_gYlyyBcP4_0;
	wire w_dff_A_gnzT7elK8_0;
	wire w_dff_A_KT063OkY9_0;
	wire w_dff_A_REvm0Ti38_0;
	wire w_dff_A_hEIdsQBR7_0;
	wire w_dff_A_lrxGnw5p6_0;
	wire w_dff_A_NksPVsVY1_0;
	wire w_dff_A_B0e1tjFT2_0;
	wire w_dff_A_wGAb6cgj5_0;
	wire w_dff_A_kOvwD4EN1_0;
	wire w_dff_A_xXh45aOw1_0;
	wire w_dff_A_F7myeWuA9_0;
	wire w_dff_A_NzAkOC3J2_0;
	wire w_dff_A_lHMY5O9U2_0;
	wire w_dff_A_WaprlTOm8_0;
	wire w_dff_A_Z9V70P7D1_0;
	wire w_dff_A_FoIMywaP6_0;
	wire w_dff_A_aUiQH5065_0;
	wire w_dff_A_UaEBNyVD6_0;
	wire w_dff_A_v8xBNfep9_0;
	wire w_dff_A_6TCBvEZt0_0;
	wire w_dff_A_UGYMim0V1_0;
	wire w_dff_A_2PjSqNPD0_0;
	wire w_dff_A_ELfXi9OM0_0;
	wire w_dff_A_ScjEGo8T7_0;
	wire w_dff_A_yLQPyHP65_0;
	wire w_dff_A_h5Z40Nx32_0;
	wire w_dff_A_e6FpgkT84_0;
	wire w_dff_A_271WHuu79_0;
	wire w_dff_A_hZJlLi9b2_0;
	wire w_dff_A_gr1AarT87_0;
	wire w_dff_A_ZsrDp5Hb4_0;
	wire w_dff_A_r7TiYwRb5_0;
	wire w_dff_A_wQc4N6F10_0;
	wire w_dff_A_w0TpfyKX6_0;
	wire w_dff_A_i00tNIAk7_0;
	wire w_dff_A_ayUQ4M2B4_0;
	wire w_dff_A_w2HyVyOp2_2;
	wire w_dff_A_dEgH3gZa5_0;
	wire w_dff_A_e3EN56Ug9_0;
	wire w_dff_A_MGsqM0QD9_0;
	wire w_dff_A_424vlOw97_0;
	wire w_dff_A_vqFXGeDc9_0;
	wire w_dff_A_fxeMHGBj1_0;
	wire w_dff_A_5eCmOOrO8_0;
	wire w_dff_A_fCnjqpdM9_0;
	wire w_dff_A_SP5xCAOO3_0;
	wire w_dff_A_nOCCSmuC9_0;
	wire w_dff_A_4y19yrRB2_0;
	wire w_dff_A_cn1xMRgu8_0;
	wire w_dff_A_lHLZynKs6_0;
	wire w_dff_A_FBWUylAB6_0;
	wire w_dff_A_hlnueaBz6_0;
	wire w_dff_A_fC7LxQrg5_0;
	wire w_dff_A_pbo0JmI97_0;
	wire w_dff_A_WtUhihMP7_0;
	wire w_dff_A_5IlrSkiZ1_0;
	wire w_dff_A_eOyP6tTM9_0;
	wire w_dff_A_wIKtdQ1K0_0;
	wire w_dff_A_cnW6YU3B0_0;
	wire w_dff_A_DNneq2c38_0;
	wire w_dff_A_vTKNXfgK2_0;
	wire w_dff_A_ETAzq8d28_0;
	wire w_dff_A_wRj2UmGg4_0;
	wire w_dff_A_TezxDVX47_0;
	wire w_dff_A_CiubDuNg1_0;
	wire w_dff_A_6839GalW5_0;
	wire w_dff_A_JZiKi63P2_0;
	wire w_dff_A_UmeOw9qz5_0;
	wire w_dff_A_om6LMqsY6_0;
	wire w_dff_A_pnKXDrFZ2_0;
	wire w_dff_A_EkvWhy9c1_0;
	wire w_dff_A_McuKVLE19_0;
	wire w_dff_A_O2c9yV886_0;
	wire w_dff_A_vmS1Tf6j7_0;
	wire w_dff_A_BcQnvUUK0_0;
	wire w_dff_A_XxhYinKL9_0;
	wire w_dff_A_jmScHiG65_0;
	wire w_dff_A_6HrDtJvH1_0;
	wire w_dff_A_EeofwH1E4_0;
	wire w_dff_A_qMNdxDAx8_0;
	wire w_dff_A_sRnl4iWS2_0;
	wire w_dff_A_Gov2DavA1_0;
	wire w_dff_A_1x2YLxUC5_0;
	wire w_dff_A_qHqQcl8L5_0;
	wire w_dff_A_AaPLH0O98_0;
	wire w_dff_A_zDreKGMw3_0;
	wire w_dff_A_1B5uHCIJ5_0;
	wire w_dff_A_obB3jffj7_0;
	wire w_dff_A_2inXgvHr5_0;
	wire w_dff_A_zMQsW4rp5_0;
	wire w_dff_A_kDzuObk15_0;
	wire w_dff_A_gM8rTyx33_0;
	wire w_dff_A_3KhK7FKk4_0;
	wire w_dff_A_YHo9eLPz9_0;
	wire w_dff_A_B3mL47Ol0_0;
	wire w_dff_A_UIose7X75_0;
	wire w_dff_A_6knHOhdi5_0;
	wire w_dff_A_ujgxaduW8_0;
	wire w_dff_A_zdrczSWU2_0;
	wire w_dff_A_nEf6vn7y6_0;
	wire w_dff_A_XuxYCQog7_0;
	wire w_dff_A_lT651o3w4_0;
	wire w_dff_A_mTAZ184J2_0;
	wire w_dff_A_NzAA6erK0_0;
	wire w_dff_A_CI7tv4nR2_0;
	wire w_dff_A_Q2dUOvdm8_0;
	wire w_dff_A_QUCKT1qY1_0;
	wire w_dff_A_XfBcr8Xc9_0;
	wire w_dff_A_0ifBWpOE0_2;
	wire w_dff_A_Rmu6IeBp3_0;
	wire w_dff_A_c13PA3Mc0_0;
	wire w_dff_A_ayPpK3iw9_0;
	wire w_dff_A_zVD5pPD83_0;
	wire w_dff_A_qhCPedcf8_0;
	wire w_dff_A_5mdW9eA25_0;
	wire w_dff_A_dL6WfK9L7_0;
	wire w_dff_A_SpbtbmWe6_0;
	wire w_dff_A_hbuPn93z3_0;
	wire w_dff_A_PMldSt8j0_0;
	wire w_dff_A_0xgDCn5z7_0;
	wire w_dff_A_c9ANKgon7_0;
	wire w_dff_A_DzYvff6t7_0;
	wire w_dff_A_dLsKJYNz0_0;
	wire w_dff_A_546VhKMd2_0;
	wire w_dff_A_2fvITQwY3_0;
	wire w_dff_A_VM0zCInD4_0;
	wire w_dff_A_qRs64vNu7_0;
	wire w_dff_A_tLRrioN56_0;
	wire w_dff_A_oLi9KfmR3_0;
	wire w_dff_A_qOumC5p46_0;
	wire w_dff_A_zc5VxotV5_0;
	wire w_dff_A_t6hlBMUT9_0;
	wire w_dff_A_4lpClHmY8_0;
	wire w_dff_A_GDcdsuGN7_0;
	wire w_dff_A_CnGQY7IH6_0;
	wire w_dff_A_IEP2ywln1_0;
	wire w_dff_A_HVl97lFC3_0;
	wire w_dff_A_9pPqOvsr4_0;
	wire w_dff_A_Ds1Iroqm5_0;
	wire w_dff_A_a4mejR9R5_0;
	wire w_dff_A_Lw9Wm6ZG2_0;
	wire w_dff_A_Qji9yAsW6_0;
	wire w_dff_A_kE8lqlHy4_0;
	wire w_dff_A_xTIwdaok7_0;
	wire w_dff_A_xLxeiD2W4_0;
	wire w_dff_A_NpK5X4pA4_0;
	wire w_dff_A_wrZW0Lw43_0;
	wire w_dff_A_iOxkUXdF8_0;
	wire w_dff_A_NSdiEKXq9_0;
	wire w_dff_A_F632qRFm3_0;
	wire w_dff_A_5oZFBbjY8_0;
	wire w_dff_A_a2vEkte32_0;
	wire w_dff_A_N7jT3wYM6_0;
	wire w_dff_A_aleX8rro6_0;
	wire w_dff_A_MsPL2tlL5_0;
	wire w_dff_A_YJjFLiKR5_0;
	wire w_dff_A_wKeEnhlP8_0;
	wire w_dff_A_5hmPO68u9_0;
	wire w_dff_A_URqIKR3N9_0;
	wire w_dff_A_b9MSUZHG0_0;
	wire w_dff_A_llSMmZCC9_0;
	wire w_dff_A_ViMwEsyT2_0;
	wire w_dff_A_6DwsPHkN2_0;
	wire w_dff_A_qjpDKxOh4_0;
	wire w_dff_A_h17dLYDX7_0;
	wire w_dff_A_qOY04Bby5_0;
	wire w_dff_A_KPm0xNmJ3_0;
	wire w_dff_A_ImRMMbb36_0;
	wire w_dff_A_l1gWUlAh7_0;
	wire w_dff_A_fJAhGCsV8_0;
	wire w_dff_A_GOtZUZXK5_0;
	wire w_dff_A_hZuXznYA9_0;
	wire w_dff_A_sL6QDJKH0_0;
	wire w_dff_A_DtTSog067_0;
	wire w_dff_A_tbGC8tld8_0;
	wire w_dff_A_64JxdCda3_0;
	wire w_dff_A_WeCI0N5o2_0;
	wire w_dff_A_mJuGf5gD4_0;
	wire w_dff_A_IvTJn8Y02_0;
	wire w_dff_A_INrlTL4v6_2;
	wire w_dff_A_dzJBt3XK3_0;
	wire w_dff_A_Vr2TkBZ93_0;
	wire w_dff_A_Flr0wM298_0;
	wire w_dff_A_Kc2qisMs5_0;
	wire w_dff_A_E2dKC4Xb7_0;
	wire w_dff_A_n5ZDpFvC7_0;
	wire w_dff_A_2R71b5u67_0;
	wire w_dff_A_Oqrq1htL2_0;
	wire w_dff_A_sHi9szqV5_0;
	wire w_dff_A_YAPjvI9S1_0;
	wire w_dff_A_nQ6HQWd80_0;
	wire w_dff_A_iXgVBlFM2_0;
	wire w_dff_A_444c1OEZ5_0;
	wire w_dff_A_JLHjEdjq5_0;
	wire w_dff_A_MUAHkjCu1_0;
	wire w_dff_A_7XJAZRSW1_0;
	wire w_dff_A_5Je0kVlb2_0;
	wire w_dff_A_UY1BCc0f6_0;
	wire w_dff_A_eQQGW6GA3_0;
	wire w_dff_A_ZxoQJk0A0_0;
	wire w_dff_A_p3P2CgPH2_0;
	wire w_dff_A_IUk9R3nt1_0;
	wire w_dff_A_Zna0LaSe0_0;
	wire w_dff_A_Y59SHbD43_0;
	wire w_dff_A_lpdVdwYS8_0;
	wire w_dff_A_wDZmmeic0_0;
	wire w_dff_A_C0U5MoLj7_0;
	wire w_dff_A_gNRhiPIO4_0;
	wire w_dff_A_lRndsGCf1_0;
	wire w_dff_A_FchBVqcv4_0;
	wire w_dff_A_xRP8DBtF8_0;
	wire w_dff_A_ySjBwn3y9_0;
	wire w_dff_A_hlCxXxgl1_0;
	wire w_dff_A_TYLYzYKD6_0;
	wire w_dff_A_YZ6lbGs56_0;
	wire w_dff_A_N3zUviHw5_0;
	wire w_dff_A_pTv2ymDG2_0;
	wire w_dff_A_265Slivm5_0;
	wire w_dff_A_YhOHnR7d2_0;
	wire w_dff_A_kPPJ7LfZ7_0;
	wire w_dff_A_bJQdLUD66_0;
	wire w_dff_A_fUKoKbHh6_0;
	wire w_dff_A_jVbtG9B81_0;
	wire w_dff_A_a3rkbpN66_0;
	wire w_dff_A_HV3QeVWQ7_0;
	wire w_dff_A_msFJJVRT6_0;
	wire w_dff_A_duC2MSQt9_0;
	wire w_dff_A_9fyzrEba9_0;
	wire w_dff_A_WfR8fa7O6_0;
	wire w_dff_A_SO0ETjHd5_0;
	wire w_dff_A_GpAnB8xc4_0;
	wire w_dff_A_oGlMQOfk5_0;
	wire w_dff_A_apJ3dJcE4_0;
	wire w_dff_A_170vd5ct5_0;
	wire w_dff_A_Tvp8A8RG7_0;
	wire w_dff_A_8Mxb0QGd8_0;
	wire w_dff_A_OFto8a2a2_0;
	wire w_dff_A_925AHoRn1_0;
	wire w_dff_A_rS0iKfSZ9_0;
	wire w_dff_A_OUfcnEjW0_0;
	wire w_dff_A_ldx1rHEh9_0;
	wire w_dff_A_PZgLZaZI0_0;
	wire w_dff_A_CInfOAQj1_0;
	wire w_dff_A_yTNymAn70_0;
	wire w_dff_A_RzedOrNj5_0;
	wire w_dff_A_GEHMCHoa3_0;
	wire w_dff_A_ddrCs4lg1_0;
	wire w_dff_A_vNi7B1Gi5_0;
	wire w_dff_A_t1ePrhYd1_0;
	wire w_dff_A_IAZs4o3E0_2;
	wire w_dff_A_ItinrNbG6_0;
	wire w_dff_A_4Abqw0o03_0;
	wire w_dff_A_RO8TXVEV8_0;
	wire w_dff_A_b4iNdPyV0_0;
	wire w_dff_A_RQdxJYaD5_0;
	wire w_dff_A_gbjOaIdn4_0;
	wire w_dff_A_64MVXsYw9_0;
	wire w_dff_A_pgHrHjs61_0;
	wire w_dff_A_bOH4RhaY2_0;
	wire w_dff_A_LBoqBJPW2_0;
	wire w_dff_A_2BYgK6QY3_0;
	wire w_dff_A_QFF96nlz6_0;
	wire w_dff_A_4H0prr0p5_0;
	wire w_dff_A_q6uyiPbh9_0;
	wire w_dff_A_g0egDFDs4_0;
	wire w_dff_A_j0XC9rSh5_0;
	wire w_dff_A_2l2u3Yf81_0;
	wire w_dff_A_oOWWJo2F3_0;
	wire w_dff_A_plnOhLod1_0;
	wire w_dff_A_oOP4xdlA8_0;
	wire w_dff_A_kjq3835h5_0;
	wire w_dff_A_Ggb9Bo7a0_0;
	wire w_dff_A_SfBCPdp25_0;
	wire w_dff_A_de5F7q3x7_0;
	wire w_dff_A_YquGHsyh8_0;
	wire w_dff_A_woFHH4tr9_0;
	wire w_dff_A_oyGr7D3X5_0;
	wire w_dff_A_Ckd77GBL9_0;
	wire w_dff_A_otg2TxFE9_0;
	wire w_dff_A_1YtZ9VoF9_0;
	wire w_dff_A_UFa0VRPK7_0;
	wire w_dff_A_y2Cpwbtj9_0;
	wire w_dff_A_z2CMdxhl6_0;
	wire w_dff_A_dsoI6mN01_0;
	wire w_dff_A_SXfYOpZi7_0;
	wire w_dff_A_VbfBQ0OQ0_0;
	wire w_dff_A_Hpj35L0u4_0;
	wire w_dff_A_pZrId7J13_0;
	wire w_dff_A_swZSLd5s3_0;
	wire w_dff_A_APbaCdFl8_0;
	wire w_dff_A_jq9MgPEF3_0;
	wire w_dff_A_bjLtbmY60_0;
	wire w_dff_A_JBBcEA4Z7_0;
	wire w_dff_A_a7ZLB98X2_0;
	wire w_dff_A_iJJYMslN2_0;
	wire w_dff_A_o1BmuXI45_0;
	wire w_dff_A_qtGxJDtF0_0;
	wire w_dff_A_7dFCxesR8_0;
	wire w_dff_A_ZY7bDPDY5_0;
	wire w_dff_A_CglyVY7S2_0;
	wire w_dff_A_OUuJVZMo4_0;
	wire w_dff_A_KeMazQGi9_0;
	wire w_dff_A_SCOSbgDQ3_0;
	wire w_dff_A_0whYsXA34_0;
	wire w_dff_A_Wj0ClU7E4_0;
	wire w_dff_A_2GVeQnEa6_0;
	wire w_dff_A_Usl54Erk1_0;
	wire w_dff_A_1wMbp6Lr0_0;
	wire w_dff_A_2UqSuI3a2_0;
	wire w_dff_A_8AN3YywG6_0;
	wire w_dff_A_Qj5uX7bo9_0;
	wire w_dff_A_zhklAO6a8_0;
	wire w_dff_A_Ld80DM2H1_0;
	wire w_dff_A_68qUDKBA9_0;
	wire w_dff_A_J5JLUTcn0_0;
	wire w_dff_A_D3oyc61M9_0;
	wire w_dff_A_MeCNDPEa6_0;
	wire w_dff_A_dFfcmXB78_0;
	wire w_dff_A_bZXjmX1T8_2;
	wire w_dff_A_J0OfzNGE4_0;
	wire w_dff_A_YxbWi1fC4_0;
	wire w_dff_A_ijb0lVcg0_0;
	wire w_dff_A_pAz3CRnI9_0;
	wire w_dff_A_RJoTSTKc7_0;
	wire w_dff_A_ojppQPfy7_0;
	wire w_dff_A_whTb4Wka5_0;
	wire w_dff_A_auNV7sAo0_0;
	wire w_dff_A_kEL4YbMu6_0;
	wire w_dff_A_rblVoy0h1_0;
	wire w_dff_A_9LhXojvx8_0;
	wire w_dff_A_iCOWJdkT5_0;
	wire w_dff_A_jJ5Qlu4Y8_0;
	wire w_dff_A_wuSrx01o9_0;
	wire w_dff_A_PmWPTiZU2_0;
	wire w_dff_A_BxlJGkPT7_0;
	wire w_dff_A_yZvDAxEX4_0;
	wire w_dff_A_bPdAc6T62_0;
	wire w_dff_A_eHi8f8rP6_0;
	wire w_dff_A_KaaP93St6_0;
	wire w_dff_A_rEQf91VJ5_0;
	wire w_dff_A_YAN38V8C2_0;
	wire w_dff_A_cZOdT8la7_0;
	wire w_dff_A_ekVHlDMz7_0;
	wire w_dff_A_gOBp3VlD1_0;
	wire w_dff_A_EIOPK32F7_0;
	wire w_dff_A_wsehX8vH1_0;
	wire w_dff_A_EXdmOgX76_0;
	wire w_dff_A_pD8UYqFN8_0;
	wire w_dff_A_5HkGXnDh4_0;
	wire w_dff_A_6mbR5O7N0_0;
	wire w_dff_A_k0MGrKmU1_0;
	wire w_dff_A_jEGbxiky3_0;
	wire w_dff_A_tYzpPAIH3_0;
	wire w_dff_A_wnoqg8Av2_0;
	wire w_dff_A_Q8slLJEZ5_0;
	wire w_dff_A_alHIAczq5_0;
	wire w_dff_A_GF0mvWa02_0;
	wire w_dff_A_f9u2wKKo3_0;
	wire w_dff_A_a6ZncgSM3_0;
	wire w_dff_A_vMU3Xfbq8_0;
	wire w_dff_A_0qqEFaxx2_0;
	wire w_dff_A_jsaQSO5d6_0;
	wire w_dff_A_DLeea00d6_0;
	wire w_dff_A_fsUUoAD81_0;
	wire w_dff_A_AFyNESGA8_0;
	wire w_dff_A_Hrp0jJln5_0;
	wire w_dff_A_M8Sx6SPF5_0;
	wire w_dff_A_P0sRalXm7_0;
	wire w_dff_A_5CAqbjeG2_0;
	wire w_dff_A_se3ZFNKb6_0;
	wire w_dff_A_93317jFh2_0;
	wire w_dff_A_D3bY47Lm8_0;
	wire w_dff_A_ezXm4KjA9_0;
	wire w_dff_A_mgudidAW3_0;
	wire w_dff_A_RXtlG59c6_0;
	wire w_dff_A_RsBttq8o1_0;
	wire w_dff_A_IFH0cgii4_0;
	wire w_dff_A_WqwQnJIn4_0;
	wire w_dff_A_EMUHb9yI1_0;
	wire w_dff_A_OaT702BY1_0;
	wire w_dff_A_MPEtOBkU2_0;
	wire w_dff_A_obS70QOw1_0;
	wire w_dff_A_mJo0oCdy0_0;
	wire w_dff_A_LXYObhyu6_0;
	wire w_dff_A_IA2TyC683_0;
	wire w_dff_A_eCTgGWm33_0;
	wire w_dff_A_73F8XiAD0_2;
	wire w_dff_A_iPKVGkco1_0;
	wire w_dff_A_6nfmMa9U8_0;
	wire w_dff_A_rLBPzbBR9_0;
	wire w_dff_A_rtDu19XC0_0;
	wire w_dff_A_XfQEC6OM4_0;
	wire w_dff_A_CB6r4lDG5_0;
	wire w_dff_A_f9s9udqi9_0;
	wire w_dff_A_0vRYqZP50_0;
	wire w_dff_A_vVkDP0P28_0;
	wire w_dff_A_61KF65Qe4_0;
	wire w_dff_A_6F1CRKmN5_0;
	wire w_dff_A_LhGzkaqS7_0;
	wire w_dff_A_P9jAgzKT0_0;
	wire w_dff_A_SWzMbmyQ7_0;
	wire w_dff_A_d1FGqUiP2_0;
	wire w_dff_A_gPVPJXCs1_0;
	wire w_dff_A_w1hs2DSQ8_0;
	wire w_dff_A_TjBlvOuY0_0;
	wire w_dff_A_HXYImnU18_0;
	wire w_dff_A_XpaLSiGt5_0;
	wire w_dff_A_PUf5IYiC5_0;
	wire w_dff_A_Mer49gxn2_0;
	wire w_dff_A_qi5lk1194_0;
	wire w_dff_A_zSOTXPk00_0;
	wire w_dff_A_w7WMnjLN2_0;
	wire w_dff_A_adGmR87B9_0;
	wire w_dff_A_KZBXlJhR1_0;
	wire w_dff_A_jjFgBrHF1_0;
	wire w_dff_A_2V4vMHZg3_0;
	wire w_dff_A_4NmUx1zy8_0;
	wire w_dff_A_f3UNqLF68_0;
	wire w_dff_A_1TkdnhK27_0;
	wire w_dff_A_7mtasAMM5_0;
	wire w_dff_A_vuUWrtzl7_0;
	wire w_dff_A_hvqVntsB3_0;
	wire w_dff_A_xn4A3gjX9_0;
	wire w_dff_A_LGA0xfO45_0;
	wire w_dff_A_xl2lWlZv4_0;
	wire w_dff_A_RyB0ER9j9_0;
	wire w_dff_A_GmkmoVbC6_0;
	wire w_dff_A_Lo3cqPBt5_0;
	wire w_dff_A_lUViqljC5_0;
	wire w_dff_A_ToIZSpra2_0;
	wire w_dff_A_xgU7Kr8u0_0;
	wire w_dff_A_ma8E5OHg5_0;
	wire w_dff_A_ga3vZeMV5_0;
	wire w_dff_A_or1Aq6e42_0;
	wire w_dff_A_96S3lsn00_0;
	wire w_dff_A_FVslTOr77_0;
	wire w_dff_A_xtPfsbII4_0;
	wire w_dff_A_b5iJ6r5u9_0;
	wire w_dff_A_BaUTZo9B0_0;
	wire w_dff_A_hy3GACAm2_0;
	wire w_dff_A_qsYpd8yx8_0;
	wire w_dff_A_lfpFRE3U9_0;
	wire w_dff_A_y67T9QrJ9_0;
	wire w_dff_A_iTEsgKpP0_0;
	wire w_dff_A_aNKI4mui0_0;
	wire w_dff_A_3z6DXO5Y2_0;
	wire w_dff_A_8S6W1afs5_0;
	wire w_dff_A_InSWDsT87_0;
	wire w_dff_A_Gw5uphno0_0;
	wire w_dff_A_3eXJ7f2T9_0;
	wire w_dff_A_CcjBL7KS9_0;
	wire w_dff_A_PQ2jiEph5_0;
	wire w_dff_A_4laSHGJN4_0;
	wire w_dff_A_cbJx3cUU7_2;
	wire w_dff_A_kN1bSLPi0_0;
	wire w_dff_A_pU53Tzbz8_0;
	wire w_dff_A_fHXVlomx4_0;
	wire w_dff_A_9lMNg9097_0;
	wire w_dff_A_r5qrXXzZ8_0;
	wire w_dff_A_NNhvWYBd5_0;
	wire w_dff_A_BW8ScAn92_0;
	wire w_dff_A_H7YuW3Io4_0;
	wire w_dff_A_jyqamt6N6_0;
	wire w_dff_A_CklLsOyq2_0;
	wire w_dff_A_6CPpkvLh9_0;
	wire w_dff_A_Wm95GZbe9_0;
	wire w_dff_A_OrJ1VE671_0;
	wire w_dff_A_O0jiO9VO5_0;
	wire w_dff_A_vDd1nOyy4_0;
	wire w_dff_A_mhtgDgWK5_0;
	wire w_dff_A_rPLaUmXr4_0;
	wire w_dff_A_Agwmk0Xn6_0;
	wire w_dff_A_YFC8JQ6b7_0;
	wire w_dff_A_ihtAkP0y8_0;
	wire w_dff_A_5BBIUexo6_0;
	wire w_dff_A_zKqflDUK0_0;
	wire w_dff_A_D3kO9vDW6_0;
	wire w_dff_A_MDB4X0DZ7_0;
	wire w_dff_A_VKvh9Ose0_0;
	wire w_dff_A_s4cSdd4I1_0;
	wire w_dff_A_nm3nGpql9_0;
	wire w_dff_A_i93jo2NR1_0;
	wire w_dff_A_fM9oUSDX1_0;
	wire w_dff_A_YzMm3uIC9_0;
	wire w_dff_A_JXKbEr9G1_0;
	wire w_dff_A_pSJFC5g39_0;
	wire w_dff_A_D1zuIqrG5_0;
	wire w_dff_A_xL28KK234_0;
	wire w_dff_A_lvTNrHnY2_0;
	wire w_dff_A_e1D8fWgY0_0;
	wire w_dff_A_3ac4XeuC1_0;
	wire w_dff_A_bKSR799b3_0;
	wire w_dff_A_PkaK4fsu9_0;
	wire w_dff_A_CD6IEukq8_0;
	wire w_dff_A_IHOJ7yki6_0;
	wire w_dff_A_vMFXKzEU7_0;
	wire w_dff_A_HPDvgGPZ5_0;
	wire w_dff_A_NE76jVWk7_0;
	wire w_dff_A_huvqzPo59_0;
	wire w_dff_A_WYyDuJiZ8_0;
	wire w_dff_A_9SEdrZrT9_0;
	wire w_dff_A_zUuFTNIx7_0;
	wire w_dff_A_IvIvHytR2_0;
	wire w_dff_A_dqathm1m8_0;
	wire w_dff_A_hKuATZ0h5_0;
	wire w_dff_A_TbdAxbTg1_0;
	wire w_dff_A_UafSs2yk8_0;
	wire w_dff_A_xejBHwc88_0;
	wire w_dff_A_npyi6nsg2_0;
	wire w_dff_A_6HR8vrRl8_0;
	wire w_dff_A_ObTwPOA53_0;
	wire w_dff_A_Gd7G0SPF3_0;
	wire w_dff_A_p921a5Ff0_0;
	wire w_dff_A_FWzLRRfM1_0;
	wire w_dff_A_7iw3XPmD2_0;
	wire w_dff_A_nMFdD3i91_0;
	wire w_dff_A_KoRukcaO3_0;
	wire w_dff_A_78UlX4T87_0;
	wire w_dff_A_XAZwDoNk6_0;
	wire w_dff_A_9pd4SMnz2_2;
	wire w_dff_A_9PfmIkxi1_0;
	wire w_dff_A_gnBGN4Av4_0;
	wire w_dff_A_tnAvPrj45_0;
	wire w_dff_A_6frgHy4c3_0;
	wire w_dff_A_UC3MrkNQ4_0;
	wire w_dff_A_jwBoS0RU2_0;
	wire w_dff_A_DAUUFlDO5_0;
	wire w_dff_A_D7LneTQU1_0;
	wire w_dff_A_GZv5SRhw9_0;
	wire w_dff_A_5ONaDWk54_0;
	wire w_dff_A_y8c5hkjk6_0;
	wire w_dff_A_DRixAHwj6_0;
	wire w_dff_A_WmqDGt3E9_0;
	wire w_dff_A_kjyaosTa3_0;
	wire w_dff_A_FLcztQVR8_0;
	wire w_dff_A_o7EYSRrV1_0;
	wire w_dff_A_k0BcLd351_0;
	wire w_dff_A_vAsdVf9t2_0;
	wire w_dff_A_Wpxldu1u5_0;
	wire w_dff_A_DsxfHCAe8_0;
	wire w_dff_A_A0VIBD6f3_0;
	wire w_dff_A_D9LoGEHc7_0;
	wire w_dff_A_3QJY9zSq4_0;
	wire w_dff_A_SHrOD7al1_0;
	wire w_dff_A_KSJ6qf754_0;
	wire w_dff_A_9R7PCgSB1_0;
	wire w_dff_A_cNqTuilG0_0;
	wire w_dff_A_ueFnkmeT1_0;
	wire w_dff_A_ItioFyrS9_0;
	wire w_dff_A_ef6IySI54_0;
	wire w_dff_A_S5c0VLsR1_0;
	wire w_dff_A_rkSGiJT10_0;
	wire w_dff_A_Rk3Hp52T3_0;
	wire w_dff_A_GU2CYuYu2_0;
	wire w_dff_A_pxNQ3lJG6_0;
	wire w_dff_A_ACfNOD8U5_0;
	wire w_dff_A_BP3jpmuq8_0;
	wire w_dff_A_o197X08U4_0;
	wire w_dff_A_IRKI83st1_0;
	wire w_dff_A_6FcKrCVq1_0;
	wire w_dff_A_hyPT4sqK1_0;
	wire w_dff_A_J4PWYUh44_0;
	wire w_dff_A_QMvEQTq83_0;
	wire w_dff_A_3B312j3m4_0;
	wire w_dff_A_ML8REE182_0;
	wire w_dff_A_JNRb510u1_0;
	wire w_dff_A_ffVbLAbd2_0;
	wire w_dff_A_1c3odY0u9_0;
	wire w_dff_A_OS0Gssdy5_0;
	wire w_dff_A_zAO9MmO81_0;
	wire w_dff_A_pRkvoXdJ9_0;
	wire w_dff_A_Ft8LhTns2_0;
	wire w_dff_A_oytcSXHT7_0;
	wire w_dff_A_mTsLmeyk1_0;
	wire w_dff_A_IeRSX9aG3_0;
	wire w_dff_A_flvMSnwk1_0;
	wire w_dff_A_4o8JhBtq6_0;
	wire w_dff_A_RLhGQEcn3_0;
	wire w_dff_A_00lUY1g44_0;
	wire w_dff_A_RAQDISZA9_0;
	wire w_dff_A_dyfR1rfK6_0;
	wire w_dff_A_mLvQVxo51_0;
	wire w_dff_A_DvKJ7lzu8_0;
	wire w_dff_A_F60rCu3e1_0;
	wire w_dff_A_was1nG0s4_2;
	wire w_dff_A_4FCaNSnF5_0;
	wire w_dff_A_sYQ3v8rF5_0;
	wire w_dff_A_qcCGrghB4_0;
	wire w_dff_A_vqWtrOhV2_0;
	wire w_dff_A_GaEtTw5l1_0;
	wire w_dff_A_nmfPLLqq2_0;
	wire w_dff_A_x4vz5G3h7_0;
	wire w_dff_A_XBV70oQG5_0;
	wire w_dff_A_swgCIWAw8_0;
	wire w_dff_A_mqJpZsjQ7_0;
	wire w_dff_A_aqiF1x5N2_0;
	wire w_dff_A_WyWQDoRG2_0;
	wire w_dff_A_lclP3gQt2_0;
	wire w_dff_A_K44fYD4X4_0;
	wire w_dff_A_9NVRQDrT2_0;
	wire w_dff_A_6eKjYWIg9_0;
	wire w_dff_A_fRvKaxiS3_0;
	wire w_dff_A_z7fDSSEg3_0;
	wire w_dff_A_02JCHMu74_0;
	wire w_dff_A_BZFTdOfS3_0;
	wire w_dff_A_cAvlbuaf4_0;
	wire w_dff_A_IzU5Us0H6_0;
	wire w_dff_A_ImNjsGOR8_0;
	wire w_dff_A_N7K6viDq1_0;
	wire w_dff_A_zNqy6v5z2_0;
	wire w_dff_A_cpJQcQWt8_0;
	wire w_dff_A_qtfGvc608_0;
	wire w_dff_A_Tsx8jgau7_0;
	wire w_dff_A_edBHmIUS6_0;
	wire w_dff_A_BmyhuMAs1_0;
	wire w_dff_A_Vq2RT1fi4_0;
	wire w_dff_A_7yvtcHVA1_0;
	wire w_dff_A_VIOSofcj5_0;
	wire w_dff_A_SWBjya4A5_0;
	wire w_dff_A_dwoItiIv1_0;
	wire w_dff_A_VnNfcXQ54_0;
	wire w_dff_A_mgEdXRmX7_0;
	wire w_dff_A_XMGpYcXb6_0;
	wire w_dff_A_eVRl7QfR7_0;
	wire w_dff_A_lz2spGC57_0;
	wire w_dff_A_Y7GSdF3e7_0;
	wire w_dff_A_7A8A5mft1_0;
	wire w_dff_A_P69w1Sok6_0;
	wire w_dff_A_Yio3Fn8R3_0;
	wire w_dff_A_cy6FQlo22_0;
	wire w_dff_A_ZMOegiTE0_0;
	wire w_dff_A_r8X4Wh9u7_0;
	wire w_dff_A_AZVzxgdu0_0;
	wire w_dff_A_2ummRGDO3_0;
	wire w_dff_A_umWVonQZ5_0;
	wire w_dff_A_bXrxUx4F1_0;
	wire w_dff_A_qP4DiCFE7_0;
	wire w_dff_A_rXVWxa8g6_0;
	wire w_dff_A_jSx6AQGo9_0;
	wire w_dff_A_4riuOLE45_0;
	wire w_dff_A_p9D2YWv37_0;
	wire w_dff_A_wzPmPtWd8_0;
	wire w_dff_A_MNTDk6jt7_0;
	wire w_dff_A_gCGFNWpA0_0;
	wire w_dff_A_VvXUNJJr1_0;
	wire w_dff_A_lwpUp4NK5_0;
	wire w_dff_A_2zudnWq70_0;
	wire w_dff_A_YGHgvoIb8_0;
	wire w_dff_A_fVeXfF3y3_2;
	wire w_dff_A_o1WbTIJ53_0;
	wire w_dff_A_4eEuNoo61_0;
	wire w_dff_A_72v3frcJ4_0;
	wire w_dff_A_kZg1QiDS8_0;
	wire w_dff_A_mednfuaS8_0;
	wire w_dff_A_sY1vGI651_0;
	wire w_dff_A_rJL7EMod6_0;
	wire w_dff_A_5MfCJlFm8_0;
	wire w_dff_A_8GWrTFld8_0;
	wire w_dff_A_gpSTQkSQ4_0;
	wire w_dff_A_lSEFbcnH4_0;
	wire w_dff_A_4SzqUtKF6_0;
	wire w_dff_A_ZI9dAyYC3_0;
	wire w_dff_A_dAmQL6R87_0;
	wire w_dff_A_D2u1fAc26_0;
	wire w_dff_A_wYVFaF601_0;
	wire w_dff_A_2fVY5uF90_0;
	wire w_dff_A_d7CVs3OQ2_0;
	wire w_dff_A_Juhqcp5p3_0;
	wire w_dff_A_jdno4zPP3_0;
	wire w_dff_A_yeIoEjSc1_0;
	wire w_dff_A_qf7H07IF0_0;
	wire w_dff_A_eIEnfp250_0;
	wire w_dff_A_pACpSUQN8_0;
	wire w_dff_A_0k2YviDZ5_0;
	wire w_dff_A_pZYcFIXx1_0;
	wire w_dff_A_yC5XCXIo3_0;
	wire w_dff_A_Oupxy7zq7_0;
	wire w_dff_A_zfJQipgK6_0;
	wire w_dff_A_PjOAOSvb3_0;
	wire w_dff_A_ZM5WpisM4_0;
	wire w_dff_A_38XLV76J4_0;
	wire w_dff_A_C0jI8AXB2_0;
	wire w_dff_A_85cmRc3R2_0;
	wire w_dff_A_50UOJVWl2_0;
	wire w_dff_A_DLG9CSI75_0;
	wire w_dff_A_sV7XXod07_0;
	wire w_dff_A_Ib9ubb7Y3_0;
	wire w_dff_A_z6Bo6U7Z8_0;
	wire w_dff_A_b2Zd016Q4_0;
	wire w_dff_A_fcRqM66B9_0;
	wire w_dff_A_ermp00R91_0;
	wire w_dff_A_WUqcmPqk2_0;
	wire w_dff_A_CwN7wier7_0;
	wire w_dff_A_c5Mig13r5_0;
	wire w_dff_A_G76WnMkG0_0;
	wire w_dff_A_NJSYByyM6_0;
	wire w_dff_A_iFj29ikR8_0;
	wire w_dff_A_SYIDHwaH8_0;
	wire w_dff_A_1CylodWj4_0;
	wire w_dff_A_zcawgL1s4_0;
	wire w_dff_A_9NCRn5P10_0;
	wire w_dff_A_a0EdeibP0_0;
	wire w_dff_A_Nw1pbC711_0;
	wire w_dff_A_3Exa6QLI5_0;
	wire w_dff_A_1Uup38GA0_0;
	wire w_dff_A_e3Y5oSoZ5_0;
	wire w_dff_A_C3SSud2Z7_0;
	wire w_dff_A_KgomdcfT8_0;
	wire w_dff_A_67JOcsvH6_0;
	wire w_dff_A_cpxzsT6Z9_0;
	wire w_dff_A_wS98UYih4_0;
	wire w_dff_A_apv54JrL0_2;
	wire w_dff_A_dBAk415Y4_0;
	wire w_dff_A_laIz5X6W5_0;
	wire w_dff_A_IRpYVF7F6_0;
	wire w_dff_A_RxKwzf739_0;
	wire w_dff_A_2S5r6X6P3_0;
	wire w_dff_A_3Us7mh066_0;
	wire w_dff_A_CvCHQFPK6_0;
	wire w_dff_A_zw0oIhC57_0;
	wire w_dff_A_h2ZRzyZK2_0;
	wire w_dff_A_AJkqN9Z77_0;
	wire w_dff_A_UW7QAg7Q5_0;
	wire w_dff_A_jXKBgfSv4_0;
	wire w_dff_A_7uW6PcDh4_0;
	wire w_dff_A_uNczXrg00_0;
	wire w_dff_A_WmkES23T9_0;
	wire w_dff_A_TCzmEIA36_0;
	wire w_dff_A_wyR3Q9Rc4_0;
	wire w_dff_A_b6xjJOkB0_0;
	wire w_dff_A_Ayg9xbJf4_0;
	wire w_dff_A_0dCwa6hS4_0;
	wire w_dff_A_9C0bhD3t7_0;
	wire w_dff_A_xUTFGiiT1_0;
	wire w_dff_A_ytRNEqYc2_0;
	wire w_dff_A_04owxQqU3_0;
	wire w_dff_A_nN3yAUis8_0;
	wire w_dff_A_0mEhRKRq8_0;
	wire w_dff_A_MTpXKLcC3_0;
	wire w_dff_A_Ydmwoqxb1_0;
	wire w_dff_A_v40fqtLM3_0;
	wire w_dff_A_CVsD3srr9_0;
	wire w_dff_A_i8WMIx4R4_0;
	wire w_dff_A_7AXU1di97_0;
	wire w_dff_A_3MNZvNFh3_0;
	wire w_dff_A_CObArfJD6_0;
	wire w_dff_A_Hi4dpTD43_0;
	wire w_dff_A_Tr95Q3F94_0;
	wire w_dff_A_o17VLYLF1_0;
	wire w_dff_A_CjEBfkaa9_0;
	wire w_dff_A_JUnIpInf4_0;
	wire w_dff_A_YF1KtEL77_0;
	wire w_dff_A_URGOLNDV3_0;
	wire w_dff_A_MMghgGcf7_0;
	wire w_dff_A_di2VmveN6_0;
	wire w_dff_A_AFgb8HMT2_0;
	wire w_dff_A_yIC4WPEG8_0;
	wire w_dff_A_yNyn99U82_0;
	wire w_dff_A_0dWn8Spw9_0;
	wire w_dff_A_FPxhwbtW1_0;
	wire w_dff_A_qatcRyM88_0;
	wire w_dff_A_F043k6ju5_0;
	wire w_dff_A_rJWNtSpD6_0;
	wire w_dff_A_uZNWG3zu3_0;
	wire w_dff_A_1DIb0yIg8_0;
	wire w_dff_A_ZPEldzRF0_0;
	wire w_dff_A_bEHjzTA55_0;
	wire w_dff_A_BrBKtJlW8_0;
	wire w_dff_A_fDLHVQoQ9_0;
	wire w_dff_A_S3Nt75zP6_0;
	wire w_dff_A_xsOYTMRG8_0;
	wire w_dff_A_YUpDGpAj9_0;
	wire w_dff_A_W18ZItLa2_0;
	wire w_dff_A_u9JR45Q39_2;
	wire w_dff_A_a7kPmvzC1_0;
	wire w_dff_A_7FNMHEa77_0;
	wire w_dff_A_Qwgnt3vg5_0;
	wire w_dff_A_p3SR5rm08_0;
	wire w_dff_A_bAfZdBgC4_0;
	wire w_dff_A_ZcmVLl2Z3_0;
	wire w_dff_A_GXhe9woH1_0;
	wire w_dff_A_iZykjJyM7_0;
	wire w_dff_A_16kHkLPy9_0;
	wire w_dff_A_saj9RMhn5_0;
	wire w_dff_A_Y3xeWqjd5_0;
	wire w_dff_A_oXRebKbp3_0;
	wire w_dff_A_4aQmSl5r0_0;
	wire w_dff_A_IGXyLNWA5_0;
	wire w_dff_A_i3ZYYbKD0_0;
	wire w_dff_A_PT6v9qWd7_0;
	wire w_dff_A_1JHiii4c8_0;
	wire w_dff_A_DVPtnxHP0_0;
	wire w_dff_A_gUQf8DSC8_0;
	wire w_dff_A_0Mnqp26m1_0;
	wire w_dff_A_rlTXzyAW9_0;
	wire w_dff_A_QfBEi23Q6_0;
	wire w_dff_A_mDtT5sAP9_0;
	wire w_dff_A_9w8IdPq26_0;
	wire w_dff_A_fhqoxttH0_0;
	wire w_dff_A_d0Uepe1X4_0;
	wire w_dff_A_WCzqahEH2_0;
	wire w_dff_A_uV48ueqp1_0;
	wire w_dff_A_OESZUosL8_0;
	wire w_dff_A_FKwp4Rvw4_0;
	wire w_dff_A_4S07OXcP6_0;
	wire w_dff_A_GinmoGLY6_0;
	wire w_dff_A_9JNqIL4L4_0;
	wire w_dff_A_wtsJNKpU2_0;
	wire w_dff_A_F1ZE7YzQ0_0;
	wire w_dff_A_mDd66k3u4_0;
	wire w_dff_A_Qt2fUqli2_0;
	wire w_dff_A_MnWZZulQ5_0;
	wire w_dff_A_ZUUa9zWM5_0;
	wire w_dff_A_5TU1mqak4_0;
	wire w_dff_A_gDAlXsIW5_0;
	wire w_dff_A_Ht03QWsm3_0;
	wire w_dff_A_DEwoiM0B5_0;
	wire w_dff_A_HnCVEyRa4_0;
	wire w_dff_A_6ACEfJDP4_0;
	wire w_dff_A_6DQffS4r7_0;
	wire w_dff_A_rX2JkSeX4_0;
	wire w_dff_A_TMJkF1bT0_0;
	wire w_dff_A_epTUJaUk7_0;
	wire w_dff_A_vLvb4JyL5_0;
	wire w_dff_A_1QrB1juE3_0;
	wire w_dff_A_NSQRscGH1_0;
	wire w_dff_A_zutMZV7w2_0;
	wire w_dff_A_xqok4ro61_0;
	wire w_dff_A_wQidtS463_0;
	wire w_dff_A_2ldpwheP1_0;
	wire w_dff_A_DzL73d7t1_0;
	wire w_dff_A_aayfAdcH5_0;
	wire w_dff_A_d3nXRxgJ1_0;
	wire w_dff_A_9ozywqgS9_0;
	wire w_dff_A_Z4pRlS9P8_2;
	wire w_dff_A_T6Ac4q6P4_0;
	wire w_dff_A_e7T8cfxq1_0;
	wire w_dff_A_IrLFQIPX6_0;
	wire w_dff_A_A4JRQDsT1_0;
	wire w_dff_A_VZFsfBxM0_0;
	wire w_dff_A_6lua5B5g5_0;
	wire w_dff_A_ql2yu8Hy8_0;
	wire w_dff_A_bhHMrDYy8_0;
	wire w_dff_A_T3eqOZBl7_0;
	wire w_dff_A_hH2QfJjq6_0;
	wire w_dff_A_9NDLG0688_0;
	wire w_dff_A_nl88IL6c8_0;
	wire w_dff_A_HxzuLJOW6_0;
	wire w_dff_A_yeY0su3y6_0;
	wire w_dff_A_8oeH0eZr5_0;
	wire w_dff_A_8qJNKg2A8_0;
	wire w_dff_A_JihLZUbE8_0;
	wire w_dff_A_SBqhS0Rm0_0;
	wire w_dff_A_CmpFw6cr6_0;
	wire w_dff_A_OKZJTjQH0_0;
	wire w_dff_A_OsKbSxXn3_0;
	wire w_dff_A_fdp4NZXr5_0;
	wire w_dff_A_3EEOslsn8_0;
	wire w_dff_A_fAtbWiGN6_0;
	wire w_dff_A_gCvvaal76_0;
	wire w_dff_A_gnFjCrWj2_0;
	wire w_dff_A_pnErWyHg1_0;
	wire w_dff_A_8B1TxZJ64_0;
	wire w_dff_A_hOBxosRT4_0;
	wire w_dff_A_wZB0b1xB6_0;
	wire w_dff_A_nXNxlDSO0_0;
	wire w_dff_A_5U1Qd4AU7_0;
	wire w_dff_A_pRm0Pu0r9_0;
	wire w_dff_A_Rq4vNT679_0;
	wire w_dff_A_odVIc5ZV1_0;
	wire w_dff_A_7BoI3UZc9_0;
	wire w_dff_A_PkAvAav43_0;
	wire w_dff_A_SWqQ5eqI6_0;
	wire w_dff_A_e3fmwp449_0;
	wire w_dff_A_MVXNSLyo2_0;
	wire w_dff_A_VnSc2x1S6_0;
	wire w_dff_A_wie0GAka4_0;
	wire w_dff_A_u7h5RBDN1_0;
	wire w_dff_A_OhoNtRXj1_0;
	wire w_dff_A_F8UnrKcz5_0;
	wire w_dff_A_0eBV2Zsm0_0;
	wire w_dff_A_klwVrK1f0_0;
	wire w_dff_A_mCCNTPrw8_0;
	wire w_dff_A_bB1MRMHH5_0;
	wire w_dff_A_ptbj28cO4_0;
	wire w_dff_A_E3KHyVyE3_0;
	wire w_dff_A_1zBUEotC4_0;
	wire w_dff_A_pm7rt7Lx9_0;
	wire w_dff_A_XRa3pBrd2_0;
	wire w_dff_A_dpu9OwYR6_0;
	wire w_dff_A_NUyaeWkZ0_0;
	wire w_dff_A_oL8BaBJh7_0;
	wire w_dff_A_Pf3ReiLo4_0;
	wire w_dff_A_4mB0fYKv9_0;
	wire w_dff_A_RBUkAX7b8_2;
	wire w_dff_A_RqmSUKBW9_0;
	wire w_dff_A_k3slauRu1_0;
	wire w_dff_A_GOpyHYSR9_0;
	wire w_dff_A_8hxzPRz46_0;
	wire w_dff_A_QQYRPL7l8_0;
	wire w_dff_A_z0ZztFCX1_0;
	wire w_dff_A_IYRw5uzD3_0;
	wire w_dff_A_hTuqk3668_0;
	wire w_dff_A_HxuQcyJS4_0;
	wire w_dff_A_DtjwSTAQ8_0;
	wire w_dff_A_91SPmLkQ8_0;
	wire w_dff_A_BgtOKDIh5_0;
	wire w_dff_A_BrDzreaM9_0;
	wire w_dff_A_6HFMtDfJ2_0;
	wire w_dff_A_RAbNNNLW2_0;
	wire w_dff_A_bukx1VUX6_0;
	wire w_dff_A_5rsQSmNv9_0;
	wire w_dff_A_fRTuTzJI9_0;
	wire w_dff_A_Yz5CW6DV2_0;
	wire w_dff_A_dhICiPAr9_0;
	wire w_dff_A_2o5QjwcZ0_0;
	wire w_dff_A_EWVIJrGP1_0;
	wire w_dff_A_b3HXEpiv9_0;
	wire w_dff_A_W0wvWbet7_0;
	wire w_dff_A_B31JlHjo7_0;
	wire w_dff_A_zLAhlYtw6_0;
	wire w_dff_A_izwGJfV66_0;
	wire w_dff_A_b9yXsjgx3_0;
	wire w_dff_A_kj1KkzTv0_0;
	wire w_dff_A_HgO7x0Lc8_0;
	wire w_dff_A_u7WqldW85_0;
	wire w_dff_A_50gaQkM69_0;
	wire w_dff_A_ZKlQ6WzA5_0;
	wire w_dff_A_KUMl4IoR8_0;
	wire w_dff_A_XgqRKVkx9_0;
	wire w_dff_A_iCEoBT3I6_0;
	wire w_dff_A_hjkRxXNl3_0;
	wire w_dff_A_GSPv2VuK4_0;
	wire w_dff_A_06bO7B0w1_0;
	wire w_dff_A_zpECHwwR8_0;
	wire w_dff_A_Shfwh0Ce9_0;
	wire w_dff_A_wu1vCQuc4_0;
	wire w_dff_A_0TV2RpM41_0;
	wire w_dff_A_pB849hJ15_0;
	wire w_dff_A_fjVHhmRR4_0;
	wire w_dff_A_5HcNXxXi3_0;
	wire w_dff_A_bTgzmGKw0_0;
	wire w_dff_A_ANew8Hpr0_0;
	wire w_dff_A_gfOrLxGB4_0;
	wire w_dff_A_gkg8OXmv0_0;
	wire w_dff_A_qDRJvr5m6_0;
	wire w_dff_A_8gqkAWhr3_0;
	wire w_dff_A_ciX2eJ1s5_0;
	wire w_dff_A_sGm9nNKc4_0;
	wire w_dff_A_Op5Zb9bh7_0;
	wire w_dff_A_rouTpG8B3_0;
	wire w_dff_A_JrVaruuE8_0;
	wire w_dff_A_PnCdcSrA3_0;
	wire w_dff_A_VF0Og0Ap9_2;
	wire w_dff_A_nXroSYXR2_0;
	wire w_dff_A_aK1T7m2b4_0;
	wire w_dff_A_qDJPqAJt3_0;
	wire w_dff_A_FWJnlYk33_0;
	wire w_dff_A_OmtCMLWa8_0;
	wire w_dff_A_H2wdNp3t5_0;
	wire w_dff_A_TGmNPq249_0;
	wire w_dff_A_wX6PvLmZ4_0;
	wire w_dff_A_Q9EfKqwD2_0;
	wire w_dff_A_EOea4nGB1_0;
	wire w_dff_A_JXFJdGuC6_0;
	wire w_dff_A_95LZ5gRE2_0;
	wire w_dff_A_VEyQvFaV5_0;
	wire w_dff_A_v4u7p8A44_0;
	wire w_dff_A_71B6alZp2_0;
	wire w_dff_A_RVmWBXHU7_0;
	wire w_dff_A_HjRXXXPB7_0;
	wire w_dff_A_0xwNUpSI0_0;
	wire w_dff_A_tbiT7czn9_0;
	wire w_dff_A_2g3snXTF8_0;
	wire w_dff_A_7LsueYe93_0;
	wire w_dff_A_cXZ7DTNB5_0;
	wire w_dff_A_rpyI8TVa0_0;
	wire w_dff_A_BUDM2W8v1_0;
	wire w_dff_A_QilB8ZQ87_0;
	wire w_dff_A_rMMBb6jS4_0;
	wire w_dff_A_axOLZP2J1_0;
	wire w_dff_A_85XXMsKB6_0;
	wire w_dff_A_cqnHyzI32_0;
	wire w_dff_A_gyDLYRcc6_0;
	wire w_dff_A_t3uaLxwH3_0;
	wire w_dff_A_3LQGQ5d49_0;
	wire w_dff_A_TmS3uBVf2_0;
	wire w_dff_A_xqstLM2H5_0;
	wire w_dff_A_CZQzgRln7_0;
	wire w_dff_A_k3Jti8gx8_0;
	wire w_dff_A_qhgXhkMW8_0;
	wire w_dff_A_2J8ko5oa0_0;
	wire w_dff_A_q4P4oeuS3_0;
	wire w_dff_A_Zg312tyK9_0;
	wire w_dff_A_NmfKAelC5_0;
	wire w_dff_A_5UUxAp4w6_0;
	wire w_dff_A_nit1TOWV1_0;
	wire w_dff_A_10If2VMj9_0;
	wire w_dff_A_KSeGRj1L7_0;
	wire w_dff_A_8I7X3FGR3_0;
	wire w_dff_A_jbfB4KMr5_0;
	wire w_dff_A_WC0wZdX67_0;
	wire w_dff_A_xLg8XN027_0;
	wire w_dff_A_TNLK19AJ3_0;
	wire w_dff_A_H8Waqkww6_0;
	wire w_dff_A_1aZCad728_0;
	wire w_dff_A_hv5F2UiU6_0;
	wire w_dff_A_MGBGWR1K2_0;
	wire w_dff_A_dowjjR7S7_0;
	wire w_dff_A_Qcl0AmRC5_0;
	wire w_dff_A_BrfBedkC6_0;
	wire w_dff_A_uaH4n4Vl7_2;
	wire w_dff_A_Hq5zPYQD9_0;
	wire w_dff_A_Pecahs0b8_0;
	wire w_dff_A_gnoytxa32_0;
	wire w_dff_A_KzdkcyGv7_0;
	wire w_dff_A_hhdyFl8l3_0;
	wire w_dff_A_a814e7N81_0;
	wire w_dff_A_dsfP5vaW0_0;
	wire w_dff_A_Ja7mqpbw9_0;
	wire w_dff_A_NV2Dn7d30_0;
	wire w_dff_A_rYk6j1yo4_0;
	wire w_dff_A_ZyjSC7Iw3_0;
	wire w_dff_A_4InucV121_0;
	wire w_dff_A_QpiFVyba8_0;
	wire w_dff_A_QTfQJtRn0_0;
	wire w_dff_A_NsEimduf1_0;
	wire w_dff_A_hwrVZa7V8_0;
	wire w_dff_A_AbMD8cxu8_0;
	wire w_dff_A_hqNDzVSf2_0;
	wire w_dff_A_uXz3jG643_0;
	wire w_dff_A_onf41rlz9_0;
	wire w_dff_A_dL6cUK7B6_0;
	wire w_dff_A_weIgDyLp5_0;
	wire w_dff_A_XRZlYPQ88_0;
	wire w_dff_A_HkakeBHP5_0;
	wire w_dff_A_KT1eTXe82_0;
	wire w_dff_A_14p1WUOo1_0;
	wire w_dff_A_MtXNWzBZ7_0;
	wire w_dff_A_E4ejwqDF9_0;
	wire w_dff_A_yYu0LAmn5_0;
	wire w_dff_A_zwhA3urF5_0;
	wire w_dff_A_y3iSHKgA9_0;
	wire w_dff_A_ElFiynBr4_0;
	wire w_dff_A_bW1f51vt8_0;
	wire w_dff_A_kszowhPr5_0;
	wire w_dff_A_mTHsZxYA7_0;
	wire w_dff_A_hu4Fzncz4_0;
	wire w_dff_A_Q1edSFGu6_0;
	wire w_dff_A_LD2x6Hs68_0;
	wire w_dff_A_27Foccp19_0;
	wire w_dff_A_SnhIeawK0_0;
	wire w_dff_A_5933i80A5_0;
	wire w_dff_A_4yDJceyl1_0;
	wire w_dff_A_banPibvB0_0;
	wire w_dff_A_VcmAb1kX0_0;
	wire w_dff_A_T4DsH9M93_0;
	wire w_dff_A_JseL2veh6_0;
	wire w_dff_A_ObIID1MB1_0;
	wire w_dff_A_jRrr0lXe2_0;
	wire w_dff_A_2QTABo543_0;
	wire w_dff_A_JkhXQLb51_0;
	wire w_dff_A_u9L4L54q2_0;
	wire w_dff_A_KK3uU43V2_0;
	wire w_dff_A_ZSPUFDMw5_0;
	wire w_dff_A_OfVv51LF4_0;
	wire w_dff_A_AMHXt1sX3_0;
	wire w_dff_A_wtn1PM5s4_0;
	wire w_dff_A_25rg4D9y4_2;
	wire w_dff_A_gMaUZ1Jh2_0;
	wire w_dff_A_QDtMMZLA4_0;
	wire w_dff_A_z3ckPqi00_0;
	wire w_dff_A_bENZVi647_0;
	wire w_dff_A_vUWQXntf0_0;
	wire w_dff_A_pmwqGBGK4_0;
	wire w_dff_A_vefyXECb7_0;
	wire w_dff_A_sPN1vKtc6_0;
	wire w_dff_A_HEiSK3Hi9_0;
	wire w_dff_A_IwfVey4W3_0;
	wire w_dff_A_bY9n5lJI0_0;
	wire w_dff_A_NnrB3y8e7_0;
	wire w_dff_A_P3m1j59o6_0;
	wire w_dff_A_FCy7iKye6_0;
	wire w_dff_A_2kk1vipH4_0;
	wire w_dff_A_RQC1bsqx4_0;
	wire w_dff_A_MbW3SaUX7_0;
	wire w_dff_A_fkQ1ghpz0_0;
	wire w_dff_A_fFssae2R6_0;
	wire w_dff_A_ZnOTxnJF5_0;
	wire w_dff_A_vC8adhUD8_0;
	wire w_dff_A_Qf1RcdE39_0;
	wire w_dff_A_aDTZ1pvD4_0;
	wire w_dff_A_eJiRy7R26_0;
	wire w_dff_A_yIJEqPa52_0;
	wire w_dff_A_fYxJTW1N1_0;
	wire w_dff_A_mAVxwpLn9_0;
	wire w_dff_A_vc5pq8HC2_0;
	wire w_dff_A_M2WDqZ791_0;
	wire w_dff_A_jLVdDsl13_0;
	wire w_dff_A_cSQmsN7w0_0;
	wire w_dff_A_f7kUYoyW4_0;
	wire w_dff_A_dWnrxnrF5_0;
	wire w_dff_A_fNU093Xm9_0;
	wire w_dff_A_L03vf5bo3_0;
	wire w_dff_A_2vfH541f0_0;
	wire w_dff_A_VilYtPz80_0;
	wire w_dff_A_ktQotUcz1_0;
	wire w_dff_A_mHBWCIWG5_0;
	wire w_dff_A_qNZugnpd2_0;
	wire w_dff_A_flTF9aTV4_0;
	wire w_dff_A_OKoF0kGo8_0;
	wire w_dff_A_Ez745p549_0;
	wire w_dff_A_dJ4jmv8Z2_0;
	wire w_dff_A_zfrwsumQ8_0;
	wire w_dff_A_H9fWrUxV1_0;
	wire w_dff_A_ODj0rsdq4_0;
	wire w_dff_A_IyOT4q7o7_0;
	wire w_dff_A_jMp5qYgI5_0;
	wire w_dff_A_glD8vUMN1_0;
	wire w_dff_A_0GrgOJQn6_0;
	wire w_dff_A_8EHSVeXd8_0;
	wire w_dff_A_EwOzXb3T5_0;
	wire w_dff_A_CbmndSSj4_0;
	wire w_dff_A_iMzLpSO62_0;
	wire w_dff_A_DAfWDgLl4_2;
	wire w_dff_A_ormSNGoe1_0;
	wire w_dff_A_A4LRAPuQ9_0;
	wire w_dff_A_82FIWrjE3_0;
	wire w_dff_A_y4UVvr3y6_0;
	wire w_dff_A_ya35myYx5_0;
	wire w_dff_A_Lz4R1lWK5_0;
	wire w_dff_A_Zhq6baI88_0;
	wire w_dff_A_5LBMkHLK3_0;
	wire w_dff_A_y1S8iZjm6_0;
	wire w_dff_A_0q7vflWe0_0;
	wire w_dff_A_kvoyxFSh5_0;
	wire w_dff_A_6rq2NHXN9_0;
	wire w_dff_A_N6H7OTw20_0;
	wire w_dff_A_4s2LNkBy1_0;
	wire w_dff_A_DBd6t99U2_0;
	wire w_dff_A_TlhoMpTp2_0;
	wire w_dff_A_sXCjoh2K5_0;
	wire w_dff_A_rVVTBUHX2_0;
	wire w_dff_A_enFI1pD69_0;
	wire w_dff_A_6kmL7lfO7_0;
	wire w_dff_A_uZ5zQV233_0;
	wire w_dff_A_74mrreFB9_0;
	wire w_dff_A_P60Qy7Dr8_0;
	wire w_dff_A_tz9aYjWz2_0;
	wire w_dff_A_VIvHBkx90_0;
	wire w_dff_A_ZHWJkbpj3_0;
	wire w_dff_A_MFwOKpof3_0;
	wire w_dff_A_i5LCXn107_0;
	wire w_dff_A_6RK1onP97_0;
	wire w_dff_A_EFtX4gxT3_0;
	wire w_dff_A_gBmXod542_0;
	wire w_dff_A_qQ4ElGug8_0;
	wire w_dff_A_2sqKCUKN9_0;
	wire w_dff_A_O333e3BQ6_0;
	wire w_dff_A_itSpDTOm5_0;
	wire w_dff_A_snOHc84O4_0;
	wire w_dff_A_SxJRLB578_0;
	wire w_dff_A_QfYySoUh0_0;
	wire w_dff_A_UErrL4eL8_0;
	wire w_dff_A_ajGKrzye8_0;
	wire w_dff_A_7tJ5UrSc9_0;
	wire w_dff_A_dZzbELHd9_0;
	wire w_dff_A_HgeQCjLO0_0;
	wire w_dff_A_7L0cfby70_0;
	wire w_dff_A_eHO7v2ZO2_0;
	wire w_dff_A_yV0xkws93_0;
	wire w_dff_A_mkQ40IJp6_0;
	wire w_dff_A_fJOoY3RV1_0;
	wire w_dff_A_sfQWWVT60_0;
	wire w_dff_A_NDhZpc6m9_0;
	wire w_dff_A_cWvrTatd2_0;
	wire w_dff_A_7FniTJ6t0_0;
	wire w_dff_A_G8Up5KFD1_0;
	wire w_dff_A_ZNGIY1Kc2_0;
	wire w_dff_A_EXeMsU4S3_2;
	wire w_dff_A_Zln0oU877_0;
	wire w_dff_A_ddoOc77z5_0;
	wire w_dff_A_OeswcQRV0_0;
	wire w_dff_A_7bPWMjHM8_0;
	wire w_dff_A_Q3UYzNZ84_0;
	wire w_dff_A_UiloeydJ2_0;
	wire w_dff_A_OJk86uQq0_0;
	wire w_dff_A_2uAwSGJB2_0;
	wire w_dff_A_P84pQi9B8_0;
	wire w_dff_A_1v0ZCuPY3_0;
	wire w_dff_A_r4WMnlBu6_0;
	wire w_dff_A_vdf4uaYD4_0;
	wire w_dff_A_2kPOqpwC0_0;
	wire w_dff_A_kJcnqBpd1_0;
	wire w_dff_A_hT9RjCqx5_0;
	wire w_dff_A_26C6OUBy8_0;
	wire w_dff_A_rHv977LH6_0;
	wire w_dff_A_8yzyMVC58_0;
	wire w_dff_A_R0f9gUP06_0;
	wire w_dff_A_vpHkwVLa3_0;
	wire w_dff_A_57Z0k43U5_0;
	wire w_dff_A_AVXp5ds75_0;
	wire w_dff_A_UrXnx3686_0;
	wire w_dff_A_vExjHH2k7_0;
	wire w_dff_A_qIxMHUAc7_0;
	wire w_dff_A_DzVIQta27_0;
	wire w_dff_A_ir2Cgy7G3_0;
	wire w_dff_A_UTSAnnYM9_0;
	wire w_dff_A_oV688GxJ2_0;
	wire w_dff_A_CU9778F21_0;
	wire w_dff_A_y8nwg7Q93_0;
	wire w_dff_A_OSuq24jR4_0;
	wire w_dff_A_jGRYtIQz1_0;
	wire w_dff_A_abtHvNhj2_0;
	wire w_dff_A_8qJ5ZTYG0_0;
	wire w_dff_A_Q9Atw7Ot1_0;
	wire w_dff_A_OzSRRr1u3_0;
	wire w_dff_A_MhGw1nBV0_0;
	wire w_dff_A_JKg0nXE20_0;
	wire w_dff_A_ioolUZBx4_0;
	wire w_dff_A_FCmgRkDz2_0;
	wire w_dff_A_VesbgQ9o3_0;
	wire w_dff_A_pIdCw4Fc9_0;
	wire w_dff_A_BYQxwySx2_0;
	wire w_dff_A_pCp4hosc2_0;
	wire w_dff_A_fxe47mxL9_0;
	wire w_dff_A_E7txir177_0;
	wire w_dff_A_qRv1pvkc8_0;
	wire w_dff_A_MHwU2F0q6_0;
	wire w_dff_A_Gkfme8RG4_0;
	wire w_dff_A_niN05KA07_0;
	wire w_dff_A_YPqapSkP7_0;
	wire w_dff_A_6q3kG0Zq9_0;
	wire w_dff_A_kBneCYEu8_2;
	wire w_dff_A_TjZ8A8ix1_0;
	wire w_dff_A_1CiS67vV3_0;
	wire w_dff_A_z3bUp2Zk4_0;
	wire w_dff_A_vak0KR2D1_0;
	wire w_dff_A_24VX1jx52_0;
	wire w_dff_A_BBODrWsH3_0;
	wire w_dff_A_QZFHM5En2_0;
	wire w_dff_A_Wqhg9N3S4_0;
	wire w_dff_A_vXutZw1S8_0;
	wire w_dff_A_iciuHiHn6_0;
	wire w_dff_A_XcqqFZXf3_0;
	wire w_dff_A_VTwqFdWs4_0;
	wire w_dff_A_0cNmxHt89_0;
	wire w_dff_A_MLzdOCKr7_0;
	wire w_dff_A_fQHa6Clv4_0;
	wire w_dff_A_RsHvLwOe4_0;
	wire w_dff_A_8SA1rCrf5_0;
	wire w_dff_A_zp4Gajy60_0;
	wire w_dff_A_ZuFX1YDI5_0;
	wire w_dff_A_kptl2weY5_0;
	wire w_dff_A_pziyDUgK7_0;
	wire w_dff_A_W0DkZNNM0_0;
	wire w_dff_A_9EVxH0J33_0;
	wire w_dff_A_KgcQRq7J0_0;
	wire w_dff_A_ne4hKc6D9_0;
	wire w_dff_A_pUAhSRLv2_0;
	wire w_dff_A_kdHeE7md9_0;
	wire w_dff_A_BnSrrkiE1_0;
	wire w_dff_A_5oIOcmNt4_0;
	wire w_dff_A_soqyhzV73_0;
	wire w_dff_A_KOeJhbke1_0;
	wire w_dff_A_e0HoVtt94_0;
	wire w_dff_A_THonSYaz8_0;
	wire w_dff_A_kE2YiNZ35_0;
	wire w_dff_A_WgHD6dXx9_0;
	wire w_dff_A_jiVWknzQ8_0;
	wire w_dff_A_9xRPcLUh0_0;
	wire w_dff_A_eENqY71f0_0;
	wire w_dff_A_1nvxvxJw7_0;
	wire w_dff_A_myuGvPEX5_0;
	wire w_dff_A_zZ8XX7Im6_0;
	wire w_dff_A_m9GsMBpB0_0;
	wire w_dff_A_h6jeR5BS2_0;
	wire w_dff_A_JQXCwFgF8_0;
	wire w_dff_A_7TUpj4h75_0;
	wire w_dff_A_CyI9Vjt95_0;
	wire w_dff_A_1aMdhNC21_0;
	wire w_dff_A_y3Sh4eqa6_0;
	wire w_dff_A_fFGGIFZt1_0;
	wire w_dff_A_UTQRMyaE7_0;
	wire w_dff_A_tf7ayJ1u7_0;
	wire w_dff_A_no3YE7WY7_0;
	wire w_dff_A_50Y8hj8Y4_2;
	wire w_dff_A_380q8mam8_0;
	wire w_dff_A_X7oXyS1x2_0;
	wire w_dff_A_wpkHACFW3_0;
	wire w_dff_A_InvMEHLe4_0;
	wire w_dff_A_F5HCMXON9_0;
	wire w_dff_A_CfyqoSyP1_0;
	wire w_dff_A_toM6jEcl8_0;
	wire w_dff_A_pwGVKEoY9_0;
	wire w_dff_A_DZHNMTCB6_0;
	wire w_dff_A_4O5YjEMr2_0;
	wire w_dff_A_l8rg3K4r0_0;
	wire w_dff_A_coYJSFtM3_0;
	wire w_dff_A_QaFodfrU7_0;
	wire w_dff_A_6eLxX7186_0;
	wire w_dff_A_JqWqSuk32_0;
	wire w_dff_A_yhKe7tuk4_0;
	wire w_dff_A_4lsRD3MB4_0;
	wire w_dff_A_xnRVGa5p6_0;
	wire w_dff_A_dE1dSX6n5_0;
	wire w_dff_A_wYYNfpNG8_0;
	wire w_dff_A_ogNIVGzk8_0;
	wire w_dff_A_4mpehFMg3_0;
	wire w_dff_A_un4NtM2z2_0;
	wire w_dff_A_0XgpDvg60_0;
	wire w_dff_A_g1mL9q8a0_0;
	wire w_dff_A_UuSyHXzk4_0;
	wire w_dff_A_kf3VfFNM8_0;
	wire w_dff_A_BAYqhi505_0;
	wire w_dff_A_qfmkJNyU5_0;
	wire w_dff_A_IsOkEG7z2_0;
	wire w_dff_A_7UcO0olk3_0;
	wire w_dff_A_MC7xgw8y3_0;
	wire w_dff_A_6ZozluVv2_0;
	wire w_dff_A_NdlSg1HD2_0;
	wire w_dff_A_mWpxkfQk3_0;
	wire w_dff_A_0DbrXdlQ5_0;
	wire w_dff_A_LRVsfhoq9_0;
	wire w_dff_A_2kNjDGHY6_0;
	wire w_dff_A_ED7W3lqk3_0;
	wire w_dff_A_5T9p8brr2_0;
	wire w_dff_A_8XdNfzqJ0_0;
	wire w_dff_A_wnWDUmlG4_0;
	wire w_dff_A_cflT37il6_0;
	wire w_dff_A_RCc5bRBT7_0;
	wire w_dff_A_cYHMH3aM1_0;
	wire w_dff_A_eeJVynR56_0;
	wire w_dff_A_tN2npZYH6_0;
	wire w_dff_A_8uOQsRJz6_0;
	wire w_dff_A_xcl1jDOn2_0;
	wire w_dff_A_kluZOFwr9_0;
	wire w_dff_A_LNISbhLH8_0;
	wire w_dff_A_uKcBLu2n9_2;
	wire w_dff_A_HvNlbdOs7_0;
	wire w_dff_A_uQeD9Zd16_0;
	wire w_dff_A_m9g9yRsp0_0;
	wire w_dff_A_YZtPaWrA2_0;
	wire w_dff_A_bXAxPrgJ7_0;
	wire w_dff_A_QtZzEh6R8_0;
	wire w_dff_A_nMPD83vr7_0;
	wire w_dff_A_901p4X1c4_0;
	wire w_dff_A_tNy2uyJd2_0;
	wire w_dff_A_Z8HE94be5_0;
	wire w_dff_A_436MqNVQ4_0;
	wire w_dff_A_yBhTrM2j2_0;
	wire w_dff_A_nVf6cY2P2_0;
	wire w_dff_A_fOnTduJx7_0;
	wire w_dff_A_ZBjk75Cn0_0;
	wire w_dff_A_2Cz1N7jj6_0;
	wire w_dff_A_3198nwiY2_0;
	wire w_dff_A_TwRnH3f17_0;
	wire w_dff_A_439zFR8x0_0;
	wire w_dff_A_8mnjl5YU9_0;
	wire w_dff_A_RzUwzywh2_0;
	wire w_dff_A_HCsF6nf21_0;
	wire w_dff_A_jkqJqvUh4_0;
	wire w_dff_A_jWjWDhNx5_0;
	wire w_dff_A_vVNBJofN9_0;
	wire w_dff_A_LVqNfCzz6_0;
	wire w_dff_A_I813dbL64_0;
	wire w_dff_A_5zUbsZL49_0;
	wire w_dff_A_emKkbmS10_0;
	wire w_dff_A_Bk4Yr6xp4_0;
	wire w_dff_A_FpDYd6Yp6_0;
	wire w_dff_A_Iu8gJkor6_0;
	wire w_dff_A_22N3g46E3_0;
	wire w_dff_A_oh8Sdo6k9_0;
	wire w_dff_A_q6da7xD82_0;
	wire w_dff_A_x6zoRZYk4_0;
	wire w_dff_A_qVpcj7jv5_0;
	wire w_dff_A_6WeRIl7A2_0;
	wire w_dff_A_1KnrDZgR5_0;
	wire w_dff_A_zLGRwzUQ5_0;
	wire w_dff_A_jHVo2UKZ5_0;
	wire w_dff_A_m1zYb7NW7_0;
	wire w_dff_A_9UOwby586_0;
	wire w_dff_A_k0PgebVk0_0;
	wire w_dff_A_OfHSRyVS1_0;
	wire w_dff_A_F4I6rUl25_0;
	wire w_dff_A_xwxd4ajW3_0;
	wire w_dff_A_XEhTiZOz8_0;
	wire w_dff_A_xENpLPdo8_0;
	wire w_dff_A_mXdx3Ypa7_0;
	wire w_dff_A_RlfpDKF12_2;
	wire w_dff_A_4DonYcxZ2_0;
	wire w_dff_A_B8HDxOQy5_0;
	wire w_dff_A_vdCQwJgC2_0;
	wire w_dff_A_vA1ZdwEd9_0;
	wire w_dff_A_ARC4LZsm0_0;
	wire w_dff_A_mWnDcfIB9_0;
	wire w_dff_A_ypgRplGv0_0;
	wire w_dff_A_lsYs4WQt0_0;
	wire w_dff_A_nnz5RsiZ8_0;
	wire w_dff_A_giFPkiTO9_0;
	wire w_dff_A_SXJ0q3Ks3_0;
	wire w_dff_A_3LmmaxXn8_0;
	wire w_dff_A_LtTDJPZR2_0;
	wire w_dff_A_foT4pxeZ4_0;
	wire w_dff_A_53QzjAf81_0;
	wire w_dff_A_ATpHjgT78_0;
	wire w_dff_A_e0VT6QzL4_0;
	wire w_dff_A_TWdJP5VH8_0;
	wire w_dff_A_q6F8wKw01_0;
	wire w_dff_A_SpF0upsw2_0;
	wire w_dff_A_YBnZHitN9_0;
	wire w_dff_A_jUQBAWXz9_0;
	wire w_dff_A_ecF1bpiO2_0;
	wire w_dff_A_cwxLrvwG9_0;
	wire w_dff_A_3Kv7FAwT0_0;
	wire w_dff_A_MBDL2fvX3_0;
	wire w_dff_A_S8ebt1Q11_0;
	wire w_dff_A_8fdtYeUp9_0;
	wire w_dff_A_mjXGhLxS5_0;
	wire w_dff_A_cmY9OMeK1_0;
	wire w_dff_A_izxOmPK24_0;
	wire w_dff_A_VBE13euG9_0;
	wire w_dff_A_YmhU2R6U4_0;
	wire w_dff_A_uFiOsNo44_0;
	wire w_dff_A_zRjKlspb3_0;
	wire w_dff_A_hFvNIyOM3_0;
	wire w_dff_A_kduNNEDK6_0;
	wire w_dff_A_wCA7ujOc8_0;
	wire w_dff_A_XyI67h5D6_0;
	wire w_dff_A_N1xKqrTB1_0;
	wire w_dff_A_OaeHKZhR1_0;
	wire w_dff_A_VqOlsUEJ2_0;
	wire w_dff_A_Wt42TrZY5_0;
	wire w_dff_A_cD2vn7133_0;
	wire w_dff_A_kINq8yqh2_0;
	wire w_dff_A_QSEBN0SL5_0;
	wire w_dff_A_l8H9QYxj0_0;
	wire w_dff_A_XD0GEFeW7_0;
	wire w_dff_A_OxCjHqpa7_0;
	wire w_dff_A_yWmtd95Z9_2;
	wire w_dff_A_qkZtBiSq1_0;
	wire w_dff_A_tScFh3Kl2_0;
	wire w_dff_A_36M7cNzF5_0;
	wire w_dff_A_CndEV1K92_0;
	wire w_dff_A_0h25dN1D6_0;
	wire w_dff_A_oHXhD8j22_0;
	wire w_dff_A_bHuRnmKC2_0;
	wire w_dff_A_F3vpQvgn6_0;
	wire w_dff_A_mZHBLTom4_0;
	wire w_dff_A_etzstDjs6_0;
	wire w_dff_A_AyGB1ZTc0_0;
	wire w_dff_A_SJUkpxY93_0;
	wire w_dff_A_mP6XtOfq4_0;
	wire w_dff_A_zfvjm2bz1_0;
	wire w_dff_A_YPoHV4Kg3_0;
	wire w_dff_A_PVCzV6Ho8_0;
	wire w_dff_A_WmuU9RFK7_0;
	wire w_dff_A_pMmWgtmU4_0;
	wire w_dff_A_RdlQZcB12_0;
	wire w_dff_A_ggR422Dh2_0;
	wire w_dff_A_ncWh2HX84_0;
	wire w_dff_A_l70S9Sxu5_0;
	wire w_dff_A_23pVAkUT1_0;
	wire w_dff_A_ib1426oH9_0;
	wire w_dff_A_b1EAwoEw3_0;
	wire w_dff_A_2zek97ag8_0;
	wire w_dff_A_oWryYxg27_0;
	wire w_dff_A_AXf38r8r6_0;
	wire w_dff_A_RQCD9r8D8_0;
	wire w_dff_A_iy1CD8ki6_0;
	wire w_dff_A_BZ7rYHzE1_0;
	wire w_dff_A_W74HFkOY5_0;
	wire w_dff_A_zdvoRqev6_0;
	wire w_dff_A_hOMlBEIg4_0;
	wire w_dff_A_PziKTnu00_0;
	wire w_dff_A_NcUkuUVK3_0;
	wire w_dff_A_KIpAsP4F0_0;
	wire w_dff_A_1PBDSoX25_0;
	wire w_dff_A_F8AbN9jj0_0;
	wire w_dff_A_bCu22zD62_0;
	wire w_dff_A_7C6icvPk2_0;
	wire w_dff_A_jMSl0l025_0;
	wire w_dff_A_FVKZY5wV7_0;
	wire w_dff_A_x7UftJps5_0;
	wire w_dff_A_MjHkPadH7_0;
	wire w_dff_A_mgVfQPcp4_0;
	wire w_dff_A_L3MUWpVP2_0;
	wire w_dff_A_ESH7nihC7_0;
	wire w_dff_A_iULoKlkx1_2;
	wire w_dff_A_hRb1WDEa6_0;
	wire w_dff_A_Lda5KRtg5_0;
	wire w_dff_A_bFIitHTF7_0;
	wire w_dff_A_XeOhAS495_0;
	wire w_dff_A_EIGSAZnU0_0;
	wire w_dff_A_suP6yMeK3_0;
	wire w_dff_A_eVjXcTaJ5_0;
	wire w_dff_A_B2RowLKo8_0;
	wire w_dff_A_u5SecGSH2_0;
	wire w_dff_A_F8FMi8VD0_0;
	wire w_dff_A_IuH4HrD66_0;
	wire w_dff_A_MXfMiRkz0_0;
	wire w_dff_A_KLf448jv9_0;
	wire w_dff_A_w2DZAeCL5_0;
	wire w_dff_A_qUQu7PYp3_0;
	wire w_dff_A_DW3tUMo90_0;
	wire w_dff_A_ml40Ebtd9_0;
	wire w_dff_A_2q0z7P6E9_0;
	wire w_dff_A_euZLH25e8_0;
	wire w_dff_A_PZ7SHKic2_0;
	wire w_dff_A_WJch9ZpO9_0;
	wire w_dff_A_quIVjniU2_0;
	wire w_dff_A_M7Q6Agcq9_0;
	wire w_dff_A_7oMQAG7l5_0;
	wire w_dff_A_dzsqJTU21_0;
	wire w_dff_A_IkcQABtj1_0;
	wire w_dff_A_GPFCbRyC3_0;
	wire w_dff_A_SX7vW9ct8_0;
	wire w_dff_A_0LazYeen7_0;
	wire w_dff_A_BoEdLu2e2_0;
	wire w_dff_A_r2SqBUtD8_0;
	wire w_dff_A_0k217cT47_0;
	wire w_dff_A_jd6fyX7m2_0;
	wire w_dff_A_oDXlhhnW8_0;
	wire w_dff_A_VzuZuzZi1_0;
	wire w_dff_A_fG4EvSUN6_0;
	wire w_dff_A_IJnyghi77_0;
	wire w_dff_A_rdCuDiAg3_0;
	wire w_dff_A_wUqX7ldH1_0;
	wire w_dff_A_q1rZZC0K4_0;
	wire w_dff_A_EHbPQLf29_0;
	wire w_dff_A_oBp2Hrva8_0;
	wire w_dff_A_0glMPIVS2_0;
	wire w_dff_A_a96g5GQv4_0;
	wire w_dff_A_8rK7WVdA8_0;
	wire w_dff_A_Td3y2RKm7_0;
	wire w_dff_A_8gHFPLMH2_0;
	wire w_dff_A_E95bjTHE6_2;
	wire w_dff_A_EkTlbwSF6_0;
	wire w_dff_A_VJtmhJed3_0;
	wire w_dff_A_ory6Rcro9_0;
	wire w_dff_A_789X5lqI1_0;
	wire w_dff_A_AWe4MnpT8_0;
	wire w_dff_A_OFWlbXqg9_0;
	wire w_dff_A_1I04ukaw6_0;
	wire w_dff_A_hjd4ZPIZ3_0;
	wire w_dff_A_bPECUQSg4_0;
	wire w_dff_A_tANPOkyx9_0;
	wire w_dff_A_5LxVsuub5_0;
	wire w_dff_A_734NZw6D6_0;
	wire w_dff_A_GuJyUhbp0_0;
	wire w_dff_A_XJkQ9pqk1_0;
	wire w_dff_A_EmnbvvHE2_0;
	wire w_dff_A_X5g9KCer4_0;
	wire w_dff_A_Q1MI5oLg1_0;
	wire w_dff_A_u5SGxHBw3_0;
	wire w_dff_A_rrICQaGk4_0;
	wire w_dff_A_pGcTZ0tE1_0;
	wire w_dff_A_7BWyScQ28_0;
	wire w_dff_A_O8l17WgZ1_0;
	wire w_dff_A_153vyNHY4_0;
	wire w_dff_A_wmySegux3_0;
	wire w_dff_A_HI40fgjV3_0;
	wire w_dff_A_1SrDlBC40_0;
	wire w_dff_A_IQzhHR6F4_0;
	wire w_dff_A_BkzKRszD2_0;
	wire w_dff_A_h04rrvJB1_0;
	wire w_dff_A_t0tkoMpx9_0;
	wire w_dff_A_bZQhJkMe0_0;
	wire w_dff_A_zaiFWFK59_0;
	wire w_dff_A_3GXMC9mH3_0;
	wire w_dff_A_aiQTVfsj5_0;
	wire w_dff_A_fvxgQ0L95_0;
	wire w_dff_A_2IzbuGBO9_0;
	wire w_dff_A_gzYSSEkJ2_0;
	wire w_dff_A_Y6FuboB72_0;
	wire w_dff_A_YLFp524t3_0;
	wire w_dff_A_deaxy2T96_0;
	wire w_dff_A_peUlOvJM1_0;
	wire w_dff_A_lB3oYaCR8_0;
	wire w_dff_A_vWLF5Wq77_0;
	wire w_dff_A_zmnA5sqz5_0;
	wire w_dff_A_AZUNBJU43_0;
	wire w_dff_A_JbtFcLIb4_0;
	wire w_dff_A_5ajlcE7V4_2;
	wire w_dff_A_yrq8RRxb6_0;
	wire w_dff_A_SRMDKckD6_0;
	wire w_dff_A_VrxVSJdl0_0;
	wire w_dff_A_RlvhMH4m9_0;
	wire w_dff_A_10ixQL8w0_0;
	wire w_dff_A_02uvXEfK9_0;
	wire w_dff_A_Y4iLZifS1_0;
	wire w_dff_A_AKZN3ET33_0;
	wire w_dff_A_L2vIkbfK1_0;
	wire w_dff_A_AUzPE6SA3_0;
	wire w_dff_A_bGLFVMNg6_0;
	wire w_dff_A_ovTPSDu90_0;
	wire w_dff_A_4jttJpBA9_0;
	wire w_dff_A_NDIwV7dc8_0;
	wire w_dff_A_CZ6Mui0E3_0;
	wire w_dff_A_Z3GL3A8L0_0;
	wire w_dff_A_1ojMFOxX6_0;
	wire w_dff_A_CbEU7rhi9_0;
	wire w_dff_A_9v7iZBZt6_0;
	wire w_dff_A_ahTrYK8P6_0;
	wire w_dff_A_1ojEdrYW0_0;
	wire w_dff_A_eIiR2u5o9_0;
	wire w_dff_A_Z1HHw6HT0_0;
	wire w_dff_A_0BLxCuJ03_0;
	wire w_dff_A_2IaUoFT26_0;
	wire w_dff_A_C1w00jop1_0;
	wire w_dff_A_P0TcQm7r4_0;
	wire w_dff_A_MTh4EHZj9_0;
	wire w_dff_A_uNYNhFHg7_0;
	wire w_dff_A_8H2zzh131_0;
	wire w_dff_A_5HtWgcmt4_0;
	wire w_dff_A_KHt6XktR9_0;
	wire w_dff_A_W1JBg2YO2_0;
	wire w_dff_A_SCF40G4p1_0;
	wire w_dff_A_Pmso16Wt4_0;
	wire w_dff_A_iBITEoki8_0;
	wire w_dff_A_w9QRzCAq2_0;
	wire w_dff_A_AxUGuuMg0_0;
	wire w_dff_A_CeEVVqsP7_0;
	wire w_dff_A_JWbKkE1b5_0;
	wire w_dff_A_GY1PQSS14_0;
	wire w_dff_A_peXopZp01_0;
	wire w_dff_A_CxEFWK3D9_0;
	wire w_dff_A_ZXdXoEhP7_0;
	wire w_dff_A_9DMIZN2c4_0;
	wire w_dff_A_Xic2Adtu8_2;
	wire w_dff_A_ae3fN4sz7_0;
	wire w_dff_A_QH3nMiW09_0;
	wire w_dff_A_8KTAWJsc8_0;
	wire w_dff_A_pwhuY45Y9_0;
	wire w_dff_A_CTN0kwmC8_0;
	wire w_dff_A_puY2T0OV1_0;
	wire w_dff_A_an8NgWan7_0;
	wire w_dff_A_zX5ZeUkR1_0;
	wire w_dff_A_E2iaVVUK0_0;
	wire w_dff_A_ZuXgAFUx9_0;
	wire w_dff_A_NGl7jE5l4_0;
	wire w_dff_A_9gwTamw38_0;
	wire w_dff_A_j7WgJTx71_0;
	wire w_dff_A_V65MCLsK6_0;
	wire w_dff_A_uSeQGyzD7_0;
	wire w_dff_A_oLANuLxA6_0;
	wire w_dff_A_kD0lhMUr7_0;
	wire w_dff_A_psXX62it7_0;
	wire w_dff_A_meDuEnw66_0;
	wire w_dff_A_sLnJVsKA3_0;
	wire w_dff_A_QsLVnZK26_0;
	wire w_dff_A_ZEWEmoHY3_0;
	wire w_dff_A_VkMBIxlN5_0;
	wire w_dff_A_UNfluSTA0_0;
	wire w_dff_A_qKZ87JSS6_0;
	wire w_dff_A_3bZjeuQH4_0;
	wire w_dff_A_AWxnT9AG4_0;
	wire w_dff_A_6cvzohV45_0;
	wire w_dff_A_UsTjmVRQ3_0;
	wire w_dff_A_rR8zS27X9_0;
	wire w_dff_A_4ZqyfDqN2_0;
	wire w_dff_A_O3GU8iZ41_0;
	wire w_dff_A_99ZTIEvf8_0;
	wire w_dff_A_8B4xFIAQ8_0;
	wire w_dff_A_JxyxPhpD7_0;
	wire w_dff_A_r7pYV3yF9_0;
	wire w_dff_A_AbmCaJOa0_0;
	wire w_dff_A_uxrj627s5_0;
	wire w_dff_A_ezZdDTRe3_0;
	wire w_dff_A_fvd9W8f35_0;
	wire w_dff_A_JZpUUvKC0_0;
	wire w_dff_A_YNha8dyU4_0;
	wire w_dff_A_MSYyxAlT7_0;
	wire w_dff_A_nfprwjxH9_0;
	wire w_dff_A_4p69wJXZ0_2;
	wire w_dff_A_w6swdRjt0_0;
	wire w_dff_A_DYyitRvE0_0;
	wire w_dff_A_kDoJtfHJ4_0;
	wire w_dff_A_hwk1w0Aw7_0;
	wire w_dff_A_WE2zlTBT3_0;
	wire w_dff_A_pj09o6s77_0;
	wire w_dff_A_PhFsf0Zp3_0;
	wire w_dff_A_QvzyRWzt3_0;
	wire w_dff_A_4VF5fkN18_0;
	wire w_dff_A_Z7Zqzz4r7_0;
	wire w_dff_A_BCFbvDCh8_0;
	wire w_dff_A_2otiWYib1_0;
	wire w_dff_A_JotKQPNE3_0;
	wire w_dff_A_r4M2cirP2_0;
	wire w_dff_A_GfUjDvhG3_0;
	wire w_dff_A_9NAaC6I83_0;
	wire w_dff_A_e32dyhpt2_0;
	wire w_dff_A_xZn3NlHG0_0;
	wire w_dff_A_Em9QqonB7_0;
	wire w_dff_A_fK589tDi0_0;
	wire w_dff_A_gGxVkSsJ6_0;
	wire w_dff_A_7dXuuxyI1_0;
	wire w_dff_A_p0Pr2fSO0_0;
	wire w_dff_A_AHH1acAs2_0;
	wire w_dff_A_0BETMRhT9_0;
	wire w_dff_A_tZHuPoOe4_0;
	wire w_dff_A_RvQ9PZEn5_0;
	wire w_dff_A_f1kVDeZt4_0;
	wire w_dff_A_DSas78eH1_0;
	wire w_dff_A_2NUdOyvW2_0;
	wire w_dff_A_lD6CANcD9_0;
	wire w_dff_A_0piiSHpC6_0;
	wire w_dff_A_1rj5URsD7_0;
	wire w_dff_A_hZ5QwYQ18_0;
	wire w_dff_A_0tirzuB48_0;
	wire w_dff_A_tQuJ6dAA6_0;
	wire w_dff_A_SNJKiRpp2_0;
	wire w_dff_A_rdkxDQHx8_0;
	wire w_dff_A_ucC8WALG7_0;
	wire w_dff_A_PWtwCDQG6_0;
	wire w_dff_A_V9eJRzxA7_0;
	wire w_dff_A_Pvlm2YmH9_0;
	wire w_dff_A_no2IkSJL9_0;
	wire w_dff_A_BzE0H6ap0_2;
	wire w_dff_A_jqXYV3io5_0;
	wire w_dff_A_iM3cI7Ek6_0;
	wire w_dff_A_iN6VqhOQ0_0;
	wire w_dff_A_k2dItjQP9_0;
	wire w_dff_A_5gdDEE0T4_0;
	wire w_dff_A_8bikkJeO1_0;
	wire w_dff_A_82vovMh69_0;
	wire w_dff_A_gxoAJqr45_0;
	wire w_dff_A_Sr6lQnSW3_0;
	wire w_dff_A_zGojD2vJ2_0;
	wire w_dff_A_4CVwlnPI9_0;
	wire w_dff_A_tYwnkX7K0_0;
	wire w_dff_A_fbUEDZNy0_0;
	wire w_dff_A_pypTNgHF6_0;
	wire w_dff_A_uP2eD7y00_0;
	wire w_dff_A_oqehDbgi8_0;
	wire w_dff_A_5woHGs6L2_0;
	wire w_dff_A_lKDEsdBe9_0;
	wire w_dff_A_j3ETKEMN7_0;
	wire w_dff_A_36FGHFrT1_0;
	wire w_dff_A_RBktoPcE9_0;
	wire w_dff_A_jP9anIDS5_0;
	wire w_dff_A_RA90Km4p2_0;
	wire w_dff_A_O9mtDMsS0_0;
	wire w_dff_A_sIaRBHlt7_0;
	wire w_dff_A_KtB7i6bB7_0;
	wire w_dff_A_BktbEgcv8_0;
	wire w_dff_A_gmnaJajv8_0;
	wire w_dff_A_X1nZomeb0_0;
	wire w_dff_A_dIw0KlYv2_0;
	wire w_dff_A_LxkoDsqn5_0;
	wire w_dff_A_noRtGyXv7_0;
	wire w_dff_A_43sNXuGm1_0;
	wire w_dff_A_6zOs2XEH1_0;
	wire w_dff_A_OM6j7uCh3_0;
	wire w_dff_A_o1R1GBQb2_0;
	wire w_dff_A_XvBrxUTX9_0;
	wire w_dff_A_XSKLV1JD8_0;
	wire w_dff_A_AsBXM55u6_0;
	wire w_dff_A_6HtQQHLd3_0;
	wire w_dff_A_vY6mp8l88_0;
	wire w_dff_A_yV6ELeiR1_0;
	wire w_dff_A_TrXEhtji4_2;
	wire w_dff_A_mpLTf4219_0;
	wire w_dff_A_TdqsOJT54_0;
	wire w_dff_A_65dX4yMa8_0;
	wire w_dff_A_1ZBM88Ll0_0;
	wire w_dff_A_izqwe0jp3_0;
	wire w_dff_A_GIYMBYEK8_0;
	wire w_dff_A_hS0PaYuw6_0;
	wire w_dff_A_0TknbbLh5_0;
	wire w_dff_A_2fCd8o253_0;
	wire w_dff_A_e8aMue1E6_0;
	wire w_dff_A_6svRrmX85_0;
	wire w_dff_A_7G0JMF6y4_0;
	wire w_dff_A_Zx36iGOO1_0;
	wire w_dff_A_LdHkQoIm5_0;
	wire w_dff_A_XF8NdbBB3_0;
	wire w_dff_A_m8NfSNeS9_0;
	wire w_dff_A_Lmimkaom8_0;
	wire w_dff_A_o23dxbw04_0;
	wire w_dff_A_WVIy7PyL2_0;
	wire w_dff_A_egOplusY3_0;
	wire w_dff_A_RphwYfE68_0;
	wire w_dff_A_kKuXQA7Z0_0;
	wire w_dff_A_KhMiOUSE8_0;
	wire w_dff_A_nQ3r0zES9_0;
	wire w_dff_A_fT2aOutz6_0;
	wire w_dff_A_nfqndw8i1_0;
	wire w_dff_A_1IWjK4N52_0;
	wire w_dff_A_ssx3bLXm1_0;
	wire w_dff_A_KtaWNVou5_0;
	wire w_dff_A_Nx4XsKVS1_0;
	wire w_dff_A_bZe6fj7x7_0;
	wire w_dff_A_P2tHqJUu4_0;
	wire w_dff_A_G27dZytw9_0;
	wire w_dff_A_rq0lcUhd8_0;
	wire w_dff_A_FNArPyWS6_0;
	wire w_dff_A_sTBbMO137_0;
	wire w_dff_A_FUmyjLvz8_0;
	wire w_dff_A_CVFYPaIh5_0;
	wire w_dff_A_wzfi7FZF1_0;
	wire w_dff_A_BfRZoENc7_0;
	wire w_dff_A_cf7dJh6C1_0;
	wire w_dff_A_HRCPkfMi4_2;
	wire w_dff_A_2rSjB1rj9_0;
	wire w_dff_A_iqMRMa617_0;
	wire w_dff_A_6Fm8woOG7_0;
	wire w_dff_A_1lyaeRjh6_0;
	wire w_dff_A_k0ULkyCV0_0;
	wire w_dff_A_Ehiqzdjb8_0;
	wire w_dff_A_qirzyIXZ2_0;
	wire w_dff_A_O4Pu32G29_0;
	wire w_dff_A_gwExHQ2I9_0;
	wire w_dff_A_JgJFqoPU0_0;
	wire w_dff_A_qXjWXTUg2_0;
	wire w_dff_A_ZQ9de3FM2_0;
	wire w_dff_A_xXRfod5m7_0;
	wire w_dff_A_mQWgElrW4_0;
	wire w_dff_A_7HuCOhJ69_0;
	wire w_dff_A_NP7LGG3o7_0;
	wire w_dff_A_l2hV5m1P4_0;
	wire w_dff_A_HfKafrgH8_0;
	wire w_dff_A_Gtybz85Q5_0;
	wire w_dff_A_s9rS4OiU4_0;
	wire w_dff_A_FDAwbgv15_0;
	wire w_dff_A_Lc4MaL958_0;
	wire w_dff_A_lA7XbW9O8_0;
	wire w_dff_A_nBj4Wp078_0;
	wire w_dff_A_MujaL6on7_0;
	wire w_dff_A_WQ6erECb2_0;
	wire w_dff_A_Ga2QGedC7_0;
	wire w_dff_A_k4aPPfJc9_0;
	wire w_dff_A_arGQulI27_0;
	wire w_dff_A_5LKyl36z9_0;
	wire w_dff_A_3dajWwuL6_0;
	wire w_dff_A_y751QZU46_0;
	wire w_dff_A_uM1C7RSr4_0;
	wire w_dff_A_piPDTxBJ9_0;
	wire w_dff_A_QaAUtGFn1_0;
	wire w_dff_A_YPwmxXCC7_0;
	wire w_dff_A_wTOgwcv32_0;
	wire w_dff_A_qn030i954_0;
	wire w_dff_A_4QHExuNR0_0;
	wire w_dff_A_eTDEE6CM9_0;
	wire w_dff_A_OCpaXqst8_2;
	wire w_dff_A_aL5mmWiS6_0;
	wire w_dff_A_bH462nvr3_0;
	wire w_dff_A_JTtXoK2j6_0;
	wire w_dff_A_pJWDczQd6_0;
	wire w_dff_A_eF43UynL5_0;
	wire w_dff_A_2F4wQ4656_0;
	wire w_dff_A_dodhWfV67_0;
	wire w_dff_A_M85m3UCZ3_0;
	wire w_dff_A_k5mq6NGH2_0;
	wire w_dff_A_45qwoUnC1_0;
	wire w_dff_A_Zm8yimOu9_0;
	wire w_dff_A_FtVypjpd1_0;
	wire w_dff_A_0NQCeKcb4_0;
	wire w_dff_A_oyOid39a5_0;
	wire w_dff_A_YS9ywHnL6_0;
	wire w_dff_A_jpXggtwh9_0;
	wire w_dff_A_dnUP1o4t7_0;
	wire w_dff_A_VcZJVNcg1_0;
	wire w_dff_A_asYK8RaT8_0;
	wire w_dff_A_g7nJLmRe3_0;
	wire w_dff_A_zaoU9vPq4_0;
	wire w_dff_A_W5OoMSxm9_0;
	wire w_dff_A_5JaNrVKA2_0;
	wire w_dff_A_2gtmGbdx0_0;
	wire w_dff_A_0J3tUHCV0_0;
	wire w_dff_A_o2qh2RJa6_0;
	wire w_dff_A_BNOrYJj89_0;
	wire w_dff_A_HUqCe9rY8_0;
	wire w_dff_A_Au62QzpP0_0;
	wire w_dff_A_nqEkH5jt7_0;
	wire w_dff_A_md8dCJji6_0;
	wire w_dff_A_YPHI7fn75_0;
	wire w_dff_A_hUAL0c5w9_0;
	wire w_dff_A_yGXTXH4b5_0;
	wire w_dff_A_scTJkbhP1_0;
	wire w_dff_A_kVrUBjav0_0;
	wire w_dff_A_ry5okceN1_0;
	wire w_dff_A_TatD4bdV2_0;
	wire w_dff_A_izocvOpF5_0;
	wire w_dff_A_LDFLxawb9_2;
	wire w_dff_A_tHuYhkTX8_0;
	wire w_dff_A_hLRD023M9_0;
	wire w_dff_A_s5yBq3Zu2_0;
	wire w_dff_A_H28RLnpR3_0;
	wire w_dff_A_fHKYOYnC1_0;
	wire w_dff_A_vASC2l875_0;
	wire w_dff_A_GL1cxy0p6_0;
	wire w_dff_A_4hgHlFrK8_0;
	wire w_dff_A_3V51jYAo2_0;
	wire w_dff_A_nYbXU8e86_0;
	wire w_dff_A_MQ1dVrCQ4_0;
	wire w_dff_A_hRaXDNNJ6_0;
	wire w_dff_A_9f2K14Wl0_0;
	wire w_dff_A_A0IN27wo8_0;
	wire w_dff_A_YAtJlaxc2_0;
	wire w_dff_A_ntlwEz2f3_0;
	wire w_dff_A_C4D9PtUC8_0;
	wire w_dff_A_kXJN3uGx6_0;
	wire w_dff_A_f2QHW6iK3_0;
	wire w_dff_A_bYB5QZVH1_0;
	wire w_dff_A_b5K3EeYA0_0;
	wire w_dff_A_LyHIUixr3_0;
	wire w_dff_A_Q5eV4ttV0_0;
	wire w_dff_A_buEUpT5x9_0;
	wire w_dff_A_a9Cq3sRo7_0;
	wire w_dff_A_O24ThT117_0;
	wire w_dff_A_K18XR8Xr6_0;
	wire w_dff_A_j2NTQjsH6_0;
	wire w_dff_A_WhluNXyf6_0;
	wire w_dff_A_9xtWOCfE8_0;
	wire w_dff_A_NvOBlU3t9_0;
	wire w_dff_A_dCFjroEQ9_0;
	wire w_dff_A_4Z7M4SiK4_0;
	wire w_dff_A_AJCKv0OJ9_0;
	wire w_dff_A_D96b6KHj4_0;
	wire w_dff_A_QHQsfEFF3_0;
	wire w_dff_A_A6Dz6kOs4_0;
	wire w_dff_A_n1lhhwon3_0;
	wire w_dff_A_6JucvmkC3_2;
	wire w_dff_A_r8Uz5tCr3_0;
	wire w_dff_A_y5A7ROmk9_0;
	wire w_dff_A_q7qUTkmZ4_0;
	wire w_dff_A_9Ba0qRj96_0;
	wire w_dff_A_mBnU1qsY4_0;
	wire w_dff_A_bJgbDpJn3_0;
	wire w_dff_A_BbDa7xMc0_0;
	wire w_dff_A_wVRommd89_0;
	wire w_dff_A_C6jrz7uf4_0;
	wire w_dff_A_VTxTo4Xn0_0;
	wire w_dff_A_909EZ1Vm2_0;
	wire w_dff_A_hHV0onUZ0_0;
	wire w_dff_A_K7gMtYAm4_0;
	wire w_dff_A_CmsjPF7W1_0;
	wire w_dff_A_nSZOk3yf3_0;
	wire w_dff_A_UyjAO2PB8_0;
	wire w_dff_A_Q0WTtCKU1_0;
	wire w_dff_A_gojJTxL90_0;
	wire w_dff_A_nDKChvTu5_0;
	wire w_dff_A_InsADXP52_0;
	wire w_dff_A_451P4qkv5_0;
	wire w_dff_A_teEmgDa31_0;
	wire w_dff_A_hW8ZtUsF5_0;
	wire w_dff_A_LCfGoxfb7_0;
	wire w_dff_A_L0Hj4WZc1_0;
	wire w_dff_A_gZ1R2zXt6_0;
	wire w_dff_A_x0XWrMoh0_0;
	wire w_dff_A_ICDD4oHo3_0;
	wire w_dff_A_vmsaB1HH5_0;
	wire w_dff_A_9mqdupKU3_0;
	wire w_dff_A_X0974R2u0_0;
	wire w_dff_A_6CNYcLKx3_0;
	wire w_dff_A_NCqyXU4Z2_0;
	wire w_dff_A_PUluDnQW3_0;
	wire w_dff_A_hQwWJGOh7_0;
	wire w_dff_A_xXVYilAv6_0;
	wire w_dff_A_kNbKvpbM7_0;
	wire w_dff_A_7kDqg9E90_2;
	wire w_dff_A_w1v5wgod7_0;
	wire w_dff_A_mrqQ34YW0_0;
	wire w_dff_A_peT6RoWX1_0;
	wire w_dff_A_zrYxOMZs0_0;
	wire w_dff_A_UIquMr658_0;
	wire w_dff_A_dAcENKSM7_0;
	wire w_dff_A_6pyLv7aY9_0;
	wire w_dff_A_4GRSAY1B4_0;
	wire w_dff_A_z7q2J3wv7_0;
	wire w_dff_A_Trh8OoQS0_0;
	wire w_dff_A_yF9MVNaO4_0;
	wire w_dff_A_arc6ByMn9_0;
	wire w_dff_A_bq6j5ewq2_0;
	wire w_dff_A_Yg9vO6lc4_0;
	wire w_dff_A_L7wIM2tI9_0;
	wire w_dff_A_megLYJw99_0;
	wire w_dff_A_c3stksiv6_0;
	wire w_dff_A_eioubO7q2_0;
	wire w_dff_A_iEdmvH551_0;
	wire w_dff_A_nltm93702_0;
	wire w_dff_A_P9jat2O28_0;
	wire w_dff_A_NpNc9lKT6_0;
	wire w_dff_A_lkLePOwx5_0;
	wire w_dff_A_KtzlBNsZ5_0;
	wire w_dff_A_Ozaj3MJi7_0;
	wire w_dff_A_r3xfQC3E5_0;
	wire w_dff_A_UELLSaGU0_0;
	wire w_dff_A_ORLJKkOG4_0;
	wire w_dff_A_HPk4UVUJ8_0;
	wire w_dff_A_qrccpb3i0_0;
	wire w_dff_A_bvv7RRTT7_0;
	wire w_dff_A_G6Ijt2045_0;
	wire w_dff_A_ZZeqKtMi4_0;
	wire w_dff_A_s2C7haa13_0;
	wire w_dff_A_oAeOVQOF6_0;
	wire w_dff_A_VDrkGpMV2_0;
	wire w_dff_A_oKzz53IO5_2;
	wire w_dff_A_lyJ8Fdoz1_0;
	wire w_dff_A_1xJrJYEB8_0;
	wire w_dff_A_xyQ40gwT1_0;
	wire w_dff_A_aI10CsNS8_0;
	wire w_dff_A_XWcZECy74_0;
	wire w_dff_A_Cys1BEmO3_0;
	wire w_dff_A_yZiay1Ra5_0;
	wire w_dff_A_CQcn7UCA4_0;
	wire w_dff_A_RXthB2Mn2_0;
	wire w_dff_A_IJfONVh88_0;
	wire w_dff_A_IdEcnlQK2_0;
	wire w_dff_A_tRJZPFQj6_0;
	wire w_dff_A_1NU2Sj192_0;
	wire w_dff_A_6NWdFAQ88_0;
	wire w_dff_A_6VZCquiV0_0;
	wire w_dff_A_2Atwsl1e8_0;
	wire w_dff_A_h7JwT59k0_0;
	wire w_dff_A_1eHLkgSZ4_0;
	wire w_dff_A_iKWKqtI07_0;
	wire w_dff_A_9jX8atez9_0;
	wire w_dff_A_x99zwbsx6_0;
	wire w_dff_A_XGMUizW88_0;
	wire w_dff_A_NgRQ9sQv0_0;
	wire w_dff_A_YdYiZ7AU3_0;
	wire w_dff_A_VJQGOMM76_0;
	wire w_dff_A_T7Z2gSsz2_0;
	wire w_dff_A_YTdbOB5J2_0;
	wire w_dff_A_MRXlh1625_0;
	wire w_dff_A_dnbNaOuy9_0;
	wire w_dff_A_5193G9Ww8_0;
	wire w_dff_A_5uSi0a8m7_0;
	wire w_dff_A_SrWgg1V45_0;
	wire w_dff_A_5J7euuBr6_0;
	wire w_dff_A_G5dtKGF12_0;
	wire w_dff_A_I4pNf0av5_0;
	wire w_dff_A_AEzxCK512_2;
	wire w_dff_A_GG2qHrda8_0;
	wire w_dff_A_HEMTRrbP5_0;
	wire w_dff_A_pmoD3Ghc4_0;
	wire w_dff_A_36qEBrI93_0;
	wire w_dff_A_9zlPCw3b3_0;
	wire w_dff_A_DjsrlyfB3_0;
	wire w_dff_A_ZKoYZQew1_0;
	wire w_dff_A_O0lCVhFz5_0;
	wire w_dff_A_7ZLbmI1O3_0;
	wire w_dff_A_2ZrH3l2z6_0;
	wire w_dff_A_y4bBXwF59_0;
	wire w_dff_A_5EqS5cp89_0;
	wire w_dff_A_pqyHQPTf7_0;
	wire w_dff_A_ZGXGSGaI8_0;
	wire w_dff_A_kk8aeY6D9_0;
	wire w_dff_A_Ym6T1lWP5_0;
	wire w_dff_A_GMReuTzS9_0;
	wire w_dff_A_xCHzNYns4_0;
	wire w_dff_A_Y0viZO0d2_0;
	wire w_dff_A_PGTCaPkD5_0;
	wire w_dff_A_FR07CoQ79_0;
	wire w_dff_A_tRN7QY4J8_0;
	wire w_dff_A_sOqrwEUk5_0;
	wire w_dff_A_FEnRIYzi5_0;
	wire w_dff_A_gVW96HaF4_0;
	wire w_dff_A_3VGk58dE0_0;
	wire w_dff_A_KSIjEYaI7_0;
	wire w_dff_A_uAg23j1w9_0;
	wire w_dff_A_4Q9byydA5_0;
	wire w_dff_A_2vk2danU6_0;
	wire w_dff_A_xFJkBUed9_0;
	wire w_dff_A_bTMQQsJo4_0;
	wire w_dff_A_gfT7eHZK6_0;
	wire w_dff_A_ha7sRvCT7_0;
	wire w_dff_A_Er2L8DHW9_2;
	wire w_dff_A_s0FhXH485_0;
	wire w_dff_A_H3KxTAOp2_0;
	wire w_dff_A_q4vYkGNi5_0;
	wire w_dff_A_27hEjulX3_0;
	wire w_dff_A_tm4LvgA97_0;
	wire w_dff_A_LcTWEY0y3_0;
	wire w_dff_A_dhjZMPjj6_0;
	wire w_dff_A_nAhy8jg97_0;
	wire w_dff_A_iZ0FBQ177_0;
	wire w_dff_A_C74O2baP2_0;
	wire w_dff_A_gurycyko8_0;
	wire w_dff_A_5hlrvbOy0_0;
	wire w_dff_A_HLpD1Wbu2_0;
	wire w_dff_A_wFI9jBks7_0;
	wire w_dff_A_jVyFTlLG6_0;
	wire w_dff_A_mVbs1mQK4_0;
	wire w_dff_A_QlmCQiEH4_0;
	wire w_dff_A_L6KSNkEp9_0;
	wire w_dff_A_j7CXxbfw8_0;
	wire w_dff_A_ZtrqJAz43_0;
	wire w_dff_A_RsvUncEq5_0;
	wire w_dff_A_0pkwwZBt8_0;
	wire w_dff_A_VpJKZxxq4_0;
	wire w_dff_A_c7ULtHPb4_0;
	wire w_dff_A_J6zzYJr99_0;
	wire w_dff_A_fEDCAqdp5_0;
	wire w_dff_A_jJz3Byz79_0;
	wire w_dff_A_6ccVvoid0_0;
	wire w_dff_A_xNjEQSO61_0;
	wire w_dff_A_uLE9o1bl6_0;
	wire w_dff_A_OeLNR1lA4_0;
	wire w_dff_A_yQAACRrt1_0;
	wire w_dff_A_GteC1O896_0;
	wire w_dff_A_XtJDEDOj6_2;
	wire w_dff_A_OyFx5A880_0;
	wire w_dff_A_KOaYgp0D9_0;
	wire w_dff_A_nkgGLMtD9_0;
	wire w_dff_A_IaiFbMsq2_0;
	wire w_dff_A_hiH3E2K55_0;
	wire w_dff_A_nFdgBBVX7_0;
	wire w_dff_A_f7KippQH5_0;
	wire w_dff_A_jZCayZcU5_0;
	wire w_dff_A_EnygtvhL5_0;
	wire w_dff_A_pTJ5ZJAZ3_0;
	wire w_dff_A_V6FZ53R40_0;
	wire w_dff_A_g6SGFTmx0_0;
	wire w_dff_A_wv7Zd7jA2_0;
	wire w_dff_A_0DkXz5Rp1_0;
	wire w_dff_A_R4ehAkps4_0;
	wire w_dff_A_wHPL78TD7_0;
	wire w_dff_A_wjbkuumn2_0;
	wire w_dff_A_87Lomuc35_0;
	wire w_dff_A_TemNoxqc6_0;
	wire w_dff_A_6feuHVrJ0_0;
	wire w_dff_A_0G0vAa8i2_0;
	wire w_dff_A_AHCT5n9d5_0;
	wire w_dff_A_mTbdqkSx3_0;
	wire w_dff_A_nrZDo8Ng2_0;
	wire w_dff_A_ftSEOCsG1_0;
	wire w_dff_A_FNAR7OHg0_0;
	wire w_dff_A_i2sXLfoG6_0;
	wire w_dff_A_Ib8X9Dm93_0;
	wire w_dff_A_4iLw99K71_0;
	wire w_dff_A_HOt6GUvs5_0;
	wire w_dff_A_3NTiZ3Yi6_0;
	wire w_dff_A_RFD5YmZp0_0;
	wire w_dff_A_AMFRU9o10_2;
	wire w_dff_A_jIVhXD069_0;
	wire w_dff_A_yTp6qN5W8_0;
	wire w_dff_A_1zUFLRwG2_0;
	wire w_dff_A_VwrrkvWe2_0;
	wire w_dff_A_sfB2jh6E7_0;
	wire w_dff_A_CBgQENVl6_0;
	wire w_dff_A_5sg1HbME6_0;
	wire w_dff_A_x8ExOody9_0;
	wire w_dff_A_21NfC90x9_0;
	wire w_dff_A_qfCcvu7Y4_0;
	wire w_dff_A_c6jxBjna5_0;
	wire w_dff_A_iGWbQu3n5_0;
	wire w_dff_A_FmNSV9Zc5_0;
	wire w_dff_A_pzOzmHdQ2_0;
	wire w_dff_A_OEUCuBTl8_0;
	wire w_dff_A_wkWBZRef1_0;
	wire w_dff_A_Fdfb4myi2_0;
	wire w_dff_A_xBzxjasY5_0;
	wire w_dff_A_K9CmqhHe0_0;
	wire w_dff_A_mVI6TKSg5_0;
	wire w_dff_A_REjKV5va8_0;
	wire w_dff_A_gIuKOqEl3_0;
	wire w_dff_A_Z2OHPcQM9_0;
	wire w_dff_A_exWGyCCJ8_0;
	wire w_dff_A_0CUD4K4l6_0;
	wire w_dff_A_Pb8O3KwZ2_0;
	wire w_dff_A_9bxlpSS61_0;
	wire w_dff_A_CCJJUVgd2_0;
	wire w_dff_A_2Xvt5aW23_0;
	wire w_dff_A_ZOVD3b5g5_0;
	wire w_dff_A_TlgeE8eC6_0;
	wire w_dff_A_4HZtpbSH1_2;
	wire w_dff_A_OzbBedJb7_0;
	wire w_dff_A_1MTZhLHc1_0;
	wire w_dff_A_ne1HhVGo4_0;
	wire w_dff_A_9qr5Z93a6_0;
	wire w_dff_A_RjQ5wP8l1_0;
	wire w_dff_A_4wBtinSQ2_0;
	wire w_dff_A_8OhVbW7t9_0;
	wire w_dff_A_x0TcEQ1t1_0;
	wire w_dff_A_E17ZPpId0_0;
	wire w_dff_A_T6bTbsre6_0;
	wire w_dff_A_m5mqXB9Y0_0;
	wire w_dff_A_QtfUI3C00_0;
	wire w_dff_A_TF6lvV6v0_0;
	wire w_dff_A_WUOT6sek2_0;
	wire w_dff_A_Cvgxm6IG7_0;
	wire w_dff_A_lC7hgAga4_0;
	wire w_dff_A_dqssucrA4_0;
	wire w_dff_A_h5Ade49L3_0;
	wire w_dff_A_bllbTu639_0;
	wire w_dff_A_WPcbLUlv7_0;
	wire w_dff_A_WezhJCRD5_0;
	wire w_dff_A_TPZG4tmn1_0;
	wire w_dff_A_AH40itoX9_0;
	wire w_dff_A_FbErS4Kj5_0;
	wire w_dff_A_oEym1vmV9_0;
	wire w_dff_A_wOnsUkqY4_0;
	wire w_dff_A_U8Ri4lTr6_0;
	wire w_dff_A_5ToOps0K2_0;
	wire w_dff_A_A1O5LbtV9_0;
	wire w_dff_A_5SZGfYla9_0;
	wire w_dff_A_LhBO705X1_2;
	wire w_dff_A_zEpGsihP7_0;
	wire w_dff_A_WRML9YSR7_0;
	wire w_dff_A_EbMEZZh34_0;
	wire w_dff_A_Jv1ane812_0;
	wire w_dff_A_0NHjkmcn2_0;
	wire w_dff_A_S8x0eCf48_0;
	wire w_dff_A_m7EI7u6d7_0;
	wire w_dff_A_0kqtpuMh4_0;
	wire w_dff_A_YOIchtsx3_0;
	wire w_dff_A_RJ6aH9HW3_0;
	wire w_dff_A_ykMiWOmd7_0;
	wire w_dff_A_r9vIpNX69_0;
	wire w_dff_A_zdj4RMZp5_0;
	wire w_dff_A_Uz5G1Hr18_0;
	wire w_dff_A_BvBDuFQC5_0;
	wire w_dff_A_H1k3tpQC5_0;
	wire w_dff_A_NR8wCoVQ3_0;
	wire w_dff_A_SOJoO6kf2_0;
	wire w_dff_A_w2pwQ2km1_0;
	wire w_dff_A_iKLN3hkd6_0;
	wire w_dff_A_oYLQsRHv3_0;
	wire w_dff_A_uL5O8sbb5_0;
	wire w_dff_A_Aurm1clF5_0;
	wire w_dff_A_mUpL9pL13_0;
	wire w_dff_A_RrdZ3eil9_0;
	wire w_dff_A_cseoMQNJ7_0;
	wire w_dff_A_tllxPUpK9_0;
	wire w_dff_A_AWDRmoyb0_0;
	wire w_dff_A_re7SjTjq8_0;
	wire w_dff_A_rQuWRbM25_2;
	wire w_dff_A_sAQW3IEU1_0;
	wire w_dff_A_p3eE2AWL6_0;
	wire w_dff_A_BMLHg5pi6_0;
	wire w_dff_A_3LVBQ0Pl4_0;
	wire w_dff_A_Dotap0Un6_0;
	wire w_dff_A_1AchSSIF2_0;
	wire w_dff_A_3f3b0Iid8_0;
	wire w_dff_A_7QRDJune4_0;
	wire w_dff_A_82QO3kuO9_0;
	wire w_dff_A_5NcD73wh4_0;
	wire w_dff_A_hY5JxQdx9_0;
	wire w_dff_A_trFWKzSG7_0;
	wire w_dff_A_TCrAfWY33_0;
	wire w_dff_A_Y5x0x0nm7_0;
	wire w_dff_A_QNGsPW584_0;
	wire w_dff_A_LoSkd3Sz7_0;
	wire w_dff_A_BWZex2k27_0;
	wire w_dff_A_ho1eOfeC8_0;
	wire w_dff_A_qd6suzrS7_0;
	wire w_dff_A_Jw6s70ey5_0;
	wire w_dff_A_cDA7P9sQ0_0;
	wire w_dff_A_ZUoVrhUy8_0;
	wire w_dff_A_WYcXydrp6_0;
	wire w_dff_A_UqF2f45e4_0;
	wire w_dff_A_052u7nYm7_0;
	wire w_dff_A_m1kegvqW0_0;
	wire w_dff_A_XYL7coZp0_0;
	wire w_dff_A_xdsG2och5_0;
	wire w_dff_A_jth7tJDE4_2;
	wire w_dff_A_V1dGsCCM7_0;
	wire w_dff_A_oqpsioch9_0;
	wire w_dff_A_FBvVIzWY2_0;
	wire w_dff_A_xbRA5X9p5_0;
	wire w_dff_A_Nm9K2iCn4_0;
	wire w_dff_A_609eHOsQ7_0;
	wire w_dff_A_LmHUcl7l8_0;
	wire w_dff_A_vR2hI2l76_0;
	wire w_dff_A_SDchV6BP6_0;
	wire w_dff_A_4RXx2lW24_0;
	wire w_dff_A_XC6hkmqM3_0;
	wire w_dff_A_DU5JkoUh6_0;
	wire w_dff_A_f7dD0e0w5_0;
	wire w_dff_A_kdfSSpBn7_0;
	wire w_dff_A_X07Dzd4B8_0;
	wire w_dff_A_TjyJTRN73_0;
	wire w_dff_A_T9LIP4ij6_0;
	wire w_dff_A_dCuIuUfN1_0;
	wire w_dff_A_2yIgaWsg8_0;
	wire w_dff_A_Ulvsk4vP0_0;
	wire w_dff_A_iheEw9AN7_0;
	wire w_dff_A_63E4zvyf8_0;
	wire w_dff_A_vBRWUc9B3_0;
	wire w_dff_A_XHOBbnYp9_0;
	wire w_dff_A_JQxkL62B2_0;
	wire w_dff_A_lMcdKPRB3_0;
	wire w_dff_A_slMcurW44_0;
	wire w_dff_A_vGnqaJJF9_2;
	wire w_dff_A_TUq5Ubjf5_0;
	wire w_dff_A_EPglFiZF0_0;
	wire w_dff_A_27Pf443e7_0;
	wire w_dff_A_CkokMeok2_0;
	wire w_dff_A_8zeaxkIn2_0;
	wire w_dff_A_u82QWup05_0;
	wire w_dff_A_gYo2DAND4_0;
	wire w_dff_A_fW51Of138_0;
	wire w_dff_A_v4W7ykMc4_0;
	wire w_dff_A_wZ7I0XZw5_0;
	wire w_dff_A_slYO8GMn1_0;
	wire w_dff_A_Bw7GPftn7_0;
	wire w_dff_A_UT8Tuj5l2_0;
	wire w_dff_A_nGZowy1a8_0;
	wire w_dff_A_JlqjK21E7_0;
	wire w_dff_A_Tx7FWKCP1_0;
	wire w_dff_A_UZ2YTpHk2_0;
	wire w_dff_A_ZXyfIqhh9_0;
	wire w_dff_A_OKIpevN61_0;
	wire w_dff_A_epiqUJjz6_0;
	wire w_dff_A_ME0a4nPr3_0;
	wire w_dff_A_zhnxk0Qq3_0;
	wire w_dff_A_2cpCqytp7_0;
	wire w_dff_A_k487bRJE0_0;
	wire w_dff_A_L5DA1Ew38_0;
	wire w_dff_A_ZN5Pv19v0_0;
	wire w_dff_A_Fj4n1Rkq2_2;
	wire w_dff_A_hXEtOOHJ7_0;
	wire w_dff_A_zPYaZlJv0_0;
	wire w_dff_A_lsstklFy5_0;
	wire w_dff_A_okMKNz337_0;
	wire w_dff_A_1sX6YB4P5_0;
	wire w_dff_A_VB2xGp2w5_0;
	wire w_dff_A_TB8mrGKu0_0;
	wire w_dff_A_6gMvx1hS4_0;
	wire w_dff_A_ntZFqKDd6_0;
	wire w_dff_A_7N4kp3X63_0;
	wire w_dff_A_bqWsk6JH0_0;
	wire w_dff_A_TYQY54Mp1_0;
	wire w_dff_A_BHPBXFJe8_0;
	wire w_dff_A_jQ0eDOjk2_0;
	wire w_dff_A_IqT8IT6l2_0;
	wire w_dff_A_cCgJvPcb8_0;
	wire w_dff_A_eovcZIHQ7_0;
	wire w_dff_A_zEDwgM0L5_0;
	wire w_dff_A_fsnrjpag8_0;
	wire w_dff_A_ST5L3gf98_0;
	wire w_dff_A_opiUc1bh3_0;
	wire w_dff_A_xl2jBpz60_0;
	wire w_dff_A_EAyseYti3_0;
	wire w_dff_A_k7kRvua23_0;
	wire w_dff_A_LEtvUaOA7_0;
	wire w_dff_A_P3vaBdYA9_2;
	wire w_dff_A_wgW0wQKP7_0;
	wire w_dff_A_TEShzEva1_0;
	wire w_dff_A_kWujKEim4_0;
	wire w_dff_A_VmhHHbww9_0;
	wire w_dff_A_JCso0TM61_0;
	wire w_dff_A_mlH8pfmY3_0;
	wire w_dff_A_y31upuPF3_0;
	wire w_dff_A_WQ5oT3ZY3_0;
	wire w_dff_A_Utd4LhlA5_0;
	wire w_dff_A_LUFoTsyR0_0;
	wire w_dff_A_7BlsdwCI3_0;
	wire w_dff_A_5JG3KtDt2_0;
	wire w_dff_A_RYwAcxiH3_0;
	wire w_dff_A_WpCQYC4I6_0;
	wire w_dff_A_fbgpJ23L3_0;
	wire w_dff_A_C0MY41l90_0;
	wire w_dff_A_dtC4Y41o0_0;
	wire w_dff_A_ztH5nZhI4_0;
	wire w_dff_A_XJ4vC2Ol1_0;
	wire w_dff_A_hTSzYaC67_0;
	wire w_dff_A_NI4DIGyU8_0;
	wire w_dff_A_7QVvKskS0_0;
	wire w_dff_A_POMwUXZ06_0;
	wire w_dff_A_mGf3FJTz7_0;
	wire w_dff_A_XMlybQoI8_2;
	wire w_dff_A_DnPGD6s15_0;
	wire w_dff_A_aLqdgAdc8_0;
	wire w_dff_A_VsMcGbNA4_0;
	wire w_dff_A_RRDLnXg30_0;
	wire w_dff_A_0RLeMwV01_0;
	wire w_dff_A_SplXach55_0;
	wire w_dff_A_Rup4IS1v6_0;
	wire w_dff_A_DUpeHa601_0;
	wire w_dff_A_gGBdJpjh0_0;
	wire w_dff_A_Dq5ar8i42_0;
	wire w_dff_A_wlDihNJk4_0;
	wire w_dff_A_qSm3hOd71_0;
	wire w_dff_A_nJg4aDGr2_0;
	wire w_dff_A_TfuZ4JPa7_0;
	wire w_dff_A_vxsUmO9G3_0;
	wire w_dff_A_y60o0Nyw9_0;
	wire w_dff_A_keigOqtW6_0;
	wire w_dff_A_G2nbdawe5_0;
	wire w_dff_A_y1NYJzuH5_0;
	wire w_dff_A_N54wXrV99_0;
	wire w_dff_A_UFL3lFAj9_0;
	wire w_dff_A_MYRBxoZT7_0;
	wire w_dff_A_vcPCwn541_0;
	wire w_dff_A_5ieeOtHr7_2;
	wire w_dff_A_zoSumTK41_0;
	wire w_dff_A_djrT8tsr0_0;
	wire w_dff_A_SW1g5nM00_0;
	wire w_dff_A_cMwlRTG65_0;
	wire w_dff_A_zzmi3HH02_0;
	wire w_dff_A_QMOoHHeL5_0;
	wire w_dff_A_gLMsXJs80_0;
	wire w_dff_A_d3b9AFFd2_0;
	wire w_dff_A_MqDIMbQG9_0;
	wire w_dff_A_xLkATVKT3_0;
	wire w_dff_A_iX2EXJGN3_0;
	wire w_dff_A_4Hojidmt9_0;
	wire w_dff_A_YiNWJ4kD9_0;
	wire w_dff_A_SxbIkGKd3_0;
	wire w_dff_A_hFFa02gQ4_0;
	wire w_dff_A_4SZg7hkt0_0;
	wire w_dff_A_2YGmEzHA8_0;
	wire w_dff_A_fbLZO0UM7_0;
	wire w_dff_A_H8mMMVgf0_0;
	wire w_dff_A_pI0NoPbT6_0;
	wire w_dff_A_MRXsOHl51_0;
	wire w_dff_A_dX5aVNW90_0;
	wire w_dff_A_ZOM6W9LV4_2;
	wire w_dff_A_mIgwi5UL9_0;
	wire w_dff_A_XFpw9E6u2_0;
	wire w_dff_A_NZF4uEZs0_0;
	wire w_dff_A_MYFDGeFq7_0;
	wire w_dff_A_0hvkPZNW7_0;
	wire w_dff_A_XyHIVfkr3_0;
	wire w_dff_A_cERMalAW1_0;
	wire w_dff_A_maQDEzpY8_0;
	wire w_dff_A_CkOgGDVh6_0;
	wire w_dff_A_hRrtdQzl4_0;
	wire w_dff_A_VhbgBBqp3_0;
	wire w_dff_A_kKmAAYk10_0;
	wire w_dff_A_Rf5lOyIV9_0;
	wire w_dff_A_HeTMY7S33_0;
	wire w_dff_A_sMpvmZLb5_0;
	wire w_dff_A_pBeQ16zq6_0;
	wire w_dff_A_k96B1frD7_0;
	wire w_dff_A_sKaCFLvi4_0;
	wire w_dff_A_JaihCoN39_0;
	wire w_dff_A_OERwHGfQ5_0;
	wire w_dff_A_6Yj68FtL3_0;
	wire w_dff_A_URhuMiJa9_2;
	wire w_dff_A_R5xOR7iw0_0;
	wire w_dff_A_AcrXoWmU0_0;
	wire w_dff_A_WIV82wZ56_0;
	wire w_dff_A_mql5OtEv4_0;
	wire w_dff_A_X14564wG4_0;
	wire w_dff_A_HRLznOIr3_0;
	wire w_dff_A_83FIooh79_0;
	wire w_dff_A_eYcdS94q2_0;
	wire w_dff_A_x0Qy0WX98_0;
	wire w_dff_A_KyRbk5do0_0;
	wire w_dff_A_gXpRIzGV1_0;
	wire w_dff_A_uFwR1n136_0;
	wire w_dff_A_Au45byRy8_0;
	wire w_dff_A_J7dGG6DA3_0;
	wire w_dff_A_yzi3vWZX4_0;
	wire w_dff_A_HVvuYU7h3_0;
	wire w_dff_A_ZuuRcs2H9_0;
	wire w_dff_A_HPNQdwgI4_0;
	wire w_dff_A_1icJqdb29_0;
	wire w_dff_A_3Lo9b6G18_0;
	wire w_dff_A_cwkY2DxV9_2;
	wire w_dff_A_QvqEaHKG4_0;
	wire w_dff_A_EjyZ383l8_0;
	wire w_dff_A_JVRc0Ru27_0;
	wire w_dff_A_Wjpi3EFy3_0;
	wire w_dff_A_svbN2EnZ7_0;
	wire w_dff_A_uq6gKeGI7_0;
	wire w_dff_A_1NPtqsrc0_0;
	wire w_dff_A_Q0YMngAh6_0;
	wire w_dff_A_IeCXc6Qg3_0;
	wire w_dff_A_64UkebS74_0;
	wire w_dff_A_d2IRJ8AP8_0;
	wire w_dff_A_nklNoIf45_0;
	wire w_dff_A_DZ28DWka4_0;
	wire w_dff_A_rdmNDJLK3_0;
	wire w_dff_A_ySSQOess4_0;
	wire w_dff_A_7eqsieVT7_0;
	wire w_dff_A_oGHixy531_0;
	wire w_dff_A_e0xhZWKO7_0;
	wire w_dff_A_0TBOmsVl5_0;
	wire w_dff_A_aQI6d3Nn2_2;
	wire w_dff_A_AzNc77CQ7_0;
	wire w_dff_A_LCM4Yejg9_0;
	wire w_dff_A_uIPLGUNv6_0;
	wire w_dff_A_YCe56c4y2_0;
	wire w_dff_A_eLLA1vKa2_0;
	wire w_dff_A_1uwtFH7b0_0;
	wire w_dff_A_zMgjeUZL0_0;
	wire w_dff_A_CMUE9ayB0_0;
	wire w_dff_A_ktuva36K9_0;
	wire w_dff_A_FyeagAyb5_0;
	wire w_dff_A_9QuLYpSU7_0;
	wire w_dff_A_I9774roP9_0;
	wire w_dff_A_woYQbONg7_0;
	wire w_dff_A_aW0JcCXM5_0;
	wire w_dff_A_7jZtU57U6_0;
	wire w_dff_A_y0zwjRrI2_0;
	wire w_dff_A_IDNxqPEX8_0;
	wire w_dff_A_QovH0nhy8_0;
	wire w_dff_A_6RAzsJrE3_2;
	wire w_dff_A_fcPJaCHr9_0;
	wire w_dff_A_Pt75JKha0_0;
	wire w_dff_A_pDrdtPCf8_0;
	wire w_dff_A_9sOSToaq3_0;
	wire w_dff_A_tats9DAT7_0;
	wire w_dff_A_xVMTakRC2_0;
	wire w_dff_A_U5svZFhj4_0;
	wire w_dff_A_qYmj0XIQ6_0;
	wire w_dff_A_j4BASZgP3_0;
	wire w_dff_A_FtrYgpAU5_0;
	wire w_dff_A_LssIE8tW7_0;
	wire w_dff_A_D23S3ID22_0;
	wire w_dff_A_6fgPjKce4_0;
	wire w_dff_A_ZSQ4I4Ui4_0;
	wire w_dff_A_jY6jEer21_0;
	wire w_dff_A_R2MXtO1e0_0;
	wire w_dff_A_apYP00tx6_0;
	wire w_dff_A_ukMTbJQ36_2;
	wire w_dff_A_wvEQ7hdg0_0;
	wire w_dff_A_VU1EFMrT3_0;
	wire w_dff_A_ZNqCzFb72_0;
	wire w_dff_A_83vQJNTY9_0;
	wire w_dff_A_Mtznnj0x6_0;
	wire w_dff_A_VFIf5r337_0;
	wire w_dff_A_yxJPLhbU3_0;
	wire w_dff_A_LKgLger15_0;
	wire w_dff_A_poO4AJMA0_0;
	wire w_dff_A_8Tl9X62H9_0;
	wire w_dff_A_4Abr1N4q3_0;
	wire w_dff_A_z9ixAAkq1_0;
	wire w_dff_A_ytJE0TKo5_0;
	wire w_dff_A_cmvhdiwe7_0;
	wire w_dff_A_bqz4TNf24_0;
	wire w_dff_A_stwvBZNp3_0;
	wire w_dff_A_kWw534XR3_2;
	wire w_dff_A_BidquCIy1_0;
	wire w_dff_A_VarZBo5k7_0;
	wire w_dff_A_bKn9TE068_0;
	wire w_dff_A_awMKTcC25_0;
	wire w_dff_A_dTG30o3B6_0;
	wire w_dff_A_Ly0DCpf35_0;
	wire w_dff_A_TcdsbM6c6_0;
	wire w_dff_A_lPHYUwfF7_0;
	wire w_dff_A_1C4UwDMw2_0;
	wire w_dff_A_wA3cx3SH3_0;
	wire w_dff_A_VYIjAtFW9_0;
	wire w_dff_A_7amHe4Bo5_0;
	wire w_dff_A_M6xb7lpj5_0;
	wire w_dff_A_tSKYmCYO7_0;
	wire w_dff_A_bHjWloGN6_0;
	wire w_dff_A_bne51yCD0_2;
	wire w_dff_A_WK6EJDtf0_0;
	wire w_dff_A_ClhUFvES4_0;
	wire w_dff_A_zqNRi1lD4_0;
	wire w_dff_A_FfOHGaCs6_0;
	wire w_dff_A_qvxSnGmK1_0;
	wire w_dff_A_BtXzz1kR5_0;
	wire w_dff_A_QIUA7GFY1_0;
	wire w_dff_A_jzqemet56_0;
	wire w_dff_A_IBAGth7O9_0;
	wire w_dff_A_B095ri797_0;
	wire w_dff_A_n2L41IjT2_0;
	wire w_dff_A_XagthY0s2_0;
	wire w_dff_A_Am07XMav3_0;
	wire w_dff_A_co00XfWT4_0;
	wire w_dff_A_3U7JlSNO5_2;
	wire w_dff_A_pnLvFod86_0;
	wire w_dff_A_aY6E5eNv5_0;
	wire w_dff_A_Y9gpwtXe4_0;
	wire w_dff_A_azWlgLyn6_0;
	wire w_dff_A_Usu1l2Kb3_0;
	wire w_dff_A_WtFxGp7T6_0;
	wire w_dff_A_AKHwbQAN1_0;
	wire w_dff_A_MfGW3Onq8_0;
	wire w_dff_A_C1MbJwYK1_0;
	wire w_dff_A_mBejUqLh8_0;
	wire w_dff_A_7LEqFVeF4_0;
	wire w_dff_A_deTQa9lE0_0;
	wire w_dff_A_fKhiDbuw8_0;
	wire w_dff_A_3VmB04UB2_2;
	wire w_dff_A_HaTQCZom3_0;
	wire w_dff_A_qzCNFlmB7_0;
	wire w_dff_A_dcPacLFt4_0;
	wire w_dff_A_HaXPQeVw0_0;
	wire w_dff_A_QHBz4jk01_0;
	wire w_dff_A_rR5VlmdJ0_0;
	wire w_dff_A_rkgx6CZI6_0;
	wire w_dff_A_ZOBgwSoD9_0;
	wire w_dff_A_qpir5nay3_0;
	wire w_dff_A_o1t3YtAy4_0;
	wire w_dff_A_ejOVAiHG2_0;
	wire w_dff_A_7RRxYpKw9_0;
	wire w_dff_A_3bA8xD5P2_2;
	wire w_dff_A_vSSzQQdW7_0;
	wire w_dff_A_M2OmrYFS7_0;
	wire w_dff_A_cZL1uRaJ3_0;
	wire w_dff_A_9yJbI2Ln9_0;
	wire w_dff_A_eSducORv0_0;
	wire w_dff_A_Pv6XwFBY6_0;
	wire w_dff_A_CLQlnbdo5_0;
	wire w_dff_A_1oBmfopY1_0;
	wire w_dff_A_FbUW3vO70_0;
	wire w_dff_A_p6zFibIm6_0;
	wire w_dff_A_8uaIeREO3_0;
	wire w_dff_A_fKN0jFwO9_2;
	wire w_dff_A_7XAfmi9u6_0;
	wire w_dff_A_OlFkYmOn2_0;
	wire w_dff_A_KCwq0QBL8_0;
	wire w_dff_A_Iz7WlUZf0_0;
	wire w_dff_A_WCk5HKwe4_0;
	wire w_dff_A_Xv5Trcx60_0;
	wire w_dff_A_SBEmuX9o8_0;
	wire w_dff_A_8dYujpQX8_0;
	wire w_dff_A_4mHypyvg4_0;
	wire w_dff_A_LBRWsrIM0_0;
	wire w_dff_A_llLQJvtS3_2;
	wire w_dff_A_xrBJtCSZ0_0;
	wire w_dff_A_UK5NQipZ2_0;
	wire w_dff_A_7JQOCkeH0_0;
	wire w_dff_A_okE5sMLk3_0;
	wire w_dff_A_mYpIoqg69_0;
	wire w_dff_A_tCCFH3Xv7_0;
	wire w_dff_A_jPfqylYA2_0;
	wire w_dff_A_zBR8Aika4_0;
	wire w_dff_A_EcfhzWiX4_0;
	wire w_dff_A_9UxeUz0e4_2;
	wire w_dff_A_ZTGYclPq4_0;
	wire w_dff_A_U7yMt1zL1_0;
	wire w_dff_A_7PxYVrBw0_0;
	wire w_dff_A_Ymx8UBmT3_0;
	wire w_dff_A_yXYCHHPO8_0;
	wire w_dff_A_JaAJ4YBp6_0;
	wire w_dff_A_gL7u1HKB1_0;
	wire w_dff_A_SaestAav7_0;
	wire w_dff_A_VEKg84Oy2_2;
	wire w_dff_A_tY6J68k74_0;
	wire w_dff_A_AasODOBE5_0;
	wire w_dff_A_7jrMCY5F3_0;
	wire w_dff_A_B81ZmGIY8_0;
	wire w_dff_A_lVdqU8uU9_0;
	wire w_dff_A_r4Mbs7zM4_0;
	wire w_dff_A_16l6xVEV2_0;
	wire w_dff_A_qLw4TMU81_2;
	wire w_dff_A_gQUcPB1M3_0;
	wire w_dff_A_gXUcJs2c8_0;
	wire w_dff_A_wFBaKcoN0_0;
	wire w_dff_A_7ieWQnUJ4_0;
	wire w_dff_A_YydnO40Y0_0;
	wire w_dff_A_l8FPsNhz8_0;
	wire w_dff_A_72ECXwuX6_2;
	wire w_dff_A_6fdH6ibw7_0;
	wire w_dff_A_V9DHNrXJ1_0;
	wire w_dff_A_YAN9LuKi3_0;
	wire w_dff_A_DIG7appW3_0;
	wire w_dff_A_l7fEUm0g5_0;
	wire w_dff_A_pUdZQfwk6_2;
	wire w_dff_A_SYV3Wbhr8_0;
	wire w_dff_A_c3di3RzO0_0;
	wire w_dff_A_HlzORNQm3_0;
	wire w_dff_A_rPEjnIGK4_0;
	wire w_dff_A_njEGwhT63_2;
	wire w_dff_A_nDWIoLhN5_0;
	wire w_dff_A_YOPuAJXX3_0;
	wire w_dff_A_YgokwFm35_0;
	wire w_dff_A_qPETohS16_2;
	wire w_dff_A_YWhCSTZH9_0;
	wire w_dff_A_Xe9XK3yk0_0;
	wire w_dff_A_Dk9V03BL7_2;
	wire w_dff_A_QYfAqV0p5_0;
	wire w_dff_A_e8TKNRw88_2;
	jxor g000(.dina(w_b0_0[1]),.dinb(w_a0_0[1]),.dout(w_dff_A_i0Y4neCV3_2),.clk(gclk));
	jand g001(.dina(w_b0_0[0]),.dinb(w_a0_0[0]),.dout(n387),.clk(gclk));
	jxor g002(.dina(w_b1_0[2]),.dinb(w_a1_0[2]),.dout(n388),.clk(gclk));
	jxor g003(.dina(n388),.dinb(w_n387_0[1]),.dout(w_dff_A_0HyOVMXh8_2),.clk(gclk));
	jand g004(.dina(w_b1_0[1]),.dinb(w_a1_0[1]),.dout(n390),.clk(gclk));
	jcb g005(.dina(w_b1_0[0]),.dinb(w_a1_0[0]),.dout(n391));
	jand g006(.dina(w_dff_B_7v1bBDjM8_0),.dinb(w_n387_0[0]),.dout(n392),.clk(gclk));
	jcb g007(.dina(n392),.dinb(w_dff_B_bq66TJJL2_1),.dout(n393));
	jxor g008(.dina(w_b2_0[2]),.dinb(w_a2_0[2]),.dout(n394),.clk(gclk));
	jxor g009(.dina(w_dff_B_y2pBBYfz5_0),.dinb(w_n393_0[1]),.dout(w_dff_A_BvD62S921_2),.clk(gclk));
	jand g010(.dina(w_b2_0[1]),.dinb(w_a2_0[1]),.dout(n396),.clk(gclk));
	jcb g011(.dina(w_b2_0[0]),.dinb(w_a2_0[0]),.dout(n397));
	jand g012(.dina(w_dff_B_MevlBocM3_0),.dinb(w_n393_0[0]),.dout(n398),.clk(gclk));
	jcb g013(.dina(n398),.dinb(w_dff_B_XC6XIR9e5_1),.dout(n399));
	jxor g014(.dina(w_b3_0[2]),.dinb(w_a3_0[2]),.dout(n400),.clk(gclk));
	jxor g015(.dina(w_dff_B_S1pCGBH96_0),.dinb(w_n399_0[1]),.dout(w_dff_A_lRUw1Ruu2_2),.clk(gclk));
	jand g016(.dina(w_b3_0[1]),.dinb(w_a3_0[1]),.dout(n402),.clk(gclk));
	jcb g017(.dina(w_b3_0[0]),.dinb(w_a3_0[0]),.dout(n403));
	jand g018(.dina(w_dff_B_tOSk0HiB9_0),.dinb(w_n399_0[0]),.dout(n404),.clk(gclk));
	jcb g019(.dina(n404),.dinb(w_dff_B_RYyduIeI2_1),.dout(n405));
	jxor g020(.dina(w_b4_0[2]),.dinb(w_a4_0[2]),.dout(n406),.clk(gclk));
	jxor g021(.dina(w_dff_B_WlKsqUMj9_0),.dinb(w_n405_0[1]),.dout(w_dff_A_1VQG7qnR4_2),.clk(gclk));
	jand g022(.dina(w_b4_0[1]),.dinb(w_a4_0[1]),.dout(n408),.clk(gclk));
	jcb g023(.dina(w_b4_0[0]),.dinb(w_a4_0[0]),.dout(n409));
	jand g024(.dina(w_dff_B_NsJlHOhQ0_0),.dinb(w_n405_0[0]),.dout(n410),.clk(gclk));
	jcb g025(.dina(n410),.dinb(w_dff_B_9DVgFh9T1_1),.dout(n411));
	jxor g026(.dina(w_b5_0[2]),.dinb(w_a5_0[2]),.dout(n412),.clk(gclk));
	jxor g027(.dina(w_dff_B_Q6vqZJ6y8_0),.dinb(w_n411_0[1]),.dout(w_dff_A_IdkFl4Xp4_2),.clk(gclk));
	jand g028(.dina(w_b5_0[1]),.dinb(w_a5_0[1]),.dout(n414),.clk(gclk));
	jcb g029(.dina(w_b5_0[0]),.dinb(w_a5_0[0]),.dout(n415));
	jand g030(.dina(w_dff_B_D2KL4nNr1_0),.dinb(w_n411_0[0]),.dout(n416),.clk(gclk));
	jcb g031(.dina(n416),.dinb(w_dff_B_IAJMsY3O3_1),.dout(n417));
	jxor g032(.dina(w_b6_0[2]),.dinb(w_a6_0[2]),.dout(n418),.clk(gclk));
	jxor g033(.dina(w_dff_B_8jJ4BMCH1_0),.dinb(w_n417_0[1]),.dout(w_dff_A_IFRtoXuS7_2),.clk(gclk));
	jand g034(.dina(w_b6_0[1]),.dinb(w_a6_0[1]),.dout(n420),.clk(gclk));
	jcb g035(.dina(w_b6_0[0]),.dinb(w_a6_0[0]),.dout(n421));
	jand g036(.dina(w_dff_B_jwfquIHg2_0),.dinb(w_n417_0[0]),.dout(n422),.clk(gclk));
	jcb g037(.dina(n422),.dinb(w_dff_B_7AXejlE29_1),.dout(n423));
	jxor g038(.dina(w_b7_0[2]),.dinb(w_a7_0[2]),.dout(n424),.clk(gclk));
	jxor g039(.dina(w_dff_B_7r08WE430_0),.dinb(w_n423_0[1]),.dout(w_dff_A_sGoHlvcX8_2),.clk(gclk));
	jand g040(.dina(w_b7_0[1]),.dinb(w_a7_0[1]),.dout(n426),.clk(gclk));
	jcb g041(.dina(w_b7_0[0]),.dinb(w_a7_0[0]),.dout(n427));
	jand g042(.dina(w_dff_B_ct1c3ZgN9_0),.dinb(w_n423_0[0]),.dout(n428),.clk(gclk));
	jcb g043(.dina(n428),.dinb(w_dff_B_hLXcHmzy9_1),.dout(n429));
	jxor g044(.dina(w_b8_0[2]),.dinb(w_a8_0[2]),.dout(n430),.clk(gclk));
	jxor g045(.dina(w_dff_B_i2DkyCua4_0),.dinb(w_n429_0[1]),.dout(w_dff_A_hqBdsfmR3_2),.clk(gclk));
	jand g046(.dina(w_b8_0[1]),.dinb(w_a8_0[1]),.dout(n432),.clk(gclk));
	jcb g047(.dina(w_b8_0[0]),.dinb(w_a8_0[0]),.dout(n433));
	jand g048(.dina(w_dff_B_mJs1Nkki5_0),.dinb(w_n429_0[0]),.dout(n434),.clk(gclk));
	jcb g049(.dina(n434),.dinb(w_dff_B_N7wdEcYt6_1),.dout(n435));
	jxor g050(.dina(w_b9_0[2]),.dinb(w_a9_0[2]),.dout(n436),.clk(gclk));
	jxor g051(.dina(w_dff_B_xJonAAGK0_0),.dinb(w_n435_0[1]),.dout(w_dff_A_TPd6RMHY6_2),.clk(gclk));
	jand g052(.dina(w_b9_0[1]),.dinb(w_a9_0[1]),.dout(n438),.clk(gclk));
	jcb g053(.dina(w_b9_0[0]),.dinb(w_a9_0[0]),.dout(n439));
	jand g054(.dina(w_dff_B_oTv1F9FH9_0),.dinb(w_n435_0[0]),.dout(n440),.clk(gclk));
	jcb g055(.dina(n440),.dinb(w_dff_B_uSgQnbDf2_1),.dout(n441));
	jxor g056(.dina(w_b10_0[2]),.dinb(w_a10_0[2]),.dout(n442),.clk(gclk));
	jxor g057(.dina(w_dff_B_KD70119c7_0),.dinb(w_n441_0[1]),.dout(w_dff_A_K99ijCAz4_2),.clk(gclk));
	jand g058(.dina(w_b10_0[1]),.dinb(w_a10_0[1]),.dout(n444),.clk(gclk));
	jcb g059(.dina(w_b10_0[0]),.dinb(w_a10_0[0]),.dout(n445));
	jand g060(.dina(w_dff_B_njqcx4ts3_0),.dinb(w_n441_0[0]),.dout(n446),.clk(gclk));
	jcb g061(.dina(n446),.dinb(w_dff_B_o5sfoxtN0_1),.dout(n447));
	jxor g062(.dina(w_b11_0[2]),.dinb(w_a11_0[2]),.dout(n448),.clk(gclk));
	jxor g063(.dina(w_dff_B_i8x4P8bS8_0),.dinb(w_n447_0[1]),.dout(w_dff_A_ZrWr9ERl4_2),.clk(gclk));
	jand g064(.dina(w_b11_0[1]),.dinb(w_a11_0[1]),.dout(n450),.clk(gclk));
	jcb g065(.dina(w_b11_0[0]),.dinb(w_a11_0[0]),.dout(n451));
	jand g066(.dina(w_dff_B_nKJsQ9ti3_0),.dinb(w_n447_0[0]),.dout(n452),.clk(gclk));
	jcb g067(.dina(n452),.dinb(w_dff_B_27LeE5x30_1),.dout(n453));
	jxor g068(.dina(w_b12_0[2]),.dinb(w_a12_0[2]),.dout(n454),.clk(gclk));
	jxor g069(.dina(w_dff_B_bSj65Sek7_0),.dinb(w_n453_0[1]),.dout(w_dff_A_fR6FTcm21_2),.clk(gclk));
	jand g070(.dina(w_b12_0[1]),.dinb(w_a12_0[1]),.dout(n456),.clk(gclk));
	jcb g071(.dina(w_b12_0[0]),.dinb(w_a12_0[0]),.dout(n457));
	jand g072(.dina(w_dff_B_PT2aeLqK8_0),.dinb(w_n453_0[0]),.dout(n458),.clk(gclk));
	jcb g073(.dina(n458),.dinb(w_dff_B_Uziv0Vnv8_1),.dout(n459));
	jxor g074(.dina(w_b13_0[2]),.dinb(w_a13_0[2]),.dout(n460),.clk(gclk));
	jxor g075(.dina(w_dff_B_YbutfiBd1_0),.dinb(w_n459_0[1]),.dout(w_dff_A_4btOcuhR0_2),.clk(gclk));
	jand g076(.dina(w_b13_0[1]),.dinb(w_a13_0[1]),.dout(n462),.clk(gclk));
	jcb g077(.dina(w_b13_0[0]),.dinb(w_a13_0[0]),.dout(n463));
	jand g078(.dina(w_dff_B_hz8fGERr9_0),.dinb(w_n459_0[0]),.dout(n464),.clk(gclk));
	jcb g079(.dina(n464),.dinb(w_dff_B_EbOdpOXS9_1),.dout(n465));
	jxor g080(.dina(w_b14_0[2]),.dinb(w_a14_0[2]),.dout(n466),.clk(gclk));
	jxor g081(.dina(w_dff_B_yvhE8Xy08_0),.dinb(w_n465_0[1]),.dout(w_dff_A_KPqmqRhW5_2),.clk(gclk));
	jand g082(.dina(w_b14_0[1]),.dinb(w_a14_0[1]),.dout(n468),.clk(gclk));
	jcb g083(.dina(w_b14_0[0]),.dinb(w_a14_0[0]),.dout(n469));
	jand g084(.dina(w_dff_B_bY5KWRW79_0),.dinb(w_n465_0[0]),.dout(n470),.clk(gclk));
	jcb g085(.dina(n470),.dinb(w_dff_B_LgXnSLIA1_1),.dout(n471));
	jxor g086(.dina(w_b15_0[2]),.dinb(w_a15_0[2]),.dout(n472),.clk(gclk));
	jxor g087(.dina(w_dff_B_0CAb5BDY8_0),.dinb(w_n471_0[1]),.dout(w_dff_A_3a83FO075_2),.clk(gclk));
	jand g088(.dina(w_b15_0[1]),.dinb(w_a15_0[1]),.dout(n474),.clk(gclk));
	jcb g089(.dina(w_b15_0[0]),.dinb(w_a15_0[0]),.dout(n475));
	jand g090(.dina(w_dff_B_Azuoeek25_0),.dinb(w_n471_0[0]),.dout(n476),.clk(gclk));
	jcb g091(.dina(n476),.dinb(w_dff_B_ORoqjfaO4_1),.dout(n477));
	jxor g092(.dina(w_b16_0[2]),.dinb(w_a16_0[2]),.dout(n478),.clk(gclk));
	jxor g093(.dina(w_dff_B_M8i2g1ka6_0),.dinb(w_n477_0[1]),.dout(w_dff_A_LnRVlKwa4_2),.clk(gclk));
	jand g094(.dina(w_b16_0[1]),.dinb(w_a16_0[1]),.dout(n480),.clk(gclk));
	jcb g095(.dina(w_b16_0[0]),.dinb(w_a16_0[0]),.dout(n481));
	jand g096(.dina(w_dff_B_Ps1HkcOR8_0),.dinb(w_n477_0[0]),.dout(n482),.clk(gclk));
	jcb g097(.dina(n482),.dinb(w_dff_B_ghzowI0M3_1),.dout(n483));
	jxor g098(.dina(w_b17_0[2]),.dinb(w_a17_0[2]),.dout(n484),.clk(gclk));
	jxor g099(.dina(w_dff_B_CPSxdA6Y0_0),.dinb(w_n483_0[1]),.dout(w_dff_A_xWMjmKJE2_2),.clk(gclk));
	jand g100(.dina(w_b17_0[1]),.dinb(w_a17_0[1]),.dout(n486),.clk(gclk));
	jcb g101(.dina(w_b17_0[0]),.dinb(w_a17_0[0]),.dout(n487));
	jand g102(.dina(w_dff_B_M2JhGCeu4_0),.dinb(w_n483_0[0]),.dout(n488),.clk(gclk));
	jcb g103(.dina(n488),.dinb(w_dff_B_LxQ84mjb0_1),.dout(n489));
	jxor g104(.dina(w_b18_0[2]),.dinb(w_a18_0[2]),.dout(n490),.clk(gclk));
	jxor g105(.dina(w_dff_B_c7YZMJgL7_0),.dinb(w_n489_0[1]),.dout(w_dff_A_0NVR8Dal9_2),.clk(gclk));
	jand g106(.dina(w_b18_0[1]),.dinb(w_a18_0[1]),.dout(n492),.clk(gclk));
	jcb g107(.dina(w_b18_0[0]),.dinb(w_a18_0[0]),.dout(n493));
	jand g108(.dina(w_dff_B_bS2zNEr15_0),.dinb(w_n489_0[0]),.dout(n494),.clk(gclk));
	jcb g109(.dina(n494),.dinb(w_dff_B_EWKSzcRm1_1),.dout(n495));
	jxor g110(.dina(w_b19_0[2]),.dinb(w_a19_0[2]),.dout(n496),.clk(gclk));
	jxor g111(.dina(w_dff_B_XC5aVfCd5_0),.dinb(w_n495_0[1]),.dout(w_dff_A_Bp4ITOiF1_2),.clk(gclk));
	jand g112(.dina(w_b19_0[1]),.dinb(w_a19_0[1]),.dout(n498),.clk(gclk));
	jcb g113(.dina(w_b19_0[0]),.dinb(w_a19_0[0]),.dout(n499));
	jand g114(.dina(w_dff_B_CcU9AiUi0_0),.dinb(w_n495_0[0]),.dout(n500),.clk(gclk));
	jcb g115(.dina(n500),.dinb(w_dff_B_eyYJitxH0_1),.dout(n501));
	jxor g116(.dina(w_b20_0[2]),.dinb(w_a20_0[2]),.dout(n502),.clk(gclk));
	jxor g117(.dina(w_dff_B_3Qs1UfWC8_0),.dinb(w_n501_0[1]),.dout(w_dff_A_UvvGn9rX2_2),.clk(gclk));
	jand g118(.dina(w_b20_0[1]),.dinb(w_a20_0[1]),.dout(n504),.clk(gclk));
	jcb g119(.dina(w_b20_0[0]),.dinb(w_a20_0[0]),.dout(n505));
	jand g120(.dina(w_dff_B_srqfiaFR0_0),.dinb(w_n501_0[0]),.dout(n506),.clk(gclk));
	jcb g121(.dina(n506),.dinb(w_dff_B_wFlt2aWE8_1),.dout(n507));
	jxor g122(.dina(w_b21_0[2]),.dinb(w_a21_0[2]),.dout(n508),.clk(gclk));
	jxor g123(.dina(w_dff_B_bBoBpv7g8_0),.dinb(w_n507_0[1]),.dout(w_dff_A_lCHLbsXY9_2),.clk(gclk));
	jand g124(.dina(w_b21_0[1]),.dinb(w_a21_0[1]),.dout(n510),.clk(gclk));
	jcb g125(.dina(w_b21_0[0]),.dinb(w_a21_0[0]),.dout(n511));
	jand g126(.dina(w_dff_B_TpJykMPA5_0),.dinb(w_n507_0[0]),.dout(n512),.clk(gclk));
	jcb g127(.dina(n512),.dinb(w_dff_B_k8b5cujs9_1),.dout(n513));
	jxor g128(.dina(w_b22_0[2]),.dinb(w_a22_0[2]),.dout(n514),.clk(gclk));
	jxor g129(.dina(w_dff_B_3eiO5ewK6_0),.dinb(w_n513_0[1]),.dout(w_dff_A_bwlIPVrT6_2),.clk(gclk));
	jand g130(.dina(w_b22_0[1]),.dinb(w_a22_0[1]),.dout(n516),.clk(gclk));
	jcb g131(.dina(w_b22_0[0]),.dinb(w_a22_0[0]),.dout(n517));
	jand g132(.dina(w_dff_B_nKZIowO61_0),.dinb(w_n513_0[0]),.dout(n518),.clk(gclk));
	jcb g133(.dina(n518),.dinb(w_dff_B_tOY8ECp76_1),.dout(n519));
	jxor g134(.dina(w_b23_0[2]),.dinb(w_a23_0[2]),.dout(n520),.clk(gclk));
	jxor g135(.dina(w_dff_B_tF6BKpIu3_0),.dinb(w_n519_0[1]),.dout(w_dff_A_SzoSoT3h7_2),.clk(gclk));
	jand g136(.dina(w_b23_0[1]),.dinb(w_a23_0[1]),.dout(n522),.clk(gclk));
	jcb g137(.dina(w_b23_0[0]),.dinb(w_a23_0[0]),.dout(n523));
	jand g138(.dina(w_dff_B_vffmUHZP1_0),.dinb(w_n519_0[0]),.dout(n524),.clk(gclk));
	jcb g139(.dina(n524),.dinb(w_dff_B_fxvTyWRy8_1),.dout(n525));
	jxor g140(.dina(w_b24_0[2]),.dinb(w_a24_0[2]),.dout(n526),.clk(gclk));
	jxor g141(.dina(w_dff_B_IxLjw79f1_0),.dinb(w_n525_0[1]),.dout(w_dff_A_ejqy7DXE0_2),.clk(gclk));
	jand g142(.dina(w_b24_0[1]),.dinb(w_a24_0[1]),.dout(n528),.clk(gclk));
	jcb g143(.dina(w_b24_0[0]),.dinb(w_a24_0[0]),.dout(n529));
	jand g144(.dina(w_dff_B_WEHr8swc1_0),.dinb(w_n525_0[0]),.dout(n530),.clk(gclk));
	jcb g145(.dina(n530),.dinb(w_dff_B_mAYLtnxH0_1),.dout(n531));
	jxor g146(.dina(w_b25_0[2]),.dinb(w_a25_0[2]),.dout(n532),.clk(gclk));
	jxor g147(.dina(w_dff_B_poGlmfvO9_0),.dinb(w_n531_0[1]),.dout(w_dff_A_0nEZ1YGf2_2),.clk(gclk));
	jand g148(.dina(w_b25_0[1]),.dinb(w_a25_0[1]),.dout(n534),.clk(gclk));
	jcb g149(.dina(w_b25_0[0]),.dinb(w_a25_0[0]),.dout(n535));
	jand g150(.dina(w_dff_B_kc8HMq882_0),.dinb(w_n531_0[0]),.dout(n536),.clk(gclk));
	jcb g151(.dina(n536),.dinb(w_dff_B_nk8Q4hzv5_1),.dout(n537));
	jxor g152(.dina(w_b26_0[2]),.dinb(w_a26_0[2]),.dout(n538),.clk(gclk));
	jxor g153(.dina(w_dff_B_aSGLFurX1_0),.dinb(w_n537_0[1]),.dout(w_dff_A_M4eemYt31_2),.clk(gclk));
	jand g154(.dina(w_b26_0[1]),.dinb(w_a26_0[1]),.dout(n540),.clk(gclk));
	jcb g155(.dina(w_b26_0[0]),.dinb(w_a26_0[0]),.dout(n541));
	jand g156(.dina(w_dff_B_bFwFmeEw7_0),.dinb(w_n537_0[0]),.dout(n542),.clk(gclk));
	jcb g157(.dina(n542),.dinb(w_dff_B_YvVPAofT6_1),.dout(n543));
	jxor g158(.dina(w_b27_0[2]),.dinb(w_a27_0[2]),.dout(n544),.clk(gclk));
	jxor g159(.dina(w_dff_B_0AYkSjrX9_0),.dinb(w_n543_0[1]),.dout(w_dff_A_JIss0YJB5_2),.clk(gclk));
	jand g160(.dina(w_b27_0[1]),.dinb(w_a27_0[1]),.dout(n546),.clk(gclk));
	jcb g161(.dina(w_b27_0[0]),.dinb(w_a27_0[0]),.dout(n547));
	jand g162(.dina(w_dff_B_d3Bc1Lmg9_0),.dinb(w_n543_0[0]),.dout(n548),.clk(gclk));
	jcb g163(.dina(n548),.dinb(w_dff_B_UIEJM1lk8_1),.dout(n549));
	jxor g164(.dina(w_b28_0[2]),.dinb(w_a28_0[2]),.dout(n550),.clk(gclk));
	jxor g165(.dina(w_dff_B_bWpvlkFu0_0),.dinb(w_n549_0[1]),.dout(w_dff_A_7BbhU6Rh4_2),.clk(gclk));
	jand g166(.dina(w_b28_0[1]),.dinb(w_a28_0[1]),.dout(n552),.clk(gclk));
	jcb g167(.dina(w_b28_0[0]),.dinb(w_a28_0[0]),.dout(n553));
	jand g168(.dina(w_dff_B_X8LY3C7p1_0),.dinb(w_n549_0[0]),.dout(n554),.clk(gclk));
	jcb g169(.dina(n554),.dinb(w_dff_B_2YMJeXnr4_1),.dout(n555));
	jxor g170(.dina(w_b29_0[2]),.dinb(w_a29_0[2]),.dout(n556),.clk(gclk));
	jxor g171(.dina(w_dff_B_OxgAFEkU9_0),.dinb(w_n555_0[1]),.dout(w_dff_A_MfypuXxv4_2),.clk(gclk));
	jand g172(.dina(w_b29_0[1]),.dinb(w_a29_0[1]),.dout(n558),.clk(gclk));
	jcb g173(.dina(w_b29_0[0]),.dinb(w_a29_0[0]),.dout(n559));
	jand g174(.dina(w_dff_B_qICniHxc5_0),.dinb(w_n555_0[0]),.dout(n560),.clk(gclk));
	jcb g175(.dina(n560),.dinb(w_dff_B_8BjQK9zd0_1),.dout(n561));
	jxor g176(.dina(w_b30_0[2]),.dinb(w_a30_0[2]),.dout(n562),.clk(gclk));
	jxor g177(.dina(w_dff_B_0NQGDTyH9_0),.dinb(w_n561_0[1]),.dout(w_dff_A_m45eyEAd4_2),.clk(gclk));
	jand g178(.dina(w_b30_0[1]),.dinb(w_a30_0[1]),.dout(n564),.clk(gclk));
	jcb g179(.dina(w_b30_0[0]),.dinb(w_a30_0[0]),.dout(n565));
	jand g180(.dina(w_dff_B_norHvl765_0),.dinb(w_n561_0[0]),.dout(n566),.clk(gclk));
	jcb g181(.dina(n566),.dinb(w_dff_B_fYp7rwhu5_1),.dout(n567));
	jxor g182(.dina(w_b31_0[2]),.dinb(w_a31_0[2]),.dout(n568),.clk(gclk));
	jxor g183(.dina(w_dff_B_yCmWmTN77_0),.dinb(w_n567_0[1]),.dout(w_dff_A_HDJk7IDG5_2),.clk(gclk));
	jand g184(.dina(w_b31_0[1]),.dinb(w_a31_0[1]),.dout(n570),.clk(gclk));
	jcb g185(.dina(w_b31_0[0]),.dinb(w_a31_0[0]),.dout(n571));
	jand g186(.dina(w_dff_B_znPY8YBC7_0),.dinb(w_n567_0[0]),.dout(n572),.clk(gclk));
	jcb g187(.dina(n572),.dinb(w_dff_B_MqGZ9eEe7_1),.dout(n573));
	jxor g188(.dina(w_b32_0[2]),.dinb(w_a32_0[2]),.dout(n574),.clk(gclk));
	jxor g189(.dina(w_dff_B_FPJBFbiz2_0),.dinb(w_n573_0[1]),.dout(w_dff_A_Vbwd5rP60_2),.clk(gclk));
	jand g190(.dina(w_b32_0[1]),.dinb(w_a32_0[1]),.dout(n576),.clk(gclk));
	jcb g191(.dina(w_b32_0[0]),.dinb(w_a32_0[0]),.dout(n577));
	jand g192(.dina(w_dff_B_cOSHsCTW4_0),.dinb(w_n573_0[0]),.dout(n578),.clk(gclk));
	jcb g193(.dina(n578),.dinb(w_dff_B_vpzfAeXc3_1),.dout(n579));
	jxor g194(.dina(w_b33_0[2]),.dinb(w_a33_0[2]),.dout(n580),.clk(gclk));
	jxor g195(.dina(w_dff_B_Qyetcsqv4_0),.dinb(w_n579_0[1]),.dout(w_dff_A_AA7idxgZ2_2),.clk(gclk));
	jand g196(.dina(w_b33_0[1]),.dinb(w_a33_0[1]),.dout(n582),.clk(gclk));
	jcb g197(.dina(w_b33_0[0]),.dinb(w_a33_0[0]),.dout(n583));
	jand g198(.dina(w_dff_B_76wrGEuj0_0),.dinb(w_n579_0[0]),.dout(n584),.clk(gclk));
	jcb g199(.dina(n584),.dinb(w_dff_B_D2kiPHXL3_1),.dout(n585));
	jxor g200(.dina(w_b34_0[2]),.dinb(w_a34_0[2]),.dout(n586),.clk(gclk));
	jxor g201(.dina(w_dff_B_WbAXqjB88_0),.dinb(w_n585_0[1]),.dout(w_dff_A_RzzGmYzn3_2),.clk(gclk));
	jand g202(.dina(w_b34_0[1]),.dinb(w_a34_0[1]),.dout(n588),.clk(gclk));
	jcb g203(.dina(w_b34_0[0]),.dinb(w_a34_0[0]),.dout(n589));
	jand g204(.dina(w_dff_B_NuWicBqk2_0),.dinb(w_n585_0[0]),.dout(n590),.clk(gclk));
	jcb g205(.dina(n590),.dinb(w_dff_B_xBRXkssz2_1),.dout(n591));
	jxor g206(.dina(w_b35_0[2]),.dinb(w_a35_0[2]),.dout(n592),.clk(gclk));
	jxor g207(.dina(w_dff_B_tTqoaoGw3_0),.dinb(w_n591_0[1]),.dout(w_dff_A_tKTU1hRn7_2),.clk(gclk));
	jand g208(.dina(w_b35_0[1]),.dinb(w_a35_0[1]),.dout(n594),.clk(gclk));
	jcb g209(.dina(w_b35_0[0]),.dinb(w_a35_0[0]),.dout(n595));
	jand g210(.dina(w_dff_B_N2n8UqAM7_0),.dinb(w_n591_0[0]),.dout(n596),.clk(gclk));
	jcb g211(.dina(n596),.dinb(w_dff_B_PbcuSyj41_1),.dout(n597));
	jxor g212(.dina(w_b36_0[2]),.dinb(w_a36_0[2]),.dout(n598),.clk(gclk));
	jxor g213(.dina(w_dff_B_OVSEBGFt8_0),.dinb(w_n597_0[1]),.dout(w_dff_A_F7Oq80ij2_2),.clk(gclk));
	jand g214(.dina(w_b36_0[1]),.dinb(w_a36_0[1]),.dout(n600),.clk(gclk));
	jcb g215(.dina(w_b36_0[0]),.dinb(w_a36_0[0]),.dout(n601));
	jand g216(.dina(w_dff_B_Giv88Gjw1_0),.dinb(w_n597_0[0]),.dout(n602),.clk(gclk));
	jcb g217(.dina(n602),.dinb(w_dff_B_ntOAyf159_1),.dout(n603));
	jxor g218(.dina(w_b37_0[2]),.dinb(w_a37_0[2]),.dout(n604),.clk(gclk));
	jxor g219(.dina(w_dff_B_hF6XnBIn6_0),.dinb(w_n603_0[1]),.dout(w_dff_A_nym5NQ194_2),.clk(gclk));
	jand g220(.dina(w_b37_0[1]),.dinb(w_a37_0[1]),.dout(n606),.clk(gclk));
	jcb g221(.dina(w_b37_0[0]),.dinb(w_a37_0[0]),.dout(n607));
	jand g222(.dina(w_dff_B_vt7Bt9w49_0),.dinb(w_n603_0[0]),.dout(n608),.clk(gclk));
	jcb g223(.dina(n608),.dinb(w_dff_B_S6RAvCjq6_1),.dout(n609));
	jxor g224(.dina(w_b38_0[2]),.dinb(w_a38_0[2]),.dout(n610),.clk(gclk));
	jxor g225(.dina(w_dff_B_oTtWTlv49_0),.dinb(w_n609_0[1]),.dout(w_dff_A_4Rn8acWn9_2),.clk(gclk));
	jand g226(.dina(w_b38_0[1]),.dinb(w_a38_0[1]),.dout(n612),.clk(gclk));
	jcb g227(.dina(w_b38_0[0]),.dinb(w_a38_0[0]),.dout(n613));
	jand g228(.dina(w_dff_B_wdau1vMx1_0),.dinb(w_n609_0[0]),.dout(n614),.clk(gclk));
	jcb g229(.dina(n614),.dinb(w_dff_B_u1eB0U854_1),.dout(n615));
	jxor g230(.dina(w_b39_0[2]),.dinb(w_a39_0[2]),.dout(n616),.clk(gclk));
	jxor g231(.dina(w_dff_B_KlorpDbQ7_0),.dinb(w_n615_0[1]),.dout(w_dff_A_f746W3Pr1_2),.clk(gclk));
	jand g232(.dina(w_b39_0[1]),.dinb(w_a39_0[1]),.dout(n618),.clk(gclk));
	jcb g233(.dina(w_b39_0[0]),.dinb(w_a39_0[0]),.dout(n619));
	jand g234(.dina(w_dff_B_GoygnPeZ7_0),.dinb(w_n615_0[0]),.dout(n620),.clk(gclk));
	jcb g235(.dina(n620),.dinb(w_dff_B_1cZChDiV8_1),.dout(n621));
	jxor g236(.dina(w_b40_0[2]),.dinb(w_a40_0[2]),.dout(n622),.clk(gclk));
	jxor g237(.dina(w_dff_B_eIHhFn8J8_0),.dinb(w_n621_0[1]),.dout(w_dff_A_m6wDD8ja6_2),.clk(gclk));
	jand g238(.dina(w_b40_0[1]),.dinb(w_a40_0[1]),.dout(n624),.clk(gclk));
	jcb g239(.dina(w_b40_0[0]),.dinb(w_a40_0[0]),.dout(n625));
	jand g240(.dina(w_dff_B_v6JmAK7j4_0),.dinb(w_n621_0[0]),.dout(n626),.clk(gclk));
	jcb g241(.dina(n626),.dinb(w_dff_B_snRizMBV3_1),.dout(n627));
	jxor g242(.dina(w_b41_0[2]),.dinb(w_a41_0[2]),.dout(n628),.clk(gclk));
	jxor g243(.dina(w_dff_B_HBMFIay39_0),.dinb(w_n627_0[1]),.dout(w_dff_A_6JBK2nPW1_2),.clk(gclk));
	jand g244(.dina(w_b41_0[1]),.dinb(w_a41_0[1]),.dout(n630),.clk(gclk));
	jcb g245(.dina(w_b41_0[0]),.dinb(w_a41_0[0]),.dout(n631));
	jand g246(.dina(w_dff_B_Vysb7cc73_0),.dinb(w_n627_0[0]),.dout(n632),.clk(gclk));
	jcb g247(.dina(n632),.dinb(w_dff_B_AyOrLbF03_1),.dout(n633));
	jxor g248(.dina(w_b42_0[2]),.dinb(w_a42_0[2]),.dout(n634),.clk(gclk));
	jxor g249(.dina(w_dff_B_UJ4VqMGy1_0),.dinb(w_n633_0[1]),.dout(w_dff_A_09ujqjlu8_2),.clk(gclk));
	jand g250(.dina(w_b42_0[1]),.dinb(w_a42_0[1]),.dout(n636),.clk(gclk));
	jcb g251(.dina(w_b42_0[0]),.dinb(w_a42_0[0]),.dout(n637));
	jand g252(.dina(w_dff_B_Fe0B8YFI0_0),.dinb(w_n633_0[0]),.dout(n638),.clk(gclk));
	jcb g253(.dina(n638),.dinb(w_dff_B_JMCouiXX8_1),.dout(n639));
	jxor g254(.dina(w_b43_0[2]),.dinb(w_a43_0[2]),.dout(n640),.clk(gclk));
	jxor g255(.dina(w_dff_B_t6QLfecs2_0),.dinb(w_n639_0[1]),.dout(w_dff_A_I2YmvXsD7_2),.clk(gclk));
	jand g256(.dina(w_b43_0[1]),.dinb(w_a43_0[1]),.dout(n642),.clk(gclk));
	jcb g257(.dina(w_b43_0[0]),.dinb(w_a43_0[0]),.dout(n643));
	jand g258(.dina(w_dff_B_O1mNMYi88_0),.dinb(w_n639_0[0]),.dout(n644),.clk(gclk));
	jcb g259(.dina(n644),.dinb(w_dff_B_OGZRqfWA9_1),.dout(n645));
	jxor g260(.dina(w_b44_0[2]),.dinb(w_a44_0[2]),.dout(n646),.clk(gclk));
	jxor g261(.dina(w_dff_B_2nixnkQN6_0),.dinb(w_n645_0[1]),.dout(w_dff_A_QwZFXhVA9_2),.clk(gclk));
	jand g262(.dina(w_b44_0[1]),.dinb(w_a44_0[1]),.dout(n648),.clk(gclk));
	jcb g263(.dina(w_b44_0[0]),.dinb(w_a44_0[0]),.dout(n649));
	jand g264(.dina(w_dff_B_XJ6b8ERc3_0),.dinb(w_n645_0[0]),.dout(n650),.clk(gclk));
	jcb g265(.dina(n650),.dinb(w_dff_B_y5N9hr4K5_1),.dout(n651));
	jxor g266(.dina(w_b45_0[2]),.dinb(w_a45_0[2]),.dout(n652),.clk(gclk));
	jxor g267(.dina(w_dff_B_9PsGZFcP4_0),.dinb(w_n651_0[1]),.dout(w_dff_A_VA8FezrL8_2),.clk(gclk));
	jand g268(.dina(w_b45_0[1]),.dinb(w_a45_0[1]),.dout(n654),.clk(gclk));
	jcb g269(.dina(w_b45_0[0]),.dinb(w_a45_0[0]),.dout(n655));
	jand g270(.dina(w_dff_B_ru1ByfvL1_0),.dinb(w_n651_0[0]),.dout(n656),.clk(gclk));
	jcb g271(.dina(n656),.dinb(w_dff_B_Fx8sXFkn9_1),.dout(n657));
	jxor g272(.dina(w_b46_0[2]),.dinb(w_a46_0[2]),.dout(n658),.clk(gclk));
	jxor g273(.dina(w_dff_B_90EtCyrN6_0),.dinb(w_n657_0[1]),.dout(w_dff_A_HG05Fu3s6_2),.clk(gclk));
	jand g274(.dina(w_b46_0[1]),.dinb(w_a46_0[1]),.dout(n660),.clk(gclk));
	jcb g275(.dina(w_b46_0[0]),.dinb(w_a46_0[0]),.dout(n661));
	jand g276(.dina(w_dff_B_ZUFZvbyO9_0),.dinb(w_n657_0[0]),.dout(n662),.clk(gclk));
	jcb g277(.dina(n662),.dinb(w_dff_B_ka8N4w5F3_1),.dout(n663));
	jxor g278(.dina(w_b47_0[2]),.dinb(w_a47_0[2]),.dout(n664),.clk(gclk));
	jxor g279(.dina(w_dff_B_mkYl9cwU3_0),.dinb(w_n663_0[1]),.dout(w_dff_A_AIhCfEsq4_2),.clk(gclk));
	jand g280(.dina(w_b47_0[1]),.dinb(w_a47_0[1]),.dout(n666),.clk(gclk));
	jcb g281(.dina(w_b47_0[0]),.dinb(w_a47_0[0]),.dout(n667));
	jand g282(.dina(w_dff_B_dL6uwy6j5_0),.dinb(w_n663_0[0]),.dout(n668),.clk(gclk));
	jcb g283(.dina(n668),.dinb(w_dff_B_HGuNeMUK0_1),.dout(n669));
	jxor g284(.dina(w_b48_0[2]),.dinb(w_a48_0[2]),.dout(n670),.clk(gclk));
	jxor g285(.dina(w_dff_B_BfaZkbuX5_0),.dinb(w_n669_0[1]),.dout(w_dff_A_aJxExRy15_2),.clk(gclk));
	jand g286(.dina(w_b48_0[1]),.dinb(w_a48_0[1]),.dout(n672),.clk(gclk));
	jcb g287(.dina(w_b48_0[0]),.dinb(w_a48_0[0]),.dout(n673));
	jand g288(.dina(w_dff_B_YAxWtq8t8_0),.dinb(w_n669_0[0]),.dout(n674),.clk(gclk));
	jcb g289(.dina(n674),.dinb(w_dff_B_jwcKYoSU1_1),.dout(n675));
	jxor g290(.dina(w_b49_0[2]),.dinb(w_a49_0[2]),.dout(n676),.clk(gclk));
	jxor g291(.dina(w_dff_B_DruCwV8I3_0),.dinb(w_n675_0[1]),.dout(w_dff_A_3mKSz1HS2_2),.clk(gclk));
	jand g292(.dina(w_b49_0[1]),.dinb(w_a49_0[1]),.dout(n678),.clk(gclk));
	jcb g293(.dina(w_b49_0[0]),.dinb(w_a49_0[0]),.dout(n679));
	jand g294(.dina(w_dff_B_CtINLd6Q5_0),.dinb(w_n675_0[0]),.dout(n680),.clk(gclk));
	jcb g295(.dina(n680),.dinb(w_dff_B_GecnHXzy9_1),.dout(n681));
	jxor g296(.dina(w_b50_0[2]),.dinb(w_a50_0[2]),.dout(n682),.clk(gclk));
	jxor g297(.dina(w_dff_B_jmJiXT5P3_0),.dinb(w_n681_0[1]),.dout(w_dff_A_s2adAl7P4_2),.clk(gclk));
	jand g298(.dina(w_b50_0[1]),.dinb(w_a50_0[1]),.dout(n684),.clk(gclk));
	jcb g299(.dina(w_b50_0[0]),.dinb(w_a50_0[0]),.dout(n685));
	jand g300(.dina(w_dff_B_puRmXWhG3_0),.dinb(w_n681_0[0]),.dout(n686),.clk(gclk));
	jcb g301(.dina(n686),.dinb(w_dff_B_YfcGYVQq4_1),.dout(n687));
	jxor g302(.dina(w_b51_0[2]),.dinb(w_a51_0[2]),.dout(n688),.clk(gclk));
	jxor g303(.dina(w_dff_B_V9qk1Xe17_0),.dinb(w_n687_0[1]),.dout(w_dff_A_FVUuRbF61_2),.clk(gclk));
	jand g304(.dina(w_b51_0[1]),.dinb(w_a51_0[1]),.dout(n690),.clk(gclk));
	jcb g305(.dina(w_b51_0[0]),.dinb(w_a51_0[0]),.dout(n691));
	jand g306(.dina(w_dff_B_pJXXJjmH2_0),.dinb(w_n687_0[0]),.dout(n692),.clk(gclk));
	jcb g307(.dina(n692),.dinb(w_dff_B_YvJN65Kw3_1),.dout(n693));
	jxor g308(.dina(w_b52_0[2]),.dinb(w_a52_0[2]),.dout(n694),.clk(gclk));
	jxor g309(.dina(w_dff_B_oLurYfyu7_0),.dinb(w_n693_0[1]),.dout(w_dff_A_G7GNSuM17_2),.clk(gclk));
	jand g310(.dina(w_b52_0[1]),.dinb(w_a52_0[1]),.dout(n696),.clk(gclk));
	jcb g311(.dina(w_b52_0[0]),.dinb(w_a52_0[0]),.dout(n697));
	jand g312(.dina(w_dff_B_YyW5ipZv0_0),.dinb(w_n693_0[0]),.dout(n698),.clk(gclk));
	jcb g313(.dina(n698),.dinb(w_dff_B_79nILaoK7_1),.dout(n699));
	jxor g314(.dina(w_b53_0[2]),.dinb(w_a53_0[2]),.dout(n700),.clk(gclk));
	jxor g315(.dina(w_dff_B_pKa8yGRz6_0),.dinb(w_n699_0[1]),.dout(w_dff_A_J9A7hwTx6_2),.clk(gclk));
	jand g316(.dina(w_b53_0[1]),.dinb(w_a53_0[1]),.dout(n702),.clk(gclk));
	jcb g317(.dina(w_b53_0[0]),.dinb(w_a53_0[0]),.dout(n703));
	jand g318(.dina(w_dff_B_PKOhVjuX2_0),.dinb(w_n699_0[0]),.dout(n704),.clk(gclk));
	jcb g319(.dina(n704),.dinb(w_dff_B_NmBOBsht4_1),.dout(n705));
	jxor g320(.dina(w_b54_0[2]),.dinb(w_a54_0[2]),.dout(n706),.clk(gclk));
	jxor g321(.dina(w_dff_B_U7KCbJ7j9_0),.dinb(w_n705_0[1]),.dout(w_dff_A_VAnnSBRN8_2),.clk(gclk));
	jand g322(.dina(w_b54_0[1]),.dinb(w_a54_0[1]),.dout(n708),.clk(gclk));
	jcb g323(.dina(w_b54_0[0]),.dinb(w_a54_0[0]),.dout(n709));
	jand g324(.dina(w_dff_B_PGiiN9Zt6_0),.dinb(w_n705_0[0]),.dout(n710),.clk(gclk));
	jcb g325(.dina(n710),.dinb(w_dff_B_o4QB8nIG6_1),.dout(n711));
	jxor g326(.dina(w_b55_0[2]),.dinb(w_a55_0[2]),.dout(n712),.clk(gclk));
	jxor g327(.dina(w_dff_B_vinPkQyy1_0),.dinb(w_n711_0[1]),.dout(w_dff_A_w2HyVyOp2_2),.clk(gclk));
	jand g328(.dina(w_b55_0[1]),.dinb(w_a55_0[1]),.dout(n714),.clk(gclk));
	jcb g329(.dina(w_b55_0[0]),.dinb(w_a55_0[0]),.dout(n715));
	jand g330(.dina(w_dff_B_krSKQ8iz1_0),.dinb(w_n711_0[0]),.dout(n716),.clk(gclk));
	jcb g331(.dina(n716),.dinb(w_dff_B_2n0kw3zB1_1),.dout(n717));
	jxor g332(.dina(w_b56_0[2]),.dinb(w_a56_0[2]),.dout(n718),.clk(gclk));
	jxor g333(.dina(w_dff_B_YzSXgHQL7_0),.dinb(w_n717_0[1]),.dout(w_dff_A_0ifBWpOE0_2),.clk(gclk));
	jand g334(.dina(w_b56_0[1]),.dinb(w_a56_0[1]),.dout(n720),.clk(gclk));
	jcb g335(.dina(w_b56_0[0]),.dinb(w_a56_0[0]),.dout(n721));
	jand g336(.dina(w_dff_B_3PM2Wo7i4_0),.dinb(w_n717_0[0]),.dout(n722),.clk(gclk));
	jcb g337(.dina(n722),.dinb(w_dff_B_7hG8iOrA5_1),.dout(n723));
	jxor g338(.dina(w_b57_0[2]),.dinb(w_a57_0[2]),.dout(n724),.clk(gclk));
	jxor g339(.dina(w_dff_B_n1rpOmAn9_0),.dinb(w_n723_0[1]),.dout(w_dff_A_INrlTL4v6_2),.clk(gclk));
	jand g340(.dina(w_b57_0[1]),.dinb(w_a57_0[1]),.dout(n726),.clk(gclk));
	jcb g341(.dina(w_b57_0[0]),.dinb(w_a57_0[0]),.dout(n727));
	jand g342(.dina(w_dff_B_y4LeRC6T7_0),.dinb(w_n723_0[0]),.dout(n728),.clk(gclk));
	jcb g343(.dina(n728),.dinb(w_dff_B_oG1alkJt9_1),.dout(n729));
	jxor g344(.dina(w_b58_0[2]),.dinb(w_a58_0[2]),.dout(n730),.clk(gclk));
	jxor g345(.dina(w_dff_B_GE2mGqKL5_0),.dinb(w_n729_0[1]),.dout(w_dff_A_IAZs4o3E0_2),.clk(gclk));
	jand g346(.dina(w_b58_0[1]),.dinb(w_a58_0[1]),.dout(n732),.clk(gclk));
	jcb g347(.dina(w_b58_0[0]),.dinb(w_a58_0[0]),.dout(n733));
	jand g348(.dina(w_dff_B_jX94jsrp1_0),.dinb(w_n729_0[0]),.dout(n734),.clk(gclk));
	jcb g349(.dina(n734),.dinb(w_dff_B_WezfSukm9_1),.dout(n735));
	jxor g350(.dina(w_b59_0[2]),.dinb(w_a59_0[2]),.dout(n736),.clk(gclk));
	jxor g351(.dina(w_dff_B_UNX9CF5n9_0),.dinb(w_n735_0[1]),.dout(w_dff_A_bZXjmX1T8_2),.clk(gclk));
	jand g352(.dina(w_b59_0[1]),.dinb(w_a59_0[1]),.dout(n738),.clk(gclk));
	jcb g353(.dina(w_b59_0[0]),.dinb(w_a59_0[0]),.dout(n739));
	jand g354(.dina(w_dff_B_pQOVSYfd7_0),.dinb(w_n735_0[0]),.dout(n740),.clk(gclk));
	jcb g355(.dina(n740),.dinb(w_dff_B_NtYVoxbX5_1),.dout(n741));
	jxor g356(.dina(w_b60_0[2]),.dinb(w_a60_0[2]),.dout(n742),.clk(gclk));
	jxor g357(.dina(w_dff_B_2Kzh4c4E2_0),.dinb(w_n741_0[1]),.dout(w_dff_A_73F8XiAD0_2),.clk(gclk));
	jand g358(.dina(w_b60_0[1]),.dinb(w_a60_0[1]),.dout(n744),.clk(gclk));
	jcb g359(.dina(w_b60_0[0]),.dinb(w_a60_0[0]),.dout(n745));
	jand g360(.dina(w_dff_B_LsprbBuG0_0),.dinb(w_n741_0[0]),.dout(n746),.clk(gclk));
	jcb g361(.dina(n746),.dinb(w_dff_B_gZ9xFATs7_1),.dout(n747));
	jxor g362(.dina(w_b61_0[2]),.dinb(w_a61_0[2]),.dout(n748),.clk(gclk));
	jxor g363(.dina(w_dff_B_OOaMoRMD8_0),.dinb(w_n747_0[1]),.dout(w_dff_A_cbJx3cUU7_2),.clk(gclk));
	jand g364(.dina(w_b61_0[1]),.dinb(w_a61_0[1]),.dout(n750),.clk(gclk));
	jcb g365(.dina(w_b61_0[0]),.dinb(w_a61_0[0]),.dout(n751));
	jand g366(.dina(w_dff_B_nUECFkPE3_0),.dinb(w_n747_0[0]),.dout(n752),.clk(gclk));
	jcb g367(.dina(n752),.dinb(w_dff_B_uGDXx6qa1_1),.dout(n753));
	jxor g368(.dina(w_b62_0[2]),.dinb(w_a62_0[2]),.dout(n754),.clk(gclk));
	jxor g369(.dina(w_dff_B_fMEyUaIT3_0),.dinb(w_n753_0[1]),.dout(w_dff_A_9pd4SMnz2_2),.clk(gclk));
	jand g370(.dina(w_b62_0[1]),.dinb(w_a62_0[1]),.dout(n756),.clk(gclk));
	jcb g371(.dina(w_b62_0[0]),.dinb(w_a62_0[0]),.dout(n757));
	jand g372(.dina(w_dff_B_fIXrmCN75_0),.dinb(w_n753_0[0]),.dout(n758),.clk(gclk));
	jcb g373(.dina(n758),.dinb(w_dff_B_cMTGAhWx0_1),.dout(n759));
	jxor g374(.dina(w_b63_0[2]),.dinb(w_a63_0[2]),.dout(n760),.clk(gclk));
	jxor g375(.dina(w_dff_B_X8L8LwPo4_0),.dinb(w_n759_0[1]),.dout(w_dff_A_was1nG0s4_2),.clk(gclk));
	jand g376(.dina(w_b63_0[1]),.dinb(w_a63_0[1]),.dout(n762),.clk(gclk));
	jcb g377(.dina(w_b63_0[0]),.dinb(w_a63_0[0]),.dout(n763));
	jand g378(.dina(w_dff_B_J5sqkVLr6_0),.dinb(w_n759_0[0]),.dout(n764),.clk(gclk));
	jcb g379(.dina(n764),.dinb(w_dff_B_HRhAL3Ck5_1),.dout(n765));
	jxor g380(.dina(w_b64_0[2]),.dinb(w_a64_0[2]),.dout(n766),.clk(gclk));
	jxor g381(.dina(w_dff_B_9ivRqQdT2_0),.dinb(w_n765_0[1]),.dout(w_dff_A_fVeXfF3y3_2),.clk(gclk));
	jand g382(.dina(w_b64_0[1]),.dinb(w_a64_0[1]),.dout(n768),.clk(gclk));
	jcb g383(.dina(w_b64_0[0]),.dinb(w_a64_0[0]),.dout(n769));
	jand g384(.dina(w_dff_B_Xj7EsTj23_0),.dinb(w_n765_0[0]),.dout(n770),.clk(gclk));
	jcb g385(.dina(n770),.dinb(w_dff_B_7KmGZ0V04_1),.dout(n771));
	jxor g386(.dina(w_b65_0[2]),.dinb(w_a65_0[2]),.dout(n772),.clk(gclk));
	jxor g387(.dina(w_dff_B_zX9xjztb5_0),.dinb(w_n771_0[1]),.dout(w_dff_A_apv54JrL0_2),.clk(gclk));
	jand g388(.dina(w_b65_0[1]),.dinb(w_a65_0[1]),.dout(n774),.clk(gclk));
	jcb g389(.dina(w_b65_0[0]),.dinb(w_a65_0[0]),.dout(n775));
	jand g390(.dina(w_dff_B_CuQ7QQJA6_0),.dinb(w_n771_0[0]),.dout(n776),.clk(gclk));
	jcb g391(.dina(n776),.dinb(w_dff_B_NsY7JH502_1),.dout(n777));
	jxor g392(.dina(w_b66_0[2]),.dinb(w_a66_0[2]),.dout(n778),.clk(gclk));
	jxor g393(.dina(w_dff_B_wTQtsp8q0_0),.dinb(w_n777_0[1]),.dout(w_dff_A_u9JR45Q39_2),.clk(gclk));
	jand g394(.dina(w_b66_0[1]),.dinb(w_a66_0[1]),.dout(n780),.clk(gclk));
	jcb g395(.dina(w_b66_0[0]),.dinb(w_a66_0[0]),.dout(n781));
	jand g396(.dina(w_dff_B_Mcr16eGs4_0),.dinb(w_n777_0[0]),.dout(n782),.clk(gclk));
	jcb g397(.dina(n782),.dinb(w_dff_B_SvQrjUup5_1),.dout(n783));
	jxor g398(.dina(w_b67_0[2]),.dinb(w_a67_0[2]),.dout(n784),.clk(gclk));
	jxor g399(.dina(w_dff_B_lE4zQQav5_0),.dinb(w_n783_0[1]),.dout(w_dff_A_Z4pRlS9P8_2),.clk(gclk));
	jand g400(.dina(w_b67_0[1]),.dinb(w_a67_0[1]),.dout(n786),.clk(gclk));
	jcb g401(.dina(w_b67_0[0]),.dinb(w_a67_0[0]),.dout(n787));
	jand g402(.dina(w_dff_B_bDbh5nUT3_0),.dinb(w_n783_0[0]),.dout(n788),.clk(gclk));
	jcb g403(.dina(n788),.dinb(w_dff_B_cSmyQJfw1_1),.dout(n789));
	jxor g404(.dina(w_b68_0[2]),.dinb(w_a68_0[2]),.dout(n790),.clk(gclk));
	jxor g405(.dina(w_dff_B_svBcB5FP3_0),.dinb(w_n789_0[1]),.dout(w_dff_A_RBUkAX7b8_2),.clk(gclk));
	jand g406(.dina(w_b68_0[1]),.dinb(w_a68_0[1]),.dout(n792),.clk(gclk));
	jcb g407(.dina(w_b68_0[0]),.dinb(w_a68_0[0]),.dout(n793));
	jand g408(.dina(w_dff_B_2OXQnYqp2_0),.dinb(w_n789_0[0]),.dout(n794),.clk(gclk));
	jcb g409(.dina(n794),.dinb(w_dff_B_qVRyJbno5_1),.dout(n795));
	jxor g410(.dina(w_b69_0[2]),.dinb(w_a69_0[2]),.dout(n796),.clk(gclk));
	jxor g411(.dina(w_dff_B_IIZIbszu3_0),.dinb(w_n795_0[1]),.dout(w_dff_A_VF0Og0Ap9_2),.clk(gclk));
	jand g412(.dina(w_b69_0[1]),.dinb(w_a69_0[1]),.dout(n798),.clk(gclk));
	jcb g413(.dina(w_b69_0[0]),.dinb(w_a69_0[0]),.dout(n799));
	jand g414(.dina(w_dff_B_iAHi3cHM6_0),.dinb(w_n795_0[0]),.dout(n800),.clk(gclk));
	jcb g415(.dina(n800),.dinb(w_dff_B_7PPvMfFA7_1),.dout(n801));
	jxor g416(.dina(w_b70_0[2]),.dinb(w_a70_0[2]),.dout(n802),.clk(gclk));
	jxor g417(.dina(w_dff_B_ikvCzPGE3_0),.dinb(w_n801_0[1]),.dout(w_dff_A_uaH4n4Vl7_2),.clk(gclk));
	jand g418(.dina(w_b70_0[1]),.dinb(w_a70_0[1]),.dout(n804),.clk(gclk));
	jcb g419(.dina(w_b70_0[0]),.dinb(w_a70_0[0]),.dout(n805));
	jand g420(.dina(w_dff_B_ok8xe67Q0_0),.dinb(w_n801_0[0]),.dout(n806),.clk(gclk));
	jcb g421(.dina(n806),.dinb(w_dff_B_pVF4M0wG0_1),.dout(n807));
	jxor g422(.dina(w_b71_0[2]),.dinb(w_a71_0[2]),.dout(n808),.clk(gclk));
	jxor g423(.dina(w_dff_B_JxWKhrsd3_0),.dinb(w_n807_0[1]),.dout(w_dff_A_25rg4D9y4_2),.clk(gclk));
	jand g424(.dina(w_b71_0[1]),.dinb(w_a71_0[1]),.dout(n810),.clk(gclk));
	jcb g425(.dina(w_b71_0[0]),.dinb(w_a71_0[0]),.dout(n811));
	jand g426(.dina(w_dff_B_opoKmvzR0_0),.dinb(w_n807_0[0]),.dout(n812),.clk(gclk));
	jcb g427(.dina(n812),.dinb(w_dff_B_2xeLz8H77_1),.dout(n813));
	jxor g428(.dina(w_b72_0[2]),.dinb(w_a72_0[2]),.dout(n814),.clk(gclk));
	jxor g429(.dina(w_dff_B_pv3sBp5K2_0),.dinb(w_n813_0[1]),.dout(w_dff_A_DAfWDgLl4_2),.clk(gclk));
	jand g430(.dina(w_b72_0[1]),.dinb(w_a72_0[1]),.dout(n816),.clk(gclk));
	jcb g431(.dina(w_b72_0[0]),.dinb(w_a72_0[0]),.dout(n817));
	jand g432(.dina(w_dff_B_FLEVHsvk5_0),.dinb(w_n813_0[0]),.dout(n818),.clk(gclk));
	jcb g433(.dina(n818),.dinb(w_dff_B_CmLHlizM1_1),.dout(n819));
	jxor g434(.dina(w_b73_0[2]),.dinb(w_a73_0[2]),.dout(n820),.clk(gclk));
	jxor g435(.dina(w_dff_B_FMC2ALGB0_0),.dinb(w_n819_0[1]),.dout(w_dff_A_EXeMsU4S3_2),.clk(gclk));
	jand g436(.dina(w_b73_0[1]),.dinb(w_a73_0[1]),.dout(n822),.clk(gclk));
	jcb g437(.dina(w_b73_0[0]),.dinb(w_a73_0[0]),.dout(n823));
	jand g438(.dina(w_dff_B_rKut0M2W1_0),.dinb(w_n819_0[0]),.dout(n824),.clk(gclk));
	jcb g439(.dina(n824),.dinb(w_dff_B_yBmv7bjw0_1),.dout(n825));
	jxor g440(.dina(w_b74_0[2]),.dinb(w_a74_0[2]),.dout(n826),.clk(gclk));
	jxor g441(.dina(w_dff_B_Zb3Aui4E2_0),.dinb(w_n825_0[1]),.dout(w_dff_A_kBneCYEu8_2),.clk(gclk));
	jand g442(.dina(w_b74_0[1]),.dinb(w_a74_0[1]),.dout(n828),.clk(gclk));
	jcb g443(.dina(w_b74_0[0]),.dinb(w_a74_0[0]),.dout(n829));
	jand g444(.dina(w_dff_B_zTdSogfq8_0),.dinb(w_n825_0[0]),.dout(n830),.clk(gclk));
	jcb g445(.dina(n830),.dinb(w_dff_B_yknhl01q3_1),.dout(n831));
	jxor g446(.dina(w_b75_0[2]),.dinb(w_a75_0[2]),.dout(n832),.clk(gclk));
	jxor g447(.dina(w_dff_B_DhOwyyt05_0),.dinb(w_n831_0[1]),.dout(w_dff_A_50Y8hj8Y4_2),.clk(gclk));
	jand g448(.dina(w_b75_0[1]),.dinb(w_a75_0[1]),.dout(n834),.clk(gclk));
	jcb g449(.dina(w_b75_0[0]),.dinb(w_a75_0[0]),.dout(n835));
	jand g450(.dina(w_dff_B_eQj5PWyb8_0),.dinb(w_n831_0[0]),.dout(n836),.clk(gclk));
	jcb g451(.dina(n836),.dinb(w_dff_B_iCcYTe8i1_1),.dout(n837));
	jxor g452(.dina(w_b76_0[2]),.dinb(w_a76_0[2]),.dout(n838),.clk(gclk));
	jxor g453(.dina(w_dff_B_djJxNpry8_0),.dinb(w_n837_0[1]),.dout(w_dff_A_uKcBLu2n9_2),.clk(gclk));
	jand g454(.dina(w_b76_0[1]),.dinb(w_a76_0[1]),.dout(n840),.clk(gclk));
	jcb g455(.dina(w_b76_0[0]),.dinb(w_a76_0[0]),.dout(n841));
	jand g456(.dina(w_dff_B_ogHkkQPV9_0),.dinb(w_n837_0[0]),.dout(n842),.clk(gclk));
	jcb g457(.dina(n842),.dinb(w_dff_B_NwsfVLEn3_1),.dout(n843));
	jxor g458(.dina(w_b77_0[2]),.dinb(w_a77_0[2]),.dout(n844),.clk(gclk));
	jxor g459(.dina(w_dff_B_uNf2OqZk3_0),.dinb(w_n843_0[1]),.dout(w_dff_A_RlfpDKF12_2),.clk(gclk));
	jand g460(.dina(w_b77_0[1]),.dinb(w_a77_0[1]),.dout(n846),.clk(gclk));
	jcb g461(.dina(w_b77_0[0]),.dinb(w_a77_0[0]),.dout(n847));
	jand g462(.dina(w_dff_B_tkkHea3i0_0),.dinb(w_n843_0[0]),.dout(n848),.clk(gclk));
	jcb g463(.dina(n848),.dinb(w_dff_B_HA2BJTtt9_1),.dout(n849));
	jxor g464(.dina(w_b78_0[2]),.dinb(w_a78_0[2]),.dout(n850),.clk(gclk));
	jxor g465(.dina(w_dff_B_F5vtCGLu7_0),.dinb(w_n849_0[1]),.dout(w_dff_A_yWmtd95Z9_2),.clk(gclk));
	jand g466(.dina(w_b78_0[1]),.dinb(w_a78_0[1]),.dout(n852),.clk(gclk));
	jcb g467(.dina(w_b78_0[0]),.dinb(w_a78_0[0]),.dout(n853));
	jand g468(.dina(w_dff_B_nx8MnoHd2_0),.dinb(w_n849_0[0]),.dout(n854),.clk(gclk));
	jcb g469(.dina(n854),.dinb(w_dff_B_PPpQ5mdn1_1),.dout(n855));
	jxor g470(.dina(w_b79_0[2]),.dinb(w_a79_0[2]),.dout(n856),.clk(gclk));
	jxor g471(.dina(w_dff_B_9rEkfsRT6_0),.dinb(w_n855_0[1]),.dout(w_dff_A_iULoKlkx1_2),.clk(gclk));
	jand g472(.dina(w_b79_0[1]),.dinb(w_a79_0[1]),.dout(n858),.clk(gclk));
	jcb g473(.dina(w_b79_0[0]),.dinb(w_a79_0[0]),.dout(n859));
	jand g474(.dina(w_dff_B_OkjULAnL9_0),.dinb(w_n855_0[0]),.dout(n860),.clk(gclk));
	jcb g475(.dina(n860),.dinb(w_dff_B_sIPXzDkp4_1),.dout(n861));
	jxor g476(.dina(w_b80_0[2]),.dinb(w_a80_0[2]),.dout(n862),.clk(gclk));
	jxor g477(.dina(w_dff_B_xD0LztTD2_0),.dinb(w_n861_0[1]),.dout(w_dff_A_E95bjTHE6_2),.clk(gclk));
	jand g478(.dina(w_b80_0[1]),.dinb(w_a80_0[1]),.dout(n864),.clk(gclk));
	jcb g479(.dina(w_b80_0[0]),.dinb(w_a80_0[0]),.dout(n865));
	jand g480(.dina(w_dff_B_MhnprG8l9_0),.dinb(w_n861_0[0]),.dout(n866),.clk(gclk));
	jcb g481(.dina(n866),.dinb(w_dff_B_e84DdMJl5_1),.dout(n867));
	jxor g482(.dina(w_b81_0[2]),.dinb(w_a81_0[2]),.dout(n868),.clk(gclk));
	jxor g483(.dina(w_dff_B_kZscPfF05_0),.dinb(w_n867_0[1]),.dout(w_dff_A_5ajlcE7V4_2),.clk(gclk));
	jand g484(.dina(w_b81_0[1]),.dinb(w_a81_0[1]),.dout(n870),.clk(gclk));
	jcb g485(.dina(w_b81_0[0]),.dinb(w_a81_0[0]),.dout(n871));
	jand g486(.dina(w_dff_B_JvDs4JAs1_0),.dinb(w_n867_0[0]),.dout(n872),.clk(gclk));
	jcb g487(.dina(n872),.dinb(w_dff_B_tvjawTBP1_1),.dout(n873));
	jxor g488(.dina(w_b82_0[2]),.dinb(w_a82_0[2]),.dout(n874),.clk(gclk));
	jxor g489(.dina(w_dff_B_pbwwiBwO7_0),.dinb(w_n873_0[1]),.dout(w_dff_A_Xic2Adtu8_2),.clk(gclk));
	jand g490(.dina(w_b82_0[1]),.dinb(w_a82_0[1]),.dout(n876),.clk(gclk));
	jcb g491(.dina(w_b82_0[0]),.dinb(w_a82_0[0]),.dout(n877));
	jand g492(.dina(w_dff_B_kq0cFdQ24_0),.dinb(w_n873_0[0]),.dout(n878),.clk(gclk));
	jcb g493(.dina(n878),.dinb(w_dff_B_GzgJUVn93_1),.dout(n879));
	jxor g494(.dina(w_b83_0[2]),.dinb(w_a83_0[2]),.dout(n880),.clk(gclk));
	jxor g495(.dina(w_dff_B_bMIFxpYM3_0),.dinb(w_n879_0[1]),.dout(w_dff_A_4p69wJXZ0_2),.clk(gclk));
	jand g496(.dina(w_b83_0[1]),.dinb(w_a83_0[1]),.dout(n882),.clk(gclk));
	jcb g497(.dina(w_b83_0[0]),.dinb(w_a83_0[0]),.dout(n883));
	jand g498(.dina(w_dff_B_XuAALr0W2_0),.dinb(w_n879_0[0]),.dout(n884),.clk(gclk));
	jcb g499(.dina(n884),.dinb(w_dff_B_pqpOHVfn2_1),.dout(n885));
	jxor g500(.dina(w_b84_0[2]),.dinb(w_a84_0[2]),.dout(n886),.clk(gclk));
	jxor g501(.dina(w_dff_B_zUsR3Qhs2_0),.dinb(w_n885_0[1]),.dout(w_dff_A_BzE0H6ap0_2),.clk(gclk));
	jand g502(.dina(w_b84_0[1]),.dinb(w_a84_0[1]),.dout(n888),.clk(gclk));
	jcb g503(.dina(w_b84_0[0]),.dinb(w_a84_0[0]),.dout(n889));
	jand g504(.dina(w_dff_B_mRYvO6bw1_0),.dinb(w_n885_0[0]),.dout(n890),.clk(gclk));
	jcb g505(.dina(n890),.dinb(w_dff_B_etx97ig43_1),.dout(n891));
	jxor g506(.dina(w_b85_0[2]),.dinb(w_a85_0[2]),.dout(n892),.clk(gclk));
	jxor g507(.dina(w_dff_B_tgwVYjIg3_0),.dinb(w_n891_0[1]),.dout(w_dff_A_TrXEhtji4_2),.clk(gclk));
	jand g508(.dina(w_b85_0[1]),.dinb(w_a85_0[1]),.dout(n894),.clk(gclk));
	jcb g509(.dina(w_b85_0[0]),.dinb(w_a85_0[0]),.dout(n895));
	jand g510(.dina(w_dff_B_LbDxoEnS2_0),.dinb(w_n891_0[0]),.dout(n896),.clk(gclk));
	jcb g511(.dina(n896),.dinb(w_dff_B_8UlPWcMp1_1),.dout(n897));
	jxor g512(.dina(w_b86_0[2]),.dinb(w_a86_0[2]),.dout(n898),.clk(gclk));
	jxor g513(.dina(w_dff_B_EZvSDj9R9_0),.dinb(w_n897_0[1]),.dout(w_dff_A_HRCPkfMi4_2),.clk(gclk));
	jand g514(.dina(w_b86_0[1]),.dinb(w_a86_0[1]),.dout(n900),.clk(gclk));
	jcb g515(.dina(w_b86_0[0]),.dinb(w_a86_0[0]),.dout(n901));
	jand g516(.dina(w_dff_B_f56FFK1t6_0),.dinb(w_n897_0[0]),.dout(n902),.clk(gclk));
	jcb g517(.dina(n902),.dinb(w_dff_B_epsTtTK93_1),.dout(n903));
	jxor g518(.dina(w_b87_0[2]),.dinb(w_a87_0[2]),.dout(n904),.clk(gclk));
	jxor g519(.dina(w_dff_B_uUkfOFQn1_0),.dinb(w_n903_0[1]),.dout(w_dff_A_OCpaXqst8_2),.clk(gclk));
	jand g520(.dina(w_b87_0[1]),.dinb(w_a87_0[1]),.dout(n906),.clk(gclk));
	jcb g521(.dina(w_b87_0[0]),.dinb(w_a87_0[0]),.dout(n907));
	jand g522(.dina(w_dff_B_dfcAYDfk0_0),.dinb(w_n903_0[0]),.dout(n908),.clk(gclk));
	jcb g523(.dina(n908),.dinb(w_dff_B_utDSKdr27_1),.dout(n909));
	jxor g524(.dina(w_b88_0[2]),.dinb(w_a88_0[2]),.dout(n910),.clk(gclk));
	jxor g525(.dina(w_dff_B_ynh2rDWK5_0),.dinb(w_n909_0[1]),.dout(w_dff_A_LDFLxawb9_2),.clk(gclk));
	jand g526(.dina(w_b88_0[1]),.dinb(w_a88_0[1]),.dout(n912),.clk(gclk));
	jcb g527(.dina(w_b88_0[0]),.dinb(w_a88_0[0]),.dout(n913));
	jand g528(.dina(w_dff_B_N7vmbMkQ0_0),.dinb(w_n909_0[0]),.dout(n914),.clk(gclk));
	jcb g529(.dina(n914),.dinb(w_dff_B_brSNaHyt4_1),.dout(n915));
	jxor g530(.dina(w_b89_0[2]),.dinb(w_a89_0[2]),.dout(n916),.clk(gclk));
	jxor g531(.dina(w_dff_B_HLQWv4eU2_0),.dinb(w_n915_0[1]),.dout(w_dff_A_6JucvmkC3_2),.clk(gclk));
	jand g532(.dina(w_b89_0[1]),.dinb(w_a89_0[1]),.dout(n918),.clk(gclk));
	jcb g533(.dina(w_b89_0[0]),.dinb(w_a89_0[0]),.dout(n919));
	jand g534(.dina(w_dff_B_AOA64WTK7_0),.dinb(w_n915_0[0]),.dout(n920),.clk(gclk));
	jcb g535(.dina(n920),.dinb(w_dff_B_fXOzDmTA4_1),.dout(n921));
	jxor g536(.dina(w_b90_0[2]),.dinb(w_a90_0[2]),.dout(n922),.clk(gclk));
	jxor g537(.dina(w_dff_B_jeAaxdpn6_0),.dinb(w_n921_0[1]),.dout(w_dff_A_7kDqg9E90_2),.clk(gclk));
	jand g538(.dina(w_b90_0[1]),.dinb(w_a90_0[1]),.dout(n924),.clk(gclk));
	jcb g539(.dina(w_b90_0[0]),.dinb(w_a90_0[0]),.dout(n925));
	jand g540(.dina(w_dff_B_wsbERzgk2_0),.dinb(w_n921_0[0]),.dout(n926),.clk(gclk));
	jcb g541(.dina(n926),.dinb(w_dff_B_8T9xx6qV1_1),.dout(n927));
	jxor g542(.dina(w_b91_0[2]),.dinb(w_a91_0[2]),.dout(n928),.clk(gclk));
	jxor g543(.dina(w_dff_B_vgkiyEAh6_0),.dinb(w_n927_0[1]),.dout(w_dff_A_oKzz53IO5_2),.clk(gclk));
	jand g544(.dina(w_b91_0[1]),.dinb(w_a91_0[1]),.dout(n930),.clk(gclk));
	jcb g545(.dina(w_b91_0[0]),.dinb(w_a91_0[0]),.dout(n931));
	jand g546(.dina(w_dff_B_yQ9eGirj0_0),.dinb(w_n927_0[0]),.dout(n932),.clk(gclk));
	jcb g547(.dina(n932),.dinb(w_dff_B_eoY4eUdu5_1),.dout(n933));
	jxor g548(.dina(w_b92_0[2]),.dinb(w_a92_0[2]),.dout(n934),.clk(gclk));
	jxor g549(.dina(w_dff_B_lJOSsY171_0),.dinb(w_n933_0[1]),.dout(w_dff_A_AEzxCK512_2),.clk(gclk));
	jand g550(.dina(w_b92_0[1]),.dinb(w_a92_0[1]),.dout(n936),.clk(gclk));
	jcb g551(.dina(w_b92_0[0]),.dinb(w_a92_0[0]),.dout(n937));
	jand g552(.dina(w_dff_B_2tpIruTy5_0),.dinb(w_n933_0[0]),.dout(n938),.clk(gclk));
	jcb g553(.dina(n938),.dinb(w_dff_B_Vnmk2IHa8_1),.dout(n939));
	jxor g554(.dina(w_b93_0[2]),.dinb(w_a93_0[2]),.dout(n940),.clk(gclk));
	jxor g555(.dina(w_dff_B_pbghLIdh4_0),.dinb(w_n939_0[1]),.dout(w_dff_A_Er2L8DHW9_2),.clk(gclk));
	jand g556(.dina(w_b93_0[1]),.dinb(w_a93_0[1]),.dout(n942),.clk(gclk));
	jcb g557(.dina(w_b93_0[0]),.dinb(w_a93_0[0]),.dout(n943));
	jand g558(.dina(w_dff_B_Z53VFgFh4_0),.dinb(w_n939_0[0]),.dout(n944),.clk(gclk));
	jcb g559(.dina(n944),.dinb(w_dff_B_qRRscppg1_1),.dout(n945));
	jxor g560(.dina(w_b94_0[2]),.dinb(w_a94_0[2]),.dout(n946),.clk(gclk));
	jxor g561(.dina(w_dff_B_NYqGAdoD6_0),.dinb(w_n945_0[1]),.dout(w_dff_A_XtJDEDOj6_2),.clk(gclk));
	jand g562(.dina(w_b94_0[1]),.dinb(w_a94_0[1]),.dout(n948),.clk(gclk));
	jcb g563(.dina(w_b94_0[0]),.dinb(w_a94_0[0]),.dout(n949));
	jand g564(.dina(w_dff_B_Tlk8jcgs4_0),.dinb(w_n945_0[0]),.dout(n950),.clk(gclk));
	jcb g565(.dina(n950),.dinb(w_dff_B_gjoULGb32_1),.dout(n951));
	jxor g566(.dina(w_b95_0[2]),.dinb(w_a95_0[2]),.dout(n952),.clk(gclk));
	jxor g567(.dina(w_dff_B_q5yKBMhs4_0),.dinb(w_n951_0[1]),.dout(w_dff_A_AMFRU9o10_2),.clk(gclk));
	jand g568(.dina(w_b95_0[1]),.dinb(w_a95_0[1]),.dout(n954),.clk(gclk));
	jcb g569(.dina(w_b95_0[0]),.dinb(w_a95_0[0]),.dout(n955));
	jand g570(.dina(w_dff_B_gF4cW8n67_0),.dinb(w_n951_0[0]),.dout(n956),.clk(gclk));
	jcb g571(.dina(n956),.dinb(w_dff_B_Jf6mJkjd5_1),.dout(n957));
	jxor g572(.dina(w_b96_0[2]),.dinb(w_a96_0[2]),.dout(n958),.clk(gclk));
	jxor g573(.dina(w_dff_B_o3ojjpxb8_0),.dinb(w_n957_0[1]),.dout(w_dff_A_4HZtpbSH1_2),.clk(gclk));
	jand g574(.dina(w_b96_0[1]),.dinb(w_a96_0[1]),.dout(n960),.clk(gclk));
	jcb g575(.dina(w_b96_0[0]),.dinb(w_a96_0[0]),.dout(n961));
	jand g576(.dina(w_dff_B_3XsPByS46_0),.dinb(w_n957_0[0]),.dout(n962),.clk(gclk));
	jcb g577(.dina(n962),.dinb(w_dff_B_i16ixeFE0_1),.dout(n963));
	jxor g578(.dina(w_b97_0[2]),.dinb(w_a97_0[2]),.dout(n964),.clk(gclk));
	jxor g579(.dina(w_dff_B_IwDOjdtB9_0),.dinb(w_n963_0[1]),.dout(w_dff_A_LhBO705X1_2),.clk(gclk));
	jand g580(.dina(w_b97_0[1]),.dinb(w_a97_0[1]),.dout(n966),.clk(gclk));
	jcb g581(.dina(w_b97_0[0]),.dinb(w_a97_0[0]),.dout(n967));
	jand g582(.dina(w_dff_B_XE2iBHU27_0),.dinb(w_n963_0[0]),.dout(n968),.clk(gclk));
	jcb g583(.dina(n968),.dinb(w_dff_B_WB80gDUQ3_1),.dout(n969));
	jxor g584(.dina(w_b98_0[2]),.dinb(w_a98_0[2]),.dout(n970),.clk(gclk));
	jxor g585(.dina(w_dff_B_vwMgjcE08_0),.dinb(w_n969_0[1]),.dout(w_dff_A_rQuWRbM25_2),.clk(gclk));
	jand g586(.dina(w_b98_0[1]),.dinb(w_a98_0[1]),.dout(n972),.clk(gclk));
	jcb g587(.dina(w_b98_0[0]),.dinb(w_a98_0[0]),.dout(n973));
	jand g588(.dina(w_dff_B_CzElqIeo4_0),.dinb(w_n969_0[0]),.dout(n974),.clk(gclk));
	jcb g589(.dina(n974),.dinb(w_dff_B_sukvz7S18_1),.dout(n975));
	jxor g590(.dina(w_b99_0[2]),.dinb(w_a99_0[2]),.dout(n976),.clk(gclk));
	jxor g591(.dina(w_dff_B_M3z591OZ9_0),.dinb(w_n975_0[1]),.dout(w_dff_A_jth7tJDE4_2),.clk(gclk));
	jand g592(.dina(w_b99_0[1]),.dinb(w_a99_0[1]),.dout(n978),.clk(gclk));
	jcb g593(.dina(w_b99_0[0]),.dinb(w_a99_0[0]),.dout(n979));
	jand g594(.dina(w_dff_B_wOyfHYTt8_0),.dinb(w_n975_0[0]),.dout(n980),.clk(gclk));
	jcb g595(.dina(n980),.dinb(w_dff_B_miF1RlLv4_1),.dout(n981));
	jxor g596(.dina(w_b100_0[2]),.dinb(w_a100_0[2]),.dout(n982),.clk(gclk));
	jxor g597(.dina(w_dff_B_hGgjVT1m4_0),.dinb(w_n981_0[1]),.dout(w_dff_A_vGnqaJJF9_2),.clk(gclk));
	jand g598(.dina(w_b100_0[1]),.dinb(w_a100_0[1]),.dout(n984),.clk(gclk));
	jcb g599(.dina(w_b100_0[0]),.dinb(w_a100_0[0]),.dout(n985));
	jand g600(.dina(w_dff_B_ZBeU3nCK4_0),.dinb(w_n981_0[0]),.dout(n986),.clk(gclk));
	jcb g601(.dina(n986),.dinb(w_dff_B_ihOKXM3G5_1),.dout(n987));
	jxor g602(.dina(w_b101_0[2]),.dinb(w_a101_0[2]),.dout(n988),.clk(gclk));
	jxor g603(.dina(w_dff_B_Rw2JWE0p7_0),.dinb(w_n987_0[1]),.dout(w_dff_A_Fj4n1Rkq2_2),.clk(gclk));
	jand g604(.dina(w_b101_0[1]),.dinb(w_a101_0[1]),.dout(n990),.clk(gclk));
	jcb g605(.dina(w_b101_0[0]),.dinb(w_a101_0[0]),.dout(n991));
	jand g606(.dina(w_dff_B_WKYHnQ064_0),.dinb(w_n987_0[0]),.dout(n992),.clk(gclk));
	jcb g607(.dina(n992),.dinb(w_dff_B_eOrMuw528_1),.dout(n993));
	jxor g608(.dina(w_b102_0[2]),.dinb(w_a102_0[2]),.dout(n994),.clk(gclk));
	jxor g609(.dina(w_dff_B_YeW3yzi12_0),.dinb(w_n993_0[1]),.dout(w_dff_A_P3vaBdYA9_2),.clk(gclk));
	jand g610(.dina(w_b102_0[1]),.dinb(w_a102_0[1]),.dout(n996),.clk(gclk));
	jcb g611(.dina(w_b102_0[0]),.dinb(w_a102_0[0]),.dout(n997));
	jand g612(.dina(w_dff_B_MNe3cJhP9_0),.dinb(w_n993_0[0]),.dout(n998),.clk(gclk));
	jcb g613(.dina(n998),.dinb(w_dff_B_CTOAbFb57_1),.dout(n999));
	jxor g614(.dina(w_b103_0[2]),.dinb(w_a103_0[2]),.dout(n1000),.clk(gclk));
	jxor g615(.dina(w_dff_B_aQY9Vmue7_0),.dinb(w_n999_0[1]),.dout(w_dff_A_XMlybQoI8_2),.clk(gclk));
	jand g616(.dina(w_b103_0[1]),.dinb(w_a103_0[1]),.dout(n1002),.clk(gclk));
	jcb g617(.dina(w_b103_0[0]),.dinb(w_a103_0[0]),.dout(n1003));
	jand g618(.dina(w_dff_B_ISBRX9kG4_0),.dinb(w_n999_0[0]),.dout(n1004),.clk(gclk));
	jcb g619(.dina(n1004),.dinb(w_dff_B_GI8cjqgr1_1),.dout(n1005));
	jxor g620(.dina(w_b104_0[2]),.dinb(w_a104_0[2]),.dout(n1006),.clk(gclk));
	jxor g621(.dina(w_dff_B_pmoeat4U0_0),.dinb(w_n1005_0[1]),.dout(w_dff_A_5ieeOtHr7_2),.clk(gclk));
	jand g622(.dina(w_b104_0[1]),.dinb(w_a104_0[1]),.dout(n1008),.clk(gclk));
	jcb g623(.dina(w_b104_0[0]),.dinb(w_a104_0[0]),.dout(n1009));
	jand g624(.dina(w_dff_B_lEwdgnFZ1_0),.dinb(w_n1005_0[0]),.dout(n1010),.clk(gclk));
	jcb g625(.dina(n1010),.dinb(w_dff_B_8BuCOaXp1_1),.dout(n1011));
	jxor g626(.dina(w_b105_0[2]),.dinb(w_a105_0[2]),.dout(n1012),.clk(gclk));
	jxor g627(.dina(w_dff_B_73IF7KRg3_0),.dinb(w_n1011_0[1]),.dout(w_dff_A_ZOM6W9LV4_2),.clk(gclk));
	jand g628(.dina(w_b105_0[1]),.dinb(w_a105_0[1]),.dout(n1014),.clk(gclk));
	jcb g629(.dina(w_b105_0[0]),.dinb(w_a105_0[0]),.dout(n1015));
	jand g630(.dina(w_dff_B_IzQy6DU01_0),.dinb(w_n1011_0[0]),.dout(n1016),.clk(gclk));
	jcb g631(.dina(n1016),.dinb(w_dff_B_opUbMGB49_1),.dout(n1017));
	jxor g632(.dina(w_b106_0[2]),.dinb(w_a106_0[2]),.dout(n1018),.clk(gclk));
	jxor g633(.dina(w_dff_B_iiL6A9U45_0),.dinb(w_n1017_0[1]),.dout(w_dff_A_URhuMiJa9_2),.clk(gclk));
	jand g634(.dina(w_b106_0[1]),.dinb(w_a106_0[1]),.dout(n1020),.clk(gclk));
	jcb g635(.dina(w_b106_0[0]),.dinb(w_a106_0[0]),.dout(n1021));
	jand g636(.dina(w_dff_B_OmEewm5z6_0),.dinb(w_n1017_0[0]),.dout(n1022),.clk(gclk));
	jcb g637(.dina(n1022),.dinb(w_dff_B_P8u9UvcR2_1),.dout(n1023));
	jxor g638(.dina(w_b107_0[2]),.dinb(w_a107_0[2]),.dout(n1024),.clk(gclk));
	jxor g639(.dina(w_dff_B_T2YmP8GL7_0),.dinb(w_n1023_0[1]),.dout(w_dff_A_cwkY2DxV9_2),.clk(gclk));
	jand g640(.dina(w_b107_0[1]),.dinb(w_a107_0[1]),.dout(n1026),.clk(gclk));
	jcb g641(.dina(w_b107_0[0]),.dinb(w_a107_0[0]),.dout(n1027));
	jand g642(.dina(w_dff_B_rQs1ywwY3_0),.dinb(w_n1023_0[0]),.dout(n1028),.clk(gclk));
	jcb g643(.dina(n1028),.dinb(w_dff_B_XTpaCHU28_1),.dout(n1029));
	jxor g644(.dina(w_b108_0[2]),.dinb(w_a108_0[2]),.dout(n1030),.clk(gclk));
	jxor g645(.dina(w_dff_B_dd0p0oAi6_0),.dinb(w_n1029_0[1]),.dout(w_dff_A_aQI6d3Nn2_2),.clk(gclk));
	jand g646(.dina(w_b108_0[1]),.dinb(w_a108_0[1]),.dout(n1032),.clk(gclk));
	jcb g647(.dina(w_b108_0[0]),.dinb(w_a108_0[0]),.dout(n1033));
	jand g648(.dina(w_dff_B_ISqqPwDn9_0),.dinb(w_n1029_0[0]),.dout(n1034),.clk(gclk));
	jcb g649(.dina(n1034),.dinb(w_dff_B_BMacVM8n4_1),.dout(n1035));
	jxor g650(.dina(w_b109_0[2]),.dinb(w_a109_0[2]),.dout(n1036),.clk(gclk));
	jxor g651(.dina(w_dff_B_k9DFeDPe2_0),.dinb(w_n1035_0[1]),.dout(w_dff_A_6RAzsJrE3_2),.clk(gclk));
	jand g652(.dina(w_b109_0[1]),.dinb(w_a109_0[1]),.dout(n1038),.clk(gclk));
	jcb g653(.dina(w_b109_0[0]),.dinb(w_a109_0[0]),.dout(n1039));
	jand g654(.dina(w_dff_B_C9QaqcpL4_0),.dinb(w_n1035_0[0]),.dout(n1040),.clk(gclk));
	jcb g655(.dina(n1040),.dinb(w_dff_B_mscM20U91_1),.dout(n1041));
	jxor g656(.dina(w_b110_0[2]),.dinb(w_a110_0[2]),.dout(n1042),.clk(gclk));
	jxor g657(.dina(w_dff_B_H2Dnf3dc2_0),.dinb(w_n1041_0[1]),.dout(w_dff_A_ukMTbJQ36_2),.clk(gclk));
	jand g658(.dina(w_b110_0[1]),.dinb(w_a110_0[1]),.dout(n1044),.clk(gclk));
	jcb g659(.dina(w_b110_0[0]),.dinb(w_a110_0[0]),.dout(n1045));
	jand g660(.dina(w_dff_B_gYw3T9cY7_0),.dinb(w_n1041_0[0]),.dout(n1046),.clk(gclk));
	jcb g661(.dina(n1046),.dinb(w_dff_B_sX8cRBX78_1),.dout(n1047));
	jxor g662(.dina(w_b111_0[2]),.dinb(w_a111_0[2]),.dout(n1048),.clk(gclk));
	jxor g663(.dina(w_dff_B_Yxb7eyNY0_0),.dinb(w_n1047_0[1]),.dout(w_dff_A_kWw534XR3_2),.clk(gclk));
	jand g664(.dina(w_b111_0[1]),.dinb(w_a111_0[1]),.dout(n1050),.clk(gclk));
	jcb g665(.dina(w_b111_0[0]),.dinb(w_a111_0[0]),.dout(n1051));
	jand g666(.dina(w_dff_B_JR5SiCzG0_0),.dinb(w_n1047_0[0]),.dout(n1052),.clk(gclk));
	jcb g667(.dina(n1052),.dinb(w_dff_B_7nEsIUQP7_1),.dout(n1053));
	jxor g668(.dina(w_b112_0[2]),.dinb(w_a112_0[2]),.dout(n1054),.clk(gclk));
	jxor g669(.dina(w_dff_B_hCzyrGpy3_0),.dinb(w_n1053_0[1]),.dout(w_dff_A_bne51yCD0_2),.clk(gclk));
	jand g670(.dina(w_b112_0[1]),.dinb(w_a112_0[1]),.dout(n1056),.clk(gclk));
	jcb g671(.dina(w_b112_0[0]),.dinb(w_a112_0[0]),.dout(n1057));
	jand g672(.dina(w_dff_B_9kk8s8Kj0_0),.dinb(w_n1053_0[0]),.dout(n1058),.clk(gclk));
	jcb g673(.dina(n1058),.dinb(w_dff_B_3fsHmRIV7_1),.dout(n1059));
	jxor g674(.dina(w_b113_0[2]),.dinb(w_a113_0[2]),.dout(n1060),.clk(gclk));
	jxor g675(.dina(w_dff_B_xwHJtFQ73_0),.dinb(w_n1059_0[1]),.dout(w_dff_A_3U7JlSNO5_2),.clk(gclk));
	jand g676(.dina(w_b113_0[1]),.dinb(w_a113_0[1]),.dout(n1062),.clk(gclk));
	jcb g677(.dina(w_b113_0[0]),.dinb(w_a113_0[0]),.dout(n1063));
	jand g678(.dina(w_dff_B_mK9qdiWp4_0),.dinb(w_n1059_0[0]),.dout(n1064),.clk(gclk));
	jcb g679(.dina(n1064),.dinb(w_dff_B_XYc0K6132_1),.dout(n1065));
	jxor g680(.dina(w_b114_0[2]),.dinb(w_a114_0[2]),.dout(n1066),.clk(gclk));
	jxor g681(.dina(w_dff_B_qONrkGfY1_0),.dinb(w_n1065_0[1]),.dout(w_dff_A_3VmB04UB2_2),.clk(gclk));
	jand g682(.dina(w_b114_0[1]),.dinb(w_a114_0[1]),.dout(n1068),.clk(gclk));
	jcb g683(.dina(w_b114_0[0]),.dinb(w_a114_0[0]),.dout(n1069));
	jand g684(.dina(w_dff_B_ImrDGPBo9_0),.dinb(w_n1065_0[0]),.dout(n1070),.clk(gclk));
	jcb g685(.dina(n1070),.dinb(w_dff_B_SjyTVPLT6_1),.dout(n1071));
	jxor g686(.dina(w_b115_0[2]),.dinb(w_a115_0[2]),.dout(n1072),.clk(gclk));
	jxor g687(.dina(w_dff_B_5DCwVdQC5_0),.dinb(w_n1071_0[1]),.dout(w_dff_A_3bA8xD5P2_2),.clk(gclk));
	jand g688(.dina(w_b115_0[1]),.dinb(w_a115_0[1]),.dout(n1074),.clk(gclk));
	jcb g689(.dina(w_b115_0[0]),.dinb(w_a115_0[0]),.dout(n1075));
	jand g690(.dina(w_dff_B_ihbYCldo3_0),.dinb(w_n1071_0[0]),.dout(n1076),.clk(gclk));
	jcb g691(.dina(n1076),.dinb(w_dff_B_DmeXqhOy3_1),.dout(n1077));
	jxor g692(.dina(w_b116_0[2]),.dinb(w_a116_0[2]),.dout(n1078),.clk(gclk));
	jxor g693(.dina(w_dff_B_t66iQooO7_0),.dinb(w_n1077_0[1]),.dout(w_dff_A_fKN0jFwO9_2),.clk(gclk));
	jand g694(.dina(w_b116_0[1]),.dinb(w_a116_0[1]),.dout(n1080),.clk(gclk));
	jcb g695(.dina(w_b116_0[0]),.dinb(w_a116_0[0]),.dout(n1081));
	jand g696(.dina(w_dff_B_k7K9XKQ61_0),.dinb(w_n1077_0[0]),.dout(n1082),.clk(gclk));
	jcb g697(.dina(n1082),.dinb(w_dff_B_0nN0BSNX5_1),.dout(n1083));
	jxor g698(.dina(w_b117_0[2]),.dinb(w_a117_0[2]),.dout(n1084),.clk(gclk));
	jxor g699(.dina(w_dff_B_Y58xZaMx0_0),.dinb(w_n1083_0[1]),.dout(w_dff_A_llLQJvtS3_2),.clk(gclk));
	jand g700(.dina(w_b117_0[1]),.dinb(w_a117_0[1]),.dout(n1086),.clk(gclk));
	jcb g701(.dina(w_b117_0[0]),.dinb(w_a117_0[0]),.dout(n1087));
	jand g702(.dina(w_dff_B_YHtR4fi00_0),.dinb(w_n1083_0[0]),.dout(n1088),.clk(gclk));
	jcb g703(.dina(n1088),.dinb(w_dff_B_Pe1iiYr60_1),.dout(n1089));
	jxor g704(.dina(w_b118_0[2]),.dinb(w_a118_0[2]),.dout(n1090),.clk(gclk));
	jxor g705(.dina(w_dff_B_M7vRvPIA2_0),.dinb(w_n1089_0[1]),.dout(w_dff_A_9UxeUz0e4_2),.clk(gclk));
	jand g706(.dina(w_b118_0[1]),.dinb(w_a118_0[1]),.dout(n1092),.clk(gclk));
	jcb g707(.dina(w_b118_0[0]),.dinb(w_a118_0[0]),.dout(n1093));
	jand g708(.dina(w_dff_B_PG2MTWyb5_0),.dinb(w_n1089_0[0]),.dout(n1094),.clk(gclk));
	jcb g709(.dina(n1094),.dinb(w_dff_B_hW63y0Sx4_1),.dout(n1095));
	jxor g710(.dina(w_b119_0[2]),.dinb(w_a119_0[2]),.dout(n1096),.clk(gclk));
	jxor g711(.dina(w_dff_B_f5k0RJ456_0),.dinb(w_n1095_0[1]),.dout(w_dff_A_VEKg84Oy2_2),.clk(gclk));
	jand g712(.dina(w_b119_0[1]),.dinb(w_a119_0[1]),.dout(n1098),.clk(gclk));
	jcb g713(.dina(w_b119_0[0]),.dinb(w_a119_0[0]),.dout(n1099));
	jand g714(.dina(w_dff_B_JSc81Qhc2_0),.dinb(w_n1095_0[0]),.dout(n1100),.clk(gclk));
	jcb g715(.dina(n1100),.dinb(w_dff_B_UxHmoAjS1_1),.dout(n1101));
	jxor g716(.dina(w_b120_0[2]),.dinb(w_a120_0[2]),.dout(n1102),.clk(gclk));
	jxor g717(.dina(w_dff_B_EPxWfQPV7_0),.dinb(w_n1101_0[1]),.dout(w_dff_A_qLw4TMU81_2),.clk(gclk));
	jand g718(.dina(w_b120_0[1]),.dinb(w_a120_0[1]),.dout(n1104),.clk(gclk));
	jcb g719(.dina(w_b120_0[0]),.dinb(w_a120_0[0]),.dout(n1105));
	jand g720(.dina(w_dff_B_urlYAJ559_0),.dinb(w_n1101_0[0]),.dout(n1106),.clk(gclk));
	jcb g721(.dina(n1106),.dinb(w_dff_B_1R6I2MTe0_1),.dout(n1107));
	jxor g722(.dina(w_b121_0[2]),.dinb(w_a121_0[2]),.dout(n1108),.clk(gclk));
	jxor g723(.dina(w_dff_B_qhYwhaxn2_0),.dinb(w_n1107_0[1]),.dout(w_dff_A_72ECXwuX6_2),.clk(gclk));
	jand g724(.dina(w_b121_0[1]),.dinb(w_a121_0[1]),.dout(n1110),.clk(gclk));
	jcb g725(.dina(w_b121_0[0]),.dinb(w_a121_0[0]),.dout(n1111));
	jand g726(.dina(w_dff_B_nEpywF7H8_0),.dinb(w_n1107_0[0]),.dout(n1112),.clk(gclk));
	jcb g727(.dina(n1112),.dinb(w_dff_B_OendyP6K5_1),.dout(n1113));
	jxor g728(.dina(w_b122_0[2]),.dinb(w_a122_0[2]),.dout(n1114),.clk(gclk));
	jxor g729(.dina(w_dff_B_sBZNRpfz4_0),.dinb(w_n1113_0[1]),.dout(w_dff_A_pUdZQfwk6_2),.clk(gclk));
	jand g730(.dina(w_b122_0[1]),.dinb(w_a122_0[1]),.dout(n1116),.clk(gclk));
	jcb g731(.dina(w_b122_0[0]),.dinb(w_a122_0[0]),.dout(n1117));
	jand g732(.dina(w_dff_B_SQmXewmR4_0),.dinb(w_n1113_0[0]),.dout(n1118),.clk(gclk));
	jcb g733(.dina(n1118),.dinb(w_dff_B_Dkr9JPcC7_1),.dout(n1119));
	jxor g734(.dina(w_b123_0[2]),.dinb(w_a123_0[2]),.dout(n1120),.clk(gclk));
	jxor g735(.dina(w_dff_B_A7qvzuar1_0),.dinb(w_n1119_0[1]),.dout(w_dff_A_njEGwhT63_2),.clk(gclk));
	jand g736(.dina(w_b123_0[1]),.dinb(w_a123_0[1]),.dout(n1122),.clk(gclk));
	jcb g737(.dina(w_b123_0[0]),.dinb(w_a123_0[0]),.dout(n1123));
	jand g738(.dina(w_dff_B_oY8pBb783_0),.dinb(w_n1119_0[0]),.dout(n1124),.clk(gclk));
	jcb g739(.dina(n1124),.dinb(w_dff_B_LkmyUViD3_1),.dout(n1125));
	jxor g740(.dina(w_b124_0[2]),.dinb(w_a124_0[2]),.dout(n1126),.clk(gclk));
	jxor g741(.dina(w_dff_B_P2qyRF8K4_0),.dinb(w_n1125_0[1]),.dout(w_dff_A_qPETohS16_2),.clk(gclk));
	jand g742(.dina(w_b124_0[1]),.dinb(w_a124_0[1]),.dout(n1128),.clk(gclk));
	jcb g743(.dina(w_b124_0[0]),.dinb(w_a124_0[0]),.dout(n1129));
	jand g744(.dina(w_dff_B_niFMbCQe5_0),.dinb(w_n1125_0[0]),.dout(n1130),.clk(gclk));
	jcb g745(.dina(n1130),.dinb(w_dff_B_WOhTpZP77_1),.dout(n1131));
	jxor g746(.dina(w_b125_0[2]),.dinb(w_a125_0[2]),.dout(n1132),.clk(gclk));
	jxor g747(.dina(w_dff_B_i84eCWYK5_0),.dinb(w_n1131_0[1]),.dout(w_dff_A_Dk9V03BL7_2),.clk(gclk));
	jand g748(.dina(w_b125_0[1]),.dinb(w_a125_0[1]),.dout(n1134),.clk(gclk));
	jcb g749(.dina(w_b125_0[0]),.dinb(w_a125_0[0]),.dout(n1135));
	jand g750(.dina(w_dff_B_B43o3NKK2_0),.dinb(w_n1131_0[0]),.dout(n1136),.clk(gclk));
	jcb g751(.dina(n1136),.dinb(w_dff_B_cdHtn6570_1),.dout(n1137));
	jxor g752(.dina(w_b126_0[2]),.dinb(w_a126_0[2]),.dout(n1138),.clk(gclk));
	jxor g753(.dina(w_dff_B_3xJzgs0k4_0),.dinb(w_n1137_0[1]),.dout(w_dff_A_e8TKNRw88_2),.clk(gclk));
	jand g754(.dina(w_b126_0[1]),.dinb(w_a126_0[1]),.dout(n1140),.clk(gclk));
	jcb g755(.dina(w_b126_0[0]),.dinb(w_a126_0[0]),.dout(n1141));
	jand g756(.dina(w_dff_B_DNEnPLV67_0),.dinb(w_n1137_0[0]),.dout(n1142),.clk(gclk));
	jcb g757(.dina(n1142),.dinb(w_dff_B_uZVHTY441_1),.dout(n1143));
	jxor g758(.dina(w_b127_0[2]),.dinb(w_a127_0[2]),.dout(n1144),.clk(gclk));
	jxor g759(.dina(w_dff_B_8Dm77OtX9_0),.dinb(w_n1143_0[1]),.dout(f127),.clk(gclk));
	jand g760(.dina(w_b127_0[1]),.dinb(w_a127_0[1]),.dout(n1146),.clk(gclk));
	jcb g761(.dina(w_b127_0[0]),.dinb(w_a127_0[0]),.dout(n1147));
	jand g762(.dina(w_dff_B_kagAjCL64_0),.dinb(w_n1143_0[0]),.dout(n1148),.clk(gclk));
	jcb g763(.dina(n1148),.dinb(w_dff_B_66p7sXjF1_1),.dout(cOut));
	jspl jspl_w_a0_0(.douta(w_a0_0[0]),.doutb(w_a0_0[1]),.din(a0));
	jspl3 jspl3_w_a1_0(.douta(w_a1_0[0]),.doutb(w_a1_0[1]),.doutc(w_a1_0[2]),.din(a1));
	jspl3 jspl3_w_a2_0(.douta(w_a2_0[0]),.doutb(w_a2_0[1]),.doutc(w_a2_0[2]),.din(a2));
	jspl3 jspl3_w_a3_0(.douta(w_a3_0[0]),.doutb(w_a3_0[1]),.doutc(w_a3_0[2]),.din(a3));
	jspl3 jspl3_w_a4_0(.douta(w_a4_0[0]),.doutb(w_a4_0[1]),.doutc(w_a4_0[2]),.din(a4));
	jspl3 jspl3_w_a5_0(.douta(w_a5_0[0]),.doutb(w_a5_0[1]),.doutc(w_a5_0[2]),.din(a5));
	jspl3 jspl3_w_a6_0(.douta(w_a6_0[0]),.doutb(w_a6_0[1]),.doutc(w_a6_0[2]),.din(a6));
	jspl3 jspl3_w_a7_0(.douta(w_a7_0[0]),.doutb(w_a7_0[1]),.doutc(w_a7_0[2]),.din(a7));
	jspl3 jspl3_w_a8_0(.douta(w_a8_0[0]),.doutb(w_a8_0[1]),.doutc(w_a8_0[2]),.din(a8));
	jspl3 jspl3_w_a9_0(.douta(w_a9_0[0]),.doutb(w_a9_0[1]),.doutc(w_a9_0[2]),.din(a9));
	jspl3 jspl3_w_a10_0(.douta(w_a10_0[0]),.doutb(w_a10_0[1]),.doutc(w_a10_0[2]),.din(a10));
	jspl3 jspl3_w_a11_0(.douta(w_a11_0[0]),.doutb(w_a11_0[1]),.doutc(w_a11_0[2]),.din(a11));
	jspl3 jspl3_w_a12_0(.douta(w_a12_0[0]),.doutb(w_a12_0[1]),.doutc(w_a12_0[2]),.din(a12));
	jspl3 jspl3_w_a13_0(.douta(w_a13_0[0]),.doutb(w_a13_0[1]),.doutc(w_a13_0[2]),.din(a13));
	jspl3 jspl3_w_a14_0(.douta(w_a14_0[0]),.doutb(w_a14_0[1]),.doutc(w_a14_0[2]),.din(a14));
	jspl3 jspl3_w_a15_0(.douta(w_a15_0[0]),.doutb(w_a15_0[1]),.doutc(w_a15_0[2]),.din(a15));
	jspl3 jspl3_w_a16_0(.douta(w_a16_0[0]),.doutb(w_a16_0[1]),.doutc(w_a16_0[2]),.din(a16));
	jspl3 jspl3_w_a17_0(.douta(w_a17_0[0]),.doutb(w_a17_0[1]),.doutc(w_a17_0[2]),.din(a17));
	jspl3 jspl3_w_a18_0(.douta(w_a18_0[0]),.doutb(w_a18_0[1]),.doutc(w_a18_0[2]),.din(a18));
	jspl3 jspl3_w_a19_0(.douta(w_a19_0[0]),.doutb(w_a19_0[1]),.doutc(w_a19_0[2]),.din(a19));
	jspl3 jspl3_w_a20_0(.douta(w_a20_0[0]),.doutb(w_a20_0[1]),.doutc(w_a20_0[2]),.din(a20));
	jspl3 jspl3_w_a21_0(.douta(w_a21_0[0]),.doutb(w_a21_0[1]),.doutc(w_a21_0[2]),.din(a21));
	jspl3 jspl3_w_a22_0(.douta(w_a22_0[0]),.doutb(w_a22_0[1]),.doutc(w_a22_0[2]),.din(a22));
	jspl3 jspl3_w_a23_0(.douta(w_a23_0[0]),.doutb(w_a23_0[1]),.doutc(w_a23_0[2]),.din(a23));
	jspl3 jspl3_w_a24_0(.douta(w_a24_0[0]),.doutb(w_a24_0[1]),.doutc(w_a24_0[2]),.din(a24));
	jspl3 jspl3_w_a25_0(.douta(w_a25_0[0]),.doutb(w_a25_0[1]),.doutc(w_a25_0[2]),.din(a25));
	jspl3 jspl3_w_a26_0(.douta(w_a26_0[0]),.doutb(w_a26_0[1]),.doutc(w_a26_0[2]),.din(a26));
	jspl3 jspl3_w_a27_0(.douta(w_a27_0[0]),.doutb(w_a27_0[1]),.doutc(w_a27_0[2]),.din(a27));
	jspl3 jspl3_w_a28_0(.douta(w_a28_0[0]),.doutb(w_a28_0[1]),.doutc(w_a28_0[2]),.din(a28));
	jspl3 jspl3_w_a29_0(.douta(w_a29_0[0]),.doutb(w_a29_0[1]),.doutc(w_a29_0[2]),.din(a29));
	jspl3 jspl3_w_a30_0(.douta(w_a30_0[0]),.doutb(w_a30_0[1]),.doutc(w_a30_0[2]),.din(a30));
	jspl3 jspl3_w_a31_0(.douta(w_a31_0[0]),.doutb(w_a31_0[1]),.doutc(w_a31_0[2]),.din(a31));
	jspl3 jspl3_w_a32_0(.douta(w_a32_0[0]),.doutb(w_a32_0[1]),.doutc(w_a32_0[2]),.din(a32));
	jspl3 jspl3_w_a33_0(.douta(w_a33_0[0]),.doutb(w_a33_0[1]),.doutc(w_a33_0[2]),.din(a33));
	jspl3 jspl3_w_a34_0(.douta(w_a34_0[0]),.doutb(w_a34_0[1]),.doutc(w_a34_0[2]),.din(a34));
	jspl3 jspl3_w_a35_0(.douta(w_a35_0[0]),.doutb(w_a35_0[1]),.doutc(w_a35_0[2]),.din(a35));
	jspl3 jspl3_w_a36_0(.douta(w_a36_0[0]),.doutb(w_a36_0[1]),.doutc(w_a36_0[2]),.din(a36));
	jspl3 jspl3_w_a37_0(.douta(w_a37_0[0]),.doutb(w_a37_0[1]),.doutc(w_a37_0[2]),.din(a37));
	jspl3 jspl3_w_a38_0(.douta(w_a38_0[0]),.doutb(w_a38_0[1]),.doutc(w_a38_0[2]),.din(a38));
	jspl3 jspl3_w_a39_0(.douta(w_a39_0[0]),.doutb(w_a39_0[1]),.doutc(w_a39_0[2]),.din(a39));
	jspl3 jspl3_w_a40_0(.douta(w_a40_0[0]),.doutb(w_a40_0[1]),.doutc(w_a40_0[2]),.din(a40));
	jspl3 jspl3_w_a41_0(.douta(w_a41_0[0]),.doutb(w_a41_0[1]),.doutc(w_a41_0[2]),.din(a41));
	jspl3 jspl3_w_a42_0(.douta(w_a42_0[0]),.doutb(w_a42_0[1]),.doutc(w_a42_0[2]),.din(a42));
	jspl3 jspl3_w_a43_0(.douta(w_a43_0[0]),.doutb(w_a43_0[1]),.doutc(w_a43_0[2]),.din(a43));
	jspl3 jspl3_w_a44_0(.douta(w_a44_0[0]),.doutb(w_a44_0[1]),.doutc(w_a44_0[2]),.din(a44));
	jspl3 jspl3_w_a45_0(.douta(w_a45_0[0]),.doutb(w_a45_0[1]),.doutc(w_a45_0[2]),.din(a45));
	jspl3 jspl3_w_a46_0(.douta(w_a46_0[0]),.doutb(w_a46_0[1]),.doutc(w_a46_0[2]),.din(a46));
	jspl3 jspl3_w_a47_0(.douta(w_a47_0[0]),.doutb(w_a47_0[1]),.doutc(w_a47_0[2]),.din(a47));
	jspl3 jspl3_w_a48_0(.douta(w_a48_0[0]),.doutb(w_a48_0[1]),.doutc(w_a48_0[2]),.din(a48));
	jspl3 jspl3_w_a49_0(.douta(w_a49_0[0]),.doutb(w_a49_0[1]),.doutc(w_a49_0[2]),.din(a49));
	jspl3 jspl3_w_a50_0(.douta(w_a50_0[0]),.doutb(w_a50_0[1]),.doutc(w_a50_0[2]),.din(a50));
	jspl3 jspl3_w_a51_0(.douta(w_a51_0[0]),.doutb(w_a51_0[1]),.doutc(w_a51_0[2]),.din(a51));
	jspl3 jspl3_w_a52_0(.douta(w_a52_0[0]),.doutb(w_a52_0[1]),.doutc(w_a52_0[2]),.din(a52));
	jspl3 jspl3_w_a53_0(.douta(w_a53_0[0]),.doutb(w_a53_0[1]),.doutc(w_a53_0[2]),.din(a53));
	jspl3 jspl3_w_a54_0(.douta(w_a54_0[0]),.doutb(w_a54_0[1]),.doutc(w_a54_0[2]),.din(a54));
	jspl3 jspl3_w_a55_0(.douta(w_a55_0[0]),.doutb(w_a55_0[1]),.doutc(w_a55_0[2]),.din(a55));
	jspl3 jspl3_w_a56_0(.douta(w_a56_0[0]),.doutb(w_a56_0[1]),.doutc(w_a56_0[2]),.din(a56));
	jspl3 jspl3_w_a57_0(.douta(w_a57_0[0]),.doutb(w_a57_0[1]),.doutc(w_a57_0[2]),.din(a57));
	jspl3 jspl3_w_a58_0(.douta(w_a58_0[0]),.doutb(w_a58_0[1]),.doutc(w_a58_0[2]),.din(a58));
	jspl3 jspl3_w_a59_0(.douta(w_a59_0[0]),.doutb(w_a59_0[1]),.doutc(w_a59_0[2]),.din(a59));
	jspl3 jspl3_w_a60_0(.douta(w_a60_0[0]),.doutb(w_a60_0[1]),.doutc(w_a60_0[2]),.din(a60));
	jspl3 jspl3_w_a61_0(.douta(w_a61_0[0]),.doutb(w_a61_0[1]),.doutc(w_a61_0[2]),.din(a61));
	jspl3 jspl3_w_a62_0(.douta(w_a62_0[0]),.doutb(w_a62_0[1]),.doutc(w_a62_0[2]),.din(a62));
	jspl3 jspl3_w_a63_0(.douta(w_a63_0[0]),.doutb(w_a63_0[1]),.doutc(w_a63_0[2]),.din(a63));
	jspl3 jspl3_w_a64_0(.douta(w_a64_0[0]),.doutb(w_a64_0[1]),.doutc(w_a64_0[2]),.din(a64));
	jspl3 jspl3_w_a65_0(.douta(w_a65_0[0]),.doutb(w_a65_0[1]),.doutc(w_a65_0[2]),.din(a65));
	jspl3 jspl3_w_a66_0(.douta(w_a66_0[0]),.doutb(w_a66_0[1]),.doutc(w_a66_0[2]),.din(a66));
	jspl3 jspl3_w_a67_0(.douta(w_a67_0[0]),.doutb(w_a67_0[1]),.doutc(w_a67_0[2]),.din(a67));
	jspl3 jspl3_w_a68_0(.douta(w_a68_0[0]),.doutb(w_a68_0[1]),.doutc(w_a68_0[2]),.din(a68));
	jspl3 jspl3_w_a69_0(.douta(w_a69_0[0]),.doutb(w_a69_0[1]),.doutc(w_a69_0[2]),.din(a69));
	jspl3 jspl3_w_a70_0(.douta(w_a70_0[0]),.doutb(w_a70_0[1]),.doutc(w_a70_0[2]),.din(a70));
	jspl3 jspl3_w_a71_0(.douta(w_a71_0[0]),.doutb(w_a71_0[1]),.doutc(w_a71_0[2]),.din(a71));
	jspl3 jspl3_w_a72_0(.douta(w_a72_0[0]),.doutb(w_a72_0[1]),.doutc(w_a72_0[2]),.din(a72));
	jspl3 jspl3_w_a73_0(.douta(w_a73_0[0]),.doutb(w_a73_0[1]),.doutc(w_a73_0[2]),.din(a73));
	jspl3 jspl3_w_a74_0(.douta(w_a74_0[0]),.doutb(w_a74_0[1]),.doutc(w_a74_0[2]),.din(a74));
	jspl3 jspl3_w_a75_0(.douta(w_a75_0[0]),.doutb(w_a75_0[1]),.doutc(w_a75_0[2]),.din(a75));
	jspl3 jspl3_w_a76_0(.douta(w_a76_0[0]),.doutb(w_a76_0[1]),.doutc(w_a76_0[2]),.din(a76));
	jspl3 jspl3_w_a77_0(.douta(w_a77_0[0]),.doutb(w_a77_0[1]),.doutc(w_a77_0[2]),.din(a77));
	jspl3 jspl3_w_a78_0(.douta(w_a78_0[0]),.doutb(w_a78_0[1]),.doutc(w_a78_0[2]),.din(a78));
	jspl3 jspl3_w_a79_0(.douta(w_a79_0[0]),.doutb(w_a79_0[1]),.doutc(w_a79_0[2]),.din(a79));
	jspl3 jspl3_w_a80_0(.douta(w_a80_0[0]),.doutb(w_a80_0[1]),.doutc(w_a80_0[2]),.din(a80));
	jspl3 jspl3_w_a81_0(.douta(w_a81_0[0]),.doutb(w_a81_0[1]),.doutc(w_a81_0[2]),.din(a81));
	jspl3 jspl3_w_a82_0(.douta(w_a82_0[0]),.doutb(w_a82_0[1]),.doutc(w_a82_0[2]),.din(a82));
	jspl3 jspl3_w_a83_0(.douta(w_a83_0[0]),.doutb(w_a83_0[1]),.doutc(w_a83_0[2]),.din(a83));
	jspl3 jspl3_w_a84_0(.douta(w_a84_0[0]),.doutb(w_a84_0[1]),.doutc(w_a84_0[2]),.din(a84));
	jspl3 jspl3_w_a85_0(.douta(w_a85_0[0]),.doutb(w_a85_0[1]),.doutc(w_a85_0[2]),.din(a85));
	jspl3 jspl3_w_a86_0(.douta(w_a86_0[0]),.doutb(w_a86_0[1]),.doutc(w_a86_0[2]),.din(a86));
	jspl3 jspl3_w_a87_0(.douta(w_a87_0[0]),.doutb(w_a87_0[1]),.doutc(w_a87_0[2]),.din(a87));
	jspl3 jspl3_w_a88_0(.douta(w_a88_0[0]),.doutb(w_a88_0[1]),.doutc(w_a88_0[2]),.din(a88));
	jspl3 jspl3_w_a89_0(.douta(w_a89_0[0]),.doutb(w_a89_0[1]),.doutc(w_a89_0[2]),.din(a89));
	jspl3 jspl3_w_a90_0(.douta(w_a90_0[0]),.doutb(w_a90_0[1]),.doutc(w_a90_0[2]),.din(a90));
	jspl3 jspl3_w_a91_0(.douta(w_a91_0[0]),.doutb(w_a91_0[1]),.doutc(w_a91_0[2]),.din(a91));
	jspl3 jspl3_w_a92_0(.douta(w_a92_0[0]),.doutb(w_a92_0[1]),.doutc(w_a92_0[2]),.din(a92));
	jspl3 jspl3_w_a93_0(.douta(w_a93_0[0]),.doutb(w_a93_0[1]),.doutc(w_a93_0[2]),.din(a93));
	jspl3 jspl3_w_a94_0(.douta(w_a94_0[0]),.doutb(w_a94_0[1]),.doutc(w_a94_0[2]),.din(a94));
	jspl3 jspl3_w_a95_0(.douta(w_a95_0[0]),.doutb(w_a95_0[1]),.doutc(w_a95_0[2]),.din(a95));
	jspl3 jspl3_w_a96_0(.douta(w_a96_0[0]),.doutb(w_a96_0[1]),.doutc(w_a96_0[2]),.din(a96));
	jspl3 jspl3_w_a97_0(.douta(w_a97_0[0]),.doutb(w_a97_0[1]),.doutc(w_a97_0[2]),.din(a97));
	jspl3 jspl3_w_a98_0(.douta(w_a98_0[0]),.doutb(w_a98_0[1]),.doutc(w_a98_0[2]),.din(a98));
	jspl3 jspl3_w_a99_0(.douta(w_a99_0[0]),.doutb(w_a99_0[1]),.doutc(w_a99_0[2]),.din(a99));
	jspl3 jspl3_w_a100_0(.douta(w_a100_0[0]),.doutb(w_a100_0[1]),.doutc(w_a100_0[2]),.din(a100));
	jspl3 jspl3_w_a101_0(.douta(w_a101_0[0]),.doutb(w_a101_0[1]),.doutc(w_a101_0[2]),.din(a101));
	jspl3 jspl3_w_a102_0(.douta(w_a102_0[0]),.doutb(w_a102_0[1]),.doutc(w_a102_0[2]),.din(a102));
	jspl3 jspl3_w_a103_0(.douta(w_a103_0[0]),.doutb(w_a103_0[1]),.doutc(w_a103_0[2]),.din(a103));
	jspl3 jspl3_w_a104_0(.douta(w_a104_0[0]),.doutb(w_a104_0[1]),.doutc(w_a104_0[2]),.din(a104));
	jspl3 jspl3_w_a105_0(.douta(w_a105_0[0]),.doutb(w_a105_0[1]),.doutc(w_a105_0[2]),.din(a105));
	jspl3 jspl3_w_a106_0(.douta(w_a106_0[0]),.doutb(w_a106_0[1]),.doutc(w_a106_0[2]),.din(a106));
	jspl3 jspl3_w_a107_0(.douta(w_a107_0[0]),.doutb(w_a107_0[1]),.doutc(w_a107_0[2]),.din(a107));
	jspl3 jspl3_w_a108_0(.douta(w_a108_0[0]),.doutb(w_a108_0[1]),.doutc(w_a108_0[2]),.din(a108));
	jspl3 jspl3_w_a109_0(.douta(w_a109_0[0]),.doutb(w_a109_0[1]),.doutc(w_a109_0[2]),.din(a109));
	jspl3 jspl3_w_a110_0(.douta(w_a110_0[0]),.doutb(w_a110_0[1]),.doutc(w_a110_0[2]),.din(a110));
	jspl3 jspl3_w_a111_0(.douta(w_a111_0[0]),.doutb(w_a111_0[1]),.doutc(w_a111_0[2]),.din(a111));
	jspl3 jspl3_w_a112_0(.douta(w_a112_0[0]),.doutb(w_a112_0[1]),.doutc(w_a112_0[2]),.din(a112));
	jspl3 jspl3_w_a113_0(.douta(w_a113_0[0]),.doutb(w_a113_0[1]),.doutc(w_a113_0[2]),.din(a113));
	jspl3 jspl3_w_a114_0(.douta(w_a114_0[0]),.doutb(w_a114_0[1]),.doutc(w_a114_0[2]),.din(a114));
	jspl3 jspl3_w_a115_0(.douta(w_a115_0[0]),.doutb(w_a115_0[1]),.doutc(w_a115_0[2]),.din(a115));
	jspl3 jspl3_w_a116_0(.douta(w_a116_0[0]),.doutb(w_a116_0[1]),.doutc(w_a116_0[2]),.din(a116));
	jspl3 jspl3_w_a117_0(.douta(w_a117_0[0]),.doutb(w_a117_0[1]),.doutc(w_a117_0[2]),.din(a117));
	jspl3 jspl3_w_a118_0(.douta(w_a118_0[0]),.doutb(w_a118_0[1]),.doutc(w_a118_0[2]),.din(a118));
	jspl3 jspl3_w_a119_0(.douta(w_a119_0[0]),.doutb(w_a119_0[1]),.doutc(w_a119_0[2]),.din(a119));
	jspl3 jspl3_w_a120_0(.douta(w_a120_0[0]),.doutb(w_a120_0[1]),.doutc(w_a120_0[2]),.din(a120));
	jspl3 jspl3_w_a121_0(.douta(w_a121_0[0]),.doutb(w_a121_0[1]),.doutc(w_a121_0[2]),.din(a121));
	jspl3 jspl3_w_a122_0(.douta(w_a122_0[0]),.doutb(w_a122_0[1]),.doutc(w_a122_0[2]),.din(a122));
	jspl3 jspl3_w_a123_0(.douta(w_a123_0[0]),.doutb(w_a123_0[1]),.doutc(w_a123_0[2]),.din(a123));
	jspl3 jspl3_w_a124_0(.douta(w_a124_0[0]),.doutb(w_a124_0[1]),.doutc(w_a124_0[2]),.din(a124));
	jspl3 jspl3_w_a125_0(.douta(w_a125_0[0]),.doutb(w_a125_0[1]),.doutc(w_a125_0[2]),.din(a125));
	jspl3 jspl3_w_a126_0(.douta(w_a126_0[0]),.doutb(w_a126_0[1]),.doutc(w_a126_0[2]),.din(a126));
	jspl3 jspl3_w_a127_0(.douta(w_a127_0[0]),.doutb(w_a127_0[1]),.doutc(w_a127_0[2]),.din(a127));
	jspl jspl_w_b0_0(.douta(w_b0_0[0]),.doutb(w_b0_0[1]),.din(b0));
	jspl3 jspl3_w_b1_0(.douta(w_b1_0[0]),.doutb(w_b1_0[1]),.doutc(w_b1_0[2]),.din(b1));
	jspl3 jspl3_w_b2_0(.douta(w_b2_0[0]),.doutb(w_b2_0[1]),.doutc(w_b2_0[2]),.din(b2));
	jspl3 jspl3_w_b3_0(.douta(w_b3_0[0]),.doutb(w_b3_0[1]),.doutc(w_b3_0[2]),.din(b3));
	jspl3 jspl3_w_b4_0(.douta(w_b4_0[0]),.doutb(w_b4_0[1]),.doutc(w_b4_0[2]),.din(b4));
	jspl3 jspl3_w_b5_0(.douta(w_b5_0[0]),.doutb(w_b5_0[1]),.doutc(w_b5_0[2]),.din(b5));
	jspl3 jspl3_w_b6_0(.douta(w_b6_0[0]),.doutb(w_b6_0[1]),.doutc(w_b6_0[2]),.din(b6));
	jspl3 jspl3_w_b7_0(.douta(w_b7_0[0]),.doutb(w_b7_0[1]),.doutc(w_b7_0[2]),.din(b7));
	jspl3 jspl3_w_b8_0(.douta(w_b8_0[0]),.doutb(w_b8_0[1]),.doutc(w_b8_0[2]),.din(b8));
	jspl3 jspl3_w_b9_0(.douta(w_b9_0[0]),.doutb(w_b9_0[1]),.doutc(w_b9_0[2]),.din(b9));
	jspl3 jspl3_w_b10_0(.douta(w_b10_0[0]),.doutb(w_b10_0[1]),.doutc(w_b10_0[2]),.din(b10));
	jspl3 jspl3_w_b11_0(.douta(w_b11_0[0]),.doutb(w_b11_0[1]),.doutc(w_b11_0[2]),.din(b11));
	jspl3 jspl3_w_b12_0(.douta(w_b12_0[0]),.doutb(w_b12_0[1]),.doutc(w_b12_0[2]),.din(b12));
	jspl3 jspl3_w_b13_0(.douta(w_b13_0[0]),.doutb(w_b13_0[1]),.doutc(w_b13_0[2]),.din(b13));
	jspl3 jspl3_w_b14_0(.douta(w_b14_0[0]),.doutb(w_b14_0[1]),.doutc(w_b14_0[2]),.din(b14));
	jspl3 jspl3_w_b15_0(.douta(w_b15_0[0]),.doutb(w_b15_0[1]),.doutc(w_b15_0[2]),.din(b15));
	jspl3 jspl3_w_b16_0(.douta(w_b16_0[0]),.doutb(w_b16_0[1]),.doutc(w_b16_0[2]),.din(b16));
	jspl3 jspl3_w_b17_0(.douta(w_b17_0[0]),.doutb(w_b17_0[1]),.doutc(w_b17_0[2]),.din(b17));
	jspl3 jspl3_w_b18_0(.douta(w_b18_0[0]),.doutb(w_b18_0[1]),.doutc(w_b18_0[2]),.din(b18));
	jspl3 jspl3_w_b19_0(.douta(w_b19_0[0]),.doutb(w_b19_0[1]),.doutc(w_b19_0[2]),.din(b19));
	jspl3 jspl3_w_b20_0(.douta(w_b20_0[0]),.doutb(w_b20_0[1]),.doutc(w_b20_0[2]),.din(b20));
	jspl3 jspl3_w_b21_0(.douta(w_b21_0[0]),.doutb(w_b21_0[1]),.doutc(w_b21_0[2]),.din(b21));
	jspl3 jspl3_w_b22_0(.douta(w_b22_0[0]),.doutb(w_b22_0[1]),.doutc(w_b22_0[2]),.din(b22));
	jspl3 jspl3_w_b23_0(.douta(w_b23_0[0]),.doutb(w_b23_0[1]),.doutc(w_b23_0[2]),.din(b23));
	jspl3 jspl3_w_b24_0(.douta(w_b24_0[0]),.doutb(w_b24_0[1]),.doutc(w_b24_0[2]),.din(b24));
	jspl3 jspl3_w_b25_0(.douta(w_b25_0[0]),.doutb(w_b25_0[1]),.doutc(w_b25_0[2]),.din(b25));
	jspl3 jspl3_w_b26_0(.douta(w_b26_0[0]),.doutb(w_b26_0[1]),.doutc(w_b26_0[2]),.din(b26));
	jspl3 jspl3_w_b27_0(.douta(w_b27_0[0]),.doutb(w_b27_0[1]),.doutc(w_b27_0[2]),.din(b27));
	jspl3 jspl3_w_b28_0(.douta(w_b28_0[0]),.doutb(w_b28_0[1]),.doutc(w_b28_0[2]),.din(b28));
	jspl3 jspl3_w_b29_0(.douta(w_b29_0[0]),.doutb(w_b29_0[1]),.doutc(w_b29_0[2]),.din(b29));
	jspl3 jspl3_w_b30_0(.douta(w_b30_0[0]),.doutb(w_b30_0[1]),.doutc(w_b30_0[2]),.din(b30));
	jspl3 jspl3_w_b31_0(.douta(w_b31_0[0]),.doutb(w_b31_0[1]),.doutc(w_b31_0[2]),.din(b31));
	jspl3 jspl3_w_b32_0(.douta(w_b32_0[0]),.doutb(w_b32_0[1]),.doutc(w_b32_0[2]),.din(b32));
	jspl3 jspl3_w_b33_0(.douta(w_b33_0[0]),.doutb(w_b33_0[1]),.doutc(w_b33_0[2]),.din(b33));
	jspl3 jspl3_w_b34_0(.douta(w_b34_0[0]),.doutb(w_b34_0[1]),.doutc(w_b34_0[2]),.din(b34));
	jspl3 jspl3_w_b35_0(.douta(w_b35_0[0]),.doutb(w_b35_0[1]),.doutc(w_b35_0[2]),.din(b35));
	jspl3 jspl3_w_b36_0(.douta(w_b36_0[0]),.doutb(w_b36_0[1]),.doutc(w_b36_0[2]),.din(b36));
	jspl3 jspl3_w_b37_0(.douta(w_b37_0[0]),.doutb(w_b37_0[1]),.doutc(w_b37_0[2]),.din(b37));
	jspl3 jspl3_w_b38_0(.douta(w_b38_0[0]),.doutb(w_b38_0[1]),.doutc(w_b38_0[2]),.din(b38));
	jspl3 jspl3_w_b39_0(.douta(w_b39_0[0]),.doutb(w_b39_0[1]),.doutc(w_b39_0[2]),.din(b39));
	jspl3 jspl3_w_b40_0(.douta(w_b40_0[0]),.doutb(w_b40_0[1]),.doutc(w_b40_0[2]),.din(b40));
	jspl3 jspl3_w_b41_0(.douta(w_b41_0[0]),.doutb(w_b41_0[1]),.doutc(w_b41_0[2]),.din(b41));
	jspl3 jspl3_w_b42_0(.douta(w_b42_0[0]),.doutb(w_b42_0[1]),.doutc(w_b42_0[2]),.din(b42));
	jspl3 jspl3_w_b43_0(.douta(w_b43_0[0]),.doutb(w_b43_0[1]),.doutc(w_b43_0[2]),.din(b43));
	jspl3 jspl3_w_b44_0(.douta(w_b44_0[0]),.doutb(w_b44_0[1]),.doutc(w_b44_0[2]),.din(b44));
	jspl3 jspl3_w_b45_0(.douta(w_b45_0[0]),.doutb(w_b45_0[1]),.doutc(w_b45_0[2]),.din(b45));
	jspl3 jspl3_w_b46_0(.douta(w_b46_0[0]),.doutb(w_b46_0[1]),.doutc(w_b46_0[2]),.din(b46));
	jspl3 jspl3_w_b47_0(.douta(w_b47_0[0]),.doutb(w_b47_0[1]),.doutc(w_b47_0[2]),.din(b47));
	jspl3 jspl3_w_b48_0(.douta(w_b48_0[0]),.doutb(w_b48_0[1]),.doutc(w_b48_0[2]),.din(b48));
	jspl3 jspl3_w_b49_0(.douta(w_b49_0[0]),.doutb(w_b49_0[1]),.doutc(w_b49_0[2]),.din(b49));
	jspl3 jspl3_w_b50_0(.douta(w_b50_0[0]),.doutb(w_b50_0[1]),.doutc(w_b50_0[2]),.din(b50));
	jspl3 jspl3_w_b51_0(.douta(w_b51_0[0]),.doutb(w_b51_0[1]),.doutc(w_b51_0[2]),.din(b51));
	jspl3 jspl3_w_b52_0(.douta(w_b52_0[0]),.doutb(w_b52_0[1]),.doutc(w_b52_0[2]),.din(b52));
	jspl3 jspl3_w_b53_0(.douta(w_b53_0[0]),.doutb(w_b53_0[1]),.doutc(w_b53_0[2]),.din(b53));
	jspl3 jspl3_w_b54_0(.douta(w_b54_0[0]),.doutb(w_b54_0[1]),.doutc(w_b54_0[2]),.din(b54));
	jspl3 jspl3_w_b55_0(.douta(w_b55_0[0]),.doutb(w_b55_0[1]),.doutc(w_b55_0[2]),.din(b55));
	jspl3 jspl3_w_b56_0(.douta(w_b56_0[0]),.doutb(w_b56_0[1]),.doutc(w_b56_0[2]),.din(b56));
	jspl3 jspl3_w_b57_0(.douta(w_b57_0[0]),.doutb(w_b57_0[1]),.doutc(w_b57_0[2]),.din(b57));
	jspl3 jspl3_w_b58_0(.douta(w_b58_0[0]),.doutb(w_b58_0[1]),.doutc(w_b58_0[2]),.din(b58));
	jspl3 jspl3_w_b59_0(.douta(w_b59_0[0]),.doutb(w_b59_0[1]),.doutc(w_b59_0[2]),.din(b59));
	jspl3 jspl3_w_b60_0(.douta(w_b60_0[0]),.doutb(w_b60_0[1]),.doutc(w_b60_0[2]),.din(b60));
	jspl3 jspl3_w_b61_0(.douta(w_b61_0[0]),.doutb(w_b61_0[1]),.doutc(w_b61_0[2]),.din(b61));
	jspl3 jspl3_w_b62_0(.douta(w_b62_0[0]),.doutb(w_b62_0[1]),.doutc(w_b62_0[2]),.din(b62));
	jspl3 jspl3_w_b63_0(.douta(w_b63_0[0]),.doutb(w_b63_0[1]),.doutc(w_b63_0[2]),.din(b63));
	jspl3 jspl3_w_b64_0(.douta(w_b64_0[0]),.doutb(w_b64_0[1]),.doutc(w_b64_0[2]),.din(b64));
	jspl3 jspl3_w_b65_0(.douta(w_b65_0[0]),.doutb(w_b65_0[1]),.doutc(w_b65_0[2]),.din(b65));
	jspl3 jspl3_w_b66_0(.douta(w_b66_0[0]),.doutb(w_b66_0[1]),.doutc(w_b66_0[2]),.din(b66));
	jspl3 jspl3_w_b67_0(.douta(w_b67_0[0]),.doutb(w_b67_0[1]),.doutc(w_b67_0[2]),.din(b67));
	jspl3 jspl3_w_b68_0(.douta(w_b68_0[0]),.doutb(w_b68_0[1]),.doutc(w_b68_0[2]),.din(b68));
	jspl3 jspl3_w_b69_0(.douta(w_b69_0[0]),.doutb(w_b69_0[1]),.doutc(w_b69_0[2]),.din(b69));
	jspl3 jspl3_w_b70_0(.douta(w_b70_0[0]),.doutb(w_b70_0[1]),.doutc(w_b70_0[2]),.din(b70));
	jspl3 jspl3_w_b71_0(.douta(w_b71_0[0]),.doutb(w_b71_0[1]),.doutc(w_b71_0[2]),.din(b71));
	jspl3 jspl3_w_b72_0(.douta(w_b72_0[0]),.doutb(w_b72_0[1]),.doutc(w_b72_0[2]),.din(b72));
	jspl3 jspl3_w_b73_0(.douta(w_b73_0[0]),.doutb(w_b73_0[1]),.doutc(w_b73_0[2]),.din(b73));
	jspl3 jspl3_w_b74_0(.douta(w_b74_0[0]),.doutb(w_b74_0[1]),.doutc(w_b74_0[2]),.din(b74));
	jspl3 jspl3_w_b75_0(.douta(w_b75_0[0]),.doutb(w_b75_0[1]),.doutc(w_b75_0[2]),.din(b75));
	jspl3 jspl3_w_b76_0(.douta(w_b76_0[0]),.doutb(w_b76_0[1]),.doutc(w_b76_0[2]),.din(b76));
	jspl3 jspl3_w_b77_0(.douta(w_b77_0[0]),.doutb(w_b77_0[1]),.doutc(w_b77_0[2]),.din(b77));
	jspl3 jspl3_w_b78_0(.douta(w_b78_0[0]),.doutb(w_b78_0[1]),.doutc(w_b78_0[2]),.din(b78));
	jspl3 jspl3_w_b79_0(.douta(w_b79_0[0]),.doutb(w_b79_0[1]),.doutc(w_b79_0[2]),.din(b79));
	jspl3 jspl3_w_b80_0(.douta(w_b80_0[0]),.doutb(w_b80_0[1]),.doutc(w_b80_0[2]),.din(b80));
	jspl3 jspl3_w_b81_0(.douta(w_b81_0[0]),.doutb(w_b81_0[1]),.doutc(w_b81_0[2]),.din(b81));
	jspl3 jspl3_w_b82_0(.douta(w_b82_0[0]),.doutb(w_b82_0[1]),.doutc(w_b82_0[2]),.din(b82));
	jspl3 jspl3_w_b83_0(.douta(w_b83_0[0]),.doutb(w_b83_0[1]),.doutc(w_b83_0[2]),.din(b83));
	jspl3 jspl3_w_b84_0(.douta(w_b84_0[0]),.doutb(w_b84_0[1]),.doutc(w_b84_0[2]),.din(b84));
	jspl3 jspl3_w_b85_0(.douta(w_b85_0[0]),.doutb(w_b85_0[1]),.doutc(w_b85_0[2]),.din(b85));
	jspl3 jspl3_w_b86_0(.douta(w_b86_0[0]),.doutb(w_b86_0[1]),.doutc(w_b86_0[2]),.din(b86));
	jspl3 jspl3_w_b87_0(.douta(w_b87_0[0]),.doutb(w_b87_0[1]),.doutc(w_b87_0[2]),.din(b87));
	jspl3 jspl3_w_b88_0(.douta(w_b88_0[0]),.doutb(w_b88_0[1]),.doutc(w_b88_0[2]),.din(b88));
	jspl3 jspl3_w_b89_0(.douta(w_b89_0[0]),.doutb(w_b89_0[1]),.doutc(w_b89_0[2]),.din(b89));
	jspl3 jspl3_w_b90_0(.douta(w_b90_0[0]),.doutb(w_b90_0[1]),.doutc(w_b90_0[2]),.din(b90));
	jspl3 jspl3_w_b91_0(.douta(w_b91_0[0]),.doutb(w_b91_0[1]),.doutc(w_b91_0[2]),.din(b91));
	jspl3 jspl3_w_b92_0(.douta(w_b92_0[0]),.doutb(w_b92_0[1]),.doutc(w_b92_0[2]),.din(b92));
	jspl3 jspl3_w_b93_0(.douta(w_b93_0[0]),.doutb(w_b93_0[1]),.doutc(w_b93_0[2]),.din(b93));
	jspl3 jspl3_w_b94_0(.douta(w_b94_0[0]),.doutb(w_b94_0[1]),.doutc(w_b94_0[2]),.din(b94));
	jspl3 jspl3_w_b95_0(.douta(w_b95_0[0]),.doutb(w_b95_0[1]),.doutc(w_b95_0[2]),.din(b95));
	jspl3 jspl3_w_b96_0(.douta(w_b96_0[0]),.doutb(w_b96_0[1]),.doutc(w_b96_0[2]),.din(b96));
	jspl3 jspl3_w_b97_0(.douta(w_b97_0[0]),.doutb(w_b97_0[1]),.doutc(w_b97_0[2]),.din(b97));
	jspl3 jspl3_w_b98_0(.douta(w_b98_0[0]),.doutb(w_b98_0[1]),.doutc(w_b98_0[2]),.din(b98));
	jspl3 jspl3_w_b99_0(.douta(w_b99_0[0]),.doutb(w_b99_0[1]),.doutc(w_b99_0[2]),.din(b99));
	jspl3 jspl3_w_b100_0(.douta(w_b100_0[0]),.doutb(w_b100_0[1]),.doutc(w_b100_0[2]),.din(b100));
	jspl3 jspl3_w_b101_0(.douta(w_b101_0[0]),.doutb(w_b101_0[1]),.doutc(w_b101_0[2]),.din(b101));
	jspl3 jspl3_w_b102_0(.douta(w_b102_0[0]),.doutb(w_b102_0[1]),.doutc(w_b102_0[2]),.din(b102));
	jspl3 jspl3_w_b103_0(.douta(w_b103_0[0]),.doutb(w_b103_0[1]),.doutc(w_b103_0[2]),.din(b103));
	jspl3 jspl3_w_b104_0(.douta(w_b104_0[0]),.doutb(w_b104_0[1]),.doutc(w_b104_0[2]),.din(b104));
	jspl3 jspl3_w_b105_0(.douta(w_b105_0[0]),.doutb(w_b105_0[1]),.doutc(w_b105_0[2]),.din(b105));
	jspl3 jspl3_w_b106_0(.douta(w_b106_0[0]),.doutb(w_b106_0[1]),.doutc(w_b106_0[2]),.din(b106));
	jspl3 jspl3_w_b107_0(.douta(w_b107_0[0]),.doutb(w_b107_0[1]),.doutc(w_b107_0[2]),.din(b107));
	jspl3 jspl3_w_b108_0(.douta(w_b108_0[0]),.doutb(w_b108_0[1]),.doutc(w_b108_0[2]),.din(b108));
	jspl3 jspl3_w_b109_0(.douta(w_b109_0[0]),.doutb(w_b109_0[1]),.doutc(w_b109_0[2]),.din(b109));
	jspl3 jspl3_w_b110_0(.douta(w_b110_0[0]),.doutb(w_b110_0[1]),.doutc(w_b110_0[2]),.din(b110));
	jspl3 jspl3_w_b111_0(.douta(w_b111_0[0]),.doutb(w_b111_0[1]),.doutc(w_b111_0[2]),.din(b111));
	jspl3 jspl3_w_b112_0(.douta(w_b112_0[0]),.doutb(w_b112_0[1]),.doutc(w_b112_0[2]),.din(b112));
	jspl3 jspl3_w_b113_0(.douta(w_b113_0[0]),.doutb(w_b113_0[1]),.doutc(w_b113_0[2]),.din(b113));
	jspl3 jspl3_w_b114_0(.douta(w_b114_0[0]),.doutb(w_b114_0[1]),.doutc(w_b114_0[2]),.din(b114));
	jspl3 jspl3_w_b115_0(.douta(w_b115_0[0]),.doutb(w_b115_0[1]),.doutc(w_b115_0[2]),.din(b115));
	jspl3 jspl3_w_b116_0(.douta(w_b116_0[0]),.doutb(w_b116_0[1]),.doutc(w_b116_0[2]),.din(b116));
	jspl3 jspl3_w_b117_0(.douta(w_b117_0[0]),.doutb(w_b117_0[1]),.doutc(w_b117_0[2]),.din(b117));
	jspl3 jspl3_w_b118_0(.douta(w_b118_0[0]),.doutb(w_b118_0[1]),.doutc(w_b118_0[2]),.din(b118));
	jspl3 jspl3_w_b119_0(.douta(w_b119_0[0]),.doutb(w_b119_0[1]),.doutc(w_b119_0[2]),.din(b119));
	jspl3 jspl3_w_b120_0(.douta(w_b120_0[0]),.doutb(w_b120_0[1]),.doutc(w_b120_0[2]),.din(b120));
	jspl3 jspl3_w_b121_0(.douta(w_b121_0[0]),.doutb(w_b121_0[1]),.doutc(w_b121_0[2]),.din(b121));
	jspl3 jspl3_w_b122_0(.douta(w_b122_0[0]),.doutb(w_b122_0[1]),.doutc(w_b122_0[2]),.din(b122));
	jspl3 jspl3_w_b123_0(.douta(w_b123_0[0]),.doutb(w_b123_0[1]),.doutc(w_b123_0[2]),.din(b123));
	jspl3 jspl3_w_b124_0(.douta(w_b124_0[0]),.doutb(w_b124_0[1]),.doutc(w_b124_0[2]),.din(b124));
	jspl3 jspl3_w_b125_0(.douta(w_b125_0[0]),.doutb(w_b125_0[1]),.doutc(w_b125_0[2]),.din(b125));
	jspl3 jspl3_w_b126_0(.douta(w_b126_0[0]),.doutb(w_b126_0[1]),.doutc(w_b126_0[2]),.din(b126));
	jspl3 jspl3_w_b127_0(.douta(w_b127_0[0]),.doutb(w_b127_0[1]),.doutc(w_b127_0[2]),.din(b127));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(n387));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n399_0(.douta(w_n399_0[0]),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(n417));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(n453));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl jspl_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.din(n495));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(n501));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl jspl_w_n525_0(.douta(w_n525_0[0]),.doutb(w_n525_0[1]),.din(n525));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n549_0(.douta(w_n549_0[0]),.doutb(w_n549_0[1]),.din(n549));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.din(n561));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(n567));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(n573));
	jspl jspl_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.din(n579));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.din(n633));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl jspl_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.din(n753));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(n783));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl jspl_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(n807));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl jspl_w_n831_0(.douta(w_n831_0[0]),.doutb(w_n831_0[1]),.din(n831));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(n837));
	jspl jspl_w_n843_0(.douta(w_n843_0[0]),.doutb(w_n843_0[1]),.din(n843));
	jspl jspl_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.din(n849));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(n861));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n873_0(.douta(w_n873_0[0]),.doutb(w_n873_0[1]),.din(n873));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(n915));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n933_0(.douta(w_n933_0[0]),.doutb(w_n933_0[1]),.din(n933));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(n939));
	jspl jspl_w_n945_0(.douta(w_n945_0[0]),.doutb(w_n945_0[1]),.din(n945));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(n951));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n963_0(.douta(w_n963_0[0]),.doutb(w_n963_0[1]),.din(n963));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n975_0(.douta(w_n975_0[0]),.doutb(w_n975_0[1]),.din(n975));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1047_0(.douta(w_n1047_0[0]),.doutb(w_n1047_0[1]),.din(n1047));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(n1053));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1065_0(.douta(w_n1065_0[0]),.doutb(w_n1065_0[1]),.din(n1065));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(n1077));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(n1083));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(n1089));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(n1095));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(n1101));
	jspl jspl_w_n1107_0(.douta(w_n1107_0[0]),.doutb(w_n1107_0[1]),.din(n1107));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.din(n1113));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(n1125));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1143_0(.douta(w_n1143_0[0]),.doutb(w_n1143_0[1]),.din(n1143));
	jdff dff_B_y2pBBYfz5_0(.din(n394),.dout(w_dff_B_y2pBBYfz5_0),.clk(gclk));
	jdff dff_B_3J0ThVUc7_0(.din(n400),.dout(w_dff_B_3J0ThVUc7_0),.clk(gclk));
	jdff dff_B_S1pCGBH96_0(.din(w_dff_B_3J0ThVUc7_0),.dout(w_dff_B_S1pCGBH96_0),.clk(gclk));
	jdff dff_B_mnbAlDI71_0(.din(n406),.dout(w_dff_B_mnbAlDI71_0),.clk(gclk));
	jdff dff_B_NzAYujON5_0(.din(w_dff_B_mnbAlDI71_0),.dout(w_dff_B_NzAYujON5_0),.clk(gclk));
	jdff dff_B_WlKsqUMj9_0(.din(w_dff_B_NzAYujON5_0),.dout(w_dff_B_WlKsqUMj9_0),.clk(gclk));
	jdff dff_B_Brc2L2JI6_0(.din(n412),.dout(w_dff_B_Brc2L2JI6_0),.clk(gclk));
	jdff dff_B_uhMTUALy6_0(.din(w_dff_B_Brc2L2JI6_0),.dout(w_dff_B_uhMTUALy6_0),.clk(gclk));
	jdff dff_B_l3Z1Mo835_0(.din(w_dff_B_uhMTUALy6_0),.dout(w_dff_B_l3Z1Mo835_0),.clk(gclk));
	jdff dff_B_Q6vqZJ6y8_0(.din(w_dff_B_l3Z1Mo835_0),.dout(w_dff_B_Q6vqZJ6y8_0),.clk(gclk));
	jdff dff_B_Vw0IBdke4_0(.din(n418),.dout(w_dff_B_Vw0IBdke4_0),.clk(gclk));
	jdff dff_B_VsIXMNjy6_0(.din(w_dff_B_Vw0IBdke4_0),.dout(w_dff_B_VsIXMNjy6_0),.clk(gclk));
	jdff dff_B_bSPwuxqp4_0(.din(w_dff_B_VsIXMNjy6_0),.dout(w_dff_B_bSPwuxqp4_0),.clk(gclk));
	jdff dff_B_s84U52Se8_0(.din(w_dff_B_bSPwuxqp4_0),.dout(w_dff_B_s84U52Se8_0),.clk(gclk));
	jdff dff_B_8jJ4BMCH1_0(.din(w_dff_B_s84U52Se8_0),.dout(w_dff_B_8jJ4BMCH1_0),.clk(gclk));
	jdff dff_B_AEPIaLck4_0(.din(n424),.dout(w_dff_B_AEPIaLck4_0),.clk(gclk));
	jdff dff_B_BPO87s3p9_0(.din(w_dff_B_AEPIaLck4_0),.dout(w_dff_B_BPO87s3p9_0),.clk(gclk));
	jdff dff_B_4zLuvkWy1_0(.din(w_dff_B_BPO87s3p9_0),.dout(w_dff_B_4zLuvkWy1_0),.clk(gclk));
	jdff dff_B_Lyc0HPPJ1_0(.din(w_dff_B_4zLuvkWy1_0),.dout(w_dff_B_Lyc0HPPJ1_0),.clk(gclk));
	jdff dff_B_1hvRqtBe9_0(.din(w_dff_B_Lyc0HPPJ1_0),.dout(w_dff_B_1hvRqtBe9_0),.clk(gclk));
	jdff dff_B_7r08WE430_0(.din(w_dff_B_1hvRqtBe9_0),.dout(w_dff_B_7r08WE430_0),.clk(gclk));
	jdff dff_B_xHIFgZia5_0(.din(n430),.dout(w_dff_B_xHIFgZia5_0),.clk(gclk));
	jdff dff_B_ENitSJQy5_0(.din(w_dff_B_xHIFgZia5_0),.dout(w_dff_B_ENitSJQy5_0),.clk(gclk));
	jdff dff_B_HCc7mr6w4_0(.din(w_dff_B_ENitSJQy5_0),.dout(w_dff_B_HCc7mr6w4_0),.clk(gclk));
	jdff dff_B_bd1c5jY57_0(.din(w_dff_B_HCc7mr6w4_0),.dout(w_dff_B_bd1c5jY57_0),.clk(gclk));
	jdff dff_B_6C0ksYw72_0(.din(w_dff_B_bd1c5jY57_0),.dout(w_dff_B_6C0ksYw72_0),.clk(gclk));
	jdff dff_B_pgqcWTDx4_0(.din(w_dff_B_6C0ksYw72_0),.dout(w_dff_B_pgqcWTDx4_0),.clk(gclk));
	jdff dff_B_i2DkyCua4_0(.din(w_dff_B_pgqcWTDx4_0),.dout(w_dff_B_i2DkyCua4_0),.clk(gclk));
	jdff dff_B_mNcyzUcq1_0(.din(n436),.dout(w_dff_B_mNcyzUcq1_0),.clk(gclk));
	jdff dff_B_DbF5kOQi0_0(.din(w_dff_B_mNcyzUcq1_0),.dout(w_dff_B_DbF5kOQi0_0),.clk(gclk));
	jdff dff_B_DYOiTE2s7_0(.din(w_dff_B_DbF5kOQi0_0),.dout(w_dff_B_DYOiTE2s7_0),.clk(gclk));
	jdff dff_B_l0i7qBUN1_0(.din(w_dff_B_DYOiTE2s7_0),.dout(w_dff_B_l0i7qBUN1_0),.clk(gclk));
	jdff dff_B_FSyTsyEj6_0(.din(w_dff_B_l0i7qBUN1_0),.dout(w_dff_B_FSyTsyEj6_0),.clk(gclk));
	jdff dff_B_BR29qnUu8_0(.din(w_dff_B_FSyTsyEj6_0),.dout(w_dff_B_BR29qnUu8_0),.clk(gclk));
	jdff dff_B_Qd56E6vg8_0(.din(w_dff_B_BR29qnUu8_0),.dout(w_dff_B_Qd56E6vg8_0),.clk(gclk));
	jdff dff_B_xJonAAGK0_0(.din(w_dff_B_Qd56E6vg8_0),.dout(w_dff_B_xJonAAGK0_0),.clk(gclk));
	jdff dff_B_BkDsgWbV3_0(.din(n442),.dout(w_dff_B_BkDsgWbV3_0),.clk(gclk));
	jdff dff_B_AnrW8w1J2_0(.din(w_dff_B_BkDsgWbV3_0),.dout(w_dff_B_AnrW8w1J2_0),.clk(gclk));
	jdff dff_B_b8mra9OC2_0(.din(w_dff_B_AnrW8w1J2_0),.dout(w_dff_B_b8mra9OC2_0),.clk(gclk));
	jdff dff_B_AkNPTd1e7_0(.din(w_dff_B_b8mra9OC2_0),.dout(w_dff_B_AkNPTd1e7_0),.clk(gclk));
	jdff dff_B_qhdODlqZ7_0(.din(w_dff_B_AkNPTd1e7_0),.dout(w_dff_B_qhdODlqZ7_0),.clk(gclk));
	jdff dff_B_Y5ecTrgg6_0(.din(w_dff_B_qhdODlqZ7_0),.dout(w_dff_B_Y5ecTrgg6_0),.clk(gclk));
	jdff dff_B_VsdGWGmT1_0(.din(w_dff_B_Y5ecTrgg6_0),.dout(w_dff_B_VsdGWGmT1_0),.clk(gclk));
	jdff dff_B_cXMlOdRu1_0(.din(w_dff_B_VsdGWGmT1_0),.dout(w_dff_B_cXMlOdRu1_0),.clk(gclk));
	jdff dff_B_KD70119c7_0(.din(w_dff_B_cXMlOdRu1_0),.dout(w_dff_B_KD70119c7_0),.clk(gclk));
	jdff dff_B_SYcaX9bI7_0(.din(n448),.dout(w_dff_B_SYcaX9bI7_0),.clk(gclk));
	jdff dff_B_VgxfLs2T1_0(.din(w_dff_B_SYcaX9bI7_0),.dout(w_dff_B_VgxfLs2T1_0),.clk(gclk));
	jdff dff_B_X0F1zZE67_0(.din(w_dff_B_VgxfLs2T1_0),.dout(w_dff_B_X0F1zZE67_0),.clk(gclk));
	jdff dff_B_cuC6wUPc7_0(.din(w_dff_B_X0F1zZE67_0),.dout(w_dff_B_cuC6wUPc7_0),.clk(gclk));
	jdff dff_B_8191GAeV7_0(.din(w_dff_B_cuC6wUPc7_0),.dout(w_dff_B_8191GAeV7_0),.clk(gclk));
	jdff dff_B_YYa4o79w2_0(.din(w_dff_B_8191GAeV7_0),.dout(w_dff_B_YYa4o79w2_0),.clk(gclk));
	jdff dff_B_GW7ply0u6_0(.din(w_dff_B_YYa4o79w2_0),.dout(w_dff_B_GW7ply0u6_0),.clk(gclk));
	jdff dff_B_8tl8GIG71_0(.din(w_dff_B_GW7ply0u6_0),.dout(w_dff_B_8tl8GIG71_0),.clk(gclk));
	jdff dff_B_u12WWdo53_0(.din(w_dff_B_8tl8GIG71_0),.dout(w_dff_B_u12WWdo53_0),.clk(gclk));
	jdff dff_B_i8x4P8bS8_0(.din(w_dff_B_u12WWdo53_0),.dout(w_dff_B_i8x4P8bS8_0),.clk(gclk));
	jdff dff_B_TzFE9tjS7_0(.din(n454),.dout(w_dff_B_TzFE9tjS7_0),.clk(gclk));
	jdff dff_B_cU72aOqo1_0(.din(w_dff_B_TzFE9tjS7_0),.dout(w_dff_B_cU72aOqo1_0),.clk(gclk));
	jdff dff_B_KZbuGsuV1_0(.din(w_dff_B_cU72aOqo1_0),.dout(w_dff_B_KZbuGsuV1_0),.clk(gclk));
	jdff dff_B_LiAiLy0l0_0(.din(w_dff_B_KZbuGsuV1_0),.dout(w_dff_B_LiAiLy0l0_0),.clk(gclk));
	jdff dff_B_s5RweoEM8_0(.din(w_dff_B_LiAiLy0l0_0),.dout(w_dff_B_s5RweoEM8_0),.clk(gclk));
	jdff dff_B_9v7STkiO0_0(.din(w_dff_B_s5RweoEM8_0),.dout(w_dff_B_9v7STkiO0_0),.clk(gclk));
	jdff dff_B_WmPJBbFW3_0(.din(w_dff_B_9v7STkiO0_0),.dout(w_dff_B_WmPJBbFW3_0),.clk(gclk));
	jdff dff_B_lAaw1exA1_0(.din(w_dff_B_WmPJBbFW3_0),.dout(w_dff_B_lAaw1exA1_0),.clk(gclk));
	jdff dff_B_DSniR09k7_0(.din(w_dff_B_lAaw1exA1_0),.dout(w_dff_B_DSniR09k7_0),.clk(gclk));
	jdff dff_B_wsiOqmRM9_0(.din(w_dff_B_DSniR09k7_0),.dout(w_dff_B_wsiOqmRM9_0),.clk(gclk));
	jdff dff_B_bSj65Sek7_0(.din(w_dff_B_wsiOqmRM9_0),.dout(w_dff_B_bSj65Sek7_0),.clk(gclk));
	jdff dff_B_utfAyrTF1_0(.din(n460),.dout(w_dff_B_utfAyrTF1_0),.clk(gclk));
	jdff dff_B_TuXlM1jX9_0(.din(w_dff_B_utfAyrTF1_0),.dout(w_dff_B_TuXlM1jX9_0),.clk(gclk));
	jdff dff_B_cLppZy5R6_0(.din(w_dff_B_TuXlM1jX9_0),.dout(w_dff_B_cLppZy5R6_0),.clk(gclk));
	jdff dff_B_UuguPchZ9_0(.din(w_dff_B_cLppZy5R6_0),.dout(w_dff_B_UuguPchZ9_0),.clk(gclk));
	jdff dff_B_Nrl2Hk9v0_0(.din(w_dff_B_UuguPchZ9_0),.dout(w_dff_B_Nrl2Hk9v0_0),.clk(gclk));
	jdff dff_B_mjt7gJjd2_0(.din(w_dff_B_Nrl2Hk9v0_0),.dout(w_dff_B_mjt7gJjd2_0),.clk(gclk));
	jdff dff_B_E3b75pyO2_0(.din(w_dff_B_mjt7gJjd2_0),.dout(w_dff_B_E3b75pyO2_0),.clk(gclk));
	jdff dff_B_qoeeGdgd2_0(.din(w_dff_B_E3b75pyO2_0),.dout(w_dff_B_qoeeGdgd2_0),.clk(gclk));
	jdff dff_B_sxe69lGc5_0(.din(w_dff_B_qoeeGdgd2_0),.dout(w_dff_B_sxe69lGc5_0),.clk(gclk));
	jdff dff_B_2raBfihI9_0(.din(w_dff_B_sxe69lGc5_0),.dout(w_dff_B_2raBfihI9_0),.clk(gclk));
	jdff dff_B_18la0t473_0(.din(w_dff_B_2raBfihI9_0),.dout(w_dff_B_18la0t473_0),.clk(gclk));
	jdff dff_B_YbutfiBd1_0(.din(w_dff_B_18la0t473_0),.dout(w_dff_B_YbutfiBd1_0),.clk(gclk));
	jdff dff_B_6urZ322P0_0(.din(n466),.dout(w_dff_B_6urZ322P0_0),.clk(gclk));
	jdff dff_B_ShgIq1m37_0(.din(w_dff_B_6urZ322P0_0),.dout(w_dff_B_ShgIq1m37_0),.clk(gclk));
	jdff dff_B_ETOlpfmb2_0(.din(w_dff_B_ShgIq1m37_0),.dout(w_dff_B_ETOlpfmb2_0),.clk(gclk));
	jdff dff_B_CEUyN6ux6_0(.din(w_dff_B_ETOlpfmb2_0),.dout(w_dff_B_CEUyN6ux6_0),.clk(gclk));
	jdff dff_B_7C2MaevD6_0(.din(w_dff_B_CEUyN6ux6_0),.dout(w_dff_B_7C2MaevD6_0),.clk(gclk));
	jdff dff_B_N6KhNZgu7_0(.din(w_dff_B_7C2MaevD6_0),.dout(w_dff_B_N6KhNZgu7_0),.clk(gclk));
	jdff dff_B_pzJrvu0e1_0(.din(w_dff_B_N6KhNZgu7_0),.dout(w_dff_B_pzJrvu0e1_0),.clk(gclk));
	jdff dff_B_A6auZr8o3_0(.din(w_dff_B_pzJrvu0e1_0),.dout(w_dff_B_A6auZr8o3_0),.clk(gclk));
	jdff dff_B_hBdeRio21_0(.din(w_dff_B_A6auZr8o3_0),.dout(w_dff_B_hBdeRio21_0),.clk(gclk));
	jdff dff_B_TKSjOwA91_0(.din(w_dff_B_hBdeRio21_0),.dout(w_dff_B_TKSjOwA91_0),.clk(gclk));
	jdff dff_B_ay9vxaw98_0(.din(w_dff_B_TKSjOwA91_0),.dout(w_dff_B_ay9vxaw98_0),.clk(gclk));
	jdff dff_B_13VDLqBe5_0(.din(w_dff_B_ay9vxaw98_0),.dout(w_dff_B_13VDLqBe5_0),.clk(gclk));
	jdff dff_B_yvhE8Xy08_0(.din(w_dff_B_13VDLqBe5_0),.dout(w_dff_B_yvhE8Xy08_0),.clk(gclk));
	jdff dff_B_PTGcPJtE0_0(.din(n472),.dout(w_dff_B_PTGcPJtE0_0),.clk(gclk));
	jdff dff_B_JpC7cviR8_0(.din(w_dff_B_PTGcPJtE0_0),.dout(w_dff_B_JpC7cviR8_0),.clk(gclk));
	jdff dff_B_H4c00HdU0_0(.din(w_dff_B_JpC7cviR8_0),.dout(w_dff_B_H4c00HdU0_0),.clk(gclk));
	jdff dff_B_upp86dzb0_0(.din(w_dff_B_H4c00HdU0_0),.dout(w_dff_B_upp86dzb0_0),.clk(gclk));
	jdff dff_B_NDnEzvqu6_0(.din(w_dff_B_upp86dzb0_0),.dout(w_dff_B_NDnEzvqu6_0),.clk(gclk));
	jdff dff_B_RpVVfcSh6_0(.din(w_dff_B_NDnEzvqu6_0),.dout(w_dff_B_RpVVfcSh6_0),.clk(gclk));
	jdff dff_B_5jursZBQ8_0(.din(w_dff_B_RpVVfcSh6_0),.dout(w_dff_B_5jursZBQ8_0),.clk(gclk));
	jdff dff_B_agPTNz1F6_0(.din(w_dff_B_5jursZBQ8_0),.dout(w_dff_B_agPTNz1F6_0),.clk(gclk));
	jdff dff_B_AvzbDx8H5_0(.din(w_dff_B_agPTNz1F6_0),.dout(w_dff_B_AvzbDx8H5_0),.clk(gclk));
	jdff dff_B_014C95Vl8_0(.din(w_dff_B_AvzbDx8H5_0),.dout(w_dff_B_014C95Vl8_0),.clk(gclk));
	jdff dff_B_kJRmBb332_0(.din(w_dff_B_014C95Vl8_0),.dout(w_dff_B_kJRmBb332_0),.clk(gclk));
	jdff dff_B_tAQ3iZIB7_0(.din(w_dff_B_kJRmBb332_0),.dout(w_dff_B_tAQ3iZIB7_0),.clk(gclk));
	jdff dff_B_cpH1PCxC9_0(.din(w_dff_B_tAQ3iZIB7_0),.dout(w_dff_B_cpH1PCxC9_0),.clk(gclk));
	jdff dff_B_0CAb5BDY8_0(.din(w_dff_B_cpH1PCxC9_0),.dout(w_dff_B_0CAb5BDY8_0),.clk(gclk));
	jdff dff_B_CVnYksQq7_0(.din(n478),.dout(w_dff_B_CVnYksQq7_0),.clk(gclk));
	jdff dff_B_LqmOP2qT4_0(.din(w_dff_B_CVnYksQq7_0),.dout(w_dff_B_LqmOP2qT4_0),.clk(gclk));
	jdff dff_B_NgxMaCRH5_0(.din(w_dff_B_LqmOP2qT4_0),.dout(w_dff_B_NgxMaCRH5_0),.clk(gclk));
	jdff dff_B_gWx6oyEi2_0(.din(w_dff_B_NgxMaCRH5_0),.dout(w_dff_B_gWx6oyEi2_0),.clk(gclk));
	jdff dff_B_Mp1NdEXh5_0(.din(w_dff_B_gWx6oyEi2_0),.dout(w_dff_B_Mp1NdEXh5_0),.clk(gclk));
	jdff dff_B_G9fjLTRe5_0(.din(w_dff_B_Mp1NdEXh5_0),.dout(w_dff_B_G9fjLTRe5_0),.clk(gclk));
	jdff dff_B_axJqJbaM2_0(.din(w_dff_B_G9fjLTRe5_0),.dout(w_dff_B_axJqJbaM2_0),.clk(gclk));
	jdff dff_B_IrnZEV9l1_0(.din(w_dff_B_axJqJbaM2_0),.dout(w_dff_B_IrnZEV9l1_0),.clk(gclk));
	jdff dff_B_0mN764PL3_0(.din(w_dff_B_IrnZEV9l1_0),.dout(w_dff_B_0mN764PL3_0),.clk(gclk));
	jdff dff_B_SqhsNIcs4_0(.din(w_dff_B_0mN764PL3_0),.dout(w_dff_B_SqhsNIcs4_0),.clk(gclk));
	jdff dff_B_4OD9xZis8_0(.din(w_dff_B_SqhsNIcs4_0),.dout(w_dff_B_4OD9xZis8_0),.clk(gclk));
	jdff dff_B_b0fr9tox6_0(.din(w_dff_B_4OD9xZis8_0),.dout(w_dff_B_b0fr9tox6_0),.clk(gclk));
	jdff dff_B_JxshsCdJ8_0(.din(w_dff_B_b0fr9tox6_0),.dout(w_dff_B_JxshsCdJ8_0),.clk(gclk));
	jdff dff_B_qiG9o07C6_0(.din(w_dff_B_JxshsCdJ8_0),.dout(w_dff_B_qiG9o07C6_0),.clk(gclk));
	jdff dff_B_M8i2g1ka6_0(.din(w_dff_B_qiG9o07C6_0),.dout(w_dff_B_M8i2g1ka6_0),.clk(gclk));
	jdff dff_B_fV77TxYs1_0(.din(n484),.dout(w_dff_B_fV77TxYs1_0),.clk(gclk));
	jdff dff_B_fksKxLpP4_0(.din(w_dff_B_fV77TxYs1_0),.dout(w_dff_B_fksKxLpP4_0),.clk(gclk));
	jdff dff_B_fCPoUfhW4_0(.din(w_dff_B_fksKxLpP4_0),.dout(w_dff_B_fCPoUfhW4_0),.clk(gclk));
	jdff dff_B_pKQ0PvID3_0(.din(w_dff_B_fCPoUfhW4_0),.dout(w_dff_B_pKQ0PvID3_0),.clk(gclk));
	jdff dff_B_jk20wsIu8_0(.din(w_dff_B_pKQ0PvID3_0),.dout(w_dff_B_jk20wsIu8_0),.clk(gclk));
	jdff dff_B_iGy5gPnm4_0(.din(w_dff_B_jk20wsIu8_0),.dout(w_dff_B_iGy5gPnm4_0),.clk(gclk));
	jdff dff_B_ZRxQ7bzK9_0(.din(w_dff_B_iGy5gPnm4_0),.dout(w_dff_B_ZRxQ7bzK9_0),.clk(gclk));
	jdff dff_B_X5bNYZFd0_0(.din(w_dff_B_ZRxQ7bzK9_0),.dout(w_dff_B_X5bNYZFd0_0),.clk(gclk));
	jdff dff_B_VFOZkSK24_0(.din(w_dff_B_X5bNYZFd0_0),.dout(w_dff_B_VFOZkSK24_0),.clk(gclk));
	jdff dff_B_QKU5NNEE8_0(.din(w_dff_B_VFOZkSK24_0),.dout(w_dff_B_QKU5NNEE8_0),.clk(gclk));
	jdff dff_B_4ZHLJ0GC2_0(.din(w_dff_B_QKU5NNEE8_0),.dout(w_dff_B_4ZHLJ0GC2_0),.clk(gclk));
	jdff dff_B_H3qk8Ngk1_0(.din(w_dff_B_4ZHLJ0GC2_0),.dout(w_dff_B_H3qk8Ngk1_0),.clk(gclk));
	jdff dff_B_sQQCfYEQ4_0(.din(w_dff_B_H3qk8Ngk1_0),.dout(w_dff_B_sQQCfYEQ4_0),.clk(gclk));
	jdff dff_B_JF1ZhYUE2_0(.din(w_dff_B_sQQCfYEQ4_0),.dout(w_dff_B_JF1ZhYUE2_0),.clk(gclk));
	jdff dff_B_F9X4gAYw8_0(.din(w_dff_B_JF1ZhYUE2_0),.dout(w_dff_B_F9X4gAYw8_0),.clk(gclk));
	jdff dff_B_CPSxdA6Y0_0(.din(w_dff_B_F9X4gAYw8_0),.dout(w_dff_B_CPSxdA6Y0_0),.clk(gclk));
	jdff dff_B_mMAUhrYt2_0(.din(n490),.dout(w_dff_B_mMAUhrYt2_0),.clk(gclk));
	jdff dff_B_2luq4joT1_0(.din(w_dff_B_mMAUhrYt2_0),.dout(w_dff_B_2luq4joT1_0),.clk(gclk));
	jdff dff_B_Pyt4EZZJ0_0(.din(w_dff_B_2luq4joT1_0),.dout(w_dff_B_Pyt4EZZJ0_0),.clk(gclk));
	jdff dff_B_Tt7ltl6B0_0(.din(w_dff_B_Pyt4EZZJ0_0),.dout(w_dff_B_Tt7ltl6B0_0),.clk(gclk));
	jdff dff_B_eOOmDQhE2_0(.din(w_dff_B_Tt7ltl6B0_0),.dout(w_dff_B_eOOmDQhE2_0),.clk(gclk));
	jdff dff_B_jEGVBdHU3_0(.din(w_dff_B_eOOmDQhE2_0),.dout(w_dff_B_jEGVBdHU3_0),.clk(gclk));
	jdff dff_B_sntaHEWZ2_0(.din(w_dff_B_jEGVBdHU3_0),.dout(w_dff_B_sntaHEWZ2_0),.clk(gclk));
	jdff dff_B_XXILh6AL2_0(.din(w_dff_B_sntaHEWZ2_0),.dout(w_dff_B_XXILh6AL2_0),.clk(gclk));
	jdff dff_B_KwalMrsG6_0(.din(w_dff_B_XXILh6AL2_0),.dout(w_dff_B_KwalMrsG6_0),.clk(gclk));
	jdff dff_B_bp4Pi2yE2_0(.din(w_dff_B_KwalMrsG6_0),.dout(w_dff_B_bp4Pi2yE2_0),.clk(gclk));
	jdff dff_B_HfK1dh8X1_0(.din(w_dff_B_bp4Pi2yE2_0),.dout(w_dff_B_HfK1dh8X1_0),.clk(gclk));
	jdff dff_B_zx6my8418_0(.din(w_dff_B_HfK1dh8X1_0),.dout(w_dff_B_zx6my8418_0),.clk(gclk));
	jdff dff_B_4KOnpXUq5_0(.din(w_dff_B_zx6my8418_0),.dout(w_dff_B_4KOnpXUq5_0),.clk(gclk));
	jdff dff_B_ZZOJ6x3S6_0(.din(w_dff_B_4KOnpXUq5_0),.dout(w_dff_B_ZZOJ6x3S6_0),.clk(gclk));
	jdff dff_B_vIxtPeBW1_0(.din(w_dff_B_ZZOJ6x3S6_0),.dout(w_dff_B_vIxtPeBW1_0),.clk(gclk));
	jdff dff_B_TRmgWZG88_0(.din(w_dff_B_vIxtPeBW1_0),.dout(w_dff_B_TRmgWZG88_0),.clk(gclk));
	jdff dff_B_c7YZMJgL7_0(.din(w_dff_B_TRmgWZG88_0),.dout(w_dff_B_c7YZMJgL7_0),.clk(gclk));
	jdff dff_B_6v93hQPr8_0(.din(n496),.dout(w_dff_B_6v93hQPr8_0),.clk(gclk));
	jdff dff_B_4hKX96Vy7_0(.din(w_dff_B_6v93hQPr8_0),.dout(w_dff_B_4hKX96Vy7_0),.clk(gclk));
	jdff dff_B_HHp5iX6Y7_0(.din(w_dff_B_4hKX96Vy7_0),.dout(w_dff_B_HHp5iX6Y7_0),.clk(gclk));
	jdff dff_B_ESPc2d4a0_0(.din(w_dff_B_HHp5iX6Y7_0),.dout(w_dff_B_ESPc2d4a0_0),.clk(gclk));
	jdff dff_B_fhX4SxUd6_0(.din(w_dff_B_ESPc2d4a0_0),.dout(w_dff_B_fhX4SxUd6_0),.clk(gclk));
	jdff dff_B_JPaywt4G5_0(.din(w_dff_B_fhX4SxUd6_0),.dout(w_dff_B_JPaywt4G5_0),.clk(gclk));
	jdff dff_B_dvfpfhKU1_0(.din(w_dff_B_JPaywt4G5_0),.dout(w_dff_B_dvfpfhKU1_0),.clk(gclk));
	jdff dff_B_jEeAVqY32_0(.din(w_dff_B_dvfpfhKU1_0),.dout(w_dff_B_jEeAVqY32_0),.clk(gclk));
	jdff dff_B_cdEo1vsy4_0(.din(w_dff_B_jEeAVqY32_0),.dout(w_dff_B_cdEo1vsy4_0),.clk(gclk));
	jdff dff_B_2wXLHRe55_0(.din(w_dff_B_cdEo1vsy4_0),.dout(w_dff_B_2wXLHRe55_0),.clk(gclk));
	jdff dff_B_4Kc4XWH48_0(.din(w_dff_B_2wXLHRe55_0),.dout(w_dff_B_4Kc4XWH48_0),.clk(gclk));
	jdff dff_B_nf5GK2AY6_0(.din(w_dff_B_4Kc4XWH48_0),.dout(w_dff_B_nf5GK2AY6_0),.clk(gclk));
	jdff dff_B_XnuqDCUM9_0(.din(w_dff_B_nf5GK2AY6_0),.dout(w_dff_B_XnuqDCUM9_0),.clk(gclk));
	jdff dff_B_xxgnqxpN8_0(.din(w_dff_B_XnuqDCUM9_0),.dout(w_dff_B_xxgnqxpN8_0),.clk(gclk));
	jdff dff_B_JbJSN1lV7_0(.din(w_dff_B_xxgnqxpN8_0),.dout(w_dff_B_JbJSN1lV7_0),.clk(gclk));
	jdff dff_B_RmSmdPOU2_0(.din(w_dff_B_JbJSN1lV7_0),.dout(w_dff_B_RmSmdPOU2_0),.clk(gclk));
	jdff dff_B_U67o42Lq5_0(.din(w_dff_B_RmSmdPOU2_0),.dout(w_dff_B_U67o42Lq5_0),.clk(gclk));
	jdff dff_B_XC5aVfCd5_0(.din(w_dff_B_U67o42Lq5_0),.dout(w_dff_B_XC5aVfCd5_0),.clk(gclk));
	jdff dff_B_G0S2GwZ09_0(.din(n502),.dout(w_dff_B_G0S2GwZ09_0),.clk(gclk));
	jdff dff_B_x62J4vje9_0(.din(w_dff_B_G0S2GwZ09_0),.dout(w_dff_B_x62J4vje9_0),.clk(gclk));
	jdff dff_B_SFRTN3Md5_0(.din(w_dff_B_x62J4vje9_0),.dout(w_dff_B_SFRTN3Md5_0),.clk(gclk));
	jdff dff_B_zkXuueZY3_0(.din(w_dff_B_SFRTN3Md5_0),.dout(w_dff_B_zkXuueZY3_0),.clk(gclk));
	jdff dff_B_ogaTn6RF0_0(.din(w_dff_B_zkXuueZY3_0),.dout(w_dff_B_ogaTn6RF0_0),.clk(gclk));
	jdff dff_B_E2Su59NV2_0(.din(w_dff_B_ogaTn6RF0_0),.dout(w_dff_B_E2Su59NV2_0),.clk(gclk));
	jdff dff_B_fRq81AU46_0(.din(w_dff_B_E2Su59NV2_0),.dout(w_dff_B_fRq81AU46_0),.clk(gclk));
	jdff dff_B_B8or83K73_0(.din(w_dff_B_fRq81AU46_0),.dout(w_dff_B_B8or83K73_0),.clk(gclk));
	jdff dff_B_BQuR4S9t9_0(.din(w_dff_B_B8or83K73_0),.dout(w_dff_B_BQuR4S9t9_0),.clk(gclk));
	jdff dff_B_dTVUfitb2_0(.din(w_dff_B_BQuR4S9t9_0),.dout(w_dff_B_dTVUfitb2_0),.clk(gclk));
	jdff dff_B_eKoNYbty9_0(.din(w_dff_B_dTVUfitb2_0),.dout(w_dff_B_eKoNYbty9_0),.clk(gclk));
	jdff dff_B_jVgOMN7k5_0(.din(w_dff_B_eKoNYbty9_0),.dout(w_dff_B_jVgOMN7k5_0),.clk(gclk));
	jdff dff_B_MVDz5b5o9_0(.din(w_dff_B_jVgOMN7k5_0),.dout(w_dff_B_MVDz5b5o9_0),.clk(gclk));
	jdff dff_B_R4DxsPjb8_0(.din(w_dff_B_MVDz5b5o9_0),.dout(w_dff_B_R4DxsPjb8_0),.clk(gclk));
	jdff dff_B_vDYeXq2q6_0(.din(w_dff_B_R4DxsPjb8_0),.dout(w_dff_B_vDYeXq2q6_0),.clk(gclk));
	jdff dff_B_R14b2tbL2_0(.din(w_dff_B_vDYeXq2q6_0),.dout(w_dff_B_R14b2tbL2_0),.clk(gclk));
	jdff dff_B_SDeuqkeB9_0(.din(w_dff_B_R14b2tbL2_0),.dout(w_dff_B_SDeuqkeB9_0),.clk(gclk));
	jdff dff_B_4GN11q8D0_0(.din(w_dff_B_SDeuqkeB9_0),.dout(w_dff_B_4GN11q8D0_0),.clk(gclk));
	jdff dff_B_3Qs1UfWC8_0(.din(w_dff_B_4GN11q8D0_0),.dout(w_dff_B_3Qs1UfWC8_0),.clk(gclk));
	jdff dff_B_MnNDT1is2_0(.din(n508),.dout(w_dff_B_MnNDT1is2_0),.clk(gclk));
	jdff dff_B_arKNd0oe8_0(.din(w_dff_B_MnNDT1is2_0),.dout(w_dff_B_arKNd0oe8_0),.clk(gclk));
	jdff dff_B_yF6uoUj18_0(.din(w_dff_B_arKNd0oe8_0),.dout(w_dff_B_yF6uoUj18_0),.clk(gclk));
	jdff dff_B_ncSfzHcb0_0(.din(w_dff_B_yF6uoUj18_0),.dout(w_dff_B_ncSfzHcb0_0),.clk(gclk));
	jdff dff_B_NxB2xmNm4_0(.din(w_dff_B_ncSfzHcb0_0),.dout(w_dff_B_NxB2xmNm4_0),.clk(gclk));
	jdff dff_B_wW0WMAum1_0(.din(w_dff_B_NxB2xmNm4_0),.dout(w_dff_B_wW0WMAum1_0),.clk(gclk));
	jdff dff_B_8bSlceo85_0(.din(w_dff_B_wW0WMAum1_0),.dout(w_dff_B_8bSlceo85_0),.clk(gclk));
	jdff dff_B_VVBAFCbw6_0(.din(w_dff_B_8bSlceo85_0),.dout(w_dff_B_VVBAFCbw6_0),.clk(gclk));
	jdff dff_B_CfV4Qxud8_0(.din(w_dff_B_VVBAFCbw6_0),.dout(w_dff_B_CfV4Qxud8_0),.clk(gclk));
	jdff dff_B_ZUkx8TLO4_0(.din(w_dff_B_CfV4Qxud8_0),.dout(w_dff_B_ZUkx8TLO4_0),.clk(gclk));
	jdff dff_B_8OWstOGa8_0(.din(w_dff_B_ZUkx8TLO4_0),.dout(w_dff_B_8OWstOGa8_0),.clk(gclk));
	jdff dff_B_mwc4vsM58_0(.din(w_dff_B_8OWstOGa8_0),.dout(w_dff_B_mwc4vsM58_0),.clk(gclk));
	jdff dff_B_LXCaRJJX6_0(.din(w_dff_B_mwc4vsM58_0),.dout(w_dff_B_LXCaRJJX6_0),.clk(gclk));
	jdff dff_B_d9dzexGR9_0(.din(w_dff_B_LXCaRJJX6_0),.dout(w_dff_B_d9dzexGR9_0),.clk(gclk));
	jdff dff_B_JSVYjlZ47_0(.din(w_dff_B_d9dzexGR9_0),.dout(w_dff_B_JSVYjlZ47_0),.clk(gclk));
	jdff dff_B_8ttyBqZq6_0(.din(w_dff_B_JSVYjlZ47_0),.dout(w_dff_B_8ttyBqZq6_0),.clk(gclk));
	jdff dff_B_Ydoe6WSr2_0(.din(w_dff_B_8ttyBqZq6_0),.dout(w_dff_B_Ydoe6WSr2_0),.clk(gclk));
	jdff dff_B_V3LACywI4_0(.din(w_dff_B_Ydoe6WSr2_0),.dout(w_dff_B_V3LACywI4_0),.clk(gclk));
	jdff dff_B_fA6vTMAx9_0(.din(w_dff_B_V3LACywI4_0),.dout(w_dff_B_fA6vTMAx9_0),.clk(gclk));
	jdff dff_B_bBoBpv7g8_0(.din(w_dff_B_fA6vTMAx9_0),.dout(w_dff_B_bBoBpv7g8_0),.clk(gclk));
	jdff dff_B_kibI2Lsn7_0(.din(n514),.dout(w_dff_B_kibI2Lsn7_0),.clk(gclk));
	jdff dff_B_1i9E8opU8_0(.din(w_dff_B_kibI2Lsn7_0),.dout(w_dff_B_1i9E8opU8_0),.clk(gclk));
	jdff dff_B_ZP0eLExa3_0(.din(w_dff_B_1i9E8opU8_0),.dout(w_dff_B_ZP0eLExa3_0),.clk(gclk));
	jdff dff_B_69jMsuV44_0(.din(w_dff_B_ZP0eLExa3_0),.dout(w_dff_B_69jMsuV44_0),.clk(gclk));
	jdff dff_B_nGUovmCT4_0(.din(w_dff_B_69jMsuV44_0),.dout(w_dff_B_nGUovmCT4_0),.clk(gclk));
	jdff dff_B_QO5EJtOg1_0(.din(w_dff_B_nGUovmCT4_0),.dout(w_dff_B_QO5EJtOg1_0),.clk(gclk));
	jdff dff_B_C6xAknTs3_0(.din(w_dff_B_QO5EJtOg1_0),.dout(w_dff_B_C6xAknTs3_0),.clk(gclk));
	jdff dff_B_UA952wVj9_0(.din(w_dff_B_C6xAknTs3_0),.dout(w_dff_B_UA952wVj9_0),.clk(gclk));
	jdff dff_B_BB5baCUN0_0(.din(w_dff_B_UA952wVj9_0),.dout(w_dff_B_BB5baCUN0_0),.clk(gclk));
	jdff dff_B_Vcl1IVhX3_0(.din(w_dff_B_BB5baCUN0_0),.dout(w_dff_B_Vcl1IVhX3_0),.clk(gclk));
	jdff dff_B_QyS5YQU86_0(.din(w_dff_B_Vcl1IVhX3_0),.dout(w_dff_B_QyS5YQU86_0),.clk(gclk));
	jdff dff_B_iZT3vNez4_0(.din(w_dff_B_QyS5YQU86_0),.dout(w_dff_B_iZT3vNez4_0),.clk(gclk));
	jdff dff_B_FmD0jpTl4_0(.din(w_dff_B_iZT3vNez4_0),.dout(w_dff_B_FmD0jpTl4_0),.clk(gclk));
	jdff dff_B_4TmnnmTU3_0(.din(w_dff_B_FmD0jpTl4_0),.dout(w_dff_B_4TmnnmTU3_0),.clk(gclk));
	jdff dff_B_uI4p7ore3_0(.din(w_dff_B_4TmnnmTU3_0),.dout(w_dff_B_uI4p7ore3_0),.clk(gclk));
	jdff dff_B_1sP5vJEI1_0(.din(w_dff_B_uI4p7ore3_0),.dout(w_dff_B_1sP5vJEI1_0),.clk(gclk));
	jdff dff_B_4hDT4OW44_0(.din(w_dff_B_1sP5vJEI1_0),.dout(w_dff_B_4hDT4OW44_0),.clk(gclk));
	jdff dff_B_DxtHLcJX3_0(.din(w_dff_B_4hDT4OW44_0),.dout(w_dff_B_DxtHLcJX3_0),.clk(gclk));
	jdff dff_B_I3FRdpeY8_0(.din(w_dff_B_DxtHLcJX3_0),.dout(w_dff_B_I3FRdpeY8_0),.clk(gclk));
	jdff dff_B_LCjZqcA51_0(.din(w_dff_B_I3FRdpeY8_0),.dout(w_dff_B_LCjZqcA51_0),.clk(gclk));
	jdff dff_B_3eiO5ewK6_0(.din(w_dff_B_LCjZqcA51_0),.dout(w_dff_B_3eiO5ewK6_0),.clk(gclk));
	jdff dff_B_bZajaUav7_0(.din(n520),.dout(w_dff_B_bZajaUav7_0),.clk(gclk));
	jdff dff_B_2ywnCjrs2_0(.din(w_dff_B_bZajaUav7_0),.dout(w_dff_B_2ywnCjrs2_0),.clk(gclk));
	jdff dff_B_cakhkuZe6_0(.din(w_dff_B_2ywnCjrs2_0),.dout(w_dff_B_cakhkuZe6_0),.clk(gclk));
	jdff dff_B_TxUsVKqT7_0(.din(w_dff_B_cakhkuZe6_0),.dout(w_dff_B_TxUsVKqT7_0),.clk(gclk));
	jdff dff_B_nQWCc0GG1_0(.din(w_dff_B_TxUsVKqT7_0),.dout(w_dff_B_nQWCc0GG1_0),.clk(gclk));
	jdff dff_B_tjUf3Qkn1_0(.din(w_dff_B_nQWCc0GG1_0),.dout(w_dff_B_tjUf3Qkn1_0),.clk(gclk));
	jdff dff_B_gl9iP9l19_0(.din(w_dff_B_tjUf3Qkn1_0),.dout(w_dff_B_gl9iP9l19_0),.clk(gclk));
	jdff dff_B_MZCl56Jb2_0(.din(w_dff_B_gl9iP9l19_0),.dout(w_dff_B_MZCl56Jb2_0),.clk(gclk));
	jdff dff_B_XQG076hP3_0(.din(w_dff_B_MZCl56Jb2_0),.dout(w_dff_B_XQG076hP3_0),.clk(gclk));
	jdff dff_B_G7z5w1fs9_0(.din(w_dff_B_XQG076hP3_0),.dout(w_dff_B_G7z5w1fs9_0),.clk(gclk));
	jdff dff_B_EiYlgQFs2_0(.din(w_dff_B_G7z5w1fs9_0),.dout(w_dff_B_EiYlgQFs2_0),.clk(gclk));
	jdff dff_B_uqHn00Cu2_0(.din(w_dff_B_EiYlgQFs2_0),.dout(w_dff_B_uqHn00Cu2_0),.clk(gclk));
	jdff dff_B_KBlSjnf81_0(.din(w_dff_B_uqHn00Cu2_0),.dout(w_dff_B_KBlSjnf81_0),.clk(gclk));
	jdff dff_B_qNnI4DkE3_0(.din(w_dff_B_KBlSjnf81_0),.dout(w_dff_B_qNnI4DkE3_0),.clk(gclk));
	jdff dff_B_QTljKgdg2_0(.din(w_dff_B_qNnI4DkE3_0),.dout(w_dff_B_QTljKgdg2_0),.clk(gclk));
	jdff dff_B_Gqcpt5RQ0_0(.din(w_dff_B_QTljKgdg2_0),.dout(w_dff_B_Gqcpt5RQ0_0),.clk(gclk));
	jdff dff_B_Mt2LI6eB8_0(.din(w_dff_B_Gqcpt5RQ0_0),.dout(w_dff_B_Mt2LI6eB8_0),.clk(gclk));
	jdff dff_B_RHnQ76dr0_0(.din(w_dff_B_Mt2LI6eB8_0),.dout(w_dff_B_RHnQ76dr0_0),.clk(gclk));
	jdff dff_B_Gv1KoaIi9_0(.din(w_dff_B_RHnQ76dr0_0),.dout(w_dff_B_Gv1KoaIi9_0),.clk(gclk));
	jdff dff_B_AxqivGkA1_0(.din(w_dff_B_Gv1KoaIi9_0),.dout(w_dff_B_AxqivGkA1_0),.clk(gclk));
	jdff dff_B_LEeGPhjq3_0(.din(w_dff_B_AxqivGkA1_0),.dout(w_dff_B_LEeGPhjq3_0),.clk(gclk));
	jdff dff_B_tF6BKpIu3_0(.din(w_dff_B_LEeGPhjq3_0),.dout(w_dff_B_tF6BKpIu3_0),.clk(gclk));
	jdff dff_B_g4pazIHh5_0(.din(n526),.dout(w_dff_B_g4pazIHh5_0),.clk(gclk));
	jdff dff_B_lpAuQVBB2_0(.din(w_dff_B_g4pazIHh5_0),.dout(w_dff_B_lpAuQVBB2_0),.clk(gclk));
	jdff dff_B_ApCAiQzs9_0(.din(w_dff_B_lpAuQVBB2_0),.dout(w_dff_B_ApCAiQzs9_0),.clk(gclk));
	jdff dff_B_SpwoBTAt1_0(.din(w_dff_B_ApCAiQzs9_0),.dout(w_dff_B_SpwoBTAt1_0),.clk(gclk));
	jdff dff_B_U96RE8xy5_0(.din(w_dff_B_SpwoBTAt1_0),.dout(w_dff_B_U96RE8xy5_0),.clk(gclk));
	jdff dff_B_eoBMukMa5_0(.din(w_dff_B_U96RE8xy5_0),.dout(w_dff_B_eoBMukMa5_0),.clk(gclk));
	jdff dff_B_4jXODQ3B9_0(.din(w_dff_B_eoBMukMa5_0),.dout(w_dff_B_4jXODQ3B9_0),.clk(gclk));
	jdff dff_B_lZcoV0uk4_0(.din(w_dff_B_4jXODQ3B9_0),.dout(w_dff_B_lZcoV0uk4_0),.clk(gclk));
	jdff dff_B_OnmiEVf42_0(.din(w_dff_B_lZcoV0uk4_0),.dout(w_dff_B_OnmiEVf42_0),.clk(gclk));
	jdff dff_B_UmPftrQi0_0(.din(w_dff_B_OnmiEVf42_0),.dout(w_dff_B_UmPftrQi0_0),.clk(gclk));
	jdff dff_B_lUONg07m6_0(.din(w_dff_B_UmPftrQi0_0),.dout(w_dff_B_lUONg07m6_0),.clk(gclk));
	jdff dff_B_3y6SCpRw2_0(.din(w_dff_B_lUONg07m6_0),.dout(w_dff_B_3y6SCpRw2_0),.clk(gclk));
	jdff dff_B_zTvh3DqS2_0(.din(w_dff_B_3y6SCpRw2_0),.dout(w_dff_B_zTvh3DqS2_0),.clk(gclk));
	jdff dff_B_5ExXoyAL2_0(.din(w_dff_B_zTvh3DqS2_0),.dout(w_dff_B_5ExXoyAL2_0),.clk(gclk));
	jdff dff_B_jT9MDiMr0_0(.din(w_dff_B_5ExXoyAL2_0),.dout(w_dff_B_jT9MDiMr0_0),.clk(gclk));
	jdff dff_B_miyIiyMV2_0(.din(w_dff_B_jT9MDiMr0_0),.dout(w_dff_B_miyIiyMV2_0),.clk(gclk));
	jdff dff_B_XvNxR3tj8_0(.din(w_dff_B_miyIiyMV2_0),.dout(w_dff_B_XvNxR3tj8_0),.clk(gclk));
	jdff dff_B_i4DJRbcS1_0(.din(w_dff_B_XvNxR3tj8_0),.dout(w_dff_B_i4DJRbcS1_0),.clk(gclk));
	jdff dff_B_eDEzBdcY7_0(.din(w_dff_B_i4DJRbcS1_0),.dout(w_dff_B_eDEzBdcY7_0),.clk(gclk));
	jdff dff_B_oJonf9lR0_0(.din(w_dff_B_eDEzBdcY7_0),.dout(w_dff_B_oJonf9lR0_0),.clk(gclk));
	jdff dff_B_9HpXUMLg0_0(.din(w_dff_B_oJonf9lR0_0),.dout(w_dff_B_9HpXUMLg0_0),.clk(gclk));
	jdff dff_B_xCoyA7NO3_0(.din(w_dff_B_9HpXUMLg0_0),.dout(w_dff_B_xCoyA7NO3_0),.clk(gclk));
	jdff dff_B_IxLjw79f1_0(.din(w_dff_B_xCoyA7NO3_0),.dout(w_dff_B_IxLjw79f1_0),.clk(gclk));
	jdff dff_B_4AYBlWCD3_0(.din(n532),.dout(w_dff_B_4AYBlWCD3_0),.clk(gclk));
	jdff dff_B_EVIdfRnr9_0(.din(w_dff_B_4AYBlWCD3_0),.dout(w_dff_B_EVIdfRnr9_0),.clk(gclk));
	jdff dff_B_M4gnDXts9_0(.din(w_dff_B_EVIdfRnr9_0),.dout(w_dff_B_M4gnDXts9_0),.clk(gclk));
	jdff dff_B_iN37gDGy2_0(.din(w_dff_B_M4gnDXts9_0),.dout(w_dff_B_iN37gDGy2_0),.clk(gclk));
	jdff dff_B_9C8KmD8m6_0(.din(w_dff_B_iN37gDGy2_0),.dout(w_dff_B_9C8KmD8m6_0),.clk(gclk));
	jdff dff_B_S5s5HRoI9_0(.din(w_dff_B_9C8KmD8m6_0),.dout(w_dff_B_S5s5HRoI9_0),.clk(gclk));
	jdff dff_B_jNAGm5og6_0(.din(w_dff_B_S5s5HRoI9_0),.dout(w_dff_B_jNAGm5og6_0),.clk(gclk));
	jdff dff_B_VG20qrEr6_0(.din(w_dff_B_jNAGm5og6_0),.dout(w_dff_B_VG20qrEr6_0),.clk(gclk));
	jdff dff_B_EwOjsB8V3_0(.din(w_dff_B_VG20qrEr6_0),.dout(w_dff_B_EwOjsB8V3_0),.clk(gclk));
	jdff dff_B_Zwux3rlQ9_0(.din(w_dff_B_EwOjsB8V3_0),.dout(w_dff_B_Zwux3rlQ9_0),.clk(gclk));
	jdff dff_B_DbvO4vQO3_0(.din(w_dff_B_Zwux3rlQ9_0),.dout(w_dff_B_DbvO4vQO3_0),.clk(gclk));
	jdff dff_B_xQjmoaY74_0(.din(w_dff_B_DbvO4vQO3_0),.dout(w_dff_B_xQjmoaY74_0),.clk(gclk));
	jdff dff_B_6a5zADIs6_0(.din(w_dff_B_xQjmoaY74_0),.dout(w_dff_B_6a5zADIs6_0),.clk(gclk));
	jdff dff_B_k2Xd6nNb8_0(.din(w_dff_B_6a5zADIs6_0),.dout(w_dff_B_k2Xd6nNb8_0),.clk(gclk));
	jdff dff_B_ms8xh3EV8_0(.din(w_dff_B_k2Xd6nNb8_0),.dout(w_dff_B_ms8xh3EV8_0),.clk(gclk));
	jdff dff_B_7kiHfSA64_0(.din(w_dff_B_ms8xh3EV8_0),.dout(w_dff_B_7kiHfSA64_0),.clk(gclk));
	jdff dff_B_chBzimeL5_0(.din(w_dff_B_7kiHfSA64_0),.dout(w_dff_B_chBzimeL5_0),.clk(gclk));
	jdff dff_B_mLe91Mmr8_0(.din(w_dff_B_chBzimeL5_0),.dout(w_dff_B_mLe91Mmr8_0),.clk(gclk));
	jdff dff_B_UeUg9eZ52_0(.din(w_dff_B_mLe91Mmr8_0),.dout(w_dff_B_UeUg9eZ52_0),.clk(gclk));
	jdff dff_B_wcqkNhM27_0(.din(w_dff_B_UeUg9eZ52_0),.dout(w_dff_B_wcqkNhM27_0),.clk(gclk));
	jdff dff_B_81f8RSgK9_0(.din(w_dff_B_wcqkNhM27_0),.dout(w_dff_B_81f8RSgK9_0),.clk(gclk));
	jdff dff_B_4pW0pTNI6_0(.din(w_dff_B_81f8RSgK9_0),.dout(w_dff_B_4pW0pTNI6_0),.clk(gclk));
	jdff dff_B_5IfrSx3F2_0(.din(w_dff_B_4pW0pTNI6_0),.dout(w_dff_B_5IfrSx3F2_0),.clk(gclk));
	jdff dff_B_poGlmfvO9_0(.din(w_dff_B_5IfrSx3F2_0),.dout(w_dff_B_poGlmfvO9_0),.clk(gclk));
	jdff dff_B_PaeZgrzM0_0(.din(n538),.dout(w_dff_B_PaeZgrzM0_0),.clk(gclk));
	jdff dff_B_OEZ0XwQM3_0(.din(w_dff_B_PaeZgrzM0_0),.dout(w_dff_B_OEZ0XwQM3_0),.clk(gclk));
	jdff dff_B_UvxWDdtn7_0(.din(w_dff_B_OEZ0XwQM3_0),.dout(w_dff_B_UvxWDdtn7_0),.clk(gclk));
	jdff dff_B_0yzfU7hL0_0(.din(w_dff_B_UvxWDdtn7_0),.dout(w_dff_B_0yzfU7hL0_0),.clk(gclk));
	jdff dff_B_bkbGC4eG6_0(.din(w_dff_B_0yzfU7hL0_0),.dout(w_dff_B_bkbGC4eG6_0),.clk(gclk));
	jdff dff_B_3RIC7VLq9_0(.din(w_dff_B_bkbGC4eG6_0),.dout(w_dff_B_3RIC7VLq9_0),.clk(gclk));
	jdff dff_B_rksoprrK5_0(.din(w_dff_B_3RIC7VLq9_0),.dout(w_dff_B_rksoprrK5_0),.clk(gclk));
	jdff dff_B_ebRdoXBX5_0(.din(w_dff_B_rksoprrK5_0),.dout(w_dff_B_ebRdoXBX5_0),.clk(gclk));
	jdff dff_B_pKVnF7wr7_0(.din(w_dff_B_ebRdoXBX5_0),.dout(w_dff_B_pKVnF7wr7_0),.clk(gclk));
	jdff dff_B_tgSJ4YhL5_0(.din(w_dff_B_pKVnF7wr7_0),.dout(w_dff_B_tgSJ4YhL5_0),.clk(gclk));
	jdff dff_B_tqmIASoO5_0(.din(w_dff_B_tgSJ4YhL5_0),.dout(w_dff_B_tqmIASoO5_0),.clk(gclk));
	jdff dff_B_1RIJh5oF4_0(.din(w_dff_B_tqmIASoO5_0),.dout(w_dff_B_1RIJh5oF4_0),.clk(gclk));
	jdff dff_B_xAhqYGbf7_0(.din(w_dff_B_1RIJh5oF4_0),.dout(w_dff_B_xAhqYGbf7_0),.clk(gclk));
	jdff dff_B_0WEnK7gQ2_0(.din(w_dff_B_xAhqYGbf7_0),.dout(w_dff_B_0WEnK7gQ2_0),.clk(gclk));
	jdff dff_B_BdA8GnSg2_0(.din(w_dff_B_0WEnK7gQ2_0),.dout(w_dff_B_BdA8GnSg2_0),.clk(gclk));
	jdff dff_B_H8v9suBR8_0(.din(w_dff_B_BdA8GnSg2_0),.dout(w_dff_B_H8v9suBR8_0),.clk(gclk));
	jdff dff_B_UriLMoYz8_0(.din(w_dff_B_H8v9suBR8_0),.dout(w_dff_B_UriLMoYz8_0),.clk(gclk));
	jdff dff_B_iL5oYczG6_0(.din(w_dff_B_UriLMoYz8_0),.dout(w_dff_B_iL5oYczG6_0),.clk(gclk));
	jdff dff_B_9HyMLtqN9_0(.din(w_dff_B_iL5oYczG6_0),.dout(w_dff_B_9HyMLtqN9_0),.clk(gclk));
	jdff dff_B_GgaWNR6y0_0(.din(w_dff_B_9HyMLtqN9_0),.dout(w_dff_B_GgaWNR6y0_0),.clk(gclk));
	jdff dff_B_WE5q7h8v2_0(.din(w_dff_B_GgaWNR6y0_0),.dout(w_dff_B_WE5q7h8v2_0),.clk(gclk));
	jdff dff_B_6VKFKMrh4_0(.din(w_dff_B_WE5q7h8v2_0),.dout(w_dff_B_6VKFKMrh4_0),.clk(gclk));
	jdff dff_B_YKUCZU4c8_0(.din(w_dff_B_6VKFKMrh4_0),.dout(w_dff_B_YKUCZU4c8_0),.clk(gclk));
	jdff dff_B_DfmVt6Xm5_0(.din(w_dff_B_YKUCZU4c8_0),.dout(w_dff_B_DfmVt6Xm5_0),.clk(gclk));
	jdff dff_B_aSGLFurX1_0(.din(w_dff_B_DfmVt6Xm5_0),.dout(w_dff_B_aSGLFurX1_0),.clk(gclk));
	jdff dff_B_RekwREfp2_0(.din(n544),.dout(w_dff_B_RekwREfp2_0),.clk(gclk));
	jdff dff_B_15CwFlLC1_0(.din(w_dff_B_RekwREfp2_0),.dout(w_dff_B_15CwFlLC1_0),.clk(gclk));
	jdff dff_B_a8rEoPRG0_0(.din(w_dff_B_15CwFlLC1_0),.dout(w_dff_B_a8rEoPRG0_0),.clk(gclk));
	jdff dff_B_vMYE1HsK1_0(.din(w_dff_B_a8rEoPRG0_0),.dout(w_dff_B_vMYE1HsK1_0),.clk(gclk));
	jdff dff_B_ovE2hrmu2_0(.din(w_dff_B_vMYE1HsK1_0),.dout(w_dff_B_ovE2hrmu2_0),.clk(gclk));
	jdff dff_B_4ZSnHJcP8_0(.din(w_dff_B_ovE2hrmu2_0),.dout(w_dff_B_4ZSnHJcP8_0),.clk(gclk));
	jdff dff_B_zgD4yy7E3_0(.din(w_dff_B_4ZSnHJcP8_0),.dout(w_dff_B_zgD4yy7E3_0),.clk(gclk));
	jdff dff_B_OYHF5RYQ2_0(.din(w_dff_B_zgD4yy7E3_0),.dout(w_dff_B_OYHF5RYQ2_0),.clk(gclk));
	jdff dff_B_LLTdxF677_0(.din(w_dff_B_OYHF5RYQ2_0),.dout(w_dff_B_LLTdxF677_0),.clk(gclk));
	jdff dff_B_eCj82QUd7_0(.din(w_dff_B_LLTdxF677_0),.dout(w_dff_B_eCj82QUd7_0),.clk(gclk));
	jdff dff_B_DFtYZ7Vw7_0(.din(w_dff_B_eCj82QUd7_0),.dout(w_dff_B_DFtYZ7Vw7_0),.clk(gclk));
	jdff dff_B_N6akSSGO5_0(.din(w_dff_B_DFtYZ7Vw7_0),.dout(w_dff_B_N6akSSGO5_0),.clk(gclk));
	jdff dff_B_bGlP83Zj6_0(.din(w_dff_B_N6akSSGO5_0),.dout(w_dff_B_bGlP83Zj6_0),.clk(gclk));
	jdff dff_B_XgB6zGjw4_0(.din(w_dff_B_bGlP83Zj6_0),.dout(w_dff_B_XgB6zGjw4_0),.clk(gclk));
	jdff dff_B_533bdWdP4_0(.din(w_dff_B_XgB6zGjw4_0),.dout(w_dff_B_533bdWdP4_0),.clk(gclk));
	jdff dff_B_GCW5oDqv4_0(.din(w_dff_B_533bdWdP4_0),.dout(w_dff_B_GCW5oDqv4_0),.clk(gclk));
	jdff dff_B_57lOSRw34_0(.din(w_dff_B_GCW5oDqv4_0),.dout(w_dff_B_57lOSRw34_0),.clk(gclk));
	jdff dff_B_CBBwr0FA9_0(.din(w_dff_B_57lOSRw34_0),.dout(w_dff_B_CBBwr0FA9_0),.clk(gclk));
	jdff dff_B_f1a1ZauG3_0(.din(w_dff_B_CBBwr0FA9_0),.dout(w_dff_B_f1a1ZauG3_0),.clk(gclk));
	jdff dff_B_ZpnRSzPu3_0(.din(w_dff_B_f1a1ZauG3_0),.dout(w_dff_B_ZpnRSzPu3_0),.clk(gclk));
	jdff dff_B_7GqLJKET8_0(.din(w_dff_B_ZpnRSzPu3_0),.dout(w_dff_B_7GqLJKET8_0),.clk(gclk));
	jdff dff_B_HcuyY8As9_0(.din(w_dff_B_7GqLJKET8_0),.dout(w_dff_B_HcuyY8As9_0),.clk(gclk));
	jdff dff_B_vBhM5tQJ7_0(.din(w_dff_B_HcuyY8As9_0),.dout(w_dff_B_vBhM5tQJ7_0),.clk(gclk));
	jdff dff_B_uJBMCCFG4_0(.din(w_dff_B_vBhM5tQJ7_0),.dout(w_dff_B_uJBMCCFG4_0),.clk(gclk));
	jdff dff_B_DbT98QkQ7_0(.din(w_dff_B_uJBMCCFG4_0),.dout(w_dff_B_DbT98QkQ7_0),.clk(gclk));
	jdff dff_B_0AYkSjrX9_0(.din(w_dff_B_DbT98QkQ7_0),.dout(w_dff_B_0AYkSjrX9_0),.clk(gclk));
	jdff dff_B_ZA1XkIpP0_0(.din(n550),.dout(w_dff_B_ZA1XkIpP0_0),.clk(gclk));
	jdff dff_B_7Cg4vMHU1_0(.din(w_dff_B_ZA1XkIpP0_0),.dout(w_dff_B_7Cg4vMHU1_0),.clk(gclk));
	jdff dff_B_br3x518c5_0(.din(w_dff_B_7Cg4vMHU1_0),.dout(w_dff_B_br3x518c5_0),.clk(gclk));
	jdff dff_B_Go7xWMxR1_0(.din(w_dff_B_br3x518c5_0),.dout(w_dff_B_Go7xWMxR1_0),.clk(gclk));
	jdff dff_B_sNH0JW9z6_0(.din(w_dff_B_Go7xWMxR1_0),.dout(w_dff_B_sNH0JW9z6_0),.clk(gclk));
	jdff dff_B_8moapIex2_0(.din(w_dff_B_sNH0JW9z6_0),.dout(w_dff_B_8moapIex2_0),.clk(gclk));
	jdff dff_B_X3q3Tuf58_0(.din(w_dff_B_8moapIex2_0),.dout(w_dff_B_X3q3Tuf58_0),.clk(gclk));
	jdff dff_B_uQpto6cv6_0(.din(w_dff_B_X3q3Tuf58_0),.dout(w_dff_B_uQpto6cv6_0),.clk(gclk));
	jdff dff_B_QH7pv2fm3_0(.din(w_dff_B_uQpto6cv6_0),.dout(w_dff_B_QH7pv2fm3_0),.clk(gclk));
	jdff dff_B_rudd1qJs9_0(.din(w_dff_B_QH7pv2fm3_0),.dout(w_dff_B_rudd1qJs9_0),.clk(gclk));
	jdff dff_B_q9N0SUOT0_0(.din(w_dff_B_rudd1qJs9_0),.dout(w_dff_B_q9N0SUOT0_0),.clk(gclk));
	jdff dff_B_c3kBIbUy9_0(.din(w_dff_B_q9N0SUOT0_0),.dout(w_dff_B_c3kBIbUy9_0),.clk(gclk));
	jdff dff_B_XWKrs8JL4_0(.din(w_dff_B_c3kBIbUy9_0),.dout(w_dff_B_XWKrs8JL4_0),.clk(gclk));
	jdff dff_B_XQAPy75b1_0(.din(w_dff_B_XWKrs8JL4_0),.dout(w_dff_B_XQAPy75b1_0),.clk(gclk));
	jdff dff_B_3xRIeh9V5_0(.din(w_dff_B_XQAPy75b1_0),.dout(w_dff_B_3xRIeh9V5_0),.clk(gclk));
	jdff dff_B_2CcKH1iZ1_0(.din(w_dff_B_3xRIeh9V5_0),.dout(w_dff_B_2CcKH1iZ1_0),.clk(gclk));
	jdff dff_B_UFIj6DOr8_0(.din(w_dff_B_2CcKH1iZ1_0),.dout(w_dff_B_UFIj6DOr8_0),.clk(gclk));
	jdff dff_B_ljBRYaAG6_0(.din(w_dff_B_UFIj6DOr8_0),.dout(w_dff_B_ljBRYaAG6_0),.clk(gclk));
	jdff dff_B_WShNyRcF1_0(.din(w_dff_B_ljBRYaAG6_0),.dout(w_dff_B_WShNyRcF1_0),.clk(gclk));
	jdff dff_B_Ift2MArW2_0(.din(w_dff_B_WShNyRcF1_0),.dout(w_dff_B_Ift2MArW2_0),.clk(gclk));
	jdff dff_B_BnUgafsP1_0(.din(w_dff_B_Ift2MArW2_0),.dout(w_dff_B_BnUgafsP1_0),.clk(gclk));
	jdff dff_B_XqJZkZQq0_0(.din(w_dff_B_BnUgafsP1_0),.dout(w_dff_B_XqJZkZQq0_0),.clk(gclk));
	jdff dff_B_8gmQCQmS9_0(.din(w_dff_B_XqJZkZQq0_0),.dout(w_dff_B_8gmQCQmS9_0),.clk(gclk));
	jdff dff_B_5C3W7TxS4_0(.din(w_dff_B_8gmQCQmS9_0),.dout(w_dff_B_5C3W7TxS4_0),.clk(gclk));
	jdff dff_B_74Scc9qY7_0(.din(w_dff_B_5C3W7TxS4_0),.dout(w_dff_B_74Scc9qY7_0),.clk(gclk));
	jdff dff_B_mgwSIloA7_0(.din(w_dff_B_74Scc9qY7_0),.dout(w_dff_B_mgwSIloA7_0),.clk(gclk));
	jdff dff_B_bWpvlkFu0_0(.din(w_dff_B_mgwSIloA7_0),.dout(w_dff_B_bWpvlkFu0_0),.clk(gclk));
	jdff dff_B_xk0VIGMy4_0(.din(n556),.dout(w_dff_B_xk0VIGMy4_0),.clk(gclk));
	jdff dff_B_OkRSIUZc4_0(.din(w_dff_B_xk0VIGMy4_0),.dout(w_dff_B_OkRSIUZc4_0),.clk(gclk));
	jdff dff_B_ZduKGcBM3_0(.din(w_dff_B_OkRSIUZc4_0),.dout(w_dff_B_ZduKGcBM3_0),.clk(gclk));
	jdff dff_B_A5WWflar5_0(.din(w_dff_B_ZduKGcBM3_0),.dout(w_dff_B_A5WWflar5_0),.clk(gclk));
	jdff dff_B_e1u8KWbN2_0(.din(w_dff_B_A5WWflar5_0),.dout(w_dff_B_e1u8KWbN2_0),.clk(gclk));
	jdff dff_B_Akd77nII6_0(.din(w_dff_B_e1u8KWbN2_0),.dout(w_dff_B_Akd77nII6_0),.clk(gclk));
	jdff dff_B_sci2xV2l0_0(.din(w_dff_B_Akd77nII6_0),.dout(w_dff_B_sci2xV2l0_0),.clk(gclk));
	jdff dff_B_ArbpdaB97_0(.din(w_dff_B_sci2xV2l0_0),.dout(w_dff_B_ArbpdaB97_0),.clk(gclk));
	jdff dff_B_uZH9Vvxy2_0(.din(w_dff_B_ArbpdaB97_0),.dout(w_dff_B_uZH9Vvxy2_0),.clk(gclk));
	jdff dff_B_5thX7RJO0_0(.din(w_dff_B_uZH9Vvxy2_0),.dout(w_dff_B_5thX7RJO0_0),.clk(gclk));
	jdff dff_B_Ip28Qx8p6_0(.din(w_dff_B_5thX7RJO0_0),.dout(w_dff_B_Ip28Qx8p6_0),.clk(gclk));
	jdff dff_B_IBiIzxcM6_0(.din(w_dff_B_Ip28Qx8p6_0),.dout(w_dff_B_IBiIzxcM6_0),.clk(gclk));
	jdff dff_B_p1vENyNf6_0(.din(w_dff_B_IBiIzxcM6_0),.dout(w_dff_B_p1vENyNf6_0),.clk(gclk));
	jdff dff_B_e6e7Efdy7_0(.din(w_dff_B_p1vENyNf6_0),.dout(w_dff_B_e6e7Efdy7_0),.clk(gclk));
	jdff dff_B_XgCxSUBy2_0(.din(w_dff_B_e6e7Efdy7_0),.dout(w_dff_B_XgCxSUBy2_0),.clk(gclk));
	jdff dff_B_4NoFRTwx4_0(.din(w_dff_B_XgCxSUBy2_0),.dout(w_dff_B_4NoFRTwx4_0),.clk(gclk));
	jdff dff_B_3QABQ9NP4_0(.din(w_dff_B_4NoFRTwx4_0),.dout(w_dff_B_3QABQ9NP4_0),.clk(gclk));
	jdff dff_B_vCI2geMr1_0(.din(w_dff_B_3QABQ9NP4_0),.dout(w_dff_B_vCI2geMr1_0),.clk(gclk));
	jdff dff_B_gfbD7nhv5_0(.din(w_dff_B_vCI2geMr1_0),.dout(w_dff_B_gfbD7nhv5_0),.clk(gclk));
	jdff dff_B_dqM3uZTx3_0(.din(w_dff_B_gfbD7nhv5_0),.dout(w_dff_B_dqM3uZTx3_0),.clk(gclk));
	jdff dff_B_tSAF1Htu7_0(.din(w_dff_B_dqM3uZTx3_0),.dout(w_dff_B_tSAF1Htu7_0),.clk(gclk));
	jdff dff_B_zdrtpEtz4_0(.din(w_dff_B_tSAF1Htu7_0),.dout(w_dff_B_zdrtpEtz4_0),.clk(gclk));
	jdff dff_B_gz9wlFdQ8_0(.din(w_dff_B_zdrtpEtz4_0),.dout(w_dff_B_gz9wlFdQ8_0),.clk(gclk));
	jdff dff_B_zr26dsR85_0(.din(w_dff_B_gz9wlFdQ8_0),.dout(w_dff_B_zr26dsR85_0),.clk(gclk));
	jdff dff_B_3xeDZl1F8_0(.din(w_dff_B_zr26dsR85_0),.dout(w_dff_B_3xeDZl1F8_0),.clk(gclk));
	jdff dff_B_UHpUPr7r5_0(.din(w_dff_B_3xeDZl1F8_0),.dout(w_dff_B_UHpUPr7r5_0),.clk(gclk));
	jdff dff_B_uaSvaVQI9_0(.din(w_dff_B_UHpUPr7r5_0),.dout(w_dff_B_uaSvaVQI9_0),.clk(gclk));
	jdff dff_B_OxgAFEkU9_0(.din(w_dff_B_uaSvaVQI9_0),.dout(w_dff_B_OxgAFEkU9_0),.clk(gclk));
	jdff dff_B_dkiH6k7t8_0(.din(n562),.dout(w_dff_B_dkiH6k7t8_0),.clk(gclk));
	jdff dff_B_z4Cbq2j73_0(.din(w_dff_B_dkiH6k7t8_0),.dout(w_dff_B_z4Cbq2j73_0),.clk(gclk));
	jdff dff_B_LPqaqJmf3_0(.din(w_dff_B_z4Cbq2j73_0),.dout(w_dff_B_LPqaqJmf3_0),.clk(gclk));
	jdff dff_B_GAEIV1Ke6_0(.din(w_dff_B_LPqaqJmf3_0),.dout(w_dff_B_GAEIV1Ke6_0),.clk(gclk));
	jdff dff_B_ZBzNic8q8_0(.din(w_dff_B_GAEIV1Ke6_0),.dout(w_dff_B_ZBzNic8q8_0),.clk(gclk));
	jdff dff_B_m43XMzew6_0(.din(w_dff_B_ZBzNic8q8_0),.dout(w_dff_B_m43XMzew6_0),.clk(gclk));
	jdff dff_B_6UDn0Zez6_0(.din(w_dff_B_m43XMzew6_0),.dout(w_dff_B_6UDn0Zez6_0),.clk(gclk));
	jdff dff_B_LCH7t6FF8_0(.din(w_dff_B_6UDn0Zez6_0),.dout(w_dff_B_LCH7t6FF8_0),.clk(gclk));
	jdff dff_B_PKAztZiL9_0(.din(w_dff_B_LCH7t6FF8_0),.dout(w_dff_B_PKAztZiL9_0),.clk(gclk));
	jdff dff_B_IN3uvrr45_0(.din(w_dff_B_PKAztZiL9_0),.dout(w_dff_B_IN3uvrr45_0),.clk(gclk));
	jdff dff_B_zbrV0bNw3_0(.din(w_dff_B_IN3uvrr45_0),.dout(w_dff_B_zbrV0bNw3_0),.clk(gclk));
	jdff dff_B_KO9pfjW92_0(.din(w_dff_B_zbrV0bNw3_0),.dout(w_dff_B_KO9pfjW92_0),.clk(gclk));
	jdff dff_B_TTIbsp2K4_0(.din(w_dff_B_KO9pfjW92_0),.dout(w_dff_B_TTIbsp2K4_0),.clk(gclk));
	jdff dff_B_72OJvSzO1_0(.din(w_dff_B_TTIbsp2K4_0),.dout(w_dff_B_72OJvSzO1_0),.clk(gclk));
	jdff dff_B_54EoEQuC5_0(.din(w_dff_B_72OJvSzO1_0),.dout(w_dff_B_54EoEQuC5_0),.clk(gclk));
	jdff dff_B_lrZU6iDG3_0(.din(w_dff_B_54EoEQuC5_0),.dout(w_dff_B_lrZU6iDG3_0),.clk(gclk));
	jdff dff_B_3GxWQUJx9_0(.din(w_dff_B_lrZU6iDG3_0),.dout(w_dff_B_3GxWQUJx9_0),.clk(gclk));
	jdff dff_B_0mxDNauX0_0(.din(w_dff_B_3GxWQUJx9_0),.dout(w_dff_B_0mxDNauX0_0),.clk(gclk));
	jdff dff_B_OynKnJcY1_0(.din(w_dff_B_0mxDNauX0_0),.dout(w_dff_B_OynKnJcY1_0),.clk(gclk));
	jdff dff_B_uNe84uCH6_0(.din(w_dff_B_OynKnJcY1_0),.dout(w_dff_B_uNe84uCH6_0),.clk(gclk));
	jdff dff_B_Jho5xa795_0(.din(w_dff_B_uNe84uCH6_0),.dout(w_dff_B_Jho5xa795_0),.clk(gclk));
	jdff dff_B_i7znTgNA4_0(.din(w_dff_B_Jho5xa795_0),.dout(w_dff_B_i7znTgNA4_0),.clk(gclk));
	jdff dff_B_KhgyE6Vj7_0(.din(w_dff_B_i7znTgNA4_0),.dout(w_dff_B_KhgyE6Vj7_0),.clk(gclk));
	jdff dff_B_0zVq1WWZ9_0(.din(w_dff_B_KhgyE6Vj7_0),.dout(w_dff_B_0zVq1WWZ9_0),.clk(gclk));
	jdff dff_B_dZKk2RTS0_0(.din(w_dff_B_0zVq1WWZ9_0),.dout(w_dff_B_dZKk2RTS0_0),.clk(gclk));
	jdff dff_B_n0Hq61xH4_0(.din(w_dff_B_dZKk2RTS0_0),.dout(w_dff_B_n0Hq61xH4_0),.clk(gclk));
	jdff dff_B_OOSrtPox1_0(.din(w_dff_B_n0Hq61xH4_0),.dout(w_dff_B_OOSrtPox1_0),.clk(gclk));
	jdff dff_B_s93P21LQ8_0(.din(w_dff_B_OOSrtPox1_0),.dout(w_dff_B_s93P21LQ8_0),.clk(gclk));
	jdff dff_B_0NQGDTyH9_0(.din(w_dff_B_s93P21LQ8_0),.dout(w_dff_B_0NQGDTyH9_0),.clk(gclk));
	jdff dff_B_CCeYgj5q7_0(.din(n568),.dout(w_dff_B_CCeYgj5q7_0),.clk(gclk));
	jdff dff_B_Gz5busOc2_0(.din(w_dff_B_CCeYgj5q7_0),.dout(w_dff_B_Gz5busOc2_0),.clk(gclk));
	jdff dff_B_hMKQex3R8_0(.din(w_dff_B_Gz5busOc2_0),.dout(w_dff_B_hMKQex3R8_0),.clk(gclk));
	jdff dff_B_k4jQfFFP9_0(.din(w_dff_B_hMKQex3R8_0),.dout(w_dff_B_k4jQfFFP9_0),.clk(gclk));
	jdff dff_B_A99Gj2sq0_0(.din(w_dff_B_k4jQfFFP9_0),.dout(w_dff_B_A99Gj2sq0_0),.clk(gclk));
	jdff dff_B_YrJgWPz39_0(.din(w_dff_B_A99Gj2sq0_0),.dout(w_dff_B_YrJgWPz39_0),.clk(gclk));
	jdff dff_B_0hPskeWw2_0(.din(w_dff_B_YrJgWPz39_0),.dout(w_dff_B_0hPskeWw2_0),.clk(gclk));
	jdff dff_B_oN2xRZGe8_0(.din(w_dff_B_0hPskeWw2_0),.dout(w_dff_B_oN2xRZGe8_0),.clk(gclk));
	jdff dff_B_ZXhiPTGj0_0(.din(w_dff_B_oN2xRZGe8_0),.dout(w_dff_B_ZXhiPTGj0_0),.clk(gclk));
	jdff dff_B_aqCZpPbu3_0(.din(w_dff_B_ZXhiPTGj0_0),.dout(w_dff_B_aqCZpPbu3_0),.clk(gclk));
	jdff dff_B_3KNPvgzG6_0(.din(w_dff_B_aqCZpPbu3_0),.dout(w_dff_B_3KNPvgzG6_0),.clk(gclk));
	jdff dff_B_tzFPXq6z6_0(.din(w_dff_B_3KNPvgzG6_0),.dout(w_dff_B_tzFPXq6z6_0),.clk(gclk));
	jdff dff_B_TYP5FPPc8_0(.din(w_dff_B_tzFPXq6z6_0),.dout(w_dff_B_TYP5FPPc8_0),.clk(gclk));
	jdff dff_B_vNHFGvCb7_0(.din(w_dff_B_TYP5FPPc8_0),.dout(w_dff_B_vNHFGvCb7_0),.clk(gclk));
	jdff dff_B_tnLjToGI0_0(.din(w_dff_B_vNHFGvCb7_0),.dout(w_dff_B_tnLjToGI0_0),.clk(gclk));
	jdff dff_B_GowKRS1P7_0(.din(w_dff_B_tnLjToGI0_0),.dout(w_dff_B_GowKRS1P7_0),.clk(gclk));
	jdff dff_B_0Sxd84Kr2_0(.din(w_dff_B_GowKRS1P7_0),.dout(w_dff_B_0Sxd84Kr2_0),.clk(gclk));
	jdff dff_B_JJ5Bdcte9_0(.din(w_dff_B_0Sxd84Kr2_0),.dout(w_dff_B_JJ5Bdcte9_0),.clk(gclk));
	jdff dff_B_6OPNAG569_0(.din(w_dff_B_JJ5Bdcte9_0),.dout(w_dff_B_6OPNAG569_0),.clk(gclk));
	jdff dff_B_DL50Llf17_0(.din(w_dff_B_6OPNAG569_0),.dout(w_dff_B_DL50Llf17_0),.clk(gclk));
	jdff dff_B_26ONQgce5_0(.din(w_dff_B_DL50Llf17_0),.dout(w_dff_B_26ONQgce5_0),.clk(gclk));
	jdff dff_B_hO1wFjem1_0(.din(w_dff_B_26ONQgce5_0),.dout(w_dff_B_hO1wFjem1_0),.clk(gclk));
	jdff dff_B_uPgWI5GI7_0(.din(w_dff_B_hO1wFjem1_0),.dout(w_dff_B_uPgWI5GI7_0),.clk(gclk));
	jdff dff_B_k9J5o1lq9_0(.din(w_dff_B_uPgWI5GI7_0),.dout(w_dff_B_k9J5o1lq9_0),.clk(gclk));
	jdff dff_B_NdhviSid4_0(.din(w_dff_B_k9J5o1lq9_0),.dout(w_dff_B_NdhviSid4_0),.clk(gclk));
	jdff dff_B_VuvCKVB06_0(.din(w_dff_B_NdhviSid4_0),.dout(w_dff_B_VuvCKVB06_0),.clk(gclk));
	jdff dff_B_QoUC1qbN7_0(.din(w_dff_B_VuvCKVB06_0),.dout(w_dff_B_QoUC1qbN7_0),.clk(gclk));
	jdff dff_B_wiC1SogH4_0(.din(w_dff_B_QoUC1qbN7_0),.dout(w_dff_B_wiC1SogH4_0),.clk(gclk));
	jdff dff_B_rcaV8e814_0(.din(w_dff_B_wiC1SogH4_0),.dout(w_dff_B_rcaV8e814_0),.clk(gclk));
	jdff dff_B_yCmWmTN77_0(.din(w_dff_B_rcaV8e814_0),.dout(w_dff_B_yCmWmTN77_0),.clk(gclk));
	jdff dff_B_A1PhRP3d7_0(.din(n574),.dout(w_dff_B_A1PhRP3d7_0),.clk(gclk));
	jdff dff_B_4hgOkIVd0_0(.din(w_dff_B_A1PhRP3d7_0),.dout(w_dff_B_4hgOkIVd0_0),.clk(gclk));
	jdff dff_B_EVbbXczU0_0(.din(w_dff_B_4hgOkIVd0_0),.dout(w_dff_B_EVbbXczU0_0),.clk(gclk));
	jdff dff_B_zQBLhk6e1_0(.din(w_dff_B_EVbbXczU0_0),.dout(w_dff_B_zQBLhk6e1_0),.clk(gclk));
	jdff dff_B_083QX3LK8_0(.din(w_dff_B_zQBLhk6e1_0),.dout(w_dff_B_083QX3LK8_0),.clk(gclk));
	jdff dff_B_ApYemFwo3_0(.din(w_dff_B_083QX3LK8_0),.dout(w_dff_B_ApYemFwo3_0),.clk(gclk));
	jdff dff_B_A8ANUUMb0_0(.din(w_dff_B_ApYemFwo3_0),.dout(w_dff_B_A8ANUUMb0_0),.clk(gclk));
	jdff dff_B_Kme2bApf0_0(.din(w_dff_B_A8ANUUMb0_0),.dout(w_dff_B_Kme2bApf0_0),.clk(gclk));
	jdff dff_B_s4c3ypYF6_0(.din(w_dff_B_Kme2bApf0_0),.dout(w_dff_B_s4c3ypYF6_0),.clk(gclk));
	jdff dff_B_CsOBqpYH6_0(.din(w_dff_B_s4c3ypYF6_0),.dout(w_dff_B_CsOBqpYH6_0),.clk(gclk));
	jdff dff_B_2B8BQQnX5_0(.din(w_dff_B_CsOBqpYH6_0),.dout(w_dff_B_2B8BQQnX5_0),.clk(gclk));
	jdff dff_B_edRF8MSF4_0(.din(w_dff_B_2B8BQQnX5_0),.dout(w_dff_B_edRF8MSF4_0),.clk(gclk));
	jdff dff_B_Qt58gf8K4_0(.din(w_dff_B_edRF8MSF4_0),.dout(w_dff_B_Qt58gf8K4_0),.clk(gclk));
	jdff dff_B_aJnvWoRe3_0(.din(w_dff_B_Qt58gf8K4_0),.dout(w_dff_B_aJnvWoRe3_0),.clk(gclk));
	jdff dff_B_WgEnrC709_0(.din(w_dff_B_aJnvWoRe3_0),.dout(w_dff_B_WgEnrC709_0),.clk(gclk));
	jdff dff_B_MKaPkcfQ1_0(.din(w_dff_B_WgEnrC709_0),.dout(w_dff_B_MKaPkcfQ1_0),.clk(gclk));
	jdff dff_B_7m3sKTyf9_0(.din(w_dff_B_MKaPkcfQ1_0),.dout(w_dff_B_7m3sKTyf9_0),.clk(gclk));
	jdff dff_B_2abs3PCw6_0(.din(w_dff_B_7m3sKTyf9_0),.dout(w_dff_B_2abs3PCw6_0),.clk(gclk));
	jdff dff_B_SJA6YXzi3_0(.din(w_dff_B_2abs3PCw6_0),.dout(w_dff_B_SJA6YXzi3_0),.clk(gclk));
	jdff dff_B_pFTfDD0O2_0(.din(w_dff_B_SJA6YXzi3_0),.dout(w_dff_B_pFTfDD0O2_0),.clk(gclk));
	jdff dff_B_GOi7Ebvm7_0(.din(w_dff_B_pFTfDD0O2_0),.dout(w_dff_B_GOi7Ebvm7_0),.clk(gclk));
	jdff dff_B_pFRLx8Ze0_0(.din(w_dff_B_GOi7Ebvm7_0),.dout(w_dff_B_pFRLx8Ze0_0),.clk(gclk));
	jdff dff_B_8TXVcxsV2_0(.din(w_dff_B_pFRLx8Ze0_0),.dout(w_dff_B_8TXVcxsV2_0),.clk(gclk));
	jdff dff_B_NVZbxlKC0_0(.din(w_dff_B_8TXVcxsV2_0),.dout(w_dff_B_NVZbxlKC0_0),.clk(gclk));
	jdff dff_B_NmIm7Vs78_0(.din(w_dff_B_NVZbxlKC0_0),.dout(w_dff_B_NmIm7Vs78_0),.clk(gclk));
	jdff dff_B_gzUCBXVb7_0(.din(w_dff_B_NmIm7Vs78_0),.dout(w_dff_B_gzUCBXVb7_0),.clk(gclk));
	jdff dff_B_TYDZLs2Y9_0(.din(w_dff_B_gzUCBXVb7_0),.dout(w_dff_B_TYDZLs2Y9_0),.clk(gclk));
	jdff dff_B_dbkJUWm80_0(.din(w_dff_B_TYDZLs2Y9_0),.dout(w_dff_B_dbkJUWm80_0),.clk(gclk));
	jdff dff_B_mLXkMxVF2_0(.din(w_dff_B_dbkJUWm80_0),.dout(w_dff_B_mLXkMxVF2_0),.clk(gclk));
	jdff dff_B_h4lQj65l7_0(.din(w_dff_B_mLXkMxVF2_0),.dout(w_dff_B_h4lQj65l7_0),.clk(gclk));
	jdff dff_B_FPJBFbiz2_0(.din(w_dff_B_h4lQj65l7_0),.dout(w_dff_B_FPJBFbiz2_0),.clk(gclk));
	jdff dff_B_46awi8rt3_0(.din(n580),.dout(w_dff_B_46awi8rt3_0),.clk(gclk));
	jdff dff_B_YxVlzGpd7_0(.din(w_dff_B_46awi8rt3_0),.dout(w_dff_B_YxVlzGpd7_0),.clk(gclk));
	jdff dff_B_R1nitSyc6_0(.din(w_dff_B_YxVlzGpd7_0),.dout(w_dff_B_R1nitSyc6_0),.clk(gclk));
	jdff dff_B_hqbYiICS9_0(.din(w_dff_B_R1nitSyc6_0),.dout(w_dff_B_hqbYiICS9_0),.clk(gclk));
	jdff dff_B_pg7DmpEf7_0(.din(w_dff_B_hqbYiICS9_0),.dout(w_dff_B_pg7DmpEf7_0),.clk(gclk));
	jdff dff_B_pjKjhEQg4_0(.din(w_dff_B_pg7DmpEf7_0),.dout(w_dff_B_pjKjhEQg4_0),.clk(gclk));
	jdff dff_B_TVag2PWB0_0(.din(w_dff_B_pjKjhEQg4_0),.dout(w_dff_B_TVag2PWB0_0),.clk(gclk));
	jdff dff_B_GnQcVHrg6_0(.din(w_dff_B_TVag2PWB0_0),.dout(w_dff_B_GnQcVHrg6_0),.clk(gclk));
	jdff dff_B_tTV78Fti3_0(.din(w_dff_B_GnQcVHrg6_0),.dout(w_dff_B_tTV78Fti3_0),.clk(gclk));
	jdff dff_B_gF7AmbBz8_0(.din(w_dff_B_tTV78Fti3_0),.dout(w_dff_B_gF7AmbBz8_0),.clk(gclk));
	jdff dff_B_Z6KugE428_0(.din(w_dff_B_gF7AmbBz8_0),.dout(w_dff_B_Z6KugE428_0),.clk(gclk));
	jdff dff_B_JM0bsTRR3_0(.din(w_dff_B_Z6KugE428_0),.dout(w_dff_B_JM0bsTRR3_0),.clk(gclk));
	jdff dff_B_vBGMu0PG3_0(.din(w_dff_B_JM0bsTRR3_0),.dout(w_dff_B_vBGMu0PG3_0),.clk(gclk));
	jdff dff_B_6oNWWjBK6_0(.din(w_dff_B_vBGMu0PG3_0),.dout(w_dff_B_6oNWWjBK6_0),.clk(gclk));
	jdff dff_B_K4cteTvu4_0(.din(w_dff_B_6oNWWjBK6_0),.dout(w_dff_B_K4cteTvu4_0),.clk(gclk));
	jdff dff_B_deVqox1S0_0(.din(w_dff_B_K4cteTvu4_0),.dout(w_dff_B_deVqox1S0_0),.clk(gclk));
	jdff dff_B_HJ0VgJV42_0(.din(w_dff_B_deVqox1S0_0),.dout(w_dff_B_HJ0VgJV42_0),.clk(gclk));
	jdff dff_B_8vVQXlFI6_0(.din(w_dff_B_HJ0VgJV42_0),.dout(w_dff_B_8vVQXlFI6_0),.clk(gclk));
	jdff dff_B_j4zovaBD6_0(.din(w_dff_B_8vVQXlFI6_0),.dout(w_dff_B_j4zovaBD6_0),.clk(gclk));
	jdff dff_B_jVByXBGy9_0(.din(w_dff_B_j4zovaBD6_0),.dout(w_dff_B_jVByXBGy9_0),.clk(gclk));
	jdff dff_B_axGXTgLD7_0(.din(w_dff_B_jVByXBGy9_0),.dout(w_dff_B_axGXTgLD7_0),.clk(gclk));
	jdff dff_B_WrhtyOD43_0(.din(w_dff_B_axGXTgLD7_0),.dout(w_dff_B_WrhtyOD43_0),.clk(gclk));
	jdff dff_B_ipdEi38z7_0(.din(w_dff_B_WrhtyOD43_0),.dout(w_dff_B_ipdEi38z7_0),.clk(gclk));
	jdff dff_B_FimWTP4Q8_0(.din(w_dff_B_ipdEi38z7_0),.dout(w_dff_B_FimWTP4Q8_0),.clk(gclk));
	jdff dff_B_sB8PY9B63_0(.din(w_dff_B_FimWTP4Q8_0),.dout(w_dff_B_sB8PY9B63_0),.clk(gclk));
	jdff dff_B_qmAnkWwJ9_0(.din(w_dff_B_sB8PY9B63_0),.dout(w_dff_B_qmAnkWwJ9_0),.clk(gclk));
	jdff dff_B_FLUg9zg23_0(.din(w_dff_B_qmAnkWwJ9_0),.dout(w_dff_B_FLUg9zg23_0),.clk(gclk));
	jdff dff_B_gsIXkc2A8_0(.din(w_dff_B_FLUg9zg23_0),.dout(w_dff_B_gsIXkc2A8_0),.clk(gclk));
	jdff dff_B_PP7MsnfQ7_0(.din(w_dff_B_gsIXkc2A8_0),.dout(w_dff_B_PP7MsnfQ7_0),.clk(gclk));
	jdff dff_B_grnNnAR75_0(.din(w_dff_B_PP7MsnfQ7_0),.dout(w_dff_B_grnNnAR75_0),.clk(gclk));
	jdff dff_B_io49pKME4_0(.din(w_dff_B_grnNnAR75_0),.dout(w_dff_B_io49pKME4_0),.clk(gclk));
	jdff dff_B_Qyetcsqv4_0(.din(w_dff_B_io49pKME4_0),.dout(w_dff_B_Qyetcsqv4_0),.clk(gclk));
	jdff dff_B_6ACmcSqa9_0(.din(n586),.dout(w_dff_B_6ACmcSqa9_0),.clk(gclk));
	jdff dff_B_1MVci1aD8_0(.din(w_dff_B_6ACmcSqa9_0),.dout(w_dff_B_1MVci1aD8_0),.clk(gclk));
	jdff dff_B_6wF6U1MK3_0(.din(w_dff_B_1MVci1aD8_0),.dout(w_dff_B_6wF6U1MK3_0),.clk(gclk));
	jdff dff_B_ek9HuBVW9_0(.din(w_dff_B_6wF6U1MK3_0),.dout(w_dff_B_ek9HuBVW9_0),.clk(gclk));
	jdff dff_B_TG8No2tq9_0(.din(w_dff_B_ek9HuBVW9_0),.dout(w_dff_B_TG8No2tq9_0),.clk(gclk));
	jdff dff_B_tLQdwva41_0(.din(w_dff_B_TG8No2tq9_0),.dout(w_dff_B_tLQdwva41_0),.clk(gclk));
	jdff dff_B_vAlmn7XW9_0(.din(w_dff_B_tLQdwva41_0),.dout(w_dff_B_vAlmn7XW9_0),.clk(gclk));
	jdff dff_B_B1g3OnwJ8_0(.din(w_dff_B_vAlmn7XW9_0),.dout(w_dff_B_B1g3OnwJ8_0),.clk(gclk));
	jdff dff_B_BpePRh142_0(.din(w_dff_B_B1g3OnwJ8_0),.dout(w_dff_B_BpePRh142_0),.clk(gclk));
	jdff dff_B_LIoqhgO00_0(.din(w_dff_B_BpePRh142_0),.dout(w_dff_B_LIoqhgO00_0),.clk(gclk));
	jdff dff_B_eRhkJaG89_0(.din(w_dff_B_LIoqhgO00_0),.dout(w_dff_B_eRhkJaG89_0),.clk(gclk));
	jdff dff_B_4dg2piZS6_0(.din(w_dff_B_eRhkJaG89_0),.dout(w_dff_B_4dg2piZS6_0),.clk(gclk));
	jdff dff_B_GLu4Oucg8_0(.din(w_dff_B_4dg2piZS6_0),.dout(w_dff_B_GLu4Oucg8_0),.clk(gclk));
	jdff dff_B_jA4rHmDX3_0(.din(w_dff_B_GLu4Oucg8_0),.dout(w_dff_B_jA4rHmDX3_0),.clk(gclk));
	jdff dff_B_oCq0iOk96_0(.din(w_dff_B_jA4rHmDX3_0),.dout(w_dff_B_oCq0iOk96_0),.clk(gclk));
	jdff dff_B_T9s7pZKK9_0(.din(w_dff_B_oCq0iOk96_0),.dout(w_dff_B_T9s7pZKK9_0),.clk(gclk));
	jdff dff_B_4lrfvYUi3_0(.din(w_dff_B_T9s7pZKK9_0),.dout(w_dff_B_4lrfvYUi3_0),.clk(gclk));
	jdff dff_B_l30poSjP7_0(.din(w_dff_B_4lrfvYUi3_0),.dout(w_dff_B_l30poSjP7_0),.clk(gclk));
	jdff dff_B_M7lWWlfJ5_0(.din(w_dff_B_l30poSjP7_0),.dout(w_dff_B_M7lWWlfJ5_0),.clk(gclk));
	jdff dff_B_BDK4HPd36_0(.din(w_dff_B_M7lWWlfJ5_0),.dout(w_dff_B_BDK4HPd36_0),.clk(gclk));
	jdff dff_B_3vTuy3Bk2_0(.din(w_dff_B_BDK4HPd36_0),.dout(w_dff_B_3vTuy3Bk2_0),.clk(gclk));
	jdff dff_B_OgM6eGew7_0(.din(w_dff_B_3vTuy3Bk2_0),.dout(w_dff_B_OgM6eGew7_0),.clk(gclk));
	jdff dff_B_5zcqJjUe4_0(.din(w_dff_B_OgM6eGew7_0),.dout(w_dff_B_5zcqJjUe4_0),.clk(gclk));
	jdff dff_B_F9Dlndwv7_0(.din(w_dff_B_5zcqJjUe4_0),.dout(w_dff_B_F9Dlndwv7_0),.clk(gclk));
	jdff dff_B_yhUe41eF5_0(.din(w_dff_B_F9Dlndwv7_0),.dout(w_dff_B_yhUe41eF5_0),.clk(gclk));
	jdff dff_B_TIbdHZ0n5_0(.din(w_dff_B_yhUe41eF5_0),.dout(w_dff_B_TIbdHZ0n5_0),.clk(gclk));
	jdff dff_B_pFCwMA4u9_0(.din(w_dff_B_TIbdHZ0n5_0),.dout(w_dff_B_pFCwMA4u9_0),.clk(gclk));
	jdff dff_B_j67cCf9n0_0(.din(w_dff_B_pFCwMA4u9_0),.dout(w_dff_B_j67cCf9n0_0),.clk(gclk));
	jdff dff_B_ZePjBeln3_0(.din(w_dff_B_j67cCf9n0_0),.dout(w_dff_B_ZePjBeln3_0),.clk(gclk));
	jdff dff_B_6lflNrwv4_0(.din(w_dff_B_ZePjBeln3_0),.dout(w_dff_B_6lflNrwv4_0),.clk(gclk));
	jdff dff_B_PxiUDOwK5_0(.din(w_dff_B_6lflNrwv4_0),.dout(w_dff_B_PxiUDOwK5_0),.clk(gclk));
	jdff dff_B_2kvT58Jr3_0(.din(w_dff_B_PxiUDOwK5_0),.dout(w_dff_B_2kvT58Jr3_0),.clk(gclk));
	jdff dff_B_WbAXqjB88_0(.din(w_dff_B_2kvT58Jr3_0),.dout(w_dff_B_WbAXqjB88_0),.clk(gclk));
	jdff dff_B_xAnXldkw5_0(.din(n592),.dout(w_dff_B_xAnXldkw5_0),.clk(gclk));
	jdff dff_B_OWT8tJf08_0(.din(w_dff_B_xAnXldkw5_0),.dout(w_dff_B_OWT8tJf08_0),.clk(gclk));
	jdff dff_B_rGvlmkGX1_0(.din(w_dff_B_OWT8tJf08_0),.dout(w_dff_B_rGvlmkGX1_0),.clk(gclk));
	jdff dff_B_coGLsrq49_0(.din(w_dff_B_rGvlmkGX1_0),.dout(w_dff_B_coGLsrq49_0),.clk(gclk));
	jdff dff_B_G9MmrI7b3_0(.din(w_dff_B_coGLsrq49_0),.dout(w_dff_B_G9MmrI7b3_0),.clk(gclk));
	jdff dff_B_S9MMtSVj8_0(.din(w_dff_B_G9MmrI7b3_0),.dout(w_dff_B_S9MMtSVj8_0),.clk(gclk));
	jdff dff_B_8tGXunFm6_0(.din(w_dff_B_S9MMtSVj8_0),.dout(w_dff_B_8tGXunFm6_0),.clk(gclk));
	jdff dff_B_0A9VS7KY5_0(.din(w_dff_B_8tGXunFm6_0),.dout(w_dff_B_0A9VS7KY5_0),.clk(gclk));
	jdff dff_B_rk3N94Bx3_0(.din(w_dff_B_0A9VS7KY5_0),.dout(w_dff_B_rk3N94Bx3_0),.clk(gclk));
	jdff dff_B_D8I1CfTd3_0(.din(w_dff_B_rk3N94Bx3_0),.dout(w_dff_B_D8I1CfTd3_0),.clk(gclk));
	jdff dff_B_7T9ullDj9_0(.din(w_dff_B_D8I1CfTd3_0),.dout(w_dff_B_7T9ullDj9_0),.clk(gclk));
	jdff dff_B_Ek0OTX2n3_0(.din(w_dff_B_7T9ullDj9_0),.dout(w_dff_B_Ek0OTX2n3_0),.clk(gclk));
	jdff dff_B_HnEY1rzJ7_0(.din(w_dff_B_Ek0OTX2n3_0),.dout(w_dff_B_HnEY1rzJ7_0),.clk(gclk));
	jdff dff_B_Pioerm9g5_0(.din(w_dff_B_HnEY1rzJ7_0),.dout(w_dff_B_Pioerm9g5_0),.clk(gclk));
	jdff dff_B_3AUJECEi4_0(.din(w_dff_B_Pioerm9g5_0),.dout(w_dff_B_3AUJECEi4_0),.clk(gclk));
	jdff dff_B_2N4y2pWX4_0(.din(w_dff_B_3AUJECEi4_0),.dout(w_dff_B_2N4y2pWX4_0),.clk(gclk));
	jdff dff_B_BA1I6UGy9_0(.din(w_dff_B_2N4y2pWX4_0),.dout(w_dff_B_BA1I6UGy9_0),.clk(gclk));
	jdff dff_B_F0uHJ1ep8_0(.din(w_dff_B_BA1I6UGy9_0),.dout(w_dff_B_F0uHJ1ep8_0),.clk(gclk));
	jdff dff_B_42e3FdGp2_0(.din(w_dff_B_F0uHJ1ep8_0),.dout(w_dff_B_42e3FdGp2_0),.clk(gclk));
	jdff dff_B_0wKyjJXR3_0(.din(w_dff_B_42e3FdGp2_0),.dout(w_dff_B_0wKyjJXR3_0),.clk(gclk));
	jdff dff_B_wyriGQ280_0(.din(w_dff_B_0wKyjJXR3_0),.dout(w_dff_B_wyriGQ280_0),.clk(gclk));
	jdff dff_B_7ZhPNr8I9_0(.din(w_dff_B_wyriGQ280_0),.dout(w_dff_B_7ZhPNr8I9_0),.clk(gclk));
	jdff dff_B_v81X9vVW2_0(.din(w_dff_B_7ZhPNr8I9_0),.dout(w_dff_B_v81X9vVW2_0),.clk(gclk));
	jdff dff_B_oErTCF311_0(.din(w_dff_B_v81X9vVW2_0),.dout(w_dff_B_oErTCF311_0),.clk(gclk));
	jdff dff_B_VWYwBy3A1_0(.din(w_dff_B_oErTCF311_0),.dout(w_dff_B_VWYwBy3A1_0),.clk(gclk));
	jdff dff_B_9zbAgTAq8_0(.din(w_dff_B_VWYwBy3A1_0),.dout(w_dff_B_9zbAgTAq8_0),.clk(gclk));
	jdff dff_B_aavi7VYB8_0(.din(w_dff_B_9zbAgTAq8_0),.dout(w_dff_B_aavi7VYB8_0),.clk(gclk));
	jdff dff_B_4ufKLp5C0_0(.din(w_dff_B_aavi7VYB8_0),.dout(w_dff_B_4ufKLp5C0_0),.clk(gclk));
	jdff dff_B_WYO79c0j5_0(.din(w_dff_B_4ufKLp5C0_0),.dout(w_dff_B_WYO79c0j5_0),.clk(gclk));
	jdff dff_B_KvlHQr7L6_0(.din(w_dff_B_WYO79c0j5_0),.dout(w_dff_B_KvlHQr7L6_0),.clk(gclk));
	jdff dff_B_UaQtGvqK4_0(.din(w_dff_B_KvlHQr7L6_0),.dout(w_dff_B_UaQtGvqK4_0),.clk(gclk));
	jdff dff_B_jkPkgNyK5_0(.din(w_dff_B_UaQtGvqK4_0),.dout(w_dff_B_jkPkgNyK5_0),.clk(gclk));
	jdff dff_B_iZCaN07y6_0(.din(w_dff_B_jkPkgNyK5_0),.dout(w_dff_B_iZCaN07y6_0),.clk(gclk));
	jdff dff_B_tTqoaoGw3_0(.din(w_dff_B_iZCaN07y6_0),.dout(w_dff_B_tTqoaoGw3_0),.clk(gclk));
	jdff dff_B_6CAW1Bi71_0(.din(n598),.dout(w_dff_B_6CAW1Bi71_0),.clk(gclk));
	jdff dff_B_EYQ4Ugbh9_0(.din(w_dff_B_6CAW1Bi71_0),.dout(w_dff_B_EYQ4Ugbh9_0),.clk(gclk));
	jdff dff_B_khqpYdj28_0(.din(w_dff_B_EYQ4Ugbh9_0),.dout(w_dff_B_khqpYdj28_0),.clk(gclk));
	jdff dff_B_BG4MiUsI7_0(.din(w_dff_B_khqpYdj28_0),.dout(w_dff_B_BG4MiUsI7_0),.clk(gclk));
	jdff dff_B_2ZdJIpg02_0(.din(w_dff_B_BG4MiUsI7_0),.dout(w_dff_B_2ZdJIpg02_0),.clk(gclk));
	jdff dff_B_LzvqDQab8_0(.din(w_dff_B_2ZdJIpg02_0),.dout(w_dff_B_LzvqDQab8_0),.clk(gclk));
	jdff dff_B_bYQSosfp4_0(.din(w_dff_B_LzvqDQab8_0),.dout(w_dff_B_bYQSosfp4_0),.clk(gclk));
	jdff dff_B_vWFugr9c6_0(.din(w_dff_B_bYQSosfp4_0),.dout(w_dff_B_vWFugr9c6_0),.clk(gclk));
	jdff dff_B_cpzefdg00_0(.din(w_dff_B_vWFugr9c6_0),.dout(w_dff_B_cpzefdg00_0),.clk(gclk));
	jdff dff_B_gTqNlWi62_0(.din(w_dff_B_cpzefdg00_0),.dout(w_dff_B_gTqNlWi62_0),.clk(gclk));
	jdff dff_B_bAB7dH8h6_0(.din(w_dff_B_gTqNlWi62_0),.dout(w_dff_B_bAB7dH8h6_0),.clk(gclk));
	jdff dff_B_tiKsYfsy3_0(.din(w_dff_B_bAB7dH8h6_0),.dout(w_dff_B_tiKsYfsy3_0),.clk(gclk));
	jdff dff_B_XwKEVTyN3_0(.din(w_dff_B_tiKsYfsy3_0),.dout(w_dff_B_XwKEVTyN3_0),.clk(gclk));
	jdff dff_B_lXZ4Dx5C8_0(.din(w_dff_B_XwKEVTyN3_0),.dout(w_dff_B_lXZ4Dx5C8_0),.clk(gclk));
	jdff dff_B_YxCaTOrB6_0(.din(w_dff_B_lXZ4Dx5C8_0),.dout(w_dff_B_YxCaTOrB6_0),.clk(gclk));
	jdff dff_B_5mJJ8JPY6_0(.din(w_dff_B_YxCaTOrB6_0),.dout(w_dff_B_5mJJ8JPY6_0),.clk(gclk));
	jdff dff_B_FofErz5J6_0(.din(w_dff_B_5mJJ8JPY6_0),.dout(w_dff_B_FofErz5J6_0),.clk(gclk));
	jdff dff_B_PguLnj7c1_0(.din(w_dff_B_FofErz5J6_0),.dout(w_dff_B_PguLnj7c1_0),.clk(gclk));
	jdff dff_B_xTbGZsq29_0(.din(w_dff_B_PguLnj7c1_0),.dout(w_dff_B_xTbGZsq29_0),.clk(gclk));
	jdff dff_B_hsHJrtbC1_0(.din(w_dff_B_xTbGZsq29_0),.dout(w_dff_B_hsHJrtbC1_0),.clk(gclk));
	jdff dff_B_uRsQPYt34_0(.din(w_dff_B_hsHJrtbC1_0),.dout(w_dff_B_uRsQPYt34_0),.clk(gclk));
	jdff dff_B_sY4gQZYM2_0(.din(w_dff_B_uRsQPYt34_0),.dout(w_dff_B_sY4gQZYM2_0),.clk(gclk));
	jdff dff_B_OGbwYld46_0(.din(w_dff_B_sY4gQZYM2_0),.dout(w_dff_B_OGbwYld46_0),.clk(gclk));
	jdff dff_B_qysdxons0_0(.din(w_dff_B_OGbwYld46_0),.dout(w_dff_B_qysdxons0_0),.clk(gclk));
	jdff dff_B_6UlW1OEO3_0(.din(w_dff_B_qysdxons0_0),.dout(w_dff_B_6UlW1OEO3_0),.clk(gclk));
	jdff dff_B_dXRCq7HD9_0(.din(w_dff_B_6UlW1OEO3_0),.dout(w_dff_B_dXRCq7HD9_0),.clk(gclk));
	jdff dff_B_TTTTHqOE9_0(.din(w_dff_B_dXRCq7HD9_0),.dout(w_dff_B_TTTTHqOE9_0),.clk(gclk));
	jdff dff_B_givM90s49_0(.din(w_dff_B_TTTTHqOE9_0),.dout(w_dff_B_givM90s49_0),.clk(gclk));
	jdff dff_B_1betfp328_0(.din(w_dff_B_givM90s49_0),.dout(w_dff_B_1betfp328_0),.clk(gclk));
	jdff dff_B_pJYiDME72_0(.din(w_dff_B_1betfp328_0),.dout(w_dff_B_pJYiDME72_0),.clk(gclk));
	jdff dff_B_noqs5PZE5_0(.din(w_dff_B_pJYiDME72_0),.dout(w_dff_B_noqs5PZE5_0),.clk(gclk));
	jdff dff_B_SyUyvPfc1_0(.din(w_dff_B_noqs5PZE5_0),.dout(w_dff_B_SyUyvPfc1_0),.clk(gclk));
	jdff dff_B_BaTwVzpv6_0(.din(w_dff_B_SyUyvPfc1_0),.dout(w_dff_B_BaTwVzpv6_0),.clk(gclk));
	jdff dff_B_9R7bTIZc0_0(.din(w_dff_B_BaTwVzpv6_0),.dout(w_dff_B_9R7bTIZc0_0),.clk(gclk));
	jdff dff_B_OVSEBGFt8_0(.din(w_dff_B_9R7bTIZc0_0),.dout(w_dff_B_OVSEBGFt8_0),.clk(gclk));
	jdff dff_B_lg7sDa4m3_0(.din(n604),.dout(w_dff_B_lg7sDa4m3_0),.clk(gclk));
	jdff dff_B_kIU5wzMk4_0(.din(w_dff_B_lg7sDa4m3_0),.dout(w_dff_B_kIU5wzMk4_0),.clk(gclk));
	jdff dff_B_oJ02hao28_0(.din(w_dff_B_kIU5wzMk4_0),.dout(w_dff_B_oJ02hao28_0),.clk(gclk));
	jdff dff_B_3s2YdROj7_0(.din(w_dff_B_oJ02hao28_0),.dout(w_dff_B_3s2YdROj7_0),.clk(gclk));
	jdff dff_B_SCoeVMVN6_0(.din(w_dff_B_3s2YdROj7_0),.dout(w_dff_B_SCoeVMVN6_0),.clk(gclk));
	jdff dff_B_cNZ24YRu3_0(.din(w_dff_B_SCoeVMVN6_0),.dout(w_dff_B_cNZ24YRu3_0),.clk(gclk));
	jdff dff_B_8ayMfOmq6_0(.din(w_dff_B_cNZ24YRu3_0),.dout(w_dff_B_8ayMfOmq6_0),.clk(gclk));
	jdff dff_B_hTGzDXm21_0(.din(w_dff_B_8ayMfOmq6_0),.dout(w_dff_B_hTGzDXm21_0),.clk(gclk));
	jdff dff_B_DjEeqKiM9_0(.din(w_dff_B_hTGzDXm21_0),.dout(w_dff_B_DjEeqKiM9_0),.clk(gclk));
	jdff dff_B_UbNdYlP46_0(.din(w_dff_B_DjEeqKiM9_0),.dout(w_dff_B_UbNdYlP46_0),.clk(gclk));
	jdff dff_B_ryaiLADL4_0(.din(w_dff_B_UbNdYlP46_0),.dout(w_dff_B_ryaiLADL4_0),.clk(gclk));
	jdff dff_B_wocJxgUa1_0(.din(w_dff_B_ryaiLADL4_0),.dout(w_dff_B_wocJxgUa1_0),.clk(gclk));
	jdff dff_B_lZ6ownHW3_0(.din(w_dff_B_wocJxgUa1_0),.dout(w_dff_B_lZ6ownHW3_0),.clk(gclk));
	jdff dff_B_zsLlWmoh9_0(.din(w_dff_B_lZ6ownHW3_0),.dout(w_dff_B_zsLlWmoh9_0),.clk(gclk));
	jdff dff_B_s6OFruit2_0(.din(w_dff_B_zsLlWmoh9_0),.dout(w_dff_B_s6OFruit2_0),.clk(gclk));
	jdff dff_B_jl4MHObG2_0(.din(w_dff_B_s6OFruit2_0),.dout(w_dff_B_jl4MHObG2_0),.clk(gclk));
	jdff dff_B_lEiK5sDf6_0(.din(w_dff_B_jl4MHObG2_0),.dout(w_dff_B_lEiK5sDf6_0),.clk(gclk));
	jdff dff_B_rleuJbWp1_0(.din(w_dff_B_lEiK5sDf6_0),.dout(w_dff_B_rleuJbWp1_0),.clk(gclk));
	jdff dff_B_mT8kbtBw0_0(.din(w_dff_B_rleuJbWp1_0),.dout(w_dff_B_mT8kbtBw0_0),.clk(gclk));
	jdff dff_B_xxSXxaR81_0(.din(w_dff_B_mT8kbtBw0_0),.dout(w_dff_B_xxSXxaR81_0),.clk(gclk));
	jdff dff_B_sTanXs5T7_0(.din(w_dff_B_xxSXxaR81_0),.dout(w_dff_B_sTanXs5T7_0),.clk(gclk));
	jdff dff_B_D0J5w3ko0_0(.din(w_dff_B_sTanXs5T7_0),.dout(w_dff_B_D0J5w3ko0_0),.clk(gclk));
	jdff dff_B_fTO4tuyx8_0(.din(w_dff_B_D0J5w3ko0_0),.dout(w_dff_B_fTO4tuyx8_0),.clk(gclk));
	jdff dff_B_sPbC4NKy2_0(.din(w_dff_B_fTO4tuyx8_0),.dout(w_dff_B_sPbC4NKy2_0),.clk(gclk));
	jdff dff_B_mUKvMdNk3_0(.din(w_dff_B_sPbC4NKy2_0),.dout(w_dff_B_mUKvMdNk3_0),.clk(gclk));
	jdff dff_B_5v9uNf036_0(.din(w_dff_B_mUKvMdNk3_0),.dout(w_dff_B_5v9uNf036_0),.clk(gclk));
	jdff dff_B_SUsZha0H6_0(.din(w_dff_B_5v9uNf036_0),.dout(w_dff_B_SUsZha0H6_0),.clk(gclk));
	jdff dff_B_JNn35Cqb3_0(.din(w_dff_B_SUsZha0H6_0),.dout(w_dff_B_JNn35Cqb3_0),.clk(gclk));
	jdff dff_B_govLfac43_0(.din(w_dff_B_JNn35Cqb3_0),.dout(w_dff_B_govLfac43_0),.clk(gclk));
	jdff dff_B_thHdjvLH8_0(.din(w_dff_B_govLfac43_0),.dout(w_dff_B_thHdjvLH8_0),.clk(gclk));
	jdff dff_B_QvoA4r4r0_0(.din(w_dff_B_thHdjvLH8_0),.dout(w_dff_B_QvoA4r4r0_0),.clk(gclk));
	jdff dff_B_e9IJL2vo2_0(.din(w_dff_B_QvoA4r4r0_0),.dout(w_dff_B_e9IJL2vo2_0),.clk(gclk));
	jdff dff_B_tNjfnhvM2_0(.din(w_dff_B_e9IJL2vo2_0),.dout(w_dff_B_tNjfnhvM2_0),.clk(gclk));
	jdff dff_B_zRB7IH6H0_0(.din(w_dff_B_tNjfnhvM2_0),.dout(w_dff_B_zRB7IH6H0_0),.clk(gclk));
	jdff dff_B_tXzk3lcN6_0(.din(w_dff_B_zRB7IH6H0_0),.dout(w_dff_B_tXzk3lcN6_0),.clk(gclk));
	jdff dff_B_hF6XnBIn6_0(.din(w_dff_B_tXzk3lcN6_0),.dout(w_dff_B_hF6XnBIn6_0),.clk(gclk));
	jdff dff_B_s6AOjeQ90_0(.din(n610),.dout(w_dff_B_s6AOjeQ90_0),.clk(gclk));
	jdff dff_B_L6wTZ6vD3_0(.din(w_dff_B_s6AOjeQ90_0),.dout(w_dff_B_L6wTZ6vD3_0),.clk(gclk));
	jdff dff_B_QB9kMdMO7_0(.din(w_dff_B_L6wTZ6vD3_0),.dout(w_dff_B_QB9kMdMO7_0),.clk(gclk));
	jdff dff_B_D3DqKLpZ9_0(.din(w_dff_B_QB9kMdMO7_0),.dout(w_dff_B_D3DqKLpZ9_0),.clk(gclk));
	jdff dff_B_DUjdZrWQ9_0(.din(w_dff_B_D3DqKLpZ9_0),.dout(w_dff_B_DUjdZrWQ9_0),.clk(gclk));
	jdff dff_B_Q97YAQfT5_0(.din(w_dff_B_DUjdZrWQ9_0),.dout(w_dff_B_Q97YAQfT5_0),.clk(gclk));
	jdff dff_B_ZS2tzXnP3_0(.din(w_dff_B_Q97YAQfT5_0),.dout(w_dff_B_ZS2tzXnP3_0),.clk(gclk));
	jdff dff_B_SrYogtzg3_0(.din(w_dff_B_ZS2tzXnP3_0),.dout(w_dff_B_SrYogtzg3_0),.clk(gclk));
	jdff dff_B_pu9WYaR28_0(.din(w_dff_B_SrYogtzg3_0),.dout(w_dff_B_pu9WYaR28_0),.clk(gclk));
	jdff dff_B_z5QIV03e6_0(.din(w_dff_B_pu9WYaR28_0),.dout(w_dff_B_z5QIV03e6_0),.clk(gclk));
	jdff dff_B_U2tAN3m88_0(.din(w_dff_B_z5QIV03e6_0),.dout(w_dff_B_U2tAN3m88_0),.clk(gclk));
	jdff dff_B_3cS8tSB59_0(.din(w_dff_B_U2tAN3m88_0),.dout(w_dff_B_3cS8tSB59_0),.clk(gclk));
	jdff dff_B_ZxrXRBFu6_0(.din(w_dff_B_3cS8tSB59_0),.dout(w_dff_B_ZxrXRBFu6_0),.clk(gclk));
	jdff dff_B_7OInyd9t9_0(.din(w_dff_B_ZxrXRBFu6_0),.dout(w_dff_B_7OInyd9t9_0),.clk(gclk));
	jdff dff_B_GB4uq2sc2_0(.din(w_dff_B_7OInyd9t9_0),.dout(w_dff_B_GB4uq2sc2_0),.clk(gclk));
	jdff dff_B_fnlH7jW21_0(.din(w_dff_B_GB4uq2sc2_0),.dout(w_dff_B_fnlH7jW21_0),.clk(gclk));
	jdff dff_B_15OWADbF9_0(.din(w_dff_B_fnlH7jW21_0),.dout(w_dff_B_15OWADbF9_0),.clk(gclk));
	jdff dff_B_g6s6WTRR0_0(.din(w_dff_B_15OWADbF9_0),.dout(w_dff_B_g6s6WTRR0_0),.clk(gclk));
	jdff dff_B_Qpf4OHly7_0(.din(w_dff_B_g6s6WTRR0_0),.dout(w_dff_B_Qpf4OHly7_0),.clk(gclk));
	jdff dff_B_CBdxbGoT2_0(.din(w_dff_B_Qpf4OHly7_0),.dout(w_dff_B_CBdxbGoT2_0),.clk(gclk));
	jdff dff_B_SBBc6YiC2_0(.din(w_dff_B_CBdxbGoT2_0),.dout(w_dff_B_SBBc6YiC2_0),.clk(gclk));
	jdff dff_B_fspb4EEp6_0(.din(w_dff_B_SBBc6YiC2_0),.dout(w_dff_B_fspb4EEp6_0),.clk(gclk));
	jdff dff_B_iF5fgSvz1_0(.din(w_dff_B_fspb4EEp6_0),.dout(w_dff_B_iF5fgSvz1_0),.clk(gclk));
	jdff dff_B_hs8zCiMD3_0(.din(w_dff_B_iF5fgSvz1_0),.dout(w_dff_B_hs8zCiMD3_0),.clk(gclk));
	jdff dff_B_HWWyhlvB1_0(.din(w_dff_B_hs8zCiMD3_0),.dout(w_dff_B_HWWyhlvB1_0),.clk(gclk));
	jdff dff_B_uc7qRFTA6_0(.din(w_dff_B_HWWyhlvB1_0),.dout(w_dff_B_uc7qRFTA6_0),.clk(gclk));
	jdff dff_B_k51Cr8G75_0(.din(w_dff_B_uc7qRFTA6_0),.dout(w_dff_B_k51Cr8G75_0),.clk(gclk));
	jdff dff_B_xdCbxJwm1_0(.din(w_dff_B_k51Cr8G75_0),.dout(w_dff_B_xdCbxJwm1_0),.clk(gclk));
	jdff dff_B_jWgQXuk67_0(.din(w_dff_B_xdCbxJwm1_0),.dout(w_dff_B_jWgQXuk67_0),.clk(gclk));
	jdff dff_B_Y9NiFqeR8_0(.din(w_dff_B_jWgQXuk67_0),.dout(w_dff_B_Y9NiFqeR8_0),.clk(gclk));
	jdff dff_B_ZX8Ch3cj2_0(.din(w_dff_B_Y9NiFqeR8_0),.dout(w_dff_B_ZX8Ch3cj2_0),.clk(gclk));
	jdff dff_B_KVHv0EiF7_0(.din(w_dff_B_ZX8Ch3cj2_0),.dout(w_dff_B_KVHv0EiF7_0),.clk(gclk));
	jdff dff_B_5g9D2yef7_0(.din(w_dff_B_KVHv0EiF7_0),.dout(w_dff_B_5g9D2yef7_0),.clk(gclk));
	jdff dff_B_2UrH3rDD2_0(.din(w_dff_B_5g9D2yef7_0),.dout(w_dff_B_2UrH3rDD2_0),.clk(gclk));
	jdff dff_B_rLtt4ApS1_0(.din(w_dff_B_2UrH3rDD2_0),.dout(w_dff_B_rLtt4ApS1_0),.clk(gclk));
	jdff dff_B_NHVH94YY0_0(.din(w_dff_B_rLtt4ApS1_0),.dout(w_dff_B_NHVH94YY0_0),.clk(gclk));
	jdff dff_B_oTtWTlv49_0(.din(w_dff_B_NHVH94YY0_0),.dout(w_dff_B_oTtWTlv49_0),.clk(gclk));
	jdff dff_B_AYUTfkV56_0(.din(n616),.dout(w_dff_B_AYUTfkV56_0),.clk(gclk));
	jdff dff_B_Jeqwa2rS2_0(.din(w_dff_B_AYUTfkV56_0),.dout(w_dff_B_Jeqwa2rS2_0),.clk(gclk));
	jdff dff_B_CmIIuVXd6_0(.din(w_dff_B_Jeqwa2rS2_0),.dout(w_dff_B_CmIIuVXd6_0),.clk(gclk));
	jdff dff_B_qeBOZr342_0(.din(w_dff_B_CmIIuVXd6_0),.dout(w_dff_B_qeBOZr342_0),.clk(gclk));
	jdff dff_B_Cd4D5MsJ2_0(.din(w_dff_B_qeBOZr342_0),.dout(w_dff_B_Cd4D5MsJ2_0),.clk(gclk));
	jdff dff_B_iVKCevZj5_0(.din(w_dff_B_Cd4D5MsJ2_0),.dout(w_dff_B_iVKCevZj5_0),.clk(gclk));
	jdff dff_B_40uHNE919_0(.din(w_dff_B_iVKCevZj5_0),.dout(w_dff_B_40uHNE919_0),.clk(gclk));
	jdff dff_B_vV7nwnsO8_0(.din(w_dff_B_40uHNE919_0),.dout(w_dff_B_vV7nwnsO8_0),.clk(gclk));
	jdff dff_B_Bz1hKt9d8_0(.din(w_dff_B_vV7nwnsO8_0),.dout(w_dff_B_Bz1hKt9d8_0),.clk(gclk));
	jdff dff_B_Lm9wk6Sc7_0(.din(w_dff_B_Bz1hKt9d8_0),.dout(w_dff_B_Lm9wk6Sc7_0),.clk(gclk));
	jdff dff_B_4UU4N0og3_0(.din(w_dff_B_Lm9wk6Sc7_0),.dout(w_dff_B_4UU4N0og3_0),.clk(gclk));
	jdff dff_B_xPZc4aF72_0(.din(w_dff_B_4UU4N0og3_0),.dout(w_dff_B_xPZc4aF72_0),.clk(gclk));
	jdff dff_B_uU69aT6S2_0(.din(w_dff_B_xPZc4aF72_0),.dout(w_dff_B_uU69aT6S2_0),.clk(gclk));
	jdff dff_B_e1LkrerN2_0(.din(w_dff_B_uU69aT6S2_0),.dout(w_dff_B_e1LkrerN2_0),.clk(gclk));
	jdff dff_B_0e0BqBiA0_0(.din(w_dff_B_e1LkrerN2_0),.dout(w_dff_B_0e0BqBiA0_0),.clk(gclk));
	jdff dff_B_ax8tszjc8_0(.din(w_dff_B_0e0BqBiA0_0),.dout(w_dff_B_ax8tszjc8_0),.clk(gclk));
	jdff dff_B_7tedKxfT2_0(.din(w_dff_B_ax8tszjc8_0),.dout(w_dff_B_7tedKxfT2_0),.clk(gclk));
	jdff dff_B_lhocc6gV7_0(.din(w_dff_B_7tedKxfT2_0),.dout(w_dff_B_lhocc6gV7_0),.clk(gclk));
	jdff dff_B_ufiuSoxG5_0(.din(w_dff_B_lhocc6gV7_0),.dout(w_dff_B_ufiuSoxG5_0),.clk(gclk));
	jdff dff_B_lWQBwcZ00_0(.din(w_dff_B_ufiuSoxG5_0),.dout(w_dff_B_lWQBwcZ00_0),.clk(gclk));
	jdff dff_B_grNQbOGn0_0(.din(w_dff_B_lWQBwcZ00_0),.dout(w_dff_B_grNQbOGn0_0),.clk(gclk));
	jdff dff_B_5OclPB0N7_0(.din(w_dff_B_grNQbOGn0_0),.dout(w_dff_B_5OclPB0N7_0),.clk(gclk));
	jdff dff_B_LSF7P0BU3_0(.din(w_dff_B_5OclPB0N7_0),.dout(w_dff_B_LSF7P0BU3_0),.clk(gclk));
	jdff dff_B_W9ILXsuc8_0(.din(w_dff_B_LSF7P0BU3_0),.dout(w_dff_B_W9ILXsuc8_0),.clk(gclk));
	jdff dff_B_fdtXQixB2_0(.din(w_dff_B_W9ILXsuc8_0),.dout(w_dff_B_fdtXQixB2_0),.clk(gclk));
	jdff dff_B_C0i8xH2k6_0(.din(w_dff_B_fdtXQixB2_0),.dout(w_dff_B_C0i8xH2k6_0),.clk(gclk));
	jdff dff_B_C8IoAg1S2_0(.din(w_dff_B_C0i8xH2k6_0),.dout(w_dff_B_C8IoAg1S2_0),.clk(gclk));
	jdff dff_B_k0MTLwlW2_0(.din(w_dff_B_C8IoAg1S2_0),.dout(w_dff_B_k0MTLwlW2_0),.clk(gclk));
	jdff dff_B_Q3Cc1CiC7_0(.din(w_dff_B_k0MTLwlW2_0),.dout(w_dff_B_Q3Cc1CiC7_0),.clk(gclk));
	jdff dff_B_RyGgbFbM5_0(.din(w_dff_B_Q3Cc1CiC7_0),.dout(w_dff_B_RyGgbFbM5_0),.clk(gclk));
	jdff dff_B_qH2NRSqL8_0(.din(w_dff_B_RyGgbFbM5_0),.dout(w_dff_B_qH2NRSqL8_0),.clk(gclk));
	jdff dff_B_rAsMQhCl6_0(.din(w_dff_B_qH2NRSqL8_0),.dout(w_dff_B_rAsMQhCl6_0),.clk(gclk));
	jdff dff_B_BioZhb744_0(.din(w_dff_B_rAsMQhCl6_0),.dout(w_dff_B_BioZhb744_0),.clk(gclk));
	jdff dff_B_teMkegph3_0(.din(w_dff_B_BioZhb744_0),.dout(w_dff_B_teMkegph3_0),.clk(gclk));
	jdff dff_B_adBxIslw7_0(.din(w_dff_B_teMkegph3_0),.dout(w_dff_B_adBxIslw7_0),.clk(gclk));
	jdff dff_B_qD5TNK5w8_0(.din(w_dff_B_adBxIslw7_0),.dout(w_dff_B_qD5TNK5w8_0),.clk(gclk));
	jdff dff_B_6kPievLc6_0(.din(w_dff_B_qD5TNK5w8_0),.dout(w_dff_B_6kPievLc6_0),.clk(gclk));
	jdff dff_B_KlorpDbQ7_0(.din(w_dff_B_6kPievLc6_0),.dout(w_dff_B_KlorpDbQ7_0),.clk(gclk));
	jdff dff_B_XM4Wf54a0_0(.din(n622),.dout(w_dff_B_XM4Wf54a0_0),.clk(gclk));
	jdff dff_B_9S0qzORT2_0(.din(w_dff_B_XM4Wf54a0_0),.dout(w_dff_B_9S0qzORT2_0),.clk(gclk));
	jdff dff_B_bxMgh0PH8_0(.din(w_dff_B_9S0qzORT2_0),.dout(w_dff_B_bxMgh0PH8_0),.clk(gclk));
	jdff dff_B_PpbC8LTR0_0(.din(w_dff_B_bxMgh0PH8_0),.dout(w_dff_B_PpbC8LTR0_0),.clk(gclk));
	jdff dff_B_nBIJ4Egf1_0(.din(w_dff_B_PpbC8LTR0_0),.dout(w_dff_B_nBIJ4Egf1_0),.clk(gclk));
	jdff dff_B_x49YZXhk0_0(.din(w_dff_B_nBIJ4Egf1_0),.dout(w_dff_B_x49YZXhk0_0),.clk(gclk));
	jdff dff_B_Vrk1oO4i9_0(.din(w_dff_B_x49YZXhk0_0),.dout(w_dff_B_Vrk1oO4i9_0),.clk(gclk));
	jdff dff_B_ZQ5NontA8_0(.din(w_dff_B_Vrk1oO4i9_0),.dout(w_dff_B_ZQ5NontA8_0),.clk(gclk));
	jdff dff_B_8bGwQLNC7_0(.din(w_dff_B_ZQ5NontA8_0),.dout(w_dff_B_8bGwQLNC7_0),.clk(gclk));
	jdff dff_B_KlX3xzeC0_0(.din(w_dff_B_8bGwQLNC7_0),.dout(w_dff_B_KlX3xzeC0_0),.clk(gclk));
	jdff dff_B_Y76ycSQN8_0(.din(w_dff_B_KlX3xzeC0_0),.dout(w_dff_B_Y76ycSQN8_0),.clk(gclk));
	jdff dff_B_Ju8ucWYV8_0(.din(w_dff_B_Y76ycSQN8_0),.dout(w_dff_B_Ju8ucWYV8_0),.clk(gclk));
	jdff dff_B_6ydS0C4u0_0(.din(w_dff_B_Ju8ucWYV8_0),.dout(w_dff_B_6ydS0C4u0_0),.clk(gclk));
	jdff dff_B_FccqzLpO7_0(.din(w_dff_B_6ydS0C4u0_0),.dout(w_dff_B_FccqzLpO7_0),.clk(gclk));
	jdff dff_B_ksDi6erO7_0(.din(w_dff_B_FccqzLpO7_0),.dout(w_dff_B_ksDi6erO7_0),.clk(gclk));
	jdff dff_B_AoPXskoG4_0(.din(w_dff_B_ksDi6erO7_0),.dout(w_dff_B_AoPXskoG4_0),.clk(gclk));
	jdff dff_B_LzZ7765N4_0(.din(w_dff_B_AoPXskoG4_0),.dout(w_dff_B_LzZ7765N4_0),.clk(gclk));
	jdff dff_B_19oxLLtM3_0(.din(w_dff_B_LzZ7765N4_0),.dout(w_dff_B_19oxLLtM3_0),.clk(gclk));
	jdff dff_B_SRRDBq9q4_0(.din(w_dff_B_19oxLLtM3_0),.dout(w_dff_B_SRRDBq9q4_0),.clk(gclk));
	jdff dff_B_FMq2Bf1y1_0(.din(w_dff_B_SRRDBq9q4_0),.dout(w_dff_B_FMq2Bf1y1_0),.clk(gclk));
	jdff dff_B_HUPcZtHT3_0(.din(w_dff_B_FMq2Bf1y1_0),.dout(w_dff_B_HUPcZtHT3_0),.clk(gclk));
	jdff dff_B_21cZmwcf1_0(.din(w_dff_B_HUPcZtHT3_0),.dout(w_dff_B_21cZmwcf1_0),.clk(gclk));
	jdff dff_B_G0Fah0Il8_0(.din(w_dff_B_21cZmwcf1_0),.dout(w_dff_B_G0Fah0Il8_0),.clk(gclk));
	jdff dff_B_CeLIn9j27_0(.din(w_dff_B_G0Fah0Il8_0),.dout(w_dff_B_CeLIn9j27_0),.clk(gclk));
	jdff dff_B_uCccFr792_0(.din(w_dff_B_CeLIn9j27_0),.dout(w_dff_B_uCccFr792_0),.clk(gclk));
	jdff dff_B_mecpBe8W0_0(.din(w_dff_B_uCccFr792_0),.dout(w_dff_B_mecpBe8W0_0),.clk(gclk));
	jdff dff_B_p6ieCHgl2_0(.din(w_dff_B_mecpBe8W0_0),.dout(w_dff_B_p6ieCHgl2_0),.clk(gclk));
	jdff dff_B_2iccKVI69_0(.din(w_dff_B_p6ieCHgl2_0),.dout(w_dff_B_2iccKVI69_0),.clk(gclk));
	jdff dff_B_EHGcNkNL6_0(.din(w_dff_B_2iccKVI69_0),.dout(w_dff_B_EHGcNkNL6_0),.clk(gclk));
	jdff dff_B_FzDe7gxx2_0(.din(w_dff_B_EHGcNkNL6_0),.dout(w_dff_B_FzDe7gxx2_0),.clk(gclk));
	jdff dff_B_zYDVsHBR5_0(.din(w_dff_B_FzDe7gxx2_0),.dout(w_dff_B_zYDVsHBR5_0),.clk(gclk));
	jdff dff_B_K1QIor8x8_0(.din(w_dff_B_zYDVsHBR5_0),.dout(w_dff_B_K1QIor8x8_0),.clk(gclk));
	jdff dff_B_U6bqcODq5_0(.din(w_dff_B_K1QIor8x8_0),.dout(w_dff_B_U6bqcODq5_0),.clk(gclk));
	jdff dff_B_YD1IGiht4_0(.din(w_dff_B_U6bqcODq5_0),.dout(w_dff_B_YD1IGiht4_0),.clk(gclk));
	jdff dff_B_bCQHAXsL2_0(.din(w_dff_B_YD1IGiht4_0),.dout(w_dff_B_bCQHAXsL2_0),.clk(gclk));
	jdff dff_B_gQ14AX0l4_0(.din(w_dff_B_bCQHAXsL2_0),.dout(w_dff_B_gQ14AX0l4_0),.clk(gclk));
	jdff dff_B_oaSy403U7_0(.din(w_dff_B_gQ14AX0l4_0),.dout(w_dff_B_oaSy403U7_0),.clk(gclk));
	jdff dff_B_d7hK51g43_0(.din(w_dff_B_oaSy403U7_0),.dout(w_dff_B_d7hK51g43_0),.clk(gclk));
	jdff dff_B_eIHhFn8J8_0(.din(w_dff_B_d7hK51g43_0),.dout(w_dff_B_eIHhFn8J8_0),.clk(gclk));
	jdff dff_B_uzwh64ZQ1_0(.din(n628),.dout(w_dff_B_uzwh64ZQ1_0),.clk(gclk));
	jdff dff_B_P26dG0r79_0(.din(w_dff_B_uzwh64ZQ1_0),.dout(w_dff_B_P26dG0r79_0),.clk(gclk));
	jdff dff_B_YrIPbXsZ4_0(.din(w_dff_B_P26dG0r79_0),.dout(w_dff_B_YrIPbXsZ4_0),.clk(gclk));
	jdff dff_B_xp16meGh1_0(.din(w_dff_B_YrIPbXsZ4_0),.dout(w_dff_B_xp16meGh1_0),.clk(gclk));
	jdff dff_B_g0c7eyZI8_0(.din(w_dff_B_xp16meGh1_0),.dout(w_dff_B_g0c7eyZI8_0),.clk(gclk));
	jdff dff_B_lWtXOHqv1_0(.din(w_dff_B_g0c7eyZI8_0),.dout(w_dff_B_lWtXOHqv1_0),.clk(gclk));
	jdff dff_B_a2r6yoBS5_0(.din(w_dff_B_lWtXOHqv1_0),.dout(w_dff_B_a2r6yoBS5_0),.clk(gclk));
	jdff dff_B_0SgxtVVo5_0(.din(w_dff_B_a2r6yoBS5_0),.dout(w_dff_B_0SgxtVVo5_0),.clk(gclk));
	jdff dff_B_4f0Wic170_0(.din(w_dff_B_0SgxtVVo5_0),.dout(w_dff_B_4f0Wic170_0),.clk(gclk));
	jdff dff_B_GZ6Jq6qm9_0(.din(w_dff_B_4f0Wic170_0),.dout(w_dff_B_GZ6Jq6qm9_0),.clk(gclk));
	jdff dff_B_gsRdRIWq7_0(.din(w_dff_B_GZ6Jq6qm9_0),.dout(w_dff_B_gsRdRIWq7_0),.clk(gclk));
	jdff dff_B_XNNavWuD4_0(.din(w_dff_B_gsRdRIWq7_0),.dout(w_dff_B_XNNavWuD4_0),.clk(gclk));
	jdff dff_B_XT8e6qB99_0(.din(w_dff_B_XNNavWuD4_0),.dout(w_dff_B_XT8e6qB99_0),.clk(gclk));
	jdff dff_B_eePq8pFt3_0(.din(w_dff_B_XT8e6qB99_0),.dout(w_dff_B_eePq8pFt3_0),.clk(gclk));
	jdff dff_B_SUABLWS71_0(.din(w_dff_B_eePq8pFt3_0),.dout(w_dff_B_SUABLWS71_0),.clk(gclk));
	jdff dff_B_8BTAbnth5_0(.din(w_dff_B_SUABLWS71_0),.dout(w_dff_B_8BTAbnth5_0),.clk(gclk));
	jdff dff_B_Ut2sz3us0_0(.din(w_dff_B_8BTAbnth5_0),.dout(w_dff_B_Ut2sz3us0_0),.clk(gclk));
	jdff dff_B_Plic3a3j8_0(.din(w_dff_B_Ut2sz3us0_0),.dout(w_dff_B_Plic3a3j8_0),.clk(gclk));
	jdff dff_B_MZEnoUNH3_0(.din(w_dff_B_Plic3a3j8_0),.dout(w_dff_B_MZEnoUNH3_0),.clk(gclk));
	jdff dff_B_DTCGJKIN6_0(.din(w_dff_B_MZEnoUNH3_0),.dout(w_dff_B_DTCGJKIN6_0),.clk(gclk));
	jdff dff_B_K5u2vD9v1_0(.din(w_dff_B_DTCGJKIN6_0),.dout(w_dff_B_K5u2vD9v1_0),.clk(gclk));
	jdff dff_B_g3h6yE2P4_0(.din(w_dff_B_K5u2vD9v1_0),.dout(w_dff_B_g3h6yE2P4_0),.clk(gclk));
	jdff dff_B_sK0uWiil3_0(.din(w_dff_B_g3h6yE2P4_0),.dout(w_dff_B_sK0uWiil3_0),.clk(gclk));
	jdff dff_B_kpCK9AYw5_0(.din(w_dff_B_sK0uWiil3_0),.dout(w_dff_B_kpCK9AYw5_0),.clk(gclk));
	jdff dff_B_fKajguko2_0(.din(w_dff_B_kpCK9AYw5_0),.dout(w_dff_B_fKajguko2_0),.clk(gclk));
	jdff dff_B_JHbXgzf36_0(.din(w_dff_B_fKajguko2_0),.dout(w_dff_B_JHbXgzf36_0),.clk(gclk));
	jdff dff_B_9DzzZAaj7_0(.din(w_dff_B_JHbXgzf36_0),.dout(w_dff_B_9DzzZAaj7_0),.clk(gclk));
	jdff dff_B_WnC1ZTp31_0(.din(w_dff_B_9DzzZAaj7_0),.dout(w_dff_B_WnC1ZTp31_0),.clk(gclk));
	jdff dff_B_NTeej0HV4_0(.din(w_dff_B_WnC1ZTp31_0),.dout(w_dff_B_NTeej0HV4_0),.clk(gclk));
	jdff dff_B_OoHRG8iE5_0(.din(w_dff_B_NTeej0HV4_0),.dout(w_dff_B_OoHRG8iE5_0),.clk(gclk));
	jdff dff_B_fwQc2M8m5_0(.din(w_dff_B_OoHRG8iE5_0),.dout(w_dff_B_fwQc2M8m5_0),.clk(gclk));
	jdff dff_B_NKGDZyvl6_0(.din(w_dff_B_fwQc2M8m5_0),.dout(w_dff_B_NKGDZyvl6_0),.clk(gclk));
	jdff dff_B_7j9CpVE68_0(.din(w_dff_B_NKGDZyvl6_0),.dout(w_dff_B_7j9CpVE68_0),.clk(gclk));
	jdff dff_B_f9MTalO10_0(.din(w_dff_B_7j9CpVE68_0),.dout(w_dff_B_f9MTalO10_0),.clk(gclk));
	jdff dff_B_bdZ8XQ5Z6_0(.din(w_dff_B_f9MTalO10_0),.dout(w_dff_B_bdZ8XQ5Z6_0),.clk(gclk));
	jdff dff_B_5Y14gjS09_0(.din(w_dff_B_bdZ8XQ5Z6_0),.dout(w_dff_B_5Y14gjS09_0),.clk(gclk));
	jdff dff_B_6Hws304o8_0(.din(w_dff_B_5Y14gjS09_0),.dout(w_dff_B_6Hws304o8_0),.clk(gclk));
	jdff dff_B_Y0kU99sb4_0(.din(w_dff_B_6Hws304o8_0),.dout(w_dff_B_Y0kU99sb4_0),.clk(gclk));
	jdff dff_B_MCBIitm02_0(.din(w_dff_B_Y0kU99sb4_0),.dout(w_dff_B_MCBIitm02_0),.clk(gclk));
	jdff dff_B_HBMFIay39_0(.din(w_dff_B_MCBIitm02_0),.dout(w_dff_B_HBMFIay39_0),.clk(gclk));
	jdff dff_B_0shDgtgi6_0(.din(n634),.dout(w_dff_B_0shDgtgi6_0),.clk(gclk));
	jdff dff_B_OwZF7A2q1_0(.din(w_dff_B_0shDgtgi6_0),.dout(w_dff_B_OwZF7A2q1_0),.clk(gclk));
	jdff dff_B_Njp67Q9q1_0(.din(w_dff_B_OwZF7A2q1_0),.dout(w_dff_B_Njp67Q9q1_0),.clk(gclk));
	jdff dff_B_knggDeZI2_0(.din(w_dff_B_Njp67Q9q1_0),.dout(w_dff_B_knggDeZI2_0),.clk(gclk));
	jdff dff_B_bijPdv523_0(.din(w_dff_B_knggDeZI2_0),.dout(w_dff_B_bijPdv523_0),.clk(gclk));
	jdff dff_B_lM6JNNjH4_0(.din(w_dff_B_bijPdv523_0),.dout(w_dff_B_lM6JNNjH4_0),.clk(gclk));
	jdff dff_B_2zNi7IL35_0(.din(w_dff_B_lM6JNNjH4_0),.dout(w_dff_B_2zNi7IL35_0),.clk(gclk));
	jdff dff_B_scuPywgt9_0(.din(w_dff_B_2zNi7IL35_0),.dout(w_dff_B_scuPywgt9_0),.clk(gclk));
	jdff dff_B_hIgJRwBa4_0(.din(w_dff_B_scuPywgt9_0),.dout(w_dff_B_hIgJRwBa4_0),.clk(gclk));
	jdff dff_B_h2i7UkD71_0(.din(w_dff_B_hIgJRwBa4_0),.dout(w_dff_B_h2i7UkD71_0),.clk(gclk));
	jdff dff_B_FhvbVRyo4_0(.din(w_dff_B_h2i7UkD71_0),.dout(w_dff_B_FhvbVRyo4_0),.clk(gclk));
	jdff dff_B_XHuxvklI3_0(.din(w_dff_B_FhvbVRyo4_0),.dout(w_dff_B_XHuxvklI3_0),.clk(gclk));
	jdff dff_B_G0qV8B3v2_0(.din(w_dff_B_XHuxvklI3_0),.dout(w_dff_B_G0qV8B3v2_0),.clk(gclk));
	jdff dff_B_5cLs7z8c3_0(.din(w_dff_B_G0qV8B3v2_0),.dout(w_dff_B_5cLs7z8c3_0),.clk(gclk));
	jdff dff_B_NtOV4SLt6_0(.din(w_dff_B_5cLs7z8c3_0),.dout(w_dff_B_NtOV4SLt6_0),.clk(gclk));
	jdff dff_B_uryy4H9k8_0(.din(w_dff_B_NtOV4SLt6_0),.dout(w_dff_B_uryy4H9k8_0),.clk(gclk));
	jdff dff_B_Au9BNQV14_0(.din(w_dff_B_uryy4H9k8_0),.dout(w_dff_B_Au9BNQV14_0),.clk(gclk));
	jdff dff_B_WfQJyuZA1_0(.din(w_dff_B_Au9BNQV14_0),.dout(w_dff_B_WfQJyuZA1_0),.clk(gclk));
	jdff dff_B_jzsr3Afh1_0(.din(w_dff_B_WfQJyuZA1_0),.dout(w_dff_B_jzsr3Afh1_0),.clk(gclk));
	jdff dff_B_xwakBVa87_0(.din(w_dff_B_jzsr3Afh1_0),.dout(w_dff_B_xwakBVa87_0),.clk(gclk));
	jdff dff_B_8FeW9SoK2_0(.din(w_dff_B_xwakBVa87_0),.dout(w_dff_B_8FeW9SoK2_0),.clk(gclk));
	jdff dff_B_BOjsym2A9_0(.din(w_dff_B_8FeW9SoK2_0),.dout(w_dff_B_BOjsym2A9_0),.clk(gclk));
	jdff dff_B_HcHVv9Zk6_0(.din(w_dff_B_BOjsym2A9_0),.dout(w_dff_B_HcHVv9Zk6_0),.clk(gclk));
	jdff dff_B_sRlJnjoU3_0(.din(w_dff_B_HcHVv9Zk6_0),.dout(w_dff_B_sRlJnjoU3_0),.clk(gclk));
	jdff dff_B_dARBkwhE0_0(.din(w_dff_B_sRlJnjoU3_0),.dout(w_dff_B_dARBkwhE0_0),.clk(gclk));
	jdff dff_B_u092cIuI7_0(.din(w_dff_B_dARBkwhE0_0),.dout(w_dff_B_u092cIuI7_0),.clk(gclk));
	jdff dff_B_WznS65yE5_0(.din(w_dff_B_u092cIuI7_0),.dout(w_dff_B_WznS65yE5_0),.clk(gclk));
	jdff dff_B_K1bWBl5p3_0(.din(w_dff_B_WznS65yE5_0),.dout(w_dff_B_K1bWBl5p3_0),.clk(gclk));
	jdff dff_B_kw6iMMN12_0(.din(w_dff_B_K1bWBl5p3_0),.dout(w_dff_B_kw6iMMN12_0),.clk(gclk));
	jdff dff_B_dZxlWiiz8_0(.din(w_dff_B_kw6iMMN12_0),.dout(w_dff_B_dZxlWiiz8_0),.clk(gclk));
	jdff dff_B_Gq1zhtW23_0(.din(w_dff_B_dZxlWiiz8_0),.dout(w_dff_B_Gq1zhtW23_0),.clk(gclk));
	jdff dff_B_2dhpKj3Z5_0(.din(w_dff_B_Gq1zhtW23_0),.dout(w_dff_B_2dhpKj3Z5_0),.clk(gclk));
	jdff dff_B_YN02L5Tb2_0(.din(w_dff_B_2dhpKj3Z5_0),.dout(w_dff_B_YN02L5Tb2_0),.clk(gclk));
	jdff dff_B_nLXJy6dc4_0(.din(w_dff_B_YN02L5Tb2_0),.dout(w_dff_B_nLXJy6dc4_0),.clk(gclk));
	jdff dff_B_UNEo6wsu4_0(.din(w_dff_B_nLXJy6dc4_0),.dout(w_dff_B_UNEo6wsu4_0),.clk(gclk));
	jdff dff_B_tdOr23mj8_0(.din(w_dff_B_UNEo6wsu4_0),.dout(w_dff_B_tdOr23mj8_0),.clk(gclk));
	jdff dff_B_4KUK3YVo4_0(.din(w_dff_B_tdOr23mj8_0),.dout(w_dff_B_4KUK3YVo4_0),.clk(gclk));
	jdff dff_B_WPrisq2B5_0(.din(w_dff_B_4KUK3YVo4_0),.dout(w_dff_B_WPrisq2B5_0),.clk(gclk));
	jdff dff_B_uohnTt1u7_0(.din(w_dff_B_WPrisq2B5_0),.dout(w_dff_B_uohnTt1u7_0),.clk(gclk));
	jdff dff_B_bPNl0kxX2_0(.din(w_dff_B_uohnTt1u7_0),.dout(w_dff_B_bPNl0kxX2_0),.clk(gclk));
	jdff dff_B_UJ4VqMGy1_0(.din(w_dff_B_bPNl0kxX2_0),.dout(w_dff_B_UJ4VqMGy1_0),.clk(gclk));
	jdff dff_B_Dw9LvKPt7_0(.din(n640),.dout(w_dff_B_Dw9LvKPt7_0),.clk(gclk));
	jdff dff_B_F3HgZvHC3_0(.din(w_dff_B_Dw9LvKPt7_0),.dout(w_dff_B_F3HgZvHC3_0),.clk(gclk));
	jdff dff_B_vpUc6sWw9_0(.din(w_dff_B_F3HgZvHC3_0),.dout(w_dff_B_vpUc6sWw9_0),.clk(gclk));
	jdff dff_B_MVoAxxd25_0(.din(w_dff_B_vpUc6sWw9_0),.dout(w_dff_B_MVoAxxd25_0),.clk(gclk));
	jdff dff_B_bG5EeO7j0_0(.din(w_dff_B_MVoAxxd25_0),.dout(w_dff_B_bG5EeO7j0_0),.clk(gclk));
	jdff dff_B_our3pX4s3_0(.din(w_dff_B_bG5EeO7j0_0),.dout(w_dff_B_our3pX4s3_0),.clk(gclk));
	jdff dff_B_SkbhW8q33_0(.din(w_dff_B_our3pX4s3_0),.dout(w_dff_B_SkbhW8q33_0),.clk(gclk));
	jdff dff_B_LBl5ZMZc8_0(.din(w_dff_B_SkbhW8q33_0),.dout(w_dff_B_LBl5ZMZc8_0),.clk(gclk));
	jdff dff_B_DFK2HWJM3_0(.din(w_dff_B_LBl5ZMZc8_0),.dout(w_dff_B_DFK2HWJM3_0),.clk(gclk));
	jdff dff_B_zoLJ1wL50_0(.din(w_dff_B_DFK2HWJM3_0),.dout(w_dff_B_zoLJ1wL50_0),.clk(gclk));
	jdff dff_B_uFCg0IJZ0_0(.din(w_dff_B_zoLJ1wL50_0),.dout(w_dff_B_uFCg0IJZ0_0),.clk(gclk));
	jdff dff_B_aQlz3YYd5_0(.din(w_dff_B_uFCg0IJZ0_0),.dout(w_dff_B_aQlz3YYd5_0),.clk(gclk));
	jdff dff_B_SlYUAo0z9_0(.din(w_dff_B_aQlz3YYd5_0),.dout(w_dff_B_SlYUAo0z9_0),.clk(gclk));
	jdff dff_B_sBBes0xc8_0(.din(w_dff_B_SlYUAo0z9_0),.dout(w_dff_B_sBBes0xc8_0),.clk(gclk));
	jdff dff_B_5njRckK90_0(.din(w_dff_B_sBBes0xc8_0),.dout(w_dff_B_5njRckK90_0),.clk(gclk));
	jdff dff_B_85bgcXBo0_0(.din(w_dff_B_5njRckK90_0),.dout(w_dff_B_85bgcXBo0_0),.clk(gclk));
	jdff dff_B_XNJW62EU4_0(.din(w_dff_B_85bgcXBo0_0),.dout(w_dff_B_XNJW62EU4_0),.clk(gclk));
	jdff dff_B_rkaCF3Ll7_0(.din(w_dff_B_XNJW62EU4_0),.dout(w_dff_B_rkaCF3Ll7_0),.clk(gclk));
	jdff dff_B_O8h5cX5Y5_0(.din(w_dff_B_rkaCF3Ll7_0),.dout(w_dff_B_O8h5cX5Y5_0),.clk(gclk));
	jdff dff_B_n87STnP53_0(.din(w_dff_B_O8h5cX5Y5_0),.dout(w_dff_B_n87STnP53_0),.clk(gclk));
	jdff dff_B_aoEp5HyJ1_0(.din(w_dff_B_n87STnP53_0),.dout(w_dff_B_aoEp5HyJ1_0),.clk(gclk));
	jdff dff_B_vkl8CucJ7_0(.din(w_dff_B_aoEp5HyJ1_0),.dout(w_dff_B_vkl8CucJ7_0),.clk(gclk));
	jdff dff_B_XSXQ0ndg2_0(.din(w_dff_B_vkl8CucJ7_0),.dout(w_dff_B_XSXQ0ndg2_0),.clk(gclk));
	jdff dff_B_qOfmuQz04_0(.din(w_dff_B_XSXQ0ndg2_0),.dout(w_dff_B_qOfmuQz04_0),.clk(gclk));
	jdff dff_B_B6IwPksD0_0(.din(w_dff_B_qOfmuQz04_0),.dout(w_dff_B_B6IwPksD0_0),.clk(gclk));
	jdff dff_B_uYunf61j5_0(.din(w_dff_B_B6IwPksD0_0),.dout(w_dff_B_uYunf61j5_0),.clk(gclk));
	jdff dff_B_ZMSEquwr8_0(.din(w_dff_B_uYunf61j5_0),.dout(w_dff_B_ZMSEquwr8_0),.clk(gclk));
	jdff dff_B_IMqFlEtW8_0(.din(w_dff_B_ZMSEquwr8_0),.dout(w_dff_B_IMqFlEtW8_0),.clk(gclk));
	jdff dff_B_fgI9Qkzi7_0(.din(w_dff_B_IMqFlEtW8_0),.dout(w_dff_B_fgI9Qkzi7_0),.clk(gclk));
	jdff dff_B_RFb61G1o8_0(.din(w_dff_B_fgI9Qkzi7_0),.dout(w_dff_B_RFb61G1o8_0),.clk(gclk));
	jdff dff_B_GTjikBJ02_0(.din(w_dff_B_RFb61G1o8_0),.dout(w_dff_B_GTjikBJ02_0),.clk(gclk));
	jdff dff_B_k8qXUAkW5_0(.din(w_dff_B_GTjikBJ02_0),.dout(w_dff_B_k8qXUAkW5_0),.clk(gclk));
	jdff dff_B_oI172RwO8_0(.din(w_dff_B_k8qXUAkW5_0),.dout(w_dff_B_oI172RwO8_0),.clk(gclk));
	jdff dff_B_rRnvMP1O8_0(.din(w_dff_B_oI172RwO8_0),.dout(w_dff_B_rRnvMP1O8_0),.clk(gclk));
	jdff dff_B_T255YwsT7_0(.din(w_dff_B_rRnvMP1O8_0),.dout(w_dff_B_T255YwsT7_0),.clk(gclk));
	jdff dff_B_42m6RJiu9_0(.din(w_dff_B_T255YwsT7_0),.dout(w_dff_B_42m6RJiu9_0),.clk(gclk));
	jdff dff_B_3xcDFFQS6_0(.din(w_dff_B_42m6RJiu9_0),.dout(w_dff_B_3xcDFFQS6_0),.clk(gclk));
	jdff dff_B_11p6Jy1p3_0(.din(w_dff_B_3xcDFFQS6_0),.dout(w_dff_B_11p6Jy1p3_0),.clk(gclk));
	jdff dff_B_WgaVymgg2_0(.din(w_dff_B_11p6Jy1p3_0),.dout(w_dff_B_WgaVymgg2_0),.clk(gclk));
	jdff dff_B_rULrk60d0_0(.din(w_dff_B_WgaVymgg2_0),.dout(w_dff_B_rULrk60d0_0),.clk(gclk));
	jdff dff_B_e5I5U3Sn2_0(.din(w_dff_B_rULrk60d0_0),.dout(w_dff_B_e5I5U3Sn2_0),.clk(gclk));
	jdff dff_B_t6QLfecs2_0(.din(w_dff_B_e5I5U3Sn2_0),.dout(w_dff_B_t6QLfecs2_0),.clk(gclk));
	jdff dff_B_ipxo879F6_0(.din(n646),.dout(w_dff_B_ipxo879F6_0),.clk(gclk));
	jdff dff_B_LSskEnMJ6_0(.din(w_dff_B_ipxo879F6_0),.dout(w_dff_B_LSskEnMJ6_0),.clk(gclk));
	jdff dff_B_kSarhR290_0(.din(w_dff_B_LSskEnMJ6_0),.dout(w_dff_B_kSarhR290_0),.clk(gclk));
	jdff dff_B_qwn9lQy21_0(.din(w_dff_B_kSarhR290_0),.dout(w_dff_B_qwn9lQy21_0),.clk(gclk));
	jdff dff_B_WKGrDndw1_0(.din(w_dff_B_qwn9lQy21_0),.dout(w_dff_B_WKGrDndw1_0),.clk(gclk));
	jdff dff_B_afJdtZAd7_0(.din(w_dff_B_WKGrDndw1_0),.dout(w_dff_B_afJdtZAd7_0),.clk(gclk));
	jdff dff_B_nNZZktFn6_0(.din(w_dff_B_afJdtZAd7_0),.dout(w_dff_B_nNZZktFn6_0),.clk(gclk));
	jdff dff_B_7MkIh2KA8_0(.din(w_dff_B_nNZZktFn6_0),.dout(w_dff_B_7MkIh2KA8_0),.clk(gclk));
	jdff dff_B_2yQ49Zkb6_0(.din(w_dff_B_7MkIh2KA8_0),.dout(w_dff_B_2yQ49Zkb6_0),.clk(gclk));
	jdff dff_B_cHmaKI156_0(.din(w_dff_B_2yQ49Zkb6_0),.dout(w_dff_B_cHmaKI156_0),.clk(gclk));
	jdff dff_B_g6wJIYSG6_0(.din(w_dff_B_cHmaKI156_0),.dout(w_dff_B_g6wJIYSG6_0),.clk(gclk));
	jdff dff_B_8QVHYHU94_0(.din(w_dff_B_g6wJIYSG6_0),.dout(w_dff_B_8QVHYHU94_0),.clk(gclk));
	jdff dff_B_OLFhO0Yd9_0(.din(w_dff_B_8QVHYHU94_0),.dout(w_dff_B_OLFhO0Yd9_0),.clk(gclk));
	jdff dff_B_PxB1hz0Q4_0(.din(w_dff_B_OLFhO0Yd9_0),.dout(w_dff_B_PxB1hz0Q4_0),.clk(gclk));
	jdff dff_B_oXVIDWno3_0(.din(w_dff_B_PxB1hz0Q4_0),.dout(w_dff_B_oXVIDWno3_0),.clk(gclk));
	jdff dff_B_PTTpeujz5_0(.din(w_dff_B_oXVIDWno3_0),.dout(w_dff_B_PTTpeujz5_0),.clk(gclk));
	jdff dff_B_Gwt3tcAo9_0(.din(w_dff_B_PTTpeujz5_0),.dout(w_dff_B_Gwt3tcAo9_0),.clk(gclk));
	jdff dff_B_GtQzg2ep8_0(.din(w_dff_B_Gwt3tcAo9_0),.dout(w_dff_B_GtQzg2ep8_0),.clk(gclk));
	jdff dff_B_2n3G3H5L4_0(.din(w_dff_B_GtQzg2ep8_0),.dout(w_dff_B_2n3G3H5L4_0),.clk(gclk));
	jdff dff_B_tsECu0FY7_0(.din(w_dff_B_2n3G3H5L4_0),.dout(w_dff_B_tsECu0FY7_0),.clk(gclk));
	jdff dff_B_VMRiwwx70_0(.din(w_dff_B_tsECu0FY7_0),.dout(w_dff_B_VMRiwwx70_0),.clk(gclk));
	jdff dff_B_XS0631CG3_0(.din(w_dff_B_VMRiwwx70_0),.dout(w_dff_B_XS0631CG3_0),.clk(gclk));
	jdff dff_B_CCSelazc3_0(.din(w_dff_B_XS0631CG3_0),.dout(w_dff_B_CCSelazc3_0),.clk(gclk));
	jdff dff_B_Bsluvwhw1_0(.din(w_dff_B_CCSelazc3_0),.dout(w_dff_B_Bsluvwhw1_0),.clk(gclk));
	jdff dff_B_51VFRWtS5_0(.din(w_dff_B_Bsluvwhw1_0),.dout(w_dff_B_51VFRWtS5_0),.clk(gclk));
	jdff dff_B_mTeLjdGv6_0(.din(w_dff_B_51VFRWtS5_0),.dout(w_dff_B_mTeLjdGv6_0),.clk(gclk));
	jdff dff_B_yGur854F1_0(.din(w_dff_B_mTeLjdGv6_0),.dout(w_dff_B_yGur854F1_0),.clk(gclk));
	jdff dff_B_QUUjOG627_0(.din(w_dff_B_yGur854F1_0),.dout(w_dff_B_QUUjOG627_0),.clk(gclk));
	jdff dff_B_yoDLszcW6_0(.din(w_dff_B_QUUjOG627_0),.dout(w_dff_B_yoDLszcW6_0),.clk(gclk));
	jdff dff_B_VIG8Z6DN4_0(.din(w_dff_B_yoDLszcW6_0),.dout(w_dff_B_VIG8Z6DN4_0),.clk(gclk));
	jdff dff_B_QJdXGEHe1_0(.din(w_dff_B_VIG8Z6DN4_0),.dout(w_dff_B_QJdXGEHe1_0),.clk(gclk));
	jdff dff_B_N4Bt5eBE8_0(.din(w_dff_B_QJdXGEHe1_0),.dout(w_dff_B_N4Bt5eBE8_0),.clk(gclk));
	jdff dff_B_e92iYarn4_0(.din(w_dff_B_N4Bt5eBE8_0),.dout(w_dff_B_e92iYarn4_0),.clk(gclk));
	jdff dff_B_X76LfSTG3_0(.din(w_dff_B_e92iYarn4_0),.dout(w_dff_B_X76LfSTG3_0),.clk(gclk));
	jdff dff_B_2xSQeiu16_0(.din(w_dff_B_X76LfSTG3_0),.dout(w_dff_B_2xSQeiu16_0),.clk(gclk));
	jdff dff_B_qvtBlUWO1_0(.din(w_dff_B_2xSQeiu16_0),.dout(w_dff_B_qvtBlUWO1_0),.clk(gclk));
	jdff dff_B_YYkGdOSP9_0(.din(w_dff_B_qvtBlUWO1_0),.dout(w_dff_B_YYkGdOSP9_0),.clk(gclk));
	jdff dff_B_j3debmty7_0(.din(w_dff_B_YYkGdOSP9_0),.dout(w_dff_B_j3debmty7_0),.clk(gclk));
	jdff dff_B_xs3cG4LX2_0(.din(w_dff_B_j3debmty7_0),.dout(w_dff_B_xs3cG4LX2_0),.clk(gclk));
	jdff dff_B_x65iNM1F9_0(.din(w_dff_B_xs3cG4LX2_0),.dout(w_dff_B_x65iNM1F9_0),.clk(gclk));
	jdff dff_B_EYuBOgii4_0(.din(w_dff_B_x65iNM1F9_0),.dout(w_dff_B_EYuBOgii4_0),.clk(gclk));
	jdff dff_B_wI3Cf3A44_0(.din(w_dff_B_EYuBOgii4_0),.dout(w_dff_B_wI3Cf3A44_0),.clk(gclk));
	jdff dff_B_2nixnkQN6_0(.din(w_dff_B_wI3Cf3A44_0),.dout(w_dff_B_2nixnkQN6_0),.clk(gclk));
	jdff dff_B_tGL8PZ947_0(.din(n652),.dout(w_dff_B_tGL8PZ947_0),.clk(gclk));
	jdff dff_B_Xu7bofGJ3_0(.din(w_dff_B_tGL8PZ947_0),.dout(w_dff_B_Xu7bofGJ3_0),.clk(gclk));
	jdff dff_B_k1reFg2Z8_0(.din(w_dff_B_Xu7bofGJ3_0),.dout(w_dff_B_k1reFg2Z8_0),.clk(gclk));
	jdff dff_B_wmCn36vi4_0(.din(w_dff_B_k1reFg2Z8_0),.dout(w_dff_B_wmCn36vi4_0),.clk(gclk));
	jdff dff_B_tqXKCHTo3_0(.din(w_dff_B_wmCn36vi4_0),.dout(w_dff_B_tqXKCHTo3_0),.clk(gclk));
	jdff dff_B_cIz092fC1_0(.din(w_dff_B_tqXKCHTo3_0),.dout(w_dff_B_cIz092fC1_0),.clk(gclk));
	jdff dff_B_Yb4ag7pK5_0(.din(w_dff_B_cIz092fC1_0),.dout(w_dff_B_Yb4ag7pK5_0),.clk(gclk));
	jdff dff_B_IGfYsjbi7_0(.din(w_dff_B_Yb4ag7pK5_0),.dout(w_dff_B_IGfYsjbi7_0),.clk(gclk));
	jdff dff_B_I9vqk8f01_0(.din(w_dff_B_IGfYsjbi7_0),.dout(w_dff_B_I9vqk8f01_0),.clk(gclk));
	jdff dff_B_ZZ7QeuFW7_0(.din(w_dff_B_I9vqk8f01_0),.dout(w_dff_B_ZZ7QeuFW7_0),.clk(gclk));
	jdff dff_B_RzKjdOXz7_0(.din(w_dff_B_ZZ7QeuFW7_0),.dout(w_dff_B_RzKjdOXz7_0),.clk(gclk));
	jdff dff_B_OTKGhE4w8_0(.din(w_dff_B_RzKjdOXz7_0),.dout(w_dff_B_OTKGhE4w8_0),.clk(gclk));
	jdff dff_B_2NqZLi6Q9_0(.din(w_dff_B_OTKGhE4w8_0),.dout(w_dff_B_2NqZLi6Q9_0),.clk(gclk));
	jdff dff_B_tWOAFbuI2_0(.din(w_dff_B_2NqZLi6Q9_0),.dout(w_dff_B_tWOAFbuI2_0),.clk(gclk));
	jdff dff_B_pmOHpTZh9_0(.din(w_dff_B_tWOAFbuI2_0),.dout(w_dff_B_pmOHpTZh9_0),.clk(gclk));
	jdff dff_B_VYgOSosZ4_0(.din(w_dff_B_pmOHpTZh9_0),.dout(w_dff_B_VYgOSosZ4_0),.clk(gclk));
	jdff dff_B_OcWz94yU5_0(.din(w_dff_B_VYgOSosZ4_0),.dout(w_dff_B_OcWz94yU5_0),.clk(gclk));
	jdff dff_B_wfURwYwy5_0(.din(w_dff_B_OcWz94yU5_0),.dout(w_dff_B_wfURwYwy5_0),.clk(gclk));
	jdff dff_B_UEbPj2ex0_0(.din(w_dff_B_wfURwYwy5_0),.dout(w_dff_B_UEbPj2ex0_0),.clk(gclk));
	jdff dff_B_7qf3MIVd5_0(.din(w_dff_B_UEbPj2ex0_0),.dout(w_dff_B_7qf3MIVd5_0),.clk(gclk));
	jdff dff_B_ZhpquE2L4_0(.din(w_dff_B_7qf3MIVd5_0),.dout(w_dff_B_ZhpquE2L4_0),.clk(gclk));
	jdff dff_B_Z1sEhCcS4_0(.din(w_dff_B_ZhpquE2L4_0),.dout(w_dff_B_Z1sEhCcS4_0),.clk(gclk));
	jdff dff_B_aEU3q0Pn6_0(.din(w_dff_B_Z1sEhCcS4_0),.dout(w_dff_B_aEU3q0Pn6_0),.clk(gclk));
	jdff dff_B_49y7Vyes8_0(.din(w_dff_B_aEU3q0Pn6_0),.dout(w_dff_B_49y7Vyes8_0),.clk(gclk));
	jdff dff_B_7UwlhvjH8_0(.din(w_dff_B_49y7Vyes8_0),.dout(w_dff_B_7UwlhvjH8_0),.clk(gclk));
	jdff dff_B_L8kWT1sg0_0(.din(w_dff_B_7UwlhvjH8_0),.dout(w_dff_B_L8kWT1sg0_0),.clk(gclk));
	jdff dff_B_XIehFfsR7_0(.din(w_dff_B_L8kWT1sg0_0),.dout(w_dff_B_XIehFfsR7_0),.clk(gclk));
	jdff dff_B_3dWOH05e9_0(.din(w_dff_B_XIehFfsR7_0),.dout(w_dff_B_3dWOH05e9_0),.clk(gclk));
	jdff dff_B_p1G72ESf6_0(.din(w_dff_B_3dWOH05e9_0),.dout(w_dff_B_p1G72ESf6_0),.clk(gclk));
	jdff dff_B_1dMPIVHc7_0(.din(w_dff_B_p1G72ESf6_0),.dout(w_dff_B_1dMPIVHc7_0),.clk(gclk));
	jdff dff_B_mgpiqFS94_0(.din(w_dff_B_1dMPIVHc7_0),.dout(w_dff_B_mgpiqFS94_0),.clk(gclk));
	jdff dff_B_BIcdm2cr2_0(.din(w_dff_B_mgpiqFS94_0),.dout(w_dff_B_BIcdm2cr2_0),.clk(gclk));
	jdff dff_B_M94wlmKC3_0(.din(w_dff_B_BIcdm2cr2_0),.dout(w_dff_B_M94wlmKC3_0),.clk(gclk));
	jdff dff_B_vcvzEnob7_0(.din(w_dff_B_M94wlmKC3_0),.dout(w_dff_B_vcvzEnob7_0),.clk(gclk));
	jdff dff_B_JORzm03B9_0(.din(w_dff_B_vcvzEnob7_0),.dout(w_dff_B_JORzm03B9_0),.clk(gclk));
	jdff dff_B_WDjfKekK6_0(.din(w_dff_B_JORzm03B9_0),.dout(w_dff_B_WDjfKekK6_0),.clk(gclk));
	jdff dff_B_H3rIGwZJ9_0(.din(w_dff_B_WDjfKekK6_0),.dout(w_dff_B_H3rIGwZJ9_0),.clk(gclk));
	jdff dff_B_PataCVEL7_0(.din(w_dff_B_H3rIGwZJ9_0),.dout(w_dff_B_PataCVEL7_0),.clk(gclk));
	jdff dff_B_rmNAAghH0_0(.din(w_dff_B_PataCVEL7_0),.dout(w_dff_B_rmNAAghH0_0),.clk(gclk));
	jdff dff_B_Xyt7SfeP9_0(.din(w_dff_B_rmNAAghH0_0),.dout(w_dff_B_Xyt7SfeP9_0),.clk(gclk));
	jdff dff_B_RW7QdTNT6_0(.din(w_dff_B_Xyt7SfeP9_0),.dout(w_dff_B_RW7QdTNT6_0),.clk(gclk));
	jdff dff_B_NOPjgN8E1_0(.din(w_dff_B_RW7QdTNT6_0),.dout(w_dff_B_NOPjgN8E1_0),.clk(gclk));
	jdff dff_B_t1FPDMuA6_0(.din(w_dff_B_NOPjgN8E1_0),.dout(w_dff_B_t1FPDMuA6_0),.clk(gclk));
	jdff dff_B_9PsGZFcP4_0(.din(w_dff_B_t1FPDMuA6_0),.dout(w_dff_B_9PsGZFcP4_0),.clk(gclk));
	jdff dff_B_trwb5HFP2_0(.din(n658),.dout(w_dff_B_trwb5HFP2_0),.clk(gclk));
	jdff dff_B_MH85wwDq2_0(.din(w_dff_B_trwb5HFP2_0),.dout(w_dff_B_MH85wwDq2_0),.clk(gclk));
	jdff dff_B_TD8lqoHM9_0(.din(w_dff_B_MH85wwDq2_0),.dout(w_dff_B_TD8lqoHM9_0),.clk(gclk));
	jdff dff_B_0zq07tCv1_0(.din(w_dff_B_TD8lqoHM9_0),.dout(w_dff_B_0zq07tCv1_0),.clk(gclk));
	jdff dff_B_W8iGleAw0_0(.din(w_dff_B_0zq07tCv1_0),.dout(w_dff_B_W8iGleAw0_0),.clk(gclk));
	jdff dff_B_nEqsQrBN6_0(.din(w_dff_B_W8iGleAw0_0),.dout(w_dff_B_nEqsQrBN6_0),.clk(gclk));
	jdff dff_B_pMmiKsav7_0(.din(w_dff_B_nEqsQrBN6_0),.dout(w_dff_B_pMmiKsav7_0),.clk(gclk));
	jdff dff_B_SAq6hZza6_0(.din(w_dff_B_pMmiKsav7_0),.dout(w_dff_B_SAq6hZza6_0),.clk(gclk));
	jdff dff_B_jPIPrOSc4_0(.din(w_dff_B_SAq6hZza6_0),.dout(w_dff_B_jPIPrOSc4_0),.clk(gclk));
	jdff dff_B_6ylCveDh5_0(.din(w_dff_B_jPIPrOSc4_0),.dout(w_dff_B_6ylCveDh5_0),.clk(gclk));
	jdff dff_B_PvWvV6dw4_0(.din(w_dff_B_6ylCveDh5_0),.dout(w_dff_B_PvWvV6dw4_0),.clk(gclk));
	jdff dff_B_TW2IQEPV5_0(.din(w_dff_B_PvWvV6dw4_0),.dout(w_dff_B_TW2IQEPV5_0),.clk(gclk));
	jdff dff_B_2QnUiGPM2_0(.din(w_dff_B_TW2IQEPV5_0),.dout(w_dff_B_2QnUiGPM2_0),.clk(gclk));
	jdff dff_B_W99afnE09_0(.din(w_dff_B_2QnUiGPM2_0),.dout(w_dff_B_W99afnE09_0),.clk(gclk));
	jdff dff_B_vzjDST0P9_0(.din(w_dff_B_W99afnE09_0),.dout(w_dff_B_vzjDST0P9_0),.clk(gclk));
	jdff dff_B_4O0hpM4s0_0(.din(w_dff_B_vzjDST0P9_0),.dout(w_dff_B_4O0hpM4s0_0),.clk(gclk));
	jdff dff_B_8xvFy2Pr7_0(.din(w_dff_B_4O0hpM4s0_0),.dout(w_dff_B_8xvFy2Pr7_0),.clk(gclk));
	jdff dff_B_thDQF12t1_0(.din(w_dff_B_8xvFy2Pr7_0),.dout(w_dff_B_thDQF12t1_0),.clk(gclk));
	jdff dff_B_wyMx9J7E2_0(.din(w_dff_B_thDQF12t1_0),.dout(w_dff_B_wyMx9J7E2_0),.clk(gclk));
	jdff dff_B_0kiQmwvd1_0(.din(w_dff_B_wyMx9J7E2_0),.dout(w_dff_B_0kiQmwvd1_0),.clk(gclk));
	jdff dff_B_Dpdunlgl8_0(.din(w_dff_B_0kiQmwvd1_0),.dout(w_dff_B_Dpdunlgl8_0),.clk(gclk));
	jdff dff_B_aZ0XF59r1_0(.din(w_dff_B_Dpdunlgl8_0),.dout(w_dff_B_aZ0XF59r1_0),.clk(gclk));
	jdff dff_B_iHqJpSWI3_0(.din(w_dff_B_aZ0XF59r1_0),.dout(w_dff_B_iHqJpSWI3_0),.clk(gclk));
	jdff dff_B_LO75H4Yn5_0(.din(w_dff_B_iHqJpSWI3_0),.dout(w_dff_B_LO75H4Yn5_0),.clk(gclk));
	jdff dff_B_x8z13wvt3_0(.din(w_dff_B_LO75H4Yn5_0),.dout(w_dff_B_x8z13wvt3_0),.clk(gclk));
	jdff dff_B_hFi1hj1w5_0(.din(w_dff_B_x8z13wvt3_0),.dout(w_dff_B_hFi1hj1w5_0),.clk(gclk));
	jdff dff_B_0QbxvLYk6_0(.din(w_dff_B_hFi1hj1w5_0),.dout(w_dff_B_0QbxvLYk6_0),.clk(gclk));
	jdff dff_B_Kpd8xOg80_0(.din(w_dff_B_0QbxvLYk6_0),.dout(w_dff_B_Kpd8xOg80_0),.clk(gclk));
	jdff dff_B_7pGZFqR42_0(.din(w_dff_B_Kpd8xOg80_0),.dout(w_dff_B_7pGZFqR42_0),.clk(gclk));
	jdff dff_B_BoQxKRqO8_0(.din(w_dff_B_7pGZFqR42_0),.dout(w_dff_B_BoQxKRqO8_0),.clk(gclk));
	jdff dff_B_nPhg2Y2v2_0(.din(w_dff_B_BoQxKRqO8_0),.dout(w_dff_B_nPhg2Y2v2_0),.clk(gclk));
	jdff dff_B_WOwpDwsM4_0(.din(w_dff_B_nPhg2Y2v2_0),.dout(w_dff_B_WOwpDwsM4_0),.clk(gclk));
	jdff dff_B_dTK5UeDT8_0(.din(w_dff_B_WOwpDwsM4_0),.dout(w_dff_B_dTK5UeDT8_0),.clk(gclk));
	jdff dff_B_Ta56FccG7_0(.din(w_dff_B_dTK5UeDT8_0),.dout(w_dff_B_Ta56FccG7_0),.clk(gclk));
	jdff dff_B_JU7qH4C10_0(.din(w_dff_B_Ta56FccG7_0),.dout(w_dff_B_JU7qH4C10_0),.clk(gclk));
	jdff dff_B_kB4Q5G4N0_0(.din(w_dff_B_JU7qH4C10_0),.dout(w_dff_B_kB4Q5G4N0_0),.clk(gclk));
	jdff dff_B_bcYDuvh83_0(.din(w_dff_B_kB4Q5G4N0_0),.dout(w_dff_B_bcYDuvh83_0),.clk(gclk));
	jdff dff_B_8PQLi2Av1_0(.din(w_dff_B_bcYDuvh83_0),.dout(w_dff_B_8PQLi2Av1_0),.clk(gclk));
	jdff dff_B_crRaYzpj9_0(.din(w_dff_B_8PQLi2Av1_0),.dout(w_dff_B_crRaYzpj9_0),.clk(gclk));
	jdff dff_B_dAp8PLhJ4_0(.din(w_dff_B_crRaYzpj9_0),.dout(w_dff_B_dAp8PLhJ4_0),.clk(gclk));
	jdff dff_B_fQ7FwhEU7_0(.din(w_dff_B_dAp8PLhJ4_0),.dout(w_dff_B_fQ7FwhEU7_0),.clk(gclk));
	jdff dff_B_UnsEc2uE7_0(.din(w_dff_B_fQ7FwhEU7_0),.dout(w_dff_B_UnsEc2uE7_0),.clk(gclk));
	jdff dff_B_pLQQcb9k9_0(.din(w_dff_B_UnsEc2uE7_0),.dout(w_dff_B_pLQQcb9k9_0),.clk(gclk));
	jdff dff_B_q1onKdbw1_0(.din(w_dff_B_pLQQcb9k9_0),.dout(w_dff_B_q1onKdbw1_0),.clk(gclk));
	jdff dff_B_90EtCyrN6_0(.din(w_dff_B_q1onKdbw1_0),.dout(w_dff_B_90EtCyrN6_0),.clk(gclk));
	jdff dff_B_tOouyl232_0(.din(n664),.dout(w_dff_B_tOouyl232_0),.clk(gclk));
	jdff dff_B_lFN408lB3_0(.din(w_dff_B_tOouyl232_0),.dout(w_dff_B_lFN408lB3_0),.clk(gclk));
	jdff dff_B_45Df4SvE2_0(.din(w_dff_B_lFN408lB3_0),.dout(w_dff_B_45Df4SvE2_0),.clk(gclk));
	jdff dff_B_U7sKnYuX5_0(.din(w_dff_B_45Df4SvE2_0),.dout(w_dff_B_U7sKnYuX5_0),.clk(gclk));
	jdff dff_B_uwZdqMql6_0(.din(w_dff_B_U7sKnYuX5_0),.dout(w_dff_B_uwZdqMql6_0),.clk(gclk));
	jdff dff_B_jKbNWyGV7_0(.din(w_dff_B_uwZdqMql6_0),.dout(w_dff_B_jKbNWyGV7_0),.clk(gclk));
	jdff dff_B_YkeJOvbQ8_0(.din(w_dff_B_jKbNWyGV7_0),.dout(w_dff_B_YkeJOvbQ8_0),.clk(gclk));
	jdff dff_B_OYCYOoLr7_0(.din(w_dff_B_YkeJOvbQ8_0),.dout(w_dff_B_OYCYOoLr7_0),.clk(gclk));
	jdff dff_B_lO2m5XBt1_0(.din(w_dff_B_OYCYOoLr7_0),.dout(w_dff_B_lO2m5XBt1_0),.clk(gclk));
	jdff dff_B_wIqwPaG54_0(.din(w_dff_B_lO2m5XBt1_0),.dout(w_dff_B_wIqwPaG54_0),.clk(gclk));
	jdff dff_B_eXa7IXzF1_0(.din(w_dff_B_wIqwPaG54_0),.dout(w_dff_B_eXa7IXzF1_0),.clk(gclk));
	jdff dff_B_zaA4lWdO2_0(.din(w_dff_B_eXa7IXzF1_0),.dout(w_dff_B_zaA4lWdO2_0),.clk(gclk));
	jdff dff_B_ynd9DkOR4_0(.din(w_dff_B_zaA4lWdO2_0),.dout(w_dff_B_ynd9DkOR4_0),.clk(gclk));
	jdff dff_B_4HGp9GPk0_0(.din(w_dff_B_ynd9DkOR4_0),.dout(w_dff_B_4HGp9GPk0_0),.clk(gclk));
	jdff dff_B_OmdS5XFl0_0(.din(w_dff_B_4HGp9GPk0_0),.dout(w_dff_B_OmdS5XFl0_0),.clk(gclk));
	jdff dff_B_nba7JulH1_0(.din(w_dff_B_OmdS5XFl0_0),.dout(w_dff_B_nba7JulH1_0),.clk(gclk));
	jdff dff_B_veUelKvJ3_0(.din(w_dff_B_nba7JulH1_0),.dout(w_dff_B_veUelKvJ3_0),.clk(gclk));
	jdff dff_B_tzpsxefS9_0(.din(w_dff_B_veUelKvJ3_0),.dout(w_dff_B_tzpsxefS9_0),.clk(gclk));
	jdff dff_B_QQFzepC22_0(.din(w_dff_B_tzpsxefS9_0),.dout(w_dff_B_QQFzepC22_0),.clk(gclk));
	jdff dff_B_186BDbZ64_0(.din(w_dff_B_QQFzepC22_0),.dout(w_dff_B_186BDbZ64_0),.clk(gclk));
	jdff dff_B_5U3yHgHO5_0(.din(w_dff_B_186BDbZ64_0),.dout(w_dff_B_5U3yHgHO5_0),.clk(gclk));
	jdff dff_B_ZMD0PT6v8_0(.din(w_dff_B_5U3yHgHO5_0),.dout(w_dff_B_ZMD0PT6v8_0),.clk(gclk));
	jdff dff_B_BlbrtC3g4_0(.din(w_dff_B_ZMD0PT6v8_0),.dout(w_dff_B_BlbrtC3g4_0),.clk(gclk));
	jdff dff_B_n153tEVi8_0(.din(w_dff_B_BlbrtC3g4_0),.dout(w_dff_B_n153tEVi8_0),.clk(gclk));
	jdff dff_B_wfbTXZfQ7_0(.din(w_dff_B_n153tEVi8_0),.dout(w_dff_B_wfbTXZfQ7_0),.clk(gclk));
	jdff dff_B_DsLZT1Gl4_0(.din(w_dff_B_wfbTXZfQ7_0),.dout(w_dff_B_DsLZT1Gl4_0),.clk(gclk));
	jdff dff_B_YSYKevg49_0(.din(w_dff_B_DsLZT1Gl4_0),.dout(w_dff_B_YSYKevg49_0),.clk(gclk));
	jdff dff_B_B6OwF0Vk7_0(.din(w_dff_B_YSYKevg49_0),.dout(w_dff_B_B6OwF0Vk7_0),.clk(gclk));
	jdff dff_B_eIv43cnw5_0(.din(w_dff_B_B6OwF0Vk7_0),.dout(w_dff_B_eIv43cnw5_0),.clk(gclk));
	jdff dff_B_FeesYoKp8_0(.din(w_dff_B_eIv43cnw5_0),.dout(w_dff_B_FeesYoKp8_0),.clk(gclk));
	jdff dff_B_Q2nhRqVk3_0(.din(w_dff_B_FeesYoKp8_0),.dout(w_dff_B_Q2nhRqVk3_0),.clk(gclk));
	jdff dff_B_6zUaJIuP2_0(.din(w_dff_B_Q2nhRqVk3_0),.dout(w_dff_B_6zUaJIuP2_0),.clk(gclk));
	jdff dff_B_EfnJsW652_0(.din(w_dff_B_6zUaJIuP2_0),.dout(w_dff_B_EfnJsW652_0),.clk(gclk));
	jdff dff_B_TVOrJfM53_0(.din(w_dff_B_EfnJsW652_0),.dout(w_dff_B_TVOrJfM53_0),.clk(gclk));
	jdff dff_B_lksUnRe12_0(.din(w_dff_B_TVOrJfM53_0),.dout(w_dff_B_lksUnRe12_0),.clk(gclk));
	jdff dff_B_kpiv2kOJ0_0(.din(w_dff_B_lksUnRe12_0),.dout(w_dff_B_kpiv2kOJ0_0),.clk(gclk));
	jdff dff_B_CJ4WeVhJ2_0(.din(w_dff_B_kpiv2kOJ0_0),.dout(w_dff_B_CJ4WeVhJ2_0),.clk(gclk));
	jdff dff_B_tWfZRAvY2_0(.din(w_dff_B_CJ4WeVhJ2_0),.dout(w_dff_B_tWfZRAvY2_0),.clk(gclk));
	jdff dff_B_LCpV3k1U4_0(.din(w_dff_B_tWfZRAvY2_0),.dout(w_dff_B_LCpV3k1U4_0),.clk(gclk));
	jdff dff_B_Gc1eLvwX5_0(.din(w_dff_B_LCpV3k1U4_0),.dout(w_dff_B_Gc1eLvwX5_0),.clk(gclk));
	jdff dff_B_ohQ0OD6A2_0(.din(w_dff_B_Gc1eLvwX5_0),.dout(w_dff_B_ohQ0OD6A2_0),.clk(gclk));
	jdff dff_B_dnOehzPz4_0(.din(w_dff_B_ohQ0OD6A2_0),.dout(w_dff_B_dnOehzPz4_0),.clk(gclk));
	jdff dff_B_h9TSedPf4_0(.din(w_dff_B_dnOehzPz4_0),.dout(w_dff_B_h9TSedPf4_0),.clk(gclk));
	jdff dff_B_fu6j3v8y6_0(.din(w_dff_B_h9TSedPf4_0),.dout(w_dff_B_fu6j3v8y6_0),.clk(gclk));
	jdff dff_B_6wxPVSvQ2_0(.din(w_dff_B_fu6j3v8y6_0),.dout(w_dff_B_6wxPVSvQ2_0),.clk(gclk));
	jdff dff_B_mkYl9cwU3_0(.din(w_dff_B_6wxPVSvQ2_0),.dout(w_dff_B_mkYl9cwU3_0),.clk(gclk));
	jdff dff_B_sekaV9lY2_0(.din(n670),.dout(w_dff_B_sekaV9lY2_0),.clk(gclk));
	jdff dff_B_s6xsKBGL4_0(.din(w_dff_B_sekaV9lY2_0),.dout(w_dff_B_s6xsKBGL4_0),.clk(gclk));
	jdff dff_B_LztGLYxd8_0(.din(w_dff_B_s6xsKBGL4_0),.dout(w_dff_B_LztGLYxd8_0),.clk(gclk));
	jdff dff_B_CiNhUuxW8_0(.din(w_dff_B_LztGLYxd8_0),.dout(w_dff_B_CiNhUuxW8_0),.clk(gclk));
	jdff dff_B_k7BLmRYR0_0(.din(w_dff_B_CiNhUuxW8_0),.dout(w_dff_B_k7BLmRYR0_0),.clk(gclk));
	jdff dff_B_dk4YZXBy8_0(.din(w_dff_B_k7BLmRYR0_0),.dout(w_dff_B_dk4YZXBy8_0),.clk(gclk));
	jdff dff_B_PfP3E5vl4_0(.din(w_dff_B_dk4YZXBy8_0),.dout(w_dff_B_PfP3E5vl4_0),.clk(gclk));
	jdff dff_B_qFKiqkCl0_0(.din(w_dff_B_PfP3E5vl4_0),.dout(w_dff_B_qFKiqkCl0_0),.clk(gclk));
	jdff dff_B_8uBRtBl74_0(.din(w_dff_B_qFKiqkCl0_0),.dout(w_dff_B_8uBRtBl74_0),.clk(gclk));
	jdff dff_B_Gw0bd02H8_0(.din(w_dff_B_8uBRtBl74_0),.dout(w_dff_B_Gw0bd02H8_0),.clk(gclk));
	jdff dff_B_WidWbth75_0(.din(w_dff_B_Gw0bd02H8_0),.dout(w_dff_B_WidWbth75_0),.clk(gclk));
	jdff dff_B_BSSA3qIB8_0(.din(w_dff_B_WidWbth75_0),.dout(w_dff_B_BSSA3qIB8_0),.clk(gclk));
	jdff dff_B_SU53ty9J8_0(.din(w_dff_B_BSSA3qIB8_0),.dout(w_dff_B_SU53ty9J8_0),.clk(gclk));
	jdff dff_B_7VIsqoqf7_0(.din(w_dff_B_SU53ty9J8_0),.dout(w_dff_B_7VIsqoqf7_0),.clk(gclk));
	jdff dff_B_nMD9NL467_0(.din(w_dff_B_7VIsqoqf7_0),.dout(w_dff_B_nMD9NL467_0),.clk(gclk));
	jdff dff_B_yBvmhV2d6_0(.din(w_dff_B_nMD9NL467_0),.dout(w_dff_B_yBvmhV2d6_0),.clk(gclk));
	jdff dff_B_VNHljr520_0(.din(w_dff_B_yBvmhV2d6_0),.dout(w_dff_B_VNHljr520_0),.clk(gclk));
	jdff dff_B_jeg0pcw54_0(.din(w_dff_B_VNHljr520_0),.dout(w_dff_B_jeg0pcw54_0),.clk(gclk));
	jdff dff_B_Ehnn5W3l9_0(.din(w_dff_B_jeg0pcw54_0),.dout(w_dff_B_Ehnn5W3l9_0),.clk(gclk));
	jdff dff_B_h6eZu3u20_0(.din(w_dff_B_Ehnn5W3l9_0),.dout(w_dff_B_h6eZu3u20_0),.clk(gclk));
	jdff dff_B_jJ915JOS1_0(.din(w_dff_B_h6eZu3u20_0),.dout(w_dff_B_jJ915JOS1_0),.clk(gclk));
	jdff dff_B_O7XTd4eo8_0(.din(w_dff_B_jJ915JOS1_0),.dout(w_dff_B_O7XTd4eo8_0),.clk(gclk));
	jdff dff_B_TBg2fwns5_0(.din(w_dff_B_O7XTd4eo8_0),.dout(w_dff_B_TBg2fwns5_0),.clk(gclk));
	jdff dff_B_Dvitz8RD4_0(.din(w_dff_B_TBg2fwns5_0),.dout(w_dff_B_Dvitz8RD4_0),.clk(gclk));
	jdff dff_B_LWByTZ2Q6_0(.din(w_dff_B_Dvitz8RD4_0),.dout(w_dff_B_LWByTZ2Q6_0),.clk(gclk));
	jdff dff_B_sxgDQVCz3_0(.din(w_dff_B_LWByTZ2Q6_0),.dout(w_dff_B_sxgDQVCz3_0),.clk(gclk));
	jdff dff_B_OgDfNBaa0_0(.din(w_dff_B_sxgDQVCz3_0),.dout(w_dff_B_OgDfNBaa0_0),.clk(gclk));
	jdff dff_B_dJodql2R1_0(.din(w_dff_B_OgDfNBaa0_0),.dout(w_dff_B_dJodql2R1_0),.clk(gclk));
	jdff dff_B_MMcPhios7_0(.din(w_dff_B_dJodql2R1_0),.dout(w_dff_B_MMcPhios7_0),.clk(gclk));
	jdff dff_B_NnBTvtU18_0(.din(w_dff_B_MMcPhios7_0),.dout(w_dff_B_NnBTvtU18_0),.clk(gclk));
	jdff dff_B_fpYlcgJ31_0(.din(w_dff_B_NnBTvtU18_0),.dout(w_dff_B_fpYlcgJ31_0),.clk(gclk));
	jdff dff_B_aUWkSl9d9_0(.din(w_dff_B_fpYlcgJ31_0),.dout(w_dff_B_aUWkSl9d9_0),.clk(gclk));
	jdff dff_B_yAb9gPcI9_0(.din(w_dff_B_aUWkSl9d9_0),.dout(w_dff_B_yAb9gPcI9_0),.clk(gclk));
	jdff dff_B_PRneCuUS5_0(.din(w_dff_B_yAb9gPcI9_0),.dout(w_dff_B_PRneCuUS5_0),.clk(gclk));
	jdff dff_B_4fwnKNCx5_0(.din(w_dff_B_PRneCuUS5_0),.dout(w_dff_B_4fwnKNCx5_0),.clk(gclk));
	jdff dff_B_tMQ513e39_0(.din(w_dff_B_4fwnKNCx5_0),.dout(w_dff_B_tMQ513e39_0),.clk(gclk));
	jdff dff_B_RjS5uZ9V2_0(.din(w_dff_B_tMQ513e39_0),.dout(w_dff_B_RjS5uZ9V2_0),.clk(gclk));
	jdff dff_B_S8ASuBaQ8_0(.din(w_dff_B_RjS5uZ9V2_0),.dout(w_dff_B_S8ASuBaQ8_0),.clk(gclk));
	jdff dff_B_OKgIkprX4_0(.din(w_dff_B_S8ASuBaQ8_0),.dout(w_dff_B_OKgIkprX4_0),.clk(gclk));
	jdff dff_B_we2ry5rk2_0(.din(w_dff_B_OKgIkprX4_0),.dout(w_dff_B_we2ry5rk2_0),.clk(gclk));
	jdff dff_B_tG45WYAK3_0(.din(w_dff_B_we2ry5rk2_0),.dout(w_dff_B_tG45WYAK3_0),.clk(gclk));
	jdff dff_B_ktByeRyp8_0(.din(w_dff_B_tG45WYAK3_0),.dout(w_dff_B_ktByeRyp8_0),.clk(gclk));
	jdff dff_B_OI0RpwXr6_0(.din(w_dff_B_ktByeRyp8_0),.dout(w_dff_B_OI0RpwXr6_0),.clk(gclk));
	jdff dff_B_7SaVDecC8_0(.din(w_dff_B_OI0RpwXr6_0),.dout(w_dff_B_7SaVDecC8_0),.clk(gclk));
	jdff dff_B_mP7mapQj4_0(.din(w_dff_B_7SaVDecC8_0),.dout(w_dff_B_mP7mapQj4_0),.clk(gclk));
	jdff dff_B_JcDN2b811_0(.din(w_dff_B_mP7mapQj4_0),.dout(w_dff_B_JcDN2b811_0),.clk(gclk));
	jdff dff_B_BfaZkbuX5_0(.din(w_dff_B_JcDN2b811_0),.dout(w_dff_B_BfaZkbuX5_0),.clk(gclk));
	jdff dff_B_yxDNEeLM8_0(.din(n676),.dout(w_dff_B_yxDNEeLM8_0),.clk(gclk));
	jdff dff_B_57i6nzTN8_0(.din(w_dff_B_yxDNEeLM8_0),.dout(w_dff_B_57i6nzTN8_0),.clk(gclk));
	jdff dff_B_2J8CZHmI3_0(.din(w_dff_B_57i6nzTN8_0),.dout(w_dff_B_2J8CZHmI3_0),.clk(gclk));
	jdff dff_B_psDzKZjJ4_0(.din(w_dff_B_2J8CZHmI3_0),.dout(w_dff_B_psDzKZjJ4_0),.clk(gclk));
	jdff dff_B_0VddD8N92_0(.din(w_dff_B_psDzKZjJ4_0),.dout(w_dff_B_0VddD8N92_0),.clk(gclk));
	jdff dff_B_L1BV0WJ00_0(.din(w_dff_B_0VddD8N92_0),.dout(w_dff_B_L1BV0WJ00_0),.clk(gclk));
	jdff dff_B_WswSo2lL0_0(.din(w_dff_B_L1BV0WJ00_0),.dout(w_dff_B_WswSo2lL0_0),.clk(gclk));
	jdff dff_B_CzFrxsGH7_0(.din(w_dff_B_WswSo2lL0_0),.dout(w_dff_B_CzFrxsGH7_0),.clk(gclk));
	jdff dff_B_5KsNWqcz0_0(.din(w_dff_B_CzFrxsGH7_0),.dout(w_dff_B_5KsNWqcz0_0),.clk(gclk));
	jdff dff_B_8sICLYOY8_0(.din(w_dff_B_5KsNWqcz0_0),.dout(w_dff_B_8sICLYOY8_0),.clk(gclk));
	jdff dff_B_p5pgjIrO1_0(.din(w_dff_B_8sICLYOY8_0),.dout(w_dff_B_p5pgjIrO1_0),.clk(gclk));
	jdff dff_B_s7QCceE05_0(.din(w_dff_B_p5pgjIrO1_0),.dout(w_dff_B_s7QCceE05_0),.clk(gclk));
	jdff dff_B_Ywwt6kAd5_0(.din(w_dff_B_s7QCceE05_0),.dout(w_dff_B_Ywwt6kAd5_0),.clk(gclk));
	jdff dff_B_IIKLaKLN3_0(.din(w_dff_B_Ywwt6kAd5_0),.dout(w_dff_B_IIKLaKLN3_0),.clk(gclk));
	jdff dff_B_OXyTg80H4_0(.din(w_dff_B_IIKLaKLN3_0),.dout(w_dff_B_OXyTg80H4_0),.clk(gclk));
	jdff dff_B_MSc4yDSg9_0(.din(w_dff_B_OXyTg80H4_0),.dout(w_dff_B_MSc4yDSg9_0),.clk(gclk));
	jdff dff_B_pqJLXFQp1_0(.din(w_dff_B_MSc4yDSg9_0),.dout(w_dff_B_pqJLXFQp1_0),.clk(gclk));
	jdff dff_B_Vfx3pym31_0(.din(w_dff_B_pqJLXFQp1_0),.dout(w_dff_B_Vfx3pym31_0),.clk(gclk));
	jdff dff_B_zt4I1oes2_0(.din(w_dff_B_Vfx3pym31_0),.dout(w_dff_B_zt4I1oes2_0),.clk(gclk));
	jdff dff_B_Yk6LgB6b9_0(.din(w_dff_B_zt4I1oes2_0),.dout(w_dff_B_Yk6LgB6b9_0),.clk(gclk));
	jdff dff_B_9aPdJM8K8_0(.din(w_dff_B_Yk6LgB6b9_0),.dout(w_dff_B_9aPdJM8K8_0),.clk(gclk));
	jdff dff_B_SmsNyQ917_0(.din(w_dff_B_9aPdJM8K8_0),.dout(w_dff_B_SmsNyQ917_0),.clk(gclk));
	jdff dff_B_Srpy44Sh5_0(.din(w_dff_B_SmsNyQ917_0),.dout(w_dff_B_Srpy44Sh5_0),.clk(gclk));
	jdff dff_B_LW8epFDI1_0(.din(w_dff_B_Srpy44Sh5_0),.dout(w_dff_B_LW8epFDI1_0),.clk(gclk));
	jdff dff_B_XtbzDpg11_0(.din(w_dff_B_LW8epFDI1_0),.dout(w_dff_B_XtbzDpg11_0),.clk(gclk));
	jdff dff_B_k2GTv2do1_0(.din(w_dff_B_XtbzDpg11_0),.dout(w_dff_B_k2GTv2do1_0),.clk(gclk));
	jdff dff_B_UBV3yPjF9_0(.din(w_dff_B_k2GTv2do1_0),.dout(w_dff_B_UBV3yPjF9_0),.clk(gclk));
	jdff dff_B_nhWUOYV77_0(.din(w_dff_B_UBV3yPjF9_0),.dout(w_dff_B_nhWUOYV77_0),.clk(gclk));
	jdff dff_B_OwAdHxPQ8_0(.din(w_dff_B_nhWUOYV77_0),.dout(w_dff_B_OwAdHxPQ8_0),.clk(gclk));
	jdff dff_B_fDafbnRY1_0(.din(w_dff_B_OwAdHxPQ8_0),.dout(w_dff_B_fDafbnRY1_0),.clk(gclk));
	jdff dff_B_RPwhy1YW9_0(.din(w_dff_B_fDafbnRY1_0),.dout(w_dff_B_RPwhy1YW9_0),.clk(gclk));
	jdff dff_B_ILpazNn41_0(.din(w_dff_B_RPwhy1YW9_0),.dout(w_dff_B_ILpazNn41_0),.clk(gclk));
	jdff dff_B_JuZidfGR8_0(.din(w_dff_B_ILpazNn41_0),.dout(w_dff_B_JuZidfGR8_0),.clk(gclk));
	jdff dff_B_TdQ3k8jt1_0(.din(w_dff_B_JuZidfGR8_0),.dout(w_dff_B_TdQ3k8jt1_0),.clk(gclk));
	jdff dff_B_TGMKnIs32_0(.din(w_dff_B_TdQ3k8jt1_0),.dout(w_dff_B_TGMKnIs32_0),.clk(gclk));
	jdff dff_B_3C1Z6RWy2_0(.din(w_dff_B_TGMKnIs32_0),.dout(w_dff_B_3C1Z6RWy2_0),.clk(gclk));
	jdff dff_B_ryw6tGTq3_0(.din(w_dff_B_3C1Z6RWy2_0),.dout(w_dff_B_ryw6tGTq3_0),.clk(gclk));
	jdff dff_B_9LLEM4Rk9_0(.din(w_dff_B_ryw6tGTq3_0),.dout(w_dff_B_9LLEM4Rk9_0),.clk(gclk));
	jdff dff_B_EutSCtWF0_0(.din(w_dff_B_9LLEM4Rk9_0),.dout(w_dff_B_EutSCtWF0_0),.clk(gclk));
	jdff dff_B_PQvP16zN4_0(.din(w_dff_B_EutSCtWF0_0),.dout(w_dff_B_PQvP16zN4_0),.clk(gclk));
	jdff dff_B_GPSvJbhD0_0(.din(w_dff_B_PQvP16zN4_0),.dout(w_dff_B_GPSvJbhD0_0),.clk(gclk));
	jdff dff_B_6BttYcdu8_0(.din(w_dff_B_GPSvJbhD0_0),.dout(w_dff_B_6BttYcdu8_0),.clk(gclk));
	jdff dff_B_169w74OF5_0(.din(w_dff_B_6BttYcdu8_0),.dout(w_dff_B_169w74OF5_0),.clk(gclk));
	jdff dff_B_v3tbDoey6_0(.din(w_dff_B_169w74OF5_0),.dout(w_dff_B_v3tbDoey6_0),.clk(gclk));
	jdff dff_B_uTo1T5Zm5_0(.din(w_dff_B_v3tbDoey6_0),.dout(w_dff_B_uTo1T5Zm5_0),.clk(gclk));
	jdff dff_B_gWZoEuR34_0(.din(w_dff_B_uTo1T5Zm5_0),.dout(w_dff_B_gWZoEuR34_0),.clk(gclk));
	jdff dff_B_E1wk1HtI2_0(.din(w_dff_B_gWZoEuR34_0),.dout(w_dff_B_E1wk1HtI2_0),.clk(gclk));
	jdff dff_B_DruCwV8I3_0(.din(w_dff_B_E1wk1HtI2_0),.dout(w_dff_B_DruCwV8I3_0),.clk(gclk));
	jdff dff_B_BUlLTBuT6_0(.din(n682),.dout(w_dff_B_BUlLTBuT6_0),.clk(gclk));
	jdff dff_B_oEbr8wJL8_0(.din(w_dff_B_BUlLTBuT6_0),.dout(w_dff_B_oEbr8wJL8_0),.clk(gclk));
	jdff dff_B_hiCdSWKo8_0(.din(w_dff_B_oEbr8wJL8_0),.dout(w_dff_B_hiCdSWKo8_0),.clk(gclk));
	jdff dff_B_rS70FZKg6_0(.din(w_dff_B_hiCdSWKo8_0),.dout(w_dff_B_rS70FZKg6_0),.clk(gclk));
	jdff dff_B_eqquUWVM5_0(.din(w_dff_B_rS70FZKg6_0),.dout(w_dff_B_eqquUWVM5_0),.clk(gclk));
	jdff dff_B_AUaRWg5r2_0(.din(w_dff_B_eqquUWVM5_0),.dout(w_dff_B_AUaRWg5r2_0),.clk(gclk));
	jdff dff_B_geFhxjpM3_0(.din(w_dff_B_AUaRWg5r2_0),.dout(w_dff_B_geFhxjpM3_0),.clk(gclk));
	jdff dff_B_owMPRISI1_0(.din(w_dff_B_geFhxjpM3_0),.dout(w_dff_B_owMPRISI1_0),.clk(gclk));
	jdff dff_B_6xRParBy0_0(.din(w_dff_B_owMPRISI1_0),.dout(w_dff_B_6xRParBy0_0),.clk(gclk));
	jdff dff_B_sdbroqEE6_0(.din(w_dff_B_6xRParBy0_0),.dout(w_dff_B_sdbroqEE6_0),.clk(gclk));
	jdff dff_B_Be2uaERX3_0(.din(w_dff_B_sdbroqEE6_0),.dout(w_dff_B_Be2uaERX3_0),.clk(gclk));
	jdff dff_B_EmFoRkGX3_0(.din(w_dff_B_Be2uaERX3_0),.dout(w_dff_B_EmFoRkGX3_0),.clk(gclk));
	jdff dff_B_6ViA2Bib7_0(.din(w_dff_B_EmFoRkGX3_0),.dout(w_dff_B_6ViA2Bib7_0),.clk(gclk));
	jdff dff_B_3eTgkbND3_0(.din(w_dff_B_6ViA2Bib7_0),.dout(w_dff_B_3eTgkbND3_0),.clk(gclk));
	jdff dff_B_3OO8t8Jy7_0(.din(w_dff_B_3eTgkbND3_0),.dout(w_dff_B_3OO8t8Jy7_0),.clk(gclk));
	jdff dff_B_F2g8Hgm21_0(.din(w_dff_B_3OO8t8Jy7_0),.dout(w_dff_B_F2g8Hgm21_0),.clk(gclk));
	jdff dff_B_wifpmEyU3_0(.din(w_dff_B_F2g8Hgm21_0),.dout(w_dff_B_wifpmEyU3_0),.clk(gclk));
	jdff dff_B_Inu1hAM00_0(.din(w_dff_B_wifpmEyU3_0),.dout(w_dff_B_Inu1hAM00_0),.clk(gclk));
	jdff dff_B_MVkbOYWV6_0(.din(w_dff_B_Inu1hAM00_0),.dout(w_dff_B_MVkbOYWV6_0),.clk(gclk));
	jdff dff_B_nYsC4c5E2_0(.din(w_dff_B_MVkbOYWV6_0),.dout(w_dff_B_nYsC4c5E2_0),.clk(gclk));
	jdff dff_B_c5HkVFLU9_0(.din(w_dff_B_nYsC4c5E2_0),.dout(w_dff_B_c5HkVFLU9_0),.clk(gclk));
	jdff dff_B_18VYH1cw3_0(.din(w_dff_B_c5HkVFLU9_0),.dout(w_dff_B_18VYH1cw3_0),.clk(gclk));
	jdff dff_B_rSnRLbSs2_0(.din(w_dff_B_18VYH1cw3_0),.dout(w_dff_B_rSnRLbSs2_0),.clk(gclk));
	jdff dff_B_eFeV68Nq8_0(.din(w_dff_B_rSnRLbSs2_0),.dout(w_dff_B_eFeV68Nq8_0),.clk(gclk));
	jdff dff_B_HW0oeEAb5_0(.din(w_dff_B_eFeV68Nq8_0),.dout(w_dff_B_HW0oeEAb5_0),.clk(gclk));
	jdff dff_B_K46a74sM1_0(.din(w_dff_B_HW0oeEAb5_0),.dout(w_dff_B_K46a74sM1_0),.clk(gclk));
	jdff dff_B_3dBMi0OY9_0(.din(w_dff_B_K46a74sM1_0),.dout(w_dff_B_3dBMi0OY9_0),.clk(gclk));
	jdff dff_B_9ev7klM63_0(.din(w_dff_B_3dBMi0OY9_0),.dout(w_dff_B_9ev7klM63_0),.clk(gclk));
	jdff dff_B_Rha8vPz39_0(.din(w_dff_B_9ev7klM63_0),.dout(w_dff_B_Rha8vPz39_0),.clk(gclk));
	jdff dff_B_wKvtrW0a8_0(.din(w_dff_B_Rha8vPz39_0),.dout(w_dff_B_wKvtrW0a8_0),.clk(gclk));
	jdff dff_B_1ruvJKk83_0(.din(w_dff_B_wKvtrW0a8_0),.dout(w_dff_B_1ruvJKk83_0),.clk(gclk));
	jdff dff_B_rd7NC96t0_0(.din(w_dff_B_1ruvJKk83_0),.dout(w_dff_B_rd7NC96t0_0),.clk(gclk));
	jdff dff_B_q8LGSXAh2_0(.din(w_dff_B_rd7NC96t0_0),.dout(w_dff_B_q8LGSXAh2_0),.clk(gclk));
	jdff dff_B_x44yHco41_0(.din(w_dff_B_q8LGSXAh2_0),.dout(w_dff_B_x44yHco41_0),.clk(gclk));
	jdff dff_B_hI0h6frj6_0(.din(w_dff_B_x44yHco41_0),.dout(w_dff_B_hI0h6frj6_0),.clk(gclk));
	jdff dff_B_iP2nRo9t5_0(.din(w_dff_B_hI0h6frj6_0),.dout(w_dff_B_iP2nRo9t5_0),.clk(gclk));
	jdff dff_B_i0z6fTE72_0(.din(w_dff_B_iP2nRo9t5_0),.dout(w_dff_B_i0z6fTE72_0),.clk(gclk));
	jdff dff_B_Sz7SJ7zR9_0(.din(w_dff_B_i0z6fTE72_0),.dout(w_dff_B_Sz7SJ7zR9_0),.clk(gclk));
	jdff dff_B_Nc7UXFJD6_0(.din(w_dff_B_Sz7SJ7zR9_0),.dout(w_dff_B_Nc7UXFJD6_0),.clk(gclk));
	jdff dff_B_gJMLFpCx6_0(.din(w_dff_B_Nc7UXFJD6_0),.dout(w_dff_B_gJMLFpCx6_0),.clk(gclk));
	jdff dff_B_Bei9iEcO9_0(.din(w_dff_B_gJMLFpCx6_0),.dout(w_dff_B_Bei9iEcO9_0),.clk(gclk));
	jdff dff_B_la3pvEnT1_0(.din(w_dff_B_Bei9iEcO9_0),.dout(w_dff_B_la3pvEnT1_0),.clk(gclk));
	jdff dff_B_K4Cen4Yd5_0(.din(w_dff_B_la3pvEnT1_0),.dout(w_dff_B_K4Cen4Yd5_0),.clk(gclk));
	jdff dff_B_LQoFq0ky3_0(.din(w_dff_B_K4Cen4Yd5_0),.dout(w_dff_B_LQoFq0ky3_0),.clk(gclk));
	jdff dff_B_ElBtdzJ98_0(.din(w_dff_B_LQoFq0ky3_0),.dout(w_dff_B_ElBtdzJ98_0),.clk(gclk));
	jdff dff_B_ZcFoxWzq4_0(.din(w_dff_B_ElBtdzJ98_0),.dout(w_dff_B_ZcFoxWzq4_0),.clk(gclk));
	jdff dff_B_lXKQqJnz9_0(.din(w_dff_B_ZcFoxWzq4_0),.dout(w_dff_B_lXKQqJnz9_0),.clk(gclk));
	jdff dff_B_kZJy5mzS5_0(.din(w_dff_B_lXKQqJnz9_0),.dout(w_dff_B_kZJy5mzS5_0),.clk(gclk));
	jdff dff_B_jmJiXT5P3_0(.din(w_dff_B_kZJy5mzS5_0),.dout(w_dff_B_jmJiXT5P3_0),.clk(gclk));
	jdff dff_B_sNAFJ17s9_0(.din(n688),.dout(w_dff_B_sNAFJ17s9_0),.clk(gclk));
	jdff dff_B_GY10BsD07_0(.din(w_dff_B_sNAFJ17s9_0),.dout(w_dff_B_GY10BsD07_0),.clk(gclk));
	jdff dff_B_4F7xIhH49_0(.din(w_dff_B_GY10BsD07_0),.dout(w_dff_B_4F7xIhH49_0),.clk(gclk));
	jdff dff_B_40TwRlPe2_0(.din(w_dff_B_4F7xIhH49_0),.dout(w_dff_B_40TwRlPe2_0),.clk(gclk));
	jdff dff_B_cnw7ZXrt7_0(.din(w_dff_B_40TwRlPe2_0),.dout(w_dff_B_cnw7ZXrt7_0),.clk(gclk));
	jdff dff_B_5wGIlZSw0_0(.din(w_dff_B_cnw7ZXrt7_0),.dout(w_dff_B_5wGIlZSw0_0),.clk(gclk));
	jdff dff_B_rUibQj4k7_0(.din(w_dff_B_5wGIlZSw0_0),.dout(w_dff_B_rUibQj4k7_0),.clk(gclk));
	jdff dff_B_JVisCbx96_0(.din(w_dff_B_rUibQj4k7_0),.dout(w_dff_B_JVisCbx96_0),.clk(gclk));
	jdff dff_B_K9bul2Ux1_0(.din(w_dff_B_JVisCbx96_0),.dout(w_dff_B_K9bul2Ux1_0),.clk(gclk));
	jdff dff_B_2K1zDfFj4_0(.din(w_dff_B_K9bul2Ux1_0),.dout(w_dff_B_2K1zDfFj4_0),.clk(gclk));
	jdff dff_B_LvzHN8Pt5_0(.din(w_dff_B_2K1zDfFj4_0),.dout(w_dff_B_LvzHN8Pt5_0),.clk(gclk));
	jdff dff_B_IsZmvvDz7_0(.din(w_dff_B_LvzHN8Pt5_0),.dout(w_dff_B_IsZmvvDz7_0),.clk(gclk));
	jdff dff_B_x6ZTmAG78_0(.din(w_dff_B_IsZmvvDz7_0),.dout(w_dff_B_x6ZTmAG78_0),.clk(gclk));
	jdff dff_B_Nnlu6zqz7_0(.din(w_dff_B_x6ZTmAG78_0),.dout(w_dff_B_Nnlu6zqz7_0),.clk(gclk));
	jdff dff_B_fl2YKFxC3_0(.din(w_dff_B_Nnlu6zqz7_0),.dout(w_dff_B_fl2YKFxC3_0),.clk(gclk));
	jdff dff_B_QafPK4mw6_0(.din(w_dff_B_fl2YKFxC3_0),.dout(w_dff_B_QafPK4mw6_0),.clk(gclk));
	jdff dff_B_aY0s1SEW5_0(.din(w_dff_B_QafPK4mw6_0),.dout(w_dff_B_aY0s1SEW5_0),.clk(gclk));
	jdff dff_B_dMpryHiW9_0(.din(w_dff_B_aY0s1SEW5_0),.dout(w_dff_B_dMpryHiW9_0),.clk(gclk));
	jdff dff_B_8jpwtIwW6_0(.din(w_dff_B_dMpryHiW9_0),.dout(w_dff_B_8jpwtIwW6_0),.clk(gclk));
	jdff dff_B_GGXDhljT5_0(.din(w_dff_B_8jpwtIwW6_0),.dout(w_dff_B_GGXDhljT5_0),.clk(gclk));
	jdff dff_B_0JOcTsYA2_0(.din(w_dff_B_GGXDhljT5_0),.dout(w_dff_B_0JOcTsYA2_0),.clk(gclk));
	jdff dff_B_zB6oGyAj9_0(.din(w_dff_B_0JOcTsYA2_0),.dout(w_dff_B_zB6oGyAj9_0),.clk(gclk));
	jdff dff_B_vBPOMeOQ3_0(.din(w_dff_B_zB6oGyAj9_0),.dout(w_dff_B_vBPOMeOQ3_0),.clk(gclk));
	jdff dff_B_IapBKDmK5_0(.din(w_dff_B_vBPOMeOQ3_0),.dout(w_dff_B_IapBKDmK5_0),.clk(gclk));
	jdff dff_B_ODRXgujl5_0(.din(w_dff_B_IapBKDmK5_0),.dout(w_dff_B_ODRXgujl5_0),.clk(gclk));
	jdff dff_B_jKPXe0550_0(.din(w_dff_B_ODRXgujl5_0),.dout(w_dff_B_jKPXe0550_0),.clk(gclk));
	jdff dff_B_Hd51AcOE8_0(.din(w_dff_B_jKPXe0550_0),.dout(w_dff_B_Hd51AcOE8_0),.clk(gclk));
	jdff dff_B_xBFkXBWB5_0(.din(w_dff_B_Hd51AcOE8_0),.dout(w_dff_B_xBFkXBWB5_0),.clk(gclk));
	jdff dff_B_dj7hx1W01_0(.din(w_dff_B_xBFkXBWB5_0),.dout(w_dff_B_dj7hx1W01_0),.clk(gclk));
	jdff dff_B_S8AfUY190_0(.din(w_dff_B_dj7hx1W01_0),.dout(w_dff_B_S8AfUY190_0),.clk(gclk));
	jdff dff_B_DXLQpCXf7_0(.din(w_dff_B_S8AfUY190_0),.dout(w_dff_B_DXLQpCXf7_0),.clk(gclk));
	jdff dff_B_JanyqvzG0_0(.din(w_dff_B_DXLQpCXf7_0),.dout(w_dff_B_JanyqvzG0_0),.clk(gclk));
	jdff dff_B_TCmfaA4x9_0(.din(w_dff_B_JanyqvzG0_0),.dout(w_dff_B_TCmfaA4x9_0),.clk(gclk));
	jdff dff_B_WvzYseF72_0(.din(w_dff_B_TCmfaA4x9_0),.dout(w_dff_B_WvzYseF72_0),.clk(gclk));
	jdff dff_B_6a4aBm4P1_0(.din(w_dff_B_WvzYseF72_0),.dout(w_dff_B_6a4aBm4P1_0),.clk(gclk));
	jdff dff_B_FtysMW8k5_0(.din(w_dff_B_6a4aBm4P1_0),.dout(w_dff_B_FtysMW8k5_0),.clk(gclk));
	jdff dff_B_Uon6fcLy0_0(.din(w_dff_B_FtysMW8k5_0),.dout(w_dff_B_Uon6fcLy0_0),.clk(gclk));
	jdff dff_B_9QZDgNNG5_0(.din(w_dff_B_Uon6fcLy0_0),.dout(w_dff_B_9QZDgNNG5_0),.clk(gclk));
	jdff dff_B_hbjWsio41_0(.din(w_dff_B_9QZDgNNG5_0),.dout(w_dff_B_hbjWsio41_0),.clk(gclk));
	jdff dff_B_OIsQTUTm0_0(.din(w_dff_B_hbjWsio41_0),.dout(w_dff_B_OIsQTUTm0_0),.clk(gclk));
	jdff dff_B_Yz3HFJhT3_0(.din(w_dff_B_OIsQTUTm0_0),.dout(w_dff_B_Yz3HFJhT3_0),.clk(gclk));
	jdff dff_B_OqAbfmLI4_0(.din(w_dff_B_Yz3HFJhT3_0),.dout(w_dff_B_OqAbfmLI4_0),.clk(gclk));
	jdff dff_B_MUt6SVHt2_0(.din(w_dff_B_OqAbfmLI4_0),.dout(w_dff_B_MUt6SVHt2_0),.clk(gclk));
	jdff dff_B_ibIrj1UC5_0(.din(w_dff_B_MUt6SVHt2_0),.dout(w_dff_B_ibIrj1UC5_0),.clk(gclk));
	jdff dff_B_IhYCeMkg9_0(.din(w_dff_B_ibIrj1UC5_0),.dout(w_dff_B_IhYCeMkg9_0),.clk(gclk));
	jdff dff_B_jZfDpBpZ8_0(.din(w_dff_B_IhYCeMkg9_0),.dout(w_dff_B_jZfDpBpZ8_0),.clk(gclk));
	jdff dff_B_fdwWzORe9_0(.din(w_dff_B_jZfDpBpZ8_0),.dout(w_dff_B_fdwWzORe9_0),.clk(gclk));
	jdff dff_B_Lls6lBYm8_0(.din(w_dff_B_fdwWzORe9_0),.dout(w_dff_B_Lls6lBYm8_0),.clk(gclk));
	jdff dff_B_3MewoJsf4_0(.din(w_dff_B_Lls6lBYm8_0),.dout(w_dff_B_3MewoJsf4_0),.clk(gclk));
	jdff dff_B_V9qk1Xe17_0(.din(w_dff_B_3MewoJsf4_0),.dout(w_dff_B_V9qk1Xe17_0),.clk(gclk));
	jdff dff_B_W0Q43Qoz4_0(.din(n694),.dout(w_dff_B_W0Q43Qoz4_0),.clk(gclk));
	jdff dff_B_sQA8Q7vv4_0(.din(w_dff_B_W0Q43Qoz4_0),.dout(w_dff_B_sQA8Q7vv4_0),.clk(gclk));
	jdff dff_B_mCg4hTSy1_0(.din(w_dff_B_sQA8Q7vv4_0),.dout(w_dff_B_mCg4hTSy1_0),.clk(gclk));
	jdff dff_B_BGPjhzNs0_0(.din(w_dff_B_mCg4hTSy1_0),.dout(w_dff_B_BGPjhzNs0_0),.clk(gclk));
	jdff dff_B_Z5d3liEd4_0(.din(w_dff_B_BGPjhzNs0_0),.dout(w_dff_B_Z5d3liEd4_0),.clk(gclk));
	jdff dff_B_JXBm3iQl2_0(.din(w_dff_B_Z5d3liEd4_0),.dout(w_dff_B_JXBm3iQl2_0),.clk(gclk));
	jdff dff_B_JA25AWF35_0(.din(w_dff_B_JXBm3iQl2_0),.dout(w_dff_B_JA25AWF35_0),.clk(gclk));
	jdff dff_B_BId30wwf6_0(.din(w_dff_B_JA25AWF35_0),.dout(w_dff_B_BId30wwf6_0),.clk(gclk));
	jdff dff_B_FqviFyMe3_0(.din(w_dff_B_BId30wwf6_0),.dout(w_dff_B_FqviFyMe3_0),.clk(gclk));
	jdff dff_B_LiFn6f3S2_0(.din(w_dff_B_FqviFyMe3_0),.dout(w_dff_B_LiFn6f3S2_0),.clk(gclk));
	jdff dff_B_XNuaHbLF9_0(.din(w_dff_B_LiFn6f3S2_0),.dout(w_dff_B_XNuaHbLF9_0),.clk(gclk));
	jdff dff_B_j4Dpw5Tz6_0(.din(w_dff_B_XNuaHbLF9_0),.dout(w_dff_B_j4Dpw5Tz6_0),.clk(gclk));
	jdff dff_B_uzC5qiMd1_0(.din(w_dff_B_j4Dpw5Tz6_0),.dout(w_dff_B_uzC5qiMd1_0),.clk(gclk));
	jdff dff_B_NmvSMw1S0_0(.din(w_dff_B_uzC5qiMd1_0),.dout(w_dff_B_NmvSMw1S0_0),.clk(gclk));
	jdff dff_B_FaiEpqTG7_0(.din(w_dff_B_NmvSMw1S0_0),.dout(w_dff_B_FaiEpqTG7_0),.clk(gclk));
	jdff dff_B_s6J6IifE4_0(.din(w_dff_B_FaiEpqTG7_0),.dout(w_dff_B_s6J6IifE4_0),.clk(gclk));
	jdff dff_B_jkLhY60Q6_0(.din(w_dff_B_s6J6IifE4_0),.dout(w_dff_B_jkLhY60Q6_0),.clk(gclk));
	jdff dff_B_plwjBdGt6_0(.din(w_dff_B_jkLhY60Q6_0),.dout(w_dff_B_plwjBdGt6_0),.clk(gclk));
	jdff dff_B_SFfPXqUT8_0(.din(w_dff_B_plwjBdGt6_0),.dout(w_dff_B_SFfPXqUT8_0),.clk(gclk));
	jdff dff_B_0OLCraVS5_0(.din(w_dff_B_SFfPXqUT8_0),.dout(w_dff_B_0OLCraVS5_0),.clk(gclk));
	jdff dff_B_E2dnobgi5_0(.din(w_dff_B_0OLCraVS5_0),.dout(w_dff_B_E2dnobgi5_0),.clk(gclk));
	jdff dff_B_3tj5RSZx6_0(.din(w_dff_B_E2dnobgi5_0),.dout(w_dff_B_3tj5RSZx6_0),.clk(gclk));
	jdff dff_B_zi1UCS4e0_0(.din(w_dff_B_3tj5RSZx6_0),.dout(w_dff_B_zi1UCS4e0_0),.clk(gclk));
	jdff dff_B_GS8UfAbF7_0(.din(w_dff_B_zi1UCS4e0_0),.dout(w_dff_B_GS8UfAbF7_0),.clk(gclk));
	jdff dff_B_by8f38tY4_0(.din(w_dff_B_GS8UfAbF7_0),.dout(w_dff_B_by8f38tY4_0),.clk(gclk));
	jdff dff_B_vvY2xB2h9_0(.din(w_dff_B_by8f38tY4_0),.dout(w_dff_B_vvY2xB2h9_0),.clk(gclk));
	jdff dff_B_r7R6QdA01_0(.din(w_dff_B_vvY2xB2h9_0),.dout(w_dff_B_r7R6QdA01_0),.clk(gclk));
	jdff dff_B_eUBIbbcW0_0(.din(w_dff_B_r7R6QdA01_0),.dout(w_dff_B_eUBIbbcW0_0),.clk(gclk));
	jdff dff_B_ZXBeAgIp8_0(.din(w_dff_B_eUBIbbcW0_0),.dout(w_dff_B_ZXBeAgIp8_0),.clk(gclk));
	jdff dff_B_FhfD9a3Z4_0(.din(w_dff_B_ZXBeAgIp8_0),.dout(w_dff_B_FhfD9a3Z4_0),.clk(gclk));
	jdff dff_B_qefyVb0a7_0(.din(w_dff_B_FhfD9a3Z4_0),.dout(w_dff_B_qefyVb0a7_0),.clk(gclk));
	jdff dff_B_peEQAwoh9_0(.din(w_dff_B_qefyVb0a7_0),.dout(w_dff_B_peEQAwoh9_0),.clk(gclk));
	jdff dff_B_egXWiJTJ1_0(.din(w_dff_B_peEQAwoh9_0),.dout(w_dff_B_egXWiJTJ1_0),.clk(gclk));
	jdff dff_B_2gX100wU4_0(.din(w_dff_B_egXWiJTJ1_0),.dout(w_dff_B_2gX100wU4_0),.clk(gclk));
	jdff dff_B_0cPouxdx1_0(.din(w_dff_B_2gX100wU4_0),.dout(w_dff_B_0cPouxdx1_0),.clk(gclk));
	jdff dff_B_9ku9ANK83_0(.din(w_dff_B_0cPouxdx1_0),.dout(w_dff_B_9ku9ANK83_0),.clk(gclk));
	jdff dff_B_g3ddMMgx6_0(.din(w_dff_B_9ku9ANK83_0),.dout(w_dff_B_g3ddMMgx6_0),.clk(gclk));
	jdff dff_B_R5L45zxX6_0(.din(w_dff_B_g3ddMMgx6_0),.dout(w_dff_B_R5L45zxX6_0),.clk(gclk));
	jdff dff_B_tZgsYkFL5_0(.din(w_dff_B_R5L45zxX6_0),.dout(w_dff_B_tZgsYkFL5_0),.clk(gclk));
	jdff dff_B_sSbbSwps5_0(.din(w_dff_B_tZgsYkFL5_0),.dout(w_dff_B_sSbbSwps5_0),.clk(gclk));
	jdff dff_B_1PFFfEyj3_0(.din(w_dff_B_sSbbSwps5_0),.dout(w_dff_B_1PFFfEyj3_0),.clk(gclk));
	jdff dff_B_vfGFsx5O2_0(.din(w_dff_B_1PFFfEyj3_0),.dout(w_dff_B_vfGFsx5O2_0),.clk(gclk));
	jdff dff_B_ziCdBN9y4_0(.din(w_dff_B_vfGFsx5O2_0),.dout(w_dff_B_ziCdBN9y4_0),.clk(gclk));
	jdff dff_B_MSvVpk5b0_0(.din(w_dff_B_ziCdBN9y4_0),.dout(w_dff_B_MSvVpk5b0_0),.clk(gclk));
	jdff dff_B_byECFDKU3_0(.din(w_dff_B_MSvVpk5b0_0),.dout(w_dff_B_byECFDKU3_0),.clk(gclk));
	jdff dff_B_nMB7fsea0_0(.din(w_dff_B_byECFDKU3_0),.dout(w_dff_B_nMB7fsea0_0),.clk(gclk));
	jdff dff_B_bzCYf9Yo1_0(.din(w_dff_B_nMB7fsea0_0),.dout(w_dff_B_bzCYf9Yo1_0),.clk(gclk));
	jdff dff_B_5O7IJApJ7_0(.din(w_dff_B_bzCYf9Yo1_0),.dout(w_dff_B_5O7IJApJ7_0),.clk(gclk));
	jdff dff_B_7HD4s21R5_0(.din(w_dff_B_5O7IJApJ7_0),.dout(w_dff_B_7HD4s21R5_0),.clk(gclk));
	jdff dff_B_ZcwQEUZV8_0(.din(w_dff_B_7HD4s21R5_0),.dout(w_dff_B_ZcwQEUZV8_0),.clk(gclk));
	jdff dff_B_oLurYfyu7_0(.din(w_dff_B_ZcwQEUZV8_0),.dout(w_dff_B_oLurYfyu7_0),.clk(gclk));
	jdff dff_B_4fMJkTpw4_0(.din(n700),.dout(w_dff_B_4fMJkTpw4_0),.clk(gclk));
	jdff dff_B_3cbsogQI9_0(.din(w_dff_B_4fMJkTpw4_0),.dout(w_dff_B_3cbsogQI9_0),.clk(gclk));
	jdff dff_B_Rbv02eXo8_0(.din(w_dff_B_3cbsogQI9_0),.dout(w_dff_B_Rbv02eXo8_0),.clk(gclk));
	jdff dff_B_nR0Dmvzw8_0(.din(w_dff_B_Rbv02eXo8_0),.dout(w_dff_B_nR0Dmvzw8_0),.clk(gclk));
	jdff dff_B_2bn6Tg174_0(.din(w_dff_B_nR0Dmvzw8_0),.dout(w_dff_B_2bn6Tg174_0),.clk(gclk));
	jdff dff_B_xyRRYFcf2_0(.din(w_dff_B_2bn6Tg174_0),.dout(w_dff_B_xyRRYFcf2_0),.clk(gclk));
	jdff dff_B_Cp6X42IN4_0(.din(w_dff_B_xyRRYFcf2_0),.dout(w_dff_B_Cp6X42IN4_0),.clk(gclk));
	jdff dff_B_Vmi8WjnT2_0(.din(w_dff_B_Cp6X42IN4_0),.dout(w_dff_B_Vmi8WjnT2_0),.clk(gclk));
	jdff dff_B_G17vDRnr2_0(.din(w_dff_B_Vmi8WjnT2_0),.dout(w_dff_B_G17vDRnr2_0),.clk(gclk));
	jdff dff_B_MvSJL1K94_0(.din(w_dff_B_G17vDRnr2_0),.dout(w_dff_B_MvSJL1K94_0),.clk(gclk));
	jdff dff_B_0cfnWS3U0_0(.din(w_dff_B_MvSJL1K94_0),.dout(w_dff_B_0cfnWS3U0_0),.clk(gclk));
	jdff dff_B_Q5WprNHv7_0(.din(w_dff_B_0cfnWS3U0_0),.dout(w_dff_B_Q5WprNHv7_0),.clk(gclk));
	jdff dff_B_IKDT7cE84_0(.din(w_dff_B_Q5WprNHv7_0),.dout(w_dff_B_IKDT7cE84_0),.clk(gclk));
	jdff dff_B_uxjXNiok6_0(.din(w_dff_B_IKDT7cE84_0),.dout(w_dff_B_uxjXNiok6_0),.clk(gclk));
	jdff dff_B_mIYGXKEz3_0(.din(w_dff_B_uxjXNiok6_0),.dout(w_dff_B_mIYGXKEz3_0),.clk(gclk));
	jdff dff_B_zs3lhyZS7_0(.din(w_dff_B_mIYGXKEz3_0),.dout(w_dff_B_zs3lhyZS7_0),.clk(gclk));
	jdff dff_B_ulKpnZJN8_0(.din(w_dff_B_zs3lhyZS7_0),.dout(w_dff_B_ulKpnZJN8_0),.clk(gclk));
	jdff dff_B_O78II1793_0(.din(w_dff_B_ulKpnZJN8_0),.dout(w_dff_B_O78II1793_0),.clk(gclk));
	jdff dff_B_UkCQW7Wl2_0(.din(w_dff_B_O78II1793_0),.dout(w_dff_B_UkCQW7Wl2_0),.clk(gclk));
	jdff dff_B_OwN5VRm39_0(.din(w_dff_B_UkCQW7Wl2_0),.dout(w_dff_B_OwN5VRm39_0),.clk(gclk));
	jdff dff_B_yxVi8SW62_0(.din(w_dff_B_OwN5VRm39_0),.dout(w_dff_B_yxVi8SW62_0),.clk(gclk));
	jdff dff_B_7YE2ABml3_0(.din(w_dff_B_yxVi8SW62_0),.dout(w_dff_B_7YE2ABml3_0),.clk(gclk));
	jdff dff_B_tu08v7UX3_0(.din(w_dff_B_7YE2ABml3_0),.dout(w_dff_B_tu08v7UX3_0),.clk(gclk));
	jdff dff_B_10M4d7Z52_0(.din(w_dff_B_tu08v7UX3_0),.dout(w_dff_B_10M4d7Z52_0),.clk(gclk));
	jdff dff_B_fRbqV2wy6_0(.din(w_dff_B_10M4d7Z52_0),.dout(w_dff_B_fRbqV2wy6_0),.clk(gclk));
	jdff dff_B_NyJsLI0T3_0(.din(w_dff_B_fRbqV2wy6_0),.dout(w_dff_B_NyJsLI0T3_0),.clk(gclk));
	jdff dff_B_XbVtB5Mq2_0(.din(w_dff_B_NyJsLI0T3_0),.dout(w_dff_B_XbVtB5Mq2_0),.clk(gclk));
	jdff dff_B_WAddHd7P2_0(.din(w_dff_B_XbVtB5Mq2_0),.dout(w_dff_B_WAddHd7P2_0),.clk(gclk));
	jdff dff_B_3sJIglB28_0(.din(w_dff_B_WAddHd7P2_0),.dout(w_dff_B_3sJIglB28_0),.clk(gclk));
	jdff dff_B_rOaV7Ugv6_0(.din(w_dff_B_3sJIglB28_0),.dout(w_dff_B_rOaV7Ugv6_0),.clk(gclk));
	jdff dff_B_bRfbUInS4_0(.din(w_dff_B_rOaV7Ugv6_0),.dout(w_dff_B_bRfbUInS4_0),.clk(gclk));
	jdff dff_B_nCKdcy2J1_0(.din(w_dff_B_bRfbUInS4_0),.dout(w_dff_B_nCKdcy2J1_0),.clk(gclk));
	jdff dff_B_dRT6h8il9_0(.din(w_dff_B_nCKdcy2J1_0),.dout(w_dff_B_dRT6h8il9_0),.clk(gclk));
	jdff dff_B_wSz2OSMi0_0(.din(w_dff_B_dRT6h8il9_0),.dout(w_dff_B_wSz2OSMi0_0),.clk(gclk));
	jdff dff_B_96zrmQzl9_0(.din(w_dff_B_wSz2OSMi0_0),.dout(w_dff_B_96zrmQzl9_0),.clk(gclk));
	jdff dff_B_ySTaNdRY2_0(.din(w_dff_B_96zrmQzl9_0),.dout(w_dff_B_ySTaNdRY2_0),.clk(gclk));
	jdff dff_B_hcLJBzb28_0(.din(w_dff_B_ySTaNdRY2_0),.dout(w_dff_B_hcLJBzb28_0),.clk(gclk));
	jdff dff_B_QmOxmh3e0_0(.din(w_dff_B_hcLJBzb28_0),.dout(w_dff_B_QmOxmh3e0_0),.clk(gclk));
	jdff dff_B_RXgXFbQm8_0(.din(w_dff_B_QmOxmh3e0_0),.dout(w_dff_B_RXgXFbQm8_0),.clk(gclk));
	jdff dff_B_43y5TZ5D9_0(.din(w_dff_B_RXgXFbQm8_0),.dout(w_dff_B_43y5TZ5D9_0),.clk(gclk));
	jdff dff_B_O25vugCd0_0(.din(w_dff_B_43y5TZ5D9_0),.dout(w_dff_B_O25vugCd0_0),.clk(gclk));
	jdff dff_B_KbCjAkss5_0(.din(w_dff_B_O25vugCd0_0),.dout(w_dff_B_KbCjAkss5_0),.clk(gclk));
	jdff dff_B_pZj7HHoE4_0(.din(w_dff_B_KbCjAkss5_0),.dout(w_dff_B_pZj7HHoE4_0),.clk(gclk));
	jdff dff_B_cU8nlsz34_0(.din(w_dff_B_pZj7HHoE4_0),.dout(w_dff_B_cU8nlsz34_0),.clk(gclk));
	jdff dff_B_uKfnj3hX2_0(.din(w_dff_B_cU8nlsz34_0),.dout(w_dff_B_uKfnj3hX2_0),.clk(gclk));
	jdff dff_B_217awbSP8_0(.din(w_dff_B_uKfnj3hX2_0),.dout(w_dff_B_217awbSP8_0),.clk(gclk));
	jdff dff_B_KjCxAh6I1_0(.din(w_dff_B_217awbSP8_0),.dout(w_dff_B_KjCxAh6I1_0),.clk(gclk));
	jdff dff_B_enEOtW2b9_0(.din(w_dff_B_KjCxAh6I1_0),.dout(w_dff_B_enEOtW2b9_0),.clk(gclk));
	jdff dff_B_9Qv9vLt90_0(.din(w_dff_B_enEOtW2b9_0),.dout(w_dff_B_9Qv9vLt90_0),.clk(gclk));
	jdff dff_B_SfvNzWud0_0(.din(w_dff_B_9Qv9vLt90_0),.dout(w_dff_B_SfvNzWud0_0),.clk(gclk));
	jdff dff_B_8Ckt47gu5_0(.din(w_dff_B_SfvNzWud0_0),.dout(w_dff_B_8Ckt47gu5_0),.clk(gclk));
	jdff dff_B_pKa8yGRz6_0(.din(w_dff_B_8Ckt47gu5_0),.dout(w_dff_B_pKa8yGRz6_0),.clk(gclk));
	jdff dff_B_19ToeBs49_0(.din(n706),.dout(w_dff_B_19ToeBs49_0),.clk(gclk));
	jdff dff_B_IPTl48vD7_0(.din(w_dff_B_19ToeBs49_0),.dout(w_dff_B_IPTl48vD7_0),.clk(gclk));
	jdff dff_B_HYG3fEyQ5_0(.din(w_dff_B_IPTl48vD7_0),.dout(w_dff_B_HYG3fEyQ5_0),.clk(gclk));
	jdff dff_B_U0anoE9b6_0(.din(w_dff_B_HYG3fEyQ5_0),.dout(w_dff_B_U0anoE9b6_0),.clk(gclk));
	jdff dff_B_IITT3hQl4_0(.din(w_dff_B_U0anoE9b6_0),.dout(w_dff_B_IITT3hQl4_0),.clk(gclk));
	jdff dff_B_zPfwqeM26_0(.din(w_dff_B_IITT3hQl4_0),.dout(w_dff_B_zPfwqeM26_0),.clk(gclk));
	jdff dff_B_dvk3k9Fa8_0(.din(w_dff_B_zPfwqeM26_0),.dout(w_dff_B_dvk3k9Fa8_0),.clk(gclk));
	jdff dff_B_1pp6wd6J6_0(.din(w_dff_B_dvk3k9Fa8_0),.dout(w_dff_B_1pp6wd6J6_0),.clk(gclk));
	jdff dff_B_bLzcn3G90_0(.din(w_dff_B_1pp6wd6J6_0),.dout(w_dff_B_bLzcn3G90_0),.clk(gclk));
	jdff dff_B_a332ttzI9_0(.din(w_dff_B_bLzcn3G90_0),.dout(w_dff_B_a332ttzI9_0),.clk(gclk));
	jdff dff_B_xUiDCcYZ3_0(.din(w_dff_B_a332ttzI9_0),.dout(w_dff_B_xUiDCcYZ3_0),.clk(gclk));
	jdff dff_B_R2YYj88I8_0(.din(w_dff_B_xUiDCcYZ3_0),.dout(w_dff_B_R2YYj88I8_0),.clk(gclk));
	jdff dff_B_GAwGDaAm2_0(.din(w_dff_B_R2YYj88I8_0),.dout(w_dff_B_GAwGDaAm2_0),.clk(gclk));
	jdff dff_B_bKAolXuJ8_0(.din(w_dff_B_GAwGDaAm2_0),.dout(w_dff_B_bKAolXuJ8_0),.clk(gclk));
	jdff dff_B_5cKWBSSc4_0(.din(w_dff_B_bKAolXuJ8_0),.dout(w_dff_B_5cKWBSSc4_0),.clk(gclk));
	jdff dff_B_z6cMncOa4_0(.din(w_dff_B_5cKWBSSc4_0),.dout(w_dff_B_z6cMncOa4_0),.clk(gclk));
	jdff dff_B_5oZj9Pw14_0(.din(w_dff_B_z6cMncOa4_0),.dout(w_dff_B_5oZj9Pw14_0),.clk(gclk));
	jdff dff_B_0VtMN9ot0_0(.din(w_dff_B_5oZj9Pw14_0),.dout(w_dff_B_0VtMN9ot0_0),.clk(gclk));
	jdff dff_B_3oBs2ErA5_0(.din(w_dff_B_0VtMN9ot0_0),.dout(w_dff_B_3oBs2ErA5_0),.clk(gclk));
	jdff dff_B_CdHiS3wE8_0(.din(w_dff_B_3oBs2ErA5_0),.dout(w_dff_B_CdHiS3wE8_0),.clk(gclk));
	jdff dff_B_X7KQmGk40_0(.din(w_dff_B_CdHiS3wE8_0),.dout(w_dff_B_X7KQmGk40_0),.clk(gclk));
	jdff dff_B_DA9hGyi26_0(.din(w_dff_B_X7KQmGk40_0),.dout(w_dff_B_DA9hGyi26_0),.clk(gclk));
	jdff dff_B_nrfe9TUa7_0(.din(w_dff_B_DA9hGyi26_0),.dout(w_dff_B_nrfe9TUa7_0),.clk(gclk));
	jdff dff_B_qm4t8A883_0(.din(w_dff_B_nrfe9TUa7_0),.dout(w_dff_B_qm4t8A883_0),.clk(gclk));
	jdff dff_B_NIzJ9Xhw8_0(.din(w_dff_B_qm4t8A883_0),.dout(w_dff_B_NIzJ9Xhw8_0),.clk(gclk));
	jdff dff_B_uapVjAvX0_0(.din(w_dff_B_NIzJ9Xhw8_0),.dout(w_dff_B_uapVjAvX0_0),.clk(gclk));
	jdff dff_B_nAQ4u5JI1_0(.din(w_dff_B_uapVjAvX0_0),.dout(w_dff_B_nAQ4u5JI1_0),.clk(gclk));
	jdff dff_B_Ibi5AWnv8_0(.din(w_dff_B_nAQ4u5JI1_0),.dout(w_dff_B_Ibi5AWnv8_0),.clk(gclk));
	jdff dff_B_nFoJi1rY6_0(.din(w_dff_B_Ibi5AWnv8_0),.dout(w_dff_B_nFoJi1rY6_0),.clk(gclk));
	jdff dff_B_WFA7gEuT7_0(.din(w_dff_B_nFoJi1rY6_0),.dout(w_dff_B_WFA7gEuT7_0),.clk(gclk));
	jdff dff_B_s9thuebF3_0(.din(w_dff_B_WFA7gEuT7_0),.dout(w_dff_B_s9thuebF3_0),.clk(gclk));
	jdff dff_B_8Qi4DYt31_0(.din(w_dff_B_s9thuebF3_0),.dout(w_dff_B_8Qi4DYt31_0),.clk(gclk));
	jdff dff_B_WGWJJZAy6_0(.din(w_dff_B_8Qi4DYt31_0),.dout(w_dff_B_WGWJJZAy6_0),.clk(gclk));
	jdff dff_B_gFYySWJQ0_0(.din(w_dff_B_WGWJJZAy6_0),.dout(w_dff_B_gFYySWJQ0_0),.clk(gclk));
	jdff dff_B_6De8olHu6_0(.din(w_dff_B_gFYySWJQ0_0),.dout(w_dff_B_6De8olHu6_0),.clk(gclk));
	jdff dff_B_KajAw35f7_0(.din(w_dff_B_6De8olHu6_0),.dout(w_dff_B_KajAw35f7_0),.clk(gclk));
	jdff dff_B_MK6rQC9c3_0(.din(w_dff_B_KajAw35f7_0),.dout(w_dff_B_MK6rQC9c3_0),.clk(gclk));
	jdff dff_B_mSydxlTZ4_0(.din(w_dff_B_MK6rQC9c3_0),.dout(w_dff_B_mSydxlTZ4_0),.clk(gclk));
	jdff dff_B_LAF4lqFX7_0(.din(w_dff_B_mSydxlTZ4_0),.dout(w_dff_B_LAF4lqFX7_0),.clk(gclk));
	jdff dff_B_yJvNFCgN8_0(.din(w_dff_B_LAF4lqFX7_0),.dout(w_dff_B_yJvNFCgN8_0),.clk(gclk));
	jdff dff_B_cIJTFFrx3_0(.din(w_dff_B_yJvNFCgN8_0),.dout(w_dff_B_cIJTFFrx3_0),.clk(gclk));
	jdff dff_B_d8Xh6XLg9_0(.din(w_dff_B_cIJTFFrx3_0),.dout(w_dff_B_d8Xh6XLg9_0),.clk(gclk));
	jdff dff_B_NDRUrUr44_0(.din(w_dff_B_d8Xh6XLg9_0),.dout(w_dff_B_NDRUrUr44_0),.clk(gclk));
	jdff dff_B_NJzcooRR5_0(.din(w_dff_B_NDRUrUr44_0),.dout(w_dff_B_NJzcooRR5_0),.clk(gclk));
	jdff dff_B_nI7y062u3_0(.din(w_dff_B_NJzcooRR5_0),.dout(w_dff_B_nI7y062u3_0),.clk(gclk));
	jdff dff_B_VeDz4Sxq6_0(.din(w_dff_B_nI7y062u3_0),.dout(w_dff_B_VeDz4Sxq6_0),.clk(gclk));
	jdff dff_B_oidi940U2_0(.din(w_dff_B_VeDz4Sxq6_0),.dout(w_dff_B_oidi940U2_0),.clk(gclk));
	jdff dff_B_jqYHvyuE2_0(.din(w_dff_B_oidi940U2_0),.dout(w_dff_B_jqYHvyuE2_0),.clk(gclk));
	jdff dff_B_fiEW4LIG5_0(.din(w_dff_B_jqYHvyuE2_0),.dout(w_dff_B_fiEW4LIG5_0),.clk(gclk));
	jdff dff_B_un4q9vJO5_0(.din(w_dff_B_fiEW4LIG5_0),.dout(w_dff_B_un4q9vJO5_0),.clk(gclk));
	jdff dff_B_4dsGElRY3_0(.din(w_dff_B_un4q9vJO5_0),.dout(w_dff_B_4dsGElRY3_0),.clk(gclk));
	jdff dff_B_PevDPDCH7_0(.din(w_dff_B_4dsGElRY3_0),.dout(w_dff_B_PevDPDCH7_0),.clk(gclk));
	jdff dff_B_U7KCbJ7j9_0(.din(w_dff_B_PevDPDCH7_0),.dout(w_dff_B_U7KCbJ7j9_0),.clk(gclk));
	jdff dff_B_5TuiCDz30_0(.din(n712),.dout(w_dff_B_5TuiCDz30_0),.clk(gclk));
	jdff dff_B_QjdKY39e7_0(.din(w_dff_B_5TuiCDz30_0),.dout(w_dff_B_QjdKY39e7_0),.clk(gclk));
	jdff dff_B_g2siNU406_0(.din(w_dff_B_QjdKY39e7_0),.dout(w_dff_B_g2siNU406_0),.clk(gclk));
	jdff dff_B_XbFs8ObF9_0(.din(w_dff_B_g2siNU406_0),.dout(w_dff_B_XbFs8ObF9_0),.clk(gclk));
	jdff dff_B_riJYA6HL1_0(.din(w_dff_B_XbFs8ObF9_0),.dout(w_dff_B_riJYA6HL1_0),.clk(gclk));
	jdff dff_B_DN2eSvy50_0(.din(w_dff_B_riJYA6HL1_0),.dout(w_dff_B_DN2eSvy50_0),.clk(gclk));
	jdff dff_B_omRn9OPr4_0(.din(w_dff_B_DN2eSvy50_0),.dout(w_dff_B_omRn9OPr4_0),.clk(gclk));
	jdff dff_B_Q9hWcdLx1_0(.din(w_dff_B_omRn9OPr4_0),.dout(w_dff_B_Q9hWcdLx1_0),.clk(gclk));
	jdff dff_B_C4A8BV2D9_0(.din(w_dff_B_Q9hWcdLx1_0),.dout(w_dff_B_C4A8BV2D9_0),.clk(gclk));
	jdff dff_B_jQlTkKXq3_0(.din(w_dff_B_C4A8BV2D9_0),.dout(w_dff_B_jQlTkKXq3_0),.clk(gclk));
	jdff dff_B_vzCeTABr8_0(.din(w_dff_B_jQlTkKXq3_0),.dout(w_dff_B_vzCeTABr8_0),.clk(gclk));
	jdff dff_B_eyEC9i7o9_0(.din(w_dff_B_vzCeTABr8_0),.dout(w_dff_B_eyEC9i7o9_0),.clk(gclk));
	jdff dff_B_Nu6GfRHJ2_0(.din(w_dff_B_eyEC9i7o9_0),.dout(w_dff_B_Nu6GfRHJ2_0),.clk(gclk));
	jdff dff_B_RoUAEUQC6_0(.din(w_dff_B_Nu6GfRHJ2_0),.dout(w_dff_B_RoUAEUQC6_0),.clk(gclk));
	jdff dff_B_V9WSAKDa9_0(.din(w_dff_B_RoUAEUQC6_0),.dout(w_dff_B_V9WSAKDa9_0),.clk(gclk));
	jdff dff_B_c19DGE9n1_0(.din(w_dff_B_V9WSAKDa9_0),.dout(w_dff_B_c19DGE9n1_0),.clk(gclk));
	jdff dff_B_lETFpnV44_0(.din(w_dff_B_c19DGE9n1_0),.dout(w_dff_B_lETFpnV44_0),.clk(gclk));
	jdff dff_B_oOk6Qdk90_0(.din(w_dff_B_lETFpnV44_0),.dout(w_dff_B_oOk6Qdk90_0),.clk(gclk));
	jdff dff_B_6O6Ff7HW3_0(.din(w_dff_B_oOk6Qdk90_0),.dout(w_dff_B_6O6Ff7HW3_0),.clk(gclk));
	jdff dff_B_3E7xKsAN8_0(.din(w_dff_B_6O6Ff7HW3_0),.dout(w_dff_B_3E7xKsAN8_0),.clk(gclk));
	jdff dff_B_qfXNonHn6_0(.din(w_dff_B_3E7xKsAN8_0),.dout(w_dff_B_qfXNonHn6_0),.clk(gclk));
	jdff dff_B_HIHTiZ7C7_0(.din(w_dff_B_qfXNonHn6_0),.dout(w_dff_B_HIHTiZ7C7_0),.clk(gclk));
	jdff dff_B_U0xETE0X2_0(.din(w_dff_B_HIHTiZ7C7_0),.dout(w_dff_B_U0xETE0X2_0),.clk(gclk));
	jdff dff_B_s7O2DkFm3_0(.din(w_dff_B_U0xETE0X2_0),.dout(w_dff_B_s7O2DkFm3_0),.clk(gclk));
	jdff dff_B_SVQM3aM76_0(.din(w_dff_B_s7O2DkFm3_0),.dout(w_dff_B_SVQM3aM76_0),.clk(gclk));
	jdff dff_B_EJoxtvbF2_0(.din(w_dff_B_SVQM3aM76_0),.dout(w_dff_B_EJoxtvbF2_0),.clk(gclk));
	jdff dff_B_gbeiSyXG1_0(.din(w_dff_B_EJoxtvbF2_0),.dout(w_dff_B_gbeiSyXG1_0),.clk(gclk));
	jdff dff_B_683DXW4G1_0(.din(w_dff_B_gbeiSyXG1_0),.dout(w_dff_B_683DXW4G1_0),.clk(gclk));
	jdff dff_B_BmhnnDgj4_0(.din(w_dff_B_683DXW4G1_0),.dout(w_dff_B_BmhnnDgj4_0),.clk(gclk));
	jdff dff_B_5bAtp4r32_0(.din(w_dff_B_BmhnnDgj4_0),.dout(w_dff_B_5bAtp4r32_0),.clk(gclk));
	jdff dff_B_CjopLBoS1_0(.din(w_dff_B_5bAtp4r32_0),.dout(w_dff_B_CjopLBoS1_0),.clk(gclk));
	jdff dff_B_ttaQeut41_0(.din(w_dff_B_CjopLBoS1_0),.dout(w_dff_B_ttaQeut41_0),.clk(gclk));
	jdff dff_B_xuig0HHX7_0(.din(w_dff_B_ttaQeut41_0),.dout(w_dff_B_xuig0HHX7_0),.clk(gclk));
	jdff dff_B_McHRGvS39_0(.din(w_dff_B_xuig0HHX7_0),.dout(w_dff_B_McHRGvS39_0),.clk(gclk));
	jdff dff_B_IDjDcG623_0(.din(w_dff_B_McHRGvS39_0),.dout(w_dff_B_IDjDcG623_0),.clk(gclk));
	jdff dff_B_XSeuToPy2_0(.din(w_dff_B_IDjDcG623_0),.dout(w_dff_B_XSeuToPy2_0),.clk(gclk));
	jdff dff_B_PDpSigoa0_0(.din(w_dff_B_XSeuToPy2_0),.dout(w_dff_B_PDpSigoa0_0),.clk(gclk));
	jdff dff_B_34pJQqSm4_0(.din(w_dff_B_PDpSigoa0_0),.dout(w_dff_B_34pJQqSm4_0),.clk(gclk));
	jdff dff_B_ikr9acNu9_0(.din(w_dff_B_34pJQqSm4_0),.dout(w_dff_B_ikr9acNu9_0),.clk(gclk));
	jdff dff_B_UA4W1WE27_0(.din(w_dff_B_ikr9acNu9_0),.dout(w_dff_B_UA4W1WE27_0),.clk(gclk));
	jdff dff_B_iBHJO64Z5_0(.din(w_dff_B_UA4W1WE27_0),.dout(w_dff_B_iBHJO64Z5_0),.clk(gclk));
	jdff dff_B_Rh4MhzGV0_0(.din(w_dff_B_iBHJO64Z5_0),.dout(w_dff_B_Rh4MhzGV0_0),.clk(gclk));
	jdff dff_B_LQXrrTHw1_0(.din(w_dff_B_Rh4MhzGV0_0),.dout(w_dff_B_LQXrrTHw1_0),.clk(gclk));
	jdff dff_B_ckVcF37S6_0(.din(w_dff_B_LQXrrTHw1_0),.dout(w_dff_B_ckVcF37S6_0),.clk(gclk));
	jdff dff_B_yOJi19wI4_0(.din(w_dff_B_ckVcF37S6_0),.dout(w_dff_B_yOJi19wI4_0),.clk(gclk));
	jdff dff_B_5hWvwEST9_0(.din(w_dff_B_yOJi19wI4_0),.dout(w_dff_B_5hWvwEST9_0),.clk(gclk));
	jdff dff_B_5QJS6uLd2_0(.din(w_dff_B_5hWvwEST9_0),.dout(w_dff_B_5QJS6uLd2_0),.clk(gclk));
	jdff dff_B_SnZrmw4R8_0(.din(w_dff_B_5QJS6uLd2_0),.dout(w_dff_B_SnZrmw4R8_0),.clk(gclk));
	jdff dff_B_ozoqehRA8_0(.din(w_dff_B_SnZrmw4R8_0),.dout(w_dff_B_ozoqehRA8_0),.clk(gclk));
	jdff dff_B_g3SxB9Dm7_0(.din(w_dff_B_ozoqehRA8_0),.dout(w_dff_B_g3SxB9Dm7_0),.clk(gclk));
	jdff dff_B_jl9lQTkz5_0(.din(w_dff_B_g3SxB9Dm7_0),.dout(w_dff_B_jl9lQTkz5_0),.clk(gclk));
	jdff dff_B_7gY3sxkf2_0(.din(w_dff_B_jl9lQTkz5_0),.dout(w_dff_B_7gY3sxkf2_0),.clk(gclk));
	jdff dff_B_bCXGpT5d5_0(.din(w_dff_B_7gY3sxkf2_0),.dout(w_dff_B_bCXGpT5d5_0),.clk(gclk));
	jdff dff_B_vinPkQyy1_0(.din(w_dff_B_bCXGpT5d5_0),.dout(w_dff_B_vinPkQyy1_0),.clk(gclk));
	jdff dff_B_RZADuqLD0_0(.din(n718),.dout(w_dff_B_RZADuqLD0_0),.clk(gclk));
	jdff dff_B_qMgMRE2O0_0(.din(w_dff_B_RZADuqLD0_0),.dout(w_dff_B_qMgMRE2O0_0),.clk(gclk));
	jdff dff_B_DMyIg8314_0(.din(w_dff_B_qMgMRE2O0_0),.dout(w_dff_B_DMyIg8314_0),.clk(gclk));
	jdff dff_B_acXU7HXC4_0(.din(w_dff_B_DMyIg8314_0),.dout(w_dff_B_acXU7HXC4_0),.clk(gclk));
	jdff dff_B_FugCq6a90_0(.din(w_dff_B_acXU7HXC4_0),.dout(w_dff_B_FugCq6a90_0),.clk(gclk));
	jdff dff_B_xzgIeZa82_0(.din(w_dff_B_FugCq6a90_0),.dout(w_dff_B_xzgIeZa82_0),.clk(gclk));
	jdff dff_B_AYtav6441_0(.din(w_dff_B_xzgIeZa82_0),.dout(w_dff_B_AYtav6441_0),.clk(gclk));
	jdff dff_B_H7tT1WGg7_0(.din(w_dff_B_AYtav6441_0),.dout(w_dff_B_H7tT1WGg7_0),.clk(gclk));
	jdff dff_B_3OyFvk4g5_0(.din(w_dff_B_H7tT1WGg7_0),.dout(w_dff_B_3OyFvk4g5_0),.clk(gclk));
	jdff dff_B_4CNIiIZT6_0(.din(w_dff_B_3OyFvk4g5_0),.dout(w_dff_B_4CNIiIZT6_0),.clk(gclk));
	jdff dff_B_aoqb0R2S4_0(.din(w_dff_B_4CNIiIZT6_0),.dout(w_dff_B_aoqb0R2S4_0),.clk(gclk));
	jdff dff_B_xwJz2MHm6_0(.din(w_dff_B_aoqb0R2S4_0),.dout(w_dff_B_xwJz2MHm6_0),.clk(gclk));
	jdff dff_B_feSsaIf44_0(.din(w_dff_B_xwJz2MHm6_0),.dout(w_dff_B_feSsaIf44_0),.clk(gclk));
	jdff dff_B_SkkzHgmv3_0(.din(w_dff_B_feSsaIf44_0),.dout(w_dff_B_SkkzHgmv3_0),.clk(gclk));
	jdff dff_B_0vsm1U1t4_0(.din(w_dff_B_SkkzHgmv3_0),.dout(w_dff_B_0vsm1U1t4_0),.clk(gclk));
	jdff dff_B_Y7ZAL5IZ0_0(.din(w_dff_B_0vsm1U1t4_0),.dout(w_dff_B_Y7ZAL5IZ0_0),.clk(gclk));
	jdff dff_B_1EBayVfX0_0(.din(w_dff_B_Y7ZAL5IZ0_0),.dout(w_dff_B_1EBayVfX0_0),.clk(gclk));
	jdff dff_B_XimjgfD55_0(.din(w_dff_B_1EBayVfX0_0),.dout(w_dff_B_XimjgfD55_0),.clk(gclk));
	jdff dff_B_VLCqTYut9_0(.din(w_dff_B_XimjgfD55_0),.dout(w_dff_B_VLCqTYut9_0),.clk(gclk));
	jdff dff_B_sARaI0Ke1_0(.din(w_dff_B_VLCqTYut9_0),.dout(w_dff_B_sARaI0Ke1_0),.clk(gclk));
	jdff dff_B_CVZrcz8n5_0(.din(w_dff_B_sARaI0Ke1_0),.dout(w_dff_B_CVZrcz8n5_0),.clk(gclk));
	jdff dff_B_HyGs87ZG4_0(.din(w_dff_B_CVZrcz8n5_0),.dout(w_dff_B_HyGs87ZG4_0),.clk(gclk));
	jdff dff_B_kv9GIGkv4_0(.din(w_dff_B_HyGs87ZG4_0),.dout(w_dff_B_kv9GIGkv4_0),.clk(gclk));
	jdff dff_B_5zy633b08_0(.din(w_dff_B_kv9GIGkv4_0),.dout(w_dff_B_5zy633b08_0),.clk(gclk));
	jdff dff_B_NaTYdP5T6_0(.din(w_dff_B_5zy633b08_0),.dout(w_dff_B_NaTYdP5T6_0),.clk(gclk));
	jdff dff_B_QTy547KM6_0(.din(w_dff_B_NaTYdP5T6_0),.dout(w_dff_B_QTy547KM6_0),.clk(gclk));
	jdff dff_B_bwENjw0O5_0(.din(w_dff_B_QTy547KM6_0),.dout(w_dff_B_bwENjw0O5_0),.clk(gclk));
	jdff dff_B_DONxhJQu0_0(.din(w_dff_B_bwENjw0O5_0),.dout(w_dff_B_DONxhJQu0_0),.clk(gclk));
	jdff dff_B_0KY7RqAv0_0(.din(w_dff_B_DONxhJQu0_0),.dout(w_dff_B_0KY7RqAv0_0),.clk(gclk));
	jdff dff_B_v2XPfulv5_0(.din(w_dff_B_0KY7RqAv0_0),.dout(w_dff_B_v2XPfulv5_0),.clk(gclk));
	jdff dff_B_iwOAdbGe8_0(.din(w_dff_B_v2XPfulv5_0),.dout(w_dff_B_iwOAdbGe8_0),.clk(gclk));
	jdff dff_B_lj5oT0lg6_0(.din(w_dff_B_iwOAdbGe8_0),.dout(w_dff_B_lj5oT0lg6_0),.clk(gclk));
	jdff dff_B_b9TMSY913_0(.din(w_dff_B_lj5oT0lg6_0),.dout(w_dff_B_b9TMSY913_0),.clk(gclk));
	jdff dff_B_DTD5nbG36_0(.din(w_dff_B_b9TMSY913_0),.dout(w_dff_B_DTD5nbG36_0),.clk(gclk));
	jdff dff_B_iTPMRVvg6_0(.din(w_dff_B_DTD5nbG36_0),.dout(w_dff_B_iTPMRVvg6_0),.clk(gclk));
	jdff dff_B_tiske0pB1_0(.din(w_dff_B_iTPMRVvg6_0),.dout(w_dff_B_tiske0pB1_0),.clk(gclk));
	jdff dff_B_KUdz2CJa8_0(.din(w_dff_B_tiske0pB1_0),.dout(w_dff_B_KUdz2CJa8_0),.clk(gclk));
	jdff dff_B_X3NPnCiV5_0(.din(w_dff_B_KUdz2CJa8_0),.dout(w_dff_B_X3NPnCiV5_0),.clk(gclk));
	jdff dff_B_n0H4Z3Uk4_0(.din(w_dff_B_X3NPnCiV5_0),.dout(w_dff_B_n0H4Z3Uk4_0),.clk(gclk));
	jdff dff_B_cCLBdCMf8_0(.din(w_dff_B_n0H4Z3Uk4_0),.dout(w_dff_B_cCLBdCMf8_0),.clk(gclk));
	jdff dff_B_BVJmrVS73_0(.din(w_dff_B_cCLBdCMf8_0),.dout(w_dff_B_BVJmrVS73_0),.clk(gclk));
	jdff dff_B_Hls79WUD8_0(.din(w_dff_B_BVJmrVS73_0),.dout(w_dff_B_Hls79WUD8_0),.clk(gclk));
	jdff dff_B_uma5x3EP1_0(.din(w_dff_B_Hls79WUD8_0),.dout(w_dff_B_uma5x3EP1_0),.clk(gclk));
	jdff dff_B_O4OgeXrX5_0(.din(w_dff_B_uma5x3EP1_0),.dout(w_dff_B_O4OgeXrX5_0),.clk(gclk));
	jdff dff_B_XFvWNnpT5_0(.din(w_dff_B_O4OgeXrX5_0),.dout(w_dff_B_XFvWNnpT5_0),.clk(gclk));
	jdff dff_B_FdDuKjM23_0(.din(w_dff_B_XFvWNnpT5_0),.dout(w_dff_B_FdDuKjM23_0),.clk(gclk));
	jdff dff_B_BpfTb8Mn0_0(.din(w_dff_B_FdDuKjM23_0),.dout(w_dff_B_BpfTb8Mn0_0),.clk(gclk));
	jdff dff_B_6YZ0MEFL6_0(.din(w_dff_B_BpfTb8Mn0_0),.dout(w_dff_B_6YZ0MEFL6_0),.clk(gclk));
	jdff dff_B_R9Rapnri9_0(.din(w_dff_B_6YZ0MEFL6_0),.dout(w_dff_B_R9Rapnri9_0),.clk(gclk));
	jdff dff_B_fjRGz4vp6_0(.din(w_dff_B_R9Rapnri9_0),.dout(w_dff_B_fjRGz4vp6_0),.clk(gclk));
	jdff dff_B_tQF2amq15_0(.din(w_dff_B_fjRGz4vp6_0),.dout(w_dff_B_tQF2amq15_0),.clk(gclk));
	jdff dff_B_DexEJ0qv7_0(.din(w_dff_B_tQF2amq15_0),.dout(w_dff_B_DexEJ0qv7_0),.clk(gclk));
	jdff dff_B_iTGijb4G3_0(.din(w_dff_B_DexEJ0qv7_0),.dout(w_dff_B_iTGijb4G3_0),.clk(gclk));
	jdff dff_B_OBMEBLRR5_0(.din(w_dff_B_iTGijb4G3_0),.dout(w_dff_B_OBMEBLRR5_0),.clk(gclk));
	jdff dff_B_YzSXgHQL7_0(.din(w_dff_B_OBMEBLRR5_0),.dout(w_dff_B_YzSXgHQL7_0),.clk(gclk));
	jdff dff_B_iLhXKM2I1_0(.din(n724),.dout(w_dff_B_iLhXKM2I1_0),.clk(gclk));
	jdff dff_B_DF3UfJ7A4_0(.din(w_dff_B_iLhXKM2I1_0),.dout(w_dff_B_DF3UfJ7A4_0),.clk(gclk));
	jdff dff_B_WBrmP0OL6_0(.din(w_dff_B_DF3UfJ7A4_0),.dout(w_dff_B_WBrmP0OL6_0),.clk(gclk));
	jdff dff_B_M32JFkM21_0(.din(w_dff_B_WBrmP0OL6_0),.dout(w_dff_B_M32JFkM21_0),.clk(gclk));
	jdff dff_B_TbxqKTGH9_0(.din(w_dff_B_M32JFkM21_0),.dout(w_dff_B_TbxqKTGH9_0),.clk(gclk));
	jdff dff_B_NtFQpDHd1_0(.din(w_dff_B_TbxqKTGH9_0),.dout(w_dff_B_NtFQpDHd1_0),.clk(gclk));
	jdff dff_B_i2ZeriDB6_0(.din(w_dff_B_NtFQpDHd1_0),.dout(w_dff_B_i2ZeriDB6_0),.clk(gclk));
	jdff dff_B_Y0i3i1aI8_0(.din(w_dff_B_i2ZeriDB6_0),.dout(w_dff_B_Y0i3i1aI8_0),.clk(gclk));
	jdff dff_B_kJ1OIEFu0_0(.din(w_dff_B_Y0i3i1aI8_0),.dout(w_dff_B_kJ1OIEFu0_0),.clk(gclk));
	jdff dff_B_515I7mq45_0(.din(w_dff_B_kJ1OIEFu0_0),.dout(w_dff_B_515I7mq45_0),.clk(gclk));
	jdff dff_B_Oeu12Ync6_0(.din(w_dff_B_515I7mq45_0),.dout(w_dff_B_Oeu12Ync6_0),.clk(gclk));
	jdff dff_B_vW9kxOqW9_0(.din(w_dff_B_Oeu12Ync6_0),.dout(w_dff_B_vW9kxOqW9_0),.clk(gclk));
	jdff dff_B_cDVxcvt91_0(.din(w_dff_B_vW9kxOqW9_0),.dout(w_dff_B_cDVxcvt91_0),.clk(gclk));
	jdff dff_B_pJtGYLR11_0(.din(w_dff_B_cDVxcvt91_0),.dout(w_dff_B_pJtGYLR11_0),.clk(gclk));
	jdff dff_B_q9r0iuA15_0(.din(w_dff_B_pJtGYLR11_0),.dout(w_dff_B_q9r0iuA15_0),.clk(gclk));
	jdff dff_B_xNHUsXCf0_0(.din(w_dff_B_q9r0iuA15_0),.dout(w_dff_B_xNHUsXCf0_0),.clk(gclk));
	jdff dff_B_CTyWitmH7_0(.din(w_dff_B_xNHUsXCf0_0),.dout(w_dff_B_CTyWitmH7_0),.clk(gclk));
	jdff dff_B_HbI5Xm1a1_0(.din(w_dff_B_CTyWitmH7_0),.dout(w_dff_B_HbI5Xm1a1_0),.clk(gclk));
	jdff dff_B_HvZTQnBa6_0(.din(w_dff_B_HbI5Xm1a1_0),.dout(w_dff_B_HvZTQnBa6_0),.clk(gclk));
	jdff dff_B_GaY4qt4a6_0(.din(w_dff_B_HvZTQnBa6_0),.dout(w_dff_B_GaY4qt4a6_0),.clk(gclk));
	jdff dff_B_K3pQ5h3w7_0(.din(w_dff_B_GaY4qt4a6_0),.dout(w_dff_B_K3pQ5h3w7_0),.clk(gclk));
	jdff dff_B_qo3EOGlQ0_0(.din(w_dff_B_K3pQ5h3w7_0),.dout(w_dff_B_qo3EOGlQ0_0),.clk(gclk));
	jdff dff_B_kMkBYx3G0_0(.din(w_dff_B_qo3EOGlQ0_0),.dout(w_dff_B_kMkBYx3G0_0),.clk(gclk));
	jdff dff_B_3D7PmEZW1_0(.din(w_dff_B_kMkBYx3G0_0),.dout(w_dff_B_3D7PmEZW1_0),.clk(gclk));
	jdff dff_B_FRZFB3478_0(.din(w_dff_B_3D7PmEZW1_0),.dout(w_dff_B_FRZFB3478_0),.clk(gclk));
	jdff dff_B_vlaHuW2B7_0(.din(w_dff_B_FRZFB3478_0),.dout(w_dff_B_vlaHuW2B7_0),.clk(gclk));
	jdff dff_B_Gf76VPPs4_0(.din(w_dff_B_vlaHuW2B7_0),.dout(w_dff_B_Gf76VPPs4_0),.clk(gclk));
	jdff dff_B_BZFvn93D9_0(.din(w_dff_B_Gf76VPPs4_0),.dout(w_dff_B_BZFvn93D9_0),.clk(gclk));
	jdff dff_B_fLKBBBCo5_0(.din(w_dff_B_BZFvn93D9_0),.dout(w_dff_B_fLKBBBCo5_0),.clk(gclk));
	jdff dff_B_cjnZ9Qlu7_0(.din(w_dff_B_fLKBBBCo5_0),.dout(w_dff_B_cjnZ9Qlu7_0),.clk(gclk));
	jdff dff_B_0qILxkjt9_0(.din(w_dff_B_cjnZ9Qlu7_0),.dout(w_dff_B_0qILxkjt9_0),.clk(gclk));
	jdff dff_B_FVAxEKMA6_0(.din(w_dff_B_0qILxkjt9_0),.dout(w_dff_B_FVAxEKMA6_0),.clk(gclk));
	jdff dff_B_ER3waTSn2_0(.din(w_dff_B_FVAxEKMA6_0),.dout(w_dff_B_ER3waTSn2_0),.clk(gclk));
	jdff dff_B_tjAPeAJ01_0(.din(w_dff_B_ER3waTSn2_0),.dout(w_dff_B_tjAPeAJ01_0),.clk(gclk));
	jdff dff_B_na8ylLxA0_0(.din(w_dff_B_tjAPeAJ01_0),.dout(w_dff_B_na8ylLxA0_0),.clk(gclk));
	jdff dff_B_fQentjdi1_0(.din(w_dff_B_na8ylLxA0_0),.dout(w_dff_B_fQentjdi1_0),.clk(gclk));
	jdff dff_B_LPOgw3ob1_0(.din(w_dff_B_fQentjdi1_0),.dout(w_dff_B_LPOgw3ob1_0),.clk(gclk));
	jdff dff_B_1xwZuAru7_0(.din(w_dff_B_LPOgw3ob1_0),.dout(w_dff_B_1xwZuAru7_0),.clk(gclk));
	jdff dff_B_rLkqJbTJ8_0(.din(w_dff_B_1xwZuAru7_0),.dout(w_dff_B_rLkqJbTJ8_0),.clk(gclk));
	jdff dff_B_4EazO7Zy9_0(.din(w_dff_B_rLkqJbTJ8_0),.dout(w_dff_B_4EazO7Zy9_0),.clk(gclk));
	jdff dff_B_8qdQpabr3_0(.din(w_dff_B_4EazO7Zy9_0),.dout(w_dff_B_8qdQpabr3_0),.clk(gclk));
	jdff dff_B_UWt7o4dv5_0(.din(w_dff_B_8qdQpabr3_0),.dout(w_dff_B_UWt7o4dv5_0),.clk(gclk));
	jdff dff_B_eaMsKA4H0_0(.din(w_dff_B_UWt7o4dv5_0),.dout(w_dff_B_eaMsKA4H0_0),.clk(gclk));
	jdff dff_B_h4aUYj344_0(.din(w_dff_B_eaMsKA4H0_0),.dout(w_dff_B_h4aUYj344_0),.clk(gclk));
	jdff dff_B_oaTA7AA74_0(.din(w_dff_B_h4aUYj344_0),.dout(w_dff_B_oaTA7AA74_0),.clk(gclk));
	jdff dff_B_AtWNkgKv1_0(.din(w_dff_B_oaTA7AA74_0),.dout(w_dff_B_AtWNkgKv1_0),.clk(gclk));
	jdff dff_B_k6zCwV8k1_0(.din(w_dff_B_AtWNkgKv1_0),.dout(w_dff_B_k6zCwV8k1_0),.clk(gclk));
	jdff dff_B_O1KolSyU1_0(.din(w_dff_B_k6zCwV8k1_0),.dout(w_dff_B_O1KolSyU1_0),.clk(gclk));
	jdff dff_B_3FVBTjde4_0(.din(w_dff_B_O1KolSyU1_0),.dout(w_dff_B_3FVBTjde4_0),.clk(gclk));
	jdff dff_B_Nn2pDx1S4_0(.din(w_dff_B_3FVBTjde4_0),.dout(w_dff_B_Nn2pDx1S4_0),.clk(gclk));
	jdff dff_B_jX7DVGGu5_0(.din(w_dff_B_Nn2pDx1S4_0),.dout(w_dff_B_jX7DVGGu5_0),.clk(gclk));
	jdff dff_B_XeWl1wDu0_0(.din(w_dff_B_jX7DVGGu5_0),.dout(w_dff_B_XeWl1wDu0_0),.clk(gclk));
	jdff dff_B_vQLxsDKn6_0(.din(w_dff_B_XeWl1wDu0_0),.dout(w_dff_B_vQLxsDKn6_0),.clk(gclk));
	jdff dff_B_txjZgmlX0_0(.din(w_dff_B_vQLxsDKn6_0),.dout(w_dff_B_txjZgmlX0_0),.clk(gclk));
	jdff dff_B_NYNGcIk41_0(.din(w_dff_B_txjZgmlX0_0),.dout(w_dff_B_NYNGcIk41_0),.clk(gclk));
	jdff dff_B_n1rpOmAn9_0(.din(w_dff_B_NYNGcIk41_0),.dout(w_dff_B_n1rpOmAn9_0),.clk(gclk));
	jdff dff_B_NIhTncFp9_0(.din(n730),.dout(w_dff_B_NIhTncFp9_0),.clk(gclk));
	jdff dff_B_HdqDu6U36_0(.din(w_dff_B_NIhTncFp9_0),.dout(w_dff_B_HdqDu6U36_0),.clk(gclk));
	jdff dff_B_RHJZsHOH9_0(.din(w_dff_B_HdqDu6U36_0),.dout(w_dff_B_RHJZsHOH9_0),.clk(gclk));
	jdff dff_B_pMSCIz955_0(.din(w_dff_B_RHJZsHOH9_0),.dout(w_dff_B_pMSCIz955_0),.clk(gclk));
	jdff dff_B_My4ZOapN3_0(.din(w_dff_B_pMSCIz955_0),.dout(w_dff_B_My4ZOapN3_0),.clk(gclk));
	jdff dff_B_gq6333Mh8_0(.din(w_dff_B_My4ZOapN3_0),.dout(w_dff_B_gq6333Mh8_0),.clk(gclk));
	jdff dff_B_ukokP1Kv3_0(.din(w_dff_B_gq6333Mh8_0),.dout(w_dff_B_ukokP1Kv3_0),.clk(gclk));
	jdff dff_B_BXBwBDdk0_0(.din(w_dff_B_ukokP1Kv3_0),.dout(w_dff_B_BXBwBDdk0_0),.clk(gclk));
	jdff dff_B_sNvwIeOx5_0(.din(w_dff_B_BXBwBDdk0_0),.dout(w_dff_B_sNvwIeOx5_0),.clk(gclk));
	jdff dff_B_OcZ9YFZp5_0(.din(w_dff_B_sNvwIeOx5_0),.dout(w_dff_B_OcZ9YFZp5_0),.clk(gclk));
	jdff dff_B_MJS4mRfO8_0(.din(w_dff_B_OcZ9YFZp5_0),.dout(w_dff_B_MJS4mRfO8_0),.clk(gclk));
	jdff dff_B_MujxiHya4_0(.din(w_dff_B_MJS4mRfO8_0),.dout(w_dff_B_MujxiHya4_0),.clk(gclk));
	jdff dff_B_yhksFV181_0(.din(w_dff_B_MujxiHya4_0),.dout(w_dff_B_yhksFV181_0),.clk(gclk));
	jdff dff_B_kyv3tfV22_0(.din(w_dff_B_yhksFV181_0),.dout(w_dff_B_kyv3tfV22_0),.clk(gclk));
	jdff dff_B_nP6cZpCl4_0(.din(w_dff_B_kyv3tfV22_0),.dout(w_dff_B_nP6cZpCl4_0),.clk(gclk));
	jdff dff_B_l9xN2bV80_0(.din(w_dff_B_nP6cZpCl4_0),.dout(w_dff_B_l9xN2bV80_0),.clk(gclk));
	jdff dff_B_Q7GsqJgO9_0(.din(w_dff_B_l9xN2bV80_0),.dout(w_dff_B_Q7GsqJgO9_0),.clk(gclk));
	jdff dff_B_Gy8x11xb5_0(.din(w_dff_B_Q7GsqJgO9_0),.dout(w_dff_B_Gy8x11xb5_0),.clk(gclk));
	jdff dff_B_akCtNz9q8_0(.din(w_dff_B_Gy8x11xb5_0),.dout(w_dff_B_akCtNz9q8_0),.clk(gclk));
	jdff dff_B_7bacJMT45_0(.din(w_dff_B_akCtNz9q8_0),.dout(w_dff_B_7bacJMT45_0),.clk(gclk));
	jdff dff_B_Mu7xJ6494_0(.din(w_dff_B_7bacJMT45_0),.dout(w_dff_B_Mu7xJ6494_0),.clk(gclk));
	jdff dff_B_aiQujMYy4_0(.din(w_dff_B_Mu7xJ6494_0),.dout(w_dff_B_aiQujMYy4_0),.clk(gclk));
	jdff dff_B_V54ZLEyd6_0(.din(w_dff_B_aiQujMYy4_0),.dout(w_dff_B_V54ZLEyd6_0),.clk(gclk));
	jdff dff_B_OpDFoOTy1_0(.din(w_dff_B_V54ZLEyd6_0),.dout(w_dff_B_OpDFoOTy1_0),.clk(gclk));
	jdff dff_B_XJOIHvXK3_0(.din(w_dff_B_OpDFoOTy1_0),.dout(w_dff_B_XJOIHvXK3_0),.clk(gclk));
	jdff dff_B_cDh3cUFn2_0(.din(w_dff_B_XJOIHvXK3_0),.dout(w_dff_B_cDh3cUFn2_0),.clk(gclk));
	jdff dff_B_CWU2bbfI4_0(.din(w_dff_B_cDh3cUFn2_0),.dout(w_dff_B_CWU2bbfI4_0),.clk(gclk));
	jdff dff_B_k043bbsw9_0(.din(w_dff_B_CWU2bbfI4_0),.dout(w_dff_B_k043bbsw9_0),.clk(gclk));
	jdff dff_B_UPHwnOKn9_0(.din(w_dff_B_k043bbsw9_0),.dout(w_dff_B_UPHwnOKn9_0),.clk(gclk));
	jdff dff_B_Ursiat8U0_0(.din(w_dff_B_UPHwnOKn9_0),.dout(w_dff_B_Ursiat8U0_0),.clk(gclk));
	jdff dff_B_WenzMoZn5_0(.din(w_dff_B_Ursiat8U0_0),.dout(w_dff_B_WenzMoZn5_0),.clk(gclk));
	jdff dff_B_Pedb5i9v1_0(.din(w_dff_B_WenzMoZn5_0),.dout(w_dff_B_Pedb5i9v1_0),.clk(gclk));
	jdff dff_B_eGWiGWuv9_0(.din(w_dff_B_Pedb5i9v1_0),.dout(w_dff_B_eGWiGWuv9_0),.clk(gclk));
	jdff dff_B_Z6tMjP6B4_0(.din(w_dff_B_eGWiGWuv9_0),.dout(w_dff_B_Z6tMjP6B4_0),.clk(gclk));
	jdff dff_B_hdhHwUwg1_0(.din(w_dff_B_Z6tMjP6B4_0),.dout(w_dff_B_hdhHwUwg1_0),.clk(gclk));
	jdff dff_B_G6vSpW5m7_0(.din(w_dff_B_hdhHwUwg1_0),.dout(w_dff_B_G6vSpW5m7_0),.clk(gclk));
	jdff dff_B_xhUP7fvG0_0(.din(w_dff_B_G6vSpW5m7_0),.dout(w_dff_B_xhUP7fvG0_0),.clk(gclk));
	jdff dff_B_ICyfZ5Ai3_0(.din(w_dff_B_xhUP7fvG0_0),.dout(w_dff_B_ICyfZ5Ai3_0),.clk(gclk));
	jdff dff_B_5y4jQn4h6_0(.din(w_dff_B_ICyfZ5Ai3_0),.dout(w_dff_B_5y4jQn4h6_0),.clk(gclk));
	jdff dff_B_fPCg0bHC7_0(.din(w_dff_B_5y4jQn4h6_0),.dout(w_dff_B_fPCg0bHC7_0),.clk(gclk));
	jdff dff_B_a656EM6I6_0(.din(w_dff_B_fPCg0bHC7_0),.dout(w_dff_B_a656EM6I6_0),.clk(gclk));
	jdff dff_B_EKqKVKYc2_0(.din(w_dff_B_a656EM6I6_0),.dout(w_dff_B_EKqKVKYc2_0),.clk(gclk));
	jdff dff_B_UWRk1O027_0(.din(w_dff_B_EKqKVKYc2_0),.dout(w_dff_B_UWRk1O027_0),.clk(gclk));
	jdff dff_B_N7DmpM2p4_0(.din(w_dff_B_UWRk1O027_0),.dout(w_dff_B_N7DmpM2p4_0),.clk(gclk));
	jdff dff_B_xN4GSsOI9_0(.din(w_dff_B_N7DmpM2p4_0),.dout(w_dff_B_xN4GSsOI9_0),.clk(gclk));
	jdff dff_B_gOmI6URF1_0(.din(w_dff_B_xN4GSsOI9_0),.dout(w_dff_B_gOmI6URF1_0),.clk(gclk));
	jdff dff_B_03uW9gTi8_0(.din(w_dff_B_gOmI6URF1_0),.dout(w_dff_B_03uW9gTi8_0),.clk(gclk));
	jdff dff_B_nqObvXTJ0_0(.din(w_dff_B_03uW9gTi8_0),.dout(w_dff_B_nqObvXTJ0_0),.clk(gclk));
	jdff dff_B_qFUYtomk5_0(.din(w_dff_B_nqObvXTJ0_0),.dout(w_dff_B_qFUYtomk5_0),.clk(gclk));
	jdff dff_B_myLaGLRL4_0(.din(w_dff_B_qFUYtomk5_0),.dout(w_dff_B_myLaGLRL4_0),.clk(gclk));
	jdff dff_B_Hdw3qxMg6_0(.din(w_dff_B_myLaGLRL4_0),.dout(w_dff_B_Hdw3qxMg6_0),.clk(gclk));
	jdff dff_B_TpAwsMsu0_0(.din(w_dff_B_Hdw3qxMg6_0),.dout(w_dff_B_TpAwsMsu0_0),.clk(gclk));
	jdff dff_B_ZhA7BnFW3_0(.din(w_dff_B_TpAwsMsu0_0),.dout(w_dff_B_ZhA7BnFW3_0),.clk(gclk));
	jdff dff_B_hL1I0h6t8_0(.din(w_dff_B_ZhA7BnFW3_0),.dout(w_dff_B_hL1I0h6t8_0),.clk(gclk));
	jdff dff_B_2xYT2Nog2_0(.din(w_dff_B_hL1I0h6t8_0),.dout(w_dff_B_2xYT2Nog2_0),.clk(gclk));
	jdff dff_B_YiiTRArl1_0(.din(w_dff_B_2xYT2Nog2_0),.dout(w_dff_B_YiiTRArl1_0),.clk(gclk));
	jdff dff_B_GE2mGqKL5_0(.din(w_dff_B_YiiTRArl1_0),.dout(w_dff_B_GE2mGqKL5_0),.clk(gclk));
	jdff dff_B_chPYLgF62_0(.din(n736),.dout(w_dff_B_chPYLgF62_0),.clk(gclk));
	jdff dff_B_T2jR5Ota3_0(.din(w_dff_B_chPYLgF62_0),.dout(w_dff_B_T2jR5Ota3_0),.clk(gclk));
	jdff dff_B_jK2apygH2_0(.din(w_dff_B_T2jR5Ota3_0),.dout(w_dff_B_jK2apygH2_0),.clk(gclk));
	jdff dff_B_VBJFopmb1_0(.din(w_dff_B_jK2apygH2_0),.dout(w_dff_B_VBJFopmb1_0),.clk(gclk));
	jdff dff_B_KAGUHmsE6_0(.din(w_dff_B_VBJFopmb1_0),.dout(w_dff_B_KAGUHmsE6_0),.clk(gclk));
	jdff dff_B_qPCq6zoJ0_0(.din(w_dff_B_KAGUHmsE6_0),.dout(w_dff_B_qPCq6zoJ0_0),.clk(gclk));
	jdff dff_B_dvXCZErz5_0(.din(w_dff_B_qPCq6zoJ0_0),.dout(w_dff_B_dvXCZErz5_0),.clk(gclk));
	jdff dff_B_bNn9kino5_0(.din(w_dff_B_dvXCZErz5_0),.dout(w_dff_B_bNn9kino5_0),.clk(gclk));
	jdff dff_B_4AzEzqTM6_0(.din(w_dff_B_bNn9kino5_0),.dout(w_dff_B_4AzEzqTM6_0),.clk(gclk));
	jdff dff_B_xZm2pGyh8_0(.din(w_dff_B_4AzEzqTM6_0),.dout(w_dff_B_xZm2pGyh8_0),.clk(gclk));
	jdff dff_B_zUUlLEYb7_0(.din(w_dff_B_xZm2pGyh8_0),.dout(w_dff_B_zUUlLEYb7_0),.clk(gclk));
	jdff dff_B_sxSxIZwr7_0(.din(w_dff_B_zUUlLEYb7_0),.dout(w_dff_B_sxSxIZwr7_0),.clk(gclk));
	jdff dff_B_cV0tdWP02_0(.din(w_dff_B_sxSxIZwr7_0),.dout(w_dff_B_cV0tdWP02_0),.clk(gclk));
	jdff dff_B_GoozpgYI0_0(.din(w_dff_B_cV0tdWP02_0),.dout(w_dff_B_GoozpgYI0_0),.clk(gclk));
	jdff dff_B_irIfkTAY9_0(.din(w_dff_B_GoozpgYI0_0),.dout(w_dff_B_irIfkTAY9_0),.clk(gclk));
	jdff dff_B_cRRE6kJz0_0(.din(w_dff_B_irIfkTAY9_0),.dout(w_dff_B_cRRE6kJz0_0),.clk(gclk));
	jdff dff_B_S0hdnirW3_0(.din(w_dff_B_cRRE6kJz0_0),.dout(w_dff_B_S0hdnirW3_0),.clk(gclk));
	jdff dff_B_AtBCkKkY5_0(.din(w_dff_B_S0hdnirW3_0),.dout(w_dff_B_AtBCkKkY5_0),.clk(gclk));
	jdff dff_B_uOxYj7qZ1_0(.din(w_dff_B_AtBCkKkY5_0),.dout(w_dff_B_uOxYj7qZ1_0),.clk(gclk));
	jdff dff_B_U4P79lTw3_0(.din(w_dff_B_uOxYj7qZ1_0),.dout(w_dff_B_U4P79lTw3_0),.clk(gclk));
	jdff dff_B_poqdFB3x7_0(.din(w_dff_B_U4P79lTw3_0),.dout(w_dff_B_poqdFB3x7_0),.clk(gclk));
	jdff dff_B_4vnyuzy01_0(.din(w_dff_B_poqdFB3x7_0),.dout(w_dff_B_4vnyuzy01_0),.clk(gclk));
	jdff dff_B_VuM2OjLO4_0(.din(w_dff_B_4vnyuzy01_0),.dout(w_dff_B_VuM2OjLO4_0),.clk(gclk));
	jdff dff_B_oYUeOmx77_0(.din(w_dff_B_VuM2OjLO4_0),.dout(w_dff_B_oYUeOmx77_0),.clk(gclk));
	jdff dff_B_uU8kckxO3_0(.din(w_dff_B_oYUeOmx77_0),.dout(w_dff_B_uU8kckxO3_0),.clk(gclk));
	jdff dff_B_mxiamplP9_0(.din(w_dff_B_uU8kckxO3_0),.dout(w_dff_B_mxiamplP9_0),.clk(gclk));
	jdff dff_B_leaqwRHk4_0(.din(w_dff_B_mxiamplP9_0),.dout(w_dff_B_leaqwRHk4_0),.clk(gclk));
	jdff dff_B_cZJonqiL8_0(.din(w_dff_B_leaqwRHk4_0),.dout(w_dff_B_cZJonqiL8_0),.clk(gclk));
	jdff dff_B_659s3U2q7_0(.din(w_dff_B_cZJonqiL8_0),.dout(w_dff_B_659s3U2q7_0),.clk(gclk));
	jdff dff_B_9YaPMIhN0_0(.din(w_dff_B_659s3U2q7_0),.dout(w_dff_B_9YaPMIhN0_0),.clk(gclk));
	jdff dff_B_uMjB28FB9_0(.din(w_dff_B_9YaPMIhN0_0),.dout(w_dff_B_uMjB28FB9_0),.clk(gclk));
	jdff dff_B_GG5sD3FW6_0(.din(w_dff_B_uMjB28FB9_0),.dout(w_dff_B_GG5sD3FW6_0),.clk(gclk));
	jdff dff_B_f08spvnV0_0(.din(w_dff_B_GG5sD3FW6_0),.dout(w_dff_B_f08spvnV0_0),.clk(gclk));
	jdff dff_B_Rc1sRFHO8_0(.din(w_dff_B_f08spvnV0_0),.dout(w_dff_B_Rc1sRFHO8_0),.clk(gclk));
	jdff dff_B_ZAgPOUSz7_0(.din(w_dff_B_Rc1sRFHO8_0),.dout(w_dff_B_ZAgPOUSz7_0),.clk(gclk));
	jdff dff_B_WRuwlgAp9_0(.din(w_dff_B_ZAgPOUSz7_0),.dout(w_dff_B_WRuwlgAp9_0),.clk(gclk));
	jdff dff_B_pTDgQpyy0_0(.din(w_dff_B_WRuwlgAp9_0),.dout(w_dff_B_pTDgQpyy0_0),.clk(gclk));
	jdff dff_B_ZEx5grzP6_0(.din(w_dff_B_pTDgQpyy0_0),.dout(w_dff_B_ZEx5grzP6_0),.clk(gclk));
	jdff dff_B_WetPrXur0_0(.din(w_dff_B_ZEx5grzP6_0),.dout(w_dff_B_WetPrXur0_0),.clk(gclk));
	jdff dff_B_tG8aemG22_0(.din(w_dff_B_WetPrXur0_0),.dout(w_dff_B_tG8aemG22_0),.clk(gclk));
	jdff dff_B_lM0srbnz1_0(.din(w_dff_B_tG8aemG22_0),.dout(w_dff_B_lM0srbnz1_0),.clk(gclk));
	jdff dff_B_c8cb8YR29_0(.din(w_dff_B_lM0srbnz1_0),.dout(w_dff_B_c8cb8YR29_0),.clk(gclk));
	jdff dff_B_QL4QL1ok3_0(.din(w_dff_B_c8cb8YR29_0),.dout(w_dff_B_QL4QL1ok3_0),.clk(gclk));
	jdff dff_B_OvwJsaxy3_0(.din(w_dff_B_QL4QL1ok3_0),.dout(w_dff_B_OvwJsaxy3_0),.clk(gclk));
	jdff dff_B_qkyB8GPw3_0(.din(w_dff_B_OvwJsaxy3_0),.dout(w_dff_B_qkyB8GPw3_0),.clk(gclk));
	jdff dff_B_gcyrlYWI8_0(.din(w_dff_B_qkyB8GPw3_0),.dout(w_dff_B_gcyrlYWI8_0),.clk(gclk));
	jdff dff_B_utaX2tZo7_0(.din(w_dff_B_gcyrlYWI8_0),.dout(w_dff_B_utaX2tZo7_0),.clk(gclk));
	jdff dff_B_3PY73daK5_0(.din(w_dff_B_utaX2tZo7_0),.dout(w_dff_B_3PY73daK5_0),.clk(gclk));
	jdff dff_B_dtl0pjpD9_0(.din(w_dff_B_3PY73daK5_0),.dout(w_dff_B_dtl0pjpD9_0),.clk(gclk));
	jdff dff_B_wGd6jGjQ2_0(.din(w_dff_B_dtl0pjpD9_0),.dout(w_dff_B_wGd6jGjQ2_0),.clk(gclk));
	jdff dff_B_W5O1D9Sp9_0(.din(w_dff_B_wGd6jGjQ2_0),.dout(w_dff_B_W5O1D9Sp9_0),.clk(gclk));
	jdff dff_B_FBhFPXnx9_0(.din(w_dff_B_W5O1D9Sp9_0),.dout(w_dff_B_FBhFPXnx9_0),.clk(gclk));
	jdff dff_B_oc2VA5YM2_0(.din(w_dff_B_FBhFPXnx9_0),.dout(w_dff_B_oc2VA5YM2_0),.clk(gclk));
	jdff dff_B_EYo8R46K4_0(.din(w_dff_B_oc2VA5YM2_0),.dout(w_dff_B_EYo8R46K4_0),.clk(gclk));
	jdff dff_B_jrRbyq497_0(.din(w_dff_B_EYo8R46K4_0),.dout(w_dff_B_jrRbyq497_0),.clk(gclk));
	jdff dff_B_WiwTm3sF9_0(.din(w_dff_B_jrRbyq497_0),.dout(w_dff_B_WiwTm3sF9_0),.clk(gclk));
	jdff dff_B_98Tylq7e8_0(.din(w_dff_B_WiwTm3sF9_0),.dout(w_dff_B_98Tylq7e8_0),.clk(gclk));
	jdff dff_B_UNX9CF5n9_0(.din(w_dff_B_98Tylq7e8_0),.dout(w_dff_B_UNX9CF5n9_0),.clk(gclk));
	jdff dff_B_wmuF7Gyw8_0(.din(n742),.dout(w_dff_B_wmuF7Gyw8_0),.clk(gclk));
	jdff dff_B_ixXLIgpD9_0(.din(w_dff_B_wmuF7Gyw8_0),.dout(w_dff_B_ixXLIgpD9_0),.clk(gclk));
	jdff dff_B_RwcTgqMI0_0(.din(w_dff_B_ixXLIgpD9_0),.dout(w_dff_B_RwcTgqMI0_0),.clk(gclk));
	jdff dff_B_oYhZq91j9_0(.din(w_dff_B_RwcTgqMI0_0),.dout(w_dff_B_oYhZq91j9_0),.clk(gclk));
	jdff dff_B_jg73UTkb8_0(.din(w_dff_B_oYhZq91j9_0),.dout(w_dff_B_jg73UTkb8_0),.clk(gclk));
	jdff dff_B_U6YufzZX2_0(.din(w_dff_B_jg73UTkb8_0),.dout(w_dff_B_U6YufzZX2_0),.clk(gclk));
	jdff dff_B_LGLrxn9n8_0(.din(w_dff_B_U6YufzZX2_0),.dout(w_dff_B_LGLrxn9n8_0),.clk(gclk));
	jdff dff_B_nzVGwEhw3_0(.din(w_dff_B_LGLrxn9n8_0),.dout(w_dff_B_nzVGwEhw3_0),.clk(gclk));
	jdff dff_B_UsWbYh5u8_0(.din(w_dff_B_nzVGwEhw3_0),.dout(w_dff_B_UsWbYh5u8_0),.clk(gclk));
	jdff dff_B_mw3sseZp8_0(.din(w_dff_B_UsWbYh5u8_0),.dout(w_dff_B_mw3sseZp8_0),.clk(gclk));
	jdff dff_B_6NZl6yYS6_0(.din(w_dff_B_mw3sseZp8_0),.dout(w_dff_B_6NZl6yYS6_0),.clk(gclk));
	jdff dff_B_3gHD8I003_0(.din(w_dff_B_6NZl6yYS6_0),.dout(w_dff_B_3gHD8I003_0),.clk(gclk));
	jdff dff_B_9MSeXjVk6_0(.din(w_dff_B_3gHD8I003_0),.dout(w_dff_B_9MSeXjVk6_0),.clk(gclk));
	jdff dff_B_USJUgjM55_0(.din(w_dff_B_9MSeXjVk6_0),.dout(w_dff_B_USJUgjM55_0),.clk(gclk));
	jdff dff_B_CyOuxERh9_0(.din(w_dff_B_USJUgjM55_0),.dout(w_dff_B_CyOuxERh9_0),.clk(gclk));
	jdff dff_B_V7Ib9fpJ1_0(.din(w_dff_B_CyOuxERh9_0),.dout(w_dff_B_V7Ib9fpJ1_0),.clk(gclk));
	jdff dff_B_UNnD9opa5_0(.din(w_dff_B_V7Ib9fpJ1_0),.dout(w_dff_B_UNnD9opa5_0),.clk(gclk));
	jdff dff_B_w4hhfaAA3_0(.din(w_dff_B_UNnD9opa5_0),.dout(w_dff_B_w4hhfaAA3_0),.clk(gclk));
	jdff dff_B_RfnKpmUW5_0(.din(w_dff_B_w4hhfaAA3_0),.dout(w_dff_B_RfnKpmUW5_0),.clk(gclk));
	jdff dff_B_QFngED6z3_0(.din(w_dff_B_RfnKpmUW5_0),.dout(w_dff_B_QFngED6z3_0),.clk(gclk));
	jdff dff_B_zhUwLWLv2_0(.din(w_dff_B_QFngED6z3_0),.dout(w_dff_B_zhUwLWLv2_0),.clk(gclk));
	jdff dff_B_js52DzsR9_0(.din(w_dff_B_zhUwLWLv2_0),.dout(w_dff_B_js52DzsR9_0),.clk(gclk));
	jdff dff_B_cQv8lHFu4_0(.din(w_dff_B_js52DzsR9_0),.dout(w_dff_B_cQv8lHFu4_0),.clk(gclk));
	jdff dff_B_ASAy6Jg10_0(.din(w_dff_B_cQv8lHFu4_0),.dout(w_dff_B_ASAy6Jg10_0),.clk(gclk));
	jdff dff_B_fV5OmoIN2_0(.din(w_dff_B_ASAy6Jg10_0),.dout(w_dff_B_fV5OmoIN2_0),.clk(gclk));
	jdff dff_B_UTK9vC4t4_0(.din(w_dff_B_fV5OmoIN2_0),.dout(w_dff_B_UTK9vC4t4_0),.clk(gclk));
	jdff dff_B_U7zIeVLj4_0(.din(w_dff_B_UTK9vC4t4_0),.dout(w_dff_B_U7zIeVLj4_0),.clk(gclk));
	jdff dff_B_mdYh0M4r5_0(.din(w_dff_B_U7zIeVLj4_0),.dout(w_dff_B_mdYh0M4r5_0),.clk(gclk));
	jdff dff_B_PgRhADgl6_0(.din(w_dff_B_mdYh0M4r5_0),.dout(w_dff_B_PgRhADgl6_0),.clk(gclk));
	jdff dff_B_ul48SBz97_0(.din(w_dff_B_PgRhADgl6_0),.dout(w_dff_B_ul48SBz97_0),.clk(gclk));
	jdff dff_B_9p7xzlIp3_0(.din(w_dff_B_ul48SBz97_0),.dout(w_dff_B_9p7xzlIp3_0),.clk(gclk));
	jdff dff_B_CdeWzgM28_0(.din(w_dff_B_9p7xzlIp3_0),.dout(w_dff_B_CdeWzgM28_0),.clk(gclk));
	jdff dff_B_5yBunGSQ8_0(.din(w_dff_B_CdeWzgM28_0),.dout(w_dff_B_5yBunGSQ8_0),.clk(gclk));
	jdff dff_B_x0WdS5e65_0(.din(w_dff_B_5yBunGSQ8_0),.dout(w_dff_B_x0WdS5e65_0),.clk(gclk));
	jdff dff_B_ZpqICiyX9_0(.din(w_dff_B_x0WdS5e65_0),.dout(w_dff_B_ZpqICiyX9_0),.clk(gclk));
	jdff dff_B_otsDwvqB3_0(.din(w_dff_B_ZpqICiyX9_0),.dout(w_dff_B_otsDwvqB3_0),.clk(gclk));
	jdff dff_B_eMqcbWqV4_0(.din(w_dff_B_otsDwvqB3_0),.dout(w_dff_B_eMqcbWqV4_0),.clk(gclk));
	jdff dff_B_BnpiaI0O1_0(.din(w_dff_B_eMqcbWqV4_0),.dout(w_dff_B_BnpiaI0O1_0),.clk(gclk));
	jdff dff_B_FInMvcY67_0(.din(w_dff_B_BnpiaI0O1_0),.dout(w_dff_B_FInMvcY67_0),.clk(gclk));
	jdff dff_B_KQX3qftb1_0(.din(w_dff_B_FInMvcY67_0),.dout(w_dff_B_KQX3qftb1_0),.clk(gclk));
	jdff dff_B_wR3EJoxe7_0(.din(w_dff_B_KQX3qftb1_0),.dout(w_dff_B_wR3EJoxe7_0),.clk(gclk));
	jdff dff_B_57uY1CXv3_0(.din(w_dff_B_wR3EJoxe7_0),.dout(w_dff_B_57uY1CXv3_0),.clk(gclk));
	jdff dff_B_1HRlSZAR2_0(.din(w_dff_B_57uY1CXv3_0),.dout(w_dff_B_1HRlSZAR2_0),.clk(gclk));
	jdff dff_B_xnyzMUxu5_0(.din(w_dff_B_1HRlSZAR2_0),.dout(w_dff_B_xnyzMUxu5_0),.clk(gclk));
	jdff dff_B_8ubBVz866_0(.din(w_dff_B_xnyzMUxu5_0),.dout(w_dff_B_8ubBVz866_0),.clk(gclk));
	jdff dff_B_9EJx8tWJ3_0(.din(w_dff_B_8ubBVz866_0),.dout(w_dff_B_9EJx8tWJ3_0),.clk(gclk));
	jdff dff_B_yjHX2iy78_0(.din(w_dff_B_9EJx8tWJ3_0),.dout(w_dff_B_yjHX2iy78_0),.clk(gclk));
	jdff dff_B_GDzeQc6Q8_0(.din(w_dff_B_yjHX2iy78_0),.dout(w_dff_B_GDzeQc6Q8_0),.clk(gclk));
	jdff dff_B_fUrlSf5P4_0(.din(w_dff_B_GDzeQc6Q8_0),.dout(w_dff_B_fUrlSf5P4_0),.clk(gclk));
	jdff dff_B_ossniog09_0(.din(w_dff_B_fUrlSf5P4_0),.dout(w_dff_B_ossniog09_0),.clk(gclk));
	jdff dff_B_7UWCIscI1_0(.din(w_dff_B_ossniog09_0),.dout(w_dff_B_7UWCIscI1_0),.clk(gclk));
	jdff dff_B_TYPlv2uD4_0(.din(w_dff_B_7UWCIscI1_0),.dout(w_dff_B_TYPlv2uD4_0),.clk(gclk));
	jdff dff_B_X86le55n6_0(.din(w_dff_B_TYPlv2uD4_0),.dout(w_dff_B_X86le55n6_0),.clk(gclk));
	jdff dff_B_DAC1g3TT6_0(.din(w_dff_B_X86le55n6_0),.dout(w_dff_B_DAC1g3TT6_0),.clk(gclk));
	jdff dff_B_ZXJBwqzf4_0(.din(w_dff_B_DAC1g3TT6_0),.dout(w_dff_B_ZXJBwqzf4_0),.clk(gclk));
	jdff dff_B_gWGVgIsu2_0(.din(w_dff_B_ZXJBwqzf4_0),.dout(w_dff_B_gWGVgIsu2_0),.clk(gclk));
	jdff dff_B_EHBKLGB74_0(.din(w_dff_B_gWGVgIsu2_0),.dout(w_dff_B_EHBKLGB74_0),.clk(gclk));
	jdff dff_B_SrGuoJOq9_0(.din(w_dff_B_EHBKLGB74_0),.dout(w_dff_B_SrGuoJOq9_0),.clk(gclk));
	jdff dff_B_2Kzh4c4E2_0(.din(w_dff_B_SrGuoJOq9_0),.dout(w_dff_B_2Kzh4c4E2_0),.clk(gclk));
	jdff dff_B_IS5Skb8y1_0(.din(n748),.dout(w_dff_B_IS5Skb8y1_0),.clk(gclk));
	jdff dff_B_ysJOZP5q0_0(.din(w_dff_B_IS5Skb8y1_0),.dout(w_dff_B_ysJOZP5q0_0),.clk(gclk));
	jdff dff_B_YbdqseU76_0(.din(w_dff_B_ysJOZP5q0_0),.dout(w_dff_B_YbdqseU76_0),.clk(gclk));
	jdff dff_B_gZ8DvZdn8_0(.din(w_dff_B_YbdqseU76_0),.dout(w_dff_B_gZ8DvZdn8_0),.clk(gclk));
	jdff dff_B_uxmgcEOt7_0(.din(w_dff_B_gZ8DvZdn8_0),.dout(w_dff_B_uxmgcEOt7_0),.clk(gclk));
	jdff dff_B_qEeD1Y121_0(.din(w_dff_B_uxmgcEOt7_0),.dout(w_dff_B_qEeD1Y121_0),.clk(gclk));
	jdff dff_B_tGyFtL8g5_0(.din(w_dff_B_qEeD1Y121_0),.dout(w_dff_B_tGyFtL8g5_0),.clk(gclk));
	jdff dff_B_ZMVjOfh13_0(.din(w_dff_B_tGyFtL8g5_0),.dout(w_dff_B_ZMVjOfh13_0),.clk(gclk));
	jdff dff_B_Yjq2hmXF0_0(.din(w_dff_B_ZMVjOfh13_0),.dout(w_dff_B_Yjq2hmXF0_0),.clk(gclk));
	jdff dff_B_WieN8Xbb0_0(.din(w_dff_B_Yjq2hmXF0_0),.dout(w_dff_B_WieN8Xbb0_0),.clk(gclk));
	jdff dff_B_HBpI1Stx1_0(.din(w_dff_B_WieN8Xbb0_0),.dout(w_dff_B_HBpI1Stx1_0),.clk(gclk));
	jdff dff_B_RnB35QRk1_0(.din(w_dff_B_HBpI1Stx1_0),.dout(w_dff_B_RnB35QRk1_0),.clk(gclk));
	jdff dff_B_mPn94spR7_0(.din(w_dff_B_RnB35QRk1_0),.dout(w_dff_B_mPn94spR7_0),.clk(gclk));
	jdff dff_B_G2fLqw7w0_0(.din(w_dff_B_mPn94spR7_0),.dout(w_dff_B_G2fLqw7w0_0),.clk(gclk));
	jdff dff_B_z7L8HmGP2_0(.din(w_dff_B_G2fLqw7w0_0),.dout(w_dff_B_z7L8HmGP2_0),.clk(gclk));
	jdff dff_B_bOYXgBcF0_0(.din(w_dff_B_z7L8HmGP2_0),.dout(w_dff_B_bOYXgBcF0_0),.clk(gclk));
	jdff dff_B_CKQVhFj62_0(.din(w_dff_B_bOYXgBcF0_0),.dout(w_dff_B_CKQVhFj62_0),.clk(gclk));
	jdff dff_B_6ASsgS4d6_0(.din(w_dff_B_CKQVhFj62_0),.dout(w_dff_B_6ASsgS4d6_0),.clk(gclk));
	jdff dff_B_AoWd7XVJ6_0(.din(w_dff_B_6ASsgS4d6_0),.dout(w_dff_B_AoWd7XVJ6_0),.clk(gclk));
	jdff dff_B_mT6luw553_0(.din(w_dff_B_AoWd7XVJ6_0),.dout(w_dff_B_mT6luw553_0),.clk(gclk));
	jdff dff_B_RYyCr0Jl8_0(.din(w_dff_B_mT6luw553_0),.dout(w_dff_B_RYyCr0Jl8_0),.clk(gclk));
	jdff dff_B_VQHeG0RE9_0(.din(w_dff_B_RYyCr0Jl8_0),.dout(w_dff_B_VQHeG0RE9_0),.clk(gclk));
	jdff dff_B_U1MaEUnW4_0(.din(w_dff_B_VQHeG0RE9_0),.dout(w_dff_B_U1MaEUnW4_0),.clk(gclk));
	jdff dff_B_7eW38oI83_0(.din(w_dff_B_U1MaEUnW4_0),.dout(w_dff_B_7eW38oI83_0),.clk(gclk));
	jdff dff_B_nMZ7Qmwa1_0(.din(w_dff_B_7eW38oI83_0),.dout(w_dff_B_nMZ7Qmwa1_0),.clk(gclk));
	jdff dff_B_pJdkeARO9_0(.din(w_dff_B_nMZ7Qmwa1_0),.dout(w_dff_B_pJdkeARO9_0),.clk(gclk));
	jdff dff_B_RWqMEuI92_0(.din(w_dff_B_pJdkeARO9_0),.dout(w_dff_B_RWqMEuI92_0),.clk(gclk));
	jdff dff_B_PeohdI955_0(.din(w_dff_B_RWqMEuI92_0),.dout(w_dff_B_PeohdI955_0),.clk(gclk));
	jdff dff_B_W1uLlMar7_0(.din(w_dff_B_PeohdI955_0),.dout(w_dff_B_W1uLlMar7_0),.clk(gclk));
	jdff dff_B_nNlo2cPj5_0(.din(w_dff_B_W1uLlMar7_0),.dout(w_dff_B_nNlo2cPj5_0),.clk(gclk));
	jdff dff_B_IQRe3tTm0_0(.din(w_dff_B_nNlo2cPj5_0),.dout(w_dff_B_IQRe3tTm0_0),.clk(gclk));
	jdff dff_B_002zxTFy5_0(.din(w_dff_B_IQRe3tTm0_0),.dout(w_dff_B_002zxTFy5_0),.clk(gclk));
	jdff dff_B_xX7EUYh51_0(.din(w_dff_B_002zxTFy5_0),.dout(w_dff_B_xX7EUYh51_0),.clk(gclk));
	jdff dff_B_rxmp0ZJd1_0(.din(w_dff_B_xX7EUYh51_0),.dout(w_dff_B_rxmp0ZJd1_0),.clk(gclk));
	jdff dff_B_ZJKUfoRx0_0(.din(w_dff_B_rxmp0ZJd1_0),.dout(w_dff_B_ZJKUfoRx0_0),.clk(gclk));
	jdff dff_B_T0Aj8f960_0(.din(w_dff_B_ZJKUfoRx0_0),.dout(w_dff_B_T0Aj8f960_0),.clk(gclk));
	jdff dff_B_9irEKkA48_0(.din(w_dff_B_T0Aj8f960_0),.dout(w_dff_B_9irEKkA48_0),.clk(gclk));
	jdff dff_B_Eztovppw0_0(.din(w_dff_B_9irEKkA48_0),.dout(w_dff_B_Eztovppw0_0),.clk(gclk));
	jdff dff_B_iTMTLhTL3_0(.din(w_dff_B_Eztovppw0_0),.dout(w_dff_B_iTMTLhTL3_0),.clk(gclk));
	jdff dff_B_ZwJF8mxF1_0(.din(w_dff_B_iTMTLhTL3_0),.dout(w_dff_B_ZwJF8mxF1_0),.clk(gclk));
	jdff dff_B_4r5E3uWs9_0(.din(w_dff_B_ZwJF8mxF1_0),.dout(w_dff_B_4r5E3uWs9_0),.clk(gclk));
	jdff dff_B_5l6h7VVR4_0(.din(w_dff_B_4r5E3uWs9_0),.dout(w_dff_B_5l6h7VVR4_0),.clk(gclk));
	jdff dff_B_Y3hWmEb72_0(.din(w_dff_B_5l6h7VVR4_0),.dout(w_dff_B_Y3hWmEb72_0),.clk(gclk));
	jdff dff_B_oK8jQHfj9_0(.din(w_dff_B_Y3hWmEb72_0),.dout(w_dff_B_oK8jQHfj9_0),.clk(gclk));
	jdff dff_B_E2MPlqZv8_0(.din(w_dff_B_oK8jQHfj9_0),.dout(w_dff_B_E2MPlqZv8_0),.clk(gclk));
	jdff dff_B_LPwPZoL92_0(.din(w_dff_B_E2MPlqZv8_0),.dout(w_dff_B_LPwPZoL92_0),.clk(gclk));
	jdff dff_B_7eD41BBB2_0(.din(w_dff_B_LPwPZoL92_0),.dout(w_dff_B_7eD41BBB2_0),.clk(gclk));
	jdff dff_B_flSfCuIw5_0(.din(w_dff_B_7eD41BBB2_0),.dout(w_dff_B_flSfCuIw5_0),.clk(gclk));
	jdff dff_B_Xp9QBovF0_0(.din(w_dff_B_flSfCuIw5_0),.dout(w_dff_B_Xp9QBovF0_0),.clk(gclk));
	jdff dff_B_CDZDHRbE1_0(.din(w_dff_B_Xp9QBovF0_0),.dout(w_dff_B_CDZDHRbE1_0),.clk(gclk));
	jdff dff_B_2LytpcSC1_0(.din(w_dff_B_CDZDHRbE1_0),.dout(w_dff_B_2LytpcSC1_0),.clk(gclk));
	jdff dff_B_txdEc3XX4_0(.din(w_dff_B_2LytpcSC1_0),.dout(w_dff_B_txdEc3XX4_0),.clk(gclk));
	jdff dff_B_24N9Dxzp9_0(.din(w_dff_B_txdEc3XX4_0),.dout(w_dff_B_24N9Dxzp9_0),.clk(gclk));
	jdff dff_B_xuLvqdrB8_0(.din(w_dff_B_24N9Dxzp9_0),.dout(w_dff_B_xuLvqdrB8_0),.clk(gclk));
	jdff dff_B_kmVvkjfY9_0(.din(w_dff_B_xuLvqdrB8_0),.dout(w_dff_B_kmVvkjfY9_0),.clk(gclk));
	jdff dff_B_vghfCz9w4_0(.din(w_dff_B_kmVvkjfY9_0),.dout(w_dff_B_vghfCz9w4_0),.clk(gclk));
	jdff dff_B_cCrAwSXp4_0(.din(w_dff_B_vghfCz9w4_0),.dout(w_dff_B_cCrAwSXp4_0),.clk(gclk));
	jdff dff_B_akSnWl4a4_0(.din(w_dff_B_cCrAwSXp4_0),.dout(w_dff_B_akSnWl4a4_0),.clk(gclk));
	jdff dff_B_g8inP2hw8_0(.din(w_dff_B_akSnWl4a4_0),.dout(w_dff_B_g8inP2hw8_0),.clk(gclk));
	jdff dff_B_OOaMoRMD8_0(.din(w_dff_B_g8inP2hw8_0),.dout(w_dff_B_OOaMoRMD8_0),.clk(gclk));
	jdff dff_B_N43TeiBD7_0(.din(n754),.dout(w_dff_B_N43TeiBD7_0),.clk(gclk));
	jdff dff_B_LkDa6SzL3_0(.din(w_dff_B_N43TeiBD7_0),.dout(w_dff_B_LkDa6SzL3_0),.clk(gclk));
	jdff dff_B_edGyBkYI7_0(.din(w_dff_B_LkDa6SzL3_0),.dout(w_dff_B_edGyBkYI7_0),.clk(gclk));
	jdff dff_B_LFmc4WlW5_0(.din(w_dff_B_edGyBkYI7_0),.dout(w_dff_B_LFmc4WlW5_0),.clk(gclk));
	jdff dff_B_dhV4u7s49_0(.din(w_dff_B_LFmc4WlW5_0),.dout(w_dff_B_dhV4u7s49_0),.clk(gclk));
	jdff dff_B_ezBkCv0e7_0(.din(w_dff_B_dhV4u7s49_0),.dout(w_dff_B_ezBkCv0e7_0),.clk(gclk));
	jdff dff_B_nTKJilRV1_0(.din(w_dff_B_ezBkCv0e7_0),.dout(w_dff_B_nTKJilRV1_0),.clk(gclk));
	jdff dff_B_ac8co5MC9_0(.din(w_dff_B_nTKJilRV1_0),.dout(w_dff_B_ac8co5MC9_0),.clk(gclk));
	jdff dff_B_Ec9Nilic5_0(.din(w_dff_B_ac8co5MC9_0),.dout(w_dff_B_Ec9Nilic5_0),.clk(gclk));
	jdff dff_B_FgwoQ8oz7_0(.din(w_dff_B_Ec9Nilic5_0),.dout(w_dff_B_FgwoQ8oz7_0),.clk(gclk));
	jdff dff_B_5U9XJDKT8_0(.din(w_dff_B_FgwoQ8oz7_0),.dout(w_dff_B_5U9XJDKT8_0),.clk(gclk));
	jdff dff_B_BHAwMt4x9_0(.din(w_dff_B_5U9XJDKT8_0),.dout(w_dff_B_BHAwMt4x9_0),.clk(gclk));
	jdff dff_B_HyKhLGrt0_0(.din(w_dff_B_BHAwMt4x9_0),.dout(w_dff_B_HyKhLGrt0_0),.clk(gclk));
	jdff dff_B_ahlsgZnF1_0(.din(w_dff_B_HyKhLGrt0_0),.dout(w_dff_B_ahlsgZnF1_0),.clk(gclk));
	jdff dff_B_dDsQNd3P2_0(.din(w_dff_B_ahlsgZnF1_0),.dout(w_dff_B_dDsQNd3P2_0),.clk(gclk));
	jdff dff_B_FtIWvVPE0_0(.din(w_dff_B_dDsQNd3P2_0),.dout(w_dff_B_FtIWvVPE0_0),.clk(gclk));
	jdff dff_B_rTIcnVp34_0(.din(w_dff_B_FtIWvVPE0_0),.dout(w_dff_B_rTIcnVp34_0),.clk(gclk));
	jdff dff_B_skcRmArv1_0(.din(w_dff_B_rTIcnVp34_0),.dout(w_dff_B_skcRmArv1_0),.clk(gclk));
	jdff dff_B_663jYFYu6_0(.din(w_dff_B_skcRmArv1_0),.dout(w_dff_B_663jYFYu6_0),.clk(gclk));
	jdff dff_B_DnYynrPR9_0(.din(w_dff_B_663jYFYu6_0),.dout(w_dff_B_DnYynrPR9_0),.clk(gclk));
	jdff dff_B_DNRvwmFk7_0(.din(w_dff_B_DnYynrPR9_0),.dout(w_dff_B_DNRvwmFk7_0),.clk(gclk));
	jdff dff_B_q2iQDC5i5_0(.din(w_dff_B_DNRvwmFk7_0),.dout(w_dff_B_q2iQDC5i5_0),.clk(gclk));
	jdff dff_B_FGpFsdqf2_0(.din(w_dff_B_q2iQDC5i5_0),.dout(w_dff_B_FGpFsdqf2_0),.clk(gclk));
	jdff dff_B_qJLgeLAP9_0(.din(w_dff_B_FGpFsdqf2_0),.dout(w_dff_B_qJLgeLAP9_0),.clk(gclk));
	jdff dff_B_DmqOkRzm7_0(.din(w_dff_B_qJLgeLAP9_0),.dout(w_dff_B_DmqOkRzm7_0),.clk(gclk));
	jdff dff_B_b182Fq3j2_0(.din(w_dff_B_DmqOkRzm7_0),.dout(w_dff_B_b182Fq3j2_0),.clk(gclk));
	jdff dff_B_xN4tYXk49_0(.din(w_dff_B_b182Fq3j2_0),.dout(w_dff_B_xN4tYXk49_0),.clk(gclk));
	jdff dff_B_9xug5xDH5_0(.din(w_dff_B_xN4tYXk49_0),.dout(w_dff_B_9xug5xDH5_0),.clk(gclk));
	jdff dff_B_B7r84Fjh7_0(.din(w_dff_B_9xug5xDH5_0),.dout(w_dff_B_B7r84Fjh7_0),.clk(gclk));
	jdff dff_B_6mQeXNux4_0(.din(w_dff_B_B7r84Fjh7_0),.dout(w_dff_B_6mQeXNux4_0),.clk(gclk));
	jdff dff_B_vmjRRzfx6_0(.din(w_dff_B_6mQeXNux4_0),.dout(w_dff_B_vmjRRzfx6_0),.clk(gclk));
	jdff dff_B_Q3Y7OAQm2_0(.din(w_dff_B_vmjRRzfx6_0),.dout(w_dff_B_Q3Y7OAQm2_0),.clk(gclk));
	jdff dff_B_5MvIazEW6_0(.din(w_dff_B_Q3Y7OAQm2_0),.dout(w_dff_B_5MvIazEW6_0),.clk(gclk));
	jdff dff_B_pbzTpi4o4_0(.din(w_dff_B_5MvIazEW6_0),.dout(w_dff_B_pbzTpi4o4_0),.clk(gclk));
	jdff dff_B_kmtiB6zx5_0(.din(w_dff_B_pbzTpi4o4_0),.dout(w_dff_B_kmtiB6zx5_0),.clk(gclk));
	jdff dff_B_Fx10VEcz9_0(.din(w_dff_B_kmtiB6zx5_0),.dout(w_dff_B_Fx10VEcz9_0),.clk(gclk));
	jdff dff_B_5wLAcNXb8_0(.din(w_dff_B_Fx10VEcz9_0),.dout(w_dff_B_5wLAcNXb8_0),.clk(gclk));
	jdff dff_B_2STa13D53_0(.din(w_dff_B_5wLAcNXb8_0),.dout(w_dff_B_2STa13D53_0),.clk(gclk));
	jdff dff_B_uyOxNtuO5_0(.din(w_dff_B_2STa13D53_0),.dout(w_dff_B_uyOxNtuO5_0),.clk(gclk));
	jdff dff_B_IrJaJ9z73_0(.din(w_dff_B_uyOxNtuO5_0),.dout(w_dff_B_IrJaJ9z73_0),.clk(gclk));
	jdff dff_B_bZqN31Th5_0(.din(w_dff_B_IrJaJ9z73_0),.dout(w_dff_B_bZqN31Th5_0),.clk(gclk));
	jdff dff_B_0qqe029j5_0(.din(w_dff_B_bZqN31Th5_0),.dout(w_dff_B_0qqe029j5_0),.clk(gclk));
	jdff dff_B_CmA98J3t2_0(.din(w_dff_B_0qqe029j5_0),.dout(w_dff_B_CmA98J3t2_0),.clk(gclk));
	jdff dff_B_4OBh7iPL5_0(.din(w_dff_B_CmA98J3t2_0),.dout(w_dff_B_4OBh7iPL5_0),.clk(gclk));
	jdff dff_B_XjSdbsaK1_0(.din(w_dff_B_4OBh7iPL5_0),.dout(w_dff_B_XjSdbsaK1_0),.clk(gclk));
	jdff dff_B_cUZt5DxM0_0(.din(w_dff_B_XjSdbsaK1_0),.dout(w_dff_B_cUZt5DxM0_0),.clk(gclk));
	jdff dff_B_Rh3ZUMp52_0(.din(w_dff_B_cUZt5DxM0_0),.dout(w_dff_B_Rh3ZUMp52_0),.clk(gclk));
	jdff dff_B_bPqCWENT8_0(.din(w_dff_B_Rh3ZUMp52_0),.dout(w_dff_B_bPqCWENT8_0),.clk(gclk));
	jdff dff_B_6JwUP94n3_0(.din(w_dff_B_bPqCWENT8_0),.dout(w_dff_B_6JwUP94n3_0),.clk(gclk));
	jdff dff_B_mHpZ10hv2_0(.din(w_dff_B_6JwUP94n3_0),.dout(w_dff_B_mHpZ10hv2_0),.clk(gclk));
	jdff dff_B_L1rg5cw88_0(.din(w_dff_B_mHpZ10hv2_0),.dout(w_dff_B_L1rg5cw88_0),.clk(gclk));
	jdff dff_B_wneQG0uC7_0(.din(w_dff_B_L1rg5cw88_0),.dout(w_dff_B_wneQG0uC7_0),.clk(gclk));
	jdff dff_B_M5p0jvDy7_0(.din(w_dff_B_wneQG0uC7_0),.dout(w_dff_B_M5p0jvDy7_0),.clk(gclk));
	jdff dff_B_DK1hHNJv9_0(.din(w_dff_B_M5p0jvDy7_0),.dout(w_dff_B_DK1hHNJv9_0),.clk(gclk));
	jdff dff_B_Ryw32P2a3_0(.din(w_dff_B_DK1hHNJv9_0),.dout(w_dff_B_Ryw32P2a3_0),.clk(gclk));
	jdff dff_B_BSSWA0AA3_0(.din(w_dff_B_Ryw32P2a3_0),.dout(w_dff_B_BSSWA0AA3_0),.clk(gclk));
	jdff dff_B_lVJ0xiQs5_0(.din(w_dff_B_BSSWA0AA3_0),.dout(w_dff_B_lVJ0xiQs5_0),.clk(gclk));
	jdff dff_B_G2lXWRYT1_0(.din(w_dff_B_lVJ0xiQs5_0),.dout(w_dff_B_G2lXWRYT1_0),.clk(gclk));
	jdff dff_B_LIAYzsse5_0(.din(w_dff_B_G2lXWRYT1_0),.dout(w_dff_B_LIAYzsse5_0),.clk(gclk));
	jdff dff_B_f4nkdD6i2_0(.din(w_dff_B_LIAYzsse5_0),.dout(w_dff_B_f4nkdD6i2_0),.clk(gclk));
	jdff dff_B_fMEyUaIT3_0(.din(w_dff_B_f4nkdD6i2_0),.dout(w_dff_B_fMEyUaIT3_0),.clk(gclk));
	jdff dff_B_MJOgI5Tc8_0(.din(n760),.dout(w_dff_B_MJOgI5Tc8_0),.clk(gclk));
	jdff dff_B_l9494gur8_0(.din(w_dff_B_MJOgI5Tc8_0),.dout(w_dff_B_l9494gur8_0),.clk(gclk));
	jdff dff_B_0xgzJT2y1_0(.din(w_dff_B_l9494gur8_0),.dout(w_dff_B_0xgzJT2y1_0),.clk(gclk));
	jdff dff_B_mnqrLOv22_0(.din(w_dff_B_0xgzJT2y1_0),.dout(w_dff_B_mnqrLOv22_0),.clk(gclk));
	jdff dff_B_oXBcbJhl3_0(.din(w_dff_B_mnqrLOv22_0),.dout(w_dff_B_oXBcbJhl3_0),.clk(gclk));
	jdff dff_B_3HCC4K1y4_0(.din(w_dff_B_oXBcbJhl3_0),.dout(w_dff_B_3HCC4K1y4_0),.clk(gclk));
	jdff dff_B_501avdZ33_0(.din(w_dff_B_3HCC4K1y4_0),.dout(w_dff_B_501avdZ33_0),.clk(gclk));
	jdff dff_B_asE3GayY1_0(.din(w_dff_B_501avdZ33_0),.dout(w_dff_B_asE3GayY1_0),.clk(gclk));
	jdff dff_B_iUDXFsaS3_0(.din(w_dff_B_asE3GayY1_0),.dout(w_dff_B_iUDXFsaS3_0),.clk(gclk));
	jdff dff_B_giK7g9yx2_0(.din(w_dff_B_iUDXFsaS3_0),.dout(w_dff_B_giK7g9yx2_0),.clk(gclk));
	jdff dff_B_6R7Dh7px6_0(.din(w_dff_B_giK7g9yx2_0),.dout(w_dff_B_6R7Dh7px6_0),.clk(gclk));
	jdff dff_B_Ifx59pLf6_0(.din(w_dff_B_6R7Dh7px6_0),.dout(w_dff_B_Ifx59pLf6_0),.clk(gclk));
	jdff dff_B_pimWYWdx2_0(.din(w_dff_B_Ifx59pLf6_0),.dout(w_dff_B_pimWYWdx2_0),.clk(gclk));
	jdff dff_B_oIFulJes4_0(.din(w_dff_B_pimWYWdx2_0),.dout(w_dff_B_oIFulJes4_0),.clk(gclk));
	jdff dff_B_WuPeaXXs8_0(.din(w_dff_B_oIFulJes4_0),.dout(w_dff_B_WuPeaXXs8_0),.clk(gclk));
	jdff dff_B_5xHWplqn2_0(.din(w_dff_B_WuPeaXXs8_0),.dout(w_dff_B_5xHWplqn2_0),.clk(gclk));
	jdff dff_B_gC55LX6C2_0(.din(w_dff_B_5xHWplqn2_0),.dout(w_dff_B_gC55LX6C2_0),.clk(gclk));
	jdff dff_B_o64XK9bE4_0(.din(w_dff_B_gC55LX6C2_0),.dout(w_dff_B_o64XK9bE4_0),.clk(gclk));
	jdff dff_B_fCQBGIZ69_0(.din(w_dff_B_o64XK9bE4_0),.dout(w_dff_B_fCQBGIZ69_0),.clk(gclk));
	jdff dff_B_0QA7Xj7o3_0(.din(w_dff_B_fCQBGIZ69_0),.dout(w_dff_B_0QA7Xj7o3_0),.clk(gclk));
	jdff dff_B_Rt9HNFXs3_0(.din(w_dff_B_0QA7Xj7o3_0),.dout(w_dff_B_Rt9HNFXs3_0),.clk(gclk));
	jdff dff_B_DPB8dIwm2_0(.din(w_dff_B_Rt9HNFXs3_0),.dout(w_dff_B_DPB8dIwm2_0),.clk(gclk));
	jdff dff_B_edIqXs2R6_0(.din(w_dff_B_DPB8dIwm2_0),.dout(w_dff_B_edIqXs2R6_0),.clk(gclk));
	jdff dff_B_dBZ8UPtm0_0(.din(w_dff_B_edIqXs2R6_0),.dout(w_dff_B_dBZ8UPtm0_0),.clk(gclk));
	jdff dff_B_eoV108Gw8_0(.din(w_dff_B_dBZ8UPtm0_0),.dout(w_dff_B_eoV108Gw8_0),.clk(gclk));
	jdff dff_B_ZURMnqwx6_0(.din(w_dff_B_eoV108Gw8_0),.dout(w_dff_B_ZURMnqwx6_0),.clk(gclk));
	jdff dff_B_bckQAAPB7_0(.din(w_dff_B_ZURMnqwx6_0),.dout(w_dff_B_bckQAAPB7_0),.clk(gclk));
	jdff dff_B_AOn8vtPx9_0(.din(w_dff_B_bckQAAPB7_0),.dout(w_dff_B_AOn8vtPx9_0),.clk(gclk));
	jdff dff_B_F2WvPzWR4_0(.din(w_dff_B_AOn8vtPx9_0),.dout(w_dff_B_F2WvPzWR4_0),.clk(gclk));
	jdff dff_B_UUF9AEbV8_0(.din(w_dff_B_F2WvPzWR4_0),.dout(w_dff_B_UUF9AEbV8_0),.clk(gclk));
	jdff dff_B_qKcTuZkc3_0(.din(w_dff_B_UUF9AEbV8_0),.dout(w_dff_B_qKcTuZkc3_0),.clk(gclk));
	jdff dff_B_PSBnQFqD2_0(.din(w_dff_B_qKcTuZkc3_0),.dout(w_dff_B_PSBnQFqD2_0),.clk(gclk));
	jdff dff_B_YwZPwZcG8_0(.din(w_dff_B_PSBnQFqD2_0),.dout(w_dff_B_YwZPwZcG8_0),.clk(gclk));
	jdff dff_B_y2YeFqmQ4_0(.din(w_dff_B_YwZPwZcG8_0),.dout(w_dff_B_y2YeFqmQ4_0),.clk(gclk));
	jdff dff_B_RnW0Gm953_0(.din(w_dff_B_y2YeFqmQ4_0),.dout(w_dff_B_RnW0Gm953_0),.clk(gclk));
	jdff dff_B_RVI3Wf2a7_0(.din(w_dff_B_RnW0Gm953_0),.dout(w_dff_B_RVI3Wf2a7_0),.clk(gclk));
	jdff dff_B_Sf5gLHx05_0(.din(w_dff_B_RVI3Wf2a7_0),.dout(w_dff_B_Sf5gLHx05_0),.clk(gclk));
	jdff dff_B_Ha4Boxhu5_0(.din(w_dff_B_Sf5gLHx05_0),.dout(w_dff_B_Ha4Boxhu5_0),.clk(gclk));
	jdff dff_B_ZzaDVEjL2_0(.din(w_dff_B_Ha4Boxhu5_0),.dout(w_dff_B_ZzaDVEjL2_0),.clk(gclk));
	jdff dff_B_9Y3EJ03L8_0(.din(w_dff_B_ZzaDVEjL2_0),.dout(w_dff_B_9Y3EJ03L8_0),.clk(gclk));
	jdff dff_B_5F1KABog7_0(.din(w_dff_B_9Y3EJ03L8_0),.dout(w_dff_B_5F1KABog7_0),.clk(gclk));
	jdff dff_B_kr0RBh2v6_0(.din(w_dff_B_5F1KABog7_0),.dout(w_dff_B_kr0RBh2v6_0),.clk(gclk));
	jdff dff_B_f6rVGAmV0_0(.din(w_dff_B_kr0RBh2v6_0),.dout(w_dff_B_f6rVGAmV0_0),.clk(gclk));
	jdff dff_B_o8aPkdjX8_0(.din(w_dff_B_f6rVGAmV0_0),.dout(w_dff_B_o8aPkdjX8_0),.clk(gclk));
	jdff dff_B_cEBpO5LL5_0(.din(w_dff_B_o8aPkdjX8_0),.dout(w_dff_B_cEBpO5LL5_0),.clk(gclk));
	jdff dff_B_G3IMKIUJ8_0(.din(w_dff_B_cEBpO5LL5_0),.dout(w_dff_B_G3IMKIUJ8_0),.clk(gclk));
	jdff dff_B_XuPlBzz87_0(.din(w_dff_B_G3IMKIUJ8_0),.dout(w_dff_B_XuPlBzz87_0),.clk(gclk));
	jdff dff_B_DKD7axMF5_0(.din(w_dff_B_XuPlBzz87_0),.dout(w_dff_B_DKD7axMF5_0),.clk(gclk));
	jdff dff_B_73KFAbEP4_0(.din(w_dff_B_DKD7axMF5_0),.dout(w_dff_B_73KFAbEP4_0),.clk(gclk));
	jdff dff_B_62dTet6S2_0(.din(w_dff_B_73KFAbEP4_0),.dout(w_dff_B_62dTet6S2_0),.clk(gclk));
	jdff dff_B_bKUQ5i801_0(.din(w_dff_B_62dTet6S2_0),.dout(w_dff_B_bKUQ5i801_0),.clk(gclk));
	jdff dff_B_0Wk2wlyL4_0(.din(w_dff_B_bKUQ5i801_0),.dout(w_dff_B_0Wk2wlyL4_0),.clk(gclk));
	jdff dff_B_2OReU4Y06_0(.din(w_dff_B_0Wk2wlyL4_0),.dout(w_dff_B_2OReU4Y06_0),.clk(gclk));
	jdff dff_B_Lv8WuXOu5_0(.din(w_dff_B_2OReU4Y06_0),.dout(w_dff_B_Lv8WuXOu5_0),.clk(gclk));
	jdff dff_B_Af5Y2zzz6_0(.din(w_dff_B_Lv8WuXOu5_0),.dout(w_dff_B_Af5Y2zzz6_0),.clk(gclk));
	jdff dff_B_XkPvtMI32_0(.din(w_dff_B_Af5Y2zzz6_0),.dout(w_dff_B_XkPvtMI32_0),.clk(gclk));
	jdff dff_B_mJ1XUryB9_0(.din(w_dff_B_XkPvtMI32_0),.dout(w_dff_B_mJ1XUryB9_0),.clk(gclk));
	jdff dff_B_gibCcTwN0_0(.din(w_dff_B_mJ1XUryB9_0),.dout(w_dff_B_gibCcTwN0_0),.clk(gclk));
	jdff dff_B_79Vh9ZuL1_0(.din(w_dff_B_gibCcTwN0_0),.dout(w_dff_B_79Vh9ZuL1_0),.clk(gclk));
	jdff dff_B_JdGYQgyg8_0(.din(w_dff_B_79Vh9ZuL1_0),.dout(w_dff_B_JdGYQgyg8_0),.clk(gclk));
	jdff dff_B_6VzbeitE7_0(.din(w_dff_B_JdGYQgyg8_0),.dout(w_dff_B_6VzbeitE7_0),.clk(gclk));
	jdff dff_B_X8L8LwPo4_0(.din(w_dff_B_6VzbeitE7_0),.dout(w_dff_B_X8L8LwPo4_0),.clk(gclk));
	jdff dff_B_cIvQSKz17_0(.din(n766),.dout(w_dff_B_cIvQSKz17_0),.clk(gclk));
	jdff dff_B_bCDgvB6u8_0(.din(w_dff_B_cIvQSKz17_0),.dout(w_dff_B_bCDgvB6u8_0),.clk(gclk));
	jdff dff_B_AZa3Ty4w1_0(.din(w_dff_B_bCDgvB6u8_0),.dout(w_dff_B_AZa3Ty4w1_0),.clk(gclk));
	jdff dff_B_awCzRtA72_0(.din(w_dff_B_AZa3Ty4w1_0),.dout(w_dff_B_awCzRtA72_0),.clk(gclk));
	jdff dff_B_MSTl2hYf1_0(.din(w_dff_B_awCzRtA72_0),.dout(w_dff_B_MSTl2hYf1_0),.clk(gclk));
	jdff dff_B_O9NJs6ZX4_0(.din(w_dff_B_MSTl2hYf1_0),.dout(w_dff_B_O9NJs6ZX4_0),.clk(gclk));
	jdff dff_B_YRxR1LVA8_0(.din(w_dff_B_O9NJs6ZX4_0),.dout(w_dff_B_YRxR1LVA8_0),.clk(gclk));
	jdff dff_B_G8PskRw15_0(.din(w_dff_B_YRxR1LVA8_0),.dout(w_dff_B_G8PskRw15_0),.clk(gclk));
	jdff dff_B_Z3WDt5Ih7_0(.din(w_dff_B_G8PskRw15_0),.dout(w_dff_B_Z3WDt5Ih7_0),.clk(gclk));
	jdff dff_B_lwby5Mh50_0(.din(w_dff_B_Z3WDt5Ih7_0),.dout(w_dff_B_lwby5Mh50_0),.clk(gclk));
	jdff dff_B_eic3tLtR8_0(.din(w_dff_B_lwby5Mh50_0),.dout(w_dff_B_eic3tLtR8_0),.clk(gclk));
	jdff dff_B_cBEC74E59_0(.din(w_dff_B_eic3tLtR8_0),.dout(w_dff_B_cBEC74E59_0),.clk(gclk));
	jdff dff_B_h9OvX51Z9_0(.din(w_dff_B_cBEC74E59_0),.dout(w_dff_B_h9OvX51Z9_0),.clk(gclk));
	jdff dff_B_OMdxyjmK4_0(.din(w_dff_B_h9OvX51Z9_0),.dout(w_dff_B_OMdxyjmK4_0),.clk(gclk));
	jdff dff_B_oGtPmaNF8_0(.din(w_dff_B_OMdxyjmK4_0),.dout(w_dff_B_oGtPmaNF8_0),.clk(gclk));
	jdff dff_B_kQsivHJf4_0(.din(w_dff_B_oGtPmaNF8_0),.dout(w_dff_B_kQsivHJf4_0),.clk(gclk));
	jdff dff_B_Qf67nob83_0(.din(w_dff_B_kQsivHJf4_0),.dout(w_dff_B_Qf67nob83_0),.clk(gclk));
	jdff dff_B_KoaiLJSL2_0(.din(w_dff_B_Qf67nob83_0),.dout(w_dff_B_KoaiLJSL2_0),.clk(gclk));
	jdff dff_B_5rTuTRhA7_0(.din(w_dff_B_KoaiLJSL2_0),.dout(w_dff_B_5rTuTRhA7_0),.clk(gclk));
	jdff dff_B_BgkCpQ985_0(.din(w_dff_B_5rTuTRhA7_0),.dout(w_dff_B_BgkCpQ985_0),.clk(gclk));
	jdff dff_B_xW01B4j49_0(.din(w_dff_B_BgkCpQ985_0),.dout(w_dff_B_xW01B4j49_0),.clk(gclk));
	jdff dff_B_mLA5TeLw9_0(.din(w_dff_B_xW01B4j49_0),.dout(w_dff_B_mLA5TeLw9_0),.clk(gclk));
	jdff dff_B_RtLE5QMn2_0(.din(w_dff_B_mLA5TeLw9_0),.dout(w_dff_B_RtLE5QMn2_0),.clk(gclk));
	jdff dff_B_1OZ8NVel5_0(.din(w_dff_B_RtLE5QMn2_0),.dout(w_dff_B_1OZ8NVel5_0),.clk(gclk));
	jdff dff_B_gGFcK9Yb2_0(.din(w_dff_B_1OZ8NVel5_0),.dout(w_dff_B_gGFcK9Yb2_0),.clk(gclk));
	jdff dff_B_BEPcJJdl5_0(.din(w_dff_B_gGFcK9Yb2_0),.dout(w_dff_B_BEPcJJdl5_0),.clk(gclk));
	jdff dff_B_OuqUwewK7_0(.din(w_dff_B_BEPcJJdl5_0),.dout(w_dff_B_OuqUwewK7_0),.clk(gclk));
	jdff dff_B_LhWWmIhT3_0(.din(w_dff_B_OuqUwewK7_0),.dout(w_dff_B_LhWWmIhT3_0),.clk(gclk));
	jdff dff_B_wrPEluAf3_0(.din(w_dff_B_LhWWmIhT3_0),.dout(w_dff_B_wrPEluAf3_0),.clk(gclk));
	jdff dff_B_v2q8aYLY4_0(.din(w_dff_B_wrPEluAf3_0),.dout(w_dff_B_v2q8aYLY4_0),.clk(gclk));
	jdff dff_B_gFOpIouM5_0(.din(w_dff_B_v2q8aYLY4_0),.dout(w_dff_B_gFOpIouM5_0),.clk(gclk));
	jdff dff_B_n03IOPfk4_0(.din(w_dff_B_gFOpIouM5_0),.dout(w_dff_B_n03IOPfk4_0),.clk(gclk));
	jdff dff_B_lILpXwza7_0(.din(w_dff_B_n03IOPfk4_0),.dout(w_dff_B_lILpXwza7_0),.clk(gclk));
	jdff dff_B_krrbxW3D4_0(.din(w_dff_B_lILpXwza7_0),.dout(w_dff_B_krrbxW3D4_0),.clk(gclk));
	jdff dff_B_uz0YGazH1_0(.din(w_dff_B_krrbxW3D4_0),.dout(w_dff_B_uz0YGazH1_0),.clk(gclk));
	jdff dff_B_oeu2xniw1_0(.din(w_dff_B_uz0YGazH1_0),.dout(w_dff_B_oeu2xniw1_0),.clk(gclk));
	jdff dff_B_fwaYqs5M7_0(.din(w_dff_B_oeu2xniw1_0),.dout(w_dff_B_fwaYqs5M7_0),.clk(gclk));
	jdff dff_B_WIdKIBsv3_0(.din(w_dff_B_fwaYqs5M7_0),.dout(w_dff_B_WIdKIBsv3_0),.clk(gclk));
	jdff dff_B_CixI2yI33_0(.din(w_dff_B_WIdKIBsv3_0),.dout(w_dff_B_CixI2yI33_0),.clk(gclk));
	jdff dff_B_ElNs0U4u4_0(.din(w_dff_B_CixI2yI33_0),.dout(w_dff_B_ElNs0U4u4_0),.clk(gclk));
	jdff dff_B_64VOXAXb8_0(.din(w_dff_B_ElNs0U4u4_0),.dout(w_dff_B_64VOXAXb8_0),.clk(gclk));
	jdff dff_B_6OTmtGd90_0(.din(w_dff_B_64VOXAXb8_0),.dout(w_dff_B_6OTmtGd90_0),.clk(gclk));
	jdff dff_B_LV1iaPcs6_0(.din(w_dff_B_6OTmtGd90_0),.dout(w_dff_B_LV1iaPcs6_0),.clk(gclk));
	jdff dff_B_C8mbCvAT8_0(.din(w_dff_B_LV1iaPcs6_0),.dout(w_dff_B_C8mbCvAT8_0),.clk(gclk));
	jdff dff_B_wBKYXJd46_0(.din(w_dff_B_C8mbCvAT8_0),.dout(w_dff_B_wBKYXJd46_0),.clk(gclk));
	jdff dff_B_0cF1byO62_0(.din(w_dff_B_wBKYXJd46_0),.dout(w_dff_B_0cF1byO62_0),.clk(gclk));
	jdff dff_B_7tBP0pSU8_0(.din(w_dff_B_0cF1byO62_0),.dout(w_dff_B_7tBP0pSU8_0),.clk(gclk));
	jdff dff_B_YFOvMl5c1_0(.din(w_dff_B_7tBP0pSU8_0),.dout(w_dff_B_YFOvMl5c1_0),.clk(gclk));
	jdff dff_B_OZSfx8AM0_0(.din(w_dff_B_YFOvMl5c1_0),.dout(w_dff_B_OZSfx8AM0_0),.clk(gclk));
	jdff dff_B_dUtt2DQQ5_0(.din(w_dff_B_OZSfx8AM0_0),.dout(w_dff_B_dUtt2DQQ5_0),.clk(gclk));
	jdff dff_B_GEwKrSO94_0(.din(w_dff_B_dUtt2DQQ5_0),.dout(w_dff_B_GEwKrSO94_0),.clk(gclk));
	jdff dff_B_bU9DLaMx5_0(.din(w_dff_B_GEwKrSO94_0),.dout(w_dff_B_bU9DLaMx5_0),.clk(gclk));
	jdff dff_B_XPR0PIQn0_0(.din(w_dff_B_bU9DLaMx5_0),.dout(w_dff_B_XPR0PIQn0_0),.clk(gclk));
	jdff dff_B_7rcaRNpq3_0(.din(w_dff_B_XPR0PIQn0_0),.dout(w_dff_B_7rcaRNpq3_0),.clk(gclk));
	jdff dff_B_BeQ7UtIn1_0(.din(w_dff_B_7rcaRNpq3_0),.dout(w_dff_B_BeQ7UtIn1_0),.clk(gclk));
	jdff dff_B_snrQQy319_0(.din(w_dff_B_BeQ7UtIn1_0),.dout(w_dff_B_snrQQy319_0),.clk(gclk));
	jdff dff_B_97akbQ6i1_0(.din(w_dff_B_snrQQy319_0),.dout(w_dff_B_97akbQ6i1_0),.clk(gclk));
	jdff dff_B_6LC8AMi52_0(.din(w_dff_B_97akbQ6i1_0),.dout(w_dff_B_6LC8AMi52_0),.clk(gclk));
	jdff dff_B_oLV1RueZ1_0(.din(w_dff_B_6LC8AMi52_0),.dout(w_dff_B_oLV1RueZ1_0),.clk(gclk));
	jdff dff_B_RdcO64tI8_0(.din(w_dff_B_oLV1RueZ1_0),.dout(w_dff_B_RdcO64tI8_0),.clk(gclk));
	jdff dff_B_ou7AWJVb2_0(.din(w_dff_B_RdcO64tI8_0),.dout(w_dff_B_ou7AWJVb2_0),.clk(gclk));
	jdff dff_B_qyexQIWU9_0(.din(w_dff_B_ou7AWJVb2_0),.dout(w_dff_B_qyexQIWU9_0),.clk(gclk));
	jdff dff_B_9ivRqQdT2_0(.din(w_dff_B_qyexQIWU9_0),.dout(w_dff_B_9ivRqQdT2_0),.clk(gclk));
	jdff dff_B_jk3ijHHm1_0(.din(n772),.dout(w_dff_B_jk3ijHHm1_0),.clk(gclk));
	jdff dff_B_H93DD0nF3_0(.din(w_dff_B_jk3ijHHm1_0),.dout(w_dff_B_H93DD0nF3_0),.clk(gclk));
	jdff dff_B_8SXtvf059_0(.din(w_dff_B_H93DD0nF3_0),.dout(w_dff_B_8SXtvf059_0),.clk(gclk));
	jdff dff_B_MYuLOHxF1_0(.din(w_dff_B_8SXtvf059_0),.dout(w_dff_B_MYuLOHxF1_0),.clk(gclk));
	jdff dff_B_0UMr1DXF2_0(.din(w_dff_B_MYuLOHxF1_0),.dout(w_dff_B_0UMr1DXF2_0),.clk(gclk));
	jdff dff_B_ByR9WVct7_0(.din(w_dff_B_0UMr1DXF2_0),.dout(w_dff_B_ByR9WVct7_0),.clk(gclk));
	jdff dff_B_DFE8za0Y6_0(.din(w_dff_B_ByR9WVct7_0),.dout(w_dff_B_DFE8za0Y6_0),.clk(gclk));
	jdff dff_B_eTO73Wi26_0(.din(w_dff_B_DFE8za0Y6_0),.dout(w_dff_B_eTO73Wi26_0),.clk(gclk));
	jdff dff_B_UgDRVKEi3_0(.din(w_dff_B_eTO73Wi26_0),.dout(w_dff_B_UgDRVKEi3_0),.clk(gclk));
	jdff dff_B_r9BUGi6K8_0(.din(w_dff_B_UgDRVKEi3_0),.dout(w_dff_B_r9BUGi6K8_0),.clk(gclk));
	jdff dff_B_ilVFZ8n37_0(.din(w_dff_B_r9BUGi6K8_0),.dout(w_dff_B_ilVFZ8n37_0),.clk(gclk));
	jdff dff_B_mUp05Keq0_0(.din(w_dff_B_ilVFZ8n37_0),.dout(w_dff_B_mUp05Keq0_0),.clk(gclk));
	jdff dff_B_7mz2ApX05_0(.din(w_dff_B_mUp05Keq0_0),.dout(w_dff_B_7mz2ApX05_0),.clk(gclk));
	jdff dff_B_uvEu02rc7_0(.din(w_dff_B_7mz2ApX05_0),.dout(w_dff_B_uvEu02rc7_0),.clk(gclk));
	jdff dff_B_yA5JL2DC2_0(.din(w_dff_B_uvEu02rc7_0),.dout(w_dff_B_yA5JL2DC2_0),.clk(gclk));
	jdff dff_B_oeXcKNM27_0(.din(w_dff_B_yA5JL2DC2_0),.dout(w_dff_B_oeXcKNM27_0),.clk(gclk));
	jdff dff_B_4RqP3Tsd3_0(.din(w_dff_B_oeXcKNM27_0),.dout(w_dff_B_4RqP3Tsd3_0),.clk(gclk));
	jdff dff_B_UsHcIBFJ8_0(.din(w_dff_B_4RqP3Tsd3_0),.dout(w_dff_B_UsHcIBFJ8_0),.clk(gclk));
	jdff dff_B_ZXKcvya14_0(.din(w_dff_B_UsHcIBFJ8_0),.dout(w_dff_B_ZXKcvya14_0),.clk(gclk));
	jdff dff_B_tYyKXsSX6_0(.din(w_dff_B_ZXKcvya14_0),.dout(w_dff_B_tYyKXsSX6_0),.clk(gclk));
	jdff dff_B_VQNZlPJU6_0(.din(w_dff_B_tYyKXsSX6_0),.dout(w_dff_B_VQNZlPJU6_0),.clk(gclk));
	jdff dff_B_H48w7ZK64_0(.din(w_dff_B_VQNZlPJU6_0),.dout(w_dff_B_H48w7ZK64_0),.clk(gclk));
	jdff dff_B_84PtJf3j8_0(.din(w_dff_B_H48w7ZK64_0),.dout(w_dff_B_84PtJf3j8_0),.clk(gclk));
	jdff dff_B_6vGDRYsK8_0(.din(w_dff_B_84PtJf3j8_0),.dout(w_dff_B_6vGDRYsK8_0),.clk(gclk));
	jdff dff_B_EmB0F3rz2_0(.din(w_dff_B_6vGDRYsK8_0),.dout(w_dff_B_EmB0F3rz2_0),.clk(gclk));
	jdff dff_B_YDxM8RvD9_0(.din(w_dff_B_EmB0F3rz2_0),.dout(w_dff_B_YDxM8RvD9_0),.clk(gclk));
	jdff dff_B_1bXMOldO3_0(.din(w_dff_B_YDxM8RvD9_0),.dout(w_dff_B_1bXMOldO3_0),.clk(gclk));
	jdff dff_B_a9yFeR9J2_0(.din(w_dff_B_1bXMOldO3_0),.dout(w_dff_B_a9yFeR9J2_0),.clk(gclk));
	jdff dff_B_yagBJeom2_0(.din(w_dff_B_a9yFeR9J2_0),.dout(w_dff_B_yagBJeom2_0),.clk(gclk));
	jdff dff_B_ZEFvyu3s1_0(.din(w_dff_B_yagBJeom2_0),.dout(w_dff_B_ZEFvyu3s1_0),.clk(gclk));
	jdff dff_B_UDWZpxXx5_0(.din(w_dff_B_ZEFvyu3s1_0),.dout(w_dff_B_UDWZpxXx5_0),.clk(gclk));
	jdff dff_B_S1OTrQt82_0(.din(w_dff_B_UDWZpxXx5_0),.dout(w_dff_B_S1OTrQt82_0),.clk(gclk));
	jdff dff_B_eNp8XkoY1_0(.din(w_dff_B_S1OTrQt82_0),.dout(w_dff_B_eNp8XkoY1_0),.clk(gclk));
	jdff dff_B_1X6NMZH98_0(.din(w_dff_B_eNp8XkoY1_0),.dout(w_dff_B_1X6NMZH98_0),.clk(gclk));
	jdff dff_B_g3LEmZ0x0_0(.din(w_dff_B_1X6NMZH98_0),.dout(w_dff_B_g3LEmZ0x0_0),.clk(gclk));
	jdff dff_B_KevCz5qh3_0(.din(w_dff_B_g3LEmZ0x0_0),.dout(w_dff_B_KevCz5qh3_0),.clk(gclk));
	jdff dff_B_7gtftLoY5_0(.din(w_dff_B_KevCz5qh3_0),.dout(w_dff_B_7gtftLoY5_0),.clk(gclk));
	jdff dff_B_BMELB3022_0(.din(w_dff_B_7gtftLoY5_0),.dout(w_dff_B_BMELB3022_0),.clk(gclk));
	jdff dff_B_m2QO5VPj0_0(.din(w_dff_B_BMELB3022_0),.dout(w_dff_B_m2QO5VPj0_0),.clk(gclk));
	jdff dff_B_B28S41fk9_0(.din(w_dff_B_m2QO5VPj0_0),.dout(w_dff_B_B28S41fk9_0),.clk(gclk));
	jdff dff_B_z5Dxn7683_0(.din(w_dff_B_B28S41fk9_0),.dout(w_dff_B_z5Dxn7683_0),.clk(gclk));
	jdff dff_B_507vvQel3_0(.din(w_dff_B_z5Dxn7683_0),.dout(w_dff_B_507vvQel3_0),.clk(gclk));
	jdff dff_B_0LW7LDP95_0(.din(w_dff_B_507vvQel3_0),.dout(w_dff_B_0LW7LDP95_0),.clk(gclk));
	jdff dff_B_Nex9M55S9_0(.din(w_dff_B_0LW7LDP95_0),.dout(w_dff_B_Nex9M55S9_0),.clk(gclk));
	jdff dff_B_CEVq4Ild6_0(.din(w_dff_B_Nex9M55S9_0),.dout(w_dff_B_CEVq4Ild6_0),.clk(gclk));
	jdff dff_B_Bj1gmevW8_0(.din(w_dff_B_CEVq4Ild6_0),.dout(w_dff_B_Bj1gmevW8_0),.clk(gclk));
	jdff dff_B_uMtHdGF47_0(.din(w_dff_B_Bj1gmevW8_0),.dout(w_dff_B_uMtHdGF47_0),.clk(gclk));
	jdff dff_B_fYF9UXz07_0(.din(w_dff_B_uMtHdGF47_0),.dout(w_dff_B_fYF9UXz07_0),.clk(gclk));
	jdff dff_B_QAeX4v7Y2_0(.din(w_dff_B_fYF9UXz07_0),.dout(w_dff_B_QAeX4v7Y2_0),.clk(gclk));
	jdff dff_B_4f3IQ6te8_0(.din(w_dff_B_QAeX4v7Y2_0),.dout(w_dff_B_4f3IQ6te8_0),.clk(gclk));
	jdff dff_B_PxVXR3hD0_0(.din(w_dff_B_4f3IQ6te8_0),.dout(w_dff_B_PxVXR3hD0_0),.clk(gclk));
	jdff dff_B_nsnTKwkU2_0(.din(w_dff_B_PxVXR3hD0_0),.dout(w_dff_B_nsnTKwkU2_0),.clk(gclk));
	jdff dff_B_6gGyzA4X6_0(.din(w_dff_B_nsnTKwkU2_0),.dout(w_dff_B_6gGyzA4X6_0),.clk(gclk));
	jdff dff_B_TaqQMqcn5_0(.din(w_dff_B_6gGyzA4X6_0),.dout(w_dff_B_TaqQMqcn5_0),.clk(gclk));
	jdff dff_B_qLRmuQ330_0(.din(w_dff_B_TaqQMqcn5_0),.dout(w_dff_B_qLRmuQ330_0),.clk(gclk));
	jdff dff_B_mRnocC4A3_0(.din(w_dff_B_qLRmuQ330_0),.dout(w_dff_B_mRnocC4A3_0),.clk(gclk));
	jdff dff_B_wNzQNQMS8_0(.din(w_dff_B_mRnocC4A3_0),.dout(w_dff_B_wNzQNQMS8_0),.clk(gclk));
	jdff dff_B_MWtU1QuQ8_0(.din(w_dff_B_wNzQNQMS8_0),.dout(w_dff_B_MWtU1QuQ8_0),.clk(gclk));
	jdff dff_B_VkLYDPww2_0(.din(w_dff_B_MWtU1QuQ8_0),.dout(w_dff_B_VkLYDPww2_0),.clk(gclk));
	jdff dff_B_sZUtHWnX4_0(.din(w_dff_B_VkLYDPww2_0),.dout(w_dff_B_sZUtHWnX4_0),.clk(gclk));
	jdff dff_B_z45pZN5j0_0(.din(w_dff_B_sZUtHWnX4_0),.dout(w_dff_B_z45pZN5j0_0),.clk(gclk));
	jdff dff_B_EA39EuGF6_0(.din(w_dff_B_z45pZN5j0_0),.dout(w_dff_B_EA39EuGF6_0),.clk(gclk));
	jdff dff_B_U0kVPIme6_0(.din(w_dff_B_EA39EuGF6_0),.dout(w_dff_B_U0kVPIme6_0),.clk(gclk));
	jdff dff_B_zX9xjztb5_0(.din(w_dff_B_U0kVPIme6_0),.dout(w_dff_B_zX9xjztb5_0),.clk(gclk));
	jdff dff_B_GwwfIdIG0_0(.din(n778),.dout(w_dff_B_GwwfIdIG0_0),.clk(gclk));
	jdff dff_B_QSc3XySm2_0(.din(w_dff_B_GwwfIdIG0_0),.dout(w_dff_B_QSc3XySm2_0),.clk(gclk));
	jdff dff_B_aOMPMwkk4_0(.din(w_dff_B_QSc3XySm2_0),.dout(w_dff_B_aOMPMwkk4_0),.clk(gclk));
	jdff dff_B_82AmGAYp6_0(.din(w_dff_B_aOMPMwkk4_0),.dout(w_dff_B_82AmGAYp6_0),.clk(gclk));
	jdff dff_B_fO2xFMpA9_0(.din(w_dff_B_82AmGAYp6_0),.dout(w_dff_B_fO2xFMpA9_0),.clk(gclk));
	jdff dff_B_odjCbIQs7_0(.din(w_dff_B_fO2xFMpA9_0),.dout(w_dff_B_odjCbIQs7_0),.clk(gclk));
	jdff dff_B_EK6QoiuF7_0(.din(w_dff_B_odjCbIQs7_0),.dout(w_dff_B_EK6QoiuF7_0),.clk(gclk));
	jdff dff_B_0sPcfCEm5_0(.din(w_dff_B_EK6QoiuF7_0),.dout(w_dff_B_0sPcfCEm5_0),.clk(gclk));
	jdff dff_B_j74OIgf71_0(.din(w_dff_B_0sPcfCEm5_0),.dout(w_dff_B_j74OIgf71_0),.clk(gclk));
	jdff dff_B_giK3ZfKT3_0(.din(w_dff_B_j74OIgf71_0),.dout(w_dff_B_giK3ZfKT3_0),.clk(gclk));
	jdff dff_B_RqpnAtEb0_0(.din(w_dff_B_giK3ZfKT3_0),.dout(w_dff_B_RqpnAtEb0_0),.clk(gclk));
	jdff dff_B_RQQx7A414_0(.din(w_dff_B_RqpnAtEb0_0),.dout(w_dff_B_RQQx7A414_0),.clk(gclk));
	jdff dff_B_SCOroRu62_0(.din(w_dff_B_RQQx7A414_0),.dout(w_dff_B_SCOroRu62_0),.clk(gclk));
	jdff dff_B_2AT6RE5v8_0(.din(w_dff_B_SCOroRu62_0),.dout(w_dff_B_2AT6RE5v8_0),.clk(gclk));
	jdff dff_B_9GLbvQK51_0(.din(w_dff_B_2AT6RE5v8_0),.dout(w_dff_B_9GLbvQK51_0),.clk(gclk));
	jdff dff_B_94ri8je74_0(.din(w_dff_B_9GLbvQK51_0),.dout(w_dff_B_94ri8je74_0),.clk(gclk));
	jdff dff_B_GHsgX6uq7_0(.din(w_dff_B_94ri8je74_0),.dout(w_dff_B_GHsgX6uq7_0),.clk(gclk));
	jdff dff_B_9jQGw9qS3_0(.din(w_dff_B_GHsgX6uq7_0),.dout(w_dff_B_9jQGw9qS3_0),.clk(gclk));
	jdff dff_B_vRSFmdnY9_0(.din(w_dff_B_9jQGw9qS3_0),.dout(w_dff_B_vRSFmdnY9_0),.clk(gclk));
	jdff dff_B_0AFXUI3J1_0(.din(w_dff_B_vRSFmdnY9_0),.dout(w_dff_B_0AFXUI3J1_0),.clk(gclk));
	jdff dff_B_YbThWPGE9_0(.din(w_dff_B_0AFXUI3J1_0),.dout(w_dff_B_YbThWPGE9_0),.clk(gclk));
	jdff dff_B_1JJ7VEFJ3_0(.din(w_dff_B_YbThWPGE9_0),.dout(w_dff_B_1JJ7VEFJ3_0),.clk(gclk));
	jdff dff_B_ph4tuA5o9_0(.din(w_dff_B_1JJ7VEFJ3_0),.dout(w_dff_B_ph4tuA5o9_0),.clk(gclk));
	jdff dff_B_PXzo0FXR5_0(.din(w_dff_B_ph4tuA5o9_0),.dout(w_dff_B_PXzo0FXR5_0),.clk(gclk));
	jdff dff_B_EI6f7HZW0_0(.din(w_dff_B_PXzo0FXR5_0),.dout(w_dff_B_EI6f7HZW0_0),.clk(gclk));
	jdff dff_B_x4x6t1UZ5_0(.din(w_dff_B_EI6f7HZW0_0),.dout(w_dff_B_x4x6t1UZ5_0),.clk(gclk));
	jdff dff_B_WQQyaq1I0_0(.din(w_dff_B_x4x6t1UZ5_0),.dout(w_dff_B_WQQyaq1I0_0),.clk(gclk));
	jdff dff_B_LJlHrdKh4_0(.din(w_dff_B_WQQyaq1I0_0),.dout(w_dff_B_LJlHrdKh4_0),.clk(gclk));
	jdff dff_B_zpJzrBeX1_0(.din(w_dff_B_LJlHrdKh4_0),.dout(w_dff_B_zpJzrBeX1_0),.clk(gclk));
	jdff dff_B_w2OrBOlf7_0(.din(w_dff_B_zpJzrBeX1_0),.dout(w_dff_B_w2OrBOlf7_0),.clk(gclk));
	jdff dff_B_MLPgA7JX5_0(.din(w_dff_B_w2OrBOlf7_0),.dout(w_dff_B_MLPgA7JX5_0),.clk(gclk));
	jdff dff_B_PPrC5dsk9_0(.din(w_dff_B_MLPgA7JX5_0),.dout(w_dff_B_PPrC5dsk9_0),.clk(gclk));
	jdff dff_B_6E3PsTwz7_0(.din(w_dff_B_PPrC5dsk9_0),.dout(w_dff_B_6E3PsTwz7_0),.clk(gclk));
	jdff dff_B_MrDsvF7h6_0(.din(w_dff_B_6E3PsTwz7_0),.dout(w_dff_B_MrDsvF7h6_0),.clk(gclk));
	jdff dff_B_r5NccNIR1_0(.din(w_dff_B_MrDsvF7h6_0),.dout(w_dff_B_r5NccNIR1_0),.clk(gclk));
	jdff dff_B_E4MrUu1v7_0(.din(w_dff_B_r5NccNIR1_0),.dout(w_dff_B_E4MrUu1v7_0),.clk(gclk));
	jdff dff_B_nW1tMMwR7_0(.din(w_dff_B_E4MrUu1v7_0),.dout(w_dff_B_nW1tMMwR7_0),.clk(gclk));
	jdff dff_B_6RU7Wz3s6_0(.din(w_dff_B_nW1tMMwR7_0),.dout(w_dff_B_6RU7Wz3s6_0),.clk(gclk));
	jdff dff_B_FBdmNrEp5_0(.din(w_dff_B_6RU7Wz3s6_0),.dout(w_dff_B_FBdmNrEp5_0),.clk(gclk));
	jdff dff_B_dQqps2ge4_0(.din(w_dff_B_FBdmNrEp5_0),.dout(w_dff_B_dQqps2ge4_0),.clk(gclk));
	jdff dff_B_u9VRLZr66_0(.din(w_dff_B_dQqps2ge4_0),.dout(w_dff_B_u9VRLZr66_0),.clk(gclk));
	jdff dff_B_P5Whr83Q3_0(.din(w_dff_B_u9VRLZr66_0),.dout(w_dff_B_P5Whr83Q3_0),.clk(gclk));
	jdff dff_B_I4nuT0x68_0(.din(w_dff_B_P5Whr83Q3_0),.dout(w_dff_B_I4nuT0x68_0),.clk(gclk));
	jdff dff_B_5BHPhDaZ7_0(.din(w_dff_B_I4nuT0x68_0),.dout(w_dff_B_5BHPhDaZ7_0),.clk(gclk));
	jdff dff_B_NZu8twoZ1_0(.din(w_dff_B_5BHPhDaZ7_0),.dout(w_dff_B_NZu8twoZ1_0),.clk(gclk));
	jdff dff_B_s825yrPp4_0(.din(w_dff_B_NZu8twoZ1_0),.dout(w_dff_B_s825yrPp4_0),.clk(gclk));
	jdff dff_B_Z3uSCLx70_0(.din(w_dff_B_s825yrPp4_0),.dout(w_dff_B_Z3uSCLx70_0),.clk(gclk));
	jdff dff_B_g2A2f35Z6_0(.din(w_dff_B_Z3uSCLx70_0),.dout(w_dff_B_g2A2f35Z6_0),.clk(gclk));
	jdff dff_B_L36zlbqn7_0(.din(w_dff_B_g2A2f35Z6_0),.dout(w_dff_B_L36zlbqn7_0),.clk(gclk));
	jdff dff_B_sFPFdYnj1_0(.din(w_dff_B_L36zlbqn7_0),.dout(w_dff_B_sFPFdYnj1_0),.clk(gclk));
	jdff dff_B_uRJN2Z1S1_0(.din(w_dff_B_sFPFdYnj1_0),.dout(w_dff_B_uRJN2Z1S1_0),.clk(gclk));
	jdff dff_B_UnriJoaA0_0(.din(w_dff_B_uRJN2Z1S1_0),.dout(w_dff_B_UnriJoaA0_0),.clk(gclk));
	jdff dff_B_V1rzDvpI3_0(.din(w_dff_B_UnriJoaA0_0),.dout(w_dff_B_V1rzDvpI3_0),.clk(gclk));
	jdff dff_B_gbFJPRZS9_0(.din(w_dff_B_V1rzDvpI3_0),.dout(w_dff_B_gbFJPRZS9_0),.clk(gclk));
	jdff dff_B_r7owaA1L1_0(.din(w_dff_B_gbFJPRZS9_0),.dout(w_dff_B_r7owaA1L1_0),.clk(gclk));
	jdff dff_B_NfOxH3mi8_0(.din(w_dff_B_r7owaA1L1_0),.dout(w_dff_B_NfOxH3mi8_0),.clk(gclk));
	jdff dff_B_e57zDC3p4_0(.din(w_dff_B_NfOxH3mi8_0),.dout(w_dff_B_e57zDC3p4_0),.clk(gclk));
	jdff dff_B_xiGkzxK49_0(.din(w_dff_B_e57zDC3p4_0),.dout(w_dff_B_xiGkzxK49_0),.clk(gclk));
	jdff dff_B_Jx6Mo8Vf4_0(.din(w_dff_B_xiGkzxK49_0),.dout(w_dff_B_Jx6Mo8Vf4_0),.clk(gclk));
	jdff dff_B_QeyU41Fr2_0(.din(w_dff_B_Jx6Mo8Vf4_0),.dout(w_dff_B_QeyU41Fr2_0),.clk(gclk));
	jdff dff_B_Jo71CWFb7_0(.din(w_dff_B_QeyU41Fr2_0),.dout(w_dff_B_Jo71CWFb7_0),.clk(gclk));
	jdff dff_B_NMNHRPtb6_0(.din(w_dff_B_Jo71CWFb7_0),.dout(w_dff_B_NMNHRPtb6_0),.clk(gclk));
	jdff dff_B_lZIL4XvH3_0(.din(w_dff_B_NMNHRPtb6_0),.dout(w_dff_B_lZIL4XvH3_0),.clk(gclk));
	jdff dff_B_NQkDBRaw2_0(.din(w_dff_B_lZIL4XvH3_0),.dout(w_dff_B_NQkDBRaw2_0),.clk(gclk));
	jdff dff_B_wTQtsp8q0_0(.din(w_dff_B_NQkDBRaw2_0),.dout(w_dff_B_wTQtsp8q0_0),.clk(gclk));
	jdff dff_B_FD61d4J13_0(.din(n784),.dout(w_dff_B_FD61d4J13_0),.clk(gclk));
	jdff dff_B_xH71X5T02_0(.din(w_dff_B_FD61d4J13_0),.dout(w_dff_B_xH71X5T02_0),.clk(gclk));
	jdff dff_B_iOAzKUIi9_0(.din(w_dff_B_xH71X5T02_0),.dout(w_dff_B_iOAzKUIi9_0),.clk(gclk));
	jdff dff_B_mSkku9xs7_0(.din(w_dff_B_iOAzKUIi9_0),.dout(w_dff_B_mSkku9xs7_0),.clk(gclk));
	jdff dff_B_AvPJCngU7_0(.din(w_dff_B_mSkku9xs7_0),.dout(w_dff_B_AvPJCngU7_0),.clk(gclk));
	jdff dff_B_yX0J0icS5_0(.din(w_dff_B_AvPJCngU7_0),.dout(w_dff_B_yX0J0icS5_0),.clk(gclk));
	jdff dff_B_a6NzBdXb7_0(.din(w_dff_B_yX0J0icS5_0),.dout(w_dff_B_a6NzBdXb7_0),.clk(gclk));
	jdff dff_B_HdgOaw0K7_0(.din(w_dff_B_a6NzBdXb7_0),.dout(w_dff_B_HdgOaw0K7_0),.clk(gclk));
	jdff dff_B_FEODvdGk4_0(.din(w_dff_B_HdgOaw0K7_0),.dout(w_dff_B_FEODvdGk4_0),.clk(gclk));
	jdff dff_B_FWlKx7Og0_0(.din(w_dff_B_FEODvdGk4_0),.dout(w_dff_B_FWlKx7Og0_0),.clk(gclk));
	jdff dff_B_oksCqqwa4_0(.din(w_dff_B_FWlKx7Og0_0),.dout(w_dff_B_oksCqqwa4_0),.clk(gclk));
	jdff dff_B_FCNovqwK4_0(.din(w_dff_B_oksCqqwa4_0),.dout(w_dff_B_FCNovqwK4_0),.clk(gclk));
	jdff dff_B_pCzqQPjj4_0(.din(w_dff_B_FCNovqwK4_0),.dout(w_dff_B_pCzqQPjj4_0),.clk(gclk));
	jdff dff_B_20WcSLIP3_0(.din(w_dff_B_pCzqQPjj4_0),.dout(w_dff_B_20WcSLIP3_0),.clk(gclk));
	jdff dff_B_h46I3nSG5_0(.din(w_dff_B_20WcSLIP3_0),.dout(w_dff_B_h46I3nSG5_0),.clk(gclk));
	jdff dff_B_gFNBuQyl4_0(.din(w_dff_B_h46I3nSG5_0),.dout(w_dff_B_gFNBuQyl4_0),.clk(gclk));
	jdff dff_B_vqACgTsP6_0(.din(w_dff_B_gFNBuQyl4_0),.dout(w_dff_B_vqACgTsP6_0),.clk(gclk));
	jdff dff_B_ifVNfQGj9_0(.din(w_dff_B_vqACgTsP6_0),.dout(w_dff_B_ifVNfQGj9_0),.clk(gclk));
	jdff dff_B_b1SK9OI79_0(.din(w_dff_B_ifVNfQGj9_0),.dout(w_dff_B_b1SK9OI79_0),.clk(gclk));
	jdff dff_B_aXx2AjZE0_0(.din(w_dff_B_b1SK9OI79_0),.dout(w_dff_B_aXx2AjZE0_0),.clk(gclk));
	jdff dff_B_ISKEB67Q8_0(.din(w_dff_B_aXx2AjZE0_0),.dout(w_dff_B_ISKEB67Q8_0),.clk(gclk));
	jdff dff_B_rkRCeR1a7_0(.din(w_dff_B_ISKEB67Q8_0),.dout(w_dff_B_rkRCeR1a7_0),.clk(gclk));
	jdff dff_B_xW2c1SZ52_0(.din(w_dff_B_rkRCeR1a7_0),.dout(w_dff_B_xW2c1SZ52_0),.clk(gclk));
	jdff dff_B_nf3ri1wv4_0(.din(w_dff_B_xW2c1SZ52_0),.dout(w_dff_B_nf3ri1wv4_0),.clk(gclk));
	jdff dff_B_vF8SRzO08_0(.din(w_dff_B_nf3ri1wv4_0),.dout(w_dff_B_vF8SRzO08_0),.clk(gclk));
	jdff dff_B_Ib2y6we34_0(.din(w_dff_B_vF8SRzO08_0),.dout(w_dff_B_Ib2y6we34_0),.clk(gclk));
	jdff dff_B_qnn6UrAm7_0(.din(w_dff_B_Ib2y6we34_0),.dout(w_dff_B_qnn6UrAm7_0),.clk(gclk));
	jdff dff_B_1Va83HTI3_0(.din(w_dff_B_qnn6UrAm7_0),.dout(w_dff_B_1Va83HTI3_0),.clk(gclk));
	jdff dff_B_m1DBBFnk4_0(.din(w_dff_B_1Va83HTI3_0),.dout(w_dff_B_m1DBBFnk4_0),.clk(gclk));
	jdff dff_B_JePJUlNE8_0(.din(w_dff_B_m1DBBFnk4_0),.dout(w_dff_B_JePJUlNE8_0),.clk(gclk));
	jdff dff_B_paCFAH7p6_0(.din(w_dff_B_JePJUlNE8_0),.dout(w_dff_B_paCFAH7p6_0),.clk(gclk));
	jdff dff_B_ZyYlB3Gf4_0(.din(w_dff_B_paCFAH7p6_0),.dout(w_dff_B_ZyYlB3Gf4_0),.clk(gclk));
	jdff dff_B_BL0604YI1_0(.din(w_dff_B_ZyYlB3Gf4_0),.dout(w_dff_B_BL0604YI1_0),.clk(gclk));
	jdff dff_B_wQwXiO6k4_0(.din(w_dff_B_BL0604YI1_0),.dout(w_dff_B_wQwXiO6k4_0),.clk(gclk));
	jdff dff_B_mOc2EWeS7_0(.din(w_dff_B_wQwXiO6k4_0),.dout(w_dff_B_mOc2EWeS7_0),.clk(gclk));
	jdff dff_B_qg03r9Uq4_0(.din(w_dff_B_mOc2EWeS7_0),.dout(w_dff_B_qg03r9Uq4_0),.clk(gclk));
	jdff dff_B_dEPqaaQ91_0(.din(w_dff_B_qg03r9Uq4_0),.dout(w_dff_B_dEPqaaQ91_0),.clk(gclk));
	jdff dff_B_amyu1Ebk7_0(.din(w_dff_B_dEPqaaQ91_0),.dout(w_dff_B_amyu1Ebk7_0),.clk(gclk));
	jdff dff_B_oAZR17Pe4_0(.din(w_dff_B_amyu1Ebk7_0),.dout(w_dff_B_oAZR17Pe4_0),.clk(gclk));
	jdff dff_B_sXxPyr587_0(.din(w_dff_B_oAZR17Pe4_0),.dout(w_dff_B_sXxPyr587_0),.clk(gclk));
	jdff dff_B_K6HNtwHg0_0(.din(w_dff_B_sXxPyr587_0),.dout(w_dff_B_K6HNtwHg0_0),.clk(gclk));
	jdff dff_B_3orl7EEY8_0(.din(w_dff_B_K6HNtwHg0_0),.dout(w_dff_B_3orl7EEY8_0),.clk(gclk));
	jdff dff_B_1YlJJ1RB6_0(.din(w_dff_B_3orl7EEY8_0),.dout(w_dff_B_1YlJJ1RB6_0),.clk(gclk));
	jdff dff_B_H4NY58EE0_0(.din(w_dff_B_1YlJJ1RB6_0),.dout(w_dff_B_H4NY58EE0_0),.clk(gclk));
	jdff dff_B_4mHE5FKx4_0(.din(w_dff_B_H4NY58EE0_0),.dout(w_dff_B_4mHE5FKx4_0),.clk(gclk));
	jdff dff_B_YYw0Pgyg2_0(.din(w_dff_B_4mHE5FKx4_0),.dout(w_dff_B_YYw0Pgyg2_0),.clk(gclk));
	jdff dff_B_Y9kCUqXx3_0(.din(w_dff_B_YYw0Pgyg2_0),.dout(w_dff_B_Y9kCUqXx3_0),.clk(gclk));
	jdff dff_B_Sm7os6q54_0(.din(w_dff_B_Y9kCUqXx3_0),.dout(w_dff_B_Sm7os6q54_0),.clk(gclk));
	jdff dff_B_XYV59m5b6_0(.din(w_dff_B_Sm7os6q54_0),.dout(w_dff_B_XYV59m5b6_0),.clk(gclk));
	jdff dff_B_vTZyJmn24_0(.din(w_dff_B_XYV59m5b6_0),.dout(w_dff_B_vTZyJmn24_0),.clk(gclk));
	jdff dff_B_qh3LR3EW9_0(.din(w_dff_B_vTZyJmn24_0),.dout(w_dff_B_qh3LR3EW9_0),.clk(gclk));
	jdff dff_B_IBTJoY8s3_0(.din(w_dff_B_qh3LR3EW9_0),.dout(w_dff_B_IBTJoY8s3_0),.clk(gclk));
	jdff dff_B_iYBVjVoJ2_0(.din(w_dff_B_IBTJoY8s3_0),.dout(w_dff_B_iYBVjVoJ2_0),.clk(gclk));
	jdff dff_B_MQB8pzWu9_0(.din(w_dff_B_iYBVjVoJ2_0),.dout(w_dff_B_MQB8pzWu9_0),.clk(gclk));
	jdff dff_B_7Irxwdwa3_0(.din(w_dff_B_MQB8pzWu9_0),.dout(w_dff_B_7Irxwdwa3_0),.clk(gclk));
	jdff dff_B_A4gxXYeT5_0(.din(w_dff_B_7Irxwdwa3_0),.dout(w_dff_B_A4gxXYeT5_0),.clk(gclk));
	jdff dff_B_L5vEnBCe4_0(.din(w_dff_B_A4gxXYeT5_0),.dout(w_dff_B_L5vEnBCe4_0),.clk(gclk));
	jdff dff_B_kjqlBjnP7_0(.din(w_dff_B_L5vEnBCe4_0),.dout(w_dff_B_kjqlBjnP7_0),.clk(gclk));
	jdff dff_B_kdk7rieD3_0(.din(w_dff_B_kjqlBjnP7_0),.dout(w_dff_B_kdk7rieD3_0),.clk(gclk));
	jdff dff_B_pz4y5f0W1_0(.din(w_dff_B_kdk7rieD3_0),.dout(w_dff_B_pz4y5f0W1_0),.clk(gclk));
	jdff dff_B_nFSDgmgh7_0(.din(w_dff_B_pz4y5f0W1_0),.dout(w_dff_B_nFSDgmgh7_0),.clk(gclk));
	jdff dff_B_Ln5O11LD0_0(.din(w_dff_B_nFSDgmgh7_0),.dout(w_dff_B_Ln5O11LD0_0),.clk(gclk));
	jdff dff_B_gMj7s1Qq5_0(.din(w_dff_B_Ln5O11LD0_0),.dout(w_dff_B_gMj7s1Qq5_0),.clk(gclk));
	jdff dff_B_AOs9NUAK2_0(.din(w_dff_B_gMj7s1Qq5_0),.dout(w_dff_B_AOs9NUAK2_0),.clk(gclk));
	jdff dff_B_KqZIl82N4_0(.din(w_dff_B_AOs9NUAK2_0),.dout(w_dff_B_KqZIl82N4_0),.clk(gclk));
	jdff dff_B_lE4zQQav5_0(.din(w_dff_B_KqZIl82N4_0),.dout(w_dff_B_lE4zQQav5_0),.clk(gclk));
	jdff dff_B_4R5fXsur6_0(.din(n790),.dout(w_dff_B_4R5fXsur6_0),.clk(gclk));
	jdff dff_B_Xwf8NQiK3_0(.din(w_dff_B_4R5fXsur6_0),.dout(w_dff_B_Xwf8NQiK3_0),.clk(gclk));
	jdff dff_B_INcZZ9du1_0(.din(w_dff_B_Xwf8NQiK3_0),.dout(w_dff_B_INcZZ9du1_0),.clk(gclk));
	jdff dff_B_0ukkx5i97_0(.din(w_dff_B_INcZZ9du1_0),.dout(w_dff_B_0ukkx5i97_0),.clk(gclk));
	jdff dff_B_ejEwZdAO5_0(.din(w_dff_B_0ukkx5i97_0),.dout(w_dff_B_ejEwZdAO5_0),.clk(gclk));
	jdff dff_B_gNkqF7ye2_0(.din(w_dff_B_ejEwZdAO5_0),.dout(w_dff_B_gNkqF7ye2_0),.clk(gclk));
	jdff dff_B_lOExTQCk0_0(.din(w_dff_B_gNkqF7ye2_0),.dout(w_dff_B_lOExTQCk0_0),.clk(gclk));
	jdff dff_B_8ilnO7ao2_0(.din(w_dff_B_lOExTQCk0_0),.dout(w_dff_B_8ilnO7ao2_0),.clk(gclk));
	jdff dff_B_mNhv8NzT0_0(.din(w_dff_B_8ilnO7ao2_0),.dout(w_dff_B_mNhv8NzT0_0),.clk(gclk));
	jdff dff_B_Vhsm7z3k9_0(.din(w_dff_B_mNhv8NzT0_0),.dout(w_dff_B_Vhsm7z3k9_0),.clk(gclk));
	jdff dff_B_x1ZgcNBL8_0(.din(w_dff_B_Vhsm7z3k9_0),.dout(w_dff_B_x1ZgcNBL8_0),.clk(gclk));
	jdff dff_B_785CZbJD3_0(.din(w_dff_B_x1ZgcNBL8_0),.dout(w_dff_B_785CZbJD3_0),.clk(gclk));
	jdff dff_B_NHxNd3fE4_0(.din(w_dff_B_785CZbJD3_0),.dout(w_dff_B_NHxNd3fE4_0),.clk(gclk));
	jdff dff_B_6oGj6A9X9_0(.din(w_dff_B_NHxNd3fE4_0),.dout(w_dff_B_6oGj6A9X9_0),.clk(gclk));
	jdff dff_B_6Ijlp6QV7_0(.din(w_dff_B_6oGj6A9X9_0),.dout(w_dff_B_6Ijlp6QV7_0),.clk(gclk));
	jdff dff_B_mJqkvpO50_0(.din(w_dff_B_6Ijlp6QV7_0),.dout(w_dff_B_mJqkvpO50_0),.clk(gclk));
	jdff dff_B_RyDPoz1Z2_0(.din(w_dff_B_mJqkvpO50_0),.dout(w_dff_B_RyDPoz1Z2_0),.clk(gclk));
	jdff dff_B_EXwwDbRq0_0(.din(w_dff_B_RyDPoz1Z2_0),.dout(w_dff_B_EXwwDbRq0_0),.clk(gclk));
	jdff dff_B_CUGELkob2_0(.din(w_dff_B_EXwwDbRq0_0),.dout(w_dff_B_CUGELkob2_0),.clk(gclk));
	jdff dff_B_5JXuxMkZ1_0(.din(w_dff_B_CUGELkob2_0),.dout(w_dff_B_5JXuxMkZ1_0),.clk(gclk));
	jdff dff_B_yelkp9xh3_0(.din(w_dff_B_5JXuxMkZ1_0),.dout(w_dff_B_yelkp9xh3_0),.clk(gclk));
	jdff dff_B_MpLxlKvI0_0(.din(w_dff_B_yelkp9xh3_0),.dout(w_dff_B_MpLxlKvI0_0),.clk(gclk));
	jdff dff_B_93Ub34Fw2_0(.din(w_dff_B_MpLxlKvI0_0),.dout(w_dff_B_93Ub34Fw2_0),.clk(gclk));
	jdff dff_B_kNmC3KVP8_0(.din(w_dff_B_93Ub34Fw2_0),.dout(w_dff_B_kNmC3KVP8_0),.clk(gclk));
	jdff dff_B_jZUSvEo03_0(.din(w_dff_B_kNmC3KVP8_0),.dout(w_dff_B_jZUSvEo03_0),.clk(gclk));
	jdff dff_B_twT26NLx5_0(.din(w_dff_B_jZUSvEo03_0),.dout(w_dff_B_twT26NLx5_0),.clk(gclk));
	jdff dff_B_ryAdrR3U8_0(.din(w_dff_B_twT26NLx5_0),.dout(w_dff_B_ryAdrR3U8_0),.clk(gclk));
	jdff dff_B_LnB9CBWC3_0(.din(w_dff_B_ryAdrR3U8_0),.dout(w_dff_B_LnB9CBWC3_0),.clk(gclk));
	jdff dff_B_1eFl5wzJ7_0(.din(w_dff_B_LnB9CBWC3_0),.dout(w_dff_B_1eFl5wzJ7_0),.clk(gclk));
	jdff dff_B_rTyNG8fO2_0(.din(w_dff_B_1eFl5wzJ7_0),.dout(w_dff_B_rTyNG8fO2_0),.clk(gclk));
	jdff dff_B_sGmwp9Yw9_0(.din(w_dff_B_rTyNG8fO2_0),.dout(w_dff_B_sGmwp9Yw9_0),.clk(gclk));
	jdff dff_B_A7pKB0Tb8_0(.din(w_dff_B_sGmwp9Yw9_0),.dout(w_dff_B_A7pKB0Tb8_0),.clk(gclk));
	jdff dff_B_BvXOgf6L3_0(.din(w_dff_B_A7pKB0Tb8_0),.dout(w_dff_B_BvXOgf6L3_0),.clk(gclk));
	jdff dff_B_MKfbWAlu6_0(.din(w_dff_B_BvXOgf6L3_0),.dout(w_dff_B_MKfbWAlu6_0),.clk(gclk));
	jdff dff_B_7rcRnx1W1_0(.din(w_dff_B_MKfbWAlu6_0),.dout(w_dff_B_7rcRnx1W1_0),.clk(gclk));
	jdff dff_B_cYQt0Qi32_0(.din(w_dff_B_7rcRnx1W1_0),.dout(w_dff_B_cYQt0Qi32_0),.clk(gclk));
	jdff dff_B_06iSBwe46_0(.din(w_dff_B_cYQt0Qi32_0),.dout(w_dff_B_06iSBwe46_0),.clk(gclk));
	jdff dff_B_wGijM75C1_0(.din(w_dff_B_06iSBwe46_0),.dout(w_dff_B_wGijM75C1_0),.clk(gclk));
	jdff dff_B_coNrT10v9_0(.din(w_dff_B_wGijM75C1_0),.dout(w_dff_B_coNrT10v9_0),.clk(gclk));
	jdff dff_B_uQ2KjSqG9_0(.din(w_dff_B_coNrT10v9_0),.dout(w_dff_B_uQ2KjSqG9_0),.clk(gclk));
	jdff dff_B_cnhrdf764_0(.din(w_dff_B_uQ2KjSqG9_0),.dout(w_dff_B_cnhrdf764_0),.clk(gclk));
	jdff dff_B_FVmLi4Tc9_0(.din(w_dff_B_cnhrdf764_0),.dout(w_dff_B_FVmLi4Tc9_0),.clk(gclk));
	jdff dff_B_Sa0d1qbJ5_0(.din(w_dff_B_FVmLi4Tc9_0),.dout(w_dff_B_Sa0d1qbJ5_0),.clk(gclk));
	jdff dff_B_7Ks559YV4_0(.din(w_dff_B_Sa0d1qbJ5_0),.dout(w_dff_B_7Ks559YV4_0),.clk(gclk));
	jdff dff_B_xGLWstaY9_0(.din(w_dff_B_7Ks559YV4_0),.dout(w_dff_B_xGLWstaY9_0),.clk(gclk));
	jdff dff_B_QpfvsARL4_0(.din(w_dff_B_xGLWstaY9_0),.dout(w_dff_B_QpfvsARL4_0),.clk(gclk));
	jdff dff_B_30CG8MC89_0(.din(w_dff_B_QpfvsARL4_0),.dout(w_dff_B_30CG8MC89_0),.clk(gclk));
	jdff dff_B_9nZW4qVC2_0(.din(w_dff_B_30CG8MC89_0),.dout(w_dff_B_9nZW4qVC2_0),.clk(gclk));
	jdff dff_B_UcgqJ7WF3_0(.din(w_dff_B_9nZW4qVC2_0),.dout(w_dff_B_UcgqJ7WF3_0),.clk(gclk));
	jdff dff_B_KA9jg2v29_0(.din(w_dff_B_UcgqJ7WF3_0),.dout(w_dff_B_KA9jg2v29_0),.clk(gclk));
	jdff dff_B_YTgPN8Ci2_0(.din(w_dff_B_KA9jg2v29_0),.dout(w_dff_B_YTgPN8Ci2_0),.clk(gclk));
	jdff dff_B_iSPnGKGf4_0(.din(w_dff_B_YTgPN8Ci2_0),.dout(w_dff_B_iSPnGKGf4_0),.clk(gclk));
	jdff dff_B_kZjuT8B68_0(.din(w_dff_B_iSPnGKGf4_0),.dout(w_dff_B_kZjuT8B68_0),.clk(gclk));
	jdff dff_B_nr9LvYBe1_0(.din(w_dff_B_kZjuT8B68_0),.dout(w_dff_B_nr9LvYBe1_0),.clk(gclk));
	jdff dff_B_17IgJkoN9_0(.din(w_dff_B_nr9LvYBe1_0),.dout(w_dff_B_17IgJkoN9_0),.clk(gclk));
	jdff dff_B_LKs6pDE20_0(.din(w_dff_B_17IgJkoN9_0),.dout(w_dff_B_LKs6pDE20_0),.clk(gclk));
	jdff dff_B_e08V3hhG5_0(.din(w_dff_B_LKs6pDE20_0),.dout(w_dff_B_e08V3hhG5_0),.clk(gclk));
	jdff dff_B_ODV3X2tf2_0(.din(w_dff_B_e08V3hhG5_0),.dout(w_dff_B_ODV3X2tf2_0),.clk(gclk));
	jdff dff_B_7jqXSN8o0_0(.din(w_dff_B_ODV3X2tf2_0),.dout(w_dff_B_7jqXSN8o0_0),.clk(gclk));
	jdff dff_B_zO1C5J2N3_0(.din(w_dff_B_7jqXSN8o0_0),.dout(w_dff_B_zO1C5J2N3_0),.clk(gclk));
	jdff dff_B_5vNkDRPz1_0(.din(w_dff_B_zO1C5J2N3_0),.dout(w_dff_B_5vNkDRPz1_0),.clk(gclk));
	jdff dff_B_yTDKng3N9_0(.din(w_dff_B_5vNkDRPz1_0),.dout(w_dff_B_yTDKng3N9_0),.clk(gclk));
	jdff dff_B_gbTIqg2C1_0(.din(w_dff_B_yTDKng3N9_0),.dout(w_dff_B_gbTIqg2C1_0),.clk(gclk));
	jdff dff_B_CgfxH41a9_0(.din(w_dff_B_gbTIqg2C1_0),.dout(w_dff_B_CgfxH41a9_0),.clk(gclk));
	jdff dff_B_UW3Tmxwx5_0(.din(w_dff_B_CgfxH41a9_0),.dout(w_dff_B_UW3Tmxwx5_0),.clk(gclk));
	jdff dff_B_dAhtKta17_0(.din(w_dff_B_UW3Tmxwx5_0),.dout(w_dff_B_dAhtKta17_0),.clk(gclk));
	jdff dff_B_svBcB5FP3_0(.din(w_dff_B_dAhtKta17_0),.dout(w_dff_B_svBcB5FP3_0),.clk(gclk));
	jdff dff_B_VggTW5wC8_0(.din(n796),.dout(w_dff_B_VggTW5wC8_0),.clk(gclk));
	jdff dff_B_aHBEsBAV9_0(.din(w_dff_B_VggTW5wC8_0),.dout(w_dff_B_aHBEsBAV9_0),.clk(gclk));
	jdff dff_B_W2ekGea47_0(.din(w_dff_B_aHBEsBAV9_0),.dout(w_dff_B_W2ekGea47_0),.clk(gclk));
	jdff dff_B_pxRZbaAB5_0(.din(w_dff_B_W2ekGea47_0),.dout(w_dff_B_pxRZbaAB5_0),.clk(gclk));
	jdff dff_B_qKzm8EVx0_0(.din(w_dff_B_pxRZbaAB5_0),.dout(w_dff_B_qKzm8EVx0_0),.clk(gclk));
	jdff dff_B_FyKgAO4j8_0(.din(w_dff_B_qKzm8EVx0_0),.dout(w_dff_B_FyKgAO4j8_0),.clk(gclk));
	jdff dff_B_0al3Uir41_0(.din(w_dff_B_FyKgAO4j8_0),.dout(w_dff_B_0al3Uir41_0),.clk(gclk));
	jdff dff_B_U8CT8aKb0_0(.din(w_dff_B_0al3Uir41_0),.dout(w_dff_B_U8CT8aKb0_0),.clk(gclk));
	jdff dff_B_dwLqq59T8_0(.din(w_dff_B_U8CT8aKb0_0),.dout(w_dff_B_dwLqq59T8_0),.clk(gclk));
	jdff dff_B_16sBN8mU4_0(.din(w_dff_B_dwLqq59T8_0),.dout(w_dff_B_16sBN8mU4_0),.clk(gclk));
	jdff dff_B_wIM70Lt96_0(.din(w_dff_B_16sBN8mU4_0),.dout(w_dff_B_wIM70Lt96_0),.clk(gclk));
	jdff dff_B_2Aa4akjp1_0(.din(w_dff_B_wIM70Lt96_0),.dout(w_dff_B_2Aa4akjp1_0),.clk(gclk));
	jdff dff_B_IZLRc0Zq7_0(.din(w_dff_B_2Aa4akjp1_0),.dout(w_dff_B_IZLRc0Zq7_0),.clk(gclk));
	jdff dff_B_GeiaIhpB2_0(.din(w_dff_B_IZLRc0Zq7_0),.dout(w_dff_B_GeiaIhpB2_0),.clk(gclk));
	jdff dff_B_uTtxsdDb0_0(.din(w_dff_B_GeiaIhpB2_0),.dout(w_dff_B_uTtxsdDb0_0),.clk(gclk));
	jdff dff_B_YZ8kRwrG8_0(.din(w_dff_B_uTtxsdDb0_0),.dout(w_dff_B_YZ8kRwrG8_0),.clk(gclk));
	jdff dff_B_bjK1uvg36_0(.din(w_dff_B_YZ8kRwrG8_0),.dout(w_dff_B_bjK1uvg36_0),.clk(gclk));
	jdff dff_B_Vm1jp9ST2_0(.din(w_dff_B_bjK1uvg36_0),.dout(w_dff_B_Vm1jp9ST2_0),.clk(gclk));
	jdff dff_B_1Xpydz3R9_0(.din(w_dff_B_Vm1jp9ST2_0),.dout(w_dff_B_1Xpydz3R9_0),.clk(gclk));
	jdff dff_B_dIqU6Kl59_0(.din(w_dff_B_1Xpydz3R9_0),.dout(w_dff_B_dIqU6Kl59_0),.clk(gclk));
	jdff dff_B_DDZo36eF4_0(.din(w_dff_B_dIqU6Kl59_0),.dout(w_dff_B_DDZo36eF4_0),.clk(gclk));
	jdff dff_B_93bkhjsh6_0(.din(w_dff_B_DDZo36eF4_0),.dout(w_dff_B_93bkhjsh6_0),.clk(gclk));
	jdff dff_B_YDXpRDLc6_0(.din(w_dff_B_93bkhjsh6_0),.dout(w_dff_B_YDXpRDLc6_0),.clk(gclk));
	jdff dff_B_dkeCP9wb0_0(.din(w_dff_B_YDXpRDLc6_0),.dout(w_dff_B_dkeCP9wb0_0),.clk(gclk));
	jdff dff_B_IDIdyPVW1_0(.din(w_dff_B_dkeCP9wb0_0),.dout(w_dff_B_IDIdyPVW1_0),.clk(gclk));
	jdff dff_B_oBtENBKi1_0(.din(w_dff_B_IDIdyPVW1_0),.dout(w_dff_B_oBtENBKi1_0),.clk(gclk));
	jdff dff_B_ukpxhzIT7_0(.din(w_dff_B_oBtENBKi1_0),.dout(w_dff_B_ukpxhzIT7_0),.clk(gclk));
	jdff dff_B_ZLlHEj7f4_0(.din(w_dff_B_ukpxhzIT7_0),.dout(w_dff_B_ZLlHEj7f4_0),.clk(gclk));
	jdff dff_B_cCMrRsyB5_0(.din(w_dff_B_ZLlHEj7f4_0),.dout(w_dff_B_cCMrRsyB5_0),.clk(gclk));
	jdff dff_B_BHgpK55x7_0(.din(w_dff_B_cCMrRsyB5_0),.dout(w_dff_B_BHgpK55x7_0),.clk(gclk));
	jdff dff_B_ahjKWMYI8_0(.din(w_dff_B_BHgpK55x7_0),.dout(w_dff_B_ahjKWMYI8_0),.clk(gclk));
	jdff dff_B_ah2lFrXF4_0(.din(w_dff_B_ahjKWMYI8_0),.dout(w_dff_B_ah2lFrXF4_0),.clk(gclk));
	jdff dff_B_funlZuGw9_0(.din(w_dff_B_ah2lFrXF4_0),.dout(w_dff_B_funlZuGw9_0),.clk(gclk));
	jdff dff_B_vmV8GutO0_0(.din(w_dff_B_funlZuGw9_0),.dout(w_dff_B_vmV8GutO0_0),.clk(gclk));
	jdff dff_B_CxiPEjsM7_0(.din(w_dff_B_vmV8GutO0_0),.dout(w_dff_B_CxiPEjsM7_0),.clk(gclk));
	jdff dff_B_UqH2Lvhu9_0(.din(w_dff_B_CxiPEjsM7_0),.dout(w_dff_B_UqH2Lvhu9_0),.clk(gclk));
	jdff dff_B_tegk8IxO0_0(.din(w_dff_B_UqH2Lvhu9_0),.dout(w_dff_B_tegk8IxO0_0),.clk(gclk));
	jdff dff_B_MfhyKy4s5_0(.din(w_dff_B_tegk8IxO0_0),.dout(w_dff_B_MfhyKy4s5_0),.clk(gclk));
	jdff dff_B_USIgyRKd7_0(.din(w_dff_B_MfhyKy4s5_0),.dout(w_dff_B_USIgyRKd7_0),.clk(gclk));
	jdff dff_B_TAMcDs7j9_0(.din(w_dff_B_USIgyRKd7_0),.dout(w_dff_B_TAMcDs7j9_0),.clk(gclk));
	jdff dff_B_QmzSZcRl3_0(.din(w_dff_B_TAMcDs7j9_0),.dout(w_dff_B_QmzSZcRl3_0),.clk(gclk));
	jdff dff_B_YNSKKBuA8_0(.din(w_dff_B_QmzSZcRl3_0),.dout(w_dff_B_YNSKKBuA8_0),.clk(gclk));
	jdff dff_B_zoZMDuln1_0(.din(w_dff_B_YNSKKBuA8_0),.dout(w_dff_B_zoZMDuln1_0),.clk(gclk));
	jdff dff_B_nuJIspEI8_0(.din(w_dff_B_zoZMDuln1_0),.dout(w_dff_B_nuJIspEI8_0),.clk(gclk));
	jdff dff_B_QvridlxU4_0(.din(w_dff_B_nuJIspEI8_0),.dout(w_dff_B_QvridlxU4_0),.clk(gclk));
	jdff dff_B_21WICGu52_0(.din(w_dff_B_QvridlxU4_0),.dout(w_dff_B_21WICGu52_0),.clk(gclk));
	jdff dff_B_4envusfo1_0(.din(w_dff_B_21WICGu52_0),.dout(w_dff_B_4envusfo1_0),.clk(gclk));
	jdff dff_B_QDFODqXv1_0(.din(w_dff_B_4envusfo1_0),.dout(w_dff_B_QDFODqXv1_0),.clk(gclk));
	jdff dff_B_5UXlMKaV7_0(.din(w_dff_B_QDFODqXv1_0),.dout(w_dff_B_5UXlMKaV7_0),.clk(gclk));
	jdff dff_B_syJO6H2N9_0(.din(w_dff_B_5UXlMKaV7_0),.dout(w_dff_B_syJO6H2N9_0),.clk(gclk));
	jdff dff_B_DlFk9U231_0(.din(w_dff_B_syJO6H2N9_0),.dout(w_dff_B_DlFk9U231_0),.clk(gclk));
	jdff dff_B_zOsfWOV19_0(.din(w_dff_B_DlFk9U231_0),.dout(w_dff_B_zOsfWOV19_0),.clk(gclk));
	jdff dff_B_8L6EIg5Q0_0(.din(w_dff_B_zOsfWOV19_0),.dout(w_dff_B_8L6EIg5Q0_0),.clk(gclk));
	jdff dff_B_mNOH6bvL0_0(.din(w_dff_B_8L6EIg5Q0_0),.dout(w_dff_B_mNOH6bvL0_0),.clk(gclk));
	jdff dff_B_X6r5gaHs0_0(.din(w_dff_B_mNOH6bvL0_0),.dout(w_dff_B_X6r5gaHs0_0),.clk(gclk));
	jdff dff_B_ay0f40Es1_0(.din(w_dff_B_X6r5gaHs0_0),.dout(w_dff_B_ay0f40Es1_0),.clk(gclk));
	jdff dff_B_aZdeldrI2_0(.din(w_dff_B_ay0f40Es1_0),.dout(w_dff_B_aZdeldrI2_0),.clk(gclk));
	jdff dff_B_4GGAXCGb2_0(.din(w_dff_B_aZdeldrI2_0),.dout(w_dff_B_4GGAXCGb2_0),.clk(gclk));
	jdff dff_B_cCak4lRB8_0(.din(w_dff_B_4GGAXCGb2_0),.dout(w_dff_B_cCak4lRB8_0),.clk(gclk));
	jdff dff_B_kY4vkloa9_0(.din(w_dff_B_cCak4lRB8_0),.dout(w_dff_B_kY4vkloa9_0),.clk(gclk));
	jdff dff_B_c1mXWdsp9_0(.din(w_dff_B_kY4vkloa9_0),.dout(w_dff_B_c1mXWdsp9_0),.clk(gclk));
	jdff dff_B_f4L9FMuC6_0(.din(w_dff_B_c1mXWdsp9_0),.dout(w_dff_B_f4L9FMuC6_0),.clk(gclk));
	jdff dff_B_QrX5sXIn5_0(.din(w_dff_B_f4L9FMuC6_0),.dout(w_dff_B_QrX5sXIn5_0),.clk(gclk));
	jdff dff_B_sLEE0XhA0_0(.din(w_dff_B_QrX5sXIn5_0),.dout(w_dff_B_sLEE0XhA0_0),.clk(gclk));
	jdff dff_B_YTVe0hl81_0(.din(w_dff_B_sLEE0XhA0_0),.dout(w_dff_B_YTVe0hl81_0),.clk(gclk));
	jdff dff_B_K7FBMU0B7_0(.din(w_dff_B_YTVe0hl81_0),.dout(w_dff_B_K7FBMU0B7_0),.clk(gclk));
	jdff dff_B_Kh1u1Frr8_0(.din(w_dff_B_K7FBMU0B7_0),.dout(w_dff_B_Kh1u1Frr8_0),.clk(gclk));
	jdff dff_B_IIZIbszu3_0(.din(w_dff_B_Kh1u1Frr8_0),.dout(w_dff_B_IIZIbszu3_0),.clk(gclk));
	jdff dff_B_0OENEO1i0_0(.din(n802),.dout(w_dff_B_0OENEO1i0_0),.clk(gclk));
	jdff dff_B_nMUnz0Bg4_0(.din(w_dff_B_0OENEO1i0_0),.dout(w_dff_B_nMUnz0Bg4_0),.clk(gclk));
	jdff dff_B_OeAAUGJF9_0(.din(w_dff_B_nMUnz0Bg4_0),.dout(w_dff_B_OeAAUGJF9_0),.clk(gclk));
	jdff dff_B_DjvEXiK80_0(.din(w_dff_B_OeAAUGJF9_0),.dout(w_dff_B_DjvEXiK80_0),.clk(gclk));
	jdff dff_B_xn03Z1tL1_0(.din(w_dff_B_DjvEXiK80_0),.dout(w_dff_B_xn03Z1tL1_0),.clk(gclk));
	jdff dff_B_QJLoltAD1_0(.din(w_dff_B_xn03Z1tL1_0),.dout(w_dff_B_QJLoltAD1_0),.clk(gclk));
	jdff dff_B_Fb8SMVIa3_0(.din(w_dff_B_QJLoltAD1_0),.dout(w_dff_B_Fb8SMVIa3_0),.clk(gclk));
	jdff dff_B_P1VHCDv58_0(.din(w_dff_B_Fb8SMVIa3_0),.dout(w_dff_B_P1VHCDv58_0),.clk(gclk));
	jdff dff_B_PAFj1S6D1_0(.din(w_dff_B_P1VHCDv58_0),.dout(w_dff_B_PAFj1S6D1_0),.clk(gclk));
	jdff dff_B_N2x4cjw34_0(.din(w_dff_B_PAFj1S6D1_0),.dout(w_dff_B_N2x4cjw34_0),.clk(gclk));
	jdff dff_B_KnV2FWR59_0(.din(w_dff_B_N2x4cjw34_0),.dout(w_dff_B_KnV2FWR59_0),.clk(gclk));
	jdff dff_B_5kCbERLf3_0(.din(w_dff_B_KnV2FWR59_0),.dout(w_dff_B_5kCbERLf3_0),.clk(gclk));
	jdff dff_B_3JMxaSLI4_0(.din(w_dff_B_5kCbERLf3_0),.dout(w_dff_B_3JMxaSLI4_0),.clk(gclk));
	jdff dff_B_ojhdoTNr5_0(.din(w_dff_B_3JMxaSLI4_0),.dout(w_dff_B_ojhdoTNr5_0),.clk(gclk));
	jdff dff_B_79hYDlnI2_0(.din(w_dff_B_ojhdoTNr5_0),.dout(w_dff_B_79hYDlnI2_0),.clk(gclk));
	jdff dff_B_hv1CnjQo8_0(.din(w_dff_B_79hYDlnI2_0),.dout(w_dff_B_hv1CnjQo8_0),.clk(gclk));
	jdff dff_B_kxzh6M3k2_0(.din(w_dff_B_hv1CnjQo8_0),.dout(w_dff_B_kxzh6M3k2_0),.clk(gclk));
	jdff dff_B_Nr5B1aJJ8_0(.din(w_dff_B_kxzh6M3k2_0),.dout(w_dff_B_Nr5B1aJJ8_0),.clk(gclk));
	jdff dff_B_5YtuNvVb7_0(.din(w_dff_B_Nr5B1aJJ8_0),.dout(w_dff_B_5YtuNvVb7_0),.clk(gclk));
	jdff dff_B_fTk6qELK8_0(.din(w_dff_B_5YtuNvVb7_0),.dout(w_dff_B_fTk6qELK8_0),.clk(gclk));
	jdff dff_B_Y9GwHcLj4_0(.din(w_dff_B_fTk6qELK8_0),.dout(w_dff_B_Y9GwHcLj4_0),.clk(gclk));
	jdff dff_B_JHsTE69f6_0(.din(w_dff_B_Y9GwHcLj4_0),.dout(w_dff_B_JHsTE69f6_0),.clk(gclk));
	jdff dff_B_0yuJfA2i9_0(.din(w_dff_B_JHsTE69f6_0),.dout(w_dff_B_0yuJfA2i9_0),.clk(gclk));
	jdff dff_B_sVYMKFjH8_0(.din(w_dff_B_0yuJfA2i9_0),.dout(w_dff_B_sVYMKFjH8_0),.clk(gclk));
	jdff dff_B_boqzDCTa7_0(.din(w_dff_B_sVYMKFjH8_0),.dout(w_dff_B_boqzDCTa7_0),.clk(gclk));
	jdff dff_B_FlQP56M19_0(.din(w_dff_B_boqzDCTa7_0),.dout(w_dff_B_FlQP56M19_0),.clk(gclk));
	jdff dff_B_pIvosuE11_0(.din(w_dff_B_FlQP56M19_0),.dout(w_dff_B_pIvosuE11_0),.clk(gclk));
	jdff dff_B_V1P11FnG5_0(.din(w_dff_B_pIvosuE11_0),.dout(w_dff_B_V1P11FnG5_0),.clk(gclk));
	jdff dff_B_ZTPMJMoB1_0(.din(w_dff_B_V1P11FnG5_0),.dout(w_dff_B_ZTPMJMoB1_0),.clk(gclk));
	jdff dff_B_vsN6OyCu7_0(.din(w_dff_B_ZTPMJMoB1_0),.dout(w_dff_B_vsN6OyCu7_0),.clk(gclk));
	jdff dff_B_RIiq7q8v4_0(.din(w_dff_B_vsN6OyCu7_0),.dout(w_dff_B_RIiq7q8v4_0),.clk(gclk));
	jdff dff_B_xxQqVvOs7_0(.din(w_dff_B_RIiq7q8v4_0),.dout(w_dff_B_xxQqVvOs7_0),.clk(gclk));
	jdff dff_B_VGi2UROn2_0(.din(w_dff_B_xxQqVvOs7_0),.dout(w_dff_B_VGi2UROn2_0),.clk(gclk));
	jdff dff_B_LfbFJvMx6_0(.din(w_dff_B_VGi2UROn2_0),.dout(w_dff_B_LfbFJvMx6_0),.clk(gclk));
	jdff dff_B_lzEq9KiS3_0(.din(w_dff_B_LfbFJvMx6_0),.dout(w_dff_B_lzEq9KiS3_0),.clk(gclk));
	jdff dff_B_51K0myhB2_0(.din(w_dff_B_lzEq9KiS3_0),.dout(w_dff_B_51K0myhB2_0),.clk(gclk));
	jdff dff_B_yVjpxSIL5_0(.din(w_dff_B_51K0myhB2_0),.dout(w_dff_B_yVjpxSIL5_0),.clk(gclk));
	jdff dff_B_u0mSMN5R4_0(.din(w_dff_B_yVjpxSIL5_0),.dout(w_dff_B_u0mSMN5R4_0),.clk(gclk));
	jdff dff_B_7Yx8Zfv35_0(.din(w_dff_B_u0mSMN5R4_0),.dout(w_dff_B_7Yx8Zfv35_0),.clk(gclk));
	jdff dff_B_Edmle6YN9_0(.din(w_dff_B_7Yx8Zfv35_0),.dout(w_dff_B_Edmle6YN9_0),.clk(gclk));
	jdff dff_B_jh9DrEGX3_0(.din(w_dff_B_Edmle6YN9_0),.dout(w_dff_B_jh9DrEGX3_0),.clk(gclk));
	jdff dff_B_uGz6KgcW3_0(.din(w_dff_B_jh9DrEGX3_0),.dout(w_dff_B_uGz6KgcW3_0),.clk(gclk));
	jdff dff_B_y4oDZyQ10_0(.din(w_dff_B_uGz6KgcW3_0),.dout(w_dff_B_y4oDZyQ10_0),.clk(gclk));
	jdff dff_B_TDBOi6gD3_0(.din(w_dff_B_y4oDZyQ10_0),.dout(w_dff_B_TDBOi6gD3_0),.clk(gclk));
	jdff dff_B_XvVdIYiY5_0(.din(w_dff_B_TDBOi6gD3_0),.dout(w_dff_B_XvVdIYiY5_0),.clk(gclk));
	jdff dff_B_EPxaUYP49_0(.din(w_dff_B_XvVdIYiY5_0),.dout(w_dff_B_EPxaUYP49_0),.clk(gclk));
	jdff dff_B_irRoFLoY9_0(.din(w_dff_B_EPxaUYP49_0),.dout(w_dff_B_irRoFLoY9_0),.clk(gclk));
	jdff dff_B_EECg9nd90_0(.din(w_dff_B_irRoFLoY9_0),.dout(w_dff_B_EECg9nd90_0),.clk(gclk));
	jdff dff_B_VgEzxSYs5_0(.din(w_dff_B_EECg9nd90_0),.dout(w_dff_B_VgEzxSYs5_0),.clk(gclk));
	jdff dff_B_7tkvVyl15_0(.din(w_dff_B_VgEzxSYs5_0),.dout(w_dff_B_7tkvVyl15_0),.clk(gclk));
	jdff dff_B_aBm5XtYk9_0(.din(w_dff_B_7tkvVyl15_0),.dout(w_dff_B_aBm5XtYk9_0),.clk(gclk));
	jdff dff_B_Go4FIk7g5_0(.din(w_dff_B_aBm5XtYk9_0),.dout(w_dff_B_Go4FIk7g5_0),.clk(gclk));
	jdff dff_B_RLqf8HKD8_0(.din(w_dff_B_Go4FIk7g5_0),.dout(w_dff_B_RLqf8HKD8_0),.clk(gclk));
	jdff dff_B_fvnQjbWl0_0(.din(w_dff_B_RLqf8HKD8_0),.dout(w_dff_B_fvnQjbWl0_0),.clk(gclk));
	jdff dff_B_TowlVJ0s3_0(.din(w_dff_B_fvnQjbWl0_0),.dout(w_dff_B_TowlVJ0s3_0),.clk(gclk));
	jdff dff_B_DDEY6Udx4_0(.din(w_dff_B_TowlVJ0s3_0),.dout(w_dff_B_DDEY6Udx4_0),.clk(gclk));
	jdff dff_B_DY0PG0Dn3_0(.din(w_dff_B_DDEY6Udx4_0),.dout(w_dff_B_DY0PG0Dn3_0),.clk(gclk));
	jdff dff_B_zfqqG6SZ4_0(.din(w_dff_B_DY0PG0Dn3_0),.dout(w_dff_B_zfqqG6SZ4_0),.clk(gclk));
	jdff dff_B_MiIHbBHu4_0(.din(w_dff_B_zfqqG6SZ4_0),.dout(w_dff_B_MiIHbBHu4_0),.clk(gclk));
	jdff dff_B_8BzBcwhQ4_0(.din(w_dff_B_MiIHbBHu4_0),.dout(w_dff_B_8BzBcwhQ4_0),.clk(gclk));
	jdff dff_B_X8rmyqlc4_0(.din(w_dff_B_8BzBcwhQ4_0),.dout(w_dff_B_X8rmyqlc4_0),.clk(gclk));
	jdff dff_B_8P2FhsK52_0(.din(w_dff_B_X8rmyqlc4_0),.dout(w_dff_B_8P2FhsK52_0),.clk(gclk));
	jdff dff_B_ziWILxZA4_0(.din(w_dff_B_8P2FhsK52_0),.dout(w_dff_B_ziWILxZA4_0),.clk(gclk));
	jdff dff_B_jJoiKGuQ9_0(.din(w_dff_B_ziWILxZA4_0),.dout(w_dff_B_jJoiKGuQ9_0),.clk(gclk));
	jdff dff_B_sERyS6cS0_0(.din(w_dff_B_jJoiKGuQ9_0),.dout(w_dff_B_sERyS6cS0_0),.clk(gclk));
	jdff dff_B_7wHWZ19s7_0(.din(w_dff_B_sERyS6cS0_0),.dout(w_dff_B_7wHWZ19s7_0),.clk(gclk));
	jdff dff_B_E2pvJraB9_0(.din(w_dff_B_7wHWZ19s7_0),.dout(w_dff_B_E2pvJraB9_0),.clk(gclk));
	jdff dff_B_tHF5p0PX1_0(.din(w_dff_B_E2pvJraB9_0),.dout(w_dff_B_tHF5p0PX1_0),.clk(gclk));
	jdff dff_B_ikvCzPGE3_0(.din(w_dff_B_tHF5p0PX1_0),.dout(w_dff_B_ikvCzPGE3_0),.clk(gclk));
	jdff dff_B_uTbkv3wM3_0(.din(n808),.dout(w_dff_B_uTbkv3wM3_0),.clk(gclk));
	jdff dff_B_nCrOTjUj5_0(.din(w_dff_B_uTbkv3wM3_0),.dout(w_dff_B_nCrOTjUj5_0),.clk(gclk));
	jdff dff_B_dWG8H5mb1_0(.din(w_dff_B_nCrOTjUj5_0),.dout(w_dff_B_dWG8H5mb1_0),.clk(gclk));
	jdff dff_B_FRzK9OWb5_0(.din(w_dff_B_dWG8H5mb1_0),.dout(w_dff_B_FRzK9OWb5_0),.clk(gclk));
	jdff dff_B_rG2duiSU8_0(.din(w_dff_B_FRzK9OWb5_0),.dout(w_dff_B_rG2duiSU8_0),.clk(gclk));
	jdff dff_B_52EbAhTZ8_0(.din(w_dff_B_rG2duiSU8_0),.dout(w_dff_B_52EbAhTZ8_0),.clk(gclk));
	jdff dff_B_iZ8uguWo3_0(.din(w_dff_B_52EbAhTZ8_0),.dout(w_dff_B_iZ8uguWo3_0),.clk(gclk));
	jdff dff_B_gHq1mxHV0_0(.din(w_dff_B_iZ8uguWo3_0),.dout(w_dff_B_gHq1mxHV0_0),.clk(gclk));
	jdff dff_B_JXVqcLXq8_0(.din(w_dff_B_gHq1mxHV0_0),.dout(w_dff_B_JXVqcLXq8_0),.clk(gclk));
	jdff dff_B_FJxIsRPF3_0(.din(w_dff_B_JXVqcLXq8_0),.dout(w_dff_B_FJxIsRPF3_0),.clk(gclk));
	jdff dff_B_mtzEfBpI2_0(.din(w_dff_B_FJxIsRPF3_0),.dout(w_dff_B_mtzEfBpI2_0),.clk(gclk));
	jdff dff_B_Ek0fZKhM6_0(.din(w_dff_B_mtzEfBpI2_0),.dout(w_dff_B_Ek0fZKhM6_0),.clk(gclk));
	jdff dff_B_MFgqODb72_0(.din(w_dff_B_Ek0fZKhM6_0),.dout(w_dff_B_MFgqODb72_0),.clk(gclk));
	jdff dff_B_E9BiMMfI4_0(.din(w_dff_B_MFgqODb72_0),.dout(w_dff_B_E9BiMMfI4_0),.clk(gclk));
	jdff dff_B_Z2B8rynr4_0(.din(w_dff_B_E9BiMMfI4_0),.dout(w_dff_B_Z2B8rynr4_0),.clk(gclk));
	jdff dff_B_qmjaMPIw1_0(.din(w_dff_B_Z2B8rynr4_0),.dout(w_dff_B_qmjaMPIw1_0),.clk(gclk));
	jdff dff_B_ECrHf2zC6_0(.din(w_dff_B_qmjaMPIw1_0),.dout(w_dff_B_ECrHf2zC6_0),.clk(gclk));
	jdff dff_B_N9Kjlmw54_0(.din(w_dff_B_ECrHf2zC6_0),.dout(w_dff_B_N9Kjlmw54_0),.clk(gclk));
	jdff dff_B_n9mxIqXi0_0(.din(w_dff_B_N9Kjlmw54_0),.dout(w_dff_B_n9mxIqXi0_0),.clk(gclk));
	jdff dff_B_EyMGRDZg7_0(.din(w_dff_B_n9mxIqXi0_0),.dout(w_dff_B_EyMGRDZg7_0),.clk(gclk));
	jdff dff_B_xU0f3KRl2_0(.din(w_dff_B_EyMGRDZg7_0),.dout(w_dff_B_xU0f3KRl2_0),.clk(gclk));
	jdff dff_B_3wEfpDUe2_0(.din(w_dff_B_xU0f3KRl2_0),.dout(w_dff_B_3wEfpDUe2_0),.clk(gclk));
	jdff dff_B_j2hspalA7_0(.din(w_dff_B_3wEfpDUe2_0),.dout(w_dff_B_j2hspalA7_0),.clk(gclk));
	jdff dff_B_8MbY1Ins3_0(.din(w_dff_B_j2hspalA7_0),.dout(w_dff_B_8MbY1Ins3_0),.clk(gclk));
	jdff dff_B_C58MuJw33_0(.din(w_dff_B_8MbY1Ins3_0),.dout(w_dff_B_C58MuJw33_0),.clk(gclk));
	jdff dff_B_it9OyEN43_0(.din(w_dff_B_C58MuJw33_0),.dout(w_dff_B_it9OyEN43_0),.clk(gclk));
	jdff dff_B_z1yQvdZP1_0(.din(w_dff_B_it9OyEN43_0),.dout(w_dff_B_z1yQvdZP1_0),.clk(gclk));
	jdff dff_B_2fj4AdYc9_0(.din(w_dff_B_z1yQvdZP1_0),.dout(w_dff_B_2fj4AdYc9_0),.clk(gclk));
	jdff dff_B_mZYvTbuO2_0(.din(w_dff_B_2fj4AdYc9_0),.dout(w_dff_B_mZYvTbuO2_0),.clk(gclk));
	jdff dff_B_hyCaKxBJ1_0(.din(w_dff_B_mZYvTbuO2_0),.dout(w_dff_B_hyCaKxBJ1_0),.clk(gclk));
	jdff dff_B_yF0xLxvP5_0(.din(w_dff_B_hyCaKxBJ1_0),.dout(w_dff_B_yF0xLxvP5_0),.clk(gclk));
	jdff dff_B_oSekbLOH3_0(.din(w_dff_B_yF0xLxvP5_0),.dout(w_dff_B_oSekbLOH3_0),.clk(gclk));
	jdff dff_B_h5XniCCh9_0(.din(w_dff_B_oSekbLOH3_0),.dout(w_dff_B_h5XniCCh9_0),.clk(gclk));
	jdff dff_B_F36HbM4L5_0(.din(w_dff_B_h5XniCCh9_0),.dout(w_dff_B_F36HbM4L5_0),.clk(gclk));
	jdff dff_B_8jbe1RDh6_0(.din(w_dff_B_F36HbM4L5_0),.dout(w_dff_B_8jbe1RDh6_0),.clk(gclk));
	jdff dff_B_MBsrpKVZ5_0(.din(w_dff_B_8jbe1RDh6_0),.dout(w_dff_B_MBsrpKVZ5_0),.clk(gclk));
	jdff dff_B_No3w8VlE4_0(.din(w_dff_B_MBsrpKVZ5_0),.dout(w_dff_B_No3w8VlE4_0),.clk(gclk));
	jdff dff_B_iTvkgpvC3_0(.din(w_dff_B_No3w8VlE4_0),.dout(w_dff_B_iTvkgpvC3_0),.clk(gclk));
	jdff dff_B_Q6i39hrm5_0(.din(w_dff_B_iTvkgpvC3_0),.dout(w_dff_B_Q6i39hrm5_0),.clk(gclk));
	jdff dff_B_jCPROOyD2_0(.din(w_dff_B_Q6i39hrm5_0),.dout(w_dff_B_jCPROOyD2_0),.clk(gclk));
	jdff dff_B_Fb065wS42_0(.din(w_dff_B_jCPROOyD2_0),.dout(w_dff_B_Fb065wS42_0),.clk(gclk));
	jdff dff_B_yX0WWuD12_0(.din(w_dff_B_Fb065wS42_0),.dout(w_dff_B_yX0WWuD12_0),.clk(gclk));
	jdff dff_B_4OnC4kUA0_0(.din(w_dff_B_yX0WWuD12_0),.dout(w_dff_B_4OnC4kUA0_0),.clk(gclk));
	jdff dff_B_NmIgjnUJ4_0(.din(w_dff_B_4OnC4kUA0_0),.dout(w_dff_B_NmIgjnUJ4_0),.clk(gclk));
	jdff dff_B_9ffK5bGL2_0(.din(w_dff_B_NmIgjnUJ4_0),.dout(w_dff_B_9ffK5bGL2_0),.clk(gclk));
	jdff dff_B_k6IMr95z9_0(.din(w_dff_B_9ffK5bGL2_0),.dout(w_dff_B_k6IMr95z9_0),.clk(gclk));
	jdff dff_B_bJdwZxlZ6_0(.din(w_dff_B_k6IMr95z9_0),.dout(w_dff_B_bJdwZxlZ6_0),.clk(gclk));
	jdff dff_B_uIoZfzIv8_0(.din(w_dff_B_bJdwZxlZ6_0),.dout(w_dff_B_uIoZfzIv8_0),.clk(gclk));
	jdff dff_B_aH30KB3z9_0(.din(w_dff_B_uIoZfzIv8_0),.dout(w_dff_B_aH30KB3z9_0),.clk(gclk));
	jdff dff_B_lHzUY87g9_0(.din(w_dff_B_aH30KB3z9_0),.dout(w_dff_B_lHzUY87g9_0),.clk(gclk));
	jdff dff_B_KUCqu5vt6_0(.din(w_dff_B_lHzUY87g9_0),.dout(w_dff_B_KUCqu5vt6_0),.clk(gclk));
	jdff dff_B_vd20wg4n1_0(.din(w_dff_B_KUCqu5vt6_0),.dout(w_dff_B_vd20wg4n1_0),.clk(gclk));
	jdff dff_B_cNHPUzQw7_0(.din(w_dff_B_vd20wg4n1_0),.dout(w_dff_B_cNHPUzQw7_0),.clk(gclk));
	jdff dff_B_EvEo9Pkn7_0(.din(w_dff_B_cNHPUzQw7_0),.dout(w_dff_B_EvEo9Pkn7_0),.clk(gclk));
	jdff dff_B_HWib5OwB6_0(.din(w_dff_B_EvEo9Pkn7_0),.dout(w_dff_B_HWib5OwB6_0),.clk(gclk));
	jdff dff_B_lsQWPwDm6_0(.din(w_dff_B_HWib5OwB6_0),.dout(w_dff_B_lsQWPwDm6_0),.clk(gclk));
	jdff dff_B_Fyj2NwWY0_0(.din(w_dff_B_lsQWPwDm6_0),.dout(w_dff_B_Fyj2NwWY0_0),.clk(gclk));
	jdff dff_B_MaksMQu45_0(.din(w_dff_B_Fyj2NwWY0_0),.dout(w_dff_B_MaksMQu45_0),.clk(gclk));
	jdff dff_B_tiLy5M3X9_0(.din(w_dff_B_MaksMQu45_0),.dout(w_dff_B_tiLy5M3X9_0),.clk(gclk));
	jdff dff_B_rEqIzkkt0_0(.din(w_dff_B_tiLy5M3X9_0),.dout(w_dff_B_rEqIzkkt0_0),.clk(gclk));
	jdff dff_B_UbiNwkFQ5_0(.din(w_dff_B_rEqIzkkt0_0),.dout(w_dff_B_UbiNwkFQ5_0),.clk(gclk));
	jdff dff_B_fLIkzIlP5_0(.din(w_dff_B_UbiNwkFQ5_0),.dout(w_dff_B_fLIkzIlP5_0),.clk(gclk));
	jdff dff_B_GKbXsgKF8_0(.din(w_dff_B_fLIkzIlP5_0),.dout(w_dff_B_GKbXsgKF8_0),.clk(gclk));
	jdff dff_B_Way09Ywm0_0(.din(w_dff_B_GKbXsgKF8_0),.dout(w_dff_B_Way09Ywm0_0),.clk(gclk));
	jdff dff_B_KUii6ckP9_0(.din(w_dff_B_Way09Ywm0_0),.dout(w_dff_B_KUii6ckP9_0),.clk(gclk));
	jdff dff_B_646MqpjW3_0(.din(w_dff_B_KUii6ckP9_0),.dout(w_dff_B_646MqpjW3_0),.clk(gclk));
	jdff dff_B_w3lR9CXB0_0(.din(w_dff_B_646MqpjW3_0),.dout(w_dff_B_w3lR9CXB0_0),.clk(gclk));
	jdff dff_B_fm8cLBpR6_0(.din(w_dff_B_w3lR9CXB0_0),.dout(w_dff_B_fm8cLBpR6_0),.clk(gclk));
	jdff dff_B_ju8l2vfT0_0(.din(w_dff_B_fm8cLBpR6_0),.dout(w_dff_B_ju8l2vfT0_0),.clk(gclk));
	jdff dff_B_JxWKhrsd3_0(.din(w_dff_B_ju8l2vfT0_0),.dout(w_dff_B_JxWKhrsd3_0),.clk(gclk));
	jdff dff_B_K8KR1v0h0_0(.din(n814),.dout(w_dff_B_K8KR1v0h0_0),.clk(gclk));
	jdff dff_B_UvqYw03W5_0(.din(w_dff_B_K8KR1v0h0_0),.dout(w_dff_B_UvqYw03W5_0),.clk(gclk));
	jdff dff_B_h9uCuHdf8_0(.din(w_dff_B_UvqYw03W5_0),.dout(w_dff_B_h9uCuHdf8_0),.clk(gclk));
	jdff dff_B_joHR6gXx1_0(.din(w_dff_B_h9uCuHdf8_0),.dout(w_dff_B_joHR6gXx1_0),.clk(gclk));
	jdff dff_B_LJCweJus4_0(.din(w_dff_B_joHR6gXx1_0),.dout(w_dff_B_LJCweJus4_0),.clk(gclk));
	jdff dff_B_6kHkPDp78_0(.din(w_dff_B_LJCweJus4_0),.dout(w_dff_B_6kHkPDp78_0),.clk(gclk));
	jdff dff_B_yQxSAM1L6_0(.din(w_dff_B_6kHkPDp78_0),.dout(w_dff_B_yQxSAM1L6_0),.clk(gclk));
	jdff dff_B_PhCI8RNz2_0(.din(w_dff_B_yQxSAM1L6_0),.dout(w_dff_B_PhCI8RNz2_0),.clk(gclk));
	jdff dff_B_SwtgvfxI4_0(.din(w_dff_B_PhCI8RNz2_0),.dout(w_dff_B_SwtgvfxI4_0),.clk(gclk));
	jdff dff_B_Ek657jhd9_0(.din(w_dff_B_SwtgvfxI4_0),.dout(w_dff_B_Ek657jhd9_0),.clk(gclk));
	jdff dff_B_6vcnl2iQ6_0(.din(w_dff_B_Ek657jhd9_0),.dout(w_dff_B_6vcnl2iQ6_0),.clk(gclk));
	jdff dff_B_5SLe2eNO3_0(.din(w_dff_B_6vcnl2iQ6_0),.dout(w_dff_B_5SLe2eNO3_0),.clk(gclk));
	jdff dff_B_CFDwVCYX8_0(.din(w_dff_B_5SLe2eNO3_0),.dout(w_dff_B_CFDwVCYX8_0),.clk(gclk));
	jdff dff_B_8XovsaSy3_0(.din(w_dff_B_CFDwVCYX8_0),.dout(w_dff_B_8XovsaSy3_0),.clk(gclk));
	jdff dff_B_Lb1t9QhG6_0(.din(w_dff_B_8XovsaSy3_0),.dout(w_dff_B_Lb1t9QhG6_0),.clk(gclk));
	jdff dff_B_1bIKvqNO8_0(.din(w_dff_B_Lb1t9QhG6_0),.dout(w_dff_B_1bIKvqNO8_0),.clk(gclk));
	jdff dff_B_HXQTeHnK9_0(.din(w_dff_B_1bIKvqNO8_0),.dout(w_dff_B_HXQTeHnK9_0),.clk(gclk));
	jdff dff_B_9xeGihgn1_0(.din(w_dff_B_HXQTeHnK9_0),.dout(w_dff_B_9xeGihgn1_0),.clk(gclk));
	jdff dff_B_rqAiToFs3_0(.din(w_dff_B_9xeGihgn1_0),.dout(w_dff_B_rqAiToFs3_0),.clk(gclk));
	jdff dff_B_30v9Th3L5_0(.din(w_dff_B_rqAiToFs3_0),.dout(w_dff_B_30v9Th3L5_0),.clk(gclk));
	jdff dff_B_a1GkOzxU4_0(.din(w_dff_B_30v9Th3L5_0),.dout(w_dff_B_a1GkOzxU4_0),.clk(gclk));
	jdff dff_B_sqLqSx5U8_0(.din(w_dff_B_a1GkOzxU4_0),.dout(w_dff_B_sqLqSx5U8_0),.clk(gclk));
	jdff dff_B_6AmJ106J1_0(.din(w_dff_B_sqLqSx5U8_0),.dout(w_dff_B_6AmJ106J1_0),.clk(gclk));
	jdff dff_B_NwqyJ2OD2_0(.din(w_dff_B_6AmJ106J1_0),.dout(w_dff_B_NwqyJ2OD2_0),.clk(gclk));
	jdff dff_B_yEk5ecGq2_0(.din(w_dff_B_NwqyJ2OD2_0),.dout(w_dff_B_yEk5ecGq2_0),.clk(gclk));
	jdff dff_B_AoKGARec0_0(.din(w_dff_B_yEk5ecGq2_0),.dout(w_dff_B_AoKGARec0_0),.clk(gclk));
	jdff dff_B_mrT4pSGv1_0(.din(w_dff_B_AoKGARec0_0),.dout(w_dff_B_mrT4pSGv1_0),.clk(gclk));
	jdff dff_B_b1mSl9DT0_0(.din(w_dff_B_mrT4pSGv1_0),.dout(w_dff_B_b1mSl9DT0_0),.clk(gclk));
	jdff dff_B_goXRnpUM6_0(.din(w_dff_B_b1mSl9DT0_0),.dout(w_dff_B_goXRnpUM6_0),.clk(gclk));
	jdff dff_B_bVBNA7wK3_0(.din(w_dff_B_goXRnpUM6_0),.dout(w_dff_B_bVBNA7wK3_0),.clk(gclk));
	jdff dff_B_R4Xup1eB1_0(.din(w_dff_B_bVBNA7wK3_0),.dout(w_dff_B_R4Xup1eB1_0),.clk(gclk));
	jdff dff_B_XdzVqCzX3_0(.din(w_dff_B_R4Xup1eB1_0),.dout(w_dff_B_XdzVqCzX3_0),.clk(gclk));
	jdff dff_B_HBiiIxZ67_0(.din(w_dff_B_XdzVqCzX3_0),.dout(w_dff_B_HBiiIxZ67_0),.clk(gclk));
	jdff dff_B_Kum9dh4r7_0(.din(w_dff_B_HBiiIxZ67_0),.dout(w_dff_B_Kum9dh4r7_0),.clk(gclk));
	jdff dff_B_u55DL7ub0_0(.din(w_dff_B_Kum9dh4r7_0),.dout(w_dff_B_u55DL7ub0_0),.clk(gclk));
	jdff dff_B_GohZT36D3_0(.din(w_dff_B_u55DL7ub0_0),.dout(w_dff_B_GohZT36D3_0),.clk(gclk));
	jdff dff_B_HvEYUVtu8_0(.din(w_dff_B_GohZT36D3_0),.dout(w_dff_B_HvEYUVtu8_0),.clk(gclk));
	jdff dff_B_zDTbwalz8_0(.din(w_dff_B_HvEYUVtu8_0),.dout(w_dff_B_zDTbwalz8_0),.clk(gclk));
	jdff dff_B_DgA6ozJq1_0(.din(w_dff_B_zDTbwalz8_0),.dout(w_dff_B_DgA6ozJq1_0),.clk(gclk));
	jdff dff_B_7b6bYiHg5_0(.din(w_dff_B_DgA6ozJq1_0),.dout(w_dff_B_7b6bYiHg5_0),.clk(gclk));
	jdff dff_B_zkA0H2TJ0_0(.din(w_dff_B_7b6bYiHg5_0),.dout(w_dff_B_zkA0H2TJ0_0),.clk(gclk));
	jdff dff_B_7A5a7cYa4_0(.din(w_dff_B_zkA0H2TJ0_0),.dout(w_dff_B_7A5a7cYa4_0),.clk(gclk));
	jdff dff_B_B0dLc4Kb9_0(.din(w_dff_B_7A5a7cYa4_0),.dout(w_dff_B_B0dLc4Kb9_0),.clk(gclk));
	jdff dff_B_geok2ODD5_0(.din(w_dff_B_B0dLc4Kb9_0),.dout(w_dff_B_geok2ODD5_0),.clk(gclk));
	jdff dff_B_TnBIMtmU7_0(.din(w_dff_B_geok2ODD5_0),.dout(w_dff_B_TnBIMtmU7_0),.clk(gclk));
	jdff dff_B_JktU5inu7_0(.din(w_dff_B_TnBIMtmU7_0),.dout(w_dff_B_JktU5inu7_0),.clk(gclk));
	jdff dff_B_Jv2UVd6g1_0(.din(w_dff_B_JktU5inu7_0),.dout(w_dff_B_Jv2UVd6g1_0),.clk(gclk));
	jdff dff_B_VkFRakZ91_0(.din(w_dff_B_Jv2UVd6g1_0),.dout(w_dff_B_VkFRakZ91_0),.clk(gclk));
	jdff dff_B_xW0kb1In4_0(.din(w_dff_B_VkFRakZ91_0),.dout(w_dff_B_xW0kb1In4_0),.clk(gclk));
	jdff dff_B_TsWlvTGw2_0(.din(w_dff_B_xW0kb1In4_0),.dout(w_dff_B_TsWlvTGw2_0),.clk(gclk));
	jdff dff_B_ghueHGkG3_0(.din(w_dff_B_TsWlvTGw2_0),.dout(w_dff_B_ghueHGkG3_0),.clk(gclk));
	jdff dff_B_csVN0p779_0(.din(w_dff_B_ghueHGkG3_0),.dout(w_dff_B_csVN0p779_0),.clk(gclk));
	jdff dff_B_Fr2XhxCO7_0(.din(w_dff_B_csVN0p779_0),.dout(w_dff_B_Fr2XhxCO7_0),.clk(gclk));
	jdff dff_B_CY5I6Dgz8_0(.din(w_dff_B_Fr2XhxCO7_0),.dout(w_dff_B_CY5I6Dgz8_0),.clk(gclk));
	jdff dff_B_pmmZEC6D4_0(.din(w_dff_B_CY5I6Dgz8_0),.dout(w_dff_B_pmmZEC6D4_0),.clk(gclk));
	jdff dff_B_WXt3uY0G0_0(.din(w_dff_B_pmmZEC6D4_0),.dout(w_dff_B_WXt3uY0G0_0),.clk(gclk));
	jdff dff_B_A0YB9WqP1_0(.din(w_dff_B_WXt3uY0G0_0),.dout(w_dff_B_A0YB9WqP1_0),.clk(gclk));
	jdff dff_B_IlM6eD5D1_0(.din(w_dff_B_A0YB9WqP1_0),.dout(w_dff_B_IlM6eD5D1_0),.clk(gclk));
	jdff dff_B_lIwnggMu4_0(.din(w_dff_B_IlM6eD5D1_0),.dout(w_dff_B_lIwnggMu4_0),.clk(gclk));
	jdff dff_B_c7NH46Op4_0(.din(w_dff_B_lIwnggMu4_0),.dout(w_dff_B_c7NH46Op4_0),.clk(gclk));
	jdff dff_B_jrvJuDlt4_0(.din(w_dff_B_c7NH46Op4_0),.dout(w_dff_B_jrvJuDlt4_0),.clk(gclk));
	jdff dff_B_Ah0VBcm17_0(.din(w_dff_B_jrvJuDlt4_0),.dout(w_dff_B_Ah0VBcm17_0),.clk(gclk));
	jdff dff_B_5orD6xrr6_0(.din(w_dff_B_Ah0VBcm17_0),.dout(w_dff_B_5orD6xrr6_0),.clk(gclk));
	jdff dff_B_JMSRNqWX5_0(.din(w_dff_B_5orD6xrr6_0),.dout(w_dff_B_JMSRNqWX5_0),.clk(gclk));
	jdff dff_B_1foiTy730_0(.din(w_dff_B_JMSRNqWX5_0),.dout(w_dff_B_1foiTy730_0),.clk(gclk));
	jdff dff_B_VrOceuR77_0(.din(w_dff_B_1foiTy730_0),.dout(w_dff_B_VrOceuR77_0),.clk(gclk));
	jdff dff_B_lsMFHzPE9_0(.din(w_dff_B_VrOceuR77_0),.dout(w_dff_B_lsMFHzPE9_0),.clk(gclk));
	jdff dff_B_pUFufnay7_0(.din(w_dff_B_lsMFHzPE9_0),.dout(w_dff_B_pUFufnay7_0),.clk(gclk));
	jdff dff_B_EUX6sfvJ6_0(.din(w_dff_B_pUFufnay7_0),.dout(w_dff_B_EUX6sfvJ6_0),.clk(gclk));
	jdff dff_B_iG9NtK4K1_0(.din(w_dff_B_EUX6sfvJ6_0),.dout(w_dff_B_iG9NtK4K1_0),.clk(gclk));
	jdff dff_B_pv3sBp5K2_0(.din(w_dff_B_iG9NtK4K1_0),.dout(w_dff_B_pv3sBp5K2_0),.clk(gclk));
	jdff dff_B_gjtWZT8u6_0(.din(n820),.dout(w_dff_B_gjtWZT8u6_0),.clk(gclk));
	jdff dff_B_U3Z9hAzM4_0(.din(w_dff_B_gjtWZT8u6_0),.dout(w_dff_B_U3Z9hAzM4_0),.clk(gclk));
	jdff dff_B_BoShgiUc7_0(.din(w_dff_B_U3Z9hAzM4_0),.dout(w_dff_B_BoShgiUc7_0),.clk(gclk));
	jdff dff_B_c9yTcfM50_0(.din(w_dff_B_BoShgiUc7_0),.dout(w_dff_B_c9yTcfM50_0),.clk(gclk));
	jdff dff_B_hD1e3CLC0_0(.din(w_dff_B_c9yTcfM50_0),.dout(w_dff_B_hD1e3CLC0_0),.clk(gclk));
	jdff dff_B_XBFHlLzf8_0(.din(w_dff_B_hD1e3CLC0_0),.dout(w_dff_B_XBFHlLzf8_0),.clk(gclk));
	jdff dff_B_bR8CSXxS3_0(.din(w_dff_B_XBFHlLzf8_0),.dout(w_dff_B_bR8CSXxS3_0),.clk(gclk));
	jdff dff_B_RYBOLw7n3_0(.din(w_dff_B_bR8CSXxS3_0),.dout(w_dff_B_RYBOLw7n3_0),.clk(gclk));
	jdff dff_B_0T3Nbega6_0(.din(w_dff_B_RYBOLw7n3_0),.dout(w_dff_B_0T3Nbega6_0),.clk(gclk));
	jdff dff_B_VB5P8UTL5_0(.din(w_dff_B_0T3Nbega6_0),.dout(w_dff_B_VB5P8UTL5_0),.clk(gclk));
	jdff dff_B_GePgwC936_0(.din(w_dff_B_VB5P8UTL5_0),.dout(w_dff_B_GePgwC936_0),.clk(gclk));
	jdff dff_B_ukDCK8Vf6_0(.din(w_dff_B_GePgwC936_0),.dout(w_dff_B_ukDCK8Vf6_0),.clk(gclk));
	jdff dff_B_KAGeyIyS6_0(.din(w_dff_B_ukDCK8Vf6_0),.dout(w_dff_B_KAGeyIyS6_0),.clk(gclk));
	jdff dff_B_QMxEWjXT3_0(.din(w_dff_B_KAGeyIyS6_0),.dout(w_dff_B_QMxEWjXT3_0),.clk(gclk));
	jdff dff_B_1DKQEo9i2_0(.din(w_dff_B_QMxEWjXT3_0),.dout(w_dff_B_1DKQEo9i2_0),.clk(gclk));
	jdff dff_B_GIOxWv5h3_0(.din(w_dff_B_1DKQEo9i2_0),.dout(w_dff_B_GIOxWv5h3_0),.clk(gclk));
	jdff dff_B_FUPMUI5t3_0(.din(w_dff_B_GIOxWv5h3_0),.dout(w_dff_B_FUPMUI5t3_0),.clk(gclk));
	jdff dff_B_lpcqvB2h3_0(.din(w_dff_B_FUPMUI5t3_0),.dout(w_dff_B_lpcqvB2h3_0),.clk(gclk));
	jdff dff_B_UUCqwFXR2_0(.din(w_dff_B_lpcqvB2h3_0),.dout(w_dff_B_UUCqwFXR2_0),.clk(gclk));
	jdff dff_B_PkJzX0Ml5_0(.din(w_dff_B_UUCqwFXR2_0),.dout(w_dff_B_PkJzX0Ml5_0),.clk(gclk));
	jdff dff_B_CWeJCeTY4_0(.din(w_dff_B_PkJzX0Ml5_0),.dout(w_dff_B_CWeJCeTY4_0),.clk(gclk));
	jdff dff_B_2A7qYmVr9_0(.din(w_dff_B_CWeJCeTY4_0),.dout(w_dff_B_2A7qYmVr9_0),.clk(gclk));
	jdff dff_B_Yx54bmGe0_0(.din(w_dff_B_2A7qYmVr9_0),.dout(w_dff_B_Yx54bmGe0_0),.clk(gclk));
	jdff dff_B_99vr0vfs6_0(.din(w_dff_B_Yx54bmGe0_0),.dout(w_dff_B_99vr0vfs6_0),.clk(gclk));
	jdff dff_B_LWpVHPFi6_0(.din(w_dff_B_99vr0vfs6_0),.dout(w_dff_B_LWpVHPFi6_0),.clk(gclk));
	jdff dff_B_LtqzSqf73_0(.din(w_dff_B_LWpVHPFi6_0),.dout(w_dff_B_LtqzSqf73_0),.clk(gclk));
	jdff dff_B_nd50uFT93_0(.din(w_dff_B_LtqzSqf73_0),.dout(w_dff_B_nd50uFT93_0),.clk(gclk));
	jdff dff_B_Sq60IGAl3_0(.din(w_dff_B_nd50uFT93_0),.dout(w_dff_B_Sq60IGAl3_0),.clk(gclk));
	jdff dff_B_WHj74Hgr6_0(.din(w_dff_B_Sq60IGAl3_0),.dout(w_dff_B_WHj74Hgr6_0),.clk(gclk));
	jdff dff_B_NKp9N87a6_0(.din(w_dff_B_WHj74Hgr6_0),.dout(w_dff_B_NKp9N87a6_0),.clk(gclk));
	jdff dff_B_KqURzsvA4_0(.din(w_dff_B_NKp9N87a6_0),.dout(w_dff_B_KqURzsvA4_0),.clk(gclk));
	jdff dff_B_XHCHRC666_0(.din(w_dff_B_KqURzsvA4_0),.dout(w_dff_B_XHCHRC666_0),.clk(gclk));
	jdff dff_B_luqQTiZz7_0(.din(w_dff_B_XHCHRC666_0),.dout(w_dff_B_luqQTiZz7_0),.clk(gclk));
	jdff dff_B_aQrUFAWZ0_0(.din(w_dff_B_luqQTiZz7_0),.dout(w_dff_B_aQrUFAWZ0_0),.clk(gclk));
	jdff dff_B_vguzv9tU7_0(.din(w_dff_B_aQrUFAWZ0_0),.dout(w_dff_B_vguzv9tU7_0),.clk(gclk));
	jdff dff_B_USkauRet9_0(.din(w_dff_B_vguzv9tU7_0),.dout(w_dff_B_USkauRet9_0),.clk(gclk));
	jdff dff_B_Ugfr3I697_0(.din(w_dff_B_USkauRet9_0),.dout(w_dff_B_Ugfr3I697_0),.clk(gclk));
	jdff dff_B_8LO3tYGd8_0(.din(w_dff_B_Ugfr3I697_0),.dout(w_dff_B_8LO3tYGd8_0),.clk(gclk));
	jdff dff_B_1Z9ckb7l5_0(.din(w_dff_B_8LO3tYGd8_0),.dout(w_dff_B_1Z9ckb7l5_0),.clk(gclk));
	jdff dff_B_bc79WY4J3_0(.din(w_dff_B_1Z9ckb7l5_0),.dout(w_dff_B_bc79WY4J3_0),.clk(gclk));
	jdff dff_B_1Yuc01Af7_0(.din(w_dff_B_bc79WY4J3_0),.dout(w_dff_B_1Yuc01Af7_0),.clk(gclk));
	jdff dff_B_zsrHNdGQ9_0(.din(w_dff_B_1Yuc01Af7_0),.dout(w_dff_B_zsrHNdGQ9_0),.clk(gclk));
	jdff dff_B_63BceWwP8_0(.din(w_dff_B_zsrHNdGQ9_0),.dout(w_dff_B_63BceWwP8_0),.clk(gclk));
	jdff dff_B_DyEX1x7T5_0(.din(w_dff_B_63BceWwP8_0),.dout(w_dff_B_DyEX1x7T5_0),.clk(gclk));
	jdff dff_B_oIFEkwfl4_0(.din(w_dff_B_DyEX1x7T5_0),.dout(w_dff_B_oIFEkwfl4_0),.clk(gclk));
	jdff dff_B_hK28HObY6_0(.din(w_dff_B_oIFEkwfl4_0),.dout(w_dff_B_hK28HObY6_0),.clk(gclk));
	jdff dff_B_73y1Gfaz3_0(.din(w_dff_B_hK28HObY6_0),.dout(w_dff_B_73y1Gfaz3_0),.clk(gclk));
	jdff dff_B_hqH6fwBA0_0(.din(w_dff_B_73y1Gfaz3_0),.dout(w_dff_B_hqH6fwBA0_0),.clk(gclk));
	jdff dff_B_CvrIixkZ0_0(.din(w_dff_B_hqH6fwBA0_0),.dout(w_dff_B_CvrIixkZ0_0),.clk(gclk));
	jdff dff_B_UWyGvAfr4_0(.din(w_dff_B_CvrIixkZ0_0),.dout(w_dff_B_UWyGvAfr4_0),.clk(gclk));
	jdff dff_B_becLxMS63_0(.din(w_dff_B_UWyGvAfr4_0),.dout(w_dff_B_becLxMS63_0),.clk(gclk));
	jdff dff_B_vlsL3pMh2_0(.din(w_dff_B_becLxMS63_0),.dout(w_dff_B_vlsL3pMh2_0),.clk(gclk));
	jdff dff_B_KApHAKxm1_0(.din(w_dff_B_vlsL3pMh2_0),.dout(w_dff_B_KApHAKxm1_0),.clk(gclk));
	jdff dff_B_mmkX4I9b6_0(.din(w_dff_B_KApHAKxm1_0),.dout(w_dff_B_mmkX4I9b6_0),.clk(gclk));
	jdff dff_B_EcdDGgM70_0(.din(w_dff_B_mmkX4I9b6_0),.dout(w_dff_B_EcdDGgM70_0),.clk(gclk));
	jdff dff_B_y1qEE1vH6_0(.din(w_dff_B_EcdDGgM70_0),.dout(w_dff_B_y1qEE1vH6_0),.clk(gclk));
	jdff dff_B_huZcUXJl1_0(.din(w_dff_B_y1qEE1vH6_0),.dout(w_dff_B_huZcUXJl1_0),.clk(gclk));
	jdff dff_B_7ys95aUX5_0(.din(w_dff_B_huZcUXJl1_0),.dout(w_dff_B_7ys95aUX5_0),.clk(gclk));
	jdff dff_B_WOH18U781_0(.din(w_dff_B_7ys95aUX5_0),.dout(w_dff_B_WOH18U781_0),.clk(gclk));
	jdff dff_B_DwoezAJJ7_0(.din(w_dff_B_WOH18U781_0),.dout(w_dff_B_DwoezAJJ7_0),.clk(gclk));
	jdff dff_B_gDS4yW2p0_0(.din(w_dff_B_DwoezAJJ7_0),.dout(w_dff_B_gDS4yW2p0_0),.clk(gclk));
	jdff dff_B_I0xZM2qy9_0(.din(w_dff_B_gDS4yW2p0_0),.dout(w_dff_B_I0xZM2qy9_0),.clk(gclk));
	jdff dff_B_LaiBGMm09_0(.din(w_dff_B_I0xZM2qy9_0),.dout(w_dff_B_LaiBGMm09_0),.clk(gclk));
	jdff dff_B_p7xA06Kb4_0(.din(w_dff_B_LaiBGMm09_0),.dout(w_dff_B_p7xA06Kb4_0),.clk(gclk));
	jdff dff_B_hwR3UXWw2_0(.din(w_dff_B_p7xA06Kb4_0),.dout(w_dff_B_hwR3UXWw2_0),.clk(gclk));
	jdff dff_B_tPJbIVE25_0(.din(w_dff_B_hwR3UXWw2_0),.dout(w_dff_B_tPJbIVE25_0),.clk(gclk));
	jdff dff_B_98rxaBb90_0(.din(w_dff_B_tPJbIVE25_0),.dout(w_dff_B_98rxaBb90_0),.clk(gclk));
	jdff dff_B_15IQasa12_0(.din(w_dff_B_98rxaBb90_0),.dout(w_dff_B_15IQasa12_0),.clk(gclk));
	jdff dff_B_FdJzxjK20_0(.din(w_dff_B_15IQasa12_0),.dout(w_dff_B_FdJzxjK20_0),.clk(gclk));
	jdff dff_B_d3OJeoQD5_0(.din(w_dff_B_FdJzxjK20_0),.dout(w_dff_B_d3OJeoQD5_0),.clk(gclk));
	jdff dff_B_mOyQaOUP6_0(.din(w_dff_B_d3OJeoQD5_0),.dout(w_dff_B_mOyQaOUP6_0),.clk(gclk));
	jdff dff_B_FMC2ALGB0_0(.din(w_dff_B_mOyQaOUP6_0),.dout(w_dff_B_FMC2ALGB0_0),.clk(gclk));
	jdff dff_B_J5hZN5sU2_0(.din(n826),.dout(w_dff_B_J5hZN5sU2_0),.clk(gclk));
	jdff dff_B_swrFznVd2_0(.din(w_dff_B_J5hZN5sU2_0),.dout(w_dff_B_swrFznVd2_0),.clk(gclk));
	jdff dff_B_V7Aqu1az5_0(.din(w_dff_B_swrFznVd2_0),.dout(w_dff_B_V7Aqu1az5_0),.clk(gclk));
	jdff dff_B_yyhY2Yw85_0(.din(w_dff_B_V7Aqu1az5_0),.dout(w_dff_B_yyhY2Yw85_0),.clk(gclk));
	jdff dff_B_Su83XJaR1_0(.din(w_dff_B_yyhY2Yw85_0),.dout(w_dff_B_Su83XJaR1_0),.clk(gclk));
	jdff dff_B_CFUw9yfu4_0(.din(w_dff_B_Su83XJaR1_0),.dout(w_dff_B_CFUw9yfu4_0),.clk(gclk));
	jdff dff_B_4pKocEiJ6_0(.din(w_dff_B_CFUw9yfu4_0),.dout(w_dff_B_4pKocEiJ6_0),.clk(gclk));
	jdff dff_B_FhqjgeKJ9_0(.din(w_dff_B_4pKocEiJ6_0),.dout(w_dff_B_FhqjgeKJ9_0),.clk(gclk));
	jdff dff_B_Cz8B2XOQ2_0(.din(w_dff_B_FhqjgeKJ9_0),.dout(w_dff_B_Cz8B2XOQ2_0),.clk(gclk));
	jdff dff_B_yZtfL8ho2_0(.din(w_dff_B_Cz8B2XOQ2_0),.dout(w_dff_B_yZtfL8ho2_0),.clk(gclk));
	jdff dff_B_AMRUMcIZ0_0(.din(w_dff_B_yZtfL8ho2_0),.dout(w_dff_B_AMRUMcIZ0_0),.clk(gclk));
	jdff dff_B_0O8dBAK65_0(.din(w_dff_B_AMRUMcIZ0_0),.dout(w_dff_B_0O8dBAK65_0),.clk(gclk));
	jdff dff_B_eeSDeSIQ4_0(.din(w_dff_B_0O8dBAK65_0),.dout(w_dff_B_eeSDeSIQ4_0),.clk(gclk));
	jdff dff_B_AieIUgmS7_0(.din(w_dff_B_eeSDeSIQ4_0),.dout(w_dff_B_AieIUgmS7_0),.clk(gclk));
	jdff dff_B_L0WXBmqO4_0(.din(w_dff_B_AieIUgmS7_0),.dout(w_dff_B_L0WXBmqO4_0),.clk(gclk));
	jdff dff_B_rKpeCilG4_0(.din(w_dff_B_L0WXBmqO4_0),.dout(w_dff_B_rKpeCilG4_0),.clk(gclk));
	jdff dff_B_aoDqEjFW7_0(.din(w_dff_B_rKpeCilG4_0),.dout(w_dff_B_aoDqEjFW7_0),.clk(gclk));
	jdff dff_B_BOz2XnWz8_0(.din(w_dff_B_aoDqEjFW7_0),.dout(w_dff_B_BOz2XnWz8_0),.clk(gclk));
	jdff dff_B_uLflUQtv0_0(.din(w_dff_B_BOz2XnWz8_0),.dout(w_dff_B_uLflUQtv0_0),.clk(gclk));
	jdff dff_B_qpYuQQtv1_0(.din(w_dff_B_uLflUQtv0_0),.dout(w_dff_B_qpYuQQtv1_0),.clk(gclk));
	jdff dff_B_sgXW8qAx8_0(.din(w_dff_B_qpYuQQtv1_0),.dout(w_dff_B_sgXW8qAx8_0),.clk(gclk));
	jdff dff_B_eSjjEMdr2_0(.din(w_dff_B_sgXW8qAx8_0),.dout(w_dff_B_eSjjEMdr2_0),.clk(gclk));
	jdff dff_B_OHrR9IVm0_0(.din(w_dff_B_eSjjEMdr2_0),.dout(w_dff_B_OHrR9IVm0_0),.clk(gclk));
	jdff dff_B_OfMJidXT3_0(.din(w_dff_B_OHrR9IVm0_0),.dout(w_dff_B_OfMJidXT3_0),.clk(gclk));
	jdff dff_B_MOLD35Y74_0(.din(w_dff_B_OfMJidXT3_0),.dout(w_dff_B_MOLD35Y74_0),.clk(gclk));
	jdff dff_B_A7lgqtib8_0(.din(w_dff_B_MOLD35Y74_0),.dout(w_dff_B_A7lgqtib8_0),.clk(gclk));
	jdff dff_B_IgoGkVoq8_0(.din(w_dff_B_A7lgqtib8_0),.dout(w_dff_B_IgoGkVoq8_0),.clk(gclk));
	jdff dff_B_5i4re2bm3_0(.din(w_dff_B_IgoGkVoq8_0),.dout(w_dff_B_5i4re2bm3_0),.clk(gclk));
	jdff dff_B_VPrzomyO6_0(.din(w_dff_B_5i4re2bm3_0),.dout(w_dff_B_VPrzomyO6_0),.clk(gclk));
	jdff dff_B_p17P0aA03_0(.din(w_dff_B_VPrzomyO6_0),.dout(w_dff_B_p17P0aA03_0),.clk(gclk));
	jdff dff_B_xsvbUtpc6_0(.din(w_dff_B_p17P0aA03_0),.dout(w_dff_B_xsvbUtpc6_0),.clk(gclk));
	jdff dff_B_em69dLqe0_0(.din(w_dff_B_xsvbUtpc6_0),.dout(w_dff_B_em69dLqe0_0),.clk(gclk));
	jdff dff_B_Gl0rW1Qn8_0(.din(w_dff_B_em69dLqe0_0),.dout(w_dff_B_Gl0rW1Qn8_0),.clk(gclk));
	jdff dff_B_PhuHTBhY4_0(.din(w_dff_B_Gl0rW1Qn8_0),.dout(w_dff_B_PhuHTBhY4_0),.clk(gclk));
	jdff dff_B_rP8ne3da3_0(.din(w_dff_B_PhuHTBhY4_0),.dout(w_dff_B_rP8ne3da3_0),.clk(gclk));
	jdff dff_B_ERrrdDkU6_0(.din(w_dff_B_rP8ne3da3_0),.dout(w_dff_B_ERrrdDkU6_0),.clk(gclk));
	jdff dff_B_qZ2VEzT82_0(.din(w_dff_B_ERrrdDkU6_0),.dout(w_dff_B_qZ2VEzT82_0),.clk(gclk));
	jdff dff_B_4HMDwuKd5_0(.din(w_dff_B_qZ2VEzT82_0),.dout(w_dff_B_4HMDwuKd5_0),.clk(gclk));
	jdff dff_B_S1Kc1tjD1_0(.din(w_dff_B_4HMDwuKd5_0),.dout(w_dff_B_S1Kc1tjD1_0),.clk(gclk));
	jdff dff_B_P6SFdFZB3_0(.din(w_dff_B_S1Kc1tjD1_0),.dout(w_dff_B_P6SFdFZB3_0),.clk(gclk));
	jdff dff_B_OMmmPeWO5_0(.din(w_dff_B_P6SFdFZB3_0),.dout(w_dff_B_OMmmPeWO5_0),.clk(gclk));
	jdff dff_B_bfp2AXte5_0(.din(w_dff_B_OMmmPeWO5_0),.dout(w_dff_B_bfp2AXte5_0),.clk(gclk));
	jdff dff_B_ux7t2bqd3_0(.din(w_dff_B_bfp2AXte5_0),.dout(w_dff_B_ux7t2bqd3_0),.clk(gclk));
	jdff dff_B_oJTqfavZ4_0(.din(w_dff_B_ux7t2bqd3_0),.dout(w_dff_B_oJTqfavZ4_0),.clk(gclk));
	jdff dff_B_sDKk6S8e7_0(.din(w_dff_B_oJTqfavZ4_0),.dout(w_dff_B_sDKk6S8e7_0),.clk(gclk));
	jdff dff_B_OfW4Jghg9_0(.din(w_dff_B_sDKk6S8e7_0),.dout(w_dff_B_OfW4Jghg9_0),.clk(gclk));
	jdff dff_B_2pB8xujb7_0(.din(w_dff_B_OfW4Jghg9_0),.dout(w_dff_B_2pB8xujb7_0),.clk(gclk));
	jdff dff_B_pz7zkUlu3_0(.din(w_dff_B_2pB8xujb7_0),.dout(w_dff_B_pz7zkUlu3_0),.clk(gclk));
	jdff dff_B_SROJpiDS2_0(.din(w_dff_B_pz7zkUlu3_0),.dout(w_dff_B_SROJpiDS2_0),.clk(gclk));
	jdff dff_B_THjixmin7_0(.din(w_dff_B_SROJpiDS2_0),.dout(w_dff_B_THjixmin7_0),.clk(gclk));
	jdff dff_B_4af4m4Ov4_0(.din(w_dff_B_THjixmin7_0),.dout(w_dff_B_4af4m4Ov4_0),.clk(gclk));
	jdff dff_B_6S96Z7S51_0(.din(w_dff_B_4af4m4Ov4_0),.dout(w_dff_B_6S96Z7S51_0),.clk(gclk));
	jdff dff_B_i6YeeLqi1_0(.din(w_dff_B_6S96Z7S51_0),.dout(w_dff_B_i6YeeLqi1_0),.clk(gclk));
	jdff dff_B_4PV1JVpJ3_0(.din(w_dff_B_i6YeeLqi1_0),.dout(w_dff_B_4PV1JVpJ3_0),.clk(gclk));
	jdff dff_B_UGsB0gXX0_0(.din(w_dff_B_4PV1JVpJ3_0),.dout(w_dff_B_UGsB0gXX0_0),.clk(gclk));
	jdff dff_B_g3aasNoc1_0(.din(w_dff_B_UGsB0gXX0_0),.dout(w_dff_B_g3aasNoc1_0),.clk(gclk));
	jdff dff_B_4FAoKlbW9_0(.din(w_dff_B_g3aasNoc1_0),.dout(w_dff_B_4FAoKlbW9_0),.clk(gclk));
	jdff dff_B_zkkXAhQn5_0(.din(w_dff_B_4FAoKlbW9_0),.dout(w_dff_B_zkkXAhQn5_0),.clk(gclk));
	jdff dff_B_OLxbQuH34_0(.din(w_dff_B_zkkXAhQn5_0),.dout(w_dff_B_OLxbQuH34_0),.clk(gclk));
	jdff dff_B_KznebfxW6_0(.din(w_dff_B_OLxbQuH34_0),.dout(w_dff_B_KznebfxW6_0),.clk(gclk));
	jdff dff_B_aRBAKbmy4_0(.din(w_dff_B_KznebfxW6_0),.dout(w_dff_B_aRBAKbmy4_0),.clk(gclk));
	jdff dff_B_bNmyuJte7_0(.din(w_dff_B_aRBAKbmy4_0),.dout(w_dff_B_bNmyuJte7_0),.clk(gclk));
	jdff dff_B_wzlBs0G79_0(.din(w_dff_B_bNmyuJte7_0),.dout(w_dff_B_wzlBs0G79_0),.clk(gclk));
	jdff dff_B_7X1cEWH71_0(.din(w_dff_B_wzlBs0G79_0),.dout(w_dff_B_7X1cEWH71_0),.clk(gclk));
	jdff dff_B_Gi5pgYEa2_0(.din(w_dff_B_7X1cEWH71_0),.dout(w_dff_B_Gi5pgYEa2_0),.clk(gclk));
	jdff dff_B_uaSauKIB2_0(.din(w_dff_B_Gi5pgYEa2_0),.dout(w_dff_B_uaSauKIB2_0),.clk(gclk));
	jdff dff_B_EB2vTghp0_0(.din(w_dff_B_uaSauKIB2_0),.dout(w_dff_B_EB2vTghp0_0),.clk(gclk));
	jdff dff_B_3V14pkZT0_0(.din(w_dff_B_EB2vTghp0_0),.dout(w_dff_B_3V14pkZT0_0),.clk(gclk));
	jdff dff_B_SloTGfGm5_0(.din(w_dff_B_3V14pkZT0_0),.dout(w_dff_B_SloTGfGm5_0),.clk(gclk));
	jdff dff_B_YVnrL50z0_0(.din(w_dff_B_SloTGfGm5_0),.dout(w_dff_B_YVnrL50z0_0),.clk(gclk));
	jdff dff_B_2IlKruwx9_0(.din(w_dff_B_YVnrL50z0_0),.dout(w_dff_B_2IlKruwx9_0),.clk(gclk));
	jdff dff_B_kVoKSRtF3_0(.din(w_dff_B_2IlKruwx9_0),.dout(w_dff_B_kVoKSRtF3_0),.clk(gclk));
	jdff dff_B_Zb3Aui4E2_0(.din(w_dff_B_kVoKSRtF3_0),.dout(w_dff_B_Zb3Aui4E2_0),.clk(gclk));
	jdff dff_B_XIBVtP5T9_0(.din(n832),.dout(w_dff_B_XIBVtP5T9_0),.clk(gclk));
	jdff dff_B_hEIbsiQx7_0(.din(w_dff_B_XIBVtP5T9_0),.dout(w_dff_B_hEIbsiQx7_0),.clk(gclk));
	jdff dff_B_vVped8t61_0(.din(w_dff_B_hEIbsiQx7_0),.dout(w_dff_B_vVped8t61_0),.clk(gclk));
	jdff dff_B_ZkDUw77u5_0(.din(w_dff_B_vVped8t61_0),.dout(w_dff_B_ZkDUw77u5_0),.clk(gclk));
	jdff dff_B_MvzMNG2t9_0(.din(w_dff_B_ZkDUw77u5_0),.dout(w_dff_B_MvzMNG2t9_0),.clk(gclk));
	jdff dff_B_Ail5uBBE2_0(.din(w_dff_B_MvzMNG2t9_0),.dout(w_dff_B_Ail5uBBE2_0),.clk(gclk));
	jdff dff_B_qV1IbSDy5_0(.din(w_dff_B_Ail5uBBE2_0),.dout(w_dff_B_qV1IbSDy5_0),.clk(gclk));
	jdff dff_B_Or6PBY1k3_0(.din(w_dff_B_qV1IbSDy5_0),.dout(w_dff_B_Or6PBY1k3_0),.clk(gclk));
	jdff dff_B_gLQI5EyF4_0(.din(w_dff_B_Or6PBY1k3_0),.dout(w_dff_B_gLQI5EyF4_0),.clk(gclk));
	jdff dff_B_VUI7xP7N1_0(.din(w_dff_B_gLQI5EyF4_0),.dout(w_dff_B_VUI7xP7N1_0),.clk(gclk));
	jdff dff_B_ZrWmxTbZ5_0(.din(w_dff_B_VUI7xP7N1_0),.dout(w_dff_B_ZrWmxTbZ5_0),.clk(gclk));
	jdff dff_B_rKXDGhNW6_0(.din(w_dff_B_ZrWmxTbZ5_0),.dout(w_dff_B_rKXDGhNW6_0),.clk(gclk));
	jdff dff_B_CVSJZ2iq8_0(.din(w_dff_B_rKXDGhNW6_0),.dout(w_dff_B_CVSJZ2iq8_0),.clk(gclk));
	jdff dff_B_rC8u444R3_0(.din(w_dff_B_CVSJZ2iq8_0),.dout(w_dff_B_rC8u444R3_0),.clk(gclk));
	jdff dff_B_cL6aYRW21_0(.din(w_dff_B_rC8u444R3_0),.dout(w_dff_B_cL6aYRW21_0),.clk(gclk));
	jdff dff_B_OGDHVhHV9_0(.din(w_dff_B_cL6aYRW21_0),.dout(w_dff_B_OGDHVhHV9_0),.clk(gclk));
	jdff dff_B_btyvR2yp6_0(.din(w_dff_B_OGDHVhHV9_0),.dout(w_dff_B_btyvR2yp6_0),.clk(gclk));
	jdff dff_B_X3Y9Qcy22_0(.din(w_dff_B_btyvR2yp6_0),.dout(w_dff_B_X3Y9Qcy22_0),.clk(gclk));
	jdff dff_B_JZJLzT7R1_0(.din(w_dff_B_X3Y9Qcy22_0),.dout(w_dff_B_JZJLzT7R1_0),.clk(gclk));
	jdff dff_B_AJ7dbya17_0(.din(w_dff_B_JZJLzT7R1_0),.dout(w_dff_B_AJ7dbya17_0),.clk(gclk));
	jdff dff_B_v3UYbTMW8_0(.din(w_dff_B_AJ7dbya17_0),.dout(w_dff_B_v3UYbTMW8_0),.clk(gclk));
	jdff dff_B_DCkNC7O52_0(.din(w_dff_B_v3UYbTMW8_0),.dout(w_dff_B_DCkNC7O52_0),.clk(gclk));
	jdff dff_B_ki1KXNyQ2_0(.din(w_dff_B_DCkNC7O52_0),.dout(w_dff_B_ki1KXNyQ2_0),.clk(gclk));
	jdff dff_B_G0kFSLcc6_0(.din(w_dff_B_ki1KXNyQ2_0),.dout(w_dff_B_G0kFSLcc6_0),.clk(gclk));
	jdff dff_B_f8cyZzge4_0(.din(w_dff_B_G0kFSLcc6_0),.dout(w_dff_B_f8cyZzge4_0),.clk(gclk));
	jdff dff_B_EzaRmUX02_0(.din(w_dff_B_f8cyZzge4_0),.dout(w_dff_B_EzaRmUX02_0),.clk(gclk));
	jdff dff_B_0f8mKj3l1_0(.din(w_dff_B_EzaRmUX02_0),.dout(w_dff_B_0f8mKj3l1_0),.clk(gclk));
	jdff dff_B_kwHn0N3C3_0(.din(w_dff_B_0f8mKj3l1_0),.dout(w_dff_B_kwHn0N3C3_0),.clk(gclk));
	jdff dff_B_GH3kbN1A4_0(.din(w_dff_B_kwHn0N3C3_0),.dout(w_dff_B_GH3kbN1A4_0),.clk(gclk));
	jdff dff_B_Up5Zwngc3_0(.din(w_dff_B_GH3kbN1A4_0),.dout(w_dff_B_Up5Zwngc3_0),.clk(gclk));
	jdff dff_B_3M6pJRuC8_0(.din(w_dff_B_Up5Zwngc3_0),.dout(w_dff_B_3M6pJRuC8_0),.clk(gclk));
	jdff dff_B_1HnMSGBx7_0(.din(w_dff_B_3M6pJRuC8_0),.dout(w_dff_B_1HnMSGBx7_0),.clk(gclk));
	jdff dff_B_iTnGCJcI5_0(.din(w_dff_B_1HnMSGBx7_0),.dout(w_dff_B_iTnGCJcI5_0),.clk(gclk));
	jdff dff_B_J8qORiw16_0(.din(w_dff_B_iTnGCJcI5_0),.dout(w_dff_B_J8qORiw16_0),.clk(gclk));
	jdff dff_B_act0EzCl1_0(.din(w_dff_B_J8qORiw16_0),.dout(w_dff_B_act0EzCl1_0),.clk(gclk));
	jdff dff_B_MPgarCf60_0(.din(w_dff_B_act0EzCl1_0),.dout(w_dff_B_MPgarCf60_0),.clk(gclk));
	jdff dff_B_Zr5e05Kd9_0(.din(w_dff_B_MPgarCf60_0),.dout(w_dff_B_Zr5e05Kd9_0),.clk(gclk));
	jdff dff_B_w7QyZyJX4_0(.din(w_dff_B_Zr5e05Kd9_0),.dout(w_dff_B_w7QyZyJX4_0),.clk(gclk));
	jdff dff_B_VQl2595z1_0(.din(w_dff_B_w7QyZyJX4_0),.dout(w_dff_B_VQl2595z1_0),.clk(gclk));
	jdff dff_B_zGWPKchG6_0(.din(w_dff_B_VQl2595z1_0),.dout(w_dff_B_zGWPKchG6_0),.clk(gclk));
	jdff dff_B_B4VkixQz7_0(.din(w_dff_B_zGWPKchG6_0),.dout(w_dff_B_B4VkixQz7_0),.clk(gclk));
	jdff dff_B_AZZAoUlg3_0(.din(w_dff_B_B4VkixQz7_0),.dout(w_dff_B_AZZAoUlg3_0),.clk(gclk));
	jdff dff_B_fcLtakTq9_0(.din(w_dff_B_AZZAoUlg3_0),.dout(w_dff_B_fcLtakTq9_0),.clk(gclk));
	jdff dff_B_GcsI27qI6_0(.din(w_dff_B_fcLtakTq9_0),.dout(w_dff_B_GcsI27qI6_0),.clk(gclk));
	jdff dff_B_79uVL9sZ7_0(.din(w_dff_B_GcsI27qI6_0),.dout(w_dff_B_79uVL9sZ7_0),.clk(gclk));
	jdff dff_B_io6zSyI37_0(.din(w_dff_B_79uVL9sZ7_0),.dout(w_dff_B_io6zSyI37_0),.clk(gclk));
	jdff dff_B_ct3BczfG9_0(.din(w_dff_B_io6zSyI37_0),.dout(w_dff_B_ct3BczfG9_0),.clk(gclk));
	jdff dff_B_NnkrXpG68_0(.din(w_dff_B_ct3BczfG9_0),.dout(w_dff_B_NnkrXpG68_0),.clk(gclk));
	jdff dff_B_82bDnHis2_0(.din(w_dff_B_NnkrXpG68_0),.dout(w_dff_B_82bDnHis2_0),.clk(gclk));
	jdff dff_B_m7a7MgSH4_0(.din(w_dff_B_82bDnHis2_0),.dout(w_dff_B_m7a7MgSH4_0),.clk(gclk));
	jdff dff_B_eMbb14EB4_0(.din(w_dff_B_m7a7MgSH4_0),.dout(w_dff_B_eMbb14EB4_0),.clk(gclk));
	jdff dff_B_AJnunAIe4_0(.din(w_dff_B_eMbb14EB4_0),.dout(w_dff_B_AJnunAIe4_0),.clk(gclk));
	jdff dff_B_mnp17btZ2_0(.din(w_dff_B_AJnunAIe4_0),.dout(w_dff_B_mnp17btZ2_0),.clk(gclk));
	jdff dff_B_Zd9dDlEE4_0(.din(w_dff_B_mnp17btZ2_0),.dout(w_dff_B_Zd9dDlEE4_0),.clk(gclk));
	jdff dff_B_24QlirJ28_0(.din(w_dff_B_Zd9dDlEE4_0),.dout(w_dff_B_24QlirJ28_0),.clk(gclk));
	jdff dff_B_p5IueDTz1_0(.din(w_dff_B_24QlirJ28_0),.dout(w_dff_B_p5IueDTz1_0),.clk(gclk));
	jdff dff_B_vbTSAZ3x6_0(.din(w_dff_B_p5IueDTz1_0),.dout(w_dff_B_vbTSAZ3x6_0),.clk(gclk));
	jdff dff_B_FmpoJySX5_0(.din(w_dff_B_vbTSAZ3x6_0),.dout(w_dff_B_FmpoJySX5_0),.clk(gclk));
	jdff dff_B_6clVDe9u5_0(.din(w_dff_B_FmpoJySX5_0),.dout(w_dff_B_6clVDe9u5_0),.clk(gclk));
	jdff dff_B_5TRClnVL4_0(.din(w_dff_B_6clVDe9u5_0),.dout(w_dff_B_5TRClnVL4_0),.clk(gclk));
	jdff dff_B_2MPg8mNX6_0(.din(w_dff_B_5TRClnVL4_0),.dout(w_dff_B_2MPg8mNX6_0),.clk(gclk));
	jdff dff_B_ipLr3u053_0(.din(w_dff_B_2MPg8mNX6_0),.dout(w_dff_B_ipLr3u053_0),.clk(gclk));
	jdff dff_B_SP6w6syZ5_0(.din(w_dff_B_ipLr3u053_0),.dout(w_dff_B_SP6w6syZ5_0),.clk(gclk));
	jdff dff_B_yk90ZYBF7_0(.din(w_dff_B_SP6w6syZ5_0),.dout(w_dff_B_yk90ZYBF7_0),.clk(gclk));
	jdff dff_B_6WPlQnjn3_0(.din(w_dff_B_yk90ZYBF7_0),.dout(w_dff_B_6WPlQnjn3_0),.clk(gclk));
	jdff dff_B_3Psgfeor4_0(.din(w_dff_B_6WPlQnjn3_0),.dout(w_dff_B_3Psgfeor4_0),.clk(gclk));
	jdff dff_B_GzQJe2hd3_0(.din(w_dff_B_3Psgfeor4_0),.dout(w_dff_B_GzQJe2hd3_0),.clk(gclk));
	jdff dff_B_fFgdS6yr2_0(.din(w_dff_B_GzQJe2hd3_0),.dout(w_dff_B_fFgdS6yr2_0),.clk(gclk));
	jdff dff_B_wCqYeAoU5_0(.din(w_dff_B_fFgdS6yr2_0),.dout(w_dff_B_wCqYeAoU5_0),.clk(gclk));
	jdff dff_B_2QkoEW2i9_0(.din(w_dff_B_wCqYeAoU5_0),.dout(w_dff_B_2QkoEW2i9_0),.clk(gclk));
	jdff dff_B_NEl2t2WK5_0(.din(w_dff_B_2QkoEW2i9_0),.dout(w_dff_B_NEl2t2WK5_0),.clk(gclk));
	jdff dff_B_jkdSfD8o0_0(.din(w_dff_B_NEl2t2WK5_0),.dout(w_dff_B_jkdSfD8o0_0),.clk(gclk));
	jdff dff_B_d9YLOmDB7_0(.din(w_dff_B_jkdSfD8o0_0),.dout(w_dff_B_d9YLOmDB7_0),.clk(gclk));
	jdff dff_B_DhOwyyt05_0(.din(w_dff_B_d9YLOmDB7_0),.dout(w_dff_B_DhOwyyt05_0),.clk(gclk));
	jdff dff_B_W0UFrXYB9_0(.din(n838),.dout(w_dff_B_W0UFrXYB9_0),.clk(gclk));
	jdff dff_B_J89MJakF3_0(.din(w_dff_B_W0UFrXYB9_0),.dout(w_dff_B_J89MJakF3_0),.clk(gclk));
	jdff dff_B_uENGzOBh2_0(.din(w_dff_B_J89MJakF3_0),.dout(w_dff_B_uENGzOBh2_0),.clk(gclk));
	jdff dff_B_Ep7ZbnL90_0(.din(w_dff_B_uENGzOBh2_0),.dout(w_dff_B_Ep7ZbnL90_0),.clk(gclk));
	jdff dff_B_MsEOaw3U3_0(.din(w_dff_B_Ep7ZbnL90_0),.dout(w_dff_B_MsEOaw3U3_0),.clk(gclk));
	jdff dff_B_Z1RMHlHD6_0(.din(w_dff_B_MsEOaw3U3_0),.dout(w_dff_B_Z1RMHlHD6_0),.clk(gclk));
	jdff dff_B_BNmrJpzO8_0(.din(w_dff_B_Z1RMHlHD6_0),.dout(w_dff_B_BNmrJpzO8_0),.clk(gclk));
	jdff dff_B_1mhdemTw3_0(.din(w_dff_B_BNmrJpzO8_0),.dout(w_dff_B_1mhdemTw3_0),.clk(gclk));
	jdff dff_B_8DX3k4f20_0(.din(w_dff_B_1mhdemTw3_0),.dout(w_dff_B_8DX3k4f20_0),.clk(gclk));
	jdff dff_B_acAylcrc9_0(.din(w_dff_B_8DX3k4f20_0),.dout(w_dff_B_acAylcrc9_0),.clk(gclk));
	jdff dff_B_setQDUl23_0(.din(w_dff_B_acAylcrc9_0),.dout(w_dff_B_setQDUl23_0),.clk(gclk));
	jdff dff_B_TC9Jipj27_0(.din(w_dff_B_setQDUl23_0),.dout(w_dff_B_TC9Jipj27_0),.clk(gclk));
	jdff dff_B_9ufmnTMV7_0(.din(w_dff_B_TC9Jipj27_0),.dout(w_dff_B_9ufmnTMV7_0),.clk(gclk));
	jdff dff_B_DMX1dXDT5_0(.din(w_dff_B_9ufmnTMV7_0),.dout(w_dff_B_DMX1dXDT5_0),.clk(gclk));
	jdff dff_B_1bnbnxWi5_0(.din(w_dff_B_DMX1dXDT5_0),.dout(w_dff_B_1bnbnxWi5_0),.clk(gclk));
	jdff dff_B_hYcRO49R2_0(.din(w_dff_B_1bnbnxWi5_0),.dout(w_dff_B_hYcRO49R2_0),.clk(gclk));
	jdff dff_B_QoNs79Ag6_0(.din(w_dff_B_hYcRO49R2_0),.dout(w_dff_B_QoNs79Ag6_0),.clk(gclk));
	jdff dff_B_7CXgmlU11_0(.din(w_dff_B_QoNs79Ag6_0),.dout(w_dff_B_7CXgmlU11_0),.clk(gclk));
	jdff dff_B_O3LNg3lQ4_0(.din(w_dff_B_7CXgmlU11_0),.dout(w_dff_B_O3LNg3lQ4_0),.clk(gclk));
	jdff dff_B_zXATzSmg4_0(.din(w_dff_B_O3LNg3lQ4_0),.dout(w_dff_B_zXATzSmg4_0),.clk(gclk));
	jdff dff_B_DbHnkhoM2_0(.din(w_dff_B_zXATzSmg4_0),.dout(w_dff_B_DbHnkhoM2_0),.clk(gclk));
	jdff dff_B_to6Tc7fS8_0(.din(w_dff_B_DbHnkhoM2_0),.dout(w_dff_B_to6Tc7fS8_0),.clk(gclk));
	jdff dff_B_r3egGGxX3_0(.din(w_dff_B_to6Tc7fS8_0),.dout(w_dff_B_r3egGGxX3_0),.clk(gclk));
	jdff dff_B_ZHEFBFy70_0(.din(w_dff_B_r3egGGxX3_0),.dout(w_dff_B_ZHEFBFy70_0),.clk(gclk));
	jdff dff_B_LGU3LcRJ3_0(.din(w_dff_B_ZHEFBFy70_0),.dout(w_dff_B_LGU3LcRJ3_0),.clk(gclk));
	jdff dff_B_BCCiiD521_0(.din(w_dff_B_LGU3LcRJ3_0),.dout(w_dff_B_BCCiiD521_0),.clk(gclk));
	jdff dff_B_BJ5MHOmb2_0(.din(w_dff_B_BCCiiD521_0),.dout(w_dff_B_BJ5MHOmb2_0),.clk(gclk));
	jdff dff_B_EiHuVkh28_0(.din(w_dff_B_BJ5MHOmb2_0),.dout(w_dff_B_EiHuVkh28_0),.clk(gclk));
	jdff dff_B_9YBHhiIi4_0(.din(w_dff_B_EiHuVkh28_0),.dout(w_dff_B_9YBHhiIi4_0),.clk(gclk));
	jdff dff_B_EzEAjWrM2_0(.din(w_dff_B_9YBHhiIi4_0),.dout(w_dff_B_EzEAjWrM2_0),.clk(gclk));
	jdff dff_B_Jt2KN0hA3_0(.din(w_dff_B_EzEAjWrM2_0),.dout(w_dff_B_Jt2KN0hA3_0),.clk(gclk));
	jdff dff_B_W4sBaM5H5_0(.din(w_dff_B_Jt2KN0hA3_0),.dout(w_dff_B_W4sBaM5H5_0),.clk(gclk));
	jdff dff_B_IIOII2UC9_0(.din(w_dff_B_W4sBaM5H5_0),.dout(w_dff_B_IIOII2UC9_0),.clk(gclk));
	jdff dff_B_JCf1MSee8_0(.din(w_dff_B_IIOII2UC9_0),.dout(w_dff_B_JCf1MSee8_0),.clk(gclk));
	jdff dff_B_Xi9YM6Iy1_0(.din(w_dff_B_JCf1MSee8_0),.dout(w_dff_B_Xi9YM6Iy1_0),.clk(gclk));
	jdff dff_B_Sg4YK8vp2_0(.din(w_dff_B_Xi9YM6Iy1_0),.dout(w_dff_B_Sg4YK8vp2_0),.clk(gclk));
	jdff dff_B_0UMBkUdK0_0(.din(w_dff_B_Sg4YK8vp2_0),.dout(w_dff_B_0UMBkUdK0_0),.clk(gclk));
	jdff dff_B_YX7CqXs84_0(.din(w_dff_B_0UMBkUdK0_0),.dout(w_dff_B_YX7CqXs84_0),.clk(gclk));
	jdff dff_B_w9rZFh0P2_0(.din(w_dff_B_YX7CqXs84_0),.dout(w_dff_B_w9rZFh0P2_0),.clk(gclk));
	jdff dff_B_nRU76yD61_0(.din(w_dff_B_w9rZFh0P2_0),.dout(w_dff_B_nRU76yD61_0),.clk(gclk));
	jdff dff_B_7QoyaaUP6_0(.din(w_dff_B_nRU76yD61_0),.dout(w_dff_B_7QoyaaUP6_0),.clk(gclk));
	jdff dff_B_xUbN0nya1_0(.din(w_dff_B_7QoyaaUP6_0),.dout(w_dff_B_xUbN0nya1_0),.clk(gclk));
	jdff dff_B_2ioswjf45_0(.din(w_dff_B_xUbN0nya1_0),.dout(w_dff_B_2ioswjf45_0),.clk(gclk));
	jdff dff_B_vKRXIBIi8_0(.din(w_dff_B_2ioswjf45_0),.dout(w_dff_B_vKRXIBIi8_0),.clk(gclk));
	jdff dff_B_0BiWx5La1_0(.din(w_dff_B_vKRXIBIi8_0),.dout(w_dff_B_0BiWx5La1_0),.clk(gclk));
	jdff dff_B_429sELnG5_0(.din(w_dff_B_0BiWx5La1_0),.dout(w_dff_B_429sELnG5_0),.clk(gclk));
	jdff dff_B_B8sF3QoZ6_0(.din(w_dff_B_429sELnG5_0),.dout(w_dff_B_B8sF3QoZ6_0),.clk(gclk));
	jdff dff_B_VVKliftS9_0(.din(w_dff_B_B8sF3QoZ6_0),.dout(w_dff_B_VVKliftS9_0),.clk(gclk));
	jdff dff_B_hC77Gjo20_0(.din(w_dff_B_VVKliftS9_0),.dout(w_dff_B_hC77Gjo20_0),.clk(gclk));
	jdff dff_B_rdLexDQC7_0(.din(w_dff_B_hC77Gjo20_0),.dout(w_dff_B_rdLexDQC7_0),.clk(gclk));
	jdff dff_B_Kab0bn8L2_0(.din(w_dff_B_rdLexDQC7_0),.dout(w_dff_B_Kab0bn8L2_0),.clk(gclk));
	jdff dff_B_yP51ITwX7_0(.din(w_dff_B_Kab0bn8L2_0),.dout(w_dff_B_yP51ITwX7_0),.clk(gclk));
	jdff dff_B_73RWRYjg9_0(.din(w_dff_B_yP51ITwX7_0),.dout(w_dff_B_73RWRYjg9_0),.clk(gclk));
	jdff dff_B_D42ptgaw7_0(.din(w_dff_B_73RWRYjg9_0),.dout(w_dff_B_D42ptgaw7_0),.clk(gclk));
	jdff dff_B_l8pJKvwU4_0(.din(w_dff_B_D42ptgaw7_0),.dout(w_dff_B_l8pJKvwU4_0),.clk(gclk));
	jdff dff_B_KbOYTM4W4_0(.din(w_dff_B_l8pJKvwU4_0),.dout(w_dff_B_KbOYTM4W4_0),.clk(gclk));
	jdff dff_B_udGSE7zz4_0(.din(w_dff_B_KbOYTM4W4_0),.dout(w_dff_B_udGSE7zz4_0),.clk(gclk));
	jdff dff_B_eBtTxwtr5_0(.din(w_dff_B_udGSE7zz4_0),.dout(w_dff_B_eBtTxwtr5_0),.clk(gclk));
	jdff dff_B_oJ7lkHKB1_0(.din(w_dff_B_eBtTxwtr5_0),.dout(w_dff_B_oJ7lkHKB1_0),.clk(gclk));
	jdff dff_B_pYbb9aiH4_0(.din(w_dff_B_oJ7lkHKB1_0),.dout(w_dff_B_pYbb9aiH4_0),.clk(gclk));
	jdff dff_B_tsHHG2pn2_0(.din(w_dff_B_pYbb9aiH4_0),.dout(w_dff_B_tsHHG2pn2_0),.clk(gclk));
	jdff dff_B_1GjYhWup4_0(.din(w_dff_B_tsHHG2pn2_0),.dout(w_dff_B_1GjYhWup4_0),.clk(gclk));
	jdff dff_B_2va0z3ho3_0(.din(w_dff_B_1GjYhWup4_0),.dout(w_dff_B_2va0z3ho3_0),.clk(gclk));
	jdff dff_B_ZzbnFaOZ9_0(.din(w_dff_B_2va0z3ho3_0),.dout(w_dff_B_ZzbnFaOZ9_0),.clk(gclk));
	jdff dff_B_Uoor99ov9_0(.din(w_dff_B_ZzbnFaOZ9_0),.dout(w_dff_B_Uoor99ov9_0),.clk(gclk));
	jdff dff_B_mwaZx1Pw1_0(.din(w_dff_B_Uoor99ov9_0),.dout(w_dff_B_mwaZx1Pw1_0),.clk(gclk));
	jdff dff_B_KE9Wtkoq3_0(.din(w_dff_B_mwaZx1Pw1_0),.dout(w_dff_B_KE9Wtkoq3_0),.clk(gclk));
	jdff dff_B_neOY6BFx7_0(.din(w_dff_B_KE9Wtkoq3_0),.dout(w_dff_B_neOY6BFx7_0),.clk(gclk));
	jdff dff_B_LXqYXlFk4_0(.din(w_dff_B_neOY6BFx7_0),.dout(w_dff_B_LXqYXlFk4_0),.clk(gclk));
	jdff dff_B_crEd0d0B0_0(.din(w_dff_B_LXqYXlFk4_0),.dout(w_dff_B_crEd0d0B0_0),.clk(gclk));
	jdff dff_B_JVQanGuL2_0(.din(w_dff_B_crEd0d0B0_0),.dout(w_dff_B_JVQanGuL2_0),.clk(gclk));
	jdff dff_B_87ABA4220_0(.din(w_dff_B_JVQanGuL2_0),.dout(w_dff_B_87ABA4220_0),.clk(gclk));
	jdff dff_B_lWIE4kdJ0_0(.din(w_dff_B_87ABA4220_0),.dout(w_dff_B_lWIE4kdJ0_0),.clk(gclk));
	jdff dff_B_uUxQQKLa1_0(.din(w_dff_B_lWIE4kdJ0_0),.dout(w_dff_B_uUxQQKLa1_0),.clk(gclk));
	jdff dff_B_djJxNpry8_0(.din(w_dff_B_uUxQQKLa1_0),.dout(w_dff_B_djJxNpry8_0),.clk(gclk));
	jdff dff_B_vM1UBh3N6_0(.din(n844),.dout(w_dff_B_vM1UBh3N6_0),.clk(gclk));
	jdff dff_B_bkQrWo0p1_0(.din(w_dff_B_vM1UBh3N6_0),.dout(w_dff_B_bkQrWo0p1_0),.clk(gclk));
	jdff dff_B_zLM4uuE45_0(.din(w_dff_B_bkQrWo0p1_0),.dout(w_dff_B_zLM4uuE45_0),.clk(gclk));
	jdff dff_B_bOWF5lqG0_0(.din(w_dff_B_zLM4uuE45_0),.dout(w_dff_B_bOWF5lqG0_0),.clk(gclk));
	jdff dff_B_LikD3aIF0_0(.din(w_dff_B_bOWF5lqG0_0),.dout(w_dff_B_LikD3aIF0_0),.clk(gclk));
	jdff dff_B_zM8ZWNiA6_0(.din(w_dff_B_LikD3aIF0_0),.dout(w_dff_B_zM8ZWNiA6_0),.clk(gclk));
	jdff dff_B_bHdvkmT64_0(.din(w_dff_B_zM8ZWNiA6_0),.dout(w_dff_B_bHdvkmT64_0),.clk(gclk));
	jdff dff_B_vcWeeyN54_0(.din(w_dff_B_bHdvkmT64_0),.dout(w_dff_B_vcWeeyN54_0),.clk(gclk));
	jdff dff_B_4JebWuIn6_0(.din(w_dff_B_vcWeeyN54_0),.dout(w_dff_B_4JebWuIn6_0),.clk(gclk));
	jdff dff_B_FdzOElnO1_0(.din(w_dff_B_4JebWuIn6_0),.dout(w_dff_B_FdzOElnO1_0),.clk(gclk));
	jdff dff_B_oJrZnA5B5_0(.din(w_dff_B_FdzOElnO1_0),.dout(w_dff_B_oJrZnA5B5_0),.clk(gclk));
	jdff dff_B_KuaKaXw61_0(.din(w_dff_B_oJrZnA5B5_0),.dout(w_dff_B_KuaKaXw61_0),.clk(gclk));
	jdff dff_B_7QB61Y7k8_0(.din(w_dff_B_KuaKaXw61_0),.dout(w_dff_B_7QB61Y7k8_0),.clk(gclk));
	jdff dff_B_6Zl32GTW5_0(.din(w_dff_B_7QB61Y7k8_0),.dout(w_dff_B_6Zl32GTW5_0),.clk(gclk));
	jdff dff_B_WiI8Ey2i9_0(.din(w_dff_B_6Zl32GTW5_0),.dout(w_dff_B_WiI8Ey2i9_0),.clk(gclk));
	jdff dff_B_Bn0J8M762_0(.din(w_dff_B_WiI8Ey2i9_0),.dout(w_dff_B_Bn0J8M762_0),.clk(gclk));
	jdff dff_B_F93XNt5i5_0(.din(w_dff_B_Bn0J8M762_0),.dout(w_dff_B_F93XNt5i5_0),.clk(gclk));
	jdff dff_B_FXkoKMnn3_0(.din(w_dff_B_F93XNt5i5_0),.dout(w_dff_B_FXkoKMnn3_0),.clk(gclk));
	jdff dff_B_7MmMkRQb7_0(.din(w_dff_B_FXkoKMnn3_0),.dout(w_dff_B_7MmMkRQb7_0),.clk(gclk));
	jdff dff_B_tmhoApgT1_0(.din(w_dff_B_7MmMkRQb7_0),.dout(w_dff_B_tmhoApgT1_0),.clk(gclk));
	jdff dff_B_IaZj5f5E6_0(.din(w_dff_B_tmhoApgT1_0),.dout(w_dff_B_IaZj5f5E6_0),.clk(gclk));
	jdff dff_B_MdaEq8cC1_0(.din(w_dff_B_IaZj5f5E6_0),.dout(w_dff_B_MdaEq8cC1_0),.clk(gclk));
	jdff dff_B_omNQpwgx2_0(.din(w_dff_B_MdaEq8cC1_0),.dout(w_dff_B_omNQpwgx2_0),.clk(gclk));
	jdff dff_B_OMXlPSJV4_0(.din(w_dff_B_omNQpwgx2_0),.dout(w_dff_B_OMXlPSJV4_0),.clk(gclk));
	jdff dff_B_DFUJyOSU3_0(.din(w_dff_B_OMXlPSJV4_0),.dout(w_dff_B_DFUJyOSU3_0),.clk(gclk));
	jdff dff_B_XhhwdUIa1_0(.din(w_dff_B_DFUJyOSU3_0),.dout(w_dff_B_XhhwdUIa1_0),.clk(gclk));
	jdff dff_B_wvHW04T62_0(.din(w_dff_B_XhhwdUIa1_0),.dout(w_dff_B_wvHW04T62_0),.clk(gclk));
	jdff dff_B_qWTm3oSy6_0(.din(w_dff_B_wvHW04T62_0),.dout(w_dff_B_qWTm3oSy6_0),.clk(gclk));
	jdff dff_B_fCIlhNPU1_0(.din(w_dff_B_qWTm3oSy6_0),.dout(w_dff_B_fCIlhNPU1_0),.clk(gclk));
	jdff dff_B_81eeMq5X9_0(.din(w_dff_B_fCIlhNPU1_0),.dout(w_dff_B_81eeMq5X9_0),.clk(gclk));
	jdff dff_B_xnChlfi34_0(.din(w_dff_B_81eeMq5X9_0),.dout(w_dff_B_xnChlfi34_0),.clk(gclk));
	jdff dff_B_Bjcvqyle8_0(.din(w_dff_B_xnChlfi34_0),.dout(w_dff_B_Bjcvqyle8_0),.clk(gclk));
	jdff dff_B_KAcvpLMI0_0(.din(w_dff_B_Bjcvqyle8_0),.dout(w_dff_B_KAcvpLMI0_0),.clk(gclk));
	jdff dff_B_c4IxKS9W8_0(.din(w_dff_B_KAcvpLMI0_0),.dout(w_dff_B_c4IxKS9W8_0),.clk(gclk));
	jdff dff_B_I6CjZlZ28_0(.din(w_dff_B_c4IxKS9W8_0),.dout(w_dff_B_I6CjZlZ28_0),.clk(gclk));
	jdff dff_B_D1jGAaK66_0(.din(w_dff_B_I6CjZlZ28_0),.dout(w_dff_B_D1jGAaK66_0),.clk(gclk));
	jdff dff_B_zDv66KOB8_0(.din(w_dff_B_D1jGAaK66_0),.dout(w_dff_B_zDv66KOB8_0),.clk(gclk));
	jdff dff_B_GGYLst9G5_0(.din(w_dff_B_zDv66KOB8_0),.dout(w_dff_B_GGYLst9G5_0),.clk(gclk));
	jdff dff_B_bfxEIaek1_0(.din(w_dff_B_GGYLst9G5_0),.dout(w_dff_B_bfxEIaek1_0),.clk(gclk));
	jdff dff_B_8UT2cDNx0_0(.din(w_dff_B_bfxEIaek1_0),.dout(w_dff_B_8UT2cDNx0_0),.clk(gclk));
	jdff dff_B_eA4AblRc4_0(.din(w_dff_B_8UT2cDNx0_0),.dout(w_dff_B_eA4AblRc4_0),.clk(gclk));
	jdff dff_B_YXCUUzBE3_0(.din(w_dff_B_eA4AblRc4_0),.dout(w_dff_B_YXCUUzBE3_0),.clk(gclk));
	jdff dff_B_RSXaTjSB4_0(.din(w_dff_B_YXCUUzBE3_0),.dout(w_dff_B_RSXaTjSB4_0),.clk(gclk));
	jdff dff_B_is0svj5R6_0(.din(w_dff_B_RSXaTjSB4_0),.dout(w_dff_B_is0svj5R6_0),.clk(gclk));
	jdff dff_B_HYzHSGIL5_0(.din(w_dff_B_is0svj5R6_0),.dout(w_dff_B_HYzHSGIL5_0),.clk(gclk));
	jdff dff_B_8axesWXT6_0(.din(w_dff_B_HYzHSGIL5_0),.dout(w_dff_B_8axesWXT6_0),.clk(gclk));
	jdff dff_B_4KtXTPat7_0(.din(w_dff_B_8axesWXT6_0),.dout(w_dff_B_4KtXTPat7_0),.clk(gclk));
	jdff dff_B_qVdVgnM63_0(.din(w_dff_B_4KtXTPat7_0),.dout(w_dff_B_qVdVgnM63_0),.clk(gclk));
	jdff dff_B_mD6PHSB68_0(.din(w_dff_B_qVdVgnM63_0),.dout(w_dff_B_mD6PHSB68_0),.clk(gclk));
	jdff dff_B_kF0Imev28_0(.din(w_dff_B_mD6PHSB68_0),.dout(w_dff_B_kF0Imev28_0),.clk(gclk));
	jdff dff_B_x7L4bWiu2_0(.din(w_dff_B_kF0Imev28_0),.dout(w_dff_B_x7L4bWiu2_0),.clk(gclk));
	jdff dff_B_DxTf15X22_0(.din(w_dff_B_x7L4bWiu2_0),.dout(w_dff_B_DxTf15X22_0),.clk(gclk));
	jdff dff_B_Spsqco3H4_0(.din(w_dff_B_DxTf15X22_0),.dout(w_dff_B_Spsqco3H4_0),.clk(gclk));
	jdff dff_B_IgtOKXGT2_0(.din(w_dff_B_Spsqco3H4_0),.dout(w_dff_B_IgtOKXGT2_0),.clk(gclk));
	jdff dff_B_qEgsXsUg9_0(.din(w_dff_B_IgtOKXGT2_0),.dout(w_dff_B_qEgsXsUg9_0),.clk(gclk));
	jdff dff_B_ov6Io3DL5_0(.din(w_dff_B_qEgsXsUg9_0),.dout(w_dff_B_ov6Io3DL5_0),.clk(gclk));
	jdff dff_B_iYpslwJ14_0(.din(w_dff_B_ov6Io3DL5_0),.dout(w_dff_B_iYpslwJ14_0),.clk(gclk));
	jdff dff_B_BOwiWPIo6_0(.din(w_dff_B_iYpslwJ14_0),.dout(w_dff_B_BOwiWPIo6_0),.clk(gclk));
	jdff dff_B_z94sYFJN8_0(.din(w_dff_B_BOwiWPIo6_0),.dout(w_dff_B_z94sYFJN8_0),.clk(gclk));
	jdff dff_B_KfH6SYsc1_0(.din(w_dff_B_z94sYFJN8_0),.dout(w_dff_B_KfH6SYsc1_0),.clk(gclk));
	jdff dff_B_IWC8jTjB4_0(.din(w_dff_B_KfH6SYsc1_0),.dout(w_dff_B_IWC8jTjB4_0),.clk(gclk));
	jdff dff_B_trIvCV9t3_0(.din(w_dff_B_IWC8jTjB4_0),.dout(w_dff_B_trIvCV9t3_0),.clk(gclk));
	jdff dff_B_7X5463831_0(.din(w_dff_B_trIvCV9t3_0),.dout(w_dff_B_7X5463831_0),.clk(gclk));
	jdff dff_B_snlhun002_0(.din(w_dff_B_7X5463831_0),.dout(w_dff_B_snlhun002_0),.clk(gclk));
	jdff dff_B_Fc8BozXS5_0(.din(w_dff_B_snlhun002_0),.dout(w_dff_B_Fc8BozXS5_0),.clk(gclk));
	jdff dff_B_znfAO9BJ3_0(.din(w_dff_B_Fc8BozXS5_0),.dout(w_dff_B_znfAO9BJ3_0),.clk(gclk));
	jdff dff_B_CcKhd9Sx9_0(.din(w_dff_B_znfAO9BJ3_0),.dout(w_dff_B_CcKhd9Sx9_0),.clk(gclk));
	jdff dff_B_nprRhfRi8_0(.din(w_dff_B_CcKhd9Sx9_0),.dout(w_dff_B_nprRhfRi8_0),.clk(gclk));
	jdff dff_B_9AY16yQp7_0(.din(w_dff_B_nprRhfRi8_0),.dout(w_dff_B_9AY16yQp7_0),.clk(gclk));
	jdff dff_B_dHVmP7kB3_0(.din(w_dff_B_9AY16yQp7_0),.dout(w_dff_B_dHVmP7kB3_0),.clk(gclk));
	jdff dff_B_uQCRUEsm3_0(.din(w_dff_B_dHVmP7kB3_0),.dout(w_dff_B_uQCRUEsm3_0),.clk(gclk));
	jdff dff_B_h1gGIhqh6_0(.din(w_dff_B_uQCRUEsm3_0),.dout(w_dff_B_h1gGIhqh6_0),.clk(gclk));
	jdff dff_B_iuEXXVGa8_0(.din(w_dff_B_h1gGIhqh6_0),.dout(w_dff_B_iuEXXVGa8_0),.clk(gclk));
	jdff dff_B_iwr7AWA66_0(.din(w_dff_B_iuEXXVGa8_0),.dout(w_dff_B_iwr7AWA66_0),.clk(gclk));
	jdff dff_B_yAqiSVRh4_0(.din(w_dff_B_iwr7AWA66_0),.dout(w_dff_B_yAqiSVRh4_0),.clk(gclk));
	jdff dff_B_uNf2OqZk3_0(.din(w_dff_B_yAqiSVRh4_0),.dout(w_dff_B_uNf2OqZk3_0),.clk(gclk));
	jdff dff_B_9HttA2JE1_0(.din(n850),.dout(w_dff_B_9HttA2JE1_0),.clk(gclk));
	jdff dff_B_00ffjm2E0_0(.din(w_dff_B_9HttA2JE1_0),.dout(w_dff_B_00ffjm2E0_0),.clk(gclk));
	jdff dff_B_8bUDF9ix8_0(.din(w_dff_B_00ffjm2E0_0),.dout(w_dff_B_8bUDF9ix8_0),.clk(gclk));
	jdff dff_B_KfswDMz35_0(.din(w_dff_B_8bUDF9ix8_0),.dout(w_dff_B_KfswDMz35_0),.clk(gclk));
	jdff dff_B_3ApTX3548_0(.din(w_dff_B_KfswDMz35_0),.dout(w_dff_B_3ApTX3548_0),.clk(gclk));
	jdff dff_B_y2TWio1J2_0(.din(w_dff_B_3ApTX3548_0),.dout(w_dff_B_y2TWio1J2_0),.clk(gclk));
	jdff dff_B_xmyoRDTp1_0(.din(w_dff_B_y2TWio1J2_0),.dout(w_dff_B_xmyoRDTp1_0),.clk(gclk));
	jdff dff_B_UijIED8f2_0(.din(w_dff_B_xmyoRDTp1_0),.dout(w_dff_B_UijIED8f2_0),.clk(gclk));
	jdff dff_B_KmQb0IHD9_0(.din(w_dff_B_UijIED8f2_0),.dout(w_dff_B_KmQb0IHD9_0),.clk(gclk));
	jdff dff_B_11gI7d5m0_0(.din(w_dff_B_KmQb0IHD9_0),.dout(w_dff_B_11gI7d5m0_0),.clk(gclk));
	jdff dff_B_QsOjsc4Y2_0(.din(w_dff_B_11gI7d5m0_0),.dout(w_dff_B_QsOjsc4Y2_0),.clk(gclk));
	jdff dff_B_LTjmnrJO1_0(.din(w_dff_B_QsOjsc4Y2_0),.dout(w_dff_B_LTjmnrJO1_0),.clk(gclk));
	jdff dff_B_zSrSj8Fp6_0(.din(w_dff_B_LTjmnrJO1_0),.dout(w_dff_B_zSrSj8Fp6_0),.clk(gclk));
	jdff dff_B_DXl8iyb68_0(.din(w_dff_B_zSrSj8Fp6_0),.dout(w_dff_B_DXl8iyb68_0),.clk(gclk));
	jdff dff_B_53UoUw6A6_0(.din(w_dff_B_DXl8iyb68_0),.dout(w_dff_B_53UoUw6A6_0),.clk(gclk));
	jdff dff_B_9Q7JBnMj2_0(.din(w_dff_B_53UoUw6A6_0),.dout(w_dff_B_9Q7JBnMj2_0),.clk(gclk));
	jdff dff_B_MPkAfAVI9_0(.din(w_dff_B_9Q7JBnMj2_0),.dout(w_dff_B_MPkAfAVI9_0),.clk(gclk));
	jdff dff_B_RjhTeT1N1_0(.din(w_dff_B_MPkAfAVI9_0),.dout(w_dff_B_RjhTeT1N1_0),.clk(gclk));
	jdff dff_B_rpzL0iEf5_0(.din(w_dff_B_RjhTeT1N1_0),.dout(w_dff_B_rpzL0iEf5_0),.clk(gclk));
	jdff dff_B_jtfNxXVo2_0(.din(w_dff_B_rpzL0iEf5_0),.dout(w_dff_B_jtfNxXVo2_0),.clk(gclk));
	jdff dff_B_epiKvRPA7_0(.din(w_dff_B_jtfNxXVo2_0),.dout(w_dff_B_epiKvRPA7_0),.clk(gclk));
	jdff dff_B_NYAa6HbO8_0(.din(w_dff_B_epiKvRPA7_0),.dout(w_dff_B_NYAa6HbO8_0),.clk(gclk));
	jdff dff_B_wrmKRBuO2_0(.din(w_dff_B_NYAa6HbO8_0),.dout(w_dff_B_wrmKRBuO2_0),.clk(gclk));
	jdff dff_B_epJUvQwS0_0(.din(w_dff_B_wrmKRBuO2_0),.dout(w_dff_B_epJUvQwS0_0),.clk(gclk));
	jdff dff_B_UkRbA1kW0_0(.din(w_dff_B_epJUvQwS0_0),.dout(w_dff_B_UkRbA1kW0_0),.clk(gclk));
	jdff dff_B_hUiR4VQm3_0(.din(w_dff_B_UkRbA1kW0_0),.dout(w_dff_B_hUiR4VQm3_0),.clk(gclk));
	jdff dff_B_eL98MWxO1_0(.din(w_dff_B_hUiR4VQm3_0),.dout(w_dff_B_eL98MWxO1_0),.clk(gclk));
	jdff dff_B_Q4DkU52J5_0(.din(w_dff_B_eL98MWxO1_0),.dout(w_dff_B_Q4DkU52J5_0),.clk(gclk));
	jdff dff_B_YV1gapoO4_0(.din(w_dff_B_Q4DkU52J5_0),.dout(w_dff_B_YV1gapoO4_0),.clk(gclk));
	jdff dff_B_OalLZ1mB6_0(.din(w_dff_B_YV1gapoO4_0),.dout(w_dff_B_OalLZ1mB6_0),.clk(gclk));
	jdff dff_B_7S2EpBCa6_0(.din(w_dff_B_OalLZ1mB6_0),.dout(w_dff_B_7S2EpBCa6_0),.clk(gclk));
	jdff dff_B_8DTpE4Zp1_0(.din(w_dff_B_7S2EpBCa6_0),.dout(w_dff_B_8DTpE4Zp1_0),.clk(gclk));
	jdff dff_B_0Vln8Pqp2_0(.din(w_dff_B_8DTpE4Zp1_0),.dout(w_dff_B_0Vln8Pqp2_0),.clk(gclk));
	jdff dff_B_AdyZIk417_0(.din(w_dff_B_0Vln8Pqp2_0),.dout(w_dff_B_AdyZIk417_0),.clk(gclk));
	jdff dff_B_iiHa9ajV1_0(.din(w_dff_B_AdyZIk417_0),.dout(w_dff_B_iiHa9ajV1_0),.clk(gclk));
	jdff dff_B_HHDt0loH9_0(.din(w_dff_B_iiHa9ajV1_0),.dout(w_dff_B_HHDt0loH9_0),.clk(gclk));
	jdff dff_B_PCcJpXXW3_0(.din(w_dff_B_HHDt0loH9_0),.dout(w_dff_B_PCcJpXXW3_0),.clk(gclk));
	jdff dff_B_8h4cd8Ej2_0(.din(w_dff_B_PCcJpXXW3_0),.dout(w_dff_B_8h4cd8Ej2_0),.clk(gclk));
	jdff dff_B_vmtII7zd4_0(.din(w_dff_B_8h4cd8Ej2_0),.dout(w_dff_B_vmtII7zd4_0),.clk(gclk));
	jdff dff_B_5GZcVb409_0(.din(w_dff_B_vmtII7zd4_0),.dout(w_dff_B_5GZcVb409_0),.clk(gclk));
	jdff dff_B_IuWpCWOI4_0(.din(w_dff_B_5GZcVb409_0),.dout(w_dff_B_IuWpCWOI4_0),.clk(gclk));
	jdff dff_B_vwhblVu44_0(.din(w_dff_B_IuWpCWOI4_0),.dout(w_dff_B_vwhblVu44_0),.clk(gclk));
	jdff dff_B_01JVspxS2_0(.din(w_dff_B_vwhblVu44_0),.dout(w_dff_B_01JVspxS2_0),.clk(gclk));
	jdff dff_B_fUUt94jj4_0(.din(w_dff_B_01JVspxS2_0),.dout(w_dff_B_fUUt94jj4_0),.clk(gclk));
	jdff dff_B_AMBEo5So0_0(.din(w_dff_B_fUUt94jj4_0),.dout(w_dff_B_AMBEo5So0_0),.clk(gclk));
	jdff dff_B_GrQU66uW6_0(.din(w_dff_B_AMBEo5So0_0),.dout(w_dff_B_GrQU66uW6_0),.clk(gclk));
	jdff dff_B_dJ0ONYrp8_0(.din(w_dff_B_GrQU66uW6_0),.dout(w_dff_B_dJ0ONYrp8_0),.clk(gclk));
	jdff dff_B_mfVQhXaw7_0(.din(w_dff_B_dJ0ONYrp8_0),.dout(w_dff_B_mfVQhXaw7_0),.clk(gclk));
	jdff dff_B_ztTZe4VO4_0(.din(w_dff_B_mfVQhXaw7_0),.dout(w_dff_B_ztTZe4VO4_0),.clk(gclk));
	jdff dff_B_UdbuoscS3_0(.din(w_dff_B_ztTZe4VO4_0),.dout(w_dff_B_UdbuoscS3_0),.clk(gclk));
	jdff dff_B_qRYVwjpB6_0(.din(w_dff_B_UdbuoscS3_0),.dout(w_dff_B_qRYVwjpB6_0),.clk(gclk));
	jdff dff_B_bI7CO9ur3_0(.din(w_dff_B_qRYVwjpB6_0),.dout(w_dff_B_bI7CO9ur3_0),.clk(gclk));
	jdff dff_B_tCIx70BC6_0(.din(w_dff_B_bI7CO9ur3_0),.dout(w_dff_B_tCIx70BC6_0),.clk(gclk));
	jdff dff_B_4X4wSKmW6_0(.din(w_dff_B_tCIx70BC6_0),.dout(w_dff_B_4X4wSKmW6_0),.clk(gclk));
	jdff dff_B_3gUUqtf63_0(.din(w_dff_B_4X4wSKmW6_0),.dout(w_dff_B_3gUUqtf63_0),.clk(gclk));
	jdff dff_B_nUY4KDfq6_0(.din(w_dff_B_3gUUqtf63_0),.dout(w_dff_B_nUY4KDfq6_0),.clk(gclk));
	jdff dff_B_POSGgnGY1_0(.din(w_dff_B_nUY4KDfq6_0),.dout(w_dff_B_POSGgnGY1_0),.clk(gclk));
	jdff dff_B_a0I8Lziu0_0(.din(w_dff_B_POSGgnGY1_0),.dout(w_dff_B_a0I8Lziu0_0),.clk(gclk));
	jdff dff_B_5Y0rdulh0_0(.din(w_dff_B_a0I8Lziu0_0),.dout(w_dff_B_5Y0rdulh0_0),.clk(gclk));
	jdff dff_B_VLP4Z1nt7_0(.din(w_dff_B_5Y0rdulh0_0),.dout(w_dff_B_VLP4Z1nt7_0),.clk(gclk));
	jdff dff_B_5FA1RMFP5_0(.din(w_dff_B_VLP4Z1nt7_0),.dout(w_dff_B_5FA1RMFP5_0),.clk(gclk));
	jdff dff_B_6SH55aU78_0(.din(w_dff_B_5FA1RMFP5_0),.dout(w_dff_B_6SH55aU78_0),.clk(gclk));
	jdff dff_B_FeHhwumd3_0(.din(w_dff_B_6SH55aU78_0),.dout(w_dff_B_FeHhwumd3_0),.clk(gclk));
	jdff dff_B_As6YPZ1T8_0(.din(w_dff_B_FeHhwumd3_0),.dout(w_dff_B_As6YPZ1T8_0),.clk(gclk));
	jdff dff_B_V85dXJTx9_0(.din(w_dff_B_As6YPZ1T8_0),.dout(w_dff_B_V85dXJTx9_0),.clk(gclk));
	jdff dff_B_lD7eShyX9_0(.din(w_dff_B_V85dXJTx9_0),.dout(w_dff_B_lD7eShyX9_0),.clk(gclk));
	jdff dff_B_18Z8L0Bs1_0(.din(w_dff_B_lD7eShyX9_0),.dout(w_dff_B_18Z8L0Bs1_0),.clk(gclk));
	jdff dff_B_wBWQwLiz3_0(.din(w_dff_B_18Z8L0Bs1_0),.dout(w_dff_B_wBWQwLiz3_0),.clk(gclk));
	jdff dff_B_XMZ24YTb2_0(.din(w_dff_B_wBWQwLiz3_0),.dout(w_dff_B_XMZ24YTb2_0),.clk(gclk));
	jdff dff_B_F7tJJUdp9_0(.din(w_dff_B_XMZ24YTb2_0),.dout(w_dff_B_F7tJJUdp9_0),.clk(gclk));
	jdff dff_B_pyH5qzWo2_0(.din(w_dff_B_F7tJJUdp9_0),.dout(w_dff_B_pyH5qzWo2_0),.clk(gclk));
	jdff dff_B_m6NqfXbK2_0(.din(w_dff_B_pyH5qzWo2_0),.dout(w_dff_B_m6NqfXbK2_0),.clk(gclk));
	jdff dff_B_71KChGh51_0(.din(w_dff_B_m6NqfXbK2_0),.dout(w_dff_B_71KChGh51_0),.clk(gclk));
	jdff dff_B_8ADYl05n4_0(.din(w_dff_B_71KChGh51_0),.dout(w_dff_B_8ADYl05n4_0),.clk(gclk));
	jdff dff_B_pFbX0ArR1_0(.din(w_dff_B_8ADYl05n4_0),.dout(w_dff_B_pFbX0ArR1_0),.clk(gclk));
	jdff dff_B_3xJwK9lW5_0(.din(w_dff_B_pFbX0ArR1_0),.dout(w_dff_B_3xJwK9lW5_0),.clk(gclk));
	jdff dff_B_F5vtCGLu7_0(.din(w_dff_B_3xJwK9lW5_0),.dout(w_dff_B_F5vtCGLu7_0),.clk(gclk));
	jdff dff_B_QF5uRPYv9_0(.din(n856),.dout(w_dff_B_QF5uRPYv9_0),.clk(gclk));
	jdff dff_B_Fxna4I119_0(.din(w_dff_B_QF5uRPYv9_0),.dout(w_dff_B_Fxna4I119_0),.clk(gclk));
	jdff dff_B_KiAsrvlZ4_0(.din(w_dff_B_Fxna4I119_0),.dout(w_dff_B_KiAsrvlZ4_0),.clk(gclk));
	jdff dff_B_RHqzMPBN8_0(.din(w_dff_B_KiAsrvlZ4_0),.dout(w_dff_B_RHqzMPBN8_0),.clk(gclk));
	jdff dff_B_C6RKWGWN4_0(.din(w_dff_B_RHqzMPBN8_0),.dout(w_dff_B_C6RKWGWN4_0),.clk(gclk));
	jdff dff_B_SGVKhsLi3_0(.din(w_dff_B_C6RKWGWN4_0),.dout(w_dff_B_SGVKhsLi3_0),.clk(gclk));
	jdff dff_B_rtGeXwMr4_0(.din(w_dff_B_SGVKhsLi3_0),.dout(w_dff_B_rtGeXwMr4_0),.clk(gclk));
	jdff dff_B_vHXhuWGI9_0(.din(w_dff_B_rtGeXwMr4_0),.dout(w_dff_B_vHXhuWGI9_0),.clk(gclk));
	jdff dff_B_kensvvsp9_0(.din(w_dff_B_vHXhuWGI9_0),.dout(w_dff_B_kensvvsp9_0),.clk(gclk));
	jdff dff_B_XKcXItV71_0(.din(w_dff_B_kensvvsp9_0),.dout(w_dff_B_XKcXItV71_0),.clk(gclk));
	jdff dff_B_7yEvBIrM2_0(.din(w_dff_B_XKcXItV71_0),.dout(w_dff_B_7yEvBIrM2_0),.clk(gclk));
	jdff dff_B_sJo82JNR4_0(.din(w_dff_B_7yEvBIrM2_0),.dout(w_dff_B_sJo82JNR4_0),.clk(gclk));
	jdff dff_B_gAOLVwCc6_0(.din(w_dff_B_sJo82JNR4_0),.dout(w_dff_B_gAOLVwCc6_0),.clk(gclk));
	jdff dff_B_pbsApzcG9_0(.din(w_dff_B_gAOLVwCc6_0),.dout(w_dff_B_pbsApzcG9_0),.clk(gclk));
	jdff dff_B_O5VqGE7U3_0(.din(w_dff_B_pbsApzcG9_0),.dout(w_dff_B_O5VqGE7U3_0),.clk(gclk));
	jdff dff_B_CBJcB2gf8_0(.din(w_dff_B_O5VqGE7U3_0),.dout(w_dff_B_CBJcB2gf8_0),.clk(gclk));
	jdff dff_B_NZ2hVoch4_0(.din(w_dff_B_CBJcB2gf8_0),.dout(w_dff_B_NZ2hVoch4_0),.clk(gclk));
	jdff dff_B_On6FOcow9_0(.din(w_dff_B_NZ2hVoch4_0),.dout(w_dff_B_On6FOcow9_0),.clk(gclk));
	jdff dff_B_9rn9yQoh0_0(.din(w_dff_B_On6FOcow9_0),.dout(w_dff_B_9rn9yQoh0_0),.clk(gclk));
	jdff dff_B_q8f9m24X0_0(.din(w_dff_B_9rn9yQoh0_0),.dout(w_dff_B_q8f9m24X0_0),.clk(gclk));
	jdff dff_B_Sjsq87yN4_0(.din(w_dff_B_q8f9m24X0_0),.dout(w_dff_B_Sjsq87yN4_0),.clk(gclk));
	jdff dff_B_L7HN03dK9_0(.din(w_dff_B_Sjsq87yN4_0),.dout(w_dff_B_L7HN03dK9_0),.clk(gclk));
	jdff dff_B_C4wOqSqZ2_0(.din(w_dff_B_L7HN03dK9_0),.dout(w_dff_B_C4wOqSqZ2_0),.clk(gclk));
	jdff dff_B_mHLvCTdP8_0(.din(w_dff_B_C4wOqSqZ2_0),.dout(w_dff_B_mHLvCTdP8_0),.clk(gclk));
	jdff dff_B_93BSnBvH2_0(.din(w_dff_B_mHLvCTdP8_0),.dout(w_dff_B_93BSnBvH2_0),.clk(gclk));
	jdff dff_B_ty1O9y3B4_0(.din(w_dff_B_93BSnBvH2_0),.dout(w_dff_B_ty1O9y3B4_0),.clk(gclk));
	jdff dff_B_bhcrfqRZ0_0(.din(w_dff_B_ty1O9y3B4_0),.dout(w_dff_B_bhcrfqRZ0_0),.clk(gclk));
	jdff dff_B_oBStXrSG2_0(.din(w_dff_B_bhcrfqRZ0_0),.dout(w_dff_B_oBStXrSG2_0),.clk(gclk));
	jdff dff_B_KkurCbps6_0(.din(w_dff_B_oBStXrSG2_0),.dout(w_dff_B_KkurCbps6_0),.clk(gclk));
	jdff dff_B_2Kk6QEAu6_0(.din(w_dff_B_KkurCbps6_0),.dout(w_dff_B_2Kk6QEAu6_0),.clk(gclk));
	jdff dff_B_Jihq6Kvy5_0(.din(w_dff_B_2Kk6QEAu6_0),.dout(w_dff_B_Jihq6Kvy5_0),.clk(gclk));
	jdff dff_B_rn1yAsyk9_0(.din(w_dff_B_Jihq6Kvy5_0),.dout(w_dff_B_rn1yAsyk9_0),.clk(gclk));
	jdff dff_B_sww4Gs9p2_0(.din(w_dff_B_rn1yAsyk9_0),.dout(w_dff_B_sww4Gs9p2_0),.clk(gclk));
	jdff dff_B_sQuyETEw9_0(.din(w_dff_B_sww4Gs9p2_0),.dout(w_dff_B_sQuyETEw9_0),.clk(gclk));
	jdff dff_B_gfYolZw20_0(.din(w_dff_B_sQuyETEw9_0),.dout(w_dff_B_gfYolZw20_0),.clk(gclk));
	jdff dff_B_tMeyRfLd1_0(.din(w_dff_B_gfYolZw20_0),.dout(w_dff_B_tMeyRfLd1_0),.clk(gclk));
	jdff dff_B_qgAHsxex2_0(.din(w_dff_B_tMeyRfLd1_0),.dout(w_dff_B_qgAHsxex2_0),.clk(gclk));
	jdff dff_B_ccFyZxub5_0(.din(w_dff_B_qgAHsxex2_0),.dout(w_dff_B_ccFyZxub5_0),.clk(gclk));
	jdff dff_B_XpilEKo69_0(.din(w_dff_B_ccFyZxub5_0),.dout(w_dff_B_XpilEKo69_0),.clk(gclk));
	jdff dff_B_UyXbQcRM5_0(.din(w_dff_B_XpilEKo69_0),.dout(w_dff_B_UyXbQcRM5_0),.clk(gclk));
	jdff dff_B_1c7ypbJ28_0(.din(w_dff_B_UyXbQcRM5_0),.dout(w_dff_B_1c7ypbJ28_0),.clk(gclk));
	jdff dff_B_quhpEhkV8_0(.din(w_dff_B_1c7ypbJ28_0),.dout(w_dff_B_quhpEhkV8_0),.clk(gclk));
	jdff dff_B_ZPMSWbcO9_0(.din(w_dff_B_quhpEhkV8_0),.dout(w_dff_B_ZPMSWbcO9_0),.clk(gclk));
	jdff dff_B_FsO2KXY16_0(.din(w_dff_B_ZPMSWbcO9_0),.dout(w_dff_B_FsO2KXY16_0),.clk(gclk));
	jdff dff_B_fK7CgUWz2_0(.din(w_dff_B_FsO2KXY16_0),.dout(w_dff_B_fK7CgUWz2_0),.clk(gclk));
	jdff dff_B_zmt3UkZY0_0(.din(w_dff_B_fK7CgUWz2_0),.dout(w_dff_B_zmt3UkZY0_0),.clk(gclk));
	jdff dff_B_jBxAI2UV6_0(.din(w_dff_B_zmt3UkZY0_0),.dout(w_dff_B_jBxAI2UV6_0),.clk(gclk));
	jdff dff_B_GgBdXz0U9_0(.din(w_dff_B_jBxAI2UV6_0),.dout(w_dff_B_GgBdXz0U9_0),.clk(gclk));
	jdff dff_B_03MzA0Kj3_0(.din(w_dff_B_GgBdXz0U9_0),.dout(w_dff_B_03MzA0Kj3_0),.clk(gclk));
	jdff dff_B_LdqzZI305_0(.din(w_dff_B_03MzA0Kj3_0),.dout(w_dff_B_LdqzZI305_0),.clk(gclk));
	jdff dff_B_o1V6vdcU0_0(.din(w_dff_B_LdqzZI305_0),.dout(w_dff_B_o1V6vdcU0_0),.clk(gclk));
	jdff dff_B_oo9mbzXF5_0(.din(w_dff_B_o1V6vdcU0_0),.dout(w_dff_B_oo9mbzXF5_0),.clk(gclk));
	jdff dff_B_UGdadZeY4_0(.din(w_dff_B_oo9mbzXF5_0),.dout(w_dff_B_UGdadZeY4_0),.clk(gclk));
	jdff dff_B_7DLzRguY7_0(.din(w_dff_B_UGdadZeY4_0),.dout(w_dff_B_7DLzRguY7_0),.clk(gclk));
	jdff dff_B_yV9B1bcm9_0(.din(w_dff_B_7DLzRguY7_0),.dout(w_dff_B_yV9B1bcm9_0),.clk(gclk));
	jdff dff_B_eqWLG71Y1_0(.din(w_dff_B_yV9B1bcm9_0),.dout(w_dff_B_eqWLG71Y1_0),.clk(gclk));
	jdff dff_B_QE3UhFth6_0(.din(w_dff_B_eqWLG71Y1_0),.dout(w_dff_B_QE3UhFth6_0),.clk(gclk));
	jdff dff_B_h6mXwqX92_0(.din(w_dff_B_QE3UhFth6_0),.dout(w_dff_B_h6mXwqX92_0),.clk(gclk));
	jdff dff_B_HMGpbvyO1_0(.din(w_dff_B_h6mXwqX92_0),.dout(w_dff_B_HMGpbvyO1_0),.clk(gclk));
	jdff dff_B_xBCyy7pN0_0(.din(w_dff_B_HMGpbvyO1_0),.dout(w_dff_B_xBCyy7pN0_0),.clk(gclk));
	jdff dff_B_W0K5zfFS9_0(.din(w_dff_B_xBCyy7pN0_0),.dout(w_dff_B_W0K5zfFS9_0),.clk(gclk));
	jdff dff_B_WlIzNb8K2_0(.din(w_dff_B_W0K5zfFS9_0),.dout(w_dff_B_WlIzNb8K2_0),.clk(gclk));
	jdff dff_B_rfckuJU06_0(.din(w_dff_B_WlIzNb8K2_0),.dout(w_dff_B_rfckuJU06_0),.clk(gclk));
	jdff dff_B_Eu8pChFF3_0(.din(w_dff_B_rfckuJU06_0),.dout(w_dff_B_Eu8pChFF3_0),.clk(gclk));
	jdff dff_B_S3pJhBGw0_0(.din(w_dff_B_Eu8pChFF3_0),.dout(w_dff_B_S3pJhBGw0_0),.clk(gclk));
	jdff dff_B_ZJUuqh130_0(.din(w_dff_B_S3pJhBGw0_0),.dout(w_dff_B_ZJUuqh130_0),.clk(gclk));
	jdff dff_B_pIrIQHYH5_0(.din(w_dff_B_ZJUuqh130_0),.dout(w_dff_B_pIrIQHYH5_0),.clk(gclk));
	jdff dff_B_ZluC5sUa1_0(.din(w_dff_B_pIrIQHYH5_0),.dout(w_dff_B_ZluC5sUa1_0),.clk(gclk));
	jdff dff_B_HWZ6xMrk3_0(.din(w_dff_B_ZluC5sUa1_0),.dout(w_dff_B_HWZ6xMrk3_0),.clk(gclk));
	jdff dff_B_ZVI1toyV6_0(.din(w_dff_B_HWZ6xMrk3_0),.dout(w_dff_B_ZVI1toyV6_0),.clk(gclk));
	jdff dff_B_e1ipzYgu1_0(.din(w_dff_B_ZVI1toyV6_0),.dout(w_dff_B_e1ipzYgu1_0),.clk(gclk));
	jdff dff_B_7P2MWAGJ5_0(.din(w_dff_B_e1ipzYgu1_0),.dout(w_dff_B_7P2MWAGJ5_0),.clk(gclk));
	jdff dff_B_eXNMIxO55_0(.din(w_dff_B_7P2MWAGJ5_0),.dout(w_dff_B_eXNMIxO55_0),.clk(gclk));
	jdff dff_B_yypIunip2_0(.din(w_dff_B_eXNMIxO55_0),.dout(w_dff_B_yypIunip2_0),.clk(gclk));
	jdff dff_B_Sy7GwzC87_0(.din(w_dff_B_yypIunip2_0),.dout(w_dff_B_Sy7GwzC87_0),.clk(gclk));
	jdff dff_B_tw0fiH2D9_0(.din(w_dff_B_Sy7GwzC87_0),.dout(w_dff_B_tw0fiH2D9_0),.clk(gclk));
	jdff dff_B_3EYGPgMO0_0(.din(w_dff_B_tw0fiH2D9_0),.dout(w_dff_B_3EYGPgMO0_0),.clk(gclk));
	jdff dff_B_9rEkfsRT6_0(.din(w_dff_B_3EYGPgMO0_0),.dout(w_dff_B_9rEkfsRT6_0),.clk(gclk));
	jdff dff_B_gKW1k3vP2_0(.din(n862),.dout(w_dff_B_gKW1k3vP2_0),.clk(gclk));
	jdff dff_B_WAKMJgJ61_0(.din(w_dff_B_gKW1k3vP2_0),.dout(w_dff_B_WAKMJgJ61_0),.clk(gclk));
	jdff dff_B_9Ci4xdAO5_0(.din(w_dff_B_WAKMJgJ61_0),.dout(w_dff_B_9Ci4xdAO5_0),.clk(gclk));
	jdff dff_B_iA0KSU5s9_0(.din(w_dff_B_9Ci4xdAO5_0),.dout(w_dff_B_iA0KSU5s9_0),.clk(gclk));
	jdff dff_B_tC36WRQz7_0(.din(w_dff_B_iA0KSU5s9_0),.dout(w_dff_B_tC36WRQz7_0),.clk(gclk));
	jdff dff_B_oiCHdwmw3_0(.din(w_dff_B_tC36WRQz7_0),.dout(w_dff_B_oiCHdwmw3_0),.clk(gclk));
	jdff dff_B_Yevv8j603_0(.din(w_dff_B_oiCHdwmw3_0),.dout(w_dff_B_Yevv8j603_0),.clk(gclk));
	jdff dff_B_rGjTU6yF8_0(.din(w_dff_B_Yevv8j603_0),.dout(w_dff_B_rGjTU6yF8_0),.clk(gclk));
	jdff dff_B_yl0RoV968_0(.din(w_dff_B_rGjTU6yF8_0),.dout(w_dff_B_yl0RoV968_0),.clk(gclk));
	jdff dff_B_1Z9pjIVe8_0(.din(w_dff_B_yl0RoV968_0),.dout(w_dff_B_1Z9pjIVe8_0),.clk(gclk));
	jdff dff_B_dQiz3B5P5_0(.din(w_dff_B_1Z9pjIVe8_0),.dout(w_dff_B_dQiz3B5P5_0),.clk(gclk));
	jdff dff_B_eiqSCjH55_0(.din(w_dff_B_dQiz3B5P5_0),.dout(w_dff_B_eiqSCjH55_0),.clk(gclk));
	jdff dff_B_CVwiXj1l3_0(.din(w_dff_B_eiqSCjH55_0),.dout(w_dff_B_CVwiXj1l3_0),.clk(gclk));
	jdff dff_B_06JyOsox7_0(.din(w_dff_B_CVwiXj1l3_0),.dout(w_dff_B_06JyOsox7_0),.clk(gclk));
	jdff dff_B_oq0Ad0me5_0(.din(w_dff_B_06JyOsox7_0),.dout(w_dff_B_oq0Ad0me5_0),.clk(gclk));
	jdff dff_B_jMoSSrJl9_0(.din(w_dff_B_oq0Ad0me5_0),.dout(w_dff_B_jMoSSrJl9_0),.clk(gclk));
	jdff dff_B_axok3U3t6_0(.din(w_dff_B_jMoSSrJl9_0),.dout(w_dff_B_axok3U3t6_0),.clk(gclk));
	jdff dff_B_ySucNKrO5_0(.din(w_dff_B_axok3U3t6_0),.dout(w_dff_B_ySucNKrO5_0),.clk(gclk));
	jdff dff_B_4ThrRtdN4_0(.din(w_dff_B_ySucNKrO5_0),.dout(w_dff_B_4ThrRtdN4_0),.clk(gclk));
	jdff dff_B_DUZzXQVu2_0(.din(w_dff_B_4ThrRtdN4_0),.dout(w_dff_B_DUZzXQVu2_0),.clk(gclk));
	jdff dff_B_okJl0APA3_0(.din(w_dff_B_DUZzXQVu2_0),.dout(w_dff_B_okJl0APA3_0),.clk(gclk));
	jdff dff_B_2lPoOPl03_0(.din(w_dff_B_okJl0APA3_0),.dout(w_dff_B_2lPoOPl03_0),.clk(gclk));
	jdff dff_B_HaoU4eN69_0(.din(w_dff_B_2lPoOPl03_0),.dout(w_dff_B_HaoU4eN69_0),.clk(gclk));
	jdff dff_B_yj6azYvT2_0(.din(w_dff_B_HaoU4eN69_0),.dout(w_dff_B_yj6azYvT2_0),.clk(gclk));
	jdff dff_B_Eu2rFSWJ1_0(.din(w_dff_B_yj6azYvT2_0),.dout(w_dff_B_Eu2rFSWJ1_0),.clk(gclk));
	jdff dff_B_PFeOYQaX8_0(.din(w_dff_B_Eu2rFSWJ1_0),.dout(w_dff_B_PFeOYQaX8_0),.clk(gclk));
	jdff dff_B_vMvenhfX3_0(.din(w_dff_B_PFeOYQaX8_0),.dout(w_dff_B_vMvenhfX3_0),.clk(gclk));
	jdff dff_B_wZ3FJX3c1_0(.din(w_dff_B_vMvenhfX3_0),.dout(w_dff_B_wZ3FJX3c1_0),.clk(gclk));
	jdff dff_B_jFOUyfxY2_0(.din(w_dff_B_wZ3FJX3c1_0),.dout(w_dff_B_jFOUyfxY2_0),.clk(gclk));
	jdff dff_B_MfeaioIt7_0(.din(w_dff_B_jFOUyfxY2_0),.dout(w_dff_B_MfeaioIt7_0),.clk(gclk));
	jdff dff_B_9kRdCrj86_0(.din(w_dff_B_MfeaioIt7_0),.dout(w_dff_B_9kRdCrj86_0),.clk(gclk));
	jdff dff_B_pwd3PH0a4_0(.din(w_dff_B_9kRdCrj86_0),.dout(w_dff_B_pwd3PH0a4_0),.clk(gclk));
	jdff dff_B_0Jx5mqXQ0_0(.din(w_dff_B_pwd3PH0a4_0),.dout(w_dff_B_0Jx5mqXQ0_0),.clk(gclk));
	jdff dff_B_VUuubfv55_0(.din(w_dff_B_0Jx5mqXQ0_0),.dout(w_dff_B_VUuubfv55_0),.clk(gclk));
	jdff dff_B_KFd18uWV7_0(.din(w_dff_B_VUuubfv55_0),.dout(w_dff_B_KFd18uWV7_0),.clk(gclk));
	jdff dff_B_K8p4uDlq8_0(.din(w_dff_B_KFd18uWV7_0),.dout(w_dff_B_K8p4uDlq8_0),.clk(gclk));
	jdff dff_B_MxdQpzyM1_0(.din(w_dff_B_K8p4uDlq8_0),.dout(w_dff_B_MxdQpzyM1_0),.clk(gclk));
	jdff dff_B_Uxw8tnbp2_0(.din(w_dff_B_MxdQpzyM1_0),.dout(w_dff_B_Uxw8tnbp2_0),.clk(gclk));
	jdff dff_B_J8jYby6L9_0(.din(w_dff_B_Uxw8tnbp2_0),.dout(w_dff_B_J8jYby6L9_0),.clk(gclk));
	jdff dff_B_1hA3Zjco7_0(.din(w_dff_B_J8jYby6L9_0),.dout(w_dff_B_1hA3Zjco7_0),.clk(gclk));
	jdff dff_B_KJK0PAH61_0(.din(w_dff_B_1hA3Zjco7_0),.dout(w_dff_B_KJK0PAH61_0),.clk(gclk));
	jdff dff_B_dJuaSdJh4_0(.din(w_dff_B_KJK0PAH61_0),.dout(w_dff_B_dJuaSdJh4_0),.clk(gclk));
	jdff dff_B_4U8x8mnJ7_0(.din(w_dff_B_dJuaSdJh4_0),.dout(w_dff_B_4U8x8mnJ7_0),.clk(gclk));
	jdff dff_B_WPojmvGb3_0(.din(w_dff_B_4U8x8mnJ7_0),.dout(w_dff_B_WPojmvGb3_0),.clk(gclk));
	jdff dff_B_eX7TXg2U3_0(.din(w_dff_B_WPojmvGb3_0),.dout(w_dff_B_eX7TXg2U3_0),.clk(gclk));
	jdff dff_B_oF2X9Cwx7_0(.din(w_dff_B_eX7TXg2U3_0),.dout(w_dff_B_oF2X9Cwx7_0),.clk(gclk));
	jdff dff_B_Gy3LbCy64_0(.din(w_dff_B_oF2X9Cwx7_0),.dout(w_dff_B_Gy3LbCy64_0),.clk(gclk));
	jdff dff_B_LHTXzUl40_0(.din(w_dff_B_Gy3LbCy64_0),.dout(w_dff_B_LHTXzUl40_0),.clk(gclk));
	jdff dff_B_5PUROoBS0_0(.din(w_dff_B_LHTXzUl40_0),.dout(w_dff_B_5PUROoBS0_0),.clk(gclk));
	jdff dff_B_l7pV1nzR2_0(.din(w_dff_B_5PUROoBS0_0),.dout(w_dff_B_l7pV1nzR2_0),.clk(gclk));
	jdff dff_B_hBR33tVC7_0(.din(w_dff_B_l7pV1nzR2_0),.dout(w_dff_B_hBR33tVC7_0),.clk(gclk));
	jdff dff_B_rxxQYZmA9_0(.din(w_dff_B_hBR33tVC7_0),.dout(w_dff_B_rxxQYZmA9_0),.clk(gclk));
	jdff dff_B_mDYmXbQU0_0(.din(w_dff_B_rxxQYZmA9_0),.dout(w_dff_B_mDYmXbQU0_0),.clk(gclk));
	jdff dff_B_mBpp0bFr9_0(.din(w_dff_B_mDYmXbQU0_0),.dout(w_dff_B_mBpp0bFr9_0),.clk(gclk));
	jdff dff_B_FjTeiGUe2_0(.din(w_dff_B_mBpp0bFr9_0),.dout(w_dff_B_FjTeiGUe2_0),.clk(gclk));
	jdff dff_B_q8d0M6PG0_0(.din(w_dff_B_FjTeiGUe2_0),.dout(w_dff_B_q8d0M6PG0_0),.clk(gclk));
	jdff dff_B_B5gUXouM3_0(.din(w_dff_B_q8d0M6PG0_0),.dout(w_dff_B_B5gUXouM3_0),.clk(gclk));
	jdff dff_B_2yOO5nOM6_0(.din(w_dff_B_B5gUXouM3_0),.dout(w_dff_B_2yOO5nOM6_0),.clk(gclk));
	jdff dff_B_sOUdE9qb5_0(.din(w_dff_B_2yOO5nOM6_0),.dout(w_dff_B_sOUdE9qb5_0),.clk(gclk));
	jdff dff_B_xcePaCNo1_0(.din(w_dff_B_sOUdE9qb5_0),.dout(w_dff_B_xcePaCNo1_0),.clk(gclk));
	jdff dff_B_63vNJJiu5_0(.din(w_dff_B_xcePaCNo1_0),.dout(w_dff_B_63vNJJiu5_0),.clk(gclk));
	jdff dff_B_2PqNYrIe4_0(.din(w_dff_B_63vNJJiu5_0),.dout(w_dff_B_2PqNYrIe4_0),.clk(gclk));
	jdff dff_B_8b1ag7og5_0(.din(w_dff_B_2PqNYrIe4_0),.dout(w_dff_B_8b1ag7og5_0),.clk(gclk));
	jdff dff_B_gdeiR5LT7_0(.din(w_dff_B_8b1ag7og5_0),.dout(w_dff_B_gdeiR5LT7_0),.clk(gclk));
	jdff dff_B_Da09Io531_0(.din(w_dff_B_gdeiR5LT7_0),.dout(w_dff_B_Da09Io531_0),.clk(gclk));
	jdff dff_B_dVmv9vHg3_0(.din(w_dff_B_Da09Io531_0),.dout(w_dff_B_dVmv9vHg3_0),.clk(gclk));
	jdff dff_B_eHQHT7xz2_0(.din(w_dff_B_dVmv9vHg3_0),.dout(w_dff_B_eHQHT7xz2_0),.clk(gclk));
	jdff dff_B_SWLTI55M8_0(.din(w_dff_B_eHQHT7xz2_0),.dout(w_dff_B_SWLTI55M8_0),.clk(gclk));
	jdff dff_B_LYXJn9qz4_0(.din(w_dff_B_SWLTI55M8_0),.dout(w_dff_B_LYXJn9qz4_0),.clk(gclk));
	jdff dff_B_KGVo2PeX0_0(.din(w_dff_B_LYXJn9qz4_0),.dout(w_dff_B_KGVo2PeX0_0),.clk(gclk));
	jdff dff_B_LAXjsAFB4_0(.din(w_dff_B_KGVo2PeX0_0),.dout(w_dff_B_LAXjsAFB4_0),.clk(gclk));
	jdff dff_B_rI9Nzwhg7_0(.din(w_dff_B_LAXjsAFB4_0),.dout(w_dff_B_rI9Nzwhg7_0),.clk(gclk));
	jdff dff_B_ugvjlxaC5_0(.din(w_dff_B_rI9Nzwhg7_0),.dout(w_dff_B_ugvjlxaC5_0),.clk(gclk));
	jdff dff_B_NANNXVAV9_0(.din(w_dff_B_ugvjlxaC5_0),.dout(w_dff_B_NANNXVAV9_0),.clk(gclk));
	jdff dff_B_j73X8DON5_0(.din(w_dff_B_NANNXVAV9_0),.dout(w_dff_B_j73X8DON5_0),.clk(gclk));
	jdff dff_B_nTtcdtcO5_0(.din(w_dff_B_j73X8DON5_0),.dout(w_dff_B_nTtcdtcO5_0),.clk(gclk));
	jdff dff_B_MXzxbtLz1_0(.din(w_dff_B_nTtcdtcO5_0),.dout(w_dff_B_MXzxbtLz1_0),.clk(gclk));
	jdff dff_B_3cPKHPvk6_0(.din(w_dff_B_MXzxbtLz1_0),.dout(w_dff_B_3cPKHPvk6_0),.clk(gclk));
	jdff dff_B_xD0LztTD2_0(.din(w_dff_B_3cPKHPvk6_0),.dout(w_dff_B_xD0LztTD2_0),.clk(gclk));
	jdff dff_B_zkxrkWd16_0(.din(n868),.dout(w_dff_B_zkxrkWd16_0),.clk(gclk));
	jdff dff_B_4dp5WdPe5_0(.din(w_dff_B_zkxrkWd16_0),.dout(w_dff_B_4dp5WdPe5_0),.clk(gclk));
	jdff dff_B_kZo5hkEK7_0(.din(w_dff_B_4dp5WdPe5_0),.dout(w_dff_B_kZo5hkEK7_0),.clk(gclk));
	jdff dff_B_hKeteD9J5_0(.din(w_dff_B_kZo5hkEK7_0),.dout(w_dff_B_hKeteD9J5_0),.clk(gclk));
	jdff dff_B_Qhoj792v0_0(.din(w_dff_B_hKeteD9J5_0),.dout(w_dff_B_Qhoj792v0_0),.clk(gclk));
	jdff dff_B_jzhPpdlh0_0(.din(w_dff_B_Qhoj792v0_0),.dout(w_dff_B_jzhPpdlh0_0),.clk(gclk));
	jdff dff_B_i1rua6Vc3_0(.din(w_dff_B_jzhPpdlh0_0),.dout(w_dff_B_i1rua6Vc3_0),.clk(gclk));
	jdff dff_B_9tkhkb5q0_0(.din(w_dff_B_i1rua6Vc3_0),.dout(w_dff_B_9tkhkb5q0_0),.clk(gclk));
	jdff dff_B_ZJ1rabc32_0(.din(w_dff_B_9tkhkb5q0_0),.dout(w_dff_B_ZJ1rabc32_0),.clk(gclk));
	jdff dff_B_s5I3v4ig9_0(.din(w_dff_B_ZJ1rabc32_0),.dout(w_dff_B_s5I3v4ig9_0),.clk(gclk));
	jdff dff_B_LkQJ95b28_0(.din(w_dff_B_s5I3v4ig9_0),.dout(w_dff_B_LkQJ95b28_0),.clk(gclk));
	jdff dff_B_sQSXIYc20_0(.din(w_dff_B_LkQJ95b28_0),.dout(w_dff_B_sQSXIYc20_0),.clk(gclk));
	jdff dff_B_rkanMmVt0_0(.din(w_dff_B_sQSXIYc20_0),.dout(w_dff_B_rkanMmVt0_0),.clk(gclk));
	jdff dff_B_QGHErctr7_0(.din(w_dff_B_rkanMmVt0_0),.dout(w_dff_B_QGHErctr7_0),.clk(gclk));
	jdff dff_B_PT7i1Ttz8_0(.din(w_dff_B_QGHErctr7_0),.dout(w_dff_B_PT7i1Ttz8_0),.clk(gclk));
	jdff dff_B_dBxtBld69_0(.din(w_dff_B_PT7i1Ttz8_0),.dout(w_dff_B_dBxtBld69_0),.clk(gclk));
	jdff dff_B_r4VKMphT6_0(.din(w_dff_B_dBxtBld69_0),.dout(w_dff_B_r4VKMphT6_0),.clk(gclk));
	jdff dff_B_31MmSSZo3_0(.din(w_dff_B_r4VKMphT6_0),.dout(w_dff_B_31MmSSZo3_0),.clk(gclk));
	jdff dff_B_5uiwG3cc4_0(.din(w_dff_B_31MmSSZo3_0),.dout(w_dff_B_5uiwG3cc4_0),.clk(gclk));
	jdff dff_B_YJlMuXGB9_0(.din(w_dff_B_5uiwG3cc4_0),.dout(w_dff_B_YJlMuXGB9_0),.clk(gclk));
	jdff dff_B_IZ6uK1A32_0(.din(w_dff_B_YJlMuXGB9_0),.dout(w_dff_B_IZ6uK1A32_0),.clk(gclk));
	jdff dff_B_878j9qzM5_0(.din(w_dff_B_IZ6uK1A32_0),.dout(w_dff_B_878j9qzM5_0),.clk(gclk));
	jdff dff_B_BIiO9j742_0(.din(w_dff_B_878j9qzM5_0),.dout(w_dff_B_BIiO9j742_0),.clk(gclk));
	jdff dff_B_Vs9rDLX22_0(.din(w_dff_B_BIiO9j742_0),.dout(w_dff_B_Vs9rDLX22_0),.clk(gclk));
	jdff dff_B_jK6Lh1E11_0(.din(w_dff_B_Vs9rDLX22_0),.dout(w_dff_B_jK6Lh1E11_0),.clk(gclk));
	jdff dff_B_xHhRv1Kb7_0(.din(w_dff_B_jK6Lh1E11_0),.dout(w_dff_B_xHhRv1Kb7_0),.clk(gclk));
	jdff dff_B_Sf1jbtGk8_0(.din(w_dff_B_xHhRv1Kb7_0),.dout(w_dff_B_Sf1jbtGk8_0),.clk(gclk));
	jdff dff_B_UhV715RX2_0(.din(w_dff_B_Sf1jbtGk8_0),.dout(w_dff_B_UhV715RX2_0),.clk(gclk));
	jdff dff_B_5YX6nJMq1_0(.din(w_dff_B_UhV715RX2_0),.dout(w_dff_B_5YX6nJMq1_0),.clk(gclk));
	jdff dff_B_5OX6T6bd1_0(.din(w_dff_B_5YX6nJMq1_0),.dout(w_dff_B_5OX6T6bd1_0),.clk(gclk));
	jdff dff_B_d5wbN7sk9_0(.din(w_dff_B_5OX6T6bd1_0),.dout(w_dff_B_d5wbN7sk9_0),.clk(gclk));
	jdff dff_B_q7YBMCvj4_0(.din(w_dff_B_d5wbN7sk9_0),.dout(w_dff_B_q7YBMCvj4_0),.clk(gclk));
	jdff dff_B_lLGCBk5P2_0(.din(w_dff_B_q7YBMCvj4_0),.dout(w_dff_B_lLGCBk5P2_0),.clk(gclk));
	jdff dff_B_yHIi2Z015_0(.din(w_dff_B_lLGCBk5P2_0),.dout(w_dff_B_yHIi2Z015_0),.clk(gclk));
	jdff dff_B_BbYLq30u9_0(.din(w_dff_B_yHIi2Z015_0),.dout(w_dff_B_BbYLq30u9_0),.clk(gclk));
	jdff dff_B_ySBxrBfl7_0(.din(w_dff_B_BbYLq30u9_0),.dout(w_dff_B_ySBxrBfl7_0),.clk(gclk));
	jdff dff_B_9gUZrYLs3_0(.din(w_dff_B_ySBxrBfl7_0),.dout(w_dff_B_9gUZrYLs3_0),.clk(gclk));
	jdff dff_B_mHreAn3l5_0(.din(w_dff_B_9gUZrYLs3_0),.dout(w_dff_B_mHreAn3l5_0),.clk(gclk));
	jdff dff_B_9LvwDiqm0_0(.din(w_dff_B_mHreAn3l5_0),.dout(w_dff_B_9LvwDiqm0_0),.clk(gclk));
	jdff dff_B_pb9bVdYe1_0(.din(w_dff_B_9LvwDiqm0_0),.dout(w_dff_B_pb9bVdYe1_0),.clk(gclk));
	jdff dff_B_LzJaCswK7_0(.din(w_dff_B_pb9bVdYe1_0),.dout(w_dff_B_LzJaCswK7_0),.clk(gclk));
	jdff dff_B_GVilGTTs0_0(.din(w_dff_B_LzJaCswK7_0),.dout(w_dff_B_GVilGTTs0_0),.clk(gclk));
	jdff dff_B_qTM2WJ6g7_0(.din(w_dff_B_GVilGTTs0_0),.dout(w_dff_B_qTM2WJ6g7_0),.clk(gclk));
	jdff dff_B_18PBxVR25_0(.din(w_dff_B_qTM2WJ6g7_0),.dout(w_dff_B_18PBxVR25_0),.clk(gclk));
	jdff dff_B_HbKJ7URU3_0(.din(w_dff_B_18PBxVR25_0),.dout(w_dff_B_HbKJ7URU3_0),.clk(gclk));
	jdff dff_B_IEfb7JRR2_0(.din(w_dff_B_HbKJ7URU3_0),.dout(w_dff_B_IEfb7JRR2_0),.clk(gclk));
	jdff dff_B_h6f9s4XF0_0(.din(w_dff_B_IEfb7JRR2_0),.dout(w_dff_B_h6f9s4XF0_0),.clk(gclk));
	jdff dff_B_QYHw80FP7_0(.din(w_dff_B_h6f9s4XF0_0),.dout(w_dff_B_QYHw80FP7_0),.clk(gclk));
	jdff dff_B_8Mtd3Naa9_0(.din(w_dff_B_QYHw80FP7_0),.dout(w_dff_B_8Mtd3Naa9_0),.clk(gclk));
	jdff dff_B_JFTcRt9D8_0(.din(w_dff_B_8Mtd3Naa9_0),.dout(w_dff_B_JFTcRt9D8_0),.clk(gclk));
	jdff dff_B_wscGVvbY9_0(.din(w_dff_B_JFTcRt9D8_0),.dout(w_dff_B_wscGVvbY9_0),.clk(gclk));
	jdff dff_B_mGCbnmdl5_0(.din(w_dff_B_wscGVvbY9_0),.dout(w_dff_B_mGCbnmdl5_0),.clk(gclk));
	jdff dff_B_sQV7d8l79_0(.din(w_dff_B_mGCbnmdl5_0),.dout(w_dff_B_sQV7d8l79_0),.clk(gclk));
	jdff dff_B_apYOr9S20_0(.din(w_dff_B_sQV7d8l79_0),.dout(w_dff_B_apYOr9S20_0),.clk(gclk));
	jdff dff_B_qnnpzRAH0_0(.din(w_dff_B_apYOr9S20_0),.dout(w_dff_B_qnnpzRAH0_0),.clk(gclk));
	jdff dff_B_U0pY4BZE9_0(.din(w_dff_B_qnnpzRAH0_0),.dout(w_dff_B_U0pY4BZE9_0),.clk(gclk));
	jdff dff_B_BHea5s6y5_0(.din(w_dff_B_U0pY4BZE9_0),.dout(w_dff_B_BHea5s6y5_0),.clk(gclk));
	jdff dff_B_tsVuorQg7_0(.din(w_dff_B_BHea5s6y5_0),.dout(w_dff_B_tsVuorQg7_0),.clk(gclk));
	jdff dff_B_3K9S219l0_0(.din(w_dff_B_tsVuorQg7_0),.dout(w_dff_B_3K9S219l0_0),.clk(gclk));
	jdff dff_B_toQCYd3N5_0(.din(w_dff_B_3K9S219l0_0),.dout(w_dff_B_toQCYd3N5_0),.clk(gclk));
	jdff dff_B_tHZmABeR8_0(.din(w_dff_B_toQCYd3N5_0),.dout(w_dff_B_tHZmABeR8_0),.clk(gclk));
	jdff dff_B_YGTEzjhz4_0(.din(w_dff_B_tHZmABeR8_0),.dout(w_dff_B_YGTEzjhz4_0),.clk(gclk));
	jdff dff_B_CLYSVPik4_0(.din(w_dff_B_YGTEzjhz4_0),.dout(w_dff_B_CLYSVPik4_0),.clk(gclk));
	jdff dff_B_DlDxpIud7_0(.din(w_dff_B_CLYSVPik4_0),.dout(w_dff_B_DlDxpIud7_0),.clk(gclk));
	jdff dff_B_wYSkosGg7_0(.din(w_dff_B_DlDxpIud7_0),.dout(w_dff_B_wYSkosGg7_0),.clk(gclk));
	jdff dff_B_jirmYym30_0(.din(w_dff_B_wYSkosGg7_0),.dout(w_dff_B_jirmYym30_0),.clk(gclk));
	jdff dff_B_w7WuqIQE6_0(.din(w_dff_B_jirmYym30_0),.dout(w_dff_B_w7WuqIQE6_0),.clk(gclk));
	jdff dff_B_ZI38D2bb7_0(.din(w_dff_B_w7WuqIQE6_0),.dout(w_dff_B_ZI38D2bb7_0),.clk(gclk));
	jdff dff_B_MTN3bQAP2_0(.din(w_dff_B_ZI38D2bb7_0),.dout(w_dff_B_MTN3bQAP2_0),.clk(gclk));
	jdff dff_B_W9tLR0IX1_0(.din(w_dff_B_MTN3bQAP2_0),.dout(w_dff_B_W9tLR0IX1_0),.clk(gclk));
	jdff dff_B_iTYTaTfQ0_0(.din(w_dff_B_W9tLR0IX1_0),.dout(w_dff_B_iTYTaTfQ0_0),.clk(gclk));
	jdff dff_B_kvU20JZV5_0(.din(w_dff_B_iTYTaTfQ0_0),.dout(w_dff_B_kvU20JZV5_0),.clk(gclk));
	jdff dff_B_E60WvHlZ6_0(.din(w_dff_B_kvU20JZV5_0),.dout(w_dff_B_E60WvHlZ6_0),.clk(gclk));
	jdff dff_B_KlI0Ouxa1_0(.din(w_dff_B_E60WvHlZ6_0),.dout(w_dff_B_KlI0Ouxa1_0),.clk(gclk));
	jdff dff_B_thqkTFDY1_0(.din(w_dff_B_KlI0Ouxa1_0),.dout(w_dff_B_thqkTFDY1_0),.clk(gclk));
	jdff dff_B_EGAh7bB19_0(.din(w_dff_B_thqkTFDY1_0),.dout(w_dff_B_EGAh7bB19_0),.clk(gclk));
	jdff dff_B_blrktEUo2_0(.din(w_dff_B_EGAh7bB19_0),.dout(w_dff_B_blrktEUo2_0),.clk(gclk));
	jdff dff_B_DYUpT7FU2_0(.din(w_dff_B_blrktEUo2_0),.dout(w_dff_B_DYUpT7FU2_0),.clk(gclk));
	jdff dff_B_pJOCtfPc7_0(.din(w_dff_B_DYUpT7FU2_0),.dout(w_dff_B_pJOCtfPc7_0),.clk(gclk));
	jdff dff_B_kZscPfF05_0(.din(w_dff_B_pJOCtfPc7_0),.dout(w_dff_B_kZscPfF05_0),.clk(gclk));
	jdff dff_B_QcZZTuIQ3_0(.din(n874),.dout(w_dff_B_QcZZTuIQ3_0),.clk(gclk));
	jdff dff_B_4Ib2ppjx9_0(.din(w_dff_B_QcZZTuIQ3_0),.dout(w_dff_B_4Ib2ppjx9_0),.clk(gclk));
	jdff dff_B_V3gwhS3V5_0(.din(w_dff_B_4Ib2ppjx9_0),.dout(w_dff_B_V3gwhS3V5_0),.clk(gclk));
	jdff dff_B_IYFP5TKO1_0(.din(w_dff_B_V3gwhS3V5_0),.dout(w_dff_B_IYFP5TKO1_0),.clk(gclk));
	jdff dff_B_X7wuqdgo1_0(.din(w_dff_B_IYFP5TKO1_0),.dout(w_dff_B_X7wuqdgo1_0),.clk(gclk));
	jdff dff_B_VnuZ65KF6_0(.din(w_dff_B_X7wuqdgo1_0),.dout(w_dff_B_VnuZ65KF6_0),.clk(gclk));
	jdff dff_B_UdcxoF2j6_0(.din(w_dff_B_VnuZ65KF6_0),.dout(w_dff_B_UdcxoF2j6_0),.clk(gclk));
	jdff dff_B_fAYQjJsa9_0(.din(w_dff_B_UdcxoF2j6_0),.dout(w_dff_B_fAYQjJsa9_0),.clk(gclk));
	jdff dff_B_CA2U5DbZ0_0(.din(w_dff_B_fAYQjJsa9_0),.dout(w_dff_B_CA2U5DbZ0_0),.clk(gclk));
	jdff dff_B_aEgfGQY88_0(.din(w_dff_B_CA2U5DbZ0_0),.dout(w_dff_B_aEgfGQY88_0),.clk(gclk));
	jdff dff_B_8cCJzAnO8_0(.din(w_dff_B_aEgfGQY88_0),.dout(w_dff_B_8cCJzAnO8_0),.clk(gclk));
	jdff dff_B_n5UIEOHW0_0(.din(w_dff_B_8cCJzAnO8_0),.dout(w_dff_B_n5UIEOHW0_0),.clk(gclk));
	jdff dff_B_yA4ojZ635_0(.din(w_dff_B_n5UIEOHW0_0),.dout(w_dff_B_yA4ojZ635_0),.clk(gclk));
	jdff dff_B_fo0qJLoY3_0(.din(w_dff_B_yA4ojZ635_0),.dout(w_dff_B_fo0qJLoY3_0),.clk(gclk));
	jdff dff_B_BQtJWMuP1_0(.din(w_dff_B_fo0qJLoY3_0),.dout(w_dff_B_BQtJWMuP1_0),.clk(gclk));
	jdff dff_B_wdKNfiWz1_0(.din(w_dff_B_BQtJWMuP1_0),.dout(w_dff_B_wdKNfiWz1_0),.clk(gclk));
	jdff dff_B_mmNYz6hq6_0(.din(w_dff_B_wdKNfiWz1_0),.dout(w_dff_B_mmNYz6hq6_0),.clk(gclk));
	jdff dff_B_B7YPRWT83_0(.din(w_dff_B_mmNYz6hq6_0),.dout(w_dff_B_B7YPRWT83_0),.clk(gclk));
	jdff dff_B_HQlYCfa04_0(.din(w_dff_B_B7YPRWT83_0),.dout(w_dff_B_HQlYCfa04_0),.clk(gclk));
	jdff dff_B_ZjO0DUm18_0(.din(w_dff_B_HQlYCfa04_0),.dout(w_dff_B_ZjO0DUm18_0),.clk(gclk));
	jdff dff_B_xGL6q3Bd5_0(.din(w_dff_B_ZjO0DUm18_0),.dout(w_dff_B_xGL6q3Bd5_0),.clk(gclk));
	jdff dff_B_GFMVAOmn4_0(.din(w_dff_B_xGL6q3Bd5_0),.dout(w_dff_B_GFMVAOmn4_0),.clk(gclk));
	jdff dff_B_WN0PGnhN3_0(.din(w_dff_B_GFMVAOmn4_0),.dout(w_dff_B_WN0PGnhN3_0),.clk(gclk));
	jdff dff_B_Fe2F91ED4_0(.din(w_dff_B_WN0PGnhN3_0),.dout(w_dff_B_Fe2F91ED4_0),.clk(gclk));
	jdff dff_B_rOptkkxL5_0(.din(w_dff_B_Fe2F91ED4_0),.dout(w_dff_B_rOptkkxL5_0),.clk(gclk));
	jdff dff_B_Aom7jxAB4_0(.din(w_dff_B_rOptkkxL5_0),.dout(w_dff_B_Aom7jxAB4_0),.clk(gclk));
	jdff dff_B_FAEDgE524_0(.din(w_dff_B_Aom7jxAB4_0),.dout(w_dff_B_FAEDgE524_0),.clk(gclk));
	jdff dff_B_VyYYL8Qt5_0(.din(w_dff_B_FAEDgE524_0),.dout(w_dff_B_VyYYL8Qt5_0),.clk(gclk));
	jdff dff_B_YlYKYX4Q4_0(.din(w_dff_B_VyYYL8Qt5_0),.dout(w_dff_B_YlYKYX4Q4_0),.clk(gclk));
	jdff dff_B_gSPGKa2r4_0(.din(w_dff_B_YlYKYX4Q4_0),.dout(w_dff_B_gSPGKa2r4_0),.clk(gclk));
	jdff dff_B_p6f5tlaT1_0(.din(w_dff_B_gSPGKa2r4_0),.dout(w_dff_B_p6f5tlaT1_0),.clk(gclk));
	jdff dff_B_vC3vzaYd9_0(.din(w_dff_B_p6f5tlaT1_0),.dout(w_dff_B_vC3vzaYd9_0),.clk(gclk));
	jdff dff_B_X1RoAtF93_0(.din(w_dff_B_vC3vzaYd9_0),.dout(w_dff_B_X1RoAtF93_0),.clk(gclk));
	jdff dff_B_vhYTa54k4_0(.din(w_dff_B_X1RoAtF93_0),.dout(w_dff_B_vhYTa54k4_0),.clk(gclk));
	jdff dff_B_Ak161OG79_0(.din(w_dff_B_vhYTa54k4_0),.dout(w_dff_B_Ak161OG79_0),.clk(gclk));
	jdff dff_B_DrnpvY3C8_0(.din(w_dff_B_Ak161OG79_0),.dout(w_dff_B_DrnpvY3C8_0),.clk(gclk));
	jdff dff_B_QrDIbC9f0_0(.din(w_dff_B_DrnpvY3C8_0),.dout(w_dff_B_QrDIbC9f0_0),.clk(gclk));
	jdff dff_B_3Bo961OP5_0(.din(w_dff_B_QrDIbC9f0_0),.dout(w_dff_B_3Bo961OP5_0),.clk(gclk));
	jdff dff_B_IshJWfsA0_0(.din(w_dff_B_3Bo961OP5_0),.dout(w_dff_B_IshJWfsA0_0),.clk(gclk));
	jdff dff_B_E3GkM9bh2_0(.din(w_dff_B_IshJWfsA0_0),.dout(w_dff_B_E3GkM9bh2_0),.clk(gclk));
	jdff dff_B_AbrcW48E5_0(.din(w_dff_B_E3GkM9bh2_0),.dout(w_dff_B_AbrcW48E5_0),.clk(gclk));
	jdff dff_B_BiVauN6W1_0(.din(w_dff_B_AbrcW48E5_0),.dout(w_dff_B_BiVauN6W1_0),.clk(gclk));
	jdff dff_B_Y8Oh2AcU8_0(.din(w_dff_B_BiVauN6W1_0),.dout(w_dff_B_Y8Oh2AcU8_0),.clk(gclk));
	jdff dff_B_TFZwZyeR2_0(.din(w_dff_B_Y8Oh2AcU8_0),.dout(w_dff_B_TFZwZyeR2_0),.clk(gclk));
	jdff dff_B_ZiNsTG490_0(.din(w_dff_B_TFZwZyeR2_0),.dout(w_dff_B_ZiNsTG490_0),.clk(gclk));
	jdff dff_B_bz2HqiGf4_0(.din(w_dff_B_ZiNsTG490_0),.dout(w_dff_B_bz2HqiGf4_0),.clk(gclk));
	jdff dff_B_1XjZcdtT3_0(.din(w_dff_B_bz2HqiGf4_0),.dout(w_dff_B_1XjZcdtT3_0),.clk(gclk));
	jdff dff_B_VmNzdaB18_0(.din(w_dff_B_1XjZcdtT3_0),.dout(w_dff_B_VmNzdaB18_0),.clk(gclk));
	jdff dff_B_O8iW6WIQ4_0(.din(w_dff_B_VmNzdaB18_0),.dout(w_dff_B_O8iW6WIQ4_0),.clk(gclk));
	jdff dff_B_dnKQIDC61_0(.din(w_dff_B_O8iW6WIQ4_0),.dout(w_dff_B_dnKQIDC61_0),.clk(gclk));
	jdff dff_B_N5uL4RCF3_0(.din(w_dff_B_dnKQIDC61_0),.dout(w_dff_B_N5uL4RCF3_0),.clk(gclk));
	jdff dff_B_gccVeE6L6_0(.din(w_dff_B_N5uL4RCF3_0),.dout(w_dff_B_gccVeE6L6_0),.clk(gclk));
	jdff dff_B_c6euSobx0_0(.din(w_dff_B_gccVeE6L6_0),.dout(w_dff_B_c6euSobx0_0),.clk(gclk));
	jdff dff_B_bZIcHaS78_0(.din(w_dff_B_c6euSobx0_0),.dout(w_dff_B_bZIcHaS78_0),.clk(gclk));
	jdff dff_B_vHG4tcom6_0(.din(w_dff_B_bZIcHaS78_0),.dout(w_dff_B_vHG4tcom6_0),.clk(gclk));
	jdff dff_B_jmbnj2jO3_0(.din(w_dff_B_vHG4tcom6_0),.dout(w_dff_B_jmbnj2jO3_0),.clk(gclk));
	jdff dff_B_6hZiz89g1_0(.din(w_dff_B_jmbnj2jO3_0),.dout(w_dff_B_6hZiz89g1_0),.clk(gclk));
	jdff dff_B_hemcgMxm7_0(.din(w_dff_B_6hZiz89g1_0),.dout(w_dff_B_hemcgMxm7_0),.clk(gclk));
	jdff dff_B_A09Z9Qnf5_0(.din(w_dff_B_hemcgMxm7_0),.dout(w_dff_B_A09Z9Qnf5_0),.clk(gclk));
	jdff dff_B_POhBay9D2_0(.din(w_dff_B_A09Z9Qnf5_0),.dout(w_dff_B_POhBay9D2_0),.clk(gclk));
	jdff dff_B_Ixb1pRGX6_0(.din(w_dff_B_POhBay9D2_0),.dout(w_dff_B_Ixb1pRGX6_0),.clk(gclk));
	jdff dff_B_wdvdLn5n6_0(.din(w_dff_B_Ixb1pRGX6_0),.dout(w_dff_B_wdvdLn5n6_0),.clk(gclk));
	jdff dff_B_TDogG1D40_0(.din(w_dff_B_wdvdLn5n6_0),.dout(w_dff_B_TDogG1D40_0),.clk(gclk));
	jdff dff_B_1owVF1lH7_0(.din(w_dff_B_TDogG1D40_0),.dout(w_dff_B_1owVF1lH7_0),.clk(gclk));
	jdff dff_B_ha0SSQzY4_0(.din(w_dff_B_1owVF1lH7_0),.dout(w_dff_B_ha0SSQzY4_0),.clk(gclk));
	jdff dff_B_2tyf0Uhe8_0(.din(w_dff_B_ha0SSQzY4_0),.dout(w_dff_B_2tyf0Uhe8_0),.clk(gclk));
	jdff dff_B_yzEFVarW7_0(.din(w_dff_B_2tyf0Uhe8_0),.dout(w_dff_B_yzEFVarW7_0),.clk(gclk));
	jdff dff_B_hNYMxaaS9_0(.din(w_dff_B_yzEFVarW7_0),.dout(w_dff_B_hNYMxaaS9_0),.clk(gclk));
	jdff dff_B_dFPTtBWq1_0(.din(w_dff_B_hNYMxaaS9_0),.dout(w_dff_B_dFPTtBWq1_0),.clk(gclk));
	jdff dff_B_cxlppIV79_0(.din(w_dff_B_dFPTtBWq1_0),.dout(w_dff_B_cxlppIV79_0),.clk(gclk));
	jdff dff_B_YVnsYMzi1_0(.din(w_dff_B_cxlppIV79_0),.dout(w_dff_B_YVnsYMzi1_0),.clk(gclk));
	jdff dff_B_HRdAuiEo4_0(.din(w_dff_B_YVnsYMzi1_0),.dout(w_dff_B_HRdAuiEo4_0),.clk(gclk));
	jdff dff_B_dVvbJW963_0(.din(w_dff_B_HRdAuiEo4_0),.dout(w_dff_B_dVvbJW963_0),.clk(gclk));
	jdff dff_B_FCutw8t22_0(.din(w_dff_B_dVvbJW963_0),.dout(w_dff_B_FCutw8t22_0),.clk(gclk));
	jdff dff_B_QClhmHSt5_0(.din(w_dff_B_FCutw8t22_0),.dout(w_dff_B_QClhmHSt5_0),.clk(gclk));
	jdff dff_B_zRyHnnjd2_0(.din(w_dff_B_QClhmHSt5_0),.dout(w_dff_B_zRyHnnjd2_0),.clk(gclk));
	jdff dff_B_kMl9yicX5_0(.din(w_dff_B_zRyHnnjd2_0),.dout(w_dff_B_kMl9yicX5_0),.clk(gclk));
	jdff dff_B_VyIGJ9183_0(.din(w_dff_B_kMl9yicX5_0),.dout(w_dff_B_VyIGJ9183_0),.clk(gclk));
	jdff dff_B_3OfqcGYA6_0(.din(w_dff_B_VyIGJ9183_0),.dout(w_dff_B_3OfqcGYA6_0),.clk(gclk));
	jdff dff_B_SxCzBEj88_0(.din(w_dff_B_3OfqcGYA6_0),.dout(w_dff_B_SxCzBEj88_0),.clk(gclk));
	jdff dff_B_pbwwiBwO7_0(.din(w_dff_B_SxCzBEj88_0),.dout(w_dff_B_pbwwiBwO7_0),.clk(gclk));
	jdff dff_B_agrR3ZMU5_0(.din(n880),.dout(w_dff_B_agrR3ZMU5_0),.clk(gclk));
	jdff dff_B_lw8QH2W58_0(.din(w_dff_B_agrR3ZMU5_0),.dout(w_dff_B_lw8QH2W58_0),.clk(gclk));
	jdff dff_B_Mnw9cP8y6_0(.din(w_dff_B_lw8QH2W58_0),.dout(w_dff_B_Mnw9cP8y6_0),.clk(gclk));
	jdff dff_B_Cnw9lZYv5_0(.din(w_dff_B_Mnw9cP8y6_0),.dout(w_dff_B_Cnw9lZYv5_0),.clk(gclk));
	jdff dff_B_ptAe97e99_0(.din(w_dff_B_Cnw9lZYv5_0),.dout(w_dff_B_ptAe97e99_0),.clk(gclk));
	jdff dff_B_A0K3CV4S3_0(.din(w_dff_B_ptAe97e99_0),.dout(w_dff_B_A0K3CV4S3_0),.clk(gclk));
	jdff dff_B_mILDGCpi8_0(.din(w_dff_B_A0K3CV4S3_0),.dout(w_dff_B_mILDGCpi8_0),.clk(gclk));
	jdff dff_B_3SwRcVo26_0(.din(w_dff_B_mILDGCpi8_0),.dout(w_dff_B_3SwRcVo26_0),.clk(gclk));
	jdff dff_B_3ImerPUB9_0(.din(w_dff_B_3SwRcVo26_0),.dout(w_dff_B_3ImerPUB9_0),.clk(gclk));
	jdff dff_B_iu3g6XT02_0(.din(w_dff_B_3ImerPUB9_0),.dout(w_dff_B_iu3g6XT02_0),.clk(gclk));
	jdff dff_B_tvgBNtyF3_0(.din(w_dff_B_iu3g6XT02_0),.dout(w_dff_B_tvgBNtyF3_0),.clk(gclk));
	jdff dff_B_DrFDeCqs3_0(.din(w_dff_B_tvgBNtyF3_0),.dout(w_dff_B_DrFDeCqs3_0),.clk(gclk));
	jdff dff_B_Z7mhA6AK0_0(.din(w_dff_B_DrFDeCqs3_0),.dout(w_dff_B_Z7mhA6AK0_0),.clk(gclk));
	jdff dff_B_a4r6e87p8_0(.din(w_dff_B_Z7mhA6AK0_0),.dout(w_dff_B_a4r6e87p8_0),.clk(gclk));
	jdff dff_B_DC1xpvVx2_0(.din(w_dff_B_a4r6e87p8_0),.dout(w_dff_B_DC1xpvVx2_0),.clk(gclk));
	jdff dff_B_JqBnzML99_0(.din(w_dff_B_DC1xpvVx2_0),.dout(w_dff_B_JqBnzML99_0),.clk(gclk));
	jdff dff_B_N6Dlo1VF8_0(.din(w_dff_B_JqBnzML99_0),.dout(w_dff_B_N6Dlo1VF8_0),.clk(gclk));
	jdff dff_B_ZNuhTeA95_0(.din(w_dff_B_N6Dlo1VF8_0),.dout(w_dff_B_ZNuhTeA95_0),.clk(gclk));
	jdff dff_B_OcH0zM7x5_0(.din(w_dff_B_ZNuhTeA95_0),.dout(w_dff_B_OcH0zM7x5_0),.clk(gclk));
	jdff dff_B_56CMJVCQ0_0(.din(w_dff_B_OcH0zM7x5_0),.dout(w_dff_B_56CMJVCQ0_0),.clk(gclk));
	jdff dff_B_WsCZY6uQ7_0(.din(w_dff_B_56CMJVCQ0_0),.dout(w_dff_B_WsCZY6uQ7_0),.clk(gclk));
	jdff dff_B_rZgtu4FG9_0(.din(w_dff_B_WsCZY6uQ7_0),.dout(w_dff_B_rZgtu4FG9_0),.clk(gclk));
	jdff dff_B_HpNBxB2c7_0(.din(w_dff_B_rZgtu4FG9_0),.dout(w_dff_B_HpNBxB2c7_0),.clk(gclk));
	jdff dff_B_gEWsEq7B9_0(.din(w_dff_B_HpNBxB2c7_0),.dout(w_dff_B_gEWsEq7B9_0),.clk(gclk));
	jdff dff_B_fUB77CFx7_0(.din(w_dff_B_gEWsEq7B9_0),.dout(w_dff_B_fUB77CFx7_0),.clk(gclk));
	jdff dff_B_xlEFsqaD2_0(.din(w_dff_B_fUB77CFx7_0),.dout(w_dff_B_xlEFsqaD2_0),.clk(gclk));
	jdff dff_B_3TpX3y4U1_0(.din(w_dff_B_xlEFsqaD2_0),.dout(w_dff_B_3TpX3y4U1_0),.clk(gclk));
	jdff dff_B_Mh8Lk0sf7_0(.din(w_dff_B_3TpX3y4U1_0),.dout(w_dff_B_Mh8Lk0sf7_0),.clk(gclk));
	jdff dff_B_nINtHQCR5_0(.din(w_dff_B_Mh8Lk0sf7_0),.dout(w_dff_B_nINtHQCR5_0),.clk(gclk));
	jdff dff_B_8RSEU8P33_0(.din(w_dff_B_nINtHQCR5_0),.dout(w_dff_B_8RSEU8P33_0),.clk(gclk));
	jdff dff_B_lmmmKN3Y3_0(.din(w_dff_B_8RSEU8P33_0),.dout(w_dff_B_lmmmKN3Y3_0),.clk(gclk));
	jdff dff_B_8rswPLN26_0(.din(w_dff_B_lmmmKN3Y3_0),.dout(w_dff_B_8rswPLN26_0),.clk(gclk));
	jdff dff_B_C0bAdgVI9_0(.din(w_dff_B_8rswPLN26_0),.dout(w_dff_B_C0bAdgVI9_0),.clk(gclk));
	jdff dff_B_rVKRJUWc9_0(.din(w_dff_B_C0bAdgVI9_0),.dout(w_dff_B_rVKRJUWc9_0),.clk(gclk));
	jdff dff_B_YRYNKleJ7_0(.din(w_dff_B_rVKRJUWc9_0),.dout(w_dff_B_YRYNKleJ7_0),.clk(gclk));
	jdff dff_B_fOXKvkXw7_0(.din(w_dff_B_YRYNKleJ7_0),.dout(w_dff_B_fOXKvkXw7_0),.clk(gclk));
	jdff dff_B_sUKwU3dg7_0(.din(w_dff_B_fOXKvkXw7_0),.dout(w_dff_B_sUKwU3dg7_0),.clk(gclk));
	jdff dff_B_HePElIVO0_0(.din(w_dff_B_sUKwU3dg7_0),.dout(w_dff_B_HePElIVO0_0),.clk(gclk));
	jdff dff_B_PFUUA1jQ0_0(.din(w_dff_B_HePElIVO0_0),.dout(w_dff_B_PFUUA1jQ0_0),.clk(gclk));
	jdff dff_B_NMYaTAso6_0(.din(w_dff_B_PFUUA1jQ0_0),.dout(w_dff_B_NMYaTAso6_0),.clk(gclk));
	jdff dff_B_n4a4ziBb1_0(.din(w_dff_B_NMYaTAso6_0),.dout(w_dff_B_n4a4ziBb1_0),.clk(gclk));
	jdff dff_B_IwOBWZwc1_0(.din(w_dff_B_n4a4ziBb1_0),.dout(w_dff_B_IwOBWZwc1_0),.clk(gclk));
	jdff dff_B_lCjMimkk7_0(.din(w_dff_B_IwOBWZwc1_0),.dout(w_dff_B_lCjMimkk7_0),.clk(gclk));
	jdff dff_B_6ns0qHdv5_0(.din(w_dff_B_lCjMimkk7_0),.dout(w_dff_B_6ns0qHdv5_0),.clk(gclk));
	jdff dff_B_D1bVyfCg7_0(.din(w_dff_B_6ns0qHdv5_0),.dout(w_dff_B_D1bVyfCg7_0),.clk(gclk));
	jdff dff_B_2dn2Sa3d9_0(.din(w_dff_B_D1bVyfCg7_0),.dout(w_dff_B_2dn2Sa3d9_0),.clk(gclk));
	jdff dff_B_P68jduJO0_0(.din(w_dff_B_2dn2Sa3d9_0),.dout(w_dff_B_P68jduJO0_0),.clk(gclk));
	jdff dff_B_6IjaQztm7_0(.din(w_dff_B_P68jduJO0_0),.dout(w_dff_B_6IjaQztm7_0),.clk(gclk));
	jdff dff_B_K1LDRKNf6_0(.din(w_dff_B_6IjaQztm7_0),.dout(w_dff_B_K1LDRKNf6_0),.clk(gclk));
	jdff dff_B_GFKdPcj02_0(.din(w_dff_B_K1LDRKNf6_0),.dout(w_dff_B_GFKdPcj02_0),.clk(gclk));
	jdff dff_B_nKk7wij81_0(.din(w_dff_B_GFKdPcj02_0),.dout(w_dff_B_nKk7wij81_0),.clk(gclk));
	jdff dff_B_MalIJpMY9_0(.din(w_dff_B_nKk7wij81_0),.dout(w_dff_B_MalIJpMY9_0),.clk(gclk));
	jdff dff_B_FVkGPY8A4_0(.din(w_dff_B_MalIJpMY9_0),.dout(w_dff_B_FVkGPY8A4_0),.clk(gclk));
	jdff dff_B_v3TbuZbB4_0(.din(w_dff_B_FVkGPY8A4_0),.dout(w_dff_B_v3TbuZbB4_0),.clk(gclk));
	jdff dff_B_ltmXst6H8_0(.din(w_dff_B_v3TbuZbB4_0),.dout(w_dff_B_ltmXst6H8_0),.clk(gclk));
	jdff dff_B_OV2vOiv01_0(.din(w_dff_B_ltmXst6H8_0),.dout(w_dff_B_OV2vOiv01_0),.clk(gclk));
	jdff dff_B_x9YPzonl1_0(.din(w_dff_B_OV2vOiv01_0),.dout(w_dff_B_x9YPzonl1_0),.clk(gclk));
	jdff dff_B_ROVXGLfr9_0(.din(w_dff_B_x9YPzonl1_0),.dout(w_dff_B_ROVXGLfr9_0),.clk(gclk));
	jdff dff_B_VNtrsrO71_0(.din(w_dff_B_ROVXGLfr9_0),.dout(w_dff_B_VNtrsrO71_0),.clk(gclk));
	jdff dff_B_BXxgX8dt2_0(.din(w_dff_B_VNtrsrO71_0),.dout(w_dff_B_BXxgX8dt2_0),.clk(gclk));
	jdff dff_B_u7Hu8Xtq8_0(.din(w_dff_B_BXxgX8dt2_0),.dout(w_dff_B_u7Hu8Xtq8_0),.clk(gclk));
	jdff dff_B_scYSoCvN2_0(.din(w_dff_B_u7Hu8Xtq8_0),.dout(w_dff_B_scYSoCvN2_0),.clk(gclk));
	jdff dff_B_Rx2TCi7i0_0(.din(w_dff_B_scYSoCvN2_0),.dout(w_dff_B_Rx2TCi7i0_0),.clk(gclk));
	jdff dff_B_YWeOlb322_0(.din(w_dff_B_Rx2TCi7i0_0),.dout(w_dff_B_YWeOlb322_0),.clk(gclk));
	jdff dff_B_m1nicARd3_0(.din(w_dff_B_YWeOlb322_0),.dout(w_dff_B_m1nicARd3_0),.clk(gclk));
	jdff dff_B_K3vHac6Q0_0(.din(w_dff_B_m1nicARd3_0),.dout(w_dff_B_K3vHac6Q0_0),.clk(gclk));
	jdff dff_B_bpZWisHi2_0(.din(w_dff_B_K3vHac6Q0_0),.dout(w_dff_B_bpZWisHi2_0),.clk(gclk));
	jdff dff_B_2WAT7UkG4_0(.din(w_dff_B_bpZWisHi2_0),.dout(w_dff_B_2WAT7UkG4_0),.clk(gclk));
	jdff dff_B_AtxdfFTw1_0(.din(w_dff_B_2WAT7UkG4_0),.dout(w_dff_B_AtxdfFTw1_0),.clk(gclk));
	jdff dff_B_WJdnsCAZ5_0(.din(w_dff_B_AtxdfFTw1_0),.dout(w_dff_B_WJdnsCAZ5_0),.clk(gclk));
	jdff dff_B_pbHjgkNb1_0(.din(w_dff_B_WJdnsCAZ5_0),.dout(w_dff_B_pbHjgkNb1_0),.clk(gclk));
	jdff dff_B_jzXi2paf6_0(.din(w_dff_B_pbHjgkNb1_0),.dout(w_dff_B_jzXi2paf6_0),.clk(gclk));
	jdff dff_B_iEMhaJPs0_0(.din(w_dff_B_jzXi2paf6_0),.dout(w_dff_B_iEMhaJPs0_0),.clk(gclk));
	jdff dff_B_xri6LWbP8_0(.din(w_dff_B_iEMhaJPs0_0),.dout(w_dff_B_xri6LWbP8_0),.clk(gclk));
	jdff dff_B_Zi36Nuu53_0(.din(w_dff_B_xri6LWbP8_0),.dout(w_dff_B_Zi36Nuu53_0),.clk(gclk));
	jdff dff_B_kP1VHHiD0_0(.din(w_dff_B_Zi36Nuu53_0),.dout(w_dff_B_kP1VHHiD0_0),.clk(gclk));
	jdff dff_B_r4NWKp934_0(.din(w_dff_B_kP1VHHiD0_0),.dout(w_dff_B_r4NWKp934_0),.clk(gclk));
	jdff dff_B_cfr2EdJo8_0(.din(w_dff_B_r4NWKp934_0),.dout(w_dff_B_cfr2EdJo8_0),.clk(gclk));
	jdff dff_B_WXj5shUv8_0(.din(w_dff_B_cfr2EdJo8_0),.dout(w_dff_B_WXj5shUv8_0),.clk(gclk));
	jdff dff_B_fHL9ewFY8_0(.din(w_dff_B_WXj5shUv8_0),.dout(w_dff_B_fHL9ewFY8_0),.clk(gclk));
	jdff dff_B_pC36Z5Il9_0(.din(w_dff_B_fHL9ewFY8_0),.dout(w_dff_B_pC36Z5Il9_0),.clk(gclk));
	jdff dff_B_bMIFxpYM3_0(.din(w_dff_B_pC36Z5Il9_0),.dout(w_dff_B_bMIFxpYM3_0),.clk(gclk));
	jdff dff_B_rKsRR8B18_0(.din(n886),.dout(w_dff_B_rKsRR8B18_0),.clk(gclk));
	jdff dff_B_vnNcVzFb2_0(.din(w_dff_B_rKsRR8B18_0),.dout(w_dff_B_vnNcVzFb2_0),.clk(gclk));
	jdff dff_B_ypXc36Wq4_0(.din(w_dff_B_vnNcVzFb2_0),.dout(w_dff_B_ypXc36Wq4_0),.clk(gclk));
	jdff dff_B_LROI9fzx7_0(.din(w_dff_B_ypXc36Wq4_0),.dout(w_dff_B_LROI9fzx7_0),.clk(gclk));
	jdff dff_B_0LUjabfV5_0(.din(w_dff_B_LROI9fzx7_0),.dout(w_dff_B_0LUjabfV5_0),.clk(gclk));
	jdff dff_B_dXjo6nTt4_0(.din(w_dff_B_0LUjabfV5_0),.dout(w_dff_B_dXjo6nTt4_0),.clk(gclk));
	jdff dff_B_Jp0UzgZy1_0(.din(w_dff_B_dXjo6nTt4_0),.dout(w_dff_B_Jp0UzgZy1_0),.clk(gclk));
	jdff dff_B_NPhRZJrd5_0(.din(w_dff_B_Jp0UzgZy1_0),.dout(w_dff_B_NPhRZJrd5_0),.clk(gclk));
	jdff dff_B_1aR2wi9I6_0(.din(w_dff_B_NPhRZJrd5_0),.dout(w_dff_B_1aR2wi9I6_0),.clk(gclk));
	jdff dff_B_P9ww9zfi6_0(.din(w_dff_B_1aR2wi9I6_0),.dout(w_dff_B_P9ww9zfi6_0),.clk(gclk));
	jdff dff_B_iwGZ0xgm9_0(.din(w_dff_B_P9ww9zfi6_0),.dout(w_dff_B_iwGZ0xgm9_0),.clk(gclk));
	jdff dff_B_WamPNYCx7_0(.din(w_dff_B_iwGZ0xgm9_0),.dout(w_dff_B_WamPNYCx7_0),.clk(gclk));
	jdff dff_B_0Dw2PQsd0_0(.din(w_dff_B_WamPNYCx7_0),.dout(w_dff_B_0Dw2PQsd0_0),.clk(gclk));
	jdff dff_B_uf1tXRsq0_0(.din(w_dff_B_0Dw2PQsd0_0),.dout(w_dff_B_uf1tXRsq0_0),.clk(gclk));
	jdff dff_B_pwH8bMZx2_0(.din(w_dff_B_uf1tXRsq0_0),.dout(w_dff_B_pwH8bMZx2_0),.clk(gclk));
	jdff dff_B_p9vSNjcF4_0(.din(w_dff_B_pwH8bMZx2_0),.dout(w_dff_B_p9vSNjcF4_0),.clk(gclk));
	jdff dff_B_gMihCNna4_0(.din(w_dff_B_p9vSNjcF4_0),.dout(w_dff_B_gMihCNna4_0),.clk(gclk));
	jdff dff_B_AnQv7iFL8_0(.din(w_dff_B_gMihCNna4_0),.dout(w_dff_B_AnQv7iFL8_0),.clk(gclk));
	jdff dff_B_6RfPHC5O5_0(.din(w_dff_B_AnQv7iFL8_0),.dout(w_dff_B_6RfPHC5O5_0),.clk(gclk));
	jdff dff_B_CNbq6GG21_0(.din(w_dff_B_6RfPHC5O5_0),.dout(w_dff_B_CNbq6GG21_0),.clk(gclk));
	jdff dff_B_cdO0cDLa8_0(.din(w_dff_B_CNbq6GG21_0),.dout(w_dff_B_cdO0cDLa8_0),.clk(gclk));
	jdff dff_B_N8p7dnMX3_0(.din(w_dff_B_cdO0cDLa8_0),.dout(w_dff_B_N8p7dnMX3_0),.clk(gclk));
	jdff dff_B_wml7S8l84_0(.din(w_dff_B_N8p7dnMX3_0),.dout(w_dff_B_wml7S8l84_0),.clk(gclk));
	jdff dff_B_M3Xd1PhB9_0(.din(w_dff_B_wml7S8l84_0),.dout(w_dff_B_M3Xd1PhB9_0),.clk(gclk));
	jdff dff_B_Gqd7YsOb9_0(.din(w_dff_B_M3Xd1PhB9_0),.dout(w_dff_B_Gqd7YsOb9_0),.clk(gclk));
	jdff dff_B_HE8KoRyj2_0(.din(w_dff_B_Gqd7YsOb9_0),.dout(w_dff_B_HE8KoRyj2_0),.clk(gclk));
	jdff dff_B_e9oF98zB1_0(.din(w_dff_B_HE8KoRyj2_0),.dout(w_dff_B_e9oF98zB1_0),.clk(gclk));
	jdff dff_B_4BEID9NH3_0(.din(w_dff_B_e9oF98zB1_0),.dout(w_dff_B_4BEID9NH3_0),.clk(gclk));
	jdff dff_B_Xcol17ju2_0(.din(w_dff_B_4BEID9NH3_0),.dout(w_dff_B_Xcol17ju2_0),.clk(gclk));
	jdff dff_B_9yfiXWsL3_0(.din(w_dff_B_Xcol17ju2_0),.dout(w_dff_B_9yfiXWsL3_0),.clk(gclk));
	jdff dff_B_dtPwKSWL7_0(.din(w_dff_B_9yfiXWsL3_0),.dout(w_dff_B_dtPwKSWL7_0),.clk(gclk));
	jdff dff_B_26hbwKBH1_0(.din(w_dff_B_dtPwKSWL7_0),.dout(w_dff_B_26hbwKBH1_0),.clk(gclk));
	jdff dff_B_2elusBl54_0(.din(w_dff_B_26hbwKBH1_0),.dout(w_dff_B_2elusBl54_0),.clk(gclk));
	jdff dff_B_hIGgbbcT3_0(.din(w_dff_B_2elusBl54_0),.dout(w_dff_B_hIGgbbcT3_0),.clk(gclk));
	jdff dff_B_RbHYZcMO1_0(.din(w_dff_B_hIGgbbcT3_0),.dout(w_dff_B_RbHYZcMO1_0),.clk(gclk));
	jdff dff_B_ugTyCguP0_0(.din(w_dff_B_RbHYZcMO1_0),.dout(w_dff_B_ugTyCguP0_0),.clk(gclk));
	jdff dff_B_Of2N23Ai3_0(.din(w_dff_B_ugTyCguP0_0),.dout(w_dff_B_Of2N23Ai3_0),.clk(gclk));
	jdff dff_B_bs1bV4Vw5_0(.din(w_dff_B_Of2N23Ai3_0),.dout(w_dff_B_bs1bV4Vw5_0),.clk(gclk));
	jdff dff_B_elqrmwr35_0(.din(w_dff_B_bs1bV4Vw5_0),.dout(w_dff_B_elqrmwr35_0),.clk(gclk));
	jdff dff_B_0Yegmpe35_0(.din(w_dff_B_elqrmwr35_0),.dout(w_dff_B_0Yegmpe35_0),.clk(gclk));
	jdff dff_B_HJwMHHa77_0(.din(w_dff_B_0Yegmpe35_0),.dout(w_dff_B_HJwMHHa77_0),.clk(gclk));
	jdff dff_B_XYONRpMX3_0(.din(w_dff_B_HJwMHHa77_0),.dout(w_dff_B_XYONRpMX3_0),.clk(gclk));
	jdff dff_B_5nRM0Uqo0_0(.din(w_dff_B_XYONRpMX3_0),.dout(w_dff_B_5nRM0Uqo0_0),.clk(gclk));
	jdff dff_B_csfMFrXb0_0(.din(w_dff_B_5nRM0Uqo0_0),.dout(w_dff_B_csfMFrXb0_0),.clk(gclk));
	jdff dff_B_gwaIQQGJ1_0(.din(w_dff_B_csfMFrXb0_0),.dout(w_dff_B_gwaIQQGJ1_0),.clk(gclk));
	jdff dff_B_IoPXxkKg5_0(.din(w_dff_B_gwaIQQGJ1_0),.dout(w_dff_B_IoPXxkKg5_0),.clk(gclk));
	jdff dff_B_Y6tCexmv9_0(.din(w_dff_B_IoPXxkKg5_0),.dout(w_dff_B_Y6tCexmv9_0),.clk(gclk));
	jdff dff_B_TbGpQ9YR5_0(.din(w_dff_B_Y6tCexmv9_0),.dout(w_dff_B_TbGpQ9YR5_0),.clk(gclk));
	jdff dff_B_V8nrYw8x2_0(.din(w_dff_B_TbGpQ9YR5_0),.dout(w_dff_B_V8nrYw8x2_0),.clk(gclk));
	jdff dff_B_4AuacWxR4_0(.din(w_dff_B_V8nrYw8x2_0),.dout(w_dff_B_4AuacWxR4_0),.clk(gclk));
	jdff dff_B_z6eD9FLQ9_0(.din(w_dff_B_4AuacWxR4_0),.dout(w_dff_B_z6eD9FLQ9_0),.clk(gclk));
	jdff dff_B_YtT6L74T6_0(.din(w_dff_B_z6eD9FLQ9_0),.dout(w_dff_B_YtT6L74T6_0),.clk(gclk));
	jdff dff_B_rQwbrXEg3_0(.din(w_dff_B_YtT6L74T6_0),.dout(w_dff_B_rQwbrXEg3_0),.clk(gclk));
	jdff dff_B_MImpxCfY7_0(.din(w_dff_B_rQwbrXEg3_0),.dout(w_dff_B_MImpxCfY7_0),.clk(gclk));
	jdff dff_B_RhWXRdSz7_0(.din(w_dff_B_MImpxCfY7_0),.dout(w_dff_B_RhWXRdSz7_0),.clk(gclk));
	jdff dff_B_e3grjneL8_0(.din(w_dff_B_RhWXRdSz7_0),.dout(w_dff_B_e3grjneL8_0),.clk(gclk));
	jdff dff_B_z6SUyQQp6_0(.din(w_dff_B_e3grjneL8_0),.dout(w_dff_B_z6SUyQQp6_0),.clk(gclk));
	jdff dff_B_wvitVInD3_0(.din(w_dff_B_z6SUyQQp6_0),.dout(w_dff_B_wvitVInD3_0),.clk(gclk));
	jdff dff_B_EJHIp3Av6_0(.din(w_dff_B_wvitVInD3_0),.dout(w_dff_B_EJHIp3Av6_0),.clk(gclk));
	jdff dff_B_fJIXlK8j6_0(.din(w_dff_B_EJHIp3Av6_0),.dout(w_dff_B_fJIXlK8j6_0),.clk(gclk));
	jdff dff_B_Ws8gdIGU2_0(.din(w_dff_B_fJIXlK8j6_0),.dout(w_dff_B_Ws8gdIGU2_0),.clk(gclk));
	jdff dff_B_rOlXoMoq9_0(.din(w_dff_B_Ws8gdIGU2_0),.dout(w_dff_B_rOlXoMoq9_0),.clk(gclk));
	jdff dff_B_rZsyBN5D7_0(.din(w_dff_B_rOlXoMoq9_0),.dout(w_dff_B_rZsyBN5D7_0),.clk(gclk));
	jdff dff_B_zadZWYrj3_0(.din(w_dff_B_rZsyBN5D7_0),.dout(w_dff_B_zadZWYrj3_0),.clk(gclk));
	jdff dff_B_dcTCKUgQ6_0(.din(w_dff_B_zadZWYrj3_0),.dout(w_dff_B_dcTCKUgQ6_0),.clk(gclk));
	jdff dff_B_Lw6x3nZ96_0(.din(w_dff_B_dcTCKUgQ6_0),.dout(w_dff_B_Lw6x3nZ96_0),.clk(gclk));
	jdff dff_B_PcOoyN266_0(.din(w_dff_B_Lw6x3nZ96_0),.dout(w_dff_B_PcOoyN266_0),.clk(gclk));
	jdff dff_B_C55CvjRy9_0(.din(w_dff_B_PcOoyN266_0),.dout(w_dff_B_C55CvjRy9_0),.clk(gclk));
	jdff dff_B_roifZn3K3_0(.din(w_dff_B_C55CvjRy9_0),.dout(w_dff_B_roifZn3K3_0),.clk(gclk));
	jdff dff_B_pwWdYu5t7_0(.din(w_dff_B_roifZn3K3_0),.dout(w_dff_B_pwWdYu5t7_0),.clk(gclk));
	jdff dff_B_5ERMbAsv8_0(.din(w_dff_B_pwWdYu5t7_0),.dout(w_dff_B_5ERMbAsv8_0),.clk(gclk));
	jdff dff_B_9IDcgHzL3_0(.din(w_dff_B_5ERMbAsv8_0),.dout(w_dff_B_9IDcgHzL3_0),.clk(gclk));
	jdff dff_B_W05GYXOh1_0(.din(w_dff_B_9IDcgHzL3_0),.dout(w_dff_B_W05GYXOh1_0),.clk(gclk));
	jdff dff_B_HeNdTa4F7_0(.din(w_dff_B_W05GYXOh1_0),.dout(w_dff_B_HeNdTa4F7_0),.clk(gclk));
	jdff dff_B_Uz6RhHJw9_0(.din(w_dff_B_HeNdTa4F7_0),.dout(w_dff_B_Uz6RhHJw9_0),.clk(gclk));
	jdff dff_B_gIlfMgXj1_0(.din(w_dff_B_Uz6RhHJw9_0),.dout(w_dff_B_gIlfMgXj1_0),.clk(gclk));
	jdff dff_B_xT417Rx08_0(.din(w_dff_B_gIlfMgXj1_0),.dout(w_dff_B_xT417Rx08_0),.clk(gclk));
	jdff dff_B_OCjNPtMl5_0(.din(w_dff_B_xT417Rx08_0),.dout(w_dff_B_OCjNPtMl5_0),.clk(gclk));
	jdff dff_B_pagZ7sfW8_0(.din(w_dff_B_OCjNPtMl5_0),.dout(w_dff_B_pagZ7sfW8_0),.clk(gclk));
	jdff dff_B_fjVtRjPI3_0(.din(w_dff_B_pagZ7sfW8_0),.dout(w_dff_B_fjVtRjPI3_0),.clk(gclk));
	jdff dff_B_zS96C8NC1_0(.din(w_dff_B_fjVtRjPI3_0),.dout(w_dff_B_zS96C8NC1_0),.clk(gclk));
	jdff dff_B_clO5nt7m5_0(.din(w_dff_B_zS96C8NC1_0),.dout(w_dff_B_clO5nt7m5_0),.clk(gclk));
	jdff dff_B_zUsR3Qhs2_0(.din(w_dff_B_clO5nt7m5_0),.dout(w_dff_B_zUsR3Qhs2_0),.clk(gclk));
	jdff dff_B_RbhAgwFf4_0(.din(n892),.dout(w_dff_B_RbhAgwFf4_0),.clk(gclk));
	jdff dff_B_gNa9njv67_0(.din(w_dff_B_RbhAgwFf4_0),.dout(w_dff_B_gNa9njv67_0),.clk(gclk));
	jdff dff_B_8M7dDNxy3_0(.din(w_dff_B_gNa9njv67_0),.dout(w_dff_B_8M7dDNxy3_0),.clk(gclk));
	jdff dff_B_q3ro8XNg6_0(.din(w_dff_B_8M7dDNxy3_0),.dout(w_dff_B_q3ro8XNg6_0),.clk(gclk));
	jdff dff_B_rkbdtrsH9_0(.din(w_dff_B_q3ro8XNg6_0),.dout(w_dff_B_rkbdtrsH9_0),.clk(gclk));
	jdff dff_B_r1GeerKW4_0(.din(w_dff_B_rkbdtrsH9_0),.dout(w_dff_B_r1GeerKW4_0),.clk(gclk));
	jdff dff_B_HwS05xRY1_0(.din(w_dff_B_r1GeerKW4_0),.dout(w_dff_B_HwS05xRY1_0),.clk(gclk));
	jdff dff_B_npdJYG3I4_0(.din(w_dff_B_HwS05xRY1_0),.dout(w_dff_B_npdJYG3I4_0),.clk(gclk));
	jdff dff_B_koDB1nkq4_0(.din(w_dff_B_npdJYG3I4_0),.dout(w_dff_B_koDB1nkq4_0),.clk(gclk));
	jdff dff_B_Q6VX4Jaw0_0(.din(w_dff_B_koDB1nkq4_0),.dout(w_dff_B_Q6VX4Jaw0_0),.clk(gclk));
	jdff dff_B_Qv1b7M2u7_0(.din(w_dff_B_Q6VX4Jaw0_0),.dout(w_dff_B_Qv1b7M2u7_0),.clk(gclk));
	jdff dff_B_VWUtoWC62_0(.din(w_dff_B_Qv1b7M2u7_0),.dout(w_dff_B_VWUtoWC62_0),.clk(gclk));
	jdff dff_B_8WOLjRNy1_0(.din(w_dff_B_VWUtoWC62_0),.dout(w_dff_B_8WOLjRNy1_0),.clk(gclk));
	jdff dff_B_0zJCpDAt8_0(.din(w_dff_B_8WOLjRNy1_0),.dout(w_dff_B_0zJCpDAt8_0),.clk(gclk));
	jdff dff_B_T6wLnEUA3_0(.din(w_dff_B_0zJCpDAt8_0),.dout(w_dff_B_T6wLnEUA3_0),.clk(gclk));
	jdff dff_B_e5rNi6qV1_0(.din(w_dff_B_T6wLnEUA3_0),.dout(w_dff_B_e5rNi6qV1_0),.clk(gclk));
	jdff dff_B_Zsje3hqI7_0(.din(w_dff_B_e5rNi6qV1_0),.dout(w_dff_B_Zsje3hqI7_0),.clk(gclk));
	jdff dff_B_88gHF54N1_0(.din(w_dff_B_Zsje3hqI7_0),.dout(w_dff_B_88gHF54N1_0),.clk(gclk));
	jdff dff_B_9lBvPZZl7_0(.din(w_dff_B_88gHF54N1_0),.dout(w_dff_B_9lBvPZZl7_0),.clk(gclk));
	jdff dff_B_QmEDQSCh9_0(.din(w_dff_B_9lBvPZZl7_0),.dout(w_dff_B_QmEDQSCh9_0),.clk(gclk));
	jdff dff_B_Fg25dwkf4_0(.din(w_dff_B_QmEDQSCh9_0),.dout(w_dff_B_Fg25dwkf4_0),.clk(gclk));
	jdff dff_B_49ZjzouG7_0(.din(w_dff_B_Fg25dwkf4_0),.dout(w_dff_B_49ZjzouG7_0),.clk(gclk));
	jdff dff_B_4M59PWGc6_0(.din(w_dff_B_49ZjzouG7_0),.dout(w_dff_B_4M59PWGc6_0),.clk(gclk));
	jdff dff_B_wSdLjt7N9_0(.din(w_dff_B_4M59PWGc6_0),.dout(w_dff_B_wSdLjt7N9_0),.clk(gclk));
	jdff dff_B_j11bFsza9_0(.din(w_dff_B_wSdLjt7N9_0),.dout(w_dff_B_j11bFsza9_0),.clk(gclk));
	jdff dff_B_OhATlEu27_0(.din(w_dff_B_j11bFsza9_0),.dout(w_dff_B_OhATlEu27_0),.clk(gclk));
	jdff dff_B_vRIIBHzo3_0(.din(w_dff_B_OhATlEu27_0),.dout(w_dff_B_vRIIBHzo3_0),.clk(gclk));
	jdff dff_B_X3atVQTg5_0(.din(w_dff_B_vRIIBHzo3_0),.dout(w_dff_B_X3atVQTg5_0),.clk(gclk));
	jdff dff_B_JrwEpjyr2_0(.din(w_dff_B_X3atVQTg5_0),.dout(w_dff_B_JrwEpjyr2_0),.clk(gclk));
	jdff dff_B_Y98Q8kZG6_0(.din(w_dff_B_JrwEpjyr2_0),.dout(w_dff_B_Y98Q8kZG6_0),.clk(gclk));
	jdff dff_B_p54lXqII9_0(.din(w_dff_B_Y98Q8kZG6_0),.dout(w_dff_B_p54lXqII9_0),.clk(gclk));
	jdff dff_B_NO92IF1B7_0(.din(w_dff_B_p54lXqII9_0),.dout(w_dff_B_NO92IF1B7_0),.clk(gclk));
	jdff dff_B_jK6mh18C6_0(.din(w_dff_B_NO92IF1B7_0),.dout(w_dff_B_jK6mh18C6_0),.clk(gclk));
	jdff dff_B_96gAZREG5_0(.din(w_dff_B_jK6mh18C6_0),.dout(w_dff_B_96gAZREG5_0),.clk(gclk));
	jdff dff_B_bwacqj0h4_0(.din(w_dff_B_96gAZREG5_0),.dout(w_dff_B_bwacqj0h4_0),.clk(gclk));
	jdff dff_B_qOsBJCSs0_0(.din(w_dff_B_bwacqj0h4_0),.dout(w_dff_B_qOsBJCSs0_0),.clk(gclk));
	jdff dff_B_ASwJeVNh8_0(.din(w_dff_B_qOsBJCSs0_0),.dout(w_dff_B_ASwJeVNh8_0),.clk(gclk));
	jdff dff_B_tu9n90Yi2_0(.din(w_dff_B_ASwJeVNh8_0),.dout(w_dff_B_tu9n90Yi2_0),.clk(gclk));
	jdff dff_B_cZXH2y5q2_0(.din(w_dff_B_tu9n90Yi2_0),.dout(w_dff_B_cZXH2y5q2_0),.clk(gclk));
	jdff dff_B_5fv9iXVj7_0(.din(w_dff_B_cZXH2y5q2_0),.dout(w_dff_B_5fv9iXVj7_0),.clk(gclk));
	jdff dff_B_HwpyzPsg3_0(.din(w_dff_B_5fv9iXVj7_0),.dout(w_dff_B_HwpyzPsg3_0),.clk(gclk));
	jdff dff_B_DWZvWsa45_0(.din(w_dff_B_HwpyzPsg3_0),.dout(w_dff_B_DWZvWsa45_0),.clk(gclk));
	jdff dff_B_aIMOrtzc2_0(.din(w_dff_B_DWZvWsa45_0),.dout(w_dff_B_aIMOrtzc2_0),.clk(gclk));
	jdff dff_B_qclTWQc92_0(.din(w_dff_B_aIMOrtzc2_0),.dout(w_dff_B_qclTWQc92_0),.clk(gclk));
	jdff dff_B_l9LFpjIh4_0(.din(w_dff_B_qclTWQc92_0),.dout(w_dff_B_l9LFpjIh4_0),.clk(gclk));
	jdff dff_B_mpEr5KH37_0(.din(w_dff_B_l9LFpjIh4_0),.dout(w_dff_B_mpEr5KH37_0),.clk(gclk));
	jdff dff_B_52FqaxSt7_0(.din(w_dff_B_mpEr5KH37_0),.dout(w_dff_B_52FqaxSt7_0),.clk(gclk));
	jdff dff_B_hvLK5edJ2_0(.din(w_dff_B_52FqaxSt7_0),.dout(w_dff_B_hvLK5edJ2_0),.clk(gclk));
	jdff dff_B_xdPZG6vH2_0(.din(w_dff_B_hvLK5edJ2_0),.dout(w_dff_B_xdPZG6vH2_0),.clk(gclk));
	jdff dff_B_ZtE1BT2l8_0(.din(w_dff_B_xdPZG6vH2_0),.dout(w_dff_B_ZtE1BT2l8_0),.clk(gclk));
	jdff dff_B_fT6YRSrD8_0(.din(w_dff_B_ZtE1BT2l8_0),.dout(w_dff_B_fT6YRSrD8_0),.clk(gclk));
	jdff dff_B_wcjQj3bN8_0(.din(w_dff_B_fT6YRSrD8_0),.dout(w_dff_B_wcjQj3bN8_0),.clk(gclk));
	jdff dff_B_bSi6h9OL1_0(.din(w_dff_B_wcjQj3bN8_0),.dout(w_dff_B_bSi6h9OL1_0),.clk(gclk));
	jdff dff_B_z2nodQ5C6_0(.din(w_dff_B_bSi6h9OL1_0),.dout(w_dff_B_z2nodQ5C6_0),.clk(gclk));
	jdff dff_B_n5fYwwXW8_0(.din(w_dff_B_z2nodQ5C6_0),.dout(w_dff_B_n5fYwwXW8_0),.clk(gclk));
	jdff dff_B_1ZNI3kEJ1_0(.din(w_dff_B_n5fYwwXW8_0),.dout(w_dff_B_1ZNI3kEJ1_0),.clk(gclk));
	jdff dff_B_LJZC9NRv6_0(.din(w_dff_B_1ZNI3kEJ1_0),.dout(w_dff_B_LJZC9NRv6_0),.clk(gclk));
	jdff dff_B_qjOYAvwg1_0(.din(w_dff_B_LJZC9NRv6_0),.dout(w_dff_B_qjOYAvwg1_0),.clk(gclk));
	jdff dff_B_U7aOzUv02_0(.din(w_dff_B_qjOYAvwg1_0),.dout(w_dff_B_U7aOzUv02_0),.clk(gclk));
	jdff dff_B_X6D9I1ru0_0(.din(w_dff_B_U7aOzUv02_0),.dout(w_dff_B_X6D9I1ru0_0),.clk(gclk));
	jdff dff_B_TnML09fW1_0(.din(w_dff_B_X6D9I1ru0_0),.dout(w_dff_B_TnML09fW1_0),.clk(gclk));
	jdff dff_B_WJrzA8LD4_0(.din(w_dff_B_TnML09fW1_0),.dout(w_dff_B_WJrzA8LD4_0),.clk(gclk));
	jdff dff_B_nAiRgwlH5_0(.din(w_dff_B_WJrzA8LD4_0),.dout(w_dff_B_nAiRgwlH5_0),.clk(gclk));
	jdff dff_B_i4A5QtzN0_0(.din(w_dff_B_nAiRgwlH5_0),.dout(w_dff_B_i4A5QtzN0_0),.clk(gclk));
	jdff dff_B_dXZMItQ46_0(.din(w_dff_B_i4A5QtzN0_0),.dout(w_dff_B_dXZMItQ46_0),.clk(gclk));
	jdff dff_B_K8ukcugw7_0(.din(w_dff_B_dXZMItQ46_0),.dout(w_dff_B_K8ukcugw7_0),.clk(gclk));
	jdff dff_B_h61f6hzY5_0(.din(w_dff_B_K8ukcugw7_0),.dout(w_dff_B_h61f6hzY5_0),.clk(gclk));
	jdff dff_B_sVa8StLI5_0(.din(w_dff_B_h61f6hzY5_0),.dout(w_dff_B_sVa8StLI5_0),.clk(gclk));
	jdff dff_B_vCxsbMFU3_0(.din(w_dff_B_sVa8StLI5_0),.dout(w_dff_B_vCxsbMFU3_0),.clk(gclk));
	jdff dff_B_9nQbLlzI0_0(.din(w_dff_B_vCxsbMFU3_0),.dout(w_dff_B_9nQbLlzI0_0),.clk(gclk));
	jdff dff_B_n1EMLMJy0_0(.din(w_dff_B_9nQbLlzI0_0),.dout(w_dff_B_n1EMLMJy0_0),.clk(gclk));
	jdff dff_B_EUPZZoSL6_0(.din(w_dff_B_n1EMLMJy0_0),.dout(w_dff_B_EUPZZoSL6_0),.clk(gclk));
	jdff dff_B_SSH81M866_0(.din(w_dff_B_EUPZZoSL6_0),.dout(w_dff_B_SSH81M866_0),.clk(gclk));
	jdff dff_B_mM8auC6O1_0(.din(w_dff_B_SSH81M866_0),.dout(w_dff_B_mM8auC6O1_0),.clk(gclk));
	jdff dff_B_x3oRt3C52_0(.din(w_dff_B_mM8auC6O1_0),.dout(w_dff_B_x3oRt3C52_0),.clk(gclk));
	jdff dff_B_KrPqwPbq3_0(.din(w_dff_B_x3oRt3C52_0),.dout(w_dff_B_KrPqwPbq3_0),.clk(gclk));
	jdff dff_B_DGGLKCV08_0(.din(w_dff_B_KrPqwPbq3_0),.dout(w_dff_B_DGGLKCV08_0),.clk(gclk));
	jdff dff_B_Sl5uAGPc7_0(.din(w_dff_B_DGGLKCV08_0),.dout(w_dff_B_Sl5uAGPc7_0),.clk(gclk));
	jdff dff_B_5CJTdA2k2_0(.din(w_dff_B_Sl5uAGPc7_0),.dout(w_dff_B_5CJTdA2k2_0),.clk(gclk));
	jdff dff_B_ku9hUzde0_0(.din(w_dff_B_5CJTdA2k2_0),.dout(w_dff_B_ku9hUzde0_0),.clk(gclk));
	jdff dff_B_YBNOgsWi6_0(.din(w_dff_B_ku9hUzde0_0),.dout(w_dff_B_YBNOgsWi6_0),.clk(gclk));
	jdff dff_B_4OTtZhrV7_0(.din(w_dff_B_YBNOgsWi6_0),.dout(w_dff_B_4OTtZhrV7_0),.clk(gclk));
	jdff dff_B_xRFEj3YO8_0(.din(w_dff_B_4OTtZhrV7_0),.dout(w_dff_B_xRFEj3YO8_0),.clk(gclk));
	jdff dff_B_tgwVYjIg3_0(.din(w_dff_B_xRFEj3YO8_0),.dout(w_dff_B_tgwVYjIg3_0),.clk(gclk));
	jdff dff_B_7fpLCNfK4_0(.din(n898),.dout(w_dff_B_7fpLCNfK4_0),.clk(gclk));
	jdff dff_B_F2e0qTWi8_0(.din(w_dff_B_7fpLCNfK4_0),.dout(w_dff_B_F2e0qTWi8_0),.clk(gclk));
	jdff dff_B_MxSY16zF0_0(.din(w_dff_B_F2e0qTWi8_0),.dout(w_dff_B_MxSY16zF0_0),.clk(gclk));
	jdff dff_B_IrsYUVUH1_0(.din(w_dff_B_MxSY16zF0_0),.dout(w_dff_B_IrsYUVUH1_0),.clk(gclk));
	jdff dff_B_MsxkzGhm3_0(.din(w_dff_B_IrsYUVUH1_0),.dout(w_dff_B_MsxkzGhm3_0),.clk(gclk));
	jdff dff_B_JFxKYQfw4_0(.din(w_dff_B_MsxkzGhm3_0),.dout(w_dff_B_JFxKYQfw4_0),.clk(gclk));
	jdff dff_B_SofAR1CR7_0(.din(w_dff_B_JFxKYQfw4_0),.dout(w_dff_B_SofAR1CR7_0),.clk(gclk));
	jdff dff_B_z3DGAngw5_0(.din(w_dff_B_SofAR1CR7_0),.dout(w_dff_B_z3DGAngw5_0),.clk(gclk));
	jdff dff_B_hPdt6xMi3_0(.din(w_dff_B_z3DGAngw5_0),.dout(w_dff_B_hPdt6xMi3_0),.clk(gclk));
	jdff dff_B_mFrJLiJ80_0(.din(w_dff_B_hPdt6xMi3_0),.dout(w_dff_B_mFrJLiJ80_0),.clk(gclk));
	jdff dff_B_bTwy420H5_0(.din(w_dff_B_mFrJLiJ80_0),.dout(w_dff_B_bTwy420H5_0),.clk(gclk));
	jdff dff_B_cLuCe9RC7_0(.din(w_dff_B_bTwy420H5_0),.dout(w_dff_B_cLuCe9RC7_0),.clk(gclk));
	jdff dff_B_jtPbMuU01_0(.din(w_dff_B_cLuCe9RC7_0),.dout(w_dff_B_jtPbMuU01_0),.clk(gclk));
	jdff dff_B_k05MxG376_0(.din(w_dff_B_jtPbMuU01_0),.dout(w_dff_B_k05MxG376_0),.clk(gclk));
	jdff dff_B_BPzy3ys37_0(.din(w_dff_B_k05MxG376_0),.dout(w_dff_B_BPzy3ys37_0),.clk(gclk));
	jdff dff_B_VqP6rJBB0_0(.din(w_dff_B_BPzy3ys37_0),.dout(w_dff_B_VqP6rJBB0_0),.clk(gclk));
	jdff dff_B_fOVkZ61s4_0(.din(w_dff_B_VqP6rJBB0_0),.dout(w_dff_B_fOVkZ61s4_0),.clk(gclk));
	jdff dff_B_DVNaRLwH1_0(.din(w_dff_B_fOVkZ61s4_0),.dout(w_dff_B_DVNaRLwH1_0),.clk(gclk));
	jdff dff_B_jmmV1UR48_0(.din(w_dff_B_DVNaRLwH1_0),.dout(w_dff_B_jmmV1UR48_0),.clk(gclk));
	jdff dff_B_Kc2Vev8J5_0(.din(w_dff_B_jmmV1UR48_0),.dout(w_dff_B_Kc2Vev8J5_0),.clk(gclk));
	jdff dff_B_StlBTWAv5_0(.din(w_dff_B_Kc2Vev8J5_0),.dout(w_dff_B_StlBTWAv5_0),.clk(gclk));
	jdff dff_B_DTWPbApp7_0(.din(w_dff_B_StlBTWAv5_0),.dout(w_dff_B_DTWPbApp7_0),.clk(gclk));
	jdff dff_B_ImRRhKX16_0(.din(w_dff_B_DTWPbApp7_0),.dout(w_dff_B_ImRRhKX16_0),.clk(gclk));
	jdff dff_B_T7cuqgKe6_0(.din(w_dff_B_ImRRhKX16_0),.dout(w_dff_B_T7cuqgKe6_0),.clk(gclk));
	jdff dff_B_26iXzTi24_0(.din(w_dff_B_T7cuqgKe6_0),.dout(w_dff_B_26iXzTi24_0),.clk(gclk));
	jdff dff_B_P5raa7iH5_0(.din(w_dff_B_26iXzTi24_0),.dout(w_dff_B_P5raa7iH5_0),.clk(gclk));
	jdff dff_B_534qgITM8_0(.din(w_dff_B_P5raa7iH5_0),.dout(w_dff_B_534qgITM8_0),.clk(gclk));
	jdff dff_B_pjy9kEid4_0(.din(w_dff_B_534qgITM8_0),.dout(w_dff_B_pjy9kEid4_0),.clk(gclk));
	jdff dff_B_IrLGOxd82_0(.din(w_dff_B_pjy9kEid4_0),.dout(w_dff_B_IrLGOxd82_0),.clk(gclk));
	jdff dff_B_LfZuWKDf0_0(.din(w_dff_B_IrLGOxd82_0),.dout(w_dff_B_LfZuWKDf0_0),.clk(gclk));
	jdff dff_B_oMjt1qKM8_0(.din(w_dff_B_LfZuWKDf0_0),.dout(w_dff_B_oMjt1qKM8_0),.clk(gclk));
	jdff dff_B_vO8bFBFu7_0(.din(w_dff_B_oMjt1qKM8_0),.dout(w_dff_B_vO8bFBFu7_0),.clk(gclk));
	jdff dff_B_RqF7z6ix8_0(.din(w_dff_B_vO8bFBFu7_0),.dout(w_dff_B_RqF7z6ix8_0),.clk(gclk));
	jdff dff_B_wboFmJWv1_0(.din(w_dff_B_RqF7z6ix8_0),.dout(w_dff_B_wboFmJWv1_0),.clk(gclk));
	jdff dff_B_9oT9nGjG2_0(.din(w_dff_B_wboFmJWv1_0),.dout(w_dff_B_9oT9nGjG2_0),.clk(gclk));
	jdff dff_B_zSCdU7MV5_0(.din(w_dff_B_9oT9nGjG2_0),.dout(w_dff_B_zSCdU7MV5_0),.clk(gclk));
	jdff dff_B_EV00l0fe4_0(.din(w_dff_B_zSCdU7MV5_0),.dout(w_dff_B_EV00l0fe4_0),.clk(gclk));
	jdff dff_B_EcNQHBKi3_0(.din(w_dff_B_EV00l0fe4_0),.dout(w_dff_B_EcNQHBKi3_0),.clk(gclk));
	jdff dff_B_ZRCvYCot5_0(.din(w_dff_B_EcNQHBKi3_0),.dout(w_dff_B_ZRCvYCot5_0),.clk(gclk));
	jdff dff_B_ptdetvH26_0(.din(w_dff_B_ZRCvYCot5_0),.dout(w_dff_B_ptdetvH26_0),.clk(gclk));
	jdff dff_B_kZfIIG5p1_0(.din(w_dff_B_ptdetvH26_0),.dout(w_dff_B_kZfIIG5p1_0),.clk(gclk));
	jdff dff_B_9E9LPpF47_0(.din(w_dff_B_kZfIIG5p1_0),.dout(w_dff_B_9E9LPpF47_0),.clk(gclk));
	jdff dff_B_cHRf4jFS6_0(.din(w_dff_B_9E9LPpF47_0),.dout(w_dff_B_cHRf4jFS6_0),.clk(gclk));
	jdff dff_B_GpbFh6gO8_0(.din(w_dff_B_cHRf4jFS6_0),.dout(w_dff_B_GpbFh6gO8_0),.clk(gclk));
	jdff dff_B_XhbPu0R95_0(.din(w_dff_B_GpbFh6gO8_0),.dout(w_dff_B_XhbPu0R95_0),.clk(gclk));
	jdff dff_B_RZJPVBIw7_0(.din(w_dff_B_XhbPu0R95_0),.dout(w_dff_B_RZJPVBIw7_0),.clk(gclk));
	jdff dff_B_e8Q3EY8E5_0(.din(w_dff_B_RZJPVBIw7_0),.dout(w_dff_B_e8Q3EY8E5_0),.clk(gclk));
	jdff dff_B_wf6N3ee44_0(.din(w_dff_B_e8Q3EY8E5_0),.dout(w_dff_B_wf6N3ee44_0),.clk(gclk));
	jdff dff_B_2dPm7vnJ7_0(.din(w_dff_B_wf6N3ee44_0),.dout(w_dff_B_2dPm7vnJ7_0),.clk(gclk));
	jdff dff_B_4J1Mwn6u0_0(.din(w_dff_B_2dPm7vnJ7_0),.dout(w_dff_B_4J1Mwn6u0_0),.clk(gclk));
	jdff dff_B_Ih6mbkCq0_0(.din(w_dff_B_4J1Mwn6u0_0),.dout(w_dff_B_Ih6mbkCq0_0),.clk(gclk));
	jdff dff_B_tnW2TgI04_0(.din(w_dff_B_Ih6mbkCq0_0),.dout(w_dff_B_tnW2TgI04_0),.clk(gclk));
	jdff dff_B_dZv1TT1s8_0(.din(w_dff_B_tnW2TgI04_0),.dout(w_dff_B_dZv1TT1s8_0),.clk(gclk));
	jdff dff_B_rNgmYX2U0_0(.din(w_dff_B_dZv1TT1s8_0),.dout(w_dff_B_rNgmYX2U0_0),.clk(gclk));
	jdff dff_B_ov8QcAIA5_0(.din(w_dff_B_rNgmYX2U0_0),.dout(w_dff_B_ov8QcAIA5_0),.clk(gclk));
	jdff dff_B_ONygDv806_0(.din(w_dff_B_ov8QcAIA5_0),.dout(w_dff_B_ONygDv806_0),.clk(gclk));
	jdff dff_B_14ddiKh63_0(.din(w_dff_B_ONygDv806_0),.dout(w_dff_B_14ddiKh63_0),.clk(gclk));
	jdff dff_B_Vqh54OtS2_0(.din(w_dff_B_14ddiKh63_0),.dout(w_dff_B_Vqh54OtS2_0),.clk(gclk));
	jdff dff_B_erkFpigz8_0(.din(w_dff_B_Vqh54OtS2_0),.dout(w_dff_B_erkFpigz8_0),.clk(gclk));
	jdff dff_B_qqggysAj0_0(.din(w_dff_B_erkFpigz8_0),.dout(w_dff_B_qqggysAj0_0),.clk(gclk));
	jdff dff_B_hsrFqxlp6_0(.din(w_dff_B_qqggysAj0_0),.dout(w_dff_B_hsrFqxlp6_0),.clk(gclk));
	jdff dff_B_DfPvFU655_0(.din(w_dff_B_hsrFqxlp6_0),.dout(w_dff_B_DfPvFU655_0),.clk(gclk));
	jdff dff_B_yB2s3Z0O7_0(.din(w_dff_B_DfPvFU655_0),.dout(w_dff_B_yB2s3Z0O7_0),.clk(gclk));
	jdff dff_B_VEuNX9yI7_0(.din(w_dff_B_yB2s3Z0O7_0),.dout(w_dff_B_VEuNX9yI7_0),.clk(gclk));
	jdff dff_B_8FKK6kC72_0(.din(w_dff_B_VEuNX9yI7_0),.dout(w_dff_B_8FKK6kC72_0),.clk(gclk));
	jdff dff_B_ON72gYPy2_0(.din(w_dff_B_8FKK6kC72_0),.dout(w_dff_B_ON72gYPy2_0),.clk(gclk));
	jdff dff_B_uFgbbB2u8_0(.din(w_dff_B_ON72gYPy2_0),.dout(w_dff_B_uFgbbB2u8_0),.clk(gclk));
	jdff dff_B_pj7MqDkE2_0(.din(w_dff_B_uFgbbB2u8_0),.dout(w_dff_B_pj7MqDkE2_0),.clk(gclk));
	jdff dff_B_FnWyRtqy7_0(.din(w_dff_B_pj7MqDkE2_0),.dout(w_dff_B_FnWyRtqy7_0),.clk(gclk));
	jdff dff_B_iLs3lp5Y6_0(.din(w_dff_B_FnWyRtqy7_0),.dout(w_dff_B_iLs3lp5Y6_0),.clk(gclk));
	jdff dff_B_Q8vJVLDZ4_0(.din(w_dff_B_iLs3lp5Y6_0),.dout(w_dff_B_Q8vJVLDZ4_0),.clk(gclk));
	jdff dff_B_aN0kJfLk4_0(.din(w_dff_B_Q8vJVLDZ4_0),.dout(w_dff_B_aN0kJfLk4_0),.clk(gclk));
	jdff dff_B_Cjr67EwA1_0(.din(w_dff_B_aN0kJfLk4_0),.dout(w_dff_B_Cjr67EwA1_0),.clk(gclk));
	jdff dff_B_RNMzg2Ln6_0(.din(w_dff_B_Cjr67EwA1_0),.dout(w_dff_B_RNMzg2Ln6_0),.clk(gclk));
	jdff dff_B_PGCdp9MW6_0(.din(w_dff_B_RNMzg2Ln6_0),.dout(w_dff_B_PGCdp9MW6_0),.clk(gclk));
	jdff dff_B_v6bMOoiR8_0(.din(w_dff_B_PGCdp9MW6_0),.dout(w_dff_B_v6bMOoiR8_0),.clk(gclk));
	jdff dff_B_a7LsIWB48_0(.din(w_dff_B_v6bMOoiR8_0),.dout(w_dff_B_a7LsIWB48_0),.clk(gclk));
	jdff dff_B_rtATlEVn0_0(.din(w_dff_B_a7LsIWB48_0),.dout(w_dff_B_rtATlEVn0_0),.clk(gclk));
	jdff dff_B_kjdSeWsF1_0(.din(w_dff_B_rtATlEVn0_0),.dout(w_dff_B_kjdSeWsF1_0),.clk(gclk));
	jdff dff_B_LOvX9Jjn0_0(.din(w_dff_B_kjdSeWsF1_0),.dout(w_dff_B_LOvX9Jjn0_0),.clk(gclk));
	jdff dff_B_T27tXn7v0_0(.din(w_dff_B_LOvX9Jjn0_0),.dout(w_dff_B_T27tXn7v0_0),.clk(gclk));
	jdff dff_B_SvjAMgLx0_0(.din(w_dff_B_T27tXn7v0_0),.dout(w_dff_B_SvjAMgLx0_0),.clk(gclk));
	jdff dff_B_ls4nVUQ24_0(.din(w_dff_B_SvjAMgLx0_0),.dout(w_dff_B_ls4nVUQ24_0),.clk(gclk));
	jdff dff_B_I7yf34Bu8_0(.din(w_dff_B_ls4nVUQ24_0),.dout(w_dff_B_I7yf34Bu8_0),.clk(gclk));
	jdff dff_B_EZvSDj9R9_0(.din(w_dff_B_I7yf34Bu8_0),.dout(w_dff_B_EZvSDj9R9_0),.clk(gclk));
	jdff dff_B_rBYNYFbH4_0(.din(n904),.dout(w_dff_B_rBYNYFbH4_0),.clk(gclk));
	jdff dff_B_RjY3VDr80_0(.din(w_dff_B_rBYNYFbH4_0),.dout(w_dff_B_RjY3VDr80_0),.clk(gclk));
	jdff dff_B_44rcrMNH1_0(.din(w_dff_B_RjY3VDr80_0),.dout(w_dff_B_44rcrMNH1_0),.clk(gclk));
	jdff dff_B_dU7m9MNj5_0(.din(w_dff_B_44rcrMNH1_0),.dout(w_dff_B_dU7m9MNj5_0),.clk(gclk));
	jdff dff_B_UmUYOyza3_0(.din(w_dff_B_dU7m9MNj5_0),.dout(w_dff_B_UmUYOyza3_0),.clk(gclk));
	jdff dff_B_VKB6AZcp7_0(.din(w_dff_B_UmUYOyza3_0),.dout(w_dff_B_VKB6AZcp7_0),.clk(gclk));
	jdff dff_B_Cx3jRaYD6_0(.din(w_dff_B_VKB6AZcp7_0),.dout(w_dff_B_Cx3jRaYD6_0),.clk(gclk));
	jdff dff_B_1DdhqPrz2_0(.din(w_dff_B_Cx3jRaYD6_0),.dout(w_dff_B_1DdhqPrz2_0),.clk(gclk));
	jdff dff_B_M6UwPZ8z2_0(.din(w_dff_B_1DdhqPrz2_0),.dout(w_dff_B_M6UwPZ8z2_0),.clk(gclk));
	jdff dff_B_mOnru5Gv3_0(.din(w_dff_B_M6UwPZ8z2_0),.dout(w_dff_B_mOnru5Gv3_0),.clk(gclk));
	jdff dff_B_CWkhzmp43_0(.din(w_dff_B_mOnru5Gv3_0),.dout(w_dff_B_CWkhzmp43_0),.clk(gclk));
	jdff dff_B_Sdq46Lib7_0(.din(w_dff_B_CWkhzmp43_0),.dout(w_dff_B_Sdq46Lib7_0),.clk(gclk));
	jdff dff_B_FGDPvwzl4_0(.din(w_dff_B_Sdq46Lib7_0),.dout(w_dff_B_FGDPvwzl4_0),.clk(gclk));
	jdff dff_B_9fRtXgjP7_0(.din(w_dff_B_FGDPvwzl4_0),.dout(w_dff_B_9fRtXgjP7_0),.clk(gclk));
	jdff dff_B_swH8lO7r2_0(.din(w_dff_B_9fRtXgjP7_0),.dout(w_dff_B_swH8lO7r2_0),.clk(gclk));
	jdff dff_B_FbfisYWQ7_0(.din(w_dff_B_swH8lO7r2_0),.dout(w_dff_B_FbfisYWQ7_0),.clk(gclk));
	jdff dff_B_VPGX3hye7_0(.din(w_dff_B_FbfisYWQ7_0),.dout(w_dff_B_VPGX3hye7_0),.clk(gclk));
	jdff dff_B_3dQSkHhr5_0(.din(w_dff_B_VPGX3hye7_0),.dout(w_dff_B_3dQSkHhr5_0),.clk(gclk));
	jdff dff_B_4749LPl88_0(.din(w_dff_B_3dQSkHhr5_0),.dout(w_dff_B_4749LPl88_0),.clk(gclk));
	jdff dff_B_Kr3St3gd4_0(.din(w_dff_B_4749LPl88_0),.dout(w_dff_B_Kr3St3gd4_0),.clk(gclk));
	jdff dff_B_HaJtJ9W44_0(.din(w_dff_B_Kr3St3gd4_0),.dout(w_dff_B_HaJtJ9W44_0),.clk(gclk));
	jdff dff_B_6KybQLdZ8_0(.din(w_dff_B_HaJtJ9W44_0),.dout(w_dff_B_6KybQLdZ8_0),.clk(gclk));
	jdff dff_B_1Nb0u8t70_0(.din(w_dff_B_6KybQLdZ8_0),.dout(w_dff_B_1Nb0u8t70_0),.clk(gclk));
	jdff dff_B_woAwXAuG2_0(.din(w_dff_B_1Nb0u8t70_0),.dout(w_dff_B_woAwXAuG2_0),.clk(gclk));
	jdff dff_B_XIdjPbaG5_0(.din(w_dff_B_woAwXAuG2_0),.dout(w_dff_B_XIdjPbaG5_0),.clk(gclk));
	jdff dff_B_KTNTSNLj0_0(.din(w_dff_B_XIdjPbaG5_0),.dout(w_dff_B_KTNTSNLj0_0),.clk(gclk));
	jdff dff_B_Y7OVtIdX1_0(.din(w_dff_B_KTNTSNLj0_0),.dout(w_dff_B_Y7OVtIdX1_0),.clk(gclk));
	jdff dff_B_Kz2tAwq64_0(.din(w_dff_B_Y7OVtIdX1_0),.dout(w_dff_B_Kz2tAwq64_0),.clk(gclk));
	jdff dff_B_84m8ypX36_0(.din(w_dff_B_Kz2tAwq64_0),.dout(w_dff_B_84m8ypX36_0),.clk(gclk));
	jdff dff_B_tWLcj1rx9_0(.din(w_dff_B_84m8ypX36_0),.dout(w_dff_B_tWLcj1rx9_0),.clk(gclk));
	jdff dff_B_rGPCty7D2_0(.din(w_dff_B_tWLcj1rx9_0),.dout(w_dff_B_rGPCty7D2_0),.clk(gclk));
	jdff dff_B_D7fCJeVx6_0(.din(w_dff_B_rGPCty7D2_0),.dout(w_dff_B_D7fCJeVx6_0),.clk(gclk));
	jdff dff_B_UwCUdrn85_0(.din(w_dff_B_D7fCJeVx6_0),.dout(w_dff_B_UwCUdrn85_0),.clk(gclk));
	jdff dff_B_Bs5fgbR58_0(.din(w_dff_B_UwCUdrn85_0),.dout(w_dff_B_Bs5fgbR58_0),.clk(gclk));
	jdff dff_B_6yx3Ua6u2_0(.din(w_dff_B_Bs5fgbR58_0),.dout(w_dff_B_6yx3Ua6u2_0),.clk(gclk));
	jdff dff_B_Wu6WLvLu6_0(.din(w_dff_B_6yx3Ua6u2_0),.dout(w_dff_B_Wu6WLvLu6_0),.clk(gclk));
	jdff dff_B_EiWb5KYS5_0(.din(w_dff_B_Wu6WLvLu6_0),.dout(w_dff_B_EiWb5KYS5_0),.clk(gclk));
	jdff dff_B_HcIa7fiQ1_0(.din(w_dff_B_EiWb5KYS5_0),.dout(w_dff_B_HcIa7fiQ1_0),.clk(gclk));
	jdff dff_B_VjETb8KY5_0(.din(w_dff_B_HcIa7fiQ1_0),.dout(w_dff_B_VjETb8KY5_0),.clk(gclk));
	jdff dff_B_HsADwHgF2_0(.din(w_dff_B_VjETb8KY5_0),.dout(w_dff_B_HsADwHgF2_0),.clk(gclk));
	jdff dff_B_TM57K66V9_0(.din(w_dff_B_HsADwHgF2_0),.dout(w_dff_B_TM57K66V9_0),.clk(gclk));
	jdff dff_B_vD6JUPlz0_0(.din(w_dff_B_TM57K66V9_0),.dout(w_dff_B_vD6JUPlz0_0),.clk(gclk));
	jdff dff_B_kAT3upPx2_0(.din(w_dff_B_vD6JUPlz0_0),.dout(w_dff_B_kAT3upPx2_0),.clk(gclk));
	jdff dff_B_krlCTgMQ1_0(.din(w_dff_B_kAT3upPx2_0),.dout(w_dff_B_krlCTgMQ1_0),.clk(gclk));
	jdff dff_B_FerMHviC0_0(.din(w_dff_B_krlCTgMQ1_0),.dout(w_dff_B_FerMHviC0_0),.clk(gclk));
	jdff dff_B_4ve86PSQ0_0(.din(w_dff_B_FerMHviC0_0),.dout(w_dff_B_4ve86PSQ0_0),.clk(gclk));
	jdff dff_B_aMV6Svoj8_0(.din(w_dff_B_4ve86PSQ0_0),.dout(w_dff_B_aMV6Svoj8_0),.clk(gclk));
	jdff dff_B_ejDlgELE4_0(.din(w_dff_B_aMV6Svoj8_0),.dout(w_dff_B_ejDlgELE4_0),.clk(gclk));
	jdff dff_B_GN0qANP52_0(.din(w_dff_B_ejDlgELE4_0),.dout(w_dff_B_GN0qANP52_0),.clk(gclk));
	jdff dff_B_c2Jq4dcx7_0(.din(w_dff_B_GN0qANP52_0),.dout(w_dff_B_c2Jq4dcx7_0),.clk(gclk));
	jdff dff_B_1BWEqvbk0_0(.din(w_dff_B_c2Jq4dcx7_0),.dout(w_dff_B_1BWEqvbk0_0),.clk(gclk));
	jdff dff_B_dWECNPgy9_0(.din(w_dff_B_1BWEqvbk0_0),.dout(w_dff_B_dWECNPgy9_0),.clk(gclk));
	jdff dff_B_rm5EmWSX5_0(.din(w_dff_B_dWECNPgy9_0),.dout(w_dff_B_rm5EmWSX5_0),.clk(gclk));
	jdff dff_B_x1BF1BUU3_0(.din(w_dff_B_rm5EmWSX5_0),.dout(w_dff_B_x1BF1BUU3_0),.clk(gclk));
	jdff dff_B_4D0e6DQI6_0(.din(w_dff_B_x1BF1BUU3_0),.dout(w_dff_B_4D0e6DQI6_0),.clk(gclk));
	jdff dff_B_PUUCstNx9_0(.din(w_dff_B_4D0e6DQI6_0),.dout(w_dff_B_PUUCstNx9_0),.clk(gclk));
	jdff dff_B_XA1RQxyR7_0(.din(w_dff_B_PUUCstNx9_0),.dout(w_dff_B_XA1RQxyR7_0),.clk(gclk));
	jdff dff_B_nAbfrSV09_0(.din(w_dff_B_XA1RQxyR7_0),.dout(w_dff_B_nAbfrSV09_0),.clk(gclk));
	jdff dff_B_Ab3IT7Dh2_0(.din(w_dff_B_nAbfrSV09_0),.dout(w_dff_B_Ab3IT7Dh2_0),.clk(gclk));
	jdff dff_B_o7WwTovS6_0(.din(w_dff_B_Ab3IT7Dh2_0),.dout(w_dff_B_o7WwTovS6_0),.clk(gclk));
	jdff dff_B_nYsULZsA3_0(.din(w_dff_B_o7WwTovS6_0),.dout(w_dff_B_nYsULZsA3_0),.clk(gclk));
	jdff dff_B_I3nbp6qU3_0(.din(w_dff_B_nYsULZsA3_0),.dout(w_dff_B_I3nbp6qU3_0),.clk(gclk));
	jdff dff_B_9biXOlce0_0(.din(w_dff_B_I3nbp6qU3_0),.dout(w_dff_B_9biXOlce0_0),.clk(gclk));
	jdff dff_B_jIivYryf8_0(.din(w_dff_B_9biXOlce0_0),.dout(w_dff_B_jIivYryf8_0),.clk(gclk));
	jdff dff_B_mwrykKhY9_0(.din(w_dff_B_jIivYryf8_0),.dout(w_dff_B_mwrykKhY9_0),.clk(gclk));
	jdff dff_B_OgruAIXJ9_0(.din(w_dff_B_mwrykKhY9_0),.dout(w_dff_B_OgruAIXJ9_0),.clk(gclk));
	jdff dff_B_YyVIEu8A4_0(.din(w_dff_B_OgruAIXJ9_0),.dout(w_dff_B_YyVIEu8A4_0),.clk(gclk));
	jdff dff_B_J4Tc4Nfx2_0(.din(w_dff_B_YyVIEu8A4_0),.dout(w_dff_B_J4Tc4Nfx2_0),.clk(gclk));
	jdff dff_B_puVG3F539_0(.din(w_dff_B_J4Tc4Nfx2_0),.dout(w_dff_B_puVG3F539_0),.clk(gclk));
	jdff dff_B_0OjSc4mg1_0(.din(w_dff_B_puVG3F539_0),.dout(w_dff_B_0OjSc4mg1_0),.clk(gclk));
	jdff dff_B_MUt2RQG45_0(.din(w_dff_B_0OjSc4mg1_0),.dout(w_dff_B_MUt2RQG45_0),.clk(gclk));
	jdff dff_B_1JLdUdCP3_0(.din(w_dff_B_MUt2RQG45_0),.dout(w_dff_B_1JLdUdCP3_0),.clk(gclk));
	jdff dff_B_o2WsywEg8_0(.din(w_dff_B_1JLdUdCP3_0),.dout(w_dff_B_o2WsywEg8_0),.clk(gclk));
	jdff dff_B_qDb9SBpR7_0(.din(w_dff_B_o2WsywEg8_0),.dout(w_dff_B_qDb9SBpR7_0),.clk(gclk));
	jdff dff_B_nRAWg75X2_0(.din(w_dff_B_qDb9SBpR7_0),.dout(w_dff_B_nRAWg75X2_0),.clk(gclk));
	jdff dff_B_muX7q6CO0_0(.din(w_dff_B_nRAWg75X2_0),.dout(w_dff_B_muX7q6CO0_0),.clk(gclk));
	jdff dff_B_JhrC8uVe4_0(.din(w_dff_B_muX7q6CO0_0),.dout(w_dff_B_JhrC8uVe4_0),.clk(gclk));
	jdff dff_B_QUTIphUX9_0(.din(w_dff_B_JhrC8uVe4_0),.dout(w_dff_B_QUTIphUX9_0),.clk(gclk));
	jdff dff_B_JrjXALgH0_0(.din(w_dff_B_QUTIphUX9_0),.dout(w_dff_B_JrjXALgH0_0),.clk(gclk));
	jdff dff_B_5Ov3MkWU4_0(.din(w_dff_B_JrjXALgH0_0),.dout(w_dff_B_5Ov3MkWU4_0),.clk(gclk));
	jdff dff_B_WOL3ufiO1_0(.din(w_dff_B_5Ov3MkWU4_0),.dout(w_dff_B_WOL3ufiO1_0),.clk(gclk));
	jdff dff_B_tWbNMCYe9_0(.din(w_dff_B_WOL3ufiO1_0),.dout(w_dff_B_tWbNMCYe9_0),.clk(gclk));
	jdff dff_B_RFIbUvxx2_0(.din(w_dff_B_tWbNMCYe9_0),.dout(w_dff_B_RFIbUvxx2_0),.clk(gclk));
	jdff dff_B_3fEKCzTR8_0(.din(w_dff_B_RFIbUvxx2_0),.dout(w_dff_B_3fEKCzTR8_0),.clk(gclk));
	jdff dff_B_pnxrMXfL6_0(.din(w_dff_B_3fEKCzTR8_0),.dout(w_dff_B_pnxrMXfL6_0),.clk(gclk));
	jdff dff_B_uUkfOFQn1_0(.din(w_dff_B_pnxrMXfL6_0),.dout(w_dff_B_uUkfOFQn1_0),.clk(gclk));
	jdff dff_B_QtSE2alq8_0(.din(n910),.dout(w_dff_B_QtSE2alq8_0),.clk(gclk));
	jdff dff_B_a60LwpbU0_0(.din(w_dff_B_QtSE2alq8_0),.dout(w_dff_B_a60LwpbU0_0),.clk(gclk));
	jdff dff_B_1xKJMbsb7_0(.din(w_dff_B_a60LwpbU0_0),.dout(w_dff_B_1xKJMbsb7_0),.clk(gclk));
	jdff dff_B_zyFmT5e05_0(.din(w_dff_B_1xKJMbsb7_0),.dout(w_dff_B_zyFmT5e05_0),.clk(gclk));
	jdff dff_B_p5DSkSea4_0(.din(w_dff_B_zyFmT5e05_0),.dout(w_dff_B_p5DSkSea4_0),.clk(gclk));
	jdff dff_B_OMwW1Zbs2_0(.din(w_dff_B_p5DSkSea4_0),.dout(w_dff_B_OMwW1Zbs2_0),.clk(gclk));
	jdff dff_B_7ean7UXY0_0(.din(w_dff_B_OMwW1Zbs2_0),.dout(w_dff_B_7ean7UXY0_0),.clk(gclk));
	jdff dff_B_oitKwxnb4_0(.din(w_dff_B_7ean7UXY0_0),.dout(w_dff_B_oitKwxnb4_0),.clk(gclk));
	jdff dff_B_PeXnXtj88_0(.din(w_dff_B_oitKwxnb4_0),.dout(w_dff_B_PeXnXtj88_0),.clk(gclk));
	jdff dff_B_t2TBwC2m4_0(.din(w_dff_B_PeXnXtj88_0),.dout(w_dff_B_t2TBwC2m4_0),.clk(gclk));
	jdff dff_B_xpfmd1fS5_0(.din(w_dff_B_t2TBwC2m4_0),.dout(w_dff_B_xpfmd1fS5_0),.clk(gclk));
	jdff dff_B_yiz34MsO2_0(.din(w_dff_B_xpfmd1fS5_0),.dout(w_dff_B_yiz34MsO2_0),.clk(gclk));
	jdff dff_B_aZrBtuQV7_0(.din(w_dff_B_yiz34MsO2_0),.dout(w_dff_B_aZrBtuQV7_0),.clk(gclk));
	jdff dff_B_hrLHjEyU9_0(.din(w_dff_B_aZrBtuQV7_0),.dout(w_dff_B_hrLHjEyU9_0),.clk(gclk));
	jdff dff_B_s3kqD9F70_0(.din(w_dff_B_hrLHjEyU9_0),.dout(w_dff_B_s3kqD9F70_0),.clk(gclk));
	jdff dff_B_MRPGm56t9_0(.din(w_dff_B_s3kqD9F70_0),.dout(w_dff_B_MRPGm56t9_0),.clk(gclk));
	jdff dff_B_idYSafC78_0(.din(w_dff_B_MRPGm56t9_0),.dout(w_dff_B_idYSafC78_0),.clk(gclk));
	jdff dff_B_mzo147uB9_0(.din(w_dff_B_idYSafC78_0),.dout(w_dff_B_mzo147uB9_0),.clk(gclk));
	jdff dff_B_wW80m5xJ7_0(.din(w_dff_B_mzo147uB9_0),.dout(w_dff_B_wW80m5xJ7_0),.clk(gclk));
	jdff dff_B_iX1elz686_0(.din(w_dff_B_wW80m5xJ7_0),.dout(w_dff_B_iX1elz686_0),.clk(gclk));
	jdff dff_B_XWi7Zoti3_0(.din(w_dff_B_iX1elz686_0),.dout(w_dff_B_XWi7Zoti3_0),.clk(gclk));
	jdff dff_B_9EyMk9Bx3_0(.din(w_dff_B_XWi7Zoti3_0),.dout(w_dff_B_9EyMk9Bx3_0),.clk(gclk));
	jdff dff_B_jg09GqFo7_0(.din(w_dff_B_9EyMk9Bx3_0),.dout(w_dff_B_jg09GqFo7_0),.clk(gclk));
	jdff dff_B_cXvUOrSZ5_0(.din(w_dff_B_jg09GqFo7_0),.dout(w_dff_B_cXvUOrSZ5_0),.clk(gclk));
	jdff dff_B_IiXRSKqj0_0(.din(w_dff_B_cXvUOrSZ5_0),.dout(w_dff_B_IiXRSKqj0_0),.clk(gclk));
	jdff dff_B_QaPpatWl3_0(.din(w_dff_B_IiXRSKqj0_0),.dout(w_dff_B_QaPpatWl3_0),.clk(gclk));
	jdff dff_B_gmU7MplD8_0(.din(w_dff_B_QaPpatWl3_0),.dout(w_dff_B_gmU7MplD8_0),.clk(gclk));
	jdff dff_B_FKgzxNck2_0(.din(w_dff_B_gmU7MplD8_0),.dout(w_dff_B_FKgzxNck2_0),.clk(gclk));
	jdff dff_B_iuRBEMsL8_0(.din(w_dff_B_FKgzxNck2_0),.dout(w_dff_B_iuRBEMsL8_0),.clk(gclk));
	jdff dff_B_zhWBGiw30_0(.din(w_dff_B_iuRBEMsL8_0),.dout(w_dff_B_zhWBGiw30_0),.clk(gclk));
	jdff dff_B_c16mnQyi5_0(.din(w_dff_B_zhWBGiw30_0),.dout(w_dff_B_c16mnQyi5_0),.clk(gclk));
	jdff dff_B_kZoiANpD2_0(.din(w_dff_B_c16mnQyi5_0),.dout(w_dff_B_kZoiANpD2_0),.clk(gclk));
	jdff dff_B_Ue9aPG913_0(.din(w_dff_B_kZoiANpD2_0),.dout(w_dff_B_Ue9aPG913_0),.clk(gclk));
	jdff dff_B_GxxhsJjw6_0(.din(w_dff_B_Ue9aPG913_0),.dout(w_dff_B_GxxhsJjw6_0),.clk(gclk));
	jdff dff_B_fviA1pj29_0(.din(w_dff_B_GxxhsJjw6_0),.dout(w_dff_B_fviA1pj29_0),.clk(gclk));
	jdff dff_B_0m1XsGUV5_0(.din(w_dff_B_fviA1pj29_0),.dout(w_dff_B_0m1XsGUV5_0),.clk(gclk));
	jdff dff_B_mFuzQE5A0_0(.din(w_dff_B_0m1XsGUV5_0),.dout(w_dff_B_mFuzQE5A0_0),.clk(gclk));
	jdff dff_B_yBF9yxPn5_0(.din(w_dff_B_mFuzQE5A0_0),.dout(w_dff_B_yBF9yxPn5_0),.clk(gclk));
	jdff dff_B_VOIcKW1j8_0(.din(w_dff_B_yBF9yxPn5_0),.dout(w_dff_B_VOIcKW1j8_0),.clk(gclk));
	jdff dff_B_SVgJJ2vo8_0(.din(w_dff_B_VOIcKW1j8_0),.dout(w_dff_B_SVgJJ2vo8_0),.clk(gclk));
	jdff dff_B_OeJl0nhT7_0(.din(w_dff_B_SVgJJ2vo8_0),.dout(w_dff_B_OeJl0nhT7_0),.clk(gclk));
	jdff dff_B_KBTawIzE0_0(.din(w_dff_B_OeJl0nhT7_0),.dout(w_dff_B_KBTawIzE0_0),.clk(gclk));
	jdff dff_B_pb8aXKb90_0(.din(w_dff_B_KBTawIzE0_0),.dout(w_dff_B_pb8aXKb90_0),.clk(gclk));
	jdff dff_B_0fImpkSC8_0(.din(w_dff_B_pb8aXKb90_0),.dout(w_dff_B_0fImpkSC8_0),.clk(gclk));
	jdff dff_B_Sq1RSOax7_0(.din(w_dff_B_0fImpkSC8_0),.dout(w_dff_B_Sq1RSOax7_0),.clk(gclk));
	jdff dff_B_iYF7zXYh2_0(.din(w_dff_B_Sq1RSOax7_0),.dout(w_dff_B_iYF7zXYh2_0),.clk(gclk));
	jdff dff_B_fl8zZlLZ3_0(.din(w_dff_B_iYF7zXYh2_0),.dout(w_dff_B_fl8zZlLZ3_0),.clk(gclk));
	jdff dff_B_cbmYB3cD6_0(.din(w_dff_B_fl8zZlLZ3_0),.dout(w_dff_B_cbmYB3cD6_0),.clk(gclk));
	jdff dff_B_JGvRZpqj5_0(.din(w_dff_B_cbmYB3cD6_0),.dout(w_dff_B_JGvRZpqj5_0),.clk(gclk));
	jdff dff_B_hrlz2aiW6_0(.din(w_dff_B_JGvRZpqj5_0),.dout(w_dff_B_hrlz2aiW6_0),.clk(gclk));
	jdff dff_B_h9Vbz6W55_0(.din(w_dff_B_hrlz2aiW6_0),.dout(w_dff_B_h9Vbz6W55_0),.clk(gclk));
	jdff dff_B_dmNLg6ON4_0(.din(w_dff_B_h9Vbz6W55_0),.dout(w_dff_B_dmNLg6ON4_0),.clk(gclk));
	jdff dff_B_DuZZPuLK1_0(.din(w_dff_B_dmNLg6ON4_0),.dout(w_dff_B_DuZZPuLK1_0),.clk(gclk));
	jdff dff_B_Cr0eBaQe4_0(.din(w_dff_B_DuZZPuLK1_0),.dout(w_dff_B_Cr0eBaQe4_0),.clk(gclk));
	jdff dff_B_4FSo0TXl9_0(.din(w_dff_B_Cr0eBaQe4_0),.dout(w_dff_B_4FSo0TXl9_0),.clk(gclk));
	jdff dff_B_3Vl08xmX6_0(.din(w_dff_B_4FSo0TXl9_0),.dout(w_dff_B_3Vl08xmX6_0),.clk(gclk));
	jdff dff_B_RGnPaSJw9_0(.din(w_dff_B_3Vl08xmX6_0),.dout(w_dff_B_RGnPaSJw9_0),.clk(gclk));
	jdff dff_B_7zZFrWzC0_0(.din(w_dff_B_RGnPaSJw9_0),.dout(w_dff_B_7zZFrWzC0_0),.clk(gclk));
	jdff dff_B_i0WlbGm57_0(.din(w_dff_B_7zZFrWzC0_0),.dout(w_dff_B_i0WlbGm57_0),.clk(gclk));
	jdff dff_B_AKFeOXCo2_0(.din(w_dff_B_i0WlbGm57_0),.dout(w_dff_B_AKFeOXCo2_0),.clk(gclk));
	jdff dff_B_rCV0ZODX8_0(.din(w_dff_B_AKFeOXCo2_0),.dout(w_dff_B_rCV0ZODX8_0),.clk(gclk));
	jdff dff_B_Y5tZFD296_0(.din(w_dff_B_rCV0ZODX8_0),.dout(w_dff_B_Y5tZFD296_0),.clk(gclk));
	jdff dff_B_dYkw7LMd5_0(.din(w_dff_B_Y5tZFD296_0),.dout(w_dff_B_dYkw7LMd5_0),.clk(gclk));
	jdff dff_B_79TJ03jF6_0(.din(w_dff_B_dYkw7LMd5_0),.dout(w_dff_B_79TJ03jF6_0),.clk(gclk));
	jdff dff_B_KoJVSAfr6_0(.din(w_dff_B_79TJ03jF6_0),.dout(w_dff_B_KoJVSAfr6_0),.clk(gclk));
	jdff dff_B_ninceOZA1_0(.din(w_dff_B_KoJVSAfr6_0),.dout(w_dff_B_ninceOZA1_0),.clk(gclk));
	jdff dff_B_ZLiEY06c5_0(.din(w_dff_B_ninceOZA1_0),.dout(w_dff_B_ZLiEY06c5_0),.clk(gclk));
	jdff dff_B_a0Wtax9k9_0(.din(w_dff_B_ZLiEY06c5_0),.dout(w_dff_B_a0Wtax9k9_0),.clk(gclk));
	jdff dff_B_KDAiu1qz2_0(.din(w_dff_B_a0Wtax9k9_0),.dout(w_dff_B_KDAiu1qz2_0),.clk(gclk));
	jdff dff_B_KvTUSNaz7_0(.din(w_dff_B_KDAiu1qz2_0),.dout(w_dff_B_KvTUSNaz7_0),.clk(gclk));
	jdff dff_B_x63XX1Ly6_0(.din(w_dff_B_KvTUSNaz7_0),.dout(w_dff_B_x63XX1Ly6_0),.clk(gclk));
	jdff dff_B_wbr0oOuf3_0(.din(w_dff_B_x63XX1Ly6_0),.dout(w_dff_B_wbr0oOuf3_0),.clk(gclk));
	jdff dff_B_87DRgOHA1_0(.din(w_dff_B_wbr0oOuf3_0),.dout(w_dff_B_87DRgOHA1_0),.clk(gclk));
	jdff dff_B_k8hJc1TX5_0(.din(w_dff_B_87DRgOHA1_0),.dout(w_dff_B_k8hJc1TX5_0),.clk(gclk));
	jdff dff_B_epM7xax95_0(.din(w_dff_B_k8hJc1TX5_0),.dout(w_dff_B_epM7xax95_0),.clk(gclk));
	jdff dff_B_IiYF23UO4_0(.din(w_dff_B_epM7xax95_0),.dout(w_dff_B_IiYF23UO4_0),.clk(gclk));
	jdff dff_B_w13Ku9pw9_0(.din(w_dff_B_IiYF23UO4_0),.dout(w_dff_B_w13Ku9pw9_0),.clk(gclk));
	jdff dff_B_nH9UmjbH6_0(.din(w_dff_B_w13Ku9pw9_0),.dout(w_dff_B_nH9UmjbH6_0),.clk(gclk));
	jdff dff_B_K5JydMTT7_0(.din(w_dff_B_nH9UmjbH6_0),.dout(w_dff_B_K5JydMTT7_0),.clk(gclk));
	jdff dff_B_QcRFm2ko6_0(.din(w_dff_B_K5JydMTT7_0),.dout(w_dff_B_QcRFm2ko6_0),.clk(gclk));
	jdff dff_B_OZsDaZDK5_0(.din(w_dff_B_QcRFm2ko6_0),.dout(w_dff_B_OZsDaZDK5_0),.clk(gclk));
	jdff dff_B_krgSRuj05_0(.din(w_dff_B_OZsDaZDK5_0),.dout(w_dff_B_krgSRuj05_0),.clk(gclk));
	jdff dff_B_VUY6y9pD5_0(.din(w_dff_B_krgSRuj05_0),.dout(w_dff_B_VUY6y9pD5_0),.clk(gclk));
	jdff dff_B_ifKdVjtU2_0(.din(w_dff_B_VUY6y9pD5_0),.dout(w_dff_B_ifKdVjtU2_0),.clk(gclk));
	jdff dff_B_YsAFealH2_0(.din(w_dff_B_ifKdVjtU2_0),.dout(w_dff_B_YsAFealH2_0),.clk(gclk));
	jdff dff_B_erm8ltah9_0(.din(w_dff_B_YsAFealH2_0),.dout(w_dff_B_erm8ltah9_0),.clk(gclk));
	jdff dff_B_ynh2rDWK5_0(.din(w_dff_B_erm8ltah9_0),.dout(w_dff_B_ynh2rDWK5_0),.clk(gclk));
	jdff dff_B_teUIUmXN2_0(.din(n916),.dout(w_dff_B_teUIUmXN2_0),.clk(gclk));
	jdff dff_B_36Nr5e4v0_0(.din(w_dff_B_teUIUmXN2_0),.dout(w_dff_B_36Nr5e4v0_0),.clk(gclk));
	jdff dff_B_evYzW6yN9_0(.din(w_dff_B_36Nr5e4v0_0),.dout(w_dff_B_evYzW6yN9_0),.clk(gclk));
	jdff dff_B_A2EaiSLS2_0(.din(w_dff_B_evYzW6yN9_0),.dout(w_dff_B_A2EaiSLS2_0),.clk(gclk));
	jdff dff_B_3WES9sEE4_0(.din(w_dff_B_A2EaiSLS2_0),.dout(w_dff_B_3WES9sEE4_0),.clk(gclk));
	jdff dff_B_i8VZmfPt2_0(.din(w_dff_B_3WES9sEE4_0),.dout(w_dff_B_i8VZmfPt2_0),.clk(gclk));
	jdff dff_B_VAXZtPOg8_0(.din(w_dff_B_i8VZmfPt2_0),.dout(w_dff_B_VAXZtPOg8_0),.clk(gclk));
	jdff dff_B_Q0AGl5hU8_0(.din(w_dff_B_VAXZtPOg8_0),.dout(w_dff_B_Q0AGl5hU8_0),.clk(gclk));
	jdff dff_B_dckM39du9_0(.din(w_dff_B_Q0AGl5hU8_0),.dout(w_dff_B_dckM39du9_0),.clk(gclk));
	jdff dff_B_IzjaZ1XN1_0(.din(w_dff_B_dckM39du9_0),.dout(w_dff_B_IzjaZ1XN1_0),.clk(gclk));
	jdff dff_B_rJRZKPlQ9_0(.din(w_dff_B_IzjaZ1XN1_0),.dout(w_dff_B_rJRZKPlQ9_0),.clk(gclk));
	jdff dff_B_ZJ7IgyKt1_0(.din(w_dff_B_rJRZKPlQ9_0),.dout(w_dff_B_ZJ7IgyKt1_0),.clk(gclk));
	jdff dff_B_GLeXHGI72_0(.din(w_dff_B_ZJ7IgyKt1_0),.dout(w_dff_B_GLeXHGI72_0),.clk(gclk));
	jdff dff_B_8orOh9oT4_0(.din(w_dff_B_GLeXHGI72_0),.dout(w_dff_B_8orOh9oT4_0),.clk(gclk));
	jdff dff_B_DCVvUxlg7_0(.din(w_dff_B_8orOh9oT4_0),.dout(w_dff_B_DCVvUxlg7_0),.clk(gclk));
	jdff dff_B_zfvIZB2u3_0(.din(w_dff_B_DCVvUxlg7_0),.dout(w_dff_B_zfvIZB2u3_0),.clk(gclk));
	jdff dff_B_alLn5dug9_0(.din(w_dff_B_zfvIZB2u3_0),.dout(w_dff_B_alLn5dug9_0),.clk(gclk));
	jdff dff_B_fNKQ5FxJ5_0(.din(w_dff_B_alLn5dug9_0),.dout(w_dff_B_fNKQ5FxJ5_0),.clk(gclk));
	jdff dff_B_zIFcmTRN6_0(.din(w_dff_B_fNKQ5FxJ5_0),.dout(w_dff_B_zIFcmTRN6_0),.clk(gclk));
	jdff dff_B_dIAPTpEE3_0(.din(w_dff_B_zIFcmTRN6_0),.dout(w_dff_B_dIAPTpEE3_0),.clk(gclk));
	jdff dff_B_SvocjBtu9_0(.din(w_dff_B_dIAPTpEE3_0),.dout(w_dff_B_SvocjBtu9_0),.clk(gclk));
	jdff dff_B_5XM7lrJ18_0(.din(w_dff_B_SvocjBtu9_0),.dout(w_dff_B_5XM7lrJ18_0),.clk(gclk));
	jdff dff_B_AvvWnsEE4_0(.din(w_dff_B_5XM7lrJ18_0),.dout(w_dff_B_AvvWnsEE4_0),.clk(gclk));
	jdff dff_B_LDPSWqN55_0(.din(w_dff_B_AvvWnsEE4_0),.dout(w_dff_B_LDPSWqN55_0),.clk(gclk));
	jdff dff_B_Ne51fv8f4_0(.din(w_dff_B_LDPSWqN55_0),.dout(w_dff_B_Ne51fv8f4_0),.clk(gclk));
	jdff dff_B_tiZ4KHiW2_0(.din(w_dff_B_Ne51fv8f4_0),.dout(w_dff_B_tiZ4KHiW2_0),.clk(gclk));
	jdff dff_B_I2jlKbNp8_0(.din(w_dff_B_tiZ4KHiW2_0),.dout(w_dff_B_I2jlKbNp8_0),.clk(gclk));
	jdff dff_B_cNBkCEVi1_0(.din(w_dff_B_I2jlKbNp8_0),.dout(w_dff_B_cNBkCEVi1_0),.clk(gclk));
	jdff dff_B_NQ03wBgH1_0(.din(w_dff_B_cNBkCEVi1_0),.dout(w_dff_B_NQ03wBgH1_0),.clk(gclk));
	jdff dff_B_Hlu0yAFh2_0(.din(w_dff_B_NQ03wBgH1_0),.dout(w_dff_B_Hlu0yAFh2_0),.clk(gclk));
	jdff dff_B_9fjo0r898_0(.din(w_dff_B_Hlu0yAFh2_0),.dout(w_dff_B_9fjo0r898_0),.clk(gclk));
	jdff dff_B_UJWMk3Z27_0(.din(w_dff_B_9fjo0r898_0),.dout(w_dff_B_UJWMk3Z27_0),.clk(gclk));
	jdff dff_B_euGD2qB86_0(.din(w_dff_B_UJWMk3Z27_0),.dout(w_dff_B_euGD2qB86_0),.clk(gclk));
	jdff dff_B_fjNKgvcU9_0(.din(w_dff_B_euGD2qB86_0),.dout(w_dff_B_fjNKgvcU9_0),.clk(gclk));
	jdff dff_B_4Vqi2sXR0_0(.din(w_dff_B_fjNKgvcU9_0),.dout(w_dff_B_4Vqi2sXR0_0),.clk(gclk));
	jdff dff_B_EyBF3q6K5_0(.din(w_dff_B_4Vqi2sXR0_0),.dout(w_dff_B_EyBF3q6K5_0),.clk(gclk));
	jdff dff_B_0JLHOIUQ5_0(.din(w_dff_B_EyBF3q6K5_0),.dout(w_dff_B_0JLHOIUQ5_0),.clk(gclk));
	jdff dff_B_PA6TGe5t5_0(.din(w_dff_B_0JLHOIUQ5_0),.dout(w_dff_B_PA6TGe5t5_0),.clk(gclk));
	jdff dff_B_LnVF8d2f1_0(.din(w_dff_B_PA6TGe5t5_0),.dout(w_dff_B_LnVF8d2f1_0),.clk(gclk));
	jdff dff_B_aPbt9GGI7_0(.din(w_dff_B_LnVF8d2f1_0),.dout(w_dff_B_aPbt9GGI7_0),.clk(gclk));
	jdff dff_B_7vk1Ogy88_0(.din(w_dff_B_aPbt9GGI7_0),.dout(w_dff_B_7vk1Ogy88_0),.clk(gclk));
	jdff dff_B_ZrbQErD96_0(.din(w_dff_B_7vk1Ogy88_0),.dout(w_dff_B_ZrbQErD96_0),.clk(gclk));
	jdff dff_B_QlkWJsah4_0(.din(w_dff_B_ZrbQErD96_0),.dout(w_dff_B_QlkWJsah4_0),.clk(gclk));
	jdff dff_B_BZuEnWnu4_0(.din(w_dff_B_QlkWJsah4_0),.dout(w_dff_B_BZuEnWnu4_0),.clk(gclk));
	jdff dff_B_QYwB1byA3_0(.din(w_dff_B_BZuEnWnu4_0),.dout(w_dff_B_QYwB1byA3_0),.clk(gclk));
	jdff dff_B_6csUr0Hr4_0(.din(w_dff_B_QYwB1byA3_0),.dout(w_dff_B_6csUr0Hr4_0),.clk(gclk));
	jdff dff_B_RA6pGNX62_0(.din(w_dff_B_6csUr0Hr4_0),.dout(w_dff_B_RA6pGNX62_0),.clk(gclk));
	jdff dff_B_hdIg99Ys2_0(.din(w_dff_B_RA6pGNX62_0),.dout(w_dff_B_hdIg99Ys2_0),.clk(gclk));
	jdff dff_B_l42FmOb26_0(.din(w_dff_B_hdIg99Ys2_0),.dout(w_dff_B_l42FmOb26_0),.clk(gclk));
	jdff dff_B_nE6sKC2a9_0(.din(w_dff_B_l42FmOb26_0),.dout(w_dff_B_nE6sKC2a9_0),.clk(gclk));
	jdff dff_B_cXEgdtn60_0(.din(w_dff_B_nE6sKC2a9_0),.dout(w_dff_B_cXEgdtn60_0),.clk(gclk));
	jdff dff_B_xrPnkjAD4_0(.din(w_dff_B_cXEgdtn60_0),.dout(w_dff_B_xrPnkjAD4_0),.clk(gclk));
	jdff dff_B_NyMCjCYC9_0(.din(w_dff_B_xrPnkjAD4_0),.dout(w_dff_B_NyMCjCYC9_0),.clk(gclk));
	jdff dff_B_FQKpehzb2_0(.din(w_dff_B_NyMCjCYC9_0),.dout(w_dff_B_FQKpehzb2_0),.clk(gclk));
	jdff dff_B_0lyI64ZE3_0(.din(w_dff_B_FQKpehzb2_0),.dout(w_dff_B_0lyI64ZE3_0),.clk(gclk));
	jdff dff_B_DVswJc5Z6_0(.din(w_dff_B_0lyI64ZE3_0),.dout(w_dff_B_DVswJc5Z6_0),.clk(gclk));
	jdff dff_B_BSKY3utX3_0(.din(w_dff_B_DVswJc5Z6_0),.dout(w_dff_B_BSKY3utX3_0),.clk(gclk));
	jdff dff_B_K9SkFrZw4_0(.din(w_dff_B_BSKY3utX3_0),.dout(w_dff_B_K9SkFrZw4_0),.clk(gclk));
	jdff dff_B_MCHK6wHv1_0(.din(w_dff_B_K9SkFrZw4_0),.dout(w_dff_B_MCHK6wHv1_0),.clk(gclk));
	jdff dff_B_PQbkRS7H2_0(.din(w_dff_B_MCHK6wHv1_0),.dout(w_dff_B_PQbkRS7H2_0),.clk(gclk));
	jdff dff_B_52sZSUvo4_0(.din(w_dff_B_PQbkRS7H2_0),.dout(w_dff_B_52sZSUvo4_0),.clk(gclk));
	jdff dff_B_679TxmNw3_0(.din(w_dff_B_52sZSUvo4_0),.dout(w_dff_B_679TxmNw3_0),.clk(gclk));
	jdff dff_B_h2KF3RLB3_0(.din(w_dff_B_679TxmNw3_0),.dout(w_dff_B_h2KF3RLB3_0),.clk(gclk));
	jdff dff_B_ILY51LBP4_0(.din(w_dff_B_h2KF3RLB3_0),.dout(w_dff_B_ILY51LBP4_0),.clk(gclk));
	jdff dff_B_cs6IY91D8_0(.din(w_dff_B_ILY51LBP4_0),.dout(w_dff_B_cs6IY91D8_0),.clk(gclk));
	jdff dff_B_qFtykAGp8_0(.din(w_dff_B_cs6IY91D8_0),.dout(w_dff_B_qFtykAGp8_0),.clk(gclk));
	jdff dff_B_knLqfLUQ0_0(.din(w_dff_B_qFtykAGp8_0),.dout(w_dff_B_knLqfLUQ0_0),.clk(gclk));
	jdff dff_B_lvEXTfsp2_0(.din(w_dff_B_knLqfLUQ0_0),.dout(w_dff_B_lvEXTfsp2_0),.clk(gclk));
	jdff dff_B_G4Gr10HC0_0(.din(w_dff_B_lvEXTfsp2_0),.dout(w_dff_B_G4Gr10HC0_0),.clk(gclk));
	jdff dff_B_vQpZ6Imv8_0(.din(w_dff_B_G4Gr10HC0_0),.dout(w_dff_B_vQpZ6Imv8_0),.clk(gclk));
	jdff dff_B_zlbjkOeu8_0(.din(w_dff_B_vQpZ6Imv8_0),.dout(w_dff_B_zlbjkOeu8_0),.clk(gclk));
	jdff dff_B_hAxxrdp33_0(.din(w_dff_B_zlbjkOeu8_0),.dout(w_dff_B_hAxxrdp33_0),.clk(gclk));
	jdff dff_B_Xe44QXIQ1_0(.din(w_dff_B_hAxxrdp33_0),.dout(w_dff_B_Xe44QXIQ1_0),.clk(gclk));
	jdff dff_B_JthLW1dC9_0(.din(w_dff_B_Xe44QXIQ1_0),.dout(w_dff_B_JthLW1dC9_0),.clk(gclk));
	jdff dff_B_AfVvE9ms4_0(.din(w_dff_B_JthLW1dC9_0),.dout(w_dff_B_AfVvE9ms4_0),.clk(gclk));
	jdff dff_B_yQndL1I96_0(.din(w_dff_B_AfVvE9ms4_0),.dout(w_dff_B_yQndL1I96_0),.clk(gclk));
	jdff dff_B_ZQpNBVcN9_0(.din(w_dff_B_yQndL1I96_0),.dout(w_dff_B_ZQpNBVcN9_0),.clk(gclk));
	jdff dff_B_yhlUcBIH5_0(.din(w_dff_B_ZQpNBVcN9_0),.dout(w_dff_B_yhlUcBIH5_0),.clk(gclk));
	jdff dff_B_CPhFAnYN7_0(.din(w_dff_B_yhlUcBIH5_0),.dout(w_dff_B_CPhFAnYN7_0),.clk(gclk));
	jdff dff_B_lbTHRrQO6_0(.din(w_dff_B_CPhFAnYN7_0),.dout(w_dff_B_lbTHRrQO6_0),.clk(gclk));
	jdff dff_B_Mx8h8HwG9_0(.din(w_dff_B_lbTHRrQO6_0),.dout(w_dff_B_Mx8h8HwG9_0),.clk(gclk));
	jdff dff_B_yZr8mdDz5_0(.din(w_dff_B_Mx8h8HwG9_0),.dout(w_dff_B_yZr8mdDz5_0),.clk(gclk));
	jdff dff_B_zsTH0Awc5_0(.din(w_dff_B_yZr8mdDz5_0),.dout(w_dff_B_zsTH0Awc5_0),.clk(gclk));
	jdff dff_B_miPfl8T48_0(.din(w_dff_B_zsTH0Awc5_0),.dout(w_dff_B_miPfl8T48_0),.clk(gclk));
	jdff dff_B_WoAWFxgM3_0(.din(w_dff_B_miPfl8T48_0),.dout(w_dff_B_WoAWFxgM3_0),.clk(gclk));
	jdff dff_B_sXDzow1e0_0(.din(w_dff_B_WoAWFxgM3_0),.dout(w_dff_B_sXDzow1e0_0),.clk(gclk));
	jdff dff_B_Yo2B737v3_0(.din(w_dff_B_sXDzow1e0_0),.dout(w_dff_B_Yo2B737v3_0),.clk(gclk));
	jdff dff_B_HLQWv4eU2_0(.din(w_dff_B_Yo2B737v3_0),.dout(w_dff_B_HLQWv4eU2_0),.clk(gclk));
	jdff dff_B_o6xCwdXu5_0(.din(n922),.dout(w_dff_B_o6xCwdXu5_0),.clk(gclk));
	jdff dff_B_tc3u8w468_0(.din(w_dff_B_o6xCwdXu5_0),.dout(w_dff_B_tc3u8w468_0),.clk(gclk));
	jdff dff_B_14EdoGIE1_0(.din(w_dff_B_tc3u8w468_0),.dout(w_dff_B_14EdoGIE1_0),.clk(gclk));
	jdff dff_B_ykoox14D0_0(.din(w_dff_B_14EdoGIE1_0),.dout(w_dff_B_ykoox14D0_0),.clk(gclk));
	jdff dff_B_V7sInmd47_0(.din(w_dff_B_ykoox14D0_0),.dout(w_dff_B_V7sInmd47_0),.clk(gclk));
	jdff dff_B_jNfKLFXS1_0(.din(w_dff_B_V7sInmd47_0),.dout(w_dff_B_jNfKLFXS1_0),.clk(gclk));
	jdff dff_B_mWjTHgVh6_0(.din(w_dff_B_jNfKLFXS1_0),.dout(w_dff_B_mWjTHgVh6_0),.clk(gclk));
	jdff dff_B_f7Ele7RO9_0(.din(w_dff_B_mWjTHgVh6_0),.dout(w_dff_B_f7Ele7RO9_0),.clk(gclk));
	jdff dff_B_piWs9FDx6_0(.din(w_dff_B_f7Ele7RO9_0),.dout(w_dff_B_piWs9FDx6_0),.clk(gclk));
	jdff dff_B_XoVzFCJj4_0(.din(w_dff_B_piWs9FDx6_0),.dout(w_dff_B_XoVzFCJj4_0),.clk(gclk));
	jdff dff_B_fLGqLtS47_0(.din(w_dff_B_XoVzFCJj4_0),.dout(w_dff_B_fLGqLtS47_0),.clk(gclk));
	jdff dff_B_Hqg8jK0B1_0(.din(w_dff_B_fLGqLtS47_0),.dout(w_dff_B_Hqg8jK0B1_0),.clk(gclk));
	jdff dff_B_vqnhZzCs2_0(.din(w_dff_B_Hqg8jK0B1_0),.dout(w_dff_B_vqnhZzCs2_0),.clk(gclk));
	jdff dff_B_E8l6wy0I3_0(.din(w_dff_B_vqnhZzCs2_0),.dout(w_dff_B_E8l6wy0I3_0),.clk(gclk));
	jdff dff_B_dvqeaSij1_0(.din(w_dff_B_E8l6wy0I3_0),.dout(w_dff_B_dvqeaSij1_0),.clk(gclk));
	jdff dff_B_wl7LBGnw1_0(.din(w_dff_B_dvqeaSij1_0),.dout(w_dff_B_wl7LBGnw1_0),.clk(gclk));
	jdff dff_B_GYR9jce80_0(.din(w_dff_B_wl7LBGnw1_0),.dout(w_dff_B_GYR9jce80_0),.clk(gclk));
	jdff dff_B_zuqBaa1S9_0(.din(w_dff_B_GYR9jce80_0),.dout(w_dff_B_zuqBaa1S9_0),.clk(gclk));
	jdff dff_B_FJzbmHpf0_0(.din(w_dff_B_zuqBaa1S9_0),.dout(w_dff_B_FJzbmHpf0_0),.clk(gclk));
	jdff dff_B_FvAWsfAE8_0(.din(w_dff_B_FJzbmHpf0_0),.dout(w_dff_B_FvAWsfAE8_0),.clk(gclk));
	jdff dff_B_tVs9R9vG9_0(.din(w_dff_B_FvAWsfAE8_0),.dout(w_dff_B_tVs9R9vG9_0),.clk(gclk));
	jdff dff_B_svSuWFHX8_0(.din(w_dff_B_tVs9R9vG9_0),.dout(w_dff_B_svSuWFHX8_0),.clk(gclk));
	jdff dff_B_DDPQKyId7_0(.din(w_dff_B_svSuWFHX8_0),.dout(w_dff_B_DDPQKyId7_0),.clk(gclk));
	jdff dff_B_wwokALGe8_0(.din(w_dff_B_DDPQKyId7_0),.dout(w_dff_B_wwokALGe8_0),.clk(gclk));
	jdff dff_B_yrfvQdy76_0(.din(w_dff_B_wwokALGe8_0),.dout(w_dff_B_yrfvQdy76_0),.clk(gclk));
	jdff dff_B_pDVPPZn74_0(.din(w_dff_B_yrfvQdy76_0),.dout(w_dff_B_pDVPPZn74_0),.clk(gclk));
	jdff dff_B_LCgeEXT91_0(.din(w_dff_B_pDVPPZn74_0),.dout(w_dff_B_LCgeEXT91_0),.clk(gclk));
	jdff dff_B_mTHEaqJk3_0(.din(w_dff_B_LCgeEXT91_0),.dout(w_dff_B_mTHEaqJk3_0),.clk(gclk));
	jdff dff_B_5tLVq2XS7_0(.din(w_dff_B_mTHEaqJk3_0),.dout(w_dff_B_5tLVq2XS7_0),.clk(gclk));
	jdff dff_B_Bb3m5DC66_0(.din(w_dff_B_5tLVq2XS7_0),.dout(w_dff_B_Bb3m5DC66_0),.clk(gclk));
	jdff dff_B_PKeVa7sH0_0(.din(w_dff_B_Bb3m5DC66_0),.dout(w_dff_B_PKeVa7sH0_0),.clk(gclk));
	jdff dff_B_zmvkgoz16_0(.din(w_dff_B_PKeVa7sH0_0),.dout(w_dff_B_zmvkgoz16_0),.clk(gclk));
	jdff dff_B_xLHrsSlh6_0(.din(w_dff_B_zmvkgoz16_0),.dout(w_dff_B_xLHrsSlh6_0),.clk(gclk));
	jdff dff_B_ZXpFUhLT6_0(.din(w_dff_B_xLHrsSlh6_0),.dout(w_dff_B_ZXpFUhLT6_0),.clk(gclk));
	jdff dff_B_Ao1UVAxz4_0(.din(w_dff_B_ZXpFUhLT6_0),.dout(w_dff_B_Ao1UVAxz4_0),.clk(gclk));
	jdff dff_B_u3YMuD0w7_0(.din(w_dff_B_Ao1UVAxz4_0),.dout(w_dff_B_u3YMuD0w7_0),.clk(gclk));
	jdff dff_B_TJU8CB1K9_0(.din(w_dff_B_u3YMuD0w7_0),.dout(w_dff_B_TJU8CB1K9_0),.clk(gclk));
	jdff dff_B_PJvjguEn8_0(.din(w_dff_B_TJU8CB1K9_0),.dout(w_dff_B_PJvjguEn8_0),.clk(gclk));
	jdff dff_B_xopPfgnR5_0(.din(w_dff_B_PJvjguEn8_0),.dout(w_dff_B_xopPfgnR5_0),.clk(gclk));
	jdff dff_B_3fx4ymWY5_0(.din(w_dff_B_xopPfgnR5_0),.dout(w_dff_B_3fx4ymWY5_0),.clk(gclk));
	jdff dff_B_ZbCqZhea4_0(.din(w_dff_B_3fx4ymWY5_0),.dout(w_dff_B_ZbCqZhea4_0),.clk(gclk));
	jdff dff_B_I8HSUCXM1_0(.din(w_dff_B_ZbCqZhea4_0),.dout(w_dff_B_I8HSUCXM1_0),.clk(gclk));
	jdff dff_B_vuPeDlkB9_0(.din(w_dff_B_I8HSUCXM1_0),.dout(w_dff_B_vuPeDlkB9_0),.clk(gclk));
	jdff dff_B_QIQQwm6M6_0(.din(w_dff_B_vuPeDlkB9_0),.dout(w_dff_B_QIQQwm6M6_0),.clk(gclk));
	jdff dff_B_3UBzza6x6_0(.din(w_dff_B_QIQQwm6M6_0),.dout(w_dff_B_3UBzza6x6_0),.clk(gclk));
	jdff dff_B_RorxNhg46_0(.din(w_dff_B_3UBzza6x6_0),.dout(w_dff_B_RorxNhg46_0),.clk(gclk));
	jdff dff_B_rr3m3kMy9_0(.din(w_dff_B_RorxNhg46_0),.dout(w_dff_B_rr3m3kMy9_0),.clk(gclk));
	jdff dff_B_u6N0CKnZ2_0(.din(w_dff_B_rr3m3kMy9_0),.dout(w_dff_B_u6N0CKnZ2_0),.clk(gclk));
	jdff dff_B_I200MfGu1_0(.din(w_dff_B_u6N0CKnZ2_0),.dout(w_dff_B_I200MfGu1_0),.clk(gclk));
	jdff dff_B_UnW3HPIw5_0(.din(w_dff_B_I200MfGu1_0),.dout(w_dff_B_UnW3HPIw5_0),.clk(gclk));
	jdff dff_B_7x7R4RIK4_0(.din(w_dff_B_UnW3HPIw5_0),.dout(w_dff_B_7x7R4RIK4_0),.clk(gclk));
	jdff dff_B_zj3vQalB8_0(.din(w_dff_B_7x7R4RIK4_0),.dout(w_dff_B_zj3vQalB8_0),.clk(gclk));
	jdff dff_B_CaCXwbVA0_0(.din(w_dff_B_zj3vQalB8_0),.dout(w_dff_B_CaCXwbVA0_0),.clk(gclk));
	jdff dff_B_KjEFd3Tr2_0(.din(w_dff_B_CaCXwbVA0_0),.dout(w_dff_B_KjEFd3Tr2_0),.clk(gclk));
	jdff dff_B_eoRU2Dig8_0(.din(w_dff_B_KjEFd3Tr2_0),.dout(w_dff_B_eoRU2Dig8_0),.clk(gclk));
	jdff dff_B_XF4TZrF18_0(.din(w_dff_B_eoRU2Dig8_0),.dout(w_dff_B_XF4TZrF18_0),.clk(gclk));
	jdff dff_B_kFIBnhRV3_0(.din(w_dff_B_XF4TZrF18_0),.dout(w_dff_B_kFIBnhRV3_0),.clk(gclk));
	jdff dff_B_bsb7w8Ld0_0(.din(w_dff_B_kFIBnhRV3_0),.dout(w_dff_B_bsb7w8Ld0_0),.clk(gclk));
	jdff dff_B_BHGtaNg47_0(.din(w_dff_B_bsb7w8Ld0_0),.dout(w_dff_B_BHGtaNg47_0),.clk(gclk));
	jdff dff_B_ENYkbVwg8_0(.din(w_dff_B_BHGtaNg47_0),.dout(w_dff_B_ENYkbVwg8_0),.clk(gclk));
	jdff dff_B_yippQWKC3_0(.din(w_dff_B_ENYkbVwg8_0),.dout(w_dff_B_yippQWKC3_0),.clk(gclk));
	jdff dff_B_vnYCDvKi3_0(.din(w_dff_B_yippQWKC3_0),.dout(w_dff_B_vnYCDvKi3_0),.clk(gclk));
	jdff dff_B_WxKeVE7v8_0(.din(w_dff_B_vnYCDvKi3_0),.dout(w_dff_B_WxKeVE7v8_0),.clk(gclk));
	jdff dff_B_0UN5UyyP6_0(.din(w_dff_B_WxKeVE7v8_0),.dout(w_dff_B_0UN5UyyP6_0),.clk(gclk));
	jdff dff_B_6h4QR3wu1_0(.din(w_dff_B_0UN5UyyP6_0),.dout(w_dff_B_6h4QR3wu1_0),.clk(gclk));
	jdff dff_B_mzldZlCK9_0(.din(w_dff_B_6h4QR3wu1_0),.dout(w_dff_B_mzldZlCK9_0),.clk(gclk));
	jdff dff_B_CjJInOFP4_0(.din(w_dff_B_mzldZlCK9_0),.dout(w_dff_B_CjJInOFP4_0),.clk(gclk));
	jdff dff_B_tg9dYumo2_0(.din(w_dff_B_CjJInOFP4_0),.dout(w_dff_B_tg9dYumo2_0),.clk(gclk));
	jdff dff_B_atYxgtNA9_0(.din(w_dff_B_tg9dYumo2_0),.dout(w_dff_B_atYxgtNA9_0),.clk(gclk));
	jdff dff_B_ZBWtA7WT3_0(.din(w_dff_B_atYxgtNA9_0),.dout(w_dff_B_ZBWtA7WT3_0),.clk(gclk));
	jdff dff_B_llTlEFUM4_0(.din(w_dff_B_ZBWtA7WT3_0),.dout(w_dff_B_llTlEFUM4_0),.clk(gclk));
	jdff dff_B_JFgWisLP9_0(.din(w_dff_B_llTlEFUM4_0),.dout(w_dff_B_JFgWisLP9_0),.clk(gclk));
	jdff dff_B_WnrB3uOv4_0(.din(w_dff_B_JFgWisLP9_0),.dout(w_dff_B_WnrB3uOv4_0),.clk(gclk));
	jdff dff_B_xl5GkG4S3_0(.din(w_dff_B_WnrB3uOv4_0),.dout(w_dff_B_xl5GkG4S3_0),.clk(gclk));
	jdff dff_B_evmwPmZp5_0(.din(w_dff_B_xl5GkG4S3_0),.dout(w_dff_B_evmwPmZp5_0),.clk(gclk));
	jdff dff_B_9v14hgE90_0(.din(w_dff_B_evmwPmZp5_0),.dout(w_dff_B_9v14hgE90_0),.clk(gclk));
	jdff dff_B_Vws8LjOK8_0(.din(w_dff_B_9v14hgE90_0),.dout(w_dff_B_Vws8LjOK8_0),.clk(gclk));
	jdff dff_B_5rb1BXV10_0(.din(w_dff_B_Vws8LjOK8_0),.dout(w_dff_B_5rb1BXV10_0),.clk(gclk));
	jdff dff_B_nKYOxuLI3_0(.din(w_dff_B_5rb1BXV10_0),.dout(w_dff_B_nKYOxuLI3_0),.clk(gclk));
	jdff dff_B_mecQYNlA7_0(.din(w_dff_B_nKYOxuLI3_0),.dout(w_dff_B_mecQYNlA7_0),.clk(gclk));
	jdff dff_B_RCFoAGTf5_0(.din(w_dff_B_mecQYNlA7_0),.dout(w_dff_B_RCFoAGTf5_0),.clk(gclk));
	jdff dff_B_hDJREAJx5_0(.din(w_dff_B_RCFoAGTf5_0),.dout(w_dff_B_hDJREAJx5_0),.clk(gclk));
	jdff dff_B_ogBL6tSm1_0(.din(w_dff_B_hDJREAJx5_0),.dout(w_dff_B_ogBL6tSm1_0),.clk(gclk));
	jdff dff_B_3Lz9qtbN5_0(.din(w_dff_B_ogBL6tSm1_0),.dout(w_dff_B_3Lz9qtbN5_0),.clk(gclk));
	jdff dff_B_rtfxgeGM8_0(.din(w_dff_B_3Lz9qtbN5_0),.dout(w_dff_B_rtfxgeGM8_0),.clk(gclk));
	jdff dff_B_0AH7p5RH7_0(.din(w_dff_B_rtfxgeGM8_0),.dout(w_dff_B_0AH7p5RH7_0),.clk(gclk));
	jdff dff_B_4x8jDMf12_0(.din(w_dff_B_0AH7p5RH7_0),.dout(w_dff_B_4x8jDMf12_0),.clk(gclk));
	jdff dff_B_hUNL9Unj1_0(.din(w_dff_B_4x8jDMf12_0),.dout(w_dff_B_hUNL9Unj1_0),.clk(gclk));
	jdff dff_B_jeAaxdpn6_0(.din(w_dff_B_hUNL9Unj1_0),.dout(w_dff_B_jeAaxdpn6_0),.clk(gclk));
	jdff dff_B_74tiN2Vz8_0(.din(n928),.dout(w_dff_B_74tiN2Vz8_0),.clk(gclk));
	jdff dff_B_krFHa4VO1_0(.din(w_dff_B_74tiN2Vz8_0),.dout(w_dff_B_krFHa4VO1_0),.clk(gclk));
	jdff dff_B_l5MegGRP7_0(.din(w_dff_B_krFHa4VO1_0),.dout(w_dff_B_l5MegGRP7_0),.clk(gclk));
	jdff dff_B_SvCz5SVf1_0(.din(w_dff_B_l5MegGRP7_0),.dout(w_dff_B_SvCz5SVf1_0),.clk(gclk));
	jdff dff_B_Ns6paOb38_0(.din(w_dff_B_SvCz5SVf1_0),.dout(w_dff_B_Ns6paOb38_0),.clk(gclk));
	jdff dff_B_Mz12lt6A9_0(.din(w_dff_B_Ns6paOb38_0),.dout(w_dff_B_Mz12lt6A9_0),.clk(gclk));
	jdff dff_B_RMoNROTT9_0(.din(w_dff_B_Mz12lt6A9_0),.dout(w_dff_B_RMoNROTT9_0),.clk(gclk));
	jdff dff_B_v0WrVMHE7_0(.din(w_dff_B_RMoNROTT9_0),.dout(w_dff_B_v0WrVMHE7_0),.clk(gclk));
	jdff dff_B_xb3SG3cp0_0(.din(w_dff_B_v0WrVMHE7_0),.dout(w_dff_B_xb3SG3cp0_0),.clk(gclk));
	jdff dff_B_YHXAcmMC2_0(.din(w_dff_B_xb3SG3cp0_0),.dout(w_dff_B_YHXAcmMC2_0),.clk(gclk));
	jdff dff_B_fVLAJgwU3_0(.din(w_dff_B_YHXAcmMC2_0),.dout(w_dff_B_fVLAJgwU3_0),.clk(gclk));
	jdff dff_B_bB01Exob1_0(.din(w_dff_B_fVLAJgwU3_0),.dout(w_dff_B_bB01Exob1_0),.clk(gclk));
	jdff dff_B_lOHYKota2_0(.din(w_dff_B_bB01Exob1_0),.dout(w_dff_B_lOHYKota2_0),.clk(gclk));
	jdff dff_B_9ql3TWyJ3_0(.din(w_dff_B_lOHYKota2_0),.dout(w_dff_B_9ql3TWyJ3_0),.clk(gclk));
	jdff dff_B_1kldjOYI8_0(.din(w_dff_B_9ql3TWyJ3_0),.dout(w_dff_B_1kldjOYI8_0),.clk(gclk));
	jdff dff_B_oIgOlh7c4_0(.din(w_dff_B_1kldjOYI8_0),.dout(w_dff_B_oIgOlh7c4_0),.clk(gclk));
	jdff dff_B_HyOB6jnY9_0(.din(w_dff_B_oIgOlh7c4_0),.dout(w_dff_B_HyOB6jnY9_0),.clk(gclk));
	jdff dff_B_jZviLZL95_0(.din(w_dff_B_HyOB6jnY9_0),.dout(w_dff_B_jZviLZL95_0),.clk(gclk));
	jdff dff_B_8MIPVDkK5_0(.din(w_dff_B_jZviLZL95_0),.dout(w_dff_B_8MIPVDkK5_0),.clk(gclk));
	jdff dff_B_gzTQnsKE7_0(.din(w_dff_B_8MIPVDkK5_0),.dout(w_dff_B_gzTQnsKE7_0),.clk(gclk));
	jdff dff_B_7gbW1flP8_0(.din(w_dff_B_gzTQnsKE7_0),.dout(w_dff_B_7gbW1flP8_0),.clk(gclk));
	jdff dff_B_NsrK7wS07_0(.din(w_dff_B_7gbW1flP8_0),.dout(w_dff_B_NsrK7wS07_0),.clk(gclk));
	jdff dff_B_7x5hpzsk3_0(.din(w_dff_B_NsrK7wS07_0),.dout(w_dff_B_7x5hpzsk3_0),.clk(gclk));
	jdff dff_B_7W05GFDH2_0(.din(w_dff_B_7x5hpzsk3_0),.dout(w_dff_B_7W05GFDH2_0),.clk(gclk));
	jdff dff_B_yNH3dqqb9_0(.din(w_dff_B_7W05GFDH2_0),.dout(w_dff_B_yNH3dqqb9_0),.clk(gclk));
	jdff dff_B_Jf7TFLmy3_0(.din(w_dff_B_yNH3dqqb9_0),.dout(w_dff_B_Jf7TFLmy3_0),.clk(gclk));
	jdff dff_B_KyJ1suCw5_0(.din(w_dff_B_Jf7TFLmy3_0),.dout(w_dff_B_KyJ1suCw5_0),.clk(gclk));
	jdff dff_B_RxOwBrzg8_0(.din(w_dff_B_KyJ1suCw5_0),.dout(w_dff_B_RxOwBrzg8_0),.clk(gclk));
	jdff dff_B_2KaLYNB77_0(.din(w_dff_B_RxOwBrzg8_0),.dout(w_dff_B_2KaLYNB77_0),.clk(gclk));
	jdff dff_B_zAQfmmks4_0(.din(w_dff_B_2KaLYNB77_0),.dout(w_dff_B_zAQfmmks4_0),.clk(gclk));
	jdff dff_B_Coi5c6uW9_0(.din(w_dff_B_zAQfmmks4_0),.dout(w_dff_B_Coi5c6uW9_0),.clk(gclk));
	jdff dff_B_xZpFUUVQ1_0(.din(w_dff_B_Coi5c6uW9_0),.dout(w_dff_B_xZpFUUVQ1_0),.clk(gclk));
	jdff dff_B_VqPChw8q9_0(.din(w_dff_B_xZpFUUVQ1_0),.dout(w_dff_B_VqPChw8q9_0),.clk(gclk));
	jdff dff_B_8cFO0wxB1_0(.din(w_dff_B_VqPChw8q9_0),.dout(w_dff_B_8cFO0wxB1_0),.clk(gclk));
	jdff dff_B_M2vePlTa1_0(.din(w_dff_B_8cFO0wxB1_0),.dout(w_dff_B_M2vePlTa1_0),.clk(gclk));
	jdff dff_B_kfcsDZEe9_0(.din(w_dff_B_M2vePlTa1_0),.dout(w_dff_B_kfcsDZEe9_0),.clk(gclk));
	jdff dff_B_4cvrNabJ5_0(.din(w_dff_B_kfcsDZEe9_0),.dout(w_dff_B_4cvrNabJ5_0),.clk(gclk));
	jdff dff_B_PeUrXRar1_0(.din(w_dff_B_4cvrNabJ5_0),.dout(w_dff_B_PeUrXRar1_0),.clk(gclk));
	jdff dff_B_KwlAvEJO9_0(.din(w_dff_B_PeUrXRar1_0),.dout(w_dff_B_KwlAvEJO9_0),.clk(gclk));
	jdff dff_B_M5Km0IC42_0(.din(w_dff_B_KwlAvEJO9_0),.dout(w_dff_B_M5Km0IC42_0),.clk(gclk));
	jdff dff_B_WbF1jP9J5_0(.din(w_dff_B_M5Km0IC42_0),.dout(w_dff_B_WbF1jP9J5_0),.clk(gclk));
	jdff dff_B_a3KQkaOj6_0(.din(w_dff_B_WbF1jP9J5_0),.dout(w_dff_B_a3KQkaOj6_0),.clk(gclk));
	jdff dff_B_YrVuElf97_0(.din(w_dff_B_a3KQkaOj6_0),.dout(w_dff_B_YrVuElf97_0),.clk(gclk));
	jdff dff_B_ZKgBPr5l0_0(.din(w_dff_B_YrVuElf97_0),.dout(w_dff_B_ZKgBPr5l0_0),.clk(gclk));
	jdff dff_B_8dWM9WLj4_0(.din(w_dff_B_ZKgBPr5l0_0),.dout(w_dff_B_8dWM9WLj4_0),.clk(gclk));
	jdff dff_B_OyaThRrB8_0(.din(w_dff_B_8dWM9WLj4_0),.dout(w_dff_B_OyaThRrB8_0),.clk(gclk));
	jdff dff_B_BYGhXWV19_0(.din(w_dff_B_OyaThRrB8_0),.dout(w_dff_B_BYGhXWV19_0),.clk(gclk));
	jdff dff_B_KMMLpX870_0(.din(w_dff_B_BYGhXWV19_0),.dout(w_dff_B_KMMLpX870_0),.clk(gclk));
	jdff dff_B_xE22n2gA2_0(.din(w_dff_B_KMMLpX870_0),.dout(w_dff_B_xE22n2gA2_0),.clk(gclk));
	jdff dff_B_eek1d2Wg1_0(.din(w_dff_B_xE22n2gA2_0),.dout(w_dff_B_eek1d2Wg1_0),.clk(gclk));
	jdff dff_B_6LtcpZ0P2_0(.din(w_dff_B_eek1d2Wg1_0),.dout(w_dff_B_6LtcpZ0P2_0),.clk(gclk));
	jdff dff_B_PlLqyFs54_0(.din(w_dff_B_6LtcpZ0P2_0),.dout(w_dff_B_PlLqyFs54_0),.clk(gclk));
	jdff dff_B_2wn8wvNT5_0(.din(w_dff_B_PlLqyFs54_0),.dout(w_dff_B_2wn8wvNT5_0),.clk(gclk));
	jdff dff_B_NJNmvW7d4_0(.din(w_dff_B_2wn8wvNT5_0),.dout(w_dff_B_NJNmvW7d4_0),.clk(gclk));
	jdff dff_B_HQtN0HWE1_0(.din(w_dff_B_NJNmvW7d4_0),.dout(w_dff_B_HQtN0HWE1_0),.clk(gclk));
	jdff dff_B_rsVJgZa16_0(.din(w_dff_B_HQtN0HWE1_0),.dout(w_dff_B_rsVJgZa16_0),.clk(gclk));
	jdff dff_B_EWG3f3tx2_0(.din(w_dff_B_rsVJgZa16_0),.dout(w_dff_B_EWG3f3tx2_0),.clk(gclk));
	jdff dff_B_cScT3Bku6_0(.din(w_dff_B_EWG3f3tx2_0),.dout(w_dff_B_cScT3Bku6_0),.clk(gclk));
	jdff dff_B_2b5Edwz26_0(.din(w_dff_B_cScT3Bku6_0),.dout(w_dff_B_2b5Edwz26_0),.clk(gclk));
	jdff dff_B_m3vZCVYd5_0(.din(w_dff_B_2b5Edwz26_0),.dout(w_dff_B_m3vZCVYd5_0),.clk(gclk));
	jdff dff_B_1WhLU8m30_0(.din(w_dff_B_m3vZCVYd5_0),.dout(w_dff_B_1WhLU8m30_0),.clk(gclk));
	jdff dff_B_6amr7AjJ7_0(.din(w_dff_B_1WhLU8m30_0),.dout(w_dff_B_6amr7AjJ7_0),.clk(gclk));
	jdff dff_B_HDFdf9d89_0(.din(w_dff_B_6amr7AjJ7_0),.dout(w_dff_B_HDFdf9d89_0),.clk(gclk));
	jdff dff_B_v7kZVRhL5_0(.din(w_dff_B_HDFdf9d89_0),.dout(w_dff_B_v7kZVRhL5_0),.clk(gclk));
	jdff dff_B_OleMdkzj5_0(.din(w_dff_B_v7kZVRhL5_0),.dout(w_dff_B_OleMdkzj5_0),.clk(gclk));
	jdff dff_B_91Mn7IRd9_0(.din(w_dff_B_OleMdkzj5_0),.dout(w_dff_B_91Mn7IRd9_0),.clk(gclk));
	jdff dff_B_IaacLBCk8_0(.din(w_dff_B_91Mn7IRd9_0),.dout(w_dff_B_IaacLBCk8_0),.clk(gclk));
	jdff dff_B_HMJx3LXH4_0(.din(w_dff_B_IaacLBCk8_0),.dout(w_dff_B_HMJx3LXH4_0),.clk(gclk));
	jdff dff_B_cYxv0T411_0(.din(w_dff_B_HMJx3LXH4_0),.dout(w_dff_B_cYxv0T411_0),.clk(gclk));
	jdff dff_B_8VYO2KIZ4_0(.din(w_dff_B_cYxv0T411_0),.dout(w_dff_B_8VYO2KIZ4_0),.clk(gclk));
	jdff dff_B_Fv0xdtCj1_0(.din(w_dff_B_8VYO2KIZ4_0),.dout(w_dff_B_Fv0xdtCj1_0),.clk(gclk));
	jdff dff_B_ei42O0my7_0(.din(w_dff_B_Fv0xdtCj1_0),.dout(w_dff_B_ei42O0my7_0),.clk(gclk));
	jdff dff_B_smcaRgdt0_0(.din(w_dff_B_ei42O0my7_0),.dout(w_dff_B_smcaRgdt0_0),.clk(gclk));
	jdff dff_B_OmXcePvN4_0(.din(w_dff_B_smcaRgdt0_0),.dout(w_dff_B_OmXcePvN4_0),.clk(gclk));
	jdff dff_B_JwZqahIm8_0(.din(w_dff_B_OmXcePvN4_0),.dout(w_dff_B_JwZqahIm8_0),.clk(gclk));
	jdff dff_B_5gDMRACq6_0(.din(w_dff_B_JwZqahIm8_0),.dout(w_dff_B_5gDMRACq6_0),.clk(gclk));
	jdff dff_B_pgIX1swX2_0(.din(w_dff_B_5gDMRACq6_0),.dout(w_dff_B_pgIX1swX2_0),.clk(gclk));
	jdff dff_B_logAA0ks9_0(.din(w_dff_B_pgIX1swX2_0),.dout(w_dff_B_logAA0ks9_0),.clk(gclk));
	jdff dff_B_BVXBqqUR5_0(.din(w_dff_B_logAA0ks9_0),.dout(w_dff_B_BVXBqqUR5_0),.clk(gclk));
	jdff dff_B_slySt0GR3_0(.din(w_dff_B_BVXBqqUR5_0),.dout(w_dff_B_slySt0GR3_0),.clk(gclk));
	jdff dff_B_zBnkBPnf2_0(.din(w_dff_B_slySt0GR3_0),.dout(w_dff_B_zBnkBPnf2_0),.clk(gclk));
	jdff dff_B_Noal6Ocm4_0(.din(w_dff_B_zBnkBPnf2_0),.dout(w_dff_B_Noal6Ocm4_0),.clk(gclk));
	jdff dff_B_2GmTQCri3_0(.din(w_dff_B_Noal6Ocm4_0),.dout(w_dff_B_2GmTQCri3_0),.clk(gclk));
	jdff dff_B_vNriQ0Vb5_0(.din(w_dff_B_2GmTQCri3_0),.dout(w_dff_B_vNriQ0Vb5_0),.clk(gclk));
	jdff dff_B_dAe9zNSK3_0(.din(w_dff_B_vNriQ0Vb5_0),.dout(w_dff_B_dAe9zNSK3_0),.clk(gclk));
	jdff dff_B_OC7rTDjS7_0(.din(w_dff_B_dAe9zNSK3_0),.dout(w_dff_B_OC7rTDjS7_0),.clk(gclk));
	jdff dff_B_kCm3iSPC2_0(.din(w_dff_B_OC7rTDjS7_0),.dout(w_dff_B_kCm3iSPC2_0),.clk(gclk));
	jdff dff_B_YgouYNVU9_0(.din(w_dff_B_kCm3iSPC2_0),.dout(w_dff_B_YgouYNVU9_0),.clk(gclk));
	jdff dff_B_oBZLviGg4_0(.din(w_dff_B_YgouYNVU9_0),.dout(w_dff_B_oBZLviGg4_0),.clk(gclk));
	jdff dff_B_vgkiyEAh6_0(.din(w_dff_B_oBZLviGg4_0),.dout(w_dff_B_vgkiyEAh6_0),.clk(gclk));
	jdff dff_B_fhcfjD9y4_0(.din(n934),.dout(w_dff_B_fhcfjD9y4_0),.clk(gclk));
	jdff dff_B_XPUb2IrR6_0(.din(w_dff_B_fhcfjD9y4_0),.dout(w_dff_B_XPUb2IrR6_0),.clk(gclk));
	jdff dff_B_Yi1rEeFd2_0(.din(w_dff_B_XPUb2IrR6_0),.dout(w_dff_B_Yi1rEeFd2_0),.clk(gclk));
	jdff dff_B_HxQvK6lw6_0(.din(w_dff_B_Yi1rEeFd2_0),.dout(w_dff_B_HxQvK6lw6_0),.clk(gclk));
	jdff dff_B_rNhTu0Fi9_0(.din(w_dff_B_HxQvK6lw6_0),.dout(w_dff_B_rNhTu0Fi9_0),.clk(gclk));
	jdff dff_B_OcI7n4Lp2_0(.din(w_dff_B_rNhTu0Fi9_0),.dout(w_dff_B_OcI7n4Lp2_0),.clk(gclk));
	jdff dff_B_RsujpwAI8_0(.din(w_dff_B_OcI7n4Lp2_0),.dout(w_dff_B_RsujpwAI8_0),.clk(gclk));
	jdff dff_B_NrE4IRjb7_0(.din(w_dff_B_RsujpwAI8_0),.dout(w_dff_B_NrE4IRjb7_0),.clk(gclk));
	jdff dff_B_Xfw0J6eh3_0(.din(w_dff_B_NrE4IRjb7_0),.dout(w_dff_B_Xfw0J6eh3_0),.clk(gclk));
	jdff dff_B_UdcaEZAD4_0(.din(w_dff_B_Xfw0J6eh3_0),.dout(w_dff_B_UdcaEZAD4_0),.clk(gclk));
	jdff dff_B_7pOuXS1g4_0(.din(w_dff_B_UdcaEZAD4_0),.dout(w_dff_B_7pOuXS1g4_0),.clk(gclk));
	jdff dff_B_QE1Q7emD3_0(.din(w_dff_B_7pOuXS1g4_0),.dout(w_dff_B_QE1Q7emD3_0),.clk(gclk));
	jdff dff_B_eA957Lio5_0(.din(w_dff_B_QE1Q7emD3_0),.dout(w_dff_B_eA957Lio5_0),.clk(gclk));
	jdff dff_B_9QEuLWPn3_0(.din(w_dff_B_eA957Lio5_0),.dout(w_dff_B_9QEuLWPn3_0),.clk(gclk));
	jdff dff_B_XVbpx3LL7_0(.din(w_dff_B_9QEuLWPn3_0),.dout(w_dff_B_XVbpx3LL7_0),.clk(gclk));
	jdff dff_B_IV28YlRB1_0(.din(w_dff_B_XVbpx3LL7_0),.dout(w_dff_B_IV28YlRB1_0),.clk(gclk));
	jdff dff_B_YWPOyVwS0_0(.din(w_dff_B_IV28YlRB1_0),.dout(w_dff_B_YWPOyVwS0_0),.clk(gclk));
	jdff dff_B_eNgZMEAZ9_0(.din(w_dff_B_YWPOyVwS0_0),.dout(w_dff_B_eNgZMEAZ9_0),.clk(gclk));
	jdff dff_B_OA6rj82y0_0(.din(w_dff_B_eNgZMEAZ9_0),.dout(w_dff_B_OA6rj82y0_0),.clk(gclk));
	jdff dff_B_mjzcpdz86_0(.din(w_dff_B_OA6rj82y0_0),.dout(w_dff_B_mjzcpdz86_0),.clk(gclk));
	jdff dff_B_YHOhW1QB9_0(.din(w_dff_B_mjzcpdz86_0),.dout(w_dff_B_YHOhW1QB9_0),.clk(gclk));
	jdff dff_B_Pdbx63Z19_0(.din(w_dff_B_YHOhW1QB9_0),.dout(w_dff_B_Pdbx63Z19_0),.clk(gclk));
	jdff dff_B_RNaotcwI3_0(.din(w_dff_B_Pdbx63Z19_0),.dout(w_dff_B_RNaotcwI3_0),.clk(gclk));
	jdff dff_B_57BS15644_0(.din(w_dff_B_RNaotcwI3_0),.dout(w_dff_B_57BS15644_0),.clk(gclk));
	jdff dff_B_55ZTfQup5_0(.din(w_dff_B_57BS15644_0),.dout(w_dff_B_55ZTfQup5_0),.clk(gclk));
	jdff dff_B_HCgo7Hcf4_0(.din(w_dff_B_55ZTfQup5_0),.dout(w_dff_B_HCgo7Hcf4_0),.clk(gclk));
	jdff dff_B_OMyKHvgZ2_0(.din(w_dff_B_HCgo7Hcf4_0),.dout(w_dff_B_OMyKHvgZ2_0),.clk(gclk));
	jdff dff_B_x9ZWGzaE2_0(.din(w_dff_B_OMyKHvgZ2_0),.dout(w_dff_B_x9ZWGzaE2_0),.clk(gclk));
	jdff dff_B_IIiexAjM3_0(.din(w_dff_B_x9ZWGzaE2_0),.dout(w_dff_B_IIiexAjM3_0),.clk(gclk));
	jdff dff_B_mB6wE1yn1_0(.din(w_dff_B_IIiexAjM3_0),.dout(w_dff_B_mB6wE1yn1_0),.clk(gclk));
	jdff dff_B_fL2y0fpg7_0(.din(w_dff_B_mB6wE1yn1_0),.dout(w_dff_B_fL2y0fpg7_0),.clk(gclk));
	jdff dff_B_0keNPwNm7_0(.din(w_dff_B_fL2y0fpg7_0),.dout(w_dff_B_0keNPwNm7_0),.clk(gclk));
	jdff dff_B_0YU51EUf1_0(.din(w_dff_B_0keNPwNm7_0),.dout(w_dff_B_0YU51EUf1_0),.clk(gclk));
	jdff dff_B_1fRvMtBU8_0(.din(w_dff_B_0YU51EUf1_0),.dout(w_dff_B_1fRvMtBU8_0),.clk(gclk));
	jdff dff_B_eNM5LHYZ1_0(.din(w_dff_B_1fRvMtBU8_0),.dout(w_dff_B_eNM5LHYZ1_0),.clk(gclk));
	jdff dff_B_mmumLB8T4_0(.din(w_dff_B_eNM5LHYZ1_0),.dout(w_dff_B_mmumLB8T4_0),.clk(gclk));
	jdff dff_B_24OWo8On2_0(.din(w_dff_B_mmumLB8T4_0),.dout(w_dff_B_24OWo8On2_0),.clk(gclk));
	jdff dff_B_Xnkv6wpE2_0(.din(w_dff_B_24OWo8On2_0),.dout(w_dff_B_Xnkv6wpE2_0),.clk(gclk));
	jdff dff_B_ClGaX7et6_0(.din(w_dff_B_Xnkv6wpE2_0),.dout(w_dff_B_ClGaX7et6_0),.clk(gclk));
	jdff dff_B_ZkimcW9H4_0(.din(w_dff_B_ClGaX7et6_0),.dout(w_dff_B_ZkimcW9H4_0),.clk(gclk));
	jdff dff_B_wuLaYuXU0_0(.din(w_dff_B_ZkimcW9H4_0),.dout(w_dff_B_wuLaYuXU0_0),.clk(gclk));
	jdff dff_B_6oRMzsHG0_0(.din(w_dff_B_wuLaYuXU0_0),.dout(w_dff_B_6oRMzsHG0_0),.clk(gclk));
	jdff dff_B_hcqYwIxD0_0(.din(w_dff_B_6oRMzsHG0_0),.dout(w_dff_B_hcqYwIxD0_0),.clk(gclk));
	jdff dff_B_GLy3QedQ0_0(.din(w_dff_B_hcqYwIxD0_0),.dout(w_dff_B_GLy3QedQ0_0),.clk(gclk));
	jdff dff_B_g7nyyOxt6_0(.din(w_dff_B_GLy3QedQ0_0),.dout(w_dff_B_g7nyyOxt6_0),.clk(gclk));
	jdff dff_B_Hj2cCQXp4_0(.din(w_dff_B_g7nyyOxt6_0),.dout(w_dff_B_Hj2cCQXp4_0),.clk(gclk));
	jdff dff_B_7qQeG4ym9_0(.din(w_dff_B_Hj2cCQXp4_0),.dout(w_dff_B_7qQeG4ym9_0),.clk(gclk));
	jdff dff_B_zj3Ax0SY9_0(.din(w_dff_B_7qQeG4ym9_0),.dout(w_dff_B_zj3Ax0SY9_0),.clk(gclk));
	jdff dff_B_JVfwb49E3_0(.din(w_dff_B_zj3Ax0SY9_0),.dout(w_dff_B_JVfwb49E3_0),.clk(gclk));
	jdff dff_B_v0Ap766Z6_0(.din(w_dff_B_JVfwb49E3_0),.dout(w_dff_B_v0Ap766Z6_0),.clk(gclk));
	jdff dff_B_OVzwgguU2_0(.din(w_dff_B_v0Ap766Z6_0),.dout(w_dff_B_OVzwgguU2_0),.clk(gclk));
	jdff dff_B_enkNNa8E7_0(.din(w_dff_B_OVzwgguU2_0),.dout(w_dff_B_enkNNa8E7_0),.clk(gclk));
	jdff dff_B_5tjnvZyx1_0(.din(w_dff_B_enkNNa8E7_0),.dout(w_dff_B_5tjnvZyx1_0),.clk(gclk));
	jdff dff_B_ldNbWkD46_0(.din(w_dff_B_5tjnvZyx1_0),.dout(w_dff_B_ldNbWkD46_0),.clk(gclk));
	jdff dff_B_razZ34i70_0(.din(w_dff_B_ldNbWkD46_0),.dout(w_dff_B_razZ34i70_0),.clk(gclk));
	jdff dff_B_iA3bsgiS9_0(.din(w_dff_B_razZ34i70_0),.dout(w_dff_B_iA3bsgiS9_0),.clk(gclk));
	jdff dff_B_WQN2CA9w4_0(.din(w_dff_B_iA3bsgiS9_0),.dout(w_dff_B_WQN2CA9w4_0),.clk(gclk));
	jdff dff_B_eqPSxxTU2_0(.din(w_dff_B_WQN2CA9w4_0),.dout(w_dff_B_eqPSxxTU2_0),.clk(gclk));
	jdff dff_B_hf3r0Hiu1_0(.din(w_dff_B_eqPSxxTU2_0),.dout(w_dff_B_hf3r0Hiu1_0),.clk(gclk));
	jdff dff_B_hiOftxfl0_0(.din(w_dff_B_hf3r0Hiu1_0),.dout(w_dff_B_hiOftxfl0_0),.clk(gclk));
	jdff dff_B_30Lb7JtM3_0(.din(w_dff_B_hiOftxfl0_0),.dout(w_dff_B_30Lb7JtM3_0),.clk(gclk));
	jdff dff_B_iU7lI2O91_0(.din(w_dff_B_30Lb7JtM3_0),.dout(w_dff_B_iU7lI2O91_0),.clk(gclk));
	jdff dff_B_0cwLrV9z8_0(.din(w_dff_B_iU7lI2O91_0),.dout(w_dff_B_0cwLrV9z8_0),.clk(gclk));
	jdff dff_B_tQitZD2H6_0(.din(w_dff_B_0cwLrV9z8_0),.dout(w_dff_B_tQitZD2H6_0),.clk(gclk));
	jdff dff_B_mbBXjP7c9_0(.din(w_dff_B_tQitZD2H6_0),.dout(w_dff_B_mbBXjP7c9_0),.clk(gclk));
	jdff dff_B_ctXXeX4L3_0(.din(w_dff_B_mbBXjP7c9_0),.dout(w_dff_B_ctXXeX4L3_0),.clk(gclk));
	jdff dff_B_aiRcMePC2_0(.din(w_dff_B_ctXXeX4L3_0),.dout(w_dff_B_aiRcMePC2_0),.clk(gclk));
	jdff dff_B_sNHO2xgZ7_0(.din(w_dff_B_aiRcMePC2_0),.dout(w_dff_B_sNHO2xgZ7_0),.clk(gclk));
	jdff dff_B_ginmtGZ63_0(.din(w_dff_B_sNHO2xgZ7_0),.dout(w_dff_B_ginmtGZ63_0),.clk(gclk));
	jdff dff_B_K9pCFAio9_0(.din(w_dff_B_ginmtGZ63_0),.dout(w_dff_B_K9pCFAio9_0),.clk(gclk));
	jdff dff_B_K67xS4pS4_0(.din(w_dff_B_K9pCFAio9_0),.dout(w_dff_B_K67xS4pS4_0),.clk(gclk));
	jdff dff_B_hVqyHXBV9_0(.din(w_dff_B_K67xS4pS4_0),.dout(w_dff_B_hVqyHXBV9_0),.clk(gclk));
	jdff dff_B_6z6HtBD57_0(.din(w_dff_B_hVqyHXBV9_0),.dout(w_dff_B_6z6HtBD57_0),.clk(gclk));
	jdff dff_B_AUHRhyGt5_0(.din(w_dff_B_6z6HtBD57_0),.dout(w_dff_B_AUHRhyGt5_0),.clk(gclk));
	jdff dff_B_TkgeNQY00_0(.din(w_dff_B_AUHRhyGt5_0),.dout(w_dff_B_TkgeNQY00_0),.clk(gclk));
	jdff dff_B_zpwJvQ515_0(.din(w_dff_B_TkgeNQY00_0),.dout(w_dff_B_zpwJvQ515_0),.clk(gclk));
	jdff dff_B_WDjhrQKW0_0(.din(w_dff_B_zpwJvQ515_0),.dout(w_dff_B_WDjhrQKW0_0),.clk(gclk));
	jdff dff_B_V270VAkB9_0(.din(w_dff_B_WDjhrQKW0_0),.dout(w_dff_B_V270VAkB9_0),.clk(gclk));
	jdff dff_B_ycw05gBQ0_0(.din(w_dff_B_V270VAkB9_0),.dout(w_dff_B_ycw05gBQ0_0),.clk(gclk));
	jdff dff_B_lcnAP0z92_0(.din(w_dff_B_ycw05gBQ0_0),.dout(w_dff_B_lcnAP0z92_0),.clk(gclk));
	jdff dff_B_DfF5ngS37_0(.din(w_dff_B_lcnAP0z92_0),.dout(w_dff_B_DfF5ngS37_0),.clk(gclk));
	jdff dff_B_NXHrwrVd0_0(.din(w_dff_B_DfF5ngS37_0),.dout(w_dff_B_NXHrwrVd0_0),.clk(gclk));
	jdff dff_B_AGThUvVk7_0(.din(w_dff_B_NXHrwrVd0_0),.dout(w_dff_B_AGThUvVk7_0),.clk(gclk));
	jdff dff_B_RNRT9YyD6_0(.din(w_dff_B_AGThUvVk7_0),.dout(w_dff_B_RNRT9YyD6_0),.clk(gclk));
	jdff dff_B_aBoh4ovx6_0(.din(w_dff_B_RNRT9YyD6_0),.dout(w_dff_B_aBoh4ovx6_0),.clk(gclk));
	jdff dff_B_JindIYki7_0(.din(w_dff_B_aBoh4ovx6_0),.dout(w_dff_B_JindIYki7_0),.clk(gclk));
	jdff dff_B_c0dpcB5P3_0(.din(w_dff_B_JindIYki7_0),.dout(w_dff_B_c0dpcB5P3_0),.clk(gclk));
	jdff dff_B_s7MyU8fC4_0(.din(w_dff_B_c0dpcB5P3_0),.dout(w_dff_B_s7MyU8fC4_0),.clk(gclk));
	jdff dff_B_MoIgWBGR4_0(.din(w_dff_B_s7MyU8fC4_0),.dout(w_dff_B_MoIgWBGR4_0),.clk(gclk));
	jdff dff_B_ub22zWvN3_0(.din(w_dff_B_MoIgWBGR4_0),.dout(w_dff_B_ub22zWvN3_0),.clk(gclk));
	jdff dff_B_lJOSsY171_0(.din(w_dff_B_ub22zWvN3_0),.dout(w_dff_B_lJOSsY171_0),.clk(gclk));
	jdff dff_B_L6XEqsQD2_0(.din(n940),.dout(w_dff_B_L6XEqsQD2_0),.clk(gclk));
	jdff dff_B_I4C07N0v0_0(.din(w_dff_B_L6XEqsQD2_0),.dout(w_dff_B_I4C07N0v0_0),.clk(gclk));
	jdff dff_B_wXsBjVto8_0(.din(w_dff_B_I4C07N0v0_0),.dout(w_dff_B_wXsBjVto8_0),.clk(gclk));
	jdff dff_B_9vfeCqXL4_0(.din(w_dff_B_wXsBjVto8_0),.dout(w_dff_B_9vfeCqXL4_0),.clk(gclk));
	jdff dff_B_cjd6mApc6_0(.din(w_dff_B_9vfeCqXL4_0),.dout(w_dff_B_cjd6mApc6_0),.clk(gclk));
	jdff dff_B_ZuhHacUi8_0(.din(w_dff_B_cjd6mApc6_0),.dout(w_dff_B_ZuhHacUi8_0),.clk(gclk));
	jdff dff_B_jqPInde50_0(.din(w_dff_B_ZuhHacUi8_0),.dout(w_dff_B_jqPInde50_0),.clk(gclk));
	jdff dff_B_ItioxTAY9_0(.din(w_dff_B_jqPInde50_0),.dout(w_dff_B_ItioxTAY9_0),.clk(gclk));
	jdff dff_B_0QPZ31Wc8_0(.din(w_dff_B_ItioxTAY9_0),.dout(w_dff_B_0QPZ31Wc8_0),.clk(gclk));
	jdff dff_B_lpUMr7ja7_0(.din(w_dff_B_0QPZ31Wc8_0),.dout(w_dff_B_lpUMr7ja7_0),.clk(gclk));
	jdff dff_B_MTK2mGuD8_0(.din(w_dff_B_lpUMr7ja7_0),.dout(w_dff_B_MTK2mGuD8_0),.clk(gclk));
	jdff dff_B_t0AoUYbB4_0(.din(w_dff_B_MTK2mGuD8_0),.dout(w_dff_B_t0AoUYbB4_0),.clk(gclk));
	jdff dff_B_LKPy1WfB0_0(.din(w_dff_B_t0AoUYbB4_0),.dout(w_dff_B_LKPy1WfB0_0),.clk(gclk));
	jdff dff_B_h8DSVQj50_0(.din(w_dff_B_LKPy1WfB0_0),.dout(w_dff_B_h8DSVQj50_0),.clk(gclk));
	jdff dff_B_ikxjbfcP3_0(.din(w_dff_B_h8DSVQj50_0),.dout(w_dff_B_ikxjbfcP3_0),.clk(gclk));
	jdff dff_B_SXAKrERt1_0(.din(w_dff_B_ikxjbfcP3_0),.dout(w_dff_B_SXAKrERt1_0),.clk(gclk));
	jdff dff_B_57EwLenK7_0(.din(w_dff_B_SXAKrERt1_0),.dout(w_dff_B_57EwLenK7_0),.clk(gclk));
	jdff dff_B_0bl1NVbR4_0(.din(w_dff_B_57EwLenK7_0),.dout(w_dff_B_0bl1NVbR4_0),.clk(gclk));
	jdff dff_B_cJmYllNu8_0(.din(w_dff_B_0bl1NVbR4_0),.dout(w_dff_B_cJmYllNu8_0),.clk(gclk));
	jdff dff_B_S0eHrJej0_0(.din(w_dff_B_cJmYllNu8_0),.dout(w_dff_B_S0eHrJej0_0),.clk(gclk));
	jdff dff_B_pjfiUR7r9_0(.din(w_dff_B_S0eHrJej0_0),.dout(w_dff_B_pjfiUR7r9_0),.clk(gclk));
	jdff dff_B_Twpr0dGv4_0(.din(w_dff_B_pjfiUR7r9_0),.dout(w_dff_B_Twpr0dGv4_0),.clk(gclk));
	jdff dff_B_eW4XODF99_0(.din(w_dff_B_Twpr0dGv4_0),.dout(w_dff_B_eW4XODF99_0),.clk(gclk));
	jdff dff_B_Jo1gIF7K4_0(.din(w_dff_B_eW4XODF99_0),.dout(w_dff_B_Jo1gIF7K4_0),.clk(gclk));
	jdff dff_B_VnSgSmds6_0(.din(w_dff_B_Jo1gIF7K4_0),.dout(w_dff_B_VnSgSmds6_0),.clk(gclk));
	jdff dff_B_z06JAgyL8_0(.din(w_dff_B_VnSgSmds6_0),.dout(w_dff_B_z06JAgyL8_0),.clk(gclk));
	jdff dff_B_f9r7QJFW6_0(.din(w_dff_B_z06JAgyL8_0),.dout(w_dff_B_f9r7QJFW6_0),.clk(gclk));
	jdff dff_B_BfgMa1Bj8_0(.din(w_dff_B_f9r7QJFW6_0),.dout(w_dff_B_BfgMa1Bj8_0),.clk(gclk));
	jdff dff_B_i5lceecz9_0(.din(w_dff_B_BfgMa1Bj8_0),.dout(w_dff_B_i5lceecz9_0),.clk(gclk));
	jdff dff_B_78vPS1tb1_0(.din(w_dff_B_i5lceecz9_0),.dout(w_dff_B_78vPS1tb1_0),.clk(gclk));
	jdff dff_B_YgGHVgip6_0(.din(w_dff_B_78vPS1tb1_0),.dout(w_dff_B_YgGHVgip6_0),.clk(gclk));
	jdff dff_B_QBbMYkpT0_0(.din(w_dff_B_YgGHVgip6_0),.dout(w_dff_B_QBbMYkpT0_0),.clk(gclk));
	jdff dff_B_V4yv1Dm83_0(.din(w_dff_B_QBbMYkpT0_0),.dout(w_dff_B_V4yv1Dm83_0),.clk(gclk));
	jdff dff_B_CPKzqgqd9_0(.din(w_dff_B_V4yv1Dm83_0),.dout(w_dff_B_CPKzqgqd9_0),.clk(gclk));
	jdff dff_B_0oeP7dUY2_0(.din(w_dff_B_CPKzqgqd9_0),.dout(w_dff_B_0oeP7dUY2_0),.clk(gclk));
	jdff dff_B_pumxgpUT7_0(.din(w_dff_B_0oeP7dUY2_0),.dout(w_dff_B_pumxgpUT7_0),.clk(gclk));
	jdff dff_B_RlP2hxfb9_0(.din(w_dff_B_pumxgpUT7_0),.dout(w_dff_B_RlP2hxfb9_0),.clk(gclk));
	jdff dff_B_H5RqFnkF4_0(.din(w_dff_B_RlP2hxfb9_0),.dout(w_dff_B_H5RqFnkF4_0),.clk(gclk));
	jdff dff_B_Vyawy5hR4_0(.din(w_dff_B_H5RqFnkF4_0),.dout(w_dff_B_Vyawy5hR4_0),.clk(gclk));
	jdff dff_B_TTvxEKge3_0(.din(w_dff_B_Vyawy5hR4_0),.dout(w_dff_B_TTvxEKge3_0),.clk(gclk));
	jdff dff_B_lgsZtvDU5_0(.din(w_dff_B_TTvxEKge3_0),.dout(w_dff_B_lgsZtvDU5_0),.clk(gclk));
	jdff dff_B_dXyKjo3Z3_0(.din(w_dff_B_lgsZtvDU5_0),.dout(w_dff_B_dXyKjo3Z3_0),.clk(gclk));
	jdff dff_B_xqNNXwyF1_0(.din(w_dff_B_dXyKjo3Z3_0),.dout(w_dff_B_xqNNXwyF1_0),.clk(gclk));
	jdff dff_B_e1hQjS0U0_0(.din(w_dff_B_xqNNXwyF1_0),.dout(w_dff_B_e1hQjS0U0_0),.clk(gclk));
	jdff dff_B_LyveZ1Xv9_0(.din(w_dff_B_e1hQjS0U0_0),.dout(w_dff_B_LyveZ1Xv9_0),.clk(gclk));
	jdff dff_B_oQyy2W5V3_0(.din(w_dff_B_LyveZ1Xv9_0),.dout(w_dff_B_oQyy2W5V3_0),.clk(gclk));
	jdff dff_B_l8okepPR3_0(.din(w_dff_B_oQyy2W5V3_0),.dout(w_dff_B_l8okepPR3_0),.clk(gclk));
	jdff dff_B_NgmasIYY3_0(.din(w_dff_B_l8okepPR3_0),.dout(w_dff_B_NgmasIYY3_0),.clk(gclk));
	jdff dff_B_ValgLkKF1_0(.din(w_dff_B_NgmasIYY3_0),.dout(w_dff_B_ValgLkKF1_0),.clk(gclk));
	jdff dff_B_9g6oaCFv5_0(.din(w_dff_B_ValgLkKF1_0),.dout(w_dff_B_9g6oaCFv5_0),.clk(gclk));
	jdff dff_B_CORAAWD78_0(.din(w_dff_B_9g6oaCFv5_0),.dout(w_dff_B_CORAAWD78_0),.clk(gclk));
	jdff dff_B_5MdrKi917_0(.din(w_dff_B_CORAAWD78_0),.dout(w_dff_B_5MdrKi917_0),.clk(gclk));
	jdff dff_B_qdA9zPt24_0(.din(w_dff_B_5MdrKi917_0),.dout(w_dff_B_qdA9zPt24_0),.clk(gclk));
	jdff dff_B_HaUILZLG0_0(.din(w_dff_B_qdA9zPt24_0),.dout(w_dff_B_HaUILZLG0_0),.clk(gclk));
	jdff dff_B_0PzgsZbI1_0(.din(w_dff_B_HaUILZLG0_0),.dout(w_dff_B_0PzgsZbI1_0),.clk(gclk));
	jdff dff_B_mpeAJpV75_0(.din(w_dff_B_0PzgsZbI1_0),.dout(w_dff_B_mpeAJpV75_0),.clk(gclk));
	jdff dff_B_zrk2oeIB9_0(.din(w_dff_B_mpeAJpV75_0),.dout(w_dff_B_zrk2oeIB9_0),.clk(gclk));
	jdff dff_B_ZSdTDVQk8_0(.din(w_dff_B_zrk2oeIB9_0),.dout(w_dff_B_ZSdTDVQk8_0),.clk(gclk));
	jdff dff_B_sGHXupt62_0(.din(w_dff_B_ZSdTDVQk8_0),.dout(w_dff_B_sGHXupt62_0),.clk(gclk));
	jdff dff_B_wDbBQEJO2_0(.din(w_dff_B_sGHXupt62_0),.dout(w_dff_B_wDbBQEJO2_0),.clk(gclk));
	jdff dff_B_ZbwhacVQ4_0(.din(w_dff_B_wDbBQEJO2_0),.dout(w_dff_B_ZbwhacVQ4_0),.clk(gclk));
	jdff dff_B_IT05QkwA1_0(.din(w_dff_B_ZbwhacVQ4_0),.dout(w_dff_B_IT05QkwA1_0),.clk(gclk));
	jdff dff_B_6lP44hqT6_0(.din(w_dff_B_IT05QkwA1_0),.dout(w_dff_B_6lP44hqT6_0),.clk(gclk));
	jdff dff_B_tNCiAupb8_0(.din(w_dff_B_6lP44hqT6_0),.dout(w_dff_B_tNCiAupb8_0),.clk(gclk));
	jdff dff_B_DdJ72lJM3_0(.din(w_dff_B_tNCiAupb8_0),.dout(w_dff_B_DdJ72lJM3_0),.clk(gclk));
	jdff dff_B_xj5rbALU6_0(.din(w_dff_B_DdJ72lJM3_0),.dout(w_dff_B_xj5rbALU6_0),.clk(gclk));
	jdff dff_B_IeLeMarR4_0(.din(w_dff_B_xj5rbALU6_0),.dout(w_dff_B_IeLeMarR4_0),.clk(gclk));
	jdff dff_B_bI9VxqpI7_0(.din(w_dff_B_IeLeMarR4_0),.dout(w_dff_B_bI9VxqpI7_0),.clk(gclk));
	jdff dff_B_CXeqhXDz3_0(.din(w_dff_B_bI9VxqpI7_0),.dout(w_dff_B_CXeqhXDz3_0),.clk(gclk));
	jdff dff_B_3yANIJ0n1_0(.din(w_dff_B_CXeqhXDz3_0),.dout(w_dff_B_3yANIJ0n1_0),.clk(gclk));
	jdff dff_B_SgKEG25y2_0(.din(w_dff_B_3yANIJ0n1_0),.dout(w_dff_B_SgKEG25y2_0),.clk(gclk));
	jdff dff_B_rtLKtDF75_0(.din(w_dff_B_SgKEG25y2_0),.dout(w_dff_B_rtLKtDF75_0),.clk(gclk));
	jdff dff_B_tsJ7SVNS7_0(.din(w_dff_B_rtLKtDF75_0),.dout(w_dff_B_tsJ7SVNS7_0),.clk(gclk));
	jdff dff_B_cR2iWGNm2_0(.din(w_dff_B_tsJ7SVNS7_0),.dout(w_dff_B_cR2iWGNm2_0),.clk(gclk));
	jdff dff_B_qXsr8YMz5_0(.din(w_dff_B_cR2iWGNm2_0),.dout(w_dff_B_qXsr8YMz5_0),.clk(gclk));
	jdff dff_B_1xXRNM1N8_0(.din(w_dff_B_qXsr8YMz5_0),.dout(w_dff_B_1xXRNM1N8_0),.clk(gclk));
	jdff dff_B_8vJgU9Pd0_0(.din(w_dff_B_1xXRNM1N8_0),.dout(w_dff_B_8vJgU9Pd0_0),.clk(gclk));
	jdff dff_B_neOEgyy66_0(.din(w_dff_B_8vJgU9Pd0_0),.dout(w_dff_B_neOEgyy66_0),.clk(gclk));
	jdff dff_B_g7yG9TCX9_0(.din(w_dff_B_neOEgyy66_0),.dout(w_dff_B_g7yG9TCX9_0),.clk(gclk));
	jdff dff_B_ObmE9enM5_0(.din(w_dff_B_g7yG9TCX9_0),.dout(w_dff_B_ObmE9enM5_0),.clk(gclk));
	jdff dff_B_xG7ijfTh9_0(.din(w_dff_B_ObmE9enM5_0),.dout(w_dff_B_xG7ijfTh9_0),.clk(gclk));
	jdff dff_B_r29RsP4F6_0(.din(w_dff_B_xG7ijfTh9_0),.dout(w_dff_B_r29RsP4F6_0),.clk(gclk));
	jdff dff_B_GC0tytrT3_0(.din(w_dff_B_r29RsP4F6_0),.dout(w_dff_B_GC0tytrT3_0),.clk(gclk));
	jdff dff_B_maDeWo187_0(.din(w_dff_B_GC0tytrT3_0),.dout(w_dff_B_maDeWo187_0),.clk(gclk));
	jdff dff_B_99vLvXpZ7_0(.din(w_dff_B_maDeWo187_0),.dout(w_dff_B_99vLvXpZ7_0),.clk(gclk));
	jdff dff_B_aOkopAdL7_0(.din(w_dff_B_99vLvXpZ7_0),.dout(w_dff_B_aOkopAdL7_0),.clk(gclk));
	jdff dff_B_iENNeByh6_0(.din(w_dff_B_aOkopAdL7_0),.dout(w_dff_B_iENNeByh6_0),.clk(gclk));
	jdff dff_B_lDGt7iS93_0(.din(w_dff_B_iENNeByh6_0),.dout(w_dff_B_lDGt7iS93_0),.clk(gclk));
	jdff dff_B_ANGAEBR29_0(.din(w_dff_B_lDGt7iS93_0),.dout(w_dff_B_ANGAEBR29_0),.clk(gclk));
	jdff dff_B_EROz8aSS0_0(.din(w_dff_B_ANGAEBR29_0),.dout(w_dff_B_EROz8aSS0_0),.clk(gclk));
	jdff dff_B_HVTuliIy6_0(.din(w_dff_B_EROz8aSS0_0),.dout(w_dff_B_HVTuliIy6_0),.clk(gclk));
	jdff dff_B_pbghLIdh4_0(.din(w_dff_B_HVTuliIy6_0),.dout(w_dff_B_pbghLIdh4_0),.clk(gclk));
	jdff dff_B_OqqO1U7D9_0(.din(n946),.dout(w_dff_B_OqqO1U7D9_0),.clk(gclk));
	jdff dff_B_JiyGNTAj4_0(.din(w_dff_B_OqqO1U7D9_0),.dout(w_dff_B_JiyGNTAj4_0),.clk(gclk));
	jdff dff_B_XUnZMClu4_0(.din(w_dff_B_JiyGNTAj4_0),.dout(w_dff_B_XUnZMClu4_0),.clk(gclk));
	jdff dff_B_DlU8PPoj8_0(.din(w_dff_B_XUnZMClu4_0),.dout(w_dff_B_DlU8PPoj8_0),.clk(gclk));
	jdff dff_B_VxUgdIIL1_0(.din(w_dff_B_DlU8PPoj8_0),.dout(w_dff_B_VxUgdIIL1_0),.clk(gclk));
	jdff dff_B_mYBB8z7y8_0(.din(w_dff_B_VxUgdIIL1_0),.dout(w_dff_B_mYBB8z7y8_0),.clk(gclk));
	jdff dff_B_HjJ4US4Q1_0(.din(w_dff_B_mYBB8z7y8_0),.dout(w_dff_B_HjJ4US4Q1_0),.clk(gclk));
	jdff dff_B_r3VVL3Wb7_0(.din(w_dff_B_HjJ4US4Q1_0),.dout(w_dff_B_r3VVL3Wb7_0),.clk(gclk));
	jdff dff_B_voI9mhzg2_0(.din(w_dff_B_r3VVL3Wb7_0),.dout(w_dff_B_voI9mhzg2_0),.clk(gclk));
	jdff dff_B_FqLqem4x5_0(.din(w_dff_B_voI9mhzg2_0),.dout(w_dff_B_FqLqem4x5_0),.clk(gclk));
	jdff dff_B_lShsHD8R7_0(.din(w_dff_B_FqLqem4x5_0),.dout(w_dff_B_lShsHD8R7_0),.clk(gclk));
	jdff dff_B_bkKN7mRm3_0(.din(w_dff_B_lShsHD8R7_0),.dout(w_dff_B_bkKN7mRm3_0),.clk(gclk));
	jdff dff_B_c3wEEVfN9_0(.din(w_dff_B_bkKN7mRm3_0),.dout(w_dff_B_c3wEEVfN9_0),.clk(gclk));
	jdff dff_B_BQqbw3445_0(.din(w_dff_B_c3wEEVfN9_0),.dout(w_dff_B_BQqbw3445_0),.clk(gclk));
	jdff dff_B_lwQ1oD6S9_0(.din(w_dff_B_BQqbw3445_0),.dout(w_dff_B_lwQ1oD6S9_0),.clk(gclk));
	jdff dff_B_y9Q5au4T4_0(.din(w_dff_B_lwQ1oD6S9_0),.dout(w_dff_B_y9Q5au4T4_0),.clk(gclk));
	jdff dff_B_DxK7zWo11_0(.din(w_dff_B_y9Q5au4T4_0),.dout(w_dff_B_DxK7zWo11_0),.clk(gclk));
	jdff dff_B_faQGBYKa9_0(.din(w_dff_B_DxK7zWo11_0),.dout(w_dff_B_faQGBYKa9_0),.clk(gclk));
	jdff dff_B_3I5pooTO7_0(.din(w_dff_B_faQGBYKa9_0),.dout(w_dff_B_3I5pooTO7_0),.clk(gclk));
	jdff dff_B_cfFB24pP0_0(.din(w_dff_B_3I5pooTO7_0),.dout(w_dff_B_cfFB24pP0_0),.clk(gclk));
	jdff dff_B_f9d0InF66_0(.din(w_dff_B_cfFB24pP0_0),.dout(w_dff_B_f9d0InF66_0),.clk(gclk));
	jdff dff_B_YbfPydN56_0(.din(w_dff_B_f9d0InF66_0),.dout(w_dff_B_YbfPydN56_0),.clk(gclk));
	jdff dff_B_K80VNsHQ9_0(.din(w_dff_B_YbfPydN56_0),.dout(w_dff_B_K80VNsHQ9_0),.clk(gclk));
	jdff dff_B_eu2N1W3a8_0(.din(w_dff_B_K80VNsHQ9_0),.dout(w_dff_B_eu2N1W3a8_0),.clk(gclk));
	jdff dff_B_h2MQXie50_0(.din(w_dff_B_eu2N1W3a8_0),.dout(w_dff_B_h2MQXie50_0),.clk(gclk));
	jdff dff_B_ikzr0D3R1_0(.din(w_dff_B_h2MQXie50_0),.dout(w_dff_B_ikzr0D3R1_0),.clk(gclk));
	jdff dff_B_8PARjvWG7_0(.din(w_dff_B_ikzr0D3R1_0),.dout(w_dff_B_8PARjvWG7_0),.clk(gclk));
	jdff dff_B_Svtva3j69_0(.din(w_dff_B_8PARjvWG7_0),.dout(w_dff_B_Svtva3j69_0),.clk(gclk));
	jdff dff_B_Q6D2xxis9_0(.din(w_dff_B_Svtva3j69_0),.dout(w_dff_B_Q6D2xxis9_0),.clk(gclk));
	jdff dff_B_Wu2J385L5_0(.din(w_dff_B_Q6D2xxis9_0),.dout(w_dff_B_Wu2J385L5_0),.clk(gclk));
	jdff dff_B_wGIDmibr0_0(.din(w_dff_B_Wu2J385L5_0),.dout(w_dff_B_wGIDmibr0_0),.clk(gclk));
	jdff dff_B_k2OEKT3Z2_0(.din(w_dff_B_wGIDmibr0_0),.dout(w_dff_B_k2OEKT3Z2_0),.clk(gclk));
	jdff dff_B_D44JhL0K2_0(.din(w_dff_B_k2OEKT3Z2_0),.dout(w_dff_B_D44JhL0K2_0),.clk(gclk));
	jdff dff_B_J0R6U13T8_0(.din(w_dff_B_D44JhL0K2_0),.dout(w_dff_B_J0R6U13T8_0),.clk(gclk));
	jdff dff_B_KaEd3tYK1_0(.din(w_dff_B_J0R6U13T8_0),.dout(w_dff_B_KaEd3tYK1_0),.clk(gclk));
	jdff dff_B_ayg7Z1Jg7_0(.din(w_dff_B_KaEd3tYK1_0),.dout(w_dff_B_ayg7Z1Jg7_0),.clk(gclk));
	jdff dff_B_7wKYrfz42_0(.din(w_dff_B_ayg7Z1Jg7_0),.dout(w_dff_B_7wKYrfz42_0),.clk(gclk));
	jdff dff_B_s1IFzW6e3_0(.din(w_dff_B_7wKYrfz42_0),.dout(w_dff_B_s1IFzW6e3_0),.clk(gclk));
	jdff dff_B_KpSIdnJ37_0(.din(w_dff_B_s1IFzW6e3_0),.dout(w_dff_B_KpSIdnJ37_0),.clk(gclk));
	jdff dff_B_h7OzLhJK2_0(.din(w_dff_B_KpSIdnJ37_0),.dout(w_dff_B_h7OzLhJK2_0),.clk(gclk));
	jdff dff_B_i0PS1ePd4_0(.din(w_dff_B_h7OzLhJK2_0),.dout(w_dff_B_i0PS1ePd4_0),.clk(gclk));
	jdff dff_B_td55wW7w2_0(.din(w_dff_B_i0PS1ePd4_0),.dout(w_dff_B_td55wW7w2_0),.clk(gclk));
	jdff dff_B_7IFs5pdC3_0(.din(w_dff_B_td55wW7w2_0),.dout(w_dff_B_7IFs5pdC3_0),.clk(gclk));
	jdff dff_B_xwjNpZHV8_0(.din(w_dff_B_7IFs5pdC3_0),.dout(w_dff_B_xwjNpZHV8_0),.clk(gclk));
	jdff dff_B_7dkg0NBF5_0(.din(w_dff_B_xwjNpZHV8_0),.dout(w_dff_B_7dkg0NBF5_0),.clk(gclk));
	jdff dff_B_4Qpql1583_0(.din(w_dff_B_7dkg0NBF5_0),.dout(w_dff_B_4Qpql1583_0),.clk(gclk));
	jdff dff_B_G0Ooledi7_0(.din(w_dff_B_4Qpql1583_0),.dout(w_dff_B_G0Ooledi7_0),.clk(gclk));
	jdff dff_B_mxh4ADsU8_0(.din(w_dff_B_G0Ooledi7_0),.dout(w_dff_B_mxh4ADsU8_0),.clk(gclk));
	jdff dff_B_8gkTUaR25_0(.din(w_dff_B_mxh4ADsU8_0),.dout(w_dff_B_8gkTUaR25_0),.clk(gclk));
	jdff dff_B_hSsav01T8_0(.din(w_dff_B_8gkTUaR25_0),.dout(w_dff_B_hSsav01T8_0),.clk(gclk));
	jdff dff_B_ExAZPzVT2_0(.din(w_dff_B_hSsav01T8_0),.dout(w_dff_B_ExAZPzVT2_0),.clk(gclk));
	jdff dff_B_NTBAdT9P8_0(.din(w_dff_B_ExAZPzVT2_0),.dout(w_dff_B_NTBAdT9P8_0),.clk(gclk));
	jdff dff_B_mqYykUGY5_0(.din(w_dff_B_NTBAdT9P8_0),.dout(w_dff_B_mqYykUGY5_0),.clk(gclk));
	jdff dff_B_NeAK7oRq0_0(.din(w_dff_B_mqYykUGY5_0),.dout(w_dff_B_NeAK7oRq0_0),.clk(gclk));
	jdff dff_B_D8ClRm555_0(.din(w_dff_B_NeAK7oRq0_0),.dout(w_dff_B_D8ClRm555_0),.clk(gclk));
	jdff dff_B_xQhJdJjm4_0(.din(w_dff_B_D8ClRm555_0),.dout(w_dff_B_xQhJdJjm4_0),.clk(gclk));
	jdff dff_B_GxAMHFJ85_0(.din(w_dff_B_xQhJdJjm4_0),.dout(w_dff_B_GxAMHFJ85_0),.clk(gclk));
	jdff dff_B_qCQkSwOJ7_0(.din(w_dff_B_GxAMHFJ85_0),.dout(w_dff_B_qCQkSwOJ7_0),.clk(gclk));
	jdff dff_B_U7lz97841_0(.din(w_dff_B_qCQkSwOJ7_0),.dout(w_dff_B_U7lz97841_0),.clk(gclk));
	jdff dff_B_bdOq4ceS9_0(.din(w_dff_B_U7lz97841_0),.dout(w_dff_B_bdOq4ceS9_0),.clk(gclk));
	jdff dff_B_2tHVEpgi4_0(.din(w_dff_B_bdOq4ceS9_0),.dout(w_dff_B_2tHVEpgi4_0),.clk(gclk));
	jdff dff_B_tQoTk3u53_0(.din(w_dff_B_2tHVEpgi4_0),.dout(w_dff_B_tQoTk3u53_0),.clk(gclk));
	jdff dff_B_k9QxEl460_0(.din(w_dff_B_tQoTk3u53_0),.dout(w_dff_B_k9QxEl460_0),.clk(gclk));
	jdff dff_B_sEuHC5Mo6_0(.din(w_dff_B_k9QxEl460_0),.dout(w_dff_B_sEuHC5Mo6_0),.clk(gclk));
	jdff dff_B_GinDUmHK9_0(.din(w_dff_B_sEuHC5Mo6_0),.dout(w_dff_B_GinDUmHK9_0),.clk(gclk));
	jdff dff_B_UZoZTpXC5_0(.din(w_dff_B_GinDUmHK9_0),.dout(w_dff_B_UZoZTpXC5_0),.clk(gclk));
	jdff dff_B_cENIvTQT9_0(.din(w_dff_B_UZoZTpXC5_0),.dout(w_dff_B_cENIvTQT9_0),.clk(gclk));
	jdff dff_B_f1xhoyIn4_0(.din(w_dff_B_cENIvTQT9_0),.dout(w_dff_B_f1xhoyIn4_0),.clk(gclk));
	jdff dff_B_gKQuFc3l4_0(.din(w_dff_B_f1xhoyIn4_0),.dout(w_dff_B_gKQuFc3l4_0),.clk(gclk));
	jdff dff_B_IklnBEV54_0(.din(w_dff_B_gKQuFc3l4_0),.dout(w_dff_B_IklnBEV54_0),.clk(gclk));
	jdff dff_B_4WXZG6qv3_0(.din(w_dff_B_IklnBEV54_0),.dout(w_dff_B_4WXZG6qv3_0),.clk(gclk));
	jdff dff_B_2QXrUTUd8_0(.din(w_dff_B_4WXZG6qv3_0),.dout(w_dff_B_2QXrUTUd8_0),.clk(gclk));
	jdff dff_B_BaobjH3z8_0(.din(w_dff_B_2QXrUTUd8_0),.dout(w_dff_B_BaobjH3z8_0),.clk(gclk));
	jdff dff_B_VbI1f1PP7_0(.din(w_dff_B_BaobjH3z8_0),.dout(w_dff_B_VbI1f1PP7_0),.clk(gclk));
	jdff dff_B_r9Uzvsxa5_0(.din(w_dff_B_VbI1f1PP7_0),.dout(w_dff_B_r9Uzvsxa5_0),.clk(gclk));
	jdff dff_B_yANSEPOJ6_0(.din(w_dff_B_r9Uzvsxa5_0),.dout(w_dff_B_yANSEPOJ6_0),.clk(gclk));
	jdff dff_B_QK4P1QL93_0(.din(w_dff_B_yANSEPOJ6_0),.dout(w_dff_B_QK4P1QL93_0),.clk(gclk));
	jdff dff_B_rtWKMnH03_0(.din(w_dff_B_QK4P1QL93_0),.dout(w_dff_B_rtWKMnH03_0),.clk(gclk));
	jdff dff_B_z2V96TGI1_0(.din(w_dff_B_rtWKMnH03_0),.dout(w_dff_B_z2V96TGI1_0),.clk(gclk));
	jdff dff_B_foUP6z4Q3_0(.din(w_dff_B_z2V96TGI1_0),.dout(w_dff_B_foUP6z4Q3_0),.clk(gclk));
	jdff dff_B_htV8mfbF1_0(.din(w_dff_B_foUP6z4Q3_0),.dout(w_dff_B_htV8mfbF1_0),.clk(gclk));
	jdff dff_B_ckD0w8RQ1_0(.din(w_dff_B_htV8mfbF1_0),.dout(w_dff_B_ckD0w8RQ1_0),.clk(gclk));
	jdff dff_B_34LSAjkY5_0(.din(w_dff_B_ckD0w8RQ1_0),.dout(w_dff_B_34LSAjkY5_0),.clk(gclk));
	jdff dff_B_I6ywWay94_0(.din(w_dff_B_34LSAjkY5_0),.dout(w_dff_B_I6ywWay94_0),.clk(gclk));
	jdff dff_B_RYCCcu415_0(.din(w_dff_B_I6ywWay94_0),.dout(w_dff_B_RYCCcu415_0),.clk(gclk));
	jdff dff_B_5VobtnOs3_0(.din(w_dff_B_RYCCcu415_0),.dout(w_dff_B_5VobtnOs3_0),.clk(gclk));
	jdff dff_B_mOQrCJ1g5_0(.din(w_dff_B_5VobtnOs3_0),.dout(w_dff_B_mOQrCJ1g5_0),.clk(gclk));
	jdff dff_B_hn22zHpw6_0(.din(w_dff_B_mOQrCJ1g5_0),.dout(w_dff_B_hn22zHpw6_0),.clk(gclk));
	jdff dff_B_OzpXqPiS3_0(.din(w_dff_B_hn22zHpw6_0),.dout(w_dff_B_OzpXqPiS3_0),.clk(gclk));
	jdff dff_B_op4UQWkT3_0(.din(w_dff_B_OzpXqPiS3_0),.dout(w_dff_B_op4UQWkT3_0),.clk(gclk));
	jdff dff_B_ropqRbhv4_0(.din(w_dff_B_op4UQWkT3_0),.dout(w_dff_B_ropqRbhv4_0),.clk(gclk));
	jdff dff_B_3oPLHGCN9_0(.din(w_dff_B_ropqRbhv4_0),.dout(w_dff_B_3oPLHGCN9_0),.clk(gclk));
	jdff dff_B_NYqGAdoD6_0(.din(w_dff_B_3oPLHGCN9_0),.dout(w_dff_B_NYqGAdoD6_0),.clk(gclk));
	jdff dff_B_woMA8ku71_0(.din(n952),.dout(w_dff_B_woMA8ku71_0),.clk(gclk));
	jdff dff_B_q0pQxjt75_0(.din(w_dff_B_woMA8ku71_0),.dout(w_dff_B_q0pQxjt75_0),.clk(gclk));
	jdff dff_B_naGqQuvO9_0(.din(w_dff_B_q0pQxjt75_0),.dout(w_dff_B_naGqQuvO9_0),.clk(gclk));
	jdff dff_B_I2oui9Xr6_0(.din(w_dff_B_naGqQuvO9_0),.dout(w_dff_B_I2oui9Xr6_0),.clk(gclk));
	jdff dff_B_SwzWSLWO7_0(.din(w_dff_B_I2oui9Xr6_0),.dout(w_dff_B_SwzWSLWO7_0),.clk(gclk));
	jdff dff_B_EpZcCx541_0(.din(w_dff_B_SwzWSLWO7_0),.dout(w_dff_B_EpZcCx541_0),.clk(gclk));
	jdff dff_B_M9fh4NkT3_0(.din(w_dff_B_EpZcCx541_0),.dout(w_dff_B_M9fh4NkT3_0),.clk(gclk));
	jdff dff_B_mHcw9xNn8_0(.din(w_dff_B_M9fh4NkT3_0),.dout(w_dff_B_mHcw9xNn8_0),.clk(gclk));
	jdff dff_B_ysMQwcks0_0(.din(w_dff_B_mHcw9xNn8_0),.dout(w_dff_B_ysMQwcks0_0),.clk(gclk));
	jdff dff_B_cIUo5hLy3_0(.din(w_dff_B_ysMQwcks0_0),.dout(w_dff_B_cIUo5hLy3_0),.clk(gclk));
	jdff dff_B_vb3gKBLM7_0(.din(w_dff_B_cIUo5hLy3_0),.dout(w_dff_B_vb3gKBLM7_0),.clk(gclk));
	jdff dff_B_gYVT3xAL8_0(.din(w_dff_B_vb3gKBLM7_0),.dout(w_dff_B_gYVT3xAL8_0),.clk(gclk));
	jdff dff_B_JGeRqTgp0_0(.din(w_dff_B_gYVT3xAL8_0),.dout(w_dff_B_JGeRqTgp0_0),.clk(gclk));
	jdff dff_B_f9vcm3833_0(.din(w_dff_B_JGeRqTgp0_0),.dout(w_dff_B_f9vcm3833_0),.clk(gclk));
	jdff dff_B_GLGQKuXA2_0(.din(w_dff_B_f9vcm3833_0),.dout(w_dff_B_GLGQKuXA2_0),.clk(gclk));
	jdff dff_B_hJxcmQD65_0(.din(w_dff_B_GLGQKuXA2_0),.dout(w_dff_B_hJxcmQD65_0),.clk(gclk));
	jdff dff_B_9KGl4FJm0_0(.din(w_dff_B_hJxcmQD65_0),.dout(w_dff_B_9KGl4FJm0_0),.clk(gclk));
	jdff dff_B_lwNpq0MP0_0(.din(w_dff_B_9KGl4FJm0_0),.dout(w_dff_B_lwNpq0MP0_0),.clk(gclk));
	jdff dff_B_teryKs1E9_0(.din(w_dff_B_lwNpq0MP0_0),.dout(w_dff_B_teryKs1E9_0),.clk(gclk));
	jdff dff_B_ROpempxJ7_0(.din(w_dff_B_teryKs1E9_0),.dout(w_dff_B_ROpempxJ7_0),.clk(gclk));
	jdff dff_B_atGRPXTu2_0(.din(w_dff_B_ROpempxJ7_0),.dout(w_dff_B_atGRPXTu2_0),.clk(gclk));
	jdff dff_B_b6Vmd6hu6_0(.din(w_dff_B_atGRPXTu2_0),.dout(w_dff_B_b6Vmd6hu6_0),.clk(gclk));
	jdff dff_B_xWQbYHu12_0(.din(w_dff_B_b6Vmd6hu6_0),.dout(w_dff_B_xWQbYHu12_0),.clk(gclk));
	jdff dff_B_MRurAhZu9_0(.din(w_dff_B_xWQbYHu12_0),.dout(w_dff_B_MRurAhZu9_0),.clk(gclk));
	jdff dff_B_KmfeMXeL1_0(.din(w_dff_B_MRurAhZu9_0),.dout(w_dff_B_KmfeMXeL1_0),.clk(gclk));
	jdff dff_B_B0RNuat01_0(.din(w_dff_B_KmfeMXeL1_0),.dout(w_dff_B_B0RNuat01_0),.clk(gclk));
	jdff dff_B_xgkKze5a9_0(.din(w_dff_B_B0RNuat01_0),.dout(w_dff_B_xgkKze5a9_0),.clk(gclk));
	jdff dff_B_LsEJxYeO3_0(.din(w_dff_B_xgkKze5a9_0),.dout(w_dff_B_LsEJxYeO3_0),.clk(gclk));
	jdff dff_B_2xberylD4_0(.din(w_dff_B_LsEJxYeO3_0),.dout(w_dff_B_2xberylD4_0),.clk(gclk));
	jdff dff_B_Wm3uww6j6_0(.din(w_dff_B_2xberylD4_0),.dout(w_dff_B_Wm3uww6j6_0),.clk(gclk));
	jdff dff_B_RdooBz740_0(.din(w_dff_B_Wm3uww6j6_0),.dout(w_dff_B_RdooBz740_0),.clk(gclk));
	jdff dff_B_rO48ehu66_0(.din(w_dff_B_RdooBz740_0),.dout(w_dff_B_rO48ehu66_0),.clk(gclk));
	jdff dff_B_AzJFvXw91_0(.din(w_dff_B_rO48ehu66_0),.dout(w_dff_B_AzJFvXw91_0),.clk(gclk));
	jdff dff_B_WrBPJO8w1_0(.din(w_dff_B_AzJFvXw91_0),.dout(w_dff_B_WrBPJO8w1_0),.clk(gclk));
	jdff dff_B_jfiZURSu5_0(.din(w_dff_B_WrBPJO8w1_0),.dout(w_dff_B_jfiZURSu5_0),.clk(gclk));
	jdff dff_B_dBqZMyST8_0(.din(w_dff_B_jfiZURSu5_0),.dout(w_dff_B_dBqZMyST8_0),.clk(gclk));
	jdff dff_B_SrYfIE7g4_0(.din(w_dff_B_dBqZMyST8_0),.dout(w_dff_B_SrYfIE7g4_0),.clk(gclk));
	jdff dff_B_6IN9eImK6_0(.din(w_dff_B_SrYfIE7g4_0),.dout(w_dff_B_6IN9eImK6_0),.clk(gclk));
	jdff dff_B_ScKd0CFw6_0(.din(w_dff_B_6IN9eImK6_0),.dout(w_dff_B_ScKd0CFw6_0),.clk(gclk));
	jdff dff_B_jN7t1Vlh5_0(.din(w_dff_B_ScKd0CFw6_0),.dout(w_dff_B_jN7t1Vlh5_0),.clk(gclk));
	jdff dff_B_9YeI7Kyf2_0(.din(w_dff_B_jN7t1Vlh5_0),.dout(w_dff_B_9YeI7Kyf2_0),.clk(gclk));
	jdff dff_B_v8tqkuBK2_0(.din(w_dff_B_9YeI7Kyf2_0),.dout(w_dff_B_v8tqkuBK2_0),.clk(gclk));
	jdff dff_B_AaTuoEnF4_0(.din(w_dff_B_v8tqkuBK2_0),.dout(w_dff_B_AaTuoEnF4_0),.clk(gclk));
	jdff dff_B_wPQSnwg69_0(.din(w_dff_B_AaTuoEnF4_0),.dout(w_dff_B_wPQSnwg69_0),.clk(gclk));
	jdff dff_B_1aNURhaJ6_0(.din(w_dff_B_wPQSnwg69_0),.dout(w_dff_B_1aNURhaJ6_0),.clk(gclk));
	jdff dff_B_7rLlObMg7_0(.din(w_dff_B_1aNURhaJ6_0),.dout(w_dff_B_7rLlObMg7_0),.clk(gclk));
	jdff dff_B_2RtrFZ1t1_0(.din(w_dff_B_7rLlObMg7_0),.dout(w_dff_B_2RtrFZ1t1_0),.clk(gclk));
	jdff dff_B_2WrZcO8O9_0(.din(w_dff_B_2RtrFZ1t1_0),.dout(w_dff_B_2WrZcO8O9_0),.clk(gclk));
	jdff dff_B_3jRpLMvD3_0(.din(w_dff_B_2WrZcO8O9_0),.dout(w_dff_B_3jRpLMvD3_0),.clk(gclk));
	jdff dff_B_hiPsxWSI4_0(.din(w_dff_B_3jRpLMvD3_0),.dout(w_dff_B_hiPsxWSI4_0),.clk(gclk));
	jdff dff_B_S7PtYfzw0_0(.din(w_dff_B_hiPsxWSI4_0),.dout(w_dff_B_S7PtYfzw0_0),.clk(gclk));
	jdff dff_B_jxVEOjI58_0(.din(w_dff_B_S7PtYfzw0_0),.dout(w_dff_B_jxVEOjI58_0),.clk(gclk));
	jdff dff_B_E1DGR5EH1_0(.din(w_dff_B_jxVEOjI58_0),.dout(w_dff_B_E1DGR5EH1_0),.clk(gclk));
	jdff dff_B_pVqGtZit6_0(.din(w_dff_B_E1DGR5EH1_0),.dout(w_dff_B_pVqGtZit6_0),.clk(gclk));
	jdff dff_B_Q5zWN9L96_0(.din(w_dff_B_pVqGtZit6_0),.dout(w_dff_B_Q5zWN9L96_0),.clk(gclk));
	jdff dff_B_hLOJOK031_0(.din(w_dff_B_Q5zWN9L96_0),.dout(w_dff_B_hLOJOK031_0),.clk(gclk));
	jdff dff_B_OBw3k05s3_0(.din(w_dff_B_hLOJOK031_0),.dout(w_dff_B_OBw3k05s3_0),.clk(gclk));
	jdff dff_B_mtmqLYXP7_0(.din(w_dff_B_OBw3k05s3_0),.dout(w_dff_B_mtmqLYXP7_0),.clk(gclk));
	jdff dff_B_nbM3Jkn44_0(.din(w_dff_B_mtmqLYXP7_0),.dout(w_dff_B_nbM3Jkn44_0),.clk(gclk));
	jdff dff_B_EMQIW3ku3_0(.din(w_dff_B_nbM3Jkn44_0),.dout(w_dff_B_EMQIW3ku3_0),.clk(gclk));
	jdff dff_B_MO27MXk02_0(.din(w_dff_B_EMQIW3ku3_0),.dout(w_dff_B_MO27MXk02_0),.clk(gclk));
	jdff dff_B_pNgJRW8u2_0(.din(w_dff_B_MO27MXk02_0),.dout(w_dff_B_pNgJRW8u2_0),.clk(gclk));
	jdff dff_B_S7QUpJyY1_0(.din(w_dff_B_pNgJRW8u2_0),.dout(w_dff_B_S7QUpJyY1_0),.clk(gclk));
	jdff dff_B_PKjSGtUM3_0(.din(w_dff_B_S7QUpJyY1_0),.dout(w_dff_B_PKjSGtUM3_0),.clk(gclk));
	jdff dff_B_S4E3W6KN6_0(.din(w_dff_B_PKjSGtUM3_0),.dout(w_dff_B_S4E3W6KN6_0),.clk(gclk));
	jdff dff_B_1nhqSAKw3_0(.din(w_dff_B_S4E3W6KN6_0),.dout(w_dff_B_1nhqSAKw3_0),.clk(gclk));
	jdff dff_B_YCGHBEaW3_0(.din(w_dff_B_1nhqSAKw3_0),.dout(w_dff_B_YCGHBEaW3_0),.clk(gclk));
	jdff dff_B_VEAuRrIs0_0(.din(w_dff_B_YCGHBEaW3_0),.dout(w_dff_B_VEAuRrIs0_0),.clk(gclk));
	jdff dff_B_1etwaut50_0(.din(w_dff_B_VEAuRrIs0_0),.dout(w_dff_B_1etwaut50_0),.clk(gclk));
	jdff dff_B_EEwoF9t74_0(.din(w_dff_B_1etwaut50_0),.dout(w_dff_B_EEwoF9t74_0),.clk(gclk));
	jdff dff_B_Cgg5vZzs0_0(.din(w_dff_B_EEwoF9t74_0),.dout(w_dff_B_Cgg5vZzs0_0),.clk(gclk));
	jdff dff_B_riVnUW115_0(.din(w_dff_B_Cgg5vZzs0_0),.dout(w_dff_B_riVnUW115_0),.clk(gclk));
	jdff dff_B_faeJll4c4_0(.din(w_dff_B_riVnUW115_0),.dout(w_dff_B_faeJll4c4_0),.clk(gclk));
	jdff dff_B_kr0Y06bI5_0(.din(w_dff_B_faeJll4c4_0),.dout(w_dff_B_kr0Y06bI5_0),.clk(gclk));
	jdff dff_B_TGDg4Fxd3_0(.din(w_dff_B_kr0Y06bI5_0),.dout(w_dff_B_TGDg4Fxd3_0),.clk(gclk));
	jdff dff_B_e7RI90VD9_0(.din(w_dff_B_TGDg4Fxd3_0),.dout(w_dff_B_e7RI90VD9_0),.clk(gclk));
	jdff dff_B_rxoS4dAY3_0(.din(w_dff_B_e7RI90VD9_0),.dout(w_dff_B_rxoS4dAY3_0),.clk(gclk));
	jdff dff_B_i0tfqvMv1_0(.din(w_dff_B_rxoS4dAY3_0),.dout(w_dff_B_i0tfqvMv1_0),.clk(gclk));
	jdff dff_B_Z1AMaSaV8_0(.din(w_dff_B_i0tfqvMv1_0),.dout(w_dff_B_Z1AMaSaV8_0),.clk(gclk));
	jdff dff_B_f6ZQH2494_0(.din(w_dff_B_Z1AMaSaV8_0),.dout(w_dff_B_f6ZQH2494_0),.clk(gclk));
	jdff dff_B_qbc8uBF02_0(.din(w_dff_B_f6ZQH2494_0),.dout(w_dff_B_qbc8uBF02_0),.clk(gclk));
	jdff dff_B_sykpQlV87_0(.din(w_dff_B_qbc8uBF02_0),.dout(w_dff_B_sykpQlV87_0),.clk(gclk));
	jdff dff_B_1vaM9zZZ1_0(.din(w_dff_B_sykpQlV87_0),.dout(w_dff_B_1vaM9zZZ1_0),.clk(gclk));
	jdff dff_B_szIUk8025_0(.din(w_dff_B_1vaM9zZZ1_0),.dout(w_dff_B_szIUk8025_0),.clk(gclk));
	jdff dff_B_xfmlBT012_0(.din(w_dff_B_szIUk8025_0),.dout(w_dff_B_xfmlBT012_0),.clk(gclk));
	jdff dff_B_qjDb8Fo38_0(.din(w_dff_B_xfmlBT012_0),.dout(w_dff_B_qjDb8Fo38_0),.clk(gclk));
	jdff dff_B_fwgvE4TM6_0(.din(w_dff_B_qjDb8Fo38_0),.dout(w_dff_B_fwgvE4TM6_0),.clk(gclk));
	jdff dff_B_VpZyQ5rH6_0(.din(w_dff_B_fwgvE4TM6_0),.dout(w_dff_B_VpZyQ5rH6_0),.clk(gclk));
	jdff dff_B_wOI1fQRM1_0(.din(w_dff_B_VpZyQ5rH6_0),.dout(w_dff_B_wOI1fQRM1_0),.clk(gclk));
	jdff dff_B_fH6asaQR3_0(.din(w_dff_B_wOI1fQRM1_0),.dout(w_dff_B_fH6asaQR3_0),.clk(gclk));
	jdff dff_B_1VBKnOCE2_0(.din(w_dff_B_fH6asaQR3_0),.dout(w_dff_B_1VBKnOCE2_0),.clk(gclk));
	jdff dff_B_4k1t9D9Y9_0(.din(w_dff_B_1VBKnOCE2_0),.dout(w_dff_B_4k1t9D9Y9_0),.clk(gclk));
	jdff dff_B_4MrxxEGB2_0(.din(w_dff_B_4k1t9D9Y9_0),.dout(w_dff_B_4MrxxEGB2_0),.clk(gclk));
	jdff dff_B_q5yKBMhs4_0(.din(w_dff_B_4MrxxEGB2_0),.dout(w_dff_B_q5yKBMhs4_0),.clk(gclk));
	jdff dff_B_2BOfN6Q42_0(.din(n958),.dout(w_dff_B_2BOfN6Q42_0),.clk(gclk));
	jdff dff_B_VBPAzVx42_0(.din(w_dff_B_2BOfN6Q42_0),.dout(w_dff_B_VBPAzVx42_0),.clk(gclk));
	jdff dff_B_ch7qP2NG1_0(.din(w_dff_B_VBPAzVx42_0),.dout(w_dff_B_ch7qP2NG1_0),.clk(gclk));
	jdff dff_B_RKgqDM6U0_0(.din(w_dff_B_ch7qP2NG1_0),.dout(w_dff_B_RKgqDM6U0_0),.clk(gclk));
	jdff dff_B_zStsKIT92_0(.din(w_dff_B_RKgqDM6U0_0),.dout(w_dff_B_zStsKIT92_0),.clk(gclk));
	jdff dff_B_iQLqDQQa3_0(.din(w_dff_B_zStsKIT92_0),.dout(w_dff_B_iQLqDQQa3_0),.clk(gclk));
	jdff dff_B_jqAhKNPr6_0(.din(w_dff_B_iQLqDQQa3_0),.dout(w_dff_B_jqAhKNPr6_0),.clk(gclk));
	jdff dff_B_vXuMHGEW4_0(.din(w_dff_B_jqAhKNPr6_0),.dout(w_dff_B_vXuMHGEW4_0),.clk(gclk));
	jdff dff_B_p9tLmpFF4_0(.din(w_dff_B_vXuMHGEW4_0),.dout(w_dff_B_p9tLmpFF4_0),.clk(gclk));
	jdff dff_B_iEAyHtIg5_0(.din(w_dff_B_p9tLmpFF4_0),.dout(w_dff_B_iEAyHtIg5_0),.clk(gclk));
	jdff dff_B_aEReYzTB6_0(.din(w_dff_B_iEAyHtIg5_0),.dout(w_dff_B_aEReYzTB6_0),.clk(gclk));
	jdff dff_B_QakGROrO1_0(.din(w_dff_B_aEReYzTB6_0),.dout(w_dff_B_QakGROrO1_0),.clk(gclk));
	jdff dff_B_HQk9F0Lb4_0(.din(w_dff_B_QakGROrO1_0),.dout(w_dff_B_HQk9F0Lb4_0),.clk(gclk));
	jdff dff_B_VWxzcZ9V8_0(.din(w_dff_B_HQk9F0Lb4_0),.dout(w_dff_B_VWxzcZ9V8_0),.clk(gclk));
	jdff dff_B_oyjkip7Q4_0(.din(w_dff_B_VWxzcZ9V8_0),.dout(w_dff_B_oyjkip7Q4_0),.clk(gclk));
	jdff dff_B_HymvBPt40_0(.din(w_dff_B_oyjkip7Q4_0),.dout(w_dff_B_HymvBPt40_0),.clk(gclk));
	jdff dff_B_V683s9sJ4_0(.din(w_dff_B_HymvBPt40_0),.dout(w_dff_B_V683s9sJ4_0),.clk(gclk));
	jdff dff_B_7p9o18fa3_0(.din(w_dff_B_V683s9sJ4_0),.dout(w_dff_B_7p9o18fa3_0),.clk(gclk));
	jdff dff_B_e7FJUkZD6_0(.din(w_dff_B_7p9o18fa3_0),.dout(w_dff_B_e7FJUkZD6_0),.clk(gclk));
	jdff dff_B_1MKuaGmE3_0(.din(w_dff_B_e7FJUkZD6_0),.dout(w_dff_B_1MKuaGmE3_0),.clk(gclk));
	jdff dff_B_t93lsMUY1_0(.din(w_dff_B_1MKuaGmE3_0),.dout(w_dff_B_t93lsMUY1_0),.clk(gclk));
	jdff dff_B_YoIkeLTo9_0(.din(w_dff_B_t93lsMUY1_0),.dout(w_dff_B_YoIkeLTo9_0),.clk(gclk));
	jdff dff_B_m7xcYI0O7_0(.din(w_dff_B_YoIkeLTo9_0),.dout(w_dff_B_m7xcYI0O7_0),.clk(gclk));
	jdff dff_B_2ZJhUVNi1_0(.din(w_dff_B_m7xcYI0O7_0),.dout(w_dff_B_2ZJhUVNi1_0),.clk(gclk));
	jdff dff_B_6UITKluf8_0(.din(w_dff_B_2ZJhUVNi1_0),.dout(w_dff_B_6UITKluf8_0),.clk(gclk));
	jdff dff_B_jJ0IIAdr6_0(.din(w_dff_B_6UITKluf8_0),.dout(w_dff_B_jJ0IIAdr6_0),.clk(gclk));
	jdff dff_B_e3sHNQI22_0(.din(w_dff_B_jJ0IIAdr6_0),.dout(w_dff_B_e3sHNQI22_0),.clk(gclk));
	jdff dff_B_rpCByu2K5_0(.din(w_dff_B_e3sHNQI22_0),.dout(w_dff_B_rpCByu2K5_0),.clk(gclk));
	jdff dff_B_UQJWJHC32_0(.din(w_dff_B_rpCByu2K5_0),.dout(w_dff_B_UQJWJHC32_0),.clk(gclk));
	jdff dff_B_9Ag1LGdL7_0(.din(w_dff_B_UQJWJHC32_0),.dout(w_dff_B_9Ag1LGdL7_0),.clk(gclk));
	jdff dff_B_DwXTjwsP2_0(.din(w_dff_B_9Ag1LGdL7_0),.dout(w_dff_B_DwXTjwsP2_0),.clk(gclk));
	jdff dff_B_aoUktpXP3_0(.din(w_dff_B_DwXTjwsP2_0),.dout(w_dff_B_aoUktpXP3_0),.clk(gclk));
	jdff dff_B_YxtDK2ns4_0(.din(w_dff_B_aoUktpXP3_0),.dout(w_dff_B_YxtDK2ns4_0),.clk(gclk));
	jdff dff_B_KzlEm6Bm6_0(.din(w_dff_B_YxtDK2ns4_0),.dout(w_dff_B_KzlEm6Bm6_0),.clk(gclk));
	jdff dff_B_ZpH52zS71_0(.din(w_dff_B_KzlEm6Bm6_0),.dout(w_dff_B_ZpH52zS71_0),.clk(gclk));
	jdff dff_B_sFUX0Vcj1_0(.din(w_dff_B_ZpH52zS71_0),.dout(w_dff_B_sFUX0Vcj1_0),.clk(gclk));
	jdff dff_B_lJORFGME9_0(.din(w_dff_B_sFUX0Vcj1_0),.dout(w_dff_B_lJORFGME9_0),.clk(gclk));
	jdff dff_B_yxViGg4Z0_0(.din(w_dff_B_lJORFGME9_0),.dout(w_dff_B_yxViGg4Z0_0),.clk(gclk));
	jdff dff_B_SLWZZrER1_0(.din(w_dff_B_yxViGg4Z0_0),.dout(w_dff_B_SLWZZrER1_0),.clk(gclk));
	jdff dff_B_n3tpDtvk4_0(.din(w_dff_B_SLWZZrER1_0),.dout(w_dff_B_n3tpDtvk4_0),.clk(gclk));
	jdff dff_B_KFl4aPQk8_0(.din(w_dff_B_n3tpDtvk4_0),.dout(w_dff_B_KFl4aPQk8_0),.clk(gclk));
	jdff dff_B_vLRY4kvG6_0(.din(w_dff_B_KFl4aPQk8_0),.dout(w_dff_B_vLRY4kvG6_0),.clk(gclk));
	jdff dff_B_vrhL2Odi7_0(.din(w_dff_B_vLRY4kvG6_0),.dout(w_dff_B_vrhL2Odi7_0),.clk(gclk));
	jdff dff_B_NZ9iKc2M8_0(.din(w_dff_B_vrhL2Odi7_0),.dout(w_dff_B_NZ9iKc2M8_0),.clk(gclk));
	jdff dff_B_DraEQZfK4_0(.din(w_dff_B_NZ9iKc2M8_0),.dout(w_dff_B_DraEQZfK4_0),.clk(gclk));
	jdff dff_B_x2KYQWpG7_0(.din(w_dff_B_DraEQZfK4_0),.dout(w_dff_B_x2KYQWpG7_0),.clk(gclk));
	jdff dff_B_RlqI4oeM9_0(.din(w_dff_B_x2KYQWpG7_0),.dout(w_dff_B_RlqI4oeM9_0),.clk(gclk));
	jdff dff_B_bAGEFQEV4_0(.din(w_dff_B_RlqI4oeM9_0),.dout(w_dff_B_bAGEFQEV4_0),.clk(gclk));
	jdff dff_B_NIXTqOCw7_0(.din(w_dff_B_bAGEFQEV4_0),.dout(w_dff_B_NIXTqOCw7_0),.clk(gclk));
	jdff dff_B_5SrNQhXs1_0(.din(w_dff_B_NIXTqOCw7_0),.dout(w_dff_B_5SrNQhXs1_0),.clk(gclk));
	jdff dff_B_82bX7yMC9_0(.din(w_dff_B_5SrNQhXs1_0),.dout(w_dff_B_82bX7yMC9_0),.clk(gclk));
	jdff dff_B_6WQrfXFa6_0(.din(w_dff_B_82bX7yMC9_0),.dout(w_dff_B_6WQrfXFa6_0),.clk(gclk));
	jdff dff_B_0KcfeBgc0_0(.din(w_dff_B_6WQrfXFa6_0),.dout(w_dff_B_0KcfeBgc0_0),.clk(gclk));
	jdff dff_B_jXUP2hUX2_0(.din(w_dff_B_0KcfeBgc0_0),.dout(w_dff_B_jXUP2hUX2_0),.clk(gclk));
	jdff dff_B_G2shiP8a3_0(.din(w_dff_B_jXUP2hUX2_0),.dout(w_dff_B_G2shiP8a3_0),.clk(gclk));
	jdff dff_B_gQgetMSG0_0(.din(w_dff_B_G2shiP8a3_0),.dout(w_dff_B_gQgetMSG0_0),.clk(gclk));
	jdff dff_B_vGY73Shj4_0(.din(w_dff_B_gQgetMSG0_0),.dout(w_dff_B_vGY73Shj4_0),.clk(gclk));
	jdff dff_B_x230VX6o2_0(.din(w_dff_B_vGY73Shj4_0),.dout(w_dff_B_x230VX6o2_0),.clk(gclk));
	jdff dff_B_ITSwtqNg0_0(.din(w_dff_B_x230VX6o2_0),.dout(w_dff_B_ITSwtqNg0_0),.clk(gclk));
	jdff dff_B_wMKWB4GX3_0(.din(w_dff_B_ITSwtqNg0_0),.dout(w_dff_B_wMKWB4GX3_0),.clk(gclk));
	jdff dff_B_PPVQVJ4W0_0(.din(w_dff_B_wMKWB4GX3_0),.dout(w_dff_B_PPVQVJ4W0_0),.clk(gclk));
	jdff dff_B_zW3vfONN5_0(.din(w_dff_B_PPVQVJ4W0_0),.dout(w_dff_B_zW3vfONN5_0),.clk(gclk));
	jdff dff_B_cQyTUBvz7_0(.din(w_dff_B_zW3vfONN5_0),.dout(w_dff_B_cQyTUBvz7_0),.clk(gclk));
	jdff dff_B_e46jy3lO4_0(.din(w_dff_B_cQyTUBvz7_0),.dout(w_dff_B_e46jy3lO4_0),.clk(gclk));
	jdff dff_B_Agii0MqL1_0(.din(w_dff_B_e46jy3lO4_0),.dout(w_dff_B_Agii0MqL1_0),.clk(gclk));
	jdff dff_B_KyY1UFWL3_0(.din(w_dff_B_Agii0MqL1_0),.dout(w_dff_B_KyY1UFWL3_0),.clk(gclk));
	jdff dff_B_MRn3By8s7_0(.din(w_dff_B_KyY1UFWL3_0),.dout(w_dff_B_MRn3By8s7_0),.clk(gclk));
	jdff dff_B_NzdugDE63_0(.din(w_dff_B_MRn3By8s7_0),.dout(w_dff_B_NzdugDE63_0),.clk(gclk));
	jdff dff_B_ds7bxBFr3_0(.din(w_dff_B_NzdugDE63_0),.dout(w_dff_B_ds7bxBFr3_0),.clk(gclk));
	jdff dff_B_Z8d4rzGQ8_0(.din(w_dff_B_ds7bxBFr3_0),.dout(w_dff_B_Z8d4rzGQ8_0),.clk(gclk));
	jdff dff_B_x7i2vxLV7_0(.din(w_dff_B_Z8d4rzGQ8_0),.dout(w_dff_B_x7i2vxLV7_0),.clk(gclk));
	jdff dff_B_0D5LiEID7_0(.din(w_dff_B_x7i2vxLV7_0),.dout(w_dff_B_0D5LiEID7_0),.clk(gclk));
	jdff dff_B_tv2RRyZy0_0(.din(w_dff_B_0D5LiEID7_0),.dout(w_dff_B_tv2RRyZy0_0),.clk(gclk));
	jdff dff_B_vIJigdPa0_0(.din(w_dff_B_tv2RRyZy0_0),.dout(w_dff_B_vIJigdPa0_0),.clk(gclk));
	jdff dff_B_N1hpe2jk4_0(.din(w_dff_B_vIJigdPa0_0),.dout(w_dff_B_N1hpe2jk4_0),.clk(gclk));
	jdff dff_B_gzoHAuVw1_0(.din(w_dff_B_N1hpe2jk4_0),.dout(w_dff_B_gzoHAuVw1_0),.clk(gclk));
	jdff dff_B_IdfMHzSF1_0(.din(w_dff_B_gzoHAuVw1_0),.dout(w_dff_B_IdfMHzSF1_0),.clk(gclk));
	jdff dff_B_8EiCbJMz0_0(.din(w_dff_B_IdfMHzSF1_0),.dout(w_dff_B_8EiCbJMz0_0),.clk(gclk));
	jdff dff_B_UQGyPA3k6_0(.din(w_dff_B_8EiCbJMz0_0),.dout(w_dff_B_UQGyPA3k6_0),.clk(gclk));
	jdff dff_B_hgTGGOc43_0(.din(w_dff_B_UQGyPA3k6_0),.dout(w_dff_B_hgTGGOc43_0),.clk(gclk));
	jdff dff_B_QpQdV85s5_0(.din(w_dff_B_hgTGGOc43_0),.dout(w_dff_B_QpQdV85s5_0),.clk(gclk));
	jdff dff_B_0Hoqw0ur1_0(.din(w_dff_B_QpQdV85s5_0),.dout(w_dff_B_0Hoqw0ur1_0),.clk(gclk));
	jdff dff_B_MwUmG7DW4_0(.din(w_dff_B_0Hoqw0ur1_0),.dout(w_dff_B_MwUmG7DW4_0),.clk(gclk));
	jdff dff_B_2zi5FKpx8_0(.din(w_dff_B_MwUmG7DW4_0),.dout(w_dff_B_2zi5FKpx8_0),.clk(gclk));
	jdff dff_B_0f1eobwe8_0(.din(w_dff_B_2zi5FKpx8_0),.dout(w_dff_B_0f1eobwe8_0),.clk(gclk));
	jdff dff_B_y052bCq92_0(.din(w_dff_B_0f1eobwe8_0),.dout(w_dff_B_y052bCq92_0),.clk(gclk));
	jdff dff_B_212jN4uS2_0(.din(w_dff_B_y052bCq92_0),.dout(w_dff_B_212jN4uS2_0),.clk(gclk));
	jdff dff_B_SwnPAFRO8_0(.din(w_dff_B_212jN4uS2_0),.dout(w_dff_B_SwnPAFRO8_0),.clk(gclk));
	jdff dff_B_eHmUQnW99_0(.din(w_dff_B_SwnPAFRO8_0),.dout(w_dff_B_eHmUQnW99_0),.clk(gclk));
	jdff dff_B_9nRjR8Ge1_0(.din(w_dff_B_eHmUQnW99_0),.dout(w_dff_B_9nRjR8Ge1_0),.clk(gclk));
	jdff dff_B_27INWU3O0_0(.din(w_dff_B_9nRjR8Ge1_0),.dout(w_dff_B_27INWU3O0_0),.clk(gclk));
	jdff dff_B_xcDE6JbJ4_0(.din(w_dff_B_27INWU3O0_0),.dout(w_dff_B_xcDE6JbJ4_0),.clk(gclk));
	jdff dff_B_35Zzwq683_0(.din(w_dff_B_xcDE6JbJ4_0),.dout(w_dff_B_35Zzwq683_0),.clk(gclk));
	jdff dff_B_tZHTz3T80_0(.din(w_dff_B_35Zzwq683_0),.dout(w_dff_B_tZHTz3T80_0),.clk(gclk));
	jdff dff_B_o3ojjpxb8_0(.din(w_dff_B_tZHTz3T80_0),.dout(w_dff_B_o3ojjpxb8_0),.clk(gclk));
	jdff dff_B_K3RS2WYq3_0(.din(n964),.dout(w_dff_B_K3RS2WYq3_0),.clk(gclk));
	jdff dff_B_4DRHh5WT2_0(.din(w_dff_B_K3RS2WYq3_0),.dout(w_dff_B_4DRHh5WT2_0),.clk(gclk));
	jdff dff_B_mSflLm8e5_0(.din(w_dff_B_4DRHh5WT2_0),.dout(w_dff_B_mSflLm8e5_0),.clk(gclk));
	jdff dff_B_DwvyECH30_0(.din(w_dff_B_mSflLm8e5_0),.dout(w_dff_B_DwvyECH30_0),.clk(gclk));
	jdff dff_B_7cyNYUos6_0(.din(w_dff_B_DwvyECH30_0),.dout(w_dff_B_7cyNYUos6_0),.clk(gclk));
	jdff dff_B_RVXe09fZ9_0(.din(w_dff_B_7cyNYUos6_0),.dout(w_dff_B_RVXe09fZ9_0),.clk(gclk));
	jdff dff_B_ShfkVBKY4_0(.din(w_dff_B_RVXe09fZ9_0),.dout(w_dff_B_ShfkVBKY4_0),.clk(gclk));
	jdff dff_B_uOBXALGU9_0(.din(w_dff_B_ShfkVBKY4_0),.dout(w_dff_B_uOBXALGU9_0),.clk(gclk));
	jdff dff_B_MGNhczvD5_0(.din(w_dff_B_uOBXALGU9_0),.dout(w_dff_B_MGNhczvD5_0),.clk(gclk));
	jdff dff_B_efcRf5aJ0_0(.din(w_dff_B_MGNhczvD5_0),.dout(w_dff_B_efcRf5aJ0_0),.clk(gclk));
	jdff dff_B_404BsHmB4_0(.din(w_dff_B_efcRf5aJ0_0),.dout(w_dff_B_404BsHmB4_0),.clk(gclk));
	jdff dff_B_ZJdyszo40_0(.din(w_dff_B_404BsHmB4_0),.dout(w_dff_B_ZJdyszo40_0),.clk(gclk));
	jdff dff_B_8zkucMzy0_0(.din(w_dff_B_ZJdyszo40_0),.dout(w_dff_B_8zkucMzy0_0),.clk(gclk));
	jdff dff_B_nrXNRODy9_0(.din(w_dff_B_8zkucMzy0_0),.dout(w_dff_B_nrXNRODy9_0),.clk(gclk));
	jdff dff_B_YTEajDhQ3_0(.din(w_dff_B_nrXNRODy9_0),.dout(w_dff_B_YTEajDhQ3_0),.clk(gclk));
	jdff dff_B_iufXdTah5_0(.din(w_dff_B_YTEajDhQ3_0),.dout(w_dff_B_iufXdTah5_0),.clk(gclk));
	jdff dff_B_wLLIM7pj7_0(.din(w_dff_B_iufXdTah5_0),.dout(w_dff_B_wLLIM7pj7_0),.clk(gclk));
	jdff dff_B_N8mw2iaZ6_0(.din(w_dff_B_wLLIM7pj7_0),.dout(w_dff_B_N8mw2iaZ6_0),.clk(gclk));
	jdff dff_B_I1xd5Q4t7_0(.din(w_dff_B_N8mw2iaZ6_0),.dout(w_dff_B_I1xd5Q4t7_0),.clk(gclk));
	jdff dff_B_OID3XpKU5_0(.din(w_dff_B_I1xd5Q4t7_0),.dout(w_dff_B_OID3XpKU5_0),.clk(gclk));
	jdff dff_B_zegGqo9K6_0(.din(w_dff_B_OID3XpKU5_0),.dout(w_dff_B_zegGqo9K6_0),.clk(gclk));
	jdff dff_B_BXAUWvT53_0(.din(w_dff_B_zegGqo9K6_0),.dout(w_dff_B_BXAUWvT53_0),.clk(gclk));
	jdff dff_B_OBBaTtj89_0(.din(w_dff_B_BXAUWvT53_0),.dout(w_dff_B_OBBaTtj89_0),.clk(gclk));
	jdff dff_B_mRCC0SPp1_0(.din(w_dff_B_OBBaTtj89_0),.dout(w_dff_B_mRCC0SPp1_0),.clk(gclk));
	jdff dff_B_0BCVMXHX7_0(.din(w_dff_B_mRCC0SPp1_0),.dout(w_dff_B_0BCVMXHX7_0),.clk(gclk));
	jdff dff_B_VD3swhdo6_0(.din(w_dff_B_0BCVMXHX7_0),.dout(w_dff_B_VD3swhdo6_0),.clk(gclk));
	jdff dff_B_aBjHiLyJ1_0(.din(w_dff_B_VD3swhdo6_0),.dout(w_dff_B_aBjHiLyJ1_0),.clk(gclk));
	jdff dff_B_ggOBYlC84_0(.din(w_dff_B_aBjHiLyJ1_0),.dout(w_dff_B_ggOBYlC84_0),.clk(gclk));
	jdff dff_B_cT2vDEWf8_0(.din(w_dff_B_ggOBYlC84_0),.dout(w_dff_B_cT2vDEWf8_0),.clk(gclk));
	jdff dff_B_ut9FwjEy7_0(.din(w_dff_B_cT2vDEWf8_0),.dout(w_dff_B_ut9FwjEy7_0),.clk(gclk));
	jdff dff_B_cK8zPTj01_0(.din(w_dff_B_ut9FwjEy7_0),.dout(w_dff_B_cK8zPTj01_0),.clk(gclk));
	jdff dff_B_RXPWPRzV5_0(.din(w_dff_B_cK8zPTj01_0),.dout(w_dff_B_RXPWPRzV5_0),.clk(gclk));
	jdff dff_B_kPeAOuBD7_0(.din(w_dff_B_RXPWPRzV5_0),.dout(w_dff_B_kPeAOuBD7_0),.clk(gclk));
	jdff dff_B_jyeDho8c0_0(.din(w_dff_B_kPeAOuBD7_0),.dout(w_dff_B_jyeDho8c0_0),.clk(gclk));
	jdff dff_B_uJdXKlai3_0(.din(w_dff_B_jyeDho8c0_0),.dout(w_dff_B_uJdXKlai3_0),.clk(gclk));
	jdff dff_B_xcaW26FH7_0(.din(w_dff_B_uJdXKlai3_0),.dout(w_dff_B_xcaW26FH7_0),.clk(gclk));
	jdff dff_B_T0Uq0v029_0(.din(w_dff_B_xcaW26FH7_0),.dout(w_dff_B_T0Uq0v029_0),.clk(gclk));
	jdff dff_B_34VbIJNH2_0(.din(w_dff_B_T0Uq0v029_0),.dout(w_dff_B_34VbIJNH2_0),.clk(gclk));
	jdff dff_B_0mp5ciba5_0(.din(w_dff_B_34VbIJNH2_0),.dout(w_dff_B_0mp5ciba5_0),.clk(gclk));
	jdff dff_B_wZxhmfKh1_0(.din(w_dff_B_0mp5ciba5_0),.dout(w_dff_B_wZxhmfKh1_0),.clk(gclk));
	jdff dff_B_oqJu9l2M4_0(.din(w_dff_B_wZxhmfKh1_0),.dout(w_dff_B_oqJu9l2M4_0),.clk(gclk));
	jdff dff_B_Yf6Y7Qkm6_0(.din(w_dff_B_oqJu9l2M4_0),.dout(w_dff_B_Yf6Y7Qkm6_0),.clk(gclk));
	jdff dff_B_VWqbhx1M7_0(.din(w_dff_B_Yf6Y7Qkm6_0),.dout(w_dff_B_VWqbhx1M7_0),.clk(gclk));
	jdff dff_B_kHA0vOpM4_0(.din(w_dff_B_VWqbhx1M7_0),.dout(w_dff_B_kHA0vOpM4_0),.clk(gclk));
	jdff dff_B_nzF5mTP21_0(.din(w_dff_B_kHA0vOpM4_0),.dout(w_dff_B_nzF5mTP21_0),.clk(gclk));
	jdff dff_B_mGRIYUKt8_0(.din(w_dff_B_nzF5mTP21_0),.dout(w_dff_B_mGRIYUKt8_0),.clk(gclk));
	jdff dff_B_FWkg8djd8_0(.din(w_dff_B_mGRIYUKt8_0),.dout(w_dff_B_FWkg8djd8_0),.clk(gclk));
	jdff dff_B_1OfimBcA7_0(.din(w_dff_B_FWkg8djd8_0),.dout(w_dff_B_1OfimBcA7_0),.clk(gclk));
	jdff dff_B_fx0rMpml0_0(.din(w_dff_B_1OfimBcA7_0),.dout(w_dff_B_fx0rMpml0_0),.clk(gclk));
	jdff dff_B_nJV9S1V85_0(.din(w_dff_B_fx0rMpml0_0),.dout(w_dff_B_nJV9S1V85_0),.clk(gclk));
	jdff dff_B_11Rp9fqm3_0(.din(w_dff_B_nJV9S1V85_0),.dout(w_dff_B_11Rp9fqm3_0),.clk(gclk));
	jdff dff_B_8m9eHZXG5_0(.din(w_dff_B_11Rp9fqm3_0),.dout(w_dff_B_8m9eHZXG5_0),.clk(gclk));
	jdff dff_B_6UM1RTYG6_0(.din(w_dff_B_8m9eHZXG5_0),.dout(w_dff_B_6UM1RTYG6_0),.clk(gclk));
	jdff dff_B_9YbEg9pz2_0(.din(w_dff_B_6UM1RTYG6_0),.dout(w_dff_B_9YbEg9pz2_0),.clk(gclk));
	jdff dff_B_Q2i4jHJO6_0(.din(w_dff_B_9YbEg9pz2_0),.dout(w_dff_B_Q2i4jHJO6_0),.clk(gclk));
	jdff dff_B_OznLmD8I1_0(.din(w_dff_B_Q2i4jHJO6_0),.dout(w_dff_B_OznLmD8I1_0),.clk(gclk));
	jdff dff_B_XKRgdknm6_0(.din(w_dff_B_OznLmD8I1_0),.dout(w_dff_B_XKRgdknm6_0),.clk(gclk));
	jdff dff_B_Ws4EjfI20_0(.din(w_dff_B_XKRgdknm6_0),.dout(w_dff_B_Ws4EjfI20_0),.clk(gclk));
	jdff dff_B_9i1h24cq5_0(.din(w_dff_B_Ws4EjfI20_0),.dout(w_dff_B_9i1h24cq5_0),.clk(gclk));
	jdff dff_B_DVy0fdLL7_0(.din(w_dff_B_9i1h24cq5_0),.dout(w_dff_B_DVy0fdLL7_0),.clk(gclk));
	jdff dff_B_JlFHpbuF3_0(.din(w_dff_B_DVy0fdLL7_0),.dout(w_dff_B_JlFHpbuF3_0),.clk(gclk));
	jdff dff_B_puJfkekU4_0(.din(w_dff_B_JlFHpbuF3_0),.dout(w_dff_B_puJfkekU4_0),.clk(gclk));
	jdff dff_B_JYGiK5QG0_0(.din(w_dff_B_puJfkekU4_0),.dout(w_dff_B_JYGiK5QG0_0),.clk(gclk));
	jdff dff_B_8yzjh6dk0_0(.din(w_dff_B_JYGiK5QG0_0),.dout(w_dff_B_8yzjh6dk0_0),.clk(gclk));
	jdff dff_B_9LrSMCjv1_0(.din(w_dff_B_8yzjh6dk0_0),.dout(w_dff_B_9LrSMCjv1_0),.clk(gclk));
	jdff dff_B_SkSkI2WZ1_0(.din(w_dff_B_9LrSMCjv1_0),.dout(w_dff_B_SkSkI2WZ1_0),.clk(gclk));
	jdff dff_B_uvsy7iJp5_0(.din(w_dff_B_SkSkI2WZ1_0),.dout(w_dff_B_uvsy7iJp5_0),.clk(gclk));
	jdff dff_B_VwIXG8d25_0(.din(w_dff_B_uvsy7iJp5_0),.dout(w_dff_B_VwIXG8d25_0),.clk(gclk));
	jdff dff_B_AkHjRKZN6_0(.din(w_dff_B_VwIXG8d25_0),.dout(w_dff_B_AkHjRKZN6_0),.clk(gclk));
	jdff dff_B_IZTrinxD5_0(.din(w_dff_B_AkHjRKZN6_0),.dout(w_dff_B_IZTrinxD5_0),.clk(gclk));
	jdff dff_B_XGyR95ZE2_0(.din(w_dff_B_IZTrinxD5_0),.dout(w_dff_B_XGyR95ZE2_0),.clk(gclk));
	jdff dff_B_leeQw8rV5_0(.din(w_dff_B_XGyR95ZE2_0),.dout(w_dff_B_leeQw8rV5_0),.clk(gclk));
	jdff dff_B_dbT628Vt1_0(.din(w_dff_B_leeQw8rV5_0),.dout(w_dff_B_dbT628Vt1_0),.clk(gclk));
	jdff dff_B_pwFhYqJa4_0(.din(w_dff_B_dbT628Vt1_0),.dout(w_dff_B_pwFhYqJa4_0),.clk(gclk));
	jdff dff_B_99DJbLNY6_0(.din(w_dff_B_pwFhYqJa4_0),.dout(w_dff_B_99DJbLNY6_0),.clk(gclk));
	jdff dff_B_BdhYscDh8_0(.din(w_dff_B_99DJbLNY6_0),.dout(w_dff_B_BdhYscDh8_0),.clk(gclk));
	jdff dff_B_fkXlF58S2_0(.din(w_dff_B_BdhYscDh8_0),.dout(w_dff_B_fkXlF58S2_0),.clk(gclk));
	jdff dff_B_fQiq6p2n4_0(.din(w_dff_B_fkXlF58S2_0),.dout(w_dff_B_fQiq6p2n4_0),.clk(gclk));
	jdff dff_B_eCA2PY434_0(.din(w_dff_B_fQiq6p2n4_0),.dout(w_dff_B_eCA2PY434_0),.clk(gclk));
	jdff dff_B_ldcyIKZa3_0(.din(w_dff_B_eCA2PY434_0),.dout(w_dff_B_ldcyIKZa3_0),.clk(gclk));
	jdff dff_B_4rXeWAsx1_0(.din(w_dff_B_ldcyIKZa3_0),.dout(w_dff_B_4rXeWAsx1_0),.clk(gclk));
	jdff dff_B_Z3uASZtT0_0(.din(w_dff_B_4rXeWAsx1_0),.dout(w_dff_B_Z3uASZtT0_0),.clk(gclk));
	jdff dff_B_gf7kSrln3_0(.din(w_dff_B_Z3uASZtT0_0),.dout(w_dff_B_gf7kSrln3_0),.clk(gclk));
	jdff dff_B_cgt4YXwf3_0(.din(w_dff_B_gf7kSrln3_0),.dout(w_dff_B_cgt4YXwf3_0),.clk(gclk));
	jdff dff_B_kjUTgarz4_0(.din(w_dff_B_cgt4YXwf3_0),.dout(w_dff_B_kjUTgarz4_0),.clk(gclk));
	jdff dff_B_DVUSMd3i4_0(.din(w_dff_B_kjUTgarz4_0),.dout(w_dff_B_DVUSMd3i4_0),.clk(gclk));
	jdff dff_B_5Er3MTwe5_0(.din(w_dff_B_DVUSMd3i4_0),.dout(w_dff_B_5Er3MTwe5_0),.clk(gclk));
	jdff dff_B_vOhFNWy42_0(.din(w_dff_B_5Er3MTwe5_0),.dout(w_dff_B_vOhFNWy42_0),.clk(gclk));
	jdff dff_B_5nUDXCC78_0(.din(w_dff_B_vOhFNWy42_0),.dout(w_dff_B_5nUDXCC78_0),.clk(gclk));
	jdff dff_B_7ldrUj3E3_0(.din(w_dff_B_5nUDXCC78_0),.dout(w_dff_B_7ldrUj3E3_0),.clk(gclk));
	jdff dff_B_Q9tuIgl56_0(.din(w_dff_B_7ldrUj3E3_0),.dout(w_dff_B_Q9tuIgl56_0),.clk(gclk));
	jdff dff_B_70D0ZeN33_0(.din(w_dff_B_Q9tuIgl56_0),.dout(w_dff_B_70D0ZeN33_0),.clk(gclk));
	jdff dff_B_IuMLLEF52_0(.din(w_dff_B_70D0ZeN33_0),.dout(w_dff_B_IuMLLEF52_0),.clk(gclk));
	jdff dff_B_rl0s45Hr5_0(.din(w_dff_B_IuMLLEF52_0),.dout(w_dff_B_rl0s45Hr5_0),.clk(gclk));
	jdff dff_B_nBOkQzRW5_0(.din(w_dff_B_rl0s45Hr5_0),.dout(w_dff_B_nBOkQzRW5_0),.clk(gclk));
	jdff dff_B_IwDOjdtB9_0(.din(w_dff_B_nBOkQzRW5_0),.dout(w_dff_B_IwDOjdtB9_0),.clk(gclk));
	jdff dff_B_zePLxlzP2_0(.din(n970),.dout(w_dff_B_zePLxlzP2_0),.clk(gclk));
	jdff dff_B_MrjC0Nsf0_0(.din(w_dff_B_zePLxlzP2_0),.dout(w_dff_B_MrjC0Nsf0_0),.clk(gclk));
	jdff dff_B_9BbWUDOQ9_0(.din(w_dff_B_MrjC0Nsf0_0),.dout(w_dff_B_9BbWUDOQ9_0),.clk(gclk));
	jdff dff_B_jkPyd1S97_0(.din(w_dff_B_9BbWUDOQ9_0),.dout(w_dff_B_jkPyd1S97_0),.clk(gclk));
	jdff dff_B_jvG7E53V9_0(.din(w_dff_B_jkPyd1S97_0),.dout(w_dff_B_jvG7E53V9_0),.clk(gclk));
	jdff dff_B_5Jo5qCoR7_0(.din(w_dff_B_jvG7E53V9_0),.dout(w_dff_B_5Jo5qCoR7_0),.clk(gclk));
	jdff dff_B_BYloEgoh5_0(.din(w_dff_B_5Jo5qCoR7_0),.dout(w_dff_B_BYloEgoh5_0),.clk(gclk));
	jdff dff_B_W53dzSHP3_0(.din(w_dff_B_BYloEgoh5_0),.dout(w_dff_B_W53dzSHP3_0),.clk(gclk));
	jdff dff_B_RzY5B0Ih6_0(.din(w_dff_B_W53dzSHP3_0),.dout(w_dff_B_RzY5B0Ih6_0),.clk(gclk));
	jdff dff_B_nXhlz6th7_0(.din(w_dff_B_RzY5B0Ih6_0),.dout(w_dff_B_nXhlz6th7_0),.clk(gclk));
	jdff dff_B_4ommtaw37_0(.din(w_dff_B_nXhlz6th7_0),.dout(w_dff_B_4ommtaw37_0),.clk(gclk));
	jdff dff_B_5QIuwX2U4_0(.din(w_dff_B_4ommtaw37_0),.dout(w_dff_B_5QIuwX2U4_0),.clk(gclk));
	jdff dff_B_qZB9Bp031_0(.din(w_dff_B_5QIuwX2U4_0),.dout(w_dff_B_qZB9Bp031_0),.clk(gclk));
	jdff dff_B_bofmnyac9_0(.din(w_dff_B_qZB9Bp031_0),.dout(w_dff_B_bofmnyac9_0),.clk(gclk));
	jdff dff_B_N6cgR2tm7_0(.din(w_dff_B_bofmnyac9_0),.dout(w_dff_B_N6cgR2tm7_0),.clk(gclk));
	jdff dff_B_OE2ZdGDa7_0(.din(w_dff_B_N6cgR2tm7_0),.dout(w_dff_B_OE2ZdGDa7_0),.clk(gclk));
	jdff dff_B_HgEHpkiR6_0(.din(w_dff_B_OE2ZdGDa7_0),.dout(w_dff_B_HgEHpkiR6_0),.clk(gclk));
	jdff dff_B_bW5lx9K62_0(.din(w_dff_B_HgEHpkiR6_0),.dout(w_dff_B_bW5lx9K62_0),.clk(gclk));
	jdff dff_B_wL4lbu5R9_0(.din(w_dff_B_bW5lx9K62_0),.dout(w_dff_B_wL4lbu5R9_0),.clk(gclk));
	jdff dff_B_2HSkl1IC8_0(.din(w_dff_B_wL4lbu5R9_0),.dout(w_dff_B_2HSkl1IC8_0),.clk(gclk));
	jdff dff_B_36IAP31z6_0(.din(w_dff_B_2HSkl1IC8_0),.dout(w_dff_B_36IAP31z6_0),.clk(gclk));
	jdff dff_B_iK5aSvpx3_0(.din(w_dff_B_36IAP31z6_0),.dout(w_dff_B_iK5aSvpx3_0),.clk(gclk));
	jdff dff_B_Gejfezgl4_0(.din(w_dff_B_iK5aSvpx3_0),.dout(w_dff_B_Gejfezgl4_0),.clk(gclk));
	jdff dff_B_dpREpI1S1_0(.din(w_dff_B_Gejfezgl4_0),.dout(w_dff_B_dpREpI1S1_0),.clk(gclk));
	jdff dff_B_xYMoj03v2_0(.din(w_dff_B_dpREpI1S1_0),.dout(w_dff_B_xYMoj03v2_0),.clk(gclk));
	jdff dff_B_x5s7SwfV5_0(.din(w_dff_B_xYMoj03v2_0),.dout(w_dff_B_x5s7SwfV5_0),.clk(gclk));
	jdff dff_B_2fiKOFhJ7_0(.din(w_dff_B_x5s7SwfV5_0),.dout(w_dff_B_2fiKOFhJ7_0),.clk(gclk));
	jdff dff_B_ozZFYezY5_0(.din(w_dff_B_2fiKOFhJ7_0),.dout(w_dff_B_ozZFYezY5_0),.clk(gclk));
	jdff dff_B_LGvLSvvD5_0(.din(w_dff_B_ozZFYezY5_0),.dout(w_dff_B_LGvLSvvD5_0),.clk(gclk));
	jdff dff_B_bZi1lRHb1_0(.din(w_dff_B_LGvLSvvD5_0),.dout(w_dff_B_bZi1lRHb1_0),.clk(gclk));
	jdff dff_B_ff5GhsKM6_0(.din(w_dff_B_bZi1lRHb1_0),.dout(w_dff_B_ff5GhsKM6_0),.clk(gclk));
	jdff dff_B_ZdVKEATP0_0(.din(w_dff_B_ff5GhsKM6_0),.dout(w_dff_B_ZdVKEATP0_0),.clk(gclk));
	jdff dff_B_UZdRAZsF9_0(.din(w_dff_B_ZdVKEATP0_0),.dout(w_dff_B_UZdRAZsF9_0),.clk(gclk));
	jdff dff_B_GsetXVEG7_0(.din(w_dff_B_UZdRAZsF9_0),.dout(w_dff_B_GsetXVEG7_0),.clk(gclk));
	jdff dff_B_38BnUpEY1_0(.din(w_dff_B_GsetXVEG7_0),.dout(w_dff_B_38BnUpEY1_0),.clk(gclk));
	jdff dff_B_vwLiHdnA7_0(.din(w_dff_B_38BnUpEY1_0),.dout(w_dff_B_vwLiHdnA7_0),.clk(gclk));
	jdff dff_B_elyoLX7k0_0(.din(w_dff_B_vwLiHdnA7_0),.dout(w_dff_B_elyoLX7k0_0),.clk(gclk));
	jdff dff_B_r45bNTik4_0(.din(w_dff_B_elyoLX7k0_0),.dout(w_dff_B_r45bNTik4_0),.clk(gclk));
	jdff dff_B_wQU9GMd80_0(.din(w_dff_B_r45bNTik4_0),.dout(w_dff_B_wQU9GMd80_0),.clk(gclk));
	jdff dff_B_9G1Awdc28_0(.din(w_dff_B_wQU9GMd80_0),.dout(w_dff_B_9G1Awdc28_0),.clk(gclk));
	jdff dff_B_yWAJKTy82_0(.din(w_dff_B_9G1Awdc28_0),.dout(w_dff_B_yWAJKTy82_0),.clk(gclk));
	jdff dff_B_x1qxu2m24_0(.din(w_dff_B_yWAJKTy82_0),.dout(w_dff_B_x1qxu2m24_0),.clk(gclk));
	jdff dff_B_sTDLdOkr7_0(.din(w_dff_B_x1qxu2m24_0),.dout(w_dff_B_sTDLdOkr7_0),.clk(gclk));
	jdff dff_B_mMr1X3771_0(.din(w_dff_B_sTDLdOkr7_0),.dout(w_dff_B_mMr1X3771_0),.clk(gclk));
	jdff dff_B_VrrlWfUi7_0(.din(w_dff_B_mMr1X3771_0),.dout(w_dff_B_VrrlWfUi7_0),.clk(gclk));
	jdff dff_B_ZOYtTr2Y4_0(.din(w_dff_B_VrrlWfUi7_0),.dout(w_dff_B_ZOYtTr2Y4_0),.clk(gclk));
	jdff dff_B_iyWXhSBQ3_0(.din(w_dff_B_ZOYtTr2Y4_0),.dout(w_dff_B_iyWXhSBQ3_0),.clk(gclk));
	jdff dff_B_D0Xw5fND1_0(.din(w_dff_B_iyWXhSBQ3_0),.dout(w_dff_B_D0Xw5fND1_0),.clk(gclk));
	jdff dff_B_3jIFMp7Q2_0(.din(w_dff_B_D0Xw5fND1_0),.dout(w_dff_B_3jIFMp7Q2_0),.clk(gclk));
	jdff dff_B_mcjqYnyk6_0(.din(w_dff_B_3jIFMp7Q2_0),.dout(w_dff_B_mcjqYnyk6_0),.clk(gclk));
	jdff dff_B_9aVcTZ3Y9_0(.din(w_dff_B_mcjqYnyk6_0),.dout(w_dff_B_9aVcTZ3Y9_0),.clk(gclk));
	jdff dff_B_FpwJ6Q869_0(.din(w_dff_B_9aVcTZ3Y9_0),.dout(w_dff_B_FpwJ6Q869_0),.clk(gclk));
	jdff dff_B_w8O0C1gR8_0(.din(w_dff_B_FpwJ6Q869_0),.dout(w_dff_B_w8O0C1gR8_0),.clk(gclk));
	jdff dff_B_StbFnvXe7_0(.din(w_dff_B_w8O0C1gR8_0),.dout(w_dff_B_StbFnvXe7_0),.clk(gclk));
	jdff dff_B_TEAACXXo2_0(.din(w_dff_B_StbFnvXe7_0),.dout(w_dff_B_TEAACXXo2_0),.clk(gclk));
	jdff dff_B_kw2VL7qC3_0(.din(w_dff_B_TEAACXXo2_0),.dout(w_dff_B_kw2VL7qC3_0),.clk(gclk));
	jdff dff_B_bnlnVv9T9_0(.din(w_dff_B_kw2VL7qC3_0),.dout(w_dff_B_bnlnVv9T9_0),.clk(gclk));
	jdff dff_B_Odk6xkZY2_0(.din(w_dff_B_bnlnVv9T9_0),.dout(w_dff_B_Odk6xkZY2_0),.clk(gclk));
	jdff dff_B_wK6zk5NY4_0(.din(w_dff_B_Odk6xkZY2_0),.dout(w_dff_B_wK6zk5NY4_0),.clk(gclk));
	jdff dff_B_4eyLIK714_0(.din(w_dff_B_wK6zk5NY4_0),.dout(w_dff_B_4eyLIK714_0),.clk(gclk));
	jdff dff_B_enxBNapu3_0(.din(w_dff_B_4eyLIK714_0),.dout(w_dff_B_enxBNapu3_0),.clk(gclk));
	jdff dff_B_ARkgyqWn6_0(.din(w_dff_B_enxBNapu3_0),.dout(w_dff_B_ARkgyqWn6_0),.clk(gclk));
	jdff dff_B_aEspfCFZ7_0(.din(w_dff_B_ARkgyqWn6_0),.dout(w_dff_B_aEspfCFZ7_0),.clk(gclk));
	jdff dff_B_tADwWlsu9_0(.din(w_dff_B_aEspfCFZ7_0),.dout(w_dff_B_tADwWlsu9_0),.clk(gclk));
	jdff dff_B_x73SyZpA3_0(.din(w_dff_B_tADwWlsu9_0),.dout(w_dff_B_x73SyZpA3_0),.clk(gclk));
	jdff dff_B_s8VjViHO6_0(.din(w_dff_B_x73SyZpA3_0),.dout(w_dff_B_s8VjViHO6_0),.clk(gclk));
	jdff dff_B_lggMrUCL2_0(.din(w_dff_B_s8VjViHO6_0),.dout(w_dff_B_lggMrUCL2_0),.clk(gclk));
	jdff dff_B_pN0pcOoO4_0(.din(w_dff_B_lggMrUCL2_0),.dout(w_dff_B_pN0pcOoO4_0),.clk(gclk));
	jdff dff_B_zAf7mVbR5_0(.din(w_dff_B_pN0pcOoO4_0),.dout(w_dff_B_zAf7mVbR5_0),.clk(gclk));
	jdff dff_B_KZq9pLel7_0(.din(w_dff_B_zAf7mVbR5_0),.dout(w_dff_B_KZq9pLel7_0),.clk(gclk));
	jdff dff_B_rzJcUxmw4_0(.din(w_dff_B_KZq9pLel7_0),.dout(w_dff_B_rzJcUxmw4_0),.clk(gclk));
	jdff dff_B_fcTx2uAt0_0(.din(w_dff_B_rzJcUxmw4_0),.dout(w_dff_B_fcTx2uAt0_0),.clk(gclk));
	jdff dff_B_sqP8r64f5_0(.din(w_dff_B_fcTx2uAt0_0),.dout(w_dff_B_sqP8r64f5_0),.clk(gclk));
	jdff dff_B_RGgWpfJX5_0(.din(w_dff_B_sqP8r64f5_0),.dout(w_dff_B_RGgWpfJX5_0),.clk(gclk));
	jdff dff_B_FGsJKvD37_0(.din(w_dff_B_RGgWpfJX5_0),.dout(w_dff_B_FGsJKvD37_0),.clk(gclk));
	jdff dff_B_AW3xLrzy1_0(.din(w_dff_B_FGsJKvD37_0),.dout(w_dff_B_AW3xLrzy1_0),.clk(gclk));
	jdff dff_B_OI2C8o5U0_0(.din(w_dff_B_AW3xLrzy1_0),.dout(w_dff_B_OI2C8o5U0_0),.clk(gclk));
	jdff dff_B_RBkikNet9_0(.din(w_dff_B_OI2C8o5U0_0),.dout(w_dff_B_RBkikNet9_0),.clk(gclk));
	jdff dff_B_n9rM7yTo3_0(.din(w_dff_B_RBkikNet9_0),.dout(w_dff_B_n9rM7yTo3_0),.clk(gclk));
	jdff dff_B_Ku1mdLTr4_0(.din(w_dff_B_n9rM7yTo3_0),.dout(w_dff_B_Ku1mdLTr4_0),.clk(gclk));
	jdff dff_B_wmDNkcw54_0(.din(w_dff_B_Ku1mdLTr4_0),.dout(w_dff_B_wmDNkcw54_0),.clk(gclk));
	jdff dff_B_ZOuSm1ZR2_0(.din(w_dff_B_wmDNkcw54_0),.dout(w_dff_B_ZOuSm1ZR2_0),.clk(gclk));
	jdff dff_B_pmPJUOSx3_0(.din(w_dff_B_ZOuSm1ZR2_0),.dout(w_dff_B_pmPJUOSx3_0),.clk(gclk));
	jdff dff_B_OHhZ9ZR25_0(.din(w_dff_B_pmPJUOSx3_0),.dout(w_dff_B_OHhZ9ZR25_0),.clk(gclk));
	jdff dff_B_PMhGhtTo9_0(.din(w_dff_B_OHhZ9ZR25_0),.dout(w_dff_B_PMhGhtTo9_0),.clk(gclk));
	jdff dff_B_kVKoFsj77_0(.din(w_dff_B_PMhGhtTo9_0),.dout(w_dff_B_kVKoFsj77_0),.clk(gclk));
	jdff dff_B_EGEXzWU93_0(.din(w_dff_B_kVKoFsj77_0),.dout(w_dff_B_EGEXzWU93_0),.clk(gclk));
	jdff dff_B_1OCYNory6_0(.din(w_dff_B_EGEXzWU93_0),.dout(w_dff_B_1OCYNory6_0),.clk(gclk));
	jdff dff_B_nr5bGOBE5_0(.din(w_dff_B_1OCYNory6_0),.dout(w_dff_B_nr5bGOBE5_0),.clk(gclk));
	jdff dff_B_ELDzrqbW5_0(.din(w_dff_B_nr5bGOBE5_0),.dout(w_dff_B_ELDzrqbW5_0),.clk(gclk));
	jdff dff_B_TQAXlIAK4_0(.din(w_dff_B_ELDzrqbW5_0),.dout(w_dff_B_TQAXlIAK4_0),.clk(gclk));
	jdff dff_B_DhS8Ndcu3_0(.din(w_dff_B_TQAXlIAK4_0),.dout(w_dff_B_DhS8Ndcu3_0),.clk(gclk));
	jdff dff_B_uh6izZ3S4_0(.din(w_dff_B_DhS8Ndcu3_0),.dout(w_dff_B_uh6izZ3S4_0),.clk(gclk));
	jdff dff_B_AYDG4Pbd6_0(.din(w_dff_B_uh6izZ3S4_0),.dout(w_dff_B_AYDG4Pbd6_0),.clk(gclk));
	jdff dff_B_fvzIQwTD7_0(.din(w_dff_B_AYDG4Pbd6_0),.dout(w_dff_B_fvzIQwTD7_0),.clk(gclk));
	jdff dff_B_ulGJImFW4_0(.din(w_dff_B_fvzIQwTD7_0),.dout(w_dff_B_ulGJImFW4_0),.clk(gclk));
	jdff dff_B_vwMgjcE08_0(.din(w_dff_B_ulGJImFW4_0),.dout(w_dff_B_vwMgjcE08_0),.clk(gclk));
	jdff dff_B_RUcxmNUm8_0(.din(n976),.dout(w_dff_B_RUcxmNUm8_0),.clk(gclk));
	jdff dff_B_uSh4msnA3_0(.din(w_dff_B_RUcxmNUm8_0),.dout(w_dff_B_uSh4msnA3_0),.clk(gclk));
	jdff dff_B_jCAhsPsG8_0(.din(w_dff_B_uSh4msnA3_0),.dout(w_dff_B_jCAhsPsG8_0),.clk(gclk));
	jdff dff_B_Q0DEtEDD9_0(.din(w_dff_B_jCAhsPsG8_0),.dout(w_dff_B_Q0DEtEDD9_0),.clk(gclk));
	jdff dff_B_xGzCzgYc1_0(.din(w_dff_B_Q0DEtEDD9_0),.dout(w_dff_B_xGzCzgYc1_0),.clk(gclk));
	jdff dff_B_47OiT29x9_0(.din(w_dff_B_xGzCzgYc1_0),.dout(w_dff_B_47OiT29x9_0),.clk(gclk));
	jdff dff_B_sjIkIasD6_0(.din(w_dff_B_47OiT29x9_0),.dout(w_dff_B_sjIkIasD6_0),.clk(gclk));
	jdff dff_B_HL4vSb0i3_0(.din(w_dff_B_sjIkIasD6_0),.dout(w_dff_B_HL4vSb0i3_0),.clk(gclk));
	jdff dff_B_GEubLeZ76_0(.din(w_dff_B_HL4vSb0i3_0),.dout(w_dff_B_GEubLeZ76_0),.clk(gclk));
	jdff dff_B_eGuVSfhE3_0(.din(w_dff_B_GEubLeZ76_0),.dout(w_dff_B_eGuVSfhE3_0),.clk(gclk));
	jdff dff_B_mWzpjlr73_0(.din(w_dff_B_eGuVSfhE3_0),.dout(w_dff_B_mWzpjlr73_0),.clk(gclk));
	jdff dff_B_pPKBXpYt4_0(.din(w_dff_B_mWzpjlr73_0),.dout(w_dff_B_pPKBXpYt4_0),.clk(gclk));
	jdff dff_B_ZKo11Bso6_0(.din(w_dff_B_pPKBXpYt4_0),.dout(w_dff_B_ZKo11Bso6_0),.clk(gclk));
	jdff dff_B_1xSGfU5p7_0(.din(w_dff_B_ZKo11Bso6_0),.dout(w_dff_B_1xSGfU5p7_0),.clk(gclk));
	jdff dff_B_oZEFHgBT9_0(.din(w_dff_B_1xSGfU5p7_0),.dout(w_dff_B_oZEFHgBT9_0),.clk(gclk));
	jdff dff_B_rizs14Rv1_0(.din(w_dff_B_oZEFHgBT9_0),.dout(w_dff_B_rizs14Rv1_0),.clk(gclk));
	jdff dff_B_3Vr6j7Op8_0(.din(w_dff_B_rizs14Rv1_0),.dout(w_dff_B_3Vr6j7Op8_0),.clk(gclk));
	jdff dff_B_rCzTFrsx2_0(.din(w_dff_B_3Vr6j7Op8_0),.dout(w_dff_B_rCzTFrsx2_0),.clk(gclk));
	jdff dff_B_SrrZ8mhG1_0(.din(w_dff_B_rCzTFrsx2_0),.dout(w_dff_B_SrrZ8mhG1_0),.clk(gclk));
	jdff dff_B_mnuMK0k33_0(.din(w_dff_B_SrrZ8mhG1_0),.dout(w_dff_B_mnuMK0k33_0),.clk(gclk));
	jdff dff_B_w3hqzGoA0_0(.din(w_dff_B_mnuMK0k33_0),.dout(w_dff_B_w3hqzGoA0_0),.clk(gclk));
	jdff dff_B_0TK6Qbt07_0(.din(w_dff_B_w3hqzGoA0_0),.dout(w_dff_B_0TK6Qbt07_0),.clk(gclk));
	jdff dff_B_pHykt49I6_0(.din(w_dff_B_0TK6Qbt07_0),.dout(w_dff_B_pHykt49I6_0),.clk(gclk));
	jdff dff_B_utkvrmZc7_0(.din(w_dff_B_pHykt49I6_0),.dout(w_dff_B_utkvrmZc7_0),.clk(gclk));
	jdff dff_B_DkLiLsCZ5_0(.din(w_dff_B_utkvrmZc7_0),.dout(w_dff_B_DkLiLsCZ5_0),.clk(gclk));
	jdff dff_B_g23GuXx38_0(.din(w_dff_B_DkLiLsCZ5_0),.dout(w_dff_B_g23GuXx38_0),.clk(gclk));
	jdff dff_B_hZb0JHan7_0(.din(w_dff_B_g23GuXx38_0),.dout(w_dff_B_hZb0JHan7_0),.clk(gclk));
	jdff dff_B_Bx7CoowZ0_0(.din(w_dff_B_hZb0JHan7_0),.dout(w_dff_B_Bx7CoowZ0_0),.clk(gclk));
	jdff dff_B_X2L28eJj8_0(.din(w_dff_B_Bx7CoowZ0_0),.dout(w_dff_B_X2L28eJj8_0),.clk(gclk));
	jdff dff_B_eRGJXM1a2_0(.din(w_dff_B_X2L28eJj8_0),.dout(w_dff_B_eRGJXM1a2_0),.clk(gclk));
	jdff dff_B_23mVQqz58_0(.din(w_dff_B_eRGJXM1a2_0),.dout(w_dff_B_23mVQqz58_0),.clk(gclk));
	jdff dff_B_xnHP6Dda9_0(.din(w_dff_B_23mVQqz58_0),.dout(w_dff_B_xnHP6Dda9_0),.clk(gclk));
	jdff dff_B_cf45dtR64_0(.din(w_dff_B_xnHP6Dda9_0),.dout(w_dff_B_cf45dtR64_0),.clk(gclk));
	jdff dff_B_lLthOjPU7_0(.din(w_dff_B_cf45dtR64_0),.dout(w_dff_B_lLthOjPU7_0),.clk(gclk));
	jdff dff_B_80iKDJKN0_0(.din(w_dff_B_lLthOjPU7_0),.dout(w_dff_B_80iKDJKN0_0),.clk(gclk));
	jdff dff_B_vC3WVPAy4_0(.din(w_dff_B_80iKDJKN0_0),.dout(w_dff_B_vC3WVPAy4_0),.clk(gclk));
	jdff dff_B_iUbw8r529_0(.din(w_dff_B_vC3WVPAy4_0),.dout(w_dff_B_iUbw8r529_0),.clk(gclk));
	jdff dff_B_qVWscI2K4_0(.din(w_dff_B_iUbw8r529_0),.dout(w_dff_B_qVWscI2K4_0),.clk(gclk));
	jdff dff_B_UiUFMzzk8_0(.din(w_dff_B_qVWscI2K4_0),.dout(w_dff_B_UiUFMzzk8_0),.clk(gclk));
	jdff dff_B_kNH1NCLK2_0(.din(w_dff_B_UiUFMzzk8_0),.dout(w_dff_B_kNH1NCLK2_0),.clk(gclk));
	jdff dff_B_NRWs1TjP5_0(.din(w_dff_B_kNH1NCLK2_0),.dout(w_dff_B_NRWs1TjP5_0),.clk(gclk));
	jdff dff_B_LOKC2fWL6_0(.din(w_dff_B_NRWs1TjP5_0),.dout(w_dff_B_LOKC2fWL6_0),.clk(gclk));
	jdff dff_B_8XA5MRG59_0(.din(w_dff_B_LOKC2fWL6_0),.dout(w_dff_B_8XA5MRG59_0),.clk(gclk));
	jdff dff_B_5hP75AeK5_0(.din(w_dff_B_8XA5MRG59_0),.dout(w_dff_B_5hP75AeK5_0),.clk(gclk));
	jdff dff_B_CpvMz4mN2_0(.din(w_dff_B_5hP75AeK5_0),.dout(w_dff_B_CpvMz4mN2_0),.clk(gclk));
	jdff dff_B_8TvSFsgr7_0(.din(w_dff_B_CpvMz4mN2_0),.dout(w_dff_B_8TvSFsgr7_0),.clk(gclk));
	jdff dff_B_skCZuw8K6_0(.din(w_dff_B_8TvSFsgr7_0),.dout(w_dff_B_skCZuw8K6_0),.clk(gclk));
	jdff dff_B_yM04tRlt4_0(.din(w_dff_B_skCZuw8K6_0),.dout(w_dff_B_yM04tRlt4_0),.clk(gclk));
	jdff dff_B_R2yF4jim3_0(.din(w_dff_B_yM04tRlt4_0),.dout(w_dff_B_R2yF4jim3_0),.clk(gclk));
	jdff dff_B_6f3dN7QN8_0(.din(w_dff_B_R2yF4jim3_0),.dout(w_dff_B_6f3dN7QN8_0),.clk(gclk));
	jdff dff_B_gDrtT0l58_0(.din(w_dff_B_6f3dN7QN8_0),.dout(w_dff_B_gDrtT0l58_0),.clk(gclk));
	jdff dff_B_3MMhsFCd0_0(.din(w_dff_B_gDrtT0l58_0),.dout(w_dff_B_3MMhsFCd0_0),.clk(gclk));
	jdff dff_B_kQ1dnboA2_0(.din(w_dff_B_3MMhsFCd0_0),.dout(w_dff_B_kQ1dnboA2_0),.clk(gclk));
	jdff dff_B_urpsbfi53_0(.din(w_dff_B_kQ1dnboA2_0),.dout(w_dff_B_urpsbfi53_0),.clk(gclk));
	jdff dff_B_MVOLU3ws7_0(.din(w_dff_B_urpsbfi53_0),.dout(w_dff_B_MVOLU3ws7_0),.clk(gclk));
	jdff dff_B_mvmwfVA57_0(.din(w_dff_B_MVOLU3ws7_0),.dout(w_dff_B_mvmwfVA57_0),.clk(gclk));
	jdff dff_B_oDDBxuIg1_0(.din(w_dff_B_mvmwfVA57_0),.dout(w_dff_B_oDDBxuIg1_0),.clk(gclk));
	jdff dff_B_fdSxHe9t4_0(.din(w_dff_B_oDDBxuIg1_0),.dout(w_dff_B_fdSxHe9t4_0),.clk(gclk));
	jdff dff_B_GFar60K43_0(.din(w_dff_B_fdSxHe9t4_0),.dout(w_dff_B_GFar60K43_0),.clk(gclk));
	jdff dff_B_e4YMGjjT1_0(.din(w_dff_B_GFar60K43_0),.dout(w_dff_B_e4YMGjjT1_0),.clk(gclk));
	jdff dff_B_WpG0zDRd4_0(.din(w_dff_B_e4YMGjjT1_0),.dout(w_dff_B_WpG0zDRd4_0),.clk(gclk));
	jdff dff_B_UtCXg2np6_0(.din(w_dff_B_WpG0zDRd4_0),.dout(w_dff_B_UtCXg2np6_0),.clk(gclk));
	jdff dff_B_D3hAIm7G6_0(.din(w_dff_B_UtCXg2np6_0),.dout(w_dff_B_D3hAIm7G6_0),.clk(gclk));
	jdff dff_B_L9ET4TqU5_0(.din(w_dff_B_D3hAIm7G6_0),.dout(w_dff_B_L9ET4TqU5_0),.clk(gclk));
	jdff dff_B_LTiPZO7K5_0(.din(w_dff_B_L9ET4TqU5_0),.dout(w_dff_B_LTiPZO7K5_0),.clk(gclk));
	jdff dff_B_LJ1iqzgF4_0(.din(w_dff_B_LTiPZO7K5_0),.dout(w_dff_B_LJ1iqzgF4_0),.clk(gclk));
	jdff dff_B_yvo7MTYZ8_0(.din(w_dff_B_LJ1iqzgF4_0),.dout(w_dff_B_yvo7MTYZ8_0),.clk(gclk));
	jdff dff_B_UqTuvFWY4_0(.din(w_dff_B_yvo7MTYZ8_0),.dout(w_dff_B_UqTuvFWY4_0),.clk(gclk));
	jdff dff_B_vUGz1A9w7_0(.din(w_dff_B_UqTuvFWY4_0),.dout(w_dff_B_vUGz1A9w7_0),.clk(gclk));
	jdff dff_B_hmjJ8dgr7_0(.din(w_dff_B_vUGz1A9w7_0),.dout(w_dff_B_hmjJ8dgr7_0),.clk(gclk));
	jdff dff_B_RrUiokRv8_0(.din(w_dff_B_hmjJ8dgr7_0),.dout(w_dff_B_RrUiokRv8_0),.clk(gclk));
	jdff dff_B_jnL9yvYN9_0(.din(w_dff_B_RrUiokRv8_0),.dout(w_dff_B_jnL9yvYN9_0),.clk(gclk));
	jdff dff_B_Ev7GUK5u2_0(.din(w_dff_B_jnL9yvYN9_0),.dout(w_dff_B_Ev7GUK5u2_0),.clk(gclk));
	jdff dff_B_3tiwEpoL1_0(.din(w_dff_B_Ev7GUK5u2_0),.dout(w_dff_B_3tiwEpoL1_0),.clk(gclk));
	jdff dff_B_VmvndDKD0_0(.din(w_dff_B_3tiwEpoL1_0),.dout(w_dff_B_VmvndDKD0_0),.clk(gclk));
	jdff dff_B_WqPYqotT9_0(.din(w_dff_B_VmvndDKD0_0),.dout(w_dff_B_WqPYqotT9_0),.clk(gclk));
	jdff dff_B_meG3HzrP3_0(.din(w_dff_B_WqPYqotT9_0),.dout(w_dff_B_meG3HzrP3_0),.clk(gclk));
	jdff dff_B_GvEgjppo1_0(.din(w_dff_B_meG3HzrP3_0),.dout(w_dff_B_GvEgjppo1_0),.clk(gclk));
	jdff dff_B_24eN53Uy1_0(.din(w_dff_B_GvEgjppo1_0),.dout(w_dff_B_24eN53Uy1_0),.clk(gclk));
	jdff dff_B_x8EtnUJm3_0(.din(w_dff_B_24eN53Uy1_0),.dout(w_dff_B_x8EtnUJm3_0),.clk(gclk));
	jdff dff_B_RBaqlklD2_0(.din(w_dff_B_x8EtnUJm3_0),.dout(w_dff_B_RBaqlklD2_0),.clk(gclk));
	jdff dff_B_qIOzllUj9_0(.din(w_dff_B_RBaqlklD2_0),.dout(w_dff_B_qIOzllUj9_0),.clk(gclk));
	jdff dff_B_rF9TcJz53_0(.din(w_dff_B_qIOzllUj9_0),.dout(w_dff_B_rF9TcJz53_0),.clk(gclk));
	jdff dff_B_R4OJcZS96_0(.din(w_dff_B_rF9TcJz53_0),.dout(w_dff_B_R4OJcZS96_0),.clk(gclk));
	jdff dff_B_mWedHaVg3_0(.din(w_dff_B_R4OJcZS96_0),.dout(w_dff_B_mWedHaVg3_0),.clk(gclk));
	jdff dff_B_8cuSA7pD9_0(.din(w_dff_B_mWedHaVg3_0),.dout(w_dff_B_8cuSA7pD9_0),.clk(gclk));
	jdff dff_B_O4Kzfig71_0(.din(w_dff_B_8cuSA7pD9_0),.dout(w_dff_B_O4Kzfig71_0),.clk(gclk));
	jdff dff_B_UNVoVzip5_0(.din(w_dff_B_O4Kzfig71_0),.dout(w_dff_B_UNVoVzip5_0),.clk(gclk));
	jdff dff_B_CSnIVTiN1_0(.din(w_dff_B_UNVoVzip5_0),.dout(w_dff_B_CSnIVTiN1_0),.clk(gclk));
	jdff dff_B_ybU4RxjG7_0(.din(w_dff_B_CSnIVTiN1_0),.dout(w_dff_B_ybU4RxjG7_0),.clk(gclk));
	jdff dff_B_HZggoPB68_0(.din(w_dff_B_ybU4RxjG7_0),.dout(w_dff_B_HZggoPB68_0),.clk(gclk));
	jdff dff_B_YQeXZEzV6_0(.din(w_dff_B_HZggoPB68_0),.dout(w_dff_B_YQeXZEzV6_0),.clk(gclk));
	jdff dff_B_DFALM1Vp0_0(.din(w_dff_B_YQeXZEzV6_0),.dout(w_dff_B_DFALM1Vp0_0),.clk(gclk));
	jdff dff_B_WRu66ThJ8_0(.din(w_dff_B_DFALM1Vp0_0),.dout(w_dff_B_WRu66ThJ8_0),.clk(gclk));
	jdff dff_B_SeIvU6JH0_0(.din(w_dff_B_WRu66ThJ8_0),.dout(w_dff_B_SeIvU6JH0_0),.clk(gclk));
	jdff dff_B_0c5FSzV43_0(.din(w_dff_B_SeIvU6JH0_0),.dout(w_dff_B_0c5FSzV43_0),.clk(gclk));
	jdff dff_B_eft00hZo3_0(.din(w_dff_B_0c5FSzV43_0),.dout(w_dff_B_eft00hZo3_0),.clk(gclk));
	jdff dff_B_M3z591OZ9_0(.din(w_dff_B_eft00hZo3_0),.dout(w_dff_B_M3z591OZ9_0),.clk(gclk));
	jdff dff_B_DAlnCixT3_0(.din(n982),.dout(w_dff_B_DAlnCixT3_0),.clk(gclk));
	jdff dff_B_480fpUpr1_0(.din(w_dff_B_DAlnCixT3_0),.dout(w_dff_B_480fpUpr1_0),.clk(gclk));
	jdff dff_B_ygXPRUIH7_0(.din(w_dff_B_480fpUpr1_0),.dout(w_dff_B_ygXPRUIH7_0),.clk(gclk));
	jdff dff_B_H3ZEg4fS0_0(.din(w_dff_B_ygXPRUIH7_0),.dout(w_dff_B_H3ZEg4fS0_0),.clk(gclk));
	jdff dff_B_OqYZB5g93_0(.din(w_dff_B_H3ZEg4fS0_0),.dout(w_dff_B_OqYZB5g93_0),.clk(gclk));
	jdff dff_B_LGS1kK4r4_0(.din(w_dff_B_OqYZB5g93_0),.dout(w_dff_B_LGS1kK4r4_0),.clk(gclk));
	jdff dff_B_PihdAonI9_0(.din(w_dff_B_LGS1kK4r4_0),.dout(w_dff_B_PihdAonI9_0),.clk(gclk));
	jdff dff_B_q4GgwZBd6_0(.din(w_dff_B_PihdAonI9_0),.dout(w_dff_B_q4GgwZBd6_0),.clk(gclk));
	jdff dff_B_nkFkux7L2_0(.din(w_dff_B_q4GgwZBd6_0),.dout(w_dff_B_nkFkux7L2_0),.clk(gclk));
	jdff dff_B_lrEKLnkW3_0(.din(w_dff_B_nkFkux7L2_0),.dout(w_dff_B_lrEKLnkW3_0),.clk(gclk));
	jdff dff_B_gNWOrdoQ1_0(.din(w_dff_B_lrEKLnkW3_0),.dout(w_dff_B_gNWOrdoQ1_0),.clk(gclk));
	jdff dff_B_Xv1sEiPb6_0(.din(w_dff_B_gNWOrdoQ1_0),.dout(w_dff_B_Xv1sEiPb6_0),.clk(gclk));
	jdff dff_B_WCh4pQGB0_0(.din(w_dff_B_Xv1sEiPb6_0),.dout(w_dff_B_WCh4pQGB0_0),.clk(gclk));
	jdff dff_B_Ujz2OuiD1_0(.din(w_dff_B_WCh4pQGB0_0),.dout(w_dff_B_Ujz2OuiD1_0),.clk(gclk));
	jdff dff_B_Hs7IZQoM5_0(.din(w_dff_B_Ujz2OuiD1_0),.dout(w_dff_B_Hs7IZQoM5_0),.clk(gclk));
	jdff dff_B_Dm54EjHG2_0(.din(w_dff_B_Hs7IZQoM5_0),.dout(w_dff_B_Dm54EjHG2_0),.clk(gclk));
	jdff dff_B_87zPumQs9_0(.din(w_dff_B_Dm54EjHG2_0),.dout(w_dff_B_87zPumQs9_0),.clk(gclk));
	jdff dff_B_xfpY7DEM9_0(.din(w_dff_B_87zPumQs9_0),.dout(w_dff_B_xfpY7DEM9_0),.clk(gclk));
	jdff dff_B_GaJW3tMO1_0(.din(w_dff_B_xfpY7DEM9_0),.dout(w_dff_B_GaJW3tMO1_0),.clk(gclk));
	jdff dff_B_xcJtpljq5_0(.din(w_dff_B_GaJW3tMO1_0),.dout(w_dff_B_xcJtpljq5_0),.clk(gclk));
	jdff dff_B_uOt7OzVK6_0(.din(w_dff_B_xcJtpljq5_0),.dout(w_dff_B_uOt7OzVK6_0),.clk(gclk));
	jdff dff_B_7qeVJBD69_0(.din(w_dff_B_uOt7OzVK6_0),.dout(w_dff_B_7qeVJBD69_0),.clk(gclk));
	jdff dff_B_yyuyMGT65_0(.din(w_dff_B_7qeVJBD69_0),.dout(w_dff_B_yyuyMGT65_0),.clk(gclk));
	jdff dff_B_zLZT0Tce6_0(.din(w_dff_B_yyuyMGT65_0),.dout(w_dff_B_zLZT0Tce6_0),.clk(gclk));
	jdff dff_B_dS418c9I0_0(.din(w_dff_B_zLZT0Tce6_0),.dout(w_dff_B_dS418c9I0_0),.clk(gclk));
	jdff dff_B_VSsCDWao5_0(.din(w_dff_B_dS418c9I0_0),.dout(w_dff_B_VSsCDWao5_0),.clk(gclk));
	jdff dff_B_RUBwzeCd5_0(.din(w_dff_B_VSsCDWao5_0),.dout(w_dff_B_RUBwzeCd5_0),.clk(gclk));
	jdff dff_B_l0PYgtk60_0(.din(w_dff_B_RUBwzeCd5_0),.dout(w_dff_B_l0PYgtk60_0),.clk(gclk));
	jdff dff_B_5ELIJgwc3_0(.din(w_dff_B_l0PYgtk60_0),.dout(w_dff_B_5ELIJgwc3_0),.clk(gclk));
	jdff dff_B_Uz8gbmkX0_0(.din(w_dff_B_5ELIJgwc3_0),.dout(w_dff_B_Uz8gbmkX0_0),.clk(gclk));
	jdff dff_B_brAe0uFP4_0(.din(w_dff_B_Uz8gbmkX0_0),.dout(w_dff_B_brAe0uFP4_0),.clk(gclk));
	jdff dff_B_OVIPcE9O7_0(.din(w_dff_B_brAe0uFP4_0),.dout(w_dff_B_OVIPcE9O7_0),.clk(gclk));
	jdff dff_B_PupL3Jnj0_0(.din(w_dff_B_OVIPcE9O7_0),.dout(w_dff_B_PupL3Jnj0_0),.clk(gclk));
	jdff dff_B_Vx2dRgeS4_0(.din(w_dff_B_PupL3Jnj0_0),.dout(w_dff_B_Vx2dRgeS4_0),.clk(gclk));
	jdff dff_B_RXjy7JkA5_0(.din(w_dff_B_Vx2dRgeS4_0),.dout(w_dff_B_RXjy7JkA5_0),.clk(gclk));
	jdff dff_B_7OIIjJiv9_0(.din(w_dff_B_RXjy7JkA5_0),.dout(w_dff_B_7OIIjJiv9_0),.clk(gclk));
	jdff dff_B_tyhbdQX67_0(.din(w_dff_B_7OIIjJiv9_0),.dout(w_dff_B_tyhbdQX67_0),.clk(gclk));
	jdff dff_B_sHGVczSf8_0(.din(w_dff_B_tyhbdQX67_0),.dout(w_dff_B_sHGVczSf8_0),.clk(gclk));
	jdff dff_B_vjNYtJUJ1_0(.din(w_dff_B_sHGVczSf8_0),.dout(w_dff_B_vjNYtJUJ1_0),.clk(gclk));
	jdff dff_B_jNUyLwVg0_0(.din(w_dff_B_vjNYtJUJ1_0),.dout(w_dff_B_jNUyLwVg0_0),.clk(gclk));
	jdff dff_B_0hXimAm42_0(.din(w_dff_B_jNUyLwVg0_0),.dout(w_dff_B_0hXimAm42_0),.clk(gclk));
	jdff dff_B_g9lvzgj05_0(.din(w_dff_B_0hXimAm42_0),.dout(w_dff_B_g9lvzgj05_0),.clk(gclk));
	jdff dff_B_nSFZB8ys0_0(.din(w_dff_B_g9lvzgj05_0),.dout(w_dff_B_nSFZB8ys0_0),.clk(gclk));
	jdff dff_B_UNfF6J3U9_0(.din(w_dff_B_nSFZB8ys0_0),.dout(w_dff_B_UNfF6J3U9_0),.clk(gclk));
	jdff dff_B_RwnIKpvb8_0(.din(w_dff_B_UNfF6J3U9_0),.dout(w_dff_B_RwnIKpvb8_0),.clk(gclk));
	jdff dff_B_7RYfViia6_0(.din(w_dff_B_RwnIKpvb8_0),.dout(w_dff_B_7RYfViia6_0),.clk(gclk));
	jdff dff_B_guqjXXO03_0(.din(w_dff_B_7RYfViia6_0),.dout(w_dff_B_guqjXXO03_0),.clk(gclk));
	jdff dff_B_wxxFjGE56_0(.din(w_dff_B_guqjXXO03_0),.dout(w_dff_B_wxxFjGE56_0),.clk(gclk));
	jdff dff_B_GPikOGZW1_0(.din(w_dff_B_wxxFjGE56_0),.dout(w_dff_B_GPikOGZW1_0),.clk(gclk));
	jdff dff_B_VdTOUKKa2_0(.din(w_dff_B_GPikOGZW1_0),.dout(w_dff_B_VdTOUKKa2_0),.clk(gclk));
	jdff dff_B_m50nFDnK3_0(.din(w_dff_B_VdTOUKKa2_0),.dout(w_dff_B_m50nFDnK3_0),.clk(gclk));
	jdff dff_B_oTXl1Gi04_0(.din(w_dff_B_m50nFDnK3_0),.dout(w_dff_B_oTXl1Gi04_0),.clk(gclk));
	jdff dff_B_GNkyk62V2_0(.din(w_dff_B_oTXl1Gi04_0),.dout(w_dff_B_GNkyk62V2_0),.clk(gclk));
	jdff dff_B_Nhts54gS1_0(.din(w_dff_B_GNkyk62V2_0),.dout(w_dff_B_Nhts54gS1_0),.clk(gclk));
	jdff dff_B_orZoKxgX9_0(.din(w_dff_B_Nhts54gS1_0),.dout(w_dff_B_orZoKxgX9_0),.clk(gclk));
	jdff dff_B_eYmwcwLz3_0(.din(w_dff_B_orZoKxgX9_0),.dout(w_dff_B_eYmwcwLz3_0),.clk(gclk));
	jdff dff_B_vxh4chKb1_0(.din(w_dff_B_eYmwcwLz3_0),.dout(w_dff_B_vxh4chKb1_0),.clk(gclk));
	jdff dff_B_O5XuocJf1_0(.din(w_dff_B_vxh4chKb1_0),.dout(w_dff_B_O5XuocJf1_0),.clk(gclk));
	jdff dff_B_qh0VNzGu2_0(.din(w_dff_B_O5XuocJf1_0),.dout(w_dff_B_qh0VNzGu2_0),.clk(gclk));
	jdff dff_B_YlgCbFom8_0(.din(w_dff_B_qh0VNzGu2_0),.dout(w_dff_B_YlgCbFom8_0),.clk(gclk));
	jdff dff_B_0JpBfqp46_0(.din(w_dff_B_YlgCbFom8_0),.dout(w_dff_B_0JpBfqp46_0),.clk(gclk));
	jdff dff_B_JyshFPPs6_0(.din(w_dff_B_0JpBfqp46_0),.dout(w_dff_B_JyshFPPs6_0),.clk(gclk));
	jdff dff_B_PPZZ7XJq1_0(.din(w_dff_B_JyshFPPs6_0),.dout(w_dff_B_PPZZ7XJq1_0),.clk(gclk));
	jdff dff_B_SbNY8Z5z6_0(.din(w_dff_B_PPZZ7XJq1_0),.dout(w_dff_B_SbNY8Z5z6_0),.clk(gclk));
	jdff dff_B_XuYarmnf2_0(.din(w_dff_B_SbNY8Z5z6_0),.dout(w_dff_B_XuYarmnf2_0),.clk(gclk));
	jdff dff_B_SgfYSBrd1_0(.din(w_dff_B_XuYarmnf2_0),.dout(w_dff_B_SgfYSBrd1_0),.clk(gclk));
	jdff dff_B_jhOqBV6g7_0(.din(w_dff_B_SgfYSBrd1_0),.dout(w_dff_B_jhOqBV6g7_0),.clk(gclk));
	jdff dff_B_l5z5e8ni8_0(.din(w_dff_B_jhOqBV6g7_0),.dout(w_dff_B_l5z5e8ni8_0),.clk(gclk));
	jdff dff_B_mUrmYZRx9_0(.din(w_dff_B_l5z5e8ni8_0),.dout(w_dff_B_mUrmYZRx9_0),.clk(gclk));
	jdff dff_B_IJW5cSVS6_0(.din(w_dff_B_mUrmYZRx9_0),.dout(w_dff_B_IJW5cSVS6_0),.clk(gclk));
	jdff dff_B_aTXPPdsk3_0(.din(w_dff_B_IJW5cSVS6_0),.dout(w_dff_B_aTXPPdsk3_0),.clk(gclk));
	jdff dff_B_OwRqrd5q0_0(.din(w_dff_B_aTXPPdsk3_0),.dout(w_dff_B_OwRqrd5q0_0),.clk(gclk));
	jdff dff_B_MXU39VTA7_0(.din(w_dff_B_OwRqrd5q0_0),.dout(w_dff_B_MXU39VTA7_0),.clk(gclk));
	jdff dff_B_zro1Avn13_0(.din(w_dff_B_MXU39VTA7_0),.dout(w_dff_B_zro1Avn13_0),.clk(gclk));
	jdff dff_B_fJl1mHSm4_0(.din(w_dff_B_zro1Avn13_0),.dout(w_dff_B_fJl1mHSm4_0),.clk(gclk));
	jdff dff_B_AxD95VGg4_0(.din(w_dff_B_fJl1mHSm4_0),.dout(w_dff_B_AxD95VGg4_0),.clk(gclk));
	jdff dff_B_vyxqTUgj3_0(.din(w_dff_B_AxD95VGg4_0),.dout(w_dff_B_vyxqTUgj3_0),.clk(gclk));
	jdff dff_B_pofWpHeK6_0(.din(w_dff_B_vyxqTUgj3_0),.dout(w_dff_B_pofWpHeK6_0),.clk(gclk));
	jdff dff_B_X7PrYFQ60_0(.din(w_dff_B_pofWpHeK6_0),.dout(w_dff_B_X7PrYFQ60_0),.clk(gclk));
	jdff dff_B_DjC3kDmD0_0(.din(w_dff_B_X7PrYFQ60_0),.dout(w_dff_B_DjC3kDmD0_0),.clk(gclk));
	jdff dff_B_oXz1HTAS4_0(.din(w_dff_B_DjC3kDmD0_0),.dout(w_dff_B_oXz1HTAS4_0),.clk(gclk));
	jdff dff_B_wMNURBNE3_0(.din(w_dff_B_oXz1HTAS4_0),.dout(w_dff_B_wMNURBNE3_0),.clk(gclk));
	jdff dff_B_6JZWmO0a8_0(.din(w_dff_B_wMNURBNE3_0),.dout(w_dff_B_6JZWmO0a8_0),.clk(gclk));
	jdff dff_B_2ZXq0dxu8_0(.din(w_dff_B_6JZWmO0a8_0),.dout(w_dff_B_2ZXq0dxu8_0),.clk(gclk));
	jdff dff_B_MxNAwhCS2_0(.din(w_dff_B_2ZXq0dxu8_0),.dout(w_dff_B_MxNAwhCS2_0),.clk(gclk));
	jdff dff_B_bCxsUiei6_0(.din(w_dff_B_MxNAwhCS2_0),.dout(w_dff_B_bCxsUiei6_0),.clk(gclk));
	jdff dff_B_9zTGPg8K3_0(.din(w_dff_B_bCxsUiei6_0),.dout(w_dff_B_9zTGPg8K3_0),.clk(gclk));
	jdff dff_B_iARsXMcr3_0(.din(w_dff_B_9zTGPg8K3_0),.dout(w_dff_B_iARsXMcr3_0),.clk(gclk));
	jdff dff_B_yT7kWIM38_0(.din(w_dff_B_iARsXMcr3_0),.dout(w_dff_B_yT7kWIM38_0),.clk(gclk));
	jdff dff_B_CRWWdflb4_0(.din(w_dff_B_yT7kWIM38_0),.dout(w_dff_B_CRWWdflb4_0),.clk(gclk));
	jdff dff_B_hZm8Mf0L9_0(.din(w_dff_B_CRWWdflb4_0),.dout(w_dff_B_hZm8Mf0L9_0),.clk(gclk));
	jdff dff_B_vz8V1pPd1_0(.din(w_dff_B_hZm8Mf0L9_0),.dout(w_dff_B_vz8V1pPd1_0),.clk(gclk));
	jdff dff_B_GL4Grb4P3_0(.din(w_dff_B_vz8V1pPd1_0),.dout(w_dff_B_GL4Grb4P3_0),.clk(gclk));
	jdff dff_B_OBczsvOg4_0(.din(w_dff_B_GL4Grb4P3_0),.dout(w_dff_B_OBczsvOg4_0),.clk(gclk));
	jdff dff_B_5KTdh6Ph9_0(.din(w_dff_B_OBczsvOg4_0),.dout(w_dff_B_5KTdh6Ph9_0),.clk(gclk));
	jdff dff_B_oeFDRw2b9_0(.din(w_dff_B_5KTdh6Ph9_0),.dout(w_dff_B_oeFDRw2b9_0),.clk(gclk));
	jdff dff_B_7MhKQS0Y9_0(.din(w_dff_B_oeFDRw2b9_0),.dout(w_dff_B_7MhKQS0Y9_0),.clk(gclk));
	jdff dff_B_7Or7W8OI3_0(.din(w_dff_B_7MhKQS0Y9_0),.dout(w_dff_B_7Or7W8OI3_0),.clk(gclk));
	jdff dff_B_hGgjVT1m4_0(.din(w_dff_B_7Or7W8OI3_0),.dout(w_dff_B_hGgjVT1m4_0),.clk(gclk));
	jdff dff_B_cxQHbRrb4_0(.din(n988),.dout(w_dff_B_cxQHbRrb4_0),.clk(gclk));
	jdff dff_B_xdSkvs3I5_0(.din(w_dff_B_cxQHbRrb4_0),.dout(w_dff_B_xdSkvs3I5_0),.clk(gclk));
	jdff dff_B_rTwRzNAk7_0(.din(w_dff_B_xdSkvs3I5_0),.dout(w_dff_B_rTwRzNAk7_0),.clk(gclk));
	jdff dff_B_lf3cti9i9_0(.din(w_dff_B_rTwRzNAk7_0),.dout(w_dff_B_lf3cti9i9_0),.clk(gclk));
	jdff dff_B_UfsG2AX90_0(.din(w_dff_B_lf3cti9i9_0),.dout(w_dff_B_UfsG2AX90_0),.clk(gclk));
	jdff dff_B_U6YoEVXG6_0(.din(w_dff_B_UfsG2AX90_0),.dout(w_dff_B_U6YoEVXG6_0),.clk(gclk));
	jdff dff_B_W24lS6cO7_0(.din(w_dff_B_U6YoEVXG6_0),.dout(w_dff_B_W24lS6cO7_0),.clk(gclk));
	jdff dff_B_yCVdShtp5_0(.din(w_dff_B_W24lS6cO7_0),.dout(w_dff_B_yCVdShtp5_0),.clk(gclk));
	jdff dff_B_a3YReHKm5_0(.din(w_dff_B_yCVdShtp5_0),.dout(w_dff_B_a3YReHKm5_0),.clk(gclk));
	jdff dff_B_H07vlX996_0(.din(w_dff_B_a3YReHKm5_0),.dout(w_dff_B_H07vlX996_0),.clk(gclk));
	jdff dff_B_p0WI3M5P7_0(.din(w_dff_B_H07vlX996_0),.dout(w_dff_B_p0WI3M5P7_0),.clk(gclk));
	jdff dff_B_D8WtqPFi1_0(.din(w_dff_B_p0WI3M5P7_0),.dout(w_dff_B_D8WtqPFi1_0),.clk(gclk));
	jdff dff_B_XveV5cCh8_0(.din(w_dff_B_D8WtqPFi1_0),.dout(w_dff_B_XveV5cCh8_0),.clk(gclk));
	jdff dff_B_tHAyiOmX3_0(.din(w_dff_B_XveV5cCh8_0),.dout(w_dff_B_tHAyiOmX3_0),.clk(gclk));
	jdff dff_B_lm6QGgng2_0(.din(w_dff_B_tHAyiOmX3_0),.dout(w_dff_B_lm6QGgng2_0),.clk(gclk));
	jdff dff_B_rJ30bGHP0_0(.din(w_dff_B_lm6QGgng2_0),.dout(w_dff_B_rJ30bGHP0_0),.clk(gclk));
	jdff dff_B_93ISU1Se1_0(.din(w_dff_B_rJ30bGHP0_0),.dout(w_dff_B_93ISU1Se1_0),.clk(gclk));
	jdff dff_B_QNtnG1XT5_0(.din(w_dff_B_93ISU1Se1_0),.dout(w_dff_B_QNtnG1XT5_0),.clk(gclk));
	jdff dff_B_mbPHK5WD0_0(.din(w_dff_B_QNtnG1XT5_0),.dout(w_dff_B_mbPHK5WD0_0),.clk(gclk));
	jdff dff_B_U9DxhiUg5_0(.din(w_dff_B_mbPHK5WD0_0),.dout(w_dff_B_U9DxhiUg5_0),.clk(gclk));
	jdff dff_B_29c6tTxp3_0(.din(w_dff_B_U9DxhiUg5_0),.dout(w_dff_B_29c6tTxp3_0),.clk(gclk));
	jdff dff_B_bGRpgUhq1_0(.din(w_dff_B_29c6tTxp3_0),.dout(w_dff_B_bGRpgUhq1_0),.clk(gclk));
	jdff dff_B_vmCGCL2L4_0(.din(w_dff_B_bGRpgUhq1_0),.dout(w_dff_B_vmCGCL2L4_0),.clk(gclk));
	jdff dff_B_6uNI6KZv2_0(.din(w_dff_B_vmCGCL2L4_0),.dout(w_dff_B_6uNI6KZv2_0),.clk(gclk));
	jdff dff_B_9qI6ZFZn9_0(.din(w_dff_B_6uNI6KZv2_0),.dout(w_dff_B_9qI6ZFZn9_0),.clk(gclk));
	jdff dff_B_9o382cXc3_0(.din(w_dff_B_9qI6ZFZn9_0),.dout(w_dff_B_9o382cXc3_0),.clk(gclk));
	jdff dff_B_h3AaYqih9_0(.din(w_dff_B_9o382cXc3_0),.dout(w_dff_B_h3AaYqih9_0),.clk(gclk));
	jdff dff_B_YaCtgqK82_0(.din(w_dff_B_h3AaYqih9_0),.dout(w_dff_B_YaCtgqK82_0),.clk(gclk));
	jdff dff_B_zanO9U3n3_0(.din(w_dff_B_YaCtgqK82_0),.dout(w_dff_B_zanO9U3n3_0),.clk(gclk));
	jdff dff_B_jBiVlFCR9_0(.din(w_dff_B_zanO9U3n3_0),.dout(w_dff_B_jBiVlFCR9_0),.clk(gclk));
	jdff dff_B_kQXg7P1b7_0(.din(w_dff_B_jBiVlFCR9_0),.dout(w_dff_B_kQXg7P1b7_0),.clk(gclk));
	jdff dff_B_s5l04Gn46_0(.din(w_dff_B_kQXg7P1b7_0),.dout(w_dff_B_s5l04Gn46_0),.clk(gclk));
	jdff dff_B_YZl2ArNk6_0(.din(w_dff_B_s5l04Gn46_0),.dout(w_dff_B_YZl2ArNk6_0),.clk(gclk));
	jdff dff_B_dPN2vdxK9_0(.din(w_dff_B_YZl2ArNk6_0),.dout(w_dff_B_dPN2vdxK9_0),.clk(gclk));
	jdff dff_B_GOisHFjS3_0(.din(w_dff_B_dPN2vdxK9_0),.dout(w_dff_B_GOisHFjS3_0),.clk(gclk));
	jdff dff_B_pg8VuWm85_0(.din(w_dff_B_GOisHFjS3_0),.dout(w_dff_B_pg8VuWm85_0),.clk(gclk));
	jdff dff_B_XFFpCov71_0(.din(w_dff_B_pg8VuWm85_0),.dout(w_dff_B_XFFpCov71_0),.clk(gclk));
	jdff dff_B_4DmOdg1F0_0(.din(w_dff_B_XFFpCov71_0),.dout(w_dff_B_4DmOdg1F0_0),.clk(gclk));
	jdff dff_B_SztyR6N21_0(.din(w_dff_B_4DmOdg1F0_0),.dout(w_dff_B_SztyR6N21_0),.clk(gclk));
	jdff dff_B_cI1t0jWd4_0(.din(w_dff_B_SztyR6N21_0),.dout(w_dff_B_cI1t0jWd4_0),.clk(gclk));
	jdff dff_B_TYj3X4Pm0_0(.din(w_dff_B_cI1t0jWd4_0),.dout(w_dff_B_TYj3X4Pm0_0),.clk(gclk));
	jdff dff_B_Ekk6QjLl5_0(.din(w_dff_B_TYj3X4Pm0_0),.dout(w_dff_B_Ekk6QjLl5_0),.clk(gclk));
	jdff dff_B_mUSciLFF7_0(.din(w_dff_B_Ekk6QjLl5_0),.dout(w_dff_B_mUSciLFF7_0),.clk(gclk));
	jdff dff_B_5TCqRFol3_0(.din(w_dff_B_mUSciLFF7_0),.dout(w_dff_B_5TCqRFol3_0),.clk(gclk));
	jdff dff_B_oQU9RbYs3_0(.din(w_dff_B_5TCqRFol3_0),.dout(w_dff_B_oQU9RbYs3_0),.clk(gclk));
	jdff dff_B_j7ga9LeB6_0(.din(w_dff_B_oQU9RbYs3_0),.dout(w_dff_B_j7ga9LeB6_0),.clk(gclk));
	jdff dff_B_ltd9MiKv9_0(.din(w_dff_B_j7ga9LeB6_0),.dout(w_dff_B_ltd9MiKv9_0),.clk(gclk));
	jdff dff_B_bb7oX1hP5_0(.din(w_dff_B_ltd9MiKv9_0),.dout(w_dff_B_bb7oX1hP5_0),.clk(gclk));
	jdff dff_B_GzIPLYZ21_0(.din(w_dff_B_bb7oX1hP5_0),.dout(w_dff_B_GzIPLYZ21_0),.clk(gclk));
	jdff dff_B_Zl28QESE7_0(.din(w_dff_B_GzIPLYZ21_0),.dout(w_dff_B_Zl28QESE7_0),.clk(gclk));
	jdff dff_B_uoX7Oait0_0(.din(w_dff_B_Zl28QESE7_0),.dout(w_dff_B_uoX7Oait0_0),.clk(gclk));
	jdff dff_B_UKPKORPl6_0(.din(w_dff_B_uoX7Oait0_0),.dout(w_dff_B_UKPKORPl6_0),.clk(gclk));
	jdff dff_B_YX7GABMR7_0(.din(w_dff_B_UKPKORPl6_0),.dout(w_dff_B_YX7GABMR7_0),.clk(gclk));
	jdff dff_B_U2ZnsQuv4_0(.din(w_dff_B_YX7GABMR7_0),.dout(w_dff_B_U2ZnsQuv4_0),.clk(gclk));
	jdff dff_B_JT82WYwF6_0(.din(w_dff_B_U2ZnsQuv4_0),.dout(w_dff_B_JT82WYwF6_0),.clk(gclk));
	jdff dff_B_apnq8xML3_0(.din(w_dff_B_JT82WYwF6_0),.dout(w_dff_B_apnq8xML3_0),.clk(gclk));
	jdff dff_B_89uhpWyp0_0(.din(w_dff_B_apnq8xML3_0),.dout(w_dff_B_89uhpWyp0_0),.clk(gclk));
	jdff dff_B_GIlVFjpc8_0(.din(w_dff_B_89uhpWyp0_0),.dout(w_dff_B_GIlVFjpc8_0),.clk(gclk));
	jdff dff_B_muW3arSx4_0(.din(w_dff_B_GIlVFjpc8_0),.dout(w_dff_B_muW3arSx4_0),.clk(gclk));
	jdff dff_B_rlyya7Q45_0(.din(w_dff_B_muW3arSx4_0),.dout(w_dff_B_rlyya7Q45_0),.clk(gclk));
	jdff dff_B_QZm4Rezf6_0(.din(w_dff_B_rlyya7Q45_0),.dout(w_dff_B_QZm4Rezf6_0),.clk(gclk));
	jdff dff_B_1c7Ow9ex5_0(.din(w_dff_B_QZm4Rezf6_0),.dout(w_dff_B_1c7Ow9ex5_0),.clk(gclk));
	jdff dff_B_1jNH5cUL4_0(.din(w_dff_B_1c7Ow9ex5_0),.dout(w_dff_B_1jNH5cUL4_0),.clk(gclk));
	jdff dff_B_qbkdhUaH2_0(.din(w_dff_B_1jNH5cUL4_0),.dout(w_dff_B_qbkdhUaH2_0),.clk(gclk));
	jdff dff_B_VcCJnFgE2_0(.din(w_dff_B_qbkdhUaH2_0),.dout(w_dff_B_VcCJnFgE2_0),.clk(gclk));
	jdff dff_B_9tz9GHYq1_0(.din(w_dff_B_VcCJnFgE2_0),.dout(w_dff_B_9tz9GHYq1_0),.clk(gclk));
	jdff dff_B_ng2nA4ap7_0(.din(w_dff_B_9tz9GHYq1_0),.dout(w_dff_B_ng2nA4ap7_0),.clk(gclk));
	jdff dff_B_Q6yt5r8u4_0(.din(w_dff_B_ng2nA4ap7_0),.dout(w_dff_B_Q6yt5r8u4_0),.clk(gclk));
	jdff dff_B_OGlxJj7O4_0(.din(w_dff_B_Q6yt5r8u4_0),.dout(w_dff_B_OGlxJj7O4_0),.clk(gclk));
	jdff dff_B_xkBpH88v2_0(.din(w_dff_B_OGlxJj7O4_0),.dout(w_dff_B_xkBpH88v2_0),.clk(gclk));
	jdff dff_B_nyNqJLOO5_0(.din(w_dff_B_xkBpH88v2_0),.dout(w_dff_B_nyNqJLOO5_0),.clk(gclk));
	jdff dff_B_pj7yDpwE5_0(.din(w_dff_B_nyNqJLOO5_0),.dout(w_dff_B_pj7yDpwE5_0),.clk(gclk));
	jdff dff_B_Aq64c9ZN5_0(.din(w_dff_B_pj7yDpwE5_0),.dout(w_dff_B_Aq64c9ZN5_0),.clk(gclk));
	jdff dff_B_XwKTvYa33_0(.din(w_dff_B_Aq64c9ZN5_0),.dout(w_dff_B_XwKTvYa33_0),.clk(gclk));
	jdff dff_B_P8lAmxvD7_0(.din(w_dff_B_XwKTvYa33_0),.dout(w_dff_B_P8lAmxvD7_0),.clk(gclk));
	jdff dff_B_lmc9HCMD2_0(.din(w_dff_B_P8lAmxvD7_0),.dout(w_dff_B_lmc9HCMD2_0),.clk(gclk));
	jdff dff_B_eH62Bknl2_0(.din(w_dff_B_lmc9HCMD2_0),.dout(w_dff_B_eH62Bknl2_0),.clk(gclk));
	jdff dff_B_m9vDMMVt4_0(.din(w_dff_B_eH62Bknl2_0),.dout(w_dff_B_m9vDMMVt4_0),.clk(gclk));
	jdff dff_B_gfGgB88U4_0(.din(w_dff_B_m9vDMMVt4_0),.dout(w_dff_B_gfGgB88U4_0),.clk(gclk));
	jdff dff_B_F95Yo3fz7_0(.din(w_dff_B_gfGgB88U4_0),.dout(w_dff_B_F95Yo3fz7_0),.clk(gclk));
	jdff dff_B_C304g7ml1_0(.din(w_dff_B_F95Yo3fz7_0),.dout(w_dff_B_C304g7ml1_0),.clk(gclk));
	jdff dff_B_VNkkN1Qm1_0(.din(w_dff_B_C304g7ml1_0),.dout(w_dff_B_VNkkN1Qm1_0),.clk(gclk));
	jdff dff_B_3k8weLLt7_0(.din(w_dff_B_VNkkN1Qm1_0),.dout(w_dff_B_3k8weLLt7_0),.clk(gclk));
	jdff dff_B_AyeCyypE6_0(.din(w_dff_B_3k8weLLt7_0),.dout(w_dff_B_AyeCyypE6_0),.clk(gclk));
	jdff dff_B_KrjLWKeI8_0(.din(w_dff_B_AyeCyypE6_0),.dout(w_dff_B_KrjLWKeI8_0),.clk(gclk));
	jdff dff_B_MfQQ1Ux78_0(.din(w_dff_B_KrjLWKeI8_0),.dout(w_dff_B_MfQQ1Ux78_0),.clk(gclk));
	jdff dff_B_3xIjYwtq8_0(.din(w_dff_B_MfQQ1Ux78_0),.dout(w_dff_B_3xIjYwtq8_0),.clk(gclk));
	jdff dff_B_Pfm1yHMo5_0(.din(w_dff_B_3xIjYwtq8_0),.dout(w_dff_B_Pfm1yHMo5_0),.clk(gclk));
	jdff dff_B_o7rBlzRd7_0(.din(w_dff_B_Pfm1yHMo5_0),.dout(w_dff_B_o7rBlzRd7_0),.clk(gclk));
	jdff dff_B_aSXVF1Rs2_0(.din(w_dff_B_o7rBlzRd7_0),.dout(w_dff_B_aSXVF1Rs2_0),.clk(gclk));
	jdff dff_B_bp9mHlMY2_0(.din(w_dff_B_aSXVF1Rs2_0),.dout(w_dff_B_bp9mHlMY2_0),.clk(gclk));
	jdff dff_B_PFpFZXWe9_0(.din(w_dff_B_bp9mHlMY2_0),.dout(w_dff_B_PFpFZXWe9_0),.clk(gclk));
	jdff dff_B_djlnkOzk7_0(.din(w_dff_B_PFpFZXWe9_0),.dout(w_dff_B_djlnkOzk7_0),.clk(gclk));
	jdff dff_B_h0WDq8K44_0(.din(w_dff_B_djlnkOzk7_0),.dout(w_dff_B_h0WDq8K44_0),.clk(gclk));
	jdff dff_B_63gHmbso9_0(.din(w_dff_B_h0WDq8K44_0),.dout(w_dff_B_63gHmbso9_0),.clk(gclk));
	jdff dff_B_xtYKZpYA4_0(.din(w_dff_B_63gHmbso9_0),.dout(w_dff_B_xtYKZpYA4_0),.clk(gclk));
	jdff dff_B_I2OCK4JD0_0(.din(w_dff_B_xtYKZpYA4_0),.dout(w_dff_B_I2OCK4JD0_0),.clk(gclk));
	jdff dff_B_pvqwtDtB6_0(.din(w_dff_B_I2OCK4JD0_0),.dout(w_dff_B_pvqwtDtB6_0),.clk(gclk));
	jdff dff_B_7vugEMsJ2_0(.din(w_dff_B_pvqwtDtB6_0),.dout(w_dff_B_7vugEMsJ2_0),.clk(gclk));
	jdff dff_B_Rw2JWE0p7_0(.din(w_dff_B_7vugEMsJ2_0),.dout(w_dff_B_Rw2JWE0p7_0),.clk(gclk));
	jdff dff_B_YpXZJu6A1_0(.din(n994),.dout(w_dff_B_YpXZJu6A1_0),.clk(gclk));
	jdff dff_B_NUMclR8m9_0(.din(w_dff_B_YpXZJu6A1_0),.dout(w_dff_B_NUMclR8m9_0),.clk(gclk));
	jdff dff_B_Ohydm42G4_0(.din(w_dff_B_NUMclR8m9_0),.dout(w_dff_B_Ohydm42G4_0),.clk(gclk));
	jdff dff_B_lfNMoP7O0_0(.din(w_dff_B_Ohydm42G4_0),.dout(w_dff_B_lfNMoP7O0_0),.clk(gclk));
	jdff dff_B_dh43NSpn4_0(.din(w_dff_B_lfNMoP7O0_0),.dout(w_dff_B_dh43NSpn4_0),.clk(gclk));
	jdff dff_B_IAtPc13h2_0(.din(w_dff_B_dh43NSpn4_0),.dout(w_dff_B_IAtPc13h2_0),.clk(gclk));
	jdff dff_B_AX0gEQ749_0(.din(w_dff_B_IAtPc13h2_0),.dout(w_dff_B_AX0gEQ749_0),.clk(gclk));
	jdff dff_B_aGKJxMg95_0(.din(w_dff_B_AX0gEQ749_0),.dout(w_dff_B_aGKJxMg95_0),.clk(gclk));
	jdff dff_B_0DOMc9m97_0(.din(w_dff_B_aGKJxMg95_0),.dout(w_dff_B_0DOMc9m97_0),.clk(gclk));
	jdff dff_B_aNkRzRjd9_0(.din(w_dff_B_0DOMc9m97_0),.dout(w_dff_B_aNkRzRjd9_0),.clk(gclk));
	jdff dff_B_FSOHVuNe4_0(.din(w_dff_B_aNkRzRjd9_0),.dout(w_dff_B_FSOHVuNe4_0),.clk(gclk));
	jdff dff_B_2fga3iRe5_0(.din(w_dff_B_FSOHVuNe4_0),.dout(w_dff_B_2fga3iRe5_0),.clk(gclk));
	jdff dff_B_BVAOB23F3_0(.din(w_dff_B_2fga3iRe5_0),.dout(w_dff_B_BVAOB23F3_0),.clk(gclk));
	jdff dff_B_cQPiGk7P6_0(.din(w_dff_B_BVAOB23F3_0),.dout(w_dff_B_cQPiGk7P6_0),.clk(gclk));
	jdff dff_B_cSBO8h2r9_0(.din(w_dff_B_cQPiGk7P6_0),.dout(w_dff_B_cSBO8h2r9_0),.clk(gclk));
	jdff dff_B_4O5uDLRc8_0(.din(w_dff_B_cSBO8h2r9_0),.dout(w_dff_B_4O5uDLRc8_0),.clk(gclk));
	jdff dff_B_mRhuBEzX7_0(.din(w_dff_B_4O5uDLRc8_0),.dout(w_dff_B_mRhuBEzX7_0),.clk(gclk));
	jdff dff_B_trsMTfJV7_0(.din(w_dff_B_mRhuBEzX7_0),.dout(w_dff_B_trsMTfJV7_0),.clk(gclk));
	jdff dff_B_hs0bIqB05_0(.din(w_dff_B_trsMTfJV7_0),.dout(w_dff_B_hs0bIqB05_0),.clk(gclk));
	jdff dff_B_YuHPHLcZ5_0(.din(w_dff_B_hs0bIqB05_0),.dout(w_dff_B_YuHPHLcZ5_0),.clk(gclk));
	jdff dff_B_CKv0lEqe8_0(.din(w_dff_B_YuHPHLcZ5_0),.dout(w_dff_B_CKv0lEqe8_0),.clk(gclk));
	jdff dff_B_0pCnJL7O1_0(.din(w_dff_B_CKv0lEqe8_0),.dout(w_dff_B_0pCnJL7O1_0),.clk(gclk));
	jdff dff_B_69MVTQxo8_0(.din(w_dff_B_0pCnJL7O1_0),.dout(w_dff_B_69MVTQxo8_0),.clk(gclk));
	jdff dff_B_yX6tNH4N1_0(.din(w_dff_B_69MVTQxo8_0),.dout(w_dff_B_yX6tNH4N1_0),.clk(gclk));
	jdff dff_B_YHoNSSNz7_0(.din(w_dff_B_yX6tNH4N1_0),.dout(w_dff_B_YHoNSSNz7_0),.clk(gclk));
	jdff dff_B_OrKrD8ZZ4_0(.din(w_dff_B_YHoNSSNz7_0),.dout(w_dff_B_OrKrD8ZZ4_0),.clk(gclk));
	jdff dff_B_kEuOdEsw4_0(.din(w_dff_B_OrKrD8ZZ4_0),.dout(w_dff_B_kEuOdEsw4_0),.clk(gclk));
	jdff dff_B_CKTaj6S72_0(.din(w_dff_B_kEuOdEsw4_0),.dout(w_dff_B_CKTaj6S72_0),.clk(gclk));
	jdff dff_B_4mjVS48m6_0(.din(w_dff_B_CKTaj6S72_0),.dout(w_dff_B_4mjVS48m6_0),.clk(gclk));
	jdff dff_B_2HaBSoxF6_0(.din(w_dff_B_4mjVS48m6_0),.dout(w_dff_B_2HaBSoxF6_0),.clk(gclk));
	jdff dff_B_OJZiK74L5_0(.din(w_dff_B_2HaBSoxF6_0),.dout(w_dff_B_OJZiK74L5_0),.clk(gclk));
	jdff dff_B_iuslrgjc1_0(.din(w_dff_B_OJZiK74L5_0),.dout(w_dff_B_iuslrgjc1_0),.clk(gclk));
	jdff dff_B_R4X4vpoZ1_0(.din(w_dff_B_iuslrgjc1_0),.dout(w_dff_B_R4X4vpoZ1_0),.clk(gclk));
	jdff dff_B_6b6Ll4sr8_0(.din(w_dff_B_R4X4vpoZ1_0),.dout(w_dff_B_6b6Ll4sr8_0),.clk(gclk));
	jdff dff_B_0nen7ZoL0_0(.din(w_dff_B_6b6Ll4sr8_0),.dout(w_dff_B_0nen7ZoL0_0),.clk(gclk));
	jdff dff_B_o5fE4GQ61_0(.din(w_dff_B_0nen7ZoL0_0),.dout(w_dff_B_o5fE4GQ61_0),.clk(gclk));
	jdff dff_B_pdB5P6nR6_0(.din(w_dff_B_o5fE4GQ61_0),.dout(w_dff_B_pdB5P6nR6_0),.clk(gclk));
	jdff dff_B_yrAlxNKZ0_0(.din(w_dff_B_pdB5P6nR6_0),.dout(w_dff_B_yrAlxNKZ0_0),.clk(gclk));
	jdff dff_B_dO9dIBhX7_0(.din(w_dff_B_yrAlxNKZ0_0),.dout(w_dff_B_dO9dIBhX7_0),.clk(gclk));
	jdff dff_B_PkSPLW072_0(.din(w_dff_B_dO9dIBhX7_0),.dout(w_dff_B_PkSPLW072_0),.clk(gclk));
	jdff dff_B_xiWc8TLK1_0(.din(w_dff_B_PkSPLW072_0),.dout(w_dff_B_xiWc8TLK1_0),.clk(gclk));
	jdff dff_B_lWhkR4ix3_0(.din(w_dff_B_xiWc8TLK1_0),.dout(w_dff_B_lWhkR4ix3_0),.clk(gclk));
	jdff dff_B_BU5Wzufg0_0(.din(w_dff_B_lWhkR4ix3_0),.dout(w_dff_B_BU5Wzufg0_0),.clk(gclk));
	jdff dff_B_J9WR5ZO72_0(.din(w_dff_B_BU5Wzufg0_0),.dout(w_dff_B_J9WR5ZO72_0),.clk(gclk));
	jdff dff_B_UosIINje5_0(.din(w_dff_B_J9WR5ZO72_0),.dout(w_dff_B_UosIINje5_0),.clk(gclk));
	jdff dff_B_Ua7JFNbw0_0(.din(w_dff_B_UosIINje5_0),.dout(w_dff_B_Ua7JFNbw0_0),.clk(gclk));
	jdff dff_B_3oYeOmZE3_0(.din(w_dff_B_Ua7JFNbw0_0),.dout(w_dff_B_3oYeOmZE3_0),.clk(gclk));
	jdff dff_B_cu7jrV3J3_0(.din(w_dff_B_3oYeOmZE3_0),.dout(w_dff_B_cu7jrV3J3_0),.clk(gclk));
	jdff dff_B_kpU3coUu6_0(.din(w_dff_B_cu7jrV3J3_0),.dout(w_dff_B_kpU3coUu6_0),.clk(gclk));
	jdff dff_B_8L7DzqaR0_0(.din(w_dff_B_kpU3coUu6_0),.dout(w_dff_B_8L7DzqaR0_0),.clk(gclk));
	jdff dff_B_esNMC7tL1_0(.din(w_dff_B_8L7DzqaR0_0),.dout(w_dff_B_esNMC7tL1_0),.clk(gclk));
	jdff dff_B_yPwD44Iu3_0(.din(w_dff_B_esNMC7tL1_0),.dout(w_dff_B_yPwD44Iu3_0),.clk(gclk));
	jdff dff_B_APOZFSFv5_0(.din(w_dff_B_yPwD44Iu3_0),.dout(w_dff_B_APOZFSFv5_0),.clk(gclk));
	jdff dff_B_CWbYvsI17_0(.din(w_dff_B_APOZFSFv5_0),.dout(w_dff_B_CWbYvsI17_0),.clk(gclk));
	jdff dff_B_bdOlm3cp4_0(.din(w_dff_B_CWbYvsI17_0),.dout(w_dff_B_bdOlm3cp4_0),.clk(gclk));
	jdff dff_B_bNXFubr90_0(.din(w_dff_B_bdOlm3cp4_0),.dout(w_dff_B_bNXFubr90_0),.clk(gclk));
	jdff dff_B_EEk01UaF8_0(.din(w_dff_B_bNXFubr90_0),.dout(w_dff_B_EEk01UaF8_0),.clk(gclk));
	jdff dff_B_5EmVVvVd1_0(.din(w_dff_B_EEk01UaF8_0),.dout(w_dff_B_5EmVVvVd1_0),.clk(gclk));
	jdff dff_B_oDm5FM826_0(.din(w_dff_B_5EmVVvVd1_0),.dout(w_dff_B_oDm5FM826_0),.clk(gclk));
	jdff dff_B_sMpz7B927_0(.din(w_dff_B_oDm5FM826_0),.dout(w_dff_B_sMpz7B927_0),.clk(gclk));
	jdff dff_B_i9iZlJfX8_0(.din(w_dff_B_sMpz7B927_0),.dout(w_dff_B_i9iZlJfX8_0),.clk(gclk));
	jdff dff_B_NFjNaAnv6_0(.din(w_dff_B_i9iZlJfX8_0),.dout(w_dff_B_NFjNaAnv6_0),.clk(gclk));
	jdff dff_B_wRkKeCvy3_0(.din(w_dff_B_NFjNaAnv6_0),.dout(w_dff_B_wRkKeCvy3_0),.clk(gclk));
	jdff dff_B_5tUusbz36_0(.din(w_dff_B_wRkKeCvy3_0),.dout(w_dff_B_5tUusbz36_0),.clk(gclk));
	jdff dff_B_PISKIqu05_0(.din(w_dff_B_5tUusbz36_0),.dout(w_dff_B_PISKIqu05_0),.clk(gclk));
	jdff dff_B_xHl8NOXM2_0(.din(w_dff_B_PISKIqu05_0),.dout(w_dff_B_xHl8NOXM2_0),.clk(gclk));
	jdff dff_B_lJWcNF2S1_0(.din(w_dff_B_xHl8NOXM2_0),.dout(w_dff_B_lJWcNF2S1_0),.clk(gclk));
	jdff dff_B_NjINS3uI3_0(.din(w_dff_B_lJWcNF2S1_0),.dout(w_dff_B_NjINS3uI3_0),.clk(gclk));
	jdff dff_B_wlpGhfkl6_0(.din(w_dff_B_NjINS3uI3_0),.dout(w_dff_B_wlpGhfkl6_0),.clk(gclk));
	jdff dff_B_v4RJQEfZ1_0(.din(w_dff_B_wlpGhfkl6_0),.dout(w_dff_B_v4RJQEfZ1_0),.clk(gclk));
	jdff dff_B_OykUYMHQ7_0(.din(w_dff_B_v4RJQEfZ1_0),.dout(w_dff_B_OykUYMHQ7_0),.clk(gclk));
	jdff dff_B_WPxIS6nV9_0(.din(w_dff_B_OykUYMHQ7_0),.dout(w_dff_B_WPxIS6nV9_0),.clk(gclk));
	jdff dff_B_y2gUNXh91_0(.din(w_dff_B_WPxIS6nV9_0),.dout(w_dff_B_y2gUNXh91_0),.clk(gclk));
	jdff dff_B_qhYrMvwl3_0(.din(w_dff_B_y2gUNXh91_0),.dout(w_dff_B_qhYrMvwl3_0),.clk(gclk));
	jdff dff_B_QibSu3MY0_0(.din(w_dff_B_qhYrMvwl3_0),.dout(w_dff_B_QibSu3MY0_0),.clk(gclk));
	jdff dff_B_CrpXcl3L2_0(.din(w_dff_B_QibSu3MY0_0),.dout(w_dff_B_CrpXcl3L2_0),.clk(gclk));
	jdff dff_B_XpzuIzld0_0(.din(w_dff_B_CrpXcl3L2_0),.dout(w_dff_B_XpzuIzld0_0),.clk(gclk));
	jdff dff_B_dAExRaPu8_0(.din(w_dff_B_XpzuIzld0_0),.dout(w_dff_B_dAExRaPu8_0),.clk(gclk));
	jdff dff_B_CbTwYaLV0_0(.din(w_dff_B_dAExRaPu8_0),.dout(w_dff_B_CbTwYaLV0_0),.clk(gclk));
	jdff dff_B_fv8mqUCh1_0(.din(w_dff_B_CbTwYaLV0_0),.dout(w_dff_B_fv8mqUCh1_0),.clk(gclk));
	jdff dff_B_89q5qkTY6_0(.din(w_dff_B_fv8mqUCh1_0),.dout(w_dff_B_89q5qkTY6_0),.clk(gclk));
	jdff dff_B_Jn5J4HWP8_0(.din(w_dff_B_89q5qkTY6_0),.dout(w_dff_B_Jn5J4HWP8_0),.clk(gclk));
	jdff dff_B_tS5qMp922_0(.din(w_dff_B_Jn5J4HWP8_0),.dout(w_dff_B_tS5qMp922_0),.clk(gclk));
	jdff dff_B_XYkhcZ5o5_0(.din(w_dff_B_tS5qMp922_0),.dout(w_dff_B_XYkhcZ5o5_0),.clk(gclk));
	jdff dff_B_5oKoSGR99_0(.din(w_dff_B_XYkhcZ5o5_0),.dout(w_dff_B_5oKoSGR99_0),.clk(gclk));
	jdff dff_B_e0jBCEhW3_0(.din(w_dff_B_5oKoSGR99_0),.dout(w_dff_B_e0jBCEhW3_0),.clk(gclk));
	jdff dff_B_4wpRwwEq3_0(.din(w_dff_B_e0jBCEhW3_0),.dout(w_dff_B_4wpRwwEq3_0),.clk(gclk));
	jdff dff_B_ymYVUOHL6_0(.din(w_dff_B_4wpRwwEq3_0),.dout(w_dff_B_ymYVUOHL6_0),.clk(gclk));
	jdff dff_B_Vw6llRE23_0(.din(w_dff_B_ymYVUOHL6_0),.dout(w_dff_B_Vw6llRE23_0),.clk(gclk));
	jdff dff_B_PGzrBREj0_0(.din(w_dff_B_Vw6llRE23_0),.dout(w_dff_B_PGzrBREj0_0),.clk(gclk));
	jdff dff_B_pNTLlTIs9_0(.din(w_dff_B_PGzrBREj0_0),.dout(w_dff_B_pNTLlTIs9_0),.clk(gclk));
	jdff dff_B_Hgrqy4jd9_0(.din(w_dff_B_pNTLlTIs9_0),.dout(w_dff_B_Hgrqy4jd9_0),.clk(gclk));
	jdff dff_B_VvfcyPt59_0(.din(w_dff_B_Hgrqy4jd9_0),.dout(w_dff_B_VvfcyPt59_0),.clk(gclk));
	jdff dff_B_eeyNjUxG1_0(.din(w_dff_B_VvfcyPt59_0),.dout(w_dff_B_eeyNjUxG1_0),.clk(gclk));
	jdff dff_B_u6K5nWz25_0(.din(w_dff_B_eeyNjUxG1_0),.dout(w_dff_B_u6K5nWz25_0),.clk(gclk));
	jdff dff_B_pHriOpf62_0(.din(w_dff_B_u6K5nWz25_0),.dout(w_dff_B_pHriOpf62_0),.clk(gclk));
	jdff dff_B_Ta2w5qNi1_0(.din(w_dff_B_pHriOpf62_0),.dout(w_dff_B_Ta2w5qNi1_0),.clk(gclk));
	jdff dff_B_pZiIGT1H6_0(.din(w_dff_B_Ta2w5qNi1_0),.dout(w_dff_B_pZiIGT1H6_0),.clk(gclk));
	jdff dff_B_hj2McUWr9_0(.din(w_dff_B_pZiIGT1H6_0),.dout(w_dff_B_hj2McUWr9_0),.clk(gclk));
	jdff dff_B_K1KhT9JZ7_0(.din(w_dff_B_hj2McUWr9_0),.dout(w_dff_B_K1KhT9JZ7_0),.clk(gclk));
	jdff dff_B_YeW3yzi12_0(.din(w_dff_B_K1KhT9JZ7_0),.dout(w_dff_B_YeW3yzi12_0),.clk(gclk));
	jdff dff_B_FHk8Cm157_0(.din(n1000),.dout(w_dff_B_FHk8Cm157_0),.clk(gclk));
	jdff dff_B_3diL9t954_0(.din(w_dff_B_FHk8Cm157_0),.dout(w_dff_B_3diL9t954_0),.clk(gclk));
	jdff dff_B_CK8pLLj75_0(.din(w_dff_B_3diL9t954_0),.dout(w_dff_B_CK8pLLj75_0),.clk(gclk));
	jdff dff_B_OWI6VM5D4_0(.din(w_dff_B_CK8pLLj75_0),.dout(w_dff_B_OWI6VM5D4_0),.clk(gclk));
	jdff dff_B_T0tTv2gd1_0(.din(w_dff_B_OWI6VM5D4_0),.dout(w_dff_B_T0tTv2gd1_0),.clk(gclk));
	jdff dff_B_GoTtdasZ9_0(.din(w_dff_B_T0tTv2gd1_0),.dout(w_dff_B_GoTtdasZ9_0),.clk(gclk));
	jdff dff_B_JZ0JOwL22_0(.din(w_dff_B_GoTtdasZ9_0),.dout(w_dff_B_JZ0JOwL22_0),.clk(gclk));
	jdff dff_B_ePoI6xiD8_0(.din(w_dff_B_JZ0JOwL22_0),.dout(w_dff_B_ePoI6xiD8_0),.clk(gclk));
	jdff dff_B_k6da1RbX4_0(.din(w_dff_B_ePoI6xiD8_0),.dout(w_dff_B_k6da1RbX4_0),.clk(gclk));
	jdff dff_B_jaMlvBPg1_0(.din(w_dff_B_k6da1RbX4_0),.dout(w_dff_B_jaMlvBPg1_0),.clk(gclk));
	jdff dff_B_fVVQV1n03_0(.din(w_dff_B_jaMlvBPg1_0),.dout(w_dff_B_fVVQV1n03_0),.clk(gclk));
	jdff dff_B_j4anH7x76_0(.din(w_dff_B_fVVQV1n03_0),.dout(w_dff_B_j4anH7x76_0),.clk(gclk));
	jdff dff_B_Wd8YoPrp2_0(.din(w_dff_B_j4anH7x76_0),.dout(w_dff_B_Wd8YoPrp2_0),.clk(gclk));
	jdff dff_B_XunoqiqL6_0(.din(w_dff_B_Wd8YoPrp2_0),.dout(w_dff_B_XunoqiqL6_0),.clk(gclk));
	jdff dff_B_zt26dltR8_0(.din(w_dff_B_XunoqiqL6_0),.dout(w_dff_B_zt26dltR8_0),.clk(gclk));
	jdff dff_B_MHc159FP6_0(.din(w_dff_B_zt26dltR8_0),.dout(w_dff_B_MHc159FP6_0),.clk(gclk));
	jdff dff_B_OlSTHSpf3_0(.din(w_dff_B_MHc159FP6_0),.dout(w_dff_B_OlSTHSpf3_0),.clk(gclk));
	jdff dff_B_4jV0ufxc0_0(.din(w_dff_B_OlSTHSpf3_0),.dout(w_dff_B_4jV0ufxc0_0),.clk(gclk));
	jdff dff_B_TG7EVUyF9_0(.din(w_dff_B_4jV0ufxc0_0),.dout(w_dff_B_TG7EVUyF9_0),.clk(gclk));
	jdff dff_B_gaWTXJfm1_0(.din(w_dff_B_TG7EVUyF9_0),.dout(w_dff_B_gaWTXJfm1_0),.clk(gclk));
	jdff dff_B_gQNYQKJR8_0(.din(w_dff_B_gaWTXJfm1_0),.dout(w_dff_B_gQNYQKJR8_0),.clk(gclk));
	jdff dff_B_FlbRwU2r1_0(.din(w_dff_B_gQNYQKJR8_0),.dout(w_dff_B_FlbRwU2r1_0),.clk(gclk));
	jdff dff_B_mX2v2CdV1_0(.din(w_dff_B_FlbRwU2r1_0),.dout(w_dff_B_mX2v2CdV1_0),.clk(gclk));
	jdff dff_B_OXjDVGjo3_0(.din(w_dff_B_mX2v2CdV1_0),.dout(w_dff_B_OXjDVGjo3_0),.clk(gclk));
	jdff dff_B_wKVifQ5f3_0(.din(w_dff_B_OXjDVGjo3_0),.dout(w_dff_B_wKVifQ5f3_0),.clk(gclk));
	jdff dff_B_1s8CBTXJ6_0(.din(w_dff_B_wKVifQ5f3_0),.dout(w_dff_B_1s8CBTXJ6_0),.clk(gclk));
	jdff dff_B_PWFs6dZC6_0(.din(w_dff_B_1s8CBTXJ6_0),.dout(w_dff_B_PWFs6dZC6_0),.clk(gclk));
	jdff dff_B_iCdOhtuk0_0(.din(w_dff_B_PWFs6dZC6_0),.dout(w_dff_B_iCdOhtuk0_0),.clk(gclk));
	jdff dff_B_EhGyXncz5_0(.din(w_dff_B_iCdOhtuk0_0),.dout(w_dff_B_EhGyXncz5_0),.clk(gclk));
	jdff dff_B_xUKp0f8C8_0(.din(w_dff_B_EhGyXncz5_0),.dout(w_dff_B_xUKp0f8C8_0),.clk(gclk));
	jdff dff_B_X80eaCwq1_0(.din(w_dff_B_xUKp0f8C8_0),.dout(w_dff_B_X80eaCwq1_0),.clk(gclk));
	jdff dff_B_jiRS4z6o0_0(.din(w_dff_B_X80eaCwq1_0),.dout(w_dff_B_jiRS4z6o0_0),.clk(gclk));
	jdff dff_B_tSNFly4b2_0(.din(w_dff_B_jiRS4z6o0_0),.dout(w_dff_B_tSNFly4b2_0),.clk(gclk));
	jdff dff_B_VghliOnV8_0(.din(w_dff_B_tSNFly4b2_0),.dout(w_dff_B_VghliOnV8_0),.clk(gclk));
	jdff dff_B_yEEv1zRe9_0(.din(w_dff_B_VghliOnV8_0),.dout(w_dff_B_yEEv1zRe9_0),.clk(gclk));
	jdff dff_B_F5HqIpao2_0(.din(w_dff_B_yEEv1zRe9_0),.dout(w_dff_B_F5HqIpao2_0),.clk(gclk));
	jdff dff_B_c52XXpUA5_0(.din(w_dff_B_F5HqIpao2_0),.dout(w_dff_B_c52XXpUA5_0),.clk(gclk));
	jdff dff_B_0cXD8FQ38_0(.din(w_dff_B_c52XXpUA5_0),.dout(w_dff_B_0cXD8FQ38_0),.clk(gclk));
	jdff dff_B_LNcVVJ9d0_0(.din(w_dff_B_0cXD8FQ38_0),.dout(w_dff_B_LNcVVJ9d0_0),.clk(gclk));
	jdff dff_B_RU6yi0Qa3_0(.din(w_dff_B_LNcVVJ9d0_0),.dout(w_dff_B_RU6yi0Qa3_0),.clk(gclk));
	jdff dff_B_q09krvnU6_0(.din(w_dff_B_RU6yi0Qa3_0),.dout(w_dff_B_q09krvnU6_0),.clk(gclk));
	jdff dff_B_0fo4sWsv3_0(.din(w_dff_B_q09krvnU6_0),.dout(w_dff_B_0fo4sWsv3_0),.clk(gclk));
	jdff dff_B_Lh9Y4DgO6_0(.din(w_dff_B_0fo4sWsv3_0),.dout(w_dff_B_Lh9Y4DgO6_0),.clk(gclk));
	jdff dff_B_fxLWi57l9_0(.din(w_dff_B_Lh9Y4DgO6_0),.dout(w_dff_B_fxLWi57l9_0),.clk(gclk));
	jdff dff_B_y3sNygWR4_0(.din(w_dff_B_fxLWi57l9_0),.dout(w_dff_B_y3sNygWR4_0),.clk(gclk));
	jdff dff_B_EGbb2BET2_0(.din(w_dff_B_y3sNygWR4_0),.dout(w_dff_B_EGbb2BET2_0),.clk(gclk));
	jdff dff_B_49lUd3Sc1_0(.din(w_dff_B_EGbb2BET2_0),.dout(w_dff_B_49lUd3Sc1_0),.clk(gclk));
	jdff dff_B_oXqwIjFO6_0(.din(w_dff_B_49lUd3Sc1_0),.dout(w_dff_B_oXqwIjFO6_0),.clk(gclk));
	jdff dff_B_2wnl7G8F9_0(.din(w_dff_B_oXqwIjFO6_0),.dout(w_dff_B_2wnl7G8F9_0),.clk(gclk));
	jdff dff_B_vPkjnst92_0(.din(w_dff_B_2wnl7G8F9_0),.dout(w_dff_B_vPkjnst92_0),.clk(gclk));
	jdff dff_B_tAmjocYI1_0(.din(w_dff_B_vPkjnst92_0),.dout(w_dff_B_tAmjocYI1_0),.clk(gclk));
	jdff dff_B_j1i98p4f2_0(.din(w_dff_B_tAmjocYI1_0),.dout(w_dff_B_j1i98p4f2_0),.clk(gclk));
	jdff dff_B_ehXNnoXo2_0(.din(w_dff_B_j1i98p4f2_0),.dout(w_dff_B_ehXNnoXo2_0),.clk(gclk));
	jdff dff_B_RcTolzv66_0(.din(w_dff_B_ehXNnoXo2_0),.dout(w_dff_B_RcTolzv66_0),.clk(gclk));
	jdff dff_B_oDb0BsKV0_0(.din(w_dff_B_RcTolzv66_0),.dout(w_dff_B_oDb0BsKV0_0),.clk(gclk));
	jdff dff_B_dcP9bSpQ5_0(.din(w_dff_B_oDb0BsKV0_0),.dout(w_dff_B_dcP9bSpQ5_0),.clk(gclk));
	jdff dff_B_FAGp2f471_0(.din(w_dff_B_dcP9bSpQ5_0),.dout(w_dff_B_FAGp2f471_0),.clk(gclk));
	jdff dff_B_eqmpm2GS2_0(.din(w_dff_B_FAGp2f471_0),.dout(w_dff_B_eqmpm2GS2_0),.clk(gclk));
	jdff dff_B_frSjzcuQ7_0(.din(w_dff_B_eqmpm2GS2_0),.dout(w_dff_B_frSjzcuQ7_0),.clk(gclk));
	jdff dff_B_vaFtvecJ7_0(.din(w_dff_B_frSjzcuQ7_0),.dout(w_dff_B_vaFtvecJ7_0),.clk(gclk));
	jdff dff_B_573kwaHL6_0(.din(w_dff_B_vaFtvecJ7_0),.dout(w_dff_B_573kwaHL6_0),.clk(gclk));
	jdff dff_B_KD4ObqjU1_0(.din(w_dff_B_573kwaHL6_0),.dout(w_dff_B_KD4ObqjU1_0),.clk(gclk));
	jdff dff_B_QA0shmqH6_0(.din(w_dff_B_KD4ObqjU1_0),.dout(w_dff_B_QA0shmqH6_0),.clk(gclk));
	jdff dff_B_R1KPK5NJ0_0(.din(w_dff_B_QA0shmqH6_0),.dout(w_dff_B_R1KPK5NJ0_0),.clk(gclk));
	jdff dff_B_lQzeQN2u2_0(.din(w_dff_B_R1KPK5NJ0_0),.dout(w_dff_B_lQzeQN2u2_0),.clk(gclk));
	jdff dff_B_XP6iymHU6_0(.din(w_dff_B_lQzeQN2u2_0),.dout(w_dff_B_XP6iymHU6_0),.clk(gclk));
	jdff dff_B_frHC1SBb8_0(.din(w_dff_B_XP6iymHU6_0),.dout(w_dff_B_frHC1SBb8_0),.clk(gclk));
	jdff dff_B_31GTaWVV9_0(.din(w_dff_B_frHC1SBb8_0),.dout(w_dff_B_31GTaWVV9_0),.clk(gclk));
	jdff dff_B_W2uokUDX2_0(.din(w_dff_B_31GTaWVV9_0),.dout(w_dff_B_W2uokUDX2_0),.clk(gclk));
	jdff dff_B_XiXwICzV1_0(.din(w_dff_B_W2uokUDX2_0),.dout(w_dff_B_XiXwICzV1_0),.clk(gclk));
	jdff dff_B_0QqotNMq2_0(.din(w_dff_B_XiXwICzV1_0),.dout(w_dff_B_0QqotNMq2_0),.clk(gclk));
	jdff dff_B_zByqVL7c6_0(.din(w_dff_B_0QqotNMq2_0),.dout(w_dff_B_zByqVL7c6_0),.clk(gclk));
	jdff dff_B_eRYks9G98_0(.din(w_dff_B_zByqVL7c6_0),.dout(w_dff_B_eRYks9G98_0),.clk(gclk));
	jdff dff_B_LdPmKlDJ3_0(.din(w_dff_B_eRYks9G98_0),.dout(w_dff_B_LdPmKlDJ3_0),.clk(gclk));
	jdff dff_B_sfLimVBe8_0(.din(w_dff_B_LdPmKlDJ3_0),.dout(w_dff_B_sfLimVBe8_0),.clk(gclk));
	jdff dff_B_VIj0WmHF4_0(.din(w_dff_B_sfLimVBe8_0),.dout(w_dff_B_VIj0WmHF4_0),.clk(gclk));
	jdff dff_B_QdNx6xj44_0(.din(w_dff_B_VIj0WmHF4_0),.dout(w_dff_B_QdNx6xj44_0),.clk(gclk));
	jdff dff_B_wEb8Cs8S4_0(.din(w_dff_B_QdNx6xj44_0),.dout(w_dff_B_wEb8Cs8S4_0),.clk(gclk));
	jdff dff_B_MTgufgRd8_0(.din(w_dff_B_wEb8Cs8S4_0),.dout(w_dff_B_MTgufgRd8_0),.clk(gclk));
	jdff dff_B_hJv1keCv8_0(.din(w_dff_B_MTgufgRd8_0),.dout(w_dff_B_hJv1keCv8_0),.clk(gclk));
	jdff dff_B_MnU9pBJ17_0(.din(w_dff_B_hJv1keCv8_0),.dout(w_dff_B_MnU9pBJ17_0),.clk(gclk));
	jdff dff_B_yJ8aqfJh2_0(.din(w_dff_B_MnU9pBJ17_0),.dout(w_dff_B_yJ8aqfJh2_0),.clk(gclk));
	jdff dff_B_prLBWnEz1_0(.din(w_dff_B_yJ8aqfJh2_0),.dout(w_dff_B_prLBWnEz1_0),.clk(gclk));
	jdff dff_B_hjICNjmV5_0(.din(w_dff_B_prLBWnEz1_0),.dout(w_dff_B_hjICNjmV5_0),.clk(gclk));
	jdff dff_B_5ZnERbT50_0(.din(w_dff_B_hjICNjmV5_0),.dout(w_dff_B_5ZnERbT50_0),.clk(gclk));
	jdff dff_B_cVKHtW8N3_0(.din(w_dff_B_5ZnERbT50_0),.dout(w_dff_B_cVKHtW8N3_0),.clk(gclk));
	jdff dff_B_UlkkA3XK1_0(.din(w_dff_B_cVKHtW8N3_0),.dout(w_dff_B_UlkkA3XK1_0),.clk(gclk));
	jdff dff_B_de56BOYi1_0(.din(w_dff_B_UlkkA3XK1_0),.dout(w_dff_B_de56BOYi1_0),.clk(gclk));
	jdff dff_B_1cD3vLbb4_0(.din(w_dff_B_de56BOYi1_0),.dout(w_dff_B_1cD3vLbb4_0),.clk(gclk));
	jdff dff_B_RYSkFlHW0_0(.din(w_dff_B_1cD3vLbb4_0),.dout(w_dff_B_RYSkFlHW0_0),.clk(gclk));
	jdff dff_B_epEwuMPm3_0(.din(w_dff_B_RYSkFlHW0_0),.dout(w_dff_B_epEwuMPm3_0),.clk(gclk));
	jdff dff_B_LKugcwPw5_0(.din(w_dff_B_epEwuMPm3_0),.dout(w_dff_B_LKugcwPw5_0),.clk(gclk));
	jdff dff_B_A71mZpmU4_0(.din(w_dff_B_LKugcwPw5_0),.dout(w_dff_B_A71mZpmU4_0),.clk(gclk));
	jdff dff_B_z3akaDy54_0(.din(w_dff_B_A71mZpmU4_0),.dout(w_dff_B_z3akaDy54_0),.clk(gclk));
	jdff dff_B_PKlVr9y60_0(.din(w_dff_B_z3akaDy54_0),.dout(w_dff_B_PKlVr9y60_0),.clk(gclk));
	jdff dff_B_H1Ismx8S3_0(.din(w_dff_B_PKlVr9y60_0),.dout(w_dff_B_H1Ismx8S3_0),.clk(gclk));
	jdff dff_B_ktnydPjl3_0(.din(w_dff_B_H1Ismx8S3_0),.dout(w_dff_B_ktnydPjl3_0),.clk(gclk));
	jdff dff_B_W3Qac7z77_0(.din(w_dff_B_ktnydPjl3_0),.dout(w_dff_B_W3Qac7z77_0),.clk(gclk));
	jdff dff_B_R9mKPtUn2_0(.din(w_dff_B_W3Qac7z77_0),.dout(w_dff_B_R9mKPtUn2_0),.clk(gclk));
	jdff dff_B_F2p7XeCT4_0(.din(w_dff_B_R9mKPtUn2_0),.dout(w_dff_B_F2p7XeCT4_0),.clk(gclk));
	jdff dff_B_m2GGTYQT1_0(.din(w_dff_B_F2p7XeCT4_0),.dout(w_dff_B_m2GGTYQT1_0),.clk(gclk));
	jdff dff_B_aQY9Vmue7_0(.din(w_dff_B_m2GGTYQT1_0),.dout(w_dff_B_aQY9Vmue7_0),.clk(gclk));
	jdff dff_B_xGN0Qqyt1_0(.din(n1006),.dout(w_dff_B_xGN0Qqyt1_0),.clk(gclk));
	jdff dff_B_fiuvY00G3_0(.din(w_dff_B_xGN0Qqyt1_0),.dout(w_dff_B_fiuvY00G3_0),.clk(gclk));
	jdff dff_B_aHO5VoQR0_0(.din(w_dff_B_fiuvY00G3_0),.dout(w_dff_B_aHO5VoQR0_0),.clk(gclk));
	jdff dff_B_xQiSzY7V8_0(.din(w_dff_B_aHO5VoQR0_0),.dout(w_dff_B_xQiSzY7V8_0),.clk(gclk));
	jdff dff_B_iZFrfk9X7_0(.din(w_dff_B_xQiSzY7V8_0),.dout(w_dff_B_iZFrfk9X7_0),.clk(gclk));
	jdff dff_B_5OkbODOr5_0(.din(w_dff_B_iZFrfk9X7_0),.dout(w_dff_B_5OkbODOr5_0),.clk(gclk));
	jdff dff_B_q7LqM9db3_0(.din(w_dff_B_5OkbODOr5_0),.dout(w_dff_B_q7LqM9db3_0),.clk(gclk));
	jdff dff_B_JYo2tjZt9_0(.din(w_dff_B_q7LqM9db3_0),.dout(w_dff_B_JYo2tjZt9_0),.clk(gclk));
	jdff dff_B_BNeCqfF61_0(.din(w_dff_B_JYo2tjZt9_0),.dout(w_dff_B_BNeCqfF61_0),.clk(gclk));
	jdff dff_B_lOIOhChm2_0(.din(w_dff_B_BNeCqfF61_0),.dout(w_dff_B_lOIOhChm2_0),.clk(gclk));
	jdff dff_B_QURScThB4_0(.din(w_dff_B_lOIOhChm2_0),.dout(w_dff_B_QURScThB4_0),.clk(gclk));
	jdff dff_B_ALmUfoUf8_0(.din(w_dff_B_QURScThB4_0),.dout(w_dff_B_ALmUfoUf8_0),.clk(gclk));
	jdff dff_B_a5BqRznn5_0(.din(w_dff_B_ALmUfoUf8_0),.dout(w_dff_B_a5BqRznn5_0),.clk(gclk));
	jdff dff_B_VE4kZJhC9_0(.din(w_dff_B_a5BqRznn5_0),.dout(w_dff_B_VE4kZJhC9_0),.clk(gclk));
	jdff dff_B_j4MSl7Rl9_0(.din(w_dff_B_VE4kZJhC9_0),.dout(w_dff_B_j4MSl7Rl9_0),.clk(gclk));
	jdff dff_B_C7b4GfIv0_0(.din(w_dff_B_j4MSl7Rl9_0),.dout(w_dff_B_C7b4GfIv0_0),.clk(gclk));
	jdff dff_B_V6i0CRwj5_0(.din(w_dff_B_C7b4GfIv0_0),.dout(w_dff_B_V6i0CRwj5_0),.clk(gclk));
	jdff dff_B_1sZ7BzvQ7_0(.din(w_dff_B_V6i0CRwj5_0),.dout(w_dff_B_1sZ7BzvQ7_0),.clk(gclk));
	jdff dff_B_ZnChadNt0_0(.din(w_dff_B_1sZ7BzvQ7_0),.dout(w_dff_B_ZnChadNt0_0),.clk(gclk));
	jdff dff_B_qQaYDmDp7_0(.din(w_dff_B_ZnChadNt0_0),.dout(w_dff_B_qQaYDmDp7_0),.clk(gclk));
	jdff dff_B_G2hJzBq82_0(.din(w_dff_B_qQaYDmDp7_0),.dout(w_dff_B_G2hJzBq82_0),.clk(gclk));
	jdff dff_B_Ycgvm1YK5_0(.din(w_dff_B_G2hJzBq82_0),.dout(w_dff_B_Ycgvm1YK5_0),.clk(gclk));
	jdff dff_B_C33CuETS7_0(.din(w_dff_B_Ycgvm1YK5_0),.dout(w_dff_B_C33CuETS7_0),.clk(gclk));
	jdff dff_B_yPPObXP35_0(.din(w_dff_B_C33CuETS7_0),.dout(w_dff_B_yPPObXP35_0),.clk(gclk));
	jdff dff_B_tn4ZeCnK3_0(.din(w_dff_B_yPPObXP35_0),.dout(w_dff_B_tn4ZeCnK3_0),.clk(gclk));
	jdff dff_B_pRYBAsFm7_0(.din(w_dff_B_tn4ZeCnK3_0),.dout(w_dff_B_pRYBAsFm7_0),.clk(gclk));
	jdff dff_B_IrTON0Rr9_0(.din(w_dff_B_pRYBAsFm7_0),.dout(w_dff_B_IrTON0Rr9_0),.clk(gclk));
	jdff dff_B_2Y63atFT6_0(.din(w_dff_B_IrTON0Rr9_0),.dout(w_dff_B_2Y63atFT6_0),.clk(gclk));
	jdff dff_B_rQNt04901_0(.din(w_dff_B_2Y63atFT6_0),.dout(w_dff_B_rQNt04901_0),.clk(gclk));
	jdff dff_B_JSfahvmV3_0(.din(w_dff_B_rQNt04901_0),.dout(w_dff_B_JSfahvmV3_0),.clk(gclk));
	jdff dff_B_IikKiVcf9_0(.din(w_dff_B_JSfahvmV3_0),.dout(w_dff_B_IikKiVcf9_0),.clk(gclk));
	jdff dff_B_ribwdkTf7_0(.din(w_dff_B_IikKiVcf9_0),.dout(w_dff_B_ribwdkTf7_0),.clk(gclk));
	jdff dff_B_pmANmI7m5_0(.din(w_dff_B_ribwdkTf7_0),.dout(w_dff_B_pmANmI7m5_0),.clk(gclk));
	jdff dff_B_37boURr84_0(.din(w_dff_B_pmANmI7m5_0),.dout(w_dff_B_37boURr84_0),.clk(gclk));
	jdff dff_B_oNmT3o6l0_0(.din(w_dff_B_37boURr84_0),.dout(w_dff_B_oNmT3o6l0_0),.clk(gclk));
	jdff dff_B_Yt4gJOsA6_0(.din(w_dff_B_oNmT3o6l0_0),.dout(w_dff_B_Yt4gJOsA6_0),.clk(gclk));
	jdff dff_B_96cPcaDV0_0(.din(w_dff_B_Yt4gJOsA6_0),.dout(w_dff_B_96cPcaDV0_0),.clk(gclk));
	jdff dff_B_JtbCCNnA0_0(.din(w_dff_B_96cPcaDV0_0),.dout(w_dff_B_JtbCCNnA0_0),.clk(gclk));
	jdff dff_B_T0jVaiTr8_0(.din(w_dff_B_JtbCCNnA0_0),.dout(w_dff_B_T0jVaiTr8_0),.clk(gclk));
	jdff dff_B_AeZXTDz20_0(.din(w_dff_B_T0jVaiTr8_0),.dout(w_dff_B_AeZXTDz20_0),.clk(gclk));
	jdff dff_B_LBHc8Nmn0_0(.din(w_dff_B_AeZXTDz20_0),.dout(w_dff_B_LBHc8Nmn0_0),.clk(gclk));
	jdff dff_B_NrqR9U6x4_0(.din(w_dff_B_LBHc8Nmn0_0),.dout(w_dff_B_NrqR9U6x4_0),.clk(gclk));
	jdff dff_B_7D8Ni5ge8_0(.din(w_dff_B_NrqR9U6x4_0),.dout(w_dff_B_7D8Ni5ge8_0),.clk(gclk));
	jdff dff_B_iV2cyu5Y3_0(.din(w_dff_B_7D8Ni5ge8_0),.dout(w_dff_B_iV2cyu5Y3_0),.clk(gclk));
	jdff dff_B_xaTPwzlo0_0(.din(w_dff_B_iV2cyu5Y3_0),.dout(w_dff_B_xaTPwzlo0_0),.clk(gclk));
	jdff dff_B_1WGYhbD68_0(.din(w_dff_B_xaTPwzlo0_0),.dout(w_dff_B_1WGYhbD68_0),.clk(gclk));
	jdff dff_B_l42Cru9g5_0(.din(w_dff_B_1WGYhbD68_0),.dout(w_dff_B_l42Cru9g5_0),.clk(gclk));
	jdff dff_B_LrX6lbra8_0(.din(w_dff_B_l42Cru9g5_0),.dout(w_dff_B_LrX6lbra8_0),.clk(gclk));
	jdff dff_B_bGSFoYhO9_0(.din(w_dff_B_LrX6lbra8_0),.dout(w_dff_B_bGSFoYhO9_0),.clk(gclk));
	jdff dff_B_saKLDtS28_0(.din(w_dff_B_bGSFoYhO9_0),.dout(w_dff_B_saKLDtS28_0),.clk(gclk));
	jdff dff_B_6A7hocPr3_0(.din(w_dff_B_saKLDtS28_0),.dout(w_dff_B_6A7hocPr3_0),.clk(gclk));
	jdff dff_B_yCU0xiTF1_0(.din(w_dff_B_6A7hocPr3_0),.dout(w_dff_B_yCU0xiTF1_0),.clk(gclk));
	jdff dff_B_TtB7TcO89_0(.din(w_dff_B_yCU0xiTF1_0),.dout(w_dff_B_TtB7TcO89_0),.clk(gclk));
	jdff dff_B_pIunSuZN1_0(.din(w_dff_B_TtB7TcO89_0),.dout(w_dff_B_pIunSuZN1_0),.clk(gclk));
	jdff dff_B_KhsCuYaB6_0(.din(w_dff_B_pIunSuZN1_0),.dout(w_dff_B_KhsCuYaB6_0),.clk(gclk));
	jdff dff_B_OcbUrppn6_0(.din(w_dff_B_KhsCuYaB6_0),.dout(w_dff_B_OcbUrppn6_0),.clk(gclk));
	jdff dff_B_PCXjid5C4_0(.din(w_dff_B_OcbUrppn6_0),.dout(w_dff_B_PCXjid5C4_0),.clk(gclk));
	jdff dff_B_y6Eorlus8_0(.din(w_dff_B_PCXjid5C4_0),.dout(w_dff_B_y6Eorlus8_0),.clk(gclk));
	jdff dff_B_owIG0yJ06_0(.din(w_dff_B_y6Eorlus8_0),.dout(w_dff_B_owIG0yJ06_0),.clk(gclk));
	jdff dff_B_Ln4sFxsX2_0(.din(w_dff_B_owIG0yJ06_0),.dout(w_dff_B_Ln4sFxsX2_0),.clk(gclk));
	jdff dff_B_eKwGPw7V8_0(.din(w_dff_B_Ln4sFxsX2_0),.dout(w_dff_B_eKwGPw7V8_0),.clk(gclk));
	jdff dff_B_OlmF5qTe4_0(.din(w_dff_B_eKwGPw7V8_0),.dout(w_dff_B_OlmF5qTe4_0),.clk(gclk));
	jdff dff_B_5SYs1ChX1_0(.din(w_dff_B_OlmF5qTe4_0),.dout(w_dff_B_5SYs1ChX1_0),.clk(gclk));
	jdff dff_B_FOkIB6aE9_0(.din(w_dff_B_5SYs1ChX1_0),.dout(w_dff_B_FOkIB6aE9_0),.clk(gclk));
	jdff dff_B_2xMjHazF1_0(.din(w_dff_B_FOkIB6aE9_0),.dout(w_dff_B_2xMjHazF1_0),.clk(gclk));
	jdff dff_B_ZrCyTODv6_0(.din(w_dff_B_2xMjHazF1_0),.dout(w_dff_B_ZrCyTODv6_0),.clk(gclk));
	jdff dff_B_de0Eltu84_0(.din(w_dff_B_ZrCyTODv6_0),.dout(w_dff_B_de0Eltu84_0),.clk(gclk));
	jdff dff_B_dNu5LnJL2_0(.din(w_dff_B_de0Eltu84_0),.dout(w_dff_B_dNu5LnJL2_0),.clk(gclk));
	jdff dff_B_mAg1Ma4N2_0(.din(w_dff_B_dNu5LnJL2_0),.dout(w_dff_B_mAg1Ma4N2_0),.clk(gclk));
	jdff dff_B_eUV9qe9P0_0(.din(w_dff_B_mAg1Ma4N2_0),.dout(w_dff_B_eUV9qe9P0_0),.clk(gclk));
	jdff dff_B_u4s8MfAV2_0(.din(w_dff_B_eUV9qe9P0_0),.dout(w_dff_B_u4s8MfAV2_0),.clk(gclk));
	jdff dff_B_QI4t88Im4_0(.din(w_dff_B_u4s8MfAV2_0),.dout(w_dff_B_QI4t88Im4_0),.clk(gclk));
	jdff dff_B_3Re7f7gr6_0(.din(w_dff_B_QI4t88Im4_0),.dout(w_dff_B_3Re7f7gr6_0),.clk(gclk));
	jdff dff_B_LrvPmcfc6_0(.din(w_dff_B_3Re7f7gr6_0),.dout(w_dff_B_LrvPmcfc6_0),.clk(gclk));
	jdff dff_B_Jpyr0i3p5_0(.din(w_dff_B_LrvPmcfc6_0),.dout(w_dff_B_Jpyr0i3p5_0),.clk(gclk));
	jdff dff_B_rgNpTVNe8_0(.din(w_dff_B_Jpyr0i3p5_0),.dout(w_dff_B_rgNpTVNe8_0),.clk(gclk));
	jdff dff_B_hRgMZVDQ0_0(.din(w_dff_B_rgNpTVNe8_0),.dout(w_dff_B_hRgMZVDQ0_0),.clk(gclk));
	jdff dff_B_8CMIGMki7_0(.din(w_dff_B_hRgMZVDQ0_0),.dout(w_dff_B_8CMIGMki7_0),.clk(gclk));
	jdff dff_B_8r5sT5Hj9_0(.din(w_dff_B_8CMIGMki7_0),.dout(w_dff_B_8r5sT5Hj9_0),.clk(gclk));
	jdff dff_B_agKJkgO88_0(.din(w_dff_B_8r5sT5Hj9_0),.dout(w_dff_B_agKJkgO88_0),.clk(gclk));
	jdff dff_B_5tUUvYSs5_0(.din(w_dff_B_agKJkgO88_0),.dout(w_dff_B_5tUUvYSs5_0),.clk(gclk));
	jdff dff_B_SUUYl2Ql6_0(.din(w_dff_B_5tUUvYSs5_0),.dout(w_dff_B_SUUYl2Ql6_0),.clk(gclk));
	jdff dff_B_2Kcfu0Ow9_0(.din(w_dff_B_SUUYl2Ql6_0),.dout(w_dff_B_2Kcfu0Ow9_0),.clk(gclk));
	jdff dff_B_V3CPQKV23_0(.din(w_dff_B_2Kcfu0Ow9_0),.dout(w_dff_B_V3CPQKV23_0),.clk(gclk));
	jdff dff_B_h8dfXeo67_0(.din(w_dff_B_V3CPQKV23_0),.dout(w_dff_B_h8dfXeo67_0),.clk(gclk));
	jdff dff_B_6fmHsrpf9_0(.din(w_dff_B_h8dfXeo67_0),.dout(w_dff_B_6fmHsrpf9_0),.clk(gclk));
	jdff dff_B_vv05b3pP6_0(.din(w_dff_B_6fmHsrpf9_0),.dout(w_dff_B_vv05b3pP6_0),.clk(gclk));
	jdff dff_B_iv0OTOHd3_0(.din(w_dff_B_vv05b3pP6_0),.dout(w_dff_B_iv0OTOHd3_0),.clk(gclk));
	jdff dff_B_Lo11yvdl1_0(.din(w_dff_B_iv0OTOHd3_0),.dout(w_dff_B_Lo11yvdl1_0),.clk(gclk));
	jdff dff_B_pCR9Yfr53_0(.din(w_dff_B_Lo11yvdl1_0),.dout(w_dff_B_pCR9Yfr53_0),.clk(gclk));
	jdff dff_B_SPDzZlbu0_0(.din(w_dff_B_pCR9Yfr53_0),.dout(w_dff_B_SPDzZlbu0_0),.clk(gclk));
	jdff dff_B_XMqaOnrd7_0(.din(w_dff_B_SPDzZlbu0_0),.dout(w_dff_B_XMqaOnrd7_0),.clk(gclk));
	jdff dff_B_2FGhGH2k2_0(.din(w_dff_B_XMqaOnrd7_0),.dout(w_dff_B_2FGhGH2k2_0),.clk(gclk));
	jdff dff_B_k6gdoh4L9_0(.din(w_dff_B_2FGhGH2k2_0),.dout(w_dff_B_k6gdoh4L9_0),.clk(gclk));
	jdff dff_B_OEcg16PF4_0(.din(w_dff_B_k6gdoh4L9_0),.dout(w_dff_B_OEcg16PF4_0),.clk(gclk));
	jdff dff_B_VuLpQPGO9_0(.din(w_dff_B_OEcg16PF4_0),.dout(w_dff_B_VuLpQPGO9_0),.clk(gclk));
	jdff dff_B_FrmXP06D2_0(.din(w_dff_B_VuLpQPGO9_0),.dout(w_dff_B_FrmXP06D2_0),.clk(gclk));
	jdff dff_B_geqgFR811_0(.din(w_dff_B_FrmXP06D2_0),.dout(w_dff_B_geqgFR811_0),.clk(gclk));
	jdff dff_B_20cXzEjq0_0(.din(w_dff_B_geqgFR811_0),.dout(w_dff_B_20cXzEjq0_0),.clk(gclk));
	jdff dff_B_moPeNJNd9_0(.din(w_dff_B_20cXzEjq0_0),.dout(w_dff_B_moPeNJNd9_0),.clk(gclk));
	jdff dff_B_N3qEAfNq3_0(.din(w_dff_B_moPeNJNd9_0),.dout(w_dff_B_N3qEAfNq3_0),.clk(gclk));
	jdff dff_B_GtfoM1uq0_0(.din(w_dff_B_N3qEAfNq3_0),.dout(w_dff_B_GtfoM1uq0_0),.clk(gclk));
	jdff dff_B_pmoeat4U0_0(.din(w_dff_B_GtfoM1uq0_0),.dout(w_dff_B_pmoeat4U0_0),.clk(gclk));
	jdff dff_B_E3ZUZcLs9_0(.din(n1012),.dout(w_dff_B_E3ZUZcLs9_0),.clk(gclk));
	jdff dff_B_ehJMKFQM6_0(.din(w_dff_B_E3ZUZcLs9_0),.dout(w_dff_B_ehJMKFQM6_0),.clk(gclk));
	jdff dff_B_3XzqoR0D2_0(.din(w_dff_B_ehJMKFQM6_0),.dout(w_dff_B_3XzqoR0D2_0),.clk(gclk));
	jdff dff_B_ajXEGd817_0(.din(w_dff_B_3XzqoR0D2_0),.dout(w_dff_B_ajXEGd817_0),.clk(gclk));
	jdff dff_B_ZStMTwQe6_0(.din(w_dff_B_ajXEGd817_0),.dout(w_dff_B_ZStMTwQe6_0),.clk(gclk));
	jdff dff_B_q9ucs9dJ6_0(.din(w_dff_B_ZStMTwQe6_0),.dout(w_dff_B_q9ucs9dJ6_0),.clk(gclk));
	jdff dff_B_22wiXwxE9_0(.din(w_dff_B_q9ucs9dJ6_0),.dout(w_dff_B_22wiXwxE9_0),.clk(gclk));
	jdff dff_B_Lk1S6Kbi7_0(.din(w_dff_B_22wiXwxE9_0),.dout(w_dff_B_Lk1S6Kbi7_0),.clk(gclk));
	jdff dff_B_66sgbL4g3_0(.din(w_dff_B_Lk1S6Kbi7_0),.dout(w_dff_B_66sgbL4g3_0),.clk(gclk));
	jdff dff_B_aTILEKEi7_0(.din(w_dff_B_66sgbL4g3_0),.dout(w_dff_B_aTILEKEi7_0),.clk(gclk));
	jdff dff_B_33JP8V1O5_0(.din(w_dff_B_aTILEKEi7_0),.dout(w_dff_B_33JP8V1O5_0),.clk(gclk));
	jdff dff_B_on5EDIln4_0(.din(w_dff_B_33JP8V1O5_0),.dout(w_dff_B_on5EDIln4_0),.clk(gclk));
	jdff dff_B_MR96iNia7_0(.din(w_dff_B_on5EDIln4_0),.dout(w_dff_B_MR96iNia7_0),.clk(gclk));
	jdff dff_B_CDWAS9cZ7_0(.din(w_dff_B_MR96iNia7_0),.dout(w_dff_B_CDWAS9cZ7_0),.clk(gclk));
	jdff dff_B_g9mHbIN76_0(.din(w_dff_B_CDWAS9cZ7_0),.dout(w_dff_B_g9mHbIN76_0),.clk(gclk));
	jdff dff_B_pXakBqg36_0(.din(w_dff_B_g9mHbIN76_0),.dout(w_dff_B_pXakBqg36_0),.clk(gclk));
	jdff dff_B_1KvY9WdL1_0(.din(w_dff_B_pXakBqg36_0),.dout(w_dff_B_1KvY9WdL1_0),.clk(gclk));
	jdff dff_B_AqTpSvBg9_0(.din(w_dff_B_1KvY9WdL1_0),.dout(w_dff_B_AqTpSvBg9_0),.clk(gclk));
	jdff dff_B_ARkWtLDg2_0(.din(w_dff_B_AqTpSvBg9_0),.dout(w_dff_B_ARkWtLDg2_0),.clk(gclk));
	jdff dff_B_RVxQSl9z2_0(.din(w_dff_B_ARkWtLDg2_0),.dout(w_dff_B_RVxQSl9z2_0),.clk(gclk));
	jdff dff_B_MXapfCiO0_0(.din(w_dff_B_RVxQSl9z2_0),.dout(w_dff_B_MXapfCiO0_0),.clk(gclk));
	jdff dff_B_NiJgqczZ6_0(.din(w_dff_B_MXapfCiO0_0),.dout(w_dff_B_NiJgqczZ6_0),.clk(gclk));
	jdff dff_B_pJBJs51D7_0(.din(w_dff_B_NiJgqczZ6_0),.dout(w_dff_B_pJBJs51D7_0),.clk(gclk));
	jdff dff_B_6VXoqg1k7_0(.din(w_dff_B_pJBJs51D7_0),.dout(w_dff_B_6VXoqg1k7_0),.clk(gclk));
	jdff dff_B_a53JGxks9_0(.din(w_dff_B_6VXoqg1k7_0),.dout(w_dff_B_a53JGxks9_0),.clk(gclk));
	jdff dff_B_EvjNB68H3_0(.din(w_dff_B_a53JGxks9_0),.dout(w_dff_B_EvjNB68H3_0),.clk(gclk));
	jdff dff_B_w96ba0o01_0(.din(w_dff_B_EvjNB68H3_0),.dout(w_dff_B_w96ba0o01_0),.clk(gclk));
	jdff dff_B_jBxV5ZP92_0(.din(w_dff_B_w96ba0o01_0),.dout(w_dff_B_jBxV5ZP92_0),.clk(gclk));
	jdff dff_B_KBm0uTY37_0(.din(w_dff_B_jBxV5ZP92_0),.dout(w_dff_B_KBm0uTY37_0),.clk(gclk));
	jdff dff_B_cu6Mvi1O3_0(.din(w_dff_B_KBm0uTY37_0),.dout(w_dff_B_cu6Mvi1O3_0),.clk(gclk));
	jdff dff_B_RHlAZacF5_0(.din(w_dff_B_cu6Mvi1O3_0),.dout(w_dff_B_RHlAZacF5_0),.clk(gclk));
	jdff dff_B_unqY8mlw0_0(.din(w_dff_B_RHlAZacF5_0),.dout(w_dff_B_unqY8mlw0_0),.clk(gclk));
	jdff dff_B_egQMpBlX8_0(.din(w_dff_B_unqY8mlw0_0),.dout(w_dff_B_egQMpBlX8_0),.clk(gclk));
	jdff dff_B_7EMz2fWV0_0(.din(w_dff_B_egQMpBlX8_0),.dout(w_dff_B_7EMz2fWV0_0),.clk(gclk));
	jdff dff_B_frwXzutk5_0(.din(w_dff_B_7EMz2fWV0_0),.dout(w_dff_B_frwXzutk5_0),.clk(gclk));
	jdff dff_B_XoAPZ96H2_0(.din(w_dff_B_frwXzutk5_0),.dout(w_dff_B_XoAPZ96H2_0),.clk(gclk));
	jdff dff_B_VxpdCQyE4_0(.din(w_dff_B_XoAPZ96H2_0),.dout(w_dff_B_VxpdCQyE4_0),.clk(gclk));
	jdff dff_B_5nGgvKrc1_0(.din(w_dff_B_VxpdCQyE4_0),.dout(w_dff_B_5nGgvKrc1_0),.clk(gclk));
	jdff dff_B_EpWcbXQC9_0(.din(w_dff_B_5nGgvKrc1_0),.dout(w_dff_B_EpWcbXQC9_0),.clk(gclk));
	jdff dff_B_ikShCIX86_0(.din(w_dff_B_EpWcbXQC9_0),.dout(w_dff_B_ikShCIX86_0),.clk(gclk));
	jdff dff_B_MDGgDhvE2_0(.din(w_dff_B_ikShCIX86_0),.dout(w_dff_B_MDGgDhvE2_0),.clk(gclk));
	jdff dff_B_uO2yOCfx7_0(.din(w_dff_B_MDGgDhvE2_0),.dout(w_dff_B_uO2yOCfx7_0),.clk(gclk));
	jdff dff_B_AFpSPMYN9_0(.din(w_dff_B_uO2yOCfx7_0),.dout(w_dff_B_AFpSPMYN9_0),.clk(gclk));
	jdff dff_B_cTffIZWH2_0(.din(w_dff_B_AFpSPMYN9_0),.dout(w_dff_B_cTffIZWH2_0),.clk(gclk));
	jdff dff_B_3ECHQIaU1_0(.din(w_dff_B_cTffIZWH2_0),.dout(w_dff_B_3ECHQIaU1_0),.clk(gclk));
	jdff dff_B_F2Lyayif5_0(.din(w_dff_B_3ECHQIaU1_0),.dout(w_dff_B_F2Lyayif5_0),.clk(gclk));
	jdff dff_B_6GcnVHFK3_0(.din(w_dff_B_F2Lyayif5_0),.dout(w_dff_B_6GcnVHFK3_0),.clk(gclk));
	jdff dff_B_z70llqHZ0_0(.din(w_dff_B_6GcnVHFK3_0),.dout(w_dff_B_z70llqHZ0_0),.clk(gclk));
	jdff dff_B_fuXnMRtv2_0(.din(w_dff_B_z70llqHZ0_0),.dout(w_dff_B_fuXnMRtv2_0),.clk(gclk));
	jdff dff_B_UkzBpdJk3_0(.din(w_dff_B_fuXnMRtv2_0),.dout(w_dff_B_UkzBpdJk3_0),.clk(gclk));
	jdff dff_B_1KN2rOI35_0(.din(w_dff_B_UkzBpdJk3_0),.dout(w_dff_B_1KN2rOI35_0),.clk(gclk));
	jdff dff_B_NDLYw4BX6_0(.din(w_dff_B_1KN2rOI35_0),.dout(w_dff_B_NDLYw4BX6_0),.clk(gclk));
	jdff dff_B_4DQBQDm09_0(.din(w_dff_B_NDLYw4BX6_0),.dout(w_dff_B_4DQBQDm09_0),.clk(gclk));
	jdff dff_B_0wTDjqhf0_0(.din(w_dff_B_4DQBQDm09_0),.dout(w_dff_B_0wTDjqhf0_0),.clk(gclk));
	jdff dff_B_wblBllOt5_0(.din(w_dff_B_0wTDjqhf0_0),.dout(w_dff_B_wblBllOt5_0),.clk(gclk));
	jdff dff_B_ZlLBXL0q4_0(.din(w_dff_B_wblBllOt5_0),.dout(w_dff_B_ZlLBXL0q4_0),.clk(gclk));
	jdff dff_B_IvDHNfVi3_0(.din(w_dff_B_ZlLBXL0q4_0),.dout(w_dff_B_IvDHNfVi3_0),.clk(gclk));
	jdff dff_B_aGRkfmxy1_0(.din(w_dff_B_IvDHNfVi3_0),.dout(w_dff_B_aGRkfmxy1_0),.clk(gclk));
	jdff dff_B_tMWeQkwK3_0(.din(w_dff_B_aGRkfmxy1_0),.dout(w_dff_B_tMWeQkwK3_0),.clk(gclk));
	jdff dff_B_7mcESinR8_0(.din(w_dff_B_tMWeQkwK3_0),.dout(w_dff_B_7mcESinR8_0),.clk(gclk));
	jdff dff_B_w75cR5T45_0(.din(w_dff_B_7mcESinR8_0),.dout(w_dff_B_w75cR5T45_0),.clk(gclk));
	jdff dff_B_JgN08Anm3_0(.din(w_dff_B_w75cR5T45_0),.dout(w_dff_B_JgN08Anm3_0),.clk(gclk));
	jdff dff_B_aFyF0oj45_0(.din(w_dff_B_JgN08Anm3_0),.dout(w_dff_B_aFyF0oj45_0),.clk(gclk));
	jdff dff_B_z4yGXYRC6_0(.din(w_dff_B_aFyF0oj45_0),.dout(w_dff_B_z4yGXYRC6_0),.clk(gclk));
	jdff dff_B_NJX6h7iV3_0(.din(w_dff_B_z4yGXYRC6_0),.dout(w_dff_B_NJX6h7iV3_0),.clk(gclk));
	jdff dff_B_jkmHeVEt0_0(.din(w_dff_B_NJX6h7iV3_0),.dout(w_dff_B_jkmHeVEt0_0),.clk(gclk));
	jdff dff_B_M1OaGsg82_0(.din(w_dff_B_jkmHeVEt0_0),.dout(w_dff_B_M1OaGsg82_0),.clk(gclk));
	jdff dff_B_n41gK4eS7_0(.din(w_dff_B_M1OaGsg82_0),.dout(w_dff_B_n41gK4eS7_0),.clk(gclk));
	jdff dff_B_UyrT6NAh6_0(.din(w_dff_B_n41gK4eS7_0),.dout(w_dff_B_UyrT6NAh6_0),.clk(gclk));
	jdff dff_B_9rc0CAUg3_0(.din(w_dff_B_UyrT6NAh6_0),.dout(w_dff_B_9rc0CAUg3_0),.clk(gclk));
	jdff dff_B_pHlugRtT4_0(.din(w_dff_B_9rc0CAUg3_0),.dout(w_dff_B_pHlugRtT4_0),.clk(gclk));
	jdff dff_B_1Nga2AzP5_0(.din(w_dff_B_pHlugRtT4_0),.dout(w_dff_B_1Nga2AzP5_0),.clk(gclk));
	jdff dff_B_m0CZFsE05_0(.din(w_dff_B_1Nga2AzP5_0),.dout(w_dff_B_m0CZFsE05_0),.clk(gclk));
	jdff dff_B_i6zH9xfd3_0(.din(w_dff_B_m0CZFsE05_0),.dout(w_dff_B_i6zH9xfd3_0),.clk(gclk));
	jdff dff_B_cOdCS9p96_0(.din(w_dff_B_i6zH9xfd3_0),.dout(w_dff_B_cOdCS9p96_0),.clk(gclk));
	jdff dff_B_bmx66jTE1_0(.din(w_dff_B_cOdCS9p96_0),.dout(w_dff_B_bmx66jTE1_0),.clk(gclk));
	jdff dff_B_5BYT7Hkh0_0(.din(w_dff_B_bmx66jTE1_0),.dout(w_dff_B_5BYT7Hkh0_0),.clk(gclk));
	jdff dff_B_iQ3YF5Pz9_0(.din(w_dff_B_5BYT7Hkh0_0),.dout(w_dff_B_iQ3YF5Pz9_0),.clk(gclk));
	jdff dff_B_vC48mWBm1_0(.din(w_dff_B_iQ3YF5Pz9_0),.dout(w_dff_B_vC48mWBm1_0),.clk(gclk));
	jdff dff_B_gwewANYg9_0(.din(w_dff_B_vC48mWBm1_0),.dout(w_dff_B_gwewANYg9_0),.clk(gclk));
	jdff dff_B_y0CcsUWT2_0(.din(w_dff_B_gwewANYg9_0),.dout(w_dff_B_y0CcsUWT2_0),.clk(gclk));
	jdff dff_B_15W38iue0_0(.din(w_dff_B_y0CcsUWT2_0),.dout(w_dff_B_15W38iue0_0),.clk(gclk));
	jdff dff_B_AlQcuCud8_0(.din(w_dff_B_15W38iue0_0),.dout(w_dff_B_AlQcuCud8_0),.clk(gclk));
	jdff dff_B_pNiayghy5_0(.din(w_dff_B_AlQcuCud8_0),.dout(w_dff_B_pNiayghy5_0),.clk(gclk));
	jdff dff_B_0QBYYCfx6_0(.din(w_dff_B_pNiayghy5_0),.dout(w_dff_B_0QBYYCfx6_0),.clk(gclk));
	jdff dff_B_kSbs4dz32_0(.din(w_dff_B_0QBYYCfx6_0),.dout(w_dff_B_kSbs4dz32_0),.clk(gclk));
	jdff dff_B_SYPE1Myu0_0(.din(w_dff_B_kSbs4dz32_0),.dout(w_dff_B_SYPE1Myu0_0),.clk(gclk));
	jdff dff_B_gjU2VSrl5_0(.din(w_dff_B_SYPE1Myu0_0),.dout(w_dff_B_gjU2VSrl5_0),.clk(gclk));
	jdff dff_B_gIhryTrY2_0(.din(w_dff_B_gjU2VSrl5_0),.dout(w_dff_B_gIhryTrY2_0),.clk(gclk));
	jdff dff_B_GGTpIqzJ3_0(.din(w_dff_B_gIhryTrY2_0),.dout(w_dff_B_GGTpIqzJ3_0),.clk(gclk));
	jdff dff_B_1sYlDTx17_0(.din(w_dff_B_GGTpIqzJ3_0),.dout(w_dff_B_1sYlDTx17_0),.clk(gclk));
	jdff dff_B_KHzhYfHX4_0(.din(w_dff_B_1sYlDTx17_0),.dout(w_dff_B_KHzhYfHX4_0),.clk(gclk));
	jdff dff_B_sVLdLstf7_0(.din(w_dff_B_KHzhYfHX4_0),.dout(w_dff_B_sVLdLstf7_0),.clk(gclk));
	jdff dff_B_aBDnNtof8_0(.din(w_dff_B_sVLdLstf7_0),.dout(w_dff_B_aBDnNtof8_0),.clk(gclk));
	jdff dff_B_rrcyax9y5_0(.din(w_dff_B_aBDnNtof8_0),.dout(w_dff_B_rrcyax9y5_0),.clk(gclk));
	jdff dff_B_iG7hTRaU5_0(.din(w_dff_B_rrcyax9y5_0),.dout(w_dff_B_iG7hTRaU5_0),.clk(gclk));
	jdff dff_B_7FQBMSLZ2_0(.din(w_dff_B_iG7hTRaU5_0),.dout(w_dff_B_7FQBMSLZ2_0),.clk(gclk));
	jdff dff_B_rrhZqAUJ7_0(.din(w_dff_B_7FQBMSLZ2_0),.dout(w_dff_B_rrhZqAUJ7_0),.clk(gclk));
	jdff dff_B_XAhX8icl7_0(.din(w_dff_B_rrhZqAUJ7_0),.dout(w_dff_B_XAhX8icl7_0),.clk(gclk));
	jdff dff_B_MHuBcaSt0_0(.din(w_dff_B_XAhX8icl7_0),.dout(w_dff_B_MHuBcaSt0_0),.clk(gclk));
	jdff dff_B_WVMFfHbY1_0(.din(w_dff_B_MHuBcaSt0_0),.dout(w_dff_B_WVMFfHbY1_0),.clk(gclk));
	jdff dff_B_o7VqJYbT7_0(.din(w_dff_B_WVMFfHbY1_0),.dout(w_dff_B_o7VqJYbT7_0),.clk(gclk));
	jdff dff_B_SmeeZ4tL6_0(.din(w_dff_B_o7VqJYbT7_0),.dout(w_dff_B_SmeeZ4tL6_0),.clk(gclk));
	jdff dff_B_73IF7KRg3_0(.din(w_dff_B_SmeeZ4tL6_0),.dout(w_dff_B_73IF7KRg3_0),.clk(gclk));
	jdff dff_B_BxbavUD39_0(.din(n1018),.dout(w_dff_B_BxbavUD39_0),.clk(gclk));
	jdff dff_B_CHIrgCrR3_0(.din(w_dff_B_BxbavUD39_0),.dout(w_dff_B_CHIrgCrR3_0),.clk(gclk));
	jdff dff_B_LYTy6ISu5_0(.din(w_dff_B_CHIrgCrR3_0),.dout(w_dff_B_LYTy6ISu5_0),.clk(gclk));
	jdff dff_B_cquNgXv40_0(.din(w_dff_B_LYTy6ISu5_0),.dout(w_dff_B_cquNgXv40_0),.clk(gclk));
	jdff dff_B_HddT7aXK1_0(.din(w_dff_B_cquNgXv40_0),.dout(w_dff_B_HddT7aXK1_0),.clk(gclk));
	jdff dff_B_9yP5DuKQ0_0(.din(w_dff_B_HddT7aXK1_0),.dout(w_dff_B_9yP5DuKQ0_0),.clk(gclk));
	jdff dff_B_PJMw2XNx9_0(.din(w_dff_B_9yP5DuKQ0_0),.dout(w_dff_B_PJMw2XNx9_0),.clk(gclk));
	jdff dff_B_xYQ7Zcz49_0(.din(w_dff_B_PJMw2XNx9_0),.dout(w_dff_B_xYQ7Zcz49_0),.clk(gclk));
	jdff dff_B_OCt7ZsUi7_0(.din(w_dff_B_xYQ7Zcz49_0),.dout(w_dff_B_OCt7ZsUi7_0),.clk(gclk));
	jdff dff_B_vtGN0D4r3_0(.din(w_dff_B_OCt7ZsUi7_0),.dout(w_dff_B_vtGN0D4r3_0),.clk(gclk));
	jdff dff_B_YOwd49Y06_0(.din(w_dff_B_vtGN0D4r3_0),.dout(w_dff_B_YOwd49Y06_0),.clk(gclk));
	jdff dff_B_XFNrNkxe1_0(.din(w_dff_B_YOwd49Y06_0),.dout(w_dff_B_XFNrNkxe1_0),.clk(gclk));
	jdff dff_B_U4mECs0r7_0(.din(w_dff_B_XFNrNkxe1_0),.dout(w_dff_B_U4mECs0r7_0),.clk(gclk));
	jdff dff_B_rXOMJpwB3_0(.din(w_dff_B_U4mECs0r7_0),.dout(w_dff_B_rXOMJpwB3_0),.clk(gclk));
	jdff dff_B_NFllEoXk6_0(.din(w_dff_B_rXOMJpwB3_0),.dout(w_dff_B_NFllEoXk6_0),.clk(gclk));
	jdff dff_B_0QsMHnpL9_0(.din(w_dff_B_NFllEoXk6_0),.dout(w_dff_B_0QsMHnpL9_0),.clk(gclk));
	jdff dff_B_Twnfa97T6_0(.din(w_dff_B_0QsMHnpL9_0),.dout(w_dff_B_Twnfa97T6_0),.clk(gclk));
	jdff dff_B_G6YcFTpg6_0(.din(w_dff_B_Twnfa97T6_0),.dout(w_dff_B_G6YcFTpg6_0),.clk(gclk));
	jdff dff_B_vZZIn7do3_0(.din(w_dff_B_G6YcFTpg6_0),.dout(w_dff_B_vZZIn7do3_0),.clk(gclk));
	jdff dff_B_9azuofPq2_0(.din(w_dff_B_vZZIn7do3_0),.dout(w_dff_B_9azuofPq2_0),.clk(gclk));
	jdff dff_B_URUsk3MO0_0(.din(w_dff_B_9azuofPq2_0),.dout(w_dff_B_URUsk3MO0_0),.clk(gclk));
	jdff dff_B_8wd0pn7A4_0(.din(w_dff_B_URUsk3MO0_0),.dout(w_dff_B_8wd0pn7A4_0),.clk(gclk));
	jdff dff_B_8HpPVXXn4_0(.din(w_dff_B_8wd0pn7A4_0),.dout(w_dff_B_8HpPVXXn4_0),.clk(gclk));
	jdff dff_B_rGoXWfzz2_0(.din(w_dff_B_8HpPVXXn4_0),.dout(w_dff_B_rGoXWfzz2_0),.clk(gclk));
	jdff dff_B_1VWRbAFr3_0(.din(w_dff_B_rGoXWfzz2_0),.dout(w_dff_B_1VWRbAFr3_0),.clk(gclk));
	jdff dff_B_YsYCyOqW2_0(.din(w_dff_B_1VWRbAFr3_0),.dout(w_dff_B_YsYCyOqW2_0),.clk(gclk));
	jdff dff_B_QcCldeJf2_0(.din(w_dff_B_YsYCyOqW2_0),.dout(w_dff_B_QcCldeJf2_0),.clk(gclk));
	jdff dff_B_REoL3ClF6_0(.din(w_dff_B_QcCldeJf2_0),.dout(w_dff_B_REoL3ClF6_0),.clk(gclk));
	jdff dff_B_rPfnGHDG2_0(.din(w_dff_B_REoL3ClF6_0),.dout(w_dff_B_rPfnGHDG2_0),.clk(gclk));
	jdff dff_B_2fmDeasB9_0(.din(w_dff_B_rPfnGHDG2_0),.dout(w_dff_B_2fmDeasB9_0),.clk(gclk));
	jdff dff_B_2I7LxLKF3_0(.din(w_dff_B_2fmDeasB9_0),.dout(w_dff_B_2I7LxLKF3_0),.clk(gclk));
	jdff dff_B_baT2ARg28_0(.din(w_dff_B_2I7LxLKF3_0),.dout(w_dff_B_baT2ARg28_0),.clk(gclk));
	jdff dff_B_i2OGFSEI6_0(.din(w_dff_B_baT2ARg28_0),.dout(w_dff_B_i2OGFSEI6_0),.clk(gclk));
	jdff dff_B_670Xcgpe5_0(.din(w_dff_B_i2OGFSEI6_0),.dout(w_dff_B_670Xcgpe5_0),.clk(gclk));
	jdff dff_B_QKAwfh3j5_0(.din(w_dff_B_670Xcgpe5_0),.dout(w_dff_B_QKAwfh3j5_0),.clk(gclk));
	jdff dff_B_ZAFVuXJo2_0(.din(w_dff_B_QKAwfh3j5_0),.dout(w_dff_B_ZAFVuXJo2_0),.clk(gclk));
	jdff dff_B_h9Owkg0i8_0(.din(w_dff_B_ZAFVuXJo2_0),.dout(w_dff_B_h9Owkg0i8_0),.clk(gclk));
	jdff dff_B_jaV6vv2Y7_0(.din(w_dff_B_h9Owkg0i8_0),.dout(w_dff_B_jaV6vv2Y7_0),.clk(gclk));
	jdff dff_B_SS39PbM01_0(.din(w_dff_B_jaV6vv2Y7_0),.dout(w_dff_B_SS39PbM01_0),.clk(gclk));
	jdff dff_B_0mdxo3WL3_0(.din(w_dff_B_SS39PbM01_0),.dout(w_dff_B_0mdxo3WL3_0),.clk(gclk));
	jdff dff_B_Dsizarx17_0(.din(w_dff_B_0mdxo3WL3_0),.dout(w_dff_B_Dsizarx17_0),.clk(gclk));
	jdff dff_B_LEMRb8hz5_0(.din(w_dff_B_Dsizarx17_0),.dout(w_dff_B_LEMRb8hz5_0),.clk(gclk));
	jdff dff_B_8WRodDgi5_0(.din(w_dff_B_LEMRb8hz5_0),.dout(w_dff_B_8WRodDgi5_0),.clk(gclk));
	jdff dff_B_2IYgpU4x5_0(.din(w_dff_B_8WRodDgi5_0),.dout(w_dff_B_2IYgpU4x5_0),.clk(gclk));
	jdff dff_B_YfZSMbct1_0(.din(w_dff_B_2IYgpU4x5_0),.dout(w_dff_B_YfZSMbct1_0),.clk(gclk));
	jdff dff_B_tJuO6fUj4_0(.din(w_dff_B_YfZSMbct1_0),.dout(w_dff_B_tJuO6fUj4_0),.clk(gclk));
	jdff dff_B_4fDFzSel4_0(.din(w_dff_B_tJuO6fUj4_0),.dout(w_dff_B_4fDFzSel4_0),.clk(gclk));
	jdff dff_B_OcSOR1jH6_0(.din(w_dff_B_4fDFzSel4_0),.dout(w_dff_B_OcSOR1jH6_0),.clk(gclk));
	jdff dff_B_ybIv3Zc71_0(.din(w_dff_B_OcSOR1jH6_0),.dout(w_dff_B_ybIv3Zc71_0),.clk(gclk));
	jdff dff_B_1BAhsGEk5_0(.din(w_dff_B_ybIv3Zc71_0),.dout(w_dff_B_1BAhsGEk5_0),.clk(gclk));
	jdff dff_B_aO7mvjEi6_0(.din(w_dff_B_1BAhsGEk5_0),.dout(w_dff_B_aO7mvjEi6_0),.clk(gclk));
	jdff dff_B_buV9XsNC1_0(.din(w_dff_B_aO7mvjEi6_0),.dout(w_dff_B_buV9XsNC1_0),.clk(gclk));
	jdff dff_B_KIVOnZwv2_0(.din(w_dff_B_buV9XsNC1_0),.dout(w_dff_B_KIVOnZwv2_0),.clk(gclk));
	jdff dff_B_6yGBRLHY8_0(.din(w_dff_B_KIVOnZwv2_0),.dout(w_dff_B_6yGBRLHY8_0),.clk(gclk));
	jdff dff_B_j58iVanm4_0(.din(w_dff_B_6yGBRLHY8_0),.dout(w_dff_B_j58iVanm4_0),.clk(gclk));
	jdff dff_B_Pot2UTII2_0(.din(w_dff_B_j58iVanm4_0),.dout(w_dff_B_Pot2UTII2_0),.clk(gclk));
	jdff dff_B_gbxrcPo36_0(.din(w_dff_B_Pot2UTII2_0),.dout(w_dff_B_gbxrcPo36_0),.clk(gclk));
	jdff dff_B_02TqhYHf2_0(.din(w_dff_B_gbxrcPo36_0),.dout(w_dff_B_02TqhYHf2_0),.clk(gclk));
	jdff dff_B_aqT3dCPg1_0(.din(w_dff_B_02TqhYHf2_0),.dout(w_dff_B_aqT3dCPg1_0),.clk(gclk));
	jdff dff_B_8cWEkuD12_0(.din(w_dff_B_aqT3dCPg1_0),.dout(w_dff_B_8cWEkuD12_0),.clk(gclk));
	jdff dff_B_71nkVB5p6_0(.din(w_dff_B_8cWEkuD12_0),.dout(w_dff_B_71nkVB5p6_0),.clk(gclk));
	jdff dff_B_KhVTjIfx9_0(.din(w_dff_B_71nkVB5p6_0),.dout(w_dff_B_KhVTjIfx9_0),.clk(gclk));
	jdff dff_B_vHLCZ4pF0_0(.din(w_dff_B_KhVTjIfx9_0),.dout(w_dff_B_vHLCZ4pF0_0),.clk(gclk));
	jdff dff_B_VBVqxeLI0_0(.din(w_dff_B_vHLCZ4pF0_0),.dout(w_dff_B_VBVqxeLI0_0),.clk(gclk));
	jdff dff_B_F4s63S5p8_0(.din(w_dff_B_VBVqxeLI0_0),.dout(w_dff_B_F4s63S5p8_0),.clk(gclk));
	jdff dff_B_CgB0dbMi4_0(.din(w_dff_B_F4s63S5p8_0),.dout(w_dff_B_CgB0dbMi4_0),.clk(gclk));
	jdff dff_B_NzYinipm2_0(.din(w_dff_B_CgB0dbMi4_0),.dout(w_dff_B_NzYinipm2_0),.clk(gclk));
	jdff dff_B_nw5wdooD7_0(.din(w_dff_B_NzYinipm2_0),.dout(w_dff_B_nw5wdooD7_0),.clk(gclk));
	jdff dff_B_Uqg6pbIw5_0(.din(w_dff_B_nw5wdooD7_0),.dout(w_dff_B_Uqg6pbIw5_0),.clk(gclk));
	jdff dff_B_MiHvLnEP0_0(.din(w_dff_B_Uqg6pbIw5_0),.dout(w_dff_B_MiHvLnEP0_0),.clk(gclk));
	jdff dff_B_FUf4G8331_0(.din(w_dff_B_MiHvLnEP0_0),.dout(w_dff_B_FUf4G8331_0),.clk(gclk));
	jdff dff_B_iwmOFbya2_0(.din(w_dff_B_FUf4G8331_0),.dout(w_dff_B_iwmOFbya2_0),.clk(gclk));
	jdff dff_B_EjbaOgTM5_0(.din(w_dff_B_iwmOFbya2_0),.dout(w_dff_B_EjbaOgTM5_0),.clk(gclk));
	jdff dff_B_qasx58sI4_0(.din(w_dff_B_EjbaOgTM5_0),.dout(w_dff_B_qasx58sI4_0),.clk(gclk));
	jdff dff_B_PTt5yt1J9_0(.din(w_dff_B_qasx58sI4_0),.dout(w_dff_B_PTt5yt1J9_0),.clk(gclk));
	jdff dff_B_Na910Bfd1_0(.din(w_dff_B_PTt5yt1J9_0),.dout(w_dff_B_Na910Bfd1_0),.clk(gclk));
	jdff dff_B_VfwFG6rv0_0(.din(w_dff_B_Na910Bfd1_0),.dout(w_dff_B_VfwFG6rv0_0),.clk(gclk));
	jdff dff_B_araAvJEA9_0(.din(w_dff_B_VfwFG6rv0_0),.dout(w_dff_B_araAvJEA9_0),.clk(gclk));
	jdff dff_B_8SlINF8p7_0(.din(w_dff_B_araAvJEA9_0),.dout(w_dff_B_8SlINF8p7_0),.clk(gclk));
	jdff dff_B_4u3RNrBc6_0(.din(w_dff_B_8SlINF8p7_0),.dout(w_dff_B_4u3RNrBc6_0),.clk(gclk));
	jdff dff_B_Fn2T9zcL1_0(.din(w_dff_B_4u3RNrBc6_0),.dout(w_dff_B_Fn2T9zcL1_0),.clk(gclk));
	jdff dff_B_HW9stFUS1_0(.din(w_dff_B_Fn2T9zcL1_0),.dout(w_dff_B_HW9stFUS1_0),.clk(gclk));
	jdff dff_B_a6v2rfvp2_0(.din(w_dff_B_HW9stFUS1_0),.dout(w_dff_B_a6v2rfvp2_0),.clk(gclk));
	jdff dff_B_sJNIWidZ7_0(.din(w_dff_B_a6v2rfvp2_0),.dout(w_dff_B_sJNIWidZ7_0),.clk(gclk));
	jdff dff_B_yqVr2DNA1_0(.din(w_dff_B_sJNIWidZ7_0),.dout(w_dff_B_yqVr2DNA1_0),.clk(gclk));
	jdff dff_B_ckxNXAPc9_0(.din(w_dff_B_yqVr2DNA1_0),.dout(w_dff_B_ckxNXAPc9_0),.clk(gclk));
	jdff dff_B_GnCUwiQs6_0(.din(w_dff_B_ckxNXAPc9_0),.dout(w_dff_B_GnCUwiQs6_0),.clk(gclk));
	jdff dff_B_TDWLEqX25_0(.din(w_dff_B_GnCUwiQs6_0),.dout(w_dff_B_TDWLEqX25_0),.clk(gclk));
	jdff dff_B_RMrYRhzl6_0(.din(w_dff_B_TDWLEqX25_0),.dout(w_dff_B_RMrYRhzl6_0),.clk(gclk));
	jdff dff_B_IVWHdDRC6_0(.din(w_dff_B_RMrYRhzl6_0),.dout(w_dff_B_IVWHdDRC6_0),.clk(gclk));
	jdff dff_B_1cZnVxff6_0(.din(w_dff_B_IVWHdDRC6_0),.dout(w_dff_B_1cZnVxff6_0),.clk(gclk));
	jdff dff_B_fQ0SBGcg6_0(.din(w_dff_B_1cZnVxff6_0),.dout(w_dff_B_fQ0SBGcg6_0),.clk(gclk));
	jdff dff_B_vtqh0Ppx6_0(.din(w_dff_B_fQ0SBGcg6_0),.dout(w_dff_B_vtqh0Ppx6_0),.clk(gclk));
	jdff dff_B_CNSv9hMK0_0(.din(w_dff_B_vtqh0Ppx6_0),.dout(w_dff_B_CNSv9hMK0_0),.clk(gclk));
	jdff dff_B_e2ljy7uB0_0(.din(w_dff_B_CNSv9hMK0_0),.dout(w_dff_B_e2ljy7uB0_0),.clk(gclk));
	jdff dff_B_xwfdHKxM6_0(.din(w_dff_B_e2ljy7uB0_0),.dout(w_dff_B_xwfdHKxM6_0),.clk(gclk));
	jdff dff_B_YljmDFe52_0(.din(w_dff_B_xwfdHKxM6_0),.dout(w_dff_B_YljmDFe52_0),.clk(gclk));
	jdff dff_B_BqZk7xP18_0(.din(w_dff_B_YljmDFe52_0),.dout(w_dff_B_BqZk7xP18_0),.clk(gclk));
	jdff dff_B_Ox9dIUWk2_0(.din(w_dff_B_BqZk7xP18_0),.dout(w_dff_B_Ox9dIUWk2_0),.clk(gclk));
	jdff dff_B_diLv3GE92_0(.din(w_dff_B_Ox9dIUWk2_0),.dout(w_dff_B_diLv3GE92_0),.clk(gclk));
	jdff dff_B_jwYYhK3T4_0(.din(w_dff_B_diLv3GE92_0),.dout(w_dff_B_jwYYhK3T4_0),.clk(gclk));
	jdff dff_B_JOmqquYs5_0(.din(w_dff_B_jwYYhK3T4_0),.dout(w_dff_B_JOmqquYs5_0),.clk(gclk));
	jdff dff_B_fTNL12B76_0(.din(w_dff_B_JOmqquYs5_0),.dout(w_dff_B_fTNL12B76_0),.clk(gclk));
	jdff dff_B_YfaYofbG5_0(.din(w_dff_B_fTNL12B76_0),.dout(w_dff_B_YfaYofbG5_0),.clk(gclk));
	jdff dff_B_iiL6A9U45_0(.din(w_dff_B_YfaYofbG5_0),.dout(w_dff_B_iiL6A9U45_0),.clk(gclk));
	jdff dff_B_6fqUfEJI2_0(.din(n1024),.dout(w_dff_B_6fqUfEJI2_0),.clk(gclk));
	jdff dff_B_A1vohAOT1_0(.din(w_dff_B_6fqUfEJI2_0),.dout(w_dff_B_A1vohAOT1_0),.clk(gclk));
	jdff dff_B_mX6zUOKX6_0(.din(w_dff_B_A1vohAOT1_0),.dout(w_dff_B_mX6zUOKX6_0),.clk(gclk));
	jdff dff_B_h1C0nFZh6_0(.din(w_dff_B_mX6zUOKX6_0),.dout(w_dff_B_h1C0nFZh6_0),.clk(gclk));
	jdff dff_B_gBJF0tbC8_0(.din(w_dff_B_h1C0nFZh6_0),.dout(w_dff_B_gBJF0tbC8_0),.clk(gclk));
	jdff dff_B_1NOccfLd7_0(.din(w_dff_B_gBJF0tbC8_0),.dout(w_dff_B_1NOccfLd7_0),.clk(gclk));
	jdff dff_B_tUimDyCa2_0(.din(w_dff_B_1NOccfLd7_0),.dout(w_dff_B_tUimDyCa2_0),.clk(gclk));
	jdff dff_B_OMh5HBhk3_0(.din(w_dff_B_tUimDyCa2_0),.dout(w_dff_B_OMh5HBhk3_0),.clk(gclk));
	jdff dff_B_7ANrYdw48_0(.din(w_dff_B_OMh5HBhk3_0),.dout(w_dff_B_7ANrYdw48_0),.clk(gclk));
	jdff dff_B_ZYkWAQb59_0(.din(w_dff_B_7ANrYdw48_0),.dout(w_dff_B_ZYkWAQb59_0),.clk(gclk));
	jdff dff_B_ay4qsUHV1_0(.din(w_dff_B_ZYkWAQb59_0),.dout(w_dff_B_ay4qsUHV1_0),.clk(gclk));
	jdff dff_B_nGVVSN2v8_0(.din(w_dff_B_ay4qsUHV1_0),.dout(w_dff_B_nGVVSN2v8_0),.clk(gclk));
	jdff dff_B_YYwv4BJ15_0(.din(w_dff_B_nGVVSN2v8_0),.dout(w_dff_B_YYwv4BJ15_0),.clk(gclk));
	jdff dff_B_bO379u7c7_0(.din(w_dff_B_YYwv4BJ15_0),.dout(w_dff_B_bO379u7c7_0),.clk(gclk));
	jdff dff_B_Y7VsG9id8_0(.din(w_dff_B_bO379u7c7_0),.dout(w_dff_B_Y7VsG9id8_0),.clk(gclk));
	jdff dff_B_63KiuyzB9_0(.din(w_dff_B_Y7VsG9id8_0),.dout(w_dff_B_63KiuyzB9_0),.clk(gclk));
	jdff dff_B_M3eWBkSk1_0(.din(w_dff_B_63KiuyzB9_0),.dout(w_dff_B_M3eWBkSk1_0),.clk(gclk));
	jdff dff_B_qNnEAjzs4_0(.din(w_dff_B_M3eWBkSk1_0),.dout(w_dff_B_qNnEAjzs4_0),.clk(gclk));
	jdff dff_B_zT7O8DQ47_0(.din(w_dff_B_qNnEAjzs4_0),.dout(w_dff_B_zT7O8DQ47_0),.clk(gclk));
	jdff dff_B_6NlwGPmf9_0(.din(w_dff_B_zT7O8DQ47_0),.dout(w_dff_B_6NlwGPmf9_0),.clk(gclk));
	jdff dff_B_UYLTsiUC7_0(.din(w_dff_B_6NlwGPmf9_0),.dout(w_dff_B_UYLTsiUC7_0),.clk(gclk));
	jdff dff_B_kWONCJSn0_0(.din(w_dff_B_UYLTsiUC7_0),.dout(w_dff_B_kWONCJSn0_0),.clk(gclk));
	jdff dff_B_MS6IPvQu3_0(.din(w_dff_B_kWONCJSn0_0),.dout(w_dff_B_MS6IPvQu3_0),.clk(gclk));
	jdff dff_B_TTOrtpJ42_0(.din(w_dff_B_MS6IPvQu3_0),.dout(w_dff_B_TTOrtpJ42_0),.clk(gclk));
	jdff dff_B_epvi4E0Y5_0(.din(w_dff_B_TTOrtpJ42_0),.dout(w_dff_B_epvi4E0Y5_0),.clk(gclk));
	jdff dff_B_jHtEUOk53_0(.din(w_dff_B_epvi4E0Y5_0),.dout(w_dff_B_jHtEUOk53_0),.clk(gclk));
	jdff dff_B_Z7NnmeeY3_0(.din(w_dff_B_jHtEUOk53_0),.dout(w_dff_B_Z7NnmeeY3_0),.clk(gclk));
	jdff dff_B_c3F1Tnwz8_0(.din(w_dff_B_Z7NnmeeY3_0),.dout(w_dff_B_c3F1Tnwz8_0),.clk(gclk));
	jdff dff_B_O2CgCM2y4_0(.din(w_dff_B_c3F1Tnwz8_0),.dout(w_dff_B_O2CgCM2y4_0),.clk(gclk));
	jdff dff_B_YueCyedn2_0(.din(w_dff_B_O2CgCM2y4_0),.dout(w_dff_B_YueCyedn2_0),.clk(gclk));
	jdff dff_B_XIit2uNM3_0(.din(w_dff_B_YueCyedn2_0),.dout(w_dff_B_XIit2uNM3_0),.clk(gclk));
	jdff dff_B_FIH0O3PE7_0(.din(w_dff_B_XIit2uNM3_0),.dout(w_dff_B_FIH0O3PE7_0),.clk(gclk));
	jdff dff_B_9QwMtVZH7_0(.din(w_dff_B_FIH0O3PE7_0),.dout(w_dff_B_9QwMtVZH7_0),.clk(gclk));
	jdff dff_B_iGBc7U835_0(.din(w_dff_B_9QwMtVZH7_0),.dout(w_dff_B_iGBc7U835_0),.clk(gclk));
	jdff dff_B_zOBFKmIG1_0(.din(w_dff_B_iGBc7U835_0),.dout(w_dff_B_zOBFKmIG1_0),.clk(gclk));
	jdff dff_B_Gv7OQc6a9_0(.din(w_dff_B_zOBFKmIG1_0),.dout(w_dff_B_Gv7OQc6a9_0),.clk(gclk));
	jdff dff_B_w0ObPVLr6_0(.din(w_dff_B_Gv7OQc6a9_0),.dout(w_dff_B_w0ObPVLr6_0),.clk(gclk));
	jdff dff_B_wB3P3ZDn1_0(.din(w_dff_B_w0ObPVLr6_0),.dout(w_dff_B_wB3P3ZDn1_0),.clk(gclk));
	jdff dff_B_QoK31wgl6_0(.din(w_dff_B_wB3P3ZDn1_0),.dout(w_dff_B_QoK31wgl6_0),.clk(gclk));
	jdff dff_B_hDGfCOUa7_0(.din(w_dff_B_QoK31wgl6_0),.dout(w_dff_B_hDGfCOUa7_0),.clk(gclk));
	jdff dff_B_rbEKOed13_0(.din(w_dff_B_hDGfCOUa7_0),.dout(w_dff_B_rbEKOed13_0),.clk(gclk));
	jdff dff_B_9w62NqoI9_0(.din(w_dff_B_rbEKOed13_0),.dout(w_dff_B_9w62NqoI9_0),.clk(gclk));
	jdff dff_B_lQ7h7CId1_0(.din(w_dff_B_9w62NqoI9_0),.dout(w_dff_B_lQ7h7CId1_0),.clk(gclk));
	jdff dff_B_q7eixNu19_0(.din(w_dff_B_lQ7h7CId1_0),.dout(w_dff_B_q7eixNu19_0),.clk(gclk));
	jdff dff_B_aVtERWWg4_0(.din(w_dff_B_q7eixNu19_0),.dout(w_dff_B_aVtERWWg4_0),.clk(gclk));
	jdff dff_B_BYV83VVI8_0(.din(w_dff_B_aVtERWWg4_0),.dout(w_dff_B_BYV83VVI8_0),.clk(gclk));
	jdff dff_B_NVMMmkC14_0(.din(w_dff_B_BYV83VVI8_0),.dout(w_dff_B_NVMMmkC14_0),.clk(gclk));
	jdff dff_B_42vFMTZd7_0(.din(w_dff_B_NVMMmkC14_0),.dout(w_dff_B_42vFMTZd7_0),.clk(gclk));
	jdff dff_B_oJnJh0Uw9_0(.din(w_dff_B_42vFMTZd7_0),.dout(w_dff_B_oJnJh0Uw9_0),.clk(gclk));
	jdff dff_B_9B4L9QN64_0(.din(w_dff_B_oJnJh0Uw9_0),.dout(w_dff_B_9B4L9QN64_0),.clk(gclk));
	jdff dff_B_8vhDov6l6_0(.din(w_dff_B_9B4L9QN64_0),.dout(w_dff_B_8vhDov6l6_0),.clk(gclk));
	jdff dff_B_eAj6qN8B3_0(.din(w_dff_B_8vhDov6l6_0),.dout(w_dff_B_eAj6qN8B3_0),.clk(gclk));
	jdff dff_B_e84rrwvS3_0(.din(w_dff_B_eAj6qN8B3_0),.dout(w_dff_B_e84rrwvS3_0),.clk(gclk));
	jdff dff_B_Q1KJMv9w1_0(.din(w_dff_B_e84rrwvS3_0),.dout(w_dff_B_Q1KJMv9w1_0),.clk(gclk));
	jdff dff_B_JfafIsUy1_0(.din(w_dff_B_Q1KJMv9w1_0),.dout(w_dff_B_JfafIsUy1_0),.clk(gclk));
	jdff dff_B_kevNxul21_0(.din(w_dff_B_JfafIsUy1_0),.dout(w_dff_B_kevNxul21_0),.clk(gclk));
	jdff dff_B_XYjokHdl6_0(.din(w_dff_B_kevNxul21_0),.dout(w_dff_B_XYjokHdl6_0),.clk(gclk));
	jdff dff_B_7U2tDgcl9_0(.din(w_dff_B_XYjokHdl6_0),.dout(w_dff_B_7U2tDgcl9_0),.clk(gclk));
	jdff dff_B_ZKGdyJ900_0(.din(w_dff_B_7U2tDgcl9_0),.dout(w_dff_B_ZKGdyJ900_0),.clk(gclk));
	jdff dff_B_U6u55A9L6_0(.din(w_dff_B_ZKGdyJ900_0),.dout(w_dff_B_U6u55A9L6_0),.clk(gclk));
	jdff dff_B_uaMqcePb5_0(.din(w_dff_B_U6u55A9L6_0),.dout(w_dff_B_uaMqcePb5_0),.clk(gclk));
	jdff dff_B_6UHE639p7_0(.din(w_dff_B_uaMqcePb5_0),.dout(w_dff_B_6UHE639p7_0),.clk(gclk));
	jdff dff_B_HPdYf0aL0_0(.din(w_dff_B_6UHE639p7_0),.dout(w_dff_B_HPdYf0aL0_0),.clk(gclk));
	jdff dff_B_RSD11qq79_0(.din(w_dff_B_HPdYf0aL0_0),.dout(w_dff_B_RSD11qq79_0),.clk(gclk));
	jdff dff_B_H7RRcInR7_0(.din(w_dff_B_RSD11qq79_0),.dout(w_dff_B_H7RRcInR7_0),.clk(gclk));
	jdff dff_B_PE1dnht06_0(.din(w_dff_B_H7RRcInR7_0),.dout(w_dff_B_PE1dnht06_0),.clk(gclk));
	jdff dff_B_CZNzxYcS2_0(.din(w_dff_B_PE1dnht06_0),.dout(w_dff_B_CZNzxYcS2_0),.clk(gclk));
	jdff dff_B_Rdfaso0W9_0(.din(w_dff_B_CZNzxYcS2_0),.dout(w_dff_B_Rdfaso0W9_0),.clk(gclk));
	jdff dff_B_DLKGojIZ2_0(.din(w_dff_B_Rdfaso0W9_0),.dout(w_dff_B_DLKGojIZ2_0),.clk(gclk));
	jdff dff_B_jSkpze7G8_0(.din(w_dff_B_DLKGojIZ2_0),.dout(w_dff_B_jSkpze7G8_0),.clk(gclk));
	jdff dff_B_oPKN4p3d5_0(.din(w_dff_B_jSkpze7G8_0),.dout(w_dff_B_oPKN4p3d5_0),.clk(gclk));
	jdff dff_B_trvscKgr9_0(.din(w_dff_B_oPKN4p3d5_0),.dout(w_dff_B_trvscKgr9_0),.clk(gclk));
	jdff dff_B_TA6RxhDI3_0(.din(w_dff_B_trvscKgr9_0),.dout(w_dff_B_TA6RxhDI3_0),.clk(gclk));
	jdff dff_B_T0eBvAu56_0(.din(w_dff_B_TA6RxhDI3_0),.dout(w_dff_B_T0eBvAu56_0),.clk(gclk));
	jdff dff_B_jQFfflpp8_0(.din(w_dff_B_T0eBvAu56_0),.dout(w_dff_B_jQFfflpp8_0),.clk(gclk));
	jdff dff_B_QLtcTgWz4_0(.din(w_dff_B_jQFfflpp8_0),.dout(w_dff_B_QLtcTgWz4_0),.clk(gclk));
	jdff dff_B_SVOxw2tu7_0(.din(w_dff_B_QLtcTgWz4_0),.dout(w_dff_B_SVOxw2tu7_0),.clk(gclk));
	jdff dff_B_vvg8Ulfn5_0(.din(w_dff_B_SVOxw2tu7_0),.dout(w_dff_B_vvg8Ulfn5_0),.clk(gclk));
	jdff dff_B_Gm9NC6fF6_0(.din(w_dff_B_vvg8Ulfn5_0),.dout(w_dff_B_Gm9NC6fF6_0),.clk(gclk));
	jdff dff_B_qpx5BBst8_0(.din(w_dff_B_Gm9NC6fF6_0),.dout(w_dff_B_qpx5BBst8_0),.clk(gclk));
	jdff dff_B_xQHFDjek1_0(.din(w_dff_B_qpx5BBst8_0),.dout(w_dff_B_xQHFDjek1_0),.clk(gclk));
	jdff dff_B_1VKNp4vS6_0(.din(w_dff_B_xQHFDjek1_0),.dout(w_dff_B_1VKNp4vS6_0),.clk(gclk));
	jdff dff_B_6cTdRamm7_0(.din(w_dff_B_1VKNp4vS6_0),.dout(w_dff_B_6cTdRamm7_0),.clk(gclk));
	jdff dff_B_Wjjk8S1x1_0(.din(w_dff_B_6cTdRamm7_0),.dout(w_dff_B_Wjjk8S1x1_0),.clk(gclk));
	jdff dff_B_9vcuXYfz0_0(.din(w_dff_B_Wjjk8S1x1_0),.dout(w_dff_B_9vcuXYfz0_0),.clk(gclk));
	jdff dff_B_Z57goe1K3_0(.din(w_dff_B_9vcuXYfz0_0),.dout(w_dff_B_Z57goe1K3_0),.clk(gclk));
	jdff dff_B_XBATHLZS6_0(.din(w_dff_B_Z57goe1K3_0),.dout(w_dff_B_XBATHLZS6_0),.clk(gclk));
	jdff dff_B_0IwsHbfy0_0(.din(w_dff_B_XBATHLZS6_0),.dout(w_dff_B_0IwsHbfy0_0),.clk(gclk));
	jdff dff_B_udcVLTQG1_0(.din(w_dff_B_0IwsHbfy0_0),.dout(w_dff_B_udcVLTQG1_0),.clk(gclk));
	jdff dff_B_67W1r02d3_0(.din(w_dff_B_udcVLTQG1_0),.dout(w_dff_B_67W1r02d3_0),.clk(gclk));
	jdff dff_B_VjDlzsGQ4_0(.din(w_dff_B_67W1r02d3_0),.dout(w_dff_B_VjDlzsGQ4_0),.clk(gclk));
	jdff dff_B_jVm8dfvb6_0(.din(w_dff_B_VjDlzsGQ4_0),.dout(w_dff_B_jVm8dfvb6_0),.clk(gclk));
	jdff dff_B_On0BB9t34_0(.din(w_dff_B_jVm8dfvb6_0),.dout(w_dff_B_On0BB9t34_0),.clk(gclk));
	jdff dff_B_plYGxNwq3_0(.din(w_dff_B_On0BB9t34_0),.dout(w_dff_B_plYGxNwq3_0),.clk(gclk));
	jdff dff_B_cDzvERom3_0(.din(w_dff_B_plYGxNwq3_0),.dout(w_dff_B_cDzvERom3_0),.clk(gclk));
	jdff dff_B_gUGUsPZu9_0(.din(w_dff_B_cDzvERom3_0),.dout(w_dff_B_gUGUsPZu9_0),.clk(gclk));
	jdff dff_B_ztDlVhTp2_0(.din(w_dff_B_gUGUsPZu9_0),.dout(w_dff_B_ztDlVhTp2_0),.clk(gclk));
	jdff dff_B_tYqDB4EN6_0(.din(w_dff_B_ztDlVhTp2_0),.dout(w_dff_B_tYqDB4EN6_0),.clk(gclk));
	jdff dff_B_3Iw6unZh7_0(.din(w_dff_B_tYqDB4EN6_0),.dout(w_dff_B_3Iw6unZh7_0),.clk(gclk));
	jdff dff_B_HqxgmXPU3_0(.din(w_dff_B_3Iw6unZh7_0),.dout(w_dff_B_HqxgmXPU3_0),.clk(gclk));
	jdff dff_B_P7HVCpYw4_0(.din(w_dff_B_HqxgmXPU3_0),.dout(w_dff_B_P7HVCpYw4_0),.clk(gclk));
	jdff dff_B_JdbqUIM05_0(.din(w_dff_B_P7HVCpYw4_0),.dout(w_dff_B_JdbqUIM05_0),.clk(gclk));
	jdff dff_B_uoTaioss2_0(.din(w_dff_B_JdbqUIM05_0),.dout(w_dff_B_uoTaioss2_0),.clk(gclk));
	jdff dff_B_xDWWmLjZ9_0(.din(w_dff_B_uoTaioss2_0),.dout(w_dff_B_xDWWmLjZ9_0),.clk(gclk));
	jdff dff_B_G5EJpep07_0(.din(w_dff_B_xDWWmLjZ9_0),.dout(w_dff_B_G5EJpep07_0),.clk(gclk));
	jdff dff_B_T2YmP8GL7_0(.din(w_dff_B_G5EJpep07_0),.dout(w_dff_B_T2YmP8GL7_0),.clk(gclk));
	jdff dff_B_nklgWzpH4_0(.din(n1030),.dout(w_dff_B_nklgWzpH4_0),.clk(gclk));
	jdff dff_B_ZXZWAm6g6_0(.din(w_dff_B_nklgWzpH4_0),.dout(w_dff_B_ZXZWAm6g6_0),.clk(gclk));
	jdff dff_B_eoEoJo673_0(.din(w_dff_B_ZXZWAm6g6_0),.dout(w_dff_B_eoEoJo673_0),.clk(gclk));
	jdff dff_B_h222w6BG3_0(.din(w_dff_B_eoEoJo673_0),.dout(w_dff_B_h222w6BG3_0),.clk(gclk));
	jdff dff_B_hdWqmTW64_0(.din(w_dff_B_h222w6BG3_0),.dout(w_dff_B_hdWqmTW64_0),.clk(gclk));
	jdff dff_B_Ysh7bVVO8_0(.din(w_dff_B_hdWqmTW64_0),.dout(w_dff_B_Ysh7bVVO8_0),.clk(gclk));
	jdff dff_B_Y1clmQ7b1_0(.din(w_dff_B_Ysh7bVVO8_0),.dout(w_dff_B_Y1clmQ7b1_0),.clk(gclk));
	jdff dff_B_ZeTPjXIe8_0(.din(w_dff_B_Y1clmQ7b1_0),.dout(w_dff_B_ZeTPjXIe8_0),.clk(gclk));
	jdff dff_B_QZq85zmY8_0(.din(w_dff_B_ZeTPjXIe8_0),.dout(w_dff_B_QZq85zmY8_0),.clk(gclk));
	jdff dff_B_XGWhxQsZ8_0(.din(w_dff_B_QZq85zmY8_0),.dout(w_dff_B_XGWhxQsZ8_0),.clk(gclk));
	jdff dff_B_IuCCrDRT4_0(.din(w_dff_B_XGWhxQsZ8_0),.dout(w_dff_B_IuCCrDRT4_0),.clk(gclk));
	jdff dff_B_0fR7u6Ys5_0(.din(w_dff_B_IuCCrDRT4_0),.dout(w_dff_B_0fR7u6Ys5_0),.clk(gclk));
	jdff dff_B_Uwelh4V23_0(.din(w_dff_B_0fR7u6Ys5_0),.dout(w_dff_B_Uwelh4V23_0),.clk(gclk));
	jdff dff_B_VLEBRs3r6_0(.din(w_dff_B_Uwelh4V23_0),.dout(w_dff_B_VLEBRs3r6_0),.clk(gclk));
	jdff dff_B_rQHQqHXQ8_0(.din(w_dff_B_VLEBRs3r6_0),.dout(w_dff_B_rQHQqHXQ8_0),.clk(gclk));
	jdff dff_B_ODsOWPSp4_0(.din(w_dff_B_rQHQqHXQ8_0),.dout(w_dff_B_ODsOWPSp4_0),.clk(gclk));
	jdff dff_B_3CI9vcSz1_0(.din(w_dff_B_ODsOWPSp4_0),.dout(w_dff_B_3CI9vcSz1_0),.clk(gclk));
	jdff dff_B_HvbPgBVb0_0(.din(w_dff_B_3CI9vcSz1_0),.dout(w_dff_B_HvbPgBVb0_0),.clk(gclk));
	jdff dff_B_DeuWbQdY2_0(.din(w_dff_B_HvbPgBVb0_0),.dout(w_dff_B_DeuWbQdY2_0),.clk(gclk));
	jdff dff_B_jpdZv3Q25_0(.din(w_dff_B_DeuWbQdY2_0),.dout(w_dff_B_jpdZv3Q25_0),.clk(gclk));
	jdff dff_B_8t2ohWji8_0(.din(w_dff_B_jpdZv3Q25_0),.dout(w_dff_B_8t2ohWji8_0),.clk(gclk));
	jdff dff_B_w6YHkdCv7_0(.din(w_dff_B_8t2ohWji8_0),.dout(w_dff_B_w6YHkdCv7_0),.clk(gclk));
	jdff dff_B_HtldMgdf0_0(.din(w_dff_B_w6YHkdCv7_0),.dout(w_dff_B_HtldMgdf0_0),.clk(gclk));
	jdff dff_B_xpuZ1OLr7_0(.din(w_dff_B_HtldMgdf0_0),.dout(w_dff_B_xpuZ1OLr7_0),.clk(gclk));
	jdff dff_B_PrRvLsxZ6_0(.din(w_dff_B_xpuZ1OLr7_0),.dout(w_dff_B_PrRvLsxZ6_0),.clk(gclk));
	jdff dff_B_gySG7fem7_0(.din(w_dff_B_PrRvLsxZ6_0),.dout(w_dff_B_gySG7fem7_0),.clk(gclk));
	jdff dff_B_IETOyFW67_0(.din(w_dff_B_gySG7fem7_0),.dout(w_dff_B_IETOyFW67_0),.clk(gclk));
	jdff dff_B_sEJhzPr62_0(.din(w_dff_B_IETOyFW67_0),.dout(w_dff_B_sEJhzPr62_0),.clk(gclk));
	jdff dff_B_nOL90Hyt4_0(.din(w_dff_B_sEJhzPr62_0),.dout(w_dff_B_nOL90Hyt4_0),.clk(gclk));
	jdff dff_B_2DN8uHtl7_0(.din(w_dff_B_nOL90Hyt4_0),.dout(w_dff_B_2DN8uHtl7_0),.clk(gclk));
	jdff dff_B_Pvyl37zS4_0(.din(w_dff_B_2DN8uHtl7_0),.dout(w_dff_B_Pvyl37zS4_0),.clk(gclk));
	jdff dff_B_jvhB9CbW7_0(.din(w_dff_B_Pvyl37zS4_0),.dout(w_dff_B_jvhB9CbW7_0),.clk(gclk));
	jdff dff_B_wSYc1CNi4_0(.din(w_dff_B_jvhB9CbW7_0),.dout(w_dff_B_wSYc1CNi4_0),.clk(gclk));
	jdff dff_B_Q3ek2Oyw4_0(.din(w_dff_B_wSYc1CNi4_0),.dout(w_dff_B_Q3ek2Oyw4_0),.clk(gclk));
	jdff dff_B_F4JkyPU58_0(.din(w_dff_B_Q3ek2Oyw4_0),.dout(w_dff_B_F4JkyPU58_0),.clk(gclk));
	jdff dff_B_SieVe3Ol3_0(.din(w_dff_B_F4JkyPU58_0),.dout(w_dff_B_SieVe3Ol3_0),.clk(gclk));
	jdff dff_B_PpvYVAPT6_0(.din(w_dff_B_SieVe3Ol3_0),.dout(w_dff_B_PpvYVAPT6_0),.clk(gclk));
	jdff dff_B_EIeNnAz38_0(.din(w_dff_B_PpvYVAPT6_0),.dout(w_dff_B_EIeNnAz38_0),.clk(gclk));
	jdff dff_B_tmuq0qS35_0(.din(w_dff_B_EIeNnAz38_0),.dout(w_dff_B_tmuq0qS35_0),.clk(gclk));
	jdff dff_B_KdnVXJbt6_0(.din(w_dff_B_tmuq0qS35_0),.dout(w_dff_B_KdnVXJbt6_0),.clk(gclk));
	jdff dff_B_Rv8hatbY5_0(.din(w_dff_B_KdnVXJbt6_0),.dout(w_dff_B_Rv8hatbY5_0),.clk(gclk));
	jdff dff_B_ZI6fjHmS7_0(.din(w_dff_B_Rv8hatbY5_0),.dout(w_dff_B_ZI6fjHmS7_0),.clk(gclk));
	jdff dff_B_Ov2dgGlC1_0(.din(w_dff_B_ZI6fjHmS7_0),.dout(w_dff_B_Ov2dgGlC1_0),.clk(gclk));
	jdff dff_B_zleW9DY09_0(.din(w_dff_B_Ov2dgGlC1_0),.dout(w_dff_B_zleW9DY09_0),.clk(gclk));
	jdff dff_B_o0Tnxdyx7_0(.din(w_dff_B_zleW9DY09_0),.dout(w_dff_B_o0Tnxdyx7_0),.clk(gclk));
	jdff dff_B_qJtkcBIK4_0(.din(w_dff_B_o0Tnxdyx7_0),.dout(w_dff_B_qJtkcBIK4_0),.clk(gclk));
	jdff dff_B_19YzJv9I1_0(.din(w_dff_B_qJtkcBIK4_0),.dout(w_dff_B_19YzJv9I1_0),.clk(gclk));
	jdff dff_B_XiworvY53_0(.din(w_dff_B_19YzJv9I1_0),.dout(w_dff_B_XiworvY53_0),.clk(gclk));
	jdff dff_B_6MPsd7W32_0(.din(w_dff_B_XiworvY53_0),.dout(w_dff_B_6MPsd7W32_0),.clk(gclk));
	jdff dff_B_yaiIkwHR2_0(.din(w_dff_B_6MPsd7W32_0),.dout(w_dff_B_yaiIkwHR2_0),.clk(gclk));
	jdff dff_B_2s1cPYZF4_0(.din(w_dff_B_yaiIkwHR2_0),.dout(w_dff_B_2s1cPYZF4_0),.clk(gclk));
	jdff dff_B_93uEfT1T0_0(.din(w_dff_B_2s1cPYZF4_0),.dout(w_dff_B_93uEfT1T0_0),.clk(gclk));
	jdff dff_B_JZXIks4y6_0(.din(w_dff_B_93uEfT1T0_0),.dout(w_dff_B_JZXIks4y6_0),.clk(gclk));
	jdff dff_B_71haXrJZ1_0(.din(w_dff_B_JZXIks4y6_0),.dout(w_dff_B_71haXrJZ1_0),.clk(gclk));
	jdff dff_B_srYQ604o0_0(.din(w_dff_B_71haXrJZ1_0),.dout(w_dff_B_srYQ604o0_0),.clk(gclk));
	jdff dff_B_tvxMLiiL9_0(.din(w_dff_B_srYQ604o0_0),.dout(w_dff_B_tvxMLiiL9_0),.clk(gclk));
	jdff dff_B_LSWn1x8e5_0(.din(w_dff_B_tvxMLiiL9_0),.dout(w_dff_B_LSWn1x8e5_0),.clk(gclk));
	jdff dff_B_hXgbemVz2_0(.din(w_dff_B_LSWn1x8e5_0),.dout(w_dff_B_hXgbemVz2_0),.clk(gclk));
	jdff dff_B_bgpFdUFS2_0(.din(w_dff_B_hXgbemVz2_0),.dout(w_dff_B_bgpFdUFS2_0),.clk(gclk));
	jdff dff_B_X4EZn1M13_0(.din(w_dff_B_bgpFdUFS2_0),.dout(w_dff_B_X4EZn1M13_0),.clk(gclk));
	jdff dff_B_eyySQIqE6_0(.din(w_dff_B_X4EZn1M13_0),.dout(w_dff_B_eyySQIqE6_0),.clk(gclk));
	jdff dff_B_JWtMNE7Q6_0(.din(w_dff_B_eyySQIqE6_0),.dout(w_dff_B_JWtMNE7Q6_0),.clk(gclk));
	jdff dff_B_2pVWTnaL9_0(.din(w_dff_B_JWtMNE7Q6_0),.dout(w_dff_B_2pVWTnaL9_0),.clk(gclk));
	jdff dff_B_0tIW24Sl2_0(.din(w_dff_B_2pVWTnaL9_0),.dout(w_dff_B_0tIW24Sl2_0),.clk(gclk));
	jdff dff_B_qmsSJ3yW5_0(.din(w_dff_B_0tIW24Sl2_0),.dout(w_dff_B_qmsSJ3yW5_0),.clk(gclk));
	jdff dff_B_0wvE8l2H8_0(.din(w_dff_B_qmsSJ3yW5_0),.dout(w_dff_B_0wvE8l2H8_0),.clk(gclk));
	jdff dff_B_QvXXgIOR5_0(.din(w_dff_B_0wvE8l2H8_0),.dout(w_dff_B_QvXXgIOR5_0),.clk(gclk));
	jdff dff_B_za769sNV7_0(.din(w_dff_B_QvXXgIOR5_0),.dout(w_dff_B_za769sNV7_0),.clk(gclk));
	jdff dff_B_HpMsnEni5_0(.din(w_dff_B_za769sNV7_0),.dout(w_dff_B_HpMsnEni5_0),.clk(gclk));
	jdff dff_B_uWMn5IYn4_0(.din(w_dff_B_HpMsnEni5_0),.dout(w_dff_B_uWMn5IYn4_0),.clk(gclk));
	jdff dff_B_DKyQyM5R7_0(.din(w_dff_B_uWMn5IYn4_0),.dout(w_dff_B_DKyQyM5R7_0),.clk(gclk));
	jdff dff_B_cl13aeGR4_0(.din(w_dff_B_DKyQyM5R7_0),.dout(w_dff_B_cl13aeGR4_0),.clk(gclk));
	jdff dff_B_Y5qPERVi0_0(.din(w_dff_B_cl13aeGR4_0),.dout(w_dff_B_Y5qPERVi0_0),.clk(gclk));
	jdff dff_B_AEjyVo2L5_0(.din(w_dff_B_Y5qPERVi0_0),.dout(w_dff_B_AEjyVo2L5_0),.clk(gclk));
	jdff dff_B_83bwYSdd1_0(.din(w_dff_B_AEjyVo2L5_0),.dout(w_dff_B_83bwYSdd1_0),.clk(gclk));
	jdff dff_B_oGYS17yU6_0(.din(w_dff_B_83bwYSdd1_0),.dout(w_dff_B_oGYS17yU6_0),.clk(gclk));
	jdff dff_B_o7cLntBr9_0(.din(w_dff_B_oGYS17yU6_0),.dout(w_dff_B_o7cLntBr9_0),.clk(gclk));
	jdff dff_B_nzpOFU7Q8_0(.din(w_dff_B_o7cLntBr9_0),.dout(w_dff_B_nzpOFU7Q8_0),.clk(gclk));
	jdff dff_B_kd2ksk6b2_0(.din(w_dff_B_nzpOFU7Q8_0),.dout(w_dff_B_kd2ksk6b2_0),.clk(gclk));
	jdff dff_B_4D1wTTfc6_0(.din(w_dff_B_kd2ksk6b2_0),.dout(w_dff_B_4D1wTTfc6_0),.clk(gclk));
	jdff dff_B_SfVIvRmZ1_0(.din(w_dff_B_4D1wTTfc6_0),.dout(w_dff_B_SfVIvRmZ1_0),.clk(gclk));
	jdff dff_B_5voHPdDr7_0(.din(w_dff_B_SfVIvRmZ1_0),.dout(w_dff_B_5voHPdDr7_0),.clk(gclk));
	jdff dff_B_968wELXU8_0(.din(w_dff_B_5voHPdDr7_0),.dout(w_dff_B_968wELXU8_0),.clk(gclk));
	jdff dff_B_lBy4Ms0D5_0(.din(w_dff_B_968wELXU8_0),.dout(w_dff_B_lBy4Ms0D5_0),.clk(gclk));
	jdff dff_B_xZski9ev2_0(.din(w_dff_B_lBy4Ms0D5_0),.dout(w_dff_B_xZski9ev2_0),.clk(gclk));
	jdff dff_B_bWWERdDD8_0(.din(w_dff_B_xZski9ev2_0),.dout(w_dff_B_bWWERdDD8_0),.clk(gclk));
	jdff dff_B_3wGUs2am8_0(.din(w_dff_B_bWWERdDD8_0),.dout(w_dff_B_3wGUs2am8_0),.clk(gclk));
	jdff dff_B_g2ZISok74_0(.din(w_dff_B_3wGUs2am8_0),.dout(w_dff_B_g2ZISok74_0),.clk(gclk));
	jdff dff_B_B7YvaD4A2_0(.din(w_dff_B_g2ZISok74_0),.dout(w_dff_B_B7YvaD4A2_0),.clk(gclk));
	jdff dff_B_2PViXef75_0(.din(w_dff_B_B7YvaD4A2_0),.dout(w_dff_B_2PViXef75_0),.clk(gclk));
	jdff dff_B_mEc9Ho3k7_0(.din(w_dff_B_2PViXef75_0),.dout(w_dff_B_mEc9Ho3k7_0),.clk(gclk));
	jdff dff_B_wgUGMa0p2_0(.din(w_dff_B_mEc9Ho3k7_0),.dout(w_dff_B_wgUGMa0p2_0),.clk(gclk));
	jdff dff_B_zAhRoE9u1_0(.din(w_dff_B_wgUGMa0p2_0),.dout(w_dff_B_zAhRoE9u1_0),.clk(gclk));
	jdff dff_B_zRVI6D4X9_0(.din(w_dff_B_zAhRoE9u1_0),.dout(w_dff_B_zRVI6D4X9_0),.clk(gclk));
	jdff dff_B_GYP6yAdF9_0(.din(w_dff_B_zRVI6D4X9_0),.dout(w_dff_B_GYP6yAdF9_0),.clk(gclk));
	jdff dff_B_ntjSw7dF6_0(.din(w_dff_B_GYP6yAdF9_0),.dout(w_dff_B_ntjSw7dF6_0),.clk(gclk));
	jdff dff_B_5Zwip4k81_0(.din(w_dff_B_ntjSw7dF6_0),.dout(w_dff_B_5Zwip4k81_0),.clk(gclk));
	jdff dff_B_jmDuG3Jx0_0(.din(w_dff_B_5Zwip4k81_0),.dout(w_dff_B_jmDuG3Jx0_0),.clk(gclk));
	jdff dff_B_DJXJUhZN3_0(.din(w_dff_B_jmDuG3Jx0_0),.dout(w_dff_B_DJXJUhZN3_0),.clk(gclk));
	jdff dff_B_GQHpvbFz1_0(.din(w_dff_B_DJXJUhZN3_0),.dout(w_dff_B_GQHpvbFz1_0),.clk(gclk));
	jdff dff_B_QHVEtMsV2_0(.din(w_dff_B_GQHpvbFz1_0),.dout(w_dff_B_QHVEtMsV2_0),.clk(gclk));
	jdff dff_B_ouP5JOAq0_0(.din(w_dff_B_QHVEtMsV2_0),.dout(w_dff_B_ouP5JOAq0_0),.clk(gclk));
	jdff dff_B_cqES8raJ6_0(.din(w_dff_B_ouP5JOAq0_0),.dout(w_dff_B_cqES8raJ6_0),.clk(gclk));
	jdff dff_B_jOXGfaj73_0(.din(w_dff_B_cqES8raJ6_0),.dout(w_dff_B_jOXGfaj73_0),.clk(gclk));
	jdff dff_B_HoMEbkSw9_0(.din(w_dff_B_jOXGfaj73_0),.dout(w_dff_B_HoMEbkSw9_0),.clk(gclk));
	jdff dff_B_bgcegKWU2_0(.din(w_dff_B_HoMEbkSw9_0),.dout(w_dff_B_bgcegKWU2_0),.clk(gclk));
	jdff dff_B_dd0p0oAi6_0(.din(w_dff_B_bgcegKWU2_0),.dout(w_dff_B_dd0p0oAi6_0),.clk(gclk));
	jdff dff_B_pusv550R7_0(.din(n1036),.dout(w_dff_B_pusv550R7_0),.clk(gclk));
	jdff dff_B_ZfxIdoRS3_0(.din(w_dff_B_pusv550R7_0),.dout(w_dff_B_ZfxIdoRS3_0),.clk(gclk));
	jdff dff_B_rZly37lq9_0(.din(w_dff_B_ZfxIdoRS3_0),.dout(w_dff_B_rZly37lq9_0),.clk(gclk));
	jdff dff_B_1QrxlgIi3_0(.din(w_dff_B_rZly37lq9_0),.dout(w_dff_B_1QrxlgIi3_0),.clk(gclk));
	jdff dff_B_EZ3bjkOA6_0(.din(w_dff_B_1QrxlgIi3_0),.dout(w_dff_B_EZ3bjkOA6_0),.clk(gclk));
	jdff dff_B_atZEI2L26_0(.din(w_dff_B_EZ3bjkOA6_0),.dout(w_dff_B_atZEI2L26_0),.clk(gclk));
	jdff dff_B_zN2WAg558_0(.din(w_dff_B_atZEI2L26_0),.dout(w_dff_B_zN2WAg558_0),.clk(gclk));
	jdff dff_B_oqDDBQ8k8_0(.din(w_dff_B_zN2WAg558_0),.dout(w_dff_B_oqDDBQ8k8_0),.clk(gclk));
	jdff dff_B_sPJWm7tm8_0(.din(w_dff_B_oqDDBQ8k8_0),.dout(w_dff_B_sPJWm7tm8_0),.clk(gclk));
	jdff dff_B_cx7ciW4N5_0(.din(w_dff_B_sPJWm7tm8_0),.dout(w_dff_B_cx7ciW4N5_0),.clk(gclk));
	jdff dff_B_8jr8A6wf2_0(.din(w_dff_B_cx7ciW4N5_0),.dout(w_dff_B_8jr8A6wf2_0),.clk(gclk));
	jdff dff_B_fKPhdPw80_0(.din(w_dff_B_8jr8A6wf2_0),.dout(w_dff_B_fKPhdPw80_0),.clk(gclk));
	jdff dff_B_ArPEip2A9_0(.din(w_dff_B_fKPhdPw80_0),.dout(w_dff_B_ArPEip2A9_0),.clk(gclk));
	jdff dff_B_w6Y4u58X5_0(.din(w_dff_B_ArPEip2A9_0),.dout(w_dff_B_w6Y4u58X5_0),.clk(gclk));
	jdff dff_B_DyWZwweL9_0(.din(w_dff_B_w6Y4u58X5_0),.dout(w_dff_B_DyWZwweL9_0),.clk(gclk));
	jdff dff_B_NTvxV2DC0_0(.din(w_dff_B_DyWZwweL9_0),.dout(w_dff_B_NTvxV2DC0_0),.clk(gclk));
	jdff dff_B_Vyjyv6Y98_0(.din(w_dff_B_NTvxV2DC0_0),.dout(w_dff_B_Vyjyv6Y98_0),.clk(gclk));
	jdff dff_B_hj3vrpnk2_0(.din(w_dff_B_Vyjyv6Y98_0),.dout(w_dff_B_hj3vrpnk2_0),.clk(gclk));
	jdff dff_B_Yx31Y2yi2_0(.din(w_dff_B_hj3vrpnk2_0),.dout(w_dff_B_Yx31Y2yi2_0),.clk(gclk));
	jdff dff_B_wzDVvkSD5_0(.din(w_dff_B_Yx31Y2yi2_0),.dout(w_dff_B_wzDVvkSD5_0),.clk(gclk));
	jdff dff_B_NkXuCfbI5_0(.din(w_dff_B_wzDVvkSD5_0),.dout(w_dff_B_NkXuCfbI5_0),.clk(gclk));
	jdff dff_B_ApEmhpxu8_0(.din(w_dff_B_NkXuCfbI5_0),.dout(w_dff_B_ApEmhpxu8_0),.clk(gclk));
	jdff dff_B_iXWoM0wB9_0(.din(w_dff_B_ApEmhpxu8_0),.dout(w_dff_B_iXWoM0wB9_0),.clk(gclk));
	jdff dff_B_FDhDBvSa8_0(.din(w_dff_B_iXWoM0wB9_0),.dout(w_dff_B_FDhDBvSa8_0),.clk(gclk));
	jdff dff_B_U9FQO6r42_0(.din(w_dff_B_FDhDBvSa8_0),.dout(w_dff_B_U9FQO6r42_0),.clk(gclk));
	jdff dff_B_AobR9bnN8_0(.din(w_dff_B_U9FQO6r42_0),.dout(w_dff_B_AobR9bnN8_0),.clk(gclk));
	jdff dff_B_DGFQE7b14_0(.din(w_dff_B_AobR9bnN8_0),.dout(w_dff_B_DGFQE7b14_0),.clk(gclk));
	jdff dff_B_z9SRrJur5_0(.din(w_dff_B_DGFQE7b14_0),.dout(w_dff_B_z9SRrJur5_0),.clk(gclk));
	jdff dff_B_VDGxEkFo7_0(.din(w_dff_B_z9SRrJur5_0),.dout(w_dff_B_VDGxEkFo7_0),.clk(gclk));
	jdff dff_B_CVH01MXj6_0(.din(w_dff_B_VDGxEkFo7_0),.dout(w_dff_B_CVH01MXj6_0),.clk(gclk));
	jdff dff_B_DGJOucNC7_0(.din(w_dff_B_CVH01MXj6_0),.dout(w_dff_B_DGJOucNC7_0),.clk(gclk));
	jdff dff_B_T0dICz7U5_0(.din(w_dff_B_DGJOucNC7_0),.dout(w_dff_B_T0dICz7U5_0),.clk(gclk));
	jdff dff_B_B1x4mKxj2_0(.din(w_dff_B_T0dICz7U5_0),.dout(w_dff_B_B1x4mKxj2_0),.clk(gclk));
	jdff dff_B_oJ9BwWfd6_0(.din(w_dff_B_B1x4mKxj2_0),.dout(w_dff_B_oJ9BwWfd6_0),.clk(gclk));
	jdff dff_B_9UTPLhqN1_0(.din(w_dff_B_oJ9BwWfd6_0),.dout(w_dff_B_9UTPLhqN1_0),.clk(gclk));
	jdff dff_B_4OocKqtL1_0(.din(w_dff_B_9UTPLhqN1_0),.dout(w_dff_B_4OocKqtL1_0),.clk(gclk));
	jdff dff_B_TA3qS7rS4_0(.din(w_dff_B_4OocKqtL1_0),.dout(w_dff_B_TA3qS7rS4_0),.clk(gclk));
	jdff dff_B_lZUXb3am7_0(.din(w_dff_B_TA3qS7rS4_0),.dout(w_dff_B_lZUXb3am7_0),.clk(gclk));
	jdff dff_B_1ztAo8ZS5_0(.din(w_dff_B_lZUXb3am7_0),.dout(w_dff_B_1ztAo8ZS5_0),.clk(gclk));
	jdff dff_B_SAc63fLB8_0(.din(w_dff_B_1ztAo8ZS5_0),.dout(w_dff_B_SAc63fLB8_0),.clk(gclk));
	jdff dff_B_anKfKQCv4_0(.din(w_dff_B_SAc63fLB8_0),.dout(w_dff_B_anKfKQCv4_0),.clk(gclk));
	jdff dff_B_P4nZcRXe7_0(.din(w_dff_B_anKfKQCv4_0),.dout(w_dff_B_P4nZcRXe7_0),.clk(gclk));
	jdff dff_B_iddLDsQe1_0(.din(w_dff_B_P4nZcRXe7_0),.dout(w_dff_B_iddLDsQe1_0),.clk(gclk));
	jdff dff_B_ac51NJ8M5_0(.din(w_dff_B_iddLDsQe1_0),.dout(w_dff_B_ac51NJ8M5_0),.clk(gclk));
	jdff dff_B_YcwgTnpQ1_0(.din(w_dff_B_ac51NJ8M5_0),.dout(w_dff_B_YcwgTnpQ1_0),.clk(gclk));
	jdff dff_B_o0JTq3177_0(.din(w_dff_B_YcwgTnpQ1_0),.dout(w_dff_B_o0JTq3177_0),.clk(gclk));
	jdff dff_B_V8yniEIl3_0(.din(w_dff_B_o0JTq3177_0),.dout(w_dff_B_V8yniEIl3_0),.clk(gclk));
	jdff dff_B_w0bV01dU2_0(.din(w_dff_B_V8yniEIl3_0),.dout(w_dff_B_w0bV01dU2_0),.clk(gclk));
	jdff dff_B_cHBo464i5_0(.din(w_dff_B_w0bV01dU2_0),.dout(w_dff_B_cHBo464i5_0),.clk(gclk));
	jdff dff_B_kzpLcWcb2_0(.din(w_dff_B_cHBo464i5_0),.dout(w_dff_B_kzpLcWcb2_0),.clk(gclk));
	jdff dff_B_R52MuZJ14_0(.din(w_dff_B_kzpLcWcb2_0),.dout(w_dff_B_R52MuZJ14_0),.clk(gclk));
	jdff dff_B_nQfUyDek2_0(.din(w_dff_B_R52MuZJ14_0),.dout(w_dff_B_nQfUyDek2_0),.clk(gclk));
	jdff dff_B_EM6Q6fXr3_0(.din(w_dff_B_nQfUyDek2_0),.dout(w_dff_B_EM6Q6fXr3_0),.clk(gclk));
	jdff dff_B_39990Mc98_0(.din(w_dff_B_EM6Q6fXr3_0),.dout(w_dff_B_39990Mc98_0),.clk(gclk));
	jdff dff_B_K8OexuYb9_0(.din(w_dff_B_39990Mc98_0),.dout(w_dff_B_K8OexuYb9_0),.clk(gclk));
	jdff dff_B_wiGiQNyH2_0(.din(w_dff_B_K8OexuYb9_0),.dout(w_dff_B_wiGiQNyH2_0),.clk(gclk));
	jdff dff_B_reHKeMie8_0(.din(w_dff_B_wiGiQNyH2_0),.dout(w_dff_B_reHKeMie8_0),.clk(gclk));
	jdff dff_B_npM5Nl0O6_0(.din(w_dff_B_reHKeMie8_0),.dout(w_dff_B_npM5Nl0O6_0),.clk(gclk));
	jdff dff_B_2OoijRqk8_0(.din(w_dff_B_npM5Nl0O6_0),.dout(w_dff_B_2OoijRqk8_0),.clk(gclk));
	jdff dff_B_mxRnyncP0_0(.din(w_dff_B_2OoijRqk8_0),.dout(w_dff_B_mxRnyncP0_0),.clk(gclk));
	jdff dff_B_u2obqZvQ8_0(.din(w_dff_B_mxRnyncP0_0),.dout(w_dff_B_u2obqZvQ8_0),.clk(gclk));
	jdff dff_B_23XQ23Vq8_0(.din(w_dff_B_u2obqZvQ8_0),.dout(w_dff_B_23XQ23Vq8_0),.clk(gclk));
	jdff dff_B_HOoJjIW81_0(.din(w_dff_B_23XQ23Vq8_0),.dout(w_dff_B_HOoJjIW81_0),.clk(gclk));
	jdff dff_B_8jGzfMY66_0(.din(w_dff_B_HOoJjIW81_0),.dout(w_dff_B_8jGzfMY66_0),.clk(gclk));
	jdff dff_B_Y5OzA62R8_0(.din(w_dff_B_8jGzfMY66_0),.dout(w_dff_B_Y5OzA62R8_0),.clk(gclk));
	jdff dff_B_x052kdxA0_0(.din(w_dff_B_Y5OzA62R8_0),.dout(w_dff_B_x052kdxA0_0),.clk(gclk));
	jdff dff_B_WvdaZn920_0(.din(w_dff_B_x052kdxA0_0),.dout(w_dff_B_WvdaZn920_0),.clk(gclk));
	jdff dff_B_gjdPgoE86_0(.din(w_dff_B_WvdaZn920_0),.dout(w_dff_B_gjdPgoE86_0),.clk(gclk));
	jdff dff_B_nzfeVEXt0_0(.din(w_dff_B_gjdPgoE86_0),.dout(w_dff_B_nzfeVEXt0_0),.clk(gclk));
	jdff dff_B_JJ9rG2Gu2_0(.din(w_dff_B_nzfeVEXt0_0),.dout(w_dff_B_JJ9rG2Gu2_0),.clk(gclk));
	jdff dff_B_ajN1aV6p4_0(.din(w_dff_B_JJ9rG2Gu2_0),.dout(w_dff_B_ajN1aV6p4_0),.clk(gclk));
	jdff dff_B_4S2NTSbc2_0(.din(w_dff_B_ajN1aV6p4_0),.dout(w_dff_B_4S2NTSbc2_0),.clk(gclk));
	jdff dff_B_XyATiomv8_0(.din(w_dff_B_4S2NTSbc2_0),.dout(w_dff_B_XyATiomv8_0),.clk(gclk));
	jdff dff_B_CctImZ677_0(.din(w_dff_B_XyATiomv8_0),.dout(w_dff_B_CctImZ677_0),.clk(gclk));
	jdff dff_B_yUO1rcyV8_0(.din(w_dff_B_CctImZ677_0),.dout(w_dff_B_yUO1rcyV8_0),.clk(gclk));
	jdff dff_B_G1nS78DA1_0(.din(w_dff_B_yUO1rcyV8_0),.dout(w_dff_B_G1nS78DA1_0),.clk(gclk));
	jdff dff_B_UWTf4VsK0_0(.din(w_dff_B_G1nS78DA1_0),.dout(w_dff_B_UWTf4VsK0_0),.clk(gclk));
	jdff dff_B_Yks2LHNj7_0(.din(w_dff_B_UWTf4VsK0_0),.dout(w_dff_B_Yks2LHNj7_0),.clk(gclk));
	jdff dff_B_fAbiPnOI4_0(.din(w_dff_B_Yks2LHNj7_0),.dout(w_dff_B_fAbiPnOI4_0),.clk(gclk));
	jdff dff_B_Eg504Qtb6_0(.din(w_dff_B_fAbiPnOI4_0),.dout(w_dff_B_Eg504Qtb6_0),.clk(gclk));
	jdff dff_B_JDOlONTx1_0(.din(w_dff_B_Eg504Qtb6_0),.dout(w_dff_B_JDOlONTx1_0),.clk(gclk));
	jdff dff_B_2tZ2TT418_0(.din(w_dff_B_JDOlONTx1_0),.dout(w_dff_B_2tZ2TT418_0),.clk(gclk));
	jdff dff_B_bQwu2pKW1_0(.din(w_dff_B_2tZ2TT418_0),.dout(w_dff_B_bQwu2pKW1_0),.clk(gclk));
	jdff dff_B_a5tYb59C2_0(.din(w_dff_B_bQwu2pKW1_0),.dout(w_dff_B_a5tYb59C2_0),.clk(gclk));
	jdff dff_B_ggmU1zId5_0(.din(w_dff_B_a5tYb59C2_0),.dout(w_dff_B_ggmU1zId5_0),.clk(gclk));
	jdff dff_B_NpqnGBF81_0(.din(w_dff_B_ggmU1zId5_0),.dout(w_dff_B_NpqnGBF81_0),.clk(gclk));
	jdff dff_B_txZuw9hH9_0(.din(w_dff_B_NpqnGBF81_0),.dout(w_dff_B_txZuw9hH9_0),.clk(gclk));
	jdff dff_B_LE2yWl298_0(.din(w_dff_B_txZuw9hH9_0),.dout(w_dff_B_LE2yWl298_0),.clk(gclk));
	jdff dff_B_Cs0dg0j89_0(.din(w_dff_B_LE2yWl298_0),.dout(w_dff_B_Cs0dg0j89_0),.clk(gclk));
	jdff dff_B_HQ0WDu3E9_0(.din(w_dff_B_Cs0dg0j89_0),.dout(w_dff_B_HQ0WDu3E9_0),.clk(gclk));
	jdff dff_B_COKo5FpP0_0(.din(w_dff_B_HQ0WDu3E9_0),.dout(w_dff_B_COKo5FpP0_0),.clk(gclk));
	jdff dff_B_nWq3XiFw8_0(.din(w_dff_B_COKo5FpP0_0),.dout(w_dff_B_nWq3XiFw8_0),.clk(gclk));
	jdff dff_B_o12N0bDT3_0(.din(w_dff_B_nWq3XiFw8_0),.dout(w_dff_B_o12N0bDT3_0),.clk(gclk));
	jdff dff_B_TY8mE9Li0_0(.din(w_dff_B_o12N0bDT3_0),.dout(w_dff_B_TY8mE9Li0_0),.clk(gclk));
	jdff dff_B_Im30cn4y5_0(.din(w_dff_B_TY8mE9Li0_0),.dout(w_dff_B_Im30cn4y5_0),.clk(gclk));
	jdff dff_B_KF5ZAWdU8_0(.din(w_dff_B_Im30cn4y5_0),.dout(w_dff_B_KF5ZAWdU8_0),.clk(gclk));
	jdff dff_B_t9e84WK16_0(.din(w_dff_B_KF5ZAWdU8_0),.dout(w_dff_B_t9e84WK16_0),.clk(gclk));
	jdff dff_B_k6pbRaNT3_0(.din(w_dff_B_t9e84WK16_0),.dout(w_dff_B_k6pbRaNT3_0),.clk(gclk));
	jdff dff_B_MKvpkoCF0_0(.din(w_dff_B_k6pbRaNT3_0),.dout(w_dff_B_MKvpkoCF0_0),.clk(gclk));
	jdff dff_B_Yf7m6c1S4_0(.din(w_dff_B_MKvpkoCF0_0),.dout(w_dff_B_Yf7m6c1S4_0),.clk(gclk));
	jdff dff_B_3rPiMYEK0_0(.din(w_dff_B_Yf7m6c1S4_0),.dout(w_dff_B_3rPiMYEK0_0),.clk(gclk));
	jdff dff_B_MtbNuX5Z5_0(.din(w_dff_B_3rPiMYEK0_0),.dout(w_dff_B_MtbNuX5Z5_0),.clk(gclk));
	jdff dff_B_8RA9EyCE0_0(.din(w_dff_B_MtbNuX5Z5_0),.dout(w_dff_B_8RA9EyCE0_0),.clk(gclk));
	jdff dff_B_1yniShmk4_0(.din(w_dff_B_8RA9EyCE0_0),.dout(w_dff_B_1yniShmk4_0),.clk(gclk));
	jdff dff_B_3j4nDcev0_0(.din(w_dff_B_1yniShmk4_0),.dout(w_dff_B_3j4nDcev0_0),.clk(gclk));
	jdff dff_B_rz3GLmFp6_0(.din(w_dff_B_3j4nDcev0_0),.dout(w_dff_B_rz3GLmFp6_0),.clk(gclk));
	jdff dff_B_Ud3Dy1Eo2_0(.din(w_dff_B_rz3GLmFp6_0),.dout(w_dff_B_Ud3Dy1Eo2_0),.clk(gclk));
	jdff dff_B_k9DFeDPe2_0(.din(w_dff_B_Ud3Dy1Eo2_0),.dout(w_dff_B_k9DFeDPe2_0),.clk(gclk));
	jdff dff_B_lZUCSA9A3_0(.din(n1042),.dout(w_dff_B_lZUCSA9A3_0),.clk(gclk));
	jdff dff_B_fDZ95RFP3_0(.din(w_dff_B_lZUCSA9A3_0),.dout(w_dff_B_fDZ95RFP3_0),.clk(gclk));
	jdff dff_B_3GgoQRQw0_0(.din(w_dff_B_fDZ95RFP3_0),.dout(w_dff_B_3GgoQRQw0_0),.clk(gclk));
	jdff dff_B_MXq7WG1f2_0(.din(w_dff_B_3GgoQRQw0_0),.dout(w_dff_B_MXq7WG1f2_0),.clk(gclk));
	jdff dff_B_I8btYOZ85_0(.din(w_dff_B_MXq7WG1f2_0),.dout(w_dff_B_I8btYOZ85_0),.clk(gclk));
	jdff dff_B_nFWX1Tk75_0(.din(w_dff_B_I8btYOZ85_0),.dout(w_dff_B_nFWX1Tk75_0),.clk(gclk));
	jdff dff_B_rLp89D2B8_0(.din(w_dff_B_nFWX1Tk75_0),.dout(w_dff_B_rLp89D2B8_0),.clk(gclk));
	jdff dff_B_L7Kwj1N42_0(.din(w_dff_B_rLp89D2B8_0),.dout(w_dff_B_L7Kwj1N42_0),.clk(gclk));
	jdff dff_B_b12LLiXT2_0(.din(w_dff_B_L7Kwj1N42_0),.dout(w_dff_B_b12LLiXT2_0),.clk(gclk));
	jdff dff_B_mwOIfAEw8_0(.din(w_dff_B_b12LLiXT2_0),.dout(w_dff_B_mwOIfAEw8_0),.clk(gclk));
	jdff dff_B_W8EQbhah2_0(.din(w_dff_B_mwOIfAEw8_0),.dout(w_dff_B_W8EQbhah2_0),.clk(gclk));
	jdff dff_B_GDLg9PZ15_0(.din(w_dff_B_W8EQbhah2_0),.dout(w_dff_B_GDLg9PZ15_0),.clk(gclk));
	jdff dff_B_QYj8j4lR1_0(.din(w_dff_B_GDLg9PZ15_0),.dout(w_dff_B_QYj8j4lR1_0),.clk(gclk));
	jdff dff_B_9L6RF8JV8_0(.din(w_dff_B_QYj8j4lR1_0),.dout(w_dff_B_9L6RF8JV8_0),.clk(gclk));
	jdff dff_B_uznJy0lY2_0(.din(w_dff_B_9L6RF8JV8_0),.dout(w_dff_B_uznJy0lY2_0),.clk(gclk));
	jdff dff_B_ziTfRZrj3_0(.din(w_dff_B_uznJy0lY2_0),.dout(w_dff_B_ziTfRZrj3_0),.clk(gclk));
	jdff dff_B_UwgeImGO4_0(.din(w_dff_B_ziTfRZrj3_0),.dout(w_dff_B_UwgeImGO4_0),.clk(gclk));
	jdff dff_B_nF1qfK8k2_0(.din(w_dff_B_UwgeImGO4_0),.dout(w_dff_B_nF1qfK8k2_0),.clk(gclk));
	jdff dff_B_7H5KW3lH4_0(.din(w_dff_B_nF1qfK8k2_0),.dout(w_dff_B_7H5KW3lH4_0),.clk(gclk));
	jdff dff_B_BvI3xdZn8_0(.din(w_dff_B_7H5KW3lH4_0),.dout(w_dff_B_BvI3xdZn8_0),.clk(gclk));
	jdff dff_B_OaUTPC2v7_0(.din(w_dff_B_BvI3xdZn8_0),.dout(w_dff_B_OaUTPC2v7_0),.clk(gclk));
	jdff dff_B_trzzL8lt6_0(.din(w_dff_B_OaUTPC2v7_0),.dout(w_dff_B_trzzL8lt6_0),.clk(gclk));
	jdff dff_B_VHdkFBLW9_0(.din(w_dff_B_trzzL8lt6_0),.dout(w_dff_B_VHdkFBLW9_0),.clk(gclk));
	jdff dff_B_ah5RcUrR1_0(.din(w_dff_B_VHdkFBLW9_0),.dout(w_dff_B_ah5RcUrR1_0),.clk(gclk));
	jdff dff_B_JPiWC0wi9_0(.din(w_dff_B_ah5RcUrR1_0),.dout(w_dff_B_JPiWC0wi9_0),.clk(gclk));
	jdff dff_B_L5Pucexw8_0(.din(w_dff_B_JPiWC0wi9_0),.dout(w_dff_B_L5Pucexw8_0),.clk(gclk));
	jdff dff_B_docg3eac9_0(.din(w_dff_B_L5Pucexw8_0),.dout(w_dff_B_docg3eac9_0),.clk(gclk));
	jdff dff_B_EttfWhTC3_0(.din(w_dff_B_docg3eac9_0),.dout(w_dff_B_EttfWhTC3_0),.clk(gclk));
	jdff dff_B_nSUBjaxG9_0(.din(w_dff_B_EttfWhTC3_0),.dout(w_dff_B_nSUBjaxG9_0),.clk(gclk));
	jdff dff_B_bdW7SarL9_0(.din(w_dff_B_nSUBjaxG9_0),.dout(w_dff_B_bdW7SarL9_0),.clk(gclk));
	jdff dff_B_Jjdj1cZ71_0(.din(w_dff_B_bdW7SarL9_0),.dout(w_dff_B_Jjdj1cZ71_0),.clk(gclk));
	jdff dff_B_BdHYiJcT4_0(.din(w_dff_B_Jjdj1cZ71_0),.dout(w_dff_B_BdHYiJcT4_0),.clk(gclk));
	jdff dff_B_3HtbydAD1_0(.din(w_dff_B_BdHYiJcT4_0),.dout(w_dff_B_3HtbydAD1_0),.clk(gclk));
	jdff dff_B_g9GROpv34_0(.din(w_dff_B_3HtbydAD1_0),.dout(w_dff_B_g9GROpv34_0),.clk(gclk));
	jdff dff_B_LrwqCsfY0_0(.din(w_dff_B_g9GROpv34_0),.dout(w_dff_B_LrwqCsfY0_0),.clk(gclk));
	jdff dff_B_Db0V13Qf3_0(.din(w_dff_B_LrwqCsfY0_0),.dout(w_dff_B_Db0V13Qf3_0),.clk(gclk));
	jdff dff_B_wAxo6ZkR6_0(.din(w_dff_B_Db0V13Qf3_0),.dout(w_dff_B_wAxo6ZkR6_0),.clk(gclk));
	jdff dff_B_hcyqwcDR8_0(.din(w_dff_B_wAxo6ZkR6_0),.dout(w_dff_B_hcyqwcDR8_0),.clk(gclk));
	jdff dff_B_ncfYkBw05_0(.din(w_dff_B_hcyqwcDR8_0),.dout(w_dff_B_ncfYkBw05_0),.clk(gclk));
	jdff dff_B_NEcMygc96_0(.din(w_dff_B_ncfYkBw05_0),.dout(w_dff_B_NEcMygc96_0),.clk(gclk));
	jdff dff_B_MnPQDsx59_0(.din(w_dff_B_NEcMygc96_0),.dout(w_dff_B_MnPQDsx59_0),.clk(gclk));
	jdff dff_B_BfVf1e9F2_0(.din(w_dff_B_MnPQDsx59_0),.dout(w_dff_B_BfVf1e9F2_0),.clk(gclk));
	jdff dff_B_Pw2BAIRZ8_0(.din(w_dff_B_BfVf1e9F2_0),.dout(w_dff_B_Pw2BAIRZ8_0),.clk(gclk));
	jdff dff_B_ciTHcdW91_0(.din(w_dff_B_Pw2BAIRZ8_0),.dout(w_dff_B_ciTHcdW91_0),.clk(gclk));
	jdff dff_B_oMPmOW1m6_0(.din(w_dff_B_ciTHcdW91_0),.dout(w_dff_B_oMPmOW1m6_0),.clk(gclk));
	jdff dff_B_0aip3RuV9_0(.din(w_dff_B_oMPmOW1m6_0),.dout(w_dff_B_0aip3RuV9_0),.clk(gclk));
	jdff dff_B_WCUJ3gjy9_0(.din(w_dff_B_0aip3RuV9_0),.dout(w_dff_B_WCUJ3gjy9_0),.clk(gclk));
	jdff dff_B_Y5Tp0Aqu1_0(.din(w_dff_B_WCUJ3gjy9_0),.dout(w_dff_B_Y5Tp0Aqu1_0),.clk(gclk));
	jdff dff_B_ZSVpoMic1_0(.din(w_dff_B_Y5Tp0Aqu1_0),.dout(w_dff_B_ZSVpoMic1_0),.clk(gclk));
	jdff dff_B_lUKJVG9c5_0(.din(w_dff_B_ZSVpoMic1_0),.dout(w_dff_B_lUKJVG9c5_0),.clk(gclk));
	jdff dff_B_53hN5EYA5_0(.din(w_dff_B_lUKJVG9c5_0),.dout(w_dff_B_53hN5EYA5_0),.clk(gclk));
	jdff dff_B_BuFh8Hxo2_0(.din(w_dff_B_53hN5EYA5_0),.dout(w_dff_B_BuFh8Hxo2_0),.clk(gclk));
	jdff dff_B_4P6ybyWZ9_0(.din(w_dff_B_BuFh8Hxo2_0),.dout(w_dff_B_4P6ybyWZ9_0),.clk(gclk));
	jdff dff_B_oBP6ETy65_0(.din(w_dff_B_4P6ybyWZ9_0),.dout(w_dff_B_oBP6ETy65_0),.clk(gclk));
	jdff dff_B_POlv0clL2_0(.din(w_dff_B_oBP6ETy65_0),.dout(w_dff_B_POlv0clL2_0),.clk(gclk));
	jdff dff_B_GQ59k3ax2_0(.din(w_dff_B_POlv0clL2_0),.dout(w_dff_B_GQ59k3ax2_0),.clk(gclk));
	jdff dff_B_q8D3XDFy9_0(.din(w_dff_B_GQ59k3ax2_0),.dout(w_dff_B_q8D3XDFy9_0),.clk(gclk));
	jdff dff_B_H4XpqHqe1_0(.din(w_dff_B_q8D3XDFy9_0),.dout(w_dff_B_H4XpqHqe1_0),.clk(gclk));
	jdff dff_B_OG2uWAfO8_0(.din(w_dff_B_H4XpqHqe1_0),.dout(w_dff_B_OG2uWAfO8_0),.clk(gclk));
	jdff dff_B_1ZXxUS0t8_0(.din(w_dff_B_OG2uWAfO8_0),.dout(w_dff_B_1ZXxUS0t8_0),.clk(gclk));
	jdff dff_B_uSbo473H4_0(.din(w_dff_B_1ZXxUS0t8_0),.dout(w_dff_B_uSbo473H4_0),.clk(gclk));
	jdff dff_B_G0PN0gDH2_0(.din(w_dff_B_uSbo473H4_0),.dout(w_dff_B_G0PN0gDH2_0),.clk(gclk));
	jdff dff_B_nVnr4XIg6_0(.din(w_dff_B_G0PN0gDH2_0),.dout(w_dff_B_nVnr4XIg6_0),.clk(gclk));
	jdff dff_B_w5tC6RVB7_0(.din(w_dff_B_nVnr4XIg6_0),.dout(w_dff_B_w5tC6RVB7_0),.clk(gclk));
	jdff dff_B_Cwao2zTs7_0(.din(w_dff_B_w5tC6RVB7_0),.dout(w_dff_B_Cwao2zTs7_0),.clk(gclk));
	jdff dff_B_IHOCXAD78_0(.din(w_dff_B_Cwao2zTs7_0),.dout(w_dff_B_IHOCXAD78_0),.clk(gclk));
	jdff dff_B_WD6Z4xBB3_0(.din(w_dff_B_IHOCXAD78_0),.dout(w_dff_B_WD6Z4xBB3_0),.clk(gclk));
	jdff dff_B_m56xR5qt0_0(.din(w_dff_B_WD6Z4xBB3_0),.dout(w_dff_B_m56xR5qt0_0),.clk(gclk));
	jdff dff_B_ceT84vat9_0(.din(w_dff_B_m56xR5qt0_0),.dout(w_dff_B_ceT84vat9_0),.clk(gclk));
	jdff dff_B_CdsB3iVe2_0(.din(w_dff_B_ceT84vat9_0),.dout(w_dff_B_CdsB3iVe2_0),.clk(gclk));
	jdff dff_B_G2vBjQl91_0(.din(w_dff_B_CdsB3iVe2_0),.dout(w_dff_B_G2vBjQl91_0),.clk(gclk));
	jdff dff_B_FzuzKVaR2_0(.din(w_dff_B_G2vBjQl91_0),.dout(w_dff_B_FzuzKVaR2_0),.clk(gclk));
	jdff dff_B_OXEH8LOc4_0(.din(w_dff_B_FzuzKVaR2_0),.dout(w_dff_B_OXEH8LOc4_0),.clk(gclk));
	jdff dff_B_phXZYXDE9_0(.din(w_dff_B_OXEH8LOc4_0),.dout(w_dff_B_phXZYXDE9_0),.clk(gclk));
	jdff dff_B_tJjvCFaF8_0(.din(w_dff_B_phXZYXDE9_0),.dout(w_dff_B_tJjvCFaF8_0),.clk(gclk));
	jdff dff_B_CG3qYiiH9_0(.din(w_dff_B_tJjvCFaF8_0),.dout(w_dff_B_CG3qYiiH9_0),.clk(gclk));
	jdff dff_B_LGaA90wP8_0(.din(w_dff_B_CG3qYiiH9_0),.dout(w_dff_B_LGaA90wP8_0),.clk(gclk));
	jdff dff_B_8qh9t5cc0_0(.din(w_dff_B_LGaA90wP8_0),.dout(w_dff_B_8qh9t5cc0_0),.clk(gclk));
	jdff dff_B_GP7jMlkS5_0(.din(w_dff_B_8qh9t5cc0_0),.dout(w_dff_B_GP7jMlkS5_0),.clk(gclk));
	jdff dff_B_QZNtyzr55_0(.din(w_dff_B_GP7jMlkS5_0),.dout(w_dff_B_QZNtyzr55_0),.clk(gclk));
	jdff dff_B_QXBGWgRV9_0(.din(w_dff_B_QZNtyzr55_0),.dout(w_dff_B_QXBGWgRV9_0),.clk(gclk));
	jdff dff_B_QjiUcXlb3_0(.din(w_dff_B_QXBGWgRV9_0),.dout(w_dff_B_QjiUcXlb3_0),.clk(gclk));
	jdff dff_B_eAL6qBVp8_0(.din(w_dff_B_QjiUcXlb3_0),.dout(w_dff_B_eAL6qBVp8_0),.clk(gclk));
	jdff dff_B_pPhVScum2_0(.din(w_dff_B_eAL6qBVp8_0),.dout(w_dff_B_pPhVScum2_0),.clk(gclk));
	jdff dff_B_Wn6DD4PA5_0(.din(w_dff_B_pPhVScum2_0),.dout(w_dff_B_Wn6DD4PA5_0),.clk(gclk));
	jdff dff_B_o5K0aP9q2_0(.din(w_dff_B_Wn6DD4PA5_0),.dout(w_dff_B_o5K0aP9q2_0),.clk(gclk));
	jdff dff_B_x1rHUAFq1_0(.din(w_dff_B_o5K0aP9q2_0),.dout(w_dff_B_x1rHUAFq1_0),.clk(gclk));
	jdff dff_B_uuZXmYkW8_0(.din(w_dff_B_x1rHUAFq1_0),.dout(w_dff_B_uuZXmYkW8_0),.clk(gclk));
	jdff dff_B_mzYG1aHG2_0(.din(w_dff_B_uuZXmYkW8_0),.dout(w_dff_B_mzYG1aHG2_0),.clk(gclk));
	jdff dff_B_9qakpVN09_0(.din(w_dff_B_mzYG1aHG2_0),.dout(w_dff_B_9qakpVN09_0),.clk(gclk));
	jdff dff_B_zUZPMoaj8_0(.din(w_dff_B_9qakpVN09_0),.dout(w_dff_B_zUZPMoaj8_0),.clk(gclk));
	jdff dff_B_28AEySVh9_0(.din(w_dff_B_zUZPMoaj8_0),.dout(w_dff_B_28AEySVh9_0),.clk(gclk));
	jdff dff_B_L4vt9y447_0(.din(w_dff_B_28AEySVh9_0),.dout(w_dff_B_L4vt9y447_0),.clk(gclk));
	jdff dff_B_cIYLqHl43_0(.din(w_dff_B_L4vt9y447_0),.dout(w_dff_B_cIYLqHl43_0),.clk(gclk));
	jdff dff_B_jV6OSf7h7_0(.din(w_dff_B_cIYLqHl43_0),.dout(w_dff_B_jV6OSf7h7_0),.clk(gclk));
	jdff dff_B_ifZD6cu69_0(.din(w_dff_B_jV6OSf7h7_0),.dout(w_dff_B_ifZD6cu69_0),.clk(gclk));
	jdff dff_B_WQMoiER83_0(.din(w_dff_B_ifZD6cu69_0),.dout(w_dff_B_WQMoiER83_0),.clk(gclk));
	jdff dff_B_pFexGzC92_0(.din(w_dff_B_WQMoiER83_0),.dout(w_dff_B_pFexGzC92_0),.clk(gclk));
	jdff dff_B_JqB01Iod7_0(.din(w_dff_B_pFexGzC92_0),.dout(w_dff_B_JqB01Iod7_0),.clk(gclk));
	jdff dff_B_p3DsJkDf3_0(.din(w_dff_B_JqB01Iod7_0),.dout(w_dff_B_p3DsJkDf3_0),.clk(gclk));
	jdff dff_B_utjsIphL0_0(.din(w_dff_B_p3DsJkDf3_0),.dout(w_dff_B_utjsIphL0_0),.clk(gclk));
	jdff dff_B_Fg3yS2qD6_0(.din(w_dff_B_utjsIphL0_0),.dout(w_dff_B_Fg3yS2qD6_0),.clk(gclk));
	jdff dff_B_TATfofGL1_0(.din(w_dff_B_Fg3yS2qD6_0),.dout(w_dff_B_TATfofGL1_0),.clk(gclk));
	jdff dff_B_mWTzbsI77_0(.din(w_dff_B_TATfofGL1_0),.dout(w_dff_B_mWTzbsI77_0),.clk(gclk));
	jdff dff_B_o03zHjcG7_0(.din(w_dff_B_mWTzbsI77_0),.dout(w_dff_B_o03zHjcG7_0),.clk(gclk));
	jdff dff_B_YY7BsTrf3_0(.din(w_dff_B_o03zHjcG7_0),.dout(w_dff_B_YY7BsTrf3_0),.clk(gclk));
	jdff dff_B_KgQKlFF93_0(.din(w_dff_B_YY7BsTrf3_0),.dout(w_dff_B_KgQKlFF93_0),.clk(gclk));
	jdff dff_B_Ttqi03tx6_0(.din(w_dff_B_KgQKlFF93_0),.dout(w_dff_B_Ttqi03tx6_0),.clk(gclk));
	jdff dff_B_H2Dnf3dc2_0(.din(w_dff_B_Ttqi03tx6_0),.dout(w_dff_B_H2Dnf3dc2_0),.clk(gclk));
	jdff dff_B_CM7jz7L08_0(.din(n1048),.dout(w_dff_B_CM7jz7L08_0),.clk(gclk));
	jdff dff_B_PGqEwNli6_0(.din(w_dff_B_CM7jz7L08_0),.dout(w_dff_B_PGqEwNli6_0),.clk(gclk));
	jdff dff_B_jZykDcjk1_0(.din(w_dff_B_PGqEwNli6_0),.dout(w_dff_B_jZykDcjk1_0),.clk(gclk));
	jdff dff_B_BGJcRS4d6_0(.din(w_dff_B_jZykDcjk1_0),.dout(w_dff_B_BGJcRS4d6_0),.clk(gclk));
	jdff dff_B_fTkniR4A9_0(.din(w_dff_B_BGJcRS4d6_0),.dout(w_dff_B_fTkniR4A9_0),.clk(gclk));
	jdff dff_B_ma8ElqK70_0(.din(w_dff_B_fTkniR4A9_0),.dout(w_dff_B_ma8ElqK70_0),.clk(gclk));
	jdff dff_B_jo4cFnr11_0(.din(w_dff_B_ma8ElqK70_0),.dout(w_dff_B_jo4cFnr11_0),.clk(gclk));
	jdff dff_B_t9ovZgvW0_0(.din(w_dff_B_jo4cFnr11_0),.dout(w_dff_B_t9ovZgvW0_0),.clk(gclk));
	jdff dff_B_meG5Ji8a6_0(.din(w_dff_B_t9ovZgvW0_0),.dout(w_dff_B_meG5Ji8a6_0),.clk(gclk));
	jdff dff_B_UpNu6R1R2_0(.din(w_dff_B_meG5Ji8a6_0),.dout(w_dff_B_UpNu6R1R2_0),.clk(gclk));
	jdff dff_B_ltHfzfbS9_0(.din(w_dff_B_UpNu6R1R2_0),.dout(w_dff_B_ltHfzfbS9_0),.clk(gclk));
	jdff dff_B_pW1NiX0c2_0(.din(w_dff_B_ltHfzfbS9_0),.dout(w_dff_B_pW1NiX0c2_0),.clk(gclk));
	jdff dff_B_5mzjNiO58_0(.din(w_dff_B_pW1NiX0c2_0),.dout(w_dff_B_5mzjNiO58_0),.clk(gclk));
	jdff dff_B_QXSd3mEE7_0(.din(w_dff_B_5mzjNiO58_0),.dout(w_dff_B_QXSd3mEE7_0),.clk(gclk));
	jdff dff_B_XQFCNxae4_0(.din(w_dff_B_QXSd3mEE7_0),.dout(w_dff_B_XQFCNxae4_0),.clk(gclk));
	jdff dff_B_E5PzlMqY3_0(.din(w_dff_B_XQFCNxae4_0),.dout(w_dff_B_E5PzlMqY3_0),.clk(gclk));
	jdff dff_B_qJ6D9iMz5_0(.din(w_dff_B_E5PzlMqY3_0),.dout(w_dff_B_qJ6D9iMz5_0),.clk(gclk));
	jdff dff_B_Uo8qwJ6z1_0(.din(w_dff_B_qJ6D9iMz5_0),.dout(w_dff_B_Uo8qwJ6z1_0),.clk(gclk));
	jdff dff_B_lf3JsRov0_0(.din(w_dff_B_Uo8qwJ6z1_0),.dout(w_dff_B_lf3JsRov0_0),.clk(gclk));
	jdff dff_B_fykQMdf01_0(.din(w_dff_B_lf3JsRov0_0),.dout(w_dff_B_fykQMdf01_0),.clk(gclk));
	jdff dff_B_neOMRHVV8_0(.din(w_dff_B_fykQMdf01_0),.dout(w_dff_B_neOMRHVV8_0),.clk(gclk));
	jdff dff_B_KXmHRlCq2_0(.din(w_dff_B_neOMRHVV8_0),.dout(w_dff_B_KXmHRlCq2_0),.clk(gclk));
	jdff dff_B_dI6UbY0n8_0(.din(w_dff_B_KXmHRlCq2_0),.dout(w_dff_B_dI6UbY0n8_0),.clk(gclk));
	jdff dff_B_xy4ZFNtu2_0(.din(w_dff_B_dI6UbY0n8_0),.dout(w_dff_B_xy4ZFNtu2_0),.clk(gclk));
	jdff dff_B_mNkORTe84_0(.din(w_dff_B_xy4ZFNtu2_0),.dout(w_dff_B_mNkORTe84_0),.clk(gclk));
	jdff dff_B_QvfpEdGf5_0(.din(w_dff_B_mNkORTe84_0),.dout(w_dff_B_QvfpEdGf5_0),.clk(gclk));
	jdff dff_B_pJs4pl4V2_0(.din(w_dff_B_QvfpEdGf5_0),.dout(w_dff_B_pJs4pl4V2_0),.clk(gclk));
	jdff dff_B_VPSKlS1d6_0(.din(w_dff_B_pJs4pl4V2_0),.dout(w_dff_B_VPSKlS1d6_0),.clk(gclk));
	jdff dff_B_PYd4ZtCy6_0(.din(w_dff_B_VPSKlS1d6_0),.dout(w_dff_B_PYd4ZtCy6_0),.clk(gclk));
	jdff dff_B_iiWokwY60_0(.din(w_dff_B_PYd4ZtCy6_0),.dout(w_dff_B_iiWokwY60_0),.clk(gclk));
	jdff dff_B_WP0JqA5K8_0(.din(w_dff_B_iiWokwY60_0),.dout(w_dff_B_WP0JqA5K8_0),.clk(gclk));
	jdff dff_B_0gnvdIXO5_0(.din(w_dff_B_WP0JqA5K8_0),.dout(w_dff_B_0gnvdIXO5_0),.clk(gclk));
	jdff dff_B_ZrazR2MC9_0(.din(w_dff_B_0gnvdIXO5_0),.dout(w_dff_B_ZrazR2MC9_0),.clk(gclk));
	jdff dff_B_Bbw3HlHC5_0(.din(w_dff_B_ZrazR2MC9_0),.dout(w_dff_B_Bbw3HlHC5_0),.clk(gclk));
	jdff dff_B_WLcoUUuU8_0(.din(w_dff_B_Bbw3HlHC5_0),.dout(w_dff_B_WLcoUUuU8_0),.clk(gclk));
	jdff dff_B_bkixuBlO8_0(.din(w_dff_B_WLcoUUuU8_0),.dout(w_dff_B_bkixuBlO8_0),.clk(gclk));
	jdff dff_B_MbqnRTuo1_0(.din(w_dff_B_bkixuBlO8_0),.dout(w_dff_B_MbqnRTuo1_0),.clk(gclk));
	jdff dff_B_expjBXjo4_0(.din(w_dff_B_MbqnRTuo1_0),.dout(w_dff_B_expjBXjo4_0),.clk(gclk));
	jdff dff_B_f3hIg0vi4_0(.din(w_dff_B_expjBXjo4_0),.dout(w_dff_B_f3hIg0vi4_0),.clk(gclk));
	jdff dff_B_J1HiIVl22_0(.din(w_dff_B_f3hIg0vi4_0),.dout(w_dff_B_J1HiIVl22_0),.clk(gclk));
	jdff dff_B_ZUkjynjR4_0(.din(w_dff_B_J1HiIVl22_0),.dout(w_dff_B_ZUkjynjR4_0),.clk(gclk));
	jdff dff_B_gDu2FW9f1_0(.din(w_dff_B_ZUkjynjR4_0),.dout(w_dff_B_gDu2FW9f1_0),.clk(gclk));
	jdff dff_B_Lz0r841V0_0(.din(w_dff_B_gDu2FW9f1_0),.dout(w_dff_B_Lz0r841V0_0),.clk(gclk));
	jdff dff_B_O4JdixWM3_0(.din(w_dff_B_Lz0r841V0_0),.dout(w_dff_B_O4JdixWM3_0),.clk(gclk));
	jdff dff_B_XSzpCLky9_0(.din(w_dff_B_O4JdixWM3_0),.dout(w_dff_B_XSzpCLky9_0),.clk(gclk));
	jdff dff_B_cCy6XunU8_0(.din(w_dff_B_XSzpCLky9_0),.dout(w_dff_B_cCy6XunU8_0),.clk(gclk));
	jdff dff_B_esXN1fYe4_0(.din(w_dff_B_cCy6XunU8_0),.dout(w_dff_B_esXN1fYe4_0),.clk(gclk));
	jdff dff_B_4464nAZJ1_0(.din(w_dff_B_esXN1fYe4_0),.dout(w_dff_B_4464nAZJ1_0),.clk(gclk));
	jdff dff_B_hfxWRCUC1_0(.din(w_dff_B_4464nAZJ1_0),.dout(w_dff_B_hfxWRCUC1_0),.clk(gclk));
	jdff dff_B_3xPxFbc54_0(.din(w_dff_B_hfxWRCUC1_0),.dout(w_dff_B_3xPxFbc54_0),.clk(gclk));
	jdff dff_B_hefYU6vU4_0(.din(w_dff_B_3xPxFbc54_0),.dout(w_dff_B_hefYU6vU4_0),.clk(gclk));
	jdff dff_B_AnswcnUc9_0(.din(w_dff_B_hefYU6vU4_0),.dout(w_dff_B_AnswcnUc9_0),.clk(gclk));
	jdff dff_B_nywxU3Bl1_0(.din(w_dff_B_AnswcnUc9_0),.dout(w_dff_B_nywxU3Bl1_0),.clk(gclk));
	jdff dff_B_t4sWVa0J3_0(.din(w_dff_B_nywxU3Bl1_0),.dout(w_dff_B_t4sWVa0J3_0),.clk(gclk));
	jdff dff_B_dC93gKEJ0_0(.din(w_dff_B_t4sWVa0J3_0),.dout(w_dff_B_dC93gKEJ0_0),.clk(gclk));
	jdff dff_B_GgBrDkta4_0(.din(w_dff_B_dC93gKEJ0_0),.dout(w_dff_B_GgBrDkta4_0),.clk(gclk));
	jdff dff_B_ATHHpgLz9_0(.din(w_dff_B_GgBrDkta4_0),.dout(w_dff_B_ATHHpgLz9_0),.clk(gclk));
	jdff dff_B_C7TWCQnK1_0(.din(w_dff_B_ATHHpgLz9_0),.dout(w_dff_B_C7TWCQnK1_0),.clk(gclk));
	jdff dff_B_RnCEMxAh9_0(.din(w_dff_B_C7TWCQnK1_0),.dout(w_dff_B_RnCEMxAh9_0),.clk(gclk));
	jdff dff_B_N56pYF8L2_0(.din(w_dff_B_RnCEMxAh9_0),.dout(w_dff_B_N56pYF8L2_0),.clk(gclk));
	jdff dff_B_4t2jEr5f5_0(.din(w_dff_B_N56pYF8L2_0),.dout(w_dff_B_4t2jEr5f5_0),.clk(gclk));
	jdff dff_B_8ausr4H82_0(.din(w_dff_B_4t2jEr5f5_0),.dout(w_dff_B_8ausr4H82_0),.clk(gclk));
	jdff dff_B_sLFdCexR5_0(.din(w_dff_B_8ausr4H82_0),.dout(w_dff_B_sLFdCexR5_0),.clk(gclk));
	jdff dff_B_wbwvO3oo7_0(.din(w_dff_B_sLFdCexR5_0),.dout(w_dff_B_wbwvO3oo7_0),.clk(gclk));
	jdff dff_B_wO1NqDRk2_0(.din(w_dff_B_wbwvO3oo7_0),.dout(w_dff_B_wO1NqDRk2_0),.clk(gclk));
	jdff dff_B_OG4wtSEy2_0(.din(w_dff_B_wO1NqDRk2_0),.dout(w_dff_B_OG4wtSEy2_0),.clk(gclk));
	jdff dff_B_CJvIfNUT8_0(.din(w_dff_B_OG4wtSEy2_0),.dout(w_dff_B_CJvIfNUT8_0),.clk(gclk));
	jdff dff_B_SuZOm4Q02_0(.din(w_dff_B_CJvIfNUT8_0),.dout(w_dff_B_SuZOm4Q02_0),.clk(gclk));
	jdff dff_B_z1ngT9Rg6_0(.din(w_dff_B_SuZOm4Q02_0),.dout(w_dff_B_z1ngT9Rg6_0),.clk(gclk));
	jdff dff_B_gObonihq8_0(.din(w_dff_B_z1ngT9Rg6_0),.dout(w_dff_B_gObonihq8_0),.clk(gclk));
	jdff dff_B_v6wFi9fD8_0(.din(w_dff_B_gObonihq8_0),.dout(w_dff_B_v6wFi9fD8_0),.clk(gclk));
	jdff dff_B_Y2LleHzL0_0(.din(w_dff_B_v6wFi9fD8_0),.dout(w_dff_B_Y2LleHzL0_0),.clk(gclk));
	jdff dff_B_7VoU9dqQ5_0(.din(w_dff_B_Y2LleHzL0_0),.dout(w_dff_B_7VoU9dqQ5_0),.clk(gclk));
	jdff dff_B_0xq9NL2h4_0(.din(w_dff_B_7VoU9dqQ5_0),.dout(w_dff_B_0xq9NL2h4_0),.clk(gclk));
	jdff dff_B_Q61pZNZz9_0(.din(w_dff_B_0xq9NL2h4_0),.dout(w_dff_B_Q61pZNZz9_0),.clk(gclk));
	jdff dff_B_OW9Ii3kI4_0(.din(w_dff_B_Q61pZNZz9_0),.dout(w_dff_B_OW9Ii3kI4_0),.clk(gclk));
	jdff dff_B_s59uKsJl0_0(.din(w_dff_B_OW9Ii3kI4_0),.dout(w_dff_B_s59uKsJl0_0),.clk(gclk));
	jdff dff_B_6njFsaYT2_0(.din(w_dff_B_s59uKsJl0_0),.dout(w_dff_B_6njFsaYT2_0),.clk(gclk));
	jdff dff_B_vmD25BkI0_0(.din(w_dff_B_6njFsaYT2_0),.dout(w_dff_B_vmD25BkI0_0),.clk(gclk));
	jdff dff_B_zz2aymKs5_0(.din(w_dff_B_vmD25BkI0_0),.dout(w_dff_B_zz2aymKs5_0),.clk(gclk));
	jdff dff_B_4ibYHJsS0_0(.din(w_dff_B_zz2aymKs5_0),.dout(w_dff_B_4ibYHJsS0_0),.clk(gclk));
	jdff dff_B_RNywH5tF7_0(.din(w_dff_B_4ibYHJsS0_0),.dout(w_dff_B_RNywH5tF7_0),.clk(gclk));
	jdff dff_B_FvakI0Qn7_0(.din(w_dff_B_RNywH5tF7_0),.dout(w_dff_B_FvakI0Qn7_0),.clk(gclk));
	jdff dff_B_REl8PntW2_0(.din(w_dff_B_FvakI0Qn7_0),.dout(w_dff_B_REl8PntW2_0),.clk(gclk));
	jdff dff_B_cUKjUDVY3_0(.din(w_dff_B_REl8PntW2_0),.dout(w_dff_B_cUKjUDVY3_0),.clk(gclk));
	jdff dff_B_wGFMoWCr4_0(.din(w_dff_B_cUKjUDVY3_0),.dout(w_dff_B_wGFMoWCr4_0),.clk(gclk));
	jdff dff_B_E6lARNtU6_0(.din(w_dff_B_wGFMoWCr4_0),.dout(w_dff_B_E6lARNtU6_0),.clk(gclk));
	jdff dff_B_d8vXLIM54_0(.din(w_dff_B_E6lARNtU6_0),.dout(w_dff_B_d8vXLIM54_0),.clk(gclk));
	jdff dff_B_I4LX4cDH5_0(.din(w_dff_B_d8vXLIM54_0),.dout(w_dff_B_I4LX4cDH5_0),.clk(gclk));
	jdff dff_B_zmexGCnF8_0(.din(w_dff_B_I4LX4cDH5_0),.dout(w_dff_B_zmexGCnF8_0),.clk(gclk));
	jdff dff_B_lxFPLiYd2_0(.din(w_dff_B_zmexGCnF8_0),.dout(w_dff_B_lxFPLiYd2_0),.clk(gclk));
	jdff dff_B_9l76CoSq6_0(.din(w_dff_B_lxFPLiYd2_0),.dout(w_dff_B_9l76CoSq6_0),.clk(gclk));
	jdff dff_B_lcFptnhE4_0(.din(w_dff_B_9l76CoSq6_0),.dout(w_dff_B_lcFptnhE4_0),.clk(gclk));
	jdff dff_B_09iEg04s5_0(.din(w_dff_B_lcFptnhE4_0),.dout(w_dff_B_09iEg04s5_0),.clk(gclk));
	jdff dff_B_xYXRn8HT4_0(.din(w_dff_B_09iEg04s5_0),.dout(w_dff_B_xYXRn8HT4_0),.clk(gclk));
	jdff dff_B_rJQqSIF11_0(.din(w_dff_B_xYXRn8HT4_0),.dout(w_dff_B_rJQqSIF11_0),.clk(gclk));
	jdff dff_B_aSuPJBe29_0(.din(w_dff_B_rJQqSIF11_0),.dout(w_dff_B_aSuPJBe29_0),.clk(gclk));
	jdff dff_B_WIH07Xkj5_0(.din(w_dff_B_aSuPJBe29_0),.dout(w_dff_B_WIH07Xkj5_0),.clk(gclk));
	jdff dff_B_PM8o8nAm7_0(.din(w_dff_B_WIH07Xkj5_0),.dout(w_dff_B_PM8o8nAm7_0),.clk(gclk));
	jdff dff_B_bWTiumqj8_0(.din(w_dff_B_PM8o8nAm7_0),.dout(w_dff_B_bWTiumqj8_0),.clk(gclk));
	jdff dff_B_nXRDLqzk4_0(.din(w_dff_B_bWTiumqj8_0),.dout(w_dff_B_nXRDLqzk4_0),.clk(gclk));
	jdff dff_B_qKmbI41y7_0(.din(w_dff_B_nXRDLqzk4_0),.dout(w_dff_B_qKmbI41y7_0),.clk(gclk));
	jdff dff_B_zr09pa7n1_0(.din(w_dff_B_qKmbI41y7_0),.dout(w_dff_B_zr09pa7n1_0),.clk(gclk));
	jdff dff_B_E4Vg84Lj1_0(.din(w_dff_B_zr09pa7n1_0),.dout(w_dff_B_E4Vg84Lj1_0),.clk(gclk));
	jdff dff_B_ZK5CgouX2_0(.din(w_dff_B_E4Vg84Lj1_0),.dout(w_dff_B_ZK5CgouX2_0),.clk(gclk));
	jdff dff_B_Kygmbtdm2_0(.din(w_dff_B_ZK5CgouX2_0),.dout(w_dff_B_Kygmbtdm2_0),.clk(gclk));
	jdff dff_B_zn43aFR24_0(.din(w_dff_B_Kygmbtdm2_0),.dout(w_dff_B_zn43aFR24_0),.clk(gclk));
	jdff dff_B_lW7n09O32_0(.din(w_dff_B_zn43aFR24_0),.dout(w_dff_B_lW7n09O32_0),.clk(gclk));
	jdff dff_B_mh8cKYwj2_0(.din(w_dff_B_lW7n09O32_0),.dout(w_dff_B_mh8cKYwj2_0),.clk(gclk));
	jdff dff_B_Yxb7eyNY0_0(.din(w_dff_B_mh8cKYwj2_0),.dout(w_dff_B_Yxb7eyNY0_0),.clk(gclk));
	jdff dff_B_i03DsB0k9_0(.din(n1054),.dout(w_dff_B_i03DsB0k9_0),.clk(gclk));
	jdff dff_B_WyresKMq8_0(.din(w_dff_B_i03DsB0k9_0),.dout(w_dff_B_WyresKMq8_0),.clk(gclk));
	jdff dff_B_JKNycuHs1_0(.din(w_dff_B_WyresKMq8_0),.dout(w_dff_B_JKNycuHs1_0),.clk(gclk));
	jdff dff_B_To6n4iMm1_0(.din(w_dff_B_JKNycuHs1_0),.dout(w_dff_B_To6n4iMm1_0),.clk(gclk));
	jdff dff_B_9nB2Bezx5_0(.din(w_dff_B_To6n4iMm1_0),.dout(w_dff_B_9nB2Bezx5_0),.clk(gclk));
	jdff dff_B_KcmTXtoY7_0(.din(w_dff_B_9nB2Bezx5_0),.dout(w_dff_B_KcmTXtoY7_0),.clk(gclk));
	jdff dff_B_ZaQbYrLH4_0(.din(w_dff_B_KcmTXtoY7_0),.dout(w_dff_B_ZaQbYrLH4_0),.clk(gclk));
	jdff dff_B_T6otSM9I4_0(.din(w_dff_B_ZaQbYrLH4_0),.dout(w_dff_B_T6otSM9I4_0),.clk(gclk));
	jdff dff_B_dCkkux5u4_0(.din(w_dff_B_T6otSM9I4_0),.dout(w_dff_B_dCkkux5u4_0),.clk(gclk));
	jdff dff_B_nzw6BVd93_0(.din(w_dff_B_dCkkux5u4_0),.dout(w_dff_B_nzw6BVd93_0),.clk(gclk));
	jdff dff_B_AaXqchK28_0(.din(w_dff_B_nzw6BVd93_0),.dout(w_dff_B_AaXqchK28_0),.clk(gclk));
	jdff dff_B_6cDGnhpg6_0(.din(w_dff_B_AaXqchK28_0),.dout(w_dff_B_6cDGnhpg6_0),.clk(gclk));
	jdff dff_B_bXGxEJQW8_0(.din(w_dff_B_6cDGnhpg6_0),.dout(w_dff_B_bXGxEJQW8_0),.clk(gclk));
	jdff dff_B_wdMnH8Ff5_0(.din(w_dff_B_bXGxEJQW8_0),.dout(w_dff_B_wdMnH8Ff5_0),.clk(gclk));
	jdff dff_B_3iKPHi4K4_0(.din(w_dff_B_wdMnH8Ff5_0),.dout(w_dff_B_3iKPHi4K4_0),.clk(gclk));
	jdff dff_B_FXQ3W1k68_0(.din(w_dff_B_3iKPHi4K4_0),.dout(w_dff_B_FXQ3W1k68_0),.clk(gclk));
	jdff dff_B_GZmZOvaj2_0(.din(w_dff_B_FXQ3W1k68_0),.dout(w_dff_B_GZmZOvaj2_0),.clk(gclk));
	jdff dff_B_RugSlYs21_0(.din(w_dff_B_GZmZOvaj2_0),.dout(w_dff_B_RugSlYs21_0),.clk(gclk));
	jdff dff_B_3vL4qTJL9_0(.din(w_dff_B_RugSlYs21_0),.dout(w_dff_B_3vL4qTJL9_0),.clk(gclk));
	jdff dff_B_N5UCnsYn8_0(.din(w_dff_B_3vL4qTJL9_0),.dout(w_dff_B_N5UCnsYn8_0),.clk(gclk));
	jdff dff_B_JS5nSguM2_0(.din(w_dff_B_N5UCnsYn8_0),.dout(w_dff_B_JS5nSguM2_0),.clk(gclk));
	jdff dff_B_XReSzSqK2_0(.din(w_dff_B_JS5nSguM2_0),.dout(w_dff_B_XReSzSqK2_0),.clk(gclk));
	jdff dff_B_xrc0AWSP3_0(.din(w_dff_B_XReSzSqK2_0),.dout(w_dff_B_xrc0AWSP3_0),.clk(gclk));
	jdff dff_B_EZTMbPfY5_0(.din(w_dff_B_xrc0AWSP3_0),.dout(w_dff_B_EZTMbPfY5_0),.clk(gclk));
	jdff dff_B_NfwtV7ar1_0(.din(w_dff_B_EZTMbPfY5_0),.dout(w_dff_B_NfwtV7ar1_0),.clk(gclk));
	jdff dff_B_U52sDTsA5_0(.din(w_dff_B_NfwtV7ar1_0),.dout(w_dff_B_U52sDTsA5_0),.clk(gclk));
	jdff dff_B_papPhMdP6_0(.din(w_dff_B_U52sDTsA5_0),.dout(w_dff_B_papPhMdP6_0),.clk(gclk));
	jdff dff_B_TdB2oZHS9_0(.din(w_dff_B_papPhMdP6_0),.dout(w_dff_B_TdB2oZHS9_0),.clk(gclk));
	jdff dff_B_jokVzOCq4_0(.din(w_dff_B_TdB2oZHS9_0),.dout(w_dff_B_jokVzOCq4_0),.clk(gclk));
	jdff dff_B_rsrwPn7Q8_0(.din(w_dff_B_jokVzOCq4_0),.dout(w_dff_B_rsrwPn7Q8_0),.clk(gclk));
	jdff dff_B_f7OWNSBZ7_0(.din(w_dff_B_rsrwPn7Q8_0),.dout(w_dff_B_f7OWNSBZ7_0),.clk(gclk));
	jdff dff_B_qb1B3slN1_0(.din(w_dff_B_f7OWNSBZ7_0),.dout(w_dff_B_qb1B3slN1_0),.clk(gclk));
	jdff dff_B_mQ6sCzV03_0(.din(w_dff_B_qb1B3slN1_0),.dout(w_dff_B_mQ6sCzV03_0),.clk(gclk));
	jdff dff_B_swq2P9Ax7_0(.din(w_dff_B_mQ6sCzV03_0),.dout(w_dff_B_swq2P9Ax7_0),.clk(gclk));
	jdff dff_B_ubxnuARn6_0(.din(w_dff_B_swq2P9Ax7_0),.dout(w_dff_B_ubxnuARn6_0),.clk(gclk));
	jdff dff_B_bZTzS0SK2_0(.din(w_dff_B_ubxnuARn6_0),.dout(w_dff_B_bZTzS0SK2_0),.clk(gclk));
	jdff dff_B_HQFZrY3k8_0(.din(w_dff_B_bZTzS0SK2_0),.dout(w_dff_B_HQFZrY3k8_0),.clk(gclk));
	jdff dff_B_amZiA1wi7_0(.din(w_dff_B_HQFZrY3k8_0),.dout(w_dff_B_amZiA1wi7_0),.clk(gclk));
	jdff dff_B_Lhi9rStt0_0(.din(w_dff_B_amZiA1wi7_0),.dout(w_dff_B_Lhi9rStt0_0),.clk(gclk));
	jdff dff_B_KvAc0izF4_0(.din(w_dff_B_Lhi9rStt0_0),.dout(w_dff_B_KvAc0izF4_0),.clk(gclk));
	jdff dff_B_l114WAU63_0(.din(w_dff_B_KvAc0izF4_0),.dout(w_dff_B_l114WAU63_0),.clk(gclk));
	jdff dff_B_IrusQLRo6_0(.din(w_dff_B_l114WAU63_0),.dout(w_dff_B_IrusQLRo6_0),.clk(gclk));
	jdff dff_B_zEafl3z17_0(.din(w_dff_B_IrusQLRo6_0),.dout(w_dff_B_zEafl3z17_0),.clk(gclk));
	jdff dff_B_Ef8Ppp8R5_0(.din(w_dff_B_zEafl3z17_0),.dout(w_dff_B_Ef8Ppp8R5_0),.clk(gclk));
	jdff dff_B_ltokuBCR5_0(.din(w_dff_B_Ef8Ppp8R5_0),.dout(w_dff_B_ltokuBCR5_0),.clk(gclk));
	jdff dff_B_RXaRnNG89_0(.din(w_dff_B_ltokuBCR5_0),.dout(w_dff_B_RXaRnNG89_0),.clk(gclk));
	jdff dff_B_lmXu2mHI5_0(.din(w_dff_B_RXaRnNG89_0),.dout(w_dff_B_lmXu2mHI5_0),.clk(gclk));
	jdff dff_B_fllAp6r39_0(.din(w_dff_B_lmXu2mHI5_0),.dout(w_dff_B_fllAp6r39_0),.clk(gclk));
	jdff dff_B_XhtHh4Cf7_0(.din(w_dff_B_fllAp6r39_0),.dout(w_dff_B_XhtHh4Cf7_0),.clk(gclk));
	jdff dff_B_49LT0sZG0_0(.din(w_dff_B_XhtHh4Cf7_0),.dout(w_dff_B_49LT0sZG0_0),.clk(gclk));
	jdff dff_B_XpAbIZSD0_0(.din(w_dff_B_49LT0sZG0_0),.dout(w_dff_B_XpAbIZSD0_0),.clk(gclk));
	jdff dff_B_Z8IhUQBi1_0(.din(w_dff_B_XpAbIZSD0_0),.dout(w_dff_B_Z8IhUQBi1_0),.clk(gclk));
	jdff dff_B_B74k7I7U6_0(.din(w_dff_B_Z8IhUQBi1_0),.dout(w_dff_B_B74k7I7U6_0),.clk(gclk));
	jdff dff_B_hPdAM3bS5_0(.din(w_dff_B_B74k7I7U6_0),.dout(w_dff_B_hPdAM3bS5_0),.clk(gclk));
	jdff dff_B_zmgDIyvg3_0(.din(w_dff_B_hPdAM3bS5_0),.dout(w_dff_B_zmgDIyvg3_0),.clk(gclk));
	jdff dff_B_xW1z9eYL7_0(.din(w_dff_B_zmgDIyvg3_0),.dout(w_dff_B_xW1z9eYL7_0),.clk(gclk));
	jdff dff_B_R6P5RagF3_0(.din(w_dff_B_xW1z9eYL7_0),.dout(w_dff_B_R6P5RagF3_0),.clk(gclk));
	jdff dff_B_VGb6Ptq23_0(.din(w_dff_B_R6P5RagF3_0),.dout(w_dff_B_VGb6Ptq23_0),.clk(gclk));
	jdff dff_B_47S8cGDP4_0(.din(w_dff_B_VGb6Ptq23_0),.dout(w_dff_B_47S8cGDP4_0),.clk(gclk));
	jdff dff_B_eF1Y3tH79_0(.din(w_dff_B_47S8cGDP4_0),.dout(w_dff_B_eF1Y3tH79_0),.clk(gclk));
	jdff dff_B_8Ib1lwHk3_0(.din(w_dff_B_eF1Y3tH79_0),.dout(w_dff_B_8Ib1lwHk3_0),.clk(gclk));
	jdff dff_B_oWJ2uPW18_0(.din(w_dff_B_8Ib1lwHk3_0),.dout(w_dff_B_oWJ2uPW18_0),.clk(gclk));
	jdff dff_B_WGZrHuMM2_0(.din(w_dff_B_oWJ2uPW18_0),.dout(w_dff_B_WGZrHuMM2_0),.clk(gclk));
	jdff dff_B_Gww81NxQ2_0(.din(w_dff_B_WGZrHuMM2_0),.dout(w_dff_B_Gww81NxQ2_0),.clk(gclk));
	jdff dff_B_z0UvKrVS2_0(.din(w_dff_B_Gww81NxQ2_0),.dout(w_dff_B_z0UvKrVS2_0),.clk(gclk));
	jdff dff_B_OhcBtwwL3_0(.din(w_dff_B_z0UvKrVS2_0),.dout(w_dff_B_OhcBtwwL3_0),.clk(gclk));
	jdff dff_B_mKRHJEaT7_0(.din(w_dff_B_OhcBtwwL3_0),.dout(w_dff_B_mKRHJEaT7_0),.clk(gclk));
	jdff dff_B_fLTydxC90_0(.din(w_dff_B_mKRHJEaT7_0),.dout(w_dff_B_fLTydxC90_0),.clk(gclk));
	jdff dff_B_SOymH8sV5_0(.din(w_dff_B_fLTydxC90_0),.dout(w_dff_B_SOymH8sV5_0),.clk(gclk));
	jdff dff_B_MkJLb7yg8_0(.din(w_dff_B_SOymH8sV5_0),.dout(w_dff_B_MkJLb7yg8_0),.clk(gclk));
	jdff dff_B_1uxv8di55_0(.din(w_dff_B_MkJLb7yg8_0),.dout(w_dff_B_1uxv8di55_0),.clk(gclk));
	jdff dff_B_lcCQC9FS8_0(.din(w_dff_B_1uxv8di55_0),.dout(w_dff_B_lcCQC9FS8_0),.clk(gclk));
	jdff dff_B_ZHC8vifY5_0(.din(w_dff_B_lcCQC9FS8_0),.dout(w_dff_B_ZHC8vifY5_0),.clk(gclk));
	jdff dff_B_3IkOFxUB6_0(.din(w_dff_B_ZHC8vifY5_0),.dout(w_dff_B_3IkOFxUB6_0),.clk(gclk));
	jdff dff_B_ncqogXVe4_0(.din(w_dff_B_3IkOFxUB6_0),.dout(w_dff_B_ncqogXVe4_0),.clk(gclk));
	jdff dff_B_3LCKPhW87_0(.din(w_dff_B_ncqogXVe4_0),.dout(w_dff_B_3LCKPhW87_0),.clk(gclk));
	jdff dff_B_ldADEgEZ5_0(.din(w_dff_B_3LCKPhW87_0),.dout(w_dff_B_ldADEgEZ5_0),.clk(gclk));
	jdff dff_B_Ti0fmlFP6_0(.din(w_dff_B_ldADEgEZ5_0),.dout(w_dff_B_Ti0fmlFP6_0),.clk(gclk));
	jdff dff_B_1EDzcKgC8_0(.din(w_dff_B_Ti0fmlFP6_0),.dout(w_dff_B_1EDzcKgC8_0),.clk(gclk));
	jdff dff_B_YkuWKzVy2_0(.din(w_dff_B_1EDzcKgC8_0),.dout(w_dff_B_YkuWKzVy2_0),.clk(gclk));
	jdff dff_B_Va3GCSV01_0(.din(w_dff_B_YkuWKzVy2_0),.dout(w_dff_B_Va3GCSV01_0),.clk(gclk));
	jdff dff_B_idmhnMSV1_0(.din(w_dff_B_Va3GCSV01_0),.dout(w_dff_B_idmhnMSV1_0),.clk(gclk));
	jdff dff_B_z1JUa0KP3_0(.din(w_dff_B_idmhnMSV1_0),.dout(w_dff_B_z1JUa0KP3_0),.clk(gclk));
	jdff dff_B_bm3uN25j4_0(.din(w_dff_B_z1JUa0KP3_0),.dout(w_dff_B_bm3uN25j4_0),.clk(gclk));
	jdff dff_B_xgu7Fjgx7_0(.din(w_dff_B_bm3uN25j4_0),.dout(w_dff_B_xgu7Fjgx7_0),.clk(gclk));
	jdff dff_B_y8TBpVZY7_0(.din(w_dff_B_xgu7Fjgx7_0),.dout(w_dff_B_y8TBpVZY7_0),.clk(gclk));
	jdff dff_B_5w3PXRDA6_0(.din(w_dff_B_y8TBpVZY7_0),.dout(w_dff_B_5w3PXRDA6_0),.clk(gclk));
	jdff dff_B_FKK7EtMa7_0(.din(w_dff_B_5w3PXRDA6_0),.dout(w_dff_B_FKK7EtMa7_0),.clk(gclk));
	jdff dff_B_tI9tqR8K8_0(.din(w_dff_B_FKK7EtMa7_0),.dout(w_dff_B_tI9tqR8K8_0),.clk(gclk));
	jdff dff_B_1A03e1BA0_0(.din(w_dff_B_tI9tqR8K8_0),.dout(w_dff_B_1A03e1BA0_0),.clk(gclk));
	jdff dff_B_l0vnjnHH8_0(.din(w_dff_B_1A03e1BA0_0),.dout(w_dff_B_l0vnjnHH8_0),.clk(gclk));
	jdff dff_B_o4NfDfSU4_0(.din(w_dff_B_l0vnjnHH8_0),.dout(w_dff_B_o4NfDfSU4_0),.clk(gclk));
	jdff dff_B_toxmDRH98_0(.din(w_dff_B_o4NfDfSU4_0),.dout(w_dff_B_toxmDRH98_0),.clk(gclk));
	jdff dff_B_8NjOG2gv0_0(.din(w_dff_B_toxmDRH98_0),.dout(w_dff_B_8NjOG2gv0_0),.clk(gclk));
	jdff dff_B_mw76b3jb4_0(.din(w_dff_B_8NjOG2gv0_0),.dout(w_dff_B_mw76b3jb4_0),.clk(gclk));
	jdff dff_B_7EhcehT73_0(.din(w_dff_B_mw76b3jb4_0),.dout(w_dff_B_7EhcehT73_0),.clk(gclk));
	jdff dff_B_IEqH6rZa1_0(.din(w_dff_B_7EhcehT73_0),.dout(w_dff_B_IEqH6rZa1_0),.clk(gclk));
	jdff dff_B_seimVXrJ4_0(.din(w_dff_B_IEqH6rZa1_0),.dout(w_dff_B_seimVXrJ4_0),.clk(gclk));
	jdff dff_B_TYRcfwl23_0(.din(w_dff_B_seimVXrJ4_0),.dout(w_dff_B_TYRcfwl23_0),.clk(gclk));
	jdff dff_B_GNfOxe4K6_0(.din(w_dff_B_TYRcfwl23_0),.dout(w_dff_B_GNfOxe4K6_0),.clk(gclk));
	jdff dff_B_ZfYPFTUU8_0(.din(w_dff_B_GNfOxe4K6_0),.dout(w_dff_B_ZfYPFTUU8_0),.clk(gclk));
	jdff dff_B_fYLTMBXi1_0(.din(w_dff_B_ZfYPFTUU8_0),.dout(w_dff_B_fYLTMBXi1_0),.clk(gclk));
	jdff dff_B_29YjHbro9_0(.din(w_dff_B_fYLTMBXi1_0),.dout(w_dff_B_29YjHbro9_0),.clk(gclk));
	jdff dff_B_JIb0ZRqE7_0(.din(w_dff_B_29YjHbro9_0),.dout(w_dff_B_JIb0ZRqE7_0),.clk(gclk));
	jdff dff_B_LyjLC9yF7_0(.din(w_dff_B_JIb0ZRqE7_0),.dout(w_dff_B_LyjLC9yF7_0),.clk(gclk));
	jdff dff_B_coRleIV87_0(.din(w_dff_B_LyjLC9yF7_0),.dout(w_dff_B_coRleIV87_0),.clk(gclk));
	jdff dff_B_1vJFv3ZA9_0(.din(w_dff_B_coRleIV87_0),.dout(w_dff_B_1vJFv3ZA9_0),.clk(gclk));
	jdff dff_B_UoItZ67J8_0(.din(w_dff_B_1vJFv3ZA9_0),.dout(w_dff_B_UoItZ67J8_0),.clk(gclk));
	jdff dff_B_9eDKA3c71_0(.din(w_dff_B_UoItZ67J8_0),.dout(w_dff_B_9eDKA3c71_0),.clk(gclk));
	jdff dff_B_WU8fFmwC2_0(.din(w_dff_B_9eDKA3c71_0),.dout(w_dff_B_WU8fFmwC2_0),.clk(gclk));
	jdff dff_B_hCzyrGpy3_0(.din(w_dff_B_WU8fFmwC2_0),.dout(w_dff_B_hCzyrGpy3_0),.clk(gclk));
	jdff dff_B_N2aM87v43_0(.din(n1060),.dout(w_dff_B_N2aM87v43_0),.clk(gclk));
	jdff dff_B_pYnbF4kV5_0(.din(w_dff_B_N2aM87v43_0),.dout(w_dff_B_pYnbF4kV5_0),.clk(gclk));
	jdff dff_B_dSTR5RCM6_0(.din(w_dff_B_pYnbF4kV5_0),.dout(w_dff_B_dSTR5RCM6_0),.clk(gclk));
	jdff dff_B_FB6kOVCH1_0(.din(w_dff_B_dSTR5RCM6_0),.dout(w_dff_B_FB6kOVCH1_0),.clk(gclk));
	jdff dff_B_GR5pGJRg3_0(.din(w_dff_B_FB6kOVCH1_0),.dout(w_dff_B_GR5pGJRg3_0),.clk(gclk));
	jdff dff_B_Dd0LCtA33_0(.din(w_dff_B_GR5pGJRg3_0),.dout(w_dff_B_Dd0LCtA33_0),.clk(gclk));
	jdff dff_B_4CsqGgUw2_0(.din(w_dff_B_Dd0LCtA33_0),.dout(w_dff_B_4CsqGgUw2_0),.clk(gclk));
	jdff dff_B_RuXI1vk84_0(.din(w_dff_B_4CsqGgUw2_0),.dout(w_dff_B_RuXI1vk84_0),.clk(gclk));
	jdff dff_B_R9eycxBg5_0(.din(w_dff_B_RuXI1vk84_0),.dout(w_dff_B_R9eycxBg5_0),.clk(gclk));
	jdff dff_B_iaVH9DLh4_0(.din(w_dff_B_R9eycxBg5_0),.dout(w_dff_B_iaVH9DLh4_0),.clk(gclk));
	jdff dff_B_W98wexpC1_0(.din(w_dff_B_iaVH9DLh4_0),.dout(w_dff_B_W98wexpC1_0),.clk(gclk));
	jdff dff_B_7OmBOugY1_0(.din(w_dff_B_W98wexpC1_0),.dout(w_dff_B_7OmBOugY1_0),.clk(gclk));
	jdff dff_B_AG6AZ9Nm4_0(.din(w_dff_B_7OmBOugY1_0),.dout(w_dff_B_AG6AZ9Nm4_0),.clk(gclk));
	jdff dff_B_eMKqIWfC0_0(.din(w_dff_B_AG6AZ9Nm4_0),.dout(w_dff_B_eMKqIWfC0_0),.clk(gclk));
	jdff dff_B_0ymKUaxh0_0(.din(w_dff_B_eMKqIWfC0_0),.dout(w_dff_B_0ymKUaxh0_0),.clk(gclk));
	jdff dff_B_7ptmFTMB5_0(.din(w_dff_B_0ymKUaxh0_0),.dout(w_dff_B_7ptmFTMB5_0),.clk(gclk));
	jdff dff_B_5WLAdz2G9_0(.din(w_dff_B_7ptmFTMB5_0),.dout(w_dff_B_5WLAdz2G9_0),.clk(gclk));
	jdff dff_B_lH9PAfsY7_0(.din(w_dff_B_5WLAdz2G9_0),.dout(w_dff_B_lH9PAfsY7_0),.clk(gclk));
	jdff dff_B_iJ9OizwH7_0(.din(w_dff_B_lH9PAfsY7_0),.dout(w_dff_B_iJ9OizwH7_0),.clk(gclk));
	jdff dff_B_uHn64dBX9_0(.din(w_dff_B_iJ9OizwH7_0),.dout(w_dff_B_uHn64dBX9_0),.clk(gclk));
	jdff dff_B_FYjWbd0t8_0(.din(w_dff_B_uHn64dBX9_0),.dout(w_dff_B_FYjWbd0t8_0),.clk(gclk));
	jdff dff_B_fk039VRl4_0(.din(w_dff_B_FYjWbd0t8_0),.dout(w_dff_B_fk039VRl4_0),.clk(gclk));
	jdff dff_B_QN6PEh9G3_0(.din(w_dff_B_fk039VRl4_0),.dout(w_dff_B_QN6PEh9G3_0),.clk(gclk));
	jdff dff_B_NYGLRl3e2_0(.din(w_dff_B_QN6PEh9G3_0),.dout(w_dff_B_NYGLRl3e2_0),.clk(gclk));
	jdff dff_B_M6pBe7jj2_0(.din(w_dff_B_NYGLRl3e2_0),.dout(w_dff_B_M6pBe7jj2_0),.clk(gclk));
	jdff dff_B_WUa0vBEc0_0(.din(w_dff_B_M6pBe7jj2_0),.dout(w_dff_B_WUa0vBEc0_0),.clk(gclk));
	jdff dff_B_mBJ7qwKY5_0(.din(w_dff_B_WUa0vBEc0_0),.dout(w_dff_B_mBJ7qwKY5_0),.clk(gclk));
	jdff dff_B_6DBQ2pi99_0(.din(w_dff_B_mBJ7qwKY5_0),.dout(w_dff_B_6DBQ2pi99_0),.clk(gclk));
	jdff dff_B_8NEJDtKE8_0(.din(w_dff_B_6DBQ2pi99_0),.dout(w_dff_B_8NEJDtKE8_0),.clk(gclk));
	jdff dff_B_KnOqWmjK0_0(.din(w_dff_B_8NEJDtKE8_0),.dout(w_dff_B_KnOqWmjK0_0),.clk(gclk));
	jdff dff_B_6n7COUYF2_0(.din(w_dff_B_KnOqWmjK0_0),.dout(w_dff_B_6n7COUYF2_0),.clk(gclk));
	jdff dff_B_FI0Lsdpt6_0(.din(w_dff_B_6n7COUYF2_0),.dout(w_dff_B_FI0Lsdpt6_0),.clk(gclk));
	jdff dff_B_QWLJXPU56_0(.din(w_dff_B_FI0Lsdpt6_0),.dout(w_dff_B_QWLJXPU56_0),.clk(gclk));
	jdff dff_B_vsx1C2pJ4_0(.din(w_dff_B_QWLJXPU56_0),.dout(w_dff_B_vsx1C2pJ4_0),.clk(gclk));
	jdff dff_B_8tXB6zb78_0(.din(w_dff_B_vsx1C2pJ4_0),.dout(w_dff_B_8tXB6zb78_0),.clk(gclk));
	jdff dff_B_T0nPAzhQ9_0(.din(w_dff_B_8tXB6zb78_0),.dout(w_dff_B_T0nPAzhQ9_0),.clk(gclk));
	jdff dff_B_B2i3kMnG5_0(.din(w_dff_B_T0nPAzhQ9_0),.dout(w_dff_B_B2i3kMnG5_0),.clk(gclk));
	jdff dff_B_dJhWv3XA1_0(.din(w_dff_B_B2i3kMnG5_0),.dout(w_dff_B_dJhWv3XA1_0),.clk(gclk));
	jdff dff_B_KxI36ckE7_0(.din(w_dff_B_dJhWv3XA1_0),.dout(w_dff_B_KxI36ckE7_0),.clk(gclk));
	jdff dff_B_s4iz3U4L5_0(.din(w_dff_B_KxI36ckE7_0),.dout(w_dff_B_s4iz3U4L5_0),.clk(gclk));
	jdff dff_B_OZxBQ9Lg8_0(.din(w_dff_B_s4iz3U4L5_0),.dout(w_dff_B_OZxBQ9Lg8_0),.clk(gclk));
	jdff dff_B_sLqxUbDO1_0(.din(w_dff_B_OZxBQ9Lg8_0),.dout(w_dff_B_sLqxUbDO1_0),.clk(gclk));
	jdff dff_B_JZ1ZxhAg2_0(.din(w_dff_B_sLqxUbDO1_0),.dout(w_dff_B_JZ1ZxhAg2_0),.clk(gclk));
	jdff dff_B_OBtaPguL1_0(.din(w_dff_B_JZ1ZxhAg2_0),.dout(w_dff_B_OBtaPguL1_0),.clk(gclk));
	jdff dff_B_jL7ZsxXN5_0(.din(w_dff_B_OBtaPguL1_0),.dout(w_dff_B_jL7ZsxXN5_0),.clk(gclk));
	jdff dff_B_6ig9KpOO3_0(.din(w_dff_B_jL7ZsxXN5_0),.dout(w_dff_B_6ig9KpOO3_0),.clk(gclk));
	jdff dff_B_bNuv0OMU7_0(.din(w_dff_B_6ig9KpOO3_0),.dout(w_dff_B_bNuv0OMU7_0),.clk(gclk));
	jdff dff_B_WTB1Tm6Y4_0(.din(w_dff_B_bNuv0OMU7_0),.dout(w_dff_B_WTB1Tm6Y4_0),.clk(gclk));
	jdff dff_B_qEcBxoGU2_0(.din(w_dff_B_WTB1Tm6Y4_0),.dout(w_dff_B_qEcBxoGU2_0),.clk(gclk));
	jdff dff_B_uMtu1fbb4_0(.din(w_dff_B_qEcBxoGU2_0),.dout(w_dff_B_uMtu1fbb4_0),.clk(gclk));
	jdff dff_B_UbU53qU97_0(.din(w_dff_B_uMtu1fbb4_0),.dout(w_dff_B_UbU53qU97_0),.clk(gclk));
	jdff dff_B_b7uIGOd70_0(.din(w_dff_B_UbU53qU97_0),.dout(w_dff_B_b7uIGOd70_0),.clk(gclk));
	jdff dff_B_fek6Kjkc8_0(.din(w_dff_B_b7uIGOd70_0),.dout(w_dff_B_fek6Kjkc8_0),.clk(gclk));
	jdff dff_B_QwJVRI1J7_0(.din(w_dff_B_fek6Kjkc8_0),.dout(w_dff_B_QwJVRI1J7_0),.clk(gclk));
	jdff dff_B_OwB2scgS6_0(.din(w_dff_B_QwJVRI1J7_0),.dout(w_dff_B_OwB2scgS6_0),.clk(gclk));
	jdff dff_B_JRmbTlP12_0(.din(w_dff_B_OwB2scgS6_0),.dout(w_dff_B_JRmbTlP12_0),.clk(gclk));
	jdff dff_B_DgPVVtDQ6_0(.din(w_dff_B_JRmbTlP12_0),.dout(w_dff_B_DgPVVtDQ6_0),.clk(gclk));
	jdff dff_B_Nog7bVeE8_0(.din(w_dff_B_DgPVVtDQ6_0),.dout(w_dff_B_Nog7bVeE8_0),.clk(gclk));
	jdff dff_B_1L36KDnF5_0(.din(w_dff_B_Nog7bVeE8_0),.dout(w_dff_B_1L36KDnF5_0),.clk(gclk));
	jdff dff_B_UpAFjjnA5_0(.din(w_dff_B_1L36KDnF5_0),.dout(w_dff_B_UpAFjjnA5_0),.clk(gclk));
	jdff dff_B_Vn54Je6Y0_0(.din(w_dff_B_UpAFjjnA5_0),.dout(w_dff_B_Vn54Je6Y0_0),.clk(gclk));
	jdff dff_B_AcNJ84GQ0_0(.din(w_dff_B_Vn54Je6Y0_0),.dout(w_dff_B_AcNJ84GQ0_0),.clk(gclk));
	jdff dff_B_cOzYuYH38_0(.din(w_dff_B_AcNJ84GQ0_0),.dout(w_dff_B_cOzYuYH38_0),.clk(gclk));
	jdff dff_B_FkT3Rce07_0(.din(w_dff_B_cOzYuYH38_0),.dout(w_dff_B_FkT3Rce07_0),.clk(gclk));
	jdff dff_B_09q1r8kV6_0(.din(w_dff_B_FkT3Rce07_0),.dout(w_dff_B_09q1r8kV6_0),.clk(gclk));
	jdff dff_B_sYCdQLvi8_0(.din(w_dff_B_09q1r8kV6_0),.dout(w_dff_B_sYCdQLvi8_0),.clk(gclk));
	jdff dff_B_GIJFw0J56_0(.din(w_dff_B_sYCdQLvi8_0),.dout(w_dff_B_GIJFw0J56_0),.clk(gclk));
	jdff dff_B_o5ByDST94_0(.din(w_dff_B_GIJFw0J56_0),.dout(w_dff_B_o5ByDST94_0),.clk(gclk));
	jdff dff_B_VudLPSsx4_0(.din(w_dff_B_o5ByDST94_0),.dout(w_dff_B_VudLPSsx4_0),.clk(gclk));
	jdff dff_B_Zi2pPeuQ7_0(.din(w_dff_B_VudLPSsx4_0),.dout(w_dff_B_Zi2pPeuQ7_0),.clk(gclk));
	jdff dff_B_aVh0GrHE4_0(.din(w_dff_B_Zi2pPeuQ7_0),.dout(w_dff_B_aVh0GrHE4_0),.clk(gclk));
	jdff dff_B_nrDSOjCU1_0(.din(w_dff_B_aVh0GrHE4_0),.dout(w_dff_B_nrDSOjCU1_0),.clk(gclk));
	jdff dff_B_kxMPYsLc4_0(.din(w_dff_B_nrDSOjCU1_0),.dout(w_dff_B_kxMPYsLc4_0),.clk(gclk));
	jdff dff_B_u3QFuncY3_0(.din(w_dff_B_kxMPYsLc4_0),.dout(w_dff_B_u3QFuncY3_0),.clk(gclk));
	jdff dff_B_MWhvCoPy3_0(.din(w_dff_B_u3QFuncY3_0),.dout(w_dff_B_MWhvCoPy3_0),.clk(gclk));
	jdff dff_B_CF887ifs5_0(.din(w_dff_B_MWhvCoPy3_0),.dout(w_dff_B_CF887ifs5_0),.clk(gclk));
	jdff dff_B_3OLCiZsM8_0(.din(w_dff_B_CF887ifs5_0),.dout(w_dff_B_3OLCiZsM8_0),.clk(gclk));
	jdff dff_B_lu049csJ5_0(.din(w_dff_B_3OLCiZsM8_0),.dout(w_dff_B_lu049csJ5_0),.clk(gclk));
	jdff dff_B_PDdhCz2h6_0(.din(w_dff_B_lu049csJ5_0),.dout(w_dff_B_PDdhCz2h6_0),.clk(gclk));
	jdff dff_B_yvif2dZq0_0(.din(w_dff_B_PDdhCz2h6_0),.dout(w_dff_B_yvif2dZq0_0),.clk(gclk));
	jdff dff_B_pZbcdhu90_0(.din(w_dff_B_yvif2dZq0_0),.dout(w_dff_B_pZbcdhu90_0),.clk(gclk));
	jdff dff_B_1bi4Tpbs2_0(.din(w_dff_B_pZbcdhu90_0),.dout(w_dff_B_1bi4Tpbs2_0),.clk(gclk));
	jdff dff_B_3UAlUXRr8_0(.din(w_dff_B_1bi4Tpbs2_0),.dout(w_dff_B_3UAlUXRr8_0),.clk(gclk));
	jdff dff_B_lCsWWIAI8_0(.din(w_dff_B_3UAlUXRr8_0),.dout(w_dff_B_lCsWWIAI8_0),.clk(gclk));
	jdff dff_B_hSBtbjYK6_0(.din(w_dff_B_lCsWWIAI8_0),.dout(w_dff_B_hSBtbjYK6_0),.clk(gclk));
	jdff dff_B_CAx6TS4B1_0(.din(w_dff_B_hSBtbjYK6_0),.dout(w_dff_B_CAx6TS4B1_0),.clk(gclk));
	jdff dff_B_agazoS5v6_0(.din(w_dff_B_CAx6TS4B1_0),.dout(w_dff_B_agazoS5v6_0),.clk(gclk));
	jdff dff_B_dd8LGRTQ5_0(.din(w_dff_B_agazoS5v6_0),.dout(w_dff_B_dd8LGRTQ5_0),.clk(gclk));
	jdff dff_B_9vgahaJ52_0(.din(w_dff_B_dd8LGRTQ5_0),.dout(w_dff_B_9vgahaJ52_0),.clk(gclk));
	jdff dff_B_TXxQZrVy5_0(.din(w_dff_B_9vgahaJ52_0),.dout(w_dff_B_TXxQZrVy5_0),.clk(gclk));
	jdff dff_B_piQYU72g2_0(.din(w_dff_B_TXxQZrVy5_0),.dout(w_dff_B_piQYU72g2_0),.clk(gclk));
	jdff dff_B_PzGOo34e2_0(.din(w_dff_B_piQYU72g2_0),.dout(w_dff_B_PzGOo34e2_0),.clk(gclk));
	jdff dff_B_qGzKW0d84_0(.din(w_dff_B_PzGOo34e2_0),.dout(w_dff_B_qGzKW0d84_0),.clk(gclk));
	jdff dff_B_PsTtP93w9_0(.din(w_dff_B_qGzKW0d84_0),.dout(w_dff_B_PsTtP93w9_0),.clk(gclk));
	jdff dff_B_wR1cEirQ8_0(.din(w_dff_B_PsTtP93w9_0),.dout(w_dff_B_wR1cEirQ8_0),.clk(gclk));
	jdff dff_B_7pacKH3a8_0(.din(w_dff_B_wR1cEirQ8_0),.dout(w_dff_B_7pacKH3a8_0),.clk(gclk));
	jdff dff_B_VY5VH9f41_0(.din(w_dff_B_7pacKH3a8_0),.dout(w_dff_B_VY5VH9f41_0),.clk(gclk));
	jdff dff_B_GFPnc5QO4_0(.din(w_dff_B_VY5VH9f41_0),.dout(w_dff_B_GFPnc5QO4_0),.clk(gclk));
	jdff dff_B_0Q3FRUhx5_0(.din(w_dff_B_GFPnc5QO4_0),.dout(w_dff_B_0Q3FRUhx5_0),.clk(gclk));
	jdff dff_B_tOzFoTvX9_0(.din(w_dff_B_0Q3FRUhx5_0),.dout(w_dff_B_tOzFoTvX9_0),.clk(gclk));
	jdff dff_B_VfmXcYWC8_0(.din(w_dff_B_tOzFoTvX9_0),.dout(w_dff_B_VfmXcYWC8_0),.clk(gclk));
	jdff dff_B_UdsshWbY0_0(.din(w_dff_B_VfmXcYWC8_0),.dout(w_dff_B_UdsshWbY0_0),.clk(gclk));
	jdff dff_B_wW5a0vz27_0(.din(w_dff_B_UdsshWbY0_0),.dout(w_dff_B_wW5a0vz27_0),.clk(gclk));
	jdff dff_B_tUgFNM0R2_0(.din(w_dff_B_wW5a0vz27_0),.dout(w_dff_B_tUgFNM0R2_0),.clk(gclk));
	jdff dff_B_F50xyKXc6_0(.din(w_dff_B_tUgFNM0R2_0),.dout(w_dff_B_F50xyKXc6_0),.clk(gclk));
	jdff dff_B_n9kt1zO44_0(.din(w_dff_B_F50xyKXc6_0),.dout(w_dff_B_n9kt1zO44_0),.clk(gclk));
	jdff dff_B_gZCxEFbs8_0(.din(w_dff_B_n9kt1zO44_0),.dout(w_dff_B_gZCxEFbs8_0),.clk(gclk));
	jdff dff_B_qXkXsSem1_0(.din(w_dff_B_gZCxEFbs8_0),.dout(w_dff_B_qXkXsSem1_0),.clk(gclk));
	jdff dff_B_AEFnbmRR7_0(.din(w_dff_B_qXkXsSem1_0),.dout(w_dff_B_AEFnbmRR7_0),.clk(gclk));
	jdff dff_B_JMkSfCVw2_0(.din(w_dff_B_AEFnbmRR7_0),.dout(w_dff_B_JMkSfCVw2_0),.clk(gclk));
	jdff dff_B_iyPTWEUJ8_0(.din(w_dff_B_JMkSfCVw2_0),.dout(w_dff_B_iyPTWEUJ8_0),.clk(gclk));
	jdff dff_B_xwHJtFQ73_0(.din(w_dff_B_iyPTWEUJ8_0),.dout(w_dff_B_xwHJtFQ73_0),.clk(gclk));
	jdff dff_B_T6cy6adT3_0(.din(n1066),.dout(w_dff_B_T6cy6adT3_0),.clk(gclk));
	jdff dff_B_YCOrLBcA4_0(.din(w_dff_B_T6cy6adT3_0),.dout(w_dff_B_YCOrLBcA4_0),.clk(gclk));
	jdff dff_B_8JBrw99v3_0(.din(w_dff_B_YCOrLBcA4_0),.dout(w_dff_B_8JBrw99v3_0),.clk(gclk));
	jdff dff_B_azvmkemw2_0(.din(w_dff_B_8JBrw99v3_0),.dout(w_dff_B_azvmkemw2_0),.clk(gclk));
	jdff dff_B_6qGfsBCE4_0(.din(w_dff_B_azvmkemw2_0),.dout(w_dff_B_6qGfsBCE4_0),.clk(gclk));
	jdff dff_B_k21MNWbT7_0(.din(w_dff_B_6qGfsBCE4_0),.dout(w_dff_B_k21MNWbT7_0),.clk(gclk));
	jdff dff_B_vAXUboMo7_0(.din(w_dff_B_k21MNWbT7_0),.dout(w_dff_B_vAXUboMo7_0),.clk(gclk));
	jdff dff_B_yZCF1dRt3_0(.din(w_dff_B_vAXUboMo7_0),.dout(w_dff_B_yZCF1dRt3_0),.clk(gclk));
	jdff dff_B_wBhNV9VT5_0(.din(w_dff_B_yZCF1dRt3_0),.dout(w_dff_B_wBhNV9VT5_0),.clk(gclk));
	jdff dff_B_Gq2Me05z8_0(.din(w_dff_B_wBhNV9VT5_0),.dout(w_dff_B_Gq2Me05z8_0),.clk(gclk));
	jdff dff_B_264E3Ppg9_0(.din(w_dff_B_Gq2Me05z8_0),.dout(w_dff_B_264E3Ppg9_0),.clk(gclk));
	jdff dff_B_XtQtJtAB7_0(.din(w_dff_B_264E3Ppg9_0),.dout(w_dff_B_XtQtJtAB7_0),.clk(gclk));
	jdff dff_B_QJcDwvRC7_0(.din(w_dff_B_XtQtJtAB7_0),.dout(w_dff_B_QJcDwvRC7_0),.clk(gclk));
	jdff dff_B_aFaLotrb9_0(.din(w_dff_B_QJcDwvRC7_0),.dout(w_dff_B_aFaLotrb9_0),.clk(gclk));
	jdff dff_B_iKLFWyxf5_0(.din(w_dff_B_aFaLotrb9_0),.dout(w_dff_B_iKLFWyxf5_0),.clk(gclk));
	jdff dff_B_CoH9D9UO9_0(.din(w_dff_B_iKLFWyxf5_0),.dout(w_dff_B_CoH9D9UO9_0),.clk(gclk));
	jdff dff_B_O4IoVMVJ8_0(.din(w_dff_B_CoH9D9UO9_0),.dout(w_dff_B_O4IoVMVJ8_0),.clk(gclk));
	jdff dff_B_iYwXAFHP3_0(.din(w_dff_B_O4IoVMVJ8_0),.dout(w_dff_B_iYwXAFHP3_0),.clk(gclk));
	jdff dff_B_DIIOGA3I4_0(.din(w_dff_B_iYwXAFHP3_0),.dout(w_dff_B_DIIOGA3I4_0),.clk(gclk));
	jdff dff_B_C6YddNUb1_0(.din(w_dff_B_DIIOGA3I4_0),.dout(w_dff_B_C6YddNUb1_0),.clk(gclk));
	jdff dff_B_wDJANGWS5_0(.din(w_dff_B_C6YddNUb1_0),.dout(w_dff_B_wDJANGWS5_0),.clk(gclk));
	jdff dff_B_NG9S8L2O4_0(.din(w_dff_B_wDJANGWS5_0),.dout(w_dff_B_NG9S8L2O4_0),.clk(gclk));
	jdff dff_B_K5VE6OX58_0(.din(w_dff_B_NG9S8L2O4_0),.dout(w_dff_B_K5VE6OX58_0),.clk(gclk));
	jdff dff_B_uFWTbJsY4_0(.din(w_dff_B_K5VE6OX58_0),.dout(w_dff_B_uFWTbJsY4_0),.clk(gclk));
	jdff dff_B_u5PZETdo0_0(.din(w_dff_B_uFWTbJsY4_0),.dout(w_dff_B_u5PZETdo0_0),.clk(gclk));
	jdff dff_B_n62NxzBo2_0(.din(w_dff_B_u5PZETdo0_0),.dout(w_dff_B_n62NxzBo2_0),.clk(gclk));
	jdff dff_B_PQuwOxuc2_0(.din(w_dff_B_n62NxzBo2_0),.dout(w_dff_B_PQuwOxuc2_0),.clk(gclk));
	jdff dff_B_aB2r7vXo0_0(.din(w_dff_B_PQuwOxuc2_0),.dout(w_dff_B_aB2r7vXo0_0),.clk(gclk));
	jdff dff_B_d9lEHOo34_0(.din(w_dff_B_aB2r7vXo0_0),.dout(w_dff_B_d9lEHOo34_0),.clk(gclk));
	jdff dff_B_eWEJ0pE03_0(.din(w_dff_B_d9lEHOo34_0),.dout(w_dff_B_eWEJ0pE03_0),.clk(gclk));
	jdff dff_B_SRTtuOkb1_0(.din(w_dff_B_eWEJ0pE03_0),.dout(w_dff_B_SRTtuOkb1_0),.clk(gclk));
	jdff dff_B_u6Kv1OwD1_0(.din(w_dff_B_SRTtuOkb1_0),.dout(w_dff_B_u6Kv1OwD1_0),.clk(gclk));
	jdff dff_B_3eRuT4Cj6_0(.din(w_dff_B_u6Kv1OwD1_0),.dout(w_dff_B_3eRuT4Cj6_0),.clk(gclk));
	jdff dff_B_Q7H5VH3Y7_0(.din(w_dff_B_3eRuT4Cj6_0),.dout(w_dff_B_Q7H5VH3Y7_0),.clk(gclk));
	jdff dff_B_C04OXU6R4_0(.din(w_dff_B_Q7H5VH3Y7_0),.dout(w_dff_B_C04OXU6R4_0),.clk(gclk));
	jdff dff_B_aCBPNTXZ4_0(.din(w_dff_B_C04OXU6R4_0),.dout(w_dff_B_aCBPNTXZ4_0),.clk(gclk));
	jdff dff_B_syBLDzeQ2_0(.din(w_dff_B_aCBPNTXZ4_0),.dout(w_dff_B_syBLDzeQ2_0),.clk(gclk));
	jdff dff_B_KdrNcJEW5_0(.din(w_dff_B_syBLDzeQ2_0),.dout(w_dff_B_KdrNcJEW5_0),.clk(gclk));
	jdff dff_B_YAiZB8iQ9_0(.din(w_dff_B_KdrNcJEW5_0),.dout(w_dff_B_YAiZB8iQ9_0),.clk(gclk));
	jdff dff_B_DaitgYX06_0(.din(w_dff_B_YAiZB8iQ9_0),.dout(w_dff_B_DaitgYX06_0),.clk(gclk));
	jdff dff_B_xsNgiLEd8_0(.din(w_dff_B_DaitgYX06_0),.dout(w_dff_B_xsNgiLEd8_0),.clk(gclk));
	jdff dff_B_qETm5rru0_0(.din(w_dff_B_xsNgiLEd8_0),.dout(w_dff_B_qETm5rru0_0),.clk(gclk));
	jdff dff_B_BGECBSbQ1_0(.din(w_dff_B_qETm5rru0_0),.dout(w_dff_B_BGECBSbQ1_0),.clk(gclk));
	jdff dff_B_NYC5UaPH9_0(.din(w_dff_B_BGECBSbQ1_0),.dout(w_dff_B_NYC5UaPH9_0),.clk(gclk));
	jdff dff_B_7Wv9h8JE6_0(.din(w_dff_B_NYC5UaPH9_0),.dout(w_dff_B_7Wv9h8JE6_0),.clk(gclk));
	jdff dff_B_2avyXCgM7_0(.din(w_dff_B_7Wv9h8JE6_0),.dout(w_dff_B_2avyXCgM7_0),.clk(gclk));
	jdff dff_B_6TgpZSP71_0(.din(w_dff_B_2avyXCgM7_0),.dout(w_dff_B_6TgpZSP71_0),.clk(gclk));
	jdff dff_B_urBmP0Nt8_0(.din(w_dff_B_6TgpZSP71_0),.dout(w_dff_B_urBmP0Nt8_0),.clk(gclk));
	jdff dff_B_KEEgq3Bz0_0(.din(w_dff_B_urBmP0Nt8_0),.dout(w_dff_B_KEEgq3Bz0_0),.clk(gclk));
	jdff dff_B_Bi0EReY61_0(.din(w_dff_B_KEEgq3Bz0_0),.dout(w_dff_B_Bi0EReY61_0),.clk(gclk));
	jdff dff_B_juAbyvRb9_0(.din(w_dff_B_Bi0EReY61_0),.dout(w_dff_B_juAbyvRb9_0),.clk(gclk));
	jdff dff_B_d4AZS7cc9_0(.din(w_dff_B_juAbyvRb9_0),.dout(w_dff_B_d4AZS7cc9_0),.clk(gclk));
	jdff dff_B_jsZ7rHLO3_0(.din(w_dff_B_d4AZS7cc9_0),.dout(w_dff_B_jsZ7rHLO3_0),.clk(gclk));
	jdff dff_B_whb7k4OF9_0(.din(w_dff_B_jsZ7rHLO3_0),.dout(w_dff_B_whb7k4OF9_0),.clk(gclk));
	jdff dff_B_HsobfZOH9_0(.din(w_dff_B_whb7k4OF9_0),.dout(w_dff_B_HsobfZOH9_0),.clk(gclk));
	jdff dff_B_CxH25B2D8_0(.din(w_dff_B_HsobfZOH9_0),.dout(w_dff_B_CxH25B2D8_0),.clk(gclk));
	jdff dff_B_z7sBEGJ62_0(.din(w_dff_B_CxH25B2D8_0),.dout(w_dff_B_z7sBEGJ62_0),.clk(gclk));
	jdff dff_B_hiOdseny2_0(.din(w_dff_B_z7sBEGJ62_0),.dout(w_dff_B_hiOdseny2_0),.clk(gclk));
	jdff dff_B_DZxoEhGy1_0(.din(w_dff_B_hiOdseny2_0),.dout(w_dff_B_DZxoEhGy1_0),.clk(gclk));
	jdff dff_B_3bixYwa48_0(.din(w_dff_B_DZxoEhGy1_0),.dout(w_dff_B_3bixYwa48_0),.clk(gclk));
	jdff dff_B_YOIBaXK64_0(.din(w_dff_B_3bixYwa48_0),.dout(w_dff_B_YOIBaXK64_0),.clk(gclk));
	jdff dff_B_rSqV4Ts16_0(.din(w_dff_B_YOIBaXK64_0),.dout(w_dff_B_rSqV4Ts16_0),.clk(gclk));
	jdff dff_B_3QdofVOX3_0(.din(w_dff_B_rSqV4Ts16_0),.dout(w_dff_B_3QdofVOX3_0),.clk(gclk));
	jdff dff_B_Vm9xGCX25_0(.din(w_dff_B_3QdofVOX3_0),.dout(w_dff_B_Vm9xGCX25_0),.clk(gclk));
	jdff dff_B_kuRuPFmE9_0(.din(w_dff_B_Vm9xGCX25_0),.dout(w_dff_B_kuRuPFmE9_0),.clk(gclk));
	jdff dff_B_k7ztCerr2_0(.din(w_dff_B_kuRuPFmE9_0),.dout(w_dff_B_k7ztCerr2_0),.clk(gclk));
	jdff dff_B_mR9z6GsX2_0(.din(w_dff_B_k7ztCerr2_0),.dout(w_dff_B_mR9z6GsX2_0),.clk(gclk));
	jdff dff_B_2MRfOOKE0_0(.din(w_dff_B_mR9z6GsX2_0),.dout(w_dff_B_2MRfOOKE0_0),.clk(gclk));
	jdff dff_B_DtUckFku0_0(.din(w_dff_B_2MRfOOKE0_0),.dout(w_dff_B_DtUckFku0_0),.clk(gclk));
	jdff dff_B_06xO03r36_0(.din(w_dff_B_DtUckFku0_0),.dout(w_dff_B_06xO03r36_0),.clk(gclk));
	jdff dff_B_LDcoyRPN9_0(.din(w_dff_B_06xO03r36_0),.dout(w_dff_B_LDcoyRPN9_0),.clk(gclk));
	jdff dff_B_ZsBkbrrA7_0(.din(w_dff_B_LDcoyRPN9_0),.dout(w_dff_B_ZsBkbrrA7_0),.clk(gclk));
	jdff dff_B_6PSJnfqR9_0(.din(w_dff_B_ZsBkbrrA7_0),.dout(w_dff_B_6PSJnfqR9_0),.clk(gclk));
	jdff dff_B_e1vuhETi1_0(.din(w_dff_B_6PSJnfqR9_0),.dout(w_dff_B_e1vuhETi1_0),.clk(gclk));
	jdff dff_B_22inKnNB2_0(.din(w_dff_B_e1vuhETi1_0),.dout(w_dff_B_22inKnNB2_0),.clk(gclk));
	jdff dff_B_1Zjtsvsj7_0(.din(w_dff_B_22inKnNB2_0),.dout(w_dff_B_1Zjtsvsj7_0),.clk(gclk));
	jdff dff_B_2g7v0kq88_0(.din(w_dff_B_1Zjtsvsj7_0),.dout(w_dff_B_2g7v0kq88_0),.clk(gclk));
	jdff dff_B_dt23Tw214_0(.din(w_dff_B_2g7v0kq88_0),.dout(w_dff_B_dt23Tw214_0),.clk(gclk));
	jdff dff_B_douDrV062_0(.din(w_dff_B_dt23Tw214_0),.dout(w_dff_B_douDrV062_0),.clk(gclk));
	jdff dff_B_bJA65jY69_0(.din(w_dff_B_douDrV062_0),.dout(w_dff_B_bJA65jY69_0),.clk(gclk));
	jdff dff_B_BocNrqby2_0(.din(w_dff_B_bJA65jY69_0),.dout(w_dff_B_BocNrqby2_0),.clk(gclk));
	jdff dff_B_4rdZMJyE1_0(.din(w_dff_B_BocNrqby2_0),.dout(w_dff_B_4rdZMJyE1_0),.clk(gclk));
	jdff dff_B_1MDfjnGS8_0(.din(w_dff_B_4rdZMJyE1_0),.dout(w_dff_B_1MDfjnGS8_0),.clk(gclk));
	jdff dff_B_19uc25ty4_0(.din(w_dff_B_1MDfjnGS8_0),.dout(w_dff_B_19uc25ty4_0),.clk(gclk));
	jdff dff_B_2sI8qR5D5_0(.din(w_dff_B_19uc25ty4_0),.dout(w_dff_B_2sI8qR5D5_0),.clk(gclk));
	jdff dff_B_iW29RgG02_0(.din(w_dff_B_2sI8qR5D5_0),.dout(w_dff_B_iW29RgG02_0),.clk(gclk));
	jdff dff_B_E0jSOTne1_0(.din(w_dff_B_iW29RgG02_0),.dout(w_dff_B_E0jSOTne1_0),.clk(gclk));
	jdff dff_B_b2KFkNXt6_0(.din(w_dff_B_E0jSOTne1_0),.dout(w_dff_B_b2KFkNXt6_0),.clk(gclk));
	jdff dff_B_3Gq8fW909_0(.din(w_dff_B_b2KFkNXt6_0),.dout(w_dff_B_3Gq8fW909_0),.clk(gclk));
	jdff dff_B_3PMSX4V41_0(.din(w_dff_B_3Gq8fW909_0),.dout(w_dff_B_3PMSX4V41_0),.clk(gclk));
	jdff dff_B_dDmiZuzD1_0(.din(w_dff_B_3PMSX4V41_0),.dout(w_dff_B_dDmiZuzD1_0),.clk(gclk));
	jdff dff_B_lKZf2caW0_0(.din(w_dff_B_dDmiZuzD1_0),.dout(w_dff_B_lKZf2caW0_0),.clk(gclk));
	jdff dff_B_SDlL0hdy8_0(.din(w_dff_B_lKZf2caW0_0),.dout(w_dff_B_SDlL0hdy8_0),.clk(gclk));
	jdff dff_B_e6Ujrzvl3_0(.din(w_dff_B_SDlL0hdy8_0),.dout(w_dff_B_e6Ujrzvl3_0),.clk(gclk));
	jdff dff_B_FrcdP5mw2_0(.din(w_dff_B_e6Ujrzvl3_0),.dout(w_dff_B_FrcdP5mw2_0),.clk(gclk));
	jdff dff_B_pDfIcIct4_0(.din(w_dff_B_FrcdP5mw2_0),.dout(w_dff_B_pDfIcIct4_0),.clk(gclk));
	jdff dff_B_qvz13JqE2_0(.din(w_dff_B_pDfIcIct4_0),.dout(w_dff_B_qvz13JqE2_0),.clk(gclk));
	jdff dff_B_iBqUaBqm5_0(.din(w_dff_B_qvz13JqE2_0),.dout(w_dff_B_iBqUaBqm5_0),.clk(gclk));
	jdff dff_B_DXCiLBRE0_0(.din(w_dff_B_iBqUaBqm5_0),.dout(w_dff_B_DXCiLBRE0_0),.clk(gclk));
	jdff dff_B_Iqv9HwlC3_0(.din(w_dff_B_DXCiLBRE0_0),.dout(w_dff_B_Iqv9HwlC3_0),.clk(gclk));
	jdff dff_B_bD4khmYF5_0(.din(w_dff_B_Iqv9HwlC3_0),.dout(w_dff_B_bD4khmYF5_0),.clk(gclk));
	jdff dff_B_5XukiGgD6_0(.din(w_dff_B_bD4khmYF5_0),.dout(w_dff_B_5XukiGgD6_0),.clk(gclk));
	jdff dff_B_1acq1Ii29_0(.din(w_dff_B_5XukiGgD6_0),.dout(w_dff_B_1acq1Ii29_0),.clk(gclk));
	jdff dff_B_4xevaueD6_0(.din(w_dff_B_1acq1Ii29_0),.dout(w_dff_B_4xevaueD6_0),.clk(gclk));
	jdff dff_B_Hx4PsOQz5_0(.din(w_dff_B_4xevaueD6_0),.dout(w_dff_B_Hx4PsOQz5_0),.clk(gclk));
	jdff dff_B_mIiTho5V0_0(.din(w_dff_B_Hx4PsOQz5_0),.dout(w_dff_B_mIiTho5V0_0),.clk(gclk));
	jdff dff_B_P2vsFb309_0(.din(w_dff_B_mIiTho5V0_0),.dout(w_dff_B_P2vsFb309_0),.clk(gclk));
	jdff dff_B_LXkLR1Fr3_0(.din(w_dff_B_P2vsFb309_0),.dout(w_dff_B_LXkLR1Fr3_0),.clk(gclk));
	jdff dff_B_sW7lNcSW5_0(.din(w_dff_B_LXkLR1Fr3_0),.dout(w_dff_B_sW7lNcSW5_0),.clk(gclk));
	jdff dff_B_xHzgBnZg4_0(.din(w_dff_B_sW7lNcSW5_0),.dout(w_dff_B_xHzgBnZg4_0),.clk(gclk));
	jdff dff_B_JpTlCLDr0_0(.din(w_dff_B_xHzgBnZg4_0),.dout(w_dff_B_JpTlCLDr0_0),.clk(gclk));
	jdff dff_B_9E4Kjc1o2_0(.din(w_dff_B_JpTlCLDr0_0),.dout(w_dff_B_9E4Kjc1o2_0),.clk(gclk));
	jdff dff_B_qONrkGfY1_0(.din(w_dff_B_9E4Kjc1o2_0),.dout(w_dff_B_qONrkGfY1_0),.clk(gclk));
	jdff dff_B_I0TawrUE3_0(.din(n1072),.dout(w_dff_B_I0TawrUE3_0),.clk(gclk));
	jdff dff_B_vDHofyhm0_0(.din(w_dff_B_I0TawrUE3_0),.dout(w_dff_B_vDHofyhm0_0),.clk(gclk));
	jdff dff_B_c7yZhhEO9_0(.din(w_dff_B_vDHofyhm0_0),.dout(w_dff_B_c7yZhhEO9_0),.clk(gclk));
	jdff dff_B_WuYUn96Y9_0(.din(w_dff_B_c7yZhhEO9_0),.dout(w_dff_B_WuYUn96Y9_0),.clk(gclk));
	jdff dff_B_Ol7JlfiZ4_0(.din(w_dff_B_WuYUn96Y9_0),.dout(w_dff_B_Ol7JlfiZ4_0),.clk(gclk));
	jdff dff_B_wSqtQmgq7_0(.din(w_dff_B_Ol7JlfiZ4_0),.dout(w_dff_B_wSqtQmgq7_0),.clk(gclk));
	jdff dff_B_bRCbm9Rl7_0(.din(w_dff_B_wSqtQmgq7_0),.dout(w_dff_B_bRCbm9Rl7_0),.clk(gclk));
	jdff dff_B_R8zKQYmx3_0(.din(w_dff_B_bRCbm9Rl7_0),.dout(w_dff_B_R8zKQYmx3_0),.clk(gclk));
	jdff dff_B_9bi76dWM7_0(.din(w_dff_B_R8zKQYmx3_0),.dout(w_dff_B_9bi76dWM7_0),.clk(gclk));
	jdff dff_B_NhSMTdg49_0(.din(w_dff_B_9bi76dWM7_0),.dout(w_dff_B_NhSMTdg49_0),.clk(gclk));
	jdff dff_B_ETzjzWvT0_0(.din(w_dff_B_NhSMTdg49_0),.dout(w_dff_B_ETzjzWvT0_0),.clk(gclk));
	jdff dff_B_wXohqQjK0_0(.din(w_dff_B_ETzjzWvT0_0),.dout(w_dff_B_wXohqQjK0_0),.clk(gclk));
	jdff dff_B_fNxdkUYc6_0(.din(w_dff_B_wXohqQjK0_0),.dout(w_dff_B_fNxdkUYc6_0),.clk(gclk));
	jdff dff_B_dplX0Cxl5_0(.din(w_dff_B_fNxdkUYc6_0),.dout(w_dff_B_dplX0Cxl5_0),.clk(gclk));
	jdff dff_B_TQvxEiMA4_0(.din(w_dff_B_dplX0Cxl5_0),.dout(w_dff_B_TQvxEiMA4_0),.clk(gclk));
	jdff dff_B_KL5N6nit9_0(.din(w_dff_B_TQvxEiMA4_0),.dout(w_dff_B_KL5N6nit9_0),.clk(gclk));
	jdff dff_B_wh4smQiZ2_0(.din(w_dff_B_KL5N6nit9_0),.dout(w_dff_B_wh4smQiZ2_0),.clk(gclk));
	jdff dff_B_tfZwkC5h7_0(.din(w_dff_B_wh4smQiZ2_0),.dout(w_dff_B_tfZwkC5h7_0),.clk(gclk));
	jdff dff_B_FDkpAuuP3_0(.din(w_dff_B_tfZwkC5h7_0),.dout(w_dff_B_FDkpAuuP3_0),.clk(gclk));
	jdff dff_B_CJRtQWYe7_0(.din(w_dff_B_FDkpAuuP3_0),.dout(w_dff_B_CJRtQWYe7_0),.clk(gclk));
	jdff dff_B_pDIF9pf89_0(.din(w_dff_B_CJRtQWYe7_0),.dout(w_dff_B_pDIF9pf89_0),.clk(gclk));
	jdff dff_B_oxDHxBc66_0(.din(w_dff_B_pDIF9pf89_0),.dout(w_dff_B_oxDHxBc66_0),.clk(gclk));
	jdff dff_B_Gq7t7FSN6_0(.din(w_dff_B_oxDHxBc66_0),.dout(w_dff_B_Gq7t7FSN6_0),.clk(gclk));
	jdff dff_B_YiUz0Nwb5_0(.din(w_dff_B_Gq7t7FSN6_0),.dout(w_dff_B_YiUz0Nwb5_0),.clk(gclk));
	jdff dff_B_18Xtw7Oy7_0(.din(w_dff_B_YiUz0Nwb5_0),.dout(w_dff_B_18Xtw7Oy7_0),.clk(gclk));
	jdff dff_B_E9kwQgXP9_0(.din(w_dff_B_18Xtw7Oy7_0),.dout(w_dff_B_E9kwQgXP9_0),.clk(gclk));
	jdff dff_B_RerU6hJo4_0(.din(w_dff_B_E9kwQgXP9_0),.dout(w_dff_B_RerU6hJo4_0),.clk(gclk));
	jdff dff_B_rl6MY5LG7_0(.din(w_dff_B_RerU6hJo4_0),.dout(w_dff_B_rl6MY5LG7_0),.clk(gclk));
	jdff dff_B_QEFc5zrY0_0(.din(w_dff_B_rl6MY5LG7_0),.dout(w_dff_B_QEFc5zrY0_0),.clk(gclk));
	jdff dff_B_JEUHMBWj4_0(.din(w_dff_B_QEFc5zrY0_0),.dout(w_dff_B_JEUHMBWj4_0),.clk(gclk));
	jdff dff_B_BsBwoum93_0(.din(w_dff_B_JEUHMBWj4_0),.dout(w_dff_B_BsBwoum93_0),.clk(gclk));
	jdff dff_B_lw6RVVWI9_0(.din(w_dff_B_BsBwoum93_0),.dout(w_dff_B_lw6RVVWI9_0),.clk(gclk));
	jdff dff_B_cHt50svL9_0(.din(w_dff_B_lw6RVVWI9_0),.dout(w_dff_B_cHt50svL9_0),.clk(gclk));
	jdff dff_B_1iwoqoe52_0(.din(w_dff_B_cHt50svL9_0),.dout(w_dff_B_1iwoqoe52_0),.clk(gclk));
	jdff dff_B_77W1sNdN3_0(.din(w_dff_B_1iwoqoe52_0),.dout(w_dff_B_77W1sNdN3_0),.clk(gclk));
	jdff dff_B_VK2ZOAJp7_0(.din(w_dff_B_77W1sNdN3_0),.dout(w_dff_B_VK2ZOAJp7_0),.clk(gclk));
	jdff dff_B_GLVqlhWB9_0(.din(w_dff_B_VK2ZOAJp7_0),.dout(w_dff_B_GLVqlhWB9_0),.clk(gclk));
	jdff dff_B_DCvC2j9c7_0(.din(w_dff_B_GLVqlhWB9_0),.dout(w_dff_B_DCvC2j9c7_0),.clk(gclk));
	jdff dff_B_bPIzqSKU1_0(.din(w_dff_B_DCvC2j9c7_0),.dout(w_dff_B_bPIzqSKU1_0),.clk(gclk));
	jdff dff_B_bkk4KhS27_0(.din(w_dff_B_bPIzqSKU1_0),.dout(w_dff_B_bkk4KhS27_0),.clk(gclk));
	jdff dff_B_MHxfriwQ6_0(.din(w_dff_B_bkk4KhS27_0),.dout(w_dff_B_MHxfriwQ6_0),.clk(gclk));
	jdff dff_B_hwvyEvxS0_0(.din(w_dff_B_MHxfriwQ6_0),.dout(w_dff_B_hwvyEvxS0_0),.clk(gclk));
	jdff dff_B_kyP5gtgY7_0(.din(w_dff_B_hwvyEvxS0_0),.dout(w_dff_B_kyP5gtgY7_0),.clk(gclk));
	jdff dff_B_HStEtvYq3_0(.din(w_dff_B_kyP5gtgY7_0),.dout(w_dff_B_HStEtvYq3_0),.clk(gclk));
	jdff dff_B_Do2DXFxA7_0(.din(w_dff_B_HStEtvYq3_0),.dout(w_dff_B_Do2DXFxA7_0),.clk(gclk));
	jdff dff_B_XfvIiYZg2_0(.din(w_dff_B_Do2DXFxA7_0),.dout(w_dff_B_XfvIiYZg2_0),.clk(gclk));
	jdff dff_B_0oGe2geI1_0(.din(w_dff_B_XfvIiYZg2_0),.dout(w_dff_B_0oGe2geI1_0),.clk(gclk));
	jdff dff_B_qyJML38p0_0(.din(w_dff_B_0oGe2geI1_0),.dout(w_dff_B_qyJML38p0_0),.clk(gclk));
	jdff dff_B_CPPLd22G2_0(.din(w_dff_B_qyJML38p0_0),.dout(w_dff_B_CPPLd22G2_0),.clk(gclk));
	jdff dff_B_I7DcFExr6_0(.din(w_dff_B_CPPLd22G2_0),.dout(w_dff_B_I7DcFExr6_0),.clk(gclk));
	jdff dff_B_pQxhO0z48_0(.din(w_dff_B_I7DcFExr6_0),.dout(w_dff_B_pQxhO0z48_0),.clk(gclk));
	jdff dff_B_o7KTXB8A8_0(.din(w_dff_B_pQxhO0z48_0),.dout(w_dff_B_o7KTXB8A8_0),.clk(gclk));
	jdff dff_B_QSbUKSIM0_0(.din(w_dff_B_o7KTXB8A8_0),.dout(w_dff_B_QSbUKSIM0_0),.clk(gclk));
	jdff dff_B_suCkceyA8_0(.din(w_dff_B_QSbUKSIM0_0),.dout(w_dff_B_suCkceyA8_0),.clk(gclk));
	jdff dff_B_m0wmeRoQ7_0(.din(w_dff_B_suCkceyA8_0),.dout(w_dff_B_m0wmeRoQ7_0),.clk(gclk));
	jdff dff_B_eMtMOVyO5_0(.din(w_dff_B_m0wmeRoQ7_0),.dout(w_dff_B_eMtMOVyO5_0),.clk(gclk));
	jdff dff_B_oWayQWxz7_0(.din(w_dff_B_eMtMOVyO5_0),.dout(w_dff_B_oWayQWxz7_0),.clk(gclk));
	jdff dff_B_XuEhrRXj2_0(.din(w_dff_B_oWayQWxz7_0),.dout(w_dff_B_XuEhrRXj2_0),.clk(gclk));
	jdff dff_B_P3abaly04_0(.din(w_dff_B_XuEhrRXj2_0),.dout(w_dff_B_P3abaly04_0),.clk(gclk));
	jdff dff_B_4oLwDK1c6_0(.din(w_dff_B_P3abaly04_0),.dout(w_dff_B_4oLwDK1c6_0),.clk(gclk));
	jdff dff_B_KRMzZgX74_0(.din(w_dff_B_4oLwDK1c6_0),.dout(w_dff_B_KRMzZgX74_0),.clk(gclk));
	jdff dff_B_tKtF7Wnt0_0(.din(w_dff_B_KRMzZgX74_0),.dout(w_dff_B_tKtF7Wnt0_0),.clk(gclk));
	jdff dff_B_iaUguIy35_0(.din(w_dff_B_tKtF7Wnt0_0),.dout(w_dff_B_iaUguIy35_0),.clk(gclk));
	jdff dff_B_5vyJka1y5_0(.din(w_dff_B_iaUguIy35_0),.dout(w_dff_B_5vyJka1y5_0),.clk(gclk));
	jdff dff_B_SncPSBPK3_0(.din(w_dff_B_5vyJka1y5_0),.dout(w_dff_B_SncPSBPK3_0),.clk(gclk));
	jdff dff_B_JCIUJa659_0(.din(w_dff_B_SncPSBPK3_0),.dout(w_dff_B_JCIUJa659_0),.clk(gclk));
	jdff dff_B_dW1k918b6_0(.din(w_dff_B_JCIUJa659_0),.dout(w_dff_B_dW1k918b6_0),.clk(gclk));
	jdff dff_B_ZCdyyF1Z7_0(.din(w_dff_B_dW1k918b6_0),.dout(w_dff_B_ZCdyyF1Z7_0),.clk(gclk));
	jdff dff_B_xUnVWRlw9_0(.din(w_dff_B_ZCdyyF1Z7_0),.dout(w_dff_B_xUnVWRlw9_0),.clk(gclk));
	jdff dff_B_ZmM808xo9_0(.din(w_dff_B_xUnVWRlw9_0),.dout(w_dff_B_ZmM808xo9_0),.clk(gclk));
	jdff dff_B_4Se8GE2H7_0(.din(w_dff_B_ZmM808xo9_0),.dout(w_dff_B_4Se8GE2H7_0),.clk(gclk));
	jdff dff_B_K4evWBVk3_0(.din(w_dff_B_4Se8GE2H7_0),.dout(w_dff_B_K4evWBVk3_0),.clk(gclk));
	jdff dff_B_tGfKGrvW6_0(.din(w_dff_B_K4evWBVk3_0),.dout(w_dff_B_tGfKGrvW6_0),.clk(gclk));
	jdff dff_B_xO6IeWhE7_0(.din(w_dff_B_tGfKGrvW6_0),.dout(w_dff_B_xO6IeWhE7_0),.clk(gclk));
	jdff dff_B_hMzYzdHY2_0(.din(w_dff_B_xO6IeWhE7_0),.dout(w_dff_B_hMzYzdHY2_0),.clk(gclk));
	jdff dff_B_9CZ7M2z41_0(.din(w_dff_B_hMzYzdHY2_0),.dout(w_dff_B_9CZ7M2z41_0),.clk(gclk));
	jdff dff_B_5PSKn6904_0(.din(w_dff_B_9CZ7M2z41_0),.dout(w_dff_B_5PSKn6904_0),.clk(gclk));
	jdff dff_B_yX6ftvJC7_0(.din(w_dff_B_5PSKn6904_0),.dout(w_dff_B_yX6ftvJC7_0),.clk(gclk));
	jdff dff_B_oasAignb1_0(.din(w_dff_B_yX6ftvJC7_0),.dout(w_dff_B_oasAignb1_0),.clk(gclk));
	jdff dff_B_GJMisELy4_0(.din(w_dff_B_oasAignb1_0),.dout(w_dff_B_GJMisELy4_0),.clk(gclk));
	jdff dff_B_LPmTurw50_0(.din(w_dff_B_GJMisELy4_0),.dout(w_dff_B_LPmTurw50_0),.clk(gclk));
	jdff dff_B_u6aglghB9_0(.din(w_dff_B_LPmTurw50_0),.dout(w_dff_B_u6aglghB9_0),.clk(gclk));
	jdff dff_B_VjkLqvdk3_0(.din(w_dff_B_u6aglghB9_0),.dout(w_dff_B_VjkLqvdk3_0),.clk(gclk));
	jdff dff_B_VlXGF5s78_0(.din(w_dff_B_VjkLqvdk3_0),.dout(w_dff_B_VlXGF5s78_0),.clk(gclk));
	jdff dff_B_MHLMp1re6_0(.din(w_dff_B_VlXGF5s78_0),.dout(w_dff_B_MHLMp1re6_0),.clk(gclk));
	jdff dff_B_d4bCQ6kf9_0(.din(w_dff_B_MHLMp1re6_0),.dout(w_dff_B_d4bCQ6kf9_0),.clk(gclk));
	jdff dff_B_RVIQ57f00_0(.din(w_dff_B_d4bCQ6kf9_0),.dout(w_dff_B_RVIQ57f00_0),.clk(gclk));
	jdff dff_B_xFHBGtJE6_0(.din(w_dff_B_RVIQ57f00_0),.dout(w_dff_B_xFHBGtJE6_0),.clk(gclk));
	jdff dff_B_JTUR309x7_0(.din(w_dff_B_xFHBGtJE6_0),.dout(w_dff_B_JTUR309x7_0),.clk(gclk));
	jdff dff_B_P52kOmzq7_0(.din(w_dff_B_JTUR309x7_0),.dout(w_dff_B_P52kOmzq7_0),.clk(gclk));
	jdff dff_B_7oXEJaj02_0(.din(w_dff_B_P52kOmzq7_0),.dout(w_dff_B_7oXEJaj02_0),.clk(gclk));
	jdff dff_B_Dk9FjoTE4_0(.din(w_dff_B_7oXEJaj02_0),.dout(w_dff_B_Dk9FjoTE4_0),.clk(gclk));
	jdff dff_B_Et4U5xZw0_0(.din(w_dff_B_Dk9FjoTE4_0),.dout(w_dff_B_Et4U5xZw0_0),.clk(gclk));
	jdff dff_B_C5dV5OGy2_0(.din(w_dff_B_Et4U5xZw0_0),.dout(w_dff_B_C5dV5OGy2_0),.clk(gclk));
	jdff dff_B_RTjt4pGP6_0(.din(w_dff_B_C5dV5OGy2_0),.dout(w_dff_B_RTjt4pGP6_0),.clk(gclk));
	jdff dff_B_46EfvZkW0_0(.din(w_dff_B_RTjt4pGP6_0),.dout(w_dff_B_46EfvZkW0_0),.clk(gclk));
	jdff dff_B_BPGfvcvo7_0(.din(w_dff_B_46EfvZkW0_0),.dout(w_dff_B_BPGfvcvo7_0),.clk(gclk));
	jdff dff_B_pIByHgSw4_0(.din(w_dff_B_BPGfvcvo7_0),.dout(w_dff_B_pIByHgSw4_0),.clk(gclk));
	jdff dff_B_NeBzaGqv9_0(.din(w_dff_B_pIByHgSw4_0),.dout(w_dff_B_NeBzaGqv9_0),.clk(gclk));
	jdff dff_B_RM4VGVsv5_0(.din(w_dff_B_NeBzaGqv9_0),.dout(w_dff_B_RM4VGVsv5_0),.clk(gclk));
	jdff dff_B_jWLrh7su1_0(.din(w_dff_B_RM4VGVsv5_0),.dout(w_dff_B_jWLrh7su1_0),.clk(gclk));
	jdff dff_B_lo2pgxl81_0(.din(w_dff_B_jWLrh7su1_0),.dout(w_dff_B_lo2pgxl81_0),.clk(gclk));
	jdff dff_B_A495pgkA5_0(.din(w_dff_B_lo2pgxl81_0),.dout(w_dff_B_A495pgkA5_0),.clk(gclk));
	jdff dff_B_VxyDIn9V8_0(.din(w_dff_B_A495pgkA5_0),.dout(w_dff_B_VxyDIn9V8_0),.clk(gclk));
	jdff dff_B_LU1BuPt49_0(.din(w_dff_B_VxyDIn9V8_0),.dout(w_dff_B_LU1BuPt49_0),.clk(gclk));
	jdff dff_B_fSaz2gyY1_0(.din(w_dff_B_LU1BuPt49_0),.dout(w_dff_B_fSaz2gyY1_0),.clk(gclk));
	jdff dff_B_rNCyxoNw2_0(.din(w_dff_B_fSaz2gyY1_0),.dout(w_dff_B_rNCyxoNw2_0),.clk(gclk));
	jdff dff_B_7k4Da50G6_0(.din(w_dff_B_rNCyxoNw2_0),.dout(w_dff_B_7k4Da50G6_0),.clk(gclk));
	jdff dff_B_Xaq2Q8Nu8_0(.din(w_dff_B_7k4Da50G6_0),.dout(w_dff_B_Xaq2Q8Nu8_0),.clk(gclk));
	jdff dff_B_NKYKeJVu9_0(.din(w_dff_B_Xaq2Q8Nu8_0),.dout(w_dff_B_NKYKeJVu9_0),.clk(gclk));
	jdff dff_B_hbroTsbw5_0(.din(w_dff_B_NKYKeJVu9_0),.dout(w_dff_B_hbroTsbw5_0),.clk(gclk));
	jdff dff_B_lbstM2MV7_0(.din(w_dff_B_hbroTsbw5_0),.dout(w_dff_B_lbstM2MV7_0),.clk(gclk));
	jdff dff_B_2RgDHNzc0_0(.din(w_dff_B_lbstM2MV7_0),.dout(w_dff_B_2RgDHNzc0_0),.clk(gclk));
	jdff dff_B_5DCwVdQC5_0(.din(w_dff_B_2RgDHNzc0_0),.dout(w_dff_B_5DCwVdQC5_0),.clk(gclk));
	jdff dff_B_mT5R6jG87_0(.din(n1078),.dout(w_dff_B_mT5R6jG87_0),.clk(gclk));
	jdff dff_B_mIhfyMt21_0(.din(w_dff_B_mT5R6jG87_0),.dout(w_dff_B_mIhfyMt21_0),.clk(gclk));
	jdff dff_B_QtSRwaCV7_0(.din(w_dff_B_mIhfyMt21_0),.dout(w_dff_B_QtSRwaCV7_0),.clk(gclk));
	jdff dff_B_CZ2aD6hQ4_0(.din(w_dff_B_QtSRwaCV7_0),.dout(w_dff_B_CZ2aD6hQ4_0),.clk(gclk));
	jdff dff_B_GFrAB78X7_0(.din(w_dff_B_CZ2aD6hQ4_0),.dout(w_dff_B_GFrAB78X7_0),.clk(gclk));
	jdff dff_B_lf7v4Nnh0_0(.din(w_dff_B_GFrAB78X7_0),.dout(w_dff_B_lf7v4Nnh0_0),.clk(gclk));
	jdff dff_B_tMnsVjYJ7_0(.din(w_dff_B_lf7v4Nnh0_0),.dout(w_dff_B_tMnsVjYJ7_0),.clk(gclk));
	jdff dff_B_p9OIkyt69_0(.din(w_dff_B_tMnsVjYJ7_0),.dout(w_dff_B_p9OIkyt69_0),.clk(gclk));
	jdff dff_B_rilLkg6K7_0(.din(w_dff_B_p9OIkyt69_0),.dout(w_dff_B_rilLkg6K7_0),.clk(gclk));
	jdff dff_B_qVUAyPpR9_0(.din(w_dff_B_rilLkg6K7_0),.dout(w_dff_B_qVUAyPpR9_0),.clk(gclk));
	jdff dff_B_KSsHrZsN1_0(.din(w_dff_B_qVUAyPpR9_0),.dout(w_dff_B_KSsHrZsN1_0),.clk(gclk));
	jdff dff_B_k7tcXP4j7_0(.din(w_dff_B_KSsHrZsN1_0),.dout(w_dff_B_k7tcXP4j7_0),.clk(gclk));
	jdff dff_B_r9Mik5vs3_0(.din(w_dff_B_k7tcXP4j7_0),.dout(w_dff_B_r9Mik5vs3_0),.clk(gclk));
	jdff dff_B_NF5QXmlA3_0(.din(w_dff_B_r9Mik5vs3_0),.dout(w_dff_B_NF5QXmlA3_0),.clk(gclk));
	jdff dff_B_jNvoTVNr1_0(.din(w_dff_B_NF5QXmlA3_0),.dout(w_dff_B_jNvoTVNr1_0),.clk(gclk));
	jdff dff_B_i0mzmYiS7_0(.din(w_dff_B_jNvoTVNr1_0),.dout(w_dff_B_i0mzmYiS7_0),.clk(gclk));
	jdff dff_B_XFSAAHqQ4_0(.din(w_dff_B_i0mzmYiS7_0),.dout(w_dff_B_XFSAAHqQ4_0),.clk(gclk));
	jdff dff_B_EhXTZVmp6_0(.din(w_dff_B_XFSAAHqQ4_0),.dout(w_dff_B_EhXTZVmp6_0),.clk(gclk));
	jdff dff_B_eCEc1y8j3_0(.din(w_dff_B_EhXTZVmp6_0),.dout(w_dff_B_eCEc1y8j3_0),.clk(gclk));
	jdff dff_B_Gmku2spy9_0(.din(w_dff_B_eCEc1y8j3_0),.dout(w_dff_B_Gmku2spy9_0),.clk(gclk));
	jdff dff_B_puhSnyon2_0(.din(w_dff_B_Gmku2spy9_0),.dout(w_dff_B_puhSnyon2_0),.clk(gclk));
	jdff dff_B_zYqCHeFc9_0(.din(w_dff_B_puhSnyon2_0),.dout(w_dff_B_zYqCHeFc9_0),.clk(gclk));
	jdff dff_B_U8RzyLka3_0(.din(w_dff_B_zYqCHeFc9_0),.dout(w_dff_B_U8RzyLka3_0),.clk(gclk));
	jdff dff_B_7q24LWYe6_0(.din(w_dff_B_U8RzyLka3_0),.dout(w_dff_B_7q24LWYe6_0),.clk(gclk));
	jdff dff_B_j10PvIAu6_0(.din(w_dff_B_7q24LWYe6_0),.dout(w_dff_B_j10PvIAu6_0),.clk(gclk));
	jdff dff_B_LycHESkq9_0(.din(w_dff_B_j10PvIAu6_0),.dout(w_dff_B_LycHESkq9_0),.clk(gclk));
	jdff dff_B_J4jM6YNu7_0(.din(w_dff_B_LycHESkq9_0),.dout(w_dff_B_J4jM6YNu7_0),.clk(gclk));
	jdff dff_B_4BdIKe0Y2_0(.din(w_dff_B_J4jM6YNu7_0),.dout(w_dff_B_4BdIKe0Y2_0),.clk(gclk));
	jdff dff_B_IT84bfga5_0(.din(w_dff_B_4BdIKe0Y2_0),.dout(w_dff_B_IT84bfga5_0),.clk(gclk));
	jdff dff_B_zuwhgRWo6_0(.din(w_dff_B_IT84bfga5_0),.dout(w_dff_B_zuwhgRWo6_0),.clk(gclk));
	jdff dff_B_tqRdfYdx0_0(.din(w_dff_B_zuwhgRWo6_0),.dout(w_dff_B_tqRdfYdx0_0),.clk(gclk));
	jdff dff_B_SZrUMgEJ2_0(.din(w_dff_B_tqRdfYdx0_0),.dout(w_dff_B_SZrUMgEJ2_0),.clk(gclk));
	jdff dff_B_kLHknRFj5_0(.din(w_dff_B_SZrUMgEJ2_0),.dout(w_dff_B_kLHknRFj5_0),.clk(gclk));
	jdff dff_B_04PfymOH4_0(.din(w_dff_B_kLHknRFj5_0),.dout(w_dff_B_04PfymOH4_0),.clk(gclk));
	jdff dff_B_Qz3IzuF57_0(.din(w_dff_B_04PfymOH4_0),.dout(w_dff_B_Qz3IzuF57_0),.clk(gclk));
	jdff dff_B_rXGf7Xad9_0(.din(w_dff_B_Qz3IzuF57_0),.dout(w_dff_B_rXGf7Xad9_0),.clk(gclk));
	jdff dff_B_dVHsq43y5_0(.din(w_dff_B_rXGf7Xad9_0),.dout(w_dff_B_dVHsq43y5_0),.clk(gclk));
	jdff dff_B_SA4ZvnlD5_0(.din(w_dff_B_dVHsq43y5_0),.dout(w_dff_B_SA4ZvnlD5_0),.clk(gclk));
	jdff dff_B_ZijGJxIu2_0(.din(w_dff_B_SA4ZvnlD5_0),.dout(w_dff_B_ZijGJxIu2_0),.clk(gclk));
	jdff dff_B_aKc547s88_0(.din(w_dff_B_ZijGJxIu2_0),.dout(w_dff_B_aKc547s88_0),.clk(gclk));
	jdff dff_B_yUzHJh7E5_0(.din(w_dff_B_aKc547s88_0),.dout(w_dff_B_yUzHJh7E5_0),.clk(gclk));
	jdff dff_B_RTeMNHTZ5_0(.din(w_dff_B_yUzHJh7E5_0),.dout(w_dff_B_RTeMNHTZ5_0),.clk(gclk));
	jdff dff_B_izNEmQzV3_0(.din(w_dff_B_RTeMNHTZ5_0),.dout(w_dff_B_izNEmQzV3_0),.clk(gclk));
	jdff dff_B_DsVZS0sS3_0(.din(w_dff_B_izNEmQzV3_0),.dout(w_dff_B_DsVZS0sS3_0),.clk(gclk));
	jdff dff_B_ZN7c288f0_0(.din(w_dff_B_DsVZS0sS3_0),.dout(w_dff_B_ZN7c288f0_0),.clk(gclk));
	jdff dff_B_SdSoa2yY1_0(.din(w_dff_B_ZN7c288f0_0),.dout(w_dff_B_SdSoa2yY1_0),.clk(gclk));
	jdff dff_B_3uBwT7VQ4_0(.din(w_dff_B_SdSoa2yY1_0),.dout(w_dff_B_3uBwT7VQ4_0),.clk(gclk));
	jdff dff_B_RCL9xhQg7_0(.din(w_dff_B_3uBwT7VQ4_0),.dout(w_dff_B_RCL9xhQg7_0),.clk(gclk));
	jdff dff_B_8MrJ8lXq4_0(.din(w_dff_B_RCL9xhQg7_0),.dout(w_dff_B_8MrJ8lXq4_0),.clk(gclk));
	jdff dff_B_vPkze0ct4_0(.din(w_dff_B_8MrJ8lXq4_0),.dout(w_dff_B_vPkze0ct4_0),.clk(gclk));
	jdff dff_B_usXJsdDZ1_0(.din(w_dff_B_vPkze0ct4_0),.dout(w_dff_B_usXJsdDZ1_0),.clk(gclk));
	jdff dff_B_BIxuUcjS6_0(.din(w_dff_B_usXJsdDZ1_0),.dout(w_dff_B_BIxuUcjS6_0),.clk(gclk));
	jdff dff_B_3JNl8jYy3_0(.din(w_dff_B_BIxuUcjS6_0),.dout(w_dff_B_3JNl8jYy3_0),.clk(gclk));
	jdff dff_B_1pR10h4d4_0(.din(w_dff_B_3JNl8jYy3_0),.dout(w_dff_B_1pR10h4d4_0),.clk(gclk));
	jdff dff_B_yH5iCWGi5_0(.din(w_dff_B_1pR10h4d4_0),.dout(w_dff_B_yH5iCWGi5_0),.clk(gclk));
	jdff dff_B_MudU0od86_0(.din(w_dff_B_yH5iCWGi5_0),.dout(w_dff_B_MudU0od86_0),.clk(gclk));
	jdff dff_B_8Tv1xEOP9_0(.din(w_dff_B_MudU0od86_0),.dout(w_dff_B_8Tv1xEOP9_0),.clk(gclk));
	jdff dff_B_Ic6ZXSpk0_0(.din(w_dff_B_8Tv1xEOP9_0),.dout(w_dff_B_Ic6ZXSpk0_0),.clk(gclk));
	jdff dff_B_hXD6z7MN7_0(.din(w_dff_B_Ic6ZXSpk0_0),.dout(w_dff_B_hXD6z7MN7_0),.clk(gclk));
	jdff dff_B_xUfZZOJ30_0(.din(w_dff_B_hXD6z7MN7_0),.dout(w_dff_B_xUfZZOJ30_0),.clk(gclk));
	jdff dff_B_LKc93ApG2_0(.din(w_dff_B_xUfZZOJ30_0),.dout(w_dff_B_LKc93ApG2_0),.clk(gclk));
	jdff dff_B_XuRZNCMp8_0(.din(w_dff_B_LKc93ApG2_0),.dout(w_dff_B_XuRZNCMp8_0),.clk(gclk));
	jdff dff_B_vOnBnEEc6_0(.din(w_dff_B_XuRZNCMp8_0),.dout(w_dff_B_vOnBnEEc6_0),.clk(gclk));
	jdff dff_B_vBjaB1Kv5_0(.din(w_dff_B_vOnBnEEc6_0),.dout(w_dff_B_vBjaB1Kv5_0),.clk(gclk));
	jdff dff_B_K8b7Wkp80_0(.din(w_dff_B_vBjaB1Kv5_0),.dout(w_dff_B_K8b7Wkp80_0),.clk(gclk));
	jdff dff_B_4sGtHFz83_0(.din(w_dff_B_K8b7Wkp80_0),.dout(w_dff_B_4sGtHFz83_0),.clk(gclk));
	jdff dff_B_D3wjCbNs9_0(.din(w_dff_B_4sGtHFz83_0),.dout(w_dff_B_D3wjCbNs9_0),.clk(gclk));
	jdff dff_B_MIEFg4NP4_0(.din(w_dff_B_D3wjCbNs9_0),.dout(w_dff_B_MIEFg4NP4_0),.clk(gclk));
	jdff dff_B_VW2R976v3_0(.din(w_dff_B_MIEFg4NP4_0),.dout(w_dff_B_VW2R976v3_0),.clk(gclk));
	jdff dff_B_e1EDcwHP2_0(.din(w_dff_B_VW2R976v3_0),.dout(w_dff_B_e1EDcwHP2_0),.clk(gclk));
	jdff dff_B_0DL2AU736_0(.din(w_dff_B_e1EDcwHP2_0),.dout(w_dff_B_0DL2AU736_0),.clk(gclk));
	jdff dff_B_pGU1PONX9_0(.din(w_dff_B_0DL2AU736_0),.dout(w_dff_B_pGU1PONX9_0),.clk(gclk));
	jdff dff_B_7vcrAh8U1_0(.din(w_dff_B_pGU1PONX9_0),.dout(w_dff_B_7vcrAh8U1_0),.clk(gclk));
	jdff dff_B_QYa9mtG04_0(.din(w_dff_B_7vcrAh8U1_0),.dout(w_dff_B_QYa9mtG04_0),.clk(gclk));
	jdff dff_B_0VzXXHas3_0(.din(w_dff_B_QYa9mtG04_0),.dout(w_dff_B_0VzXXHas3_0),.clk(gclk));
	jdff dff_B_heA6ovfd9_0(.din(w_dff_B_0VzXXHas3_0),.dout(w_dff_B_heA6ovfd9_0),.clk(gclk));
	jdff dff_B_WGCSYcQp2_0(.din(w_dff_B_heA6ovfd9_0),.dout(w_dff_B_WGCSYcQp2_0),.clk(gclk));
	jdff dff_B_TepX1mJy4_0(.din(w_dff_B_WGCSYcQp2_0),.dout(w_dff_B_TepX1mJy4_0),.clk(gclk));
	jdff dff_B_h8NG1vhQ1_0(.din(w_dff_B_TepX1mJy4_0),.dout(w_dff_B_h8NG1vhQ1_0),.clk(gclk));
	jdff dff_B_liZh6P9O6_0(.din(w_dff_B_h8NG1vhQ1_0),.dout(w_dff_B_liZh6P9O6_0),.clk(gclk));
	jdff dff_B_t7m5dmNK3_0(.din(w_dff_B_liZh6P9O6_0),.dout(w_dff_B_t7m5dmNK3_0),.clk(gclk));
	jdff dff_B_jY8FVxd07_0(.din(w_dff_B_t7m5dmNK3_0),.dout(w_dff_B_jY8FVxd07_0),.clk(gclk));
	jdff dff_B_ltuIUQgE2_0(.din(w_dff_B_jY8FVxd07_0),.dout(w_dff_B_ltuIUQgE2_0),.clk(gclk));
	jdff dff_B_OijgP3js1_0(.din(w_dff_B_ltuIUQgE2_0),.dout(w_dff_B_OijgP3js1_0),.clk(gclk));
	jdff dff_B_J9gvKhVz0_0(.din(w_dff_B_OijgP3js1_0),.dout(w_dff_B_J9gvKhVz0_0),.clk(gclk));
	jdff dff_B_sA4odH6z4_0(.din(w_dff_B_J9gvKhVz0_0),.dout(w_dff_B_sA4odH6z4_0),.clk(gclk));
	jdff dff_B_KKQcqHFT5_0(.din(w_dff_B_sA4odH6z4_0),.dout(w_dff_B_KKQcqHFT5_0),.clk(gclk));
	jdff dff_B_iBJsnuCg0_0(.din(w_dff_B_KKQcqHFT5_0),.dout(w_dff_B_iBJsnuCg0_0),.clk(gclk));
	jdff dff_B_nRwV1o3D6_0(.din(w_dff_B_iBJsnuCg0_0),.dout(w_dff_B_nRwV1o3D6_0),.clk(gclk));
	jdff dff_B_NE8vMLC30_0(.din(w_dff_B_nRwV1o3D6_0),.dout(w_dff_B_NE8vMLC30_0),.clk(gclk));
	jdff dff_B_jTuWiCzY7_0(.din(w_dff_B_NE8vMLC30_0),.dout(w_dff_B_jTuWiCzY7_0),.clk(gclk));
	jdff dff_B_ruBSvo7p8_0(.din(w_dff_B_jTuWiCzY7_0),.dout(w_dff_B_ruBSvo7p8_0),.clk(gclk));
	jdff dff_B_5GLQo37P4_0(.din(w_dff_B_ruBSvo7p8_0),.dout(w_dff_B_5GLQo37P4_0),.clk(gclk));
	jdff dff_B_G4SMXkX32_0(.din(w_dff_B_5GLQo37P4_0),.dout(w_dff_B_G4SMXkX32_0),.clk(gclk));
	jdff dff_B_Qus7NFco4_0(.din(w_dff_B_G4SMXkX32_0),.dout(w_dff_B_Qus7NFco4_0),.clk(gclk));
	jdff dff_B_6dujABMS3_0(.din(w_dff_B_Qus7NFco4_0),.dout(w_dff_B_6dujABMS3_0),.clk(gclk));
	jdff dff_B_J6S3xhdH7_0(.din(w_dff_B_6dujABMS3_0),.dout(w_dff_B_J6S3xhdH7_0),.clk(gclk));
	jdff dff_B_Ld0uTr3D8_0(.din(w_dff_B_J6S3xhdH7_0),.dout(w_dff_B_Ld0uTr3D8_0),.clk(gclk));
	jdff dff_B_8XdTk8ch5_0(.din(w_dff_B_Ld0uTr3D8_0),.dout(w_dff_B_8XdTk8ch5_0),.clk(gclk));
	jdff dff_B_jfc1YHB47_0(.din(w_dff_B_8XdTk8ch5_0),.dout(w_dff_B_jfc1YHB47_0),.clk(gclk));
	jdff dff_B_6vJjOm7R7_0(.din(w_dff_B_jfc1YHB47_0),.dout(w_dff_B_6vJjOm7R7_0),.clk(gclk));
	jdff dff_B_kzx7Qa7Z2_0(.din(w_dff_B_6vJjOm7R7_0),.dout(w_dff_B_kzx7Qa7Z2_0),.clk(gclk));
	jdff dff_B_QvU9Dc3X3_0(.din(w_dff_B_kzx7Qa7Z2_0),.dout(w_dff_B_QvU9Dc3X3_0),.clk(gclk));
	jdff dff_B_6yz624wj1_0(.din(w_dff_B_QvU9Dc3X3_0),.dout(w_dff_B_6yz624wj1_0),.clk(gclk));
	jdff dff_B_zEJtToqs3_0(.din(w_dff_B_6yz624wj1_0),.dout(w_dff_B_zEJtToqs3_0),.clk(gclk));
	jdff dff_B_p2OEjJJb5_0(.din(w_dff_B_zEJtToqs3_0),.dout(w_dff_B_p2OEjJJb5_0),.clk(gclk));
	jdff dff_B_pPzyjyLF1_0(.din(w_dff_B_p2OEjJJb5_0),.dout(w_dff_B_pPzyjyLF1_0),.clk(gclk));
	jdff dff_B_dvlsUwcj9_0(.din(w_dff_B_pPzyjyLF1_0),.dout(w_dff_B_dvlsUwcj9_0),.clk(gclk));
	jdff dff_B_IBM8fJMC1_0(.din(w_dff_B_dvlsUwcj9_0),.dout(w_dff_B_IBM8fJMC1_0),.clk(gclk));
	jdff dff_B_irXSsmDw9_0(.din(w_dff_B_IBM8fJMC1_0),.dout(w_dff_B_irXSsmDw9_0),.clk(gclk));
	jdff dff_B_y4jpDxnt1_0(.din(w_dff_B_irXSsmDw9_0),.dout(w_dff_B_y4jpDxnt1_0),.clk(gclk));
	jdff dff_B_WrHyyegD7_0(.din(w_dff_B_y4jpDxnt1_0),.dout(w_dff_B_WrHyyegD7_0),.clk(gclk));
	jdff dff_B_FAYirqBa0_0(.din(w_dff_B_WrHyyegD7_0),.dout(w_dff_B_FAYirqBa0_0),.clk(gclk));
	jdff dff_B_3eMcAsGG5_0(.din(w_dff_B_FAYirqBa0_0),.dout(w_dff_B_3eMcAsGG5_0),.clk(gclk));
	jdff dff_B_t66iQooO7_0(.din(w_dff_B_3eMcAsGG5_0),.dout(w_dff_B_t66iQooO7_0),.clk(gclk));
	jdff dff_B_OgbsSv5y6_0(.din(n1084),.dout(w_dff_B_OgbsSv5y6_0),.clk(gclk));
	jdff dff_B_bj17yU8k5_0(.din(w_dff_B_OgbsSv5y6_0),.dout(w_dff_B_bj17yU8k5_0),.clk(gclk));
	jdff dff_B_DOU5GeaM0_0(.din(w_dff_B_bj17yU8k5_0),.dout(w_dff_B_DOU5GeaM0_0),.clk(gclk));
	jdff dff_B_QJPgP2Ii8_0(.din(w_dff_B_DOU5GeaM0_0),.dout(w_dff_B_QJPgP2Ii8_0),.clk(gclk));
	jdff dff_B_dvTrZ2uC7_0(.din(w_dff_B_QJPgP2Ii8_0),.dout(w_dff_B_dvTrZ2uC7_0),.clk(gclk));
	jdff dff_B_1J0CQA1T1_0(.din(w_dff_B_dvTrZ2uC7_0),.dout(w_dff_B_1J0CQA1T1_0),.clk(gclk));
	jdff dff_B_O5pd8KNF2_0(.din(w_dff_B_1J0CQA1T1_0),.dout(w_dff_B_O5pd8KNF2_0),.clk(gclk));
	jdff dff_B_xKyJSnvx9_0(.din(w_dff_B_O5pd8KNF2_0),.dout(w_dff_B_xKyJSnvx9_0),.clk(gclk));
	jdff dff_B_xUxwdEOO4_0(.din(w_dff_B_xKyJSnvx9_0),.dout(w_dff_B_xUxwdEOO4_0),.clk(gclk));
	jdff dff_B_WvWxvWzg8_0(.din(w_dff_B_xUxwdEOO4_0),.dout(w_dff_B_WvWxvWzg8_0),.clk(gclk));
	jdff dff_B_4JurAnWO1_0(.din(w_dff_B_WvWxvWzg8_0),.dout(w_dff_B_4JurAnWO1_0),.clk(gclk));
	jdff dff_B_1PywuMYM8_0(.din(w_dff_B_4JurAnWO1_0),.dout(w_dff_B_1PywuMYM8_0),.clk(gclk));
	jdff dff_B_qQK6xdmP0_0(.din(w_dff_B_1PywuMYM8_0),.dout(w_dff_B_qQK6xdmP0_0),.clk(gclk));
	jdff dff_B_yHbwg9zI7_0(.din(w_dff_B_qQK6xdmP0_0),.dout(w_dff_B_yHbwg9zI7_0),.clk(gclk));
	jdff dff_B_e35l5UNQ1_0(.din(w_dff_B_yHbwg9zI7_0),.dout(w_dff_B_e35l5UNQ1_0),.clk(gclk));
	jdff dff_B_cdkBYG2h0_0(.din(w_dff_B_e35l5UNQ1_0),.dout(w_dff_B_cdkBYG2h0_0),.clk(gclk));
	jdff dff_B_IG7pST6V5_0(.din(w_dff_B_cdkBYG2h0_0),.dout(w_dff_B_IG7pST6V5_0),.clk(gclk));
	jdff dff_B_EPH60IHt3_0(.din(w_dff_B_IG7pST6V5_0),.dout(w_dff_B_EPH60IHt3_0),.clk(gclk));
	jdff dff_B_l5qyYNxV1_0(.din(w_dff_B_EPH60IHt3_0),.dout(w_dff_B_l5qyYNxV1_0),.clk(gclk));
	jdff dff_B_IAiQbhVG9_0(.din(w_dff_B_l5qyYNxV1_0),.dout(w_dff_B_IAiQbhVG9_0),.clk(gclk));
	jdff dff_B_fnq00r5f8_0(.din(w_dff_B_IAiQbhVG9_0),.dout(w_dff_B_fnq00r5f8_0),.clk(gclk));
	jdff dff_B_hAq0AFvq7_0(.din(w_dff_B_fnq00r5f8_0),.dout(w_dff_B_hAq0AFvq7_0),.clk(gclk));
	jdff dff_B_rwtN9Dwa0_0(.din(w_dff_B_hAq0AFvq7_0),.dout(w_dff_B_rwtN9Dwa0_0),.clk(gclk));
	jdff dff_B_e8jJu26v3_0(.din(w_dff_B_rwtN9Dwa0_0),.dout(w_dff_B_e8jJu26v3_0),.clk(gclk));
	jdff dff_B_eHsvm46h3_0(.din(w_dff_B_e8jJu26v3_0),.dout(w_dff_B_eHsvm46h3_0),.clk(gclk));
	jdff dff_B_TtgmAGTn0_0(.din(w_dff_B_eHsvm46h3_0),.dout(w_dff_B_TtgmAGTn0_0),.clk(gclk));
	jdff dff_B_4EMNny3E5_0(.din(w_dff_B_TtgmAGTn0_0),.dout(w_dff_B_4EMNny3E5_0),.clk(gclk));
	jdff dff_B_u2LK2WNV2_0(.din(w_dff_B_4EMNny3E5_0),.dout(w_dff_B_u2LK2WNV2_0),.clk(gclk));
	jdff dff_B_BfiVhUQz3_0(.din(w_dff_B_u2LK2WNV2_0),.dout(w_dff_B_BfiVhUQz3_0),.clk(gclk));
	jdff dff_B_7KHaRl9h8_0(.din(w_dff_B_BfiVhUQz3_0),.dout(w_dff_B_7KHaRl9h8_0),.clk(gclk));
	jdff dff_B_4ZgDo9038_0(.din(w_dff_B_7KHaRl9h8_0),.dout(w_dff_B_4ZgDo9038_0),.clk(gclk));
	jdff dff_B_7vLfPSF12_0(.din(w_dff_B_4ZgDo9038_0),.dout(w_dff_B_7vLfPSF12_0),.clk(gclk));
	jdff dff_B_qwfiJ8jA7_0(.din(w_dff_B_7vLfPSF12_0),.dout(w_dff_B_qwfiJ8jA7_0),.clk(gclk));
	jdff dff_B_Gn6RKfnD8_0(.din(w_dff_B_qwfiJ8jA7_0),.dout(w_dff_B_Gn6RKfnD8_0),.clk(gclk));
	jdff dff_B_VoKB9te33_0(.din(w_dff_B_Gn6RKfnD8_0),.dout(w_dff_B_VoKB9te33_0),.clk(gclk));
	jdff dff_B_i5Ln6cRk3_0(.din(w_dff_B_VoKB9te33_0),.dout(w_dff_B_i5Ln6cRk3_0),.clk(gclk));
	jdff dff_B_dRIK55IK4_0(.din(w_dff_B_i5Ln6cRk3_0),.dout(w_dff_B_dRIK55IK4_0),.clk(gclk));
	jdff dff_B_yHwN6seX7_0(.din(w_dff_B_dRIK55IK4_0),.dout(w_dff_B_yHwN6seX7_0),.clk(gclk));
	jdff dff_B_1hYcPsh28_0(.din(w_dff_B_yHwN6seX7_0),.dout(w_dff_B_1hYcPsh28_0),.clk(gclk));
	jdff dff_B_iQdA0oYB7_0(.din(w_dff_B_1hYcPsh28_0),.dout(w_dff_B_iQdA0oYB7_0),.clk(gclk));
	jdff dff_B_ONiY33U54_0(.din(w_dff_B_iQdA0oYB7_0),.dout(w_dff_B_ONiY33U54_0),.clk(gclk));
	jdff dff_B_SsvILKT16_0(.din(w_dff_B_ONiY33U54_0),.dout(w_dff_B_SsvILKT16_0),.clk(gclk));
	jdff dff_B_DPy1PlS17_0(.din(w_dff_B_SsvILKT16_0),.dout(w_dff_B_DPy1PlS17_0),.clk(gclk));
	jdff dff_B_dQL4cCvp1_0(.din(w_dff_B_DPy1PlS17_0),.dout(w_dff_B_dQL4cCvp1_0),.clk(gclk));
	jdff dff_B_zHY7OdU13_0(.din(w_dff_B_dQL4cCvp1_0),.dout(w_dff_B_zHY7OdU13_0),.clk(gclk));
	jdff dff_B_EpjFEFeS6_0(.din(w_dff_B_zHY7OdU13_0),.dout(w_dff_B_EpjFEFeS6_0),.clk(gclk));
	jdff dff_B_M9AbqevZ7_0(.din(w_dff_B_EpjFEFeS6_0),.dout(w_dff_B_M9AbqevZ7_0),.clk(gclk));
	jdff dff_B_N3uT70rS9_0(.din(w_dff_B_M9AbqevZ7_0),.dout(w_dff_B_N3uT70rS9_0),.clk(gclk));
	jdff dff_B_Kzc4vf1Y8_0(.din(w_dff_B_N3uT70rS9_0),.dout(w_dff_B_Kzc4vf1Y8_0),.clk(gclk));
	jdff dff_B_qeU1Jg9J3_0(.din(w_dff_B_Kzc4vf1Y8_0),.dout(w_dff_B_qeU1Jg9J3_0),.clk(gclk));
	jdff dff_B_YxVz6JQl8_0(.din(w_dff_B_qeU1Jg9J3_0),.dout(w_dff_B_YxVz6JQl8_0),.clk(gclk));
	jdff dff_B_FoBnzwng2_0(.din(w_dff_B_YxVz6JQl8_0),.dout(w_dff_B_FoBnzwng2_0),.clk(gclk));
	jdff dff_B_ydFqt54R5_0(.din(w_dff_B_FoBnzwng2_0),.dout(w_dff_B_ydFqt54R5_0),.clk(gclk));
	jdff dff_B_0Yk60AUn4_0(.din(w_dff_B_ydFqt54R5_0),.dout(w_dff_B_0Yk60AUn4_0),.clk(gclk));
	jdff dff_B_KWjZkP2Z7_0(.din(w_dff_B_0Yk60AUn4_0),.dout(w_dff_B_KWjZkP2Z7_0),.clk(gclk));
	jdff dff_B_jaK0c1Xn0_0(.din(w_dff_B_KWjZkP2Z7_0),.dout(w_dff_B_jaK0c1Xn0_0),.clk(gclk));
	jdff dff_B_7EiIuLxG6_0(.din(w_dff_B_jaK0c1Xn0_0),.dout(w_dff_B_7EiIuLxG6_0),.clk(gclk));
	jdff dff_B_yzxG5pAF8_0(.din(w_dff_B_7EiIuLxG6_0),.dout(w_dff_B_yzxG5pAF8_0),.clk(gclk));
	jdff dff_B_m2cDGtgO7_0(.din(w_dff_B_yzxG5pAF8_0),.dout(w_dff_B_m2cDGtgO7_0),.clk(gclk));
	jdff dff_B_KXAHi7d68_0(.din(w_dff_B_m2cDGtgO7_0),.dout(w_dff_B_KXAHi7d68_0),.clk(gclk));
	jdff dff_B_OwyZ7XQu4_0(.din(w_dff_B_KXAHi7d68_0),.dout(w_dff_B_OwyZ7XQu4_0),.clk(gclk));
	jdff dff_B_8nhSkh2d0_0(.din(w_dff_B_OwyZ7XQu4_0),.dout(w_dff_B_8nhSkh2d0_0),.clk(gclk));
	jdff dff_B_doTWgxu09_0(.din(w_dff_B_8nhSkh2d0_0),.dout(w_dff_B_doTWgxu09_0),.clk(gclk));
	jdff dff_B_DfJVRy199_0(.din(w_dff_B_doTWgxu09_0),.dout(w_dff_B_DfJVRy199_0),.clk(gclk));
	jdff dff_B_YryYg53B0_0(.din(w_dff_B_DfJVRy199_0),.dout(w_dff_B_YryYg53B0_0),.clk(gclk));
	jdff dff_B_tDNBPcBN1_0(.din(w_dff_B_YryYg53B0_0),.dout(w_dff_B_tDNBPcBN1_0),.clk(gclk));
	jdff dff_B_VYbjiQVo0_0(.din(w_dff_B_tDNBPcBN1_0),.dout(w_dff_B_VYbjiQVo0_0),.clk(gclk));
	jdff dff_B_SvvQIaor6_0(.din(w_dff_B_VYbjiQVo0_0),.dout(w_dff_B_SvvQIaor6_0),.clk(gclk));
	jdff dff_B_Mbm0k7Ty0_0(.din(w_dff_B_SvvQIaor6_0),.dout(w_dff_B_Mbm0k7Ty0_0),.clk(gclk));
	jdff dff_B_KNGBHHix8_0(.din(w_dff_B_Mbm0k7Ty0_0),.dout(w_dff_B_KNGBHHix8_0),.clk(gclk));
	jdff dff_B_liyVAZm50_0(.din(w_dff_B_KNGBHHix8_0),.dout(w_dff_B_liyVAZm50_0),.clk(gclk));
	jdff dff_B_tmovH3rI1_0(.din(w_dff_B_liyVAZm50_0),.dout(w_dff_B_tmovH3rI1_0),.clk(gclk));
	jdff dff_B_vLltUVYY5_0(.din(w_dff_B_tmovH3rI1_0),.dout(w_dff_B_vLltUVYY5_0),.clk(gclk));
	jdff dff_B_AKb6EvBO0_0(.din(w_dff_B_vLltUVYY5_0),.dout(w_dff_B_AKb6EvBO0_0),.clk(gclk));
	jdff dff_B_OCrwxUvx1_0(.din(w_dff_B_AKb6EvBO0_0),.dout(w_dff_B_OCrwxUvx1_0),.clk(gclk));
	jdff dff_B_w7pQ7NKj8_0(.din(w_dff_B_OCrwxUvx1_0),.dout(w_dff_B_w7pQ7NKj8_0),.clk(gclk));
	jdff dff_B_k1aDtxx55_0(.din(w_dff_B_w7pQ7NKj8_0),.dout(w_dff_B_k1aDtxx55_0),.clk(gclk));
	jdff dff_B_NtITRMw89_0(.din(w_dff_B_k1aDtxx55_0),.dout(w_dff_B_NtITRMw89_0),.clk(gclk));
	jdff dff_B_RvtWyrLH0_0(.din(w_dff_B_NtITRMw89_0),.dout(w_dff_B_RvtWyrLH0_0),.clk(gclk));
	jdff dff_B_9vinJAyS7_0(.din(w_dff_B_RvtWyrLH0_0),.dout(w_dff_B_9vinJAyS7_0),.clk(gclk));
	jdff dff_B_hbD1bP0Y2_0(.din(w_dff_B_9vinJAyS7_0),.dout(w_dff_B_hbD1bP0Y2_0),.clk(gclk));
	jdff dff_B_KOeHJObt7_0(.din(w_dff_B_hbD1bP0Y2_0),.dout(w_dff_B_KOeHJObt7_0),.clk(gclk));
	jdff dff_B_ZlvCaaZo4_0(.din(w_dff_B_KOeHJObt7_0),.dout(w_dff_B_ZlvCaaZo4_0),.clk(gclk));
	jdff dff_B_aLUVpM9m6_0(.din(w_dff_B_ZlvCaaZo4_0),.dout(w_dff_B_aLUVpM9m6_0),.clk(gclk));
	jdff dff_B_UwlWFzeN5_0(.din(w_dff_B_aLUVpM9m6_0),.dout(w_dff_B_UwlWFzeN5_0),.clk(gclk));
	jdff dff_B_UEFFLVhB1_0(.din(w_dff_B_UwlWFzeN5_0),.dout(w_dff_B_UEFFLVhB1_0),.clk(gclk));
	jdff dff_B_0LkHLgGP3_0(.din(w_dff_B_UEFFLVhB1_0),.dout(w_dff_B_0LkHLgGP3_0),.clk(gclk));
	jdff dff_B_G9OQg0hk8_0(.din(w_dff_B_0LkHLgGP3_0),.dout(w_dff_B_G9OQg0hk8_0),.clk(gclk));
	jdff dff_B_fZJ5prOr5_0(.din(w_dff_B_G9OQg0hk8_0),.dout(w_dff_B_fZJ5prOr5_0),.clk(gclk));
	jdff dff_B_MGTlem011_0(.din(w_dff_B_fZJ5prOr5_0),.dout(w_dff_B_MGTlem011_0),.clk(gclk));
	jdff dff_B_P2bGgnOC2_0(.din(w_dff_B_MGTlem011_0),.dout(w_dff_B_P2bGgnOC2_0),.clk(gclk));
	jdff dff_B_gKKZ7ijG5_0(.din(w_dff_B_P2bGgnOC2_0),.dout(w_dff_B_gKKZ7ijG5_0),.clk(gclk));
	jdff dff_B_GZS0JPIc8_0(.din(w_dff_B_gKKZ7ijG5_0),.dout(w_dff_B_GZS0JPIc8_0),.clk(gclk));
	jdff dff_B_BfDKFQb51_0(.din(w_dff_B_GZS0JPIc8_0),.dout(w_dff_B_BfDKFQb51_0),.clk(gclk));
	jdff dff_B_TiIBP8De2_0(.din(w_dff_B_BfDKFQb51_0),.dout(w_dff_B_TiIBP8De2_0),.clk(gclk));
	jdff dff_B_ahi47YUR1_0(.din(w_dff_B_TiIBP8De2_0),.dout(w_dff_B_ahi47YUR1_0),.clk(gclk));
	jdff dff_B_2L9c7xNO9_0(.din(w_dff_B_ahi47YUR1_0),.dout(w_dff_B_2L9c7xNO9_0),.clk(gclk));
	jdff dff_B_cirpKDKK6_0(.din(w_dff_B_2L9c7xNO9_0),.dout(w_dff_B_cirpKDKK6_0),.clk(gclk));
	jdff dff_B_YTaqmtxP4_0(.din(w_dff_B_cirpKDKK6_0),.dout(w_dff_B_YTaqmtxP4_0),.clk(gclk));
	jdff dff_B_pbCKghN20_0(.din(w_dff_B_YTaqmtxP4_0),.dout(w_dff_B_pbCKghN20_0),.clk(gclk));
	jdff dff_B_5ypTpoPi5_0(.din(w_dff_B_pbCKghN20_0),.dout(w_dff_B_5ypTpoPi5_0),.clk(gclk));
	jdff dff_B_z4G8Pj2d1_0(.din(w_dff_B_5ypTpoPi5_0),.dout(w_dff_B_z4G8Pj2d1_0),.clk(gclk));
	jdff dff_B_jCrwUYlh1_0(.din(w_dff_B_z4G8Pj2d1_0),.dout(w_dff_B_jCrwUYlh1_0),.clk(gclk));
	jdff dff_B_3jsugFd75_0(.din(w_dff_B_jCrwUYlh1_0),.dout(w_dff_B_3jsugFd75_0),.clk(gclk));
	jdff dff_B_h3kS9t0a5_0(.din(w_dff_B_3jsugFd75_0),.dout(w_dff_B_h3kS9t0a5_0),.clk(gclk));
	jdff dff_B_ZQaquU432_0(.din(w_dff_B_h3kS9t0a5_0),.dout(w_dff_B_ZQaquU432_0),.clk(gclk));
	jdff dff_B_LtIRXA7N4_0(.din(w_dff_B_ZQaquU432_0),.dout(w_dff_B_LtIRXA7N4_0),.clk(gclk));
	jdff dff_B_zsf56dpY7_0(.din(w_dff_B_LtIRXA7N4_0),.dout(w_dff_B_zsf56dpY7_0),.clk(gclk));
	jdff dff_B_I6JZrKXq3_0(.din(w_dff_B_zsf56dpY7_0),.dout(w_dff_B_I6JZrKXq3_0),.clk(gclk));
	jdff dff_B_euQRbziA8_0(.din(w_dff_B_I6JZrKXq3_0),.dout(w_dff_B_euQRbziA8_0),.clk(gclk));
	jdff dff_B_mGH4Jypu5_0(.din(w_dff_B_euQRbziA8_0),.dout(w_dff_B_mGH4Jypu5_0),.clk(gclk));
	jdff dff_B_4iPpF1Tk3_0(.din(w_dff_B_mGH4Jypu5_0),.dout(w_dff_B_4iPpF1Tk3_0),.clk(gclk));
	jdff dff_B_mlscRo030_0(.din(w_dff_B_4iPpF1Tk3_0),.dout(w_dff_B_mlscRo030_0),.clk(gclk));
	jdff dff_B_ZTDC1JDE7_0(.din(w_dff_B_mlscRo030_0),.dout(w_dff_B_ZTDC1JDE7_0),.clk(gclk));
	jdff dff_B_TERbME9F8_0(.din(w_dff_B_ZTDC1JDE7_0),.dout(w_dff_B_TERbME9F8_0),.clk(gclk));
	jdff dff_B_Y58xZaMx0_0(.din(w_dff_B_TERbME9F8_0),.dout(w_dff_B_Y58xZaMx0_0),.clk(gclk));
	jdff dff_B_U0SaqLbB5_0(.din(n1090),.dout(w_dff_B_U0SaqLbB5_0),.clk(gclk));
	jdff dff_B_nlS8FHBj7_0(.din(w_dff_B_U0SaqLbB5_0),.dout(w_dff_B_nlS8FHBj7_0),.clk(gclk));
	jdff dff_B_6jrtoveD4_0(.din(w_dff_B_nlS8FHBj7_0),.dout(w_dff_B_6jrtoveD4_0),.clk(gclk));
	jdff dff_B_nrJpjEzB0_0(.din(w_dff_B_6jrtoveD4_0),.dout(w_dff_B_nrJpjEzB0_0),.clk(gclk));
	jdff dff_B_VCHSalno5_0(.din(w_dff_B_nrJpjEzB0_0),.dout(w_dff_B_VCHSalno5_0),.clk(gclk));
	jdff dff_B_sw1P9WON5_0(.din(w_dff_B_VCHSalno5_0),.dout(w_dff_B_sw1P9WON5_0),.clk(gclk));
	jdff dff_B_mqJ7AQMa2_0(.din(w_dff_B_sw1P9WON5_0),.dout(w_dff_B_mqJ7AQMa2_0),.clk(gclk));
	jdff dff_B_0Eyj2soR8_0(.din(w_dff_B_mqJ7AQMa2_0),.dout(w_dff_B_0Eyj2soR8_0),.clk(gclk));
	jdff dff_B_x8wOIjQS5_0(.din(w_dff_B_0Eyj2soR8_0),.dout(w_dff_B_x8wOIjQS5_0),.clk(gclk));
	jdff dff_B_T1tXy2XH0_0(.din(w_dff_B_x8wOIjQS5_0),.dout(w_dff_B_T1tXy2XH0_0),.clk(gclk));
	jdff dff_B_NQAJivaY7_0(.din(w_dff_B_T1tXy2XH0_0),.dout(w_dff_B_NQAJivaY7_0),.clk(gclk));
	jdff dff_B_Hbnqvyz66_0(.din(w_dff_B_NQAJivaY7_0),.dout(w_dff_B_Hbnqvyz66_0),.clk(gclk));
	jdff dff_B_wd0ZXQVw3_0(.din(w_dff_B_Hbnqvyz66_0),.dout(w_dff_B_wd0ZXQVw3_0),.clk(gclk));
	jdff dff_B_yKICTire7_0(.din(w_dff_B_wd0ZXQVw3_0),.dout(w_dff_B_yKICTire7_0),.clk(gclk));
	jdff dff_B_YNYFKqvT1_0(.din(w_dff_B_yKICTire7_0),.dout(w_dff_B_YNYFKqvT1_0),.clk(gclk));
	jdff dff_B_pzm6NvQh4_0(.din(w_dff_B_YNYFKqvT1_0),.dout(w_dff_B_pzm6NvQh4_0),.clk(gclk));
	jdff dff_B_yi97ZAmR0_0(.din(w_dff_B_pzm6NvQh4_0),.dout(w_dff_B_yi97ZAmR0_0),.clk(gclk));
	jdff dff_B_NysdbI4B7_0(.din(w_dff_B_yi97ZAmR0_0),.dout(w_dff_B_NysdbI4B7_0),.clk(gclk));
	jdff dff_B_Z8oEXEOq5_0(.din(w_dff_B_NysdbI4B7_0),.dout(w_dff_B_Z8oEXEOq5_0),.clk(gclk));
	jdff dff_B_PrvvhIbo1_0(.din(w_dff_B_Z8oEXEOq5_0),.dout(w_dff_B_PrvvhIbo1_0),.clk(gclk));
	jdff dff_B_0oklccaG4_0(.din(w_dff_B_PrvvhIbo1_0),.dout(w_dff_B_0oklccaG4_0),.clk(gclk));
	jdff dff_B_uiSXcZUB4_0(.din(w_dff_B_0oklccaG4_0),.dout(w_dff_B_uiSXcZUB4_0),.clk(gclk));
	jdff dff_B_mDeIGuJ43_0(.din(w_dff_B_uiSXcZUB4_0),.dout(w_dff_B_mDeIGuJ43_0),.clk(gclk));
	jdff dff_B_bPjvRbd34_0(.din(w_dff_B_mDeIGuJ43_0),.dout(w_dff_B_bPjvRbd34_0),.clk(gclk));
	jdff dff_B_ENEpxAde1_0(.din(w_dff_B_bPjvRbd34_0),.dout(w_dff_B_ENEpxAde1_0),.clk(gclk));
	jdff dff_B_YYh6OEfL0_0(.din(w_dff_B_ENEpxAde1_0),.dout(w_dff_B_YYh6OEfL0_0),.clk(gclk));
	jdff dff_B_m2uiIz561_0(.din(w_dff_B_YYh6OEfL0_0),.dout(w_dff_B_m2uiIz561_0),.clk(gclk));
	jdff dff_B_kNSsNfC44_0(.din(w_dff_B_m2uiIz561_0),.dout(w_dff_B_kNSsNfC44_0),.clk(gclk));
	jdff dff_B_LiqLZPqr6_0(.din(w_dff_B_kNSsNfC44_0),.dout(w_dff_B_LiqLZPqr6_0),.clk(gclk));
	jdff dff_B_17rldnQW9_0(.din(w_dff_B_LiqLZPqr6_0),.dout(w_dff_B_17rldnQW9_0),.clk(gclk));
	jdff dff_B_whrCssj15_0(.din(w_dff_B_17rldnQW9_0),.dout(w_dff_B_whrCssj15_0),.clk(gclk));
	jdff dff_B_7HpG867R3_0(.din(w_dff_B_whrCssj15_0),.dout(w_dff_B_7HpG867R3_0),.clk(gclk));
	jdff dff_B_3qU7Pgnd1_0(.din(w_dff_B_7HpG867R3_0),.dout(w_dff_B_3qU7Pgnd1_0),.clk(gclk));
	jdff dff_B_VasuzH687_0(.din(w_dff_B_3qU7Pgnd1_0),.dout(w_dff_B_VasuzH687_0),.clk(gclk));
	jdff dff_B_jTSAjFIp4_0(.din(w_dff_B_VasuzH687_0),.dout(w_dff_B_jTSAjFIp4_0),.clk(gclk));
	jdff dff_B_szxPUmwE9_0(.din(w_dff_B_jTSAjFIp4_0),.dout(w_dff_B_szxPUmwE9_0),.clk(gclk));
	jdff dff_B_wILe7lwQ1_0(.din(w_dff_B_szxPUmwE9_0),.dout(w_dff_B_wILe7lwQ1_0),.clk(gclk));
	jdff dff_B_jxkLKYS50_0(.din(w_dff_B_wILe7lwQ1_0),.dout(w_dff_B_jxkLKYS50_0),.clk(gclk));
	jdff dff_B_FDORIHlv4_0(.din(w_dff_B_jxkLKYS50_0),.dout(w_dff_B_FDORIHlv4_0),.clk(gclk));
	jdff dff_B_aAOVCfFw2_0(.din(w_dff_B_FDORIHlv4_0),.dout(w_dff_B_aAOVCfFw2_0),.clk(gclk));
	jdff dff_B_xzNnsrPZ7_0(.din(w_dff_B_aAOVCfFw2_0),.dout(w_dff_B_xzNnsrPZ7_0),.clk(gclk));
	jdff dff_B_DvZpfQh54_0(.din(w_dff_B_xzNnsrPZ7_0),.dout(w_dff_B_DvZpfQh54_0),.clk(gclk));
	jdff dff_B_81zvE9Ef0_0(.din(w_dff_B_DvZpfQh54_0),.dout(w_dff_B_81zvE9Ef0_0),.clk(gclk));
	jdff dff_B_bNJMmZSS0_0(.din(w_dff_B_81zvE9Ef0_0),.dout(w_dff_B_bNJMmZSS0_0),.clk(gclk));
	jdff dff_B_WEjQ75Xz2_0(.din(w_dff_B_bNJMmZSS0_0),.dout(w_dff_B_WEjQ75Xz2_0),.clk(gclk));
	jdff dff_B_od168AOs0_0(.din(w_dff_B_WEjQ75Xz2_0),.dout(w_dff_B_od168AOs0_0),.clk(gclk));
	jdff dff_B_hkNZmOeF6_0(.din(w_dff_B_od168AOs0_0),.dout(w_dff_B_hkNZmOeF6_0),.clk(gclk));
	jdff dff_B_0HABUdRj6_0(.din(w_dff_B_hkNZmOeF6_0),.dout(w_dff_B_0HABUdRj6_0),.clk(gclk));
	jdff dff_B_1Ox4RIbi2_0(.din(w_dff_B_0HABUdRj6_0),.dout(w_dff_B_1Ox4RIbi2_0),.clk(gclk));
	jdff dff_B_urGQZy9D3_0(.din(w_dff_B_1Ox4RIbi2_0),.dout(w_dff_B_urGQZy9D3_0),.clk(gclk));
	jdff dff_B_Et0Ae4xm4_0(.din(w_dff_B_urGQZy9D3_0),.dout(w_dff_B_Et0Ae4xm4_0),.clk(gclk));
	jdff dff_B_eNc3Quge2_0(.din(w_dff_B_Et0Ae4xm4_0),.dout(w_dff_B_eNc3Quge2_0),.clk(gclk));
	jdff dff_B_nRcI7H9Q4_0(.din(w_dff_B_eNc3Quge2_0),.dout(w_dff_B_nRcI7H9Q4_0),.clk(gclk));
	jdff dff_B_kJjiz5uG4_0(.din(w_dff_B_nRcI7H9Q4_0),.dout(w_dff_B_kJjiz5uG4_0),.clk(gclk));
	jdff dff_B_u2z4JjPk5_0(.din(w_dff_B_kJjiz5uG4_0),.dout(w_dff_B_u2z4JjPk5_0),.clk(gclk));
	jdff dff_B_aUXWCfaT5_0(.din(w_dff_B_u2z4JjPk5_0),.dout(w_dff_B_aUXWCfaT5_0),.clk(gclk));
	jdff dff_B_vSmmTJWj6_0(.din(w_dff_B_aUXWCfaT5_0),.dout(w_dff_B_vSmmTJWj6_0),.clk(gclk));
	jdff dff_B_4GQKI0Wq5_0(.din(w_dff_B_vSmmTJWj6_0),.dout(w_dff_B_4GQKI0Wq5_0),.clk(gclk));
	jdff dff_B_l749LOFF5_0(.din(w_dff_B_4GQKI0Wq5_0),.dout(w_dff_B_l749LOFF5_0),.clk(gclk));
	jdff dff_B_aRd4vaSr9_0(.din(w_dff_B_l749LOFF5_0),.dout(w_dff_B_aRd4vaSr9_0),.clk(gclk));
	jdff dff_B_vPSmcQff2_0(.din(w_dff_B_aRd4vaSr9_0),.dout(w_dff_B_vPSmcQff2_0),.clk(gclk));
	jdff dff_B_kNchVSOD4_0(.din(w_dff_B_vPSmcQff2_0),.dout(w_dff_B_kNchVSOD4_0),.clk(gclk));
	jdff dff_B_qYjdLf3P0_0(.din(w_dff_B_kNchVSOD4_0),.dout(w_dff_B_qYjdLf3P0_0),.clk(gclk));
	jdff dff_B_F0FQD6cg9_0(.din(w_dff_B_qYjdLf3P0_0),.dout(w_dff_B_F0FQD6cg9_0),.clk(gclk));
	jdff dff_B_hJIGDIrz4_0(.din(w_dff_B_F0FQD6cg9_0),.dout(w_dff_B_hJIGDIrz4_0),.clk(gclk));
	jdff dff_B_AR2FvIXN8_0(.din(w_dff_B_hJIGDIrz4_0),.dout(w_dff_B_AR2FvIXN8_0),.clk(gclk));
	jdff dff_B_d50zOTAp5_0(.din(w_dff_B_AR2FvIXN8_0),.dout(w_dff_B_d50zOTAp5_0),.clk(gclk));
	jdff dff_B_k7v2pxiZ3_0(.din(w_dff_B_d50zOTAp5_0),.dout(w_dff_B_k7v2pxiZ3_0),.clk(gclk));
	jdff dff_B_lRwxMITQ8_0(.din(w_dff_B_k7v2pxiZ3_0),.dout(w_dff_B_lRwxMITQ8_0),.clk(gclk));
	jdff dff_B_zex4fiO20_0(.din(w_dff_B_lRwxMITQ8_0),.dout(w_dff_B_zex4fiO20_0),.clk(gclk));
	jdff dff_B_97cjC2gG3_0(.din(w_dff_B_zex4fiO20_0),.dout(w_dff_B_97cjC2gG3_0),.clk(gclk));
	jdff dff_B_ubt9NPi78_0(.din(w_dff_B_97cjC2gG3_0),.dout(w_dff_B_ubt9NPi78_0),.clk(gclk));
	jdff dff_B_Y2DU5Z5c3_0(.din(w_dff_B_ubt9NPi78_0),.dout(w_dff_B_Y2DU5Z5c3_0),.clk(gclk));
	jdff dff_B_VULUXgp86_0(.din(w_dff_B_Y2DU5Z5c3_0),.dout(w_dff_B_VULUXgp86_0),.clk(gclk));
	jdff dff_B_Hg2syQxk9_0(.din(w_dff_B_VULUXgp86_0),.dout(w_dff_B_Hg2syQxk9_0),.clk(gclk));
	jdff dff_B_JB3M4uWh1_0(.din(w_dff_B_Hg2syQxk9_0),.dout(w_dff_B_JB3M4uWh1_0),.clk(gclk));
	jdff dff_B_aBle1NC62_0(.din(w_dff_B_JB3M4uWh1_0),.dout(w_dff_B_aBle1NC62_0),.clk(gclk));
	jdff dff_B_zM0TcW941_0(.din(w_dff_B_aBle1NC62_0),.dout(w_dff_B_zM0TcW941_0),.clk(gclk));
	jdff dff_B_n0oxOqpK1_0(.din(w_dff_B_zM0TcW941_0),.dout(w_dff_B_n0oxOqpK1_0),.clk(gclk));
	jdff dff_B_N8XFtalI6_0(.din(w_dff_B_n0oxOqpK1_0),.dout(w_dff_B_N8XFtalI6_0),.clk(gclk));
	jdff dff_B_OaRocCCV1_0(.din(w_dff_B_N8XFtalI6_0),.dout(w_dff_B_OaRocCCV1_0),.clk(gclk));
	jdff dff_B_Bha0PZ8T5_0(.din(w_dff_B_OaRocCCV1_0),.dout(w_dff_B_Bha0PZ8T5_0),.clk(gclk));
	jdff dff_B_bdyIpRd64_0(.din(w_dff_B_Bha0PZ8T5_0),.dout(w_dff_B_bdyIpRd64_0),.clk(gclk));
	jdff dff_B_PayoqlsK8_0(.din(w_dff_B_bdyIpRd64_0),.dout(w_dff_B_PayoqlsK8_0),.clk(gclk));
	jdff dff_B_cJe2QCEx9_0(.din(w_dff_B_PayoqlsK8_0),.dout(w_dff_B_cJe2QCEx9_0),.clk(gclk));
	jdff dff_B_OvBXG0gx8_0(.din(w_dff_B_cJe2QCEx9_0),.dout(w_dff_B_OvBXG0gx8_0),.clk(gclk));
	jdff dff_B_Dls3IOzT3_0(.din(w_dff_B_OvBXG0gx8_0),.dout(w_dff_B_Dls3IOzT3_0),.clk(gclk));
	jdff dff_B_gRUP5ac66_0(.din(w_dff_B_Dls3IOzT3_0),.dout(w_dff_B_gRUP5ac66_0),.clk(gclk));
	jdff dff_B_JWa0fYzz7_0(.din(w_dff_B_gRUP5ac66_0),.dout(w_dff_B_JWa0fYzz7_0),.clk(gclk));
	jdff dff_B_gfnlPPgT8_0(.din(w_dff_B_JWa0fYzz7_0),.dout(w_dff_B_gfnlPPgT8_0),.clk(gclk));
	jdff dff_B_X5fasANi6_0(.din(w_dff_B_gfnlPPgT8_0),.dout(w_dff_B_X5fasANi6_0),.clk(gclk));
	jdff dff_B_gELEVP791_0(.din(w_dff_B_X5fasANi6_0),.dout(w_dff_B_gELEVP791_0),.clk(gclk));
	jdff dff_B_4FyXF39X4_0(.din(w_dff_B_gELEVP791_0),.dout(w_dff_B_4FyXF39X4_0),.clk(gclk));
	jdff dff_B_JzUETrMd5_0(.din(w_dff_B_4FyXF39X4_0),.dout(w_dff_B_JzUETrMd5_0),.clk(gclk));
	jdff dff_B_ZMSgl2eg8_0(.din(w_dff_B_JzUETrMd5_0),.dout(w_dff_B_ZMSgl2eg8_0),.clk(gclk));
	jdff dff_B_arvvqOuV6_0(.din(w_dff_B_ZMSgl2eg8_0),.dout(w_dff_B_arvvqOuV6_0),.clk(gclk));
	jdff dff_B_IJFnLUlT7_0(.din(w_dff_B_arvvqOuV6_0),.dout(w_dff_B_IJFnLUlT7_0),.clk(gclk));
	jdff dff_B_OZzL7Krh5_0(.din(w_dff_B_IJFnLUlT7_0),.dout(w_dff_B_OZzL7Krh5_0),.clk(gclk));
	jdff dff_B_j68Ib33U5_0(.din(w_dff_B_OZzL7Krh5_0),.dout(w_dff_B_j68Ib33U5_0),.clk(gclk));
	jdff dff_B_6zFH5uQN4_0(.din(w_dff_B_j68Ib33U5_0),.dout(w_dff_B_6zFH5uQN4_0),.clk(gclk));
	jdff dff_B_hQxUX1WK5_0(.din(w_dff_B_6zFH5uQN4_0),.dout(w_dff_B_hQxUX1WK5_0),.clk(gclk));
	jdff dff_B_8itDHIDq3_0(.din(w_dff_B_hQxUX1WK5_0),.dout(w_dff_B_8itDHIDq3_0),.clk(gclk));
	jdff dff_B_oIn76kGK6_0(.din(w_dff_B_8itDHIDq3_0),.dout(w_dff_B_oIn76kGK6_0),.clk(gclk));
	jdff dff_B_xRqNo4PA0_0(.din(w_dff_B_oIn76kGK6_0),.dout(w_dff_B_xRqNo4PA0_0),.clk(gclk));
	jdff dff_B_UgChdVzk8_0(.din(w_dff_B_xRqNo4PA0_0),.dout(w_dff_B_UgChdVzk8_0),.clk(gclk));
	jdff dff_B_enyuX2n99_0(.din(w_dff_B_UgChdVzk8_0),.dout(w_dff_B_enyuX2n99_0),.clk(gclk));
	jdff dff_B_weeMWlHm2_0(.din(w_dff_B_enyuX2n99_0),.dout(w_dff_B_weeMWlHm2_0),.clk(gclk));
	jdff dff_B_Cp0yVbP13_0(.din(w_dff_B_weeMWlHm2_0),.dout(w_dff_B_Cp0yVbP13_0),.clk(gclk));
	jdff dff_B_SBebaV8n2_0(.din(w_dff_B_Cp0yVbP13_0),.dout(w_dff_B_SBebaV8n2_0),.clk(gclk));
	jdff dff_B_oqHghBrO3_0(.din(w_dff_B_SBebaV8n2_0),.dout(w_dff_B_oqHghBrO3_0),.clk(gclk));
	jdff dff_B_F0e8169s2_0(.din(w_dff_B_oqHghBrO3_0),.dout(w_dff_B_F0e8169s2_0),.clk(gclk));
	jdff dff_B_csu2yVde3_0(.din(w_dff_B_F0e8169s2_0),.dout(w_dff_B_csu2yVde3_0),.clk(gclk));
	jdff dff_B_Z7PCXxEK1_0(.din(w_dff_B_csu2yVde3_0),.dout(w_dff_B_Z7PCXxEK1_0),.clk(gclk));
	jdff dff_B_XMyPOCWG6_0(.din(w_dff_B_Z7PCXxEK1_0),.dout(w_dff_B_XMyPOCWG6_0),.clk(gclk));
	jdff dff_B_VlgJaTYI1_0(.din(w_dff_B_XMyPOCWG6_0),.dout(w_dff_B_VlgJaTYI1_0),.clk(gclk));
	jdff dff_B_rWJ1jfPs7_0(.din(w_dff_B_VlgJaTYI1_0),.dout(w_dff_B_rWJ1jfPs7_0),.clk(gclk));
	jdff dff_B_M7vRvPIA2_0(.din(w_dff_B_rWJ1jfPs7_0),.dout(w_dff_B_M7vRvPIA2_0),.clk(gclk));
	jdff dff_B_H52zktDU8_0(.din(n1096),.dout(w_dff_B_H52zktDU8_0),.clk(gclk));
	jdff dff_B_jXczRxPA9_0(.din(w_dff_B_H52zktDU8_0),.dout(w_dff_B_jXczRxPA9_0),.clk(gclk));
	jdff dff_B_qUOG4h1x1_0(.din(w_dff_B_jXczRxPA9_0),.dout(w_dff_B_qUOG4h1x1_0),.clk(gclk));
	jdff dff_B_o2BsuHd70_0(.din(w_dff_B_qUOG4h1x1_0),.dout(w_dff_B_o2BsuHd70_0),.clk(gclk));
	jdff dff_B_Uy391QM83_0(.din(w_dff_B_o2BsuHd70_0),.dout(w_dff_B_Uy391QM83_0),.clk(gclk));
	jdff dff_B_yWsdAQQN4_0(.din(w_dff_B_Uy391QM83_0),.dout(w_dff_B_yWsdAQQN4_0),.clk(gclk));
	jdff dff_B_hSS5iuJ31_0(.din(w_dff_B_yWsdAQQN4_0),.dout(w_dff_B_hSS5iuJ31_0),.clk(gclk));
	jdff dff_B_QRoVHLTH5_0(.din(w_dff_B_hSS5iuJ31_0),.dout(w_dff_B_QRoVHLTH5_0),.clk(gclk));
	jdff dff_B_asFz572A4_0(.din(w_dff_B_QRoVHLTH5_0),.dout(w_dff_B_asFz572A4_0),.clk(gclk));
	jdff dff_B_Q17GLZcN7_0(.din(w_dff_B_asFz572A4_0),.dout(w_dff_B_Q17GLZcN7_0),.clk(gclk));
	jdff dff_B_enQSSbSI4_0(.din(w_dff_B_Q17GLZcN7_0),.dout(w_dff_B_enQSSbSI4_0),.clk(gclk));
	jdff dff_B_7HO00lui4_0(.din(w_dff_B_enQSSbSI4_0),.dout(w_dff_B_7HO00lui4_0),.clk(gclk));
	jdff dff_B_GRsMJyys5_0(.din(w_dff_B_7HO00lui4_0),.dout(w_dff_B_GRsMJyys5_0),.clk(gclk));
	jdff dff_B_oYeez4Mp4_0(.din(w_dff_B_GRsMJyys5_0),.dout(w_dff_B_oYeez4Mp4_0),.clk(gclk));
	jdff dff_B_OCCOYnUR6_0(.din(w_dff_B_oYeez4Mp4_0),.dout(w_dff_B_OCCOYnUR6_0),.clk(gclk));
	jdff dff_B_XykJq9xE8_0(.din(w_dff_B_OCCOYnUR6_0),.dout(w_dff_B_XykJq9xE8_0),.clk(gclk));
	jdff dff_B_pSQIn4d31_0(.din(w_dff_B_XykJq9xE8_0),.dout(w_dff_B_pSQIn4d31_0),.clk(gclk));
	jdff dff_B_mrE4b4hj0_0(.din(w_dff_B_pSQIn4d31_0),.dout(w_dff_B_mrE4b4hj0_0),.clk(gclk));
	jdff dff_B_FEC12HEQ4_0(.din(w_dff_B_mrE4b4hj0_0),.dout(w_dff_B_FEC12HEQ4_0),.clk(gclk));
	jdff dff_B_UkKKrox99_0(.din(w_dff_B_FEC12HEQ4_0),.dout(w_dff_B_UkKKrox99_0),.clk(gclk));
	jdff dff_B_rBIY3iHI6_0(.din(w_dff_B_UkKKrox99_0),.dout(w_dff_B_rBIY3iHI6_0),.clk(gclk));
	jdff dff_B_akrvIWaH5_0(.din(w_dff_B_rBIY3iHI6_0),.dout(w_dff_B_akrvIWaH5_0),.clk(gclk));
	jdff dff_B_axc63lYQ5_0(.din(w_dff_B_akrvIWaH5_0),.dout(w_dff_B_axc63lYQ5_0),.clk(gclk));
	jdff dff_B_jgXX1eQ82_0(.din(w_dff_B_axc63lYQ5_0),.dout(w_dff_B_jgXX1eQ82_0),.clk(gclk));
	jdff dff_B_PcGZrH3T8_0(.din(w_dff_B_jgXX1eQ82_0),.dout(w_dff_B_PcGZrH3T8_0),.clk(gclk));
	jdff dff_B_f3795ANB1_0(.din(w_dff_B_PcGZrH3T8_0),.dout(w_dff_B_f3795ANB1_0),.clk(gclk));
	jdff dff_B_FvBLlsaI2_0(.din(w_dff_B_f3795ANB1_0),.dout(w_dff_B_FvBLlsaI2_0),.clk(gclk));
	jdff dff_B_eAwVNVwG9_0(.din(w_dff_B_FvBLlsaI2_0),.dout(w_dff_B_eAwVNVwG9_0),.clk(gclk));
	jdff dff_B_ziZwOSYL3_0(.din(w_dff_B_eAwVNVwG9_0),.dout(w_dff_B_ziZwOSYL3_0),.clk(gclk));
	jdff dff_B_yPdosjHg9_0(.din(w_dff_B_ziZwOSYL3_0),.dout(w_dff_B_yPdosjHg9_0),.clk(gclk));
	jdff dff_B_wymPk2af8_0(.din(w_dff_B_yPdosjHg9_0),.dout(w_dff_B_wymPk2af8_0),.clk(gclk));
	jdff dff_B_R0WSs6Kl2_0(.din(w_dff_B_wymPk2af8_0),.dout(w_dff_B_R0WSs6Kl2_0),.clk(gclk));
	jdff dff_B_pvkvl9fo4_0(.din(w_dff_B_R0WSs6Kl2_0),.dout(w_dff_B_pvkvl9fo4_0),.clk(gclk));
	jdff dff_B_aitfsw0Y0_0(.din(w_dff_B_pvkvl9fo4_0),.dout(w_dff_B_aitfsw0Y0_0),.clk(gclk));
	jdff dff_B_7g7gUE3u9_0(.din(w_dff_B_aitfsw0Y0_0),.dout(w_dff_B_7g7gUE3u9_0),.clk(gclk));
	jdff dff_B_tPg7xZrw4_0(.din(w_dff_B_7g7gUE3u9_0),.dout(w_dff_B_tPg7xZrw4_0),.clk(gclk));
	jdff dff_B_iBS0wxeZ6_0(.din(w_dff_B_tPg7xZrw4_0),.dout(w_dff_B_iBS0wxeZ6_0),.clk(gclk));
	jdff dff_B_jjVcmA4s4_0(.din(w_dff_B_iBS0wxeZ6_0),.dout(w_dff_B_jjVcmA4s4_0),.clk(gclk));
	jdff dff_B_WQjdV6h15_0(.din(w_dff_B_jjVcmA4s4_0),.dout(w_dff_B_WQjdV6h15_0),.clk(gclk));
	jdff dff_B_CZLR0oVD8_0(.din(w_dff_B_WQjdV6h15_0),.dout(w_dff_B_CZLR0oVD8_0),.clk(gclk));
	jdff dff_B_OySqiWIz0_0(.din(w_dff_B_CZLR0oVD8_0),.dout(w_dff_B_OySqiWIz0_0),.clk(gclk));
	jdff dff_B_LEjgoI5o0_0(.din(w_dff_B_OySqiWIz0_0),.dout(w_dff_B_LEjgoI5o0_0),.clk(gclk));
	jdff dff_B_4WD5y66k1_0(.din(w_dff_B_LEjgoI5o0_0),.dout(w_dff_B_4WD5y66k1_0),.clk(gclk));
	jdff dff_B_skvqbat10_0(.din(w_dff_B_4WD5y66k1_0),.dout(w_dff_B_skvqbat10_0),.clk(gclk));
	jdff dff_B_058xrlB73_0(.din(w_dff_B_skvqbat10_0),.dout(w_dff_B_058xrlB73_0),.clk(gclk));
	jdff dff_B_C1xAoHo36_0(.din(w_dff_B_058xrlB73_0),.dout(w_dff_B_C1xAoHo36_0),.clk(gclk));
	jdff dff_B_SP7zVPQj4_0(.din(w_dff_B_C1xAoHo36_0),.dout(w_dff_B_SP7zVPQj4_0),.clk(gclk));
	jdff dff_B_eIXA1Ojg3_0(.din(w_dff_B_SP7zVPQj4_0),.dout(w_dff_B_eIXA1Ojg3_0),.clk(gclk));
	jdff dff_B_VZFoyD096_0(.din(w_dff_B_eIXA1Ojg3_0),.dout(w_dff_B_VZFoyD096_0),.clk(gclk));
	jdff dff_B_UXRrNooA3_0(.din(w_dff_B_VZFoyD096_0),.dout(w_dff_B_UXRrNooA3_0),.clk(gclk));
	jdff dff_B_mx6QzdhE8_0(.din(w_dff_B_UXRrNooA3_0),.dout(w_dff_B_mx6QzdhE8_0),.clk(gclk));
	jdff dff_B_lo3ftZGt8_0(.din(w_dff_B_mx6QzdhE8_0),.dout(w_dff_B_lo3ftZGt8_0),.clk(gclk));
	jdff dff_B_wJjz88Px4_0(.din(w_dff_B_lo3ftZGt8_0),.dout(w_dff_B_wJjz88Px4_0),.clk(gclk));
	jdff dff_B_RcaFbYO23_0(.din(w_dff_B_wJjz88Px4_0),.dout(w_dff_B_RcaFbYO23_0),.clk(gclk));
	jdff dff_B_2dC1oWKF0_0(.din(w_dff_B_RcaFbYO23_0),.dout(w_dff_B_2dC1oWKF0_0),.clk(gclk));
	jdff dff_B_9Syh3jcY8_0(.din(w_dff_B_2dC1oWKF0_0),.dout(w_dff_B_9Syh3jcY8_0),.clk(gclk));
	jdff dff_B_RGCJIKH71_0(.din(w_dff_B_9Syh3jcY8_0),.dout(w_dff_B_RGCJIKH71_0),.clk(gclk));
	jdff dff_B_Ysl7iKtY3_0(.din(w_dff_B_RGCJIKH71_0),.dout(w_dff_B_Ysl7iKtY3_0),.clk(gclk));
	jdff dff_B_6dFmWfct1_0(.din(w_dff_B_Ysl7iKtY3_0),.dout(w_dff_B_6dFmWfct1_0),.clk(gclk));
	jdff dff_B_Ctcu9det7_0(.din(w_dff_B_6dFmWfct1_0),.dout(w_dff_B_Ctcu9det7_0),.clk(gclk));
	jdff dff_B_rdyuhxwe7_0(.din(w_dff_B_Ctcu9det7_0),.dout(w_dff_B_rdyuhxwe7_0),.clk(gclk));
	jdff dff_B_o6lmB5kz9_0(.din(w_dff_B_rdyuhxwe7_0),.dout(w_dff_B_o6lmB5kz9_0),.clk(gclk));
	jdff dff_B_7igJX8uc5_0(.din(w_dff_B_o6lmB5kz9_0),.dout(w_dff_B_7igJX8uc5_0),.clk(gclk));
	jdff dff_B_J1cj6hri7_0(.din(w_dff_B_7igJX8uc5_0),.dout(w_dff_B_J1cj6hri7_0),.clk(gclk));
	jdff dff_B_vqBhSY1U0_0(.din(w_dff_B_J1cj6hri7_0),.dout(w_dff_B_vqBhSY1U0_0),.clk(gclk));
	jdff dff_B_2pDodbty5_0(.din(w_dff_B_vqBhSY1U0_0),.dout(w_dff_B_2pDodbty5_0),.clk(gclk));
	jdff dff_B_r6L3mB699_0(.din(w_dff_B_2pDodbty5_0),.dout(w_dff_B_r6L3mB699_0),.clk(gclk));
	jdff dff_B_hUioI3XI0_0(.din(w_dff_B_r6L3mB699_0),.dout(w_dff_B_hUioI3XI0_0),.clk(gclk));
	jdff dff_B_h7a50YUe6_0(.din(w_dff_B_hUioI3XI0_0),.dout(w_dff_B_h7a50YUe6_0),.clk(gclk));
	jdff dff_B_R39OpCJ14_0(.din(w_dff_B_h7a50YUe6_0),.dout(w_dff_B_R39OpCJ14_0),.clk(gclk));
	jdff dff_B_R1MBCPqW0_0(.din(w_dff_B_R39OpCJ14_0),.dout(w_dff_B_R1MBCPqW0_0),.clk(gclk));
	jdff dff_B_ayKbiZxB8_0(.din(w_dff_B_R1MBCPqW0_0),.dout(w_dff_B_ayKbiZxB8_0),.clk(gclk));
	jdff dff_B_mI9qiqLD3_0(.din(w_dff_B_ayKbiZxB8_0),.dout(w_dff_B_mI9qiqLD3_0),.clk(gclk));
	jdff dff_B_XQ5VNEIN0_0(.din(w_dff_B_mI9qiqLD3_0),.dout(w_dff_B_XQ5VNEIN0_0),.clk(gclk));
	jdff dff_B_olB7Nf1l5_0(.din(w_dff_B_XQ5VNEIN0_0),.dout(w_dff_B_olB7Nf1l5_0),.clk(gclk));
	jdff dff_B_Z8bPN8lA7_0(.din(w_dff_B_olB7Nf1l5_0),.dout(w_dff_B_Z8bPN8lA7_0),.clk(gclk));
	jdff dff_B_a4ImkX0F1_0(.din(w_dff_B_Z8bPN8lA7_0),.dout(w_dff_B_a4ImkX0F1_0),.clk(gclk));
	jdff dff_B_lDMaNvAY8_0(.din(w_dff_B_a4ImkX0F1_0),.dout(w_dff_B_lDMaNvAY8_0),.clk(gclk));
	jdff dff_B_PPVk8cTU1_0(.din(w_dff_B_lDMaNvAY8_0),.dout(w_dff_B_PPVk8cTU1_0),.clk(gclk));
	jdff dff_B_f06G2IVk1_0(.din(w_dff_B_PPVk8cTU1_0),.dout(w_dff_B_f06G2IVk1_0),.clk(gclk));
	jdff dff_B_4G0r33FD6_0(.din(w_dff_B_f06G2IVk1_0),.dout(w_dff_B_4G0r33FD6_0),.clk(gclk));
	jdff dff_B_Uo9sTI2d6_0(.din(w_dff_B_4G0r33FD6_0),.dout(w_dff_B_Uo9sTI2d6_0),.clk(gclk));
	jdff dff_B_ceXLxFiL2_0(.din(w_dff_B_Uo9sTI2d6_0),.dout(w_dff_B_ceXLxFiL2_0),.clk(gclk));
	jdff dff_B_3McNI1BL0_0(.din(w_dff_B_ceXLxFiL2_0),.dout(w_dff_B_3McNI1BL0_0),.clk(gclk));
	jdff dff_B_zDAuNtQN3_0(.din(w_dff_B_3McNI1BL0_0),.dout(w_dff_B_zDAuNtQN3_0),.clk(gclk));
	jdff dff_B_YzTcwtiy2_0(.din(w_dff_B_zDAuNtQN3_0),.dout(w_dff_B_YzTcwtiy2_0),.clk(gclk));
	jdff dff_B_JGsJ6wVA3_0(.din(w_dff_B_YzTcwtiy2_0),.dout(w_dff_B_JGsJ6wVA3_0),.clk(gclk));
	jdff dff_B_8Y8lLYyy9_0(.din(w_dff_B_JGsJ6wVA3_0),.dout(w_dff_B_8Y8lLYyy9_0),.clk(gclk));
	jdff dff_B_D5b77H9w0_0(.din(w_dff_B_8Y8lLYyy9_0),.dout(w_dff_B_D5b77H9w0_0),.clk(gclk));
	jdff dff_B_1B8zarzA9_0(.din(w_dff_B_D5b77H9w0_0),.dout(w_dff_B_1B8zarzA9_0),.clk(gclk));
	jdff dff_B_TEwD6oFa2_0(.din(w_dff_B_1B8zarzA9_0),.dout(w_dff_B_TEwD6oFa2_0),.clk(gclk));
	jdff dff_B_uBe9ALIw3_0(.din(w_dff_B_TEwD6oFa2_0),.dout(w_dff_B_uBe9ALIw3_0),.clk(gclk));
	jdff dff_B_g89ZXUxF9_0(.din(w_dff_B_uBe9ALIw3_0),.dout(w_dff_B_g89ZXUxF9_0),.clk(gclk));
	jdff dff_B_HQ3uB9VM1_0(.din(w_dff_B_g89ZXUxF9_0),.dout(w_dff_B_HQ3uB9VM1_0),.clk(gclk));
	jdff dff_B_mtJwnctp2_0(.din(w_dff_B_HQ3uB9VM1_0),.dout(w_dff_B_mtJwnctp2_0),.clk(gclk));
	jdff dff_B_aCmArjJb1_0(.din(w_dff_B_mtJwnctp2_0),.dout(w_dff_B_aCmArjJb1_0),.clk(gclk));
	jdff dff_B_sQImK0oE6_0(.din(w_dff_B_aCmArjJb1_0),.dout(w_dff_B_sQImK0oE6_0),.clk(gclk));
	jdff dff_B_yvHaVn4I2_0(.din(w_dff_B_sQImK0oE6_0),.dout(w_dff_B_yvHaVn4I2_0),.clk(gclk));
	jdff dff_B_2adiK2LN7_0(.din(w_dff_B_yvHaVn4I2_0),.dout(w_dff_B_2adiK2LN7_0),.clk(gclk));
	jdff dff_B_pTGyYuFZ4_0(.din(w_dff_B_2adiK2LN7_0),.dout(w_dff_B_pTGyYuFZ4_0),.clk(gclk));
	jdff dff_B_7LYmdE161_0(.din(w_dff_B_pTGyYuFZ4_0),.dout(w_dff_B_7LYmdE161_0),.clk(gclk));
	jdff dff_B_gH0gpuAR2_0(.din(w_dff_B_7LYmdE161_0),.dout(w_dff_B_gH0gpuAR2_0),.clk(gclk));
	jdff dff_B_5l3KvKCB6_0(.din(w_dff_B_gH0gpuAR2_0),.dout(w_dff_B_5l3KvKCB6_0),.clk(gclk));
	jdff dff_B_ONbJNmru1_0(.din(w_dff_B_5l3KvKCB6_0),.dout(w_dff_B_ONbJNmru1_0),.clk(gclk));
	jdff dff_B_8YOxLtd12_0(.din(w_dff_B_ONbJNmru1_0),.dout(w_dff_B_8YOxLtd12_0),.clk(gclk));
	jdff dff_B_bda9rMd55_0(.din(w_dff_B_8YOxLtd12_0),.dout(w_dff_B_bda9rMd55_0),.clk(gclk));
	jdff dff_B_zBiJ20cc7_0(.din(w_dff_B_bda9rMd55_0),.dout(w_dff_B_zBiJ20cc7_0),.clk(gclk));
	jdff dff_B_yw4Ht0p46_0(.din(w_dff_B_zBiJ20cc7_0),.dout(w_dff_B_yw4Ht0p46_0),.clk(gclk));
	jdff dff_B_QKXuQfY94_0(.din(w_dff_B_yw4Ht0p46_0),.dout(w_dff_B_QKXuQfY94_0),.clk(gclk));
	jdff dff_B_xkcW9Ldj2_0(.din(w_dff_B_QKXuQfY94_0),.dout(w_dff_B_xkcW9Ldj2_0),.clk(gclk));
	jdff dff_B_YSC6YNxi9_0(.din(w_dff_B_xkcW9Ldj2_0),.dout(w_dff_B_YSC6YNxi9_0),.clk(gclk));
	jdff dff_B_ht3ZNn0X2_0(.din(w_dff_B_YSC6YNxi9_0),.dout(w_dff_B_ht3ZNn0X2_0),.clk(gclk));
	jdff dff_B_2y13gvOT4_0(.din(w_dff_B_ht3ZNn0X2_0),.dout(w_dff_B_2y13gvOT4_0),.clk(gclk));
	jdff dff_B_WHfWUouE0_0(.din(w_dff_B_2y13gvOT4_0),.dout(w_dff_B_WHfWUouE0_0),.clk(gclk));
	jdff dff_B_VaxtxZZ68_0(.din(w_dff_B_WHfWUouE0_0),.dout(w_dff_B_VaxtxZZ68_0),.clk(gclk));
	jdff dff_B_8kTQRZpM2_0(.din(w_dff_B_VaxtxZZ68_0),.dout(w_dff_B_8kTQRZpM2_0),.clk(gclk));
	jdff dff_B_sLqCAoEz9_0(.din(w_dff_B_8kTQRZpM2_0),.dout(w_dff_B_sLqCAoEz9_0),.clk(gclk));
	jdff dff_B_f5k0RJ456_0(.din(w_dff_B_sLqCAoEz9_0),.dout(w_dff_B_f5k0RJ456_0),.clk(gclk));
	jdff dff_B_uvwQYYe33_0(.din(n1102),.dout(w_dff_B_uvwQYYe33_0),.clk(gclk));
	jdff dff_B_PRHQDVjY9_0(.din(w_dff_B_uvwQYYe33_0),.dout(w_dff_B_PRHQDVjY9_0),.clk(gclk));
	jdff dff_B_NfGs6jPv4_0(.din(w_dff_B_PRHQDVjY9_0),.dout(w_dff_B_NfGs6jPv4_0),.clk(gclk));
	jdff dff_B_br24ce4R8_0(.din(w_dff_B_NfGs6jPv4_0),.dout(w_dff_B_br24ce4R8_0),.clk(gclk));
	jdff dff_B_PfkViLOG8_0(.din(w_dff_B_br24ce4R8_0),.dout(w_dff_B_PfkViLOG8_0),.clk(gclk));
	jdff dff_B_M3EDA1xX7_0(.din(w_dff_B_PfkViLOG8_0),.dout(w_dff_B_M3EDA1xX7_0),.clk(gclk));
	jdff dff_B_Dv7mLFTF0_0(.din(w_dff_B_M3EDA1xX7_0),.dout(w_dff_B_Dv7mLFTF0_0),.clk(gclk));
	jdff dff_B_lWCsIlXA3_0(.din(w_dff_B_Dv7mLFTF0_0),.dout(w_dff_B_lWCsIlXA3_0),.clk(gclk));
	jdff dff_B_b6Ptx8On0_0(.din(w_dff_B_lWCsIlXA3_0),.dout(w_dff_B_b6Ptx8On0_0),.clk(gclk));
	jdff dff_B_JqoYJHNx4_0(.din(w_dff_B_b6Ptx8On0_0),.dout(w_dff_B_JqoYJHNx4_0),.clk(gclk));
	jdff dff_B_QUgVbbHD2_0(.din(w_dff_B_JqoYJHNx4_0),.dout(w_dff_B_QUgVbbHD2_0),.clk(gclk));
	jdff dff_B_tAlzt0PE9_0(.din(w_dff_B_QUgVbbHD2_0),.dout(w_dff_B_tAlzt0PE9_0),.clk(gclk));
	jdff dff_B_zFlF74da1_0(.din(w_dff_B_tAlzt0PE9_0),.dout(w_dff_B_zFlF74da1_0),.clk(gclk));
	jdff dff_B_KfmETYUc9_0(.din(w_dff_B_zFlF74da1_0),.dout(w_dff_B_KfmETYUc9_0),.clk(gclk));
	jdff dff_B_h9TbfxFo9_0(.din(w_dff_B_KfmETYUc9_0),.dout(w_dff_B_h9TbfxFo9_0),.clk(gclk));
	jdff dff_B_8yg7ndMK2_0(.din(w_dff_B_h9TbfxFo9_0),.dout(w_dff_B_8yg7ndMK2_0),.clk(gclk));
	jdff dff_B_3MpH5j2X5_0(.din(w_dff_B_8yg7ndMK2_0),.dout(w_dff_B_3MpH5j2X5_0),.clk(gclk));
	jdff dff_B_EWl41ZHf9_0(.din(w_dff_B_3MpH5j2X5_0),.dout(w_dff_B_EWl41ZHf9_0),.clk(gclk));
	jdff dff_B_XInmM5uu3_0(.din(w_dff_B_EWl41ZHf9_0),.dout(w_dff_B_XInmM5uu3_0),.clk(gclk));
	jdff dff_B_dIrbEeRa3_0(.din(w_dff_B_XInmM5uu3_0),.dout(w_dff_B_dIrbEeRa3_0),.clk(gclk));
	jdff dff_B_gBbA07bB9_0(.din(w_dff_B_dIrbEeRa3_0),.dout(w_dff_B_gBbA07bB9_0),.clk(gclk));
	jdff dff_B_pghgJ4ba8_0(.din(w_dff_B_gBbA07bB9_0),.dout(w_dff_B_pghgJ4ba8_0),.clk(gclk));
	jdff dff_B_Q37UsApI4_0(.din(w_dff_B_pghgJ4ba8_0),.dout(w_dff_B_Q37UsApI4_0),.clk(gclk));
	jdff dff_B_yQhmpA628_0(.din(w_dff_B_Q37UsApI4_0),.dout(w_dff_B_yQhmpA628_0),.clk(gclk));
	jdff dff_B_viVkT27L6_0(.din(w_dff_B_yQhmpA628_0),.dout(w_dff_B_viVkT27L6_0),.clk(gclk));
	jdff dff_B_XxWJ1Jxq1_0(.din(w_dff_B_viVkT27L6_0),.dout(w_dff_B_XxWJ1Jxq1_0),.clk(gclk));
	jdff dff_B_qJ6EI6jf5_0(.din(w_dff_B_XxWJ1Jxq1_0),.dout(w_dff_B_qJ6EI6jf5_0),.clk(gclk));
	jdff dff_B_OrBgQSXt0_0(.din(w_dff_B_qJ6EI6jf5_0),.dout(w_dff_B_OrBgQSXt0_0),.clk(gclk));
	jdff dff_B_949NfNXB3_0(.din(w_dff_B_OrBgQSXt0_0),.dout(w_dff_B_949NfNXB3_0),.clk(gclk));
	jdff dff_B_EZeSEKlo9_0(.din(w_dff_B_949NfNXB3_0),.dout(w_dff_B_EZeSEKlo9_0),.clk(gclk));
	jdff dff_B_RkqjMSOq9_0(.din(w_dff_B_EZeSEKlo9_0),.dout(w_dff_B_RkqjMSOq9_0),.clk(gclk));
	jdff dff_B_Mh3FBitm2_0(.din(w_dff_B_RkqjMSOq9_0),.dout(w_dff_B_Mh3FBitm2_0),.clk(gclk));
	jdff dff_B_Na2H7pV40_0(.din(w_dff_B_Mh3FBitm2_0),.dout(w_dff_B_Na2H7pV40_0),.clk(gclk));
	jdff dff_B_YtrVJamn6_0(.din(w_dff_B_Na2H7pV40_0),.dout(w_dff_B_YtrVJamn6_0),.clk(gclk));
	jdff dff_B_YYP0CtYA1_0(.din(w_dff_B_YtrVJamn6_0),.dout(w_dff_B_YYP0CtYA1_0),.clk(gclk));
	jdff dff_B_d6p7MoRg9_0(.din(w_dff_B_YYP0CtYA1_0),.dout(w_dff_B_d6p7MoRg9_0),.clk(gclk));
	jdff dff_B_8kAJQYO34_0(.din(w_dff_B_d6p7MoRg9_0),.dout(w_dff_B_8kAJQYO34_0),.clk(gclk));
	jdff dff_B_qH5oY8uJ3_0(.din(w_dff_B_8kAJQYO34_0),.dout(w_dff_B_qH5oY8uJ3_0),.clk(gclk));
	jdff dff_B_D5Uc1jHX5_0(.din(w_dff_B_qH5oY8uJ3_0),.dout(w_dff_B_D5Uc1jHX5_0),.clk(gclk));
	jdff dff_B_oFWzUzBP3_0(.din(w_dff_B_D5Uc1jHX5_0),.dout(w_dff_B_oFWzUzBP3_0),.clk(gclk));
	jdff dff_B_xqY3nI2K4_0(.din(w_dff_B_oFWzUzBP3_0),.dout(w_dff_B_xqY3nI2K4_0),.clk(gclk));
	jdff dff_B_OdI2Kmp07_0(.din(w_dff_B_xqY3nI2K4_0),.dout(w_dff_B_OdI2Kmp07_0),.clk(gclk));
	jdff dff_B_hjy5hvL31_0(.din(w_dff_B_OdI2Kmp07_0),.dout(w_dff_B_hjy5hvL31_0),.clk(gclk));
	jdff dff_B_tO9ZQHds9_0(.din(w_dff_B_hjy5hvL31_0),.dout(w_dff_B_tO9ZQHds9_0),.clk(gclk));
	jdff dff_B_XQ6nkice2_0(.din(w_dff_B_tO9ZQHds9_0),.dout(w_dff_B_XQ6nkice2_0),.clk(gclk));
	jdff dff_B_255O0Gm10_0(.din(w_dff_B_XQ6nkice2_0),.dout(w_dff_B_255O0Gm10_0),.clk(gclk));
	jdff dff_B_xkVcMmOa7_0(.din(w_dff_B_255O0Gm10_0),.dout(w_dff_B_xkVcMmOa7_0),.clk(gclk));
	jdff dff_B_3AGfhD7j7_0(.din(w_dff_B_xkVcMmOa7_0),.dout(w_dff_B_3AGfhD7j7_0),.clk(gclk));
	jdff dff_B_iAB8pE324_0(.din(w_dff_B_3AGfhD7j7_0),.dout(w_dff_B_iAB8pE324_0),.clk(gclk));
	jdff dff_B_0R0K3Tct8_0(.din(w_dff_B_iAB8pE324_0),.dout(w_dff_B_0R0K3Tct8_0),.clk(gclk));
	jdff dff_B_myEnWWZf3_0(.din(w_dff_B_0R0K3Tct8_0),.dout(w_dff_B_myEnWWZf3_0),.clk(gclk));
	jdff dff_B_ALKRB9Qx1_0(.din(w_dff_B_myEnWWZf3_0),.dout(w_dff_B_ALKRB9Qx1_0),.clk(gclk));
	jdff dff_B_w5qCJn1V6_0(.din(w_dff_B_ALKRB9Qx1_0),.dout(w_dff_B_w5qCJn1V6_0),.clk(gclk));
	jdff dff_B_4vYjZtvV4_0(.din(w_dff_B_w5qCJn1V6_0),.dout(w_dff_B_4vYjZtvV4_0),.clk(gclk));
	jdff dff_B_JW8XbCeJ8_0(.din(w_dff_B_4vYjZtvV4_0),.dout(w_dff_B_JW8XbCeJ8_0),.clk(gclk));
	jdff dff_B_1NVcs1eF0_0(.din(w_dff_B_JW8XbCeJ8_0),.dout(w_dff_B_1NVcs1eF0_0),.clk(gclk));
	jdff dff_B_XpuqO2R07_0(.din(w_dff_B_1NVcs1eF0_0),.dout(w_dff_B_XpuqO2R07_0),.clk(gclk));
	jdff dff_B_9YuaLM9C6_0(.din(w_dff_B_XpuqO2R07_0),.dout(w_dff_B_9YuaLM9C6_0),.clk(gclk));
	jdff dff_B_MXoq1Ttp7_0(.din(w_dff_B_9YuaLM9C6_0),.dout(w_dff_B_MXoq1Ttp7_0),.clk(gclk));
	jdff dff_B_qGiSvxQb7_0(.din(w_dff_B_MXoq1Ttp7_0),.dout(w_dff_B_qGiSvxQb7_0),.clk(gclk));
	jdff dff_B_ENTmt6wu3_0(.din(w_dff_B_qGiSvxQb7_0),.dout(w_dff_B_ENTmt6wu3_0),.clk(gclk));
	jdff dff_B_LEA0bSTb9_0(.din(w_dff_B_ENTmt6wu3_0),.dout(w_dff_B_LEA0bSTb9_0),.clk(gclk));
	jdff dff_B_hy3o6oGJ7_0(.din(w_dff_B_LEA0bSTb9_0),.dout(w_dff_B_hy3o6oGJ7_0),.clk(gclk));
	jdff dff_B_bOmHALdH6_0(.din(w_dff_B_hy3o6oGJ7_0),.dout(w_dff_B_bOmHALdH6_0),.clk(gclk));
	jdff dff_B_lEZK15qY6_0(.din(w_dff_B_bOmHALdH6_0),.dout(w_dff_B_lEZK15qY6_0),.clk(gclk));
	jdff dff_B_qSxc1DSk1_0(.din(w_dff_B_lEZK15qY6_0),.dout(w_dff_B_qSxc1DSk1_0),.clk(gclk));
	jdff dff_B_ctoUowCc3_0(.din(w_dff_B_qSxc1DSk1_0),.dout(w_dff_B_ctoUowCc3_0),.clk(gclk));
	jdff dff_B_m3x6gj4X9_0(.din(w_dff_B_ctoUowCc3_0),.dout(w_dff_B_m3x6gj4X9_0),.clk(gclk));
	jdff dff_B_Uo2YVoss8_0(.din(w_dff_B_m3x6gj4X9_0),.dout(w_dff_B_Uo2YVoss8_0),.clk(gclk));
	jdff dff_B_GjpHOfA39_0(.din(w_dff_B_Uo2YVoss8_0),.dout(w_dff_B_GjpHOfA39_0),.clk(gclk));
	jdff dff_B_XejYHmwb3_0(.din(w_dff_B_GjpHOfA39_0),.dout(w_dff_B_XejYHmwb3_0),.clk(gclk));
	jdff dff_B_q3JTuYo19_0(.din(w_dff_B_XejYHmwb3_0),.dout(w_dff_B_q3JTuYo19_0),.clk(gclk));
	jdff dff_B_3NMrET7T2_0(.din(w_dff_B_q3JTuYo19_0),.dout(w_dff_B_3NMrET7T2_0),.clk(gclk));
	jdff dff_B_Q3ZifXet2_0(.din(w_dff_B_3NMrET7T2_0),.dout(w_dff_B_Q3ZifXet2_0),.clk(gclk));
	jdff dff_B_zd7nAWJf9_0(.din(w_dff_B_Q3ZifXet2_0),.dout(w_dff_B_zd7nAWJf9_0),.clk(gclk));
	jdff dff_B_B7UsuSFP8_0(.din(w_dff_B_zd7nAWJf9_0),.dout(w_dff_B_B7UsuSFP8_0),.clk(gclk));
	jdff dff_B_xds5KlN45_0(.din(w_dff_B_B7UsuSFP8_0),.dout(w_dff_B_xds5KlN45_0),.clk(gclk));
	jdff dff_B_Xk0JZCvB8_0(.din(w_dff_B_xds5KlN45_0),.dout(w_dff_B_Xk0JZCvB8_0),.clk(gclk));
	jdff dff_B_J7YFGtA00_0(.din(w_dff_B_Xk0JZCvB8_0),.dout(w_dff_B_J7YFGtA00_0),.clk(gclk));
	jdff dff_B_bv29g9Jy1_0(.din(w_dff_B_J7YFGtA00_0),.dout(w_dff_B_bv29g9Jy1_0),.clk(gclk));
	jdff dff_B_lZGlEFem2_0(.din(w_dff_B_bv29g9Jy1_0),.dout(w_dff_B_lZGlEFem2_0),.clk(gclk));
	jdff dff_B_FQSNxKtS7_0(.din(w_dff_B_lZGlEFem2_0),.dout(w_dff_B_FQSNxKtS7_0),.clk(gclk));
	jdff dff_B_Hvq6Grez2_0(.din(w_dff_B_FQSNxKtS7_0),.dout(w_dff_B_Hvq6Grez2_0),.clk(gclk));
	jdff dff_B_TcFL9nsw1_0(.din(w_dff_B_Hvq6Grez2_0),.dout(w_dff_B_TcFL9nsw1_0),.clk(gclk));
	jdff dff_B_xRZ7eL2I9_0(.din(w_dff_B_TcFL9nsw1_0),.dout(w_dff_B_xRZ7eL2I9_0),.clk(gclk));
	jdff dff_B_4uVeLXgT1_0(.din(w_dff_B_xRZ7eL2I9_0),.dout(w_dff_B_4uVeLXgT1_0),.clk(gclk));
	jdff dff_B_S1hPxKk54_0(.din(w_dff_B_4uVeLXgT1_0),.dout(w_dff_B_S1hPxKk54_0),.clk(gclk));
	jdff dff_B_pQEcvPJv2_0(.din(w_dff_B_S1hPxKk54_0),.dout(w_dff_B_pQEcvPJv2_0),.clk(gclk));
	jdff dff_B_NHJIqKwT4_0(.din(w_dff_B_pQEcvPJv2_0),.dout(w_dff_B_NHJIqKwT4_0),.clk(gclk));
	jdff dff_B_64vqJbq99_0(.din(w_dff_B_NHJIqKwT4_0),.dout(w_dff_B_64vqJbq99_0),.clk(gclk));
	jdff dff_B_zcyh6tyj7_0(.din(w_dff_B_64vqJbq99_0),.dout(w_dff_B_zcyh6tyj7_0),.clk(gclk));
	jdff dff_B_OGYbucAE2_0(.din(w_dff_B_zcyh6tyj7_0),.dout(w_dff_B_OGYbucAE2_0),.clk(gclk));
	jdff dff_B_5soQjnSu7_0(.din(w_dff_B_OGYbucAE2_0),.dout(w_dff_B_5soQjnSu7_0),.clk(gclk));
	jdff dff_B_Tfb2awxR8_0(.din(w_dff_B_5soQjnSu7_0),.dout(w_dff_B_Tfb2awxR8_0),.clk(gclk));
	jdff dff_B_QW5uwTx62_0(.din(w_dff_B_Tfb2awxR8_0),.dout(w_dff_B_QW5uwTx62_0),.clk(gclk));
	jdff dff_B_J79DAcIc8_0(.din(w_dff_B_QW5uwTx62_0),.dout(w_dff_B_J79DAcIc8_0),.clk(gclk));
	jdff dff_B_sYWKG7EC6_0(.din(w_dff_B_J79DAcIc8_0),.dout(w_dff_B_sYWKG7EC6_0),.clk(gclk));
	jdff dff_B_VQvPcADU8_0(.din(w_dff_B_sYWKG7EC6_0),.dout(w_dff_B_VQvPcADU8_0),.clk(gclk));
	jdff dff_B_AL82UpN57_0(.din(w_dff_B_VQvPcADU8_0),.dout(w_dff_B_AL82UpN57_0),.clk(gclk));
	jdff dff_B_ZdleOjl17_0(.din(w_dff_B_AL82UpN57_0),.dout(w_dff_B_ZdleOjl17_0),.clk(gclk));
	jdff dff_B_1R7ICl8B5_0(.din(w_dff_B_ZdleOjl17_0),.dout(w_dff_B_1R7ICl8B5_0),.clk(gclk));
	jdff dff_B_6j3JQ2Ye1_0(.din(w_dff_B_1R7ICl8B5_0),.dout(w_dff_B_6j3JQ2Ye1_0),.clk(gclk));
	jdff dff_B_GwRlqcdt9_0(.din(w_dff_B_6j3JQ2Ye1_0),.dout(w_dff_B_GwRlqcdt9_0),.clk(gclk));
	jdff dff_B_aFU78AoU4_0(.din(w_dff_B_GwRlqcdt9_0),.dout(w_dff_B_aFU78AoU4_0),.clk(gclk));
	jdff dff_B_k7Sv53oC8_0(.din(w_dff_B_aFU78AoU4_0),.dout(w_dff_B_k7Sv53oC8_0),.clk(gclk));
	jdff dff_B_zNXCch063_0(.din(w_dff_B_k7Sv53oC8_0),.dout(w_dff_B_zNXCch063_0),.clk(gclk));
	jdff dff_B_06188mbO7_0(.din(w_dff_B_zNXCch063_0),.dout(w_dff_B_06188mbO7_0),.clk(gclk));
	jdff dff_B_0T21YHHZ5_0(.din(w_dff_B_06188mbO7_0),.dout(w_dff_B_0T21YHHZ5_0),.clk(gclk));
	jdff dff_B_4MTCsF4h5_0(.din(w_dff_B_0T21YHHZ5_0),.dout(w_dff_B_4MTCsF4h5_0),.clk(gclk));
	jdff dff_B_Z2ZYBYoe5_0(.din(w_dff_B_4MTCsF4h5_0),.dout(w_dff_B_Z2ZYBYoe5_0),.clk(gclk));
	jdff dff_B_9NJc5g0k8_0(.din(w_dff_B_Z2ZYBYoe5_0),.dout(w_dff_B_9NJc5g0k8_0),.clk(gclk));
	jdff dff_B_tsUyjEzS5_0(.din(w_dff_B_9NJc5g0k8_0),.dout(w_dff_B_tsUyjEzS5_0),.clk(gclk));
	jdff dff_B_dRJvOagH5_0(.din(w_dff_B_tsUyjEzS5_0),.dout(w_dff_B_dRJvOagH5_0),.clk(gclk));
	jdff dff_B_X1ffWE3Q5_0(.din(w_dff_B_dRJvOagH5_0),.dout(w_dff_B_X1ffWE3Q5_0),.clk(gclk));
	jdff dff_B_rTAMs7736_0(.din(w_dff_B_X1ffWE3Q5_0),.dout(w_dff_B_rTAMs7736_0),.clk(gclk));
	jdff dff_B_m05ehC0M4_0(.din(w_dff_B_rTAMs7736_0),.dout(w_dff_B_m05ehC0M4_0),.clk(gclk));
	jdff dff_B_R0ah8XUb0_0(.din(w_dff_B_m05ehC0M4_0),.dout(w_dff_B_R0ah8XUb0_0),.clk(gclk));
	jdff dff_B_R9A4UXxW7_0(.din(w_dff_B_R0ah8XUb0_0),.dout(w_dff_B_R9A4UXxW7_0),.clk(gclk));
	jdff dff_B_EPxWfQPV7_0(.din(w_dff_B_R9A4UXxW7_0),.dout(w_dff_B_EPxWfQPV7_0),.clk(gclk));
	jdff dff_B_Mf4bGIIs7_0(.din(n1108),.dout(w_dff_B_Mf4bGIIs7_0),.clk(gclk));
	jdff dff_B_QaQNlswz9_0(.din(w_dff_B_Mf4bGIIs7_0),.dout(w_dff_B_QaQNlswz9_0),.clk(gclk));
	jdff dff_B_EuzV3vtZ1_0(.din(w_dff_B_QaQNlswz9_0),.dout(w_dff_B_EuzV3vtZ1_0),.clk(gclk));
	jdff dff_B_QNasHvvk5_0(.din(w_dff_B_EuzV3vtZ1_0),.dout(w_dff_B_QNasHvvk5_0),.clk(gclk));
	jdff dff_B_y4hAOaeC8_0(.din(w_dff_B_QNasHvvk5_0),.dout(w_dff_B_y4hAOaeC8_0),.clk(gclk));
	jdff dff_B_DW7Hd0zZ4_0(.din(w_dff_B_y4hAOaeC8_0),.dout(w_dff_B_DW7Hd0zZ4_0),.clk(gclk));
	jdff dff_B_pEIU1tti0_0(.din(w_dff_B_DW7Hd0zZ4_0),.dout(w_dff_B_pEIU1tti0_0),.clk(gclk));
	jdff dff_B_ansSb8I39_0(.din(w_dff_B_pEIU1tti0_0),.dout(w_dff_B_ansSb8I39_0),.clk(gclk));
	jdff dff_B_fAjzcvNj6_0(.din(w_dff_B_ansSb8I39_0),.dout(w_dff_B_fAjzcvNj6_0),.clk(gclk));
	jdff dff_B_QLIZezVG4_0(.din(w_dff_B_fAjzcvNj6_0),.dout(w_dff_B_QLIZezVG4_0),.clk(gclk));
	jdff dff_B_Qg9q82gk7_0(.din(w_dff_B_QLIZezVG4_0),.dout(w_dff_B_Qg9q82gk7_0),.clk(gclk));
	jdff dff_B_dRcAfLlT1_0(.din(w_dff_B_Qg9q82gk7_0),.dout(w_dff_B_dRcAfLlT1_0),.clk(gclk));
	jdff dff_B_03kc00be7_0(.din(w_dff_B_dRcAfLlT1_0),.dout(w_dff_B_03kc00be7_0),.clk(gclk));
	jdff dff_B_tTmkozGb2_0(.din(w_dff_B_03kc00be7_0),.dout(w_dff_B_tTmkozGb2_0),.clk(gclk));
	jdff dff_B_mvqwZPIt5_0(.din(w_dff_B_tTmkozGb2_0),.dout(w_dff_B_mvqwZPIt5_0),.clk(gclk));
	jdff dff_B_fsFWWfRn4_0(.din(w_dff_B_mvqwZPIt5_0),.dout(w_dff_B_fsFWWfRn4_0),.clk(gclk));
	jdff dff_B_ryLtxjvR4_0(.din(w_dff_B_fsFWWfRn4_0),.dout(w_dff_B_ryLtxjvR4_0),.clk(gclk));
	jdff dff_B_Zi7Kn8s95_0(.din(w_dff_B_ryLtxjvR4_0),.dout(w_dff_B_Zi7Kn8s95_0),.clk(gclk));
	jdff dff_B_ewEgondB9_0(.din(w_dff_B_Zi7Kn8s95_0),.dout(w_dff_B_ewEgondB9_0),.clk(gclk));
	jdff dff_B_s8fARmAD6_0(.din(w_dff_B_ewEgondB9_0),.dout(w_dff_B_s8fARmAD6_0),.clk(gclk));
	jdff dff_B_eeDG3VW25_0(.din(w_dff_B_s8fARmAD6_0),.dout(w_dff_B_eeDG3VW25_0),.clk(gclk));
	jdff dff_B_DxlMODMl8_0(.din(w_dff_B_eeDG3VW25_0),.dout(w_dff_B_DxlMODMl8_0),.clk(gclk));
	jdff dff_B_ZaOHtoZ17_0(.din(w_dff_B_DxlMODMl8_0),.dout(w_dff_B_ZaOHtoZ17_0),.clk(gclk));
	jdff dff_B_f7st35aB7_0(.din(w_dff_B_ZaOHtoZ17_0),.dout(w_dff_B_f7st35aB7_0),.clk(gclk));
	jdff dff_B_gX65ix2R6_0(.din(w_dff_B_f7st35aB7_0),.dout(w_dff_B_gX65ix2R6_0),.clk(gclk));
	jdff dff_B_XaPkAPXA9_0(.din(w_dff_B_gX65ix2R6_0),.dout(w_dff_B_XaPkAPXA9_0),.clk(gclk));
	jdff dff_B_YvAd3XN95_0(.din(w_dff_B_XaPkAPXA9_0),.dout(w_dff_B_YvAd3XN95_0),.clk(gclk));
	jdff dff_B_If53B8Lr3_0(.din(w_dff_B_YvAd3XN95_0),.dout(w_dff_B_If53B8Lr3_0),.clk(gclk));
	jdff dff_B_3qhl4UMJ7_0(.din(w_dff_B_If53B8Lr3_0),.dout(w_dff_B_3qhl4UMJ7_0),.clk(gclk));
	jdff dff_B_FjrUDAfU4_0(.din(w_dff_B_3qhl4UMJ7_0),.dout(w_dff_B_FjrUDAfU4_0),.clk(gclk));
	jdff dff_B_99w7Z6TT5_0(.din(w_dff_B_FjrUDAfU4_0),.dout(w_dff_B_99w7Z6TT5_0),.clk(gclk));
	jdff dff_B_gGSxsUmt7_0(.din(w_dff_B_99w7Z6TT5_0),.dout(w_dff_B_gGSxsUmt7_0),.clk(gclk));
	jdff dff_B_oHLn4Y4u5_0(.din(w_dff_B_gGSxsUmt7_0),.dout(w_dff_B_oHLn4Y4u5_0),.clk(gclk));
	jdff dff_B_m1lKuX0E8_0(.din(w_dff_B_oHLn4Y4u5_0),.dout(w_dff_B_m1lKuX0E8_0),.clk(gclk));
	jdff dff_B_FoVXwOim6_0(.din(w_dff_B_m1lKuX0E8_0),.dout(w_dff_B_FoVXwOim6_0),.clk(gclk));
	jdff dff_B_Ci8weqxh9_0(.din(w_dff_B_FoVXwOim6_0),.dout(w_dff_B_Ci8weqxh9_0),.clk(gclk));
	jdff dff_B_dvfqsnxx7_0(.din(w_dff_B_Ci8weqxh9_0),.dout(w_dff_B_dvfqsnxx7_0),.clk(gclk));
	jdff dff_B_uaufbcCs8_0(.din(w_dff_B_dvfqsnxx7_0),.dout(w_dff_B_uaufbcCs8_0),.clk(gclk));
	jdff dff_B_VwnMBN5V0_0(.din(w_dff_B_uaufbcCs8_0),.dout(w_dff_B_VwnMBN5V0_0),.clk(gclk));
	jdff dff_B_PAFSZUxB2_0(.din(w_dff_B_VwnMBN5V0_0),.dout(w_dff_B_PAFSZUxB2_0),.clk(gclk));
	jdff dff_B_fTJkyqac6_0(.din(w_dff_B_PAFSZUxB2_0),.dout(w_dff_B_fTJkyqac6_0),.clk(gclk));
	jdff dff_B_Z5KanTJ08_0(.din(w_dff_B_fTJkyqac6_0),.dout(w_dff_B_Z5KanTJ08_0),.clk(gclk));
	jdff dff_B_sumWS9Vf1_0(.din(w_dff_B_Z5KanTJ08_0),.dout(w_dff_B_sumWS9Vf1_0),.clk(gclk));
	jdff dff_B_Hs5hme0D4_0(.din(w_dff_B_sumWS9Vf1_0),.dout(w_dff_B_Hs5hme0D4_0),.clk(gclk));
	jdff dff_B_aUHOxU028_0(.din(w_dff_B_Hs5hme0D4_0),.dout(w_dff_B_aUHOxU028_0),.clk(gclk));
	jdff dff_B_bDPtbaLa9_0(.din(w_dff_B_aUHOxU028_0),.dout(w_dff_B_bDPtbaLa9_0),.clk(gclk));
	jdff dff_B_LWzBJ1wn8_0(.din(w_dff_B_bDPtbaLa9_0),.dout(w_dff_B_LWzBJ1wn8_0),.clk(gclk));
	jdff dff_B_K9EmdHoN5_0(.din(w_dff_B_LWzBJ1wn8_0),.dout(w_dff_B_K9EmdHoN5_0),.clk(gclk));
	jdff dff_B_VUr17GFe9_0(.din(w_dff_B_K9EmdHoN5_0),.dout(w_dff_B_VUr17GFe9_0),.clk(gclk));
	jdff dff_B_Am7rY1bk0_0(.din(w_dff_B_VUr17GFe9_0),.dout(w_dff_B_Am7rY1bk0_0),.clk(gclk));
	jdff dff_B_U4RWagem4_0(.din(w_dff_B_Am7rY1bk0_0),.dout(w_dff_B_U4RWagem4_0),.clk(gclk));
	jdff dff_B_xMv1cFCZ6_0(.din(w_dff_B_U4RWagem4_0),.dout(w_dff_B_xMv1cFCZ6_0),.clk(gclk));
	jdff dff_B_iJ80qHxz8_0(.din(w_dff_B_xMv1cFCZ6_0),.dout(w_dff_B_iJ80qHxz8_0),.clk(gclk));
	jdff dff_B_ZyQYSZ7M0_0(.din(w_dff_B_iJ80qHxz8_0),.dout(w_dff_B_ZyQYSZ7M0_0),.clk(gclk));
	jdff dff_B_vqi0rSWK0_0(.din(w_dff_B_ZyQYSZ7M0_0),.dout(w_dff_B_vqi0rSWK0_0),.clk(gclk));
	jdff dff_B_JNlauO5R2_0(.din(w_dff_B_vqi0rSWK0_0),.dout(w_dff_B_JNlauO5R2_0),.clk(gclk));
	jdff dff_B_q8wKsiWr7_0(.din(w_dff_B_JNlauO5R2_0),.dout(w_dff_B_q8wKsiWr7_0),.clk(gclk));
	jdff dff_B_BT95v4uZ1_0(.din(w_dff_B_q8wKsiWr7_0),.dout(w_dff_B_BT95v4uZ1_0),.clk(gclk));
	jdff dff_B_zUs7LGxC3_0(.din(w_dff_B_BT95v4uZ1_0),.dout(w_dff_B_zUs7LGxC3_0),.clk(gclk));
	jdff dff_B_dERnxNsj3_0(.din(w_dff_B_zUs7LGxC3_0),.dout(w_dff_B_dERnxNsj3_0),.clk(gclk));
	jdff dff_B_5xRsFM2h0_0(.din(w_dff_B_dERnxNsj3_0),.dout(w_dff_B_5xRsFM2h0_0),.clk(gclk));
	jdff dff_B_SVtCOT2J2_0(.din(w_dff_B_5xRsFM2h0_0),.dout(w_dff_B_SVtCOT2J2_0),.clk(gclk));
	jdff dff_B_HZqNBcJf9_0(.din(w_dff_B_SVtCOT2J2_0),.dout(w_dff_B_HZqNBcJf9_0),.clk(gclk));
	jdff dff_B_Pf0M2pUw5_0(.din(w_dff_B_HZqNBcJf9_0),.dout(w_dff_B_Pf0M2pUw5_0),.clk(gclk));
	jdff dff_B_oft0TmF22_0(.din(w_dff_B_Pf0M2pUw5_0),.dout(w_dff_B_oft0TmF22_0),.clk(gclk));
	jdff dff_B_MeInrIck5_0(.din(w_dff_B_oft0TmF22_0),.dout(w_dff_B_MeInrIck5_0),.clk(gclk));
	jdff dff_B_D7IZ15Xj8_0(.din(w_dff_B_MeInrIck5_0),.dout(w_dff_B_D7IZ15Xj8_0),.clk(gclk));
	jdff dff_B_lex8LvAY0_0(.din(w_dff_B_D7IZ15Xj8_0),.dout(w_dff_B_lex8LvAY0_0),.clk(gclk));
	jdff dff_B_0EacPJrC4_0(.din(w_dff_B_lex8LvAY0_0),.dout(w_dff_B_0EacPJrC4_0),.clk(gclk));
	jdff dff_B_K6gDg8ps6_0(.din(w_dff_B_0EacPJrC4_0),.dout(w_dff_B_K6gDg8ps6_0),.clk(gclk));
	jdff dff_B_R6jgogip4_0(.din(w_dff_B_K6gDg8ps6_0),.dout(w_dff_B_R6jgogip4_0),.clk(gclk));
	jdff dff_B_UxC2HckD4_0(.din(w_dff_B_R6jgogip4_0),.dout(w_dff_B_UxC2HckD4_0),.clk(gclk));
	jdff dff_B_tTc713Uj8_0(.din(w_dff_B_UxC2HckD4_0),.dout(w_dff_B_tTc713Uj8_0),.clk(gclk));
	jdff dff_B_oRHtQbeD3_0(.din(w_dff_B_tTc713Uj8_0),.dout(w_dff_B_oRHtQbeD3_0),.clk(gclk));
	jdff dff_B_9xMQN7mS8_0(.din(w_dff_B_oRHtQbeD3_0),.dout(w_dff_B_9xMQN7mS8_0),.clk(gclk));
	jdff dff_B_ywF9zxmX0_0(.din(w_dff_B_9xMQN7mS8_0),.dout(w_dff_B_ywF9zxmX0_0),.clk(gclk));
	jdff dff_B_b2mL7x6g3_0(.din(w_dff_B_ywF9zxmX0_0),.dout(w_dff_B_b2mL7x6g3_0),.clk(gclk));
	jdff dff_B_QA871eee6_0(.din(w_dff_B_b2mL7x6g3_0),.dout(w_dff_B_QA871eee6_0),.clk(gclk));
	jdff dff_B_pyQmjL5f4_0(.din(w_dff_B_QA871eee6_0),.dout(w_dff_B_pyQmjL5f4_0),.clk(gclk));
	jdff dff_B_Kz5OZ4SS3_0(.din(w_dff_B_pyQmjL5f4_0),.dout(w_dff_B_Kz5OZ4SS3_0),.clk(gclk));
	jdff dff_B_GX8upgfY9_0(.din(w_dff_B_Kz5OZ4SS3_0),.dout(w_dff_B_GX8upgfY9_0),.clk(gclk));
	jdff dff_B_7KiseVrI1_0(.din(w_dff_B_GX8upgfY9_0),.dout(w_dff_B_7KiseVrI1_0),.clk(gclk));
	jdff dff_B_USkwMxb58_0(.din(w_dff_B_7KiseVrI1_0),.dout(w_dff_B_USkwMxb58_0),.clk(gclk));
	jdff dff_B_1PbrWO2m0_0(.din(w_dff_B_USkwMxb58_0),.dout(w_dff_B_1PbrWO2m0_0),.clk(gclk));
	jdff dff_B_YL5KE44k3_0(.din(w_dff_B_1PbrWO2m0_0),.dout(w_dff_B_YL5KE44k3_0),.clk(gclk));
	jdff dff_B_jr9TK7yz0_0(.din(w_dff_B_YL5KE44k3_0),.dout(w_dff_B_jr9TK7yz0_0),.clk(gclk));
	jdff dff_B_YE7lnPud9_0(.din(w_dff_B_jr9TK7yz0_0),.dout(w_dff_B_YE7lnPud9_0),.clk(gclk));
	jdff dff_B_6SYbh95w9_0(.din(w_dff_B_YE7lnPud9_0),.dout(w_dff_B_6SYbh95w9_0),.clk(gclk));
	jdff dff_B_BZZufOtI5_0(.din(w_dff_B_6SYbh95w9_0),.dout(w_dff_B_BZZufOtI5_0),.clk(gclk));
	jdff dff_B_yqvkyrSA5_0(.din(w_dff_B_BZZufOtI5_0),.dout(w_dff_B_yqvkyrSA5_0),.clk(gclk));
	jdff dff_B_SsVTULxg1_0(.din(w_dff_B_yqvkyrSA5_0),.dout(w_dff_B_SsVTULxg1_0),.clk(gclk));
	jdff dff_B_tWhdsU6j2_0(.din(w_dff_B_SsVTULxg1_0),.dout(w_dff_B_tWhdsU6j2_0),.clk(gclk));
	jdff dff_B_ZMiI4tSI8_0(.din(w_dff_B_tWhdsU6j2_0),.dout(w_dff_B_ZMiI4tSI8_0),.clk(gclk));
	jdff dff_B_28DVf9vj6_0(.din(w_dff_B_ZMiI4tSI8_0),.dout(w_dff_B_28DVf9vj6_0),.clk(gclk));
	jdff dff_B_WEwKMJx30_0(.din(w_dff_B_28DVf9vj6_0),.dout(w_dff_B_WEwKMJx30_0),.clk(gclk));
	jdff dff_B_EpwZydaA5_0(.din(w_dff_B_WEwKMJx30_0),.dout(w_dff_B_EpwZydaA5_0),.clk(gclk));
	jdff dff_B_eYXoIjyu2_0(.din(w_dff_B_EpwZydaA5_0),.dout(w_dff_B_eYXoIjyu2_0),.clk(gclk));
	jdff dff_B_jrLI29pl5_0(.din(w_dff_B_eYXoIjyu2_0),.dout(w_dff_B_jrLI29pl5_0),.clk(gclk));
	jdff dff_B_JG8DkIUd7_0(.din(w_dff_B_jrLI29pl5_0),.dout(w_dff_B_JG8DkIUd7_0),.clk(gclk));
	jdff dff_B_OxKsOoDk2_0(.din(w_dff_B_JG8DkIUd7_0),.dout(w_dff_B_OxKsOoDk2_0),.clk(gclk));
	jdff dff_B_gSM54LjO2_0(.din(w_dff_B_OxKsOoDk2_0),.dout(w_dff_B_gSM54LjO2_0),.clk(gclk));
	jdff dff_B_DW3JjsXk5_0(.din(w_dff_B_gSM54LjO2_0),.dout(w_dff_B_DW3JjsXk5_0),.clk(gclk));
	jdff dff_B_bMYepiXd0_0(.din(w_dff_B_DW3JjsXk5_0),.dout(w_dff_B_bMYepiXd0_0),.clk(gclk));
	jdff dff_B_RxDlKpGR1_0(.din(w_dff_B_bMYepiXd0_0),.dout(w_dff_B_RxDlKpGR1_0),.clk(gclk));
	jdff dff_B_jgeBD7LJ0_0(.din(w_dff_B_RxDlKpGR1_0),.dout(w_dff_B_jgeBD7LJ0_0),.clk(gclk));
	jdff dff_B_lSnu0hEj7_0(.din(w_dff_B_jgeBD7LJ0_0),.dout(w_dff_B_lSnu0hEj7_0),.clk(gclk));
	jdff dff_B_voGnUNqX6_0(.din(w_dff_B_lSnu0hEj7_0),.dout(w_dff_B_voGnUNqX6_0),.clk(gclk));
	jdff dff_B_RiP2rXi55_0(.din(w_dff_B_voGnUNqX6_0),.dout(w_dff_B_RiP2rXi55_0),.clk(gclk));
	jdff dff_B_Xj5IwNDZ3_0(.din(w_dff_B_RiP2rXi55_0),.dout(w_dff_B_Xj5IwNDZ3_0),.clk(gclk));
	jdff dff_B_DreSfcaI6_0(.din(w_dff_B_Xj5IwNDZ3_0),.dout(w_dff_B_DreSfcaI6_0),.clk(gclk));
	jdff dff_B_sKqGZVVb5_0(.din(w_dff_B_DreSfcaI6_0),.dout(w_dff_B_sKqGZVVb5_0),.clk(gclk));
	jdff dff_B_c9qoYoWt5_0(.din(w_dff_B_sKqGZVVb5_0),.dout(w_dff_B_c9qoYoWt5_0),.clk(gclk));
	jdff dff_B_45FinX8J8_0(.din(w_dff_B_c9qoYoWt5_0),.dout(w_dff_B_45FinX8J8_0),.clk(gclk));
	jdff dff_B_QXacbdg74_0(.din(w_dff_B_45FinX8J8_0),.dout(w_dff_B_QXacbdg74_0),.clk(gclk));
	jdff dff_B_UhqzJBa99_0(.din(w_dff_B_QXacbdg74_0),.dout(w_dff_B_UhqzJBa99_0),.clk(gclk));
	jdff dff_B_Ize3D40m1_0(.din(w_dff_B_UhqzJBa99_0),.dout(w_dff_B_Ize3D40m1_0),.clk(gclk));
	jdff dff_B_ddhj3QHk2_0(.din(w_dff_B_Ize3D40m1_0),.dout(w_dff_B_ddhj3QHk2_0),.clk(gclk));
	jdff dff_B_8W09mOKq3_0(.din(w_dff_B_ddhj3QHk2_0),.dout(w_dff_B_8W09mOKq3_0),.clk(gclk));
	jdff dff_B_em62HQD64_0(.din(w_dff_B_8W09mOKq3_0),.dout(w_dff_B_em62HQD64_0),.clk(gclk));
	jdff dff_B_qhYwhaxn2_0(.din(w_dff_B_em62HQD64_0),.dout(w_dff_B_qhYwhaxn2_0),.clk(gclk));
	jdff dff_B_MI6HC4ki4_0(.din(n1114),.dout(w_dff_B_MI6HC4ki4_0),.clk(gclk));
	jdff dff_B_hCdq7GtP3_0(.din(w_dff_B_MI6HC4ki4_0),.dout(w_dff_B_hCdq7GtP3_0),.clk(gclk));
	jdff dff_B_XsNGDlmV1_0(.din(w_dff_B_hCdq7GtP3_0),.dout(w_dff_B_XsNGDlmV1_0),.clk(gclk));
	jdff dff_B_yKkBc2z46_0(.din(w_dff_B_XsNGDlmV1_0),.dout(w_dff_B_yKkBc2z46_0),.clk(gclk));
	jdff dff_B_snxZhQFr4_0(.din(w_dff_B_yKkBc2z46_0),.dout(w_dff_B_snxZhQFr4_0),.clk(gclk));
	jdff dff_B_8ObNGCI84_0(.din(w_dff_B_snxZhQFr4_0),.dout(w_dff_B_8ObNGCI84_0),.clk(gclk));
	jdff dff_B_HG9Vk3OM7_0(.din(w_dff_B_8ObNGCI84_0),.dout(w_dff_B_HG9Vk3OM7_0),.clk(gclk));
	jdff dff_B_r0rT2Is62_0(.din(w_dff_B_HG9Vk3OM7_0),.dout(w_dff_B_r0rT2Is62_0),.clk(gclk));
	jdff dff_B_5PrLCwF72_0(.din(w_dff_B_r0rT2Is62_0),.dout(w_dff_B_5PrLCwF72_0),.clk(gclk));
	jdff dff_B_lU5TZhx31_0(.din(w_dff_B_5PrLCwF72_0),.dout(w_dff_B_lU5TZhx31_0),.clk(gclk));
	jdff dff_B_gIvtSsaY3_0(.din(w_dff_B_lU5TZhx31_0),.dout(w_dff_B_gIvtSsaY3_0),.clk(gclk));
	jdff dff_B_Io6IhENr2_0(.din(w_dff_B_gIvtSsaY3_0),.dout(w_dff_B_Io6IhENr2_0),.clk(gclk));
	jdff dff_B_j2B6MhCB5_0(.din(w_dff_B_Io6IhENr2_0),.dout(w_dff_B_j2B6MhCB5_0),.clk(gclk));
	jdff dff_B_1YfhAhGF9_0(.din(w_dff_B_j2B6MhCB5_0),.dout(w_dff_B_1YfhAhGF9_0),.clk(gclk));
	jdff dff_B_VGPns6hT5_0(.din(w_dff_B_1YfhAhGF9_0),.dout(w_dff_B_VGPns6hT5_0),.clk(gclk));
	jdff dff_B_sW6nfMfl4_0(.din(w_dff_B_VGPns6hT5_0),.dout(w_dff_B_sW6nfMfl4_0),.clk(gclk));
	jdff dff_B_dUGc9UGL1_0(.din(w_dff_B_sW6nfMfl4_0),.dout(w_dff_B_dUGc9UGL1_0),.clk(gclk));
	jdff dff_B_ssziijg54_0(.din(w_dff_B_dUGc9UGL1_0),.dout(w_dff_B_ssziijg54_0),.clk(gclk));
	jdff dff_B_qBqDYGex6_0(.din(w_dff_B_ssziijg54_0),.dout(w_dff_B_qBqDYGex6_0),.clk(gclk));
	jdff dff_B_bvcHLzuZ9_0(.din(w_dff_B_qBqDYGex6_0),.dout(w_dff_B_bvcHLzuZ9_0),.clk(gclk));
	jdff dff_B_BdjdFfqJ5_0(.din(w_dff_B_bvcHLzuZ9_0),.dout(w_dff_B_BdjdFfqJ5_0),.clk(gclk));
	jdff dff_B_Lcy99c6n0_0(.din(w_dff_B_BdjdFfqJ5_0),.dout(w_dff_B_Lcy99c6n0_0),.clk(gclk));
	jdff dff_B_8T58l3zu0_0(.din(w_dff_B_Lcy99c6n0_0),.dout(w_dff_B_8T58l3zu0_0),.clk(gclk));
	jdff dff_B_MKoIYWEN1_0(.din(w_dff_B_8T58l3zu0_0),.dout(w_dff_B_MKoIYWEN1_0),.clk(gclk));
	jdff dff_B_sFYOgUgD2_0(.din(w_dff_B_MKoIYWEN1_0),.dout(w_dff_B_sFYOgUgD2_0),.clk(gclk));
	jdff dff_B_iqj7Ez2z2_0(.din(w_dff_B_sFYOgUgD2_0),.dout(w_dff_B_iqj7Ez2z2_0),.clk(gclk));
	jdff dff_B_1VTFtqw26_0(.din(w_dff_B_iqj7Ez2z2_0),.dout(w_dff_B_1VTFtqw26_0),.clk(gclk));
	jdff dff_B_QFCS8o9h9_0(.din(w_dff_B_1VTFtqw26_0),.dout(w_dff_B_QFCS8o9h9_0),.clk(gclk));
	jdff dff_B_qCbSgFBQ9_0(.din(w_dff_B_QFCS8o9h9_0),.dout(w_dff_B_qCbSgFBQ9_0),.clk(gclk));
	jdff dff_B_NCSjtdzZ5_0(.din(w_dff_B_qCbSgFBQ9_0),.dout(w_dff_B_NCSjtdzZ5_0),.clk(gclk));
	jdff dff_B_t0LAegjI5_0(.din(w_dff_B_NCSjtdzZ5_0),.dout(w_dff_B_t0LAegjI5_0),.clk(gclk));
	jdff dff_B_lGbTRTlI6_0(.din(w_dff_B_t0LAegjI5_0),.dout(w_dff_B_lGbTRTlI6_0),.clk(gclk));
	jdff dff_B_2Mau76xd5_0(.din(w_dff_B_lGbTRTlI6_0),.dout(w_dff_B_2Mau76xd5_0),.clk(gclk));
	jdff dff_B_ZYiFP1Iv4_0(.din(w_dff_B_2Mau76xd5_0),.dout(w_dff_B_ZYiFP1Iv4_0),.clk(gclk));
	jdff dff_B_ESvanhO48_0(.din(w_dff_B_ZYiFP1Iv4_0),.dout(w_dff_B_ESvanhO48_0),.clk(gclk));
	jdff dff_B_mStUFvyr1_0(.din(w_dff_B_ESvanhO48_0),.dout(w_dff_B_mStUFvyr1_0),.clk(gclk));
	jdff dff_B_qjSeEygS7_0(.din(w_dff_B_mStUFvyr1_0),.dout(w_dff_B_qjSeEygS7_0),.clk(gclk));
	jdff dff_B_NvsNP2829_0(.din(w_dff_B_qjSeEygS7_0),.dout(w_dff_B_NvsNP2829_0),.clk(gclk));
	jdff dff_B_VDy8bCyP8_0(.din(w_dff_B_NvsNP2829_0),.dout(w_dff_B_VDy8bCyP8_0),.clk(gclk));
	jdff dff_B_o1pTnOrf9_0(.din(w_dff_B_VDy8bCyP8_0),.dout(w_dff_B_o1pTnOrf9_0),.clk(gclk));
	jdff dff_B_AOv7yzLK2_0(.din(w_dff_B_o1pTnOrf9_0),.dout(w_dff_B_AOv7yzLK2_0),.clk(gclk));
	jdff dff_B_UjFyqUbx8_0(.din(w_dff_B_AOv7yzLK2_0),.dout(w_dff_B_UjFyqUbx8_0),.clk(gclk));
	jdff dff_B_dZRukDxF5_0(.din(w_dff_B_UjFyqUbx8_0),.dout(w_dff_B_dZRukDxF5_0),.clk(gclk));
	jdff dff_B_GfOiaw6Q0_0(.din(w_dff_B_dZRukDxF5_0),.dout(w_dff_B_GfOiaw6Q0_0),.clk(gclk));
	jdff dff_B_85W6pltF8_0(.din(w_dff_B_GfOiaw6Q0_0),.dout(w_dff_B_85W6pltF8_0),.clk(gclk));
	jdff dff_B_c6d7m3HU2_0(.din(w_dff_B_85W6pltF8_0),.dout(w_dff_B_c6d7m3HU2_0),.clk(gclk));
	jdff dff_B_uZzhl7WP6_0(.din(w_dff_B_c6d7m3HU2_0),.dout(w_dff_B_uZzhl7WP6_0),.clk(gclk));
	jdff dff_B_NWbI1MMV8_0(.din(w_dff_B_uZzhl7WP6_0),.dout(w_dff_B_NWbI1MMV8_0),.clk(gclk));
	jdff dff_B_UEfEi3w39_0(.din(w_dff_B_NWbI1MMV8_0),.dout(w_dff_B_UEfEi3w39_0),.clk(gclk));
	jdff dff_B_wiPKtVAr4_0(.din(w_dff_B_UEfEi3w39_0),.dout(w_dff_B_wiPKtVAr4_0),.clk(gclk));
	jdff dff_B_DzQbWtaQ8_0(.din(w_dff_B_wiPKtVAr4_0),.dout(w_dff_B_DzQbWtaQ8_0),.clk(gclk));
	jdff dff_B_U0D9RSqn3_0(.din(w_dff_B_DzQbWtaQ8_0),.dout(w_dff_B_U0D9RSqn3_0),.clk(gclk));
	jdff dff_B_5Pb8sBBf1_0(.din(w_dff_B_U0D9RSqn3_0),.dout(w_dff_B_5Pb8sBBf1_0),.clk(gclk));
	jdff dff_B_CovSE80Y8_0(.din(w_dff_B_5Pb8sBBf1_0),.dout(w_dff_B_CovSE80Y8_0),.clk(gclk));
	jdff dff_B_1Zq4LUxj6_0(.din(w_dff_B_CovSE80Y8_0),.dout(w_dff_B_1Zq4LUxj6_0),.clk(gclk));
	jdff dff_B_ISTrKf4C6_0(.din(w_dff_B_1Zq4LUxj6_0),.dout(w_dff_B_ISTrKf4C6_0),.clk(gclk));
	jdff dff_B_JDhcM3W96_0(.din(w_dff_B_ISTrKf4C6_0),.dout(w_dff_B_JDhcM3W96_0),.clk(gclk));
	jdff dff_B_sQoUExAW5_0(.din(w_dff_B_JDhcM3W96_0),.dout(w_dff_B_sQoUExAW5_0),.clk(gclk));
	jdff dff_B_ogw97NAZ1_0(.din(w_dff_B_sQoUExAW5_0),.dout(w_dff_B_ogw97NAZ1_0),.clk(gclk));
	jdff dff_B_VQv6UVHk6_0(.din(w_dff_B_ogw97NAZ1_0),.dout(w_dff_B_VQv6UVHk6_0),.clk(gclk));
	jdff dff_B_QBMXYK116_0(.din(w_dff_B_VQv6UVHk6_0),.dout(w_dff_B_QBMXYK116_0),.clk(gclk));
	jdff dff_B_YHtLDvGi4_0(.din(w_dff_B_QBMXYK116_0),.dout(w_dff_B_YHtLDvGi4_0),.clk(gclk));
	jdff dff_B_DVQi1o885_0(.din(w_dff_B_YHtLDvGi4_0),.dout(w_dff_B_DVQi1o885_0),.clk(gclk));
	jdff dff_B_PP84ZHW99_0(.din(w_dff_B_DVQi1o885_0),.dout(w_dff_B_PP84ZHW99_0),.clk(gclk));
	jdff dff_B_1SGkRLQA4_0(.din(w_dff_B_PP84ZHW99_0),.dout(w_dff_B_1SGkRLQA4_0),.clk(gclk));
	jdff dff_B_qNjiej5C5_0(.din(w_dff_B_1SGkRLQA4_0),.dout(w_dff_B_qNjiej5C5_0),.clk(gclk));
	jdff dff_B_ByIazu2g6_0(.din(w_dff_B_qNjiej5C5_0),.dout(w_dff_B_ByIazu2g6_0),.clk(gclk));
	jdff dff_B_zUO80eUi9_0(.din(w_dff_B_ByIazu2g6_0),.dout(w_dff_B_zUO80eUi9_0),.clk(gclk));
	jdff dff_B_5g0mg10I0_0(.din(w_dff_B_zUO80eUi9_0),.dout(w_dff_B_5g0mg10I0_0),.clk(gclk));
	jdff dff_B_xLNxPQP56_0(.din(w_dff_B_5g0mg10I0_0),.dout(w_dff_B_xLNxPQP56_0),.clk(gclk));
	jdff dff_B_BDrDtfkc8_0(.din(w_dff_B_xLNxPQP56_0),.dout(w_dff_B_BDrDtfkc8_0),.clk(gclk));
	jdff dff_B_ZS5RtR481_0(.din(w_dff_B_BDrDtfkc8_0),.dout(w_dff_B_ZS5RtR481_0),.clk(gclk));
	jdff dff_B_LEyHzAeA3_0(.din(w_dff_B_ZS5RtR481_0),.dout(w_dff_B_LEyHzAeA3_0),.clk(gclk));
	jdff dff_B_zrSZD4I47_0(.din(w_dff_B_LEyHzAeA3_0),.dout(w_dff_B_zrSZD4I47_0),.clk(gclk));
	jdff dff_B_gJ9PIjdI8_0(.din(w_dff_B_zrSZD4I47_0),.dout(w_dff_B_gJ9PIjdI8_0),.clk(gclk));
	jdff dff_B_HOTVZBKz6_0(.din(w_dff_B_gJ9PIjdI8_0),.dout(w_dff_B_HOTVZBKz6_0),.clk(gclk));
	jdff dff_B_ka6z1FoH1_0(.din(w_dff_B_HOTVZBKz6_0),.dout(w_dff_B_ka6z1FoH1_0),.clk(gclk));
	jdff dff_B_8I44RRvp5_0(.din(w_dff_B_ka6z1FoH1_0),.dout(w_dff_B_8I44RRvp5_0),.clk(gclk));
	jdff dff_B_atTc2hgQ9_0(.din(w_dff_B_8I44RRvp5_0),.dout(w_dff_B_atTc2hgQ9_0),.clk(gclk));
	jdff dff_B_joWKk9zU8_0(.din(w_dff_B_atTc2hgQ9_0),.dout(w_dff_B_joWKk9zU8_0),.clk(gclk));
	jdff dff_B_pzth4bdp0_0(.din(w_dff_B_joWKk9zU8_0),.dout(w_dff_B_pzth4bdp0_0),.clk(gclk));
	jdff dff_B_284155wq5_0(.din(w_dff_B_pzth4bdp0_0),.dout(w_dff_B_284155wq5_0),.clk(gclk));
	jdff dff_B_1vZ8lB9m6_0(.din(w_dff_B_284155wq5_0),.dout(w_dff_B_1vZ8lB9m6_0),.clk(gclk));
	jdff dff_B_0X0LIAop1_0(.din(w_dff_B_1vZ8lB9m6_0),.dout(w_dff_B_0X0LIAop1_0),.clk(gclk));
	jdff dff_B_XZ0A7KtN8_0(.din(w_dff_B_0X0LIAop1_0),.dout(w_dff_B_XZ0A7KtN8_0),.clk(gclk));
	jdff dff_B_mnnh0AzY7_0(.din(w_dff_B_XZ0A7KtN8_0),.dout(w_dff_B_mnnh0AzY7_0),.clk(gclk));
	jdff dff_B_MKKp3jhp1_0(.din(w_dff_B_mnnh0AzY7_0),.dout(w_dff_B_MKKp3jhp1_0),.clk(gclk));
	jdff dff_B_RZoLLbOj0_0(.din(w_dff_B_MKKp3jhp1_0),.dout(w_dff_B_RZoLLbOj0_0),.clk(gclk));
	jdff dff_B_ENFkvwC06_0(.din(w_dff_B_RZoLLbOj0_0),.dout(w_dff_B_ENFkvwC06_0),.clk(gclk));
	jdff dff_B_9mEdzbOZ5_0(.din(w_dff_B_ENFkvwC06_0),.dout(w_dff_B_9mEdzbOZ5_0),.clk(gclk));
	jdff dff_B_AgmQJTh00_0(.din(w_dff_B_9mEdzbOZ5_0),.dout(w_dff_B_AgmQJTh00_0),.clk(gclk));
	jdff dff_B_fToZhYKv6_0(.din(w_dff_B_AgmQJTh00_0),.dout(w_dff_B_fToZhYKv6_0),.clk(gclk));
	jdff dff_B_p9ed42J71_0(.din(w_dff_B_fToZhYKv6_0),.dout(w_dff_B_p9ed42J71_0),.clk(gclk));
	jdff dff_B_GoAFN8DH7_0(.din(w_dff_B_p9ed42J71_0),.dout(w_dff_B_GoAFN8DH7_0),.clk(gclk));
	jdff dff_B_jQkod9A81_0(.din(w_dff_B_GoAFN8DH7_0),.dout(w_dff_B_jQkod9A81_0),.clk(gclk));
	jdff dff_B_Hgt3bEnx2_0(.din(w_dff_B_jQkod9A81_0),.dout(w_dff_B_Hgt3bEnx2_0),.clk(gclk));
	jdff dff_B_C7skC0hb3_0(.din(w_dff_B_Hgt3bEnx2_0),.dout(w_dff_B_C7skC0hb3_0),.clk(gclk));
	jdff dff_B_V65TL54Q8_0(.din(w_dff_B_C7skC0hb3_0),.dout(w_dff_B_V65TL54Q8_0),.clk(gclk));
	jdff dff_B_IZRQj2473_0(.din(w_dff_B_V65TL54Q8_0),.dout(w_dff_B_IZRQj2473_0),.clk(gclk));
	jdff dff_B_4eavRGSr6_0(.din(w_dff_B_IZRQj2473_0),.dout(w_dff_B_4eavRGSr6_0),.clk(gclk));
	jdff dff_B_rZoTZyJt8_0(.din(w_dff_B_4eavRGSr6_0),.dout(w_dff_B_rZoTZyJt8_0),.clk(gclk));
	jdff dff_B_3v5VLc1J9_0(.din(w_dff_B_rZoTZyJt8_0),.dout(w_dff_B_3v5VLc1J9_0),.clk(gclk));
	jdff dff_B_REMF3GuW0_0(.din(w_dff_B_3v5VLc1J9_0),.dout(w_dff_B_REMF3GuW0_0),.clk(gclk));
	jdff dff_B_YL8zTHVl5_0(.din(w_dff_B_REMF3GuW0_0),.dout(w_dff_B_YL8zTHVl5_0),.clk(gclk));
	jdff dff_B_9thUzuR96_0(.din(w_dff_B_YL8zTHVl5_0),.dout(w_dff_B_9thUzuR96_0),.clk(gclk));
	jdff dff_B_19GLMtJm4_0(.din(w_dff_B_9thUzuR96_0),.dout(w_dff_B_19GLMtJm4_0),.clk(gclk));
	jdff dff_B_EbqXdmSo3_0(.din(w_dff_B_19GLMtJm4_0),.dout(w_dff_B_EbqXdmSo3_0),.clk(gclk));
	jdff dff_B_6UmJmk6w2_0(.din(w_dff_B_EbqXdmSo3_0),.dout(w_dff_B_6UmJmk6w2_0),.clk(gclk));
	jdff dff_B_PPxofY7O6_0(.din(w_dff_B_6UmJmk6w2_0),.dout(w_dff_B_PPxofY7O6_0),.clk(gclk));
	jdff dff_B_c4gdAp6b7_0(.din(w_dff_B_PPxofY7O6_0),.dout(w_dff_B_c4gdAp6b7_0),.clk(gclk));
	jdff dff_B_vpmjKDyh7_0(.din(w_dff_B_c4gdAp6b7_0),.dout(w_dff_B_vpmjKDyh7_0),.clk(gclk));
	jdff dff_B_j2nwwKNV3_0(.din(w_dff_B_vpmjKDyh7_0),.dout(w_dff_B_j2nwwKNV3_0),.clk(gclk));
	jdff dff_B_rnPYDQLn4_0(.din(w_dff_B_j2nwwKNV3_0),.dout(w_dff_B_rnPYDQLn4_0),.clk(gclk));
	jdff dff_B_tcacvOZJ7_0(.din(w_dff_B_rnPYDQLn4_0),.dout(w_dff_B_tcacvOZJ7_0),.clk(gclk));
	jdff dff_B_w68Wzjw10_0(.din(w_dff_B_tcacvOZJ7_0),.dout(w_dff_B_w68Wzjw10_0),.clk(gclk));
	jdff dff_B_8yU9wllU8_0(.din(w_dff_B_w68Wzjw10_0),.dout(w_dff_B_8yU9wllU8_0),.clk(gclk));
	jdff dff_B_FdVK2dLW7_0(.din(w_dff_B_8yU9wllU8_0),.dout(w_dff_B_FdVK2dLW7_0),.clk(gclk));
	jdff dff_B_QI4Zre4z6_0(.din(w_dff_B_FdVK2dLW7_0),.dout(w_dff_B_QI4Zre4z6_0),.clk(gclk));
	jdff dff_B_0lZtMVcn2_0(.din(w_dff_B_QI4Zre4z6_0),.dout(w_dff_B_0lZtMVcn2_0),.clk(gclk));
	jdff dff_B_uFUJ54ht2_0(.din(w_dff_B_0lZtMVcn2_0),.dout(w_dff_B_uFUJ54ht2_0),.clk(gclk));
	jdff dff_B_sBZNRpfz4_0(.din(w_dff_B_uFUJ54ht2_0),.dout(w_dff_B_sBZNRpfz4_0),.clk(gclk));
	jdff dff_B_2QRWqBTN5_0(.din(n1120),.dout(w_dff_B_2QRWqBTN5_0),.clk(gclk));
	jdff dff_B_smbicmKF2_0(.din(w_dff_B_2QRWqBTN5_0),.dout(w_dff_B_smbicmKF2_0),.clk(gclk));
	jdff dff_B_mdCtVYWR7_0(.din(w_dff_B_smbicmKF2_0),.dout(w_dff_B_mdCtVYWR7_0),.clk(gclk));
	jdff dff_B_HgspKiik1_0(.din(w_dff_B_mdCtVYWR7_0),.dout(w_dff_B_HgspKiik1_0),.clk(gclk));
	jdff dff_B_9Ky0V8JL3_0(.din(w_dff_B_HgspKiik1_0),.dout(w_dff_B_9Ky0V8JL3_0),.clk(gclk));
	jdff dff_B_SeDHYRt34_0(.din(w_dff_B_9Ky0V8JL3_0),.dout(w_dff_B_SeDHYRt34_0),.clk(gclk));
	jdff dff_B_P7kR7Qdy5_0(.din(w_dff_B_SeDHYRt34_0),.dout(w_dff_B_P7kR7Qdy5_0),.clk(gclk));
	jdff dff_B_6G9lhlBa7_0(.din(w_dff_B_P7kR7Qdy5_0),.dout(w_dff_B_6G9lhlBa7_0),.clk(gclk));
	jdff dff_B_pbLhd0ZI9_0(.din(w_dff_B_6G9lhlBa7_0),.dout(w_dff_B_pbLhd0ZI9_0),.clk(gclk));
	jdff dff_B_m8tgTlRz8_0(.din(w_dff_B_pbLhd0ZI9_0),.dout(w_dff_B_m8tgTlRz8_0),.clk(gclk));
	jdff dff_B_BKRcikdw8_0(.din(w_dff_B_m8tgTlRz8_0),.dout(w_dff_B_BKRcikdw8_0),.clk(gclk));
	jdff dff_B_j67ywXjT4_0(.din(w_dff_B_BKRcikdw8_0),.dout(w_dff_B_j67ywXjT4_0),.clk(gclk));
	jdff dff_B_5Ra9CF982_0(.din(w_dff_B_j67ywXjT4_0),.dout(w_dff_B_5Ra9CF982_0),.clk(gclk));
	jdff dff_B_FiLo6R6S7_0(.din(w_dff_B_5Ra9CF982_0),.dout(w_dff_B_FiLo6R6S7_0),.clk(gclk));
	jdff dff_B_5bEhIJ632_0(.din(w_dff_B_FiLo6R6S7_0),.dout(w_dff_B_5bEhIJ632_0),.clk(gclk));
	jdff dff_B_jeXDElwt5_0(.din(w_dff_B_5bEhIJ632_0),.dout(w_dff_B_jeXDElwt5_0),.clk(gclk));
	jdff dff_B_bCG1tQmS9_0(.din(w_dff_B_jeXDElwt5_0),.dout(w_dff_B_bCG1tQmS9_0),.clk(gclk));
	jdff dff_B_IjR9ApJg5_0(.din(w_dff_B_bCG1tQmS9_0),.dout(w_dff_B_IjR9ApJg5_0),.clk(gclk));
	jdff dff_B_7rPX4sM22_0(.din(w_dff_B_IjR9ApJg5_0),.dout(w_dff_B_7rPX4sM22_0),.clk(gclk));
	jdff dff_B_sGrvLns29_0(.din(w_dff_B_7rPX4sM22_0),.dout(w_dff_B_sGrvLns29_0),.clk(gclk));
	jdff dff_B_2OtMJ1Xt4_0(.din(w_dff_B_sGrvLns29_0),.dout(w_dff_B_2OtMJ1Xt4_0),.clk(gclk));
	jdff dff_B_68K6qTvt9_0(.din(w_dff_B_2OtMJ1Xt4_0),.dout(w_dff_B_68K6qTvt9_0),.clk(gclk));
	jdff dff_B_eeev1QQd4_0(.din(w_dff_B_68K6qTvt9_0),.dout(w_dff_B_eeev1QQd4_0),.clk(gclk));
	jdff dff_B_hjcSyLNg5_0(.din(w_dff_B_eeev1QQd4_0),.dout(w_dff_B_hjcSyLNg5_0),.clk(gclk));
	jdff dff_B_6M3CObuF1_0(.din(w_dff_B_hjcSyLNg5_0),.dout(w_dff_B_6M3CObuF1_0),.clk(gclk));
	jdff dff_B_9eMXsrWy4_0(.din(w_dff_B_6M3CObuF1_0),.dout(w_dff_B_9eMXsrWy4_0),.clk(gclk));
	jdff dff_B_Mh3FSkp80_0(.din(w_dff_B_9eMXsrWy4_0),.dout(w_dff_B_Mh3FSkp80_0),.clk(gclk));
	jdff dff_B_yWARzmpv9_0(.din(w_dff_B_Mh3FSkp80_0),.dout(w_dff_B_yWARzmpv9_0),.clk(gclk));
	jdff dff_B_RxGkl3gm1_0(.din(w_dff_B_yWARzmpv9_0),.dout(w_dff_B_RxGkl3gm1_0),.clk(gclk));
	jdff dff_B_qTLKcbfh6_0(.din(w_dff_B_RxGkl3gm1_0),.dout(w_dff_B_qTLKcbfh6_0),.clk(gclk));
	jdff dff_B_6KdzJKNr2_0(.din(w_dff_B_qTLKcbfh6_0),.dout(w_dff_B_6KdzJKNr2_0),.clk(gclk));
	jdff dff_B_Fbuael3j4_0(.din(w_dff_B_6KdzJKNr2_0),.dout(w_dff_B_Fbuael3j4_0),.clk(gclk));
	jdff dff_B_QkoZ85Tr4_0(.din(w_dff_B_Fbuael3j4_0),.dout(w_dff_B_QkoZ85Tr4_0),.clk(gclk));
	jdff dff_B_1VDCeoYA1_0(.din(w_dff_B_QkoZ85Tr4_0),.dout(w_dff_B_1VDCeoYA1_0),.clk(gclk));
	jdff dff_B_TxOxlGYx1_0(.din(w_dff_B_1VDCeoYA1_0),.dout(w_dff_B_TxOxlGYx1_0),.clk(gclk));
	jdff dff_B_g7IHH28r6_0(.din(w_dff_B_TxOxlGYx1_0),.dout(w_dff_B_g7IHH28r6_0),.clk(gclk));
	jdff dff_B_OOLDaeKM9_0(.din(w_dff_B_g7IHH28r6_0),.dout(w_dff_B_OOLDaeKM9_0),.clk(gclk));
	jdff dff_B_U5FsKTUb8_0(.din(w_dff_B_OOLDaeKM9_0),.dout(w_dff_B_U5FsKTUb8_0),.clk(gclk));
	jdff dff_B_bRcugeFv7_0(.din(w_dff_B_U5FsKTUb8_0),.dout(w_dff_B_bRcugeFv7_0),.clk(gclk));
	jdff dff_B_oBKVmUkv2_0(.din(w_dff_B_bRcugeFv7_0),.dout(w_dff_B_oBKVmUkv2_0),.clk(gclk));
	jdff dff_B_1uR9BjNH7_0(.din(w_dff_B_oBKVmUkv2_0),.dout(w_dff_B_1uR9BjNH7_0),.clk(gclk));
	jdff dff_B_3GpbkWYZ1_0(.din(w_dff_B_1uR9BjNH7_0),.dout(w_dff_B_3GpbkWYZ1_0),.clk(gclk));
	jdff dff_B_yKw6r9jY3_0(.din(w_dff_B_3GpbkWYZ1_0),.dout(w_dff_B_yKw6r9jY3_0),.clk(gclk));
	jdff dff_B_hHaX25Fb6_0(.din(w_dff_B_yKw6r9jY3_0),.dout(w_dff_B_hHaX25Fb6_0),.clk(gclk));
	jdff dff_B_qju38gGh4_0(.din(w_dff_B_hHaX25Fb6_0),.dout(w_dff_B_qju38gGh4_0),.clk(gclk));
	jdff dff_B_QE9vSeWv1_0(.din(w_dff_B_qju38gGh4_0),.dout(w_dff_B_QE9vSeWv1_0),.clk(gclk));
	jdff dff_B_jjYXaImP1_0(.din(w_dff_B_QE9vSeWv1_0),.dout(w_dff_B_jjYXaImP1_0),.clk(gclk));
	jdff dff_B_javhpdaP0_0(.din(w_dff_B_jjYXaImP1_0),.dout(w_dff_B_javhpdaP0_0),.clk(gclk));
	jdff dff_B_3cYRPfB37_0(.din(w_dff_B_javhpdaP0_0),.dout(w_dff_B_3cYRPfB37_0),.clk(gclk));
	jdff dff_B_cfrql63o5_0(.din(w_dff_B_3cYRPfB37_0),.dout(w_dff_B_cfrql63o5_0),.clk(gclk));
	jdff dff_B_JybZEV0g6_0(.din(w_dff_B_cfrql63o5_0),.dout(w_dff_B_JybZEV0g6_0),.clk(gclk));
	jdff dff_B_3lg6fRCH6_0(.din(w_dff_B_JybZEV0g6_0),.dout(w_dff_B_3lg6fRCH6_0),.clk(gclk));
	jdff dff_B_fMZ9bkJ64_0(.din(w_dff_B_3lg6fRCH6_0),.dout(w_dff_B_fMZ9bkJ64_0),.clk(gclk));
	jdff dff_B_aMrycb0I8_0(.din(w_dff_B_fMZ9bkJ64_0),.dout(w_dff_B_aMrycb0I8_0),.clk(gclk));
	jdff dff_B_ErX8eh0w8_0(.din(w_dff_B_aMrycb0I8_0),.dout(w_dff_B_ErX8eh0w8_0),.clk(gclk));
	jdff dff_B_fz9SrC2q4_0(.din(w_dff_B_ErX8eh0w8_0),.dout(w_dff_B_fz9SrC2q4_0),.clk(gclk));
	jdff dff_B_UOrXbJRB7_0(.din(w_dff_B_fz9SrC2q4_0),.dout(w_dff_B_UOrXbJRB7_0),.clk(gclk));
	jdff dff_B_FdPiqGdg7_0(.din(w_dff_B_UOrXbJRB7_0),.dout(w_dff_B_FdPiqGdg7_0),.clk(gclk));
	jdff dff_B_8Sw8H5AL9_0(.din(w_dff_B_FdPiqGdg7_0),.dout(w_dff_B_8Sw8H5AL9_0),.clk(gclk));
	jdff dff_B_Kk8YkuMB3_0(.din(w_dff_B_8Sw8H5AL9_0),.dout(w_dff_B_Kk8YkuMB3_0),.clk(gclk));
	jdff dff_B_v4AOX7le2_0(.din(w_dff_B_Kk8YkuMB3_0),.dout(w_dff_B_v4AOX7le2_0),.clk(gclk));
	jdff dff_B_1OpR2KMz8_0(.din(w_dff_B_v4AOX7le2_0),.dout(w_dff_B_1OpR2KMz8_0),.clk(gclk));
	jdff dff_B_b9FCcMva1_0(.din(w_dff_B_1OpR2KMz8_0),.dout(w_dff_B_b9FCcMva1_0),.clk(gclk));
	jdff dff_B_TkMiZdKv2_0(.din(w_dff_B_b9FCcMva1_0),.dout(w_dff_B_TkMiZdKv2_0),.clk(gclk));
	jdff dff_B_yXx7r8rJ8_0(.din(w_dff_B_TkMiZdKv2_0),.dout(w_dff_B_yXx7r8rJ8_0),.clk(gclk));
	jdff dff_B_HDJXbPwf3_0(.din(w_dff_B_yXx7r8rJ8_0),.dout(w_dff_B_HDJXbPwf3_0),.clk(gclk));
	jdff dff_B_NfgRmekj8_0(.din(w_dff_B_HDJXbPwf3_0),.dout(w_dff_B_NfgRmekj8_0),.clk(gclk));
	jdff dff_B_8szD1fQj3_0(.din(w_dff_B_NfgRmekj8_0),.dout(w_dff_B_8szD1fQj3_0),.clk(gclk));
	jdff dff_B_XTu2tx6K5_0(.din(w_dff_B_8szD1fQj3_0),.dout(w_dff_B_XTu2tx6K5_0),.clk(gclk));
	jdff dff_B_1Cp3Xlu70_0(.din(w_dff_B_XTu2tx6K5_0),.dout(w_dff_B_1Cp3Xlu70_0),.clk(gclk));
	jdff dff_B_4i5xBvOj4_0(.din(w_dff_B_1Cp3Xlu70_0),.dout(w_dff_B_4i5xBvOj4_0),.clk(gclk));
	jdff dff_B_sFCzxq8x1_0(.din(w_dff_B_4i5xBvOj4_0),.dout(w_dff_B_sFCzxq8x1_0),.clk(gclk));
	jdff dff_B_phmHkO1L6_0(.din(w_dff_B_sFCzxq8x1_0),.dout(w_dff_B_phmHkO1L6_0),.clk(gclk));
	jdff dff_B_pUjW3O9p8_0(.din(w_dff_B_phmHkO1L6_0),.dout(w_dff_B_pUjW3O9p8_0),.clk(gclk));
	jdff dff_B_anFKiTtd6_0(.din(w_dff_B_pUjW3O9p8_0),.dout(w_dff_B_anFKiTtd6_0),.clk(gclk));
	jdff dff_B_H6faowjM1_0(.din(w_dff_B_anFKiTtd6_0),.dout(w_dff_B_H6faowjM1_0),.clk(gclk));
	jdff dff_B_UMLMKIGX4_0(.din(w_dff_B_H6faowjM1_0),.dout(w_dff_B_UMLMKIGX4_0),.clk(gclk));
	jdff dff_B_3nIU2xaG7_0(.din(w_dff_B_UMLMKIGX4_0),.dout(w_dff_B_3nIU2xaG7_0),.clk(gclk));
	jdff dff_B_WuVoAzyj4_0(.din(w_dff_B_3nIU2xaG7_0),.dout(w_dff_B_WuVoAzyj4_0),.clk(gclk));
	jdff dff_B_B6fpBHaI4_0(.din(w_dff_B_WuVoAzyj4_0),.dout(w_dff_B_B6fpBHaI4_0),.clk(gclk));
	jdff dff_B_PCtYaWD78_0(.din(w_dff_B_B6fpBHaI4_0),.dout(w_dff_B_PCtYaWD78_0),.clk(gclk));
	jdff dff_B_4nyGGiF76_0(.din(w_dff_B_PCtYaWD78_0),.dout(w_dff_B_4nyGGiF76_0),.clk(gclk));
	jdff dff_B_v7S6j6CY4_0(.din(w_dff_B_4nyGGiF76_0),.dout(w_dff_B_v7S6j6CY4_0),.clk(gclk));
	jdff dff_B_9Q9O6KN22_0(.din(w_dff_B_v7S6j6CY4_0),.dout(w_dff_B_9Q9O6KN22_0),.clk(gclk));
	jdff dff_B_Ha3Ou0wu8_0(.din(w_dff_B_9Q9O6KN22_0),.dout(w_dff_B_Ha3Ou0wu8_0),.clk(gclk));
	jdff dff_B_1qy6kROB1_0(.din(w_dff_B_Ha3Ou0wu8_0),.dout(w_dff_B_1qy6kROB1_0),.clk(gclk));
	jdff dff_B_kEvV7k6J1_0(.din(w_dff_B_1qy6kROB1_0),.dout(w_dff_B_kEvV7k6J1_0),.clk(gclk));
	jdff dff_B_BziCGQdg9_0(.din(w_dff_B_kEvV7k6J1_0),.dout(w_dff_B_BziCGQdg9_0),.clk(gclk));
	jdff dff_B_0mJkoMhS3_0(.din(w_dff_B_BziCGQdg9_0),.dout(w_dff_B_0mJkoMhS3_0),.clk(gclk));
	jdff dff_B_IMvfyqJ12_0(.din(w_dff_B_0mJkoMhS3_0),.dout(w_dff_B_IMvfyqJ12_0),.clk(gclk));
	jdff dff_B_1yjF3upI3_0(.din(w_dff_B_IMvfyqJ12_0),.dout(w_dff_B_1yjF3upI3_0),.clk(gclk));
	jdff dff_B_hU2xvfoD7_0(.din(w_dff_B_1yjF3upI3_0),.dout(w_dff_B_hU2xvfoD7_0),.clk(gclk));
	jdff dff_B_jH1vbdlj8_0(.din(w_dff_B_hU2xvfoD7_0),.dout(w_dff_B_jH1vbdlj8_0),.clk(gclk));
	jdff dff_B_Q4Iyc5pC2_0(.din(w_dff_B_jH1vbdlj8_0),.dout(w_dff_B_Q4Iyc5pC2_0),.clk(gclk));
	jdff dff_B_GZusmrKV4_0(.din(w_dff_B_Q4Iyc5pC2_0),.dout(w_dff_B_GZusmrKV4_0),.clk(gclk));
	jdff dff_B_kdLNS5yS3_0(.din(w_dff_B_GZusmrKV4_0),.dout(w_dff_B_kdLNS5yS3_0),.clk(gclk));
	jdff dff_B_WHZpE7LF3_0(.din(w_dff_B_kdLNS5yS3_0),.dout(w_dff_B_WHZpE7LF3_0),.clk(gclk));
	jdff dff_B_3JNz2vpY1_0(.din(w_dff_B_WHZpE7LF3_0),.dout(w_dff_B_3JNz2vpY1_0),.clk(gclk));
	jdff dff_B_Gblky7394_0(.din(w_dff_B_3JNz2vpY1_0),.dout(w_dff_B_Gblky7394_0),.clk(gclk));
	jdff dff_B_yf4HX0u41_0(.din(w_dff_B_Gblky7394_0),.dout(w_dff_B_yf4HX0u41_0),.clk(gclk));
	jdff dff_B_nvu97efN1_0(.din(w_dff_B_yf4HX0u41_0),.dout(w_dff_B_nvu97efN1_0),.clk(gclk));
	jdff dff_B_qwVr1rC41_0(.din(w_dff_B_nvu97efN1_0),.dout(w_dff_B_qwVr1rC41_0),.clk(gclk));
	jdff dff_B_2w3gAkD51_0(.din(w_dff_B_qwVr1rC41_0),.dout(w_dff_B_2w3gAkD51_0),.clk(gclk));
	jdff dff_B_GhXrqSip5_0(.din(w_dff_B_2w3gAkD51_0),.dout(w_dff_B_GhXrqSip5_0),.clk(gclk));
	jdff dff_B_Zt6Razf06_0(.din(w_dff_B_GhXrqSip5_0),.dout(w_dff_B_Zt6Razf06_0),.clk(gclk));
	jdff dff_B_sOUg29rq1_0(.din(w_dff_B_Zt6Razf06_0),.dout(w_dff_B_sOUg29rq1_0),.clk(gclk));
	jdff dff_B_iIcRMXxs5_0(.din(w_dff_B_sOUg29rq1_0),.dout(w_dff_B_iIcRMXxs5_0),.clk(gclk));
	jdff dff_B_BUHZyAWR0_0(.din(w_dff_B_iIcRMXxs5_0),.dout(w_dff_B_BUHZyAWR0_0),.clk(gclk));
	jdff dff_B_FLyeW2pl1_0(.din(w_dff_B_BUHZyAWR0_0),.dout(w_dff_B_FLyeW2pl1_0),.clk(gclk));
	jdff dff_B_wWRlteQQ2_0(.din(w_dff_B_FLyeW2pl1_0),.dout(w_dff_B_wWRlteQQ2_0),.clk(gclk));
	jdff dff_B_PTeZlwlE6_0(.din(w_dff_B_wWRlteQQ2_0),.dout(w_dff_B_PTeZlwlE6_0),.clk(gclk));
	jdff dff_B_lHTRrGFV1_0(.din(w_dff_B_PTeZlwlE6_0),.dout(w_dff_B_lHTRrGFV1_0),.clk(gclk));
	jdff dff_B_ecVL8fmo2_0(.din(w_dff_B_lHTRrGFV1_0),.dout(w_dff_B_ecVL8fmo2_0),.clk(gclk));
	jdff dff_B_jVlAcpZ07_0(.din(w_dff_B_ecVL8fmo2_0),.dout(w_dff_B_jVlAcpZ07_0),.clk(gclk));
	jdff dff_B_KhIlBopL1_0(.din(w_dff_B_jVlAcpZ07_0),.dout(w_dff_B_KhIlBopL1_0),.clk(gclk));
	jdff dff_B_eyergLvU9_0(.din(w_dff_B_KhIlBopL1_0),.dout(w_dff_B_eyergLvU9_0),.clk(gclk));
	jdff dff_B_5meeMWcj3_0(.din(w_dff_B_eyergLvU9_0),.dout(w_dff_B_5meeMWcj3_0),.clk(gclk));
	jdff dff_B_Xh6h7Du88_0(.din(w_dff_B_5meeMWcj3_0),.dout(w_dff_B_Xh6h7Du88_0),.clk(gclk));
	jdff dff_B_bcVvLfRG8_0(.din(w_dff_B_Xh6h7Du88_0),.dout(w_dff_B_bcVvLfRG8_0),.clk(gclk));
	jdff dff_B_FSoIWlHL6_0(.din(w_dff_B_bcVvLfRG8_0),.dout(w_dff_B_FSoIWlHL6_0),.clk(gclk));
	jdff dff_B_xEbicrAq0_0(.din(w_dff_B_FSoIWlHL6_0),.dout(w_dff_B_xEbicrAq0_0),.clk(gclk));
	jdff dff_B_A7qvzuar1_0(.din(w_dff_B_xEbicrAq0_0),.dout(w_dff_B_A7qvzuar1_0),.clk(gclk));
	jdff dff_B_aPcMadu43_0(.din(n1126),.dout(w_dff_B_aPcMadu43_0),.clk(gclk));
	jdff dff_B_Oy2qUmD86_0(.din(w_dff_B_aPcMadu43_0),.dout(w_dff_B_Oy2qUmD86_0),.clk(gclk));
	jdff dff_B_DtXJgLC54_0(.din(w_dff_B_Oy2qUmD86_0),.dout(w_dff_B_DtXJgLC54_0),.clk(gclk));
	jdff dff_B_3WtYBPXV5_0(.din(w_dff_B_DtXJgLC54_0),.dout(w_dff_B_3WtYBPXV5_0),.clk(gclk));
	jdff dff_B_4eYAOaTo8_0(.din(w_dff_B_3WtYBPXV5_0),.dout(w_dff_B_4eYAOaTo8_0),.clk(gclk));
	jdff dff_B_T0S1fxii1_0(.din(w_dff_B_4eYAOaTo8_0),.dout(w_dff_B_T0S1fxii1_0),.clk(gclk));
	jdff dff_B_b1Ymardl7_0(.din(w_dff_B_T0S1fxii1_0),.dout(w_dff_B_b1Ymardl7_0),.clk(gclk));
	jdff dff_B_pqJMNoT86_0(.din(w_dff_B_b1Ymardl7_0),.dout(w_dff_B_pqJMNoT86_0),.clk(gclk));
	jdff dff_B_NfLNTYs39_0(.din(w_dff_B_pqJMNoT86_0),.dout(w_dff_B_NfLNTYs39_0),.clk(gclk));
	jdff dff_B_KyDhcp9D5_0(.din(w_dff_B_NfLNTYs39_0),.dout(w_dff_B_KyDhcp9D5_0),.clk(gclk));
	jdff dff_B_LCasklDP8_0(.din(w_dff_B_KyDhcp9D5_0),.dout(w_dff_B_LCasklDP8_0),.clk(gclk));
	jdff dff_B_MMDUX33q7_0(.din(w_dff_B_LCasklDP8_0),.dout(w_dff_B_MMDUX33q7_0),.clk(gclk));
	jdff dff_B_An18KtIF3_0(.din(w_dff_B_MMDUX33q7_0),.dout(w_dff_B_An18KtIF3_0),.clk(gclk));
	jdff dff_B_RAJSq0ts6_0(.din(w_dff_B_An18KtIF3_0),.dout(w_dff_B_RAJSq0ts6_0),.clk(gclk));
	jdff dff_B_HuWpDLE56_0(.din(w_dff_B_RAJSq0ts6_0),.dout(w_dff_B_HuWpDLE56_0),.clk(gclk));
	jdff dff_B_NhwbHhev1_0(.din(w_dff_B_HuWpDLE56_0),.dout(w_dff_B_NhwbHhev1_0),.clk(gclk));
	jdff dff_B_YRI7OsJv7_0(.din(w_dff_B_NhwbHhev1_0),.dout(w_dff_B_YRI7OsJv7_0),.clk(gclk));
	jdff dff_B_IL0XQ2Gf9_0(.din(w_dff_B_YRI7OsJv7_0),.dout(w_dff_B_IL0XQ2Gf9_0),.clk(gclk));
	jdff dff_B_ZSWQYgik1_0(.din(w_dff_B_IL0XQ2Gf9_0),.dout(w_dff_B_ZSWQYgik1_0),.clk(gclk));
	jdff dff_B_3UeKj0wI6_0(.din(w_dff_B_ZSWQYgik1_0),.dout(w_dff_B_3UeKj0wI6_0),.clk(gclk));
	jdff dff_B_td0aycKm9_0(.din(w_dff_B_3UeKj0wI6_0),.dout(w_dff_B_td0aycKm9_0),.clk(gclk));
	jdff dff_B_RtpiBDq05_0(.din(w_dff_B_td0aycKm9_0),.dout(w_dff_B_RtpiBDq05_0),.clk(gclk));
	jdff dff_B_7OGDhqiW4_0(.din(w_dff_B_RtpiBDq05_0),.dout(w_dff_B_7OGDhqiW4_0),.clk(gclk));
	jdff dff_B_eBH4Nj4a2_0(.din(w_dff_B_7OGDhqiW4_0),.dout(w_dff_B_eBH4Nj4a2_0),.clk(gclk));
	jdff dff_B_bXyXzKVd9_0(.din(w_dff_B_eBH4Nj4a2_0),.dout(w_dff_B_bXyXzKVd9_0),.clk(gclk));
	jdff dff_B_QDR0W5Gu0_0(.din(w_dff_B_bXyXzKVd9_0),.dout(w_dff_B_QDR0W5Gu0_0),.clk(gclk));
	jdff dff_B_6u9PMJ075_0(.din(w_dff_B_QDR0W5Gu0_0),.dout(w_dff_B_6u9PMJ075_0),.clk(gclk));
	jdff dff_B_s74rdd5T0_0(.din(w_dff_B_6u9PMJ075_0),.dout(w_dff_B_s74rdd5T0_0),.clk(gclk));
	jdff dff_B_rLBFfNfn7_0(.din(w_dff_B_s74rdd5T0_0),.dout(w_dff_B_rLBFfNfn7_0),.clk(gclk));
	jdff dff_B_ES4MEgR89_0(.din(w_dff_B_rLBFfNfn7_0),.dout(w_dff_B_ES4MEgR89_0),.clk(gclk));
	jdff dff_B_T2zANDhP2_0(.din(w_dff_B_ES4MEgR89_0),.dout(w_dff_B_T2zANDhP2_0),.clk(gclk));
	jdff dff_B_2jSCno820_0(.din(w_dff_B_T2zANDhP2_0),.dout(w_dff_B_2jSCno820_0),.clk(gclk));
	jdff dff_B_vqvVnJq35_0(.din(w_dff_B_2jSCno820_0),.dout(w_dff_B_vqvVnJq35_0),.clk(gclk));
	jdff dff_B_jIGXsslq5_0(.din(w_dff_B_vqvVnJq35_0),.dout(w_dff_B_jIGXsslq5_0),.clk(gclk));
	jdff dff_B_KiDbaGfZ6_0(.din(w_dff_B_jIGXsslq5_0),.dout(w_dff_B_KiDbaGfZ6_0),.clk(gclk));
	jdff dff_B_fpRKzTs10_0(.din(w_dff_B_KiDbaGfZ6_0),.dout(w_dff_B_fpRKzTs10_0),.clk(gclk));
	jdff dff_B_sIING38w8_0(.din(w_dff_B_fpRKzTs10_0),.dout(w_dff_B_sIING38w8_0),.clk(gclk));
	jdff dff_B_ZsY46qQz4_0(.din(w_dff_B_sIING38w8_0),.dout(w_dff_B_ZsY46qQz4_0),.clk(gclk));
	jdff dff_B_ErAW2XY51_0(.din(w_dff_B_ZsY46qQz4_0),.dout(w_dff_B_ErAW2XY51_0),.clk(gclk));
	jdff dff_B_gEFk0bmc1_0(.din(w_dff_B_ErAW2XY51_0),.dout(w_dff_B_gEFk0bmc1_0),.clk(gclk));
	jdff dff_B_3xKuW1hJ6_0(.din(w_dff_B_gEFk0bmc1_0),.dout(w_dff_B_3xKuW1hJ6_0),.clk(gclk));
	jdff dff_B_HhkzoLIB2_0(.din(w_dff_B_3xKuW1hJ6_0),.dout(w_dff_B_HhkzoLIB2_0),.clk(gclk));
	jdff dff_B_MuZniDyC9_0(.din(w_dff_B_HhkzoLIB2_0),.dout(w_dff_B_MuZniDyC9_0),.clk(gclk));
	jdff dff_B_KuwhWxoR5_0(.din(w_dff_B_MuZniDyC9_0),.dout(w_dff_B_KuwhWxoR5_0),.clk(gclk));
	jdff dff_B_fhhbusxU7_0(.din(w_dff_B_KuwhWxoR5_0),.dout(w_dff_B_fhhbusxU7_0),.clk(gclk));
	jdff dff_B_hDHP5zhU4_0(.din(w_dff_B_fhhbusxU7_0),.dout(w_dff_B_hDHP5zhU4_0),.clk(gclk));
	jdff dff_B_nzYEIVwr7_0(.din(w_dff_B_hDHP5zhU4_0),.dout(w_dff_B_nzYEIVwr7_0),.clk(gclk));
	jdff dff_B_46uvAGbh6_0(.din(w_dff_B_nzYEIVwr7_0),.dout(w_dff_B_46uvAGbh6_0),.clk(gclk));
	jdff dff_B_AHKtGtyA9_0(.din(w_dff_B_46uvAGbh6_0),.dout(w_dff_B_AHKtGtyA9_0),.clk(gclk));
	jdff dff_B_2ghRHon87_0(.din(w_dff_B_AHKtGtyA9_0),.dout(w_dff_B_2ghRHon87_0),.clk(gclk));
	jdff dff_B_bhSZisTk0_0(.din(w_dff_B_2ghRHon87_0),.dout(w_dff_B_bhSZisTk0_0),.clk(gclk));
	jdff dff_B_p3naK36l8_0(.din(w_dff_B_bhSZisTk0_0),.dout(w_dff_B_p3naK36l8_0),.clk(gclk));
	jdff dff_B_FVbAlllk6_0(.din(w_dff_B_p3naK36l8_0),.dout(w_dff_B_FVbAlllk6_0),.clk(gclk));
	jdff dff_B_Dn0jecqQ2_0(.din(w_dff_B_FVbAlllk6_0),.dout(w_dff_B_Dn0jecqQ2_0),.clk(gclk));
	jdff dff_B_ohuDVRCW4_0(.din(w_dff_B_Dn0jecqQ2_0),.dout(w_dff_B_ohuDVRCW4_0),.clk(gclk));
	jdff dff_B_2IA0E61U7_0(.din(w_dff_B_ohuDVRCW4_0),.dout(w_dff_B_2IA0E61U7_0),.clk(gclk));
	jdff dff_B_Up3ANdop7_0(.din(w_dff_B_2IA0E61U7_0),.dout(w_dff_B_Up3ANdop7_0),.clk(gclk));
	jdff dff_B_yeLqkkRE2_0(.din(w_dff_B_Up3ANdop7_0),.dout(w_dff_B_yeLqkkRE2_0),.clk(gclk));
	jdff dff_B_SVmc92bt7_0(.din(w_dff_B_yeLqkkRE2_0),.dout(w_dff_B_SVmc92bt7_0),.clk(gclk));
	jdff dff_B_WJJ7y8Tu3_0(.din(w_dff_B_SVmc92bt7_0),.dout(w_dff_B_WJJ7y8Tu3_0),.clk(gclk));
	jdff dff_B_C0Lb6Ahd1_0(.din(w_dff_B_WJJ7y8Tu3_0),.dout(w_dff_B_C0Lb6Ahd1_0),.clk(gclk));
	jdff dff_B_YuupTCKx4_0(.din(w_dff_B_C0Lb6Ahd1_0),.dout(w_dff_B_YuupTCKx4_0),.clk(gclk));
	jdff dff_B_uDFyPzGp7_0(.din(w_dff_B_YuupTCKx4_0),.dout(w_dff_B_uDFyPzGp7_0),.clk(gclk));
	jdff dff_B_ZhgGiEm79_0(.din(w_dff_B_uDFyPzGp7_0),.dout(w_dff_B_ZhgGiEm79_0),.clk(gclk));
	jdff dff_B_3WmfKVE20_0(.din(w_dff_B_ZhgGiEm79_0),.dout(w_dff_B_3WmfKVE20_0),.clk(gclk));
	jdff dff_B_kz2WX4gh7_0(.din(w_dff_B_3WmfKVE20_0),.dout(w_dff_B_kz2WX4gh7_0),.clk(gclk));
	jdff dff_B_n6Brr1eb3_0(.din(w_dff_B_kz2WX4gh7_0),.dout(w_dff_B_n6Brr1eb3_0),.clk(gclk));
	jdff dff_B_m9yS7dMG9_0(.din(w_dff_B_n6Brr1eb3_0),.dout(w_dff_B_m9yS7dMG9_0),.clk(gclk));
	jdff dff_B_LkM9bzTO1_0(.din(w_dff_B_m9yS7dMG9_0),.dout(w_dff_B_LkM9bzTO1_0),.clk(gclk));
	jdff dff_B_XA6Jgvc14_0(.din(w_dff_B_LkM9bzTO1_0),.dout(w_dff_B_XA6Jgvc14_0),.clk(gclk));
	jdff dff_B_ZvEhLFv78_0(.din(w_dff_B_XA6Jgvc14_0),.dout(w_dff_B_ZvEhLFv78_0),.clk(gclk));
	jdff dff_B_45o3fjhQ8_0(.din(w_dff_B_ZvEhLFv78_0),.dout(w_dff_B_45o3fjhQ8_0),.clk(gclk));
	jdff dff_B_EATydhzE5_0(.din(w_dff_B_45o3fjhQ8_0),.dout(w_dff_B_EATydhzE5_0),.clk(gclk));
	jdff dff_B_gVXHyWQB0_0(.din(w_dff_B_EATydhzE5_0),.dout(w_dff_B_gVXHyWQB0_0),.clk(gclk));
	jdff dff_B_DmkAllKZ6_0(.din(w_dff_B_gVXHyWQB0_0),.dout(w_dff_B_DmkAllKZ6_0),.clk(gclk));
	jdff dff_B_jn1ccoQw8_0(.din(w_dff_B_DmkAllKZ6_0),.dout(w_dff_B_jn1ccoQw8_0),.clk(gclk));
	jdff dff_B_G7wQ0CCE4_0(.din(w_dff_B_jn1ccoQw8_0),.dout(w_dff_B_G7wQ0CCE4_0),.clk(gclk));
	jdff dff_B_HlSrfZPG6_0(.din(w_dff_B_G7wQ0CCE4_0),.dout(w_dff_B_HlSrfZPG6_0),.clk(gclk));
	jdff dff_B_3yoVrpNn1_0(.din(w_dff_B_HlSrfZPG6_0),.dout(w_dff_B_3yoVrpNn1_0),.clk(gclk));
	jdff dff_B_6VPqM88X8_0(.din(w_dff_B_3yoVrpNn1_0),.dout(w_dff_B_6VPqM88X8_0),.clk(gclk));
	jdff dff_B_ZmveveaH3_0(.din(w_dff_B_6VPqM88X8_0),.dout(w_dff_B_ZmveveaH3_0),.clk(gclk));
	jdff dff_B_FUMUhn2t4_0(.din(w_dff_B_ZmveveaH3_0),.dout(w_dff_B_FUMUhn2t4_0),.clk(gclk));
	jdff dff_B_DRGqoQst1_0(.din(w_dff_B_FUMUhn2t4_0),.dout(w_dff_B_DRGqoQst1_0),.clk(gclk));
	jdff dff_B_t56nAR5Z5_0(.din(w_dff_B_DRGqoQst1_0),.dout(w_dff_B_t56nAR5Z5_0),.clk(gclk));
	jdff dff_B_bvUpw8fz1_0(.din(w_dff_B_t56nAR5Z5_0),.dout(w_dff_B_bvUpw8fz1_0),.clk(gclk));
	jdff dff_B_AGsYW8xa2_0(.din(w_dff_B_bvUpw8fz1_0),.dout(w_dff_B_AGsYW8xa2_0),.clk(gclk));
	jdff dff_B_rtt6Mkn48_0(.din(w_dff_B_AGsYW8xa2_0),.dout(w_dff_B_rtt6Mkn48_0),.clk(gclk));
	jdff dff_B_HLpB3qmL5_0(.din(w_dff_B_rtt6Mkn48_0),.dout(w_dff_B_HLpB3qmL5_0),.clk(gclk));
	jdff dff_B_9YJnsIyF7_0(.din(w_dff_B_HLpB3qmL5_0),.dout(w_dff_B_9YJnsIyF7_0),.clk(gclk));
	jdff dff_B_baHvFq3V2_0(.din(w_dff_B_9YJnsIyF7_0),.dout(w_dff_B_baHvFq3V2_0),.clk(gclk));
	jdff dff_B_XFUunqJn0_0(.din(w_dff_B_baHvFq3V2_0),.dout(w_dff_B_XFUunqJn0_0),.clk(gclk));
	jdff dff_B_nlEza59P2_0(.din(w_dff_B_XFUunqJn0_0),.dout(w_dff_B_nlEza59P2_0),.clk(gclk));
	jdff dff_B_5iTdFiWG2_0(.din(w_dff_B_nlEza59P2_0),.dout(w_dff_B_5iTdFiWG2_0),.clk(gclk));
	jdff dff_B_5ik7dOD48_0(.din(w_dff_B_5iTdFiWG2_0),.dout(w_dff_B_5ik7dOD48_0),.clk(gclk));
	jdff dff_B_PaVAueOx8_0(.din(w_dff_B_5ik7dOD48_0),.dout(w_dff_B_PaVAueOx8_0),.clk(gclk));
	jdff dff_B_Y4t0NgXz6_0(.din(w_dff_B_PaVAueOx8_0),.dout(w_dff_B_Y4t0NgXz6_0),.clk(gclk));
	jdff dff_B_qsS8u5Pp1_0(.din(w_dff_B_Y4t0NgXz6_0),.dout(w_dff_B_qsS8u5Pp1_0),.clk(gclk));
	jdff dff_B_BRhErMvA7_0(.din(w_dff_B_qsS8u5Pp1_0),.dout(w_dff_B_BRhErMvA7_0),.clk(gclk));
	jdff dff_B_pHw6SCC42_0(.din(w_dff_B_BRhErMvA7_0),.dout(w_dff_B_pHw6SCC42_0),.clk(gclk));
	jdff dff_B_14qw1mBa3_0(.din(w_dff_B_pHw6SCC42_0),.dout(w_dff_B_14qw1mBa3_0),.clk(gclk));
	jdff dff_B_TE2W0Imk6_0(.din(w_dff_B_14qw1mBa3_0),.dout(w_dff_B_TE2W0Imk6_0),.clk(gclk));
	jdff dff_B_MgAJtuB17_0(.din(w_dff_B_TE2W0Imk6_0),.dout(w_dff_B_MgAJtuB17_0),.clk(gclk));
	jdff dff_B_XGT53Xsq2_0(.din(w_dff_B_MgAJtuB17_0),.dout(w_dff_B_XGT53Xsq2_0),.clk(gclk));
	jdff dff_B_5TxQLPZP6_0(.din(w_dff_B_XGT53Xsq2_0),.dout(w_dff_B_5TxQLPZP6_0),.clk(gclk));
	jdff dff_B_YvLwp3Ut5_0(.din(w_dff_B_5TxQLPZP6_0),.dout(w_dff_B_YvLwp3Ut5_0),.clk(gclk));
	jdff dff_B_ol8bmYDi8_0(.din(w_dff_B_YvLwp3Ut5_0),.dout(w_dff_B_ol8bmYDi8_0),.clk(gclk));
	jdff dff_B_xKAiLwJm3_0(.din(w_dff_B_ol8bmYDi8_0),.dout(w_dff_B_xKAiLwJm3_0),.clk(gclk));
	jdff dff_B_bgj8K81M1_0(.din(w_dff_B_xKAiLwJm3_0),.dout(w_dff_B_bgj8K81M1_0),.clk(gclk));
	jdff dff_B_uxuYl4C17_0(.din(w_dff_B_bgj8K81M1_0),.dout(w_dff_B_uxuYl4C17_0),.clk(gclk));
	jdff dff_B_qSlEKpkG6_0(.din(w_dff_B_uxuYl4C17_0),.dout(w_dff_B_qSlEKpkG6_0),.clk(gclk));
	jdff dff_B_LsxtOyh74_0(.din(w_dff_B_qSlEKpkG6_0),.dout(w_dff_B_LsxtOyh74_0),.clk(gclk));
	jdff dff_B_pa6Wo2BO4_0(.din(w_dff_B_LsxtOyh74_0),.dout(w_dff_B_pa6Wo2BO4_0),.clk(gclk));
	jdff dff_B_OfLeGgiB6_0(.din(w_dff_B_pa6Wo2BO4_0),.dout(w_dff_B_OfLeGgiB6_0),.clk(gclk));
	jdff dff_B_zCGL2FI74_0(.din(w_dff_B_OfLeGgiB6_0),.dout(w_dff_B_zCGL2FI74_0),.clk(gclk));
	jdff dff_B_AnGKKJt33_0(.din(w_dff_B_zCGL2FI74_0),.dout(w_dff_B_AnGKKJt33_0),.clk(gclk));
	jdff dff_B_w6bDZ4HN5_0(.din(w_dff_B_AnGKKJt33_0),.dout(w_dff_B_w6bDZ4HN5_0),.clk(gclk));
	jdff dff_B_Z5lumHrF3_0(.din(w_dff_B_w6bDZ4HN5_0),.dout(w_dff_B_Z5lumHrF3_0),.clk(gclk));
	jdff dff_B_NqhsmJQc3_0(.din(w_dff_B_Z5lumHrF3_0),.dout(w_dff_B_NqhsmJQc3_0),.clk(gclk));
	jdff dff_B_2I9oic4J2_0(.din(w_dff_B_NqhsmJQc3_0),.dout(w_dff_B_2I9oic4J2_0),.clk(gclk));
	jdff dff_B_jE3gGIn46_0(.din(w_dff_B_2I9oic4J2_0),.dout(w_dff_B_jE3gGIn46_0),.clk(gclk));
	jdff dff_B_QmriqQQA9_0(.din(w_dff_B_jE3gGIn46_0),.dout(w_dff_B_QmriqQQA9_0),.clk(gclk));
	jdff dff_B_E02EDSMt1_0(.din(w_dff_B_QmriqQQA9_0),.dout(w_dff_B_E02EDSMt1_0),.clk(gclk));
	jdff dff_B_P2qyRF8K4_0(.din(w_dff_B_E02EDSMt1_0),.dout(w_dff_B_P2qyRF8K4_0),.clk(gclk));
	jdff dff_B_AnUBsgCg0_0(.din(n1132),.dout(w_dff_B_AnUBsgCg0_0),.clk(gclk));
	jdff dff_B_ciRIYHl29_0(.din(w_dff_B_AnUBsgCg0_0),.dout(w_dff_B_ciRIYHl29_0),.clk(gclk));
	jdff dff_B_bjaqF0ZD9_0(.din(w_dff_B_ciRIYHl29_0),.dout(w_dff_B_bjaqF0ZD9_0),.clk(gclk));
	jdff dff_B_7k9h5O3k6_0(.din(w_dff_B_bjaqF0ZD9_0),.dout(w_dff_B_7k9h5O3k6_0),.clk(gclk));
	jdff dff_B_BNluhNy42_0(.din(w_dff_B_7k9h5O3k6_0),.dout(w_dff_B_BNluhNy42_0),.clk(gclk));
	jdff dff_B_QIT3SBBW6_0(.din(w_dff_B_BNluhNy42_0),.dout(w_dff_B_QIT3SBBW6_0),.clk(gclk));
	jdff dff_B_JQzpuMXS8_0(.din(w_dff_B_QIT3SBBW6_0),.dout(w_dff_B_JQzpuMXS8_0),.clk(gclk));
	jdff dff_B_bqCTjpcL9_0(.din(w_dff_B_JQzpuMXS8_0),.dout(w_dff_B_bqCTjpcL9_0),.clk(gclk));
	jdff dff_B_uX9IqRB81_0(.din(w_dff_B_bqCTjpcL9_0),.dout(w_dff_B_uX9IqRB81_0),.clk(gclk));
	jdff dff_B_mzA3Cg8J6_0(.din(w_dff_B_uX9IqRB81_0),.dout(w_dff_B_mzA3Cg8J6_0),.clk(gclk));
	jdff dff_B_xO3KsHO66_0(.din(w_dff_B_mzA3Cg8J6_0),.dout(w_dff_B_xO3KsHO66_0),.clk(gclk));
	jdff dff_B_4SmdUwi71_0(.din(w_dff_B_xO3KsHO66_0),.dout(w_dff_B_4SmdUwi71_0),.clk(gclk));
	jdff dff_B_H8oqT6J93_0(.din(w_dff_B_4SmdUwi71_0),.dout(w_dff_B_H8oqT6J93_0),.clk(gclk));
	jdff dff_B_4XzJK8Gg6_0(.din(w_dff_B_H8oqT6J93_0),.dout(w_dff_B_4XzJK8Gg6_0),.clk(gclk));
	jdff dff_B_1XX0WgBP1_0(.din(w_dff_B_4XzJK8Gg6_0),.dout(w_dff_B_1XX0WgBP1_0),.clk(gclk));
	jdff dff_B_R6YUz3z28_0(.din(w_dff_B_1XX0WgBP1_0),.dout(w_dff_B_R6YUz3z28_0),.clk(gclk));
	jdff dff_B_8yFHfUiN2_0(.din(w_dff_B_R6YUz3z28_0),.dout(w_dff_B_8yFHfUiN2_0),.clk(gclk));
	jdff dff_B_FeM8thi53_0(.din(w_dff_B_8yFHfUiN2_0),.dout(w_dff_B_FeM8thi53_0),.clk(gclk));
	jdff dff_B_F4p0snYn0_0(.din(w_dff_B_FeM8thi53_0),.dout(w_dff_B_F4p0snYn0_0),.clk(gclk));
	jdff dff_B_AU3wcHUQ1_0(.din(w_dff_B_F4p0snYn0_0),.dout(w_dff_B_AU3wcHUQ1_0),.clk(gclk));
	jdff dff_B_3vKBcR4y2_0(.din(w_dff_B_AU3wcHUQ1_0),.dout(w_dff_B_3vKBcR4y2_0),.clk(gclk));
	jdff dff_B_XevCGRFb7_0(.din(w_dff_B_3vKBcR4y2_0),.dout(w_dff_B_XevCGRFb7_0),.clk(gclk));
	jdff dff_B_b9l9YqWJ8_0(.din(w_dff_B_XevCGRFb7_0),.dout(w_dff_B_b9l9YqWJ8_0),.clk(gclk));
	jdff dff_B_3JKDk23U9_0(.din(w_dff_B_b9l9YqWJ8_0),.dout(w_dff_B_3JKDk23U9_0),.clk(gclk));
	jdff dff_B_GdCBevGf7_0(.din(w_dff_B_3JKDk23U9_0),.dout(w_dff_B_GdCBevGf7_0),.clk(gclk));
	jdff dff_B_fjQdDwis8_0(.din(w_dff_B_GdCBevGf7_0),.dout(w_dff_B_fjQdDwis8_0),.clk(gclk));
	jdff dff_B_iOjoLuk30_0(.din(w_dff_B_fjQdDwis8_0),.dout(w_dff_B_iOjoLuk30_0),.clk(gclk));
	jdff dff_B_yVtB9mxq8_0(.din(w_dff_B_iOjoLuk30_0),.dout(w_dff_B_yVtB9mxq8_0),.clk(gclk));
	jdff dff_B_y1DUNIKE2_0(.din(w_dff_B_yVtB9mxq8_0),.dout(w_dff_B_y1DUNIKE2_0),.clk(gclk));
	jdff dff_B_ktNdov5X8_0(.din(w_dff_B_y1DUNIKE2_0),.dout(w_dff_B_ktNdov5X8_0),.clk(gclk));
	jdff dff_B_BKRWFx523_0(.din(w_dff_B_ktNdov5X8_0),.dout(w_dff_B_BKRWFx523_0),.clk(gclk));
	jdff dff_B_EI038q2N7_0(.din(w_dff_B_BKRWFx523_0),.dout(w_dff_B_EI038q2N7_0),.clk(gclk));
	jdff dff_B_b1QayugI9_0(.din(w_dff_B_EI038q2N7_0),.dout(w_dff_B_b1QayugI9_0),.clk(gclk));
	jdff dff_B_gtdu5Yxn6_0(.din(w_dff_B_b1QayugI9_0),.dout(w_dff_B_gtdu5Yxn6_0),.clk(gclk));
	jdff dff_B_7ZLA1AEU3_0(.din(w_dff_B_gtdu5Yxn6_0),.dout(w_dff_B_7ZLA1AEU3_0),.clk(gclk));
	jdff dff_B_kmfv2In99_0(.din(w_dff_B_7ZLA1AEU3_0),.dout(w_dff_B_kmfv2In99_0),.clk(gclk));
	jdff dff_B_qYy2l2GS4_0(.din(w_dff_B_kmfv2In99_0),.dout(w_dff_B_qYy2l2GS4_0),.clk(gclk));
	jdff dff_B_4QyGyHa53_0(.din(w_dff_B_qYy2l2GS4_0),.dout(w_dff_B_4QyGyHa53_0),.clk(gclk));
	jdff dff_B_z3YLYRms7_0(.din(w_dff_B_4QyGyHa53_0),.dout(w_dff_B_z3YLYRms7_0),.clk(gclk));
	jdff dff_B_uq6nkgFO0_0(.din(w_dff_B_z3YLYRms7_0),.dout(w_dff_B_uq6nkgFO0_0),.clk(gclk));
	jdff dff_B_EVYUVjSW2_0(.din(w_dff_B_uq6nkgFO0_0),.dout(w_dff_B_EVYUVjSW2_0),.clk(gclk));
	jdff dff_B_Yyrez7Fi4_0(.din(w_dff_B_EVYUVjSW2_0),.dout(w_dff_B_Yyrez7Fi4_0),.clk(gclk));
	jdff dff_B_bkkM4V7I5_0(.din(w_dff_B_Yyrez7Fi4_0),.dout(w_dff_B_bkkM4V7I5_0),.clk(gclk));
	jdff dff_B_SSO2b7TT0_0(.din(w_dff_B_bkkM4V7I5_0),.dout(w_dff_B_SSO2b7TT0_0),.clk(gclk));
	jdff dff_B_4ybstWh80_0(.din(w_dff_B_SSO2b7TT0_0),.dout(w_dff_B_4ybstWh80_0),.clk(gclk));
	jdff dff_B_2xbCP0oy1_0(.din(w_dff_B_4ybstWh80_0),.dout(w_dff_B_2xbCP0oy1_0),.clk(gclk));
	jdff dff_B_6wLIYx6m8_0(.din(w_dff_B_2xbCP0oy1_0),.dout(w_dff_B_6wLIYx6m8_0),.clk(gclk));
	jdff dff_B_Dj6JnDZ11_0(.din(w_dff_B_6wLIYx6m8_0),.dout(w_dff_B_Dj6JnDZ11_0),.clk(gclk));
	jdff dff_B_lHMxqmMG1_0(.din(w_dff_B_Dj6JnDZ11_0),.dout(w_dff_B_lHMxqmMG1_0),.clk(gclk));
	jdff dff_B_Lu0eTXOt5_0(.din(w_dff_B_lHMxqmMG1_0),.dout(w_dff_B_Lu0eTXOt5_0),.clk(gclk));
	jdff dff_B_M8n3SWsm2_0(.din(w_dff_B_Lu0eTXOt5_0),.dout(w_dff_B_M8n3SWsm2_0),.clk(gclk));
	jdff dff_B_QFKVtpy08_0(.din(w_dff_B_M8n3SWsm2_0),.dout(w_dff_B_QFKVtpy08_0),.clk(gclk));
	jdff dff_B_W9RkfTyR1_0(.din(w_dff_B_QFKVtpy08_0),.dout(w_dff_B_W9RkfTyR1_0),.clk(gclk));
	jdff dff_B_WqYsR6aj0_0(.din(w_dff_B_W9RkfTyR1_0),.dout(w_dff_B_WqYsR6aj0_0),.clk(gclk));
	jdff dff_B_JG6RM1k87_0(.din(w_dff_B_WqYsR6aj0_0),.dout(w_dff_B_JG6RM1k87_0),.clk(gclk));
	jdff dff_B_rtgGt7my7_0(.din(w_dff_B_JG6RM1k87_0),.dout(w_dff_B_rtgGt7my7_0),.clk(gclk));
	jdff dff_B_QlndlzQS4_0(.din(w_dff_B_rtgGt7my7_0),.dout(w_dff_B_QlndlzQS4_0),.clk(gclk));
	jdff dff_B_du85iw1C5_0(.din(w_dff_B_QlndlzQS4_0),.dout(w_dff_B_du85iw1C5_0),.clk(gclk));
	jdff dff_B_s14OcBtD5_0(.din(w_dff_B_du85iw1C5_0),.dout(w_dff_B_s14OcBtD5_0),.clk(gclk));
	jdff dff_B_tidPtZPJ4_0(.din(w_dff_B_s14OcBtD5_0),.dout(w_dff_B_tidPtZPJ4_0),.clk(gclk));
	jdff dff_B_VZw7honL6_0(.din(w_dff_B_tidPtZPJ4_0),.dout(w_dff_B_VZw7honL6_0),.clk(gclk));
	jdff dff_B_TT45QkOS2_0(.din(w_dff_B_VZw7honL6_0),.dout(w_dff_B_TT45QkOS2_0),.clk(gclk));
	jdff dff_B_bjiHRgdS3_0(.din(w_dff_B_TT45QkOS2_0),.dout(w_dff_B_bjiHRgdS3_0),.clk(gclk));
	jdff dff_B_Ss7i2Bw90_0(.din(w_dff_B_bjiHRgdS3_0),.dout(w_dff_B_Ss7i2Bw90_0),.clk(gclk));
	jdff dff_B_0zDidFUn2_0(.din(w_dff_B_Ss7i2Bw90_0),.dout(w_dff_B_0zDidFUn2_0),.clk(gclk));
	jdff dff_B_Qek5J5k80_0(.din(w_dff_B_0zDidFUn2_0),.dout(w_dff_B_Qek5J5k80_0),.clk(gclk));
	jdff dff_B_0QfYaqb86_0(.din(w_dff_B_Qek5J5k80_0),.dout(w_dff_B_0QfYaqb86_0),.clk(gclk));
	jdff dff_B_o9yTFobN5_0(.din(w_dff_B_0QfYaqb86_0),.dout(w_dff_B_o9yTFobN5_0),.clk(gclk));
	jdff dff_B_n0xpXh2y6_0(.din(w_dff_B_o9yTFobN5_0),.dout(w_dff_B_n0xpXh2y6_0),.clk(gclk));
	jdff dff_B_Ajd5YtvK8_0(.din(w_dff_B_n0xpXh2y6_0),.dout(w_dff_B_Ajd5YtvK8_0),.clk(gclk));
	jdff dff_B_FskJtOUr8_0(.din(w_dff_B_Ajd5YtvK8_0),.dout(w_dff_B_FskJtOUr8_0),.clk(gclk));
	jdff dff_B_b30rvFHq0_0(.din(w_dff_B_FskJtOUr8_0),.dout(w_dff_B_b30rvFHq0_0),.clk(gclk));
	jdff dff_B_pGdrETgs8_0(.din(w_dff_B_b30rvFHq0_0),.dout(w_dff_B_pGdrETgs8_0),.clk(gclk));
	jdff dff_B_7icUPGR23_0(.din(w_dff_B_pGdrETgs8_0),.dout(w_dff_B_7icUPGR23_0),.clk(gclk));
	jdff dff_B_L2IWobFb8_0(.din(w_dff_B_7icUPGR23_0),.dout(w_dff_B_L2IWobFb8_0),.clk(gclk));
	jdff dff_B_0t8LD5oz6_0(.din(w_dff_B_L2IWobFb8_0),.dout(w_dff_B_0t8LD5oz6_0),.clk(gclk));
	jdff dff_B_YvoUw0471_0(.din(w_dff_B_0t8LD5oz6_0),.dout(w_dff_B_YvoUw0471_0),.clk(gclk));
	jdff dff_B_f7FrN3YU6_0(.din(w_dff_B_YvoUw0471_0),.dout(w_dff_B_f7FrN3YU6_0),.clk(gclk));
	jdff dff_B_Y1DsgdCH2_0(.din(w_dff_B_f7FrN3YU6_0),.dout(w_dff_B_Y1DsgdCH2_0),.clk(gclk));
	jdff dff_B_aESggMQI6_0(.din(w_dff_B_Y1DsgdCH2_0),.dout(w_dff_B_aESggMQI6_0),.clk(gclk));
	jdff dff_B_SsLNApqS7_0(.din(w_dff_B_aESggMQI6_0),.dout(w_dff_B_SsLNApqS7_0),.clk(gclk));
	jdff dff_B_aBvX1duK8_0(.din(w_dff_B_SsLNApqS7_0),.dout(w_dff_B_aBvX1duK8_0),.clk(gclk));
	jdff dff_B_MuOTdBbz6_0(.din(w_dff_B_aBvX1duK8_0),.dout(w_dff_B_MuOTdBbz6_0),.clk(gclk));
	jdff dff_B_sui8Kq456_0(.din(w_dff_B_MuOTdBbz6_0),.dout(w_dff_B_sui8Kq456_0),.clk(gclk));
	jdff dff_B_PcdbTwvc7_0(.din(w_dff_B_sui8Kq456_0),.dout(w_dff_B_PcdbTwvc7_0),.clk(gclk));
	jdff dff_B_aNnGcEt09_0(.din(w_dff_B_PcdbTwvc7_0),.dout(w_dff_B_aNnGcEt09_0),.clk(gclk));
	jdff dff_B_PU1wLCQP7_0(.din(w_dff_B_aNnGcEt09_0),.dout(w_dff_B_PU1wLCQP7_0),.clk(gclk));
	jdff dff_B_n7s0thyv7_0(.din(w_dff_B_PU1wLCQP7_0),.dout(w_dff_B_n7s0thyv7_0),.clk(gclk));
	jdff dff_B_3QDAHMmj4_0(.din(w_dff_B_n7s0thyv7_0),.dout(w_dff_B_3QDAHMmj4_0),.clk(gclk));
	jdff dff_B_QlbG0Nm58_0(.din(w_dff_B_3QDAHMmj4_0),.dout(w_dff_B_QlbG0Nm58_0),.clk(gclk));
	jdff dff_B_kdyOUyGn4_0(.din(w_dff_B_QlbG0Nm58_0),.dout(w_dff_B_kdyOUyGn4_0),.clk(gclk));
	jdff dff_B_RZbOA3Em1_0(.din(w_dff_B_kdyOUyGn4_0),.dout(w_dff_B_RZbOA3Em1_0),.clk(gclk));
	jdff dff_B_TSji5Tyv4_0(.din(w_dff_B_RZbOA3Em1_0),.dout(w_dff_B_TSji5Tyv4_0),.clk(gclk));
	jdff dff_B_DB401HXm8_0(.din(w_dff_B_TSji5Tyv4_0),.dout(w_dff_B_DB401HXm8_0),.clk(gclk));
	jdff dff_B_eFVXScsq6_0(.din(w_dff_B_DB401HXm8_0),.dout(w_dff_B_eFVXScsq6_0),.clk(gclk));
	jdff dff_B_sEGwsu4a0_0(.din(w_dff_B_eFVXScsq6_0),.dout(w_dff_B_sEGwsu4a0_0),.clk(gclk));
	jdff dff_B_AF3T9QpX6_0(.din(w_dff_B_sEGwsu4a0_0),.dout(w_dff_B_AF3T9QpX6_0),.clk(gclk));
	jdff dff_B_i4xc8eaS5_0(.din(w_dff_B_AF3T9QpX6_0),.dout(w_dff_B_i4xc8eaS5_0),.clk(gclk));
	jdff dff_B_YZX0D7ZM2_0(.din(w_dff_B_i4xc8eaS5_0),.dout(w_dff_B_YZX0D7ZM2_0),.clk(gclk));
	jdff dff_B_07X3RyDd9_0(.din(w_dff_B_YZX0D7ZM2_0),.dout(w_dff_B_07X3RyDd9_0),.clk(gclk));
	jdff dff_B_Q8QjIA982_0(.din(w_dff_B_07X3RyDd9_0),.dout(w_dff_B_Q8QjIA982_0),.clk(gclk));
	jdff dff_B_0ji4sAsF1_0(.din(w_dff_B_Q8QjIA982_0),.dout(w_dff_B_0ji4sAsF1_0),.clk(gclk));
	jdff dff_B_caf0nWoP4_0(.din(w_dff_B_0ji4sAsF1_0),.dout(w_dff_B_caf0nWoP4_0),.clk(gclk));
	jdff dff_B_cEKkY6bt2_0(.din(w_dff_B_caf0nWoP4_0),.dout(w_dff_B_cEKkY6bt2_0),.clk(gclk));
	jdff dff_B_hTmF8Qd97_0(.din(w_dff_B_cEKkY6bt2_0),.dout(w_dff_B_hTmF8Qd97_0),.clk(gclk));
	jdff dff_B_38UupXcB0_0(.din(w_dff_B_hTmF8Qd97_0),.dout(w_dff_B_38UupXcB0_0),.clk(gclk));
	jdff dff_B_rHs3VIWw9_0(.din(w_dff_B_38UupXcB0_0),.dout(w_dff_B_rHs3VIWw9_0),.clk(gclk));
	jdff dff_B_DsdfOOoK5_0(.din(w_dff_B_rHs3VIWw9_0),.dout(w_dff_B_DsdfOOoK5_0),.clk(gclk));
	jdff dff_B_LWTCzuch2_0(.din(w_dff_B_DsdfOOoK5_0),.dout(w_dff_B_LWTCzuch2_0),.clk(gclk));
	jdff dff_B_wNh2ztIJ3_0(.din(w_dff_B_LWTCzuch2_0),.dout(w_dff_B_wNh2ztIJ3_0),.clk(gclk));
	jdff dff_B_d7f7UIjm7_0(.din(w_dff_B_wNh2ztIJ3_0),.dout(w_dff_B_d7f7UIjm7_0),.clk(gclk));
	jdff dff_B_OQgYeVkg6_0(.din(w_dff_B_d7f7UIjm7_0),.dout(w_dff_B_OQgYeVkg6_0),.clk(gclk));
	jdff dff_B_GKypNqJd2_0(.din(w_dff_B_OQgYeVkg6_0),.dout(w_dff_B_GKypNqJd2_0),.clk(gclk));
	jdff dff_B_qvwEj2Hf4_0(.din(w_dff_B_GKypNqJd2_0),.dout(w_dff_B_qvwEj2Hf4_0),.clk(gclk));
	jdff dff_B_YpJDZxaE6_0(.din(w_dff_B_qvwEj2Hf4_0),.dout(w_dff_B_YpJDZxaE6_0),.clk(gclk));
	jdff dff_B_Ucig1agG3_0(.din(w_dff_B_YpJDZxaE6_0),.dout(w_dff_B_Ucig1agG3_0),.clk(gclk));
	jdff dff_B_u9OY4RPb0_0(.din(w_dff_B_Ucig1agG3_0),.dout(w_dff_B_u9OY4RPb0_0),.clk(gclk));
	jdff dff_B_uNC1l8Z80_0(.din(w_dff_B_u9OY4RPb0_0),.dout(w_dff_B_uNC1l8Z80_0),.clk(gclk));
	jdff dff_B_8U7G98lZ4_0(.din(w_dff_B_uNC1l8Z80_0),.dout(w_dff_B_8U7G98lZ4_0),.clk(gclk));
	jdff dff_B_YEsUQv1B3_0(.din(w_dff_B_8U7G98lZ4_0),.dout(w_dff_B_YEsUQv1B3_0),.clk(gclk));
	jdff dff_B_VxjKO3032_0(.din(w_dff_B_YEsUQv1B3_0),.dout(w_dff_B_VxjKO3032_0),.clk(gclk));
	jdff dff_B_KCv9h0wh2_0(.din(w_dff_B_VxjKO3032_0),.dout(w_dff_B_KCv9h0wh2_0),.clk(gclk));
	jdff dff_B_XuMixnZF9_0(.din(w_dff_B_KCv9h0wh2_0),.dout(w_dff_B_XuMixnZF9_0),.clk(gclk));
	jdff dff_B_i84eCWYK5_0(.din(w_dff_B_XuMixnZF9_0),.dout(w_dff_B_i84eCWYK5_0),.clk(gclk));
	jdff dff_B_U6iwCUZI0_0(.din(n1138),.dout(w_dff_B_U6iwCUZI0_0),.clk(gclk));
	jdff dff_B_a5doqkpu9_0(.din(w_dff_B_U6iwCUZI0_0),.dout(w_dff_B_a5doqkpu9_0),.clk(gclk));
	jdff dff_B_57llpIob9_0(.din(w_dff_B_a5doqkpu9_0),.dout(w_dff_B_57llpIob9_0),.clk(gclk));
	jdff dff_B_7vRhbgR89_0(.din(w_dff_B_57llpIob9_0),.dout(w_dff_B_7vRhbgR89_0),.clk(gclk));
	jdff dff_B_oEK9mALP8_0(.din(w_dff_B_7vRhbgR89_0),.dout(w_dff_B_oEK9mALP8_0),.clk(gclk));
	jdff dff_B_vIkxOLPx8_0(.din(w_dff_B_oEK9mALP8_0),.dout(w_dff_B_vIkxOLPx8_0),.clk(gclk));
	jdff dff_B_E6iKKrI60_0(.din(w_dff_B_vIkxOLPx8_0),.dout(w_dff_B_E6iKKrI60_0),.clk(gclk));
	jdff dff_B_Uyuf2mfa0_0(.din(w_dff_B_E6iKKrI60_0),.dout(w_dff_B_Uyuf2mfa0_0),.clk(gclk));
	jdff dff_B_1Xzww8T78_0(.din(w_dff_B_Uyuf2mfa0_0),.dout(w_dff_B_1Xzww8T78_0),.clk(gclk));
	jdff dff_B_njK3vFMj2_0(.din(w_dff_B_1Xzww8T78_0),.dout(w_dff_B_njK3vFMj2_0),.clk(gclk));
	jdff dff_B_HhC6SGrG6_0(.din(w_dff_B_njK3vFMj2_0),.dout(w_dff_B_HhC6SGrG6_0),.clk(gclk));
	jdff dff_B_TMD9qqX40_0(.din(w_dff_B_HhC6SGrG6_0),.dout(w_dff_B_TMD9qqX40_0),.clk(gclk));
	jdff dff_B_sGe1J2sr6_0(.din(w_dff_B_TMD9qqX40_0),.dout(w_dff_B_sGe1J2sr6_0),.clk(gclk));
	jdff dff_B_WgXCP8oB1_0(.din(w_dff_B_sGe1J2sr6_0),.dout(w_dff_B_WgXCP8oB1_0),.clk(gclk));
	jdff dff_B_WOjvGSCr8_0(.din(w_dff_B_WgXCP8oB1_0),.dout(w_dff_B_WOjvGSCr8_0),.clk(gclk));
	jdff dff_B_zakEMstQ7_0(.din(w_dff_B_WOjvGSCr8_0),.dout(w_dff_B_zakEMstQ7_0),.clk(gclk));
	jdff dff_B_ss1rzqcX8_0(.din(w_dff_B_zakEMstQ7_0),.dout(w_dff_B_ss1rzqcX8_0),.clk(gclk));
	jdff dff_B_6NJbhcMc8_0(.din(w_dff_B_ss1rzqcX8_0),.dout(w_dff_B_6NJbhcMc8_0),.clk(gclk));
	jdff dff_B_gEKVGIrr0_0(.din(w_dff_B_6NJbhcMc8_0),.dout(w_dff_B_gEKVGIrr0_0),.clk(gclk));
	jdff dff_B_TeeUhAJH4_0(.din(w_dff_B_gEKVGIrr0_0),.dout(w_dff_B_TeeUhAJH4_0),.clk(gclk));
	jdff dff_B_pwRMvVCF2_0(.din(w_dff_B_TeeUhAJH4_0),.dout(w_dff_B_pwRMvVCF2_0),.clk(gclk));
	jdff dff_B_0Btbh8ue2_0(.din(w_dff_B_pwRMvVCF2_0),.dout(w_dff_B_0Btbh8ue2_0),.clk(gclk));
	jdff dff_B_REEkhnWJ6_0(.din(w_dff_B_0Btbh8ue2_0),.dout(w_dff_B_REEkhnWJ6_0),.clk(gclk));
	jdff dff_B_osRhnc4L7_0(.din(w_dff_B_REEkhnWJ6_0),.dout(w_dff_B_osRhnc4L7_0),.clk(gclk));
	jdff dff_B_urmRmVsn4_0(.din(w_dff_B_osRhnc4L7_0),.dout(w_dff_B_urmRmVsn4_0),.clk(gclk));
	jdff dff_B_DyS7xSXY7_0(.din(w_dff_B_urmRmVsn4_0),.dout(w_dff_B_DyS7xSXY7_0),.clk(gclk));
	jdff dff_B_NRtyQ9LL2_0(.din(w_dff_B_DyS7xSXY7_0),.dout(w_dff_B_NRtyQ9LL2_0),.clk(gclk));
	jdff dff_B_pSYE8h1n8_0(.din(w_dff_B_NRtyQ9LL2_0),.dout(w_dff_B_pSYE8h1n8_0),.clk(gclk));
	jdff dff_B_CWAAsrHB5_0(.din(w_dff_B_pSYE8h1n8_0),.dout(w_dff_B_CWAAsrHB5_0),.clk(gclk));
	jdff dff_B_j4qLCyvR0_0(.din(w_dff_B_CWAAsrHB5_0),.dout(w_dff_B_j4qLCyvR0_0),.clk(gclk));
	jdff dff_B_AfDCJyYt4_0(.din(w_dff_B_j4qLCyvR0_0),.dout(w_dff_B_AfDCJyYt4_0),.clk(gclk));
	jdff dff_B_Rrv7Kelz8_0(.din(w_dff_B_AfDCJyYt4_0),.dout(w_dff_B_Rrv7Kelz8_0),.clk(gclk));
	jdff dff_B_qX4CVjCr3_0(.din(w_dff_B_Rrv7Kelz8_0),.dout(w_dff_B_qX4CVjCr3_0),.clk(gclk));
	jdff dff_B_CAupgnU25_0(.din(w_dff_B_qX4CVjCr3_0),.dout(w_dff_B_CAupgnU25_0),.clk(gclk));
	jdff dff_B_0a5auGct7_0(.din(w_dff_B_CAupgnU25_0),.dout(w_dff_B_0a5auGct7_0),.clk(gclk));
	jdff dff_B_OstfHIGV8_0(.din(w_dff_B_0a5auGct7_0),.dout(w_dff_B_OstfHIGV8_0),.clk(gclk));
	jdff dff_B_JlgY5HaC6_0(.din(w_dff_B_OstfHIGV8_0),.dout(w_dff_B_JlgY5HaC6_0),.clk(gclk));
	jdff dff_B_CArRZfBW6_0(.din(w_dff_B_JlgY5HaC6_0),.dout(w_dff_B_CArRZfBW6_0),.clk(gclk));
	jdff dff_B_LhDuKVVU8_0(.din(w_dff_B_CArRZfBW6_0),.dout(w_dff_B_LhDuKVVU8_0),.clk(gclk));
	jdff dff_B_5FrZBA1s4_0(.din(w_dff_B_LhDuKVVU8_0),.dout(w_dff_B_5FrZBA1s4_0),.clk(gclk));
	jdff dff_B_XQ9Rjv7h6_0(.din(w_dff_B_5FrZBA1s4_0),.dout(w_dff_B_XQ9Rjv7h6_0),.clk(gclk));
	jdff dff_B_a8gC8uVN9_0(.din(w_dff_B_XQ9Rjv7h6_0),.dout(w_dff_B_a8gC8uVN9_0),.clk(gclk));
	jdff dff_B_483hyO8g4_0(.din(w_dff_B_a8gC8uVN9_0),.dout(w_dff_B_483hyO8g4_0),.clk(gclk));
	jdff dff_B_qEAYffRl1_0(.din(w_dff_B_483hyO8g4_0),.dout(w_dff_B_qEAYffRl1_0),.clk(gclk));
	jdff dff_B_kcLCUR772_0(.din(w_dff_B_qEAYffRl1_0),.dout(w_dff_B_kcLCUR772_0),.clk(gclk));
	jdff dff_B_7szMmokO0_0(.din(w_dff_B_kcLCUR772_0),.dout(w_dff_B_7szMmokO0_0),.clk(gclk));
	jdff dff_B_KMCHcUBV0_0(.din(w_dff_B_7szMmokO0_0),.dout(w_dff_B_KMCHcUBV0_0),.clk(gclk));
	jdff dff_B_heNREE0Y6_0(.din(w_dff_B_KMCHcUBV0_0),.dout(w_dff_B_heNREE0Y6_0),.clk(gclk));
	jdff dff_B_H6bPQElY1_0(.din(w_dff_B_heNREE0Y6_0),.dout(w_dff_B_H6bPQElY1_0),.clk(gclk));
	jdff dff_B_gz2OrYPI9_0(.din(w_dff_B_H6bPQElY1_0),.dout(w_dff_B_gz2OrYPI9_0),.clk(gclk));
	jdff dff_B_nAxAlxz78_0(.din(w_dff_B_gz2OrYPI9_0),.dout(w_dff_B_nAxAlxz78_0),.clk(gclk));
	jdff dff_B_5wyFce4n6_0(.din(w_dff_B_nAxAlxz78_0),.dout(w_dff_B_5wyFce4n6_0),.clk(gclk));
	jdff dff_B_quUKTcuk1_0(.din(w_dff_B_5wyFce4n6_0),.dout(w_dff_B_quUKTcuk1_0),.clk(gclk));
	jdff dff_B_oPL44UVW6_0(.din(w_dff_B_quUKTcuk1_0),.dout(w_dff_B_oPL44UVW6_0),.clk(gclk));
	jdff dff_B_iE6Jz1SW3_0(.din(w_dff_B_oPL44UVW6_0),.dout(w_dff_B_iE6Jz1SW3_0),.clk(gclk));
	jdff dff_B_DE3XsQ635_0(.din(w_dff_B_iE6Jz1SW3_0),.dout(w_dff_B_DE3XsQ635_0),.clk(gclk));
	jdff dff_B_jnOUUyph7_0(.din(w_dff_B_DE3XsQ635_0),.dout(w_dff_B_jnOUUyph7_0),.clk(gclk));
	jdff dff_B_nn041RUC8_0(.din(w_dff_B_jnOUUyph7_0),.dout(w_dff_B_nn041RUC8_0),.clk(gclk));
	jdff dff_B_Ott5IRF98_0(.din(w_dff_B_nn041RUC8_0),.dout(w_dff_B_Ott5IRF98_0),.clk(gclk));
	jdff dff_B_abhOlZYA7_0(.din(w_dff_B_Ott5IRF98_0),.dout(w_dff_B_abhOlZYA7_0),.clk(gclk));
	jdff dff_B_lQFKS9cz2_0(.din(w_dff_B_abhOlZYA7_0),.dout(w_dff_B_lQFKS9cz2_0),.clk(gclk));
	jdff dff_B_M9azyQZp9_0(.din(w_dff_B_lQFKS9cz2_0),.dout(w_dff_B_M9azyQZp9_0),.clk(gclk));
	jdff dff_B_0H2INgDW0_0(.din(w_dff_B_M9azyQZp9_0),.dout(w_dff_B_0H2INgDW0_0),.clk(gclk));
	jdff dff_B_ZiTnUagd1_0(.din(w_dff_B_0H2INgDW0_0),.dout(w_dff_B_ZiTnUagd1_0),.clk(gclk));
	jdff dff_B_CbJ52ZMk7_0(.din(w_dff_B_ZiTnUagd1_0),.dout(w_dff_B_CbJ52ZMk7_0),.clk(gclk));
	jdff dff_B_PQxVaC210_0(.din(w_dff_B_CbJ52ZMk7_0),.dout(w_dff_B_PQxVaC210_0),.clk(gclk));
	jdff dff_B_OR5nETYs0_0(.din(w_dff_B_PQxVaC210_0),.dout(w_dff_B_OR5nETYs0_0),.clk(gclk));
	jdff dff_B_T319vpfa4_0(.din(w_dff_B_OR5nETYs0_0),.dout(w_dff_B_T319vpfa4_0),.clk(gclk));
	jdff dff_B_f8akAoUd3_0(.din(w_dff_B_T319vpfa4_0),.dout(w_dff_B_f8akAoUd3_0),.clk(gclk));
	jdff dff_B_qyLKJi1A2_0(.din(w_dff_B_f8akAoUd3_0),.dout(w_dff_B_qyLKJi1A2_0),.clk(gclk));
	jdff dff_B_aC6sKNmO2_0(.din(w_dff_B_qyLKJi1A2_0),.dout(w_dff_B_aC6sKNmO2_0),.clk(gclk));
	jdff dff_B_8d2RFYTT9_0(.din(w_dff_B_aC6sKNmO2_0),.dout(w_dff_B_8d2RFYTT9_0),.clk(gclk));
	jdff dff_B_i0l3dmF45_0(.din(w_dff_B_8d2RFYTT9_0),.dout(w_dff_B_i0l3dmF45_0),.clk(gclk));
	jdff dff_B_byNuTY3P8_0(.din(w_dff_B_i0l3dmF45_0),.dout(w_dff_B_byNuTY3P8_0),.clk(gclk));
	jdff dff_B_XmlN3y7k5_0(.din(w_dff_B_byNuTY3P8_0),.dout(w_dff_B_XmlN3y7k5_0),.clk(gclk));
	jdff dff_B_kTjdueIQ1_0(.din(w_dff_B_XmlN3y7k5_0),.dout(w_dff_B_kTjdueIQ1_0),.clk(gclk));
	jdff dff_B_1psdxSCW2_0(.din(w_dff_B_kTjdueIQ1_0),.dout(w_dff_B_1psdxSCW2_0),.clk(gclk));
	jdff dff_B_WdQRaDsG6_0(.din(w_dff_B_1psdxSCW2_0),.dout(w_dff_B_WdQRaDsG6_0),.clk(gclk));
	jdff dff_B_t91WNSGm1_0(.din(w_dff_B_WdQRaDsG6_0),.dout(w_dff_B_t91WNSGm1_0),.clk(gclk));
	jdff dff_B_IEwWzTiz3_0(.din(w_dff_B_t91WNSGm1_0),.dout(w_dff_B_IEwWzTiz3_0),.clk(gclk));
	jdff dff_B_mf48kb8J1_0(.din(w_dff_B_IEwWzTiz3_0),.dout(w_dff_B_mf48kb8J1_0),.clk(gclk));
	jdff dff_B_AeV4wvcd9_0(.din(w_dff_B_mf48kb8J1_0),.dout(w_dff_B_AeV4wvcd9_0),.clk(gclk));
	jdff dff_B_PJyJoXTf0_0(.din(w_dff_B_AeV4wvcd9_0),.dout(w_dff_B_PJyJoXTf0_0),.clk(gclk));
	jdff dff_B_t74qSl9a8_0(.din(w_dff_B_PJyJoXTf0_0),.dout(w_dff_B_t74qSl9a8_0),.clk(gclk));
	jdff dff_B_IZc4wbgh8_0(.din(w_dff_B_t74qSl9a8_0),.dout(w_dff_B_IZc4wbgh8_0),.clk(gclk));
	jdff dff_B_KbFwBhXd3_0(.din(w_dff_B_IZc4wbgh8_0),.dout(w_dff_B_KbFwBhXd3_0),.clk(gclk));
	jdff dff_B_oV4kSYUM3_0(.din(w_dff_B_KbFwBhXd3_0),.dout(w_dff_B_oV4kSYUM3_0),.clk(gclk));
	jdff dff_B_71zA2kTt4_0(.din(w_dff_B_oV4kSYUM3_0),.dout(w_dff_B_71zA2kTt4_0),.clk(gclk));
	jdff dff_B_3ieDKJEX2_0(.din(w_dff_B_71zA2kTt4_0),.dout(w_dff_B_3ieDKJEX2_0),.clk(gclk));
	jdff dff_B_goPzpxyf9_0(.din(w_dff_B_3ieDKJEX2_0),.dout(w_dff_B_goPzpxyf9_0),.clk(gclk));
	jdff dff_B_8fhEuSZk1_0(.din(w_dff_B_goPzpxyf9_0),.dout(w_dff_B_8fhEuSZk1_0),.clk(gclk));
	jdff dff_B_QdgWjF0B1_0(.din(w_dff_B_8fhEuSZk1_0),.dout(w_dff_B_QdgWjF0B1_0),.clk(gclk));
	jdff dff_B_9spmQcSQ7_0(.din(w_dff_B_QdgWjF0B1_0),.dout(w_dff_B_9spmQcSQ7_0),.clk(gclk));
	jdff dff_B_wvt8aCLK8_0(.din(w_dff_B_9spmQcSQ7_0),.dout(w_dff_B_wvt8aCLK8_0),.clk(gclk));
	jdff dff_B_LHvcpfcj5_0(.din(w_dff_B_wvt8aCLK8_0),.dout(w_dff_B_LHvcpfcj5_0),.clk(gclk));
	jdff dff_B_MkSo5soc6_0(.din(w_dff_B_LHvcpfcj5_0),.dout(w_dff_B_MkSo5soc6_0),.clk(gclk));
	jdff dff_B_Z36m5uF72_0(.din(w_dff_B_MkSo5soc6_0),.dout(w_dff_B_Z36m5uF72_0),.clk(gclk));
	jdff dff_B_4RoGkf3r2_0(.din(w_dff_B_Z36m5uF72_0),.dout(w_dff_B_4RoGkf3r2_0),.clk(gclk));
	jdff dff_B_hFDQBF8z9_0(.din(w_dff_B_4RoGkf3r2_0),.dout(w_dff_B_hFDQBF8z9_0),.clk(gclk));
	jdff dff_B_AeXMupvd9_0(.din(w_dff_B_hFDQBF8z9_0),.dout(w_dff_B_AeXMupvd9_0),.clk(gclk));
	jdff dff_B_B3apuCFj8_0(.din(w_dff_B_AeXMupvd9_0),.dout(w_dff_B_B3apuCFj8_0),.clk(gclk));
	jdff dff_B_prjaBGQ89_0(.din(w_dff_B_B3apuCFj8_0),.dout(w_dff_B_prjaBGQ89_0),.clk(gclk));
	jdff dff_B_OMpeXpLq6_0(.din(w_dff_B_prjaBGQ89_0),.dout(w_dff_B_OMpeXpLq6_0),.clk(gclk));
	jdff dff_B_g1TsJgxk4_0(.din(w_dff_B_OMpeXpLq6_0),.dout(w_dff_B_g1TsJgxk4_0),.clk(gclk));
	jdff dff_B_mUKxOZ513_0(.din(w_dff_B_g1TsJgxk4_0),.dout(w_dff_B_mUKxOZ513_0),.clk(gclk));
	jdff dff_B_SeZRqgZB9_0(.din(w_dff_B_mUKxOZ513_0),.dout(w_dff_B_SeZRqgZB9_0),.clk(gclk));
	jdff dff_B_wSkievnF8_0(.din(w_dff_B_SeZRqgZB9_0),.dout(w_dff_B_wSkievnF8_0),.clk(gclk));
	jdff dff_B_s2zO63RE6_0(.din(w_dff_B_wSkievnF8_0),.dout(w_dff_B_s2zO63RE6_0),.clk(gclk));
	jdff dff_B_tyiABXnk7_0(.din(w_dff_B_s2zO63RE6_0),.dout(w_dff_B_tyiABXnk7_0),.clk(gclk));
	jdff dff_B_PkwEA4Rc9_0(.din(w_dff_B_tyiABXnk7_0),.dout(w_dff_B_PkwEA4Rc9_0),.clk(gclk));
	jdff dff_B_gVaUN1NU5_0(.din(w_dff_B_PkwEA4Rc9_0),.dout(w_dff_B_gVaUN1NU5_0),.clk(gclk));
	jdff dff_B_9P7yv7Ye7_0(.din(w_dff_B_gVaUN1NU5_0),.dout(w_dff_B_9P7yv7Ye7_0),.clk(gclk));
	jdff dff_B_Vr9tWKYM4_0(.din(w_dff_B_9P7yv7Ye7_0),.dout(w_dff_B_Vr9tWKYM4_0),.clk(gclk));
	jdff dff_B_yp9b0hnF4_0(.din(w_dff_B_Vr9tWKYM4_0),.dout(w_dff_B_yp9b0hnF4_0),.clk(gclk));
	jdff dff_B_1D79UTZf5_0(.din(w_dff_B_yp9b0hnF4_0),.dout(w_dff_B_1D79UTZf5_0),.clk(gclk));
	jdff dff_B_VAj705Ce6_0(.din(w_dff_B_1D79UTZf5_0),.dout(w_dff_B_VAj705Ce6_0),.clk(gclk));
	jdff dff_B_qTwxy58w0_0(.din(w_dff_B_VAj705Ce6_0),.dout(w_dff_B_qTwxy58w0_0),.clk(gclk));
	jdff dff_B_e8dfjaRZ9_0(.din(w_dff_B_qTwxy58w0_0),.dout(w_dff_B_e8dfjaRZ9_0),.clk(gclk));
	jdff dff_B_FJS06Muv8_0(.din(w_dff_B_e8dfjaRZ9_0),.dout(w_dff_B_FJS06Muv8_0),.clk(gclk));
	jdff dff_B_eMzPEEbX4_0(.din(w_dff_B_FJS06Muv8_0),.dout(w_dff_B_eMzPEEbX4_0),.clk(gclk));
	jdff dff_B_gXpXSEfj8_0(.din(w_dff_B_eMzPEEbX4_0),.dout(w_dff_B_gXpXSEfj8_0),.clk(gclk));
	jdff dff_B_lewfv43k5_0(.din(w_dff_B_gXpXSEfj8_0),.dout(w_dff_B_lewfv43k5_0),.clk(gclk));
	jdff dff_B_xIRT4pZK3_0(.din(w_dff_B_lewfv43k5_0),.dout(w_dff_B_xIRT4pZK3_0),.clk(gclk));
	jdff dff_B_MT6YAPpC5_0(.din(w_dff_B_xIRT4pZK3_0),.dout(w_dff_B_MT6YAPpC5_0),.clk(gclk));
	jdff dff_B_3xJzgs0k4_0(.din(w_dff_B_MT6YAPpC5_0),.dout(w_dff_B_3xJzgs0k4_0),.clk(gclk));
	jdff dff_B_HjcxW1gs6_0(.din(n1144),.dout(w_dff_B_HjcxW1gs6_0),.clk(gclk));
	jdff dff_B_EzdcUTXM9_0(.din(w_dff_B_HjcxW1gs6_0),.dout(w_dff_B_EzdcUTXM9_0),.clk(gclk));
	jdff dff_B_jx9QqAFk1_0(.din(w_dff_B_EzdcUTXM9_0),.dout(w_dff_B_jx9QqAFk1_0),.clk(gclk));
	jdff dff_B_pYIFf5wj1_0(.din(w_dff_B_jx9QqAFk1_0),.dout(w_dff_B_pYIFf5wj1_0),.clk(gclk));
	jdff dff_B_C8hsQ1t99_0(.din(w_dff_B_pYIFf5wj1_0),.dout(w_dff_B_C8hsQ1t99_0),.clk(gclk));
	jdff dff_B_um4WyG5E7_0(.din(w_dff_B_C8hsQ1t99_0),.dout(w_dff_B_um4WyG5E7_0),.clk(gclk));
	jdff dff_B_Mh8g19Sk5_0(.din(w_dff_B_um4WyG5E7_0),.dout(w_dff_B_Mh8g19Sk5_0),.clk(gclk));
	jdff dff_B_eh7BWXtk3_0(.din(w_dff_B_Mh8g19Sk5_0),.dout(w_dff_B_eh7BWXtk3_0),.clk(gclk));
	jdff dff_B_RRKtcs4q6_0(.din(w_dff_B_eh7BWXtk3_0),.dout(w_dff_B_RRKtcs4q6_0),.clk(gclk));
	jdff dff_B_MueYSLX36_0(.din(w_dff_B_RRKtcs4q6_0),.dout(w_dff_B_MueYSLX36_0),.clk(gclk));
	jdff dff_B_wooc5c0P3_0(.din(w_dff_B_MueYSLX36_0),.dout(w_dff_B_wooc5c0P3_0),.clk(gclk));
	jdff dff_B_ziaGA0rp2_0(.din(w_dff_B_wooc5c0P3_0),.dout(w_dff_B_ziaGA0rp2_0),.clk(gclk));
	jdff dff_B_WXptrmNp1_0(.din(w_dff_B_ziaGA0rp2_0),.dout(w_dff_B_WXptrmNp1_0),.clk(gclk));
	jdff dff_B_3zbQGrC62_0(.din(w_dff_B_WXptrmNp1_0),.dout(w_dff_B_3zbQGrC62_0),.clk(gclk));
	jdff dff_B_y6XPv0xv4_0(.din(w_dff_B_3zbQGrC62_0),.dout(w_dff_B_y6XPv0xv4_0),.clk(gclk));
	jdff dff_B_ci8m6xmH5_0(.din(w_dff_B_y6XPv0xv4_0),.dout(w_dff_B_ci8m6xmH5_0),.clk(gclk));
	jdff dff_B_DbwP4hdC4_0(.din(w_dff_B_ci8m6xmH5_0),.dout(w_dff_B_DbwP4hdC4_0),.clk(gclk));
	jdff dff_B_XE6q6rOO0_0(.din(w_dff_B_DbwP4hdC4_0),.dout(w_dff_B_XE6q6rOO0_0),.clk(gclk));
	jdff dff_B_5DMJKqlB4_0(.din(w_dff_B_XE6q6rOO0_0),.dout(w_dff_B_5DMJKqlB4_0),.clk(gclk));
	jdff dff_B_eCn7Nu3a1_0(.din(w_dff_B_5DMJKqlB4_0),.dout(w_dff_B_eCn7Nu3a1_0),.clk(gclk));
	jdff dff_B_JolXBKwI8_0(.din(w_dff_B_eCn7Nu3a1_0),.dout(w_dff_B_JolXBKwI8_0),.clk(gclk));
	jdff dff_B_Bq8QRUuD3_0(.din(w_dff_B_JolXBKwI8_0),.dout(w_dff_B_Bq8QRUuD3_0),.clk(gclk));
	jdff dff_B_ck9hUul88_0(.din(w_dff_B_Bq8QRUuD3_0),.dout(w_dff_B_ck9hUul88_0),.clk(gclk));
	jdff dff_B_WIJZ78gw8_0(.din(w_dff_B_ck9hUul88_0),.dout(w_dff_B_WIJZ78gw8_0),.clk(gclk));
	jdff dff_B_oZAz2n0E1_0(.din(w_dff_B_WIJZ78gw8_0),.dout(w_dff_B_oZAz2n0E1_0),.clk(gclk));
	jdff dff_B_3xVA9W6i1_0(.din(w_dff_B_oZAz2n0E1_0),.dout(w_dff_B_3xVA9W6i1_0),.clk(gclk));
	jdff dff_B_XQPE7p0h1_0(.din(w_dff_B_3xVA9W6i1_0),.dout(w_dff_B_XQPE7p0h1_0),.clk(gclk));
	jdff dff_B_cd2KeBby1_0(.din(w_dff_B_XQPE7p0h1_0),.dout(w_dff_B_cd2KeBby1_0),.clk(gclk));
	jdff dff_B_1uRJoPpO1_0(.din(w_dff_B_cd2KeBby1_0),.dout(w_dff_B_1uRJoPpO1_0),.clk(gclk));
	jdff dff_B_jTqEqb1H4_0(.din(w_dff_B_1uRJoPpO1_0),.dout(w_dff_B_jTqEqb1H4_0),.clk(gclk));
	jdff dff_B_hbt8k0ef1_0(.din(w_dff_B_jTqEqb1H4_0),.dout(w_dff_B_hbt8k0ef1_0),.clk(gclk));
	jdff dff_B_MYelRpm85_0(.din(w_dff_B_hbt8k0ef1_0),.dout(w_dff_B_MYelRpm85_0),.clk(gclk));
	jdff dff_B_pTlWKZ6x2_0(.din(w_dff_B_MYelRpm85_0),.dout(w_dff_B_pTlWKZ6x2_0),.clk(gclk));
	jdff dff_B_d8VofKpQ0_0(.din(w_dff_B_pTlWKZ6x2_0),.dout(w_dff_B_d8VofKpQ0_0),.clk(gclk));
	jdff dff_B_wbZG7QoE8_0(.din(w_dff_B_d8VofKpQ0_0),.dout(w_dff_B_wbZG7QoE8_0),.clk(gclk));
	jdff dff_B_phoMujdh2_0(.din(w_dff_B_wbZG7QoE8_0),.dout(w_dff_B_phoMujdh2_0),.clk(gclk));
	jdff dff_B_jVs3W3jJ7_0(.din(w_dff_B_phoMujdh2_0),.dout(w_dff_B_jVs3W3jJ7_0),.clk(gclk));
	jdff dff_B_qI0VCpAH7_0(.din(w_dff_B_jVs3W3jJ7_0),.dout(w_dff_B_qI0VCpAH7_0),.clk(gclk));
	jdff dff_B_GWSHrsgV9_0(.din(w_dff_B_qI0VCpAH7_0),.dout(w_dff_B_GWSHrsgV9_0),.clk(gclk));
	jdff dff_B_Qg6BnTtV9_0(.din(w_dff_B_GWSHrsgV9_0),.dout(w_dff_B_Qg6BnTtV9_0),.clk(gclk));
	jdff dff_B_6hzz9GG38_0(.din(w_dff_B_Qg6BnTtV9_0),.dout(w_dff_B_6hzz9GG38_0),.clk(gclk));
	jdff dff_B_sbZw3v7L2_0(.din(w_dff_B_6hzz9GG38_0),.dout(w_dff_B_sbZw3v7L2_0),.clk(gclk));
	jdff dff_B_BjYlc2CB4_0(.din(w_dff_B_sbZw3v7L2_0),.dout(w_dff_B_BjYlc2CB4_0),.clk(gclk));
	jdff dff_B_LXw0OWrp3_0(.din(w_dff_B_BjYlc2CB4_0),.dout(w_dff_B_LXw0OWrp3_0),.clk(gclk));
	jdff dff_B_UDcq6OOm5_0(.din(w_dff_B_LXw0OWrp3_0),.dout(w_dff_B_UDcq6OOm5_0),.clk(gclk));
	jdff dff_B_WuYhmjkv6_0(.din(w_dff_B_UDcq6OOm5_0),.dout(w_dff_B_WuYhmjkv6_0),.clk(gclk));
	jdff dff_B_oHjSdhyP1_0(.din(w_dff_B_WuYhmjkv6_0),.dout(w_dff_B_oHjSdhyP1_0),.clk(gclk));
	jdff dff_B_DvEsZjMl7_0(.din(w_dff_B_oHjSdhyP1_0),.dout(w_dff_B_DvEsZjMl7_0),.clk(gclk));
	jdff dff_B_AgOf2Dca6_0(.din(w_dff_B_DvEsZjMl7_0),.dout(w_dff_B_AgOf2Dca6_0),.clk(gclk));
	jdff dff_B_kaMqvGnX4_0(.din(w_dff_B_AgOf2Dca6_0),.dout(w_dff_B_kaMqvGnX4_0),.clk(gclk));
	jdff dff_B_LMcbZJOa8_0(.din(w_dff_B_kaMqvGnX4_0),.dout(w_dff_B_LMcbZJOa8_0),.clk(gclk));
	jdff dff_B_D4G1r1cU8_0(.din(w_dff_B_LMcbZJOa8_0),.dout(w_dff_B_D4G1r1cU8_0),.clk(gclk));
	jdff dff_B_6vOmPyiY1_0(.din(w_dff_B_D4G1r1cU8_0),.dout(w_dff_B_6vOmPyiY1_0),.clk(gclk));
	jdff dff_B_aeNsupF99_0(.din(w_dff_B_6vOmPyiY1_0),.dout(w_dff_B_aeNsupF99_0),.clk(gclk));
	jdff dff_B_T4j0H2KR2_0(.din(w_dff_B_aeNsupF99_0),.dout(w_dff_B_T4j0H2KR2_0),.clk(gclk));
	jdff dff_B_fphVRBL66_0(.din(w_dff_B_T4j0H2KR2_0),.dout(w_dff_B_fphVRBL66_0),.clk(gclk));
	jdff dff_B_2c6vUZbK5_0(.din(w_dff_B_fphVRBL66_0),.dout(w_dff_B_2c6vUZbK5_0),.clk(gclk));
	jdff dff_B_ZEmVIxwi4_0(.din(w_dff_B_2c6vUZbK5_0),.dout(w_dff_B_ZEmVIxwi4_0),.clk(gclk));
	jdff dff_B_HnKcbF1T8_0(.din(w_dff_B_ZEmVIxwi4_0),.dout(w_dff_B_HnKcbF1T8_0),.clk(gclk));
	jdff dff_B_9wjeYoBY6_0(.din(w_dff_B_HnKcbF1T8_0),.dout(w_dff_B_9wjeYoBY6_0),.clk(gclk));
	jdff dff_B_nWqcM3FS5_0(.din(w_dff_B_9wjeYoBY6_0),.dout(w_dff_B_nWqcM3FS5_0),.clk(gclk));
	jdff dff_B_7QFPOCrV6_0(.din(w_dff_B_nWqcM3FS5_0),.dout(w_dff_B_7QFPOCrV6_0),.clk(gclk));
	jdff dff_B_TgiI1lZR5_0(.din(w_dff_B_7QFPOCrV6_0),.dout(w_dff_B_TgiI1lZR5_0),.clk(gclk));
	jdff dff_B_ClKSzvHU7_0(.din(w_dff_B_TgiI1lZR5_0),.dout(w_dff_B_ClKSzvHU7_0),.clk(gclk));
	jdff dff_B_IfW2Sv7q7_0(.din(w_dff_B_ClKSzvHU7_0),.dout(w_dff_B_IfW2Sv7q7_0),.clk(gclk));
	jdff dff_B_NeD4Nn9y8_0(.din(w_dff_B_IfW2Sv7q7_0),.dout(w_dff_B_NeD4Nn9y8_0),.clk(gclk));
	jdff dff_B_UPVdnHXy5_0(.din(w_dff_B_NeD4Nn9y8_0),.dout(w_dff_B_UPVdnHXy5_0),.clk(gclk));
	jdff dff_B_6zU42Z0I9_0(.din(w_dff_B_UPVdnHXy5_0),.dout(w_dff_B_6zU42Z0I9_0),.clk(gclk));
	jdff dff_B_cAeYRSUq6_0(.din(w_dff_B_6zU42Z0I9_0),.dout(w_dff_B_cAeYRSUq6_0),.clk(gclk));
	jdff dff_B_rkqSrGhN4_0(.din(w_dff_B_cAeYRSUq6_0),.dout(w_dff_B_rkqSrGhN4_0),.clk(gclk));
	jdff dff_B_uw8WfP724_0(.din(w_dff_B_rkqSrGhN4_0),.dout(w_dff_B_uw8WfP724_0),.clk(gclk));
	jdff dff_B_SkhbmHSz9_0(.din(w_dff_B_uw8WfP724_0),.dout(w_dff_B_SkhbmHSz9_0),.clk(gclk));
	jdff dff_B_9rgiGrKw2_0(.din(w_dff_B_SkhbmHSz9_0),.dout(w_dff_B_9rgiGrKw2_0),.clk(gclk));
	jdff dff_B_DyeB2vL03_0(.din(w_dff_B_9rgiGrKw2_0),.dout(w_dff_B_DyeB2vL03_0),.clk(gclk));
	jdff dff_B_mcwkPAkL2_0(.din(w_dff_B_DyeB2vL03_0),.dout(w_dff_B_mcwkPAkL2_0),.clk(gclk));
	jdff dff_B_XuY9E4Ou4_0(.din(w_dff_B_mcwkPAkL2_0),.dout(w_dff_B_XuY9E4Ou4_0),.clk(gclk));
	jdff dff_B_BppOGXt43_0(.din(w_dff_B_XuY9E4Ou4_0),.dout(w_dff_B_BppOGXt43_0),.clk(gclk));
	jdff dff_B_pZ6P6bM07_0(.din(w_dff_B_BppOGXt43_0),.dout(w_dff_B_pZ6P6bM07_0),.clk(gclk));
	jdff dff_B_uuKE7prV9_0(.din(w_dff_B_pZ6P6bM07_0),.dout(w_dff_B_uuKE7prV9_0),.clk(gclk));
	jdff dff_B_YFkhXDhi0_0(.din(w_dff_B_uuKE7prV9_0),.dout(w_dff_B_YFkhXDhi0_0),.clk(gclk));
	jdff dff_B_ofaTlYyf5_0(.din(w_dff_B_YFkhXDhi0_0),.dout(w_dff_B_ofaTlYyf5_0),.clk(gclk));
	jdff dff_B_l1BQO1Bu9_0(.din(w_dff_B_ofaTlYyf5_0),.dout(w_dff_B_l1BQO1Bu9_0),.clk(gclk));
	jdff dff_B_87RqLrR94_0(.din(w_dff_B_l1BQO1Bu9_0),.dout(w_dff_B_87RqLrR94_0),.clk(gclk));
	jdff dff_B_BohxU8tM5_0(.din(w_dff_B_87RqLrR94_0),.dout(w_dff_B_BohxU8tM5_0),.clk(gclk));
	jdff dff_B_FT6qOtrS4_0(.din(w_dff_B_BohxU8tM5_0),.dout(w_dff_B_FT6qOtrS4_0),.clk(gclk));
	jdff dff_B_EuTOQkN66_0(.din(w_dff_B_FT6qOtrS4_0),.dout(w_dff_B_EuTOQkN66_0),.clk(gclk));
	jdff dff_B_Kr4Saxpw5_0(.din(w_dff_B_EuTOQkN66_0),.dout(w_dff_B_Kr4Saxpw5_0),.clk(gclk));
	jdff dff_B_aN2YQPxw9_0(.din(w_dff_B_Kr4Saxpw5_0),.dout(w_dff_B_aN2YQPxw9_0),.clk(gclk));
	jdff dff_B_lvOHKtlw4_0(.din(w_dff_B_aN2YQPxw9_0),.dout(w_dff_B_lvOHKtlw4_0),.clk(gclk));
	jdff dff_B_Bh5TkV9c9_0(.din(w_dff_B_lvOHKtlw4_0),.dout(w_dff_B_Bh5TkV9c9_0),.clk(gclk));
	jdff dff_B_yBY6zIKE7_0(.din(w_dff_B_Bh5TkV9c9_0),.dout(w_dff_B_yBY6zIKE7_0),.clk(gclk));
	jdff dff_B_OktgxKr12_0(.din(w_dff_B_yBY6zIKE7_0),.dout(w_dff_B_OktgxKr12_0),.clk(gclk));
	jdff dff_B_jXu0gceh6_0(.din(w_dff_B_OktgxKr12_0),.dout(w_dff_B_jXu0gceh6_0),.clk(gclk));
	jdff dff_B_RdfHookR8_0(.din(w_dff_B_jXu0gceh6_0),.dout(w_dff_B_RdfHookR8_0),.clk(gclk));
	jdff dff_B_H0luIVyz1_0(.din(w_dff_B_RdfHookR8_0),.dout(w_dff_B_H0luIVyz1_0),.clk(gclk));
	jdff dff_B_zzFl00kT8_0(.din(w_dff_B_H0luIVyz1_0),.dout(w_dff_B_zzFl00kT8_0),.clk(gclk));
	jdff dff_B_Mpjw50Ap0_0(.din(w_dff_B_zzFl00kT8_0),.dout(w_dff_B_Mpjw50Ap0_0),.clk(gclk));
	jdff dff_B_IY2l35Pl2_0(.din(w_dff_B_Mpjw50Ap0_0),.dout(w_dff_B_IY2l35Pl2_0),.clk(gclk));
	jdff dff_B_WO4CwQt12_0(.din(w_dff_B_IY2l35Pl2_0),.dout(w_dff_B_WO4CwQt12_0),.clk(gclk));
	jdff dff_B_vTtcFnaX1_0(.din(w_dff_B_WO4CwQt12_0),.dout(w_dff_B_vTtcFnaX1_0),.clk(gclk));
	jdff dff_B_Ov5Jfpqt1_0(.din(w_dff_B_vTtcFnaX1_0),.dout(w_dff_B_Ov5Jfpqt1_0),.clk(gclk));
	jdff dff_B_9CkXA9AG3_0(.din(w_dff_B_Ov5Jfpqt1_0),.dout(w_dff_B_9CkXA9AG3_0),.clk(gclk));
	jdff dff_B_gVkbTBwR4_0(.din(w_dff_B_9CkXA9AG3_0),.dout(w_dff_B_gVkbTBwR4_0),.clk(gclk));
	jdff dff_B_vlndYaxx5_0(.din(w_dff_B_gVkbTBwR4_0),.dout(w_dff_B_vlndYaxx5_0),.clk(gclk));
	jdff dff_B_r3RtS4sf5_0(.din(w_dff_B_vlndYaxx5_0),.dout(w_dff_B_r3RtS4sf5_0),.clk(gclk));
	jdff dff_B_20S2Q5oJ1_0(.din(w_dff_B_r3RtS4sf5_0),.dout(w_dff_B_20S2Q5oJ1_0),.clk(gclk));
	jdff dff_B_ZaARAyP08_0(.din(w_dff_B_20S2Q5oJ1_0),.dout(w_dff_B_ZaARAyP08_0),.clk(gclk));
	jdff dff_B_aG5BVySM7_0(.din(w_dff_B_ZaARAyP08_0),.dout(w_dff_B_aG5BVySM7_0),.clk(gclk));
	jdff dff_B_vqfDjWX14_0(.din(w_dff_B_aG5BVySM7_0),.dout(w_dff_B_vqfDjWX14_0),.clk(gclk));
	jdff dff_B_lx4KyX9J6_0(.din(w_dff_B_vqfDjWX14_0),.dout(w_dff_B_lx4KyX9J6_0),.clk(gclk));
	jdff dff_B_G6kldeH14_0(.din(w_dff_B_lx4KyX9J6_0),.dout(w_dff_B_G6kldeH14_0),.clk(gclk));
	jdff dff_B_v8aBzas02_0(.din(w_dff_B_G6kldeH14_0),.dout(w_dff_B_v8aBzas02_0),.clk(gclk));
	jdff dff_B_uVItd6s24_0(.din(w_dff_B_v8aBzas02_0),.dout(w_dff_B_uVItd6s24_0),.clk(gclk));
	jdff dff_B_ZLMwJtYI1_0(.din(w_dff_B_uVItd6s24_0),.dout(w_dff_B_ZLMwJtYI1_0),.clk(gclk));
	jdff dff_B_1FVKKcoT6_0(.din(w_dff_B_ZLMwJtYI1_0),.dout(w_dff_B_1FVKKcoT6_0),.clk(gclk));
	jdff dff_B_SRgO1VNq5_0(.din(w_dff_B_1FVKKcoT6_0),.dout(w_dff_B_SRgO1VNq5_0),.clk(gclk));
	jdff dff_B_TSH1xZyN5_0(.din(w_dff_B_SRgO1VNq5_0),.dout(w_dff_B_TSH1xZyN5_0),.clk(gclk));
	jdff dff_B_Vt8WOKXG1_0(.din(w_dff_B_TSH1xZyN5_0),.dout(w_dff_B_Vt8WOKXG1_0),.clk(gclk));
	jdff dff_B_xOmJmBh08_0(.din(w_dff_B_Vt8WOKXG1_0),.dout(w_dff_B_xOmJmBh08_0),.clk(gclk));
	jdff dff_B_yMpw4ghJ6_0(.din(w_dff_B_xOmJmBh08_0),.dout(w_dff_B_yMpw4ghJ6_0),.clk(gclk));
	jdff dff_B_E0UEn0QU0_0(.din(w_dff_B_yMpw4ghJ6_0),.dout(w_dff_B_E0UEn0QU0_0),.clk(gclk));
	jdff dff_B_lIfmeSyV2_0(.din(w_dff_B_E0UEn0QU0_0),.dout(w_dff_B_lIfmeSyV2_0),.clk(gclk));
	jdff dff_B_hcdQaGWh9_0(.din(w_dff_B_lIfmeSyV2_0),.dout(w_dff_B_hcdQaGWh9_0),.clk(gclk));
	jdff dff_B_GZvz9KB76_0(.din(w_dff_B_hcdQaGWh9_0),.dout(w_dff_B_GZvz9KB76_0),.clk(gclk));
	jdff dff_B_Q2Hc1GQB1_0(.din(w_dff_B_GZvz9KB76_0),.dout(w_dff_B_Q2Hc1GQB1_0),.clk(gclk));
	jdff dff_B_8Dm77OtX9_0(.din(w_dff_B_Q2Hc1GQB1_0),.dout(w_dff_B_8Dm77OtX9_0),.clk(gclk));
	jdff dff_B_atmx5RPm8_1(.din(n1146),.dout(w_dff_B_atmx5RPm8_1),.clk(gclk));
	jdff dff_B_RFADscL76_1(.din(w_dff_B_atmx5RPm8_1),.dout(w_dff_B_RFADscL76_1),.clk(gclk));
	jdff dff_B_rj31xIls3_1(.din(w_dff_B_RFADscL76_1),.dout(w_dff_B_rj31xIls3_1),.clk(gclk));
	jdff dff_B_9RGDo8fL4_1(.din(w_dff_B_rj31xIls3_1),.dout(w_dff_B_9RGDo8fL4_1),.clk(gclk));
	jdff dff_B_oeDww5zt9_1(.din(w_dff_B_9RGDo8fL4_1),.dout(w_dff_B_oeDww5zt9_1),.clk(gclk));
	jdff dff_B_RPTgCTBP0_1(.din(w_dff_B_oeDww5zt9_1),.dout(w_dff_B_RPTgCTBP0_1),.clk(gclk));
	jdff dff_B_x6gtpROe7_1(.din(w_dff_B_RPTgCTBP0_1),.dout(w_dff_B_x6gtpROe7_1),.clk(gclk));
	jdff dff_B_4EzZvJGs4_1(.din(w_dff_B_x6gtpROe7_1),.dout(w_dff_B_4EzZvJGs4_1),.clk(gclk));
	jdff dff_B_AmluzxDU4_1(.din(w_dff_B_4EzZvJGs4_1),.dout(w_dff_B_AmluzxDU4_1),.clk(gclk));
	jdff dff_B_tv8mwf8P2_1(.din(w_dff_B_AmluzxDU4_1),.dout(w_dff_B_tv8mwf8P2_1),.clk(gclk));
	jdff dff_B_igS4eQLx5_1(.din(w_dff_B_tv8mwf8P2_1),.dout(w_dff_B_igS4eQLx5_1),.clk(gclk));
	jdff dff_B_U48KMSgO0_1(.din(w_dff_B_igS4eQLx5_1),.dout(w_dff_B_U48KMSgO0_1),.clk(gclk));
	jdff dff_B_NczshOmV4_1(.din(w_dff_B_U48KMSgO0_1),.dout(w_dff_B_NczshOmV4_1),.clk(gclk));
	jdff dff_B_THkn9HEh5_1(.din(w_dff_B_NczshOmV4_1),.dout(w_dff_B_THkn9HEh5_1),.clk(gclk));
	jdff dff_B_9wMpNnnR9_1(.din(w_dff_B_THkn9HEh5_1),.dout(w_dff_B_9wMpNnnR9_1),.clk(gclk));
	jdff dff_B_79Q61mpM9_1(.din(w_dff_B_9wMpNnnR9_1),.dout(w_dff_B_79Q61mpM9_1),.clk(gclk));
	jdff dff_B_9PuQADfm2_1(.din(w_dff_B_79Q61mpM9_1),.dout(w_dff_B_9PuQADfm2_1),.clk(gclk));
	jdff dff_B_okaXoeu12_1(.din(w_dff_B_9PuQADfm2_1),.dout(w_dff_B_okaXoeu12_1),.clk(gclk));
	jdff dff_B_JFAqEzkK9_1(.din(w_dff_B_okaXoeu12_1),.dout(w_dff_B_JFAqEzkK9_1),.clk(gclk));
	jdff dff_B_Z5PLn4Da1_1(.din(w_dff_B_JFAqEzkK9_1),.dout(w_dff_B_Z5PLn4Da1_1),.clk(gclk));
	jdff dff_B_6CiEtYja6_1(.din(w_dff_B_Z5PLn4Da1_1),.dout(w_dff_B_6CiEtYja6_1),.clk(gclk));
	jdff dff_B_2vwo12f40_1(.din(w_dff_B_6CiEtYja6_1),.dout(w_dff_B_2vwo12f40_1),.clk(gclk));
	jdff dff_B_rqpUrkEP4_1(.din(w_dff_B_2vwo12f40_1),.dout(w_dff_B_rqpUrkEP4_1),.clk(gclk));
	jdff dff_B_zt1VhDA51_1(.din(w_dff_B_rqpUrkEP4_1),.dout(w_dff_B_zt1VhDA51_1),.clk(gclk));
	jdff dff_B_bd1VUPjf7_1(.din(w_dff_B_zt1VhDA51_1),.dout(w_dff_B_bd1VUPjf7_1),.clk(gclk));
	jdff dff_B_HGpO0FUN8_1(.din(w_dff_B_bd1VUPjf7_1),.dout(w_dff_B_HGpO0FUN8_1),.clk(gclk));
	jdff dff_B_GsGj0xnB0_1(.din(w_dff_B_HGpO0FUN8_1),.dout(w_dff_B_GsGj0xnB0_1),.clk(gclk));
	jdff dff_B_WBxiJ5p85_1(.din(w_dff_B_GsGj0xnB0_1),.dout(w_dff_B_WBxiJ5p85_1),.clk(gclk));
	jdff dff_B_M7puSxrt0_1(.din(w_dff_B_WBxiJ5p85_1),.dout(w_dff_B_M7puSxrt0_1),.clk(gclk));
	jdff dff_B_5OJSG2Qz4_1(.din(w_dff_B_M7puSxrt0_1),.dout(w_dff_B_5OJSG2Qz4_1),.clk(gclk));
	jdff dff_B_JJKXNAmW8_1(.din(w_dff_B_5OJSG2Qz4_1),.dout(w_dff_B_JJKXNAmW8_1),.clk(gclk));
	jdff dff_B_XLWcYd4j3_1(.din(w_dff_B_JJKXNAmW8_1),.dout(w_dff_B_XLWcYd4j3_1),.clk(gclk));
	jdff dff_B_72ROqm773_1(.din(w_dff_B_XLWcYd4j3_1),.dout(w_dff_B_72ROqm773_1),.clk(gclk));
	jdff dff_B_p25PetQz4_1(.din(w_dff_B_72ROqm773_1),.dout(w_dff_B_p25PetQz4_1),.clk(gclk));
	jdff dff_B_67EOdVvO7_1(.din(w_dff_B_p25PetQz4_1),.dout(w_dff_B_67EOdVvO7_1),.clk(gclk));
	jdff dff_B_AYhQO0aq8_1(.din(w_dff_B_67EOdVvO7_1),.dout(w_dff_B_AYhQO0aq8_1),.clk(gclk));
	jdff dff_B_76oJad779_1(.din(w_dff_B_AYhQO0aq8_1),.dout(w_dff_B_76oJad779_1),.clk(gclk));
	jdff dff_B_rP15x5Rj0_1(.din(w_dff_B_76oJad779_1),.dout(w_dff_B_rP15x5Rj0_1),.clk(gclk));
	jdff dff_B_up7mT3Jm8_1(.din(w_dff_B_rP15x5Rj0_1),.dout(w_dff_B_up7mT3Jm8_1),.clk(gclk));
	jdff dff_B_KFzFLXDC0_1(.din(w_dff_B_up7mT3Jm8_1),.dout(w_dff_B_KFzFLXDC0_1),.clk(gclk));
	jdff dff_B_VY05avO17_1(.din(w_dff_B_KFzFLXDC0_1),.dout(w_dff_B_VY05avO17_1),.clk(gclk));
	jdff dff_B_S5uGMGjZ9_1(.din(w_dff_B_VY05avO17_1),.dout(w_dff_B_S5uGMGjZ9_1),.clk(gclk));
	jdff dff_B_jCQhqh0Q3_1(.din(w_dff_B_S5uGMGjZ9_1),.dout(w_dff_B_jCQhqh0Q3_1),.clk(gclk));
	jdff dff_B_w0dy3pmO6_1(.din(w_dff_B_jCQhqh0Q3_1),.dout(w_dff_B_w0dy3pmO6_1),.clk(gclk));
	jdff dff_B_T6It8k2d6_1(.din(w_dff_B_w0dy3pmO6_1),.dout(w_dff_B_T6It8k2d6_1),.clk(gclk));
	jdff dff_B_rtoXt2Is2_1(.din(w_dff_B_T6It8k2d6_1),.dout(w_dff_B_rtoXt2Is2_1),.clk(gclk));
	jdff dff_B_g2MJLP8o2_1(.din(w_dff_B_rtoXt2Is2_1),.dout(w_dff_B_g2MJLP8o2_1),.clk(gclk));
	jdff dff_B_whyfvX1e7_1(.din(w_dff_B_g2MJLP8o2_1),.dout(w_dff_B_whyfvX1e7_1),.clk(gclk));
	jdff dff_B_HZYjyU0U5_1(.din(w_dff_B_whyfvX1e7_1),.dout(w_dff_B_HZYjyU0U5_1),.clk(gclk));
	jdff dff_B_oQqu21dV9_1(.din(w_dff_B_HZYjyU0U5_1),.dout(w_dff_B_oQqu21dV9_1),.clk(gclk));
	jdff dff_B_DRUxcFe53_1(.din(w_dff_B_oQqu21dV9_1),.dout(w_dff_B_DRUxcFe53_1),.clk(gclk));
	jdff dff_B_WzSQX1Jb5_1(.din(w_dff_B_DRUxcFe53_1),.dout(w_dff_B_WzSQX1Jb5_1),.clk(gclk));
	jdff dff_B_v9ivZ9ad6_1(.din(w_dff_B_WzSQX1Jb5_1),.dout(w_dff_B_v9ivZ9ad6_1),.clk(gclk));
	jdff dff_B_gYpFQRhC0_1(.din(w_dff_B_v9ivZ9ad6_1),.dout(w_dff_B_gYpFQRhC0_1),.clk(gclk));
	jdff dff_B_6w1SuZ9p1_1(.din(w_dff_B_gYpFQRhC0_1),.dout(w_dff_B_6w1SuZ9p1_1),.clk(gclk));
	jdff dff_B_3p7OZ9v27_1(.din(w_dff_B_6w1SuZ9p1_1),.dout(w_dff_B_3p7OZ9v27_1),.clk(gclk));
	jdff dff_B_dMb07bMO2_1(.din(w_dff_B_3p7OZ9v27_1),.dout(w_dff_B_dMb07bMO2_1),.clk(gclk));
	jdff dff_B_pItQfPMm5_1(.din(w_dff_B_dMb07bMO2_1),.dout(w_dff_B_pItQfPMm5_1),.clk(gclk));
	jdff dff_B_HX5bYkUY3_1(.din(w_dff_B_pItQfPMm5_1),.dout(w_dff_B_HX5bYkUY3_1),.clk(gclk));
	jdff dff_B_1FMtGHUR4_1(.din(w_dff_B_HX5bYkUY3_1),.dout(w_dff_B_1FMtGHUR4_1),.clk(gclk));
	jdff dff_B_cYrW1LaP2_1(.din(w_dff_B_1FMtGHUR4_1),.dout(w_dff_B_cYrW1LaP2_1),.clk(gclk));
	jdff dff_B_XzpDLXSC2_1(.din(w_dff_B_cYrW1LaP2_1),.dout(w_dff_B_XzpDLXSC2_1),.clk(gclk));
	jdff dff_B_LfM2WKy50_1(.din(w_dff_B_XzpDLXSC2_1),.dout(w_dff_B_LfM2WKy50_1),.clk(gclk));
	jdff dff_B_V5Hlthry0_1(.din(w_dff_B_LfM2WKy50_1),.dout(w_dff_B_V5Hlthry0_1),.clk(gclk));
	jdff dff_B_Y42FY6WM1_1(.din(w_dff_B_V5Hlthry0_1),.dout(w_dff_B_Y42FY6WM1_1),.clk(gclk));
	jdff dff_B_4gytCVG11_1(.din(w_dff_B_Y42FY6WM1_1),.dout(w_dff_B_4gytCVG11_1),.clk(gclk));
	jdff dff_B_G4aqjBaa6_1(.din(w_dff_B_4gytCVG11_1),.dout(w_dff_B_G4aqjBaa6_1),.clk(gclk));
	jdff dff_B_Wnrjcml20_1(.din(w_dff_B_G4aqjBaa6_1),.dout(w_dff_B_Wnrjcml20_1),.clk(gclk));
	jdff dff_B_94XqCZLk3_1(.din(w_dff_B_Wnrjcml20_1),.dout(w_dff_B_94XqCZLk3_1),.clk(gclk));
	jdff dff_B_PfKSA2qF1_1(.din(w_dff_B_94XqCZLk3_1),.dout(w_dff_B_PfKSA2qF1_1),.clk(gclk));
	jdff dff_B_KgBkMctq7_1(.din(w_dff_B_PfKSA2qF1_1),.dout(w_dff_B_KgBkMctq7_1),.clk(gclk));
	jdff dff_B_OjoujAV64_1(.din(w_dff_B_KgBkMctq7_1),.dout(w_dff_B_OjoujAV64_1),.clk(gclk));
	jdff dff_B_HynhC1Us7_1(.din(w_dff_B_OjoujAV64_1),.dout(w_dff_B_HynhC1Us7_1),.clk(gclk));
	jdff dff_B_NQC4b47e6_1(.din(w_dff_B_HynhC1Us7_1),.dout(w_dff_B_NQC4b47e6_1),.clk(gclk));
	jdff dff_B_1tKqnsoN1_1(.din(w_dff_B_NQC4b47e6_1),.dout(w_dff_B_1tKqnsoN1_1),.clk(gclk));
	jdff dff_B_uGDjLqrh9_1(.din(w_dff_B_1tKqnsoN1_1),.dout(w_dff_B_uGDjLqrh9_1),.clk(gclk));
	jdff dff_B_Vl6FtdEh6_1(.din(w_dff_B_uGDjLqrh9_1),.dout(w_dff_B_Vl6FtdEh6_1),.clk(gclk));
	jdff dff_B_C6bW0Lci0_1(.din(w_dff_B_Vl6FtdEh6_1),.dout(w_dff_B_C6bW0Lci0_1),.clk(gclk));
	jdff dff_B_ZkHqpgI72_1(.din(w_dff_B_C6bW0Lci0_1),.dout(w_dff_B_ZkHqpgI72_1),.clk(gclk));
	jdff dff_B_G8a6zfWg1_1(.din(w_dff_B_ZkHqpgI72_1),.dout(w_dff_B_G8a6zfWg1_1),.clk(gclk));
	jdff dff_B_4LuSDWLC6_1(.din(w_dff_B_G8a6zfWg1_1),.dout(w_dff_B_4LuSDWLC6_1),.clk(gclk));
	jdff dff_B_9mDyfVzL3_1(.din(w_dff_B_4LuSDWLC6_1),.dout(w_dff_B_9mDyfVzL3_1),.clk(gclk));
	jdff dff_B_YPSKTM3S9_1(.din(w_dff_B_9mDyfVzL3_1),.dout(w_dff_B_YPSKTM3S9_1),.clk(gclk));
	jdff dff_B_PRKFr2OB3_1(.din(w_dff_B_YPSKTM3S9_1),.dout(w_dff_B_PRKFr2OB3_1),.clk(gclk));
	jdff dff_B_3jV6T0em6_1(.din(w_dff_B_PRKFr2OB3_1),.dout(w_dff_B_3jV6T0em6_1),.clk(gclk));
	jdff dff_B_RFINkQKi6_1(.din(w_dff_B_3jV6T0em6_1),.dout(w_dff_B_RFINkQKi6_1),.clk(gclk));
	jdff dff_B_reVxmV880_1(.din(w_dff_B_RFINkQKi6_1),.dout(w_dff_B_reVxmV880_1),.clk(gclk));
	jdff dff_B_2zQ7FImu0_1(.din(w_dff_B_reVxmV880_1),.dout(w_dff_B_2zQ7FImu0_1),.clk(gclk));
	jdff dff_B_dh03SZt34_1(.din(w_dff_B_2zQ7FImu0_1),.dout(w_dff_B_dh03SZt34_1),.clk(gclk));
	jdff dff_B_ldiTaqoA7_1(.din(w_dff_B_dh03SZt34_1),.dout(w_dff_B_ldiTaqoA7_1),.clk(gclk));
	jdff dff_B_C5rcPgpM8_1(.din(w_dff_B_ldiTaqoA7_1),.dout(w_dff_B_C5rcPgpM8_1),.clk(gclk));
	jdff dff_B_QPQLq1Oy9_1(.din(w_dff_B_C5rcPgpM8_1),.dout(w_dff_B_QPQLq1Oy9_1),.clk(gclk));
	jdff dff_B_lvX0xXKI8_1(.din(w_dff_B_QPQLq1Oy9_1),.dout(w_dff_B_lvX0xXKI8_1),.clk(gclk));
	jdff dff_B_rgz1z64h0_1(.din(w_dff_B_lvX0xXKI8_1),.dout(w_dff_B_rgz1z64h0_1),.clk(gclk));
	jdff dff_B_PyqAeOa11_1(.din(w_dff_B_rgz1z64h0_1),.dout(w_dff_B_PyqAeOa11_1),.clk(gclk));
	jdff dff_B_wOfb5myz5_1(.din(w_dff_B_PyqAeOa11_1),.dout(w_dff_B_wOfb5myz5_1),.clk(gclk));
	jdff dff_B_xNcuImkN8_1(.din(w_dff_B_wOfb5myz5_1),.dout(w_dff_B_xNcuImkN8_1),.clk(gclk));
	jdff dff_B_t6eym27f6_1(.din(w_dff_B_xNcuImkN8_1),.dout(w_dff_B_t6eym27f6_1),.clk(gclk));
	jdff dff_B_53l1Clmq1_1(.din(w_dff_B_t6eym27f6_1),.dout(w_dff_B_53l1Clmq1_1),.clk(gclk));
	jdff dff_B_fCkwkyjV4_1(.din(w_dff_B_53l1Clmq1_1),.dout(w_dff_B_fCkwkyjV4_1),.clk(gclk));
	jdff dff_B_DJ7IG5Eh6_1(.din(w_dff_B_fCkwkyjV4_1),.dout(w_dff_B_DJ7IG5Eh6_1),.clk(gclk));
	jdff dff_B_l3OTR7B54_1(.din(w_dff_B_DJ7IG5Eh6_1),.dout(w_dff_B_l3OTR7B54_1),.clk(gclk));
	jdff dff_B_qMaKviYj5_1(.din(w_dff_B_l3OTR7B54_1),.dout(w_dff_B_qMaKviYj5_1),.clk(gclk));
	jdff dff_B_KaLZeSy47_1(.din(w_dff_B_qMaKviYj5_1),.dout(w_dff_B_KaLZeSy47_1),.clk(gclk));
	jdff dff_B_mv5YzRGw0_1(.din(w_dff_B_KaLZeSy47_1),.dout(w_dff_B_mv5YzRGw0_1),.clk(gclk));
	jdff dff_B_e5DQr9QO4_1(.din(w_dff_B_mv5YzRGw0_1),.dout(w_dff_B_e5DQr9QO4_1),.clk(gclk));
	jdff dff_B_n6QN3WIB6_1(.din(w_dff_B_e5DQr9QO4_1),.dout(w_dff_B_n6QN3WIB6_1),.clk(gclk));
	jdff dff_B_x0BLhzmH2_1(.din(w_dff_B_n6QN3WIB6_1),.dout(w_dff_B_x0BLhzmH2_1),.clk(gclk));
	jdff dff_B_QdGEdET97_1(.din(w_dff_B_x0BLhzmH2_1),.dout(w_dff_B_QdGEdET97_1),.clk(gclk));
	jdff dff_B_4mX8BWrB6_1(.din(w_dff_B_QdGEdET97_1),.dout(w_dff_B_4mX8BWrB6_1),.clk(gclk));
	jdff dff_B_UigGvA6R5_1(.din(w_dff_B_4mX8BWrB6_1),.dout(w_dff_B_UigGvA6R5_1),.clk(gclk));
	jdff dff_B_8QcYi2eM7_1(.din(w_dff_B_UigGvA6R5_1),.dout(w_dff_B_8QcYi2eM7_1),.clk(gclk));
	jdff dff_B_QJqq90ea5_1(.din(w_dff_B_8QcYi2eM7_1),.dout(w_dff_B_QJqq90ea5_1),.clk(gclk));
	jdff dff_B_9bOUD3e91_1(.din(w_dff_B_QJqq90ea5_1),.dout(w_dff_B_9bOUD3e91_1),.clk(gclk));
	jdff dff_B_LP806dpe2_1(.din(w_dff_B_9bOUD3e91_1),.dout(w_dff_B_LP806dpe2_1),.clk(gclk));
	jdff dff_B_FTExwWGv4_1(.din(w_dff_B_LP806dpe2_1),.dout(w_dff_B_FTExwWGv4_1),.clk(gclk));
	jdff dff_B_RCPZkv7G0_1(.din(w_dff_B_FTExwWGv4_1),.dout(w_dff_B_RCPZkv7G0_1),.clk(gclk));
	jdff dff_B_NaKG4y3Z2_1(.din(w_dff_B_RCPZkv7G0_1),.dout(w_dff_B_NaKG4y3Z2_1),.clk(gclk));
	jdff dff_B_HRz2cCEW6_1(.din(w_dff_B_NaKG4y3Z2_1),.dout(w_dff_B_HRz2cCEW6_1),.clk(gclk));
	jdff dff_B_WC60V9Pu8_1(.din(w_dff_B_HRz2cCEW6_1),.dout(w_dff_B_WC60V9Pu8_1),.clk(gclk));
	jdff dff_B_gzY9tO7N6_1(.din(w_dff_B_WC60V9Pu8_1),.dout(w_dff_B_gzY9tO7N6_1),.clk(gclk));
	jdff dff_B_6uRnwMLP0_1(.din(w_dff_B_gzY9tO7N6_1),.dout(w_dff_B_6uRnwMLP0_1),.clk(gclk));
	jdff dff_B_5QD35np92_1(.din(w_dff_B_6uRnwMLP0_1),.dout(w_dff_B_5QD35np92_1),.clk(gclk));
	jdff dff_B_d1nf5OLW0_1(.din(w_dff_B_5QD35np92_1),.dout(w_dff_B_d1nf5OLW0_1),.clk(gclk));
	jdff dff_B_cokVGotX5_1(.din(w_dff_B_d1nf5OLW0_1),.dout(w_dff_B_cokVGotX5_1),.clk(gclk));
	jdff dff_B_tpBuigwr1_1(.din(w_dff_B_cokVGotX5_1),.dout(w_dff_B_tpBuigwr1_1),.clk(gclk));
	jdff dff_B_66p7sXjF1_1(.din(w_dff_B_tpBuigwr1_1),.dout(w_dff_B_66p7sXjF1_1),.clk(gclk));
	jdff dff_B_ZhSybxxK6_0(.din(n1147),.dout(w_dff_B_ZhSybxxK6_0),.clk(gclk));
	jdff dff_B_HR6ojHVk8_0(.din(w_dff_B_ZhSybxxK6_0),.dout(w_dff_B_HR6ojHVk8_0),.clk(gclk));
	jdff dff_B_7v69VILJ0_0(.din(w_dff_B_HR6ojHVk8_0),.dout(w_dff_B_7v69VILJ0_0),.clk(gclk));
	jdff dff_B_pxZt5sZd2_0(.din(w_dff_B_7v69VILJ0_0),.dout(w_dff_B_pxZt5sZd2_0),.clk(gclk));
	jdff dff_B_CTEC44q93_0(.din(w_dff_B_pxZt5sZd2_0),.dout(w_dff_B_CTEC44q93_0),.clk(gclk));
	jdff dff_B_tUSTaSsl3_0(.din(w_dff_B_CTEC44q93_0),.dout(w_dff_B_tUSTaSsl3_0),.clk(gclk));
	jdff dff_B_T9b8DQA04_0(.din(w_dff_B_tUSTaSsl3_0),.dout(w_dff_B_T9b8DQA04_0),.clk(gclk));
	jdff dff_B_rGAOrHRK2_0(.din(w_dff_B_T9b8DQA04_0),.dout(w_dff_B_rGAOrHRK2_0),.clk(gclk));
	jdff dff_B_fCOsxztJ2_0(.din(w_dff_B_rGAOrHRK2_0),.dout(w_dff_B_fCOsxztJ2_0),.clk(gclk));
	jdff dff_B_r98hkcrQ3_0(.din(w_dff_B_fCOsxztJ2_0),.dout(w_dff_B_r98hkcrQ3_0),.clk(gclk));
	jdff dff_B_Ah5Lmctq4_0(.din(w_dff_B_r98hkcrQ3_0),.dout(w_dff_B_Ah5Lmctq4_0),.clk(gclk));
	jdff dff_B_JiODjbEz2_0(.din(w_dff_B_Ah5Lmctq4_0),.dout(w_dff_B_JiODjbEz2_0),.clk(gclk));
	jdff dff_B_U6Q9QYTM3_0(.din(w_dff_B_JiODjbEz2_0),.dout(w_dff_B_U6Q9QYTM3_0),.clk(gclk));
	jdff dff_B_ERbzeH3g0_0(.din(w_dff_B_U6Q9QYTM3_0),.dout(w_dff_B_ERbzeH3g0_0),.clk(gclk));
	jdff dff_B_ia2eZ6ML2_0(.din(w_dff_B_ERbzeH3g0_0),.dout(w_dff_B_ia2eZ6ML2_0),.clk(gclk));
	jdff dff_B_iVplwo8H9_0(.din(w_dff_B_ia2eZ6ML2_0),.dout(w_dff_B_iVplwo8H9_0),.clk(gclk));
	jdff dff_B_yUEcPzMJ8_0(.din(w_dff_B_iVplwo8H9_0),.dout(w_dff_B_yUEcPzMJ8_0),.clk(gclk));
	jdff dff_B_t1A2hG7x9_0(.din(w_dff_B_yUEcPzMJ8_0),.dout(w_dff_B_t1A2hG7x9_0),.clk(gclk));
	jdff dff_B_QdtDZF1S8_0(.din(w_dff_B_t1A2hG7x9_0),.dout(w_dff_B_QdtDZF1S8_0),.clk(gclk));
	jdff dff_B_EVcLzrgm9_0(.din(w_dff_B_QdtDZF1S8_0),.dout(w_dff_B_EVcLzrgm9_0),.clk(gclk));
	jdff dff_B_slC5Nc3n2_0(.din(w_dff_B_EVcLzrgm9_0),.dout(w_dff_B_slC5Nc3n2_0),.clk(gclk));
	jdff dff_B_XXcTucB50_0(.din(w_dff_B_slC5Nc3n2_0),.dout(w_dff_B_XXcTucB50_0),.clk(gclk));
	jdff dff_B_2D1X5yUO2_0(.din(w_dff_B_XXcTucB50_0),.dout(w_dff_B_2D1X5yUO2_0),.clk(gclk));
	jdff dff_B_K180yQkN7_0(.din(w_dff_B_2D1X5yUO2_0),.dout(w_dff_B_K180yQkN7_0),.clk(gclk));
	jdff dff_B_qWhpoLDA6_0(.din(w_dff_B_K180yQkN7_0),.dout(w_dff_B_qWhpoLDA6_0),.clk(gclk));
	jdff dff_B_aT2LDygW3_0(.din(w_dff_B_qWhpoLDA6_0),.dout(w_dff_B_aT2LDygW3_0),.clk(gclk));
	jdff dff_B_vXRpq0DC2_0(.din(w_dff_B_aT2LDygW3_0),.dout(w_dff_B_vXRpq0DC2_0),.clk(gclk));
	jdff dff_B_V1JEaggK4_0(.din(w_dff_B_vXRpq0DC2_0),.dout(w_dff_B_V1JEaggK4_0),.clk(gclk));
	jdff dff_B_izUq2Um46_0(.din(w_dff_B_V1JEaggK4_0),.dout(w_dff_B_izUq2Um46_0),.clk(gclk));
	jdff dff_B_I0K9myuV1_0(.din(w_dff_B_izUq2Um46_0),.dout(w_dff_B_I0K9myuV1_0),.clk(gclk));
	jdff dff_B_sTaUWHyB2_0(.din(w_dff_B_I0K9myuV1_0),.dout(w_dff_B_sTaUWHyB2_0),.clk(gclk));
	jdff dff_B_fGAkXdOh0_0(.din(w_dff_B_sTaUWHyB2_0),.dout(w_dff_B_fGAkXdOh0_0),.clk(gclk));
	jdff dff_B_XO1po3HH2_0(.din(w_dff_B_fGAkXdOh0_0),.dout(w_dff_B_XO1po3HH2_0),.clk(gclk));
	jdff dff_B_9tav4sVA3_0(.din(w_dff_B_XO1po3HH2_0),.dout(w_dff_B_9tav4sVA3_0),.clk(gclk));
	jdff dff_B_dFPmVX9Y9_0(.din(w_dff_B_9tav4sVA3_0),.dout(w_dff_B_dFPmVX9Y9_0),.clk(gclk));
	jdff dff_B_Wed9gell2_0(.din(w_dff_B_dFPmVX9Y9_0),.dout(w_dff_B_Wed9gell2_0),.clk(gclk));
	jdff dff_B_Vwnu2Rxe2_0(.din(w_dff_B_Wed9gell2_0),.dout(w_dff_B_Vwnu2Rxe2_0),.clk(gclk));
	jdff dff_B_C9l0aCj93_0(.din(w_dff_B_Vwnu2Rxe2_0),.dout(w_dff_B_C9l0aCj93_0),.clk(gclk));
	jdff dff_B_h369j09H8_0(.din(w_dff_B_C9l0aCj93_0),.dout(w_dff_B_h369j09H8_0),.clk(gclk));
	jdff dff_B_TAuZZkPz3_0(.din(w_dff_B_h369j09H8_0),.dout(w_dff_B_TAuZZkPz3_0),.clk(gclk));
	jdff dff_B_HlRPPLr95_0(.din(w_dff_B_TAuZZkPz3_0),.dout(w_dff_B_HlRPPLr95_0),.clk(gclk));
	jdff dff_B_QnUObPUF9_0(.din(w_dff_B_HlRPPLr95_0),.dout(w_dff_B_QnUObPUF9_0),.clk(gclk));
	jdff dff_B_Z1hgLreU2_0(.din(w_dff_B_QnUObPUF9_0),.dout(w_dff_B_Z1hgLreU2_0),.clk(gclk));
	jdff dff_B_qv50o4BA2_0(.din(w_dff_B_Z1hgLreU2_0),.dout(w_dff_B_qv50o4BA2_0),.clk(gclk));
	jdff dff_B_o0Xx4yWp2_0(.din(w_dff_B_qv50o4BA2_0),.dout(w_dff_B_o0Xx4yWp2_0),.clk(gclk));
	jdff dff_B_U0qfYNmh5_0(.din(w_dff_B_o0Xx4yWp2_0),.dout(w_dff_B_U0qfYNmh5_0),.clk(gclk));
	jdff dff_B_ChDSmj630_0(.din(w_dff_B_U0qfYNmh5_0),.dout(w_dff_B_ChDSmj630_0),.clk(gclk));
	jdff dff_B_oFOHarpP0_0(.din(w_dff_B_ChDSmj630_0),.dout(w_dff_B_oFOHarpP0_0),.clk(gclk));
	jdff dff_B_99EVfNFn0_0(.din(w_dff_B_oFOHarpP0_0),.dout(w_dff_B_99EVfNFn0_0),.clk(gclk));
	jdff dff_B_d3FmXBNv1_0(.din(w_dff_B_99EVfNFn0_0),.dout(w_dff_B_d3FmXBNv1_0),.clk(gclk));
	jdff dff_B_P0Yr2uRG2_0(.din(w_dff_B_d3FmXBNv1_0),.dout(w_dff_B_P0Yr2uRG2_0),.clk(gclk));
	jdff dff_B_1Va7SEkL2_0(.din(w_dff_B_P0Yr2uRG2_0),.dout(w_dff_B_1Va7SEkL2_0),.clk(gclk));
	jdff dff_B_2fTAI0Us1_0(.din(w_dff_B_1Va7SEkL2_0),.dout(w_dff_B_2fTAI0Us1_0),.clk(gclk));
	jdff dff_B_6Eg9timZ0_0(.din(w_dff_B_2fTAI0Us1_0),.dout(w_dff_B_6Eg9timZ0_0),.clk(gclk));
	jdff dff_B_1pfZkSI01_0(.din(w_dff_B_6Eg9timZ0_0),.dout(w_dff_B_1pfZkSI01_0),.clk(gclk));
	jdff dff_B_TibFc1XT8_0(.din(w_dff_B_1pfZkSI01_0),.dout(w_dff_B_TibFc1XT8_0),.clk(gclk));
	jdff dff_B_SR7b3DuN5_0(.din(w_dff_B_TibFc1XT8_0),.dout(w_dff_B_SR7b3DuN5_0),.clk(gclk));
	jdff dff_B_Yj5jmHab9_0(.din(w_dff_B_SR7b3DuN5_0),.dout(w_dff_B_Yj5jmHab9_0),.clk(gclk));
	jdff dff_B_WOyGo2ic5_0(.din(w_dff_B_Yj5jmHab9_0),.dout(w_dff_B_WOyGo2ic5_0),.clk(gclk));
	jdff dff_B_ABWPYzyd1_0(.din(w_dff_B_WOyGo2ic5_0),.dout(w_dff_B_ABWPYzyd1_0),.clk(gclk));
	jdff dff_B_Clj5FDQq8_0(.din(w_dff_B_ABWPYzyd1_0),.dout(w_dff_B_Clj5FDQq8_0),.clk(gclk));
	jdff dff_B_DmpqHqSc8_0(.din(w_dff_B_Clj5FDQq8_0),.dout(w_dff_B_DmpqHqSc8_0),.clk(gclk));
	jdff dff_B_J1aLXGbI4_0(.din(w_dff_B_DmpqHqSc8_0),.dout(w_dff_B_J1aLXGbI4_0),.clk(gclk));
	jdff dff_B_N8wg7laN4_0(.din(w_dff_B_J1aLXGbI4_0),.dout(w_dff_B_N8wg7laN4_0),.clk(gclk));
	jdff dff_B_GP5vLHyv2_0(.din(w_dff_B_N8wg7laN4_0),.dout(w_dff_B_GP5vLHyv2_0),.clk(gclk));
	jdff dff_B_Be2Ysxib5_0(.din(w_dff_B_GP5vLHyv2_0),.dout(w_dff_B_Be2Ysxib5_0),.clk(gclk));
	jdff dff_B_gPsQtPnN3_0(.din(w_dff_B_Be2Ysxib5_0),.dout(w_dff_B_gPsQtPnN3_0),.clk(gclk));
	jdff dff_B_A36AN5835_0(.din(w_dff_B_gPsQtPnN3_0),.dout(w_dff_B_A36AN5835_0),.clk(gclk));
	jdff dff_B_My5FkOem5_0(.din(w_dff_B_A36AN5835_0),.dout(w_dff_B_My5FkOem5_0),.clk(gclk));
	jdff dff_B_AErbHNx32_0(.din(w_dff_B_My5FkOem5_0),.dout(w_dff_B_AErbHNx32_0),.clk(gclk));
	jdff dff_B_3lw6lXpq4_0(.din(w_dff_B_AErbHNx32_0),.dout(w_dff_B_3lw6lXpq4_0),.clk(gclk));
	jdff dff_B_e5kn9bDL4_0(.din(w_dff_B_3lw6lXpq4_0),.dout(w_dff_B_e5kn9bDL4_0),.clk(gclk));
	jdff dff_B_WOXC58xL9_0(.din(w_dff_B_e5kn9bDL4_0),.dout(w_dff_B_WOXC58xL9_0),.clk(gclk));
	jdff dff_B_MBNxqEwQ0_0(.din(w_dff_B_WOXC58xL9_0),.dout(w_dff_B_MBNxqEwQ0_0),.clk(gclk));
	jdff dff_B_5wamTYmW5_0(.din(w_dff_B_MBNxqEwQ0_0),.dout(w_dff_B_5wamTYmW5_0),.clk(gclk));
	jdff dff_B_RdYtaUpK3_0(.din(w_dff_B_5wamTYmW5_0),.dout(w_dff_B_RdYtaUpK3_0),.clk(gclk));
	jdff dff_B_nqSKNmyc3_0(.din(w_dff_B_RdYtaUpK3_0),.dout(w_dff_B_nqSKNmyc3_0),.clk(gclk));
	jdff dff_B_7h0FUDYy4_0(.din(w_dff_B_nqSKNmyc3_0),.dout(w_dff_B_7h0FUDYy4_0),.clk(gclk));
	jdff dff_B_QRFl5BpH5_0(.din(w_dff_B_7h0FUDYy4_0),.dout(w_dff_B_QRFl5BpH5_0),.clk(gclk));
	jdff dff_B_lHKGjeth2_0(.din(w_dff_B_QRFl5BpH5_0),.dout(w_dff_B_lHKGjeth2_0),.clk(gclk));
	jdff dff_B_DzG9wZ8R8_0(.din(w_dff_B_lHKGjeth2_0),.dout(w_dff_B_DzG9wZ8R8_0),.clk(gclk));
	jdff dff_B_OetR8HtG3_0(.din(w_dff_B_DzG9wZ8R8_0),.dout(w_dff_B_OetR8HtG3_0),.clk(gclk));
	jdff dff_B_QD3eN4qy0_0(.din(w_dff_B_OetR8HtG3_0),.dout(w_dff_B_QD3eN4qy0_0),.clk(gclk));
	jdff dff_B_xcOhM3897_0(.din(w_dff_B_QD3eN4qy0_0),.dout(w_dff_B_xcOhM3897_0),.clk(gclk));
	jdff dff_B_nsrOx64v5_0(.din(w_dff_B_xcOhM3897_0),.dout(w_dff_B_nsrOx64v5_0),.clk(gclk));
	jdff dff_B_Lw4EMmik2_0(.din(w_dff_B_nsrOx64v5_0),.dout(w_dff_B_Lw4EMmik2_0),.clk(gclk));
	jdff dff_B_vaPzb9Lh3_0(.din(w_dff_B_Lw4EMmik2_0),.dout(w_dff_B_vaPzb9Lh3_0),.clk(gclk));
	jdff dff_B_twdsDPhj4_0(.din(w_dff_B_vaPzb9Lh3_0),.dout(w_dff_B_twdsDPhj4_0),.clk(gclk));
	jdff dff_B_2BgPyPxL1_0(.din(w_dff_B_twdsDPhj4_0),.dout(w_dff_B_2BgPyPxL1_0),.clk(gclk));
	jdff dff_B_cdmP6FRm8_0(.din(w_dff_B_2BgPyPxL1_0),.dout(w_dff_B_cdmP6FRm8_0),.clk(gclk));
	jdff dff_B_3MLd8POT7_0(.din(w_dff_B_cdmP6FRm8_0),.dout(w_dff_B_3MLd8POT7_0),.clk(gclk));
	jdff dff_B_Q6N4BjUs1_0(.din(w_dff_B_3MLd8POT7_0),.dout(w_dff_B_Q6N4BjUs1_0),.clk(gclk));
	jdff dff_B_ZwTS8L4J5_0(.din(w_dff_B_Q6N4BjUs1_0),.dout(w_dff_B_ZwTS8L4J5_0),.clk(gclk));
	jdff dff_B_5eT1uxPd5_0(.din(w_dff_B_ZwTS8L4J5_0),.dout(w_dff_B_5eT1uxPd5_0),.clk(gclk));
	jdff dff_B_1znjDKfO1_0(.din(w_dff_B_5eT1uxPd5_0),.dout(w_dff_B_1znjDKfO1_0),.clk(gclk));
	jdff dff_B_k7saA5fi9_0(.din(w_dff_B_1znjDKfO1_0),.dout(w_dff_B_k7saA5fi9_0),.clk(gclk));
	jdff dff_B_ScYLCaw14_0(.din(w_dff_B_k7saA5fi9_0),.dout(w_dff_B_ScYLCaw14_0),.clk(gclk));
	jdff dff_B_DGImIhA32_0(.din(w_dff_B_ScYLCaw14_0),.dout(w_dff_B_DGImIhA32_0),.clk(gclk));
	jdff dff_B_XVsxPe4A7_0(.din(w_dff_B_DGImIhA32_0),.dout(w_dff_B_XVsxPe4A7_0),.clk(gclk));
	jdff dff_B_ZywCeo2z8_0(.din(w_dff_B_XVsxPe4A7_0),.dout(w_dff_B_ZywCeo2z8_0),.clk(gclk));
	jdff dff_B_lWlKqLvt3_0(.din(w_dff_B_ZywCeo2z8_0),.dout(w_dff_B_lWlKqLvt3_0),.clk(gclk));
	jdff dff_B_YtYriMyZ3_0(.din(w_dff_B_lWlKqLvt3_0),.dout(w_dff_B_YtYriMyZ3_0),.clk(gclk));
	jdff dff_B_IythJWoj7_0(.din(w_dff_B_YtYriMyZ3_0),.dout(w_dff_B_IythJWoj7_0),.clk(gclk));
	jdff dff_B_2877Msfg5_0(.din(w_dff_B_IythJWoj7_0),.dout(w_dff_B_2877Msfg5_0),.clk(gclk));
	jdff dff_B_JRRpibkr5_0(.din(w_dff_B_2877Msfg5_0),.dout(w_dff_B_JRRpibkr5_0),.clk(gclk));
	jdff dff_B_q1Ka5dt06_0(.din(w_dff_B_JRRpibkr5_0),.dout(w_dff_B_q1Ka5dt06_0),.clk(gclk));
	jdff dff_B_LbHYiKyu6_0(.din(w_dff_B_q1Ka5dt06_0),.dout(w_dff_B_LbHYiKyu6_0),.clk(gclk));
	jdff dff_B_8K7Rwd960_0(.din(w_dff_B_LbHYiKyu6_0),.dout(w_dff_B_8K7Rwd960_0),.clk(gclk));
	jdff dff_B_UkkkbCyZ2_0(.din(w_dff_B_8K7Rwd960_0),.dout(w_dff_B_UkkkbCyZ2_0),.clk(gclk));
	jdff dff_B_V6CDGR0q8_0(.din(w_dff_B_UkkkbCyZ2_0),.dout(w_dff_B_V6CDGR0q8_0),.clk(gclk));
	jdff dff_B_pTlsvhYO1_0(.din(w_dff_B_V6CDGR0q8_0),.dout(w_dff_B_pTlsvhYO1_0),.clk(gclk));
	jdff dff_B_QExLkNpv5_0(.din(w_dff_B_pTlsvhYO1_0),.dout(w_dff_B_QExLkNpv5_0),.clk(gclk));
	jdff dff_B_XiOn47WN8_0(.din(w_dff_B_QExLkNpv5_0),.dout(w_dff_B_XiOn47WN8_0),.clk(gclk));
	jdff dff_B_l2bArXxB7_0(.din(w_dff_B_XiOn47WN8_0),.dout(w_dff_B_l2bArXxB7_0),.clk(gclk));
	jdff dff_B_Q93H77K29_0(.din(w_dff_B_l2bArXxB7_0),.dout(w_dff_B_Q93H77K29_0),.clk(gclk));
	jdff dff_B_9qSwlpjO1_0(.din(w_dff_B_Q93H77K29_0),.dout(w_dff_B_9qSwlpjO1_0),.clk(gclk));
	jdff dff_B_x5VFf4df8_0(.din(w_dff_B_9qSwlpjO1_0),.dout(w_dff_B_x5VFf4df8_0),.clk(gclk));
	jdff dff_B_htIWiGFV0_0(.din(w_dff_B_x5VFf4df8_0),.dout(w_dff_B_htIWiGFV0_0),.clk(gclk));
	jdff dff_B_rp9vt6i54_0(.din(w_dff_B_htIWiGFV0_0),.dout(w_dff_B_rp9vt6i54_0),.clk(gclk));
	jdff dff_B_qK05uAH65_0(.din(w_dff_B_rp9vt6i54_0),.dout(w_dff_B_qK05uAH65_0),.clk(gclk));
	jdff dff_B_PLXBpS6r1_0(.din(w_dff_B_qK05uAH65_0),.dout(w_dff_B_PLXBpS6r1_0),.clk(gclk));
	jdff dff_B_lW1mhuSE7_0(.din(w_dff_B_PLXBpS6r1_0),.dout(w_dff_B_lW1mhuSE7_0),.clk(gclk));
	jdff dff_B_HMySgqvW9_0(.din(w_dff_B_lW1mhuSE7_0),.dout(w_dff_B_HMySgqvW9_0),.clk(gclk));
	jdff dff_B_chQOsgIx4_0(.din(w_dff_B_HMySgqvW9_0),.dout(w_dff_B_chQOsgIx4_0),.clk(gclk));
	jdff dff_B_Ld72VMUp9_0(.din(w_dff_B_chQOsgIx4_0),.dout(w_dff_B_Ld72VMUp9_0),.clk(gclk));
	jdff dff_B_LAftCvl50_0(.din(w_dff_B_Ld72VMUp9_0),.dout(w_dff_B_LAftCvl50_0),.clk(gclk));
	jdff dff_B_kagAjCL64_0(.din(w_dff_B_LAftCvl50_0),.dout(w_dff_B_kagAjCL64_0),.clk(gclk));
	jdff dff_B_qjFwTGxP1_1(.din(n1140),.dout(w_dff_B_qjFwTGxP1_1),.clk(gclk));
	jdff dff_B_LtZsPGh25_1(.din(w_dff_B_qjFwTGxP1_1),.dout(w_dff_B_LtZsPGh25_1),.clk(gclk));
	jdff dff_B_dW92EnaZ1_1(.din(w_dff_B_LtZsPGh25_1),.dout(w_dff_B_dW92EnaZ1_1),.clk(gclk));
	jdff dff_B_rDobrcMO9_1(.din(w_dff_B_dW92EnaZ1_1),.dout(w_dff_B_rDobrcMO9_1),.clk(gclk));
	jdff dff_B_TaIFXNXn5_1(.din(w_dff_B_rDobrcMO9_1),.dout(w_dff_B_TaIFXNXn5_1),.clk(gclk));
	jdff dff_B_fTXL76RH1_1(.din(w_dff_B_TaIFXNXn5_1),.dout(w_dff_B_fTXL76RH1_1),.clk(gclk));
	jdff dff_B_SWO1VNoZ6_1(.din(w_dff_B_fTXL76RH1_1),.dout(w_dff_B_SWO1VNoZ6_1),.clk(gclk));
	jdff dff_B_qtwiTqLc8_1(.din(w_dff_B_SWO1VNoZ6_1),.dout(w_dff_B_qtwiTqLc8_1),.clk(gclk));
	jdff dff_B_MyLOtbVu5_1(.din(w_dff_B_qtwiTqLc8_1),.dout(w_dff_B_MyLOtbVu5_1),.clk(gclk));
	jdff dff_B_iTtCN6C14_1(.din(w_dff_B_MyLOtbVu5_1),.dout(w_dff_B_iTtCN6C14_1),.clk(gclk));
	jdff dff_B_9xGNOBzr6_1(.din(w_dff_B_iTtCN6C14_1),.dout(w_dff_B_9xGNOBzr6_1),.clk(gclk));
	jdff dff_B_TYMDtaDg2_1(.din(w_dff_B_9xGNOBzr6_1),.dout(w_dff_B_TYMDtaDg2_1),.clk(gclk));
	jdff dff_B_HpHI2JVg1_1(.din(w_dff_B_TYMDtaDg2_1),.dout(w_dff_B_HpHI2JVg1_1),.clk(gclk));
	jdff dff_B_yY55FNfD7_1(.din(w_dff_B_HpHI2JVg1_1),.dout(w_dff_B_yY55FNfD7_1),.clk(gclk));
	jdff dff_B_IqeghPMR8_1(.din(w_dff_B_yY55FNfD7_1),.dout(w_dff_B_IqeghPMR8_1),.clk(gclk));
	jdff dff_B_keFfFJ6t8_1(.din(w_dff_B_IqeghPMR8_1),.dout(w_dff_B_keFfFJ6t8_1),.clk(gclk));
	jdff dff_B_wsQ3WbNG3_1(.din(w_dff_B_keFfFJ6t8_1),.dout(w_dff_B_wsQ3WbNG3_1),.clk(gclk));
	jdff dff_B_oboScFUG6_1(.din(w_dff_B_wsQ3WbNG3_1),.dout(w_dff_B_oboScFUG6_1),.clk(gclk));
	jdff dff_B_xe0Kf96f6_1(.din(w_dff_B_oboScFUG6_1),.dout(w_dff_B_xe0Kf96f6_1),.clk(gclk));
	jdff dff_B_CGzX8wAP5_1(.din(w_dff_B_xe0Kf96f6_1),.dout(w_dff_B_CGzX8wAP5_1),.clk(gclk));
	jdff dff_B_ZSzkqT5D6_1(.din(w_dff_B_CGzX8wAP5_1),.dout(w_dff_B_ZSzkqT5D6_1),.clk(gclk));
	jdff dff_B_LglLR6kE2_1(.din(w_dff_B_ZSzkqT5D6_1),.dout(w_dff_B_LglLR6kE2_1),.clk(gclk));
	jdff dff_B_QTPQCk5J0_1(.din(w_dff_B_LglLR6kE2_1),.dout(w_dff_B_QTPQCk5J0_1),.clk(gclk));
	jdff dff_B_c8PZR3jf8_1(.din(w_dff_B_QTPQCk5J0_1),.dout(w_dff_B_c8PZR3jf8_1),.clk(gclk));
	jdff dff_B_K09zfacP0_1(.din(w_dff_B_c8PZR3jf8_1),.dout(w_dff_B_K09zfacP0_1),.clk(gclk));
	jdff dff_B_T5fnkjyI2_1(.din(w_dff_B_K09zfacP0_1),.dout(w_dff_B_T5fnkjyI2_1),.clk(gclk));
	jdff dff_B_v5OMq2pA1_1(.din(w_dff_B_T5fnkjyI2_1),.dout(w_dff_B_v5OMq2pA1_1),.clk(gclk));
	jdff dff_B_C0kMhk337_1(.din(w_dff_B_v5OMq2pA1_1),.dout(w_dff_B_C0kMhk337_1),.clk(gclk));
	jdff dff_B_7Mvjc0O61_1(.din(w_dff_B_C0kMhk337_1),.dout(w_dff_B_7Mvjc0O61_1),.clk(gclk));
	jdff dff_B_XM4TILbz7_1(.din(w_dff_B_7Mvjc0O61_1),.dout(w_dff_B_XM4TILbz7_1),.clk(gclk));
	jdff dff_B_QpGGAeox1_1(.din(w_dff_B_XM4TILbz7_1),.dout(w_dff_B_QpGGAeox1_1),.clk(gclk));
	jdff dff_B_WeuonUrS6_1(.din(w_dff_B_QpGGAeox1_1),.dout(w_dff_B_WeuonUrS6_1),.clk(gclk));
	jdff dff_B_B7L9MCGb4_1(.din(w_dff_B_WeuonUrS6_1),.dout(w_dff_B_B7L9MCGb4_1),.clk(gclk));
	jdff dff_B_ycXMBjR54_1(.din(w_dff_B_B7L9MCGb4_1),.dout(w_dff_B_ycXMBjR54_1),.clk(gclk));
	jdff dff_B_KAGggqh48_1(.din(w_dff_B_ycXMBjR54_1),.dout(w_dff_B_KAGggqh48_1),.clk(gclk));
	jdff dff_B_FoMRjuHa9_1(.din(w_dff_B_KAGggqh48_1),.dout(w_dff_B_FoMRjuHa9_1),.clk(gclk));
	jdff dff_B_TyMT8Oai1_1(.din(w_dff_B_FoMRjuHa9_1),.dout(w_dff_B_TyMT8Oai1_1),.clk(gclk));
	jdff dff_B_QThEvbVe3_1(.din(w_dff_B_TyMT8Oai1_1),.dout(w_dff_B_QThEvbVe3_1),.clk(gclk));
	jdff dff_B_2qV6bWAY7_1(.din(w_dff_B_QThEvbVe3_1),.dout(w_dff_B_2qV6bWAY7_1),.clk(gclk));
	jdff dff_B_QhCdLOFK5_1(.din(w_dff_B_2qV6bWAY7_1),.dout(w_dff_B_QhCdLOFK5_1),.clk(gclk));
	jdff dff_B_BlA5O6cd2_1(.din(w_dff_B_QhCdLOFK5_1),.dout(w_dff_B_BlA5O6cd2_1),.clk(gclk));
	jdff dff_B_KFzOiraL5_1(.din(w_dff_B_BlA5O6cd2_1),.dout(w_dff_B_KFzOiraL5_1),.clk(gclk));
	jdff dff_B_7JGkfJtD3_1(.din(w_dff_B_KFzOiraL5_1),.dout(w_dff_B_7JGkfJtD3_1),.clk(gclk));
	jdff dff_B_XV0pEo2l3_1(.din(w_dff_B_7JGkfJtD3_1),.dout(w_dff_B_XV0pEo2l3_1),.clk(gclk));
	jdff dff_B_LKNlVyBz8_1(.din(w_dff_B_XV0pEo2l3_1),.dout(w_dff_B_LKNlVyBz8_1),.clk(gclk));
	jdff dff_B_WNu5eXCK1_1(.din(w_dff_B_LKNlVyBz8_1),.dout(w_dff_B_WNu5eXCK1_1),.clk(gclk));
	jdff dff_B_gObKPTmG6_1(.din(w_dff_B_WNu5eXCK1_1),.dout(w_dff_B_gObKPTmG6_1),.clk(gclk));
	jdff dff_B_cNENFW5t7_1(.din(w_dff_B_gObKPTmG6_1),.dout(w_dff_B_cNENFW5t7_1),.clk(gclk));
	jdff dff_B_0vsjRolz6_1(.din(w_dff_B_cNENFW5t7_1),.dout(w_dff_B_0vsjRolz6_1),.clk(gclk));
	jdff dff_B_Fxvm5vPZ1_1(.din(w_dff_B_0vsjRolz6_1),.dout(w_dff_B_Fxvm5vPZ1_1),.clk(gclk));
	jdff dff_B_sFpfKT8X7_1(.din(w_dff_B_Fxvm5vPZ1_1),.dout(w_dff_B_sFpfKT8X7_1),.clk(gclk));
	jdff dff_B_pFdDnQGj7_1(.din(w_dff_B_sFpfKT8X7_1),.dout(w_dff_B_pFdDnQGj7_1),.clk(gclk));
	jdff dff_B_GNmagbj10_1(.din(w_dff_B_pFdDnQGj7_1),.dout(w_dff_B_GNmagbj10_1),.clk(gclk));
	jdff dff_B_VaZwxek65_1(.din(w_dff_B_GNmagbj10_1),.dout(w_dff_B_VaZwxek65_1),.clk(gclk));
	jdff dff_B_T70BR5b65_1(.din(w_dff_B_VaZwxek65_1),.dout(w_dff_B_T70BR5b65_1),.clk(gclk));
	jdff dff_B_nPV2hRap2_1(.din(w_dff_B_T70BR5b65_1),.dout(w_dff_B_nPV2hRap2_1),.clk(gclk));
	jdff dff_B_BalEm5O52_1(.din(w_dff_B_nPV2hRap2_1),.dout(w_dff_B_BalEm5O52_1),.clk(gclk));
	jdff dff_B_Rhqgx9ps7_1(.din(w_dff_B_BalEm5O52_1),.dout(w_dff_B_Rhqgx9ps7_1),.clk(gclk));
	jdff dff_B_8yRd9DR00_1(.din(w_dff_B_Rhqgx9ps7_1),.dout(w_dff_B_8yRd9DR00_1),.clk(gclk));
	jdff dff_B_aiH2UxQ45_1(.din(w_dff_B_8yRd9DR00_1),.dout(w_dff_B_aiH2UxQ45_1),.clk(gclk));
	jdff dff_B_0j3WZ4HX0_1(.din(w_dff_B_aiH2UxQ45_1),.dout(w_dff_B_0j3WZ4HX0_1),.clk(gclk));
	jdff dff_B_DrP1uDhV9_1(.din(w_dff_B_0j3WZ4HX0_1),.dout(w_dff_B_DrP1uDhV9_1),.clk(gclk));
	jdff dff_B_txnh3JSb9_1(.din(w_dff_B_DrP1uDhV9_1),.dout(w_dff_B_txnh3JSb9_1),.clk(gclk));
	jdff dff_B_ACmiHmq19_1(.din(w_dff_B_txnh3JSb9_1),.dout(w_dff_B_ACmiHmq19_1),.clk(gclk));
	jdff dff_B_yiv7h9zv4_1(.din(w_dff_B_ACmiHmq19_1),.dout(w_dff_B_yiv7h9zv4_1),.clk(gclk));
	jdff dff_B_5SoWRpiD4_1(.din(w_dff_B_yiv7h9zv4_1),.dout(w_dff_B_5SoWRpiD4_1),.clk(gclk));
	jdff dff_B_MpXvo99k6_1(.din(w_dff_B_5SoWRpiD4_1),.dout(w_dff_B_MpXvo99k6_1),.clk(gclk));
	jdff dff_B_FUFG53Ln1_1(.din(w_dff_B_MpXvo99k6_1),.dout(w_dff_B_FUFG53Ln1_1),.clk(gclk));
	jdff dff_B_cwwQTsWZ7_1(.din(w_dff_B_FUFG53Ln1_1),.dout(w_dff_B_cwwQTsWZ7_1),.clk(gclk));
	jdff dff_B_UD1By94n0_1(.din(w_dff_B_cwwQTsWZ7_1),.dout(w_dff_B_UD1By94n0_1),.clk(gclk));
	jdff dff_B_O3NfOOfO1_1(.din(w_dff_B_UD1By94n0_1),.dout(w_dff_B_O3NfOOfO1_1),.clk(gclk));
	jdff dff_B_5Oq74Rxk8_1(.din(w_dff_B_O3NfOOfO1_1),.dout(w_dff_B_5Oq74Rxk8_1),.clk(gclk));
	jdff dff_B_XsxOnK867_1(.din(w_dff_B_5Oq74Rxk8_1),.dout(w_dff_B_XsxOnK867_1),.clk(gclk));
	jdff dff_B_mN8OCDtM7_1(.din(w_dff_B_XsxOnK867_1),.dout(w_dff_B_mN8OCDtM7_1),.clk(gclk));
	jdff dff_B_nS57dSDL7_1(.din(w_dff_B_mN8OCDtM7_1),.dout(w_dff_B_nS57dSDL7_1),.clk(gclk));
	jdff dff_B_BmHiU5VO6_1(.din(w_dff_B_nS57dSDL7_1),.dout(w_dff_B_BmHiU5VO6_1),.clk(gclk));
	jdff dff_B_3VNwujLj4_1(.din(w_dff_B_BmHiU5VO6_1),.dout(w_dff_B_3VNwujLj4_1),.clk(gclk));
	jdff dff_B_Q0alDEF74_1(.din(w_dff_B_3VNwujLj4_1),.dout(w_dff_B_Q0alDEF74_1),.clk(gclk));
	jdff dff_B_sa97GCRl4_1(.din(w_dff_B_Q0alDEF74_1),.dout(w_dff_B_sa97GCRl4_1),.clk(gclk));
	jdff dff_B_szP7HnQ50_1(.din(w_dff_B_sa97GCRl4_1),.dout(w_dff_B_szP7HnQ50_1),.clk(gclk));
	jdff dff_B_u3ipOcjU8_1(.din(w_dff_B_szP7HnQ50_1),.dout(w_dff_B_u3ipOcjU8_1),.clk(gclk));
	jdff dff_B_kn1vR85C7_1(.din(w_dff_B_u3ipOcjU8_1),.dout(w_dff_B_kn1vR85C7_1),.clk(gclk));
	jdff dff_B_G7DdSTmA4_1(.din(w_dff_B_kn1vR85C7_1),.dout(w_dff_B_G7DdSTmA4_1),.clk(gclk));
	jdff dff_B_3nYI5KG06_1(.din(w_dff_B_G7DdSTmA4_1),.dout(w_dff_B_3nYI5KG06_1),.clk(gclk));
	jdff dff_B_fBlOQnWp2_1(.din(w_dff_B_3nYI5KG06_1),.dout(w_dff_B_fBlOQnWp2_1),.clk(gclk));
	jdff dff_B_94aJhMqB6_1(.din(w_dff_B_fBlOQnWp2_1),.dout(w_dff_B_94aJhMqB6_1),.clk(gclk));
	jdff dff_B_KHP2p4OH7_1(.din(w_dff_B_94aJhMqB6_1),.dout(w_dff_B_KHP2p4OH7_1),.clk(gclk));
	jdff dff_B_Ytc35zPu3_1(.din(w_dff_B_KHP2p4OH7_1),.dout(w_dff_B_Ytc35zPu3_1),.clk(gclk));
	jdff dff_B_JVQ57C7i9_1(.din(w_dff_B_Ytc35zPu3_1),.dout(w_dff_B_JVQ57C7i9_1),.clk(gclk));
	jdff dff_B_0s0dPjLj1_1(.din(w_dff_B_JVQ57C7i9_1),.dout(w_dff_B_0s0dPjLj1_1),.clk(gclk));
	jdff dff_B_t1GTVvN16_1(.din(w_dff_B_0s0dPjLj1_1),.dout(w_dff_B_t1GTVvN16_1),.clk(gclk));
	jdff dff_B_0chOpwD94_1(.din(w_dff_B_t1GTVvN16_1),.dout(w_dff_B_0chOpwD94_1),.clk(gclk));
	jdff dff_B_JawOBCjj5_1(.din(w_dff_B_0chOpwD94_1),.dout(w_dff_B_JawOBCjj5_1),.clk(gclk));
	jdff dff_B_U16ejgIK9_1(.din(w_dff_B_JawOBCjj5_1),.dout(w_dff_B_U16ejgIK9_1),.clk(gclk));
	jdff dff_B_EGczAVq93_1(.din(w_dff_B_U16ejgIK9_1),.dout(w_dff_B_EGczAVq93_1),.clk(gclk));
	jdff dff_B_uV8QYM7I5_1(.din(w_dff_B_EGczAVq93_1),.dout(w_dff_B_uV8QYM7I5_1),.clk(gclk));
	jdff dff_B_0KbJmfYC1_1(.din(w_dff_B_uV8QYM7I5_1),.dout(w_dff_B_0KbJmfYC1_1),.clk(gclk));
	jdff dff_B_OScwFDyr0_1(.din(w_dff_B_0KbJmfYC1_1),.dout(w_dff_B_OScwFDyr0_1),.clk(gclk));
	jdff dff_B_j3dgmtwS6_1(.din(w_dff_B_OScwFDyr0_1),.dout(w_dff_B_j3dgmtwS6_1),.clk(gclk));
	jdff dff_B_9LeGDpeM8_1(.din(w_dff_B_j3dgmtwS6_1),.dout(w_dff_B_9LeGDpeM8_1),.clk(gclk));
	jdff dff_B_Au9YUNtD6_1(.din(w_dff_B_9LeGDpeM8_1),.dout(w_dff_B_Au9YUNtD6_1),.clk(gclk));
	jdff dff_B_iTtZdKQ85_1(.din(w_dff_B_Au9YUNtD6_1),.dout(w_dff_B_iTtZdKQ85_1),.clk(gclk));
	jdff dff_B_3SuEsW770_1(.din(w_dff_B_iTtZdKQ85_1),.dout(w_dff_B_3SuEsW770_1),.clk(gclk));
	jdff dff_B_I7tw9qDa5_1(.din(w_dff_B_3SuEsW770_1),.dout(w_dff_B_I7tw9qDa5_1),.clk(gclk));
	jdff dff_B_LaZLcbmA8_1(.din(w_dff_B_I7tw9qDa5_1),.dout(w_dff_B_LaZLcbmA8_1),.clk(gclk));
	jdff dff_B_PXYmFUcf2_1(.din(w_dff_B_LaZLcbmA8_1),.dout(w_dff_B_PXYmFUcf2_1),.clk(gclk));
	jdff dff_B_vqCGRPoq9_1(.din(w_dff_B_PXYmFUcf2_1),.dout(w_dff_B_vqCGRPoq9_1),.clk(gclk));
	jdff dff_B_C5nm0R890_1(.din(w_dff_B_vqCGRPoq9_1),.dout(w_dff_B_C5nm0R890_1),.clk(gclk));
	jdff dff_B_jDEcKhfV6_1(.din(w_dff_B_C5nm0R890_1),.dout(w_dff_B_jDEcKhfV6_1),.clk(gclk));
	jdff dff_B_vbK5iP3S2_1(.din(w_dff_B_jDEcKhfV6_1),.dout(w_dff_B_vbK5iP3S2_1),.clk(gclk));
	jdff dff_B_fF9qNdta0_1(.din(w_dff_B_vbK5iP3S2_1),.dout(w_dff_B_fF9qNdta0_1),.clk(gclk));
	jdff dff_B_fJF763LR9_1(.din(w_dff_B_fF9qNdta0_1),.dout(w_dff_B_fJF763LR9_1),.clk(gclk));
	jdff dff_B_130cv7473_1(.din(w_dff_B_fJF763LR9_1),.dout(w_dff_B_130cv7473_1),.clk(gclk));
	jdff dff_B_JzjrsjBu9_1(.din(w_dff_B_130cv7473_1),.dout(w_dff_B_JzjrsjBu9_1),.clk(gclk));
	jdff dff_B_mJD14FKk0_1(.din(w_dff_B_JzjrsjBu9_1),.dout(w_dff_B_mJD14FKk0_1),.clk(gclk));
	jdff dff_B_Qux1WfCy1_1(.din(w_dff_B_mJD14FKk0_1),.dout(w_dff_B_Qux1WfCy1_1),.clk(gclk));
	jdff dff_B_YuEZvZoQ4_1(.din(w_dff_B_Qux1WfCy1_1),.dout(w_dff_B_YuEZvZoQ4_1),.clk(gclk));
	jdff dff_B_N12tJPel7_1(.din(w_dff_B_YuEZvZoQ4_1),.dout(w_dff_B_N12tJPel7_1),.clk(gclk));
	jdff dff_B_VtuFAYEw0_1(.din(w_dff_B_N12tJPel7_1),.dout(w_dff_B_VtuFAYEw0_1),.clk(gclk));
	jdff dff_B_es37bXV36_1(.din(w_dff_B_VtuFAYEw0_1),.dout(w_dff_B_es37bXV36_1),.clk(gclk));
	jdff dff_B_VPzNwCch5_1(.din(w_dff_B_es37bXV36_1),.dout(w_dff_B_VPzNwCch5_1),.clk(gclk));
	jdff dff_B_QoliabzH9_1(.din(w_dff_B_VPzNwCch5_1),.dout(w_dff_B_QoliabzH9_1),.clk(gclk));
	jdff dff_B_7vxyjbbi2_1(.din(w_dff_B_QoliabzH9_1),.dout(w_dff_B_7vxyjbbi2_1),.clk(gclk));
	jdff dff_B_xndqxWZN7_1(.din(w_dff_B_7vxyjbbi2_1),.dout(w_dff_B_xndqxWZN7_1),.clk(gclk));
	jdff dff_B_DkDpKM995_1(.din(w_dff_B_xndqxWZN7_1),.dout(w_dff_B_DkDpKM995_1),.clk(gclk));
	jdff dff_B_uZVHTY441_1(.din(w_dff_B_DkDpKM995_1),.dout(w_dff_B_uZVHTY441_1),.clk(gclk));
	jdff dff_B_UIfRMMo17_0(.din(n1141),.dout(w_dff_B_UIfRMMo17_0),.clk(gclk));
	jdff dff_B_sEYm1PnX8_0(.din(w_dff_B_UIfRMMo17_0),.dout(w_dff_B_sEYm1PnX8_0),.clk(gclk));
	jdff dff_B_8KdiZ2Z47_0(.din(w_dff_B_sEYm1PnX8_0),.dout(w_dff_B_8KdiZ2Z47_0),.clk(gclk));
	jdff dff_B_OIU4Vtun3_0(.din(w_dff_B_8KdiZ2Z47_0),.dout(w_dff_B_OIU4Vtun3_0),.clk(gclk));
	jdff dff_B_vcMhgbVm8_0(.din(w_dff_B_OIU4Vtun3_0),.dout(w_dff_B_vcMhgbVm8_0),.clk(gclk));
	jdff dff_B_BDBknKSh5_0(.din(w_dff_B_vcMhgbVm8_0),.dout(w_dff_B_BDBknKSh5_0),.clk(gclk));
	jdff dff_B_K4cpapNp1_0(.din(w_dff_B_BDBknKSh5_0),.dout(w_dff_B_K4cpapNp1_0),.clk(gclk));
	jdff dff_B_gh47d6QV4_0(.din(w_dff_B_K4cpapNp1_0),.dout(w_dff_B_gh47d6QV4_0),.clk(gclk));
	jdff dff_B_gYxJyOCt7_0(.din(w_dff_B_gh47d6QV4_0),.dout(w_dff_B_gYxJyOCt7_0),.clk(gclk));
	jdff dff_B_nQcCXD8u0_0(.din(w_dff_B_gYxJyOCt7_0),.dout(w_dff_B_nQcCXD8u0_0),.clk(gclk));
	jdff dff_B_ehj63xts3_0(.din(w_dff_B_nQcCXD8u0_0),.dout(w_dff_B_ehj63xts3_0),.clk(gclk));
	jdff dff_B_7PaJGfIE5_0(.din(w_dff_B_ehj63xts3_0),.dout(w_dff_B_7PaJGfIE5_0),.clk(gclk));
	jdff dff_B_NWKKcmph6_0(.din(w_dff_B_7PaJGfIE5_0),.dout(w_dff_B_NWKKcmph6_0),.clk(gclk));
	jdff dff_B_hJuN2ovf5_0(.din(w_dff_B_NWKKcmph6_0),.dout(w_dff_B_hJuN2ovf5_0),.clk(gclk));
	jdff dff_B_SJH1WdSV3_0(.din(w_dff_B_hJuN2ovf5_0),.dout(w_dff_B_SJH1WdSV3_0),.clk(gclk));
	jdff dff_B_2OKllxAE7_0(.din(w_dff_B_SJH1WdSV3_0),.dout(w_dff_B_2OKllxAE7_0),.clk(gclk));
	jdff dff_B_TAYlzFfb9_0(.din(w_dff_B_2OKllxAE7_0),.dout(w_dff_B_TAYlzFfb9_0),.clk(gclk));
	jdff dff_B_wE5QgV1g8_0(.din(w_dff_B_TAYlzFfb9_0),.dout(w_dff_B_wE5QgV1g8_0),.clk(gclk));
	jdff dff_B_7KhKfUyC7_0(.din(w_dff_B_wE5QgV1g8_0),.dout(w_dff_B_7KhKfUyC7_0),.clk(gclk));
	jdff dff_B_HoSP0Or07_0(.din(w_dff_B_7KhKfUyC7_0),.dout(w_dff_B_HoSP0Or07_0),.clk(gclk));
	jdff dff_B_Cn1zECOW4_0(.din(w_dff_B_HoSP0Or07_0),.dout(w_dff_B_Cn1zECOW4_0),.clk(gclk));
	jdff dff_B_GfXPN2PZ0_0(.din(w_dff_B_Cn1zECOW4_0),.dout(w_dff_B_GfXPN2PZ0_0),.clk(gclk));
	jdff dff_B_tTPtnnub5_0(.din(w_dff_B_GfXPN2PZ0_0),.dout(w_dff_B_tTPtnnub5_0),.clk(gclk));
	jdff dff_B_G10VaWMB6_0(.din(w_dff_B_tTPtnnub5_0),.dout(w_dff_B_G10VaWMB6_0),.clk(gclk));
	jdff dff_B_8T7Deinj5_0(.din(w_dff_B_G10VaWMB6_0),.dout(w_dff_B_8T7Deinj5_0),.clk(gclk));
	jdff dff_B_Wd5Ui0yN3_0(.din(w_dff_B_8T7Deinj5_0),.dout(w_dff_B_Wd5Ui0yN3_0),.clk(gclk));
	jdff dff_B_0sixEjbQ6_0(.din(w_dff_B_Wd5Ui0yN3_0),.dout(w_dff_B_0sixEjbQ6_0),.clk(gclk));
	jdff dff_B_GDVSf4dv0_0(.din(w_dff_B_0sixEjbQ6_0),.dout(w_dff_B_GDVSf4dv0_0),.clk(gclk));
	jdff dff_B_mKPcTAxu1_0(.din(w_dff_B_GDVSf4dv0_0),.dout(w_dff_B_mKPcTAxu1_0),.clk(gclk));
	jdff dff_B_OlPObljC3_0(.din(w_dff_B_mKPcTAxu1_0),.dout(w_dff_B_OlPObljC3_0),.clk(gclk));
	jdff dff_B_oAcq70lk2_0(.din(w_dff_B_OlPObljC3_0),.dout(w_dff_B_oAcq70lk2_0),.clk(gclk));
	jdff dff_B_XkINiefj9_0(.din(w_dff_B_oAcq70lk2_0),.dout(w_dff_B_XkINiefj9_0),.clk(gclk));
	jdff dff_B_8bxpsKze5_0(.din(w_dff_B_XkINiefj9_0),.dout(w_dff_B_8bxpsKze5_0),.clk(gclk));
	jdff dff_B_SF4PPvlF0_0(.din(w_dff_B_8bxpsKze5_0),.dout(w_dff_B_SF4PPvlF0_0),.clk(gclk));
	jdff dff_B_CbEzOaUY6_0(.din(w_dff_B_SF4PPvlF0_0),.dout(w_dff_B_CbEzOaUY6_0),.clk(gclk));
	jdff dff_B_5EOOx0lr4_0(.din(w_dff_B_CbEzOaUY6_0),.dout(w_dff_B_5EOOx0lr4_0),.clk(gclk));
	jdff dff_B_A1tBblZP1_0(.din(w_dff_B_5EOOx0lr4_0),.dout(w_dff_B_A1tBblZP1_0),.clk(gclk));
	jdff dff_B_Mat87lFi1_0(.din(w_dff_B_A1tBblZP1_0),.dout(w_dff_B_Mat87lFi1_0),.clk(gclk));
	jdff dff_B_mcHp6r683_0(.din(w_dff_B_Mat87lFi1_0),.dout(w_dff_B_mcHp6r683_0),.clk(gclk));
	jdff dff_B_KU7I6zKP9_0(.din(w_dff_B_mcHp6r683_0),.dout(w_dff_B_KU7I6zKP9_0),.clk(gclk));
	jdff dff_B_QnzTMJqT8_0(.din(w_dff_B_KU7I6zKP9_0),.dout(w_dff_B_QnzTMJqT8_0),.clk(gclk));
	jdff dff_B_NMAoaklK0_0(.din(w_dff_B_QnzTMJqT8_0),.dout(w_dff_B_NMAoaklK0_0),.clk(gclk));
	jdff dff_B_wdNxyA832_0(.din(w_dff_B_NMAoaklK0_0),.dout(w_dff_B_wdNxyA832_0),.clk(gclk));
	jdff dff_B_3toypXCa5_0(.din(w_dff_B_wdNxyA832_0),.dout(w_dff_B_3toypXCa5_0),.clk(gclk));
	jdff dff_B_YKASeoiX4_0(.din(w_dff_B_3toypXCa5_0),.dout(w_dff_B_YKASeoiX4_0),.clk(gclk));
	jdff dff_B_qAHBOJ486_0(.din(w_dff_B_YKASeoiX4_0),.dout(w_dff_B_qAHBOJ486_0),.clk(gclk));
	jdff dff_B_pzGJ38Re2_0(.din(w_dff_B_qAHBOJ486_0),.dout(w_dff_B_pzGJ38Re2_0),.clk(gclk));
	jdff dff_B_2exID8Tl9_0(.din(w_dff_B_pzGJ38Re2_0),.dout(w_dff_B_2exID8Tl9_0),.clk(gclk));
	jdff dff_B_Y6E4ZdBX8_0(.din(w_dff_B_2exID8Tl9_0),.dout(w_dff_B_Y6E4ZdBX8_0),.clk(gclk));
	jdff dff_B_2s67h5uY5_0(.din(w_dff_B_Y6E4ZdBX8_0),.dout(w_dff_B_2s67h5uY5_0),.clk(gclk));
	jdff dff_B_pbRwGNh50_0(.din(w_dff_B_2s67h5uY5_0),.dout(w_dff_B_pbRwGNh50_0),.clk(gclk));
	jdff dff_B_ReqN87sL7_0(.din(w_dff_B_pbRwGNh50_0),.dout(w_dff_B_ReqN87sL7_0),.clk(gclk));
	jdff dff_B_6FhJ5evS2_0(.din(w_dff_B_ReqN87sL7_0),.dout(w_dff_B_6FhJ5evS2_0),.clk(gclk));
	jdff dff_B_3dqMHn1g2_0(.din(w_dff_B_6FhJ5evS2_0),.dout(w_dff_B_3dqMHn1g2_0),.clk(gclk));
	jdff dff_B_APLbVDTH9_0(.din(w_dff_B_3dqMHn1g2_0),.dout(w_dff_B_APLbVDTH9_0),.clk(gclk));
	jdff dff_B_lMhO8JRY7_0(.din(w_dff_B_APLbVDTH9_0),.dout(w_dff_B_lMhO8JRY7_0),.clk(gclk));
	jdff dff_B_2jCeuxHF1_0(.din(w_dff_B_lMhO8JRY7_0),.dout(w_dff_B_2jCeuxHF1_0),.clk(gclk));
	jdff dff_B_dXUYhB749_0(.din(w_dff_B_2jCeuxHF1_0),.dout(w_dff_B_dXUYhB749_0),.clk(gclk));
	jdff dff_B_W48yjts62_0(.din(w_dff_B_dXUYhB749_0),.dout(w_dff_B_W48yjts62_0),.clk(gclk));
	jdff dff_B_p7p98mYh4_0(.din(w_dff_B_W48yjts62_0),.dout(w_dff_B_p7p98mYh4_0),.clk(gclk));
	jdff dff_B_j7c3tMRw0_0(.din(w_dff_B_p7p98mYh4_0),.dout(w_dff_B_j7c3tMRw0_0),.clk(gclk));
	jdff dff_B_p5TH6L823_0(.din(w_dff_B_j7c3tMRw0_0),.dout(w_dff_B_p5TH6L823_0),.clk(gclk));
	jdff dff_B_6Xmhg7f57_0(.din(w_dff_B_p5TH6L823_0),.dout(w_dff_B_6Xmhg7f57_0),.clk(gclk));
	jdff dff_B_kT7l4loP3_0(.din(w_dff_B_6Xmhg7f57_0),.dout(w_dff_B_kT7l4loP3_0),.clk(gclk));
	jdff dff_B_J1bnMWc63_0(.din(w_dff_B_kT7l4loP3_0),.dout(w_dff_B_J1bnMWc63_0),.clk(gclk));
	jdff dff_B_UAfeS6Mu0_0(.din(w_dff_B_J1bnMWc63_0),.dout(w_dff_B_UAfeS6Mu0_0),.clk(gclk));
	jdff dff_B_rdW3g0p80_0(.din(w_dff_B_UAfeS6Mu0_0),.dout(w_dff_B_rdW3g0p80_0),.clk(gclk));
	jdff dff_B_8m3f4Rrq7_0(.din(w_dff_B_rdW3g0p80_0),.dout(w_dff_B_8m3f4Rrq7_0),.clk(gclk));
	jdff dff_B_IOD82zOu5_0(.din(w_dff_B_8m3f4Rrq7_0),.dout(w_dff_B_IOD82zOu5_0),.clk(gclk));
	jdff dff_B_0uvycL3x0_0(.din(w_dff_B_IOD82zOu5_0),.dout(w_dff_B_0uvycL3x0_0),.clk(gclk));
	jdff dff_B_ZBjdw3w07_0(.din(w_dff_B_0uvycL3x0_0),.dout(w_dff_B_ZBjdw3w07_0),.clk(gclk));
	jdff dff_B_oxf2Vwjv0_0(.din(w_dff_B_ZBjdw3w07_0),.dout(w_dff_B_oxf2Vwjv0_0),.clk(gclk));
	jdff dff_B_DnBCThME5_0(.din(w_dff_B_oxf2Vwjv0_0),.dout(w_dff_B_DnBCThME5_0),.clk(gclk));
	jdff dff_B_FdPlqoNF3_0(.din(w_dff_B_DnBCThME5_0),.dout(w_dff_B_FdPlqoNF3_0),.clk(gclk));
	jdff dff_B_NMFWkd9N5_0(.din(w_dff_B_FdPlqoNF3_0),.dout(w_dff_B_NMFWkd9N5_0),.clk(gclk));
	jdff dff_B_fTphxSUS6_0(.din(w_dff_B_NMFWkd9N5_0),.dout(w_dff_B_fTphxSUS6_0),.clk(gclk));
	jdff dff_B_U7uYyPWd0_0(.din(w_dff_B_fTphxSUS6_0),.dout(w_dff_B_U7uYyPWd0_0),.clk(gclk));
	jdff dff_B_FnDkmIOv6_0(.din(w_dff_B_U7uYyPWd0_0),.dout(w_dff_B_FnDkmIOv6_0),.clk(gclk));
	jdff dff_B_IzXv99gG7_0(.din(w_dff_B_FnDkmIOv6_0),.dout(w_dff_B_IzXv99gG7_0),.clk(gclk));
	jdff dff_B_uW34HRL47_0(.din(w_dff_B_IzXv99gG7_0),.dout(w_dff_B_uW34HRL47_0),.clk(gclk));
	jdff dff_B_pUcGSPB91_0(.din(w_dff_B_uW34HRL47_0),.dout(w_dff_B_pUcGSPB91_0),.clk(gclk));
	jdff dff_B_PYBMFpUb9_0(.din(w_dff_B_pUcGSPB91_0),.dout(w_dff_B_PYBMFpUb9_0),.clk(gclk));
	jdff dff_B_jm6gE8V13_0(.din(w_dff_B_PYBMFpUb9_0),.dout(w_dff_B_jm6gE8V13_0),.clk(gclk));
	jdff dff_B_iF8OvDmU2_0(.din(w_dff_B_jm6gE8V13_0),.dout(w_dff_B_iF8OvDmU2_0),.clk(gclk));
	jdff dff_B_TE85hIov6_0(.din(w_dff_B_iF8OvDmU2_0),.dout(w_dff_B_TE85hIov6_0),.clk(gclk));
	jdff dff_B_XETMNRd40_0(.din(w_dff_B_TE85hIov6_0),.dout(w_dff_B_XETMNRd40_0),.clk(gclk));
	jdff dff_B_YSZ4SavV4_0(.din(w_dff_B_XETMNRd40_0),.dout(w_dff_B_YSZ4SavV4_0),.clk(gclk));
	jdff dff_B_lji79BQR2_0(.din(w_dff_B_YSZ4SavV4_0),.dout(w_dff_B_lji79BQR2_0),.clk(gclk));
	jdff dff_B_gLPIv3Ty4_0(.din(w_dff_B_lji79BQR2_0),.dout(w_dff_B_gLPIv3Ty4_0),.clk(gclk));
	jdff dff_B_ksQmPqfu1_0(.din(w_dff_B_gLPIv3Ty4_0),.dout(w_dff_B_ksQmPqfu1_0),.clk(gclk));
	jdff dff_B_6x9ub2bx4_0(.din(w_dff_B_ksQmPqfu1_0),.dout(w_dff_B_6x9ub2bx4_0),.clk(gclk));
	jdff dff_B_Cl8mEKel8_0(.din(w_dff_B_6x9ub2bx4_0),.dout(w_dff_B_Cl8mEKel8_0),.clk(gclk));
	jdff dff_B_A4SJWYP19_0(.din(w_dff_B_Cl8mEKel8_0),.dout(w_dff_B_A4SJWYP19_0),.clk(gclk));
	jdff dff_B_mTnZeH0p7_0(.din(w_dff_B_A4SJWYP19_0),.dout(w_dff_B_mTnZeH0p7_0),.clk(gclk));
	jdff dff_B_fB6MDpEm1_0(.din(w_dff_B_mTnZeH0p7_0),.dout(w_dff_B_fB6MDpEm1_0),.clk(gclk));
	jdff dff_B_cqAod1e78_0(.din(w_dff_B_fB6MDpEm1_0),.dout(w_dff_B_cqAod1e78_0),.clk(gclk));
	jdff dff_B_W8rLN8me8_0(.din(w_dff_B_cqAod1e78_0),.dout(w_dff_B_W8rLN8me8_0),.clk(gclk));
	jdff dff_B_PmHIsatk6_0(.din(w_dff_B_W8rLN8me8_0),.dout(w_dff_B_PmHIsatk6_0),.clk(gclk));
	jdff dff_B_8FhigV8A8_0(.din(w_dff_B_PmHIsatk6_0),.dout(w_dff_B_8FhigV8A8_0),.clk(gclk));
	jdff dff_B_3CUW0Tyv3_0(.din(w_dff_B_8FhigV8A8_0),.dout(w_dff_B_3CUW0Tyv3_0),.clk(gclk));
	jdff dff_B_agaIgjiY5_0(.din(w_dff_B_3CUW0Tyv3_0),.dout(w_dff_B_agaIgjiY5_0),.clk(gclk));
	jdff dff_B_5QoASS2s3_0(.din(w_dff_B_agaIgjiY5_0),.dout(w_dff_B_5QoASS2s3_0),.clk(gclk));
	jdff dff_B_F6829vpX1_0(.din(w_dff_B_5QoASS2s3_0),.dout(w_dff_B_F6829vpX1_0),.clk(gclk));
	jdff dff_B_CTLNycMm9_0(.din(w_dff_B_F6829vpX1_0),.dout(w_dff_B_CTLNycMm9_0),.clk(gclk));
	jdff dff_B_UkIALfw99_0(.din(w_dff_B_CTLNycMm9_0),.dout(w_dff_B_UkIALfw99_0),.clk(gclk));
	jdff dff_B_DEayxWl14_0(.din(w_dff_B_UkIALfw99_0),.dout(w_dff_B_DEayxWl14_0),.clk(gclk));
	jdff dff_B_6i5RghSa5_0(.din(w_dff_B_DEayxWl14_0),.dout(w_dff_B_6i5RghSa5_0),.clk(gclk));
	jdff dff_B_e2MUULoz3_0(.din(w_dff_B_6i5RghSa5_0),.dout(w_dff_B_e2MUULoz3_0),.clk(gclk));
	jdff dff_B_GUJnZhVb8_0(.din(w_dff_B_e2MUULoz3_0),.dout(w_dff_B_GUJnZhVb8_0),.clk(gclk));
	jdff dff_B_qOClIXxQ1_0(.din(w_dff_B_GUJnZhVb8_0),.dout(w_dff_B_qOClIXxQ1_0),.clk(gclk));
	jdff dff_B_pllzwnu44_0(.din(w_dff_B_qOClIXxQ1_0),.dout(w_dff_B_pllzwnu44_0),.clk(gclk));
	jdff dff_B_7vzSVvY71_0(.din(w_dff_B_pllzwnu44_0),.dout(w_dff_B_7vzSVvY71_0),.clk(gclk));
	jdff dff_B_RZx1FXN96_0(.din(w_dff_B_7vzSVvY71_0),.dout(w_dff_B_RZx1FXN96_0),.clk(gclk));
	jdff dff_B_K9G9WEws1_0(.din(w_dff_B_RZx1FXN96_0),.dout(w_dff_B_K9G9WEws1_0),.clk(gclk));
	jdff dff_B_dlKyWSjy4_0(.din(w_dff_B_K9G9WEws1_0),.dout(w_dff_B_dlKyWSjy4_0),.clk(gclk));
	jdff dff_B_I3zJEqxf4_0(.din(w_dff_B_dlKyWSjy4_0),.dout(w_dff_B_I3zJEqxf4_0),.clk(gclk));
	jdff dff_B_bNbjF7No7_0(.din(w_dff_B_I3zJEqxf4_0),.dout(w_dff_B_bNbjF7No7_0),.clk(gclk));
	jdff dff_B_yB78cJMU8_0(.din(w_dff_B_bNbjF7No7_0),.dout(w_dff_B_yB78cJMU8_0),.clk(gclk));
	jdff dff_B_05sQ1YAL9_0(.din(w_dff_B_yB78cJMU8_0),.dout(w_dff_B_05sQ1YAL9_0),.clk(gclk));
	jdff dff_B_HurN6bGI8_0(.din(w_dff_B_05sQ1YAL9_0),.dout(w_dff_B_HurN6bGI8_0),.clk(gclk));
	jdff dff_B_dXaR3gRJ0_0(.din(w_dff_B_HurN6bGI8_0),.dout(w_dff_B_dXaR3gRJ0_0),.clk(gclk));
	jdff dff_B_N9gTvttA7_0(.din(w_dff_B_dXaR3gRJ0_0),.dout(w_dff_B_N9gTvttA7_0),.clk(gclk));
	jdff dff_B_lrDVgVsa3_0(.din(w_dff_B_N9gTvttA7_0),.dout(w_dff_B_lrDVgVsa3_0),.clk(gclk));
	jdff dff_B_t6WIj8CJ3_0(.din(w_dff_B_lrDVgVsa3_0),.dout(w_dff_B_t6WIj8CJ3_0),.clk(gclk));
	jdff dff_B_3yjLCZJr2_0(.din(w_dff_B_t6WIj8CJ3_0),.dout(w_dff_B_3yjLCZJr2_0),.clk(gclk));
	jdff dff_B_DNEnPLV67_0(.din(w_dff_B_3yjLCZJr2_0),.dout(w_dff_B_DNEnPLV67_0),.clk(gclk));
	jdff dff_B_PeJMRXYm7_1(.din(n1134),.dout(w_dff_B_PeJMRXYm7_1),.clk(gclk));
	jdff dff_B_Wiq7zt4W4_1(.din(w_dff_B_PeJMRXYm7_1),.dout(w_dff_B_Wiq7zt4W4_1),.clk(gclk));
	jdff dff_B_2gazRcPi3_1(.din(w_dff_B_Wiq7zt4W4_1),.dout(w_dff_B_2gazRcPi3_1),.clk(gclk));
	jdff dff_B_sT1NyVZW5_1(.din(w_dff_B_2gazRcPi3_1),.dout(w_dff_B_sT1NyVZW5_1),.clk(gclk));
	jdff dff_B_xeKHbRBE2_1(.din(w_dff_B_sT1NyVZW5_1),.dout(w_dff_B_xeKHbRBE2_1),.clk(gclk));
	jdff dff_B_MsoxdLTO7_1(.din(w_dff_B_xeKHbRBE2_1),.dout(w_dff_B_MsoxdLTO7_1),.clk(gclk));
	jdff dff_B_HA2m0Zgv2_1(.din(w_dff_B_MsoxdLTO7_1),.dout(w_dff_B_HA2m0Zgv2_1),.clk(gclk));
	jdff dff_B_uZln1uGt9_1(.din(w_dff_B_HA2m0Zgv2_1),.dout(w_dff_B_uZln1uGt9_1),.clk(gclk));
	jdff dff_B_TfEDFa7M4_1(.din(w_dff_B_uZln1uGt9_1),.dout(w_dff_B_TfEDFa7M4_1),.clk(gclk));
	jdff dff_B_VBNbnLRv9_1(.din(w_dff_B_TfEDFa7M4_1),.dout(w_dff_B_VBNbnLRv9_1),.clk(gclk));
	jdff dff_B_NMbhZqF13_1(.din(w_dff_B_VBNbnLRv9_1),.dout(w_dff_B_NMbhZqF13_1),.clk(gclk));
	jdff dff_B_GRKZgOnA9_1(.din(w_dff_B_NMbhZqF13_1),.dout(w_dff_B_GRKZgOnA9_1),.clk(gclk));
	jdff dff_B_fgWc8n1X0_1(.din(w_dff_B_GRKZgOnA9_1),.dout(w_dff_B_fgWc8n1X0_1),.clk(gclk));
	jdff dff_B_Y4Lnimlj8_1(.din(w_dff_B_fgWc8n1X0_1),.dout(w_dff_B_Y4Lnimlj8_1),.clk(gclk));
	jdff dff_B_dW8iRuQT6_1(.din(w_dff_B_Y4Lnimlj8_1),.dout(w_dff_B_dW8iRuQT6_1),.clk(gclk));
	jdff dff_B_3SXHIxi50_1(.din(w_dff_B_dW8iRuQT6_1),.dout(w_dff_B_3SXHIxi50_1),.clk(gclk));
	jdff dff_B_tZaEXAva8_1(.din(w_dff_B_3SXHIxi50_1),.dout(w_dff_B_tZaEXAva8_1),.clk(gclk));
	jdff dff_B_ZYlAkPz61_1(.din(w_dff_B_tZaEXAva8_1),.dout(w_dff_B_ZYlAkPz61_1),.clk(gclk));
	jdff dff_B_cLYFJyYG0_1(.din(w_dff_B_ZYlAkPz61_1),.dout(w_dff_B_cLYFJyYG0_1),.clk(gclk));
	jdff dff_B_y5VyVXjM1_1(.din(w_dff_B_cLYFJyYG0_1),.dout(w_dff_B_y5VyVXjM1_1),.clk(gclk));
	jdff dff_B_lZ3nBqQK4_1(.din(w_dff_B_y5VyVXjM1_1),.dout(w_dff_B_lZ3nBqQK4_1),.clk(gclk));
	jdff dff_B_j5JC0dDh6_1(.din(w_dff_B_lZ3nBqQK4_1),.dout(w_dff_B_j5JC0dDh6_1),.clk(gclk));
	jdff dff_B_dWwtbhsU4_1(.din(w_dff_B_j5JC0dDh6_1),.dout(w_dff_B_dWwtbhsU4_1),.clk(gclk));
	jdff dff_B_wQxpwdh25_1(.din(w_dff_B_dWwtbhsU4_1),.dout(w_dff_B_wQxpwdh25_1),.clk(gclk));
	jdff dff_B_c6XBPG3H8_1(.din(w_dff_B_wQxpwdh25_1),.dout(w_dff_B_c6XBPG3H8_1),.clk(gclk));
	jdff dff_B_YP6fwQ929_1(.din(w_dff_B_c6XBPG3H8_1),.dout(w_dff_B_YP6fwQ929_1),.clk(gclk));
	jdff dff_B_ZTkp6LO53_1(.din(w_dff_B_YP6fwQ929_1),.dout(w_dff_B_ZTkp6LO53_1),.clk(gclk));
	jdff dff_B_gXu6JrfR9_1(.din(w_dff_B_ZTkp6LO53_1),.dout(w_dff_B_gXu6JrfR9_1),.clk(gclk));
	jdff dff_B_9iLnkI9X5_1(.din(w_dff_B_gXu6JrfR9_1),.dout(w_dff_B_9iLnkI9X5_1),.clk(gclk));
	jdff dff_B_yBBxLciN0_1(.din(w_dff_B_9iLnkI9X5_1),.dout(w_dff_B_yBBxLciN0_1),.clk(gclk));
	jdff dff_B_Gz5WVE5l6_1(.din(w_dff_B_yBBxLciN0_1),.dout(w_dff_B_Gz5WVE5l6_1),.clk(gclk));
	jdff dff_B_Ce3V9bNW4_1(.din(w_dff_B_Gz5WVE5l6_1),.dout(w_dff_B_Ce3V9bNW4_1),.clk(gclk));
	jdff dff_B_GnAuJlnv8_1(.din(w_dff_B_Ce3V9bNW4_1),.dout(w_dff_B_GnAuJlnv8_1),.clk(gclk));
	jdff dff_B_ehn53vEQ9_1(.din(w_dff_B_GnAuJlnv8_1),.dout(w_dff_B_ehn53vEQ9_1),.clk(gclk));
	jdff dff_B_iiv3RP1D2_1(.din(w_dff_B_ehn53vEQ9_1),.dout(w_dff_B_iiv3RP1D2_1),.clk(gclk));
	jdff dff_B_FxNAlomB1_1(.din(w_dff_B_iiv3RP1D2_1),.dout(w_dff_B_FxNAlomB1_1),.clk(gclk));
	jdff dff_B_u2AVdzzZ3_1(.din(w_dff_B_FxNAlomB1_1),.dout(w_dff_B_u2AVdzzZ3_1),.clk(gclk));
	jdff dff_B_3sFZ7W2j9_1(.din(w_dff_B_u2AVdzzZ3_1),.dout(w_dff_B_3sFZ7W2j9_1),.clk(gclk));
	jdff dff_B_EXsJSvgH9_1(.din(w_dff_B_3sFZ7W2j9_1),.dout(w_dff_B_EXsJSvgH9_1),.clk(gclk));
	jdff dff_B_ntYIyMmg4_1(.din(w_dff_B_EXsJSvgH9_1),.dout(w_dff_B_ntYIyMmg4_1),.clk(gclk));
	jdff dff_B_Eskgs0l44_1(.din(w_dff_B_ntYIyMmg4_1),.dout(w_dff_B_Eskgs0l44_1),.clk(gclk));
	jdff dff_B_fSiQxdSn4_1(.din(w_dff_B_Eskgs0l44_1),.dout(w_dff_B_fSiQxdSn4_1),.clk(gclk));
	jdff dff_B_r5W895SF3_1(.din(w_dff_B_fSiQxdSn4_1),.dout(w_dff_B_r5W895SF3_1),.clk(gclk));
	jdff dff_B_B4JZwX4C6_1(.din(w_dff_B_r5W895SF3_1),.dout(w_dff_B_B4JZwX4C6_1),.clk(gclk));
	jdff dff_B_oI7yG2Ov5_1(.din(w_dff_B_B4JZwX4C6_1),.dout(w_dff_B_oI7yG2Ov5_1),.clk(gclk));
	jdff dff_B_tw7DQOUz7_1(.din(w_dff_B_oI7yG2Ov5_1),.dout(w_dff_B_tw7DQOUz7_1),.clk(gclk));
	jdff dff_B_vhFocqyv4_1(.din(w_dff_B_tw7DQOUz7_1),.dout(w_dff_B_vhFocqyv4_1),.clk(gclk));
	jdff dff_B_NkncWFJK2_1(.din(w_dff_B_vhFocqyv4_1),.dout(w_dff_B_NkncWFJK2_1),.clk(gclk));
	jdff dff_B_rZ8NEeaP6_1(.din(w_dff_B_NkncWFJK2_1),.dout(w_dff_B_rZ8NEeaP6_1),.clk(gclk));
	jdff dff_B_OfHGrOCt1_1(.din(w_dff_B_rZ8NEeaP6_1),.dout(w_dff_B_OfHGrOCt1_1),.clk(gclk));
	jdff dff_B_woq8m1pW8_1(.din(w_dff_B_OfHGrOCt1_1),.dout(w_dff_B_woq8m1pW8_1),.clk(gclk));
	jdff dff_B_lCWMDEcX7_1(.din(w_dff_B_woq8m1pW8_1),.dout(w_dff_B_lCWMDEcX7_1),.clk(gclk));
	jdff dff_B_mxIvtezJ4_1(.din(w_dff_B_lCWMDEcX7_1),.dout(w_dff_B_mxIvtezJ4_1),.clk(gclk));
	jdff dff_B_HLDupKPU2_1(.din(w_dff_B_mxIvtezJ4_1),.dout(w_dff_B_HLDupKPU2_1),.clk(gclk));
	jdff dff_B_73FFJ3sa5_1(.din(w_dff_B_HLDupKPU2_1),.dout(w_dff_B_73FFJ3sa5_1),.clk(gclk));
	jdff dff_B_CgV9igpK7_1(.din(w_dff_B_73FFJ3sa5_1),.dout(w_dff_B_CgV9igpK7_1),.clk(gclk));
	jdff dff_B_Cj5fSiLs3_1(.din(w_dff_B_CgV9igpK7_1),.dout(w_dff_B_Cj5fSiLs3_1),.clk(gclk));
	jdff dff_B_9AuY64Sa9_1(.din(w_dff_B_Cj5fSiLs3_1),.dout(w_dff_B_9AuY64Sa9_1),.clk(gclk));
	jdff dff_B_Q8xiu3zP2_1(.din(w_dff_B_9AuY64Sa9_1),.dout(w_dff_B_Q8xiu3zP2_1),.clk(gclk));
	jdff dff_B_QZGKarUy1_1(.din(w_dff_B_Q8xiu3zP2_1),.dout(w_dff_B_QZGKarUy1_1),.clk(gclk));
	jdff dff_B_vClkgFhS3_1(.din(w_dff_B_QZGKarUy1_1),.dout(w_dff_B_vClkgFhS3_1),.clk(gclk));
	jdff dff_B_YT8xm2Iy4_1(.din(w_dff_B_vClkgFhS3_1),.dout(w_dff_B_YT8xm2Iy4_1),.clk(gclk));
	jdff dff_B_TO3BQIx44_1(.din(w_dff_B_YT8xm2Iy4_1),.dout(w_dff_B_TO3BQIx44_1),.clk(gclk));
	jdff dff_B_bz3EMpQq3_1(.din(w_dff_B_TO3BQIx44_1),.dout(w_dff_B_bz3EMpQq3_1),.clk(gclk));
	jdff dff_B_moqXD66n7_1(.din(w_dff_B_bz3EMpQq3_1),.dout(w_dff_B_moqXD66n7_1),.clk(gclk));
	jdff dff_B_b5S2fOyC0_1(.din(w_dff_B_moqXD66n7_1),.dout(w_dff_B_b5S2fOyC0_1),.clk(gclk));
	jdff dff_B_ok1ZS0Ps8_1(.din(w_dff_B_b5S2fOyC0_1),.dout(w_dff_B_ok1ZS0Ps8_1),.clk(gclk));
	jdff dff_B_MrONCrF44_1(.din(w_dff_B_ok1ZS0Ps8_1),.dout(w_dff_B_MrONCrF44_1),.clk(gclk));
	jdff dff_B_kE4BFMRr0_1(.din(w_dff_B_MrONCrF44_1),.dout(w_dff_B_kE4BFMRr0_1),.clk(gclk));
	jdff dff_B_FgS4MFPD2_1(.din(w_dff_B_kE4BFMRr0_1),.dout(w_dff_B_FgS4MFPD2_1),.clk(gclk));
	jdff dff_B_q2OKyHLx5_1(.din(w_dff_B_FgS4MFPD2_1),.dout(w_dff_B_q2OKyHLx5_1),.clk(gclk));
	jdff dff_B_6KYO2uzd1_1(.din(w_dff_B_q2OKyHLx5_1),.dout(w_dff_B_6KYO2uzd1_1),.clk(gclk));
	jdff dff_B_GR044DAE2_1(.din(w_dff_B_6KYO2uzd1_1),.dout(w_dff_B_GR044DAE2_1),.clk(gclk));
	jdff dff_B_XcQe7W8l6_1(.din(w_dff_B_GR044DAE2_1),.dout(w_dff_B_XcQe7W8l6_1),.clk(gclk));
	jdff dff_B_OtRXcKN75_1(.din(w_dff_B_XcQe7W8l6_1),.dout(w_dff_B_OtRXcKN75_1),.clk(gclk));
	jdff dff_B_vOTZvkpf8_1(.din(w_dff_B_OtRXcKN75_1),.dout(w_dff_B_vOTZvkpf8_1),.clk(gclk));
	jdff dff_B_vKoWYKZv4_1(.din(w_dff_B_vOTZvkpf8_1),.dout(w_dff_B_vKoWYKZv4_1),.clk(gclk));
	jdff dff_B_djybVx9m5_1(.din(w_dff_B_vKoWYKZv4_1),.dout(w_dff_B_djybVx9m5_1),.clk(gclk));
	jdff dff_B_8fq1QfUs8_1(.din(w_dff_B_djybVx9m5_1),.dout(w_dff_B_8fq1QfUs8_1),.clk(gclk));
	jdff dff_B_cCfbTfJ69_1(.din(w_dff_B_8fq1QfUs8_1),.dout(w_dff_B_cCfbTfJ69_1),.clk(gclk));
	jdff dff_B_e1CJdju65_1(.din(w_dff_B_cCfbTfJ69_1),.dout(w_dff_B_e1CJdju65_1),.clk(gclk));
	jdff dff_B_q7oS9qaI6_1(.din(w_dff_B_e1CJdju65_1),.dout(w_dff_B_q7oS9qaI6_1),.clk(gclk));
	jdff dff_B_5fD5dJ1C8_1(.din(w_dff_B_q7oS9qaI6_1),.dout(w_dff_B_5fD5dJ1C8_1),.clk(gclk));
	jdff dff_B_vlqhbnTp1_1(.din(w_dff_B_5fD5dJ1C8_1),.dout(w_dff_B_vlqhbnTp1_1),.clk(gclk));
	jdff dff_B_1baSNXil2_1(.din(w_dff_B_vlqhbnTp1_1),.dout(w_dff_B_1baSNXil2_1),.clk(gclk));
	jdff dff_B_YyUQP1Yz7_1(.din(w_dff_B_1baSNXil2_1),.dout(w_dff_B_YyUQP1Yz7_1),.clk(gclk));
	jdff dff_B_CgvCYpeL9_1(.din(w_dff_B_YyUQP1Yz7_1),.dout(w_dff_B_CgvCYpeL9_1),.clk(gclk));
	jdff dff_B_KWmywiR21_1(.din(w_dff_B_CgvCYpeL9_1),.dout(w_dff_B_KWmywiR21_1),.clk(gclk));
	jdff dff_B_fA0kqpSB9_1(.din(w_dff_B_KWmywiR21_1),.dout(w_dff_B_fA0kqpSB9_1),.clk(gclk));
	jdff dff_B_jkzuCscJ6_1(.din(w_dff_B_fA0kqpSB9_1),.dout(w_dff_B_jkzuCscJ6_1),.clk(gclk));
	jdff dff_B_yP5rpBqu2_1(.din(w_dff_B_jkzuCscJ6_1),.dout(w_dff_B_yP5rpBqu2_1),.clk(gclk));
	jdff dff_B_iikdZxSv7_1(.din(w_dff_B_yP5rpBqu2_1),.dout(w_dff_B_iikdZxSv7_1),.clk(gclk));
	jdff dff_B_W0jaPUOG6_1(.din(w_dff_B_iikdZxSv7_1),.dout(w_dff_B_W0jaPUOG6_1),.clk(gclk));
	jdff dff_B_PXAohauM5_1(.din(w_dff_B_W0jaPUOG6_1),.dout(w_dff_B_PXAohauM5_1),.clk(gclk));
	jdff dff_B_j7qJ5wGm2_1(.din(w_dff_B_PXAohauM5_1),.dout(w_dff_B_j7qJ5wGm2_1),.clk(gclk));
	jdff dff_B_TTGlPZDV5_1(.din(w_dff_B_j7qJ5wGm2_1),.dout(w_dff_B_TTGlPZDV5_1),.clk(gclk));
	jdff dff_B_ZynYgw6A7_1(.din(w_dff_B_TTGlPZDV5_1),.dout(w_dff_B_ZynYgw6A7_1),.clk(gclk));
	jdff dff_B_bmzlTLMw4_1(.din(w_dff_B_ZynYgw6A7_1),.dout(w_dff_B_bmzlTLMw4_1),.clk(gclk));
	jdff dff_B_Uh1CetYi7_1(.din(w_dff_B_bmzlTLMw4_1),.dout(w_dff_B_Uh1CetYi7_1),.clk(gclk));
	jdff dff_B_LVp9OJPG9_1(.din(w_dff_B_Uh1CetYi7_1),.dout(w_dff_B_LVp9OJPG9_1),.clk(gclk));
	jdff dff_B_OTRMn5AT1_1(.din(w_dff_B_LVp9OJPG9_1),.dout(w_dff_B_OTRMn5AT1_1),.clk(gclk));
	jdff dff_B_XNx55mJc4_1(.din(w_dff_B_OTRMn5AT1_1),.dout(w_dff_B_XNx55mJc4_1),.clk(gclk));
	jdff dff_B_WCVQQn2Z4_1(.din(w_dff_B_XNx55mJc4_1),.dout(w_dff_B_WCVQQn2Z4_1),.clk(gclk));
	jdff dff_B_8xeGuheq1_1(.din(w_dff_B_WCVQQn2Z4_1),.dout(w_dff_B_8xeGuheq1_1),.clk(gclk));
	jdff dff_B_8rWM0NSK2_1(.din(w_dff_B_8xeGuheq1_1),.dout(w_dff_B_8rWM0NSK2_1),.clk(gclk));
	jdff dff_B_DpVfeCqn9_1(.din(w_dff_B_8rWM0NSK2_1),.dout(w_dff_B_DpVfeCqn9_1),.clk(gclk));
	jdff dff_B_FLooi0u00_1(.din(w_dff_B_DpVfeCqn9_1),.dout(w_dff_B_FLooi0u00_1),.clk(gclk));
	jdff dff_B_NxsP3JOE5_1(.din(w_dff_B_FLooi0u00_1),.dout(w_dff_B_NxsP3JOE5_1),.clk(gclk));
	jdff dff_B_xSyMuwPc9_1(.din(w_dff_B_NxsP3JOE5_1),.dout(w_dff_B_xSyMuwPc9_1),.clk(gclk));
	jdff dff_B_YPjSjgan5_1(.din(w_dff_B_xSyMuwPc9_1),.dout(w_dff_B_YPjSjgan5_1),.clk(gclk));
	jdff dff_B_zHcoyCFp8_1(.din(w_dff_B_YPjSjgan5_1),.dout(w_dff_B_zHcoyCFp8_1),.clk(gclk));
	jdff dff_B_GY0f20Nd8_1(.din(w_dff_B_zHcoyCFp8_1),.dout(w_dff_B_GY0f20Nd8_1),.clk(gclk));
	jdff dff_B_qZte3hRw7_1(.din(w_dff_B_GY0f20Nd8_1),.dout(w_dff_B_qZte3hRw7_1),.clk(gclk));
	jdff dff_B_8PR18gDU6_1(.din(w_dff_B_qZte3hRw7_1),.dout(w_dff_B_8PR18gDU6_1),.clk(gclk));
	jdff dff_B_GtqqI2B20_1(.din(w_dff_B_8PR18gDU6_1),.dout(w_dff_B_GtqqI2B20_1),.clk(gclk));
	jdff dff_B_I3zmRXlp5_1(.din(w_dff_B_GtqqI2B20_1),.dout(w_dff_B_I3zmRXlp5_1),.clk(gclk));
	jdff dff_B_qgE89aah3_1(.din(w_dff_B_I3zmRXlp5_1),.dout(w_dff_B_qgE89aah3_1),.clk(gclk));
	jdff dff_B_nj5brqWu0_1(.din(w_dff_B_qgE89aah3_1),.dout(w_dff_B_nj5brqWu0_1),.clk(gclk));
	jdff dff_B_NmWQJAZR7_1(.din(w_dff_B_nj5brqWu0_1),.dout(w_dff_B_NmWQJAZR7_1),.clk(gclk));
	jdff dff_B_yTS1F6IJ9_1(.din(w_dff_B_NmWQJAZR7_1),.dout(w_dff_B_yTS1F6IJ9_1),.clk(gclk));
	jdff dff_B_ZVxn8VaI5_1(.din(w_dff_B_yTS1F6IJ9_1),.dout(w_dff_B_ZVxn8VaI5_1),.clk(gclk));
	jdff dff_B_zUudwbrL0_1(.din(w_dff_B_ZVxn8VaI5_1),.dout(w_dff_B_zUudwbrL0_1),.clk(gclk));
	jdff dff_B_19MZpVs95_1(.din(w_dff_B_zUudwbrL0_1),.dout(w_dff_B_19MZpVs95_1),.clk(gclk));
	jdff dff_B_lUBrKJW10_1(.din(w_dff_B_19MZpVs95_1),.dout(w_dff_B_lUBrKJW10_1),.clk(gclk));
	jdff dff_B_cdHtn6570_1(.din(w_dff_B_lUBrKJW10_1),.dout(w_dff_B_cdHtn6570_1),.clk(gclk));
	jdff dff_B_IMnVun0Q4_0(.din(n1135),.dout(w_dff_B_IMnVun0Q4_0),.clk(gclk));
	jdff dff_B_VAjhsi152_0(.din(w_dff_B_IMnVun0Q4_0),.dout(w_dff_B_VAjhsi152_0),.clk(gclk));
	jdff dff_B_Ixsoupfq3_0(.din(w_dff_B_VAjhsi152_0),.dout(w_dff_B_Ixsoupfq3_0),.clk(gclk));
	jdff dff_B_EQRSAtTk3_0(.din(w_dff_B_Ixsoupfq3_0),.dout(w_dff_B_EQRSAtTk3_0),.clk(gclk));
	jdff dff_B_TLcepq6k1_0(.din(w_dff_B_EQRSAtTk3_0),.dout(w_dff_B_TLcepq6k1_0),.clk(gclk));
	jdff dff_B_fQZLxhSm3_0(.din(w_dff_B_TLcepq6k1_0),.dout(w_dff_B_fQZLxhSm3_0),.clk(gclk));
	jdff dff_B_4uq5uk1e2_0(.din(w_dff_B_fQZLxhSm3_0),.dout(w_dff_B_4uq5uk1e2_0),.clk(gclk));
	jdff dff_B_ntVLpPRX3_0(.din(w_dff_B_4uq5uk1e2_0),.dout(w_dff_B_ntVLpPRX3_0),.clk(gclk));
	jdff dff_B_z1gylA3Q9_0(.din(w_dff_B_ntVLpPRX3_0),.dout(w_dff_B_z1gylA3Q9_0),.clk(gclk));
	jdff dff_B_OrwUJUdw2_0(.din(w_dff_B_z1gylA3Q9_0),.dout(w_dff_B_OrwUJUdw2_0),.clk(gclk));
	jdff dff_B_edf8jYCF8_0(.din(w_dff_B_OrwUJUdw2_0),.dout(w_dff_B_edf8jYCF8_0),.clk(gclk));
	jdff dff_B_PnV34B7w1_0(.din(w_dff_B_edf8jYCF8_0),.dout(w_dff_B_PnV34B7w1_0),.clk(gclk));
	jdff dff_B_8DldS5Cp0_0(.din(w_dff_B_PnV34B7w1_0),.dout(w_dff_B_8DldS5Cp0_0),.clk(gclk));
	jdff dff_B_oW1zYRmF0_0(.din(w_dff_B_8DldS5Cp0_0),.dout(w_dff_B_oW1zYRmF0_0),.clk(gclk));
	jdff dff_B_tgWlweE71_0(.din(w_dff_B_oW1zYRmF0_0),.dout(w_dff_B_tgWlweE71_0),.clk(gclk));
	jdff dff_B_J6Y7qPpE9_0(.din(w_dff_B_tgWlweE71_0),.dout(w_dff_B_J6Y7qPpE9_0),.clk(gclk));
	jdff dff_B_qjzBuBzg3_0(.din(w_dff_B_J6Y7qPpE9_0),.dout(w_dff_B_qjzBuBzg3_0),.clk(gclk));
	jdff dff_B_oqchZ6051_0(.din(w_dff_B_qjzBuBzg3_0),.dout(w_dff_B_oqchZ6051_0),.clk(gclk));
	jdff dff_B_V3QrYPJO2_0(.din(w_dff_B_oqchZ6051_0),.dout(w_dff_B_V3QrYPJO2_0),.clk(gclk));
	jdff dff_B_rjdoaBX81_0(.din(w_dff_B_V3QrYPJO2_0),.dout(w_dff_B_rjdoaBX81_0),.clk(gclk));
	jdff dff_B_zAWkoLjI6_0(.din(w_dff_B_rjdoaBX81_0),.dout(w_dff_B_zAWkoLjI6_0),.clk(gclk));
	jdff dff_B_JsKDRV3C8_0(.din(w_dff_B_zAWkoLjI6_0),.dout(w_dff_B_JsKDRV3C8_0),.clk(gclk));
	jdff dff_B_WhF391KJ4_0(.din(w_dff_B_JsKDRV3C8_0),.dout(w_dff_B_WhF391KJ4_0),.clk(gclk));
	jdff dff_B_sB3hWUCX2_0(.din(w_dff_B_WhF391KJ4_0),.dout(w_dff_B_sB3hWUCX2_0),.clk(gclk));
	jdff dff_B_66SgVw1a1_0(.din(w_dff_B_sB3hWUCX2_0),.dout(w_dff_B_66SgVw1a1_0),.clk(gclk));
	jdff dff_B_kZMA0rtj5_0(.din(w_dff_B_66SgVw1a1_0),.dout(w_dff_B_kZMA0rtj5_0),.clk(gclk));
	jdff dff_B_gdCCQYfR3_0(.din(w_dff_B_kZMA0rtj5_0),.dout(w_dff_B_gdCCQYfR3_0),.clk(gclk));
	jdff dff_B_4lD30sUO7_0(.din(w_dff_B_gdCCQYfR3_0),.dout(w_dff_B_4lD30sUO7_0),.clk(gclk));
	jdff dff_B_wpCC2XWU0_0(.din(w_dff_B_4lD30sUO7_0),.dout(w_dff_B_wpCC2XWU0_0),.clk(gclk));
	jdff dff_B_F6QzjSia3_0(.din(w_dff_B_wpCC2XWU0_0),.dout(w_dff_B_F6QzjSia3_0),.clk(gclk));
	jdff dff_B_IEIK7X0Y5_0(.din(w_dff_B_F6QzjSia3_0),.dout(w_dff_B_IEIK7X0Y5_0),.clk(gclk));
	jdff dff_B_pG3rpEGJ8_0(.din(w_dff_B_IEIK7X0Y5_0),.dout(w_dff_B_pG3rpEGJ8_0),.clk(gclk));
	jdff dff_B_BGA3TmS48_0(.din(w_dff_B_pG3rpEGJ8_0),.dout(w_dff_B_BGA3TmS48_0),.clk(gclk));
	jdff dff_B_GU0xIJok8_0(.din(w_dff_B_BGA3TmS48_0),.dout(w_dff_B_GU0xIJok8_0),.clk(gclk));
	jdff dff_B_FDmijpER7_0(.din(w_dff_B_GU0xIJok8_0),.dout(w_dff_B_FDmijpER7_0),.clk(gclk));
	jdff dff_B_7AEMpKiG2_0(.din(w_dff_B_FDmijpER7_0),.dout(w_dff_B_7AEMpKiG2_0),.clk(gclk));
	jdff dff_B_wJ749GZi2_0(.din(w_dff_B_7AEMpKiG2_0),.dout(w_dff_B_wJ749GZi2_0),.clk(gclk));
	jdff dff_B_Rf01G3uW1_0(.din(w_dff_B_wJ749GZi2_0),.dout(w_dff_B_Rf01G3uW1_0),.clk(gclk));
	jdff dff_B_WMy4NIXB7_0(.din(w_dff_B_Rf01G3uW1_0),.dout(w_dff_B_WMy4NIXB7_0),.clk(gclk));
	jdff dff_B_G4MNqFtJ3_0(.din(w_dff_B_WMy4NIXB7_0),.dout(w_dff_B_G4MNqFtJ3_0),.clk(gclk));
	jdff dff_B_J9bsXzV72_0(.din(w_dff_B_G4MNqFtJ3_0),.dout(w_dff_B_J9bsXzV72_0),.clk(gclk));
	jdff dff_B_yX6gfEQc1_0(.din(w_dff_B_J9bsXzV72_0),.dout(w_dff_B_yX6gfEQc1_0),.clk(gclk));
	jdff dff_B_lmlGSbUF3_0(.din(w_dff_B_yX6gfEQc1_0),.dout(w_dff_B_lmlGSbUF3_0),.clk(gclk));
	jdff dff_B_tT4OUdiy7_0(.din(w_dff_B_lmlGSbUF3_0),.dout(w_dff_B_tT4OUdiy7_0),.clk(gclk));
	jdff dff_B_MPcLLEvy5_0(.din(w_dff_B_tT4OUdiy7_0),.dout(w_dff_B_MPcLLEvy5_0),.clk(gclk));
	jdff dff_B_8sGAn65s6_0(.din(w_dff_B_MPcLLEvy5_0),.dout(w_dff_B_8sGAn65s6_0),.clk(gclk));
	jdff dff_B_ZQuoN1vj4_0(.din(w_dff_B_8sGAn65s6_0),.dout(w_dff_B_ZQuoN1vj4_0),.clk(gclk));
	jdff dff_B_K7JEPbt00_0(.din(w_dff_B_ZQuoN1vj4_0),.dout(w_dff_B_K7JEPbt00_0),.clk(gclk));
	jdff dff_B_sO04ZVAK5_0(.din(w_dff_B_K7JEPbt00_0),.dout(w_dff_B_sO04ZVAK5_0),.clk(gclk));
	jdff dff_B_9bIks27h4_0(.din(w_dff_B_sO04ZVAK5_0),.dout(w_dff_B_9bIks27h4_0),.clk(gclk));
	jdff dff_B_PGSfgcW68_0(.din(w_dff_B_9bIks27h4_0),.dout(w_dff_B_PGSfgcW68_0),.clk(gclk));
	jdff dff_B_86JATPbA0_0(.din(w_dff_B_PGSfgcW68_0),.dout(w_dff_B_86JATPbA0_0),.clk(gclk));
	jdff dff_B_QTuAey3s3_0(.din(w_dff_B_86JATPbA0_0),.dout(w_dff_B_QTuAey3s3_0),.clk(gclk));
	jdff dff_B_UHWEwQSi7_0(.din(w_dff_B_QTuAey3s3_0),.dout(w_dff_B_UHWEwQSi7_0),.clk(gclk));
	jdff dff_B_OcX2W1w95_0(.din(w_dff_B_UHWEwQSi7_0),.dout(w_dff_B_OcX2W1w95_0),.clk(gclk));
	jdff dff_B_UAiq6hR03_0(.din(w_dff_B_OcX2W1w95_0),.dout(w_dff_B_UAiq6hR03_0),.clk(gclk));
	jdff dff_B_6ylJCuaV5_0(.din(w_dff_B_UAiq6hR03_0),.dout(w_dff_B_6ylJCuaV5_0),.clk(gclk));
	jdff dff_B_MOSNjWBY3_0(.din(w_dff_B_6ylJCuaV5_0),.dout(w_dff_B_MOSNjWBY3_0),.clk(gclk));
	jdff dff_B_w3VS5xRg5_0(.din(w_dff_B_MOSNjWBY3_0),.dout(w_dff_B_w3VS5xRg5_0),.clk(gclk));
	jdff dff_B_1NVCE82i5_0(.din(w_dff_B_w3VS5xRg5_0),.dout(w_dff_B_1NVCE82i5_0),.clk(gclk));
	jdff dff_B_8KX8VFWz4_0(.din(w_dff_B_1NVCE82i5_0),.dout(w_dff_B_8KX8VFWz4_0),.clk(gclk));
	jdff dff_B_Cg23HPDG3_0(.din(w_dff_B_8KX8VFWz4_0),.dout(w_dff_B_Cg23HPDG3_0),.clk(gclk));
	jdff dff_B_mliKyHbN2_0(.din(w_dff_B_Cg23HPDG3_0),.dout(w_dff_B_mliKyHbN2_0),.clk(gclk));
	jdff dff_B_V1byI0Ol4_0(.din(w_dff_B_mliKyHbN2_0),.dout(w_dff_B_V1byI0Ol4_0),.clk(gclk));
	jdff dff_B_TMNy6PmX6_0(.din(w_dff_B_V1byI0Ol4_0),.dout(w_dff_B_TMNy6PmX6_0),.clk(gclk));
	jdff dff_B_Gew0W3Sr4_0(.din(w_dff_B_TMNy6PmX6_0),.dout(w_dff_B_Gew0W3Sr4_0),.clk(gclk));
	jdff dff_B_a1U805450_0(.din(w_dff_B_Gew0W3Sr4_0),.dout(w_dff_B_a1U805450_0),.clk(gclk));
	jdff dff_B_6f6WCIrx7_0(.din(w_dff_B_a1U805450_0),.dout(w_dff_B_6f6WCIrx7_0),.clk(gclk));
	jdff dff_B_vv5kaedV9_0(.din(w_dff_B_6f6WCIrx7_0),.dout(w_dff_B_vv5kaedV9_0),.clk(gclk));
	jdff dff_B_n79wEXfz3_0(.din(w_dff_B_vv5kaedV9_0),.dout(w_dff_B_n79wEXfz3_0),.clk(gclk));
	jdff dff_B_6uJn5AC98_0(.din(w_dff_B_n79wEXfz3_0),.dout(w_dff_B_6uJn5AC98_0),.clk(gclk));
	jdff dff_B_o4nmDaC89_0(.din(w_dff_B_6uJn5AC98_0),.dout(w_dff_B_o4nmDaC89_0),.clk(gclk));
	jdff dff_B_OZuFnDnY0_0(.din(w_dff_B_o4nmDaC89_0),.dout(w_dff_B_OZuFnDnY0_0),.clk(gclk));
	jdff dff_B_JXaLon864_0(.din(w_dff_B_OZuFnDnY0_0),.dout(w_dff_B_JXaLon864_0),.clk(gclk));
	jdff dff_B_iOrtRVcg5_0(.din(w_dff_B_JXaLon864_0),.dout(w_dff_B_iOrtRVcg5_0),.clk(gclk));
	jdff dff_B_ge1i3KHv5_0(.din(w_dff_B_iOrtRVcg5_0),.dout(w_dff_B_ge1i3KHv5_0),.clk(gclk));
	jdff dff_B_vcgDCCJj4_0(.din(w_dff_B_ge1i3KHv5_0),.dout(w_dff_B_vcgDCCJj4_0),.clk(gclk));
	jdff dff_B_LOUOG8p22_0(.din(w_dff_B_vcgDCCJj4_0),.dout(w_dff_B_LOUOG8p22_0),.clk(gclk));
	jdff dff_B_MToH7Jdj3_0(.din(w_dff_B_LOUOG8p22_0),.dout(w_dff_B_MToH7Jdj3_0),.clk(gclk));
	jdff dff_B_jHXk46My1_0(.din(w_dff_B_MToH7Jdj3_0),.dout(w_dff_B_jHXk46My1_0),.clk(gclk));
	jdff dff_B_pDBIaVaB3_0(.din(w_dff_B_jHXk46My1_0),.dout(w_dff_B_pDBIaVaB3_0),.clk(gclk));
	jdff dff_B_b9itHejq2_0(.din(w_dff_B_pDBIaVaB3_0),.dout(w_dff_B_b9itHejq2_0),.clk(gclk));
	jdff dff_B_sK6nx3kW4_0(.din(w_dff_B_b9itHejq2_0),.dout(w_dff_B_sK6nx3kW4_0),.clk(gclk));
	jdff dff_B_0NHkqqYB9_0(.din(w_dff_B_sK6nx3kW4_0),.dout(w_dff_B_0NHkqqYB9_0),.clk(gclk));
	jdff dff_B_Vw1HvXim9_0(.din(w_dff_B_0NHkqqYB9_0),.dout(w_dff_B_Vw1HvXim9_0),.clk(gclk));
	jdff dff_B_CEp2nxG80_0(.din(w_dff_B_Vw1HvXim9_0),.dout(w_dff_B_CEp2nxG80_0),.clk(gclk));
	jdff dff_B_CQZJfCA03_0(.din(w_dff_B_CEp2nxG80_0),.dout(w_dff_B_CQZJfCA03_0),.clk(gclk));
	jdff dff_B_ciFCD8mz4_0(.din(w_dff_B_CQZJfCA03_0),.dout(w_dff_B_ciFCD8mz4_0),.clk(gclk));
	jdff dff_B_vSHuAQsA7_0(.din(w_dff_B_ciFCD8mz4_0),.dout(w_dff_B_vSHuAQsA7_0),.clk(gclk));
	jdff dff_B_1PWnsKMM0_0(.din(w_dff_B_vSHuAQsA7_0),.dout(w_dff_B_1PWnsKMM0_0),.clk(gclk));
	jdff dff_B_VcH6Qt5e8_0(.din(w_dff_B_1PWnsKMM0_0),.dout(w_dff_B_VcH6Qt5e8_0),.clk(gclk));
	jdff dff_B_ADb1uOCp2_0(.din(w_dff_B_VcH6Qt5e8_0),.dout(w_dff_B_ADb1uOCp2_0),.clk(gclk));
	jdff dff_B_iVlYBZ2r1_0(.din(w_dff_B_ADb1uOCp2_0),.dout(w_dff_B_iVlYBZ2r1_0),.clk(gclk));
	jdff dff_B_vjwpUNmO4_0(.din(w_dff_B_iVlYBZ2r1_0),.dout(w_dff_B_vjwpUNmO4_0),.clk(gclk));
	jdff dff_B_LWLymFrt1_0(.din(w_dff_B_vjwpUNmO4_0),.dout(w_dff_B_LWLymFrt1_0),.clk(gclk));
	jdff dff_B_G8sbiDlD9_0(.din(w_dff_B_LWLymFrt1_0),.dout(w_dff_B_G8sbiDlD9_0),.clk(gclk));
	jdff dff_B_blWbO9755_0(.din(w_dff_B_G8sbiDlD9_0),.dout(w_dff_B_blWbO9755_0),.clk(gclk));
	jdff dff_B_u6Rv9ZsP2_0(.din(w_dff_B_blWbO9755_0),.dout(w_dff_B_u6Rv9ZsP2_0),.clk(gclk));
	jdff dff_B_n0eQyWeG0_0(.din(w_dff_B_u6Rv9ZsP2_0),.dout(w_dff_B_n0eQyWeG0_0),.clk(gclk));
	jdff dff_B_kwMRE6wA3_0(.din(w_dff_B_n0eQyWeG0_0),.dout(w_dff_B_kwMRE6wA3_0),.clk(gclk));
	jdff dff_B_FWLe1q7S2_0(.din(w_dff_B_kwMRE6wA3_0),.dout(w_dff_B_FWLe1q7S2_0),.clk(gclk));
	jdff dff_B_1ugbiaKb4_0(.din(w_dff_B_FWLe1q7S2_0),.dout(w_dff_B_1ugbiaKb4_0),.clk(gclk));
	jdff dff_B_cm9WZrdO1_0(.din(w_dff_B_1ugbiaKb4_0),.dout(w_dff_B_cm9WZrdO1_0),.clk(gclk));
	jdff dff_B_CbHCSJUA3_0(.din(w_dff_B_cm9WZrdO1_0),.dout(w_dff_B_CbHCSJUA3_0),.clk(gclk));
	jdff dff_B_DTokUmuG5_0(.din(w_dff_B_CbHCSJUA3_0),.dout(w_dff_B_DTokUmuG5_0),.clk(gclk));
	jdff dff_B_0vreo1EL3_0(.din(w_dff_B_DTokUmuG5_0),.dout(w_dff_B_0vreo1EL3_0),.clk(gclk));
	jdff dff_B_cRzaImJV4_0(.din(w_dff_B_0vreo1EL3_0),.dout(w_dff_B_cRzaImJV4_0),.clk(gclk));
	jdff dff_B_A2ESqh3h9_0(.din(w_dff_B_cRzaImJV4_0),.dout(w_dff_B_A2ESqh3h9_0),.clk(gclk));
	jdff dff_B_YrV7BLld1_0(.din(w_dff_B_A2ESqh3h9_0),.dout(w_dff_B_YrV7BLld1_0),.clk(gclk));
	jdff dff_B_lJAXRhCf6_0(.din(w_dff_B_YrV7BLld1_0),.dout(w_dff_B_lJAXRhCf6_0),.clk(gclk));
	jdff dff_B_OkhOkxN08_0(.din(w_dff_B_lJAXRhCf6_0),.dout(w_dff_B_OkhOkxN08_0),.clk(gclk));
	jdff dff_B_DzyeuD2h9_0(.din(w_dff_B_OkhOkxN08_0),.dout(w_dff_B_DzyeuD2h9_0),.clk(gclk));
	jdff dff_B_aMON1cWP4_0(.din(w_dff_B_DzyeuD2h9_0),.dout(w_dff_B_aMON1cWP4_0),.clk(gclk));
	jdff dff_B_zdX2rrMt1_0(.din(w_dff_B_aMON1cWP4_0),.dout(w_dff_B_zdX2rrMt1_0),.clk(gclk));
	jdff dff_B_JNK6Lsyf7_0(.din(w_dff_B_zdX2rrMt1_0),.dout(w_dff_B_JNK6Lsyf7_0),.clk(gclk));
	jdff dff_B_Roaq9tY26_0(.din(w_dff_B_JNK6Lsyf7_0),.dout(w_dff_B_Roaq9tY26_0),.clk(gclk));
	jdff dff_B_pUvYqRzk6_0(.din(w_dff_B_Roaq9tY26_0),.dout(w_dff_B_pUvYqRzk6_0),.clk(gclk));
	jdff dff_B_o4kFetsG5_0(.din(w_dff_B_pUvYqRzk6_0),.dout(w_dff_B_o4kFetsG5_0),.clk(gclk));
	jdff dff_B_fTvzuKQH5_0(.din(w_dff_B_o4kFetsG5_0),.dout(w_dff_B_fTvzuKQH5_0),.clk(gclk));
	jdff dff_B_bDPP2thR9_0(.din(w_dff_B_fTvzuKQH5_0),.dout(w_dff_B_bDPP2thR9_0),.clk(gclk));
	jdff dff_B_s4dAHRDt0_0(.din(w_dff_B_bDPP2thR9_0),.dout(w_dff_B_s4dAHRDt0_0),.clk(gclk));
	jdff dff_B_c2ue1IU29_0(.din(w_dff_B_s4dAHRDt0_0),.dout(w_dff_B_c2ue1IU29_0),.clk(gclk));
	jdff dff_B_sfOAAu5Y1_0(.din(w_dff_B_c2ue1IU29_0),.dout(w_dff_B_sfOAAu5Y1_0),.clk(gclk));
	jdff dff_B_Q63QvkbE0_0(.din(w_dff_B_sfOAAu5Y1_0),.dout(w_dff_B_Q63QvkbE0_0),.clk(gclk));
	jdff dff_B_B43o3NKK2_0(.din(w_dff_B_Q63QvkbE0_0),.dout(w_dff_B_B43o3NKK2_0),.clk(gclk));
	jdff dff_B_oqYIPTeU4_1(.din(n1128),.dout(w_dff_B_oqYIPTeU4_1),.clk(gclk));
	jdff dff_B_tczRxsH46_1(.din(w_dff_B_oqYIPTeU4_1),.dout(w_dff_B_tczRxsH46_1),.clk(gclk));
	jdff dff_B_94Gh0IAv1_1(.din(w_dff_B_tczRxsH46_1),.dout(w_dff_B_94Gh0IAv1_1),.clk(gclk));
	jdff dff_B_XvVnduTm9_1(.din(w_dff_B_94Gh0IAv1_1),.dout(w_dff_B_XvVnduTm9_1),.clk(gclk));
	jdff dff_B_rNTs7xoz3_1(.din(w_dff_B_XvVnduTm9_1),.dout(w_dff_B_rNTs7xoz3_1),.clk(gclk));
	jdff dff_B_6JR2JrYa2_1(.din(w_dff_B_rNTs7xoz3_1),.dout(w_dff_B_6JR2JrYa2_1),.clk(gclk));
	jdff dff_B_sQjGRBF71_1(.din(w_dff_B_6JR2JrYa2_1),.dout(w_dff_B_sQjGRBF71_1),.clk(gclk));
	jdff dff_B_EDAuk2Xe2_1(.din(w_dff_B_sQjGRBF71_1),.dout(w_dff_B_EDAuk2Xe2_1),.clk(gclk));
	jdff dff_B_FgnK8xl14_1(.din(w_dff_B_EDAuk2Xe2_1),.dout(w_dff_B_FgnK8xl14_1),.clk(gclk));
	jdff dff_B_uBHNsLnf1_1(.din(w_dff_B_FgnK8xl14_1),.dout(w_dff_B_uBHNsLnf1_1),.clk(gclk));
	jdff dff_B_INXEK2Sg7_1(.din(w_dff_B_uBHNsLnf1_1),.dout(w_dff_B_INXEK2Sg7_1),.clk(gclk));
	jdff dff_B_GmlP5Xla5_1(.din(w_dff_B_INXEK2Sg7_1),.dout(w_dff_B_GmlP5Xla5_1),.clk(gclk));
	jdff dff_B_MnxEDMVB5_1(.din(w_dff_B_GmlP5Xla5_1),.dout(w_dff_B_MnxEDMVB5_1),.clk(gclk));
	jdff dff_B_MTCX9mng9_1(.din(w_dff_B_MnxEDMVB5_1),.dout(w_dff_B_MTCX9mng9_1),.clk(gclk));
	jdff dff_B_qYZaejB08_1(.din(w_dff_B_MTCX9mng9_1),.dout(w_dff_B_qYZaejB08_1),.clk(gclk));
	jdff dff_B_cMZ91g1w8_1(.din(w_dff_B_qYZaejB08_1),.dout(w_dff_B_cMZ91g1w8_1),.clk(gclk));
	jdff dff_B_oMOrSPYN7_1(.din(w_dff_B_cMZ91g1w8_1),.dout(w_dff_B_oMOrSPYN7_1),.clk(gclk));
	jdff dff_B_BXYP1xeg3_1(.din(w_dff_B_oMOrSPYN7_1),.dout(w_dff_B_BXYP1xeg3_1),.clk(gclk));
	jdff dff_B_AHH63meh4_1(.din(w_dff_B_BXYP1xeg3_1),.dout(w_dff_B_AHH63meh4_1),.clk(gclk));
	jdff dff_B_d9kr3czF9_1(.din(w_dff_B_AHH63meh4_1),.dout(w_dff_B_d9kr3czF9_1),.clk(gclk));
	jdff dff_B_UtVzCpwt7_1(.din(w_dff_B_d9kr3czF9_1),.dout(w_dff_B_UtVzCpwt7_1),.clk(gclk));
	jdff dff_B_0WpDxjBa2_1(.din(w_dff_B_UtVzCpwt7_1),.dout(w_dff_B_0WpDxjBa2_1),.clk(gclk));
	jdff dff_B_ZcROiVMY9_1(.din(w_dff_B_0WpDxjBa2_1),.dout(w_dff_B_ZcROiVMY9_1),.clk(gclk));
	jdff dff_B_ufTqqo5U5_1(.din(w_dff_B_ZcROiVMY9_1),.dout(w_dff_B_ufTqqo5U5_1),.clk(gclk));
	jdff dff_B_CDvLvOWq8_1(.din(w_dff_B_ufTqqo5U5_1),.dout(w_dff_B_CDvLvOWq8_1),.clk(gclk));
	jdff dff_B_nvs7VNKf2_1(.din(w_dff_B_CDvLvOWq8_1),.dout(w_dff_B_nvs7VNKf2_1),.clk(gclk));
	jdff dff_B_FplUPSm90_1(.din(w_dff_B_nvs7VNKf2_1),.dout(w_dff_B_FplUPSm90_1),.clk(gclk));
	jdff dff_B_MahhnMRB5_1(.din(w_dff_B_FplUPSm90_1),.dout(w_dff_B_MahhnMRB5_1),.clk(gclk));
	jdff dff_B_DFKLVSkq8_1(.din(w_dff_B_MahhnMRB5_1),.dout(w_dff_B_DFKLVSkq8_1),.clk(gclk));
	jdff dff_B_txR1o5Zc9_1(.din(w_dff_B_DFKLVSkq8_1),.dout(w_dff_B_txR1o5Zc9_1),.clk(gclk));
	jdff dff_B_fyi9rg8v3_1(.din(w_dff_B_txR1o5Zc9_1),.dout(w_dff_B_fyi9rg8v3_1),.clk(gclk));
	jdff dff_B_LV0zw84p6_1(.din(w_dff_B_fyi9rg8v3_1),.dout(w_dff_B_LV0zw84p6_1),.clk(gclk));
	jdff dff_B_FWEQGw1X9_1(.din(w_dff_B_LV0zw84p6_1),.dout(w_dff_B_FWEQGw1X9_1),.clk(gclk));
	jdff dff_B_ZxzevGlQ1_1(.din(w_dff_B_FWEQGw1X9_1),.dout(w_dff_B_ZxzevGlQ1_1),.clk(gclk));
	jdff dff_B_9ql3iZh97_1(.din(w_dff_B_ZxzevGlQ1_1),.dout(w_dff_B_9ql3iZh97_1),.clk(gclk));
	jdff dff_B_XVc5QF827_1(.din(w_dff_B_9ql3iZh97_1),.dout(w_dff_B_XVc5QF827_1),.clk(gclk));
	jdff dff_B_fjNElSGi8_1(.din(w_dff_B_XVc5QF827_1),.dout(w_dff_B_fjNElSGi8_1),.clk(gclk));
	jdff dff_B_vsWrkZtp1_1(.din(w_dff_B_fjNElSGi8_1),.dout(w_dff_B_vsWrkZtp1_1),.clk(gclk));
	jdff dff_B_X9CsLi1a8_1(.din(w_dff_B_vsWrkZtp1_1),.dout(w_dff_B_X9CsLi1a8_1),.clk(gclk));
	jdff dff_B_hKtTLNWx7_1(.din(w_dff_B_X9CsLi1a8_1),.dout(w_dff_B_hKtTLNWx7_1),.clk(gclk));
	jdff dff_B_WPMBjTXD5_1(.din(w_dff_B_hKtTLNWx7_1),.dout(w_dff_B_WPMBjTXD5_1),.clk(gclk));
	jdff dff_B_ybwBwObn5_1(.din(w_dff_B_WPMBjTXD5_1),.dout(w_dff_B_ybwBwObn5_1),.clk(gclk));
	jdff dff_B_dG6QAN7L1_1(.din(w_dff_B_ybwBwObn5_1),.dout(w_dff_B_dG6QAN7L1_1),.clk(gclk));
	jdff dff_B_PUCooeSz0_1(.din(w_dff_B_dG6QAN7L1_1),.dout(w_dff_B_PUCooeSz0_1),.clk(gclk));
	jdff dff_B_1jMSfx4V9_1(.din(w_dff_B_PUCooeSz0_1),.dout(w_dff_B_1jMSfx4V9_1),.clk(gclk));
	jdff dff_B_j0u58wpI3_1(.din(w_dff_B_1jMSfx4V9_1),.dout(w_dff_B_j0u58wpI3_1),.clk(gclk));
	jdff dff_B_w58al6FC3_1(.din(w_dff_B_j0u58wpI3_1),.dout(w_dff_B_w58al6FC3_1),.clk(gclk));
	jdff dff_B_SmpS2Qz92_1(.din(w_dff_B_w58al6FC3_1),.dout(w_dff_B_SmpS2Qz92_1),.clk(gclk));
	jdff dff_B_ETZ2rAul2_1(.din(w_dff_B_SmpS2Qz92_1),.dout(w_dff_B_ETZ2rAul2_1),.clk(gclk));
	jdff dff_B_akscmYcW3_1(.din(w_dff_B_ETZ2rAul2_1),.dout(w_dff_B_akscmYcW3_1),.clk(gclk));
	jdff dff_B_b6lpjkdW7_1(.din(w_dff_B_akscmYcW3_1),.dout(w_dff_B_b6lpjkdW7_1),.clk(gclk));
	jdff dff_B_7jBWCWQc8_1(.din(w_dff_B_b6lpjkdW7_1),.dout(w_dff_B_7jBWCWQc8_1),.clk(gclk));
	jdff dff_B_1MyMxmme0_1(.din(w_dff_B_7jBWCWQc8_1),.dout(w_dff_B_1MyMxmme0_1),.clk(gclk));
	jdff dff_B_A48oSovy9_1(.din(w_dff_B_1MyMxmme0_1),.dout(w_dff_B_A48oSovy9_1),.clk(gclk));
	jdff dff_B_f3QWxPvS1_1(.din(w_dff_B_A48oSovy9_1),.dout(w_dff_B_f3QWxPvS1_1),.clk(gclk));
	jdff dff_B_FdaaEdc90_1(.din(w_dff_B_f3QWxPvS1_1),.dout(w_dff_B_FdaaEdc90_1),.clk(gclk));
	jdff dff_B_WX9EqciO9_1(.din(w_dff_B_FdaaEdc90_1),.dout(w_dff_B_WX9EqciO9_1),.clk(gclk));
	jdff dff_B_JlDiXBcc5_1(.din(w_dff_B_WX9EqciO9_1),.dout(w_dff_B_JlDiXBcc5_1),.clk(gclk));
	jdff dff_B_uJZLxMzu9_1(.din(w_dff_B_JlDiXBcc5_1),.dout(w_dff_B_uJZLxMzu9_1),.clk(gclk));
	jdff dff_B_ewjeKkt57_1(.din(w_dff_B_uJZLxMzu9_1),.dout(w_dff_B_ewjeKkt57_1),.clk(gclk));
	jdff dff_B_zNb99BgK9_1(.din(w_dff_B_ewjeKkt57_1),.dout(w_dff_B_zNb99BgK9_1),.clk(gclk));
	jdff dff_B_yCb8gJMo4_1(.din(w_dff_B_zNb99BgK9_1),.dout(w_dff_B_yCb8gJMo4_1),.clk(gclk));
	jdff dff_B_GwhiUGWz6_1(.din(w_dff_B_yCb8gJMo4_1),.dout(w_dff_B_GwhiUGWz6_1),.clk(gclk));
	jdff dff_B_PyafcMaX9_1(.din(w_dff_B_GwhiUGWz6_1),.dout(w_dff_B_PyafcMaX9_1),.clk(gclk));
	jdff dff_B_1NTTxpba1_1(.din(w_dff_B_PyafcMaX9_1),.dout(w_dff_B_1NTTxpba1_1),.clk(gclk));
	jdff dff_B_TmiynQBN1_1(.din(w_dff_B_1NTTxpba1_1),.dout(w_dff_B_TmiynQBN1_1),.clk(gclk));
	jdff dff_B_ZCOOpv8o9_1(.din(w_dff_B_TmiynQBN1_1),.dout(w_dff_B_ZCOOpv8o9_1),.clk(gclk));
	jdff dff_B_W6zwAjlI8_1(.din(w_dff_B_ZCOOpv8o9_1),.dout(w_dff_B_W6zwAjlI8_1),.clk(gclk));
	jdff dff_B_7T53m27X3_1(.din(w_dff_B_W6zwAjlI8_1),.dout(w_dff_B_7T53m27X3_1),.clk(gclk));
	jdff dff_B_JgzDgTE35_1(.din(w_dff_B_7T53m27X3_1),.dout(w_dff_B_JgzDgTE35_1),.clk(gclk));
	jdff dff_B_voazf92t0_1(.din(w_dff_B_JgzDgTE35_1),.dout(w_dff_B_voazf92t0_1),.clk(gclk));
	jdff dff_B_tpLLy3Nz5_1(.din(w_dff_B_voazf92t0_1),.dout(w_dff_B_tpLLy3Nz5_1),.clk(gclk));
	jdff dff_B_yqCccnhz8_1(.din(w_dff_B_tpLLy3Nz5_1),.dout(w_dff_B_yqCccnhz8_1),.clk(gclk));
	jdff dff_B_dNhs6sjE3_1(.din(w_dff_B_yqCccnhz8_1),.dout(w_dff_B_dNhs6sjE3_1),.clk(gclk));
	jdff dff_B_qs6ENmwM9_1(.din(w_dff_B_dNhs6sjE3_1),.dout(w_dff_B_qs6ENmwM9_1),.clk(gclk));
	jdff dff_B_FTFsp5691_1(.din(w_dff_B_qs6ENmwM9_1),.dout(w_dff_B_FTFsp5691_1),.clk(gclk));
	jdff dff_B_YgFGocW31_1(.din(w_dff_B_FTFsp5691_1),.dout(w_dff_B_YgFGocW31_1),.clk(gclk));
	jdff dff_B_alByZtzp2_1(.din(w_dff_B_YgFGocW31_1),.dout(w_dff_B_alByZtzp2_1),.clk(gclk));
	jdff dff_B_IRMbgUJC1_1(.din(w_dff_B_alByZtzp2_1),.dout(w_dff_B_IRMbgUJC1_1),.clk(gclk));
	jdff dff_B_v9XqOznu2_1(.din(w_dff_B_IRMbgUJC1_1),.dout(w_dff_B_v9XqOznu2_1),.clk(gclk));
	jdff dff_B_0n6r3ASl7_1(.din(w_dff_B_v9XqOznu2_1),.dout(w_dff_B_0n6r3ASl7_1),.clk(gclk));
	jdff dff_B_z25WlsvQ2_1(.din(w_dff_B_0n6r3ASl7_1),.dout(w_dff_B_z25WlsvQ2_1),.clk(gclk));
	jdff dff_B_pnGvleuN1_1(.din(w_dff_B_z25WlsvQ2_1),.dout(w_dff_B_pnGvleuN1_1),.clk(gclk));
	jdff dff_B_diEdI7F51_1(.din(w_dff_B_pnGvleuN1_1),.dout(w_dff_B_diEdI7F51_1),.clk(gclk));
	jdff dff_B_ZNS5qQJ09_1(.din(w_dff_B_diEdI7F51_1),.dout(w_dff_B_ZNS5qQJ09_1),.clk(gclk));
	jdff dff_B_FIuPFV7o8_1(.din(w_dff_B_ZNS5qQJ09_1),.dout(w_dff_B_FIuPFV7o8_1),.clk(gclk));
	jdff dff_B_nrVoCE1H5_1(.din(w_dff_B_FIuPFV7o8_1),.dout(w_dff_B_nrVoCE1H5_1),.clk(gclk));
	jdff dff_B_0DsO1CXd1_1(.din(w_dff_B_nrVoCE1H5_1),.dout(w_dff_B_0DsO1CXd1_1),.clk(gclk));
	jdff dff_B_YUEfFZ5L7_1(.din(w_dff_B_0DsO1CXd1_1),.dout(w_dff_B_YUEfFZ5L7_1),.clk(gclk));
	jdff dff_B_v2mJS4Ls8_1(.din(w_dff_B_YUEfFZ5L7_1),.dout(w_dff_B_v2mJS4Ls8_1),.clk(gclk));
	jdff dff_B_wtPgOPWs2_1(.din(w_dff_B_v2mJS4Ls8_1),.dout(w_dff_B_wtPgOPWs2_1),.clk(gclk));
	jdff dff_B_9ALlXqTx1_1(.din(w_dff_B_wtPgOPWs2_1),.dout(w_dff_B_9ALlXqTx1_1),.clk(gclk));
	jdff dff_B_G452Aqi41_1(.din(w_dff_B_9ALlXqTx1_1),.dout(w_dff_B_G452Aqi41_1),.clk(gclk));
	jdff dff_B_RMo9ksG02_1(.din(w_dff_B_G452Aqi41_1),.dout(w_dff_B_RMo9ksG02_1),.clk(gclk));
	jdff dff_B_PvgHgzWU1_1(.din(w_dff_B_RMo9ksG02_1),.dout(w_dff_B_PvgHgzWU1_1),.clk(gclk));
	jdff dff_B_p1QddroD8_1(.din(w_dff_B_PvgHgzWU1_1),.dout(w_dff_B_p1QddroD8_1),.clk(gclk));
	jdff dff_B_RS4PnBFr1_1(.din(w_dff_B_p1QddroD8_1),.dout(w_dff_B_RS4PnBFr1_1),.clk(gclk));
	jdff dff_B_33mC7kB02_1(.din(w_dff_B_RS4PnBFr1_1),.dout(w_dff_B_33mC7kB02_1),.clk(gclk));
	jdff dff_B_1NxulKpu3_1(.din(w_dff_B_33mC7kB02_1),.dout(w_dff_B_1NxulKpu3_1),.clk(gclk));
	jdff dff_B_ONvdAm0F7_1(.din(w_dff_B_1NxulKpu3_1),.dout(w_dff_B_ONvdAm0F7_1),.clk(gclk));
	jdff dff_B_LYWOGmNa2_1(.din(w_dff_B_ONvdAm0F7_1),.dout(w_dff_B_LYWOGmNa2_1),.clk(gclk));
	jdff dff_B_umajNF3R8_1(.din(w_dff_B_LYWOGmNa2_1),.dout(w_dff_B_umajNF3R8_1),.clk(gclk));
	jdff dff_B_VeU5RgRJ8_1(.din(w_dff_B_umajNF3R8_1),.dout(w_dff_B_VeU5RgRJ8_1),.clk(gclk));
	jdff dff_B_s8eJBhyK0_1(.din(w_dff_B_VeU5RgRJ8_1),.dout(w_dff_B_s8eJBhyK0_1),.clk(gclk));
	jdff dff_B_UWk2V1Pd2_1(.din(w_dff_B_s8eJBhyK0_1),.dout(w_dff_B_UWk2V1Pd2_1),.clk(gclk));
	jdff dff_B_5evCLscw5_1(.din(w_dff_B_UWk2V1Pd2_1),.dout(w_dff_B_5evCLscw5_1),.clk(gclk));
	jdff dff_B_T1nghpIG3_1(.din(w_dff_B_5evCLscw5_1),.dout(w_dff_B_T1nghpIG3_1),.clk(gclk));
	jdff dff_B_e1tHOO0X9_1(.din(w_dff_B_T1nghpIG3_1),.dout(w_dff_B_e1tHOO0X9_1),.clk(gclk));
	jdff dff_B_5bCn8Jlu3_1(.din(w_dff_B_e1tHOO0X9_1),.dout(w_dff_B_5bCn8Jlu3_1),.clk(gclk));
	jdff dff_B_xE3dXEMe3_1(.din(w_dff_B_5bCn8Jlu3_1),.dout(w_dff_B_xE3dXEMe3_1),.clk(gclk));
	jdff dff_B_peXNoHOm5_1(.din(w_dff_B_xE3dXEMe3_1),.dout(w_dff_B_peXNoHOm5_1),.clk(gclk));
	jdff dff_B_9YhTGdo50_1(.din(w_dff_B_peXNoHOm5_1),.dout(w_dff_B_9YhTGdo50_1),.clk(gclk));
	jdff dff_B_ZJIp1DiE6_1(.din(w_dff_B_9YhTGdo50_1),.dout(w_dff_B_ZJIp1DiE6_1),.clk(gclk));
	jdff dff_B_Ro3hG1000_1(.din(w_dff_B_ZJIp1DiE6_1),.dout(w_dff_B_Ro3hG1000_1),.clk(gclk));
	jdff dff_B_IOCsQ4RV2_1(.din(w_dff_B_Ro3hG1000_1),.dout(w_dff_B_IOCsQ4RV2_1),.clk(gclk));
	jdff dff_B_604l9mpP4_1(.din(w_dff_B_IOCsQ4RV2_1),.dout(w_dff_B_604l9mpP4_1),.clk(gclk));
	jdff dff_B_UO7xfXY45_1(.din(w_dff_B_604l9mpP4_1),.dout(w_dff_B_UO7xfXY45_1),.clk(gclk));
	jdff dff_B_beTjcDsf8_1(.din(w_dff_B_UO7xfXY45_1),.dout(w_dff_B_beTjcDsf8_1),.clk(gclk));
	jdff dff_B_6TPkIcMj8_1(.din(w_dff_B_beTjcDsf8_1),.dout(w_dff_B_6TPkIcMj8_1),.clk(gclk));
	jdff dff_B_dHP4styR0_1(.din(w_dff_B_6TPkIcMj8_1),.dout(w_dff_B_dHP4styR0_1),.clk(gclk));
	jdff dff_B_PKoAfIOJ3_1(.din(w_dff_B_dHP4styR0_1),.dout(w_dff_B_PKoAfIOJ3_1),.clk(gclk));
	jdff dff_B_BiApeeNs4_1(.din(w_dff_B_PKoAfIOJ3_1),.dout(w_dff_B_BiApeeNs4_1),.clk(gclk));
	jdff dff_B_tBVIKrr45_1(.din(w_dff_B_BiApeeNs4_1),.dout(w_dff_B_tBVIKrr45_1),.clk(gclk));
	jdff dff_B_WOhTpZP77_1(.din(w_dff_B_tBVIKrr45_1),.dout(w_dff_B_WOhTpZP77_1),.clk(gclk));
	jdff dff_B_w2UCqheB3_0(.din(n1129),.dout(w_dff_B_w2UCqheB3_0),.clk(gclk));
	jdff dff_B_HpGTHQgg6_0(.din(w_dff_B_w2UCqheB3_0),.dout(w_dff_B_HpGTHQgg6_0),.clk(gclk));
	jdff dff_B_CvmUCDRx5_0(.din(w_dff_B_HpGTHQgg6_0),.dout(w_dff_B_CvmUCDRx5_0),.clk(gclk));
	jdff dff_B_AujreAjX9_0(.din(w_dff_B_CvmUCDRx5_0),.dout(w_dff_B_AujreAjX9_0),.clk(gclk));
	jdff dff_B_R1Cc6msq6_0(.din(w_dff_B_AujreAjX9_0),.dout(w_dff_B_R1Cc6msq6_0),.clk(gclk));
	jdff dff_B_Xegf7MA70_0(.din(w_dff_B_R1Cc6msq6_0),.dout(w_dff_B_Xegf7MA70_0),.clk(gclk));
	jdff dff_B_bxDlTe5U9_0(.din(w_dff_B_Xegf7MA70_0),.dout(w_dff_B_bxDlTe5U9_0),.clk(gclk));
	jdff dff_B_ORPkQi6C5_0(.din(w_dff_B_bxDlTe5U9_0),.dout(w_dff_B_ORPkQi6C5_0),.clk(gclk));
	jdff dff_B_uufp58WE3_0(.din(w_dff_B_ORPkQi6C5_0),.dout(w_dff_B_uufp58WE3_0),.clk(gclk));
	jdff dff_B_DPYAbrse2_0(.din(w_dff_B_uufp58WE3_0),.dout(w_dff_B_DPYAbrse2_0),.clk(gclk));
	jdff dff_B_jiF5o9EO0_0(.din(w_dff_B_DPYAbrse2_0),.dout(w_dff_B_jiF5o9EO0_0),.clk(gclk));
	jdff dff_B_CgGeWtOV6_0(.din(w_dff_B_jiF5o9EO0_0),.dout(w_dff_B_CgGeWtOV6_0),.clk(gclk));
	jdff dff_B_u4tJx7aG3_0(.din(w_dff_B_CgGeWtOV6_0),.dout(w_dff_B_u4tJx7aG3_0),.clk(gclk));
	jdff dff_B_0GuDs4pM9_0(.din(w_dff_B_u4tJx7aG3_0),.dout(w_dff_B_0GuDs4pM9_0),.clk(gclk));
	jdff dff_B_UYsi4ikq6_0(.din(w_dff_B_0GuDs4pM9_0),.dout(w_dff_B_UYsi4ikq6_0),.clk(gclk));
	jdff dff_B_2MQqjAKP6_0(.din(w_dff_B_UYsi4ikq6_0),.dout(w_dff_B_2MQqjAKP6_0),.clk(gclk));
	jdff dff_B_Nwen2Gf48_0(.din(w_dff_B_2MQqjAKP6_0),.dout(w_dff_B_Nwen2Gf48_0),.clk(gclk));
	jdff dff_B_Oc2ksfoM5_0(.din(w_dff_B_Nwen2Gf48_0),.dout(w_dff_B_Oc2ksfoM5_0),.clk(gclk));
	jdff dff_B_DEh6uNc78_0(.din(w_dff_B_Oc2ksfoM5_0),.dout(w_dff_B_DEh6uNc78_0),.clk(gclk));
	jdff dff_B_0bHlZmKc5_0(.din(w_dff_B_DEh6uNc78_0),.dout(w_dff_B_0bHlZmKc5_0),.clk(gclk));
	jdff dff_B_i1XNPAwE8_0(.din(w_dff_B_0bHlZmKc5_0),.dout(w_dff_B_i1XNPAwE8_0),.clk(gclk));
	jdff dff_B_hasKDMsR0_0(.din(w_dff_B_i1XNPAwE8_0),.dout(w_dff_B_hasKDMsR0_0),.clk(gclk));
	jdff dff_B_DEsPVo3N8_0(.din(w_dff_B_hasKDMsR0_0),.dout(w_dff_B_DEsPVo3N8_0),.clk(gclk));
	jdff dff_B_HVt6udWA8_0(.din(w_dff_B_DEsPVo3N8_0),.dout(w_dff_B_HVt6udWA8_0),.clk(gclk));
	jdff dff_B_NESNjduk9_0(.din(w_dff_B_HVt6udWA8_0),.dout(w_dff_B_NESNjduk9_0),.clk(gclk));
	jdff dff_B_AMT9FJqQ7_0(.din(w_dff_B_NESNjduk9_0),.dout(w_dff_B_AMT9FJqQ7_0),.clk(gclk));
	jdff dff_B_KnOO89J35_0(.din(w_dff_B_AMT9FJqQ7_0),.dout(w_dff_B_KnOO89J35_0),.clk(gclk));
	jdff dff_B_2uodiFBb9_0(.din(w_dff_B_KnOO89J35_0),.dout(w_dff_B_2uodiFBb9_0),.clk(gclk));
	jdff dff_B_GLG2pbkc1_0(.din(w_dff_B_2uodiFBb9_0),.dout(w_dff_B_GLG2pbkc1_0),.clk(gclk));
	jdff dff_B_Bk5mbJEd8_0(.din(w_dff_B_GLG2pbkc1_0),.dout(w_dff_B_Bk5mbJEd8_0),.clk(gclk));
	jdff dff_B_uioYmElR4_0(.din(w_dff_B_Bk5mbJEd8_0),.dout(w_dff_B_uioYmElR4_0),.clk(gclk));
	jdff dff_B_gwao8SRb2_0(.din(w_dff_B_uioYmElR4_0),.dout(w_dff_B_gwao8SRb2_0),.clk(gclk));
	jdff dff_B_NXEfhIWO4_0(.din(w_dff_B_gwao8SRb2_0),.dout(w_dff_B_NXEfhIWO4_0),.clk(gclk));
	jdff dff_B_I6JWxblv6_0(.din(w_dff_B_NXEfhIWO4_0),.dout(w_dff_B_I6JWxblv6_0),.clk(gclk));
	jdff dff_B_P1MrBnLi0_0(.din(w_dff_B_I6JWxblv6_0),.dout(w_dff_B_P1MrBnLi0_0),.clk(gclk));
	jdff dff_B_rn3dF23u3_0(.din(w_dff_B_P1MrBnLi0_0),.dout(w_dff_B_rn3dF23u3_0),.clk(gclk));
	jdff dff_B_fHEgJ9xt0_0(.din(w_dff_B_rn3dF23u3_0),.dout(w_dff_B_fHEgJ9xt0_0),.clk(gclk));
	jdff dff_B_WvEAAH396_0(.din(w_dff_B_fHEgJ9xt0_0),.dout(w_dff_B_WvEAAH396_0),.clk(gclk));
	jdff dff_B_Or6unfsz9_0(.din(w_dff_B_WvEAAH396_0),.dout(w_dff_B_Or6unfsz9_0),.clk(gclk));
	jdff dff_B_ZQ79dYv42_0(.din(w_dff_B_Or6unfsz9_0),.dout(w_dff_B_ZQ79dYv42_0),.clk(gclk));
	jdff dff_B_VgMkRi0F4_0(.din(w_dff_B_ZQ79dYv42_0),.dout(w_dff_B_VgMkRi0F4_0),.clk(gclk));
	jdff dff_B_c1la2naF7_0(.din(w_dff_B_VgMkRi0F4_0),.dout(w_dff_B_c1la2naF7_0),.clk(gclk));
	jdff dff_B_8BlCHmGs9_0(.din(w_dff_B_c1la2naF7_0),.dout(w_dff_B_8BlCHmGs9_0),.clk(gclk));
	jdff dff_B_RTuFv2jB9_0(.din(w_dff_B_8BlCHmGs9_0),.dout(w_dff_B_RTuFv2jB9_0),.clk(gclk));
	jdff dff_B_NMI6u2Vm1_0(.din(w_dff_B_RTuFv2jB9_0),.dout(w_dff_B_NMI6u2Vm1_0),.clk(gclk));
	jdff dff_B_bA1aj1Ja5_0(.din(w_dff_B_NMI6u2Vm1_0),.dout(w_dff_B_bA1aj1Ja5_0),.clk(gclk));
	jdff dff_B_mzhRBYUq3_0(.din(w_dff_B_bA1aj1Ja5_0),.dout(w_dff_B_mzhRBYUq3_0),.clk(gclk));
	jdff dff_B_H5VpTsS30_0(.din(w_dff_B_mzhRBYUq3_0),.dout(w_dff_B_H5VpTsS30_0),.clk(gclk));
	jdff dff_B_bxObI4uX7_0(.din(w_dff_B_H5VpTsS30_0),.dout(w_dff_B_bxObI4uX7_0),.clk(gclk));
	jdff dff_B_RK0TCsYA3_0(.din(w_dff_B_bxObI4uX7_0),.dout(w_dff_B_RK0TCsYA3_0),.clk(gclk));
	jdff dff_B_eqjkK41L5_0(.din(w_dff_B_RK0TCsYA3_0),.dout(w_dff_B_eqjkK41L5_0),.clk(gclk));
	jdff dff_B_n171pwKy9_0(.din(w_dff_B_eqjkK41L5_0),.dout(w_dff_B_n171pwKy9_0),.clk(gclk));
	jdff dff_B_kYJw0nya1_0(.din(w_dff_B_n171pwKy9_0),.dout(w_dff_B_kYJw0nya1_0),.clk(gclk));
	jdff dff_B_Vku1k3N08_0(.din(w_dff_B_kYJw0nya1_0),.dout(w_dff_B_Vku1k3N08_0),.clk(gclk));
	jdff dff_B_6k4dRwQa8_0(.din(w_dff_B_Vku1k3N08_0),.dout(w_dff_B_6k4dRwQa8_0),.clk(gclk));
	jdff dff_B_I7H3BmAH6_0(.din(w_dff_B_6k4dRwQa8_0),.dout(w_dff_B_I7H3BmAH6_0),.clk(gclk));
	jdff dff_B_zsz0bKgE1_0(.din(w_dff_B_I7H3BmAH6_0),.dout(w_dff_B_zsz0bKgE1_0),.clk(gclk));
	jdff dff_B_4k8l3izr5_0(.din(w_dff_B_zsz0bKgE1_0),.dout(w_dff_B_4k8l3izr5_0),.clk(gclk));
	jdff dff_B_5SfkRjzQ9_0(.din(w_dff_B_4k8l3izr5_0),.dout(w_dff_B_5SfkRjzQ9_0),.clk(gclk));
	jdff dff_B_aRzmjmHw2_0(.din(w_dff_B_5SfkRjzQ9_0),.dout(w_dff_B_aRzmjmHw2_0),.clk(gclk));
	jdff dff_B_YBWHNTm40_0(.din(w_dff_B_aRzmjmHw2_0),.dout(w_dff_B_YBWHNTm40_0),.clk(gclk));
	jdff dff_B_3YExAsal2_0(.din(w_dff_B_YBWHNTm40_0),.dout(w_dff_B_3YExAsal2_0),.clk(gclk));
	jdff dff_B_cTy98Or30_0(.din(w_dff_B_3YExAsal2_0),.dout(w_dff_B_cTy98Or30_0),.clk(gclk));
	jdff dff_B_jXru8UAN5_0(.din(w_dff_B_cTy98Or30_0),.dout(w_dff_B_jXru8UAN5_0),.clk(gclk));
	jdff dff_B_j4fPjshF6_0(.din(w_dff_B_jXru8UAN5_0),.dout(w_dff_B_j4fPjshF6_0),.clk(gclk));
	jdff dff_B_BcVUBeY14_0(.din(w_dff_B_j4fPjshF6_0),.dout(w_dff_B_BcVUBeY14_0),.clk(gclk));
	jdff dff_B_nodnidlk9_0(.din(w_dff_B_BcVUBeY14_0),.dout(w_dff_B_nodnidlk9_0),.clk(gclk));
	jdff dff_B_Mo6z9htM5_0(.din(w_dff_B_nodnidlk9_0),.dout(w_dff_B_Mo6z9htM5_0),.clk(gclk));
	jdff dff_B_5lfFUUGb7_0(.din(w_dff_B_Mo6z9htM5_0),.dout(w_dff_B_5lfFUUGb7_0),.clk(gclk));
	jdff dff_B_HNKWwTdp5_0(.din(w_dff_B_5lfFUUGb7_0),.dout(w_dff_B_HNKWwTdp5_0),.clk(gclk));
	jdff dff_B_tgMHmLvg7_0(.din(w_dff_B_HNKWwTdp5_0),.dout(w_dff_B_tgMHmLvg7_0),.clk(gclk));
	jdff dff_B_yGx9XO0y1_0(.din(w_dff_B_tgMHmLvg7_0),.dout(w_dff_B_yGx9XO0y1_0),.clk(gclk));
	jdff dff_B_7wOukHDP7_0(.din(w_dff_B_yGx9XO0y1_0),.dout(w_dff_B_7wOukHDP7_0),.clk(gclk));
	jdff dff_B_3mCMrSM53_0(.din(w_dff_B_7wOukHDP7_0),.dout(w_dff_B_3mCMrSM53_0),.clk(gclk));
	jdff dff_B_EjhPv0Ue1_0(.din(w_dff_B_3mCMrSM53_0),.dout(w_dff_B_EjhPv0Ue1_0),.clk(gclk));
	jdff dff_B_586AmrHn1_0(.din(w_dff_B_EjhPv0Ue1_0),.dout(w_dff_B_586AmrHn1_0),.clk(gclk));
	jdff dff_B_sVeiOpTv3_0(.din(w_dff_B_586AmrHn1_0),.dout(w_dff_B_sVeiOpTv3_0),.clk(gclk));
	jdff dff_B_mHJk5P6P4_0(.din(w_dff_B_sVeiOpTv3_0),.dout(w_dff_B_mHJk5P6P4_0),.clk(gclk));
	jdff dff_B_SQy7amcp8_0(.din(w_dff_B_mHJk5P6P4_0),.dout(w_dff_B_SQy7amcp8_0),.clk(gclk));
	jdff dff_B_JqvLh42k3_0(.din(w_dff_B_SQy7amcp8_0),.dout(w_dff_B_JqvLh42k3_0),.clk(gclk));
	jdff dff_B_kvx9Yotb4_0(.din(w_dff_B_JqvLh42k3_0),.dout(w_dff_B_kvx9Yotb4_0),.clk(gclk));
	jdff dff_B_lvO8LczQ8_0(.din(w_dff_B_kvx9Yotb4_0),.dout(w_dff_B_lvO8LczQ8_0),.clk(gclk));
	jdff dff_B_iXWmVun97_0(.din(w_dff_B_lvO8LczQ8_0),.dout(w_dff_B_iXWmVun97_0),.clk(gclk));
	jdff dff_B_mQHMMDY13_0(.din(w_dff_B_iXWmVun97_0),.dout(w_dff_B_mQHMMDY13_0),.clk(gclk));
	jdff dff_B_VeaFra8e0_0(.din(w_dff_B_mQHMMDY13_0),.dout(w_dff_B_VeaFra8e0_0),.clk(gclk));
	jdff dff_B_1oDJRiut2_0(.din(w_dff_B_VeaFra8e0_0),.dout(w_dff_B_1oDJRiut2_0),.clk(gclk));
	jdff dff_B_JOP3wQKt7_0(.din(w_dff_B_1oDJRiut2_0),.dout(w_dff_B_JOP3wQKt7_0),.clk(gclk));
	jdff dff_B_QO7hosX06_0(.din(w_dff_B_JOP3wQKt7_0),.dout(w_dff_B_QO7hosX06_0),.clk(gclk));
	jdff dff_B_30HJfyvr3_0(.din(w_dff_B_QO7hosX06_0),.dout(w_dff_B_30HJfyvr3_0),.clk(gclk));
	jdff dff_B_t5TBYdXg2_0(.din(w_dff_B_30HJfyvr3_0),.dout(w_dff_B_t5TBYdXg2_0),.clk(gclk));
	jdff dff_B_hiulta0n9_0(.din(w_dff_B_t5TBYdXg2_0),.dout(w_dff_B_hiulta0n9_0),.clk(gclk));
	jdff dff_B_a0ANJVWH8_0(.din(w_dff_B_hiulta0n9_0),.dout(w_dff_B_a0ANJVWH8_0),.clk(gclk));
	jdff dff_B_eQDhJaQr8_0(.din(w_dff_B_a0ANJVWH8_0),.dout(w_dff_B_eQDhJaQr8_0),.clk(gclk));
	jdff dff_B_jblAHUSy8_0(.din(w_dff_B_eQDhJaQr8_0),.dout(w_dff_B_jblAHUSy8_0),.clk(gclk));
	jdff dff_B_TeqD7gin4_0(.din(w_dff_B_jblAHUSy8_0),.dout(w_dff_B_TeqD7gin4_0),.clk(gclk));
	jdff dff_B_h49672xp6_0(.din(w_dff_B_TeqD7gin4_0),.dout(w_dff_B_h49672xp6_0),.clk(gclk));
	jdff dff_B_RPfYOhkB3_0(.din(w_dff_B_h49672xp6_0),.dout(w_dff_B_RPfYOhkB3_0),.clk(gclk));
	jdff dff_B_NGWKogmw0_0(.din(w_dff_B_RPfYOhkB3_0),.dout(w_dff_B_NGWKogmw0_0),.clk(gclk));
	jdff dff_B_Wk4KetGe0_0(.din(w_dff_B_NGWKogmw0_0),.dout(w_dff_B_Wk4KetGe0_0),.clk(gclk));
	jdff dff_B_uTflJdG17_0(.din(w_dff_B_Wk4KetGe0_0),.dout(w_dff_B_uTflJdG17_0),.clk(gclk));
	jdff dff_B_UXItrIjW6_0(.din(w_dff_B_uTflJdG17_0),.dout(w_dff_B_UXItrIjW6_0),.clk(gclk));
	jdff dff_B_EOLcdZNy0_0(.din(w_dff_B_UXItrIjW6_0),.dout(w_dff_B_EOLcdZNy0_0),.clk(gclk));
	jdff dff_B_WiSVbLIf7_0(.din(w_dff_B_EOLcdZNy0_0),.dout(w_dff_B_WiSVbLIf7_0),.clk(gclk));
	jdff dff_B_YSwUJrZg9_0(.din(w_dff_B_WiSVbLIf7_0),.dout(w_dff_B_YSwUJrZg9_0),.clk(gclk));
	jdff dff_B_NDXc5CgD3_0(.din(w_dff_B_YSwUJrZg9_0),.dout(w_dff_B_NDXc5CgD3_0),.clk(gclk));
	jdff dff_B_oQb1CUJZ6_0(.din(w_dff_B_NDXc5CgD3_0),.dout(w_dff_B_oQb1CUJZ6_0),.clk(gclk));
	jdff dff_B_yTiXYGqt9_0(.din(w_dff_B_oQb1CUJZ6_0),.dout(w_dff_B_yTiXYGqt9_0),.clk(gclk));
	jdff dff_B_7QWeiGtI1_0(.din(w_dff_B_yTiXYGqt9_0),.dout(w_dff_B_7QWeiGtI1_0),.clk(gclk));
	jdff dff_B_zVUTpR733_0(.din(w_dff_B_7QWeiGtI1_0),.dout(w_dff_B_zVUTpR733_0),.clk(gclk));
	jdff dff_B_ErcSPY5p9_0(.din(w_dff_B_zVUTpR733_0),.dout(w_dff_B_ErcSPY5p9_0),.clk(gclk));
	jdff dff_B_Lso0hCi86_0(.din(w_dff_B_ErcSPY5p9_0),.dout(w_dff_B_Lso0hCi86_0),.clk(gclk));
	jdff dff_B_oj9BPdGt0_0(.din(w_dff_B_Lso0hCi86_0),.dout(w_dff_B_oj9BPdGt0_0),.clk(gclk));
	jdff dff_B_pETxBHAB6_0(.din(w_dff_B_oj9BPdGt0_0),.dout(w_dff_B_pETxBHAB6_0),.clk(gclk));
	jdff dff_B_9oeEatje8_0(.din(w_dff_B_pETxBHAB6_0),.dout(w_dff_B_9oeEatje8_0),.clk(gclk));
	jdff dff_B_CDVe9Lni1_0(.din(w_dff_B_9oeEatje8_0),.dout(w_dff_B_CDVe9Lni1_0),.clk(gclk));
	jdff dff_B_5AJeGuG53_0(.din(w_dff_B_CDVe9Lni1_0),.dout(w_dff_B_5AJeGuG53_0),.clk(gclk));
	jdff dff_B_mD9JOMR65_0(.din(w_dff_B_5AJeGuG53_0),.dout(w_dff_B_mD9JOMR65_0),.clk(gclk));
	jdff dff_B_tAMSHKno7_0(.din(w_dff_B_mD9JOMR65_0),.dout(w_dff_B_tAMSHKno7_0),.clk(gclk));
	jdff dff_B_FE4voPy93_0(.din(w_dff_B_tAMSHKno7_0),.dout(w_dff_B_FE4voPy93_0),.clk(gclk));
	jdff dff_B_3BlTFiyi6_0(.din(w_dff_B_FE4voPy93_0),.dout(w_dff_B_3BlTFiyi6_0),.clk(gclk));
	jdff dff_B_qlKuB7PC5_0(.din(w_dff_B_3BlTFiyi6_0),.dout(w_dff_B_qlKuB7PC5_0),.clk(gclk));
	jdff dff_B_w0Xu8MMm0_0(.din(w_dff_B_qlKuB7PC5_0),.dout(w_dff_B_w0Xu8MMm0_0),.clk(gclk));
	jdff dff_B_yYEBiORo3_0(.din(w_dff_B_w0Xu8MMm0_0),.dout(w_dff_B_yYEBiORo3_0),.clk(gclk));
	jdff dff_B_niFMbCQe5_0(.din(w_dff_B_yYEBiORo3_0),.dout(w_dff_B_niFMbCQe5_0),.clk(gclk));
	jdff dff_B_xlvf58vQ1_1(.din(n1122),.dout(w_dff_B_xlvf58vQ1_1),.clk(gclk));
	jdff dff_B_TTyx2DR68_1(.din(w_dff_B_xlvf58vQ1_1),.dout(w_dff_B_TTyx2DR68_1),.clk(gclk));
	jdff dff_B_adBEQpWH4_1(.din(w_dff_B_TTyx2DR68_1),.dout(w_dff_B_adBEQpWH4_1),.clk(gclk));
	jdff dff_B_T9SsQlCm4_1(.din(w_dff_B_adBEQpWH4_1),.dout(w_dff_B_T9SsQlCm4_1),.clk(gclk));
	jdff dff_B_YZTMGZrP2_1(.din(w_dff_B_T9SsQlCm4_1),.dout(w_dff_B_YZTMGZrP2_1),.clk(gclk));
	jdff dff_B_aqGz3X2U2_1(.din(w_dff_B_YZTMGZrP2_1),.dout(w_dff_B_aqGz3X2U2_1),.clk(gclk));
	jdff dff_B_1T0xIEXj0_1(.din(w_dff_B_aqGz3X2U2_1),.dout(w_dff_B_1T0xIEXj0_1),.clk(gclk));
	jdff dff_B_j4Qr55xX6_1(.din(w_dff_B_1T0xIEXj0_1),.dout(w_dff_B_j4Qr55xX6_1),.clk(gclk));
	jdff dff_B_X9ys2ipn3_1(.din(w_dff_B_j4Qr55xX6_1),.dout(w_dff_B_X9ys2ipn3_1),.clk(gclk));
	jdff dff_B_MZTRSDSN5_1(.din(w_dff_B_X9ys2ipn3_1),.dout(w_dff_B_MZTRSDSN5_1),.clk(gclk));
	jdff dff_B_wKjbdVkK8_1(.din(w_dff_B_MZTRSDSN5_1),.dout(w_dff_B_wKjbdVkK8_1),.clk(gclk));
	jdff dff_B_K65fyst61_1(.din(w_dff_B_wKjbdVkK8_1),.dout(w_dff_B_K65fyst61_1),.clk(gclk));
	jdff dff_B_naMSC7bd7_1(.din(w_dff_B_K65fyst61_1),.dout(w_dff_B_naMSC7bd7_1),.clk(gclk));
	jdff dff_B_mFpoFg8w0_1(.din(w_dff_B_naMSC7bd7_1),.dout(w_dff_B_mFpoFg8w0_1),.clk(gclk));
	jdff dff_B_ZNTO9vlu6_1(.din(w_dff_B_mFpoFg8w0_1),.dout(w_dff_B_ZNTO9vlu6_1),.clk(gclk));
	jdff dff_B_JiBjjnmS5_1(.din(w_dff_B_ZNTO9vlu6_1),.dout(w_dff_B_JiBjjnmS5_1),.clk(gclk));
	jdff dff_B_PGJdhn066_1(.din(w_dff_B_JiBjjnmS5_1),.dout(w_dff_B_PGJdhn066_1),.clk(gclk));
	jdff dff_B_g9jBuuxl1_1(.din(w_dff_B_PGJdhn066_1),.dout(w_dff_B_g9jBuuxl1_1),.clk(gclk));
	jdff dff_B_IORxOFa64_1(.din(w_dff_B_g9jBuuxl1_1),.dout(w_dff_B_IORxOFa64_1),.clk(gclk));
	jdff dff_B_EkBj8YK36_1(.din(w_dff_B_IORxOFa64_1),.dout(w_dff_B_EkBj8YK36_1),.clk(gclk));
	jdff dff_B_JlYTub2w1_1(.din(w_dff_B_EkBj8YK36_1),.dout(w_dff_B_JlYTub2w1_1),.clk(gclk));
	jdff dff_B_tTXzqfwP3_1(.din(w_dff_B_JlYTub2w1_1),.dout(w_dff_B_tTXzqfwP3_1),.clk(gclk));
	jdff dff_B_YCcPspPj9_1(.din(w_dff_B_tTXzqfwP3_1),.dout(w_dff_B_YCcPspPj9_1),.clk(gclk));
	jdff dff_B_anQ1ieDQ0_1(.din(w_dff_B_YCcPspPj9_1),.dout(w_dff_B_anQ1ieDQ0_1),.clk(gclk));
	jdff dff_B_zHkaOqPY2_1(.din(w_dff_B_anQ1ieDQ0_1),.dout(w_dff_B_zHkaOqPY2_1),.clk(gclk));
	jdff dff_B_xcwH6Zn87_1(.din(w_dff_B_zHkaOqPY2_1),.dout(w_dff_B_xcwH6Zn87_1),.clk(gclk));
	jdff dff_B_qRV4VmrB4_1(.din(w_dff_B_xcwH6Zn87_1),.dout(w_dff_B_qRV4VmrB4_1),.clk(gclk));
	jdff dff_B_7AeT5CL99_1(.din(w_dff_B_qRV4VmrB4_1),.dout(w_dff_B_7AeT5CL99_1),.clk(gclk));
	jdff dff_B_wnJwFzY71_1(.din(w_dff_B_7AeT5CL99_1),.dout(w_dff_B_wnJwFzY71_1),.clk(gclk));
	jdff dff_B_Eli4ENS49_1(.din(w_dff_B_wnJwFzY71_1),.dout(w_dff_B_Eli4ENS49_1),.clk(gclk));
	jdff dff_B_8z4rXfXo1_1(.din(w_dff_B_Eli4ENS49_1),.dout(w_dff_B_8z4rXfXo1_1),.clk(gclk));
	jdff dff_B_Q71ONbxz9_1(.din(w_dff_B_8z4rXfXo1_1),.dout(w_dff_B_Q71ONbxz9_1),.clk(gclk));
	jdff dff_B_so9NQCV50_1(.din(w_dff_B_Q71ONbxz9_1),.dout(w_dff_B_so9NQCV50_1),.clk(gclk));
	jdff dff_B_qF4M63Kt9_1(.din(w_dff_B_so9NQCV50_1),.dout(w_dff_B_qF4M63Kt9_1),.clk(gclk));
	jdff dff_B_WRQBdW015_1(.din(w_dff_B_qF4M63Kt9_1),.dout(w_dff_B_WRQBdW015_1),.clk(gclk));
	jdff dff_B_dpIq37uP5_1(.din(w_dff_B_WRQBdW015_1),.dout(w_dff_B_dpIq37uP5_1),.clk(gclk));
	jdff dff_B_n7rxVgFO2_1(.din(w_dff_B_dpIq37uP5_1),.dout(w_dff_B_n7rxVgFO2_1),.clk(gclk));
	jdff dff_B_EKVtwnh58_1(.din(w_dff_B_n7rxVgFO2_1),.dout(w_dff_B_EKVtwnh58_1),.clk(gclk));
	jdff dff_B_RlNahTF76_1(.din(w_dff_B_EKVtwnh58_1),.dout(w_dff_B_RlNahTF76_1),.clk(gclk));
	jdff dff_B_J8BvEfSI5_1(.din(w_dff_B_RlNahTF76_1),.dout(w_dff_B_J8BvEfSI5_1),.clk(gclk));
	jdff dff_B_MyWIFJO38_1(.din(w_dff_B_J8BvEfSI5_1),.dout(w_dff_B_MyWIFJO38_1),.clk(gclk));
	jdff dff_B_nr4Ulwcs3_1(.din(w_dff_B_MyWIFJO38_1),.dout(w_dff_B_nr4Ulwcs3_1),.clk(gclk));
	jdff dff_B_CD4EsmfM2_1(.din(w_dff_B_nr4Ulwcs3_1),.dout(w_dff_B_CD4EsmfM2_1),.clk(gclk));
	jdff dff_B_VZOseP6H2_1(.din(w_dff_B_CD4EsmfM2_1),.dout(w_dff_B_VZOseP6H2_1),.clk(gclk));
	jdff dff_B_xH6WR0Bc1_1(.din(w_dff_B_VZOseP6H2_1),.dout(w_dff_B_xH6WR0Bc1_1),.clk(gclk));
	jdff dff_B_PXmMgz7r5_1(.din(w_dff_B_xH6WR0Bc1_1),.dout(w_dff_B_PXmMgz7r5_1),.clk(gclk));
	jdff dff_B_B8ucmhgy9_1(.din(w_dff_B_PXmMgz7r5_1),.dout(w_dff_B_B8ucmhgy9_1),.clk(gclk));
	jdff dff_B_kSGBWEoK7_1(.din(w_dff_B_B8ucmhgy9_1),.dout(w_dff_B_kSGBWEoK7_1),.clk(gclk));
	jdff dff_B_8FwmaDCC8_1(.din(w_dff_B_kSGBWEoK7_1),.dout(w_dff_B_8FwmaDCC8_1),.clk(gclk));
	jdff dff_B_yHBsplJU6_1(.din(w_dff_B_8FwmaDCC8_1),.dout(w_dff_B_yHBsplJU6_1),.clk(gclk));
	jdff dff_B_lEUKQ5Jh8_1(.din(w_dff_B_yHBsplJU6_1),.dout(w_dff_B_lEUKQ5Jh8_1),.clk(gclk));
	jdff dff_B_GfxfQfyG5_1(.din(w_dff_B_lEUKQ5Jh8_1),.dout(w_dff_B_GfxfQfyG5_1),.clk(gclk));
	jdff dff_B_8nnEb4cf0_1(.din(w_dff_B_GfxfQfyG5_1),.dout(w_dff_B_8nnEb4cf0_1),.clk(gclk));
	jdff dff_B_0pJFpHVi2_1(.din(w_dff_B_8nnEb4cf0_1),.dout(w_dff_B_0pJFpHVi2_1),.clk(gclk));
	jdff dff_B_V243fT3F8_1(.din(w_dff_B_0pJFpHVi2_1),.dout(w_dff_B_V243fT3F8_1),.clk(gclk));
	jdff dff_B_H85nIkPZ7_1(.din(w_dff_B_V243fT3F8_1),.dout(w_dff_B_H85nIkPZ7_1),.clk(gclk));
	jdff dff_B_mBuljhDl0_1(.din(w_dff_B_H85nIkPZ7_1),.dout(w_dff_B_mBuljhDl0_1),.clk(gclk));
	jdff dff_B_EPJKOdEc2_1(.din(w_dff_B_mBuljhDl0_1),.dout(w_dff_B_EPJKOdEc2_1),.clk(gclk));
	jdff dff_B_25L9GQSA6_1(.din(w_dff_B_EPJKOdEc2_1),.dout(w_dff_B_25L9GQSA6_1),.clk(gclk));
	jdff dff_B_35sVY74G7_1(.din(w_dff_B_25L9GQSA6_1),.dout(w_dff_B_35sVY74G7_1),.clk(gclk));
	jdff dff_B_YzfdV7da7_1(.din(w_dff_B_35sVY74G7_1),.dout(w_dff_B_YzfdV7da7_1),.clk(gclk));
	jdff dff_B_md59xA725_1(.din(w_dff_B_YzfdV7da7_1),.dout(w_dff_B_md59xA725_1),.clk(gclk));
	jdff dff_B_U6lud0nQ2_1(.din(w_dff_B_md59xA725_1),.dout(w_dff_B_U6lud0nQ2_1),.clk(gclk));
	jdff dff_B_Q0IpHpA16_1(.din(w_dff_B_U6lud0nQ2_1),.dout(w_dff_B_Q0IpHpA16_1),.clk(gclk));
	jdff dff_B_hDsqDcpX3_1(.din(w_dff_B_Q0IpHpA16_1),.dout(w_dff_B_hDsqDcpX3_1),.clk(gclk));
	jdff dff_B_56ZfvXFK9_1(.din(w_dff_B_hDsqDcpX3_1),.dout(w_dff_B_56ZfvXFK9_1),.clk(gclk));
	jdff dff_B_cbNCLpXx7_1(.din(w_dff_B_56ZfvXFK9_1),.dout(w_dff_B_cbNCLpXx7_1),.clk(gclk));
	jdff dff_B_wiLcXbuD1_1(.din(w_dff_B_cbNCLpXx7_1),.dout(w_dff_B_wiLcXbuD1_1),.clk(gclk));
	jdff dff_B_wOYgkfWA2_1(.din(w_dff_B_wiLcXbuD1_1),.dout(w_dff_B_wOYgkfWA2_1),.clk(gclk));
	jdff dff_B_VenL9k034_1(.din(w_dff_B_wOYgkfWA2_1),.dout(w_dff_B_VenL9k034_1),.clk(gclk));
	jdff dff_B_adRC1Spb7_1(.din(w_dff_B_VenL9k034_1),.dout(w_dff_B_adRC1Spb7_1),.clk(gclk));
	jdff dff_B_HWwsSvMW8_1(.din(w_dff_B_adRC1Spb7_1),.dout(w_dff_B_HWwsSvMW8_1),.clk(gclk));
	jdff dff_B_yH7bPvti5_1(.din(w_dff_B_HWwsSvMW8_1),.dout(w_dff_B_yH7bPvti5_1),.clk(gclk));
	jdff dff_B_teslDa011_1(.din(w_dff_B_yH7bPvti5_1),.dout(w_dff_B_teslDa011_1),.clk(gclk));
	jdff dff_B_z5Xic96G8_1(.din(w_dff_B_teslDa011_1),.dout(w_dff_B_z5Xic96G8_1),.clk(gclk));
	jdff dff_B_ZdRgUDh58_1(.din(w_dff_B_z5Xic96G8_1),.dout(w_dff_B_ZdRgUDh58_1),.clk(gclk));
	jdff dff_B_YOC3YxSe5_1(.din(w_dff_B_ZdRgUDh58_1),.dout(w_dff_B_YOC3YxSe5_1),.clk(gclk));
	jdff dff_B_9Oysk1De1_1(.din(w_dff_B_YOC3YxSe5_1),.dout(w_dff_B_9Oysk1De1_1),.clk(gclk));
	jdff dff_B_svYgorby7_1(.din(w_dff_B_9Oysk1De1_1),.dout(w_dff_B_svYgorby7_1),.clk(gclk));
	jdff dff_B_orUwcZHc5_1(.din(w_dff_B_svYgorby7_1),.dout(w_dff_B_orUwcZHc5_1),.clk(gclk));
	jdff dff_B_bZOTdtDJ1_1(.din(w_dff_B_orUwcZHc5_1),.dout(w_dff_B_bZOTdtDJ1_1),.clk(gclk));
	jdff dff_B_E0o0jsJD4_1(.din(w_dff_B_bZOTdtDJ1_1),.dout(w_dff_B_E0o0jsJD4_1),.clk(gclk));
	jdff dff_B_7Xb5Yn1W7_1(.din(w_dff_B_E0o0jsJD4_1),.dout(w_dff_B_7Xb5Yn1W7_1),.clk(gclk));
	jdff dff_B_qfEGJUMP1_1(.din(w_dff_B_7Xb5Yn1W7_1),.dout(w_dff_B_qfEGJUMP1_1),.clk(gclk));
	jdff dff_B_uaPWsuno6_1(.din(w_dff_B_qfEGJUMP1_1),.dout(w_dff_B_uaPWsuno6_1),.clk(gclk));
	jdff dff_B_PTdKFq1Z2_1(.din(w_dff_B_uaPWsuno6_1),.dout(w_dff_B_PTdKFq1Z2_1),.clk(gclk));
	jdff dff_B_sE6Z9dCs6_1(.din(w_dff_B_PTdKFq1Z2_1),.dout(w_dff_B_sE6Z9dCs6_1),.clk(gclk));
	jdff dff_B_vvcFx5Je0_1(.din(w_dff_B_sE6Z9dCs6_1),.dout(w_dff_B_vvcFx5Je0_1),.clk(gclk));
	jdff dff_B_SLYAROsV1_1(.din(w_dff_B_vvcFx5Je0_1),.dout(w_dff_B_SLYAROsV1_1),.clk(gclk));
	jdff dff_B_meIXkeyV2_1(.din(w_dff_B_SLYAROsV1_1),.dout(w_dff_B_meIXkeyV2_1),.clk(gclk));
	jdff dff_B_A7VceNDg4_1(.din(w_dff_B_meIXkeyV2_1),.dout(w_dff_B_A7VceNDg4_1),.clk(gclk));
	jdff dff_B_GzoORZZi1_1(.din(w_dff_B_A7VceNDg4_1),.dout(w_dff_B_GzoORZZi1_1),.clk(gclk));
	jdff dff_B_n6pIe9V38_1(.din(w_dff_B_GzoORZZi1_1),.dout(w_dff_B_n6pIe9V38_1),.clk(gclk));
	jdff dff_B_mlFwG6D14_1(.din(w_dff_B_n6pIe9V38_1),.dout(w_dff_B_mlFwG6D14_1),.clk(gclk));
	jdff dff_B_UVzWyeGm8_1(.din(w_dff_B_mlFwG6D14_1),.dout(w_dff_B_UVzWyeGm8_1),.clk(gclk));
	jdff dff_B_i0Hw55dn2_1(.din(w_dff_B_UVzWyeGm8_1),.dout(w_dff_B_i0Hw55dn2_1),.clk(gclk));
	jdff dff_B_1K9eH9dv7_1(.din(w_dff_B_i0Hw55dn2_1),.dout(w_dff_B_1K9eH9dv7_1),.clk(gclk));
	jdff dff_B_XjxpKpjw4_1(.din(w_dff_B_1K9eH9dv7_1),.dout(w_dff_B_XjxpKpjw4_1),.clk(gclk));
	jdff dff_B_9QPXdl4i0_1(.din(w_dff_B_XjxpKpjw4_1),.dout(w_dff_B_9QPXdl4i0_1),.clk(gclk));
	jdff dff_B_NocTdLFw2_1(.din(w_dff_B_9QPXdl4i0_1),.dout(w_dff_B_NocTdLFw2_1),.clk(gclk));
	jdff dff_B_tmehyRQF0_1(.din(w_dff_B_NocTdLFw2_1),.dout(w_dff_B_tmehyRQF0_1),.clk(gclk));
	jdff dff_B_jvRcFlPW4_1(.din(w_dff_B_tmehyRQF0_1),.dout(w_dff_B_jvRcFlPW4_1),.clk(gclk));
	jdff dff_B_GpQlljSz4_1(.din(w_dff_B_jvRcFlPW4_1),.dout(w_dff_B_GpQlljSz4_1),.clk(gclk));
	jdff dff_B_DJBJuvdo1_1(.din(w_dff_B_GpQlljSz4_1),.dout(w_dff_B_DJBJuvdo1_1),.clk(gclk));
	jdff dff_B_RVAyDpQT0_1(.din(w_dff_B_DJBJuvdo1_1),.dout(w_dff_B_RVAyDpQT0_1),.clk(gclk));
	jdff dff_B_6tPjsgCX7_1(.din(w_dff_B_RVAyDpQT0_1),.dout(w_dff_B_6tPjsgCX7_1),.clk(gclk));
	jdff dff_B_F9qXrrgj8_1(.din(w_dff_B_6tPjsgCX7_1),.dout(w_dff_B_F9qXrrgj8_1),.clk(gclk));
	jdff dff_B_rjefnjaQ8_1(.din(w_dff_B_F9qXrrgj8_1),.dout(w_dff_B_rjefnjaQ8_1),.clk(gclk));
	jdff dff_B_gFjkcwoc6_1(.din(w_dff_B_rjefnjaQ8_1),.dout(w_dff_B_gFjkcwoc6_1),.clk(gclk));
	jdff dff_B_QTmH9Rgb2_1(.din(w_dff_B_gFjkcwoc6_1),.dout(w_dff_B_QTmH9Rgb2_1),.clk(gclk));
	jdff dff_B_FNn87wEo1_1(.din(w_dff_B_QTmH9Rgb2_1),.dout(w_dff_B_FNn87wEo1_1),.clk(gclk));
	jdff dff_B_0wPVGqB70_1(.din(w_dff_B_FNn87wEo1_1),.dout(w_dff_B_0wPVGqB70_1),.clk(gclk));
	jdff dff_B_wyrOMR8X2_1(.din(w_dff_B_0wPVGqB70_1),.dout(w_dff_B_wyrOMR8X2_1),.clk(gclk));
	jdff dff_B_0ShiLpUC5_1(.din(w_dff_B_wyrOMR8X2_1),.dout(w_dff_B_0ShiLpUC5_1),.clk(gclk));
	jdff dff_B_CPSFP8od5_1(.din(w_dff_B_0ShiLpUC5_1),.dout(w_dff_B_CPSFP8od5_1),.clk(gclk));
	jdff dff_B_XFU1OhDk3_1(.din(w_dff_B_CPSFP8od5_1),.dout(w_dff_B_XFU1OhDk3_1),.clk(gclk));
	jdff dff_B_7EmC7Be77_1(.din(w_dff_B_XFU1OhDk3_1),.dout(w_dff_B_7EmC7Be77_1),.clk(gclk));
	jdff dff_B_5lYm1sbU4_1(.din(w_dff_B_7EmC7Be77_1),.dout(w_dff_B_5lYm1sbU4_1),.clk(gclk));
	jdff dff_B_T057vtT76_1(.din(w_dff_B_5lYm1sbU4_1),.dout(w_dff_B_T057vtT76_1),.clk(gclk));
	jdff dff_B_v0qgbIni3_1(.din(w_dff_B_T057vtT76_1),.dout(w_dff_B_v0qgbIni3_1),.clk(gclk));
	jdff dff_B_OXDQLYQM0_1(.din(w_dff_B_v0qgbIni3_1),.dout(w_dff_B_OXDQLYQM0_1),.clk(gclk));
	jdff dff_B_R2r5urwW2_1(.din(w_dff_B_OXDQLYQM0_1),.dout(w_dff_B_R2r5urwW2_1),.clk(gclk));
	jdff dff_B_LkmyUViD3_1(.din(w_dff_B_R2r5urwW2_1),.dout(w_dff_B_LkmyUViD3_1),.clk(gclk));
	jdff dff_B_ihlUGtXO8_0(.din(n1123),.dout(w_dff_B_ihlUGtXO8_0),.clk(gclk));
	jdff dff_B_NkOGzgBJ9_0(.din(w_dff_B_ihlUGtXO8_0),.dout(w_dff_B_NkOGzgBJ9_0),.clk(gclk));
	jdff dff_B_p09xVsVY1_0(.din(w_dff_B_NkOGzgBJ9_0),.dout(w_dff_B_p09xVsVY1_0),.clk(gclk));
	jdff dff_B_0x2a8bzk6_0(.din(w_dff_B_p09xVsVY1_0),.dout(w_dff_B_0x2a8bzk6_0),.clk(gclk));
	jdff dff_B_2D9RksV12_0(.din(w_dff_B_0x2a8bzk6_0),.dout(w_dff_B_2D9RksV12_0),.clk(gclk));
	jdff dff_B_Jl3mnOkw2_0(.din(w_dff_B_2D9RksV12_0),.dout(w_dff_B_Jl3mnOkw2_0),.clk(gclk));
	jdff dff_B_XjypEmla5_0(.din(w_dff_B_Jl3mnOkw2_0),.dout(w_dff_B_XjypEmla5_0),.clk(gclk));
	jdff dff_B_tKy7lzpq7_0(.din(w_dff_B_XjypEmla5_0),.dout(w_dff_B_tKy7lzpq7_0),.clk(gclk));
	jdff dff_B_83FZHCaX8_0(.din(w_dff_B_tKy7lzpq7_0),.dout(w_dff_B_83FZHCaX8_0),.clk(gclk));
	jdff dff_B_5bmOblIn6_0(.din(w_dff_B_83FZHCaX8_0),.dout(w_dff_B_5bmOblIn6_0),.clk(gclk));
	jdff dff_B_nYDAu46E0_0(.din(w_dff_B_5bmOblIn6_0),.dout(w_dff_B_nYDAu46E0_0),.clk(gclk));
	jdff dff_B_IoIH5eRg8_0(.din(w_dff_B_nYDAu46E0_0),.dout(w_dff_B_IoIH5eRg8_0),.clk(gclk));
	jdff dff_B_sVYv0QnC7_0(.din(w_dff_B_IoIH5eRg8_0),.dout(w_dff_B_sVYv0QnC7_0),.clk(gclk));
	jdff dff_B_rLBMJeiD5_0(.din(w_dff_B_sVYv0QnC7_0),.dout(w_dff_B_rLBMJeiD5_0),.clk(gclk));
	jdff dff_B_FQUOScfA3_0(.din(w_dff_B_rLBMJeiD5_0),.dout(w_dff_B_FQUOScfA3_0),.clk(gclk));
	jdff dff_B_s0pUiaCh4_0(.din(w_dff_B_FQUOScfA3_0),.dout(w_dff_B_s0pUiaCh4_0),.clk(gclk));
	jdff dff_B_wUX6OwdT6_0(.din(w_dff_B_s0pUiaCh4_0),.dout(w_dff_B_wUX6OwdT6_0),.clk(gclk));
	jdff dff_B_mBlZF68n9_0(.din(w_dff_B_wUX6OwdT6_0),.dout(w_dff_B_mBlZF68n9_0),.clk(gclk));
	jdff dff_B_xqzbBVX38_0(.din(w_dff_B_mBlZF68n9_0),.dout(w_dff_B_xqzbBVX38_0),.clk(gclk));
	jdff dff_B_0I10pM2n0_0(.din(w_dff_B_xqzbBVX38_0),.dout(w_dff_B_0I10pM2n0_0),.clk(gclk));
	jdff dff_B_mhdMjQlu8_0(.din(w_dff_B_0I10pM2n0_0),.dout(w_dff_B_mhdMjQlu8_0),.clk(gclk));
	jdff dff_B_a4Wax3J05_0(.din(w_dff_B_mhdMjQlu8_0),.dout(w_dff_B_a4Wax3J05_0),.clk(gclk));
	jdff dff_B_tTbJZN4b2_0(.din(w_dff_B_a4Wax3J05_0),.dout(w_dff_B_tTbJZN4b2_0),.clk(gclk));
	jdff dff_B_5grlECEy6_0(.din(w_dff_B_tTbJZN4b2_0),.dout(w_dff_B_5grlECEy6_0),.clk(gclk));
	jdff dff_B_9ahz7QzT3_0(.din(w_dff_B_5grlECEy6_0),.dout(w_dff_B_9ahz7QzT3_0),.clk(gclk));
	jdff dff_B_qpkKpWaP2_0(.din(w_dff_B_9ahz7QzT3_0),.dout(w_dff_B_qpkKpWaP2_0),.clk(gclk));
	jdff dff_B_vEA4YN229_0(.din(w_dff_B_qpkKpWaP2_0),.dout(w_dff_B_vEA4YN229_0),.clk(gclk));
	jdff dff_B_SfiivDl58_0(.din(w_dff_B_vEA4YN229_0),.dout(w_dff_B_SfiivDl58_0),.clk(gclk));
	jdff dff_B_XhnCNJfe9_0(.din(w_dff_B_SfiivDl58_0),.dout(w_dff_B_XhnCNJfe9_0),.clk(gclk));
	jdff dff_B_Yae4X7aV0_0(.din(w_dff_B_XhnCNJfe9_0),.dout(w_dff_B_Yae4X7aV0_0),.clk(gclk));
	jdff dff_B_Lmsr50hD4_0(.din(w_dff_B_Yae4X7aV0_0),.dout(w_dff_B_Lmsr50hD4_0),.clk(gclk));
	jdff dff_B_o0rAgbcO7_0(.din(w_dff_B_Lmsr50hD4_0),.dout(w_dff_B_o0rAgbcO7_0),.clk(gclk));
	jdff dff_B_sMgtRZuH6_0(.din(w_dff_B_o0rAgbcO7_0),.dout(w_dff_B_sMgtRZuH6_0),.clk(gclk));
	jdff dff_B_BwpORKUs8_0(.din(w_dff_B_sMgtRZuH6_0),.dout(w_dff_B_BwpORKUs8_0),.clk(gclk));
	jdff dff_B_1Ba3HmeU4_0(.din(w_dff_B_BwpORKUs8_0),.dout(w_dff_B_1Ba3HmeU4_0),.clk(gclk));
	jdff dff_B_Tqt3ylUe4_0(.din(w_dff_B_1Ba3HmeU4_0),.dout(w_dff_B_Tqt3ylUe4_0),.clk(gclk));
	jdff dff_B_O4Aey8852_0(.din(w_dff_B_Tqt3ylUe4_0),.dout(w_dff_B_O4Aey8852_0),.clk(gclk));
	jdff dff_B_OaP1z9Xp8_0(.din(w_dff_B_O4Aey8852_0),.dout(w_dff_B_OaP1z9Xp8_0),.clk(gclk));
	jdff dff_B_s9IXb4lF0_0(.din(w_dff_B_OaP1z9Xp8_0),.dout(w_dff_B_s9IXb4lF0_0),.clk(gclk));
	jdff dff_B_Y4AE17Yg8_0(.din(w_dff_B_s9IXb4lF0_0),.dout(w_dff_B_Y4AE17Yg8_0),.clk(gclk));
	jdff dff_B_zj0fm7Vz6_0(.din(w_dff_B_Y4AE17Yg8_0),.dout(w_dff_B_zj0fm7Vz6_0),.clk(gclk));
	jdff dff_B_TtMNznxo2_0(.din(w_dff_B_zj0fm7Vz6_0),.dout(w_dff_B_TtMNznxo2_0),.clk(gclk));
	jdff dff_B_LIHsrAjx8_0(.din(w_dff_B_TtMNznxo2_0),.dout(w_dff_B_LIHsrAjx8_0),.clk(gclk));
	jdff dff_B_VzGHiERh0_0(.din(w_dff_B_LIHsrAjx8_0),.dout(w_dff_B_VzGHiERh0_0),.clk(gclk));
	jdff dff_B_7h1ZVCIE7_0(.din(w_dff_B_VzGHiERh0_0),.dout(w_dff_B_7h1ZVCIE7_0),.clk(gclk));
	jdff dff_B_63WDjKph8_0(.din(w_dff_B_7h1ZVCIE7_0),.dout(w_dff_B_63WDjKph8_0),.clk(gclk));
	jdff dff_B_OFGWtzhD9_0(.din(w_dff_B_63WDjKph8_0),.dout(w_dff_B_OFGWtzhD9_0),.clk(gclk));
	jdff dff_B_x9UyrlZa1_0(.din(w_dff_B_OFGWtzhD9_0),.dout(w_dff_B_x9UyrlZa1_0),.clk(gclk));
	jdff dff_B_MjH3lbxJ4_0(.din(w_dff_B_x9UyrlZa1_0),.dout(w_dff_B_MjH3lbxJ4_0),.clk(gclk));
	jdff dff_B_k478VyFo3_0(.din(w_dff_B_MjH3lbxJ4_0),.dout(w_dff_B_k478VyFo3_0),.clk(gclk));
	jdff dff_B_qz2r93Fu4_0(.din(w_dff_B_k478VyFo3_0),.dout(w_dff_B_qz2r93Fu4_0),.clk(gclk));
	jdff dff_B_69GanfH85_0(.din(w_dff_B_qz2r93Fu4_0),.dout(w_dff_B_69GanfH85_0),.clk(gclk));
	jdff dff_B_lEHpw3uC9_0(.din(w_dff_B_69GanfH85_0),.dout(w_dff_B_lEHpw3uC9_0),.clk(gclk));
	jdff dff_B_MBR4Bqag1_0(.din(w_dff_B_lEHpw3uC9_0),.dout(w_dff_B_MBR4Bqag1_0),.clk(gclk));
	jdff dff_B_uMesbX2l8_0(.din(w_dff_B_MBR4Bqag1_0),.dout(w_dff_B_uMesbX2l8_0),.clk(gclk));
	jdff dff_B_lcmLEtLN4_0(.din(w_dff_B_uMesbX2l8_0),.dout(w_dff_B_lcmLEtLN4_0),.clk(gclk));
	jdff dff_B_1cJYQPYZ4_0(.din(w_dff_B_lcmLEtLN4_0),.dout(w_dff_B_1cJYQPYZ4_0),.clk(gclk));
	jdff dff_B_lbqFqpCt7_0(.din(w_dff_B_1cJYQPYZ4_0),.dout(w_dff_B_lbqFqpCt7_0),.clk(gclk));
	jdff dff_B_voKNSnEL7_0(.din(w_dff_B_lbqFqpCt7_0),.dout(w_dff_B_voKNSnEL7_0),.clk(gclk));
	jdff dff_B_MeW3wqjq1_0(.din(w_dff_B_voKNSnEL7_0),.dout(w_dff_B_MeW3wqjq1_0),.clk(gclk));
	jdff dff_B_Zr6U3pSh6_0(.din(w_dff_B_MeW3wqjq1_0),.dout(w_dff_B_Zr6U3pSh6_0),.clk(gclk));
	jdff dff_B_ZpdeBxHt9_0(.din(w_dff_B_Zr6U3pSh6_0),.dout(w_dff_B_ZpdeBxHt9_0),.clk(gclk));
	jdff dff_B_JNmQcTox4_0(.din(w_dff_B_ZpdeBxHt9_0),.dout(w_dff_B_JNmQcTox4_0),.clk(gclk));
	jdff dff_B_wccacKVF9_0(.din(w_dff_B_JNmQcTox4_0),.dout(w_dff_B_wccacKVF9_0),.clk(gclk));
	jdff dff_B_kj4qZUcD2_0(.din(w_dff_B_wccacKVF9_0),.dout(w_dff_B_kj4qZUcD2_0),.clk(gclk));
	jdff dff_B_87nUqp621_0(.din(w_dff_B_kj4qZUcD2_0),.dout(w_dff_B_87nUqp621_0),.clk(gclk));
	jdff dff_B_tg6XyGZ03_0(.din(w_dff_B_87nUqp621_0),.dout(w_dff_B_tg6XyGZ03_0),.clk(gclk));
	jdff dff_B_SHyb2bd79_0(.din(w_dff_B_tg6XyGZ03_0),.dout(w_dff_B_SHyb2bd79_0),.clk(gclk));
	jdff dff_B_Yt7Y0Cxy4_0(.din(w_dff_B_SHyb2bd79_0),.dout(w_dff_B_Yt7Y0Cxy4_0),.clk(gclk));
	jdff dff_B_rfBshHXY2_0(.din(w_dff_B_Yt7Y0Cxy4_0),.dout(w_dff_B_rfBshHXY2_0),.clk(gclk));
	jdff dff_B_Mr0V7Xre1_0(.din(w_dff_B_rfBshHXY2_0),.dout(w_dff_B_Mr0V7Xre1_0),.clk(gclk));
	jdff dff_B_NDj991vz6_0(.din(w_dff_B_Mr0V7Xre1_0),.dout(w_dff_B_NDj991vz6_0),.clk(gclk));
	jdff dff_B_dGrQ0FDj8_0(.din(w_dff_B_NDj991vz6_0),.dout(w_dff_B_dGrQ0FDj8_0),.clk(gclk));
	jdff dff_B_E5uY0JtH1_0(.din(w_dff_B_dGrQ0FDj8_0),.dout(w_dff_B_E5uY0JtH1_0),.clk(gclk));
	jdff dff_B_ylzSd0Ly2_0(.din(w_dff_B_E5uY0JtH1_0),.dout(w_dff_B_ylzSd0Ly2_0),.clk(gclk));
	jdff dff_B_PJUHQmdO7_0(.din(w_dff_B_ylzSd0Ly2_0),.dout(w_dff_B_PJUHQmdO7_0),.clk(gclk));
	jdff dff_B_timsz4Qi5_0(.din(w_dff_B_PJUHQmdO7_0),.dout(w_dff_B_timsz4Qi5_0),.clk(gclk));
	jdff dff_B_DHMhyWsv2_0(.din(w_dff_B_timsz4Qi5_0),.dout(w_dff_B_DHMhyWsv2_0),.clk(gclk));
	jdff dff_B_MWCuFCjn1_0(.din(w_dff_B_DHMhyWsv2_0),.dout(w_dff_B_MWCuFCjn1_0),.clk(gclk));
	jdff dff_B_hqSiKuxP5_0(.din(w_dff_B_MWCuFCjn1_0),.dout(w_dff_B_hqSiKuxP5_0),.clk(gclk));
	jdff dff_B_ASvLsKR52_0(.din(w_dff_B_hqSiKuxP5_0),.dout(w_dff_B_ASvLsKR52_0),.clk(gclk));
	jdff dff_B_4EYPuryV6_0(.din(w_dff_B_ASvLsKR52_0),.dout(w_dff_B_4EYPuryV6_0),.clk(gclk));
	jdff dff_B_bfXD3M9V8_0(.din(w_dff_B_4EYPuryV6_0),.dout(w_dff_B_bfXD3M9V8_0),.clk(gclk));
	jdff dff_B_E8z8KThg7_0(.din(w_dff_B_bfXD3M9V8_0),.dout(w_dff_B_E8z8KThg7_0),.clk(gclk));
	jdff dff_B_ARYa9xKC7_0(.din(w_dff_B_E8z8KThg7_0),.dout(w_dff_B_ARYa9xKC7_0),.clk(gclk));
	jdff dff_B_XnBYhEer7_0(.din(w_dff_B_ARYa9xKC7_0),.dout(w_dff_B_XnBYhEer7_0),.clk(gclk));
	jdff dff_B_39n8ryt86_0(.din(w_dff_B_XnBYhEer7_0),.dout(w_dff_B_39n8ryt86_0),.clk(gclk));
	jdff dff_B_mFbzyEFd7_0(.din(w_dff_B_39n8ryt86_0),.dout(w_dff_B_mFbzyEFd7_0),.clk(gclk));
	jdff dff_B_mPsRocZH1_0(.din(w_dff_B_mFbzyEFd7_0),.dout(w_dff_B_mPsRocZH1_0),.clk(gclk));
	jdff dff_B_H2ouOVSo6_0(.din(w_dff_B_mPsRocZH1_0),.dout(w_dff_B_H2ouOVSo6_0),.clk(gclk));
	jdff dff_B_zqeayftb6_0(.din(w_dff_B_H2ouOVSo6_0),.dout(w_dff_B_zqeayftb6_0),.clk(gclk));
	jdff dff_B_1OcOLfLf1_0(.din(w_dff_B_zqeayftb6_0),.dout(w_dff_B_1OcOLfLf1_0),.clk(gclk));
	jdff dff_B_hLBaU4Vj8_0(.din(w_dff_B_1OcOLfLf1_0),.dout(w_dff_B_hLBaU4Vj8_0),.clk(gclk));
	jdff dff_B_FSI0gpRE5_0(.din(w_dff_B_hLBaU4Vj8_0),.dout(w_dff_B_FSI0gpRE5_0),.clk(gclk));
	jdff dff_B_QyQe0UJL1_0(.din(w_dff_B_FSI0gpRE5_0),.dout(w_dff_B_QyQe0UJL1_0),.clk(gclk));
	jdff dff_B_GPWikoaz1_0(.din(w_dff_B_QyQe0UJL1_0),.dout(w_dff_B_GPWikoaz1_0),.clk(gclk));
	jdff dff_B_WA7ccQy34_0(.din(w_dff_B_GPWikoaz1_0),.dout(w_dff_B_WA7ccQy34_0),.clk(gclk));
	jdff dff_B_DiQtJIPr7_0(.din(w_dff_B_WA7ccQy34_0),.dout(w_dff_B_DiQtJIPr7_0),.clk(gclk));
	jdff dff_B_wYuGZ2Ig5_0(.din(w_dff_B_DiQtJIPr7_0),.dout(w_dff_B_wYuGZ2Ig5_0),.clk(gclk));
	jdff dff_B_LEg1aN8I1_0(.din(w_dff_B_wYuGZ2Ig5_0),.dout(w_dff_B_LEg1aN8I1_0),.clk(gclk));
	jdff dff_B_OkPLZWAi8_0(.din(w_dff_B_LEg1aN8I1_0),.dout(w_dff_B_OkPLZWAi8_0),.clk(gclk));
	jdff dff_B_DufBxwSX9_0(.din(w_dff_B_OkPLZWAi8_0),.dout(w_dff_B_DufBxwSX9_0),.clk(gclk));
	jdff dff_B_70nLApIG0_0(.din(w_dff_B_DufBxwSX9_0),.dout(w_dff_B_70nLApIG0_0),.clk(gclk));
	jdff dff_B_TX9Xt2la9_0(.din(w_dff_B_70nLApIG0_0),.dout(w_dff_B_TX9Xt2la9_0),.clk(gclk));
	jdff dff_B_GapYUI1h5_0(.din(w_dff_B_TX9Xt2la9_0),.dout(w_dff_B_GapYUI1h5_0),.clk(gclk));
	jdff dff_B_9svg7rmL1_0(.din(w_dff_B_GapYUI1h5_0),.dout(w_dff_B_9svg7rmL1_0),.clk(gclk));
	jdff dff_B_tWWdQgtJ4_0(.din(w_dff_B_9svg7rmL1_0),.dout(w_dff_B_tWWdQgtJ4_0),.clk(gclk));
	jdff dff_B_0CQMMybI4_0(.din(w_dff_B_tWWdQgtJ4_0),.dout(w_dff_B_0CQMMybI4_0),.clk(gclk));
	jdff dff_B_cYfT9H400_0(.din(w_dff_B_0CQMMybI4_0),.dout(w_dff_B_cYfT9H400_0),.clk(gclk));
	jdff dff_B_aqla3uee8_0(.din(w_dff_B_cYfT9H400_0),.dout(w_dff_B_aqla3uee8_0),.clk(gclk));
	jdff dff_B_Idkb6SYB6_0(.din(w_dff_B_aqla3uee8_0),.dout(w_dff_B_Idkb6SYB6_0),.clk(gclk));
	jdff dff_B_se6qxCOK7_0(.din(w_dff_B_Idkb6SYB6_0),.dout(w_dff_B_se6qxCOK7_0),.clk(gclk));
	jdff dff_B_a1OSw7zZ0_0(.din(w_dff_B_se6qxCOK7_0),.dout(w_dff_B_a1OSw7zZ0_0),.clk(gclk));
	jdff dff_B_O6ZXWT2t0_0(.din(w_dff_B_a1OSw7zZ0_0),.dout(w_dff_B_O6ZXWT2t0_0),.clk(gclk));
	jdff dff_B_4rJmYiWA4_0(.din(w_dff_B_O6ZXWT2t0_0),.dout(w_dff_B_4rJmYiWA4_0),.clk(gclk));
	jdff dff_B_JXHIGKBh9_0(.din(w_dff_B_4rJmYiWA4_0),.dout(w_dff_B_JXHIGKBh9_0),.clk(gclk));
	jdff dff_B_zTMJ1CSA8_0(.din(w_dff_B_JXHIGKBh9_0),.dout(w_dff_B_zTMJ1CSA8_0),.clk(gclk));
	jdff dff_B_r5wJPKfA1_0(.din(w_dff_B_zTMJ1CSA8_0),.dout(w_dff_B_r5wJPKfA1_0),.clk(gclk));
	jdff dff_B_T0elTxmH8_0(.din(w_dff_B_r5wJPKfA1_0),.dout(w_dff_B_T0elTxmH8_0),.clk(gclk));
	jdff dff_B_RHjZapdP3_0(.din(w_dff_B_T0elTxmH8_0),.dout(w_dff_B_RHjZapdP3_0),.clk(gclk));
	jdff dff_B_ziihU3C56_0(.din(w_dff_B_RHjZapdP3_0),.dout(w_dff_B_ziihU3C56_0),.clk(gclk));
	jdff dff_B_kb0qb4o00_0(.din(w_dff_B_ziihU3C56_0),.dout(w_dff_B_kb0qb4o00_0),.clk(gclk));
	jdff dff_B_oY8pBb783_0(.din(w_dff_B_kb0qb4o00_0),.dout(w_dff_B_oY8pBb783_0),.clk(gclk));
	jdff dff_B_z01nDMwv4_1(.din(n1116),.dout(w_dff_B_z01nDMwv4_1),.clk(gclk));
	jdff dff_B_6EtclvnV9_1(.din(w_dff_B_z01nDMwv4_1),.dout(w_dff_B_6EtclvnV9_1),.clk(gclk));
	jdff dff_B_ZBcu8scr0_1(.din(w_dff_B_6EtclvnV9_1),.dout(w_dff_B_ZBcu8scr0_1),.clk(gclk));
	jdff dff_B_LqkFspZw1_1(.din(w_dff_B_ZBcu8scr0_1),.dout(w_dff_B_LqkFspZw1_1),.clk(gclk));
	jdff dff_B_tXP1X49f7_1(.din(w_dff_B_LqkFspZw1_1),.dout(w_dff_B_tXP1X49f7_1),.clk(gclk));
	jdff dff_B_eCcyG9jT8_1(.din(w_dff_B_tXP1X49f7_1),.dout(w_dff_B_eCcyG9jT8_1),.clk(gclk));
	jdff dff_B_Uv9PxNtF9_1(.din(w_dff_B_eCcyG9jT8_1),.dout(w_dff_B_Uv9PxNtF9_1),.clk(gclk));
	jdff dff_B_HpBrX3Se1_1(.din(w_dff_B_Uv9PxNtF9_1),.dout(w_dff_B_HpBrX3Se1_1),.clk(gclk));
	jdff dff_B_MRgkquuw9_1(.din(w_dff_B_HpBrX3Se1_1),.dout(w_dff_B_MRgkquuw9_1),.clk(gclk));
	jdff dff_B_HOA0lw9V2_1(.din(w_dff_B_MRgkquuw9_1),.dout(w_dff_B_HOA0lw9V2_1),.clk(gclk));
	jdff dff_B_ONoDfZCu1_1(.din(w_dff_B_HOA0lw9V2_1),.dout(w_dff_B_ONoDfZCu1_1),.clk(gclk));
	jdff dff_B_MEYCNacy8_1(.din(w_dff_B_ONoDfZCu1_1),.dout(w_dff_B_MEYCNacy8_1),.clk(gclk));
	jdff dff_B_WPOUJTJr9_1(.din(w_dff_B_MEYCNacy8_1),.dout(w_dff_B_WPOUJTJr9_1),.clk(gclk));
	jdff dff_B_ppgNypcU2_1(.din(w_dff_B_WPOUJTJr9_1),.dout(w_dff_B_ppgNypcU2_1),.clk(gclk));
	jdff dff_B_AVKslCmw2_1(.din(w_dff_B_ppgNypcU2_1),.dout(w_dff_B_AVKslCmw2_1),.clk(gclk));
	jdff dff_B_TgzzxENF2_1(.din(w_dff_B_AVKslCmw2_1),.dout(w_dff_B_TgzzxENF2_1),.clk(gclk));
	jdff dff_B_3PUyYZIX2_1(.din(w_dff_B_TgzzxENF2_1),.dout(w_dff_B_3PUyYZIX2_1),.clk(gclk));
	jdff dff_B_DNpmCXYj4_1(.din(w_dff_B_3PUyYZIX2_1),.dout(w_dff_B_DNpmCXYj4_1),.clk(gclk));
	jdff dff_B_67KCkxOw9_1(.din(w_dff_B_DNpmCXYj4_1),.dout(w_dff_B_67KCkxOw9_1),.clk(gclk));
	jdff dff_B_CUHpFrCa8_1(.din(w_dff_B_67KCkxOw9_1),.dout(w_dff_B_CUHpFrCa8_1),.clk(gclk));
	jdff dff_B_zmYC0MD74_1(.din(w_dff_B_CUHpFrCa8_1),.dout(w_dff_B_zmYC0MD74_1),.clk(gclk));
	jdff dff_B_gmcrlBtl9_1(.din(w_dff_B_zmYC0MD74_1),.dout(w_dff_B_gmcrlBtl9_1),.clk(gclk));
	jdff dff_B_NesNbuze8_1(.din(w_dff_B_gmcrlBtl9_1),.dout(w_dff_B_NesNbuze8_1),.clk(gclk));
	jdff dff_B_cIPg8KD27_1(.din(w_dff_B_NesNbuze8_1),.dout(w_dff_B_cIPg8KD27_1),.clk(gclk));
	jdff dff_B_2JZ92O8j0_1(.din(w_dff_B_cIPg8KD27_1),.dout(w_dff_B_2JZ92O8j0_1),.clk(gclk));
	jdff dff_B_fVztKYZX7_1(.din(w_dff_B_2JZ92O8j0_1),.dout(w_dff_B_fVztKYZX7_1),.clk(gclk));
	jdff dff_B_IzdbYgxG7_1(.din(w_dff_B_fVztKYZX7_1),.dout(w_dff_B_IzdbYgxG7_1),.clk(gclk));
	jdff dff_B_1hjlMMYl6_1(.din(w_dff_B_IzdbYgxG7_1),.dout(w_dff_B_1hjlMMYl6_1),.clk(gclk));
	jdff dff_B_GLxaCAdr4_1(.din(w_dff_B_1hjlMMYl6_1),.dout(w_dff_B_GLxaCAdr4_1),.clk(gclk));
	jdff dff_B_MsmGbAwv0_1(.din(w_dff_B_GLxaCAdr4_1),.dout(w_dff_B_MsmGbAwv0_1),.clk(gclk));
	jdff dff_B_olb9qy8G0_1(.din(w_dff_B_MsmGbAwv0_1),.dout(w_dff_B_olb9qy8G0_1),.clk(gclk));
	jdff dff_B_sBQ2Plh99_1(.din(w_dff_B_olb9qy8G0_1),.dout(w_dff_B_sBQ2Plh99_1),.clk(gclk));
	jdff dff_B_sUg2zMX23_1(.din(w_dff_B_sBQ2Plh99_1),.dout(w_dff_B_sUg2zMX23_1),.clk(gclk));
	jdff dff_B_M4JPRDYr3_1(.din(w_dff_B_sUg2zMX23_1),.dout(w_dff_B_M4JPRDYr3_1),.clk(gclk));
	jdff dff_B_C4vEU0F57_1(.din(w_dff_B_M4JPRDYr3_1),.dout(w_dff_B_C4vEU0F57_1),.clk(gclk));
	jdff dff_B_pBcnD1kN2_1(.din(w_dff_B_C4vEU0F57_1),.dout(w_dff_B_pBcnD1kN2_1),.clk(gclk));
	jdff dff_B_YpoTIwnV5_1(.din(w_dff_B_pBcnD1kN2_1),.dout(w_dff_B_YpoTIwnV5_1),.clk(gclk));
	jdff dff_B_ecaywQ3W4_1(.din(w_dff_B_YpoTIwnV5_1),.dout(w_dff_B_ecaywQ3W4_1),.clk(gclk));
	jdff dff_B_SNpKsaVS6_1(.din(w_dff_B_ecaywQ3W4_1),.dout(w_dff_B_SNpKsaVS6_1),.clk(gclk));
	jdff dff_B_xDU3utD33_1(.din(w_dff_B_SNpKsaVS6_1),.dout(w_dff_B_xDU3utD33_1),.clk(gclk));
	jdff dff_B_IOoVO09q8_1(.din(w_dff_B_xDU3utD33_1),.dout(w_dff_B_IOoVO09q8_1),.clk(gclk));
	jdff dff_B_r7OxnRq26_1(.din(w_dff_B_IOoVO09q8_1),.dout(w_dff_B_r7OxnRq26_1),.clk(gclk));
	jdff dff_B_ncp8gaxD0_1(.din(w_dff_B_r7OxnRq26_1),.dout(w_dff_B_ncp8gaxD0_1),.clk(gclk));
	jdff dff_B_5AKjTN8n2_1(.din(w_dff_B_ncp8gaxD0_1),.dout(w_dff_B_5AKjTN8n2_1),.clk(gclk));
	jdff dff_B_KUJBXrMG0_1(.din(w_dff_B_5AKjTN8n2_1),.dout(w_dff_B_KUJBXrMG0_1),.clk(gclk));
	jdff dff_B_YREIpQpD8_1(.din(w_dff_B_KUJBXrMG0_1),.dout(w_dff_B_YREIpQpD8_1),.clk(gclk));
	jdff dff_B_t3AX2Ue72_1(.din(w_dff_B_YREIpQpD8_1),.dout(w_dff_B_t3AX2Ue72_1),.clk(gclk));
	jdff dff_B_la8TEb3D4_1(.din(w_dff_B_t3AX2Ue72_1),.dout(w_dff_B_la8TEb3D4_1),.clk(gclk));
	jdff dff_B_xjVI8tzM6_1(.din(w_dff_B_la8TEb3D4_1),.dout(w_dff_B_xjVI8tzM6_1),.clk(gclk));
	jdff dff_B_kkNod70o8_1(.din(w_dff_B_xjVI8tzM6_1),.dout(w_dff_B_kkNod70o8_1),.clk(gclk));
	jdff dff_B_bmzszsJ56_1(.din(w_dff_B_kkNod70o8_1),.dout(w_dff_B_bmzszsJ56_1),.clk(gclk));
	jdff dff_B_o6lofO308_1(.din(w_dff_B_bmzszsJ56_1),.dout(w_dff_B_o6lofO308_1),.clk(gclk));
	jdff dff_B_kYVXWfTh4_1(.din(w_dff_B_o6lofO308_1),.dout(w_dff_B_kYVXWfTh4_1),.clk(gclk));
	jdff dff_B_vLlqJdbV1_1(.din(w_dff_B_kYVXWfTh4_1),.dout(w_dff_B_vLlqJdbV1_1),.clk(gclk));
	jdff dff_B_K7P2meAE5_1(.din(w_dff_B_vLlqJdbV1_1),.dout(w_dff_B_K7P2meAE5_1),.clk(gclk));
	jdff dff_B_XAzC2BvG2_1(.din(w_dff_B_K7P2meAE5_1),.dout(w_dff_B_XAzC2BvG2_1),.clk(gclk));
	jdff dff_B_ip7Lp4sn8_1(.din(w_dff_B_XAzC2BvG2_1),.dout(w_dff_B_ip7Lp4sn8_1),.clk(gclk));
	jdff dff_B_0OQMVJdH3_1(.din(w_dff_B_ip7Lp4sn8_1),.dout(w_dff_B_0OQMVJdH3_1),.clk(gclk));
	jdff dff_B_anGpywdC9_1(.din(w_dff_B_0OQMVJdH3_1),.dout(w_dff_B_anGpywdC9_1),.clk(gclk));
	jdff dff_B_6oxiMOGB8_1(.din(w_dff_B_anGpywdC9_1),.dout(w_dff_B_6oxiMOGB8_1),.clk(gclk));
	jdff dff_B_NGvF5hsp6_1(.din(w_dff_B_6oxiMOGB8_1),.dout(w_dff_B_NGvF5hsp6_1),.clk(gclk));
	jdff dff_B_DHufxwt50_1(.din(w_dff_B_NGvF5hsp6_1),.dout(w_dff_B_DHufxwt50_1),.clk(gclk));
	jdff dff_B_rotnroWx9_1(.din(w_dff_B_DHufxwt50_1),.dout(w_dff_B_rotnroWx9_1),.clk(gclk));
	jdff dff_B_6vbS29bj1_1(.din(w_dff_B_rotnroWx9_1),.dout(w_dff_B_6vbS29bj1_1),.clk(gclk));
	jdff dff_B_Jw6tLjP76_1(.din(w_dff_B_6vbS29bj1_1),.dout(w_dff_B_Jw6tLjP76_1),.clk(gclk));
	jdff dff_B_oZMBEcqh6_1(.din(w_dff_B_Jw6tLjP76_1),.dout(w_dff_B_oZMBEcqh6_1),.clk(gclk));
	jdff dff_B_jTWHkSJH5_1(.din(w_dff_B_oZMBEcqh6_1),.dout(w_dff_B_jTWHkSJH5_1),.clk(gclk));
	jdff dff_B_6FxYUHsi9_1(.din(w_dff_B_jTWHkSJH5_1),.dout(w_dff_B_6FxYUHsi9_1),.clk(gclk));
	jdff dff_B_IlitXWrR5_1(.din(w_dff_B_6FxYUHsi9_1),.dout(w_dff_B_IlitXWrR5_1),.clk(gclk));
	jdff dff_B_CKCoXO692_1(.din(w_dff_B_IlitXWrR5_1),.dout(w_dff_B_CKCoXO692_1),.clk(gclk));
	jdff dff_B_SNgoNgaX4_1(.din(w_dff_B_CKCoXO692_1),.dout(w_dff_B_SNgoNgaX4_1),.clk(gclk));
	jdff dff_B_eriyZy030_1(.din(w_dff_B_SNgoNgaX4_1),.dout(w_dff_B_eriyZy030_1),.clk(gclk));
	jdff dff_B_wNtVVCzX3_1(.din(w_dff_B_eriyZy030_1),.dout(w_dff_B_wNtVVCzX3_1),.clk(gclk));
	jdff dff_B_KVFVZLHq7_1(.din(w_dff_B_wNtVVCzX3_1),.dout(w_dff_B_KVFVZLHq7_1),.clk(gclk));
	jdff dff_B_8KVgezxO5_1(.din(w_dff_B_KVFVZLHq7_1),.dout(w_dff_B_8KVgezxO5_1),.clk(gclk));
	jdff dff_B_gFiwlnzb6_1(.din(w_dff_B_8KVgezxO5_1),.dout(w_dff_B_gFiwlnzb6_1),.clk(gclk));
	jdff dff_B_sNmxpQxx6_1(.din(w_dff_B_gFiwlnzb6_1),.dout(w_dff_B_sNmxpQxx6_1),.clk(gclk));
	jdff dff_B_924ILho16_1(.din(w_dff_B_sNmxpQxx6_1),.dout(w_dff_B_924ILho16_1),.clk(gclk));
	jdff dff_B_9LdlSj4V6_1(.din(w_dff_B_924ILho16_1),.dout(w_dff_B_9LdlSj4V6_1),.clk(gclk));
	jdff dff_B_DFKto3wA5_1(.din(w_dff_B_9LdlSj4V6_1),.dout(w_dff_B_DFKto3wA5_1),.clk(gclk));
	jdff dff_B_UWXbKLbW8_1(.din(w_dff_B_DFKto3wA5_1),.dout(w_dff_B_UWXbKLbW8_1),.clk(gclk));
	jdff dff_B_trU4JIUl8_1(.din(w_dff_B_UWXbKLbW8_1),.dout(w_dff_B_trU4JIUl8_1),.clk(gclk));
	jdff dff_B_Knj0R4De6_1(.din(w_dff_B_trU4JIUl8_1),.dout(w_dff_B_Knj0R4De6_1),.clk(gclk));
	jdff dff_B_yNA9Lu6y2_1(.din(w_dff_B_Knj0R4De6_1),.dout(w_dff_B_yNA9Lu6y2_1),.clk(gclk));
	jdff dff_B_4lLcYCez9_1(.din(w_dff_B_yNA9Lu6y2_1),.dout(w_dff_B_4lLcYCez9_1),.clk(gclk));
	jdff dff_B_HuepJOaS9_1(.din(w_dff_B_4lLcYCez9_1),.dout(w_dff_B_HuepJOaS9_1),.clk(gclk));
	jdff dff_B_2BHqe7X89_1(.din(w_dff_B_HuepJOaS9_1),.dout(w_dff_B_2BHqe7X89_1),.clk(gclk));
	jdff dff_B_itN1NFKy7_1(.din(w_dff_B_2BHqe7X89_1),.dout(w_dff_B_itN1NFKy7_1),.clk(gclk));
	jdff dff_B_oSek1iaI0_1(.din(w_dff_B_itN1NFKy7_1),.dout(w_dff_B_oSek1iaI0_1),.clk(gclk));
	jdff dff_B_YMziUT3Y2_1(.din(w_dff_B_oSek1iaI0_1),.dout(w_dff_B_YMziUT3Y2_1),.clk(gclk));
	jdff dff_B_3rqvSSHv2_1(.din(w_dff_B_YMziUT3Y2_1),.dout(w_dff_B_3rqvSSHv2_1),.clk(gclk));
	jdff dff_B_ttCYVUMl4_1(.din(w_dff_B_3rqvSSHv2_1),.dout(w_dff_B_ttCYVUMl4_1),.clk(gclk));
	jdff dff_B_HD3rvZxt5_1(.din(w_dff_B_ttCYVUMl4_1),.dout(w_dff_B_HD3rvZxt5_1),.clk(gclk));
	jdff dff_B_zmpdtUQ97_1(.din(w_dff_B_HD3rvZxt5_1),.dout(w_dff_B_zmpdtUQ97_1),.clk(gclk));
	jdff dff_B_rManAGOy5_1(.din(w_dff_B_zmpdtUQ97_1),.dout(w_dff_B_rManAGOy5_1),.clk(gclk));
	jdff dff_B_UEUloay98_1(.din(w_dff_B_rManAGOy5_1),.dout(w_dff_B_UEUloay98_1),.clk(gclk));
	jdff dff_B_SpQZ42fl5_1(.din(w_dff_B_UEUloay98_1),.dout(w_dff_B_SpQZ42fl5_1),.clk(gclk));
	jdff dff_B_SeLCNm5T1_1(.din(w_dff_B_SpQZ42fl5_1),.dout(w_dff_B_SeLCNm5T1_1),.clk(gclk));
	jdff dff_B_jMmJiZJx6_1(.din(w_dff_B_SeLCNm5T1_1),.dout(w_dff_B_jMmJiZJx6_1),.clk(gclk));
	jdff dff_B_bNTJcCDt2_1(.din(w_dff_B_jMmJiZJx6_1),.dout(w_dff_B_bNTJcCDt2_1),.clk(gclk));
	jdff dff_B_6BHKAgrd5_1(.din(w_dff_B_bNTJcCDt2_1),.dout(w_dff_B_6BHKAgrd5_1),.clk(gclk));
	jdff dff_B_jxo5zOz77_1(.din(w_dff_B_6BHKAgrd5_1),.dout(w_dff_B_jxo5zOz77_1),.clk(gclk));
	jdff dff_B_lbhvHxMg9_1(.din(w_dff_B_jxo5zOz77_1),.dout(w_dff_B_lbhvHxMg9_1),.clk(gclk));
	jdff dff_B_xqOVZdHf7_1(.din(w_dff_B_lbhvHxMg9_1),.dout(w_dff_B_xqOVZdHf7_1),.clk(gclk));
	jdff dff_B_Jgzy3lKO9_1(.din(w_dff_B_xqOVZdHf7_1),.dout(w_dff_B_Jgzy3lKO9_1),.clk(gclk));
	jdff dff_B_AJU9a7Vx9_1(.din(w_dff_B_Jgzy3lKO9_1),.dout(w_dff_B_AJU9a7Vx9_1),.clk(gclk));
	jdff dff_B_gS8sz9dN8_1(.din(w_dff_B_AJU9a7Vx9_1),.dout(w_dff_B_gS8sz9dN8_1),.clk(gclk));
	jdff dff_B_uyZpVk0P3_1(.din(w_dff_B_gS8sz9dN8_1),.dout(w_dff_B_uyZpVk0P3_1),.clk(gclk));
	jdff dff_B_xGhH23sQ3_1(.din(w_dff_B_uyZpVk0P3_1),.dout(w_dff_B_xGhH23sQ3_1),.clk(gclk));
	jdff dff_B_nUbtSo662_1(.din(w_dff_B_xGhH23sQ3_1),.dout(w_dff_B_nUbtSo662_1),.clk(gclk));
	jdff dff_B_lx2Ms7HH6_1(.din(w_dff_B_nUbtSo662_1),.dout(w_dff_B_lx2Ms7HH6_1),.clk(gclk));
	jdff dff_B_aTskClIk1_1(.din(w_dff_B_lx2Ms7HH6_1),.dout(w_dff_B_aTskClIk1_1),.clk(gclk));
	jdff dff_B_q4H6WhDe7_1(.din(w_dff_B_aTskClIk1_1),.dout(w_dff_B_q4H6WhDe7_1),.clk(gclk));
	jdff dff_B_ac2BNYvd5_1(.din(w_dff_B_q4H6WhDe7_1),.dout(w_dff_B_ac2BNYvd5_1),.clk(gclk));
	jdff dff_B_P3pcQVXZ3_1(.din(w_dff_B_ac2BNYvd5_1),.dout(w_dff_B_P3pcQVXZ3_1),.clk(gclk));
	jdff dff_B_qTfinytC8_1(.din(w_dff_B_P3pcQVXZ3_1),.dout(w_dff_B_qTfinytC8_1),.clk(gclk));
	jdff dff_B_T4KtDsWT1_1(.din(w_dff_B_qTfinytC8_1),.dout(w_dff_B_T4KtDsWT1_1),.clk(gclk));
	jdff dff_B_Jt2yUwxU0_1(.din(w_dff_B_T4KtDsWT1_1),.dout(w_dff_B_Jt2yUwxU0_1),.clk(gclk));
	jdff dff_B_72b234om0_1(.din(w_dff_B_Jt2yUwxU0_1),.dout(w_dff_B_72b234om0_1),.clk(gclk));
	jdff dff_B_uyXBKvGh3_1(.din(w_dff_B_72b234om0_1),.dout(w_dff_B_uyXBKvGh3_1),.clk(gclk));
	jdff dff_B_QDVmiuHX6_1(.din(w_dff_B_uyXBKvGh3_1),.dout(w_dff_B_QDVmiuHX6_1),.clk(gclk));
	jdff dff_B_Dkr9JPcC7_1(.din(w_dff_B_QDVmiuHX6_1),.dout(w_dff_B_Dkr9JPcC7_1),.clk(gclk));
	jdff dff_B_2QfVLIYH5_0(.din(n1117),.dout(w_dff_B_2QfVLIYH5_0),.clk(gclk));
	jdff dff_B_Wes1Bi1r1_0(.din(w_dff_B_2QfVLIYH5_0),.dout(w_dff_B_Wes1Bi1r1_0),.clk(gclk));
	jdff dff_B_UIsyTEMs9_0(.din(w_dff_B_Wes1Bi1r1_0),.dout(w_dff_B_UIsyTEMs9_0),.clk(gclk));
	jdff dff_B_4BfkN1Pp6_0(.din(w_dff_B_UIsyTEMs9_0),.dout(w_dff_B_4BfkN1Pp6_0),.clk(gclk));
	jdff dff_B_BrBkJX9S6_0(.din(w_dff_B_4BfkN1Pp6_0),.dout(w_dff_B_BrBkJX9S6_0),.clk(gclk));
	jdff dff_B_XQSODnrH6_0(.din(w_dff_B_BrBkJX9S6_0),.dout(w_dff_B_XQSODnrH6_0),.clk(gclk));
	jdff dff_B_95JaTi651_0(.din(w_dff_B_XQSODnrH6_0),.dout(w_dff_B_95JaTi651_0),.clk(gclk));
	jdff dff_B_0hjvQMEF6_0(.din(w_dff_B_95JaTi651_0),.dout(w_dff_B_0hjvQMEF6_0),.clk(gclk));
	jdff dff_B_LI958ltJ2_0(.din(w_dff_B_0hjvQMEF6_0),.dout(w_dff_B_LI958ltJ2_0),.clk(gclk));
	jdff dff_B_2Gtl6xCK7_0(.din(w_dff_B_LI958ltJ2_0),.dout(w_dff_B_2Gtl6xCK7_0),.clk(gclk));
	jdff dff_B_In46HT6Z1_0(.din(w_dff_B_2Gtl6xCK7_0),.dout(w_dff_B_In46HT6Z1_0),.clk(gclk));
	jdff dff_B_rxc7WBZp7_0(.din(w_dff_B_In46HT6Z1_0),.dout(w_dff_B_rxc7WBZp7_0),.clk(gclk));
	jdff dff_B_5QllazsF0_0(.din(w_dff_B_rxc7WBZp7_0),.dout(w_dff_B_5QllazsF0_0),.clk(gclk));
	jdff dff_B_pd7me7DP9_0(.din(w_dff_B_5QllazsF0_0),.dout(w_dff_B_pd7me7DP9_0),.clk(gclk));
	jdff dff_B_Ng3dVv7L3_0(.din(w_dff_B_pd7me7DP9_0),.dout(w_dff_B_Ng3dVv7L3_0),.clk(gclk));
	jdff dff_B_paORnNy44_0(.din(w_dff_B_Ng3dVv7L3_0),.dout(w_dff_B_paORnNy44_0),.clk(gclk));
	jdff dff_B_tYW6IXLz0_0(.din(w_dff_B_paORnNy44_0),.dout(w_dff_B_tYW6IXLz0_0),.clk(gclk));
	jdff dff_B_PNkgAw1z0_0(.din(w_dff_B_tYW6IXLz0_0),.dout(w_dff_B_PNkgAw1z0_0),.clk(gclk));
	jdff dff_B_jFxQUTmn4_0(.din(w_dff_B_PNkgAw1z0_0),.dout(w_dff_B_jFxQUTmn4_0),.clk(gclk));
	jdff dff_B_KOUcbzYt3_0(.din(w_dff_B_jFxQUTmn4_0),.dout(w_dff_B_KOUcbzYt3_0),.clk(gclk));
	jdff dff_B_c4kYWWfy1_0(.din(w_dff_B_KOUcbzYt3_0),.dout(w_dff_B_c4kYWWfy1_0),.clk(gclk));
	jdff dff_B_E8XILlGk4_0(.din(w_dff_B_c4kYWWfy1_0),.dout(w_dff_B_E8XILlGk4_0),.clk(gclk));
	jdff dff_B_uirCvuzF7_0(.din(w_dff_B_E8XILlGk4_0),.dout(w_dff_B_uirCvuzF7_0),.clk(gclk));
	jdff dff_B_qr4s4FB56_0(.din(w_dff_B_uirCvuzF7_0),.dout(w_dff_B_qr4s4FB56_0),.clk(gclk));
	jdff dff_B_X7dPO1SY9_0(.din(w_dff_B_qr4s4FB56_0),.dout(w_dff_B_X7dPO1SY9_0),.clk(gclk));
	jdff dff_B_bLwAzQAS1_0(.din(w_dff_B_X7dPO1SY9_0),.dout(w_dff_B_bLwAzQAS1_0),.clk(gclk));
	jdff dff_B_NQR8LqCj4_0(.din(w_dff_B_bLwAzQAS1_0),.dout(w_dff_B_NQR8LqCj4_0),.clk(gclk));
	jdff dff_B_gx2VO75d9_0(.din(w_dff_B_NQR8LqCj4_0),.dout(w_dff_B_gx2VO75d9_0),.clk(gclk));
	jdff dff_B_e80M7d9g1_0(.din(w_dff_B_gx2VO75d9_0),.dout(w_dff_B_e80M7d9g1_0),.clk(gclk));
	jdff dff_B_0dzIYKbP7_0(.din(w_dff_B_e80M7d9g1_0),.dout(w_dff_B_0dzIYKbP7_0),.clk(gclk));
	jdff dff_B_kY197Etg9_0(.din(w_dff_B_0dzIYKbP7_0),.dout(w_dff_B_kY197Etg9_0),.clk(gclk));
	jdff dff_B_i7ozsX6s0_0(.din(w_dff_B_kY197Etg9_0),.dout(w_dff_B_i7ozsX6s0_0),.clk(gclk));
	jdff dff_B_9KdxYw2t2_0(.din(w_dff_B_i7ozsX6s0_0),.dout(w_dff_B_9KdxYw2t2_0),.clk(gclk));
	jdff dff_B_xoD3q1Lo0_0(.din(w_dff_B_9KdxYw2t2_0),.dout(w_dff_B_xoD3q1Lo0_0),.clk(gclk));
	jdff dff_B_h0i9s6pm8_0(.din(w_dff_B_xoD3q1Lo0_0),.dout(w_dff_B_h0i9s6pm8_0),.clk(gclk));
	jdff dff_B_gyFCuJcJ4_0(.din(w_dff_B_h0i9s6pm8_0),.dout(w_dff_B_gyFCuJcJ4_0),.clk(gclk));
	jdff dff_B_dZZslLEA1_0(.din(w_dff_B_gyFCuJcJ4_0),.dout(w_dff_B_dZZslLEA1_0),.clk(gclk));
	jdff dff_B_zcoK2CbP8_0(.din(w_dff_B_dZZslLEA1_0),.dout(w_dff_B_zcoK2CbP8_0),.clk(gclk));
	jdff dff_B_LtYDAigb7_0(.din(w_dff_B_zcoK2CbP8_0),.dout(w_dff_B_LtYDAigb7_0),.clk(gclk));
	jdff dff_B_xC8rs0ZH0_0(.din(w_dff_B_LtYDAigb7_0),.dout(w_dff_B_xC8rs0ZH0_0),.clk(gclk));
	jdff dff_B_97RnY4z27_0(.din(w_dff_B_xC8rs0ZH0_0),.dout(w_dff_B_97RnY4z27_0),.clk(gclk));
	jdff dff_B_wwrpkPNY5_0(.din(w_dff_B_97RnY4z27_0),.dout(w_dff_B_wwrpkPNY5_0),.clk(gclk));
	jdff dff_B_KPx9lQ8r3_0(.din(w_dff_B_wwrpkPNY5_0),.dout(w_dff_B_KPx9lQ8r3_0),.clk(gclk));
	jdff dff_B_qHUuajeQ1_0(.din(w_dff_B_KPx9lQ8r3_0),.dout(w_dff_B_qHUuajeQ1_0),.clk(gclk));
	jdff dff_B_Pm4eCqHe4_0(.din(w_dff_B_qHUuajeQ1_0),.dout(w_dff_B_Pm4eCqHe4_0),.clk(gclk));
	jdff dff_B_wI1OGoCG9_0(.din(w_dff_B_Pm4eCqHe4_0),.dout(w_dff_B_wI1OGoCG9_0),.clk(gclk));
	jdff dff_B_3RujAxvW8_0(.din(w_dff_B_wI1OGoCG9_0),.dout(w_dff_B_3RujAxvW8_0),.clk(gclk));
	jdff dff_B_Uoqk2gai7_0(.din(w_dff_B_3RujAxvW8_0),.dout(w_dff_B_Uoqk2gai7_0),.clk(gclk));
	jdff dff_B_lQMt7VwU9_0(.din(w_dff_B_Uoqk2gai7_0),.dout(w_dff_B_lQMt7VwU9_0),.clk(gclk));
	jdff dff_B_DlHCO0Au0_0(.din(w_dff_B_lQMt7VwU9_0),.dout(w_dff_B_DlHCO0Au0_0),.clk(gclk));
	jdff dff_B_qOQepiXU5_0(.din(w_dff_B_DlHCO0Au0_0),.dout(w_dff_B_qOQepiXU5_0),.clk(gclk));
	jdff dff_B_MKtVx2j64_0(.din(w_dff_B_qOQepiXU5_0),.dout(w_dff_B_MKtVx2j64_0),.clk(gclk));
	jdff dff_B_1HUQQNxE1_0(.din(w_dff_B_MKtVx2j64_0),.dout(w_dff_B_1HUQQNxE1_0),.clk(gclk));
	jdff dff_B_9n9MJrX61_0(.din(w_dff_B_1HUQQNxE1_0),.dout(w_dff_B_9n9MJrX61_0),.clk(gclk));
	jdff dff_B_HoqXpdaz5_0(.din(w_dff_B_9n9MJrX61_0),.dout(w_dff_B_HoqXpdaz5_0),.clk(gclk));
	jdff dff_B_t6nFwwmc3_0(.din(w_dff_B_HoqXpdaz5_0),.dout(w_dff_B_t6nFwwmc3_0),.clk(gclk));
	jdff dff_B_nKknmpYo9_0(.din(w_dff_B_t6nFwwmc3_0),.dout(w_dff_B_nKknmpYo9_0),.clk(gclk));
	jdff dff_B_rKedzUXh7_0(.din(w_dff_B_nKknmpYo9_0),.dout(w_dff_B_rKedzUXh7_0),.clk(gclk));
	jdff dff_B_V7vZN6FK0_0(.din(w_dff_B_rKedzUXh7_0),.dout(w_dff_B_V7vZN6FK0_0),.clk(gclk));
	jdff dff_B_lQpIsANE1_0(.din(w_dff_B_V7vZN6FK0_0),.dout(w_dff_B_lQpIsANE1_0),.clk(gclk));
	jdff dff_B_7aoBpfmz5_0(.din(w_dff_B_lQpIsANE1_0),.dout(w_dff_B_7aoBpfmz5_0),.clk(gclk));
	jdff dff_B_g49WO7MT8_0(.din(w_dff_B_7aoBpfmz5_0),.dout(w_dff_B_g49WO7MT8_0),.clk(gclk));
	jdff dff_B_MMDdDQD77_0(.din(w_dff_B_g49WO7MT8_0),.dout(w_dff_B_MMDdDQD77_0),.clk(gclk));
	jdff dff_B_nmYTSN6j2_0(.din(w_dff_B_MMDdDQD77_0),.dout(w_dff_B_nmYTSN6j2_0),.clk(gclk));
	jdff dff_B_d8TqjGOz3_0(.din(w_dff_B_nmYTSN6j2_0),.dout(w_dff_B_d8TqjGOz3_0),.clk(gclk));
	jdff dff_B_IcaMaKP03_0(.din(w_dff_B_d8TqjGOz3_0),.dout(w_dff_B_IcaMaKP03_0),.clk(gclk));
	jdff dff_B_yGQm8Yee8_0(.din(w_dff_B_IcaMaKP03_0),.dout(w_dff_B_yGQm8Yee8_0),.clk(gclk));
	jdff dff_B_QtqRXhAW0_0(.din(w_dff_B_yGQm8Yee8_0),.dout(w_dff_B_QtqRXhAW0_0),.clk(gclk));
	jdff dff_B_QeyUCVkz9_0(.din(w_dff_B_QtqRXhAW0_0),.dout(w_dff_B_QeyUCVkz9_0),.clk(gclk));
	jdff dff_B_ZqSRhkFK7_0(.din(w_dff_B_QeyUCVkz9_0),.dout(w_dff_B_ZqSRhkFK7_0),.clk(gclk));
	jdff dff_B_luahPtJk9_0(.din(w_dff_B_ZqSRhkFK7_0),.dout(w_dff_B_luahPtJk9_0),.clk(gclk));
	jdff dff_B_onDud58R2_0(.din(w_dff_B_luahPtJk9_0),.dout(w_dff_B_onDud58R2_0),.clk(gclk));
	jdff dff_B_MLyS5MlY8_0(.din(w_dff_B_onDud58R2_0),.dout(w_dff_B_MLyS5MlY8_0),.clk(gclk));
	jdff dff_B_BhJ4dnG18_0(.din(w_dff_B_MLyS5MlY8_0),.dout(w_dff_B_BhJ4dnG18_0),.clk(gclk));
	jdff dff_B_ldVdQmma7_0(.din(w_dff_B_BhJ4dnG18_0),.dout(w_dff_B_ldVdQmma7_0),.clk(gclk));
	jdff dff_B_1aJlZVpr2_0(.din(w_dff_B_ldVdQmma7_0),.dout(w_dff_B_1aJlZVpr2_0),.clk(gclk));
	jdff dff_B_upfcGmyu1_0(.din(w_dff_B_1aJlZVpr2_0),.dout(w_dff_B_upfcGmyu1_0),.clk(gclk));
	jdff dff_B_xV9BH7HW1_0(.din(w_dff_B_upfcGmyu1_0),.dout(w_dff_B_xV9BH7HW1_0),.clk(gclk));
	jdff dff_B_kVcx0yfU9_0(.din(w_dff_B_xV9BH7HW1_0),.dout(w_dff_B_kVcx0yfU9_0),.clk(gclk));
	jdff dff_B_T9G1J35g1_0(.din(w_dff_B_kVcx0yfU9_0),.dout(w_dff_B_T9G1J35g1_0),.clk(gclk));
	jdff dff_B_EybFPoWC5_0(.din(w_dff_B_T9G1J35g1_0),.dout(w_dff_B_EybFPoWC5_0),.clk(gclk));
	jdff dff_B_1xv37al60_0(.din(w_dff_B_EybFPoWC5_0),.dout(w_dff_B_1xv37al60_0),.clk(gclk));
	jdff dff_B_YOXAaZZZ7_0(.din(w_dff_B_1xv37al60_0),.dout(w_dff_B_YOXAaZZZ7_0),.clk(gclk));
	jdff dff_B_Mg0wGt1V0_0(.din(w_dff_B_YOXAaZZZ7_0),.dout(w_dff_B_Mg0wGt1V0_0),.clk(gclk));
	jdff dff_B_POLVBjgc3_0(.din(w_dff_B_Mg0wGt1V0_0),.dout(w_dff_B_POLVBjgc3_0),.clk(gclk));
	jdff dff_B_ZQprZfvQ5_0(.din(w_dff_B_POLVBjgc3_0),.dout(w_dff_B_ZQprZfvQ5_0),.clk(gclk));
	jdff dff_B_DqUs78GW9_0(.din(w_dff_B_ZQprZfvQ5_0),.dout(w_dff_B_DqUs78GW9_0),.clk(gclk));
	jdff dff_B_BszbWXgZ0_0(.din(w_dff_B_DqUs78GW9_0),.dout(w_dff_B_BszbWXgZ0_0),.clk(gclk));
	jdff dff_B_1umRlSl88_0(.din(w_dff_B_BszbWXgZ0_0),.dout(w_dff_B_1umRlSl88_0),.clk(gclk));
	jdff dff_B_rm6x90Wr2_0(.din(w_dff_B_1umRlSl88_0),.dout(w_dff_B_rm6x90Wr2_0),.clk(gclk));
	jdff dff_B_FeSijBGi5_0(.din(w_dff_B_rm6x90Wr2_0),.dout(w_dff_B_FeSijBGi5_0),.clk(gclk));
	jdff dff_B_9B6tyNHQ4_0(.din(w_dff_B_FeSijBGi5_0),.dout(w_dff_B_9B6tyNHQ4_0),.clk(gclk));
	jdff dff_B_HpvtjtJC5_0(.din(w_dff_B_9B6tyNHQ4_0),.dout(w_dff_B_HpvtjtJC5_0),.clk(gclk));
	jdff dff_B_uIwZqBG17_0(.din(w_dff_B_HpvtjtJC5_0),.dout(w_dff_B_uIwZqBG17_0),.clk(gclk));
	jdff dff_B_QpDocHiI5_0(.din(w_dff_B_uIwZqBG17_0),.dout(w_dff_B_QpDocHiI5_0),.clk(gclk));
	jdff dff_B_9Wsz7g1n1_0(.din(w_dff_B_QpDocHiI5_0),.dout(w_dff_B_9Wsz7g1n1_0),.clk(gclk));
	jdff dff_B_QWohCsaE2_0(.din(w_dff_B_9Wsz7g1n1_0),.dout(w_dff_B_QWohCsaE2_0),.clk(gclk));
	jdff dff_B_DxydY4YS6_0(.din(w_dff_B_QWohCsaE2_0),.dout(w_dff_B_DxydY4YS6_0),.clk(gclk));
	jdff dff_B_HSoN7PQp5_0(.din(w_dff_B_DxydY4YS6_0),.dout(w_dff_B_HSoN7PQp5_0),.clk(gclk));
	jdff dff_B_d291vfqe6_0(.din(w_dff_B_HSoN7PQp5_0),.dout(w_dff_B_d291vfqe6_0),.clk(gclk));
	jdff dff_B_jGs1Z1vX5_0(.din(w_dff_B_d291vfqe6_0),.dout(w_dff_B_jGs1Z1vX5_0),.clk(gclk));
	jdff dff_B_MK4eVmub9_0(.din(w_dff_B_jGs1Z1vX5_0),.dout(w_dff_B_MK4eVmub9_0),.clk(gclk));
	jdff dff_B_TfcBQnjB7_0(.din(w_dff_B_MK4eVmub9_0),.dout(w_dff_B_TfcBQnjB7_0),.clk(gclk));
	jdff dff_B_gjEZsume5_0(.din(w_dff_B_TfcBQnjB7_0),.dout(w_dff_B_gjEZsume5_0),.clk(gclk));
	jdff dff_B_aGv1906U0_0(.din(w_dff_B_gjEZsume5_0),.dout(w_dff_B_aGv1906U0_0),.clk(gclk));
	jdff dff_B_JIAURANF6_0(.din(w_dff_B_aGv1906U0_0),.dout(w_dff_B_JIAURANF6_0),.clk(gclk));
	jdff dff_B_0v4CG99s9_0(.din(w_dff_B_JIAURANF6_0),.dout(w_dff_B_0v4CG99s9_0),.clk(gclk));
	jdff dff_B_zhjxi2Ld9_0(.din(w_dff_B_0v4CG99s9_0),.dout(w_dff_B_zhjxi2Ld9_0),.clk(gclk));
	jdff dff_B_RArV20Il7_0(.din(w_dff_B_zhjxi2Ld9_0),.dout(w_dff_B_RArV20Il7_0),.clk(gclk));
	jdff dff_B_kHjcuUnU5_0(.din(w_dff_B_RArV20Il7_0),.dout(w_dff_B_kHjcuUnU5_0),.clk(gclk));
	jdff dff_B_tR6hnRcF9_0(.din(w_dff_B_kHjcuUnU5_0),.dout(w_dff_B_tR6hnRcF9_0),.clk(gclk));
	jdff dff_B_X4yn2Anp8_0(.din(w_dff_B_tR6hnRcF9_0),.dout(w_dff_B_X4yn2Anp8_0),.clk(gclk));
	jdff dff_B_wtkyyWPf7_0(.din(w_dff_B_X4yn2Anp8_0),.dout(w_dff_B_wtkyyWPf7_0),.clk(gclk));
	jdff dff_B_Sl9F6Et71_0(.din(w_dff_B_wtkyyWPf7_0),.dout(w_dff_B_Sl9F6Et71_0),.clk(gclk));
	jdff dff_B_jTE3N4Z76_0(.din(w_dff_B_Sl9F6Et71_0),.dout(w_dff_B_jTE3N4Z76_0),.clk(gclk));
	jdff dff_B_4rxem5xX4_0(.din(w_dff_B_jTE3N4Z76_0),.dout(w_dff_B_4rxem5xX4_0),.clk(gclk));
	jdff dff_B_sqISUf5R2_0(.din(w_dff_B_4rxem5xX4_0),.dout(w_dff_B_sqISUf5R2_0),.clk(gclk));
	jdff dff_B_aHDWCnpi6_0(.din(w_dff_B_sqISUf5R2_0),.dout(w_dff_B_aHDWCnpi6_0),.clk(gclk));
	jdff dff_B_r5P8x6jF2_0(.din(w_dff_B_aHDWCnpi6_0),.dout(w_dff_B_r5P8x6jF2_0),.clk(gclk));
	jdff dff_B_zb1bl7zN4_0(.din(w_dff_B_r5P8x6jF2_0),.dout(w_dff_B_zb1bl7zN4_0),.clk(gclk));
	jdff dff_B_cidGYdUa6_0(.din(w_dff_B_zb1bl7zN4_0),.dout(w_dff_B_cidGYdUa6_0),.clk(gclk));
	jdff dff_B_SQmXewmR4_0(.din(w_dff_B_cidGYdUa6_0),.dout(w_dff_B_SQmXewmR4_0),.clk(gclk));
	jdff dff_B_f8qTgXte9_1(.din(n1110),.dout(w_dff_B_f8qTgXte9_1),.clk(gclk));
	jdff dff_B_wA3ayJKz9_1(.din(w_dff_B_f8qTgXte9_1),.dout(w_dff_B_wA3ayJKz9_1),.clk(gclk));
	jdff dff_B_WyYKA7pW5_1(.din(w_dff_B_wA3ayJKz9_1),.dout(w_dff_B_WyYKA7pW5_1),.clk(gclk));
	jdff dff_B_DAvIUI0Y4_1(.din(w_dff_B_WyYKA7pW5_1),.dout(w_dff_B_DAvIUI0Y4_1),.clk(gclk));
	jdff dff_B_NMD9kh3O2_1(.din(w_dff_B_DAvIUI0Y4_1),.dout(w_dff_B_NMD9kh3O2_1),.clk(gclk));
	jdff dff_B_eqxDkH0O8_1(.din(w_dff_B_NMD9kh3O2_1),.dout(w_dff_B_eqxDkH0O8_1),.clk(gclk));
	jdff dff_B_QNlR3t9x8_1(.din(w_dff_B_eqxDkH0O8_1),.dout(w_dff_B_QNlR3t9x8_1),.clk(gclk));
	jdff dff_B_Pi83P7Jj1_1(.din(w_dff_B_QNlR3t9x8_1),.dout(w_dff_B_Pi83P7Jj1_1),.clk(gclk));
	jdff dff_B_yLelrGJg4_1(.din(w_dff_B_Pi83P7Jj1_1),.dout(w_dff_B_yLelrGJg4_1),.clk(gclk));
	jdff dff_B_265rvvmm7_1(.din(w_dff_B_yLelrGJg4_1),.dout(w_dff_B_265rvvmm7_1),.clk(gclk));
	jdff dff_B_VIpU8MEZ7_1(.din(w_dff_B_265rvvmm7_1),.dout(w_dff_B_VIpU8MEZ7_1),.clk(gclk));
	jdff dff_B_IR4m8D4z1_1(.din(w_dff_B_VIpU8MEZ7_1),.dout(w_dff_B_IR4m8D4z1_1),.clk(gclk));
	jdff dff_B_kR8xyHfm8_1(.din(w_dff_B_IR4m8D4z1_1),.dout(w_dff_B_kR8xyHfm8_1),.clk(gclk));
	jdff dff_B_xJsZXO0B1_1(.din(w_dff_B_kR8xyHfm8_1),.dout(w_dff_B_xJsZXO0B1_1),.clk(gclk));
	jdff dff_B_d532XBxq9_1(.din(w_dff_B_xJsZXO0B1_1),.dout(w_dff_B_d532XBxq9_1),.clk(gclk));
	jdff dff_B_lBPAWRUn6_1(.din(w_dff_B_d532XBxq9_1),.dout(w_dff_B_lBPAWRUn6_1),.clk(gclk));
	jdff dff_B_lAZCmoHB9_1(.din(w_dff_B_lBPAWRUn6_1),.dout(w_dff_B_lAZCmoHB9_1),.clk(gclk));
	jdff dff_B_s2oQhqpx5_1(.din(w_dff_B_lAZCmoHB9_1),.dout(w_dff_B_s2oQhqpx5_1),.clk(gclk));
	jdff dff_B_LwVyTjA67_1(.din(w_dff_B_s2oQhqpx5_1),.dout(w_dff_B_LwVyTjA67_1),.clk(gclk));
	jdff dff_B_KxcTmLCk6_1(.din(w_dff_B_LwVyTjA67_1),.dout(w_dff_B_KxcTmLCk6_1),.clk(gclk));
	jdff dff_B_ojx8xbw63_1(.din(w_dff_B_KxcTmLCk6_1),.dout(w_dff_B_ojx8xbw63_1),.clk(gclk));
	jdff dff_B_pxnZdb897_1(.din(w_dff_B_ojx8xbw63_1),.dout(w_dff_B_pxnZdb897_1),.clk(gclk));
	jdff dff_B_yrZG7lNJ0_1(.din(w_dff_B_pxnZdb897_1),.dout(w_dff_B_yrZG7lNJ0_1),.clk(gclk));
	jdff dff_B_pXzA0Phq4_1(.din(w_dff_B_yrZG7lNJ0_1),.dout(w_dff_B_pXzA0Phq4_1),.clk(gclk));
	jdff dff_B_FyDdRiCH4_1(.din(w_dff_B_pXzA0Phq4_1),.dout(w_dff_B_FyDdRiCH4_1),.clk(gclk));
	jdff dff_B_GsYgYjUL2_1(.din(w_dff_B_FyDdRiCH4_1),.dout(w_dff_B_GsYgYjUL2_1),.clk(gclk));
	jdff dff_B_Y6rFuYd22_1(.din(w_dff_B_GsYgYjUL2_1),.dout(w_dff_B_Y6rFuYd22_1),.clk(gclk));
	jdff dff_B_dcMSza5I3_1(.din(w_dff_B_Y6rFuYd22_1),.dout(w_dff_B_dcMSza5I3_1),.clk(gclk));
	jdff dff_B_6kx3AJcv9_1(.din(w_dff_B_dcMSza5I3_1),.dout(w_dff_B_6kx3AJcv9_1),.clk(gclk));
	jdff dff_B_b3YpRzjt5_1(.din(w_dff_B_6kx3AJcv9_1),.dout(w_dff_B_b3YpRzjt5_1),.clk(gclk));
	jdff dff_B_oUWhOode7_1(.din(w_dff_B_b3YpRzjt5_1),.dout(w_dff_B_oUWhOode7_1),.clk(gclk));
	jdff dff_B_wjF3NDpp9_1(.din(w_dff_B_oUWhOode7_1),.dout(w_dff_B_wjF3NDpp9_1),.clk(gclk));
	jdff dff_B_6gLk7Eoc2_1(.din(w_dff_B_wjF3NDpp9_1),.dout(w_dff_B_6gLk7Eoc2_1),.clk(gclk));
	jdff dff_B_eFZlryEr7_1(.din(w_dff_B_6gLk7Eoc2_1),.dout(w_dff_B_eFZlryEr7_1),.clk(gclk));
	jdff dff_B_Wj3Se4Si7_1(.din(w_dff_B_eFZlryEr7_1),.dout(w_dff_B_Wj3Se4Si7_1),.clk(gclk));
	jdff dff_B_6C6wDDRI7_1(.din(w_dff_B_Wj3Se4Si7_1),.dout(w_dff_B_6C6wDDRI7_1),.clk(gclk));
	jdff dff_B_ULOEeAsr5_1(.din(w_dff_B_6C6wDDRI7_1),.dout(w_dff_B_ULOEeAsr5_1),.clk(gclk));
	jdff dff_B_dhJpIDDa4_1(.din(w_dff_B_ULOEeAsr5_1),.dout(w_dff_B_dhJpIDDa4_1),.clk(gclk));
	jdff dff_B_z7DTt5rD6_1(.din(w_dff_B_dhJpIDDa4_1),.dout(w_dff_B_z7DTt5rD6_1),.clk(gclk));
	jdff dff_B_KlTVUsek4_1(.din(w_dff_B_z7DTt5rD6_1),.dout(w_dff_B_KlTVUsek4_1),.clk(gclk));
	jdff dff_B_cBByDh8p3_1(.din(w_dff_B_KlTVUsek4_1),.dout(w_dff_B_cBByDh8p3_1),.clk(gclk));
	jdff dff_B_2z1bpdKs2_1(.din(w_dff_B_cBByDh8p3_1),.dout(w_dff_B_2z1bpdKs2_1),.clk(gclk));
	jdff dff_B_z7AfpNzJ1_1(.din(w_dff_B_2z1bpdKs2_1),.dout(w_dff_B_z7AfpNzJ1_1),.clk(gclk));
	jdff dff_B_Za6DAwDP4_1(.din(w_dff_B_z7AfpNzJ1_1),.dout(w_dff_B_Za6DAwDP4_1),.clk(gclk));
	jdff dff_B_rLMbyeqU8_1(.din(w_dff_B_Za6DAwDP4_1),.dout(w_dff_B_rLMbyeqU8_1),.clk(gclk));
	jdff dff_B_fhjaWZTg6_1(.din(w_dff_B_rLMbyeqU8_1),.dout(w_dff_B_fhjaWZTg6_1),.clk(gclk));
	jdff dff_B_7jtK5JmY3_1(.din(w_dff_B_fhjaWZTg6_1),.dout(w_dff_B_7jtK5JmY3_1),.clk(gclk));
	jdff dff_B_omyDYBd36_1(.din(w_dff_B_7jtK5JmY3_1),.dout(w_dff_B_omyDYBd36_1),.clk(gclk));
	jdff dff_B_hnAAJgEf7_1(.din(w_dff_B_omyDYBd36_1),.dout(w_dff_B_hnAAJgEf7_1),.clk(gclk));
	jdff dff_B_QoQ55iHQ4_1(.din(w_dff_B_hnAAJgEf7_1),.dout(w_dff_B_QoQ55iHQ4_1),.clk(gclk));
	jdff dff_B_E5bJ3CFB0_1(.din(w_dff_B_QoQ55iHQ4_1),.dout(w_dff_B_E5bJ3CFB0_1),.clk(gclk));
	jdff dff_B_mOjoM2Lg9_1(.din(w_dff_B_E5bJ3CFB0_1),.dout(w_dff_B_mOjoM2Lg9_1),.clk(gclk));
	jdff dff_B_DQsGlLso2_1(.din(w_dff_B_mOjoM2Lg9_1),.dout(w_dff_B_DQsGlLso2_1),.clk(gclk));
	jdff dff_B_Cdfil6tL6_1(.din(w_dff_B_DQsGlLso2_1),.dout(w_dff_B_Cdfil6tL6_1),.clk(gclk));
	jdff dff_B_o8JT9GyU6_1(.din(w_dff_B_Cdfil6tL6_1),.dout(w_dff_B_o8JT9GyU6_1),.clk(gclk));
	jdff dff_B_6bKoZvuP1_1(.din(w_dff_B_o8JT9GyU6_1),.dout(w_dff_B_6bKoZvuP1_1),.clk(gclk));
	jdff dff_B_PxObT3Vs6_1(.din(w_dff_B_6bKoZvuP1_1),.dout(w_dff_B_PxObT3Vs6_1),.clk(gclk));
	jdff dff_B_3dBdoVri1_1(.din(w_dff_B_PxObT3Vs6_1),.dout(w_dff_B_3dBdoVri1_1),.clk(gclk));
	jdff dff_B_vBOC7GO92_1(.din(w_dff_B_3dBdoVri1_1),.dout(w_dff_B_vBOC7GO92_1),.clk(gclk));
	jdff dff_B_IFAYAUit5_1(.din(w_dff_B_vBOC7GO92_1),.dout(w_dff_B_IFAYAUit5_1),.clk(gclk));
	jdff dff_B_yXVD7yRc9_1(.din(w_dff_B_IFAYAUit5_1),.dout(w_dff_B_yXVD7yRc9_1),.clk(gclk));
	jdff dff_B_U7bVR98W5_1(.din(w_dff_B_yXVD7yRc9_1),.dout(w_dff_B_U7bVR98W5_1),.clk(gclk));
	jdff dff_B_unEQqwuE6_1(.din(w_dff_B_U7bVR98W5_1),.dout(w_dff_B_unEQqwuE6_1),.clk(gclk));
	jdff dff_B_d8TCTVuy2_1(.din(w_dff_B_unEQqwuE6_1),.dout(w_dff_B_d8TCTVuy2_1),.clk(gclk));
	jdff dff_B_ET6JeDMn7_1(.din(w_dff_B_d8TCTVuy2_1),.dout(w_dff_B_ET6JeDMn7_1),.clk(gclk));
	jdff dff_B_wDNmYvA14_1(.din(w_dff_B_ET6JeDMn7_1),.dout(w_dff_B_wDNmYvA14_1),.clk(gclk));
	jdff dff_B_xt6JAc2B0_1(.din(w_dff_B_wDNmYvA14_1),.dout(w_dff_B_xt6JAc2B0_1),.clk(gclk));
	jdff dff_B_60AoPMW41_1(.din(w_dff_B_xt6JAc2B0_1),.dout(w_dff_B_60AoPMW41_1),.clk(gclk));
	jdff dff_B_t8sMV8DN2_1(.din(w_dff_B_60AoPMW41_1),.dout(w_dff_B_t8sMV8DN2_1),.clk(gclk));
	jdff dff_B_R85AbA0R6_1(.din(w_dff_B_t8sMV8DN2_1),.dout(w_dff_B_R85AbA0R6_1),.clk(gclk));
	jdff dff_B_HIYxCD2f2_1(.din(w_dff_B_R85AbA0R6_1),.dout(w_dff_B_HIYxCD2f2_1),.clk(gclk));
	jdff dff_B_B2eYx8Q56_1(.din(w_dff_B_HIYxCD2f2_1),.dout(w_dff_B_B2eYx8Q56_1),.clk(gclk));
	jdff dff_B_uf7oa47w9_1(.din(w_dff_B_B2eYx8Q56_1),.dout(w_dff_B_uf7oa47w9_1),.clk(gclk));
	jdff dff_B_YPJ9nDUz1_1(.din(w_dff_B_uf7oa47w9_1),.dout(w_dff_B_YPJ9nDUz1_1),.clk(gclk));
	jdff dff_B_nMc59K3H8_1(.din(w_dff_B_YPJ9nDUz1_1),.dout(w_dff_B_nMc59K3H8_1),.clk(gclk));
	jdff dff_B_bCwx0H6p0_1(.din(w_dff_B_nMc59K3H8_1),.dout(w_dff_B_bCwx0H6p0_1),.clk(gclk));
	jdff dff_B_gu03SAMI3_1(.din(w_dff_B_bCwx0H6p0_1),.dout(w_dff_B_gu03SAMI3_1),.clk(gclk));
	jdff dff_B_zt312RzB2_1(.din(w_dff_B_gu03SAMI3_1),.dout(w_dff_B_zt312RzB2_1),.clk(gclk));
	jdff dff_B_UM1NDhb67_1(.din(w_dff_B_zt312RzB2_1),.dout(w_dff_B_UM1NDhb67_1),.clk(gclk));
	jdff dff_B_hYu6J6jU6_1(.din(w_dff_B_UM1NDhb67_1),.dout(w_dff_B_hYu6J6jU6_1),.clk(gclk));
	jdff dff_B_mhyCqDbY7_1(.din(w_dff_B_hYu6J6jU6_1),.dout(w_dff_B_mhyCqDbY7_1),.clk(gclk));
	jdff dff_B_FRFxtHCR1_1(.din(w_dff_B_mhyCqDbY7_1),.dout(w_dff_B_FRFxtHCR1_1),.clk(gclk));
	jdff dff_B_VuOuJlF88_1(.din(w_dff_B_FRFxtHCR1_1),.dout(w_dff_B_VuOuJlF88_1),.clk(gclk));
	jdff dff_B_17FqGLs39_1(.din(w_dff_B_VuOuJlF88_1),.dout(w_dff_B_17FqGLs39_1),.clk(gclk));
	jdff dff_B_OOADEoCA0_1(.din(w_dff_B_17FqGLs39_1),.dout(w_dff_B_OOADEoCA0_1),.clk(gclk));
	jdff dff_B_x4DAf78o5_1(.din(w_dff_B_OOADEoCA0_1),.dout(w_dff_B_x4DAf78o5_1),.clk(gclk));
	jdff dff_B_ATNpuaLy3_1(.din(w_dff_B_x4DAf78o5_1),.dout(w_dff_B_ATNpuaLy3_1),.clk(gclk));
	jdff dff_B_pCOqBZ5a6_1(.din(w_dff_B_ATNpuaLy3_1),.dout(w_dff_B_pCOqBZ5a6_1),.clk(gclk));
	jdff dff_B_7JFpEUAY0_1(.din(w_dff_B_pCOqBZ5a6_1),.dout(w_dff_B_7JFpEUAY0_1),.clk(gclk));
	jdff dff_B_oZIYArVl3_1(.din(w_dff_B_7JFpEUAY0_1),.dout(w_dff_B_oZIYArVl3_1),.clk(gclk));
	jdff dff_B_D8FKC54r8_1(.din(w_dff_B_oZIYArVl3_1),.dout(w_dff_B_D8FKC54r8_1),.clk(gclk));
	jdff dff_B_5f3WTAVR3_1(.din(w_dff_B_D8FKC54r8_1),.dout(w_dff_B_5f3WTAVR3_1),.clk(gclk));
	jdff dff_B_qkFObSEu1_1(.din(w_dff_B_5f3WTAVR3_1),.dout(w_dff_B_qkFObSEu1_1),.clk(gclk));
	jdff dff_B_oGDOMs2B4_1(.din(w_dff_B_qkFObSEu1_1),.dout(w_dff_B_oGDOMs2B4_1),.clk(gclk));
	jdff dff_B_QvyQniSd7_1(.din(w_dff_B_oGDOMs2B4_1),.dout(w_dff_B_QvyQniSd7_1),.clk(gclk));
	jdff dff_B_yLWVVCBF6_1(.din(w_dff_B_QvyQniSd7_1),.dout(w_dff_B_yLWVVCBF6_1),.clk(gclk));
	jdff dff_B_RJLZJt0h9_1(.din(w_dff_B_yLWVVCBF6_1),.dout(w_dff_B_RJLZJt0h9_1),.clk(gclk));
	jdff dff_B_N1hPepM65_1(.din(w_dff_B_RJLZJt0h9_1),.dout(w_dff_B_N1hPepM65_1),.clk(gclk));
	jdff dff_B_0OGwauoM3_1(.din(w_dff_B_N1hPepM65_1),.dout(w_dff_B_0OGwauoM3_1),.clk(gclk));
	jdff dff_B_PnYoe6II7_1(.din(w_dff_B_0OGwauoM3_1),.dout(w_dff_B_PnYoe6II7_1),.clk(gclk));
	jdff dff_B_SCCLtmRc5_1(.din(w_dff_B_PnYoe6II7_1),.dout(w_dff_B_SCCLtmRc5_1),.clk(gclk));
	jdff dff_B_zEYqtAP65_1(.din(w_dff_B_SCCLtmRc5_1),.dout(w_dff_B_zEYqtAP65_1),.clk(gclk));
	jdff dff_B_AMsAyZTz4_1(.din(w_dff_B_zEYqtAP65_1),.dout(w_dff_B_AMsAyZTz4_1),.clk(gclk));
	jdff dff_B_oi0tPcgv1_1(.din(w_dff_B_AMsAyZTz4_1),.dout(w_dff_B_oi0tPcgv1_1),.clk(gclk));
	jdff dff_B_IGwUYizm5_1(.din(w_dff_B_oi0tPcgv1_1),.dout(w_dff_B_IGwUYizm5_1),.clk(gclk));
	jdff dff_B_vP1BvdZd9_1(.din(w_dff_B_IGwUYizm5_1),.dout(w_dff_B_vP1BvdZd9_1),.clk(gclk));
	jdff dff_B_nSQTaVBp1_1(.din(w_dff_B_vP1BvdZd9_1),.dout(w_dff_B_nSQTaVBp1_1),.clk(gclk));
	jdff dff_B_yVI5i3fN6_1(.din(w_dff_B_nSQTaVBp1_1),.dout(w_dff_B_yVI5i3fN6_1),.clk(gclk));
	jdff dff_B_B88AtstK2_1(.din(w_dff_B_yVI5i3fN6_1),.dout(w_dff_B_B88AtstK2_1),.clk(gclk));
	jdff dff_B_Tc3infSS9_1(.din(w_dff_B_B88AtstK2_1),.dout(w_dff_B_Tc3infSS9_1),.clk(gclk));
	jdff dff_B_BM859FES4_1(.din(w_dff_B_Tc3infSS9_1),.dout(w_dff_B_BM859FES4_1),.clk(gclk));
	jdff dff_B_3BFB0Ztv8_1(.din(w_dff_B_BM859FES4_1),.dout(w_dff_B_3BFB0Ztv8_1),.clk(gclk));
	jdff dff_B_SM8s8saF5_1(.din(w_dff_B_3BFB0Ztv8_1),.dout(w_dff_B_SM8s8saF5_1),.clk(gclk));
	jdff dff_B_sICl1CVE1_1(.din(w_dff_B_SM8s8saF5_1),.dout(w_dff_B_sICl1CVE1_1),.clk(gclk));
	jdff dff_B_DSAnUEkB6_1(.din(w_dff_B_sICl1CVE1_1),.dout(w_dff_B_DSAnUEkB6_1),.clk(gclk));
	jdff dff_B_ComdkNfQ3_1(.din(w_dff_B_DSAnUEkB6_1),.dout(w_dff_B_ComdkNfQ3_1),.clk(gclk));
	jdff dff_B_XXu7XgUA8_1(.din(w_dff_B_ComdkNfQ3_1),.dout(w_dff_B_XXu7XgUA8_1),.clk(gclk));
	jdff dff_B_9RfZLfa71_1(.din(w_dff_B_XXu7XgUA8_1),.dout(w_dff_B_9RfZLfa71_1),.clk(gclk));
	jdff dff_B_ksM03QlX8_1(.din(w_dff_B_9RfZLfa71_1),.dout(w_dff_B_ksM03QlX8_1),.clk(gclk));
	jdff dff_B_MPBIqVyH9_1(.din(w_dff_B_ksM03QlX8_1),.dout(w_dff_B_MPBIqVyH9_1),.clk(gclk));
	jdff dff_B_OendyP6K5_1(.din(w_dff_B_MPBIqVyH9_1),.dout(w_dff_B_OendyP6K5_1),.clk(gclk));
	jdff dff_B_tM9vMwNR4_0(.din(n1111),.dout(w_dff_B_tM9vMwNR4_0),.clk(gclk));
	jdff dff_B_uhfXwzUK0_0(.din(w_dff_B_tM9vMwNR4_0),.dout(w_dff_B_uhfXwzUK0_0),.clk(gclk));
	jdff dff_B_XHOQ2RTY8_0(.din(w_dff_B_uhfXwzUK0_0),.dout(w_dff_B_XHOQ2RTY8_0),.clk(gclk));
	jdff dff_B_73KsFIbG8_0(.din(w_dff_B_XHOQ2RTY8_0),.dout(w_dff_B_73KsFIbG8_0),.clk(gclk));
	jdff dff_B_SxANcsW96_0(.din(w_dff_B_73KsFIbG8_0),.dout(w_dff_B_SxANcsW96_0),.clk(gclk));
	jdff dff_B_ppFd768R0_0(.din(w_dff_B_SxANcsW96_0),.dout(w_dff_B_ppFd768R0_0),.clk(gclk));
	jdff dff_B_lpXl7YPL9_0(.din(w_dff_B_ppFd768R0_0),.dout(w_dff_B_lpXl7YPL9_0),.clk(gclk));
	jdff dff_B_J9MsiBFx0_0(.din(w_dff_B_lpXl7YPL9_0),.dout(w_dff_B_J9MsiBFx0_0),.clk(gclk));
	jdff dff_B_C60neQfg4_0(.din(w_dff_B_J9MsiBFx0_0),.dout(w_dff_B_C60neQfg4_0),.clk(gclk));
	jdff dff_B_NgVd2CZr6_0(.din(w_dff_B_C60neQfg4_0),.dout(w_dff_B_NgVd2CZr6_0),.clk(gclk));
	jdff dff_B_2JwzRc4A8_0(.din(w_dff_B_NgVd2CZr6_0),.dout(w_dff_B_2JwzRc4A8_0),.clk(gclk));
	jdff dff_B_w5pizpHP7_0(.din(w_dff_B_2JwzRc4A8_0),.dout(w_dff_B_w5pizpHP7_0),.clk(gclk));
	jdff dff_B_EuSPMpIl3_0(.din(w_dff_B_w5pizpHP7_0),.dout(w_dff_B_EuSPMpIl3_0),.clk(gclk));
	jdff dff_B_um4AIsXm5_0(.din(w_dff_B_EuSPMpIl3_0),.dout(w_dff_B_um4AIsXm5_0),.clk(gclk));
	jdff dff_B_6MmOjB9R5_0(.din(w_dff_B_um4AIsXm5_0),.dout(w_dff_B_6MmOjB9R5_0),.clk(gclk));
	jdff dff_B_9XSbfqsG5_0(.din(w_dff_B_6MmOjB9R5_0),.dout(w_dff_B_9XSbfqsG5_0),.clk(gclk));
	jdff dff_B_Bp5qn2KU0_0(.din(w_dff_B_9XSbfqsG5_0),.dout(w_dff_B_Bp5qn2KU0_0),.clk(gclk));
	jdff dff_B_Kh6MxY7r6_0(.din(w_dff_B_Bp5qn2KU0_0),.dout(w_dff_B_Kh6MxY7r6_0),.clk(gclk));
	jdff dff_B_Sqbvxk8B1_0(.din(w_dff_B_Kh6MxY7r6_0),.dout(w_dff_B_Sqbvxk8B1_0),.clk(gclk));
	jdff dff_B_GhAuJcPK3_0(.din(w_dff_B_Sqbvxk8B1_0),.dout(w_dff_B_GhAuJcPK3_0),.clk(gclk));
	jdff dff_B_BulXm3oD5_0(.din(w_dff_B_GhAuJcPK3_0),.dout(w_dff_B_BulXm3oD5_0),.clk(gclk));
	jdff dff_B_UtNuC4Me2_0(.din(w_dff_B_BulXm3oD5_0),.dout(w_dff_B_UtNuC4Me2_0),.clk(gclk));
	jdff dff_B_VvVgAdlR8_0(.din(w_dff_B_UtNuC4Me2_0),.dout(w_dff_B_VvVgAdlR8_0),.clk(gclk));
	jdff dff_B_xlFP8uDR4_0(.din(w_dff_B_VvVgAdlR8_0),.dout(w_dff_B_xlFP8uDR4_0),.clk(gclk));
	jdff dff_B_MwNB2qsV2_0(.din(w_dff_B_xlFP8uDR4_0),.dout(w_dff_B_MwNB2qsV2_0),.clk(gclk));
	jdff dff_B_J9oGn0sy9_0(.din(w_dff_B_MwNB2qsV2_0),.dout(w_dff_B_J9oGn0sy9_0),.clk(gclk));
	jdff dff_B_M22xxVJq7_0(.din(w_dff_B_J9oGn0sy9_0),.dout(w_dff_B_M22xxVJq7_0),.clk(gclk));
	jdff dff_B_emQo0S9V2_0(.din(w_dff_B_M22xxVJq7_0),.dout(w_dff_B_emQo0S9V2_0),.clk(gclk));
	jdff dff_B_gj13ySDt2_0(.din(w_dff_B_emQo0S9V2_0),.dout(w_dff_B_gj13ySDt2_0),.clk(gclk));
	jdff dff_B_SdpwCDWy9_0(.din(w_dff_B_gj13ySDt2_0),.dout(w_dff_B_SdpwCDWy9_0),.clk(gclk));
	jdff dff_B_PXt43aUE0_0(.din(w_dff_B_SdpwCDWy9_0),.dout(w_dff_B_PXt43aUE0_0),.clk(gclk));
	jdff dff_B_PQZUbu0R6_0(.din(w_dff_B_PXt43aUE0_0),.dout(w_dff_B_PQZUbu0R6_0),.clk(gclk));
	jdff dff_B_okE9LWUO4_0(.din(w_dff_B_PQZUbu0R6_0),.dout(w_dff_B_okE9LWUO4_0),.clk(gclk));
	jdff dff_B_aFeTWQFj3_0(.din(w_dff_B_okE9LWUO4_0),.dout(w_dff_B_aFeTWQFj3_0),.clk(gclk));
	jdff dff_B_lGd3crRN0_0(.din(w_dff_B_aFeTWQFj3_0),.dout(w_dff_B_lGd3crRN0_0),.clk(gclk));
	jdff dff_B_03Ua75Cb7_0(.din(w_dff_B_lGd3crRN0_0),.dout(w_dff_B_03Ua75Cb7_0),.clk(gclk));
	jdff dff_B_nL371TK89_0(.din(w_dff_B_03Ua75Cb7_0),.dout(w_dff_B_nL371TK89_0),.clk(gclk));
	jdff dff_B_vMAzRO376_0(.din(w_dff_B_nL371TK89_0),.dout(w_dff_B_vMAzRO376_0),.clk(gclk));
	jdff dff_B_Sfu57Pet3_0(.din(w_dff_B_vMAzRO376_0),.dout(w_dff_B_Sfu57Pet3_0),.clk(gclk));
	jdff dff_B_Vfxkiga97_0(.din(w_dff_B_Sfu57Pet3_0),.dout(w_dff_B_Vfxkiga97_0),.clk(gclk));
	jdff dff_B_0Du4hO558_0(.din(w_dff_B_Vfxkiga97_0),.dout(w_dff_B_0Du4hO558_0),.clk(gclk));
	jdff dff_B_FQwcILQr1_0(.din(w_dff_B_0Du4hO558_0),.dout(w_dff_B_FQwcILQr1_0),.clk(gclk));
	jdff dff_B_7deU1YPm7_0(.din(w_dff_B_FQwcILQr1_0),.dout(w_dff_B_7deU1YPm7_0),.clk(gclk));
	jdff dff_B_U6WaxnyG7_0(.din(w_dff_B_7deU1YPm7_0),.dout(w_dff_B_U6WaxnyG7_0),.clk(gclk));
	jdff dff_B_IE4XmMqO1_0(.din(w_dff_B_U6WaxnyG7_0),.dout(w_dff_B_IE4XmMqO1_0),.clk(gclk));
	jdff dff_B_XIDhGfYe4_0(.din(w_dff_B_IE4XmMqO1_0),.dout(w_dff_B_XIDhGfYe4_0),.clk(gclk));
	jdff dff_B_BbSW8EG01_0(.din(w_dff_B_XIDhGfYe4_0),.dout(w_dff_B_BbSW8EG01_0),.clk(gclk));
	jdff dff_B_01j2suE16_0(.din(w_dff_B_BbSW8EG01_0),.dout(w_dff_B_01j2suE16_0),.clk(gclk));
	jdff dff_B_ZQNxCRW28_0(.din(w_dff_B_01j2suE16_0),.dout(w_dff_B_ZQNxCRW28_0),.clk(gclk));
	jdff dff_B_qs0z4ASg3_0(.din(w_dff_B_ZQNxCRW28_0),.dout(w_dff_B_qs0z4ASg3_0),.clk(gclk));
	jdff dff_B_Hb5oaEBn9_0(.din(w_dff_B_qs0z4ASg3_0),.dout(w_dff_B_Hb5oaEBn9_0),.clk(gclk));
	jdff dff_B_aIXkLAfO7_0(.din(w_dff_B_Hb5oaEBn9_0),.dout(w_dff_B_aIXkLAfO7_0),.clk(gclk));
	jdff dff_B_hzIHzoj10_0(.din(w_dff_B_aIXkLAfO7_0),.dout(w_dff_B_hzIHzoj10_0),.clk(gclk));
	jdff dff_B_S9no621i9_0(.din(w_dff_B_hzIHzoj10_0),.dout(w_dff_B_S9no621i9_0),.clk(gclk));
	jdff dff_B_zdSxhAjc0_0(.din(w_dff_B_S9no621i9_0),.dout(w_dff_B_zdSxhAjc0_0),.clk(gclk));
	jdff dff_B_Ihpyj1898_0(.din(w_dff_B_zdSxhAjc0_0),.dout(w_dff_B_Ihpyj1898_0),.clk(gclk));
	jdff dff_B_djmgujPx9_0(.din(w_dff_B_Ihpyj1898_0),.dout(w_dff_B_djmgujPx9_0),.clk(gclk));
	jdff dff_B_HHXF1L2n9_0(.din(w_dff_B_djmgujPx9_0),.dout(w_dff_B_HHXF1L2n9_0),.clk(gclk));
	jdff dff_B_pfSse2or9_0(.din(w_dff_B_HHXF1L2n9_0),.dout(w_dff_B_pfSse2or9_0),.clk(gclk));
	jdff dff_B_yoLIBYJa9_0(.din(w_dff_B_pfSse2or9_0),.dout(w_dff_B_yoLIBYJa9_0),.clk(gclk));
	jdff dff_B_t3JcdQsG3_0(.din(w_dff_B_yoLIBYJa9_0),.dout(w_dff_B_t3JcdQsG3_0),.clk(gclk));
	jdff dff_B_s6VMMbPr3_0(.din(w_dff_B_t3JcdQsG3_0),.dout(w_dff_B_s6VMMbPr3_0),.clk(gclk));
	jdff dff_B_ZrFR8mMC6_0(.din(w_dff_B_s6VMMbPr3_0),.dout(w_dff_B_ZrFR8mMC6_0),.clk(gclk));
	jdff dff_B_bd95D6VF7_0(.din(w_dff_B_ZrFR8mMC6_0),.dout(w_dff_B_bd95D6VF7_0),.clk(gclk));
	jdff dff_B_VOdgSkbG9_0(.din(w_dff_B_bd95D6VF7_0),.dout(w_dff_B_VOdgSkbG9_0),.clk(gclk));
	jdff dff_B_ghxMdhcM0_0(.din(w_dff_B_VOdgSkbG9_0),.dout(w_dff_B_ghxMdhcM0_0),.clk(gclk));
	jdff dff_B_Oa236skM5_0(.din(w_dff_B_ghxMdhcM0_0),.dout(w_dff_B_Oa236skM5_0),.clk(gclk));
	jdff dff_B_VA5Wc4EH5_0(.din(w_dff_B_Oa236skM5_0),.dout(w_dff_B_VA5Wc4EH5_0),.clk(gclk));
	jdff dff_B_LpvTUo541_0(.din(w_dff_B_VA5Wc4EH5_0),.dout(w_dff_B_LpvTUo541_0),.clk(gclk));
	jdff dff_B_1BZtxsHt4_0(.din(w_dff_B_LpvTUo541_0),.dout(w_dff_B_1BZtxsHt4_0),.clk(gclk));
	jdff dff_B_4nt7qEs50_0(.din(w_dff_B_1BZtxsHt4_0),.dout(w_dff_B_4nt7qEs50_0),.clk(gclk));
	jdff dff_B_0aC17Nfq2_0(.din(w_dff_B_4nt7qEs50_0),.dout(w_dff_B_0aC17Nfq2_0),.clk(gclk));
	jdff dff_B_DiQQ739I5_0(.din(w_dff_B_0aC17Nfq2_0),.dout(w_dff_B_DiQQ739I5_0),.clk(gclk));
	jdff dff_B_6ecbn7gn4_0(.din(w_dff_B_DiQQ739I5_0),.dout(w_dff_B_6ecbn7gn4_0),.clk(gclk));
	jdff dff_B_lMrzd39c6_0(.din(w_dff_B_6ecbn7gn4_0),.dout(w_dff_B_lMrzd39c6_0),.clk(gclk));
	jdff dff_B_1DV4jHEs3_0(.din(w_dff_B_lMrzd39c6_0),.dout(w_dff_B_1DV4jHEs3_0),.clk(gclk));
	jdff dff_B_nBgWTI0J3_0(.din(w_dff_B_1DV4jHEs3_0),.dout(w_dff_B_nBgWTI0J3_0),.clk(gclk));
	jdff dff_B_OhnaNYWH1_0(.din(w_dff_B_nBgWTI0J3_0),.dout(w_dff_B_OhnaNYWH1_0),.clk(gclk));
	jdff dff_B_64tDrTxv7_0(.din(w_dff_B_OhnaNYWH1_0),.dout(w_dff_B_64tDrTxv7_0),.clk(gclk));
	jdff dff_B_2LR4zyBv1_0(.din(w_dff_B_64tDrTxv7_0),.dout(w_dff_B_2LR4zyBv1_0),.clk(gclk));
	jdff dff_B_K8ptnSmK4_0(.din(w_dff_B_2LR4zyBv1_0),.dout(w_dff_B_K8ptnSmK4_0),.clk(gclk));
	jdff dff_B_LwH556Dk7_0(.din(w_dff_B_K8ptnSmK4_0),.dout(w_dff_B_LwH556Dk7_0),.clk(gclk));
	jdff dff_B_z0aXwVt17_0(.din(w_dff_B_LwH556Dk7_0),.dout(w_dff_B_z0aXwVt17_0),.clk(gclk));
	jdff dff_B_tDRux8yC0_0(.din(w_dff_B_z0aXwVt17_0),.dout(w_dff_B_tDRux8yC0_0),.clk(gclk));
	jdff dff_B_GM9gKOZD0_0(.din(w_dff_B_tDRux8yC0_0),.dout(w_dff_B_GM9gKOZD0_0),.clk(gclk));
	jdff dff_B_ICeIw2zD9_0(.din(w_dff_B_GM9gKOZD0_0),.dout(w_dff_B_ICeIw2zD9_0),.clk(gclk));
	jdff dff_B_DvyPNxlV8_0(.din(w_dff_B_ICeIw2zD9_0),.dout(w_dff_B_DvyPNxlV8_0),.clk(gclk));
	jdff dff_B_4awwGqWm6_0(.din(w_dff_B_DvyPNxlV8_0),.dout(w_dff_B_4awwGqWm6_0),.clk(gclk));
	jdff dff_B_wmcfKzZl8_0(.din(w_dff_B_4awwGqWm6_0),.dout(w_dff_B_wmcfKzZl8_0),.clk(gclk));
	jdff dff_B_2TFoYEKO8_0(.din(w_dff_B_wmcfKzZl8_0),.dout(w_dff_B_2TFoYEKO8_0),.clk(gclk));
	jdff dff_B_PQZmsKa46_0(.din(w_dff_B_2TFoYEKO8_0),.dout(w_dff_B_PQZmsKa46_0),.clk(gclk));
	jdff dff_B_n73NktSA9_0(.din(w_dff_B_PQZmsKa46_0),.dout(w_dff_B_n73NktSA9_0),.clk(gclk));
	jdff dff_B_50ryWj8f7_0(.din(w_dff_B_n73NktSA9_0),.dout(w_dff_B_50ryWj8f7_0),.clk(gclk));
	jdff dff_B_e8KebvRU4_0(.din(w_dff_B_50ryWj8f7_0),.dout(w_dff_B_e8KebvRU4_0),.clk(gclk));
	jdff dff_B_HoUCemaA0_0(.din(w_dff_B_e8KebvRU4_0),.dout(w_dff_B_HoUCemaA0_0),.clk(gclk));
	jdff dff_B_YrOPCbeR4_0(.din(w_dff_B_HoUCemaA0_0),.dout(w_dff_B_YrOPCbeR4_0),.clk(gclk));
	jdff dff_B_WDW6ZdUQ4_0(.din(w_dff_B_YrOPCbeR4_0),.dout(w_dff_B_WDW6ZdUQ4_0),.clk(gclk));
	jdff dff_B_yjJ4ndBe6_0(.din(w_dff_B_WDW6ZdUQ4_0),.dout(w_dff_B_yjJ4ndBe6_0),.clk(gclk));
	jdff dff_B_kPdv9fzy6_0(.din(w_dff_B_yjJ4ndBe6_0),.dout(w_dff_B_kPdv9fzy6_0),.clk(gclk));
	jdff dff_B_ZQHcXbS85_0(.din(w_dff_B_kPdv9fzy6_0),.dout(w_dff_B_ZQHcXbS85_0),.clk(gclk));
	jdff dff_B_XgwZm5Cj9_0(.din(w_dff_B_ZQHcXbS85_0),.dout(w_dff_B_XgwZm5Cj9_0),.clk(gclk));
	jdff dff_B_uClfECq68_0(.din(w_dff_B_XgwZm5Cj9_0),.dout(w_dff_B_uClfECq68_0),.clk(gclk));
	jdff dff_B_MTcd4K5W2_0(.din(w_dff_B_uClfECq68_0),.dout(w_dff_B_MTcd4K5W2_0),.clk(gclk));
	jdff dff_B_RHYhS3Pp0_0(.din(w_dff_B_MTcd4K5W2_0),.dout(w_dff_B_RHYhS3Pp0_0),.clk(gclk));
	jdff dff_B_l6aiJ5Rp7_0(.din(w_dff_B_RHYhS3Pp0_0),.dout(w_dff_B_l6aiJ5Rp7_0),.clk(gclk));
	jdff dff_B_uRpD9wvm9_0(.din(w_dff_B_l6aiJ5Rp7_0),.dout(w_dff_B_uRpD9wvm9_0),.clk(gclk));
	jdff dff_B_189KW5Mw0_0(.din(w_dff_B_uRpD9wvm9_0),.dout(w_dff_B_189KW5Mw0_0),.clk(gclk));
	jdff dff_B_1gXPrIcA9_0(.din(w_dff_B_189KW5Mw0_0),.dout(w_dff_B_1gXPrIcA9_0),.clk(gclk));
	jdff dff_B_YJ3IFZiO7_0(.din(w_dff_B_1gXPrIcA9_0),.dout(w_dff_B_YJ3IFZiO7_0),.clk(gclk));
	jdff dff_B_PEAcNf6L2_0(.din(w_dff_B_YJ3IFZiO7_0),.dout(w_dff_B_PEAcNf6L2_0),.clk(gclk));
	jdff dff_B_brIu6GOx4_0(.din(w_dff_B_PEAcNf6L2_0),.dout(w_dff_B_brIu6GOx4_0),.clk(gclk));
	jdff dff_B_Kxq0iqGR4_0(.din(w_dff_B_brIu6GOx4_0),.dout(w_dff_B_Kxq0iqGR4_0),.clk(gclk));
	jdff dff_B_rUdkOYQS7_0(.din(w_dff_B_Kxq0iqGR4_0),.dout(w_dff_B_rUdkOYQS7_0),.clk(gclk));
	jdff dff_B_Qmh2opri7_0(.din(w_dff_B_rUdkOYQS7_0),.dout(w_dff_B_Qmh2opri7_0),.clk(gclk));
	jdff dff_B_0yt44FnY0_0(.din(w_dff_B_Qmh2opri7_0),.dout(w_dff_B_0yt44FnY0_0),.clk(gclk));
	jdff dff_B_TVVClLn13_0(.din(w_dff_B_0yt44FnY0_0),.dout(w_dff_B_TVVClLn13_0),.clk(gclk));
	jdff dff_B_dw3rFMsF8_0(.din(w_dff_B_TVVClLn13_0),.dout(w_dff_B_dw3rFMsF8_0),.clk(gclk));
	jdff dff_B_iNsE2v409_0(.din(w_dff_B_dw3rFMsF8_0),.dout(w_dff_B_iNsE2v409_0),.clk(gclk));
	jdff dff_B_QOuDUobD7_0(.din(w_dff_B_iNsE2v409_0),.dout(w_dff_B_QOuDUobD7_0),.clk(gclk));
	jdff dff_B_6CFEKehx6_0(.din(w_dff_B_QOuDUobD7_0),.dout(w_dff_B_6CFEKehx6_0),.clk(gclk));
	jdff dff_B_nEpywF7H8_0(.din(w_dff_B_6CFEKehx6_0),.dout(w_dff_B_nEpywF7H8_0),.clk(gclk));
	jdff dff_B_hcPXkUGE1_1(.din(n1104),.dout(w_dff_B_hcPXkUGE1_1),.clk(gclk));
	jdff dff_B_XavnPH2f0_1(.din(w_dff_B_hcPXkUGE1_1),.dout(w_dff_B_XavnPH2f0_1),.clk(gclk));
	jdff dff_B_NiDlEVIN3_1(.din(w_dff_B_XavnPH2f0_1),.dout(w_dff_B_NiDlEVIN3_1),.clk(gclk));
	jdff dff_B_tsdEwm0t4_1(.din(w_dff_B_NiDlEVIN3_1),.dout(w_dff_B_tsdEwm0t4_1),.clk(gclk));
	jdff dff_B_FCy9SeUg6_1(.din(w_dff_B_tsdEwm0t4_1),.dout(w_dff_B_FCy9SeUg6_1),.clk(gclk));
	jdff dff_B_0Exq71OG3_1(.din(w_dff_B_FCy9SeUg6_1),.dout(w_dff_B_0Exq71OG3_1),.clk(gclk));
	jdff dff_B_NPApAPev3_1(.din(w_dff_B_0Exq71OG3_1),.dout(w_dff_B_NPApAPev3_1),.clk(gclk));
	jdff dff_B_sBpTzv4r9_1(.din(w_dff_B_NPApAPev3_1),.dout(w_dff_B_sBpTzv4r9_1),.clk(gclk));
	jdff dff_B_G4lqCRRS9_1(.din(w_dff_B_sBpTzv4r9_1),.dout(w_dff_B_G4lqCRRS9_1),.clk(gclk));
	jdff dff_B_7IAmLvla7_1(.din(w_dff_B_G4lqCRRS9_1),.dout(w_dff_B_7IAmLvla7_1),.clk(gclk));
	jdff dff_B_GPatByqn8_1(.din(w_dff_B_7IAmLvla7_1),.dout(w_dff_B_GPatByqn8_1),.clk(gclk));
	jdff dff_B_ZKEP9MCn9_1(.din(w_dff_B_GPatByqn8_1),.dout(w_dff_B_ZKEP9MCn9_1),.clk(gclk));
	jdff dff_B_D3tTMyic2_1(.din(w_dff_B_ZKEP9MCn9_1),.dout(w_dff_B_D3tTMyic2_1),.clk(gclk));
	jdff dff_B_IBo4gq5x8_1(.din(w_dff_B_D3tTMyic2_1),.dout(w_dff_B_IBo4gq5x8_1),.clk(gclk));
	jdff dff_B_0icHqgb25_1(.din(w_dff_B_IBo4gq5x8_1),.dout(w_dff_B_0icHqgb25_1),.clk(gclk));
	jdff dff_B_n2e5uGBN9_1(.din(w_dff_B_0icHqgb25_1),.dout(w_dff_B_n2e5uGBN9_1),.clk(gclk));
	jdff dff_B_hRxZAZiG2_1(.din(w_dff_B_n2e5uGBN9_1),.dout(w_dff_B_hRxZAZiG2_1),.clk(gclk));
	jdff dff_B_Rd3qvTtt0_1(.din(w_dff_B_hRxZAZiG2_1),.dout(w_dff_B_Rd3qvTtt0_1),.clk(gclk));
	jdff dff_B_Jep5mWU60_1(.din(w_dff_B_Rd3qvTtt0_1),.dout(w_dff_B_Jep5mWU60_1),.clk(gclk));
	jdff dff_B_hZbkHOKL3_1(.din(w_dff_B_Jep5mWU60_1),.dout(w_dff_B_hZbkHOKL3_1),.clk(gclk));
	jdff dff_B_qszaWM906_1(.din(w_dff_B_hZbkHOKL3_1),.dout(w_dff_B_qszaWM906_1),.clk(gclk));
	jdff dff_B_49zXDCoS0_1(.din(w_dff_B_qszaWM906_1),.dout(w_dff_B_49zXDCoS0_1),.clk(gclk));
	jdff dff_B_7ofKzIcq7_1(.din(w_dff_B_49zXDCoS0_1),.dout(w_dff_B_7ofKzIcq7_1),.clk(gclk));
	jdff dff_B_8fFQuj1P1_1(.din(w_dff_B_7ofKzIcq7_1),.dout(w_dff_B_8fFQuj1P1_1),.clk(gclk));
	jdff dff_B_fAzq0rhf7_1(.din(w_dff_B_8fFQuj1P1_1),.dout(w_dff_B_fAzq0rhf7_1),.clk(gclk));
	jdff dff_B_ggWrBE816_1(.din(w_dff_B_fAzq0rhf7_1),.dout(w_dff_B_ggWrBE816_1),.clk(gclk));
	jdff dff_B_LfEh797H2_1(.din(w_dff_B_ggWrBE816_1),.dout(w_dff_B_LfEh797H2_1),.clk(gclk));
	jdff dff_B_veqfGzta2_1(.din(w_dff_B_LfEh797H2_1),.dout(w_dff_B_veqfGzta2_1),.clk(gclk));
	jdff dff_B_GbvyUG1R8_1(.din(w_dff_B_veqfGzta2_1),.dout(w_dff_B_GbvyUG1R8_1),.clk(gclk));
	jdff dff_B_8VBbc0aR6_1(.din(w_dff_B_GbvyUG1R8_1),.dout(w_dff_B_8VBbc0aR6_1),.clk(gclk));
	jdff dff_B_Zs2b4iHb1_1(.din(w_dff_B_8VBbc0aR6_1),.dout(w_dff_B_Zs2b4iHb1_1),.clk(gclk));
	jdff dff_B_EZVwhznK9_1(.din(w_dff_B_Zs2b4iHb1_1),.dout(w_dff_B_EZVwhznK9_1),.clk(gclk));
	jdff dff_B_PoMe8pHi9_1(.din(w_dff_B_EZVwhznK9_1),.dout(w_dff_B_PoMe8pHi9_1),.clk(gclk));
	jdff dff_B_LeNXRqvp5_1(.din(w_dff_B_PoMe8pHi9_1),.dout(w_dff_B_LeNXRqvp5_1),.clk(gclk));
	jdff dff_B_mZf2a6280_1(.din(w_dff_B_LeNXRqvp5_1),.dout(w_dff_B_mZf2a6280_1),.clk(gclk));
	jdff dff_B_WCvTiAP60_1(.din(w_dff_B_mZf2a6280_1),.dout(w_dff_B_WCvTiAP60_1),.clk(gclk));
	jdff dff_B_sbOnY7HQ4_1(.din(w_dff_B_WCvTiAP60_1),.dout(w_dff_B_sbOnY7HQ4_1),.clk(gclk));
	jdff dff_B_ZKH5Vzcn5_1(.din(w_dff_B_sbOnY7HQ4_1),.dout(w_dff_B_ZKH5Vzcn5_1),.clk(gclk));
	jdff dff_B_bntmMVLk9_1(.din(w_dff_B_ZKH5Vzcn5_1),.dout(w_dff_B_bntmMVLk9_1),.clk(gclk));
	jdff dff_B_QJYQALB37_1(.din(w_dff_B_bntmMVLk9_1),.dout(w_dff_B_QJYQALB37_1),.clk(gclk));
	jdff dff_B_meGUUGBf9_1(.din(w_dff_B_QJYQALB37_1),.dout(w_dff_B_meGUUGBf9_1),.clk(gclk));
	jdff dff_B_000zO23n4_1(.din(w_dff_B_meGUUGBf9_1),.dout(w_dff_B_000zO23n4_1),.clk(gclk));
	jdff dff_B_TBAxneeS1_1(.din(w_dff_B_000zO23n4_1),.dout(w_dff_B_TBAxneeS1_1),.clk(gclk));
	jdff dff_B_73HDM3X21_1(.din(w_dff_B_TBAxneeS1_1),.dout(w_dff_B_73HDM3X21_1),.clk(gclk));
	jdff dff_B_pknlHcXd7_1(.din(w_dff_B_73HDM3X21_1),.dout(w_dff_B_pknlHcXd7_1),.clk(gclk));
	jdff dff_B_Znt4o8t94_1(.din(w_dff_B_pknlHcXd7_1),.dout(w_dff_B_Znt4o8t94_1),.clk(gclk));
	jdff dff_B_9EbzWdIs4_1(.din(w_dff_B_Znt4o8t94_1),.dout(w_dff_B_9EbzWdIs4_1),.clk(gclk));
	jdff dff_B_ujnXSU5j3_1(.din(w_dff_B_9EbzWdIs4_1),.dout(w_dff_B_ujnXSU5j3_1),.clk(gclk));
	jdff dff_B_9v9Cnyda0_1(.din(w_dff_B_ujnXSU5j3_1),.dout(w_dff_B_9v9Cnyda0_1),.clk(gclk));
	jdff dff_B_yMQhW0og4_1(.din(w_dff_B_9v9Cnyda0_1),.dout(w_dff_B_yMQhW0og4_1),.clk(gclk));
	jdff dff_B_A97W2rSp1_1(.din(w_dff_B_yMQhW0og4_1),.dout(w_dff_B_A97W2rSp1_1),.clk(gclk));
	jdff dff_B_NNlyL4r45_1(.din(w_dff_B_A97W2rSp1_1),.dout(w_dff_B_NNlyL4r45_1),.clk(gclk));
	jdff dff_B_jb6OiXs53_1(.din(w_dff_B_NNlyL4r45_1),.dout(w_dff_B_jb6OiXs53_1),.clk(gclk));
	jdff dff_B_bh6ScHfj7_1(.din(w_dff_B_jb6OiXs53_1),.dout(w_dff_B_bh6ScHfj7_1),.clk(gclk));
	jdff dff_B_i73NuGwF8_1(.din(w_dff_B_bh6ScHfj7_1),.dout(w_dff_B_i73NuGwF8_1),.clk(gclk));
	jdff dff_B_3oSRHMcu2_1(.din(w_dff_B_i73NuGwF8_1),.dout(w_dff_B_3oSRHMcu2_1),.clk(gclk));
	jdff dff_B_MY1TNxua8_1(.din(w_dff_B_3oSRHMcu2_1),.dout(w_dff_B_MY1TNxua8_1),.clk(gclk));
	jdff dff_B_Gpy4nZj66_1(.din(w_dff_B_MY1TNxua8_1),.dout(w_dff_B_Gpy4nZj66_1),.clk(gclk));
	jdff dff_B_M8iJ3Vjo0_1(.din(w_dff_B_Gpy4nZj66_1),.dout(w_dff_B_M8iJ3Vjo0_1),.clk(gclk));
	jdff dff_B_9GKw9ZeA2_1(.din(w_dff_B_M8iJ3Vjo0_1),.dout(w_dff_B_9GKw9ZeA2_1),.clk(gclk));
	jdff dff_B_C6w6ReHm6_1(.din(w_dff_B_9GKw9ZeA2_1),.dout(w_dff_B_C6w6ReHm6_1),.clk(gclk));
	jdff dff_B_Gejv70dY2_1(.din(w_dff_B_C6w6ReHm6_1),.dout(w_dff_B_Gejv70dY2_1),.clk(gclk));
	jdff dff_B_DMNb6yXX3_1(.din(w_dff_B_Gejv70dY2_1),.dout(w_dff_B_DMNb6yXX3_1),.clk(gclk));
	jdff dff_B_iASjosPi7_1(.din(w_dff_B_DMNb6yXX3_1),.dout(w_dff_B_iASjosPi7_1),.clk(gclk));
	jdff dff_B_SqGZmNoZ8_1(.din(w_dff_B_iASjosPi7_1),.dout(w_dff_B_SqGZmNoZ8_1),.clk(gclk));
	jdff dff_B_BxmfDQnp5_1(.din(w_dff_B_SqGZmNoZ8_1),.dout(w_dff_B_BxmfDQnp5_1),.clk(gclk));
	jdff dff_B_aYsRzhlY7_1(.din(w_dff_B_BxmfDQnp5_1),.dout(w_dff_B_aYsRzhlY7_1),.clk(gclk));
	jdff dff_B_dPkQc1ws0_1(.din(w_dff_B_aYsRzhlY7_1),.dout(w_dff_B_dPkQc1ws0_1),.clk(gclk));
	jdff dff_B_6joKHa8G6_1(.din(w_dff_B_dPkQc1ws0_1),.dout(w_dff_B_6joKHa8G6_1),.clk(gclk));
	jdff dff_B_Tmao4VgQ4_1(.din(w_dff_B_6joKHa8G6_1),.dout(w_dff_B_Tmao4VgQ4_1),.clk(gclk));
	jdff dff_B_aMb3kUaa9_1(.din(w_dff_B_Tmao4VgQ4_1),.dout(w_dff_B_aMb3kUaa9_1),.clk(gclk));
	jdff dff_B_rLZvEJYF1_1(.din(w_dff_B_aMb3kUaa9_1),.dout(w_dff_B_rLZvEJYF1_1),.clk(gclk));
	jdff dff_B_6xpklti30_1(.din(w_dff_B_rLZvEJYF1_1),.dout(w_dff_B_6xpklti30_1),.clk(gclk));
	jdff dff_B_2CwzFqti7_1(.din(w_dff_B_6xpklti30_1),.dout(w_dff_B_2CwzFqti7_1),.clk(gclk));
	jdff dff_B_OznFFY1o0_1(.din(w_dff_B_2CwzFqti7_1),.dout(w_dff_B_OznFFY1o0_1),.clk(gclk));
	jdff dff_B_EW07CUuS2_1(.din(w_dff_B_OznFFY1o0_1),.dout(w_dff_B_EW07CUuS2_1),.clk(gclk));
	jdff dff_B_6FfilXMI5_1(.din(w_dff_B_EW07CUuS2_1),.dout(w_dff_B_6FfilXMI5_1),.clk(gclk));
	jdff dff_B_94zh6EBI2_1(.din(w_dff_B_6FfilXMI5_1),.dout(w_dff_B_94zh6EBI2_1),.clk(gclk));
	jdff dff_B_mkwV1cs23_1(.din(w_dff_B_94zh6EBI2_1),.dout(w_dff_B_mkwV1cs23_1),.clk(gclk));
	jdff dff_B_TDFNha2V0_1(.din(w_dff_B_mkwV1cs23_1),.dout(w_dff_B_TDFNha2V0_1),.clk(gclk));
	jdff dff_B_kJuc7Mag6_1(.din(w_dff_B_TDFNha2V0_1),.dout(w_dff_B_kJuc7Mag6_1),.clk(gclk));
	jdff dff_B_idxkDdah9_1(.din(w_dff_B_kJuc7Mag6_1),.dout(w_dff_B_idxkDdah9_1),.clk(gclk));
	jdff dff_B_EEKgkwFg3_1(.din(w_dff_B_idxkDdah9_1),.dout(w_dff_B_EEKgkwFg3_1),.clk(gclk));
	jdff dff_B_64Zi7aej0_1(.din(w_dff_B_EEKgkwFg3_1),.dout(w_dff_B_64Zi7aej0_1),.clk(gclk));
	jdff dff_B_0JplkbLq1_1(.din(w_dff_B_64Zi7aej0_1),.dout(w_dff_B_0JplkbLq1_1),.clk(gclk));
	jdff dff_B_K6GtJeIq1_1(.din(w_dff_B_0JplkbLq1_1),.dout(w_dff_B_K6GtJeIq1_1),.clk(gclk));
	jdff dff_B_YkZSwbtn1_1(.din(w_dff_B_K6GtJeIq1_1),.dout(w_dff_B_YkZSwbtn1_1),.clk(gclk));
	jdff dff_B_cj0DCRd02_1(.din(w_dff_B_YkZSwbtn1_1),.dout(w_dff_B_cj0DCRd02_1),.clk(gclk));
	jdff dff_B_rbMxRyTo5_1(.din(w_dff_B_cj0DCRd02_1),.dout(w_dff_B_rbMxRyTo5_1),.clk(gclk));
	jdff dff_B_5tzGr4sn5_1(.din(w_dff_B_rbMxRyTo5_1),.dout(w_dff_B_5tzGr4sn5_1),.clk(gclk));
	jdff dff_B_rHvzfJJ14_1(.din(w_dff_B_5tzGr4sn5_1),.dout(w_dff_B_rHvzfJJ14_1),.clk(gclk));
	jdff dff_B_i8VpmdVF1_1(.din(w_dff_B_rHvzfJJ14_1),.dout(w_dff_B_i8VpmdVF1_1),.clk(gclk));
	jdff dff_B_MAneHMCi1_1(.din(w_dff_B_i8VpmdVF1_1),.dout(w_dff_B_MAneHMCi1_1),.clk(gclk));
	jdff dff_B_SpCXiGba5_1(.din(w_dff_B_MAneHMCi1_1),.dout(w_dff_B_SpCXiGba5_1),.clk(gclk));
	jdff dff_B_H16gR1LR8_1(.din(w_dff_B_SpCXiGba5_1),.dout(w_dff_B_H16gR1LR8_1),.clk(gclk));
	jdff dff_B_EtPlqHiY4_1(.din(w_dff_B_H16gR1LR8_1),.dout(w_dff_B_EtPlqHiY4_1),.clk(gclk));
	jdff dff_B_mCInpfKO7_1(.din(w_dff_B_EtPlqHiY4_1),.dout(w_dff_B_mCInpfKO7_1),.clk(gclk));
	jdff dff_B_3bP3hiG91_1(.din(w_dff_B_mCInpfKO7_1),.dout(w_dff_B_3bP3hiG91_1),.clk(gclk));
	jdff dff_B_X5cDXw4r7_1(.din(w_dff_B_3bP3hiG91_1),.dout(w_dff_B_X5cDXw4r7_1),.clk(gclk));
	jdff dff_B_OJL8zPrG4_1(.din(w_dff_B_X5cDXw4r7_1),.dout(w_dff_B_OJL8zPrG4_1),.clk(gclk));
	jdff dff_B_hBHzNRVd9_1(.din(w_dff_B_OJL8zPrG4_1),.dout(w_dff_B_hBHzNRVd9_1),.clk(gclk));
	jdff dff_B_dwQb54sa4_1(.din(w_dff_B_hBHzNRVd9_1),.dout(w_dff_B_dwQb54sa4_1),.clk(gclk));
	jdff dff_B_RJCOAlA64_1(.din(w_dff_B_dwQb54sa4_1),.dout(w_dff_B_RJCOAlA64_1),.clk(gclk));
	jdff dff_B_vwzyujkD1_1(.din(w_dff_B_RJCOAlA64_1),.dout(w_dff_B_vwzyujkD1_1),.clk(gclk));
	jdff dff_B_9l6upuw68_1(.din(w_dff_B_vwzyujkD1_1),.dout(w_dff_B_9l6upuw68_1),.clk(gclk));
	jdff dff_B_7ltLWsBY1_1(.din(w_dff_B_9l6upuw68_1),.dout(w_dff_B_7ltLWsBY1_1),.clk(gclk));
	jdff dff_B_iQBBJXrU8_1(.din(w_dff_B_7ltLWsBY1_1),.dout(w_dff_B_iQBBJXrU8_1),.clk(gclk));
	jdff dff_B_VXYiMtsS7_1(.din(w_dff_B_iQBBJXrU8_1),.dout(w_dff_B_VXYiMtsS7_1),.clk(gclk));
	jdff dff_B_b0te6clD6_1(.din(w_dff_B_VXYiMtsS7_1),.dout(w_dff_B_b0te6clD6_1),.clk(gclk));
	jdff dff_B_dPftqRX89_1(.din(w_dff_B_b0te6clD6_1),.dout(w_dff_B_dPftqRX89_1),.clk(gclk));
	jdff dff_B_Zmadsj9k4_1(.din(w_dff_B_dPftqRX89_1),.dout(w_dff_B_Zmadsj9k4_1),.clk(gclk));
	jdff dff_B_Ix7BLOaU6_1(.din(w_dff_B_Zmadsj9k4_1),.dout(w_dff_B_Ix7BLOaU6_1),.clk(gclk));
	jdff dff_B_VFrBBxDi6_1(.din(w_dff_B_Ix7BLOaU6_1),.dout(w_dff_B_VFrBBxDi6_1),.clk(gclk));
	jdff dff_B_CozY5rtY7_1(.din(w_dff_B_VFrBBxDi6_1),.dout(w_dff_B_CozY5rtY7_1),.clk(gclk));
	jdff dff_B_CK5ljyiq2_1(.din(w_dff_B_CozY5rtY7_1),.dout(w_dff_B_CK5ljyiq2_1),.clk(gclk));
	jdff dff_B_wckZfDj72_1(.din(w_dff_B_CK5ljyiq2_1),.dout(w_dff_B_wckZfDj72_1),.clk(gclk));
	jdff dff_B_ElPFh7Of1_1(.din(w_dff_B_wckZfDj72_1),.dout(w_dff_B_ElPFh7Of1_1),.clk(gclk));
	jdff dff_B_cixnBFfE0_1(.din(w_dff_B_ElPFh7Of1_1),.dout(w_dff_B_cixnBFfE0_1),.clk(gclk));
	jdff dff_B_sKL4thCY2_1(.din(w_dff_B_cixnBFfE0_1),.dout(w_dff_B_sKL4thCY2_1),.clk(gclk));
	jdff dff_B_1R6I2MTe0_1(.din(w_dff_B_sKL4thCY2_1),.dout(w_dff_B_1R6I2MTe0_1),.clk(gclk));
	jdff dff_B_DmiS8B3L6_0(.din(n1105),.dout(w_dff_B_DmiS8B3L6_0),.clk(gclk));
	jdff dff_B_xM345Y5V1_0(.din(w_dff_B_DmiS8B3L6_0),.dout(w_dff_B_xM345Y5V1_0),.clk(gclk));
	jdff dff_B_oSVMpu7v5_0(.din(w_dff_B_xM345Y5V1_0),.dout(w_dff_B_oSVMpu7v5_0),.clk(gclk));
	jdff dff_B_KouUV3Fd1_0(.din(w_dff_B_oSVMpu7v5_0),.dout(w_dff_B_KouUV3Fd1_0),.clk(gclk));
	jdff dff_B_Yy1fBsMj8_0(.din(w_dff_B_KouUV3Fd1_0),.dout(w_dff_B_Yy1fBsMj8_0),.clk(gclk));
	jdff dff_B_nAvb8QQy7_0(.din(w_dff_B_Yy1fBsMj8_0),.dout(w_dff_B_nAvb8QQy7_0),.clk(gclk));
	jdff dff_B_wkengbpg0_0(.din(w_dff_B_nAvb8QQy7_0),.dout(w_dff_B_wkengbpg0_0),.clk(gclk));
	jdff dff_B_dfED2d4k5_0(.din(w_dff_B_wkengbpg0_0),.dout(w_dff_B_dfED2d4k5_0),.clk(gclk));
	jdff dff_B_dJHgZWeo9_0(.din(w_dff_B_dfED2d4k5_0),.dout(w_dff_B_dJHgZWeo9_0),.clk(gclk));
	jdff dff_B_ljmptqht0_0(.din(w_dff_B_dJHgZWeo9_0),.dout(w_dff_B_ljmptqht0_0),.clk(gclk));
	jdff dff_B_Kyq8mKWQ1_0(.din(w_dff_B_ljmptqht0_0),.dout(w_dff_B_Kyq8mKWQ1_0),.clk(gclk));
	jdff dff_B_s1mHkyUz2_0(.din(w_dff_B_Kyq8mKWQ1_0),.dout(w_dff_B_s1mHkyUz2_0),.clk(gclk));
	jdff dff_B_0loYNIRv6_0(.din(w_dff_B_s1mHkyUz2_0),.dout(w_dff_B_0loYNIRv6_0),.clk(gclk));
	jdff dff_B_jdQ8jHyh8_0(.din(w_dff_B_0loYNIRv6_0),.dout(w_dff_B_jdQ8jHyh8_0),.clk(gclk));
	jdff dff_B_E1V2KQSA9_0(.din(w_dff_B_jdQ8jHyh8_0),.dout(w_dff_B_E1V2KQSA9_0),.clk(gclk));
	jdff dff_B_zMfk9k0r8_0(.din(w_dff_B_E1V2KQSA9_0),.dout(w_dff_B_zMfk9k0r8_0),.clk(gclk));
	jdff dff_B_3RRmFZWD3_0(.din(w_dff_B_zMfk9k0r8_0),.dout(w_dff_B_3RRmFZWD3_0),.clk(gclk));
	jdff dff_B_2c5LqGLI7_0(.din(w_dff_B_3RRmFZWD3_0),.dout(w_dff_B_2c5LqGLI7_0),.clk(gclk));
	jdff dff_B_lViASZIE5_0(.din(w_dff_B_2c5LqGLI7_0),.dout(w_dff_B_lViASZIE5_0),.clk(gclk));
	jdff dff_B_mPEnpJo82_0(.din(w_dff_B_lViASZIE5_0),.dout(w_dff_B_mPEnpJo82_0),.clk(gclk));
	jdff dff_B_nNwMIVFG9_0(.din(w_dff_B_mPEnpJo82_0),.dout(w_dff_B_nNwMIVFG9_0),.clk(gclk));
	jdff dff_B_7ktKAge17_0(.din(w_dff_B_nNwMIVFG9_0),.dout(w_dff_B_7ktKAge17_0),.clk(gclk));
	jdff dff_B_xsGop4tW1_0(.din(w_dff_B_7ktKAge17_0),.dout(w_dff_B_xsGop4tW1_0),.clk(gclk));
	jdff dff_B_MPpvUto57_0(.din(w_dff_B_xsGop4tW1_0),.dout(w_dff_B_MPpvUto57_0),.clk(gclk));
	jdff dff_B_W9XfOpxT6_0(.din(w_dff_B_MPpvUto57_0),.dout(w_dff_B_W9XfOpxT6_0),.clk(gclk));
	jdff dff_B_hZWpFjNb3_0(.din(w_dff_B_W9XfOpxT6_0),.dout(w_dff_B_hZWpFjNb3_0),.clk(gclk));
	jdff dff_B_x1rojjt17_0(.din(w_dff_B_hZWpFjNb3_0),.dout(w_dff_B_x1rojjt17_0),.clk(gclk));
	jdff dff_B_dNqLqrhV5_0(.din(w_dff_B_x1rojjt17_0),.dout(w_dff_B_dNqLqrhV5_0),.clk(gclk));
	jdff dff_B_T3qWaSKq3_0(.din(w_dff_B_dNqLqrhV5_0),.dout(w_dff_B_T3qWaSKq3_0),.clk(gclk));
	jdff dff_B_Xm1Erx5e7_0(.din(w_dff_B_T3qWaSKq3_0),.dout(w_dff_B_Xm1Erx5e7_0),.clk(gclk));
	jdff dff_B_wHWGp6hT9_0(.din(w_dff_B_Xm1Erx5e7_0),.dout(w_dff_B_wHWGp6hT9_0),.clk(gclk));
	jdff dff_B_bW9oJaLB3_0(.din(w_dff_B_wHWGp6hT9_0),.dout(w_dff_B_bW9oJaLB3_0),.clk(gclk));
	jdff dff_B_wu9PpQbf9_0(.din(w_dff_B_bW9oJaLB3_0),.dout(w_dff_B_wu9PpQbf9_0),.clk(gclk));
	jdff dff_B_iBx7VdQm5_0(.din(w_dff_B_wu9PpQbf9_0),.dout(w_dff_B_iBx7VdQm5_0),.clk(gclk));
	jdff dff_B_N72PAhuE2_0(.din(w_dff_B_iBx7VdQm5_0),.dout(w_dff_B_N72PAhuE2_0),.clk(gclk));
	jdff dff_B_FFOjzuJe2_0(.din(w_dff_B_N72PAhuE2_0),.dout(w_dff_B_FFOjzuJe2_0),.clk(gclk));
	jdff dff_B_slu5ZbCq0_0(.din(w_dff_B_FFOjzuJe2_0),.dout(w_dff_B_slu5ZbCq0_0),.clk(gclk));
	jdff dff_B_v9KEctaI6_0(.din(w_dff_B_slu5ZbCq0_0),.dout(w_dff_B_v9KEctaI6_0),.clk(gclk));
	jdff dff_B_KBKTvPqe1_0(.din(w_dff_B_v9KEctaI6_0),.dout(w_dff_B_KBKTvPqe1_0),.clk(gclk));
	jdff dff_B_mCLtrh4K2_0(.din(w_dff_B_KBKTvPqe1_0),.dout(w_dff_B_mCLtrh4K2_0),.clk(gclk));
	jdff dff_B_w7nRcUPN4_0(.din(w_dff_B_mCLtrh4K2_0),.dout(w_dff_B_w7nRcUPN4_0),.clk(gclk));
	jdff dff_B_m7SxjzDl7_0(.din(w_dff_B_w7nRcUPN4_0),.dout(w_dff_B_m7SxjzDl7_0),.clk(gclk));
	jdff dff_B_ZKKb9tCi2_0(.din(w_dff_B_m7SxjzDl7_0),.dout(w_dff_B_ZKKb9tCi2_0),.clk(gclk));
	jdff dff_B_kR8FmrOM0_0(.din(w_dff_B_ZKKb9tCi2_0),.dout(w_dff_B_kR8FmrOM0_0),.clk(gclk));
	jdff dff_B_tBfkhtXm6_0(.din(w_dff_B_kR8FmrOM0_0),.dout(w_dff_B_tBfkhtXm6_0),.clk(gclk));
	jdff dff_B_pLKwh8m85_0(.din(w_dff_B_tBfkhtXm6_0),.dout(w_dff_B_pLKwh8m85_0),.clk(gclk));
	jdff dff_B_guDWjVXa2_0(.din(w_dff_B_pLKwh8m85_0),.dout(w_dff_B_guDWjVXa2_0),.clk(gclk));
	jdff dff_B_tw7DMU3u7_0(.din(w_dff_B_guDWjVXa2_0),.dout(w_dff_B_tw7DMU3u7_0),.clk(gclk));
	jdff dff_B_AZ7Okffn0_0(.din(w_dff_B_tw7DMU3u7_0),.dout(w_dff_B_AZ7Okffn0_0),.clk(gclk));
	jdff dff_B_ppIKGOWx6_0(.din(w_dff_B_AZ7Okffn0_0),.dout(w_dff_B_ppIKGOWx6_0),.clk(gclk));
	jdff dff_B_uvX2sCY46_0(.din(w_dff_B_ppIKGOWx6_0),.dout(w_dff_B_uvX2sCY46_0),.clk(gclk));
	jdff dff_B_obRL9Nk68_0(.din(w_dff_B_uvX2sCY46_0),.dout(w_dff_B_obRL9Nk68_0),.clk(gclk));
	jdff dff_B_qWD0E8fM5_0(.din(w_dff_B_obRL9Nk68_0),.dout(w_dff_B_qWD0E8fM5_0),.clk(gclk));
	jdff dff_B_z0aR4dFB1_0(.din(w_dff_B_qWD0E8fM5_0),.dout(w_dff_B_z0aR4dFB1_0),.clk(gclk));
	jdff dff_B_0DOth7S28_0(.din(w_dff_B_z0aR4dFB1_0),.dout(w_dff_B_0DOth7S28_0),.clk(gclk));
	jdff dff_B_xeLSmYp20_0(.din(w_dff_B_0DOth7S28_0),.dout(w_dff_B_xeLSmYp20_0),.clk(gclk));
	jdff dff_B_c2xrgluw2_0(.din(w_dff_B_xeLSmYp20_0),.dout(w_dff_B_c2xrgluw2_0),.clk(gclk));
	jdff dff_B_d6r4A8FF6_0(.din(w_dff_B_c2xrgluw2_0),.dout(w_dff_B_d6r4A8FF6_0),.clk(gclk));
	jdff dff_B_JEvOvgSL6_0(.din(w_dff_B_d6r4A8FF6_0),.dout(w_dff_B_JEvOvgSL6_0),.clk(gclk));
	jdff dff_B_xYXnW7nk7_0(.din(w_dff_B_JEvOvgSL6_0),.dout(w_dff_B_xYXnW7nk7_0),.clk(gclk));
	jdff dff_B_SOqUhn952_0(.din(w_dff_B_xYXnW7nk7_0),.dout(w_dff_B_SOqUhn952_0),.clk(gclk));
	jdff dff_B_SAxdX41Y0_0(.din(w_dff_B_SOqUhn952_0),.dout(w_dff_B_SAxdX41Y0_0),.clk(gclk));
	jdff dff_B_Hcbg1YCr6_0(.din(w_dff_B_SAxdX41Y0_0),.dout(w_dff_B_Hcbg1YCr6_0),.clk(gclk));
	jdff dff_B_PGV85OmQ9_0(.din(w_dff_B_Hcbg1YCr6_0),.dout(w_dff_B_PGV85OmQ9_0),.clk(gclk));
	jdff dff_B_j54TmuRa9_0(.din(w_dff_B_PGV85OmQ9_0),.dout(w_dff_B_j54TmuRa9_0),.clk(gclk));
	jdff dff_B_bztkgWoP0_0(.din(w_dff_B_j54TmuRa9_0),.dout(w_dff_B_bztkgWoP0_0),.clk(gclk));
	jdff dff_B_qjPM2jJE8_0(.din(w_dff_B_bztkgWoP0_0),.dout(w_dff_B_qjPM2jJE8_0),.clk(gclk));
	jdff dff_B_okt0GNZc0_0(.din(w_dff_B_qjPM2jJE8_0),.dout(w_dff_B_okt0GNZc0_0),.clk(gclk));
	jdff dff_B_25Fh1sIl3_0(.din(w_dff_B_okt0GNZc0_0),.dout(w_dff_B_25Fh1sIl3_0),.clk(gclk));
	jdff dff_B_EKVjkUM46_0(.din(w_dff_B_25Fh1sIl3_0),.dout(w_dff_B_EKVjkUM46_0),.clk(gclk));
	jdff dff_B_q9JfqPeX9_0(.din(w_dff_B_EKVjkUM46_0),.dout(w_dff_B_q9JfqPeX9_0),.clk(gclk));
	jdff dff_B_uPnr1PXO2_0(.din(w_dff_B_q9JfqPeX9_0),.dout(w_dff_B_uPnr1PXO2_0),.clk(gclk));
	jdff dff_B_Ase3oQJF2_0(.din(w_dff_B_uPnr1PXO2_0),.dout(w_dff_B_Ase3oQJF2_0),.clk(gclk));
	jdff dff_B_ELk0EIzV2_0(.din(w_dff_B_Ase3oQJF2_0),.dout(w_dff_B_ELk0EIzV2_0),.clk(gclk));
	jdff dff_B_I3pdV6ZQ7_0(.din(w_dff_B_ELk0EIzV2_0),.dout(w_dff_B_I3pdV6ZQ7_0),.clk(gclk));
	jdff dff_B_VMtiRCuB4_0(.din(w_dff_B_I3pdV6ZQ7_0),.dout(w_dff_B_VMtiRCuB4_0),.clk(gclk));
	jdff dff_B_69LrehmD4_0(.din(w_dff_B_VMtiRCuB4_0),.dout(w_dff_B_69LrehmD4_0),.clk(gclk));
	jdff dff_B_FVWarx0c0_0(.din(w_dff_B_69LrehmD4_0),.dout(w_dff_B_FVWarx0c0_0),.clk(gclk));
	jdff dff_B_WkrqLDnN7_0(.din(w_dff_B_FVWarx0c0_0),.dout(w_dff_B_WkrqLDnN7_0),.clk(gclk));
	jdff dff_B_i0uWrgGi7_0(.din(w_dff_B_WkrqLDnN7_0),.dout(w_dff_B_i0uWrgGi7_0),.clk(gclk));
	jdff dff_B_YesU9k7I7_0(.din(w_dff_B_i0uWrgGi7_0),.dout(w_dff_B_YesU9k7I7_0),.clk(gclk));
	jdff dff_B_e4Q0tUh28_0(.din(w_dff_B_YesU9k7I7_0),.dout(w_dff_B_e4Q0tUh28_0),.clk(gclk));
	jdff dff_B_49iqi9vY3_0(.din(w_dff_B_e4Q0tUh28_0),.dout(w_dff_B_49iqi9vY3_0),.clk(gclk));
	jdff dff_B_i0V7VUL25_0(.din(w_dff_B_49iqi9vY3_0),.dout(w_dff_B_i0V7VUL25_0),.clk(gclk));
	jdff dff_B_wU6ltCAi4_0(.din(w_dff_B_i0V7VUL25_0),.dout(w_dff_B_wU6ltCAi4_0),.clk(gclk));
	jdff dff_B_mGSRjdud1_0(.din(w_dff_B_wU6ltCAi4_0),.dout(w_dff_B_mGSRjdud1_0),.clk(gclk));
	jdff dff_B_iUAbyBWy9_0(.din(w_dff_B_mGSRjdud1_0),.dout(w_dff_B_iUAbyBWy9_0),.clk(gclk));
	jdff dff_B_bZgMucZP1_0(.din(w_dff_B_iUAbyBWy9_0),.dout(w_dff_B_bZgMucZP1_0),.clk(gclk));
	jdff dff_B_nRGCw61o8_0(.din(w_dff_B_bZgMucZP1_0),.dout(w_dff_B_nRGCw61o8_0),.clk(gclk));
	jdff dff_B_81XXrLxH6_0(.din(w_dff_B_nRGCw61o8_0),.dout(w_dff_B_81XXrLxH6_0),.clk(gclk));
	jdff dff_B_WFX7lA4x4_0(.din(w_dff_B_81XXrLxH6_0),.dout(w_dff_B_WFX7lA4x4_0),.clk(gclk));
	jdff dff_B_ADdjmPg34_0(.din(w_dff_B_WFX7lA4x4_0),.dout(w_dff_B_ADdjmPg34_0),.clk(gclk));
	jdff dff_B_xiMQvOmp7_0(.din(w_dff_B_ADdjmPg34_0),.dout(w_dff_B_xiMQvOmp7_0),.clk(gclk));
	jdff dff_B_XHdonrsG8_0(.din(w_dff_B_xiMQvOmp7_0),.dout(w_dff_B_XHdonrsG8_0),.clk(gclk));
	jdff dff_B_oQaVnIZW9_0(.din(w_dff_B_XHdonrsG8_0),.dout(w_dff_B_oQaVnIZW9_0),.clk(gclk));
	jdff dff_B_wu6hGo3Y6_0(.din(w_dff_B_oQaVnIZW9_0),.dout(w_dff_B_wu6hGo3Y6_0),.clk(gclk));
	jdff dff_B_wC10m9iq3_0(.din(w_dff_B_wu6hGo3Y6_0),.dout(w_dff_B_wC10m9iq3_0),.clk(gclk));
	jdff dff_B_5A8lEkG11_0(.din(w_dff_B_wC10m9iq3_0),.dout(w_dff_B_5A8lEkG11_0),.clk(gclk));
	jdff dff_B_ZQ3O21mD6_0(.din(w_dff_B_5A8lEkG11_0),.dout(w_dff_B_ZQ3O21mD6_0),.clk(gclk));
	jdff dff_B_oFzw8wIp7_0(.din(w_dff_B_ZQ3O21mD6_0),.dout(w_dff_B_oFzw8wIp7_0),.clk(gclk));
	jdff dff_B_oVB96x231_0(.din(w_dff_B_oFzw8wIp7_0),.dout(w_dff_B_oVB96x231_0),.clk(gclk));
	jdff dff_B_s6kolGIt8_0(.din(w_dff_B_oVB96x231_0),.dout(w_dff_B_s6kolGIt8_0),.clk(gclk));
	jdff dff_B_QmsGdkTE8_0(.din(w_dff_B_s6kolGIt8_0),.dout(w_dff_B_QmsGdkTE8_0),.clk(gclk));
	jdff dff_B_IkOAgSwj0_0(.din(w_dff_B_QmsGdkTE8_0),.dout(w_dff_B_IkOAgSwj0_0),.clk(gclk));
	jdff dff_B_hRaer5xI2_0(.din(w_dff_B_IkOAgSwj0_0),.dout(w_dff_B_hRaer5xI2_0),.clk(gclk));
	jdff dff_B_rwRBUbz36_0(.din(w_dff_B_hRaer5xI2_0),.dout(w_dff_B_rwRBUbz36_0),.clk(gclk));
	jdff dff_B_9ykGo8Rk9_0(.din(w_dff_B_rwRBUbz36_0),.dout(w_dff_B_9ykGo8Rk9_0),.clk(gclk));
	jdff dff_B_901ryyiL2_0(.din(w_dff_B_9ykGo8Rk9_0),.dout(w_dff_B_901ryyiL2_0),.clk(gclk));
	jdff dff_B_kvAOLe5b5_0(.din(w_dff_B_901ryyiL2_0),.dout(w_dff_B_kvAOLe5b5_0),.clk(gclk));
	jdff dff_B_0gEsQm253_0(.din(w_dff_B_kvAOLe5b5_0),.dout(w_dff_B_0gEsQm253_0),.clk(gclk));
	jdff dff_B_gCBSyele0_0(.din(w_dff_B_0gEsQm253_0),.dout(w_dff_B_gCBSyele0_0),.clk(gclk));
	jdff dff_B_fToHlPGI9_0(.din(w_dff_B_gCBSyele0_0),.dout(w_dff_B_fToHlPGI9_0),.clk(gclk));
	jdff dff_B_8veaDZvP9_0(.din(w_dff_B_fToHlPGI9_0),.dout(w_dff_B_8veaDZvP9_0),.clk(gclk));
	jdff dff_B_rYFOO46L8_0(.din(w_dff_B_8veaDZvP9_0),.dout(w_dff_B_rYFOO46L8_0),.clk(gclk));
	jdff dff_B_RXU664dX3_0(.din(w_dff_B_rYFOO46L8_0),.dout(w_dff_B_RXU664dX3_0),.clk(gclk));
	jdff dff_B_GeyrJEWw2_0(.din(w_dff_B_RXU664dX3_0),.dout(w_dff_B_GeyrJEWw2_0),.clk(gclk));
	jdff dff_B_Xua6oPfC8_0(.din(w_dff_B_GeyrJEWw2_0),.dout(w_dff_B_Xua6oPfC8_0),.clk(gclk));
	jdff dff_B_f4y5YBEj1_0(.din(w_dff_B_Xua6oPfC8_0),.dout(w_dff_B_f4y5YBEj1_0),.clk(gclk));
	jdff dff_B_VUdKXJJA4_0(.din(w_dff_B_f4y5YBEj1_0),.dout(w_dff_B_VUdKXJJA4_0),.clk(gclk));
	jdff dff_B_urlYAJ559_0(.din(w_dff_B_VUdKXJJA4_0),.dout(w_dff_B_urlYAJ559_0),.clk(gclk));
	jdff dff_B_6ZJ2B90F4_1(.din(n1098),.dout(w_dff_B_6ZJ2B90F4_1),.clk(gclk));
	jdff dff_B_XgC1VJGa5_1(.din(w_dff_B_6ZJ2B90F4_1),.dout(w_dff_B_XgC1VJGa5_1),.clk(gclk));
	jdff dff_B_WmFTPlty5_1(.din(w_dff_B_XgC1VJGa5_1),.dout(w_dff_B_WmFTPlty5_1),.clk(gclk));
	jdff dff_B_8EtGIwQl3_1(.din(w_dff_B_WmFTPlty5_1),.dout(w_dff_B_8EtGIwQl3_1),.clk(gclk));
	jdff dff_B_wkSUwda18_1(.din(w_dff_B_8EtGIwQl3_1),.dout(w_dff_B_wkSUwda18_1),.clk(gclk));
	jdff dff_B_VwBccq4w1_1(.din(w_dff_B_wkSUwda18_1),.dout(w_dff_B_VwBccq4w1_1),.clk(gclk));
	jdff dff_B_M7KbPZg11_1(.din(w_dff_B_VwBccq4w1_1),.dout(w_dff_B_M7KbPZg11_1),.clk(gclk));
	jdff dff_B_C1gAATUa6_1(.din(w_dff_B_M7KbPZg11_1),.dout(w_dff_B_C1gAATUa6_1),.clk(gclk));
	jdff dff_B_qeGtAeP11_1(.din(w_dff_B_C1gAATUa6_1),.dout(w_dff_B_qeGtAeP11_1),.clk(gclk));
	jdff dff_B_20oawz8w8_1(.din(w_dff_B_qeGtAeP11_1),.dout(w_dff_B_20oawz8w8_1),.clk(gclk));
	jdff dff_B_4brz1GLZ3_1(.din(w_dff_B_20oawz8w8_1),.dout(w_dff_B_4brz1GLZ3_1),.clk(gclk));
	jdff dff_B_zrub0edS1_1(.din(w_dff_B_4brz1GLZ3_1),.dout(w_dff_B_zrub0edS1_1),.clk(gclk));
	jdff dff_B_sM48ITAY0_1(.din(w_dff_B_zrub0edS1_1),.dout(w_dff_B_sM48ITAY0_1),.clk(gclk));
	jdff dff_B_Xu8dHqAK3_1(.din(w_dff_B_sM48ITAY0_1),.dout(w_dff_B_Xu8dHqAK3_1),.clk(gclk));
	jdff dff_B_fL4r92p34_1(.din(w_dff_B_Xu8dHqAK3_1),.dout(w_dff_B_fL4r92p34_1),.clk(gclk));
	jdff dff_B_WfLpBtFN7_1(.din(w_dff_B_fL4r92p34_1),.dout(w_dff_B_WfLpBtFN7_1),.clk(gclk));
	jdff dff_B_iz6GKrWj5_1(.din(w_dff_B_WfLpBtFN7_1),.dout(w_dff_B_iz6GKrWj5_1),.clk(gclk));
	jdff dff_B_wyixcF4B0_1(.din(w_dff_B_iz6GKrWj5_1),.dout(w_dff_B_wyixcF4B0_1),.clk(gclk));
	jdff dff_B_AO8gYpzD9_1(.din(w_dff_B_wyixcF4B0_1),.dout(w_dff_B_AO8gYpzD9_1),.clk(gclk));
	jdff dff_B_uOiJMq6z7_1(.din(w_dff_B_AO8gYpzD9_1),.dout(w_dff_B_uOiJMq6z7_1),.clk(gclk));
	jdff dff_B_WO3mDd509_1(.din(w_dff_B_uOiJMq6z7_1),.dout(w_dff_B_WO3mDd509_1),.clk(gclk));
	jdff dff_B_EDFrqSX08_1(.din(w_dff_B_WO3mDd509_1),.dout(w_dff_B_EDFrqSX08_1),.clk(gclk));
	jdff dff_B_4SwMoBnw2_1(.din(w_dff_B_EDFrqSX08_1),.dout(w_dff_B_4SwMoBnw2_1),.clk(gclk));
	jdff dff_B_YdzkRIGQ2_1(.din(w_dff_B_4SwMoBnw2_1),.dout(w_dff_B_YdzkRIGQ2_1),.clk(gclk));
	jdff dff_B_e1ZjCM265_1(.din(w_dff_B_YdzkRIGQ2_1),.dout(w_dff_B_e1ZjCM265_1),.clk(gclk));
	jdff dff_B_LPgF5hbc9_1(.din(w_dff_B_e1ZjCM265_1),.dout(w_dff_B_LPgF5hbc9_1),.clk(gclk));
	jdff dff_B_6dyapKtA8_1(.din(w_dff_B_LPgF5hbc9_1),.dout(w_dff_B_6dyapKtA8_1),.clk(gclk));
	jdff dff_B_0QxXBDYG7_1(.din(w_dff_B_6dyapKtA8_1),.dout(w_dff_B_0QxXBDYG7_1),.clk(gclk));
	jdff dff_B_98SYshbP6_1(.din(w_dff_B_0QxXBDYG7_1),.dout(w_dff_B_98SYshbP6_1),.clk(gclk));
	jdff dff_B_urFNhsEF8_1(.din(w_dff_B_98SYshbP6_1),.dout(w_dff_B_urFNhsEF8_1),.clk(gclk));
	jdff dff_B_PIt4L3yH5_1(.din(w_dff_B_urFNhsEF8_1),.dout(w_dff_B_PIt4L3yH5_1),.clk(gclk));
	jdff dff_B_EPL9IKN54_1(.din(w_dff_B_PIt4L3yH5_1),.dout(w_dff_B_EPL9IKN54_1),.clk(gclk));
	jdff dff_B_Of9cqFmO5_1(.din(w_dff_B_EPL9IKN54_1),.dout(w_dff_B_Of9cqFmO5_1),.clk(gclk));
	jdff dff_B_GISs8RJ51_1(.din(w_dff_B_Of9cqFmO5_1),.dout(w_dff_B_GISs8RJ51_1),.clk(gclk));
	jdff dff_B_dYhzJzpb8_1(.din(w_dff_B_GISs8RJ51_1),.dout(w_dff_B_dYhzJzpb8_1),.clk(gclk));
	jdff dff_B_8Ly5VTXd8_1(.din(w_dff_B_dYhzJzpb8_1),.dout(w_dff_B_8Ly5VTXd8_1),.clk(gclk));
	jdff dff_B_DbFJDAab5_1(.din(w_dff_B_8Ly5VTXd8_1),.dout(w_dff_B_DbFJDAab5_1),.clk(gclk));
	jdff dff_B_ZG6E00pS5_1(.din(w_dff_B_DbFJDAab5_1),.dout(w_dff_B_ZG6E00pS5_1),.clk(gclk));
	jdff dff_B_V9E5ZCbc0_1(.din(w_dff_B_ZG6E00pS5_1),.dout(w_dff_B_V9E5ZCbc0_1),.clk(gclk));
	jdff dff_B_zPKZP7zU2_1(.din(w_dff_B_V9E5ZCbc0_1),.dout(w_dff_B_zPKZP7zU2_1),.clk(gclk));
	jdff dff_B_BrVhiL6R4_1(.din(w_dff_B_zPKZP7zU2_1),.dout(w_dff_B_BrVhiL6R4_1),.clk(gclk));
	jdff dff_B_VutLSd6n2_1(.din(w_dff_B_BrVhiL6R4_1),.dout(w_dff_B_VutLSd6n2_1),.clk(gclk));
	jdff dff_B_JFCPEFzO0_1(.din(w_dff_B_VutLSd6n2_1),.dout(w_dff_B_JFCPEFzO0_1),.clk(gclk));
	jdff dff_B_30izPVSv6_1(.din(w_dff_B_JFCPEFzO0_1),.dout(w_dff_B_30izPVSv6_1),.clk(gclk));
	jdff dff_B_Wk0fSFGf1_1(.din(w_dff_B_30izPVSv6_1),.dout(w_dff_B_Wk0fSFGf1_1),.clk(gclk));
	jdff dff_B_SXk16agu8_1(.din(w_dff_B_Wk0fSFGf1_1),.dout(w_dff_B_SXk16agu8_1),.clk(gclk));
	jdff dff_B_PvVYcDLX3_1(.din(w_dff_B_SXk16agu8_1),.dout(w_dff_B_PvVYcDLX3_1),.clk(gclk));
	jdff dff_B_qoCEinwP9_1(.din(w_dff_B_PvVYcDLX3_1),.dout(w_dff_B_qoCEinwP9_1),.clk(gclk));
	jdff dff_B_o1h7roaU7_1(.din(w_dff_B_qoCEinwP9_1),.dout(w_dff_B_o1h7roaU7_1),.clk(gclk));
	jdff dff_B_JB3fTzTe2_1(.din(w_dff_B_o1h7roaU7_1),.dout(w_dff_B_JB3fTzTe2_1),.clk(gclk));
	jdff dff_B_jm7fkLfB0_1(.din(w_dff_B_JB3fTzTe2_1),.dout(w_dff_B_jm7fkLfB0_1),.clk(gclk));
	jdff dff_B_XNEXT1Yz7_1(.din(w_dff_B_jm7fkLfB0_1),.dout(w_dff_B_XNEXT1Yz7_1),.clk(gclk));
	jdff dff_B_YRJHmesp2_1(.din(w_dff_B_XNEXT1Yz7_1),.dout(w_dff_B_YRJHmesp2_1),.clk(gclk));
	jdff dff_B_SqtNvor55_1(.din(w_dff_B_YRJHmesp2_1),.dout(w_dff_B_SqtNvor55_1),.clk(gclk));
	jdff dff_B_iPznLBaZ5_1(.din(w_dff_B_SqtNvor55_1),.dout(w_dff_B_iPznLBaZ5_1),.clk(gclk));
	jdff dff_B_mMYuIlKN1_1(.din(w_dff_B_iPznLBaZ5_1),.dout(w_dff_B_mMYuIlKN1_1),.clk(gclk));
	jdff dff_B_2NAZTEHk9_1(.din(w_dff_B_mMYuIlKN1_1),.dout(w_dff_B_2NAZTEHk9_1),.clk(gclk));
	jdff dff_B_9Ww78L353_1(.din(w_dff_B_2NAZTEHk9_1),.dout(w_dff_B_9Ww78L353_1),.clk(gclk));
	jdff dff_B_kRLCanVC8_1(.din(w_dff_B_9Ww78L353_1),.dout(w_dff_B_kRLCanVC8_1),.clk(gclk));
	jdff dff_B_HZqQIV0C5_1(.din(w_dff_B_kRLCanVC8_1),.dout(w_dff_B_HZqQIV0C5_1),.clk(gclk));
	jdff dff_B_M1Si2zLj9_1(.din(w_dff_B_HZqQIV0C5_1),.dout(w_dff_B_M1Si2zLj9_1),.clk(gclk));
	jdff dff_B_2Y7KoNG93_1(.din(w_dff_B_M1Si2zLj9_1),.dout(w_dff_B_2Y7KoNG93_1),.clk(gclk));
	jdff dff_B_3cnDEG7O2_1(.din(w_dff_B_2Y7KoNG93_1),.dout(w_dff_B_3cnDEG7O2_1),.clk(gclk));
	jdff dff_B_NQ50Ym6f1_1(.din(w_dff_B_3cnDEG7O2_1),.dout(w_dff_B_NQ50Ym6f1_1),.clk(gclk));
	jdff dff_B_PYA67cGF4_1(.din(w_dff_B_NQ50Ym6f1_1),.dout(w_dff_B_PYA67cGF4_1),.clk(gclk));
	jdff dff_B_nayPBG5B4_1(.din(w_dff_B_PYA67cGF4_1),.dout(w_dff_B_nayPBG5B4_1),.clk(gclk));
	jdff dff_B_4ulNaD3g2_1(.din(w_dff_B_nayPBG5B4_1),.dout(w_dff_B_4ulNaD3g2_1),.clk(gclk));
	jdff dff_B_kDmaarHJ3_1(.din(w_dff_B_4ulNaD3g2_1),.dout(w_dff_B_kDmaarHJ3_1),.clk(gclk));
	jdff dff_B_Bnr84nrE0_1(.din(w_dff_B_kDmaarHJ3_1),.dout(w_dff_B_Bnr84nrE0_1),.clk(gclk));
	jdff dff_B_pq6LVOGV7_1(.din(w_dff_B_Bnr84nrE0_1),.dout(w_dff_B_pq6LVOGV7_1),.clk(gclk));
	jdff dff_B_drpfdpA27_1(.din(w_dff_B_pq6LVOGV7_1),.dout(w_dff_B_drpfdpA27_1),.clk(gclk));
	jdff dff_B_PJuHsV6V7_1(.din(w_dff_B_drpfdpA27_1),.dout(w_dff_B_PJuHsV6V7_1),.clk(gclk));
	jdff dff_B_fa5dLJkX3_1(.din(w_dff_B_PJuHsV6V7_1),.dout(w_dff_B_fa5dLJkX3_1),.clk(gclk));
	jdff dff_B_RTmzCHU50_1(.din(w_dff_B_fa5dLJkX3_1),.dout(w_dff_B_RTmzCHU50_1),.clk(gclk));
	jdff dff_B_OLvzY3yV7_1(.din(w_dff_B_RTmzCHU50_1),.dout(w_dff_B_OLvzY3yV7_1),.clk(gclk));
	jdff dff_B_n24jqsHS5_1(.din(w_dff_B_OLvzY3yV7_1),.dout(w_dff_B_n24jqsHS5_1),.clk(gclk));
	jdff dff_B_PdbcKl9C7_1(.din(w_dff_B_n24jqsHS5_1),.dout(w_dff_B_PdbcKl9C7_1),.clk(gclk));
	jdff dff_B_hsnAgIWa7_1(.din(w_dff_B_PdbcKl9C7_1),.dout(w_dff_B_hsnAgIWa7_1),.clk(gclk));
	jdff dff_B_ym7hkXN32_1(.din(w_dff_B_hsnAgIWa7_1),.dout(w_dff_B_ym7hkXN32_1),.clk(gclk));
	jdff dff_B_7L1oB9EE3_1(.din(w_dff_B_ym7hkXN32_1),.dout(w_dff_B_7L1oB9EE3_1),.clk(gclk));
	jdff dff_B_ApfBJJJa7_1(.din(w_dff_B_7L1oB9EE3_1),.dout(w_dff_B_ApfBJJJa7_1),.clk(gclk));
	jdff dff_B_q6X1lfWl7_1(.din(w_dff_B_ApfBJJJa7_1),.dout(w_dff_B_q6X1lfWl7_1),.clk(gclk));
	jdff dff_B_YTRcjFPY5_1(.din(w_dff_B_q6X1lfWl7_1),.dout(w_dff_B_YTRcjFPY5_1),.clk(gclk));
	jdff dff_B_Gcy5hbj28_1(.din(w_dff_B_YTRcjFPY5_1),.dout(w_dff_B_Gcy5hbj28_1),.clk(gclk));
	jdff dff_B_CZQncF1E6_1(.din(w_dff_B_Gcy5hbj28_1),.dout(w_dff_B_CZQncF1E6_1),.clk(gclk));
	jdff dff_B_JBLnxQhL5_1(.din(w_dff_B_CZQncF1E6_1),.dout(w_dff_B_JBLnxQhL5_1),.clk(gclk));
	jdff dff_B_VoUNmmqo6_1(.din(w_dff_B_JBLnxQhL5_1),.dout(w_dff_B_VoUNmmqo6_1),.clk(gclk));
	jdff dff_B_63FwWgcJ4_1(.din(w_dff_B_VoUNmmqo6_1),.dout(w_dff_B_63FwWgcJ4_1),.clk(gclk));
	jdff dff_B_pXt3VUrN4_1(.din(w_dff_B_63FwWgcJ4_1),.dout(w_dff_B_pXt3VUrN4_1),.clk(gclk));
	jdff dff_B_ybk2Lthi7_1(.din(w_dff_B_pXt3VUrN4_1),.dout(w_dff_B_ybk2Lthi7_1),.clk(gclk));
	jdff dff_B_sEFt6puM4_1(.din(w_dff_B_ybk2Lthi7_1),.dout(w_dff_B_sEFt6puM4_1),.clk(gclk));
	jdff dff_B_InfOptXn7_1(.din(w_dff_B_sEFt6puM4_1),.dout(w_dff_B_InfOptXn7_1),.clk(gclk));
	jdff dff_B_GJsT1EFX3_1(.din(w_dff_B_InfOptXn7_1),.dout(w_dff_B_GJsT1EFX3_1),.clk(gclk));
	jdff dff_B_KFZzT8EC1_1(.din(w_dff_B_GJsT1EFX3_1),.dout(w_dff_B_KFZzT8EC1_1),.clk(gclk));
	jdff dff_B_zeegFoI83_1(.din(w_dff_B_KFZzT8EC1_1),.dout(w_dff_B_zeegFoI83_1),.clk(gclk));
	jdff dff_B_oNZa8tcN5_1(.din(w_dff_B_zeegFoI83_1),.dout(w_dff_B_oNZa8tcN5_1),.clk(gclk));
	jdff dff_B_wEZ7oaDq3_1(.din(w_dff_B_oNZa8tcN5_1),.dout(w_dff_B_wEZ7oaDq3_1),.clk(gclk));
	jdff dff_B_kdT267tF2_1(.din(w_dff_B_wEZ7oaDq3_1),.dout(w_dff_B_kdT267tF2_1),.clk(gclk));
	jdff dff_B_ByNyOFpy6_1(.din(w_dff_B_kdT267tF2_1),.dout(w_dff_B_ByNyOFpy6_1),.clk(gclk));
	jdff dff_B_9P3BuhQo2_1(.din(w_dff_B_ByNyOFpy6_1),.dout(w_dff_B_9P3BuhQo2_1),.clk(gclk));
	jdff dff_B_vN3PQZCt4_1(.din(w_dff_B_9P3BuhQo2_1),.dout(w_dff_B_vN3PQZCt4_1),.clk(gclk));
	jdff dff_B_Gai0xEha7_1(.din(w_dff_B_vN3PQZCt4_1),.dout(w_dff_B_Gai0xEha7_1),.clk(gclk));
	jdff dff_B_7UDU43za0_1(.din(w_dff_B_Gai0xEha7_1),.dout(w_dff_B_7UDU43za0_1),.clk(gclk));
	jdff dff_B_2VUUf3kt9_1(.din(w_dff_B_7UDU43za0_1),.dout(w_dff_B_2VUUf3kt9_1),.clk(gclk));
	jdff dff_B_rZOacF6j8_1(.din(w_dff_B_2VUUf3kt9_1),.dout(w_dff_B_rZOacF6j8_1),.clk(gclk));
	jdff dff_B_FPE0Tijx2_1(.din(w_dff_B_rZOacF6j8_1),.dout(w_dff_B_FPE0Tijx2_1),.clk(gclk));
	jdff dff_B_ThiYQWt53_1(.din(w_dff_B_FPE0Tijx2_1),.dout(w_dff_B_ThiYQWt53_1),.clk(gclk));
	jdff dff_B_VJrSGc3j8_1(.din(w_dff_B_ThiYQWt53_1),.dout(w_dff_B_VJrSGc3j8_1),.clk(gclk));
	jdff dff_B_mddY9Gl86_1(.din(w_dff_B_VJrSGc3j8_1),.dout(w_dff_B_mddY9Gl86_1),.clk(gclk));
	jdff dff_B_j3h3KUec4_1(.din(w_dff_B_mddY9Gl86_1),.dout(w_dff_B_j3h3KUec4_1),.clk(gclk));
	jdff dff_B_NSTQJrwo2_1(.din(w_dff_B_j3h3KUec4_1),.dout(w_dff_B_NSTQJrwo2_1),.clk(gclk));
	jdff dff_B_o2gN1zCD0_1(.din(w_dff_B_NSTQJrwo2_1),.dout(w_dff_B_o2gN1zCD0_1),.clk(gclk));
	jdff dff_B_XTp20tg52_1(.din(w_dff_B_o2gN1zCD0_1),.dout(w_dff_B_XTp20tg52_1),.clk(gclk));
	jdff dff_B_Pv7emCxc2_1(.din(w_dff_B_XTp20tg52_1),.dout(w_dff_B_Pv7emCxc2_1),.clk(gclk));
	jdff dff_B_phve4e6S7_1(.din(w_dff_B_Pv7emCxc2_1),.dout(w_dff_B_phve4e6S7_1),.clk(gclk));
	jdff dff_B_2HboaWI04_1(.din(w_dff_B_phve4e6S7_1),.dout(w_dff_B_2HboaWI04_1),.clk(gclk));
	jdff dff_B_Gbt3fbkn3_1(.din(w_dff_B_2HboaWI04_1),.dout(w_dff_B_Gbt3fbkn3_1),.clk(gclk));
	jdff dff_B_ClWslrlp8_1(.din(w_dff_B_Gbt3fbkn3_1),.dout(w_dff_B_ClWslrlp8_1),.clk(gclk));
	jdff dff_B_UxHmoAjS1_1(.din(w_dff_B_ClWslrlp8_1),.dout(w_dff_B_UxHmoAjS1_1),.clk(gclk));
	jdff dff_B_OBvIyR2T2_0(.din(n1099),.dout(w_dff_B_OBvIyR2T2_0),.clk(gclk));
	jdff dff_B_eWmltQAJ2_0(.din(w_dff_B_OBvIyR2T2_0),.dout(w_dff_B_eWmltQAJ2_0),.clk(gclk));
	jdff dff_B_Y72cGf7J8_0(.din(w_dff_B_eWmltQAJ2_0),.dout(w_dff_B_Y72cGf7J8_0),.clk(gclk));
	jdff dff_B_BC3x89br9_0(.din(w_dff_B_Y72cGf7J8_0),.dout(w_dff_B_BC3x89br9_0),.clk(gclk));
	jdff dff_B_MEM72NPB9_0(.din(w_dff_B_BC3x89br9_0),.dout(w_dff_B_MEM72NPB9_0),.clk(gclk));
	jdff dff_B_Rxh12fnE0_0(.din(w_dff_B_MEM72NPB9_0),.dout(w_dff_B_Rxh12fnE0_0),.clk(gclk));
	jdff dff_B_UoFrLTCG1_0(.din(w_dff_B_Rxh12fnE0_0),.dout(w_dff_B_UoFrLTCG1_0),.clk(gclk));
	jdff dff_B_3OINwGFg5_0(.din(w_dff_B_UoFrLTCG1_0),.dout(w_dff_B_3OINwGFg5_0),.clk(gclk));
	jdff dff_B_mUYbJReH6_0(.din(w_dff_B_3OINwGFg5_0),.dout(w_dff_B_mUYbJReH6_0),.clk(gclk));
	jdff dff_B_TNRdxHUH4_0(.din(w_dff_B_mUYbJReH6_0),.dout(w_dff_B_TNRdxHUH4_0),.clk(gclk));
	jdff dff_B_4YzXJCMG6_0(.din(w_dff_B_TNRdxHUH4_0),.dout(w_dff_B_4YzXJCMG6_0),.clk(gclk));
	jdff dff_B_1EZGvYVA3_0(.din(w_dff_B_4YzXJCMG6_0),.dout(w_dff_B_1EZGvYVA3_0),.clk(gclk));
	jdff dff_B_rVw9kkY29_0(.din(w_dff_B_1EZGvYVA3_0),.dout(w_dff_B_rVw9kkY29_0),.clk(gclk));
	jdff dff_B_5xkRPJOT0_0(.din(w_dff_B_rVw9kkY29_0),.dout(w_dff_B_5xkRPJOT0_0),.clk(gclk));
	jdff dff_B_euOwuYcp1_0(.din(w_dff_B_5xkRPJOT0_0),.dout(w_dff_B_euOwuYcp1_0),.clk(gclk));
	jdff dff_B_3s9L8Xct4_0(.din(w_dff_B_euOwuYcp1_0),.dout(w_dff_B_3s9L8Xct4_0),.clk(gclk));
	jdff dff_B_k7W7nsZ06_0(.din(w_dff_B_3s9L8Xct4_0),.dout(w_dff_B_k7W7nsZ06_0),.clk(gclk));
	jdff dff_B_7NcmlQOG5_0(.din(w_dff_B_k7W7nsZ06_0),.dout(w_dff_B_7NcmlQOG5_0),.clk(gclk));
	jdff dff_B_xTQDePxT7_0(.din(w_dff_B_7NcmlQOG5_0),.dout(w_dff_B_xTQDePxT7_0),.clk(gclk));
	jdff dff_B_e5nEBnQ64_0(.din(w_dff_B_xTQDePxT7_0),.dout(w_dff_B_e5nEBnQ64_0),.clk(gclk));
	jdff dff_B_Cf6qzudz3_0(.din(w_dff_B_e5nEBnQ64_0),.dout(w_dff_B_Cf6qzudz3_0),.clk(gclk));
	jdff dff_B_QXgl2pq38_0(.din(w_dff_B_Cf6qzudz3_0),.dout(w_dff_B_QXgl2pq38_0),.clk(gclk));
	jdff dff_B_i3mZi5lB3_0(.din(w_dff_B_QXgl2pq38_0),.dout(w_dff_B_i3mZi5lB3_0),.clk(gclk));
	jdff dff_B_8JW7Ni1S3_0(.din(w_dff_B_i3mZi5lB3_0),.dout(w_dff_B_8JW7Ni1S3_0),.clk(gclk));
	jdff dff_B_LKO01fNs5_0(.din(w_dff_B_8JW7Ni1S3_0),.dout(w_dff_B_LKO01fNs5_0),.clk(gclk));
	jdff dff_B_eMsTXzsS2_0(.din(w_dff_B_LKO01fNs5_0),.dout(w_dff_B_eMsTXzsS2_0),.clk(gclk));
	jdff dff_B_YuiZujfi8_0(.din(w_dff_B_eMsTXzsS2_0),.dout(w_dff_B_YuiZujfi8_0),.clk(gclk));
	jdff dff_B_6eZnYLSU0_0(.din(w_dff_B_YuiZujfi8_0),.dout(w_dff_B_6eZnYLSU0_0),.clk(gclk));
	jdff dff_B_dUlwXxJt7_0(.din(w_dff_B_6eZnYLSU0_0),.dout(w_dff_B_dUlwXxJt7_0),.clk(gclk));
	jdff dff_B_ymEwlZYF7_0(.din(w_dff_B_dUlwXxJt7_0),.dout(w_dff_B_ymEwlZYF7_0),.clk(gclk));
	jdff dff_B_3G7ikQ5o6_0(.din(w_dff_B_ymEwlZYF7_0),.dout(w_dff_B_3G7ikQ5o6_0),.clk(gclk));
	jdff dff_B_pQvlhuLM9_0(.din(w_dff_B_3G7ikQ5o6_0),.dout(w_dff_B_pQvlhuLM9_0),.clk(gclk));
	jdff dff_B_ufgw2k0D4_0(.din(w_dff_B_pQvlhuLM9_0),.dout(w_dff_B_ufgw2k0D4_0),.clk(gclk));
	jdff dff_B_SGEmeXaY1_0(.din(w_dff_B_ufgw2k0D4_0),.dout(w_dff_B_SGEmeXaY1_0),.clk(gclk));
	jdff dff_B_dClj0k4s2_0(.din(w_dff_B_SGEmeXaY1_0),.dout(w_dff_B_dClj0k4s2_0),.clk(gclk));
	jdff dff_B_Jq6PPaxS6_0(.din(w_dff_B_dClj0k4s2_0),.dout(w_dff_B_Jq6PPaxS6_0),.clk(gclk));
	jdff dff_B_lRd8Bw9X9_0(.din(w_dff_B_Jq6PPaxS6_0),.dout(w_dff_B_lRd8Bw9X9_0),.clk(gclk));
	jdff dff_B_ZMqTcW402_0(.din(w_dff_B_lRd8Bw9X9_0),.dout(w_dff_B_ZMqTcW402_0),.clk(gclk));
	jdff dff_B_IZ6xCIZG4_0(.din(w_dff_B_ZMqTcW402_0),.dout(w_dff_B_IZ6xCIZG4_0),.clk(gclk));
	jdff dff_B_0GZFFMdT6_0(.din(w_dff_B_IZ6xCIZG4_0),.dout(w_dff_B_0GZFFMdT6_0),.clk(gclk));
	jdff dff_B_6EBpYBOK9_0(.din(w_dff_B_0GZFFMdT6_0),.dout(w_dff_B_6EBpYBOK9_0),.clk(gclk));
	jdff dff_B_dUEPX3IQ8_0(.din(w_dff_B_6EBpYBOK9_0),.dout(w_dff_B_dUEPX3IQ8_0),.clk(gclk));
	jdff dff_B_4EUFmaEt2_0(.din(w_dff_B_dUEPX3IQ8_0),.dout(w_dff_B_4EUFmaEt2_0),.clk(gclk));
	jdff dff_B_EXZkEsnB0_0(.din(w_dff_B_4EUFmaEt2_0),.dout(w_dff_B_EXZkEsnB0_0),.clk(gclk));
	jdff dff_B_nNv8vYer8_0(.din(w_dff_B_EXZkEsnB0_0),.dout(w_dff_B_nNv8vYer8_0),.clk(gclk));
	jdff dff_B_OtnZcrah8_0(.din(w_dff_B_nNv8vYer8_0),.dout(w_dff_B_OtnZcrah8_0),.clk(gclk));
	jdff dff_B_rLGjJ4bu1_0(.din(w_dff_B_OtnZcrah8_0),.dout(w_dff_B_rLGjJ4bu1_0),.clk(gclk));
	jdff dff_B_b07krKOj1_0(.din(w_dff_B_rLGjJ4bu1_0),.dout(w_dff_B_b07krKOj1_0),.clk(gclk));
	jdff dff_B_0kuo0w8A7_0(.din(w_dff_B_b07krKOj1_0),.dout(w_dff_B_0kuo0w8A7_0),.clk(gclk));
	jdff dff_B_bzSXEorl7_0(.din(w_dff_B_0kuo0w8A7_0),.dout(w_dff_B_bzSXEorl7_0),.clk(gclk));
	jdff dff_B_ujWic2xz4_0(.din(w_dff_B_bzSXEorl7_0),.dout(w_dff_B_ujWic2xz4_0),.clk(gclk));
	jdff dff_B_JqlrhBWN9_0(.din(w_dff_B_ujWic2xz4_0),.dout(w_dff_B_JqlrhBWN9_0),.clk(gclk));
	jdff dff_B_edZwPy4H8_0(.din(w_dff_B_JqlrhBWN9_0),.dout(w_dff_B_edZwPy4H8_0),.clk(gclk));
	jdff dff_B_fXIJTsZQ2_0(.din(w_dff_B_edZwPy4H8_0),.dout(w_dff_B_fXIJTsZQ2_0),.clk(gclk));
	jdff dff_B_atBFjTsy7_0(.din(w_dff_B_fXIJTsZQ2_0),.dout(w_dff_B_atBFjTsy7_0),.clk(gclk));
	jdff dff_B_sVCfwL192_0(.din(w_dff_B_atBFjTsy7_0),.dout(w_dff_B_sVCfwL192_0),.clk(gclk));
	jdff dff_B_KZGo2XtR5_0(.din(w_dff_B_sVCfwL192_0),.dout(w_dff_B_KZGo2XtR5_0),.clk(gclk));
	jdff dff_B_uDWde4n81_0(.din(w_dff_B_KZGo2XtR5_0),.dout(w_dff_B_uDWde4n81_0),.clk(gclk));
	jdff dff_B_njBhggTg5_0(.din(w_dff_B_uDWde4n81_0),.dout(w_dff_B_njBhggTg5_0),.clk(gclk));
	jdff dff_B_P5Hzo2Zp1_0(.din(w_dff_B_njBhggTg5_0),.dout(w_dff_B_P5Hzo2Zp1_0),.clk(gclk));
	jdff dff_B_4BfguwV94_0(.din(w_dff_B_P5Hzo2Zp1_0),.dout(w_dff_B_4BfguwV94_0),.clk(gclk));
	jdff dff_B_HkBAUb3b0_0(.din(w_dff_B_4BfguwV94_0),.dout(w_dff_B_HkBAUb3b0_0),.clk(gclk));
	jdff dff_B_ngRyoD7x8_0(.din(w_dff_B_HkBAUb3b0_0),.dout(w_dff_B_ngRyoD7x8_0),.clk(gclk));
	jdff dff_B_oEZXVowk2_0(.din(w_dff_B_ngRyoD7x8_0),.dout(w_dff_B_oEZXVowk2_0),.clk(gclk));
	jdff dff_B_8K6VsHfA3_0(.din(w_dff_B_oEZXVowk2_0),.dout(w_dff_B_8K6VsHfA3_0),.clk(gclk));
	jdff dff_B_l6DYfbgB3_0(.din(w_dff_B_8K6VsHfA3_0),.dout(w_dff_B_l6DYfbgB3_0),.clk(gclk));
	jdff dff_B_mwtPgu9c0_0(.din(w_dff_B_l6DYfbgB3_0),.dout(w_dff_B_mwtPgu9c0_0),.clk(gclk));
	jdff dff_B_xFbV3PoU2_0(.din(w_dff_B_mwtPgu9c0_0),.dout(w_dff_B_xFbV3PoU2_0),.clk(gclk));
	jdff dff_B_AgqJIlai1_0(.din(w_dff_B_xFbV3PoU2_0),.dout(w_dff_B_AgqJIlai1_0),.clk(gclk));
	jdff dff_B_1nPrVcnp2_0(.din(w_dff_B_AgqJIlai1_0),.dout(w_dff_B_1nPrVcnp2_0),.clk(gclk));
	jdff dff_B_5zKXETA53_0(.din(w_dff_B_1nPrVcnp2_0),.dout(w_dff_B_5zKXETA53_0),.clk(gclk));
	jdff dff_B_8epVmzz87_0(.din(w_dff_B_5zKXETA53_0),.dout(w_dff_B_8epVmzz87_0),.clk(gclk));
	jdff dff_B_N5cJ9LNb5_0(.din(w_dff_B_8epVmzz87_0),.dout(w_dff_B_N5cJ9LNb5_0),.clk(gclk));
	jdff dff_B_afPq0GAY8_0(.din(w_dff_B_N5cJ9LNb5_0),.dout(w_dff_B_afPq0GAY8_0),.clk(gclk));
	jdff dff_B_5XU8T3Mw8_0(.din(w_dff_B_afPq0GAY8_0),.dout(w_dff_B_5XU8T3Mw8_0),.clk(gclk));
	jdff dff_B_XQ2xL5tM2_0(.din(w_dff_B_5XU8T3Mw8_0),.dout(w_dff_B_XQ2xL5tM2_0),.clk(gclk));
	jdff dff_B_vzYWFa9T8_0(.din(w_dff_B_XQ2xL5tM2_0),.dout(w_dff_B_vzYWFa9T8_0),.clk(gclk));
	jdff dff_B_nMCaWRfT6_0(.din(w_dff_B_vzYWFa9T8_0),.dout(w_dff_B_nMCaWRfT6_0),.clk(gclk));
	jdff dff_B_m2LfiuhB0_0(.din(w_dff_B_nMCaWRfT6_0),.dout(w_dff_B_m2LfiuhB0_0),.clk(gclk));
	jdff dff_B_RrwnGvqr5_0(.din(w_dff_B_m2LfiuhB0_0),.dout(w_dff_B_RrwnGvqr5_0),.clk(gclk));
	jdff dff_B_unXnc3AO8_0(.din(w_dff_B_RrwnGvqr5_0),.dout(w_dff_B_unXnc3AO8_0),.clk(gclk));
	jdff dff_B_Hu2gvB395_0(.din(w_dff_B_unXnc3AO8_0),.dout(w_dff_B_Hu2gvB395_0),.clk(gclk));
	jdff dff_B_mWU2Bni57_0(.din(w_dff_B_Hu2gvB395_0),.dout(w_dff_B_mWU2Bni57_0),.clk(gclk));
	jdff dff_B_qxljZjVO0_0(.din(w_dff_B_mWU2Bni57_0),.dout(w_dff_B_qxljZjVO0_0),.clk(gclk));
	jdff dff_B_CNui0XvE3_0(.din(w_dff_B_qxljZjVO0_0),.dout(w_dff_B_CNui0XvE3_0),.clk(gclk));
	jdff dff_B_Eo4JERnf8_0(.din(w_dff_B_CNui0XvE3_0),.dout(w_dff_B_Eo4JERnf8_0),.clk(gclk));
	jdff dff_B_d8B3KVR47_0(.din(w_dff_B_Eo4JERnf8_0),.dout(w_dff_B_d8B3KVR47_0),.clk(gclk));
	jdff dff_B_P1cmW4xQ4_0(.din(w_dff_B_d8B3KVR47_0),.dout(w_dff_B_P1cmW4xQ4_0),.clk(gclk));
	jdff dff_B_LBXBeSez1_0(.din(w_dff_B_P1cmW4xQ4_0),.dout(w_dff_B_LBXBeSez1_0),.clk(gclk));
	jdff dff_B_8KmYPTae8_0(.din(w_dff_B_LBXBeSez1_0),.dout(w_dff_B_8KmYPTae8_0),.clk(gclk));
	jdff dff_B_14oMNk0D7_0(.din(w_dff_B_8KmYPTae8_0),.dout(w_dff_B_14oMNk0D7_0),.clk(gclk));
	jdff dff_B_Rnhj953L7_0(.din(w_dff_B_14oMNk0D7_0),.dout(w_dff_B_Rnhj953L7_0),.clk(gclk));
	jdff dff_B_ZvnWeP999_0(.din(w_dff_B_Rnhj953L7_0),.dout(w_dff_B_ZvnWeP999_0),.clk(gclk));
	jdff dff_B_3fAtqGT09_0(.din(w_dff_B_ZvnWeP999_0),.dout(w_dff_B_3fAtqGT09_0),.clk(gclk));
	jdff dff_B_aAhtehik0_0(.din(w_dff_B_3fAtqGT09_0),.dout(w_dff_B_aAhtehik0_0),.clk(gclk));
	jdff dff_B_o6Rq3phW0_0(.din(w_dff_B_aAhtehik0_0),.dout(w_dff_B_o6Rq3phW0_0),.clk(gclk));
	jdff dff_B_cnh7sGxs4_0(.din(w_dff_B_o6Rq3phW0_0),.dout(w_dff_B_cnh7sGxs4_0),.clk(gclk));
	jdff dff_B_UhYaz45r0_0(.din(w_dff_B_cnh7sGxs4_0),.dout(w_dff_B_UhYaz45r0_0),.clk(gclk));
	jdff dff_B_heSdbbWs5_0(.din(w_dff_B_UhYaz45r0_0),.dout(w_dff_B_heSdbbWs5_0),.clk(gclk));
	jdff dff_B_L3uyP2X62_0(.din(w_dff_B_heSdbbWs5_0),.dout(w_dff_B_L3uyP2X62_0),.clk(gclk));
	jdff dff_B_zIWosCQc7_0(.din(w_dff_B_L3uyP2X62_0),.dout(w_dff_B_zIWosCQc7_0),.clk(gclk));
	jdff dff_B_ZNc4ox7c3_0(.din(w_dff_B_zIWosCQc7_0),.dout(w_dff_B_ZNc4ox7c3_0),.clk(gclk));
	jdff dff_B_ZOLbvdtG2_0(.din(w_dff_B_ZNc4ox7c3_0),.dout(w_dff_B_ZOLbvdtG2_0),.clk(gclk));
	jdff dff_B_x1mt1XC68_0(.din(w_dff_B_ZOLbvdtG2_0),.dout(w_dff_B_x1mt1XC68_0),.clk(gclk));
	jdff dff_B_oIFa4bEX1_0(.din(w_dff_B_x1mt1XC68_0),.dout(w_dff_B_oIFa4bEX1_0),.clk(gclk));
	jdff dff_B_iQmPgdEz3_0(.din(w_dff_B_oIFa4bEX1_0),.dout(w_dff_B_iQmPgdEz3_0),.clk(gclk));
	jdff dff_B_Ch1LW24n7_0(.din(w_dff_B_iQmPgdEz3_0),.dout(w_dff_B_Ch1LW24n7_0),.clk(gclk));
	jdff dff_B_rOyHgDks8_0(.din(w_dff_B_Ch1LW24n7_0),.dout(w_dff_B_rOyHgDks8_0),.clk(gclk));
	jdff dff_B_kGDwxasu3_0(.din(w_dff_B_rOyHgDks8_0),.dout(w_dff_B_kGDwxasu3_0),.clk(gclk));
	jdff dff_B_wHLiDIXZ9_0(.din(w_dff_B_kGDwxasu3_0),.dout(w_dff_B_wHLiDIXZ9_0),.clk(gclk));
	jdff dff_B_j1x5kQTT0_0(.din(w_dff_B_wHLiDIXZ9_0),.dout(w_dff_B_j1x5kQTT0_0),.clk(gclk));
	jdff dff_B_uAUjPAjr6_0(.din(w_dff_B_j1x5kQTT0_0),.dout(w_dff_B_uAUjPAjr6_0),.clk(gclk));
	jdff dff_B_rXf4j4Y44_0(.din(w_dff_B_uAUjPAjr6_0),.dout(w_dff_B_rXf4j4Y44_0),.clk(gclk));
	jdff dff_B_nEavyAKv3_0(.din(w_dff_B_rXf4j4Y44_0),.dout(w_dff_B_nEavyAKv3_0),.clk(gclk));
	jdff dff_B_QcxVJFj87_0(.din(w_dff_B_nEavyAKv3_0),.dout(w_dff_B_QcxVJFj87_0),.clk(gclk));
	jdff dff_B_LrzuCVep6_0(.din(w_dff_B_QcxVJFj87_0),.dout(w_dff_B_LrzuCVep6_0),.clk(gclk));
	jdff dff_B_J9zqpGSM3_0(.din(w_dff_B_LrzuCVep6_0),.dout(w_dff_B_J9zqpGSM3_0),.clk(gclk));
	jdff dff_B_mAq3ZGyQ2_0(.din(w_dff_B_J9zqpGSM3_0),.dout(w_dff_B_mAq3ZGyQ2_0),.clk(gclk));
	jdff dff_B_JSc81Qhc2_0(.din(w_dff_B_mAq3ZGyQ2_0),.dout(w_dff_B_JSc81Qhc2_0),.clk(gclk));
	jdff dff_B_sYq6oIB27_1(.din(n1092),.dout(w_dff_B_sYq6oIB27_1),.clk(gclk));
	jdff dff_B_Mc2PPan17_1(.din(w_dff_B_sYq6oIB27_1),.dout(w_dff_B_Mc2PPan17_1),.clk(gclk));
	jdff dff_B_4qKbGJTO6_1(.din(w_dff_B_Mc2PPan17_1),.dout(w_dff_B_4qKbGJTO6_1),.clk(gclk));
	jdff dff_B_14xh7Ujc8_1(.din(w_dff_B_4qKbGJTO6_1),.dout(w_dff_B_14xh7Ujc8_1),.clk(gclk));
	jdff dff_B_xwiTDYel3_1(.din(w_dff_B_14xh7Ujc8_1),.dout(w_dff_B_xwiTDYel3_1),.clk(gclk));
	jdff dff_B_rTuSd1994_1(.din(w_dff_B_xwiTDYel3_1),.dout(w_dff_B_rTuSd1994_1),.clk(gclk));
	jdff dff_B_8cR0rBkV4_1(.din(w_dff_B_rTuSd1994_1),.dout(w_dff_B_8cR0rBkV4_1),.clk(gclk));
	jdff dff_B_5JI2EuHq8_1(.din(w_dff_B_8cR0rBkV4_1),.dout(w_dff_B_5JI2EuHq8_1),.clk(gclk));
	jdff dff_B_DZkDuAc95_1(.din(w_dff_B_5JI2EuHq8_1),.dout(w_dff_B_DZkDuAc95_1),.clk(gclk));
	jdff dff_B_ATEK1pgC7_1(.din(w_dff_B_DZkDuAc95_1),.dout(w_dff_B_ATEK1pgC7_1),.clk(gclk));
	jdff dff_B_U5pTLMyQ0_1(.din(w_dff_B_ATEK1pgC7_1),.dout(w_dff_B_U5pTLMyQ0_1),.clk(gclk));
	jdff dff_B_S9U0rcYm5_1(.din(w_dff_B_U5pTLMyQ0_1),.dout(w_dff_B_S9U0rcYm5_1),.clk(gclk));
	jdff dff_B_cfPrY5Fi9_1(.din(w_dff_B_S9U0rcYm5_1),.dout(w_dff_B_cfPrY5Fi9_1),.clk(gclk));
	jdff dff_B_aXfLR1ZS2_1(.din(w_dff_B_cfPrY5Fi9_1),.dout(w_dff_B_aXfLR1ZS2_1),.clk(gclk));
	jdff dff_B_IKfIb25a1_1(.din(w_dff_B_aXfLR1ZS2_1),.dout(w_dff_B_IKfIb25a1_1),.clk(gclk));
	jdff dff_B_389xdMPT9_1(.din(w_dff_B_IKfIb25a1_1),.dout(w_dff_B_389xdMPT9_1),.clk(gclk));
	jdff dff_B_3VHdWk4Q2_1(.din(w_dff_B_389xdMPT9_1),.dout(w_dff_B_3VHdWk4Q2_1),.clk(gclk));
	jdff dff_B_5nYmQITp2_1(.din(w_dff_B_3VHdWk4Q2_1),.dout(w_dff_B_5nYmQITp2_1),.clk(gclk));
	jdff dff_B_oxm5N6Bn3_1(.din(w_dff_B_5nYmQITp2_1),.dout(w_dff_B_oxm5N6Bn3_1),.clk(gclk));
	jdff dff_B_qWa1F2rv8_1(.din(w_dff_B_oxm5N6Bn3_1),.dout(w_dff_B_qWa1F2rv8_1),.clk(gclk));
	jdff dff_B_repZVBIo9_1(.din(w_dff_B_qWa1F2rv8_1),.dout(w_dff_B_repZVBIo9_1),.clk(gclk));
	jdff dff_B_TmJcs3DT1_1(.din(w_dff_B_repZVBIo9_1),.dout(w_dff_B_TmJcs3DT1_1),.clk(gclk));
	jdff dff_B_cyz57FfY7_1(.din(w_dff_B_TmJcs3DT1_1),.dout(w_dff_B_cyz57FfY7_1),.clk(gclk));
	jdff dff_B_55ap0eZ79_1(.din(w_dff_B_cyz57FfY7_1),.dout(w_dff_B_55ap0eZ79_1),.clk(gclk));
	jdff dff_B_qv9xgGOe2_1(.din(w_dff_B_55ap0eZ79_1),.dout(w_dff_B_qv9xgGOe2_1),.clk(gclk));
	jdff dff_B_GUSy8BVL6_1(.din(w_dff_B_qv9xgGOe2_1),.dout(w_dff_B_GUSy8BVL6_1),.clk(gclk));
	jdff dff_B_Tfg8qDL46_1(.din(w_dff_B_GUSy8BVL6_1),.dout(w_dff_B_Tfg8qDL46_1),.clk(gclk));
	jdff dff_B_QRI6PbSb5_1(.din(w_dff_B_Tfg8qDL46_1),.dout(w_dff_B_QRI6PbSb5_1),.clk(gclk));
	jdff dff_B_xAuy5jje1_1(.din(w_dff_B_QRI6PbSb5_1),.dout(w_dff_B_xAuy5jje1_1),.clk(gclk));
	jdff dff_B_dmKlRpZe2_1(.din(w_dff_B_xAuy5jje1_1),.dout(w_dff_B_dmKlRpZe2_1),.clk(gclk));
	jdff dff_B_64Fs2Iib3_1(.din(w_dff_B_dmKlRpZe2_1),.dout(w_dff_B_64Fs2Iib3_1),.clk(gclk));
	jdff dff_B_2K2x6IeT6_1(.din(w_dff_B_64Fs2Iib3_1),.dout(w_dff_B_2K2x6IeT6_1),.clk(gclk));
	jdff dff_B_SAKsbJUN6_1(.din(w_dff_B_2K2x6IeT6_1),.dout(w_dff_B_SAKsbJUN6_1),.clk(gclk));
	jdff dff_B_E07jwBMe0_1(.din(w_dff_B_SAKsbJUN6_1),.dout(w_dff_B_E07jwBMe0_1),.clk(gclk));
	jdff dff_B_kMxHPedC1_1(.din(w_dff_B_E07jwBMe0_1),.dout(w_dff_B_kMxHPedC1_1),.clk(gclk));
	jdff dff_B_JYngolCI4_1(.din(w_dff_B_kMxHPedC1_1),.dout(w_dff_B_JYngolCI4_1),.clk(gclk));
	jdff dff_B_ODzATTYR9_1(.din(w_dff_B_JYngolCI4_1),.dout(w_dff_B_ODzATTYR9_1),.clk(gclk));
	jdff dff_B_GnLQI6qe3_1(.din(w_dff_B_ODzATTYR9_1),.dout(w_dff_B_GnLQI6qe3_1),.clk(gclk));
	jdff dff_B_Z0zr7KT67_1(.din(w_dff_B_GnLQI6qe3_1),.dout(w_dff_B_Z0zr7KT67_1),.clk(gclk));
	jdff dff_B_ExfL3PUW8_1(.din(w_dff_B_Z0zr7KT67_1),.dout(w_dff_B_ExfL3PUW8_1),.clk(gclk));
	jdff dff_B_GNT1NYBN3_1(.din(w_dff_B_ExfL3PUW8_1),.dout(w_dff_B_GNT1NYBN3_1),.clk(gclk));
	jdff dff_B_uomdK2v57_1(.din(w_dff_B_GNT1NYBN3_1),.dout(w_dff_B_uomdK2v57_1),.clk(gclk));
	jdff dff_B_qRHjwwew8_1(.din(w_dff_B_uomdK2v57_1),.dout(w_dff_B_qRHjwwew8_1),.clk(gclk));
	jdff dff_B_nB5crXne1_1(.din(w_dff_B_qRHjwwew8_1),.dout(w_dff_B_nB5crXne1_1),.clk(gclk));
	jdff dff_B_kZAoHPhN5_1(.din(w_dff_B_nB5crXne1_1),.dout(w_dff_B_kZAoHPhN5_1),.clk(gclk));
	jdff dff_B_cxsi7iuI6_1(.din(w_dff_B_kZAoHPhN5_1),.dout(w_dff_B_cxsi7iuI6_1),.clk(gclk));
	jdff dff_B_pf5jKgF90_1(.din(w_dff_B_cxsi7iuI6_1),.dout(w_dff_B_pf5jKgF90_1),.clk(gclk));
	jdff dff_B_VPlu4Mi47_1(.din(w_dff_B_pf5jKgF90_1),.dout(w_dff_B_VPlu4Mi47_1),.clk(gclk));
	jdff dff_B_H3zG7Jxj5_1(.din(w_dff_B_VPlu4Mi47_1),.dout(w_dff_B_H3zG7Jxj5_1),.clk(gclk));
	jdff dff_B_VEUU7NPZ3_1(.din(w_dff_B_H3zG7Jxj5_1),.dout(w_dff_B_VEUU7NPZ3_1),.clk(gclk));
	jdff dff_B_oIkXknC90_1(.din(w_dff_B_VEUU7NPZ3_1),.dout(w_dff_B_oIkXknC90_1),.clk(gclk));
	jdff dff_B_6s7AcXor9_1(.din(w_dff_B_oIkXknC90_1),.dout(w_dff_B_6s7AcXor9_1),.clk(gclk));
	jdff dff_B_SwbCaKMk0_1(.din(w_dff_B_6s7AcXor9_1),.dout(w_dff_B_SwbCaKMk0_1),.clk(gclk));
	jdff dff_B_S9QDlWnx4_1(.din(w_dff_B_SwbCaKMk0_1),.dout(w_dff_B_S9QDlWnx4_1),.clk(gclk));
	jdff dff_B_pdKY1lxM4_1(.din(w_dff_B_S9QDlWnx4_1),.dout(w_dff_B_pdKY1lxM4_1),.clk(gclk));
	jdff dff_B_u3lptrnf8_1(.din(w_dff_B_pdKY1lxM4_1),.dout(w_dff_B_u3lptrnf8_1),.clk(gclk));
	jdff dff_B_GbBouQ5h7_1(.din(w_dff_B_u3lptrnf8_1),.dout(w_dff_B_GbBouQ5h7_1),.clk(gclk));
	jdff dff_B_EI245wFH6_1(.din(w_dff_B_GbBouQ5h7_1),.dout(w_dff_B_EI245wFH6_1),.clk(gclk));
	jdff dff_B_ETIGfcFn8_1(.din(w_dff_B_EI245wFH6_1),.dout(w_dff_B_ETIGfcFn8_1),.clk(gclk));
	jdff dff_B_2AMTPYFz5_1(.din(w_dff_B_ETIGfcFn8_1),.dout(w_dff_B_2AMTPYFz5_1),.clk(gclk));
	jdff dff_B_1HLApl003_1(.din(w_dff_B_2AMTPYFz5_1),.dout(w_dff_B_1HLApl003_1),.clk(gclk));
	jdff dff_B_8JnTbCBE4_1(.din(w_dff_B_1HLApl003_1),.dout(w_dff_B_8JnTbCBE4_1),.clk(gclk));
	jdff dff_B_N5jV3Jlw4_1(.din(w_dff_B_8JnTbCBE4_1),.dout(w_dff_B_N5jV3Jlw4_1),.clk(gclk));
	jdff dff_B_34Yuk4Sg7_1(.din(w_dff_B_N5jV3Jlw4_1),.dout(w_dff_B_34Yuk4Sg7_1),.clk(gclk));
	jdff dff_B_E7KxLBXn5_1(.din(w_dff_B_34Yuk4Sg7_1),.dout(w_dff_B_E7KxLBXn5_1),.clk(gclk));
	jdff dff_B_HAqv7guS4_1(.din(w_dff_B_E7KxLBXn5_1),.dout(w_dff_B_HAqv7guS4_1),.clk(gclk));
	jdff dff_B_ZEdYL15L5_1(.din(w_dff_B_HAqv7guS4_1),.dout(w_dff_B_ZEdYL15L5_1),.clk(gclk));
	jdff dff_B_z2K6vSV76_1(.din(w_dff_B_ZEdYL15L5_1),.dout(w_dff_B_z2K6vSV76_1),.clk(gclk));
	jdff dff_B_EbPlB7874_1(.din(w_dff_B_z2K6vSV76_1),.dout(w_dff_B_EbPlB7874_1),.clk(gclk));
	jdff dff_B_aene9t648_1(.din(w_dff_B_EbPlB7874_1),.dout(w_dff_B_aene9t648_1),.clk(gclk));
	jdff dff_B_8Henj0RT7_1(.din(w_dff_B_aene9t648_1),.dout(w_dff_B_8Henj0RT7_1),.clk(gclk));
	jdff dff_B_lSUaYgkw1_1(.din(w_dff_B_8Henj0RT7_1),.dout(w_dff_B_lSUaYgkw1_1),.clk(gclk));
	jdff dff_B_W1RGT3kX4_1(.din(w_dff_B_lSUaYgkw1_1),.dout(w_dff_B_W1RGT3kX4_1),.clk(gclk));
	jdff dff_B_L2Yyhw4X1_1(.din(w_dff_B_W1RGT3kX4_1),.dout(w_dff_B_L2Yyhw4X1_1),.clk(gclk));
	jdff dff_B_OAK4GISu9_1(.din(w_dff_B_L2Yyhw4X1_1),.dout(w_dff_B_OAK4GISu9_1),.clk(gclk));
	jdff dff_B_n6MpM0oR2_1(.din(w_dff_B_OAK4GISu9_1),.dout(w_dff_B_n6MpM0oR2_1),.clk(gclk));
	jdff dff_B_WgCHhUfe4_1(.din(w_dff_B_n6MpM0oR2_1),.dout(w_dff_B_WgCHhUfe4_1),.clk(gclk));
	jdff dff_B_V24btCTU1_1(.din(w_dff_B_WgCHhUfe4_1),.dout(w_dff_B_V24btCTU1_1),.clk(gclk));
	jdff dff_B_46iaAK8d8_1(.din(w_dff_B_V24btCTU1_1),.dout(w_dff_B_46iaAK8d8_1),.clk(gclk));
	jdff dff_B_GRRWWKgJ3_1(.din(w_dff_B_46iaAK8d8_1),.dout(w_dff_B_GRRWWKgJ3_1),.clk(gclk));
	jdff dff_B_LSoTwvbM4_1(.din(w_dff_B_GRRWWKgJ3_1),.dout(w_dff_B_LSoTwvbM4_1),.clk(gclk));
	jdff dff_B_5H1TghRK9_1(.din(w_dff_B_LSoTwvbM4_1),.dout(w_dff_B_5H1TghRK9_1),.clk(gclk));
	jdff dff_B_nYUPnOY41_1(.din(w_dff_B_5H1TghRK9_1),.dout(w_dff_B_nYUPnOY41_1),.clk(gclk));
	jdff dff_B_WFoDYRVC3_1(.din(w_dff_B_nYUPnOY41_1),.dout(w_dff_B_WFoDYRVC3_1),.clk(gclk));
	jdff dff_B_m5g4kFHf0_1(.din(w_dff_B_WFoDYRVC3_1),.dout(w_dff_B_m5g4kFHf0_1),.clk(gclk));
	jdff dff_B_uYMdIVgf0_1(.din(w_dff_B_m5g4kFHf0_1),.dout(w_dff_B_uYMdIVgf0_1),.clk(gclk));
	jdff dff_B_SVUFnekn2_1(.din(w_dff_B_uYMdIVgf0_1),.dout(w_dff_B_SVUFnekn2_1),.clk(gclk));
	jdff dff_B_6OfZvN8s7_1(.din(w_dff_B_SVUFnekn2_1),.dout(w_dff_B_6OfZvN8s7_1),.clk(gclk));
	jdff dff_B_ac5b9gd27_1(.din(w_dff_B_6OfZvN8s7_1),.dout(w_dff_B_ac5b9gd27_1),.clk(gclk));
	jdff dff_B_9oCCIevO5_1(.din(w_dff_B_ac5b9gd27_1),.dout(w_dff_B_9oCCIevO5_1),.clk(gclk));
	jdff dff_B_6rRwW7Ws4_1(.din(w_dff_B_9oCCIevO5_1),.dout(w_dff_B_6rRwW7Ws4_1),.clk(gclk));
	jdff dff_B_tY1rLmmh2_1(.din(w_dff_B_6rRwW7Ws4_1),.dout(w_dff_B_tY1rLmmh2_1),.clk(gclk));
	jdff dff_B_OCEhKZzF9_1(.din(w_dff_B_tY1rLmmh2_1),.dout(w_dff_B_OCEhKZzF9_1),.clk(gclk));
	jdff dff_B_Et1lDeqa9_1(.din(w_dff_B_OCEhKZzF9_1),.dout(w_dff_B_Et1lDeqa9_1),.clk(gclk));
	jdff dff_B_1VOxYzwg9_1(.din(w_dff_B_Et1lDeqa9_1),.dout(w_dff_B_1VOxYzwg9_1),.clk(gclk));
	jdff dff_B_64aPibxn5_1(.din(w_dff_B_1VOxYzwg9_1),.dout(w_dff_B_64aPibxn5_1),.clk(gclk));
	jdff dff_B_eKWjpM350_1(.din(w_dff_B_64aPibxn5_1),.dout(w_dff_B_eKWjpM350_1),.clk(gclk));
	jdff dff_B_V500e5aP3_1(.din(w_dff_B_eKWjpM350_1),.dout(w_dff_B_V500e5aP3_1),.clk(gclk));
	jdff dff_B_U74oms4w5_1(.din(w_dff_B_V500e5aP3_1),.dout(w_dff_B_U74oms4w5_1),.clk(gclk));
	jdff dff_B_p8i8DXbS3_1(.din(w_dff_B_U74oms4w5_1),.dout(w_dff_B_p8i8DXbS3_1),.clk(gclk));
	jdff dff_B_bSrTy1ev8_1(.din(w_dff_B_p8i8DXbS3_1),.dout(w_dff_B_bSrTy1ev8_1),.clk(gclk));
	jdff dff_B_aBlLHLBO6_1(.din(w_dff_B_bSrTy1ev8_1),.dout(w_dff_B_aBlLHLBO6_1),.clk(gclk));
	jdff dff_B_Bs4WsX2g9_1(.din(w_dff_B_aBlLHLBO6_1),.dout(w_dff_B_Bs4WsX2g9_1),.clk(gclk));
	jdff dff_B_4JDGpC0g4_1(.din(w_dff_B_Bs4WsX2g9_1),.dout(w_dff_B_4JDGpC0g4_1),.clk(gclk));
	jdff dff_B_p2Dyonl82_1(.din(w_dff_B_4JDGpC0g4_1),.dout(w_dff_B_p2Dyonl82_1),.clk(gclk));
	jdff dff_B_BBY7MKTB9_1(.din(w_dff_B_p2Dyonl82_1),.dout(w_dff_B_BBY7MKTB9_1),.clk(gclk));
	jdff dff_B_r2RFdo4Y5_1(.din(w_dff_B_BBY7MKTB9_1),.dout(w_dff_B_r2RFdo4Y5_1),.clk(gclk));
	jdff dff_B_LIENfJEl4_1(.din(w_dff_B_r2RFdo4Y5_1),.dout(w_dff_B_LIENfJEl4_1),.clk(gclk));
	jdff dff_B_ZHJlxTIa7_1(.din(w_dff_B_LIENfJEl4_1),.dout(w_dff_B_ZHJlxTIa7_1),.clk(gclk));
	jdff dff_B_dGDIGRuM0_1(.din(w_dff_B_ZHJlxTIa7_1),.dout(w_dff_B_dGDIGRuM0_1),.clk(gclk));
	jdff dff_B_TeLvXY2Y6_1(.din(w_dff_B_dGDIGRuM0_1),.dout(w_dff_B_TeLvXY2Y6_1),.clk(gclk));
	jdff dff_B_Izmrb4xg5_1(.din(w_dff_B_TeLvXY2Y6_1),.dout(w_dff_B_Izmrb4xg5_1),.clk(gclk));
	jdff dff_B_tuOP7eqL8_1(.din(w_dff_B_Izmrb4xg5_1),.dout(w_dff_B_tuOP7eqL8_1),.clk(gclk));
	jdff dff_B_dMzdyEiI6_1(.din(w_dff_B_tuOP7eqL8_1),.dout(w_dff_B_dMzdyEiI6_1),.clk(gclk));
	jdff dff_B_hB0Mxx1g3_1(.din(w_dff_B_dMzdyEiI6_1),.dout(w_dff_B_hB0Mxx1g3_1),.clk(gclk));
	jdff dff_B_hhejUK2T5_1(.din(w_dff_B_hB0Mxx1g3_1),.dout(w_dff_B_hhejUK2T5_1),.clk(gclk));
	jdff dff_B_W6b68rBH3_1(.din(w_dff_B_hhejUK2T5_1),.dout(w_dff_B_W6b68rBH3_1),.clk(gclk));
	jdff dff_B_hW63y0Sx4_1(.din(w_dff_B_W6b68rBH3_1),.dout(w_dff_B_hW63y0Sx4_1),.clk(gclk));
	jdff dff_B_syFTwmB93_0(.din(n1093),.dout(w_dff_B_syFTwmB93_0),.clk(gclk));
	jdff dff_B_rGkd5r7P5_0(.din(w_dff_B_syFTwmB93_0),.dout(w_dff_B_rGkd5r7P5_0),.clk(gclk));
	jdff dff_B_OlmzySVc6_0(.din(w_dff_B_rGkd5r7P5_0),.dout(w_dff_B_OlmzySVc6_0),.clk(gclk));
	jdff dff_B_Ut9vB0XY6_0(.din(w_dff_B_OlmzySVc6_0),.dout(w_dff_B_Ut9vB0XY6_0),.clk(gclk));
	jdff dff_B_EoLinNfp9_0(.din(w_dff_B_Ut9vB0XY6_0),.dout(w_dff_B_EoLinNfp9_0),.clk(gclk));
	jdff dff_B_6j2dYUEX7_0(.din(w_dff_B_EoLinNfp9_0),.dout(w_dff_B_6j2dYUEX7_0),.clk(gclk));
	jdff dff_B_z2173c6s1_0(.din(w_dff_B_6j2dYUEX7_0),.dout(w_dff_B_z2173c6s1_0),.clk(gclk));
	jdff dff_B_On7zB16x4_0(.din(w_dff_B_z2173c6s1_0),.dout(w_dff_B_On7zB16x4_0),.clk(gclk));
	jdff dff_B_biyyJnSh6_0(.din(w_dff_B_On7zB16x4_0),.dout(w_dff_B_biyyJnSh6_0),.clk(gclk));
	jdff dff_B_TezYp0Ra8_0(.din(w_dff_B_biyyJnSh6_0),.dout(w_dff_B_TezYp0Ra8_0),.clk(gclk));
	jdff dff_B_braLNV6O5_0(.din(w_dff_B_TezYp0Ra8_0),.dout(w_dff_B_braLNV6O5_0),.clk(gclk));
	jdff dff_B_ZeUtcFsF7_0(.din(w_dff_B_braLNV6O5_0),.dout(w_dff_B_ZeUtcFsF7_0),.clk(gclk));
	jdff dff_B_zC3DyTHw6_0(.din(w_dff_B_ZeUtcFsF7_0),.dout(w_dff_B_zC3DyTHw6_0),.clk(gclk));
	jdff dff_B_SvOZJ9Gi3_0(.din(w_dff_B_zC3DyTHw6_0),.dout(w_dff_B_SvOZJ9Gi3_0),.clk(gclk));
	jdff dff_B_ky4sKzd06_0(.din(w_dff_B_SvOZJ9Gi3_0),.dout(w_dff_B_ky4sKzd06_0),.clk(gclk));
	jdff dff_B_gE3zK0w63_0(.din(w_dff_B_ky4sKzd06_0),.dout(w_dff_B_gE3zK0w63_0),.clk(gclk));
	jdff dff_B_YAnSMdnK3_0(.din(w_dff_B_gE3zK0w63_0),.dout(w_dff_B_YAnSMdnK3_0),.clk(gclk));
	jdff dff_B_9Q80FKWm6_0(.din(w_dff_B_YAnSMdnK3_0),.dout(w_dff_B_9Q80FKWm6_0),.clk(gclk));
	jdff dff_B_TR0D03kd1_0(.din(w_dff_B_9Q80FKWm6_0),.dout(w_dff_B_TR0D03kd1_0),.clk(gclk));
	jdff dff_B_GRLNTJPk4_0(.din(w_dff_B_TR0D03kd1_0),.dout(w_dff_B_GRLNTJPk4_0),.clk(gclk));
	jdff dff_B_22X2GU6B4_0(.din(w_dff_B_GRLNTJPk4_0),.dout(w_dff_B_22X2GU6B4_0),.clk(gclk));
	jdff dff_B_b5lIMHw38_0(.din(w_dff_B_22X2GU6B4_0),.dout(w_dff_B_b5lIMHw38_0),.clk(gclk));
	jdff dff_B_K1i8waze1_0(.din(w_dff_B_b5lIMHw38_0),.dout(w_dff_B_K1i8waze1_0),.clk(gclk));
	jdff dff_B_XFLWQoGc7_0(.din(w_dff_B_K1i8waze1_0),.dout(w_dff_B_XFLWQoGc7_0),.clk(gclk));
	jdff dff_B_GSByVAd25_0(.din(w_dff_B_XFLWQoGc7_0),.dout(w_dff_B_GSByVAd25_0),.clk(gclk));
	jdff dff_B_MtzmmXRR6_0(.din(w_dff_B_GSByVAd25_0),.dout(w_dff_B_MtzmmXRR6_0),.clk(gclk));
	jdff dff_B_cbNpikyc7_0(.din(w_dff_B_MtzmmXRR6_0),.dout(w_dff_B_cbNpikyc7_0),.clk(gclk));
	jdff dff_B_YNm8l35B3_0(.din(w_dff_B_cbNpikyc7_0),.dout(w_dff_B_YNm8l35B3_0),.clk(gclk));
	jdff dff_B_7apRK40L8_0(.din(w_dff_B_YNm8l35B3_0),.dout(w_dff_B_7apRK40L8_0),.clk(gclk));
	jdff dff_B_XIt328QY0_0(.din(w_dff_B_7apRK40L8_0),.dout(w_dff_B_XIt328QY0_0),.clk(gclk));
	jdff dff_B_7l6hmQ2M6_0(.din(w_dff_B_XIt328QY0_0),.dout(w_dff_B_7l6hmQ2M6_0),.clk(gclk));
	jdff dff_B_pfmQUzfS4_0(.din(w_dff_B_7l6hmQ2M6_0),.dout(w_dff_B_pfmQUzfS4_0),.clk(gclk));
	jdff dff_B_IPy17bNt9_0(.din(w_dff_B_pfmQUzfS4_0),.dout(w_dff_B_IPy17bNt9_0),.clk(gclk));
	jdff dff_B_1Et8djZy2_0(.din(w_dff_B_IPy17bNt9_0),.dout(w_dff_B_1Et8djZy2_0),.clk(gclk));
	jdff dff_B_fCD8ZvnQ2_0(.din(w_dff_B_1Et8djZy2_0),.dout(w_dff_B_fCD8ZvnQ2_0),.clk(gclk));
	jdff dff_B_l3TqqqL40_0(.din(w_dff_B_fCD8ZvnQ2_0),.dout(w_dff_B_l3TqqqL40_0),.clk(gclk));
	jdff dff_B_5UKu6m229_0(.din(w_dff_B_l3TqqqL40_0),.dout(w_dff_B_5UKu6m229_0),.clk(gclk));
	jdff dff_B_FHMUvI1i3_0(.din(w_dff_B_5UKu6m229_0),.dout(w_dff_B_FHMUvI1i3_0),.clk(gclk));
	jdff dff_B_tH7rGPYO5_0(.din(w_dff_B_FHMUvI1i3_0),.dout(w_dff_B_tH7rGPYO5_0),.clk(gclk));
	jdff dff_B_Lj3TNSSx7_0(.din(w_dff_B_tH7rGPYO5_0),.dout(w_dff_B_Lj3TNSSx7_0),.clk(gclk));
	jdff dff_B_zviujcVA6_0(.din(w_dff_B_Lj3TNSSx7_0),.dout(w_dff_B_zviujcVA6_0),.clk(gclk));
	jdff dff_B_rWTKYZYJ1_0(.din(w_dff_B_zviujcVA6_0),.dout(w_dff_B_rWTKYZYJ1_0),.clk(gclk));
	jdff dff_B_6WqjrJA54_0(.din(w_dff_B_rWTKYZYJ1_0),.dout(w_dff_B_6WqjrJA54_0),.clk(gclk));
	jdff dff_B_ZHDe1QPz3_0(.din(w_dff_B_6WqjrJA54_0),.dout(w_dff_B_ZHDe1QPz3_0),.clk(gclk));
	jdff dff_B_Q4rko9hu3_0(.din(w_dff_B_ZHDe1QPz3_0),.dout(w_dff_B_Q4rko9hu3_0),.clk(gclk));
	jdff dff_B_2O1AmU713_0(.din(w_dff_B_Q4rko9hu3_0),.dout(w_dff_B_2O1AmU713_0),.clk(gclk));
	jdff dff_B_NFRIOZh67_0(.din(w_dff_B_2O1AmU713_0),.dout(w_dff_B_NFRIOZh67_0),.clk(gclk));
	jdff dff_B_lo9ZQOI16_0(.din(w_dff_B_NFRIOZh67_0),.dout(w_dff_B_lo9ZQOI16_0),.clk(gclk));
	jdff dff_B_ofOAyfxh7_0(.din(w_dff_B_lo9ZQOI16_0),.dout(w_dff_B_ofOAyfxh7_0),.clk(gclk));
	jdff dff_B_fzgk1dLt9_0(.din(w_dff_B_ofOAyfxh7_0),.dout(w_dff_B_fzgk1dLt9_0),.clk(gclk));
	jdff dff_B_HS7BREav1_0(.din(w_dff_B_fzgk1dLt9_0),.dout(w_dff_B_HS7BREav1_0),.clk(gclk));
	jdff dff_B_uD5oK2bF2_0(.din(w_dff_B_HS7BREav1_0),.dout(w_dff_B_uD5oK2bF2_0),.clk(gclk));
	jdff dff_B_eOv37QLa0_0(.din(w_dff_B_uD5oK2bF2_0),.dout(w_dff_B_eOv37QLa0_0),.clk(gclk));
	jdff dff_B_8bTL8iVs7_0(.din(w_dff_B_eOv37QLa0_0),.dout(w_dff_B_8bTL8iVs7_0),.clk(gclk));
	jdff dff_B_Yn0zx3027_0(.din(w_dff_B_8bTL8iVs7_0),.dout(w_dff_B_Yn0zx3027_0),.clk(gclk));
	jdff dff_B_z5vT4OBK5_0(.din(w_dff_B_Yn0zx3027_0),.dout(w_dff_B_z5vT4OBK5_0),.clk(gclk));
	jdff dff_B_g87oetmx9_0(.din(w_dff_B_z5vT4OBK5_0),.dout(w_dff_B_g87oetmx9_0),.clk(gclk));
	jdff dff_B_gzj3X2n83_0(.din(w_dff_B_g87oetmx9_0),.dout(w_dff_B_gzj3X2n83_0),.clk(gclk));
	jdff dff_B_xICX0ZDl7_0(.din(w_dff_B_gzj3X2n83_0),.dout(w_dff_B_xICX0ZDl7_0),.clk(gclk));
	jdff dff_B_sBJqN9m51_0(.din(w_dff_B_xICX0ZDl7_0),.dout(w_dff_B_sBJqN9m51_0),.clk(gclk));
	jdff dff_B_VH8U2p3E4_0(.din(w_dff_B_sBJqN9m51_0),.dout(w_dff_B_VH8U2p3E4_0),.clk(gclk));
	jdff dff_B_SZttFc7V6_0(.din(w_dff_B_VH8U2p3E4_0),.dout(w_dff_B_SZttFc7V6_0),.clk(gclk));
	jdff dff_B_JjBTIVlq7_0(.din(w_dff_B_SZttFc7V6_0),.dout(w_dff_B_JjBTIVlq7_0),.clk(gclk));
	jdff dff_B_k8niOOyu4_0(.din(w_dff_B_JjBTIVlq7_0),.dout(w_dff_B_k8niOOyu4_0),.clk(gclk));
	jdff dff_B_XnQzF0iA4_0(.din(w_dff_B_k8niOOyu4_0),.dout(w_dff_B_XnQzF0iA4_0),.clk(gclk));
	jdff dff_B_RegjiEZj8_0(.din(w_dff_B_XnQzF0iA4_0),.dout(w_dff_B_RegjiEZj8_0),.clk(gclk));
	jdff dff_B_NybTSBVG7_0(.din(w_dff_B_RegjiEZj8_0),.dout(w_dff_B_NybTSBVG7_0),.clk(gclk));
	jdff dff_B_3WTVIihh4_0(.din(w_dff_B_NybTSBVG7_0),.dout(w_dff_B_3WTVIihh4_0),.clk(gclk));
	jdff dff_B_T8lG7MNp5_0(.din(w_dff_B_3WTVIihh4_0),.dout(w_dff_B_T8lG7MNp5_0),.clk(gclk));
	jdff dff_B_5ZteBW1k8_0(.din(w_dff_B_T8lG7MNp5_0),.dout(w_dff_B_5ZteBW1k8_0),.clk(gclk));
	jdff dff_B_TldflRhm2_0(.din(w_dff_B_5ZteBW1k8_0),.dout(w_dff_B_TldflRhm2_0),.clk(gclk));
	jdff dff_B_r1gEPlLE9_0(.din(w_dff_B_TldflRhm2_0),.dout(w_dff_B_r1gEPlLE9_0),.clk(gclk));
	jdff dff_B_yjFeG0Ie1_0(.din(w_dff_B_r1gEPlLE9_0),.dout(w_dff_B_yjFeG0Ie1_0),.clk(gclk));
	jdff dff_B_pvQFLMEh1_0(.din(w_dff_B_yjFeG0Ie1_0),.dout(w_dff_B_pvQFLMEh1_0),.clk(gclk));
	jdff dff_B_tN67ZL9p9_0(.din(w_dff_B_pvQFLMEh1_0),.dout(w_dff_B_tN67ZL9p9_0),.clk(gclk));
	jdff dff_B_2y2p9ZtR8_0(.din(w_dff_B_tN67ZL9p9_0),.dout(w_dff_B_2y2p9ZtR8_0),.clk(gclk));
	jdff dff_B_oCxJMgs76_0(.din(w_dff_B_2y2p9ZtR8_0),.dout(w_dff_B_oCxJMgs76_0),.clk(gclk));
	jdff dff_B_QWiCdKsj9_0(.din(w_dff_B_oCxJMgs76_0),.dout(w_dff_B_QWiCdKsj9_0),.clk(gclk));
	jdff dff_B_yaSwftAH4_0(.din(w_dff_B_QWiCdKsj9_0),.dout(w_dff_B_yaSwftAH4_0),.clk(gclk));
	jdff dff_B_tpsQhyHM6_0(.din(w_dff_B_yaSwftAH4_0),.dout(w_dff_B_tpsQhyHM6_0),.clk(gclk));
	jdff dff_B_TU5WsVp09_0(.din(w_dff_B_tpsQhyHM6_0),.dout(w_dff_B_TU5WsVp09_0),.clk(gclk));
	jdff dff_B_VATC0ZSr1_0(.din(w_dff_B_TU5WsVp09_0),.dout(w_dff_B_VATC0ZSr1_0),.clk(gclk));
	jdff dff_B_QbGTHADZ6_0(.din(w_dff_B_VATC0ZSr1_0),.dout(w_dff_B_QbGTHADZ6_0),.clk(gclk));
	jdff dff_B_sT7RScMQ8_0(.din(w_dff_B_QbGTHADZ6_0),.dout(w_dff_B_sT7RScMQ8_0),.clk(gclk));
	jdff dff_B_yKyhJFUi5_0(.din(w_dff_B_sT7RScMQ8_0),.dout(w_dff_B_yKyhJFUi5_0),.clk(gclk));
	jdff dff_B_fFXzhb695_0(.din(w_dff_B_yKyhJFUi5_0),.dout(w_dff_B_fFXzhb695_0),.clk(gclk));
	jdff dff_B_pYbeUMXS7_0(.din(w_dff_B_fFXzhb695_0),.dout(w_dff_B_pYbeUMXS7_0),.clk(gclk));
	jdff dff_B_P25KHeJ97_0(.din(w_dff_B_pYbeUMXS7_0),.dout(w_dff_B_P25KHeJ97_0),.clk(gclk));
	jdff dff_B_4ghMgmNn1_0(.din(w_dff_B_P25KHeJ97_0),.dout(w_dff_B_4ghMgmNn1_0),.clk(gclk));
	jdff dff_B_FaRzaNcD9_0(.din(w_dff_B_4ghMgmNn1_0),.dout(w_dff_B_FaRzaNcD9_0),.clk(gclk));
	jdff dff_B_v7bfzJ8b8_0(.din(w_dff_B_FaRzaNcD9_0),.dout(w_dff_B_v7bfzJ8b8_0),.clk(gclk));
	jdff dff_B_ndlISqRV8_0(.din(w_dff_B_v7bfzJ8b8_0),.dout(w_dff_B_ndlISqRV8_0),.clk(gclk));
	jdff dff_B_wAapW3Cd0_0(.din(w_dff_B_ndlISqRV8_0),.dout(w_dff_B_wAapW3Cd0_0),.clk(gclk));
	jdff dff_B_2a2fGktN2_0(.din(w_dff_B_wAapW3Cd0_0),.dout(w_dff_B_2a2fGktN2_0),.clk(gclk));
	jdff dff_B_SUJAiTxQ9_0(.din(w_dff_B_2a2fGktN2_0),.dout(w_dff_B_SUJAiTxQ9_0),.clk(gclk));
	jdff dff_B_fvMxO81f6_0(.din(w_dff_B_SUJAiTxQ9_0),.dout(w_dff_B_fvMxO81f6_0),.clk(gclk));
	jdff dff_B_8XPyocbv2_0(.din(w_dff_B_fvMxO81f6_0),.dout(w_dff_B_8XPyocbv2_0),.clk(gclk));
	jdff dff_B_bnveSGRw9_0(.din(w_dff_B_8XPyocbv2_0),.dout(w_dff_B_bnveSGRw9_0),.clk(gclk));
	jdff dff_B_FmRSMsMy7_0(.din(w_dff_B_bnveSGRw9_0),.dout(w_dff_B_FmRSMsMy7_0),.clk(gclk));
	jdff dff_B_ZkNNlGdm5_0(.din(w_dff_B_FmRSMsMy7_0),.dout(w_dff_B_ZkNNlGdm5_0),.clk(gclk));
	jdff dff_B_vv73V3B65_0(.din(w_dff_B_ZkNNlGdm5_0),.dout(w_dff_B_vv73V3B65_0),.clk(gclk));
	jdff dff_B_go8YdW1i5_0(.din(w_dff_B_vv73V3B65_0),.dout(w_dff_B_go8YdW1i5_0),.clk(gclk));
	jdff dff_B_blbbGZV41_0(.din(w_dff_B_go8YdW1i5_0),.dout(w_dff_B_blbbGZV41_0),.clk(gclk));
	jdff dff_B_0b0N0YCK5_0(.din(w_dff_B_blbbGZV41_0),.dout(w_dff_B_0b0N0YCK5_0),.clk(gclk));
	jdff dff_B_kQMGscL80_0(.din(w_dff_B_0b0N0YCK5_0),.dout(w_dff_B_kQMGscL80_0),.clk(gclk));
	jdff dff_B_xXGtxy0E0_0(.din(w_dff_B_kQMGscL80_0),.dout(w_dff_B_xXGtxy0E0_0),.clk(gclk));
	jdff dff_B_sSzFJBc48_0(.din(w_dff_B_xXGtxy0E0_0),.dout(w_dff_B_sSzFJBc48_0),.clk(gclk));
	jdff dff_B_L0Gow7Jz5_0(.din(w_dff_B_sSzFJBc48_0),.dout(w_dff_B_L0Gow7Jz5_0),.clk(gclk));
	jdff dff_B_OSMMiefa9_0(.din(w_dff_B_L0Gow7Jz5_0),.dout(w_dff_B_OSMMiefa9_0),.clk(gclk));
	jdff dff_B_7v4lYdnc4_0(.din(w_dff_B_OSMMiefa9_0),.dout(w_dff_B_7v4lYdnc4_0),.clk(gclk));
	jdff dff_B_XfwMWNn70_0(.din(w_dff_B_7v4lYdnc4_0),.dout(w_dff_B_XfwMWNn70_0),.clk(gclk));
	jdff dff_B_wkxq2Bkn0_0(.din(w_dff_B_XfwMWNn70_0),.dout(w_dff_B_wkxq2Bkn0_0),.clk(gclk));
	jdff dff_B_59cngZlb0_0(.din(w_dff_B_wkxq2Bkn0_0),.dout(w_dff_B_59cngZlb0_0),.clk(gclk));
	jdff dff_B_UHQtzWZl8_0(.din(w_dff_B_59cngZlb0_0),.dout(w_dff_B_UHQtzWZl8_0),.clk(gclk));
	jdff dff_B_vgJcCKrd6_0(.din(w_dff_B_UHQtzWZl8_0),.dout(w_dff_B_vgJcCKrd6_0),.clk(gclk));
	jdff dff_B_e0HN5Sku6_0(.din(w_dff_B_vgJcCKrd6_0),.dout(w_dff_B_e0HN5Sku6_0),.clk(gclk));
	jdff dff_B_xoZojuwa7_0(.din(w_dff_B_e0HN5Sku6_0),.dout(w_dff_B_xoZojuwa7_0),.clk(gclk));
	jdff dff_B_PG2MTWyb5_0(.din(w_dff_B_xoZojuwa7_0),.dout(w_dff_B_PG2MTWyb5_0),.clk(gclk));
	jdff dff_B_VHn9TJQs4_1(.din(n1086),.dout(w_dff_B_VHn9TJQs4_1),.clk(gclk));
	jdff dff_B_weU0RXLM5_1(.din(w_dff_B_VHn9TJQs4_1),.dout(w_dff_B_weU0RXLM5_1),.clk(gclk));
	jdff dff_B_mXLpm9LL5_1(.din(w_dff_B_weU0RXLM5_1),.dout(w_dff_B_mXLpm9LL5_1),.clk(gclk));
	jdff dff_B_QQvrlayg6_1(.din(w_dff_B_mXLpm9LL5_1),.dout(w_dff_B_QQvrlayg6_1),.clk(gclk));
	jdff dff_B_7yNumaUC6_1(.din(w_dff_B_QQvrlayg6_1),.dout(w_dff_B_7yNumaUC6_1),.clk(gclk));
	jdff dff_B_g2vZiXYP5_1(.din(w_dff_B_7yNumaUC6_1),.dout(w_dff_B_g2vZiXYP5_1),.clk(gclk));
	jdff dff_B_8FnJnD3z7_1(.din(w_dff_B_g2vZiXYP5_1),.dout(w_dff_B_8FnJnD3z7_1),.clk(gclk));
	jdff dff_B_8d4CFpGF3_1(.din(w_dff_B_8FnJnD3z7_1),.dout(w_dff_B_8d4CFpGF3_1),.clk(gclk));
	jdff dff_B_FZaX2W3d6_1(.din(w_dff_B_8d4CFpGF3_1),.dout(w_dff_B_FZaX2W3d6_1),.clk(gclk));
	jdff dff_B_Ba1mraEJ8_1(.din(w_dff_B_FZaX2W3d6_1),.dout(w_dff_B_Ba1mraEJ8_1),.clk(gclk));
	jdff dff_B_CvJGr1j23_1(.din(w_dff_B_Ba1mraEJ8_1),.dout(w_dff_B_CvJGr1j23_1),.clk(gclk));
	jdff dff_B_VrLSQstI7_1(.din(w_dff_B_CvJGr1j23_1),.dout(w_dff_B_VrLSQstI7_1),.clk(gclk));
	jdff dff_B_yp0kKRyi6_1(.din(w_dff_B_VrLSQstI7_1),.dout(w_dff_B_yp0kKRyi6_1),.clk(gclk));
	jdff dff_B_alNwLkmM0_1(.din(w_dff_B_yp0kKRyi6_1),.dout(w_dff_B_alNwLkmM0_1),.clk(gclk));
	jdff dff_B_M1rMyHoL3_1(.din(w_dff_B_alNwLkmM0_1),.dout(w_dff_B_M1rMyHoL3_1),.clk(gclk));
	jdff dff_B_T6NVnOqK7_1(.din(w_dff_B_M1rMyHoL3_1),.dout(w_dff_B_T6NVnOqK7_1),.clk(gclk));
	jdff dff_B_TKF9hkmS6_1(.din(w_dff_B_T6NVnOqK7_1),.dout(w_dff_B_TKF9hkmS6_1),.clk(gclk));
	jdff dff_B_DfttxFvS3_1(.din(w_dff_B_TKF9hkmS6_1),.dout(w_dff_B_DfttxFvS3_1),.clk(gclk));
	jdff dff_B_hz3xGkkH4_1(.din(w_dff_B_DfttxFvS3_1),.dout(w_dff_B_hz3xGkkH4_1),.clk(gclk));
	jdff dff_B_mlrtrj4I8_1(.din(w_dff_B_hz3xGkkH4_1),.dout(w_dff_B_mlrtrj4I8_1),.clk(gclk));
	jdff dff_B_Z9uRKsnt5_1(.din(w_dff_B_mlrtrj4I8_1),.dout(w_dff_B_Z9uRKsnt5_1),.clk(gclk));
	jdff dff_B_tbdN8ecb3_1(.din(w_dff_B_Z9uRKsnt5_1),.dout(w_dff_B_tbdN8ecb3_1),.clk(gclk));
	jdff dff_B_8vwSmKNJ9_1(.din(w_dff_B_tbdN8ecb3_1),.dout(w_dff_B_8vwSmKNJ9_1),.clk(gclk));
	jdff dff_B_IioFGClq1_1(.din(w_dff_B_8vwSmKNJ9_1),.dout(w_dff_B_IioFGClq1_1),.clk(gclk));
	jdff dff_B_P91aLeGR0_1(.din(w_dff_B_IioFGClq1_1),.dout(w_dff_B_P91aLeGR0_1),.clk(gclk));
	jdff dff_B_72K5SKWg9_1(.din(w_dff_B_P91aLeGR0_1),.dout(w_dff_B_72K5SKWg9_1),.clk(gclk));
	jdff dff_B_gMB6IRLs1_1(.din(w_dff_B_72K5SKWg9_1),.dout(w_dff_B_gMB6IRLs1_1),.clk(gclk));
	jdff dff_B_Z6f4XFcB3_1(.din(w_dff_B_gMB6IRLs1_1),.dout(w_dff_B_Z6f4XFcB3_1),.clk(gclk));
	jdff dff_B_hfhOpRUK7_1(.din(w_dff_B_Z6f4XFcB3_1),.dout(w_dff_B_hfhOpRUK7_1),.clk(gclk));
	jdff dff_B_xOxumTwj5_1(.din(w_dff_B_hfhOpRUK7_1),.dout(w_dff_B_xOxumTwj5_1),.clk(gclk));
	jdff dff_B_0GcyFVx43_1(.din(w_dff_B_xOxumTwj5_1),.dout(w_dff_B_0GcyFVx43_1),.clk(gclk));
	jdff dff_B_uzSnaecV0_1(.din(w_dff_B_0GcyFVx43_1),.dout(w_dff_B_uzSnaecV0_1),.clk(gclk));
	jdff dff_B_WSTVPVVF3_1(.din(w_dff_B_uzSnaecV0_1),.dout(w_dff_B_WSTVPVVF3_1),.clk(gclk));
	jdff dff_B_QVr6NXvU1_1(.din(w_dff_B_WSTVPVVF3_1),.dout(w_dff_B_QVr6NXvU1_1),.clk(gclk));
	jdff dff_B_2X7izOS41_1(.din(w_dff_B_QVr6NXvU1_1),.dout(w_dff_B_2X7izOS41_1),.clk(gclk));
	jdff dff_B_rkbMdsOO8_1(.din(w_dff_B_2X7izOS41_1),.dout(w_dff_B_rkbMdsOO8_1),.clk(gclk));
	jdff dff_B_yph8wovY1_1(.din(w_dff_B_rkbMdsOO8_1),.dout(w_dff_B_yph8wovY1_1),.clk(gclk));
	jdff dff_B_tzqPMpLH0_1(.din(w_dff_B_yph8wovY1_1),.dout(w_dff_B_tzqPMpLH0_1),.clk(gclk));
	jdff dff_B_4iMasuAT4_1(.din(w_dff_B_tzqPMpLH0_1),.dout(w_dff_B_4iMasuAT4_1),.clk(gclk));
	jdff dff_B_7BewOAbz1_1(.din(w_dff_B_4iMasuAT4_1),.dout(w_dff_B_7BewOAbz1_1),.clk(gclk));
	jdff dff_B_0wCuhX9P9_1(.din(w_dff_B_7BewOAbz1_1),.dout(w_dff_B_0wCuhX9P9_1),.clk(gclk));
	jdff dff_B_HxRmiiOV9_1(.din(w_dff_B_0wCuhX9P9_1),.dout(w_dff_B_HxRmiiOV9_1),.clk(gclk));
	jdff dff_B_Legzqtl65_1(.din(w_dff_B_HxRmiiOV9_1),.dout(w_dff_B_Legzqtl65_1),.clk(gclk));
	jdff dff_B_9i2TSU313_1(.din(w_dff_B_Legzqtl65_1),.dout(w_dff_B_9i2TSU313_1),.clk(gclk));
	jdff dff_B_ORN53I3K0_1(.din(w_dff_B_9i2TSU313_1),.dout(w_dff_B_ORN53I3K0_1),.clk(gclk));
	jdff dff_B_8DFnl29K3_1(.din(w_dff_B_ORN53I3K0_1),.dout(w_dff_B_8DFnl29K3_1),.clk(gclk));
	jdff dff_B_eQXs7xZY4_1(.din(w_dff_B_8DFnl29K3_1),.dout(w_dff_B_eQXs7xZY4_1),.clk(gclk));
	jdff dff_B_QWKKtUMY4_1(.din(w_dff_B_eQXs7xZY4_1),.dout(w_dff_B_QWKKtUMY4_1),.clk(gclk));
	jdff dff_B_Pu7APPQZ1_1(.din(w_dff_B_QWKKtUMY4_1),.dout(w_dff_B_Pu7APPQZ1_1),.clk(gclk));
	jdff dff_B_pUrO5l0j5_1(.din(w_dff_B_Pu7APPQZ1_1),.dout(w_dff_B_pUrO5l0j5_1),.clk(gclk));
	jdff dff_B_zAqgsTp33_1(.din(w_dff_B_pUrO5l0j5_1),.dout(w_dff_B_zAqgsTp33_1),.clk(gclk));
	jdff dff_B_NeOthQYI5_1(.din(w_dff_B_zAqgsTp33_1),.dout(w_dff_B_NeOthQYI5_1),.clk(gclk));
	jdff dff_B_OFPMgZrs6_1(.din(w_dff_B_NeOthQYI5_1),.dout(w_dff_B_OFPMgZrs6_1),.clk(gclk));
	jdff dff_B_5qdPJeJF5_1(.din(w_dff_B_OFPMgZrs6_1),.dout(w_dff_B_5qdPJeJF5_1),.clk(gclk));
	jdff dff_B_9YZ0tzTb7_1(.din(w_dff_B_5qdPJeJF5_1),.dout(w_dff_B_9YZ0tzTb7_1),.clk(gclk));
	jdff dff_B_dxokdYOo3_1(.din(w_dff_B_9YZ0tzTb7_1),.dout(w_dff_B_dxokdYOo3_1),.clk(gclk));
	jdff dff_B_BAh8xJSH5_1(.din(w_dff_B_dxokdYOo3_1),.dout(w_dff_B_BAh8xJSH5_1),.clk(gclk));
	jdff dff_B_wUKF8ogW1_1(.din(w_dff_B_BAh8xJSH5_1),.dout(w_dff_B_wUKF8ogW1_1),.clk(gclk));
	jdff dff_B_3cFsxSls8_1(.din(w_dff_B_wUKF8ogW1_1),.dout(w_dff_B_3cFsxSls8_1),.clk(gclk));
	jdff dff_B_MJ8qJrJc7_1(.din(w_dff_B_3cFsxSls8_1),.dout(w_dff_B_MJ8qJrJc7_1),.clk(gclk));
	jdff dff_B_YJ9BY6258_1(.din(w_dff_B_MJ8qJrJc7_1),.dout(w_dff_B_YJ9BY6258_1),.clk(gclk));
	jdff dff_B_IbaBSp9K6_1(.din(w_dff_B_YJ9BY6258_1),.dout(w_dff_B_IbaBSp9K6_1),.clk(gclk));
	jdff dff_B_gphZL0c48_1(.din(w_dff_B_IbaBSp9K6_1),.dout(w_dff_B_gphZL0c48_1),.clk(gclk));
	jdff dff_B_zjBEs5kK9_1(.din(w_dff_B_gphZL0c48_1),.dout(w_dff_B_zjBEs5kK9_1),.clk(gclk));
	jdff dff_B_RCtKRZoy9_1(.din(w_dff_B_zjBEs5kK9_1),.dout(w_dff_B_RCtKRZoy9_1),.clk(gclk));
	jdff dff_B_CWTtPHLv0_1(.din(w_dff_B_RCtKRZoy9_1),.dout(w_dff_B_CWTtPHLv0_1),.clk(gclk));
	jdff dff_B_9vygHb7i0_1(.din(w_dff_B_CWTtPHLv0_1),.dout(w_dff_B_9vygHb7i0_1),.clk(gclk));
	jdff dff_B_zrbP7GxY7_1(.din(w_dff_B_9vygHb7i0_1),.dout(w_dff_B_zrbP7GxY7_1),.clk(gclk));
	jdff dff_B_vlgOJ9V45_1(.din(w_dff_B_zrbP7GxY7_1),.dout(w_dff_B_vlgOJ9V45_1),.clk(gclk));
	jdff dff_B_lQdenUxA3_1(.din(w_dff_B_vlgOJ9V45_1),.dout(w_dff_B_lQdenUxA3_1),.clk(gclk));
	jdff dff_B_T9S4j88q1_1(.din(w_dff_B_lQdenUxA3_1),.dout(w_dff_B_T9S4j88q1_1),.clk(gclk));
	jdff dff_B_YMHPHOGC7_1(.din(w_dff_B_T9S4j88q1_1),.dout(w_dff_B_YMHPHOGC7_1),.clk(gclk));
	jdff dff_B_e3vPg3aK4_1(.din(w_dff_B_YMHPHOGC7_1),.dout(w_dff_B_e3vPg3aK4_1),.clk(gclk));
	jdff dff_B_3haVZqPq3_1(.din(w_dff_B_e3vPg3aK4_1),.dout(w_dff_B_3haVZqPq3_1),.clk(gclk));
	jdff dff_B_XWeteEXP6_1(.din(w_dff_B_3haVZqPq3_1),.dout(w_dff_B_XWeteEXP6_1),.clk(gclk));
	jdff dff_B_smQYrNTu9_1(.din(w_dff_B_XWeteEXP6_1),.dout(w_dff_B_smQYrNTu9_1),.clk(gclk));
	jdff dff_B_ubSYQkAp4_1(.din(w_dff_B_smQYrNTu9_1),.dout(w_dff_B_ubSYQkAp4_1),.clk(gclk));
	jdff dff_B_S1mvOlBs1_1(.din(w_dff_B_ubSYQkAp4_1),.dout(w_dff_B_S1mvOlBs1_1),.clk(gclk));
	jdff dff_B_sVsR5Bib1_1(.din(w_dff_B_S1mvOlBs1_1),.dout(w_dff_B_sVsR5Bib1_1),.clk(gclk));
	jdff dff_B_THBBGuER1_1(.din(w_dff_B_sVsR5Bib1_1),.dout(w_dff_B_THBBGuER1_1),.clk(gclk));
	jdff dff_B_Fvn1pcjV7_1(.din(w_dff_B_THBBGuER1_1),.dout(w_dff_B_Fvn1pcjV7_1),.clk(gclk));
	jdff dff_B_6kjFu5kD2_1(.din(w_dff_B_Fvn1pcjV7_1),.dout(w_dff_B_6kjFu5kD2_1),.clk(gclk));
	jdff dff_B_QQqIqfzG1_1(.din(w_dff_B_6kjFu5kD2_1),.dout(w_dff_B_QQqIqfzG1_1),.clk(gclk));
	jdff dff_B_JUYeebX73_1(.din(w_dff_B_QQqIqfzG1_1),.dout(w_dff_B_JUYeebX73_1),.clk(gclk));
	jdff dff_B_ZcZAQ4h83_1(.din(w_dff_B_JUYeebX73_1),.dout(w_dff_B_ZcZAQ4h83_1),.clk(gclk));
	jdff dff_B_KasNIBlK6_1(.din(w_dff_B_ZcZAQ4h83_1),.dout(w_dff_B_KasNIBlK6_1),.clk(gclk));
	jdff dff_B_PxF00urH7_1(.din(w_dff_B_KasNIBlK6_1),.dout(w_dff_B_PxF00urH7_1),.clk(gclk));
	jdff dff_B_AhfhLbtx1_1(.din(w_dff_B_PxF00urH7_1),.dout(w_dff_B_AhfhLbtx1_1),.clk(gclk));
	jdff dff_B_6jqm9QDu1_1(.din(w_dff_B_AhfhLbtx1_1),.dout(w_dff_B_6jqm9QDu1_1),.clk(gclk));
	jdff dff_B_RAzeX9Ee3_1(.din(w_dff_B_6jqm9QDu1_1),.dout(w_dff_B_RAzeX9Ee3_1),.clk(gclk));
	jdff dff_B_h5ZmYzif9_1(.din(w_dff_B_RAzeX9Ee3_1),.dout(w_dff_B_h5ZmYzif9_1),.clk(gclk));
	jdff dff_B_Gq98wQqv7_1(.din(w_dff_B_h5ZmYzif9_1),.dout(w_dff_B_Gq98wQqv7_1),.clk(gclk));
	jdff dff_B_LJPx6NS17_1(.din(w_dff_B_Gq98wQqv7_1),.dout(w_dff_B_LJPx6NS17_1),.clk(gclk));
	jdff dff_B_4wHqYd5m9_1(.din(w_dff_B_LJPx6NS17_1),.dout(w_dff_B_4wHqYd5m9_1),.clk(gclk));
	jdff dff_B_TzECuIlT0_1(.din(w_dff_B_4wHqYd5m9_1),.dout(w_dff_B_TzECuIlT0_1),.clk(gclk));
	jdff dff_B_CYelCk5L1_1(.din(w_dff_B_TzECuIlT0_1),.dout(w_dff_B_CYelCk5L1_1),.clk(gclk));
	jdff dff_B_MJQcLT6M0_1(.din(w_dff_B_CYelCk5L1_1),.dout(w_dff_B_MJQcLT6M0_1),.clk(gclk));
	jdff dff_B_ES7KtxQN2_1(.din(w_dff_B_MJQcLT6M0_1),.dout(w_dff_B_ES7KtxQN2_1),.clk(gclk));
	jdff dff_B_BqWfWFbi0_1(.din(w_dff_B_ES7KtxQN2_1),.dout(w_dff_B_BqWfWFbi0_1),.clk(gclk));
	jdff dff_B_07dyed016_1(.din(w_dff_B_BqWfWFbi0_1),.dout(w_dff_B_07dyed016_1),.clk(gclk));
	jdff dff_B_F5vh5ikl9_1(.din(w_dff_B_07dyed016_1),.dout(w_dff_B_F5vh5ikl9_1),.clk(gclk));
	jdff dff_B_pqau9lx39_1(.din(w_dff_B_F5vh5ikl9_1),.dout(w_dff_B_pqau9lx39_1),.clk(gclk));
	jdff dff_B_71rkZhAP6_1(.din(w_dff_B_pqau9lx39_1),.dout(w_dff_B_71rkZhAP6_1),.clk(gclk));
	jdff dff_B_GhOmgY1E2_1(.din(w_dff_B_71rkZhAP6_1),.dout(w_dff_B_GhOmgY1E2_1),.clk(gclk));
	jdff dff_B_suawknRD1_1(.din(w_dff_B_GhOmgY1E2_1),.dout(w_dff_B_suawknRD1_1),.clk(gclk));
	jdff dff_B_J6ckBTzW4_1(.din(w_dff_B_suawknRD1_1),.dout(w_dff_B_J6ckBTzW4_1),.clk(gclk));
	jdff dff_B_GWvrKgw21_1(.din(w_dff_B_J6ckBTzW4_1),.dout(w_dff_B_GWvrKgw21_1),.clk(gclk));
	jdff dff_B_20TtFKlF8_1(.din(w_dff_B_GWvrKgw21_1),.dout(w_dff_B_20TtFKlF8_1),.clk(gclk));
	jdff dff_B_dguU4IQa4_1(.din(w_dff_B_20TtFKlF8_1),.dout(w_dff_B_dguU4IQa4_1),.clk(gclk));
	jdff dff_B_0Xx7iimN3_1(.din(w_dff_B_dguU4IQa4_1),.dout(w_dff_B_0Xx7iimN3_1),.clk(gclk));
	jdff dff_B_UiQkJDS42_1(.din(w_dff_B_0Xx7iimN3_1),.dout(w_dff_B_UiQkJDS42_1),.clk(gclk));
	jdff dff_B_KQYMATR73_1(.din(w_dff_B_UiQkJDS42_1),.dout(w_dff_B_KQYMATR73_1),.clk(gclk));
	jdff dff_B_Tm6JEVns6_1(.din(w_dff_B_KQYMATR73_1),.dout(w_dff_B_Tm6JEVns6_1),.clk(gclk));
	jdff dff_B_QmP3Pabd6_1(.din(w_dff_B_Tm6JEVns6_1),.dout(w_dff_B_QmP3Pabd6_1),.clk(gclk));
	jdff dff_B_I3kkLVVQ0_1(.din(w_dff_B_QmP3Pabd6_1),.dout(w_dff_B_I3kkLVVQ0_1),.clk(gclk));
	jdff dff_B_rs3vVlKB5_1(.din(w_dff_B_I3kkLVVQ0_1),.dout(w_dff_B_rs3vVlKB5_1),.clk(gclk));
	jdff dff_B_Pe1iiYr60_1(.din(w_dff_B_rs3vVlKB5_1),.dout(w_dff_B_Pe1iiYr60_1),.clk(gclk));
	jdff dff_B_M7EI9SW90_0(.din(n1087),.dout(w_dff_B_M7EI9SW90_0),.clk(gclk));
	jdff dff_B_5DlrnuB45_0(.din(w_dff_B_M7EI9SW90_0),.dout(w_dff_B_5DlrnuB45_0),.clk(gclk));
	jdff dff_B_4NvbCU4G1_0(.din(w_dff_B_5DlrnuB45_0),.dout(w_dff_B_4NvbCU4G1_0),.clk(gclk));
	jdff dff_B_ifBdqo8a5_0(.din(w_dff_B_4NvbCU4G1_0),.dout(w_dff_B_ifBdqo8a5_0),.clk(gclk));
	jdff dff_B_oAaGdQqR9_0(.din(w_dff_B_ifBdqo8a5_0),.dout(w_dff_B_oAaGdQqR9_0),.clk(gclk));
	jdff dff_B_IeYAlWuO9_0(.din(w_dff_B_oAaGdQqR9_0),.dout(w_dff_B_IeYAlWuO9_0),.clk(gclk));
	jdff dff_B_JqH1fp9I9_0(.din(w_dff_B_IeYAlWuO9_0),.dout(w_dff_B_JqH1fp9I9_0),.clk(gclk));
	jdff dff_B_P673onFb5_0(.din(w_dff_B_JqH1fp9I9_0),.dout(w_dff_B_P673onFb5_0),.clk(gclk));
	jdff dff_B_AgSz4TSZ3_0(.din(w_dff_B_P673onFb5_0),.dout(w_dff_B_AgSz4TSZ3_0),.clk(gclk));
	jdff dff_B_OZ0h0jjA9_0(.din(w_dff_B_AgSz4TSZ3_0),.dout(w_dff_B_OZ0h0jjA9_0),.clk(gclk));
	jdff dff_B_xxaRuZgU2_0(.din(w_dff_B_OZ0h0jjA9_0),.dout(w_dff_B_xxaRuZgU2_0),.clk(gclk));
	jdff dff_B_bPA1eVCN6_0(.din(w_dff_B_xxaRuZgU2_0),.dout(w_dff_B_bPA1eVCN6_0),.clk(gclk));
	jdff dff_B_QiiZuJe62_0(.din(w_dff_B_bPA1eVCN6_0),.dout(w_dff_B_QiiZuJe62_0),.clk(gclk));
	jdff dff_B_rSHWIbpy0_0(.din(w_dff_B_QiiZuJe62_0),.dout(w_dff_B_rSHWIbpy0_0),.clk(gclk));
	jdff dff_B_5nrxxgvh5_0(.din(w_dff_B_rSHWIbpy0_0),.dout(w_dff_B_5nrxxgvh5_0),.clk(gclk));
	jdff dff_B_ytaZtXJp0_0(.din(w_dff_B_5nrxxgvh5_0),.dout(w_dff_B_ytaZtXJp0_0),.clk(gclk));
	jdff dff_B_5RqGnWwl9_0(.din(w_dff_B_ytaZtXJp0_0),.dout(w_dff_B_5RqGnWwl9_0),.clk(gclk));
	jdff dff_B_PYHhmXPH4_0(.din(w_dff_B_5RqGnWwl9_0),.dout(w_dff_B_PYHhmXPH4_0),.clk(gclk));
	jdff dff_B_4eOcVJVv8_0(.din(w_dff_B_PYHhmXPH4_0),.dout(w_dff_B_4eOcVJVv8_0),.clk(gclk));
	jdff dff_B_wSv5OMIn7_0(.din(w_dff_B_4eOcVJVv8_0),.dout(w_dff_B_wSv5OMIn7_0),.clk(gclk));
	jdff dff_B_rCGn6ZpC6_0(.din(w_dff_B_wSv5OMIn7_0),.dout(w_dff_B_rCGn6ZpC6_0),.clk(gclk));
	jdff dff_B_FDrzNFow4_0(.din(w_dff_B_rCGn6ZpC6_0),.dout(w_dff_B_FDrzNFow4_0),.clk(gclk));
	jdff dff_B_nM0r0Jkc4_0(.din(w_dff_B_FDrzNFow4_0),.dout(w_dff_B_nM0r0Jkc4_0),.clk(gclk));
	jdff dff_B_JZkn5b0e9_0(.din(w_dff_B_nM0r0Jkc4_0),.dout(w_dff_B_JZkn5b0e9_0),.clk(gclk));
	jdff dff_B_n0IIdDsi3_0(.din(w_dff_B_JZkn5b0e9_0),.dout(w_dff_B_n0IIdDsi3_0),.clk(gclk));
	jdff dff_B_JYv0oRdD6_0(.din(w_dff_B_n0IIdDsi3_0),.dout(w_dff_B_JYv0oRdD6_0),.clk(gclk));
	jdff dff_B_tMe3Qlhx6_0(.din(w_dff_B_JYv0oRdD6_0),.dout(w_dff_B_tMe3Qlhx6_0),.clk(gclk));
	jdff dff_B_YAvOovI92_0(.din(w_dff_B_tMe3Qlhx6_0),.dout(w_dff_B_YAvOovI92_0),.clk(gclk));
	jdff dff_B_mhDkDj2e1_0(.din(w_dff_B_YAvOovI92_0),.dout(w_dff_B_mhDkDj2e1_0),.clk(gclk));
	jdff dff_B_iPZzOWWJ1_0(.din(w_dff_B_mhDkDj2e1_0),.dout(w_dff_B_iPZzOWWJ1_0),.clk(gclk));
	jdff dff_B_oWM6jmUt7_0(.din(w_dff_B_iPZzOWWJ1_0),.dout(w_dff_B_oWM6jmUt7_0),.clk(gclk));
	jdff dff_B_cN3zvUzP9_0(.din(w_dff_B_oWM6jmUt7_0),.dout(w_dff_B_cN3zvUzP9_0),.clk(gclk));
	jdff dff_B_Jd1DXDNY2_0(.din(w_dff_B_cN3zvUzP9_0),.dout(w_dff_B_Jd1DXDNY2_0),.clk(gclk));
	jdff dff_B_ReW7hyrU9_0(.din(w_dff_B_Jd1DXDNY2_0),.dout(w_dff_B_ReW7hyrU9_0),.clk(gclk));
	jdff dff_B_kPvfq4EU7_0(.din(w_dff_B_ReW7hyrU9_0),.dout(w_dff_B_kPvfq4EU7_0),.clk(gclk));
	jdff dff_B_eNJRRZPe3_0(.din(w_dff_B_kPvfq4EU7_0),.dout(w_dff_B_eNJRRZPe3_0),.clk(gclk));
	jdff dff_B_0JaJ4R4P9_0(.din(w_dff_B_eNJRRZPe3_0),.dout(w_dff_B_0JaJ4R4P9_0),.clk(gclk));
	jdff dff_B_yQhDGsuU4_0(.din(w_dff_B_0JaJ4R4P9_0),.dout(w_dff_B_yQhDGsuU4_0),.clk(gclk));
	jdff dff_B_whvYdmgG3_0(.din(w_dff_B_yQhDGsuU4_0),.dout(w_dff_B_whvYdmgG3_0),.clk(gclk));
	jdff dff_B_sJQDvEHQ2_0(.din(w_dff_B_whvYdmgG3_0),.dout(w_dff_B_sJQDvEHQ2_0),.clk(gclk));
	jdff dff_B_hLcmAr003_0(.din(w_dff_B_sJQDvEHQ2_0),.dout(w_dff_B_hLcmAr003_0),.clk(gclk));
	jdff dff_B_N5ZZWG9P9_0(.din(w_dff_B_hLcmAr003_0),.dout(w_dff_B_N5ZZWG9P9_0),.clk(gclk));
	jdff dff_B_E9XpuREw2_0(.din(w_dff_B_N5ZZWG9P9_0),.dout(w_dff_B_E9XpuREw2_0),.clk(gclk));
	jdff dff_B_tHJtXSo34_0(.din(w_dff_B_E9XpuREw2_0),.dout(w_dff_B_tHJtXSo34_0),.clk(gclk));
	jdff dff_B_pvKd1m2w5_0(.din(w_dff_B_tHJtXSo34_0),.dout(w_dff_B_pvKd1m2w5_0),.clk(gclk));
	jdff dff_B_unjXOp8p0_0(.din(w_dff_B_pvKd1m2w5_0),.dout(w_dff_B_unjXOp8p0_0),.clk(gclk));
	jdff dff_B_ZI0RRKRl2_0(.din(w_dff_B_unjXOp8p0_0),.dout(w_dff_B_ZI0RRKRl2_0),.clk(gclk));
	jdff dff_B_CnP0slgD6_0(.din(w_dff_B_ZI0RRKRl2_0),.dout(w_dff_B_CnP0slgD6_0),.clk(gclk));
	jdff dff_B_Pu8KmmXN5_0(.din(w_dff_B_CnP0slgD6_0),.dout(w_dff_B_Pu8KmmXN5_0),.clk(gclk));
	jdff dff_B_IzNaHN1V0_0(.din(w_dff_B_Pu8KmmXN5_0),.dout(w_dff_B_IzNaHN1V0_0),.clk(gclk));
	jdff dff_B_8ejwgIiy8_0(.din(w_dff_B_IzNaHN1V0_0),.dout(w_dff_B_8ejwgIiy8_0),.clk(gclk));
	jdff dff_B_maSwbOzT1_0(.din(w_dff_B_8ejwgIiy8_0),.dout(w_dff_B_maSwbOzT1_0),.clk(gclk));
	jdff dff_B_HiyVQhUE9_0(.din(w_dff_B_maSwbOzT1_0),.dout(w_dff_B_HiyVQhUE9_0),.clk(gclk));
	jdff dff_B_OreHujBm1_0(.din(w_dff_B_HiyVQhUE9_0),.dout(w_dff_B_OreHujBm1_0),.clk(gclk));
	jdff dff_B_snYMKc227_0(.din(w_dff_B_OreHujBm1_0),.dout(w_dff_B_snYMKc227_0),.clk(gclk));
	jdff dff_B_hv0woxsA1_0(.din(w_dff_B_snYMKc227_0),.dout(w_dff_B_hv0woxsA1_0),.clk(gclk));
	jdff dff_B_mC0dDsO84_0(.din(w_dff_B_hv0woxsA1_0),.dout(w_dff_B_mC0dDsO84_0),.clk(gclk));
	jdff dff_B_gFIsGDk84_0(.din(w_dff_B_mC0dDsO84_0),.dout(w_dff_B_gFIsGDk84_0),.clk(gclk));
	jdff dff_B_A5aTERoy1_0(.din(w_dff_B_gFIsGDk84_0),.dout(w_dff_B_A5aTERoy1_0),.clk(gclk));
	jdff dff_B_2gLOA8Ld4_0(.din(w_dff_B_A5aTERoy1_0),.dout(w_dff_B_2gLOA8Ld4_0),.clk(gclk));
	jdff dff_B_IT5vkL4H7_0(.din(w_dff_B_2gLOA8Ld4_0),.dout(w_dff_B_IT5vkL4H7_0),.clk(gclk));
	jdff dff_B_qO9ITuGd6_0(.din(w_dff_B_IT5vkL4H7_0),.dout(w_dff_B_qO9ITuGd6_0),.clk(gclk));
	jdff dff_B_1nPCrTZm5_0(.din(w_dff_B_qO9ITuGd6_0),.dout(w_dff_B_1nPCrTZm5_0),.clk(gclk));
	jdff dff_B_6iS57Xmq5_0(.din(w_dff_B_1nPCrTZm5_0),.dout(w_dff_B_6iS57Xmq5_0),.clk(gclk));
	jdff dff_B_YHJplSgl9_0(.din(w_dff_B_6iS57Xmq5_0),.dout(w_dff_B_YHJplSgl9_0),.clk(gclk));
	jdff dff_B_12qGtThZ1_0(.din(w_dff_B_YHJplSgl9_0),.dout(w_dff_B_12qGtThZ1_0),.clk(gclk));
	jdff dff_B_NxXlxi6j0_0(.din(w_dff_B_12qGtThZ1_0),.dout(w_dff_B_NxXlxi6j0_0),.clk(gclk));
	jdff dff_B_iVAxyb5X0_0(.din(w_dff_B_NxXlxi6j0_0),.dout(w_dff_B_iVAxyb5X0_0),.clk(gclk));
	jdff dff_B_kZAyKJ1V6_0(.din(w_dff_B_iVAxyb5X0_0),.dout(w_dff_B_kZAyKJ1V6_0),.clk(gclk));
	jdff dff_B_CPMIU3Et0_0(.din(w_dff_B_kZAyKJ1V6_0),.dout(w_dff_B_CPMIU3Et0_0),.clk(gclk));
	jdff dff_B_yKLMkLdr5_0(.din(w_dff_B_CPMIU3Et0_0),.dout(w_dff_B_yKLMkLdr5_0),.clk(gclk));
	jdff dff_B_t9ulnEnL3_0(.din(w_dff_B_yKLMkLdr5_0),.dout(w_dff_B_t9ulnEnL3_0),.clk(gclk));
	jdff dff_B_ZYEy1BOh6_0(.din(w_dff_B_t9ulnEnL3_0),.dout(w_dff_B_ZYEy1BOh6_0),.clk(gclk));
	jdff dff_B_1eWsj6Xp4_0(.din(w_dff_B_ZYEy1BOh6_0),.dout(w_dff_B_1eWsj6Xp4_0),.clk(gclk));
	jdff dff_B_PNx1tVtz4_0(.din(w_dff_B_1eWsj6Xp4_0),.dout(w_dff_B_PNx1tVtz4_0),.clk(gclk));
	jdff dff_B_25zsk5Pn9_0(.din(w_dff_B_PNx1tVtz4_0),.dout(w_dff_B_25zsk5Pn9_0),.clk(gclk));
	jdff dff_B_Kqqn8YoK4_0(.din(w_dff_B_25zsk5Pn9_0),.dout(w_dff_B_Kqqn8YoK4_0),.clk(gclk));
	jdff dff_B_H6KRydry6_0(.din(w_dff_B_Kqqn8YoK4_0),.dout(w_dff_B_H6KRydry6_0),.clk(gclk));
	jdff dff_B_Zbe0OBqx2_0(.din(w_dff_B_H6KRydry6_0),.dout(w_dff_B_Zbe0OBqx2_0),.clk(gclk));
	jdff dff_B_h6ThyQlb0_0(.din(w_dff_B_Zbe0OBqx2_0),.dout(w_dff_B_h6ThyQlb0_0),.clk(gclk));
	jdff dff_B_LDP8luwg1_0(.din(w_dff_B_h6ThyQlb0_0),.dout(w_dff_B_LDP8luwg1_0),.clk(gclk));
	jdff dff_B_Rfes5znt0_0(.din(w_dff_B_LDP8luwg1_0),.dout(w_dff_B_Rfes5znt0_0),.clk(gclk));
	jdff dff_B_h0BAPlbY7_0(.din(w_dff_B_Rfes5znt0_0),.dout(w_dff_B_h0BAPlbY7_0),.clk(gclk));
	jdff dff_B_2pwfBrSc6_0(.din(w_dff_B_h0BAPlbY7_0),.dout(w_dff_B_2pwfBrSc6_0),.clk(gclk));
	jdff dff_B_zIGcAts16_0(.din(w_dff_B_2pwfBrSc6_0),.dout(w_dff_B_zIGcAts16_0),.clk(gclk));
	jdff dff_B_WwPZX7ES5_0(.din(w_dff_B_zIGcAts16_0),.dout(w_dff_B_WwPZX7ES5_0),.clk(gclk));
	jdff dff_B_v3N7St3I6_0(.din(w_dff_B_WwPZX7ES5_0),.dout(w_dff_B_v3N7St3I6_0),.clk(gclk));
	jdff dff_B_lpQCQZH77_0(.din(w_dff_B_v3N7St3I6_0),.dout(w_dff_B_lpQCQZH77_0),.clk(gclk));
	jdff dff_B_Zoxst3704_0(.din(w_dff_B_lpQCQZH77_0),.dout(w_dff_B_Zoxst3704_0),.clk(gclk));
	jdff dff_B_T8aQEHVr2_0(.din(w_dff_B_Zoxst3704_0),.dout(w_dff_B_T8aQEHVr2_0),.clk(gclk));
	jdff dff_B_qxcsQPKH3_0(.din(w_dff_B_T8aQEHVr2_0),.dout(w_dff_B_qxcsQPKH3_0),.clk(gclk));
	jdff dff_B_WFv9DYoH8_0(.din(w_dff_B_qxcsQPKH3_0),.dout(w_dff_B_WFv9DYoH8_0),.clk(gclk));
	jdff dff_B_tWf3XB4i8_0(.din(w_dff_B_WFv9DYoH8_0),.dout(w_dff_B_tWf3XB4i8_0),.clk(gclk));
	jdff dff_B_iJS4LuBa1_0(.din(w_dff_B_tWf3XB4i8_0),.dout(w_dff_B_iJS4LuBa1_0),.clk(gclk));
	jdff dff_B_P2oTfjLT0_0(.din(w_dff_B_iJS4LuBa1_0),.dout(w_dff_B_P2oTfjLT0_0),.clk(gclk));
	jdff dff_B_V9TZ42Uf4_0(.din(w_dff_B_P2oTfjLT0_0),.dout(w_dff_B_V9TZ42Uf4_0),.clk(gclk));
	jdff dff_B_JKBWP2Ai8_0(.din(w_dff_B_V9TZ42Uf4_0),.dout(w_dff_B_JKBWP2Ai8_0),.clk(gclk));
	jdff dff_B_UjaNzp175_0(.din(w_dff_B_JKBWP2Ai8_0),.dout(w_dff_B_UjaNzp175_0),.clk(gclk));
	jdff dff_B_m9DS1XgK6_0(.din(w_dff_B_UjaNzp175_0),.dout(w_dff_B_m9DS1XgK6_0),.clk(gclk));
	jdff dff_B_CaNEwa7s6_0(.din(w_dff_B_m9DS1XgK6_0),.dout(w_dff_B_CaNEwa7s6_0),.clk(gclk));
	jdff dff_B_huh2ku8H8_0(.din(w_dff_B_CaNEwa7s6_0),.dout(w_dff_B_huh2ku8H8_0),.clk(gclk));
	jdff dff_B_Z6mUNCq97_0(.din(w_dff_B_huh2ku8H8_0),.dout(w_dff_B_Z6mUNCq97_0),.clk(gclk));
	jdff dff_B_znD4ty7R5_0(.din(w_dff_B_Z6mUNCq97_0),.dout(w_dff_B_znD4ty7R5_0),.clk(gclk));
	jdff dff_B_TnCyVnkM8_0(.din(w_dff_B_znD4ty7R5_0),.dout(w_dff_B_TnCyVnkM8_0),.clk(gclk));
	jdff dff_B_kNPdqaCW7_0(.din(w_dff_B_TnCyVnkM8_0),.dout(w_dff_B_kNPdqaCW7_0),.clk(gclk));
	jdff dff_B_nRrdxhvB4_0(.din(w_dff_B_kNPdqaCW7_0),.dout(w_dff_B_nRrdxhvB4_0),.clk(gclk));
	jdff dff_B_u4rFfE759_0(.din(w_dff_B_nRrdxhvB4_0),.dout(w_dff_B_u4rFfE759_0),.clk(gclk));
	jdff dff_B_jRJlZfOd8_0(.din(w_dff_B_u4rFfE759_0),.dout(w_dff_B_jRJlZfOd8_0),.clk(gclk));
	jdff dff_B_7SiybSqA8_0(.din(w_dff_B_jRJlZfOd8_0),.dout(w_dff_B_7SiybSqA8_0),.clk(gclk));
	jdff dff_B_0oAT4Rev5_0(.din(w_dff_B_7SiybSqA8_0),.dout(w_dff_B_0oAT4Rev5_0),.clk(gclk));
	jdff dff_B_s2gsltDL7_0(.din(w_dff_B_0oAT4Rev5_0),.dout(w_dff_B_s2gsltDL7_0),.clk(gclk));
	jdff dff_B_Va5VyfBr5_0(.din(w_dff_B_s2gsltDL7_0),.dout(w_dff_B_Va5VyfBr5_0),.clk(gclk));
	jdff dff_B_YEIBzdqU3_0(.din(w_dff_B_Va5VyfBr5_0),.dout(w_dff_B_YEIBzdqU3_0),.clk(gclk));
	jdff dff_B_1330L5tP0_0(.din(w_dff_B_YEIBzdqU3_0),.dout(w_dff_B_1330L5tP0_0),.clk(gclk));
	jdff dff_B_7DRwlRO77_0(.din(w_dff_B_1330L5tP0_0),.dout(w_dff_B_7DRwlRO77_0),.clk(gclk));
	jdff dff_B_kLMAFHjd5_0(.din(w_dff_B_7DRwlRO77_0),.dout(w_dff_B_kLMAFHjd5_0),.clk(gclk));
	jdff dff_B_YHtR4fi00_0(.din(w_dff_B_kLMAFHjd5_0),.dout(w_dff_B_YHtR4fi00_0),.clk(gclk));
	jdff dff_B_Mva6TcQC3_1(.din(n1080),.dout(w_dff_B_Mva6TcQC3_1),.clk(gclk));
	jdff dff_B_kokxEdVW1_1(.din(w_dff_B_Mva6TcQC3_1),.dout(w_dff_B_kokxEdVW1_1),.clk(gclk));
	jdff dff_B_DuHvCeXp9_1(.din(w_dff_B_kokxEdVW1_1),.dout(w_dff_B_DuHvCeXp9_1),.clk(gclk));
	jdff dff_B_8HTLUvlt4_1(.din(w_dff_B_DuHvCeXp9_1),.dout(w_dff_B_8HTLUvlt4_1),.clk(gclk));
	jdff dff_B_IVq4IGff9_1(.din(w_dff_B_8HTLUvlt4_1),.dout(w_dff_B_IVq4IGff9_1),.clk(gclk));
	jdff dff_B_X4mKLp5N4_1(.din(w_dff_B_IVq4IGff9_1),.dout(w_dff_B_X4mKLp5N4_1),.clk(gclk));
	jdff dff_B_KmwrLEB03_1(.din(w_dff_B_X4mKLp5N4_1),.dout(w_dff_B_KmwrLEB03_1),.clk(gclk));
	jdff dff_B_0esGfP8z2_1(.din(w_dff_B_KmwrLEB03_1),.dout(w_dff_B_0esGfP8z2_1),.clk(gclk));
	jdff dff_B_f7vGlDzW6_1(.din(w_dff_B_0esGfP8z2_1),.dout(w_dff_B_f7vGlDzW6_1),.clk(gclk));
	jdff dff_B_DasWWJJw4_1(.din(w_dff_B_f7vGlDzW6_1),.dout(w_dff_B_DasWWJJw4_1),.clk(gclk));
	jdff dff_B_mWMed6LW1_1(.din(w_dff_B_DasWWJJw4_1),.dout(w_dff_B_mWMed6LW1_1),.clk(gclk));
	jdff dff_B_fOpm9S0e6_1(.din(w_dff_B_mWMed6LW1_1),.dout(w_dff_B_fOpm9S0e6_1),.clk(gclk));
	jdff dff_B_QMMBpxF42_1(.din(w_dff_B_fOpm9S0e6_1),.dout(w_dff_B_QMMBpxF42_1),.clk(gclk));
	jdff dff_B_rRAhMiLx1_1(.din(w_dff_B_QMMBpxF42_1),.dout(w_dff_B_rRAhMiLx1_1),.clk(gclk));
	jdff dff_B_Iogz5Cyt4_1(.din(w_dff_B_rRAhMiLx1_1),.dout(w_dff_B_Iogz5Cyt4_1),.clk(gclk));
	jdff dff_B_eMcL5tkk0_1(.din(w_dff_B_Iogz5Cyt4_1),.dout(w_dff_B_eMcL5tkk0_1),.clk(gclk));
	jdff dff_B_5UlNxpAs9_1(.din(w_dff_B_eMcL5tkk0_1),.dout(w_dff_B_5UlNxpAs9_1),.clk(gclk));
	jdff dff_B_2jjWzCxk8_1(.din(w_dff_B_5UlNxpAs9_1),.dout(w_dff_B_2jjWzCxk8_1),.clk(gclk));
	jdff dff_B_9SLRow335_1(.din(w_dff_B_2jjWzCxk8_1),.dout(w_dff_B_9SLRow335_1),.clk(gclk));
	jdff dff_B_7LXNU9WD0_1(.din(w_dff_B_9SLRow335_1),.dout(w_dff_B_7LXNU9WD0_1),.clk(gclk));
	jdff dff_B_YPTKF3bv0_1(.din(w_dff_B_7LXNU9WD0_1),.dout(w_dff_B_YPTKF3bv0_1),.clk(gclk));
	jdff dff_B_8YfUqkGs4_1(.din(w_dff_B_YPTKF3bv0_1),.dout(w_dff_B_8YfUqkGs4_1),.clk(gclk));
	jdff dff_B_RvV3B9Lk6_1(.din(w_dff_B_8YfUqkGs4_1),.dout(w_dff_B_RvV3B9Lk6_1),.clk(gclk));
	jdff dff_B_16YwknhO5_1(.din(w_dff_B_RvV3B9Lk6_1),.dout(w_dff_B_16YwknhO5_1),.clk(gclk));
	jdff dff_B_pCxzE4MB2_1(.din(w_dff_B_16YwknhO5_1),.dout(w_dff_B_pCxzE4MB2_1),.clk(gclk));
	jdff dff_B_80BoNJFi1_1(.din(w_dff_B_pCxzE4MB2_1),.dout(w_dff_B_80BoNJFi1_1),.clk(gclk));
	jdff dff_B_pm0YsuEi7_1(.din(w_dff_B_80BoNJFi1_1),.dout(w_dff_B_pm0YsuEi7_1),.clk(gclk));
	jdff dff_B_jh7lPzj90_1(.din(w_dff_B_pm0YsuEi7_1),.dout(w_dff_B_jh7lPzj90_1),.clk(gclk));
	jdff dff_B_XJpTwJ1N0_1(.din(w_dff_B_jh7lPzj90_1),.dout(w_dff_B_XJpTwJ1N0_1),.clk(gclk));
	jdff dff_B_TgmkPTjJ5_1(.din(w_dff_B_XJpTwJ1N0_1),.dout(w_dff_B_TgmkPTjJ5_1),.clk(gclk));
	jdff dff_B_MlefUiER5_1(.din(w_dff_B_TgmkPTjJ5_1),.dout(w_dff_B_MlefUiER5_1),.clk(gclk));
	jdff dff_B_BQFQkRKn1_1(.din(w_dff_B_MlefUiER5_1),.dout(w_dff_B_BQFQkRKn1_1),.clk(gclk));
	jdff dff_B_uKilCTj05_1(.din(w_dff_B_BQFQkRKn1_1),.dout(w_dff_B_uKilCTj05_1),.clk(gclk));
	jdff dff_B_rfi7v14r4_1(.din(w_dff_B_uKilCTj05_1),.dout(w_dff_B_rfi7v14r4_1),.clk(gclk));
	jdff dff_B_wOr8EqwB9_1(.din(w_dff_B_rfi7v14r4_1),.dout(w_dff_B_wOr8EqwB9_1),.clk(gclk));
	jdff dff_B_Y5ha6kkK4_1(.din(w_dff_B_wOr8EqwB9_1),.dout(w_dff_B_Y5ha6kkK4_1),.clk(gclk));
	jdff dff_B_agJMqJbA9_1(.din(w_dff_B_Y5ha6kkK4_1),.dout(w_dff_B_agJMqJbA9_1),.clk(gclk));
	jdff dff_B_7cWnK8Ja1_1(.din(w_dff_B_agJMqJbA9_1),.dout(w_dff_B_7cWnK8Ja1_1),.clk(gclk));
	jdff dff_B_lJyKqemu5_1(.din(w_dff_B_7cWnK8Ja1_1),.dout(w_dff_B_lJyKqemu5_1),.clk(gclk));
	jdff dff_B_gFAVYVfM6_1(.din(w_dff_B_lJyKqemu5_1),.dout(w_dff_B_gFAVYVfM6_1),.clk(gclk));
	jdff dff_B_wpEhMsoK1_1(.din(w_dff_B_gFAVYVfM6_1),.dout(w_dff_B_wpEhMsoK1_1),.clk(gclk));
	jdff dff_B_pMpQUgLF2_1(.din(w_dff_B_wpEhMsoK1_1),.dout(w_dff_B_pMpQUgLF2_1),.clk(gclk));
	jdff dff_B_R5Emixij0_1(.din(w_dff_B_pMpQUgLF2_1),.dout(w_dff_B_R5Emixij0_1),.clk(gclk));
	jdff dff_B_gAskS9d85_1(.din(w_dff_B_R5Emixij0_1),.dout(w_dff_B_gAskS9d85_1),.clk(gclk));
	jdff dff_B_SO7QG9tp3_1(.din(w_dff_B_gAskS9d85_1),.dout(w_dff_B_SO7QG9tp3_1),.clk(gclk));
	jdff dff_B_0LAQqcji3_1(.din(w_dff_B_SO7QG9tp3_1),.dout(w_dff_B_0LAQqcji3_1),.clk(gclk));
	jdff dff_B_wjK4LdHO2_1(.din(w_dff_B_0LAQqcji3_1),.dout(w_dff_B_wjK4LdHO2_1),.clk(gclk));
	jdff dff_B_m3Z1pYuz1_1(.din(w_dff_B_wjK4LdHO2_1),.dout(w_dff_B_m3Z1pYuz1_1),.clk(gclk));
	jdff dff_B_40pTdnTV4_1(.din(w_dff_B_m3Z1pYuz1_1),.dout(w_dff_B_40pTdnTV4_1),.clk(gclk));
	jdff dff_B_9cYSHblH7_1(.din(w_dff_B_40pTdnTV4_1),.dout(w_dff_B_9cYSHblH7_1),.clk(gclk));
	jdff dff_B_R0KXtrdP2_1(.din(w_dff_B_9cYSHblH7_1),.dout(w_dff_B_R0KXtrdP2_1),.clk(gclk));
	jdff dff_B_haSwwdUt8_1(.din(w_dff_B_R0KXtrdP2_1),.dout(w_dff_B_haSwwdUt8_1),.clk(gclk));
	jdff dff_B_vwQnEUg09_1(.din(w_dff_B_haSwwdUt8_1),.dout(w_dff_B_vwQnEUg09_1),.clk(gclk));
	jdff dff_B_IzzOXkwY4_1(.din(w_dff_B_vwQnEUg09_1),.dout(w_dff_B_IzzOXkwY4_1),.clk(gclk));
	jdff dff_B_OxkcOqHu1_1(.din(w_dff_B_IzzOXkwY4_1),.dout(w_dff_B_OxkcOqHu1_1),.clk(gclk));
	jdff dff_B_oGgbXCnT8_1(.din(w_dff_B_OxkcOqHu1_1),.dout(w_dff_B_oGgbXCnT8_1),.clk(gclk));
	jdff dff_B_7AuRGt5N5_1(.din(w_dff_B_oGgbXCnT8_1),.dout(w_dff_B_7AuRGt5N5_1),.clk(gclk));
	jdff dff_B_5r4wPzZq0_1(.din(w_dff_B_7AuRGt5N5_1),.dout(w_dff_B_5r4wPzZq0_1),.clk(gclk));
	jdff dff_B_yJ5n5j3l9_1(.din(w_dff_B_5r4wPzZq0_1),.dout(w_dff_B_yJ5n5j3l9_1),.clk(gclk));
	jdff dff_B_nFZjQded9_1(.din(w_dff_B_yJ5n5j3l9_1),.dout(w_dff_B_nFZjQded9_1),.clk(gclk));
	jdff dff_B_dUut2OlH6_1(.din(w_dff_B_nFZjQded9_1),.dout(w_dff_B_dUut2OlH6_1),.clk(gclk));
	jdff dff_B_oAvWXRvp2_1(.din(w_dff_B_dUut2OlH6_1),.dout(w_dff_B_oAvWXRvp2_1),.clk(gclk));
	jdff dff_B_9eImSTrN9_1(.din(w_dff_B_oAvWXRvp2_1),.dout(w_dff_B_9eImSTrN9_1),.clk(gclk));
	jdff dff_B_j3wGZEew6_1(.din(w_dff_B_9eImSTrN9_1),.dout(w_dff_B_j3wGZEew6_1),.clk(gclk));
	jdff dff_B_S52isB6i7_1(.din(w_dff_B_j3wGZEew6_1),.dout(w_dff_B_S52isB6i7_1),.clk(gclk));
	jdff dff_B_5RxK6jmr7_1(.din(w_dff_B_S52isB6i7_1),.dout(w_dff_B_5RxK6jmr7_1),.clk(gclk));
	jdff dff_B_SGuEypJX3_1(.din(w_dff_B_5RxK6jmr7_1),.dout(w_dff_B_SGuEypJX3_1),.clk(gclk));
	jdff dff_B_6HNUGjpl2_1(.din(w_dff_B_SGuEypJX3_1),.dout(w_dff_B_6HNUGjpl2_1),.clk(gclk));
	jdff dff_B_X2BqJM3K4_1(.din(w_dff_B_6HNUGjpl2_1),.dout(w_dff_B_X2BqJM3K4_1),.clk(gclk));
	jdff dff_B_2LKZDNeI3_1(.din(w_dff_B_X2BqJM3K4_1),.dout(w_dff_B_2LKZDNeI3_1),.clk(gclk));
	jdff dff_B_QhYOYsAE4_1(.din(w_dff_B_2LKZDNeI3_1),.dout(w_dff_B_QhYOYsAE4_1),.clk(gclk));
	jdff dff_B_zuJZW8bC6_1(.din(w_dff_B_QhYOYsAE4_1),.dout(w_dff_B_zuJZW8bC6_1),.clk(gclk));
	jdff dff_B_idOx3eYX8_1(.din(w_dff_B_zuJZW8bC6_1),.dout(w_dff_B_idOx3eYX8_1),.clk(gclk));
	jdff dff_B_7Tzfi5aE0_1(.din(w_dff_B_idOx3eYX8_1),.dout(w_dff_B_7Tzfi5aE0_1),.clk(gclk));
	jdff dff_B_Nee9REeW2_1(.din(w_dff_B_7Tzfi5aE0_1),.dout(w_dff_B_Nee9REeW2_1),.clk(gclk));
	jdff dff_B_a6PbQl1x4_1(.din(w_dff_B_Nee9REeW2_1),.dout(w_dff_B_a6PbQl1x4_1),.clk(gclk));
	jdff dff_B_kpwezgEs1_1(.din(w_dff_B_a6PbQl1x4_1),.dout(w_dff_B_kpwezgEs1_1),.clk(gclk));
	jdff dff_B_WKnQEFf81_1(.din(w_dff_B_kpwezgEs1_1),.dout(w_dff_B_WKnQEFf81_1),.clk(gclk));
	jdff dff_B_tN7muEOo9_1(.din(w_dff_B_WKnQEFf81_1),.dout(w_dff_B_tN7muEOo9_1),.clk(gclk));
	jdff dff_B_pj5Q2XNi2_1(.din(w_dff_B_tN7muEOo9_1),.dout(w_dff_B_pj5Q2XNi2_1),.clk(gclk));
	jdff dff_B_glfGUBZ16_1(.din(w_dff_B_pj5Q2XNi2_1),.dout(w_dff_B_glfGUBZ16_1),.clk(gclk));
	jdff dff_B_nXjSbwsS7_1(.din(w_dff_B_glfGUBZ16_1),.dout(w_dff_B_nXjSbwsS7_1),.clk(gclk));
	jdff dff_B_Gz2BeENo0_1(.din(w_dff_B_nXjSbwsS7_1),.dout(w_dff_B_Gz2BeENo0_1),.clk(gclk));
	jdff dff_B_8nUXdlyh2_1(.din(w_dff_B_Gz2BeENo0_1),.dout(w_dff_B_8nUXdlyh2_1),.clk(gclk));
	jdff dff_B_ECD4Emfb9_1(.din(w_dff_B_8nUXdlyh2_1),.dout(w_dff_B_ECD4Emfb9_1),.clk(gclk));
	jdff dff_B_1XgQn9YC1_1(.din(w_dff_B_ECD4Emfb9_1),.dout(w_dff_B_1XgQn9YC1_1),.clk(gclk));
	jdff dff_B_lUQjkxGn7_1(.din(w_dff_B_1XgQn9YC1_1),.dout(w_dff_B_lUQjkxGn7_1),.clk(gclk));
	jdff dff_B_qUO7qdcq1_1(.din(w_dff_B_lUQjkxGn7_1),.dout(w_dff_B_qUO7qdcq1_1),.clk(gclk));
	jdff dff_B_ZwrzRpIa0_1(.din(w_dff_B_qUO7qdcq1_1),.dout(w_dff_B_ZwrzRpIa0_1),.clk(gclk));
	jdff dff_B_r2zxWOiQ3_1(.din(w_dff_B_ZwrzRpIa0_1),.dout(w_dff_B_r2zxWOiQ3_1),.clk(gclk));
	jdff dff_B_wjrD4Gba7_1(.din(w_dff_B_r2zxWOiQ3_1),.dout(w_dff_B_wjrD4Gba7_1),.clk(gclk));
	jdff dff_B_omgaa8xX0_1(.din(w_dff_B_wjrD4Gba7_1),.dout(w_dff_B_omgaa8xX0_1),.clk(gclk));
	jdff dff_B_vpfARLRc8_1(.din(w_dff_B_omgaa8xX0_1),.dout(w_dff_B_vpfARLRc8_1),.clk(gclk));
	jdff dff_B_fFrIurs99_1(.din(w_dff_B_vpfARLRc8_1),.dout(w_dff_B_fFrIurs99_1),.clk(gclk));
	jdff dff_B_oO9qGIbb9_1(.din(w_dff_B_fFrIurs99_1),.dout(w_dff_B_oO9qGIbb9_1),.clk(gclk));
	jdff dff_B_kq1FULtz0_1(.din(w_dff_B_oO9qGIbb9_1),.dout(w_dff_B_kq1FULtz0_1),.clk(gclk));
	jdff dff_B_vzduoSy73_1(.din(w_dff_B_kq1FULtz0_1),.dout(w_dff_B_vzduoSy73_1),.clk(gclk));
	jdff dff_B_CSU5Exqh4_1(.din(w_dff_B_vzduoSy73_1),.dout(w_dff_B_CSU5Exqh4_1),.clk(gclk));
	jdff dff_B_eGVwxzAz7_1(.din(w_dff_B_CSU5Exqh4_1),.dout(w_dff_B_eGVwxzAz7_1),.clk(gclk));
	jdff dff_B_NhGUpUZd7_1(.din(w_dff_B_eGVwxzAz7_1),.dout(w_dff_B_NhGUpUZd7_1),.clk(gclk));
	jdff dff_B_Ymc7dSyE2_1(.din(w_dff_B_NhGUpUZd7_1),.dout(w_dff_B_Ymc7dSyE2_1),.clk(gclk));
	jdff dff_B_3aAy86DJ0_1(.din(w_dff_B_Ymc7dSyE2_1),.dout(w_dff_B_3aAy86DJ0_1),.clk(gclk));
	jdff dff_B_HLeWyBgG7_1(.din(w_dff_B_3aAy86DJ0_1),.dout(w_dff_B_HLeWyBgG7_1),.clk(gclk));
	jdff dff_B_k9kLOO4a2_1(.din(w_dff_B_HLeWyBgG7_1),.dout(w_dff_B_k9kLOO4a2_1),.clk(gclk));
	jdff dff_B_qEvwrYGp8_1(.din(w_dff_B_k9kLOO4a2_1),.dout(w_dff_B_qEvwrYGp8_1),.clk(gclk));
	jdff dff_B_P4oizCHC4_1(.din(w_dff_B_qEvwrYGp8_1),.dout(w_dff_B_P4oizCHC4_1),.clk(gclk));
	jdff dff_B_MvLDE62y9_1(.din(w_dff_B_P4oizCHC4_1),.dout(w_dff_B_MvLDE62y9_1),.clk(gclk));
	jdff dff_B_c8t4eMk40_1(.din(w_dff_B_MvLDE62y9_1),.dout(w_dff_B_c8t4eMk40_1),.clk(gclk));
	jdff dff_B_ST0q4Qjd2_1(.din(w_dff_B_c8t4eMk40_1),.dout(w_dff_B_ST0q4Qjd2_1),.clk(gclk));
	jdff dff_B_XxBlAudr6_1(.din(w_dff_B_ST0q4Qjd2_1),.dout(w_dff_B_XxBlAudr6_1),.clk(gclk));
	jdff dff_B_YGBlSZ3u7_1(.din(w_dff_B_XxBlAudr6_1),.dout(w_dff_B_YGBlSZ3u7_1),.clk(gclk));
	jdff dff_B_7Z2MS1fk0_1(.din(w_dff_B_YGBlSZ3u7_1),.dout(w_dff_B_7Z2MS1fk0_1),.clk(gclk));
	jdff dff_B_drTDZiCu1_1(.din(w_dff_B_7Z2MS1fk0_1),.dout(w_dff_B_drTDZiCu1_1),.clk(gclk));
	jdff dff_B_3iG0t9it0_1(.din(w_dff_B_drTDZiCu1_1),.dout(w_dff_B_3iG0t9it0_1),.clk(gclk));
	jdff dff_B_y9BNTbnt8_1(.din(w_dff_B_3iG0t9it0_1),.dout(w_dff_B_y9BNTbnt8_1),.clk(gclk));
	jdff dff_B_0nN0BSNX5_1(.din(w_dff_B_y9BNTbnt8_1),.dout(w_dff_B_0nN0BSNX5_1),.clk(gclk));
	jdff dff_B_CEcVRHjZ2_0(.din(n1081),.dout(w_dff_B_CEcVRHjZ2_0),.clk(gclk));
	jdff dff_B_rtlwDItD9_0(.din(w_dff_B_CEcVRHjZ2_0),.dout(w_dff_B_rtlwDItD9_0),.clk(gclk));
	jdff dff_B_of6DTMrQ5_0(.din(w_dff_B_rtlwDItD9_0),.dout(w_dff_B_of6DTMrQ5_0),.clk(gclk));
	jdff dff_B_aGCFd8mm2_0(.din(w_dff_B_of6DTMrQ5_0),.dout(w_dff_B_aGCFd8mm2_0),.clk(gclk));
	jdff dff_B_yZyw2owQ2_0(.din(w_dff_B_aGCFd8mm2_0),.dout(w_dff_B_yZyw2owQ2_0),.clk(gclk));
	jdff dff_B_Dlo29GBj3_0(.din(w_dff_B_yZyw2owQ2_0),.dout(w_dff_B_Dlo29GBj3_0),.clk(gclk));
	jdff dff_B_zbDTd6015_0(.din(w_dff_B_Dlo29GBj3_0),.dout(w_dff_B_zbDTd6015_0),.clk(gclk));
	jdff dff_B_eR62aRzx5_0(.din(w_dff_B_zbDTd6015_0),.dout(w_dff_B_eR62aRzx5_0),.clk(gclk));
	jdff dff_B_PZtNmySa7_0(.din(w_dff_B_eR62aRzx5_0),.dout(w_dff_B_PZtNmySa7_0),.clk(gclk));
	jdff dff_B_Rfo3o5cV2_0(.din(w_dff_B_PZtNmySa7_0),.dout(w_dff_B_Rfo3o5cV2_0),.clk(gclk));
	jdff dff_B_uSCRDwjQ9_0(.din(w_dff_B_Rfo3o5cV2_0),.dout(w_dff_B_uSCRDwjQ9_0),.clk(gclk));
	jdff dff_B_ctbF1Ulq7_0(.din(w_dff_B_uSCRDwjQ9_0),.dout(w_dff_B_ctbF1Ulq7_0),.clk(gclk));
	jdff dff_B_D07dR8wm2_0(.din(w_dff_B_ctbF1Ulq7_0),.dout(w_dff_B_D07dR8wm2_0),.clk(gclk));
	jdff dff_B_XaUGYvOY0_0(.din(w_dff_B_D07dR8wm2_0),.dout(w_dff_B_XaUGYvOY0_0),.clk(gclk));
	jdff dff_B_rVRna2Hg5_0(.din(w_dff_B_XaUGYvOY0_0),.dout(w_dff_B_rVRna2Hg5_0),.clk(gclk));
	jdff dff_B_xJHVUlZX9_0(.din(w_dff_B_rVRna2Hg5_0),.dout(w_dff_B_xJHVUlZX9_0),.clk(gclk));
	jdff dff_B_G8boljKA9_0(.din(w_dff_B_xJHVUlZX9_0),.dout(w_dff_B_G8boljKA9_0),.clk(gclk));
	jdff dff_B_d1IG8QGg3_0(.din(w_dff_B_G8boljKA9_0),.dout(w_dff_B_d1IG8QGg3_0),.clk(gclk));
	jdff dff_B_sr4Fp0DC8_0(.din(w_dff_B_d1IG8QGg3_0),.dout(w_dff_B_sr4Fp0DC8_0),.clk(gclk));
	jdff dff_B_AQh94kD40_0(.din(w_dff_B_sr4Fp0DC8_0),.dout(w_dff_B_AQh94kD40_0),.clk(gclk));
	jdff dff_B_Lp8ee4nw7_0(.din(w_dff_B_AQh94kD40_0),.dout(w_dff_B_Lp8ee4nw7_0),.clk(gclk));
	jdff dff_B_HYqQiyx82_0(.din(w_dff_B_Lp8ee4nw7_0),.dout(w_dff_B_HYqQiyx82_0),.clk(gclk));
	jdff dff_B_aQcdx7hr4_0(.din(w_dff_B_HYqQiyx82_0),.dout(w_dff_B_aQcdx7hr4_0),.clk(gclk));
	jdff dff_B_S2Wl7Q1L0_0(.din(w_dff_B_aQcdx7hr4_0),.dout(w_dff_B_S2Wl7Q1L0_0),.clk(gclk));
	jdff dff_B_nWgaLhR66_0(.din(w_dff_B_S2Wl7Q1L0_0),.dout(w_dff_B_nWgaLhR66_0),.clk(gclk));
	jdff dff_B_aXF9oQJA9_0(.din(w_dff_B_nWgaLhR66_0),.dout(w_dff_B_aXF9oQJA9_0),.clk(gclk));
	jdff dff_B_24trkB455_0(.din(w_dff_B_aXF9oQJA9_0),.dout(w_dff_B_24trkB455_0),.clk(gclk));
	jdff dff_B_I1UaNswh3_0(.din(w_dff_B_24trkB455_0),.dout(w_dff_B_I1UaNswh3_0),.clk(gclk));
	jdff dff_B_kBbz9s5V5_0(.din(w_dff_B_I1UaNswh3_0),.dout(w_dff_B_kBbz9s5V5_0),.clk(gclk));
	jdff dff_B_OaRGEu4p4_0(.din(w_dff_B_kBbz9s5V5_0),.dout(w_dff_B_OaRGEu4p4_0),.clk(gclk));
	jdff dff_B_3jpsfhIq4_0(.din(w_dff_B_OaRGEu4p4_0),.dout(w_dff_B_3jpsfhIq4_0),.clk(gclk));
	jdff dff_B_hb446n6I6_0(.din(w_dff_B_3jpsfhIq4_0),.dout(w_dff_B_hb446n6I6_0),.clk(gclk));
	jdff dff_B_vD5iaqfe1_0(.din(w_dff_B_hb446n6I6_0),.dout(w_dff_B_vD5iaqfe1_0),.clk(gclk));
	jdff dff_B_dbx7uHRZ9_0(.din(w_dff_B_vD5iaqfe1_0),.dout(w_dff_B_dbx7uHRZ9_0),.clk(gclk));
	jdff dff_B_2hUrxHKo4_0(.din(w_dff_B_dbx7uHRZ9_0),.dout(w_dff_B_2hUrxHKo4_0),.clk(gclk));
	jdff dff_B_hGpOnTPN3_0(.din(w_dff_B_2hUrxHKo4_0),.dout(w_dff_B_hGpOnTPN3_0),.clk(gclk));
	jdff dff_B_O15gnHGa9_0(.din(w_dff_B_hGpOnTPN3_0),.dout(w_dff_B_O15gnHGa9_0),.clk(gclk));
	jdff dff_B_dKN9ee4Y3_0(.din(w_dff_B_O15gnHGa9_0),.dout(w_dff_B_dKN9ee4Y3_0),.clk(gclk));
	jdff dff_B_yTcj7qUT3_0(.din(w_dff_B_dKN9ee4Y3_0),.dout(w_dff_B_yTcj7qUT3_0),.clk(gclk));
	jdff dff_B_ib5h5OsW0_0(.din(w_dff_B_yTcj7qUT3_0),.dout(w_dff_B_ib5h5OsW0_0),.clk(gclk));
	jdff dff_B_ddup17tU2_0(.din(w_dff_B_ib5h5OsW0_0),.dout(w_dff_B_ddup17tU2_0),.clk(gclk));
	jdff dff_B_2UOiuz2B8_0(.din(w_dff_B_ddup17tU2_0),.dout(w_dff_B_2UOiuz2B8_0),.clk(gclk));
	jdff dff_B_LUjfoTF04_0(.din(w_dff_B_2UOiuz2B8_0),.dout(w_dff_B_LUjfoTF04_0),.clk(gclk));
	jdff dff_B_GtbWfExF2_0(.din(w_dff_B_LUjfoTF04_0),.dout(w_dff_B_GtbWfExF2_0),.clk(gclk));
	jdff dff_B_HBYounN53_0(.din(w_dff_B_GtbWfExF2_0),.dout(w_dff_B_HBYounN53_0),.clk(gclk));
	jdff dff_B_mzyMEDLv4_0(.din(w_dff_B_HBYounN53_0),.dout(w_dff_B_mzyMEDLv4_0),.clk(gclk));
	jdff dff_B_MbtIKZL59_0(.din(w_dff_B_mzyMEDLv4_0),.dout(w_dff_B_MbtIKZL59_0),.clk(gclk));
	jdff dff_B_Pj03Arrf8_0(.din(w_dff_B_MbtIKZL59_0),.dout(w_dff_B_Pj03Arrf8_0),.clk(gclk));
	jdff dff_B_IyBTYlXi1_0(.din(w_dff_B_Pj03Arrf8_0),.dout(w_dff_B_IyBTYlXi1_0),.clk(gclk));
	jdff dff_B_8FEiPlDW9_0(.din(w_dff_B_IyBTYlXi1_0),.dout(w_dff_B_8FEiPlDW9_0),.clk(gclk));
	jdff dff_B_pqfQ7txp5_0(.din(w_dff_B_8FEiPlDW9_0),.dout(w_dff_B_pqfQ7txp5_0),.clk(gclk));
	jdff dff_B_dtxSjQuc6_0(.din(w_dff_B_pqfQ7txp5_0),.dout(w_dff_B_dtxSjQuc6_0),.clk(gclk));
	jdff dff_B_wifl28q81_0(.din(w_dff_B_dtxSjQuc6_0),.dout(w_dff_B_wifl28q81_0),.clk(gclk));
	jdff dff_B_SHW4TUzh0_0(.din(w_dff_B_wifl28q81_0),.dout(w_dff_B_SHW4TUzh0_0),.clk(gclk));
	jdff dff_B_selpxYZT2_0(.din(w_dff_B_SHW4TUzh0_0),.dout(w_dff_B_selpxYZT2_0),.clk(gclk));
	jdff dff_B_VBGAhItr7_0(.din(w_dff_B_selpxYZT2_0),.dout(w_dff_B_VBGAhItr7_0),.clk(gclk));
	jdff dff_B_HW5IhkaJ7_0(.din(w_dff_B_VBGAhItr7_0),.dout(w_dff_B_HW5IhkaJ7_0),.clk(gclk));
	jdff dff_B_iQMTKuhs4_0(.din(w_dff_B_HW5IhkaJ7_0),.dout(w_dff_B_iQMTKuhs4_0),.clk(gclk));
	jdff dff_B_TqCDsnul8_0(.din(w_dff_B_iQMTKuhs4_0),.dout(w_dff_B_TqCDsnul8_0),.clk(gclk));
	jdff dff_B_GBPh6MQS4_0(.din(w_dff_B_TqCDsnul8_0),.dout(w_dff_B_GBPh6MQS4_0),.clk(gclk));
	jdff dff_B_QI3oEd8p6_0(.din(w_dff_B_GBPh6MQS4_0),.dout(w_dff_B_QI3oEd8p6_0),.clk(gclk));
	jdff dff_B_LfXWihqg3_0(.din(w_dff_B_QI3oEd8p6_0),.dout(w_dff_B_LfXWihqg3_0),.clk(gclk));
	jdff dff_B_iM4xOC2P8_0(.din(w_dff_B_LfXWihqg3_0),.dout(w_dff_B_iM4xOC2P8_0),.clk(gclk));
	jdff dff_B_q8o5KloS6_0(.din(w_dff_B_iM4xOC2P8_0),.dout(w_dff_B_q8o5KloS6_0),.clk(gclk));
	jdff dff_B_Xtx4G3vh9_0(.din(w_dff_B_q8o5KloS6_0),.dout(w_dff_B_Xtx4G3vh9_0),.clk(gclk));
	jdff dff_B_OlsHckU21_0(.din(w_dff_B_Xtx4G3vh9_0),.dout(w_dff_B_OlsHckU21_0),.clk(gclk));
	jdff dff_B_fiU3edQc3_0(.din(w_dff_B_OlsHckU21_0),.dout(w_dff_B_fiU3edQc3_0),.clk(gclk));
	jdff dff_B_TfRCJYOG4_0(.din(w_dff_B_fiU3edQc3_0),.dout(w_dff_B_TfRCJYOG4_0),.clk(gclk));
	jdff dff_B_im0ifTAi2_0(.din(w_dff_B_TfRCJYOG4_0),.dout(w_dff_B_im0ifTAi2_0),.clk(gclk));
	jdff dff_B_G0vFep251_0(.din(w_dff_B_im0ifTAi2_0),.dout(w_dff_B_G0vFep251_0),.clk(gclk));
	jdff dff_B_RGRYrxUn1_0(.din(w_dff_B_G0vFep251_0),.dout(w_dff_B_RGRYrxUn1_0),.clk(gclk));
	jdff dff_B_hC79WNhS4_0(.din(w_dff_B_RGRYrxUn1_0),.dout(w_dff_B_hC79WNhS4_0),.clk(gclk));
	jdff dff_B_dZ5dLyHX5_0(.din(w_dff_B_hC79WNhS4_0),.dout(w_dff_B_dZ5dLyHX5_0),.clk(gclk));
	jdff dff_B_52nLrKKd8_0(.din(w_dff_B_dZ5dLyHX5_0),.dout(w_dff_B_52nLrKKd8_0),.clk(gclk));
	jdff dff_B_4bzjMXpP9_0(.din(w_dff_B_52nLrKKd8_0),.dout(w_dff_B_4bzjMXpP9_0),.clk(gclk));
	jdff dff_B_U0vtRxJ48_0(.din(w_dff_B_4bzjMXpP9_0),.dout(w_dff_B_U0vtRxJ48_0),.clk(gclk));
	jdff dff_B_TJG1b6v82_0(.din(w_dff_B_U0vtRxJ48_0),.dout(w_dff_B_TJG1b6v82_0),.clk(gclk));
	jdff dff_B_AQV777Rz8_0(.din(w_dff_B_TJG1b6v82_0),.dout(w_dff_B_AQV777Rz8_0),.clk(gclk));
	jdff dff_B_20FlKqlq1_0(.din(w_dff_B_AQV777Rz8_0),.dout(w_dff_B_20FlKqlq1_0),.clk(gclk));
	jdff dff_B_pAha6tjz5_0(.din(w_dff_B_20FlKqlq1_0),.dout(w_dff_B_pAha6tjz5_0),.clk(gclk));
	jdff dff_B_PvD6pQJi1_0(.din(w_dff_B_pAha6tjz5_0),.dout(w_dff_B_PvD6pQJi1_0),.clk(gclk));
	jdff dff_B_hN9yoSho4_0(.din(w_dff_B_PvD6pQJi1_0),.dout(w_dff_B_hN9yoSho4_0),.clk(gclk));
	jdff dff_B_yKt2x2n35_0(.din(w_dff_B_hN9yoSho4_0),.dout(w_dff_B_yKt2x2n35_0),.clk(gclk));
	jdff dff_B_fzOSd82d7_0(.din(w_dff_B_yKt2x2n35_0),.dout(w_dff_B_fzOSd82d7_0),.clk(gclk));
	jdff dff_B_nxMiRQsR4_0(.din(w_dff_B_fzOSd82d7_0),.dout(w_dff_B_nxMiRQsR4_0),.clk(gclk));
	jdff dff_B_jWjuFFjz3_0(.din(w_dff_B_nxMiRQsR4_0),.dout(w_dff_B_jWjuFFjz3_0),.clk(gclk));
	jdff dff_B_QUhzDHYV7_0(.din(w_dff_B_jWjuFFjz3_0),.dout(w_dff_B_QUhzDHYV7_0),.clk(gclk));
	jdff dff_B_UhNmhSVy5_0(.din(w_dff_B_QUhzDHYV7_0),.dout(w_dff_B_UhNmhSVy5_0),.clk(gclk));
	jdff dff_B_FWBfXhrK8_0(.din(w_dff_B_UhNmhSVy5_0),.dout(w_dff_B_FWBfXhrK8_0),.clk(gclk));
	jdff dff_B_8b2KP5PT2_0(.din(w_dff_B_FWBfXhrK8_0),.dout(w_dff_B_8b2KP5PT2_0),.clk(gclk));
	jdff dff_B_WnWnmiv69_0(.din(w_dff_B_8b2KP5PT2_0),.dout(w_dff_B_WnWnmiv69_0),.clk(gclk));
	jdff dff_B_QJWQ2UHw3_0(.din(w_dff_B_WnWnmiv69_0),.dout(w_dff_B_QJWQ2UHw3_0),.clk(gclk));
	jdff dff_B_RhzAqGUo2_0(.din(w_dff_B_QJWQ2UHw3_0),.dout(w_dff_B_RhzAqGUo2_0),.clk(gclk));
	jdff dff_B_objedPYf6_0(.din(w_dff_B_RhzAqGUo2_0),.dout(w_dff_B_objedPYf6_0),.clk(gclk));
	jdff dff_B_6keo17Jm9_0(.din(w_dff_B_objedPYf6_0),.dout(w_dff_B_6keo17Jm9_0),.clk(gclk));
	jdff dff_B_e7wX5awP2_0(.din(w_dff_B_6keo17Jm9_0),.dout(w_dff_B_e7wX5awP2_0),.clk(gclk));
	jdff dff_B_3m9OCgPF3_0(.din(w_dff_B_e7wX5awP2_0),.dout(w_dff_B_3m9OCgPF3_0),.clk(gclk));
	jdff dff_B_4N8ppNo25_0(.din(w_dff_B_3m9OCgPF3_0),.dout(w_dff_B_4N8ppNo25_0),.clk(gclk));
	jdff dff_B_FTJBg4vB8_0(.din(w_dff_B_4N8ppNo25_0),.dout(w_dff_B_FTJBg4vB8_0),.clk(gclk));
	jdff dff_B_5vL8vtHN2_0(.din(w_dff_B_FTJBg4vB8_0),.dout(w_dff_B_5vL8vtHN2_0),.clk(gclk));
	jdff dff_B_jTacgAvb5_0(.din(w_dff_B_5vL8vtHN2_0),.dout(w_dff_B_jTacgAvb5_0),.clk(gclk));
	jdff dff_B_KxjvUQzK3_0(.din(w_dff_B_jTacgAvb5_0),.dout(w_dff_B_KxjvUQzK3_0),.clk(gclk));
	jdff dff_B_mtt3OAM07_0(.din(w_dff_B_KxjvUQzK3_0),.dout(w_dff_B_mtt3OAM07_0),.clk(gclk));
	jdff dff_B_JNEE5kdi4_0(.din(w_dff_B_mtt3OAM07_0),.dout(w_dff_B_JNEE5kdi4_0),.clk(gclk));
	jdff dff_B_qZNb5GWQ4_0(.din(w_dff_B_JNEE5kdi4_0),.dout(w_dff_B_qZNb5GWQ4_0),.clk(gclk));
	jdff dff_B_w9DRzh0n4_0(.din(w_dff_B_qZNb5GWQ4_0),.dout(w_dff_B_w9DRzh0n4_0),.clk(gclk));
	jdff dff_B_YHspHjoT1_0(.din(w_dff_B_w9DRzh0n4_0),.dout(w_dff_B_YHspHjoT1_0),.clk(gclk));
	jdff dff_B_2BPQpjbO1_0(.din(w_dff_B_YHspHjoT1_0),.dout(w_dff_B_2BPQpjbO1_0),.clk(gclk));
	jdff dff_B_kA9YYPZO5_0(.din(w_dff_B_2BPQpjbO1_0),.dout(w_dff_B_kA9YYPZO5_0),.clk(gclk));
	jdff dff_B_vtBo1Mg96_0(.din(w_dff_B_kA9YYPZO5_0),.dout(w_dff_B_vtBo1Mg96_0),.clk(gclk));
	jdff dff_B_6X3X32i51_0(.din(w_dff_B_vtBo1Mg96_0),.dout(w_dff_B_6X3X32i51_0),.clk(gclk));
	jdff dff_B_mMX3SkrN1_0(.din(w_dff_B_6X3X32i51_0),.dout(w_dff_B_mMX3SkrN1_0),.clk(gclk));
	jdff dff_B_ImCUCeM42_0(.din(w_dff_B_mMX3SkrN1_0),.dout(w_dff_B_ImCUCeM42_0),.clk(gclk));
	jdff dff_B_GTZSpFw73_0(.din(w_dff_B_ImCUCeM42_0),.dout(w_dff_B_GTZSpFw73_0),.clk(gclk));
	jdff dff_B_QRImenJk5_0(.din(w_dff_B_GTZSpFw73_0),.dout(w_dff_B_QRImenJk5_0),.clk(gclk));
	jdff dff_B_k7K9XKQ61_0(.din(w_dff_B_QRImenJk5_0),.dout(w_dff_B_k7K9XKQ61_0),.clk(gclk));
	jdff dff_B_J6E6OeuB3_1(.din(n1074),.dout(w_dff_B_J6E6OeuB3_1),.clk(gclk));
	jdff dff_B_ekydRNRm6_1(.din(w_dff_B_J6E6OeuB3_1),.dout(w_dff_B_ekydRNRm6_1),.clk(gclk));
	jdff dff_B_suaHM4gB9_1(.din(w_dff_B_ekydRNRm6_1),.dout(w_dff_B_suaHM4gB9_1),.clk(gclk));
	jdff dff_B_5EltmYY89_1(.din(w_dff_B_suaHM4gB9_1),.dout(w_dff_B_5EltmYY89_1),.clk(gclk));
	jdff dff_B_lD71pSi28_1(.din(w_dff_B_5EltmYY89_1),.dout(w_dff_B_lD71pSi28_1),.clk(gclk));
	jdff dff_B_u8T8jq7S0_1(.din(w_dff_B_lD71pSi28_1),.dout(w_dff_B_u8T8jq7S0_1),.clk(gclk));
	jdff dff_B_NE17rn8J7_1(.din(w_dff_B_u8T8jq7S0_1),.dout(w_dff_B_NE17rn8J7_1),.clk(gclk));
	jdff dff_B_yBgVfDsw0_1(.din(w_dff_B_NE17rn8J7_1),.dout(w_dff_B_yBgVfDsw0_1),.clk(gclk));
	jdff dff_B_AATsKAgO0_1(.din(w_dff_B_yBgVfDsw0_1),.dout(w_dff_B_AATsKAgO0_1),.clk(gclk));
	jdff dff_B_GiCsjwu04_1(.din(w_dff_B_AATsKAgO0_1),.dout(w_dff_B_GiCsjwu04_1),.clk(gclk));
	jdff dff_B_qlHzmWSj8_1(.din(w_dff_B_GiCsjwu04_1),.dout(w_dff_B_qlHzmWSj8_1),.clk(gclk));
	jdff dff_B_Gx5ECXYr8_1(.din(w_dff_B_qlHzmWSj8_1),.dout(w_dff_B_Gx5ECXYr8_1),.clk(gclk));
	jdff dff_B_poKQ7djP9_1(.din(w_dff_B_Gx5ECXYr8_1),.dout(w_dff_B_poKQ7djP9_1),.clk(gclk));
	jdff dff_B_vTuWXpzW1_1(.din(w_dff_B_poKQ7djP9_1),.dout(w_dff_B_vTuWXpzW1_1),.clk(gclk));
	jdff dff_B_aims8asC2_1(.din(w_dff_B_vTuWXpzW1_1),.dout(w_dff_B_aims8asC2_1),.clk(gclk));
	jdff dff_B_ET657AIj5_1(.din(w_dff_B_aims8asC2_1),.dout(w_dff_B_ET657AIj5_1),.clk(gclk));
	jdff dff_B_ahSjjnQt0_1(.din(w_dff_B_ET657AIj5_1),.dout(w_dff_B_ahSjjnQt0_1),.clk(gclk));
	jdff dff_B_5Nle80dz1_1(.din(w_dff_B_ahSjjnQt0_1),.dout(w_dff_B_5Nle80dz1_1),.clk(gclk));
	jdff dff_B_tPvJuUk45_1(.din(w_dff_B_5Nle80dz1_1),.dout(w_dff_B_tPvJuUk45_1),.clk(gclk));
	jdff dff_B_BVn2FPyB8_1(.din(w_dff_B_tPvJuUk45_1),.dout(w_dff_B_BVn2FPyB8_1),.clk(gclk));
	jdff dff_B_HlVO66GQ5_1(.din(w_dff_B_BVn2FPyB8_1),.dout(w_dff_B_HlVO66GQ5_1),.clk(gclk));
	jdff dff_B_u0lvtJJE5_1(.din(w_dff_B_HlVO66GQ5_1),.dout(w_dff_B_u0lvtJJE5_1),.clk(gclk));
	jdff dff_B_RVNTHlCb6_1(.din(w_dff_B_u0lvtJJE5_1),.dout(w_dff_B_RVNTHlCb6_1),.clk(gclk));
	jdff dff_B_SuN8QHy73_1(.din(w_dff_B_RVNTHlCb6_1),.dout(w_dff_B_SuN8QHy73_1),.clk(gclk));
	jdff dff_B_TUfV9tun7_1(.din(w_dff_B_SuN8QHy73_1),.dout(w_dff_B_TUfV9tun7_1),.clk(gclk));
	jdff dff_B_E6WB9u2o6_1(.din(w_dff_B_TUfV9tun7_1),.dout(w_dff_B_E6WB9u2o6_1),.clk(gclk));
	jdff dff_B_KUEmSiAk1_1(.din(w_dff_B_E6WB9u2o6_1),.dout(w_dff_B_KUEmSiAk1_1),.clk(gclk));
	jdff dff_B_BQQkszUf4_1(.din(w_dff_B_KUEmSiAk1_1),.dout(w_dff_B_BQQkszUf4_1),.clk(gclk));
	jdff dff_B_BtVFA8sJ2_1(.din(w_dff_B_BQQkszUf4_1),.dout(w_dff_B_BtVFA8sJ2_1),.clk(gclk));
	jdff dff_B_crFtoYkU7_1(.din(w_dff_B_BtVFA8sJ2_1),.dout(w_dff_B_crFtoYkU7_1),.clk(gclk));
	jdff dff_B_DN9HcD6v8_1(.din(w_dff_B_crFtoYkU7_1),.dout(w_dff_B_DN9HcD6v8_1),.clk(gclk));
	jdff dff_B_oXzvce9N8_1(.din(w_dff_B_DN9HcD6v8_1),.dout(w_dff_B_oXzvce9N8_1),.clk(gclk));
	jdff dff_B_sQSF0xzh9_1(.din(w_dff_B_oXzvce9N8_1),.dout(w_dff_B_sQSF0xzh9_1),.clk(gclk));
	jdff dff_B_CXs5HuYa5_1(.din(w_dff_B_sQSF0xzh9_1),.dout(w_dff_B_CXs5HuYa5_1),.clk(gclk));
	jdff dff_B_vbxfDsLv8_1(.din(w_dff_B_CXs5HuYa5_1),.dout(w_dff_B_vbxfDsLv8_1),.clk(gclk));
	jdff dff_B_NBisfOiF6_1(.din(w_dff_B_vbxfDsLv8_1),.dout(w_dff_B_NBisfOiF6_1),.clk(gclk));
	jdff dff_B_SjS2hqwN4_1(.din(w_dff_B_NBisfOiF6_1),.dout(w_dff_B_SjS2hqwN4_1),.clk(gclk));
	jdff dff_B_pCJ7e4FS0_1(.din(w_dff_B_SjS2hqwN4_1),.dout(w_dff_B_pCJ7e4FS0_1),.clk(gclk));
	jdff dff_B_zTB39jfD1_1(.din(w_dff_B_pCJ7e4FS0_1),.dout(w_dff_B_zTB39jfD1_1),.clk(gclk));
	jdff dff_B_c9y4j0191_1(.din(w_dff_B_zTB39jfD1_1),.dout(w_dff_B_c9y4j0191_1),.clk(gclk));
	jdff dff_B_VQULySjX2_1(.din(w_dff_B_c9y4j0191_1),.dout(w_dff_B_VQULySjX2_1),.clk(gclk));
	jdff dff_B_2RLTwiEG8_1(.din(w_dff_B_VQULySjX2_1),.dout(w_dff_B_2RLTwiEG8_1),.clk(gclk));
	jdff dff_B_xP8l1tt87_1(.din(w_dff_B_2RLTwiEG8_1),.dout(w_dff_B_xP8l1tt87_1),.clk(gclk));
	jdff dff_B_qId6cRTo7_1(.din(w_dff_B_xP8l1tt87_1),.dout(w_dff_B_qId6cRTo7_1),.clk(gclk));
	jdff dff_B_2STgaVi67_1(.din(w_dff_B_qId6cRTo7_1),.dout(w_dff_B_2STgaVi67_1),.clk(gclk));
	jdff dff_B_KDy1Bz6A2_1(.din(w_dff_B_2STgaVi67_1),.dout(w_dff_B_KDy1Bz6A2_1),.clk(gclk));
	jdff dff_B_IpbddDJP9_1(.din(w_dff_B_KDy1Bz6A2_1),.dout(w_dff_B_IpbddDJP9_1),.clk(gclk));
	jdff dff_B_P0XRYMY91_1(.din(w_dff_B_IpbddDJP9_1),.dout(w_dff_B_P0XRYMY91_1),.clk(gclk));
	jdff dff_B_RHvkn7l22_1(.din(w_dff_B_P0XRYMY91_1),.dout(w_dff_B_RHvkn7l22_1),.clk(gclk));
	jdff dff_B_08w6AZx02_1(.din(w_dff_B_RHvkn7l22_1),.dout(w_dff_B_08w6AZx02_1),.clk(gclk));
	jdff dff_B_5pmxiRyR9_1(.din(w_dff_B_08w6AZx02_1),.dout(w_dff_B_5pmxiRyR9_1),.clk(gclk));
	jdff dff_B_L6DvscGH8_1(.din(w_dff_B_5pmxiRyR9_1),.dout(w_dff_B_L6DvscGH8_1),.clk(gclk));
	jdff dff_B_pupEmGhs4_1(.din(w_dff_B_L6DvscGH8_1),.dout(w_dff_B_pupEmGhs4_1),.clk(gclk));
	jdff dff_B_DeJ34ZzK6_1(.din(w_dff_B_pupEmGhs4_1),.dout(w_dff_B_DeJ34ZzK6_1),.clk(gclk));
	jdff dff_B_GIgX8GWm1_1(.din(w_dff_B_DeJ34ZzK6_1),.dout(w_dff_B_GIgX8GWm1_1),.clk(gclk));
	jdff dff_B_xCUqtNJg5_1(.din(w_dff_B_GIgX8GWm1_1),.dout(w_dff_B_xCUqtNJg5_1),.clk(gclk));
	jdff dff_B_Jcg7lNh85_1(.din(w_dff_B_xCUqtNJg5_1),.dout(w_dff_B_Jcg7lNh85_1),.clk(gclk));
	jdff dff_B_EqrXVh3y8_1(.din(w_dff_B_Jcg7lNh85_1),.dout(w_dff_B_EqrXVh3y8_1),.clk(gclk));
	jdff dff_B_LbTHXGcd5_1(.din(w_dff_B_EqrXVh3y8_1),.dout(w_dff_B_LbTHXGcd5_1),.clk(gclk));
	jdff dff_B_FjYwjX1l2_1(.din(w_dff_B_LbTHXGcd5_1),.dout(w_dff_B_FjYwjX1l2_1),.clk(gclk));
	jdff dff_B_Wtk5BMNj5_1(.din(w_dff_B_FjYwjX1l2_1),.dout(w_dff_B_Wtk5BMNj5_1),.clk(gclk));
	jdff dff_B_5yVe6hZN7_1(.din(w_dff_B_Wtk5BMNj5_1),.dout(w_dff_B_5yVe6hZN7_1),.clk(gclk));
	jdff dff_B_56GWUrSm9_1(.din(w_dff_B_5yVe6hZN7_1),.dout(w_dff_B_56GWUrSm9_1),.clk(gclk));
	jdff dff_B_8R9OaSo16_1(.din(w_dff_B_56GWUrSm9_1),.dout(w_dff_B_8R9OaSo16_1),.clk(gclk));
	jdff dff_B_81DG4xZv0_1(.din(w_dff_B_8R9OaSo16_1),.dout(w_dff_B_81DG4xZv0_1),.clk(gclk));
	jdff dff_B_hvsfi7SJ6_1(.din(w_dff_B_81DG4xZv0_1),.dout(w_dff_B_hvsfi7SJ6_1),.clk(gclk));
	jdff dff_B_HLXjHnPc8_1(.din(w_dff_B_hvsfi7SJ6_1),.dout(w_dff_B_HLXjHnPc8_1),.clk(gclk));
	jdff dff_B_xDhUz0eA5_1(.din(w_dff_B_HLXjHnPc8_1),.dout(w_dff_B_xDhUz0eA5_1),.clk(gclk));
	jdff dff_B_23oKKmbI4_1(.din(w_dff_B_xDhUz0eA5_1),.dout(w_dff_B_23oKKmbI4_1),.clk(gclk));
	jdff dff_B_2emqIVQY5_1(.din(w_dff_B_23oKKmbI4_1),.dout(w_dff_B_2emqIVQY5_1),.clk(gclk));
	jdff dff_B_JKcatsSO6_1(.din(w_dff_B_2emqIVQY5_1),.dout(w_dff_B_JKcatsSO6_1),.clk(gclk));
	jdff dff_B_LghcBRfS2_1(.din(w_dff_B_JKcatsSO6_1),.dout(w_dff_B_LghcBRfS2_1),.clk(gclk));
	jdff dff_B_JpVDBtyl4_1(.din(w_dff_B_LghcBRfS2_1),.dout(w_dff_B_JpVDBtyl4_1),.clk(gclk));
	jdff dff_B_pA2MZHhR0_1(.din(w_dff_B_JpVDBtyl4_1),.dout(w_dff_B_pA2MZHhR0_1),.clk(gclk));
	jdff dff_B_JtLkvqGU5_1(.din(w_dff_B_pA2MZHhR0_1),.dout(w_dff_B_JtLkvqGU5_1),.clk(gclk));
	jdff dff_B_fzcsPpco2_1(.din(w_dff_B_JtLkvqGU5_1),.dout(w_dff_B_fzcsPpco2_1),.clk(gclk));
	jdff dff_B_aEjRS6Me4_1(.din(w_dff_B_fzcsPpco2_1),.dout(w_dff_B_aEjRS6Me4_1),.clk(gclk));
	jdff dff_B_SXLNZ0VT1_1(.din(w_dff_B_aEjRS6Me4_1),.dout(w_dff_B_SXLNZ0VT1_1),.clk(gclk));
	jdff dff_B_AMj6Dc9L6_1(.din(w_dff_B_SXLNZ0VT1_1),.dout(w_dff_B_AMj6Dc9L6_1),.clk(gclk));
	jdff dff_B_pLuib1cd8_1(.din(w_dff_B_AMj6Dc9L6_1),.dout(w_dff_B_pLuib1cd8_1),.clk(gclk));
	jdff dff_B_1JDqF20i7_1(.din(w_dff_B_pLuib1cd8_1),.dout(w_dff_B_1JDqF20i7_1),.clk(gclk));
	jdff dff_B_kGF785tx7_1(.din(w_dff_B_1JDqF20i7_1),.dout(w_dff_B_kGF785tx7_1),.clk(gclk));
	jdff dff_B_i3F51tK17_1(.din(w_dff_B_kGF785tx7_1),.dout(w_dff_B_i3F51tK17_1),.clk(gclk));
	jdff dff_B_EoSNBCoy9_1(.din(w_dff_B_i3F51tK17_1),.dout(w_dff_B_EoSNBCoy9_1),.clk(gclk));
	jdff dff_B_L6UfDWSe7_1(.din(w_dff_B_EoSNBCoy9_1),.dout(w_dff_B_L6UfDWSe7_1),.clk(gclk));
	jdff dff_B_iePPLRq35_1(.din(w_dff_B_L6UfDWSe7_1),.dout(w_dff_B_iePPLRq35_1),.clk(gclk));
	jdff dff_B_qD8wQudE5_1(.din(w_dff_B_iePPLRq35_1),.dout(w_dff_B_qD8wQudE5_1),.clk(gclk));
	jdff dff_B_MxFvXjqI2_1(.din(w_dff_B_qD8wQudE5_1),.dout(w_dff_B_MxFvXjqI2_1),.clk(gclk));
	jdff dff_B_ghFUSEBb1_1(.din(w_dff_B_MxFvXjqI2_1),.dout(w_dff_B_ghFUSEBb1_1),.clk(gclk));
	jdff dff_B_nsOANQZh1_1(.din(w_dff_B_ghFUSEBb1_1),.dout(w_dff_B_nsOANQZh1_1),.clk(gclk));
	jdff dff_B_DE0PeJcg4_1(.din(w_dff_B_nsOANQZh1_1),.dout(w_dff_B_DE0PeJcg4_1),.clk(gclk));
	jdff dff_B_i4sfX0Pi6_1(.din(w_dff_B_DE0PeJcg4_1),.dout(w_dff_B_i4sfX0Pi6_1),.clk(gclk));
	jdff dff_B_S3nrAXFr5_1(.din(w_dff_B_i4sfX0Pi6_1),.dout(w_dff_B_S3nrAXFr5_1),.clk(gclk));
	jdff dff_B_u6tmZq4Y7_1(.din(w_dff_B_S3nrAXFr5_1),.dout(w_dff_B_u6tmZq4Y7_1),.clk(gclk));
	jdff dff_B_pyCIjXkf4_1(.din(w_dff_B_u6tmZq4Y7_1),.dout(w_dff_B_pyCIjXkf4_1),.clk(gclk));
	jdff dff_B_QnA1DRYy5_1(.din(w_dff_B_pyCIjXkf4_1),.dout(w_dff_B_QnA1DRYy5_1),.clk(gclk));
	jdff dff_B_9MMvWxuV1_1(.din(w_dff_B_QnA1DRYy5_1),.dout(w_dff_B_9MMvWxuV1_1),.clk(gclk));
	jdff dff_B_sxf07jmx3_1(.din(w_dff_B_9MMvWxuV1_1),.dout(w_dff_B_sxf07jmx3_1),.clk(gclk));
	jdff dff_B_I6aAMcYr7_1(.din(w_dff_B_sxf07jmx3_1),.dout(w_dff_B_I6aAMcYr7_1),.clk(gclk));
	jdff dff_B_TOH2blfR3_1(.din(w_dff_B_I6aAMcYr7_1),.dout(w_dff_B_TOH2blfR3_1),.clk(gclk));
	jdff dff_B_sJRHqjKW8_1(.din(w_dff_B_TOH2blfR3_1),.dout(w_dff_B_sJRHqjKW8_1),.clk(gclk));
	jdff dff_B_DMXGwRS08_1(.din(w_dff_B_sJRHqjKW8_1),.dout(w_dff_B_DMXGwRS08_1),.clk(gclk));
	jdff dff_B_3ppe9bG11_1(.din(w_dff_B_DMXGwRS08_1),.dout(w_dff_B_3ppe9bG11_1),.clk(gclk));
	jdff dff_B_GVRlRWhZ4_1(.din(w_dff_B_3ppe9bG11_1),.dout(w_dff_B_GVRlRWhZ4_1),.clk(gclk));
	jdff dff_B_SEb04kH37_1(.din(w_dff_B_GVRlRWhZ4_1),.dout(w_dff_B_SEb04kH37_1),.clk(gclk));
	jdff dff_B_V6SJyvHn0_1(.din(w_dff_B_SEb04kH37_1),.dout(w_dff_B_V6SJyvHn0_1),.clk(gclk));
	jdff dff_B_brRxbKFR7_1(.din(w_dff_B_V6SJyvHn0_1),.dout(w_dff_B_brRxbKFR7_1),.clk(gclk));
	jdff dff_B_ME5l3UJt3_1(.din(w_dff_B_brRxbKFR7_1),.dout(w_dff_B_ME5l3UJt3_1),.clk(gclk));
	jdff dff_B_mvUyxB3H1_1(.din(w_dff_B_ME5l3UJt3_1),.dout(w_dff_B_mvUyxB3H1_1),.clk(gclk));
	jdff dff_B_Wa3rStW03_1(.din(w_dff_B_mvUyxB3H1_1),.dout(w_dff_B_Wa3rStW03_1),.clk(gclk));
	jdff dff_B_P9Er4em07_1(.din(w_dff_B_Wa3rStW03_1),.dout(w_dff_B_P9Er4em07_1),.clk(gclk));
	jdff dff_B_TUvV9uPf5_1(.din(w_dff_B_P9Er4em07_1),.dout(w_dff_B_TUvV9uPf5_1),.clk(gclk));
	jdff dff_B_XqHKqY9F6_1(.din(w_dff_B_TUvV9uPf5_1),.dout(w_dff_B_XqHKqY9F6_1),.clk(gclk));
	jdff dff_B_Calt62xu3_1(.din(w_dff_B_XqHKqY9F6_1),.dout(w_dff_B_Calt62xu3_1),.clk(gclk));
	jdff dff_B_DmeXqhOy3_1(.din(w_dff_B_Calt62xu3_1),.dout(w_dff_B_DmeXqhOy3_1),.clk(gclk));
	jdff dff_B_pfbTqXXG1_0(.din(n1075),.dout(w_dff_B_pfbTqXXG1_0),.clk(gclk));
	jdff dff_B_Uw8Pseyl7_0(.din(w_dff_B_pfbTqXXG1_0),.dout(w_dff_B_Uw8Pseyl7_0),.clk(gclk));
	jdff dff_B_7fLCgk2S3_0(.din(w_dff_B_Uw8Pseyl7_0),.dout(w_dff_B_7fLCgk2S3_0),.clk(gclk));
	jdff dff_B_MmQqyFOf1_0(.din(w_dff_B_7fLCgk2S3_0),.dout(w_dff_B_MmQqyFOf1_0),.clk(gclk));
	jdff dff_B_itpXekh08_0(.din(w_dff_B_MmQqyFOf1_0),.dout(w_dff_B_itpXekh08_0),.clk(gclk));
	jdff dff_B_h23wqXfC7_0(.din(w_dff_B_itpXekh08_0),.dout(w_dff_B_h23wqXfC7_0),.clk(gclk));
	jdff dff_B_DOUJuvoL0_0(.din(w_dff_B_h23wqXfC7_0),.dout(w_dff_B_DOUJuvoL0_0),.clk(gclk));
	jdff dff_B_2j34fPCF0_0(.din(w_dff_B_DOUJuvoL0_0),.dout(w_dff_B_2j34fPCF0_0),.clk(gclk));
	jdff dff_B_QHYXr5C66_0(.din(w_dff_B_2j34fPCF0_0),.dout(w_dff_B_QHYXr5C66_0),.clk(gclk));
	jdff dff_B_ABtQpvYU0_0(.din(w_dff_B_QHYXr5C66_0),.dout(w_dff_B_ABtQpvYU0_0),.clk(gclk));
	jdff dff_B_nL1OYnUx2_0(.din(w_dff_B_ABtQpvYU0_0),.dout(w_dff_B_nL1OYnUx2_0),.clk(gclk));
	jdff dff_B_XzTRCcCo3_0(.din(w_dff_B_nL1OYnUx2_0),.dout(w_dff_B_XzTRCcCo3_0),.clk(gclk));
	jdff dff_B_b9FQ16xm8_0(.din(w_dff_B_XzTRCcCo3_0),.dout(w_dff_B_b9FQ16xm8_0),.clk(gclk));
	jdff dff_B_4vLICp688_0(.din(w_dff_B_b9FQ16xm8_0),.dout(w_dff_B_4vLICp688_0),.clk(gclk));
	jdff dff_B_Yv3JoQzG6_0(.din(w_dff_B_4vLICp688_0),.dout(w_dff_B_Yv3JoQzG6_0),.clk(gclk));
	jdff dff_B_QQNqunm91_0(.din(w_dff_B_Yv3JoQzG6_0),.dout(w_dff_B_QQNqunm91_0),.clk(gclk));
	jdff dff_B_pZb2KrV00_0(.din(w_dff_B_QQNqunm91_0),.dout(w_dff_B_pZb2KrV00_0),.clk(gclk));
	jdff dff_B_Q4ztJBHL6_0(.din(w_dff_B_pZb2KrV00_0),.dout(w_dff_B_Q4ztJBHL6_0),.clk(gclk));
	jdff dff_B_SmBl1Bcb9_0(.din(w_dff_B_Q4ztJBHL6_0),.dout(w_dff_B_SmBl1Bcb9_0),.clk(gclk));
	jdff dff_B_hFgz3um19_0(.din(w_dff_B_SmBl1Bcb9_0),.dout(w_dff_B_hFgz3um19_0),.clk(gclk));
	jdff dff_B_tOH1vVKL3_0(.din(w_dff_B_hFgz3um19_0),.dout(w_dff_B_tOH1vVKL3_0),.clk(gclk));
	jdff dff_B_5Ws8UyBA0_0(.din(w_dff_B_tOH1vVKL3_0),.dout(w_dff_B_5Ws8UyBA0_0),.clk(gclk));
	jdff dff_B_HszMZe0m8_0(.din(w_dff_B_5Ws8UyBA0_0),.dout(w_dff_B_HszMZe0m8_0),.clk(gclk));
	jdff dff_B_MVLtSCjV3_0(.din(w_dff_B_HszMZe0m8_0),.dout(w_dff_B_MVLtSCjV3_0),.clk(gclk));
	jdff dff_B_bOnyNOFe7_0(.din(w_dff_B_MVLtSCjV3_0),.dout(w_dff_B_bOnyNOFe7_0),.clk(gclk));
	jdff dff_B_fkoJ5Jjw0_0(.din(w_dff_B_bOnyNOFe7_0),.dout(w_dff_B_fkoJ5Jjw0_0),.clk(gclk));
	jdff dff_B_Q90IWg9Q2_0(.din(w_dff_B_fkoJ5Jjw0_0),.dout(w_dff_B_Q90IWg9Q2_0),.clk(gclk));
	jdff dff_B_KN1fh3TJ9_0(.din(w_dff_B_Q90IWg9Q2_0),.dout(w_dff_B_KN1fh3TJ9_0),.clk(gclk));
	jdff dff_B_rqRohDcD8_0(.din(w_dff_B_KN1fh3TJ9_0),.dout(w_dff_B_rqRohDcD8_0),.clk(gclk));
	jdff dff_B_aH8b8GyH8_0(.din(w_dff_B_rqRohDcD8_0),.dout(w_dff_B_aH8b8GyH8_0),.clk(gclk));
	jdff dff_B_qrJMhkEn0_0(.din(w_dff_B_aH8b8GyH8_0),.dout(w_dff_B_qrJMhkEn0_0),.clk(gclk));
	jdff dff_B_gpbDAU8f9_0(.din(w_dff_B_qrJMhkEn0_0),.dout(w_dff_B_gpbDAU8f9_0),.clk(gclk));
	jdff dff_B_rPBKxsxN2_0(.din(w_dff_B_gpbDAU8f9_0),.dout(w_dff_B_rPBKxsxN2_0),.clk(gclk));
	jdff dff_B_MjESDd3Q7_0(.din(w_dff_B_rPBKxsxN2_0),.dout(w_dff_B_MjESDd3Q7_0),.clk(gclk));
	jdff dff_B_RycHrpEV1_0(.din(w_dff_B_MjESDd3Q7_0),.dout(w_dff_B_RycHrpEV1_0),.clk(gclk));
	jdff dff_B_nhS8BPsd1_0(.din(w_dff_B_RycHrpEV1_0),.dout(w_dff_B_nhS8BPsd1_0),.clk(gclk));
	jdff dff_B_ZIVdhz7i0_0(.din(w_dff_B_nhS8BPsd1_0),.dout(w_dff_B_ZIVdhz7i0_0),.clk(gclk));
	jdff dff_B_vjqSo6t65_0(.din(w_dff_B_ZIVdhz7i0_0),.dout(w_dff_B_vjqSo6t65_0),.clk(gclk));
	jdff dff_B_v4lwbTeb6_0(.din(w_dff_B_vjqSo6t65_0),.dout(w_dff_B_v4lwbTeb6_0),.clk(gclk));
	jdff dff_B_xXxxeBEB6_0(.din(w_dff_B_v4lwbTeb6_0),.dout(w_dff_B_xXxxeBEB6_0),.clk(gclk));
	jdff dff_B_xX9ZufBE2_0(.din(w_dff_B_xXxxeBEB6_0),.dout(w_dff_B_xX9ZufBE2_0),.clk(gclk));
	jdff dff_B_WYln5OOG2_0(.din(w_dff_B_xX9ZufBE2_0),.dout(w_dff_B_WYln5OOG2_0),.clk(gclk));
	jdff dff_B_TQay20PG3_0(.din(w_dff_B_WYln5OOG2_0),.dout(w_dff_B_TQay20PG3_0),.clk(gclk));
	jdff dff_B_9EfsfU6D7_0(.din(w_dff_B_TQay20PG3_0),.dout(w_dff_B_9EfsfU6D7_0),.clk(gclk));
	jdff dff_B_bEE8t4SK3_0(.din(w_dff_B_9EfsfU6D7_0),.dout(w_dff_B_bEE8t4SK3_0),.clk(gclk));
	jdff dff_B_vWmN97LW1_0(.din(w_dff_B_bEE8t4SK3_0),.dout(w_dff_B_vWmN97LW1_0),.clk(gclk));
	jdff dff_B_m5khuecM8_0(.din(w_dff_B_vWmN97LW1_0),.dout(w_dff_B_m5khuecM8_0),.clk(gclk));
	jdff dff_B_shrIfdo19_0(.din(w_dff_B_m5khuecM8_0),.dout(w_dff_B_shrIfdo19_0),.clk(gclk));
	jdff dff_B_Q7YSl3iw1_0(.din(w_dff_B_shrIfdo19_0),.dout(w_dff_B_Q7YSl3iw1_0),.clk(gclk));
	jdff dff_B_m0afCjyx2_0(.din(w_dff_B_Q7YSl3iw1_0),.dout(w_dff_B_m0afCjyx2_0),.clk(gclk));
	jdff dff_B_s8DUX3p31_0(.din(w_dff_B_m0afCjyx2_0),.dout(w_dff_B_s8DUX3p31_0),.clk(gclk));
	jdff dff_B_eVwcYOHQ0_0(.din(w_dff_B_s8DUX3p31_0),.dout(w_dff_B_eVwcYOHQ0_0),.clk(gclk));
	jdff dff_B_sfgFyjIt5_0(.din(w_dff_B_eVwcYOHQ0_0),.dout(w_dff_B_sfgFyjIt5_0),.clk(gclk));
	jdff dff_B_LhS3JG1z7_0(.din(w_dff_B_sfgFyjIt5_0),.dout(w_dff_B_LhS3JG1z7_0),.clk(gclk));
	jdff dff_B_bSNws27A1_0(.din(w_dff_B_LhS3JG1z7_0),.dout(w_dff_B_bSNws27A1_0),.clk(gclk));
	jdff dff_B_11pDVKuv4_0(.din(w_dff_B_bSNws27A1_0),.dout(w_dff_B_11pDVKuv4_0),.clk(gclk));
	jdff dff_B_wV4uZ5Sm8_0(.din(w_dff_B_11pDVKuv4_0),.dout(w_dff_B_wV4uZ5Sm8_0),.clk(gclk));
	jdff dff_B_oV9dxKqX1_0(.din(w_dff_B_wV4uZ5Sm8_0),.dout(w_dff_B_oV9dxKqX1_0),.clk(gclk));
	jdff dff_B_VBE0HBhG1_0(.din(w_dff_B_oV9dxKqX1_0),.dout(w_dff_B_VBE0HBhG1_0),.clk(gclk));
	jdff dff_B_6fngLBZU7_0(.din(w_dff_B_VBE0HBhG1_0),.dout(w_dff_B_6fngLBZU7_0),.clk(gclk));
	jdff dff_B_VQwpoh080_0(.din(w_dff_B_6fngLBZU7_0),.dout(w_dff_B_VQwpoh080_0),.clk(gclk));
	jdff dff_B_YEKvAFMu1_0(.din(w_dff_B_VQwpoh080_0),.dout(w_dff_B_YEKvAFMu1_0),.clk(gclk));
	jdff dff_B_cbIx5wA74_0(.din(w_dff_B_YEKvAFMu1_0),.dout(w_dff_B_cbIx5wA74_0),.clk(gclk));
	jdff dff_B_t0Hsi3QP9_0(.din(w_dff_B_cbIx5wA74_0),.dout(w_dff_B_t0Hsi3QP9_0),.clk(gclk));
	jdff dff_B_eJSab3Vq4_0(.din(w_dff_B_t0Hsi3QP9_0),.dout(w_dff_B_eJSab3Vq4_0),.clk(gclk));
	jdff dff_B_rie5fYW03_0(.din(w_dff_B_eJSab3Vq4_0),.dout(w_dff_B_rie5fYW03_0),.clk(gclk));
	jdff dff_B_vmrkeYnu7_0(.din(w_dff_B_rie5fYW03_0),.dout(w_dff_B_vmrkeYnu7_0),.clk(gclk));
	jdff dff_B_2oe3zhVW3_0(.din(w_dff_B_vmrkeYnu7_0),.dout(w_dff_B_2oe3zhVW3_0),.clk(gclk));
	jdff dff_B_DLgEEcHe4_0(.din(w_dff_B_2oe3zhVW3_0),.dout(w_dff_B_DLgEEcHe4_0),.clk(gclk));
	jdff dff_B_Wgfequ1T0_0(.din(w_dff_B_DLgEEcHe4_0),.dout(w_dff_B_Wgfequ1T0_0),.clk(gclk));
	jdff dff_B_gtK7CO3B1_0(.din(w_dff_B_Wgfequ1T0_0),.dout(w_dff_B_gtK7CO3B1_0),.clk(gclk));
	jdff dff_B_freIDPdd8_0(.din(w_dff_B_gtK7CO3B1_0),.dout(w_dff_B_freIDPdd8_0),.clk(gclk));
	jdff dff_B_bKzCqqpN1_0(.din(w_dff_B_freIDPdd8_0),.dout(w_dff_B_bKzCqqpN1_0),.clk(gclk));
	jdff dff_B_MAeA0RML4_0(.din(w_dff_B_bKzCqqpN1_0),.dout(w_dff_B_MAeA0RML4_0),.clk(gclk));
	jdff dff_B_YQAMhp5n0_0(.din(w_dff_B_MAeA0RML4_0),.dout(w_dff_B_YQAMhp5n0_0),.clk(gclk));
	jdff dff_B_wapMKsOJ8_0(.din(w_dff_B_YQAMhp5n0_0),.dout(w_dff_B_wapMKsOJ8_0),.clk(gclk));
	jdff dff_B_Lo3ItOgO2_0(.din(w_dff_B_wapMKsOJ8_0),.dout(w_dff_B_Lo3ItOgO2_0),.clk(gclk));
	jdff dff_B_pXkKd7Kz1_0(.din(w_dff_B_Lo3ItOgO2_0),.dout(w_dff_B_pXkKd7Kz1_0),.clk(gclk));
	jdff dff_B_b5IQTnp33_0(.din(w_dff_B_pXkKd7Kz1_0),.dout(w_dff_B_b5IQTnp33_0),.clk(gclk));
	jdff dff_B_D9rd5KXP6_0(.din(w_dff_B_b5IQTnp33_0),.dout(w_dff_B_D9rd5KXP6_0),.clk(gclk));
	jdff dff_B_lkMRwUoy4_0(.din(w_dff_B_D9rd5KXP6_0),.dout(w_dff_B_lkMRwUoy4_0),.clk(gclk));
	jdff dff_B_UOZ77J6s6_0(.din(w_dff_B_lkMRwUoy4_0),.dout(w_dff_B_UOZ77J6s6_0),.clk(gclk));
	jdff dff_B_4dmaQakO5_0(.din(w_dff_B_UOZ77J6s6_0),.dout(w_dff_B_4dmaQakO5_0),.clk(gclk));
	jdff dff_B_HfHV0p9z3_0(.din(w_dff_B_4dmaQakO5_0),.dout(w_dff_B_HfHV0p9z3_0),.clk(gclk));
	jdff dff_B_2h1MaLiM2_0(.din(w_dff_B_HfHV0p9z3_0),.dout(w_dff_B_2h1MaLiM2_0),.clk(gclk));
	jdff dff_B_RU2aNEET8_0(.din(w_dff_B_2h1MaLiM2_0),.dout(w_dff_B_RU2aNEET8_0),.clk(gclk));
	jdff dff_B_l5c4V3iN3_0(.din(w_dff_B_RU2aNEET8_0),.dout(w_dff_B_l5c4V3iN3_0),.clk(gclk));
	jdff dff_B_w1tZACVk8_0(.din(w_dff_B_l5c4V3iN3_0),.dout(w_dff_B_w1tZACVk8_0),.clk(gclk));
	jdff dff_B_Fl7D7wAm4_0(.din(w_dff_B_w1tZACVk8_0),.dout(w_dff_B_Fl7D7wAm4_0),.clk(gclk));
	jdff dff_B_pshJjRMi3_0(.din(w_dff_B_Fl7D7wAm4_0),.dout(w_dff_B_pshJjRMi3_0),.clk(gclk));
	jdff dff_B_aQv0bGNk7_0(.din(w_dff_B_pshJjRMi3_0),.dout(w_dff_B_aQv0bGNk7_0),.clk(gclk));
	jdff dff_B_ae7OEHZp0_0(.din(w_dff_B_aQv0bGNk7_0),.dout(w_dff_B_ae7OEHZp0_0),.clk(gclk));
	jdff dff_B_kvtzmL0r4_0(.din(w_dff_B_ae7OEHZp0_0),.dout(w_dff_B_kvtzmL0r4_0),.clk(gclk));
	jdff dff_B_oDI3aSF29_0(.din(w_dff_B_kvtzmL0r4_0),.dout(w_dff_B_oDI3aSF29_0),.clk(gclk));
	jdff dff_B_mqkx78xk3_0(.din(w_dff_B_oDI3aSF29_0),.dout(w_dff_B_mqkx78xk3_0),.clk(gclk));
	jdff dff_B_0seXyGFE9_0(.din(w_dff_B_mqkx78xk3_0),.dout(w_dff_B_0seXyGFE9_0),.clk(gclk));
	jdff dff_B_lR7n1kre2_0(.din(w_dff_B_0seXyGFE9_0),.dout(w_dff_B_lR7n1kre2_0),.clk(gclk));
	jdff dff_B_q9sw8fpB1_0(.din(w_dff_B_lR7n1kre2_0),.dout(w_dff_B_q9sw8fpB1_0),.clk(gclk));
	jdff dff_B_pDiftYiS6_0(.din(w_dff_B_q9sw8fpB1_0),.dout(w_dff_B_pDiftYiS6_0),.clk(gclk));
	jdff dff_B_4Mik9kMM2_0(.din(w_dff_B_pDiftYiS6_0),.dout(w_dff_B_4Mik9kMM2_0),.clk(gclk));
	jdff dff_B_2Gw5om041_0(.din(w_dff_B_4Mik9kMM2_0),.dout(w_dff_B_2Gw5om041_0),.clk(gclk));
	jdff dff_B_0xMzr56d5_0(.din(w_dff_B_2Gw5om041_0),.dout(w_dff_B_0xMzr56d5_0),.clk(gclk));
	jdff dff_B_Bc3aEgHa3_0(.din(w_dff_B_0xMzr56d5_0),.dout(w_dff_B_Bc3aEgHa3_0),.clk(gclk));
	jdff dff_B_Jr5rAzQK1_0(.din(w_dff_B_Bc3aEgHa3_0),.dout(w_dff_B_Jr5rAzQK1_0),.clk(gclk));
	jdff dff_B_Z0Qj2PC29_0(.din(w_dff_B_Jr5rAzQK1_0),.dout(w_dff_B_Z0Qj2PC29_0),.clk(gclk));
	jdff dff_B_5Iw6WGuZ5_0(.din(w_dff_B_Z0Qj2PC29_0),.dout(w_dff_B_5Iw6WGuZ5_0),.clk(gclk));
	jdff dff_B_M4XffYyu2_0(.din(w_dff_B_5Iw6WGuZ5_0),.dout(w_dff_B_M4XffYyu2_0),.clk(gclk));
	jdff dff_B_sOSJEZFe8_0(.din(w_dff_B_M4XffYyu2_0),.dout(w_dff_B_sOSJEZFe8_0),.clk(gclk));
	jdff dff_B_Fiym9kQc9_0(.din(w_dff_B_sOSJEZFe8_0),.dout(w_dff_B_Fiym9kQc9_0),.clk(gclk));
	jdff dff_B_4gkEbQSM5_0(.din(w_dff_B_Fiym9kQc9_0),.dout(w_dff_B_4gkEbQSM5_0),.clk(gclk));
	jdff dff_B_ekHpHopO6_0(.din(w_dff_B_4gkEbQSM5_0),.dout(w_dff_B_ekHpHopO6_0),.clk(gclk));
	jdff dff_B_t9WZNTWu4_0(.din(w_dff_B_ekHpHopO6_0),.dout(w_dff_B_t9WZNTWu4_0),.clk(gclk));
	jdff dff_B_tAY2Yj6h5_0(.din(w_dff_B_t9WZNTWu4_0),.dout(w_dff_B_tAY2Yj6h5_0),.clk(gclk));
	jdff dff_B_EYJkHRuW1_0(.din(w_dff_B_tAY2Yj6h5_0),.dout(w_dff_B_EYJkHRuW1_0),.clk(gclk));
	jdff dff_B_ihbYCldo3_0(.din(w_dff_B_EYJkHRuW1_0),.dout(w_dff_B_ihbYCldo3_0),.clk(gclk));
	jdff dff_B_MCq281UY6_1(.din(n1068),.dout(w_dff_B_MCq281UY6_1),.clk(gclk));
	jdff dff_B_1ADqnZNQ4_1(.din(w_dff_B_MCq281UY6_1),.dout(w_dff_B_1ADqnZNQ4_1),.clk(gclk));
	jdff dff_B_7t9HJ7sx2_1(.din(w_dff_B_1ADqnZNQ4_1),.dout(w_dff_B_7t9HJ7sx2_1),.clk(gclk));
	jdff dff_B_tkwL7lN16_1(.din(w_dff_B_7t9HJ7sx2_1),.dout(w_dff_B_tkwL7lN16_1),.clk(gclk));
	jdff dff_B_LS2fiSKH2_1(.din(w_dff_B_tkwL7lN16_1),.dout(w_dff_B_LS2fiSKH2_1),.clk(gclk));
	jdff dff_B_TcM1PmAn2_1(.din(w_dff_B_LS2fiSKH2_1),.dout(w_dff_B_TcM1PmAn2_1),.clk(gclk));
	jdff dff_B_4uTXGvEq7_1(.din(w_dff_B_TcM1PmAn2_1),.dout(w_dff_B_4uTXGvEq7_1),.clk(gclk));
	jdff dff_B_dWw8OsXj0_1(.din(w_dff_B_4uTXGvEq7_1),.dout(w_dff_B_dWw8OsXj0_1),.clk(gclk));
	jdff dff_B_JbviCirz7_1(.din(w_dff_B_dWw8OsXj0_1),.dout(w_dff_B_JbviCirz7_1),.clk(gclk));
	jdff dff_B_aYarJ7CU1_1(.din(w_dff_B_JbviCirz7_1),.dout(w_dff_B_aYarJ7CU1_1),.clk(gclk));
	jdff dff_B_FSEIA4MW4_1(.din(w_dff_B_aYarJ7CU1_1),.dout(w_dff_B_FSEIA4MW4_1),.clk(gclk));
	jdff dff_B_aoJppHH29_1(.din(w_dff_B_FSEIA4MW4_1),.dout(w_dff_B_aoJppHH29_1),.clk(gclk));
	jdff dff_B_QLFHExor6_1(.din(w_dff_B_aoJppHH29_1),.dout(w_dff_B_QLFHExor6_1),.clk(gclk));
	jdff dff_B_zFQXqWL58_1(.din(w_dff_B_QLFHExor6_1),.dout(w_dff_B_zFQXqWL58_1),.clk(gclk));
	jdff dff_B_7QDYzYvG2_1(.din(w_dff_B_zFQXqWL58_1),.dout(w_dff_B_7QDYzYvG2_1),.clk(gclk));
	jdff dff_B_Mp43LeOg9_1(.din(w_dff_B_7QDYzYvG2_1),.dout(w_dff_B_Mp43LeOg9_1),.clk(gclk));
	jdff dff_B_F1SHhpCQ7_1(.din(w_dff_B_Mp43LeOg9_1),.dout(w_dff_B_F1SHhpCQ7_1),.clk(gclk));
	jdff dff_B_VQv64JSq9_1(.din(w_dff_B_F1SHhpCQ7_1),.dout(w_dff_B_VQv64JSq9_1),.clk(gclk));
	jdff dff_B_3wJaWl3d6_1(.din(w_dff_B_VQv64JSq9_1),.dout(w_dff_B_3wJaWl3d6_1),.clk(gclk));
	jdff dff_B_B1q10AOM0_1(.din(w_dff_B_3wJaWl3d6_1),.dout(w_dff_B_B1q10AOM0_1),.clk(gclk));
	jdff dff_B_clg6xez41_1(.din(w_dff_B_B1q10AOM0_1),.dout(w_dff_B_clg6xez41_1),.clk(gclk));
	jdff dff_B_xDt5lsgj7_1(.din(w_dff_B_clg6xez41_1),.dout(w_dff_B_xDt5lsgj7_1),.clk(gclk));
	jdff dff_B_8pKmFt6G3_1(.din(w_dff_B_xDt5lsgj7_1),.dout(w_dff_B_8pKmFt6G3_1),.clk(gclk));
	jdff dff_B_kmhcdLiB8_1(.din(w_dff_B_8pKmFt6G3_1),.dout(w_dff_B_kmhcdLiB8_1),.clk(gclk));
	jdff dff_B_PyKYIiaX0_1(.din(w_dff_B_kmhcdLiB8_1),.dout(w_dff_B_PyKYIiaX0_1),.clk(gclk));
	jdff dff_B_d0BVUFZ00_1(.din(w_dff_B_PyKYIiaX0_1),.dout(w_dff_B_d0BVUFZ00_1),.clk(gclk));
	jdff dff_B_JZeDEizN3_1(.din(w_dff_B_d0BVUFZ00_1),.dout(w_dff_B_JZeDEizN3_1),.clk(gclk));
	jdff dff_B_6V9OAOSy1_1(.din(w_dff_B_JZeDEizN3_1),.dout(w_dff_B_6V9OAOSy1_1),.clk(gclk));
	jdff dff_B_AOGEX5kr0_1(.din(w_dff_B_6V9OAOSy1_1),.dout(w_dff_B_AOGEX5kr0_1),.clk(gclk));
	jdff dff_B_cl58WqLZ2_1(.din(w_dff_B_AOGEX5kr0_1),.dout(w_dff_B_cl58WqLZ2_1),.clk(gclk));
	jdff dff_B_bzBy4IcZ8_1(.din(w_dff_B_cl58WqLZ2_1),.dout(w_dff_B_bzBy4IcZ8_1),.clk(gclk));
	jdff dff_B_D3X6rZeS0_1(.din(w_dff_B_bzBy4IcZ8_1),.dout(w_dff_B_D3X6rZeS0_1),.clk(gclk));
	jdff dff_B_cAPbxwEv0_1(.din(w_dff_B_D3X6rZeS0_1),.dout(w_dff_B_cAPbxwEv0_1),.clk(gclk));
	jdff dff_B_rhVk8whC4_1(.din(w_dff_B_cAPbxwEv0_1),.dout(w_dff_B_rhVk8whC4_1),.clk(gclk));
	jdff dff_B_mhBkypJF1_1(.din(w_dff_B_rhVk8whC4_1),.dout(w_dff_B_mhBkypJF1_1),.clk(gclk));
	jdff dff_B_rTK8PBFd5_1(.din(w_dff_B_mhBkypJF1_1),.dout(w_dff_B_rTK8PBFd5_1),.clk(gclk));
	jdff dff_B_8YIYuS5L0_1(.din(w_dff_B_rTK8PBFd5_1),.dout(w_dff_B_8YIYuS5L0_1),.clk(gclk));
	jdff dff_B_d7sc9C9q5_1(.din(w_dff_B_8YIYuS5L0_1),.dout(w_dff_B_d7sc9C9q5_1),.clk(gclk));
	jdff dff_B_AEfYuPVR1_1(.din(w_dff_B_d7sc9C9q5_1),.dout(w_dff_B_AEfYuPVR1_1),.clk(gclk));
	jdff dff_B_1mAkaiIM9_1(.din(w_dff_B_AEfYuPVR1_1),.dout(w_dff_B_1mAkaiIM9_1),.clk(gclk));
	jdff dff_B_1dwby9fs1_1(.din(w_dff_B_1mAkaiIM9_1),.dout(w_dff_B_1dwby9fs1_1),.clk(gclk));
	jdff dff_B_6zeCK66Z0_1(.din(w_dff_B_1dwby9fs1_1),.dout(w_dff_B_6zeCK66Z0_1),.clk(gclk));
	jdff dff_B_ScERKzgl5_1(.din(w_dff_B_6zeCK66Z0_1),.dout(w_dff_B_ScERKzgl5_1),.clk(gclk));
	jdff dff_B_vIYE3bUe5_1(.din(w_dff_B_ScERKzgl5_1),.dout(w_dff_B_vIYE3bUe5_1),.clk(gclk));
	jdff dff_B_kIQ57ik54_1(.din(w_dff_B_vIYE3bUe5_1),.dout(w_dff_B_kIQ57ik54_1),.clk(gclk));
	jdff dff_B_hVvEonaG5_1(.din(w_dff_B_kIQ57ik54_1),.dout(w_dff_B_hVvEonaG5_1),.clk(gclk));
	jdff dff_B_PcC3HCUZ7_1(.din(w_dff_B_hVvEonaG5_1),.dout(w_dff_B_PcC3HCUZ7_1),.clk(gclk));
	jdff dff_B_uAN9qSbH8_1(.din(w_dff_B_PcC3HCUZ7_1),.dout(w_dff_B_uAN9qSbH8_1),.clk(gclk));
	jdff dff_B_v2YTIsda9_1(.din(w_dff_B_uAN9qSbH8_1),.dout(w_dff_B_v2YTIsda9_1),.clk(gclk));
	jdff dff_B_iAVuv22D1_1(.din(w_dff_B_v2YTIsda9_1),.dout(w_dff_B_iAVuv22D1_1),.clk(gclk));
	jdff dff_B_d1gWu6fs3_1(.din(w_dff_B_iAVuv22D1_1),.dout(w_dff_B_d1gWu6fs3_1),.clk(gclk));
	jdff dff_B_vpO54gNf1_1(.din(w_dff_B_d1gWu6fs3_1),.dout(w_dff_B_vpO54gNf1_1),.clk(gclk));
	jdff dff_B_2e7ZQvDb0_1(.din(w_dff_B_vpO54gNf1_1),.dout(w_dff_B_2e7ZQvDb0_1),.clk(gclk));
	jdff dff_B_mx0LxQZu7_1(.din(w_dff_B_2e7ZQvDb0_1),.dout(w_dff_B_mx0LxQZu7_1),.clk(gclk));
	jdff dff_B_0Ugtxr3R0_1(.din(w_dff_B_mx0LxQZu7_1),.dout(w_dff_B_0Ugtxr3R0_1),.clk(gclk));
	jdff dff_B_1WfTxDNM8_1(.din(w_dff_B_0Ugtxr3R0_1),.dout(w_dff_B_1WfTxDNM8_1),.clk(gclk));
	jdff dff_B_5HYuIW3Y0_1(.din(w_dff_B_1WfTxDNM8_1),.dout(w_dff_B_5HYuIW3Y0_1),.clk(gclk));
	jdff dff_B_l6t5TALj6_1(.din(w_dff_B_5HYuIW3Y0_1),.dout(w_dff_B_l6t5TALj6_1),.clk(gclk));
	jdff dff_B_GzfykcJo7_1(.din(w_dff_B_l6t5TALj6_1),.dout(w_dff_B_GzfykcJo7_1),.clk(gclk));
	jdff dff_B_JGt70JuB2_1(.din(w_dff_B_GzfykcJo7_1),.dout(w_dff_B_JGt70JuB2_1),.clk(gclk));
	jdff dff_B_AdA6CQ5C8_1(.din(w_dff_B_JGt70JuB2_1),.dout(w_dff_B_AdA6CQ5C8_1),.clk(gclk));
	jdff dff_B_ykauX71l3_1(.din(w_dff_B_AdA6CQ5C8_1),.dout(w_dff_B_ykauX71l3_1),.clk(gclk));
	jdff dff_B_A1KMzE375_1(.din(w_dff_B_ykauX71l3_1),.dout(w_dff_B_A1KMzE375_1),.clk(gclk));
	jdff dff_B_C60JWqCY9_1(.din(w_dff_B_A1KMzE375_1),.dout(w_dff_B_C60JWqCY9_1),.clk(gclk));
	jdff dff_B_guAiUpl23_1(.din(w_dff_B_C60JWqCY9_1),.dout(w_dff_B_guAiUpl23_1),.clk(gclk));
	jdff dff_B_Qgnwv9a00_1(.din(w_dff_B_guAiUpl23_1),.dout(w_dff_B_Qgnwv9a00_1),.clk(gclk));
	jdff dff_B_wp7I8PDh1_1(.din(w_dff_B_Qgnwv9a00_1),.dout(w_dff_B_wp7I8PDh1_1),.clk(gclk));
	jdff dff_B_PGq0nBXZ0_1(.din(w_dff_B_wp7I8PDh1_1),.dout(w_dff_B_PGq0nBXZ0_1),.clk(gclk));
	jdff dff_B_Jt5JYBMu5_1(.din(w_dff_B_PGq0nBXZ0_1),.dout(w_dff_B_Jt5JYBMu5_1),.clk(gclk));
	jdff dff_B_aVZHfeaP9_1(.din(w_dff_B_Jt5JYBMu5_1),.dout(w_dff_B_aVZHfeaP9_1),.clk(gclk));
	jdff dff_B_uT9UZBIX0_1(.din(w_dff_B_aVZHfeaP9_1),.dout(w_dff_B_uT9UZBIX0_1),.clk(gclk));
	jdff dff_B_L5Bx4XHE3_1(.din(w_dff_B_uT9UZBIX0_1),.dout(w_dff_B_L5Bx4XHE3_1),.clk(gclk));
	jdff dff_B_T9MpUjrF1_1(.din(w_dff_B_L5Bx4XHE3_1),.dout(w_dff_B_T9MpUjrF1_1),.clk(gclk));
	jdff dff_B_btAq2qi01_1(.din(w_dff_B_T9MpUjrF1_1),.dout(w_dff_B_btAq2qi01_1),.clk(gclk));
	jdff dff_B_nyAcjzIt9_1(.din(w_dff_B_btAq2qi01_1),.dout(w_dff_B_nyAcjzIt9_1),.clk(gclk));
	jdff dff_B_EBQj51um8_1(.din(w_dff_B_nyAcjzIt9_1),.dout(w_dff_B_EBQj51um8_1),.clk(gclk));
	jdff dff_B_eoCRFH6e6_1(.din(w_dff_B_EBQj51um8_1),.dout(w_dff_B_eoCRFH6e6_1),.clk(gclk));
	jdff dff_B_QM9cp9qm2_1(.din(w_dff_B_eoCRFH6e6_1),.dout(w_dff_B_QM9cp9qm2_1),.clk(gclk));
	jdff dff_B_MSkuuZ4p9_1(.din(w_dff_B_QM9cp9qm2_1),.dout(w_dff_B_MSkuuZ4p9_1),.clk(gclk));
	jdff dff_B_crHZNiH82_1(.din(w_dff_B_MSkuuZ4p9_1),.dout(w_dff_B_crHZNiH82_1),.clk(gclk));
	jdff dff_B_Y3HQ5Wur3_1(.din(w_dff_B_crHZNiH82_1),.dout(w_dff_B_Y3HQ5Wur3_1),.clk(gclk));
	jdff dff_B_0SguyIlg0_1(.din(w_dff_B_Y3HQ5Wur3_1),.dout(w_dff_B_0SguyIlg0_1),.clk(gclk));
	jdff dff_B_06qyFdKf7_1(.din(w_dff_B_0SguyIlg0_1),.dout(w_dff_B_06qyFdKf7_1),.clk(gclk));
	jdff dff_B_6xfsC01k5_1(.din(w_dff_B_06qyFdKf7_1),.dout(w_dff_B_6xfsC01k5_1),.clk(gclk));
	jdff dff_B_VBOUQcis4_1(.din(w_dff_B_6xfsC01k5_1),.dout(w_dff_B_VBOUQcis4_1),.clk(gclk));
	jdff dff_B_crKgyBc98_1(.din(w_dff_B_VBOUQcis4_1),.dout(w_dff_B_crKgyBc98_1),.clk(gclk));
	jdff dff_B_mCFwTzhf3_1(.din(w_dff_B_crKgyBc98_1),.dout(w_dff_B_mCFwTzhf3_1),.clk(gclk));
	jdff dff_B_XuCysnJ71_1(.din(w_dff_B_mCFwTzhf3_1),.dout(w_dff_B_XuCysnJ71_1),.clk(gclk));
	jdff dff_B_iLbXeH9p5_1(.din(w_dff_B_XuCysnJ71_1),.dout(w_dff_B_iLbXeH9p5_1),.clk(gclk));
	jdff dff_B_FwauJUrI0_1(.din(w_dff_B_iLbXeH9p5_1),.dout(w_dff_B_FwauJUrI0_1),.clk(gclk));
	jdff dff_B_iB5XbIjn2_1(.din(w_dff_B_FwauJUrI0_1),.dout(w_dff_B_iB5XbIjn2_1),.clk(gclk));
	jdff dff_B_lSJMyNrK1_1(.din(w_dff_B_iB5XbIjn2_1),.dout(w_dff_B_lSJMyNrK1_1),.clk(gclk));
	jdff dff_B_WsG7DlL11_1(.din(w_dff_B_lSJMyNrK1_1),.dout(w_dff_B_WsG7DlL11_1),.clk(gclk));
	jdff dff_B_VUxvO5sy1_1(.din(w_dff_B_WsG7DlL11_1),.dout(w_dff_B_VUxvO5sy1_1),.clk(gclk));
	jdff dff_B_Eypraqwc0_1(.din(w_dff_B_VUxvO5sy1_1),.dout(w_dff_B_Eypraqwc0_1),.clk(gclk));
	jdff dff_B_66VSaaGL4_1(.din(w_dff_B_Eypraqwc0_1),.dout(w_dff_B_66VSaaGL4_1),.clk(gclk));
	jdff dff_B_cAtCcmj90_1(.din(w_dff_B_66VSaaGL4_1),.dout(w_dff_B_cAtCcmj90_1),.clk(gclk));
	jdff dff_B_Lh9aLFRP8_1(.din(w_dff_B_cAtCcmj90_1),.dout(w_dff_B_Lh9aLFRP8_1),.clk(gclk));
	jdff dff_B_Hh59ncTe1_1(.din(w_dff_B_Lh9aLFRP8_1),.dout(w_dff_B_Hh59ncTe1_1),.clk(gclk));
	jdff dff_B_5KD1EUHe7_1(.din(w_dff_B_Hh59ncTe1_1),.dout(w_dff_B_5KD1EUHe7_1),.clk(gclk));
	jdff dff_B_yRZwIymy7_1(.din(w_dff_B_5KD1EUHe7_1),.dout(w_dff_B_yRZwIymy7_1),.clk(gclk));
	jdff dff_B_Gpc3FdUr1_1(.din(w_dff_B_yRZwIymy7_1),.dout(w_dff_B_Gpc3FdUr1_1),.clk(gclk));
	jdff dff_B_ZdtaE59g7_1(.din(w_dff_B_Gpc3FdUr1_1),.dout(w_dff_B_ZdtaE59g7_1),.clk(gclk));
	jdff dff_B_uJ1qSNMa2_1(.din(w_dff_B_ZdtaE59g7_1),.dout(w_dff_B_uJ1qSNMa2_1),.clk(gclk));
	jdff dff_B_Ipw2d4wE4_1(.din(w_dff_B_uJ1qSNMa2_1),.dout(w_dff_B_Ipw2d4wE4_1),.clk(gclk));
	jdff dff_B_1SY2ypEI3_1(.din(w_dff_B_Ipw2d4wE4_1),.dout(w_dff_B_1SY2ypEI3_1),.clk(gclk));
	jdff dff_B_nUFQeGhJ8_1(.din(w_dff_B_1SY2ypEI3_1),.dout(w_dff_B_nUFQeGhJ8_1),.clk(gclk));
	jdff dff_B_HllRApmp6_1(.din(w_dff_B_nUFQeGhJ8_1),.dout(w_dff_B_HllRApmp6_1),.clk(gclk));
	jdff dff_B_Th2DnWdp4_1(.din(w_dff_B_HllRApmp6_1),.dout(w_dff_B_Th2DnWdp4_1),.clk(gclk));
	jdff dff_B_ZsBjt1bw8_1(.din(w_dff_B_Th2DnWdp4_1),.dout(w_dff_B_ZsBjt1bw8_1),.clk(gclk));
	jdff dff_B_vDC3FAL36_1(.din(w_dff_B_ZsBjt1bw8_1),.dout(w_dff_B_vDC3FAL36_1),.clk(gclk));
	jdff dff_B_dBiYiSsG8_1(.din(w_dff_B_vDC3FAL36_1),.dout(w_dff_B_dBiYiSsG8_1),.clk(gclk));
	jdff dff_B_N3sp0qOL9_1(.din(w_dff_B_dBiYiSsG8_1),.dout(w_dff_B_N3sp0qOL9_1),.clk(gclk));
	jdff dff_B_SjyTVPLT6_1(.din(w_dff_B_N3sp0qOL9_1),.dout(w_dff_B_SjyTVPLT6_1),.clk(gclk));
	jdff dff_B_rg3QJQk22_0(.din(n1069),.dout(w_dff_B_rg3QJQk22_0),.clk(gclk));
	jdff dff_B_Nx6dgmj31_0(.din(w_dff_B_rg3QJQk22_0),.dout(w_dff_B_Nx6dgmj31_0),.clk(gclk));
	jdff dff_B_KysPl3gz9_0(.din(w_dff_B_Nx6dgmj31_0),.dout(w_dff_B_KysPl3gz9_0),.clk(gclk));
	jdff dff_B_SeUWHHwM7_0(.din(w_dff_B_KysPl3gz9_0),.dout(w_dff_B_SeUWHHwM7_0),.clk(gclk));
	jdff dff_B_eGxZdXiI3_0(.din(w_dff_B_SeUWHHwM7_0),.dout(w_dff_B_eGxZdXiI3_0),.clk(gclk));
	jdff dff_B_Ep13Dq9T0_0(.din(w_dff_B_eGxZdXiI3_0),.dout(w_dff_B_Ep13Dq9T0_0),.clk(gclk));
	jdff dff_B_ceXWccHN8_0(.din(w_dff_B_Ep13Dq9T0_0),.dout(w_dff_B_ceXWccHN8_0),.clk(gclk));
	jdff dff_B_zj6XrN4j8_0(.din(w_dff_B_ceXWccHN8_0),.dout(w_dff_B_zj6XrN4j8_0),.clk(gclk));
	jdff dff_B_gMo14vJs2_0(.din(w_dff_B_zj6XrN4j8_0),.dout(w_dff_B_gMo14vJs2_0),.clk(gclk));
	jdff dff_B_PDxzq8wM0_0(.din(w_dff_B_gMo14vJs2_0),.dout(w_dff_B_PDxzq8wM0_0),.clk(gclk));
	jdff dff_B_K4PqtKp17_0(.din(w_dff_B_PDxzq8wM0_0),.dout(w_dff_B_K4PqtKp17_0),.clk(gclk));
	jdff dff_B_B7TEkhld6_0(.din(w_dff_B_K4PqtKp17_0),.dout(w_dff_B_B7TEkhld6_0),.clk(gclk));
	jdff dff_B_jcJlavc00_0(.din(w_dff_B_B7TEkhld6_0),.dout(w_dff_B_jcJlavc00_0),.clk(gclk));
	jdff dff_B_NnIjIV0h6_0(.din(w_dff_B_jcJlavc00_0),.dout(w_dff_B_NnIjIV0h6_0),.clk(gclk));
	jdff dff_B_6Fdzq0SK4_0(.din(w_dff_B_NnIjIV0h6_0),.dout(w_dff_B_6Fdzq0SK4_0),.clk(gclk));
	jdff dff_B_l1raEnt12_0(.din(w_dff_B_6Fdzq0SK4_0),.dout(w_dff_B_l1raEnt12_0),.clk(gclk));
	jdff dff_B_aDh62mhu6_0(.din(w_dff_B_l1raEnt12_0),.dout(w_dff_B_aDh62mhu6_0),.clk(gclk));
	jdff dff_B_7Ee6opFT4_0(.din(w_dff_B_aDh62mhu6_0),.dout(w_dff_B_7Ee6opFT4_0),.clk(gclk));
	jdff dff_B_siN5GXkT0_0(.din(w_dff_B_7Ee6opFT4_0),.dout(w_dff_B_siN5GXkT0_0),.clk(gclk));
	jdff dff_B_b6AujLj70_0(.din(w_dff_B_siN5GXkT0_0),.dout(w_dff_B_b6AujLj70_0),.clk(gclk));
	jdff dff_B_kXQa8VgV0_0(.din(w_dff_B_b6AujLj70_0),.dout(w_dff_B_kXQa8VgV0_0),.clk(gclk));
	jdff dff_B_z3JHWaLb1_0(.din(w_dff_B_kXQa8VgV0_0),.dout(w_dff_B_z3JHWaLb1_0),.clk(gclk));
	jdff dff_B_k3kLrxQj5_0(.din(w_dff_B_z3JHWaLb1_0),.dout(w_dff_B_k3kLrxQj5_0),.clk(gclk));
	jdff dff_B_Bwpn8EZg4_0(.din(w_dff_B_k3kLrxQj5_0),.dout(w_dff_B_Bwpn8EZg4_0),.clk(gclk));
	jdff dff_B_c0DkvoDH8_0(.din(w_dff_B_Bwpn8EZg4_0),.dout(w_dff_B_c0DkvoDH8_0),.clk(gclk));
	jdff dff_B_lflksyiR1_0(.din(w_dff_B_c0DkvoDH8_0),.dout(w_dff_B_lflksyiR1_0),.clk(gclk));
	jdff dff_B_U5P7Atke3_0(.din(w_dff_B_lflksyiR1_0),.dout(w_dff_B_U5P7Atke3_0),.clk(gclk));
	jdff dff_B_NjVlTxqN8_0(.din(w_dff_B_U5P7Atke3_0),.dout(w_dff_B_NjVlTxqN8_0),.clk(gclk));
	jdff dff_B_LtIpXpqa0_0(.din(w_dff_B_NjVlTxqN8_0),.dout(w_dff_B_LtIpXpqa0_0),.clk(gclk));
	jdff dff_B_JeA7Omf62_0(.din(w_dff_B_LtIpXpqa0_0),.dout(w_dff_B_JeA7Omf62_0),.clk(gclk));
	jdff dff_B_hkxHifVD3_0(.din(w_dff_B_JeA7Omf62_0),.dout(w_dff_B_hkxHifVD3_0),.clk(gclk));
	jdff dff_B_1InYddIc5_0(.din(w_dff_B_hkxHifVD3_0),.dout(w_dff_B_1InYddIc5_0),.clk(gclk));
	jdff dff_B_YbkFbB3G2_0(.din(w_dff_B_1InYddIc5_0),.dout(w_dff_B_YbkFbB3G2_0),.clk(gclk));
	jdff dff_B_bWMHe5lm3_0(.din(w_dff_B_YbkFbB3G2_0),.dout(w_dff_B_bWMHe5lm3_0),.clk(gclk));
	jdff dff_B_brMV1ppe7_0(.din(w_dff_B_bWMHe5lm3_0),.dout(w_dff_B_brMV1ppe7_0),.clk(gclk));
	jdff dff_B_168MpKru2_0(.din(w_dff_B_brMV1ppe7_0),.dout(w_dff_B_168MpKru2_0),.clk(gclk));
	jdff dff_B_7HhTAQmD7_0(.din(w_dff_B_168MpKru2_0),.dout(w_dff_B_7HhTAQmD7_0),.clk(gclk));
	jdff dff_B_aMaKUyGa1_0(.din(w_dff_B_7HhTAQmD7_0),.dout(w_dff_B_aMaKUyGa1_0),.clk(gclk));
	jdff dff_B_KYvt7k1M0_0(.din(w_dff_B_aMaKUyGa1_0),.dout(w_dff_B_KYvt7k1M0_0),.clk(gclk));
	jdff dff_B_eDN03dgm5_0(.din(w_dff_B_KYvt7k1M0_0),.dout(w_dff_B_eDN03dgm5_0),.clk(gclk));
	jdff dff_B_5IxD8TV83_0(.din(w_dff_B_eDN03dgm5_0),.dout(w_dff_B_5IxD8TV83_0),.clk(gclk));
	jdff dff_B_dcqs8CCV5_0(.din(w_dff_B_5IxD8TV83_0),.dout(w_dff_B_dcqs8CCV5_0),.clk(gclk));
	jdff dff_B_oDmOby2X9_0(.din(w_dff_B_dcqs8CCV5_0),.dout(w_dff_B_oDmOby2X9_0),.clk(gclk));
	jdff dff_B_c6WqCTZd7_0(.din(w_dff_B_oDmOby2X9_0),.dout(w_dff_B_c6WqCTZd7_0),.clk(gclk));
	jdff dff_B_acMX1Wc62_0(.din(w_dff_B_c6WqCTZd7_0),.dout(w_dff_B_acMX1Wc62_0),.clk(gclk));
	jdff dff_B_6PQFdLeR0_0(.din(w_dff_B_acMX1Wc62_0),.dout(w_dff_B_6PQFdLeR0_0),.clk(gclk));
	jdff dff_B_uhdn1nIl4_0(.din(w_dff_B_6PQFdLeR0_0),.dout(w_dff_B_uhdn1nIl4_0),.clk(gclk));
	jdff dff_B_8LyOA8hz0_0(.din(w_dff_B_uhdn1nIl4_0),.dout(w_dff_B_8LyOA8hz0_0),.clk(gclk));
	jdff dff_B_uNcXXOMv4_0(.din(w_dff_B_8LyOA8hz0_0),.dout(w_dff_B_uNcXXOMv4_0),.clk(gclk));
	jdff dff_B_3J9Fc0WC8_0(.din(w_dff_B_uNcXXOMv4_0),.dout(w_dff_B_3J9Fc0WC8_0),.clk(gclk));
	jdff dff_B_3zEPpAuD4_0(.din(w_dff_B_3J9Fc0WC8_0),.dout(w_dff_B_3zEPpAuD4_0),.clk(gclk));
	jdff dff_B_1k8uGg8o9_0(.din(w_dff_B_3zEPpAuD4_0),.dout(w_dff_B_1k8uGg8o9_0),.clk(gclk));
	jdff dff_B_JmP4pRMn8_0(.din(w_dff_B_1k8uGg8o9_0),.dout(w_dff_B_JmP4pRMn8_0),.clk(gclk));
	jdff dff_B_ue8z7mek9_0(.din(w_dff_B_JmP4pRMn8_0),.dout(w_dff_B_ue8z7mek9_0),.clk(gclk));
	jdff dff_B_ObduV78a6_0(.din(w_dff_B_ue8z7mek9_0),.dout(w_dff_B_ObduV78a6_0),.clk(gclk));
	jdff dff_B_13KbV9xF6_0(.din(w_dff_B_ObduV78a6_0),.dout(w_dff_B_13KbV9xF6_0),.clk(gclk));
	jdff dff_B_Kx3hxUf32_0(.din(w_dff_B_13KbV9xF6_0),.dout(w_dff_B_Kx3hxUf32_0),.clk(gclk));
	jdff dff_B_ZLSlyOH09_0(.din(w_dff_B_Kx3hxUf32_0),.dout(w_dff_B_ZLSlyOH09_0),.clk(gclk));
	jdff dff_B_M2jtz1wW7_0(.din(w_dff_B_ZLSlyOH09_0),.dout(w_dff_B_M2jtz1wW7_0),.clk(gclk));
	jdff dff_B_0Ko6pMOz6_0(.din(w_dff_B_M2jtz1wW7_0),.dout(w_dff_B_0Ko6pMOz6_0),.clk(gclk));
	jdff dff_B_hkrtPrUb0_0(.din(w_dff_B_0Ko6pMOz6_0),.dout(w_dff_B_hkrtPrUb0_0),.clk(gclk));
	jdff dff_B_kL9ZBm5j1_0(.din(w_dff_B_hkrtPrUb0_0),.dout(w_dff_B_kL9ZBm5j1_0),.clk(gclk));
	jdff dff_B_mMhx6LXN6_0(.din(w_dff_B_kL9ZBm5j1_0),.dout(w_dff_B_mMhx6LXN6_0),.clk(gclk));
	jdff dff_B_4bl9Za4H4_0(.din(w_dff_B_mMhx6LXN6_0),.dout(w_dff_B_4bl9Za4H4_0),.clk(gclk));
	jdff dff_B_3sapSiPS0_0(.din(w_dff_B_4bl9Za4H4_0),.dout(w_dff_B_3sapSiPS0_0),.clk(gclk));
	jdff dff_B_KhuvoFix5_0(.din(w_dff_B_3sapSiPS0_0),.dout(w_dff_B_KhuvoFix5_0),.clk(gclk));
	jdff dff_B_lMUXr4I70_0(.din(w_dff_B_KhuvoFix5_0),.dout(w_dff_B_lMUXr4I70_0),.clk(gclk));
	jdff dff_B_f6r8Q5kc6_0(.din(w_dff_B_lMUXr4I70_0),.dout(w_dff_B_f6r8Q5kc6_0),.clk(gclk));
	jdff dff_B_oLrwJps75_0(.din(w_dff_B_f6r8Q5kc6_0),.dout(w_dff_B_oLrwJps75_0),.clk(gclk));
	jdff dff_B_t9Iu0MLT7_0(.din(w_dff_B_oLrwJps75_0),.dout(w_dff_B_t9Iu0MLT7_0),.clk(gclk));
	jdff dff_B_sez2YKZZ9_0(.din(w_dff_B_t9Iu0MLT7_0),.dout(w_dff_B_sez2YKZZ9_0),.clk(gclk));
	jdff dff_B_NamGkoJa6_0(.din(w_dff_B_sez2YKZZ9_0),.dout(w_dff_B_NamGkoJa6_0),.clk(gclk));
	jdff dff_B_xBEy1UkH8_0(.din(w_dff_B_NamGkoJa6_0),.dout(w_dff_B_xBEy1UkH8_0),.clk(gclk));
	jdff dff_B_FkU27wbF6_0(.din(w_dff_B_xBEy1UkH8_0),.dout(w_dff_B_FkU27wbF6_0),.clk(gclk));
	jdff dff_B_pBSIRIN01_0(.din(w_dff_B_FkU27wbF6_0),.dout(w_dff_B_pBSIRIN01_0),.clk(gclk));
	jdff dff_B_9nAlsUlr3_0(.din(w_dff_B_pBSIRIN01_0),.dout(w_dff_B_9nAlsUlr3_0),.clk(gclk));
	jdff dff_B_u4rYNDtK3_0(.din(w_dff_B_9nAlsUlr3_0),.dout(w_dff_B_u4rYNDtK3_0),.clk(gclk));
	jdff dff_B_PSnlgtFe9_0(.din(w_dff_B_u4rYNDtK3_0),.dout(w_dff_B_PSnlgtFe9_0),.clk(gclk));
	jdff dff_B_kkT2CKVd4_0(.din(w_dff_B_PSnlgtFe9_0),.dout(w_dff_B_kkT2CKVd4_0),.clk(gclk));
	jdff dff_B_GPuOuC477_0(.din(w_dff_B_kkT2CKVd4_0),.dout(w_dff_B_GPuOuC477_0),.clk(gclk));
	jdff dff_B_QVnjppW31_0(.din(w_dff_B_GPuOuC477_0),.dout(w_dff_B_QVnjppW31_0),.clk(gclk));
	jdff dff_B_KVxzluwI4_0(.din(w_dff_B_QVnjppW31_0),.dout(w_dff_B_KVxzluwI4_0),.clk(gclk));
	jdff dff_B_4luu63Vb9_0(.din(w_dff_B_KVxzluwI4_0),.dout(w_dff_B_4luu63Vb9_0),.clk(gclk));
	jdff dff_B_TiySji0B7_0(.din(w_dff_B_4luu63Vb9_0),.dout(w_dff_B_TiySji0B7_0),.clk(gclk));
	jdff dff_B_Px9S1YhM1_0(.din(w_dff_B_TiySji0B7_0),.dout(w_dff_B_Px9S1YhM1_0),.clk(gclk));
	jdff dff_B_rAMLmSKL9_0(.din(w_dff_B_Px9S1YhM1_0),.dout(w_dff_B_rAMLmSKL9_0),.clk(gclk));
	jdff dff_B_tY4ONek58_0(.din(w_dff_B_rAMLmSKL9_0),.dout(w_dff_B_tY4ONek58_0),.clk(gclk));
	jdff dff_B_8PiApWfS9_0(.din(w_dff_B_tY4ONek58_0),.dout(w_dff_B_8PiApWfS9_0),.clk(gclk));
	jdff dff_B_N3vIpLre2_0(.din(w_dff_B_8PiApWfS9_0),.dout(w_dff_B_N3vIpLre2_0),.clk(gclk));
	jdff dff_B_Cr822LdL2_0(.din(w_dff_B_N3vIpLre2_0),.dout(w_dff_B_Cr822LdL2_0),.clk(gclk));
	jdff dff_B_6oH8S5ZE0_0(.din(w_dff_B_Cr822LdL2_0),.dout(w_dff_B_6oH8S5ZE0_0),.clk(gclk));
	jdff dff_B_f1r3VukZ1_0(.din(w_dff_B_6oH8S5ZE0_0),.dout(w_dff_B_f1r3VukZ1_0),.clk(gclk));
	jdff dff_B_10cwXiW89_0(.din(w_dff_B_f1r3VukZ1_0),.dout(w_dff_B_10cwXiW89_0),.clk(gclk));
	jdff dff_B_5xQYjxiu8_0(.din(w_dff_B_10cwXiW89_0),.dout(w_dff_B_5xQYjxiu8_0),.clk(gclk));
	jdff dff_B_QUlRPTPT1_0(.din(w_dff_B_5xQYjxiu8_0),.dout(w_dff_B_QUlRPTPT1_0),.clk(gclk));
	jdff dff_B_umu8oH3l7_0(.din(w_dff_B_QUlRPTPT1_0),.dout(w_dff_B_umu8oH3l7_0),.clk(gclk));
	jdff dff_B_xDl0uCko9_0(.din(w_dff_B_umu8oH3l7_0),.dout(w_dff_B_xDl0uCko9_0),.clk(gclk));
	jdff dff_B_wldbdp9X1_0(.din(w_dff_B_xDl0uCko9_0),.dout(w_dff_B_wldbdp9X1_0),.clk(gclk));
	jdff dff_B_DEzZXAY44_0(.din(w_dff_B_wldbdp9X1_0),.dout(w_dff_B_DEzZXAY44_0),.clk(gclk));
	jdff dff_B_fgFgXz0K2_0(.din(w_dff_B_DEzZXAY44_0),.dout(w_dff_B_fgFgXz0K2_0),.clk(gclk));
	jdff dff_B_TJfmdXyR9_0(.din(w_dff_B_fgFgXz0K2_0),.dout(w_dff_B_TJfmdXyR9_0),.clk(gclk));
	jdff dff_B_jITTrzJr3_0(.din(w_dff_B_TJfmdXyR9_0),.dout(w_dff_B_jITTrzJr3_0),.clk(gclk));
	jdff dff_B_dfkGlCKW3_0(.din(w_dff_B_jITTrzJr3_0),.dout(w_dff_B_dfkGlCKW3_0),.clk(gclk));
	jdff dff_B_2HsMWCV05_0(.din(w_dff_B_dfkGlCKW3_0),.dout(w_dff_B_2HsMWCV05_0),.clk(gclk));
	jdff dff_B_IGnLiNoR8_0(.din(w_dff_B_2HsMWCV05_0),.dout(w_dff_B_IGnLiNoR8_0),.clk(gclk));
	jdff dff_B_Ee0N77Yf4_0(.din(w_dff_B_IGnLiNoR8_0),.dout(w_dff_B_Ee0N77Yf4_0),.clk(gclk));
	jdff dff_B_2yz6TJGX7_0(.din(w_dff_B_Ee0N77Yf4_0),.dout(w_dff_B_2yz6TJGX7_0),.clk(gclk));
	jdff dff_B_B35LWGEU2_0(.din(w_dff_B_2yz6TJGX7_0),.dout(w_dff_B_B35LWGEU2_0),.clk(gclk));
	jdff dff_B_CQUcic3R1_0(.din(w_dff_B_B35LWGEU2_0),.dout(w_dff_B_CQUcic3R1_0),.clk(gclk));
	jdff dff_B_T7Gd17DH7_0(.din(w_dff_B_CQUcic3R1_0),.dout(w_dff_B_T7Gd17DH7_0),.clk(gclk));
	jdff dff_B_ujDnUcL90_0(.din(w_dff_B_T7Gd17DH7_0),.dout(w_dff_B_ujDnUcL90_0),.clk(gclk));
	jdff dff_B_MNUzXlcS1_0(.din(w_dff_B_ujDnUcL90_0),.dout(w_dff_B_MNUzXlcS1_0),.clk(gclk));
	jdff dff_B_niRhq5lk6_0(.din(w_dff_B_MNUzXlcS1_0),.dout(w_dff_B_niRhq5lk6_0),.clk(gclk));
	jdff dff_B_ImrDGPBo9_0(.din(w_dff_B_niRhq5lk6_0),.dout(w_dff_B_ImrDGPBo9_0),.clk(gclk));
	jdff dff_B_3YQA7GhO9_1(.din(n1062),.dout(w_dff_B_3YQA7GhO9_1),.clk(gclk));
	jdff dff_B_7EGcvmRq3_1(.din(w_dff_B_3YQA7GhO9_1),.dout(w_dff_B_7EGcvmRq3_1),.clk(gclk));
	jdff dff_B_pUnIl0Xh3_1(.din(w_dff_B_7EGcvmRq3_1),.dout(w_dff_B_pUnIl0Xh3_1),.clk(gclk));
	jdff dff_B_5gwzeTxg7_1(.din(w_dff_B_pUnIl0Xh3_1),.dout(w_dff_B_5gwzeTxg7_1),.clk(gclk));
	jdff dff_B_6jaL3z8x1_1(.din(w_dff_B_5gwzeTxg7_1),.dout(w_dff_B_6jaL3z8x1_1),.clk(gclk));
	jdff dff_B_NvKWCXoq0_1(.din(w_dff_B_6jaL3z8x1_1),.dout(w_dff_B_NvKWCXoq0_1),.clk(gclk));
	jdff dff_B_znCzwP0g0_1(.din(w_dff_B_NvKWCXoq0_1),.dout(w_dff_B_znCzwP0g0_1),.clk(gclk));
	jdff dff_B_cbogA8Uf5_1(.din(w_dff_B_znCzwP0g0_1),.dout(w_dff_B_cbogA8Uf5_1),.clk(gclk));
	jdff dff_B_s9dFUFog4_1(.din(w_dff_B_cbogA8Uf5_1),.dout(w_dff_B_s9dFUFog4_1),.clk(gclk));
	jdff dff_B_B9SRpaRN6_1(.din(w_dff_B_s9dFUFog4_1),.dout(w_dff_B_B9SRpaRN6_1),.clk(gclk));
	jdff dff_B_nCnhwQNR3_1(.din(w_dff_B_B9SRpaRN6_1),.dout(w_dff_B_nCnhwQNR3_1),.clk(gclk));
	jdff dff_B_FOYIMpm94_1(.din(w_dff_B_nCnhwQNR3_1),.dout(w_dff_B_FOYIMpm94_1),.clk(gclk));
	jdff dff_B_M6mVhZ1P9_1(.din(w_dff_B_FOYIMpm94_1),.dout(w_dff_B_M6mVhZ1P9_1),.clk(gclk));
	jdff dff_B_KdElwcez9_1(.din(w_dff_B_M6mVhZ1P9_1),.dout(w_dff_B_KdElwcez9_1),.clk(gclk));
	jdff dff_B_yQ7FiiUG3_1(.din(w_dff_B_KdElwcez9_1),.dout(w_dff_B_yQ7FiiUG3_1),.clk(gclk));
	jdff dff_B_vq1MESMN7_1(.din(w_dff_B_yQ7FiiUG3_1),.dout(w_dff_B_vq1MESMN7_1),.clk(gclk));
	jdff dff_B_uRYvc69a5_1(.din(w_dff_B_vq1MESMN7_1),.dout(w_dff_B_uRYvc69a5_1),.clk(gclk));
	jdff dff_B_FurXDm5T5_1(.din(w_dff_B_uRYvc69a5_1),.dout(w_dff_B_FurXDm5T5_1),.clk(gclk));
	jdff dff_B_YZp21Yuy0_1(.din(w_dff_B_FurXDm5T5_1),.dout(w_dff_B_YZp21Yuy0_1),.clk(gclk));
	jdff dff_B_d6l3VUG36_1(.din(w_dff_B_YZp21Yuy0_1),.dout(w_dff_B_d6l3VUG36_1),.clk(gclk));
	jdff dff_B_fcZjSejq7_1(.din(w_dff_B_d6l3VUG36_1),.dout(w_dff_B_fcZjSejq7_1),.clk(gclk));
	jdff dff_B_NNZYOxKS1_1(.din(w_dff_B_fcZjSejq7_1),.dout(w_dff_B_NNZYOxKS1_1),.clk(gclk));
	jdff dff_B_spvH7CPH3_1(.din(w_dff_B_NNZYOxKS1_1),.dout(w_dff_B_spvH7CPH3_1),.clk(gclk));
	jdff dff_B_I2keuj8g4_1(.din(w_dff_B_spvH7CPH3_1),.dout(w_dff_B_I2keuj8g4_1),.clk(gclk));
	jdff dff_B_hdTPNeFH5_1(.din(w_dff_B_I2keuj8g4_1),.dout(w_dff_B_hdTPNeFH5_1),.clk(gclk));
	jdff dff_B_3uxEPy1t5_1(.din(w_dff_B_hdTPNeFH5_1),.dout(w_dff_B_3uxEPy1t5_1),.clk(gclk));
	jdff dff_B_hdaFrKyw2_1(.din(w_dff_B_3uxEPy1t5_1),.dout(w_dff_B_hdaFrKyw2_1),.clk(gclk));
	jdff dff_B_7CmvGMNf7_1(.din(w_dff_B_hdaFrKyw2_1),.dout(w_dff_B_7CmvGMNf7_1),.clk(gclk));
	jdff dff_B_IQOONsFh7_1(.din(w_dff_B_7CmvGMNf7_1),.dout(w_dff_B_IQOONsFh7_1),.clk(gclk));
	jdff dff_B_VtDU580u3_1(.din(w_dff_B_IQOONsFh7_1),.dout(w_dff_B_VtDU580u3_1),.clk(gclk));
	jdff dff_B_FSdbyO547_1(.din(w_dff_B_VtDU580u3_1),.dout(w_dff_B_FSdbyO547_1),.clk(gclk));
	jdff dff_B_AVrF9Nqd9_1(.din(w_dff_B_FSdbyO547_1),.dout(w_dff_B_AVrF9Nqd9_1),.clk(gclk));
	jdff dff_B_ETEiR65W2_1(.din(w_dff_B_AVrF9Nqd9_1),.dout(w_dff_B_ETEiR65W2_1),.clk(gclk));
	jdff dff_B_j3AUtkRy7_1(.din(w_dff_B_ETEiR65W2_1),.dout(w_dff_B_j3AUtkRy7_1),.clk(gclk));
	jdff dff_B_aOgU4ELB6_1(.din(w_dff_B_j3AUtkRy7_1),.dout(w_dff_B_aOgU4ELB6_1),.clk(gclk));
	jdff dff_B_jBp8iQ3Q9_1(.din(w_dff_B_aOgU4ELB6_1),.dout(w_dff_B_jBp8iQ3Q9_1),.clk(gclk));
	jdff dff_B_g0i2eiEM2_1(.din(w_dff_B_jBp8iQ3Q9_1),.dout(w_dff_B_g0i2eiEM2_1),.clk(gclk));
	jdff dff_B_naq7KaiY9_1(.din(w_dff_B_g0i2eiEM2_1),.dout(w_dff_B_naq7KaiY9_1),.clk(gclk));
	jdff dff_B_m4BD1M7t1_1(.din(w_dff_B_naq7KaiY9_1),.dout(w_dff_B_m4BD1M7t1_1),.clk(gclk));
	jdff dff_B_qFC3XSkr0_1(.din(w_dff_B_m4BD1M7t1_1),.dout(w_dff_B_qFC3XSkr0_1),.clk(gclk));
	jdff dff_B_2H7MoZBm6_1(.din(w_dff_B_qFC3XSkr0_1),.dout(w_dff_B_2H7MoZBm6_1),.clk(gclk));
	jdff dff_B_4ffmlxfy8_1(.din(w_dff_B_2H7MoZBm6_1),.dout(w_dff_B_4ffmlxfy8_1),.clk(gclk));
	jdff dff_B_qkn14MKe0_1(.din(w_dff_B_4ffmlxfy8_1),.dout(w_dff_B_qkn14MKe0_1),.clk(gclk));
	jdff dff_B_GV0mab0N4_1(.din(w_dff_B_qkn14MKe0_1),.dout(w_dff_B_GV0mab0N4_1),.clk(gclk));
	jdff dff_B_fzBtasrw2_1(.din(w_dff_B_GV0mab0N4_1),.dout(w_dff_B_fzBtasrw2_1),.clk(gclk));
	jdff dff_B_5dTKk3Gk5_1(.din(w_dff_B_fzBtasrw2_1),.dout(w_dff_B_5dTKk3Gk5_1),.clk(gclk));
	jdff dff_B_5rHczfM12_1(.din(w_dff_B_5dTKk3Gk5_1),.dout(w_dff_B_5rHczfM12_1),.clk(gclk));
	jdff dff_B_BARQITdw4_1(.din(w_dff_B_5rHczfM12_1),.dout(w_dff_B_BARQITdw4_1),.clk(gclk));
	jdff dff_B_S6Xp7R9T7_1(.din(w_dff_B_BARQITdw4_1),.dout(w_dff_B_S6Xp7R9T7_1),.clk(gclk));
	jdff dff_B_CJy5Xudd4_1(.din(w_dff_B_S6Xp7R9T7_1),.dout(w_dff_B_CJy5Xudd4_1),.clk(gclk));
	jdff dff_B_UYfj7fOI1_1(.din(w_dff_B_CJy5Xudd4_1),.dout(w_dff_B_UYfj7fOI1_1),.clk(gclk));
	jdff dff_B_yS4atw2d4_1(.din(w_dff_B_UYfj7fOI1_1),.dout(w_dff_B_yS4atw2d4_1),.clk(gclk));
	jdff dff_B_NswG0Ans4_1(.din(w_dff_B_yS4atw2d4_1),.dout(w_dff_B_NswG0Ans4_1),.clk(gclk));
	jdff dff_B_un6YYT3w5_1(.din(w_dff_B_NswG0Ans4_1),.dout(w_dff_B_un6YYT3w5_1),.clk(gclk));
	jdff dff_B_cd3W0sKe7_1(.din(w_dff_B_un6YYT3w5_1),.dout(w_dff_B_cd3W0sKe7_1),.clk(gclk));
	jdff dff_B_PxnsfXQZ8_1(.din(w_dff_B_cd3W0sKe7_1),.dout(w_dff_B_PxnsfXQZ8_1),.clk(gclk));
	jdff dff_B_s8ZLoxsW1_1(.din(w_dff_B_PxnsfXQZ8_1),.dout(w_dff_B_s8ZLoxsW1_1),.clk(gclk));
	jdff dff_B_68u018ga6_1(.din(w_dff_B_s8ZLoxsW1_1),.dout(w_dff_B_68u018ga6_1),.clk(gclk));
	jdff dff_B_FqSwABMJ7_1(.din(w_dff_B_68u018ga6_1),.dout(w_dff_B_FqSwABMJ7_1),.clk(gclk));
	jdff dff_B_DQBQpGpU6_1(.din(w_dff_B_FqSwABMJ7_1),.dout(w_dff_B_DQBQpGpU6_1),.clk(gclk));
	jdff dff_B_c6elk3rw8_1(.din(w_dff_B_DQBQpGpU6_1),.dout(w_dff_B_c6elk3rw8_1),.clk(gclk));
	jdff dff_B_2LS1FMrT4_1(.din(w_dff_B_c6elk3rw8_1),.dout(w_dff_B_2LS1FMrT4_1),.clk(gclk));
	jdff dff_B_J0Fw0MuX7_1(.din(w_dff_B_2LS1FMrT4_1),.dout(w_dff_B_J0Fw0MuX7_1),.clk(gclk));
	jdff dff_B_TjlvXwnq4_1(.din(w_dff_B_J0Fw0MuX7_1),.dout(w_dff_B_TjlvXwnq4_1),.clk(gclk));
	jdff dff_B_svhjiGLW0_1(.din(w_dff_B_TjlvXwnq4_1),.dout(w_dff_B_svhjiGLW0_1),.clk(gclk));
	jdff dff_B_y1tLFf3b4_1(.din(w_dff_B_svhjiGLW0_1),.dout(w_dff_B_y1tLFf3b4_1),.clk(gclk));
	jdff dff_B_dXwZTh0u6_1(.din(w_dff_B_y1tLFf3b4_1),.dout(w_dff_B_dXwZTh0u6_1),.clk(gclk));
	jdff dff_B_2MiLxxwT9_1(.din(w_dff_B_dXwZTh0u6_1),.dout(w_dff_B_2MiLxxwT9_1),.clk(gclk));
	jdff dff_B_5h9EYBja3_1(.din(w_dff_B_2MiLxxwT9_1),.dout(w_dff_B_5h9EYBja3_1),.clk(gclk));
	jdff dff_B_uuDfBczC4_1(.din(w_dff_B_5h9EYBja3_1),.dout(w_dff_B_uuDfBczC4_1),.clk(gclk));
	jdff dff_B_bodVyx9Q6_1(.din(w_dff_B_uuDfBczC4_1),.dout(w_dff_B_bodVyx9Q6_1),.clk(gclk));
	jdff dff_B_0YEbGJsP3_1(.din(w_dff_B_bodVyx9Q6_1),.dout(w_dff_B_0YEbGJsP3_1),.clk(gclk));
	jdff dff_B_mKcGy4RO9_1(.din(w_dff_B_0YEbGJsP3_1),.dout(w_dff_B_mKcGy4RO9_1),.clk(gclk));
	jdff dff_B_Zofr1Qmk2_1(.din(w_dff_B_mKcGy4RO9_1),.dout(w_dff_B_Zofr1Qmk2_1),.clk(gclk));
	jdff dff_B_UCeFjkBI3_1(.din(w_dff_B_Zofr1Qmk2_1),.dout(w_dff_B_UCeFjkBI3_1),.clk(gclk));
	jdff dff_B_Bi5E5g4R2_1(.din(w_dff_B_UCeFjkBI3_1),.dout(w_dff_B_Bi5E5g4R2_1),.clk(gclk));
	jdff dff_B_HWGdJFXr9_1(.din(w_dff_B_Bi5E5g4R2_1),.dout(w_dff_B_HWGdJFXr9_1),.clk(gclk));
	jdff dff_B_Y3aalqrp4_1(.din(w_dff_B_HWGdJFXr9_1),.dout(w_dff_B_Y3aalqrp4_1),.clk(gclk));
	jdff dff_B_694Nfgxd3_1(.din(w_dff_B_Y3aalqrp4_1),.dout(w_dff_B_694Nfgxd3_1),.clk(gclk));
	jdff dff_B_5nkSaVSg7_1(.din(w_dff_B_694Nfgxd3_1),.dout(w_dff_B_5nkSaVSg7_1),.clk(gclk));
	jdff dff_B_3ae3CVYA4_1(.din(w_dff_B_5nkSaVSg7_1),.dout(w_dff_B_3ae3CVYA4_1),.clk(gclk));
	jdff dff_B_qwKXXEMs6_1(.din(w_dff_B_3ae3CVYA4_1),.dout(w_dff_B_qwKXXEMs6_1),.clk(gclk));
	jdff dff_B_vwIKYOXo0_1(.din(w_dff_B_qwKXXEMs6_1),.dout(w_dff_B_vwIKYOXo0_1),.clk(gclk));
	jdff dff_B_EkvemZGx2_1(.din(w_dff_B_vwIKYOXo0_1),.dout(w_dff_B_EkvemZGx2_1),.clk(gclk));
	jdff dff_B_GWiituuR1_1(.din(w_dff_B_EkvemZGx2_1),.dout(w_dff_B_GWiituuR1_1),.clk(gclk));
	jdff dff_B_cAicZc2D5_1(.din(w_dff_B_GWiituuR1_1),.dout(w_dff_B_cAicZc2D5_1),.clk(gclk));
	jdff dff_B_EJZE4J9r1_1(.din(w_dff_B_cAicZc2D5_1),.dout(w_dff_B_EJZE4J9r1_1),.clk(gclk));
	jdff dff_B_h1oZradx8_1(.din(w_dff_B_EJZE4J9r1_1),.dout(w_dff_B_h1oZradx8_1),.clk(gclk));
	jdff dff_B_1yxZmgRd1_1(.din(w_dff_B_h1oZradx8_1),.dout(w_dff_B_1yxZmgRd1_1),.clk(gclk));
	jdff dff_B_uDLlYtDu1_1(.din(w_dff_B_1yxZmgRd1_1),.dout(w_dff_B_uDLlYtDu1_1),.clk(gclk));
	jdff dff_B_leKrtHrF3_1(.din(w_dff_B_uDLlYtDu1_1),.dout(w_dff_B_leKrtHrF3_1),.clk(gclk));
	jdff dff_B_oAT0uDd04_1(.din(w_dff_B_leKrtHrF3_1),.dout(w_dff_B_oAT0uDd04_1),.clk(gclk));
	jdff dff_B_LBcou8w18_1(.din(w_dff_B_oAT0uDd04_1),.dout(w_dff_B_LBcou8w18_1),.clk(gclk));
	jdff dff_B_edF1hDSZ5_1(.din(w_dff_B_LBcou8w18_1),.dout(w_dff_B_edF1hDSZ5_1),.clk(gclk));
	jdff dff_B_trYikcLE6_1(.din(w_dff_B_edF1hDSZ5_1),.dout(w_dff_B_trYikcLE6_1),.clk(gclk));
	jdff dff_B_2ijSUluq4_1(.din(w_dff_B_trYikcLE6_1),.dout(w_dff_B_2ijSUluq4_1),.clk(gclk));
	jdff dff_B_cK3bqB2z0_1(.din(w_dff_B_2ijSUluq4_1),.dout(w_dff_B_cK3bqB2z0_1),.clk(gclk));
	jdff dff_B_X3eQIbMu3_1(.din(w_dff_B_cK3bqB2z0_1),.dout(w_dff_B_X3eQIbMu3_1),.clk(gclk));
	jdff dff_B_1wTGGqE21_1(.din(w_dff_B_X3eQIbMu3_1),.dout(w_dff_B_1wTGGqE21_1),.clk(gclk));
	jdff dff_B_RChdCOTh8_1(.din(w_dff_B_1wTGGqE21_1),.dout(w_dff_B_RChdCOTh8_1),.clk(gclk));
	jdff dff_B_wh6kJdJV9_1(.din(w_dff_B_RChdCOTh8_1),.dout(w_dff_B_wh6kJdJV9_1),.clk(gclk));
	jdff dff_B_YNnywHuL3_1(.din(w_dff_B_wh6kJdJV9_1),.dout(w_dff_B_YNnywHuL3_1),.clk(gclk));
	jdff dff_B_V2jjIySG7_1(.din(w_dff_B_YNnywHuL3_1),.dout(w_dff_B_V2jjIySG7_1),.clk(gclk));
	jdff dff_B_JXQfFvYb1_1(.din(w_dff_B_V2jjIySG7_1),.dout(w_dff_B_JXQfFvYb1_1),.clk(gclk));
	jdff dff_B_ktrX3pFw7_1(.din(w_dff_B_JXQfFvYb1_1),.dout(w_dff_B_ktrX3pFw7_1),.clk(gclk));
	jdff dff_B_g5pGDcfh4_1(.din(w_dff_B_ktrX3pFw7_1),.dout(w_dff_B_g5pGDcfh4_1),.clk(gclk));
	jdff dff_B_ls9plk3d3_1(.din(w_dff_B_g5pGDcfh4_1),.dout(w_dff_B_ls9plk3d3_1),.clk(gclk));
	jdff dff_B_Wtb0mdY08_1(.din(w_dff_B_ls9plk3d3_1),.dout(w_dff_B_Wtb0mdY08_1),.clk(gclk));
	jdff dff_B_TtFRaT1f7_1(.din(w_dff_B_Wtb0mdY08_1),.dout(w_dff_B_TtFRaT1f7_1),.clk(gclk));
	jdff dff_B_bcnFMOvs1_1(.din(w_dff_B_TtFRaT1f7_1),.dout(w_dff_B_bcnFMOvs1_1),.clk(gclk));
	jdff dff_B_kx5kWE2b9_1(.din(w_dff_B_bcnFMOvs1_1),.dout(w_dff_B_kx5kWE2b9_1),.clk(gclk));
	jdff dff_B_VQf37a1h2_1(.din(w_dff_B_kx5kWE2b9_1),.dout(w_dff_B_VQf37a1h2_1),.clk(gclk));
	jdff dff_B_XYc0K6132_1(.din(w_dff_B_VQf37a1h2_1),.dout(w_dff_B_XYc0K6132_1),.clk(gclk));
	jdff dff_B_EzaJodqS8_0(.din(n1063),.dout(w_dff_B_EzaJodqS8_0),.clk(gclk));
	jdff dff_B_zP9IFLva5_0(.din(w_dff_B_EzaJodqS8_0),.dout(w_dff_B_zP9IFLva5_0),.clk(gclk));
	jdff dff_B_Tbfqh9zA3_0(.din(w_dff_B_zP9IFLva5_0),.dout(w_dff_B_Tbfqh9zA3_0),.clk(gclk));
	jdff dff_B_Cwt730ap3_0(.din(w_dff_B_Tbfqh9zA3_0),.dout(w_dff_B_Cwt730ap3_0),.clk(gclk));
	jdff dff_B_cy1KuHkc1_0(.din(w_dff_B_Cwt730ap3_0),.dout(w_dff_B_cy1KuHkc1_0),.clk(gclk));
	jdff dff_B_CSikebnx7_0(.din(w_dff_B_cy1KuHkc1_0),.dout(w_dff_B_CSikebnx7_0),.clk(gclk));
	jdff dff_B_t9C8YF5G1_0(.din(w_dff_B_CSikebnx7_0),.dout(w_dff_B_t9C8YF5G1_0),.clk(gclk));
	jdff dff_B_s8yVXaTS5_0(.din(w_dff_B_t9C8YF5G1_0),.dout(w_dff_B_s8yVXaTS5_0),.clk(gclk));
	jdff dff_B_aJeEXzM93_0(.din(w_dff_B_s8yVXaTS5_0),.dout(w_dff_B_aJeEXzM93_0),.clk(gclk));
	jdff dff_B_QdFdyFSq2_0(.din(w_dff_B_aJeEXzM93_0),.dout(w_dff_B_QdFdyFSq2_0),.clk(gclk));
	jdff dff_B_jdvTHacl8_0(.din(w_dff_B_QdFdyFSq2_0),.dout(w_dff_B_jdvTHacl8_0),.clk(gclk));
	jdff dff_B_wDvCAyRX8_0(.din(w_dff_B_jdvTHacl8_0),.dout(w_dff_B_wDvCAyRX8_0),.clk(gclk));
	jdff dff_B_RMSbwqqE2_0(.din(w_dff_B_wDvCAyRX8_0),.dout(w_dff_B_RMSbwqqE2_0),.clk(gclk));
	jdff dff_B_xDL61mur8_0(.din(w_dff_B_RMSbwqqE2_0),.dout(w_dff_B_xDL61mur8_0),.clk(gclk));
	jdff dff_B_ZO8MFldP8_0(.din(w_dff_B_xDL61mur8_0),.dout(w_dff_B_ZO8MFldP8_0),.clk(gclk));
	jdff dff_B_X0KhYbQ66_0(.din(w_dff_B_ZO8MFldP8_0),.dout(w_dff_B_X0KhYbQ66_0),.clk(gclk));
	jdff dff_B_dVn7ltZl7_0(.din(w_dff_B_X0KhYbQ66_0),.dout(w_dff_B_dVn7ltZl7_0),.clk(gclk));
	jdff dff_B_vxWHWu4e2_0(.din(w_dff_B_dVn7ltZl7_0),.dout(w_dff_B_vxWHWu4e2_0),.clk(gclk));
	jdff dff_B_W9yqDw8o0_0(.din(w_dff_B_vxWHWu4e2_0),.dout(w_dff_B_W9yqDw8o0_0),.clk(gclk));
	jdff dff_B_CjTMqDBl6_0(.din(w_dff_B_W9yqDw8o0_0),.dout(w_dff_B_CjTMqDBl6_0),.clk(gclk));
	jdff dff_B_hInJTAAg2_0(.din(w_dff_B_CjTMqDBl6_0),.dout(w_dff_B_hInJTAAg2_0),.clk(gclk));
	jdff dff_B_HXswUPXO0_0(.din(w_dff_B_hInJTAAg2_0),.dout(w_dff_B_HXswUPXO0_0),.clk(gclk));
	jdff dff_B_1Rl8B2Dz8_0(.din(w_dff_B_HXswUPXO0_0),.dout(w_dff_B_1Rl8B2Dz8_0),.clk(gclk));
	jdff dff_B_v0oqxoB94_0(.din(w_dff_B_1Rl8B2Dz8_0),.dout(w_dff_B_v0oqxoB94_0),.clk(gclk));
	jdff dff_B_MIFTPmTL7_0(.din(w_dff_B_v0oqxoB94_0),.dout(w_dff_B_MIFTPmTL7_0),.clk(gclk));
	jdff dff_B_bBDwxaEU5_0(.din(w_dff_B_MIFTPmTL7_0),.dout(w_dff_B_bBDwxaEU5_0),.clk(gclk));
	jdff dff_B_WXLUjImo9_0(.din(w_dff_B_bBDwxaEU5_0),.dout(w_dff_B_WXLUjImo9_0),.clk(gclk));
	jdff dff_B_NK50IKiS3_0(.din(w_dff_B_WXLUjImo9_0),.dout(w_dff_B_NK50IKiS3_0),.clk(gclk));
	jdff dff_B_2YiMrnQS0_0(.din(w_dff_B_NK50IKiS3_0),.dout(w_dff_B_2YiMrnQS0_0),.clk(gclk));
	jdff dff_B_tVBaLwx42_0(.din(w_dff_B_2YiMrnQS0_0),.dout(w_dff_B_tVBaLwx42_0),.clk(gclk));
	jdff dff_B_fLtHDs0x3_0(.din(w_dff_B_tVBaLwx42_0),.dout(w_dff_B_fLtHDs0x3_0),.clk(gclk));
	jdff dff_B_Xjiu6Mnu7_0(.din(w_dff_B_fLtHDs0x3_0),.dout(w_dff_B_Xjiu6Mnu7_0),.clk(gclk));
	jdff dff_B_XFhThrOF0_0(.din(w_dff_B_Xjiu6Mnu7_0),.dout(w_dff_B_XFhThrOF0_0),.clk(gclk));
	jdff dff_B_FA6HpplW5_0(.din(w_dff_B_XFhThrOF0_0),.dout(w_dff_B_FA6HpplW5_0),.clk(gclk));
	jdff dff_B_ojhXwi681_0(.din(w_dff_B_FA6HpplW5_0),.dout(w_dff_B_ojhXwi681_0),.clk(gclk));
	jdff dff_B_9NYK3v9Z0_0(.din(w_dff_B_ojhXwi681_0),.dout(w_dff_B_9NYK3v9Z0_0),.clk(gclk));
	jdff dff_B_MCt5C8fh3_0(.din(w_dff_B_9NYK3v9Z0_0),.dout(w_dff_B_MCt5C8fh3_0),.clk(gclk));
	jdff dff_B_bCCKn63x3_0(.din(w_dff_B_MCt5C8fh3_0),.dout(w_dff_B_bCCKn63x3_0),.clk(gclk));
	jdff dff_B_q0ybYMd12_0(.din(w_dff_B_bCCKn63x3_0),.dout(w_dff_B_q0ybYMd12_0),.clk(gclk));
	jdff dff_B_euud8xNN7_0(.din(w_dff_B_q0ybYMd12_0),.dout(w_dff_B_euud8xNN7_0),.clk(gclk));
	jdff dff_B_Y2Vo3erM5_0(.din(w_dff_B_euud8xNN7_0),.dout(w_dff_B_Y2Vo3erM5_0),.clk(gclk));
	jdff dff_B_qhJxRSJ44_0(.din(w_dff_B_Y2Vo3erM5_0),.dout(w_dff_B_qhJxRSJ44_0),.clk(gclk));
	jdff dff_B_EBNT5MeV9_0(.din(w_dff_B_qhJxRSJ44_0),.dout(w_dff_B_EBNT5MeV9_0),.clk(gclk));
	jdff dff_B_YnX8SGd08_0(.din(w_dff_B_EBNT5MeV9_0),.dout(w_dff_B_YnX8SGd08_0),.clk(gclk));
	jdff dff_B_2kQGa55j6_0(.din(w_dff_B_YnX8SGd08_0),.dout(w_dff_B_2kQGa55j6_0),.clk(gclk));
	jdff dff_B_obwXsIGL8_0(.din(w_dff_B_2kQGa55j6_0),.dout(w_dff_B_obwXsIGL8_0),.clk(gclk));
	jdff dff_B_gdTSAvy01_0(.din(w_dff_B_obwXsIGL8_0),.dout(w_dff_B_gdTSAvy01_0),.clk(gclk));
	jdff dff_B_mHLn9DCy3_0(.din(w_dff_B_gdTSAvy01_0),.dout(w_dff_B_mHLn9DCy3_0),.clk(gclk));
	jdff dff_B_A1Djr5mL5_0(.din(w_dff_B_mHLn9DCy3_0),.dout(w_dff_B_A1Djr5mL5_0),.clk(gclk));
	jdff dff_B_Vp1hRAYR3_0(.din(w_dff_B_A1Djr5mL5_0),.dout(w_dff_B_Vp1hRAYR3_0),.clk(gclk));
	jdff dff_B_YtUm7cWw3_0(.din(w_dff_B_Vp1hRAYR3_0),.dout(w_dff_B_YtUm7cWw3_0),.clk(gclk));
	jdff dff_B_snbSRhzY7_0(.din(w_dff_B_YtUm7cWw3_0),.dout(w_dff_B_snbSRhzY7_0),.clk(gclk));
	jdff dff_B_7mOYbSHb8_0(.din(w_dff_B_snbSRhzY7_0),.dout(w_dff_B_7mOYbSHb8_0),.clk(gclk));
	jdff dff_B_RxgRsp3S6_0(.din(w_dff_B_7mOYbSHb8_0),.dout(w_dff_B_RxgRsp3S6_0),.clk(gclk));
	jdff dff_B_TTEbFWa84_0(.din(w_dff_B_RxgRsp3S6_0),.dout(w_dff_B_TTEbFWa84_0),.clk(gclk));
	jdff dff_B_pJYDz0MA3_0(.din(w_dff_B_TTEbFWa84_0),.dout(w_dff_B_pJYDz0MA3_0),.clk(gclk));
	jdff dff_B_W5BfMJYa0_0(.din(w_dff_B_pJYDz0MA3_0),.dout(w_dff_B_W5BfMJYa0_0),.clk(gclk));
	jdff dff_B_Zd3kwPHU1_0(.din(w_dff_B_W5BfMJYa0_0),.dout(w_dff_B_Zd3kwPHU1_0),.clk(gclk));
	jdff dff_B_SFBUncDH0_0(.din(w_dff_B_Zd3kwPHU1_0),.dout(w_dff_B_SFBUncDH0_0),.clk(gclk));
	jdff dff_B_Dp1BL3Ip1_0(.din(w_dff_B_SFBUncDH0_0),.dout(w_dff_B_Dp1BL3Ip1_0),.clk(gclk));
	jdff dff_B_KlGlmZea4_0(.din(w_dff_B_Dp1BL3Ip1_0),.dout(w_dff_B_KlGlmZea4_0),.clk(gclk));
	jdff dff_B_8bIsnR6f2_0(.din(w_dff_B_KlGlmZea4_0),.dout(w_dff_B_8bIsnR6f2_0),.clk(gclk));
	jdff dff_B_VwcpeNwQ2_0(.din(w_dff_B_8bIsnR6f2_0),.dout(w_dff_B_VwcpeNwQ2_0),.clk(gclk));
	jdff dff_B_zjprAQc92_0(.din(w_dff_B_VwcpeNwQ2_0),.dout(w_dff_B_zjprAQc92_0),.clk(gclk));
	jdff dff_B_zlkwCEOt7_0(.din(w_dff_B_zjprAQc92_0),.dout(w_dff_B_zlkwCEOt7_0),.clk(gclk));
	jdff dff_B_jGVr0YIp3_0(.din(w_dff_B_zlkwCEOt7_0),.dout(w_dff_B_jGVr0YIp3_0),.clk(gclk));
	jdff dff_B_IlVMj93h0_0(.din(w_dff_B_jGVr0YIp3_0),.dout(w_dff_B_IlVMj93h0_0),.clk(gclk));
	jdff dff_B_rWdFK9hF0_0(.din(w_dff_B_IlVMj93h0_0),.dout(w_dff_B_rWdFK9hF0_0),.clk(gclk));
	jdff dff_B_ViOOoSv25_0(.din(w_dff_B_rWdFK9hF0_0),.dout(w_dff_B_ViOOoSv25_0),.clk(gclk));
	jdff dff_B_8nK4QXOd6_0(.din(w_dff_B_ViOOoSv25_0),.dout(w_dff_B_8nK4QXOd6_0),.clk(gclk));
	jdff dff_B_gxbzngQU7_0(.din(w_dff_B_8nK4QXOd6_0),.dout(w_dff_B_gxbzngQU7_0),.clk(gclk));
	jdff dff_B_NSLytmao5_0(.din(w_dff_B_gxbzngQU7_0),.dout(w_dff_B_NSLytmao5_0),.clk(gclk));
	jdff dff_B_7hn2KMY03_0(.din(w_dff_B_NSLytmao5_0),.dout(w_dff_B_7hn2KMY03_0),.clk(gclk));
	jdff dff_B_avi2Sthf6_0(.din(w_dff_B_7hn2KMY03_0),.dout(w_dff_B_avi2Sthf6_0),.clk(gclk));
	jdff dff_B_Z6X1g8iq5_0(.din(w_dff_B_avi2Sthf6_0),.dout(w_dff_B_Z6X1g8iq5_0),.clk(gclk));
	jdff dff_B_i4Og4My66_0(.din(w_dff_B_Z6X1g8iq5_0),.dout(w_dff_B_i4Og4My66_0),.clk(gclk));
	jdff dff_B_mdAtJWfp1_0(.din(w_dff_B_i4Og4My66_0),.dout(w_dff_B_mdAtJWfp1_0),.clk(gclk));
	jdff dff_B_v8vyGl5N8_0(.din(w_dff_B_mdAtJWfp1_0),.dout(w_dff_B_v8vyGl5N8_0),.clk(gclk));
	jdff dff_B_0QReq4ua6_0(.din(w_dff_B_v8vyGl5N8_0),.dout(w_dff_B_0QReq4ua6_0),.clk(gclk));
	jdff dff_B_W21oVGa69_0(.din(w_dff_B_0QReq4ua6_0),.dout(w_dff_B_W21oVGa69_0),.clk(gclk));
	jdff dff_B_AI11iYyS8_0(.din(w_dff_B_W21oVGa69_0),.dout(w_dff_B_AI11iYyS8_0),.clk(gclk));
	jdff dff_B_1cVDvt215_0(.din(w_dff_B_AI11iYyS8_0),.dout(w_dff_B_1cVDvt215_0),.clk(gclk));
	jdff dff_B_5L1xQX1p4_0(.din(w_dff_B_1cVDvt215_0),.dout(w_dff_B_5L1xQX1p4_0),.clk(gclk));
	jdff dff_B_TlSqn3Pj0_0(.din(w_dff_B_5L1xQX1p4_0),.dout(w_dff_B_TlSqn3Pj0_0),.clk(gclk));
	jdff dff_B_swBtowFI2_0(.din(w_dff_B_TlSqn3Pj0_0),.dout(w_dff_B_swBtowFI2_0),.clk(gclk));
	jdff dff_B_T8dJDN1p1_0(.din(w_dff_B_swBtowFI2_0),.dout(w_dff_B_T8dJDN1p1_0),.clk(gclk));
	jdff dff_B_8Z3eKigZ2_0(.din(w_dff_B_T8dJDN1p1_0),.dout(w_dff_B_8Z3eKigZ2_0),.clk(gclk));
	jdff dff_B_fihr9Zdv1_0(.din(w_dff_B_8Z3eKigZ2_0),.dout(w_dff_B_fihr9Zdv1_0),.clk(gclk));
	jdff dff_B_rSXCiBYb8_0(.din(w_dff_B_fihr9Zdv1_0),.dout(w_dff_B_rSXCiBYb8_0),.clk(gclk));
	jdff dff_B_Cb0KbrkC5_0(.din(w_dff_B_rSXCiBYb8_0),.dout(w_dff_B_Cb0KbrkC5_0),.clk(gclk));
	jdff dff_B_c9NF1VNd0_0(.din(w_dff_B_Cb0KbrkC5_0),.dout(w_dff_B_c9NF1VNd0_0),.clk(gclk));
	jdff dff_B_hg4UEku54_0(.din(w_dff_B_c9NF1VNd0_0),.dout(w_dff_B_hg4UEku54_0),.clk(gclk));
	jdff dff_B_ZAsXg52V5_0(.din(w_dff_B_hg4UEku54_0),.dout(w_dff_B_ZAsXg52V5_0),.clk(gclk));
	jdff dff_B_L3vW8Ise2_0(.din(w_dff_B_ZAsXg52V5_0),.dout(w_dff_B_L3vW8Ise2_0),.clk(gclk));
	jdff dff_B_ODlMj3Lr1_0(.din(w_dff_B_L3vW8Ise2_0),.dout(w_dff_B_ODlMj3Lr1_0),.clk(gclk));
	jdff dff_B_LYbrjwl59_0(.din(w_dff_B_ODlMj3Lr1_0),.dout(w_dff_B_LYbrjwl59_0),.clk(gclk));
	jdff dff_B_Eipc1ETl2_0(.din(w_dff_B_LYbrjwl59_0),.dout(w_dff_B_Eipc1ETl2_0),.clk(gclk));
	jdff dff_B_Xt1ZESqP2_0(.din(w_dff_B_Eipc1ETl2_0),.dout(w_dff_B_Xt1ZESqP2_0),.clk(gclk));
	jdff dff_B_NKXseSeN5_0(.din(w_dff_B_Xt1ZESqP2_0),.dout(w_dff_B_NKXseSeN5_0),.clk(gclk));
	jdff dff_B_05y7fX6B6_0(.din(w_dff_B_NKXseSeN5_0),.dout(w_dff_B_05y7fX6B6_0),.clk(gclk));
	jdff dff_B_aRt1Bn6g6_0(.din(w_dff_B_05y7fX6B6_0),.dout(w_dff_B_aRt1Bn6g6_0),.clk(gclk));
	jdff dff_B_opvjvs1u1_0(.din(w_dff_B_aRt1Bn6g6_0),.dout(w_dff_B_opvjvs1u1_0),.clk(gclk));
	jdff dff_B_kAHZOL9x7_0(.din(w_dff_B_opvjvs1u1_0),.dout(w_dff_B_kAHZOL9x7_0),.clk(gclk));
	jdff dff_B_sAfaT4qB9_0(.din(w_dff_B_kAHZOL9x7_0),.dout(w_dff_B_sAfaT4qB9_0),.clk(gclk));
	jdff dff_B_INXXsf2p8_0(.din(w_dff_B_sAfaT4qB9_0),.dout(w_dff_B_INXXsf2p8_0),.clk(gclk));
	jdff dff_B_mv8K2Y7q9_0(.din(w_dff_B_INXXsf2p8_0),.dout(w_dff_B_mv8K2Y7q9_0),.clk(gclk));
	jdff dff_B_F9qpmOda1_0(.din(w_dff_B_mv8K2Y7q9_0),.dout(w_dff_B_F9qpmOda1_0),.clk(gclk));
	jdff dff_B_yF8jyCHj7_0(.din(w_dff_B_F9qpmOda1_0),.dout(w_dff_B_yF8jyCHj7_0),.clk(gclk));
	jdff dff_B_cCpjDktR2_0(.din(w_dff_B_yF8jyCHj7_0),.dout(w_dff_B_cCpjDktR2_0),.clk(gclk));
	jdff dff_B_SjSOfdQk3_0(.din(w_dff_B_cCpjDktR2_0),.dout(w_dff_B_SjSOfdQk3_0),.clk(gclk));
	jdff dff_B_RljpaGqd9_0(.din(w_dff_B_SjSOfdQk3_0),.dout(w_dff_B_RljpaGqd9_0),.clk(gclk));
	jdff dff_B_9stgRsss9_0(.din(w_dff_B_RljpaGqd9_0),.dout(w_dff_B_9stgRsss9_0),.clk(gclk));
	jdff dff_B_mK9qdiWp4_0(.din(w_dff_B_9stgRsss9_0),.dout(w_dff_B_mK9qdiWp4_0),.clk(gclk));
	jdff dff_B_6gTBK1EM9_1(.din(n1056),.dout(w_dff_B_6gTBK1EM9_1),.clk(gclk));
	jdff dff_B_uO3UTTnK8_1(.din(w_dff_B_6gTBK1EM9_1),.dout(w_dff_B_uO3UTTnK8_1),.clk(gclk));
	jdff dff_B_5EwD6ijE8_1(.din(w_dff_B_uO3UTTnK8_1),.dout(w_dff_B_5EwD6ijE8_1),.clk(gclk));
	jdff dff_B_SS19RUqy0_1(.din(w_dff_B_5EwD6ijE8_1),.dout(w_dff_B_SS19RUqy0_1),.clk(gclk));
	jdff dff_B_3Auiu3ZY0_1(.din(w_dff_B_SS19RUqy0_1),.dout(w_dff_B_3Auiu3ZY0_1),.clk(gclk));
	jdff dff_B_PyWlXHIR0_1(.din(w_dff_B_3Auiu3ZY0_1),.dout(w_dff_B_PyWlXHIR0_1),.clk(gclk));
	jdff dff_B_8YIlveUk2_1(.din(w_dff_B_PyWlXHIR0_1),.dout(w_dff_B_8YIlveUk2_1),.clk(gclk));
	jdff dff_B_1irRMUgK8_1(.din(w_dff_B_8YIlveUk2_1),.dout(w_dff_B_1irRMUgK8_1),.clk(gclk));
	jdff dff_B_KABtyeGH4_1(.din(w_dff_B_1irRMUgK8_1),.dout(w_dff_B_KABtyeGH4_1),.clk(gclk));
	jdff dff_B_OuEdJBBJ2_1(.din(w_dff_B_KABtyeGH4_1),.dout(w_dff_B_OuEdJBBJ2_1),.clk(gclk));
	jdff dff_B_s25cA4pm4_1(.din(w_dff_B_OuEdJBBJ2_1),.dout(w_dff_B_s25cA4pm4_1),.clk(gclk));
	jdff dff_B_On2QhlCc3_1(.din(w_dff_B_s25cA4pm4_1),.dout(w_dff_B_On2QhlCc3_1),.clk(gclk));
	jdff dff_B_WgDPmVKq6_1(.din(w_dff_B_On2QhlCc3_1),.dout(w_dff_B_WgDPmVKq6_1),.clk(gclk));
	jdff dff_B_oespMl3E3_1(.din(w_dff_B_WgDPmVKq6_1),.dout(w_dff_B_oespMl3E3_1),.clk(gclk));
	jdff dff_B_JtFFY2kH1_1(.din(w_dff_B_oespMl3E3_1),.dout(w_dff_B_JtFFY2kH1_1),.clk(gclk));
	jdff dff_B_Ywq9y5Pz7_1(.din(w_dff_B_JtFFY2kH1_1),.dout(w_dff_B_Ywq9y5Pz7_1),.clk(gclk));
	jdff dff_B_ShCw1KZ54_1(.din(w_dff_B_Ywq9y5Pz7_1),.dout(w_dff_B_ShCw1KZ54_1),.clk(gclk));
	jdff dff_B_I1gBqC4w6_1(.din(w_dff_B_ShCw1KZ54_1),.dout(w_dff_B_I1gBqC4w6_1),.clk(gclk));
	jdff dff_B_M9LTqsTF1_1(.din(w_dff_B_I1gBqC4w6_1),.dout(w_dff_B_M9LTqsTF1_1),.clk(gclk));
	jdff dff_B_rTrhKZFH4_1(.din(w_dff_B_M9LTqsTF1_1),.dout(w_dff_B_rTrhKZFH4_1),.clk(gclk));
	jdff dff_B_3C1foqNi2_1(.din(w_dff_B_rTrhKZFH4_1),.dout(w_dff_B_3C1foqNi2_1),.clk(gclk));
	jdff dff_B_6gFS1gOo3_1(.din(w_dff_B_3C1foqNi2_1),.dout(w_dff_B_6gFS1gOo3_1),.clk(gclk));
	jdff dff_B_shiMa7fG2_1(.din(w_dff_B_6gFS1gOo3_1),.dout(w_dff_B_shiMa7fG2_1),.clk(gclk));
	jdff dff_B_rVLoYAcl3_1(.din(w_dff_B_shiMa7fG2_1),.dout(w_dff_B_rVLoYAcl3_1),.clk(gclk));
	jdff dff_B_no7Scwuv7_1(.din(w_dff_B_rVLoYAcl3_1),.dout(w_dff_B_no7Scwuv7_1),.clk(gclk));
	jdff dff_B_EiUnT0Xk6_1(.din(w_dff_B_no7Scwuv7_1),.dout(w_dff_B_EiUnT0Xk6_1),.clk(gclk));
	jdff dff_B_gMfcn3ey0_1(.din(w_dff_B_EiUnT0Xk6_1),.dout(w_dff_B_gMfcn3ey0_1),.clk(gclk));
	jdff dff_B_ZJad3ImK8_1(.din(w_dff_B_gMfcn3ey0_1),.dout(w_dff_B_ZJad3ImK8_1),.clk(gclk));
	jdff dff_B_Zx9Qqb762_1(.din(w_dff_B_ZJad3ImK8_1),.dout(w_dff_B_Zx9Qqb762_1),.clk(gclk));
	jdff dff_B_aFJm5bRw2_1(.din(w_dff_B_Zx9Qqb762_1),.dout(w_dff_B_aFJm5bRw2_1),.clk(gclk));
	jdff dff_B_OPZyebUE7_1(.din(w_dff_B_aFJm5bRw2_1),.dout(w_dff_B_OPZyebUE7_1),.clk(gclk));
	jdff dff_B_1dzxiVp58_1(.din(w_dff_B_OPZyebUE7_1),.dout(w_dff_B_1dzxiVp58_1),.clk(gclk));
	jdff dff_B_xz3eF4Kt5_1(.din(w_dff_B_1dzxiVp58_1),.dout(w_dff_B_xz3eF4Kt5_1),.clk(gclk));
	jdff dff_B_1ISlxlMM6_1(.din(w_dff_B_xz3eF4Kt5_1),.dout(w_dff_B_1ISlxlMM6_1),.clk(gclk));
	jdff dff_B_fUyMmErb8_1(.din(w_dff_B_1ISlxlMM6_1),.dout(w_dff_B_fUyMmErb8_1),.clk(gclk));
	jdff dff_B_IqkULnpB5_1(.din(w_dff_B_fUyMmErb8_1),.dout(w_dff_B_IqkULnpB5_1),.clk(gclk));
	jdff dff_B_UvgY0M8H1_1(.din(w_dff_B_IqkULnpB5_1),.dout(w_dff_B_UvgY0M8H1_1),.clk(gclk));
	jdff dff_B_21IILwOy6_1(.din(w_dff_B_UvgY0M8H1_1),.dout(w_dff_B_21IILwOy6_1),.clk(gclk));
	jdff dff_B_JpGOYLhV7_1(.din(w_dff_B_21IILwOy6_1),.dout(w_dff_B_JpGOYLhV7_1),.clk(gclk));
	jdff dff_B_kNQKgbCZ1_1(.din(w_dff_B_JpGOYLhV7_1),.dout(w_dff_B_kNQKgbCZ1_1),.clk(gclk));
	jdff dff_B_x22SxgCY9_1(.din(w_dff_B_kNQKgbCZ1_1),.dout(w_dff_B_x22SxgCY9_1),.clk(gclk));
	jdff dff_B_qnhqOrjf0_1(.din(w_dff_B_x22SxgCY9_1),.dout(w_dff_B_qnhqOrjf0_1),.clk(gclk));
	jdff dff_B_nW3xrQnc4_1(.din(w_dff_B_qnhqOrjf0_1),.dout(w_dff_B_nW3xrQnc4_1),.clk(gclk));
	jdff dff_B_yil0NI7m4_1(.din(w_dff_B_nW3xrQnc4_1),.dout(w_dff_B_yil0NI7m4_1),.clk(gclk));
	jdff dff_B_ViHlSzoC8_1(.din(w_dff_B_yil0NI7m4_1),.dout(w_dff_B_ViHlSzoC8_1),.clk(gclk));
	jdff dff_B_SHNQ3Gih2_1(.din(w_dff_B_ViHlSzoC8_1),.dout(w_dff_B_SHNQ3Gih2_1),.clk(gclk));
	jdff dff_B_WBZVi2Sp6_1(.din(w_dff_B_SHNQ3Gih2_1),.dout(w_dff_B_WBZVi2Sp6_1),.clk(gclk));
	jdff dff_B_fhZXCH4n9_1(.din(w_dff_B_WBZVi2Sp6_1),.dout(w_dff_B_fhZXCH4n9_1),.clk(gclk));
	jdff dff_B_OxdEpg1X7_1(.din(w_dff_B_fhZXCH4n9_1),.dout(w_dff_B_OxdEpg1X7_1),.clk(gclk));
	jdff dff_B_rTh80AY43_1(.din(w_dff_B_OxdEpg1X7_1),.dout(w_dff_B_rTh80AY43_1),.clk(gclk));
	jdff dff_B_KCrW0SRh0_1(.din(w_dff_B_rTh80AY43_1),.dout(w_dff_B_KCrW0SRh0_1),.clk(gclk));
	jdff dff_B_4SdYkNW89_1(.din(w_dff_B_KCrW0SRh0_1),.dout(w_dff_B_4SdYkNW89_1),.clk(gclk));
	jdff dff_B_rQo4x9RC5_1(.din(w_dff_B_4SdYkNW89_1),.dout(w_dff_B_rQo4x9RC5_1),.clk(gclk));
	jdff dff_B_4Y1khT4L6_1(.din(w_dff_B_rQo4x9RC5_1),.dout(w_dff_B_4Y1khT4L6_1),.clk(gclk));
	jdff dff_B_uvutIR678_1(.din(w_dff_B_4Y1khT4L6_1),.dout(w_dff_B_uvutIR678_1),.clk(gclk));
	jdff dff_B_igaI8JiZ5_1(.din(w_dff_B_uvutIR678_1),.dout(w_dff_B_igaI8JiZ5_1),.clk(gclk));
	jdff dff_B_SOzl5xTF5_1(.din(w_dff_B_igaI8JiZ5_1),.dout(w_dff_B_SOzl5xTF5_1),.clk(gclk));
	jdff dff_B_IxxP0Bnh6_1(.din(w_dff_B_SOzl5xTF5_1),.dout(w_dff_B_IxxP0Bnh6_1),.clk(gclk));
	jdff dff_B_kXPR3RWX8_1(.din(w_dff_B_IxxP0Bnh6_1),.dout(w_dff_B_kXPR3RWX8_1),.clk(gclk));
	jdff dff_B_pF9ZeJ1X1_1(.din(w_dff_B_kXPR3RWX8_1),.dout(w_dff_B_pF9ZeJ1X1_1),.clk(gclk));
	jdff dff_B_Q7o9wOw31_1(.din(w_dff_B_pF9ZeJ1X1_1),.dout(w_dff_B_Q7o9wOw31_1),.clk(gclk));
	jdff dff_B_zUheRpOz1_1(.din(w_dff_B_Q7o9wOw31_1),.dout(w_dff_B_zUheRpOz1_1),.clk(gclk));
	jdff dff_B_tlrv0vL40_1(.din(w_dff_B_zUheRpOz1_1),.dout(w_dff_B_tlrv0vL40_1),.clk(gclk));
	jdff dff_B_3vKfztKj3_1(.din(w_dff_B_tlrv0vL40_1),.dout(w_dff_B_3vKfztKj3_1),.clk(gclk));
	jdff dff_B_lNyLmvjt8_1(.din(w_dff_B_3vKfztKj3_1),.dout(w_dff_B_lNyLmvjt8_1),.clk(gclk));
	jdff dff_B_EFXnHh7B1_1(.din(w_dff_B_lNyLmvjt8_1),.dout(w_dff_B_EFXnHh7B1_1),.clk(gclk));
	jdff dff_B_hJto8FeZ3_1(.din(w_dff_B_EFXnHh7B1_1),.dout(w_dff_B_hJto8FeZ3_1),.clk(gclk));
	jdff dff_B_YJbujVQj7_1(.din(w_dff_B_hJto8FeZ3_1),.dout(w_dff_B_YJbujVQj7_1),.clk(gclk));
	jdff dff_B_wcygeEKr6_1(.din(w_dff_B_YJbujVQj7_1),.dout(w_dff_B_wcygeEKr6_1),.clk(gclk));
	jdff dff_B_EmmdnPCY9_1(.din(w_dff_B_wcygeEKr6_1),.dout(w_dff_B_EmmdnPCY9_1),.clk(gclk));
	jdff dff_B_5W2tTDgZ9_1(.din(w_dff_B_EmmdnPCY9_1),.dout(w_dff_B_5W2tTDgZ9_1),.clk(gclk));
	jdff dff_B_iAO25kjD1_1(.din(w_dff_B_5W2tTDgZ9_1),.dout(w_dff_B_iAO25kjD1_1),.clk(gclk));
	jdff dff_B_mK9JxwEz8_1(.din(w_dff_B_iAO25kjD1_1),.dout(w_dff_B_mK9JxwEz8_1),.clk(gclk));
	jdff dff_B_bLpnqNvP2_1(.din(w_dff_B_mK9JxwEz8_1),.dout(w_dff_B_bLpnqNvP2_1),.clk(gclk));
	jdff dff_B_yDw2jqZu1_1(.din(w_dff_B_bLpnqNvP2_1),.dout(w_dff_B_yDw2jqZu1_1),.clk(gclk));
	jdff dff_B_zNwX4zva2_1(.din(w_dff_B_yDw2jqZu1_1),.dout(w_dff_B_zNwX4zva2_1),.clk(gclk));
	jdff dff_B_jd7v22GO3_1(.din(w_dff_B_zNwX4zva2_1),.dout(w_dff_B_jd7v22GO3_1),.clk(gclk));
	jdff dff_B_GAORwh6C2_1(.din(w_dff_B_jd7v22GO3_1),.dout(w_dff_B_GAORwh6C2_1),.clk(gclk));
	jdff dff_B_EFQ4ScXG5_1(.din(w_dff_B_GAORwh6C2_1),.dout(w_dff_B_EFQ4ScXG5_1),.clk(gclk));
	jdff dff_B_b6GgD02e2_1(.din(w_dff_B_EFQ4ScXG5_1),.dout(w_dff_B_b6GgD02e2_1),.clk(gclk));
	jdff dff_B_MManmxoV8_1(.din(w_dff_B_b6GgD02e2_1),.dout(w_dff_B_MManmxoV8_1),.clk(gclk));
	jdff dff_B_iqZtTlaH8_1(.din(w_dff_B_MManmxoV8_1),.dout(w_dff_B_iqZtTlaH8_1),.clk(gclk));
	jdff dff_B_8WEQ1V9L1_1(.din(w_dff_B_iqZtTlaH8_1),.dout(w_dff_B_8WEQ1V9L1_1),.clk(gclk));
	jdff dff_B_srh5O0R77_1(.din(w_dff_B_8WEQ1V9L1_1),.dout(w_dff_B_srh5O0R77_1),.clk(gclk));
	jdff dff_B_iMUG4Dhp3_1(.din(w_dff_B_srh5O0R77_1),.dout(w_dff_B_iMUG4Dhp3_1),.clk(gclk));
	jdff dff_B_8u58h2Jp6_1(.din(w_dff_B_iMUG4Dhp3_1),.dout(w_dff_B_8u58h2Jp6_1),.clk(gclk));
	jdff dff_B_KPr0hUaE8_1(.din(w_dff_B_8u58h2Jp6_1),.dout(w_dff_B_KPr0hUaE8_1),.clk(gclk));
	jdff dff_B_nbLOdoHx7_1(.din(w_dff_B_KPr0hUaE8_1),.dout(w_dff_B_nbLOdoHx7_1),.clk(gclk));
	jdff dff_B_vyLBmnSz8_1(.din(w_dff_B_nbLOdoHx7_1),.dout(w_dff_B_vyLBmnSz8_1),.clk(gclk));
	jdff dff_B_BKCZKVgF8_1(.din(w_dff_B_vyLBmnSz8_1),.dout(w_dff_B_BKCZKVgF8_1),.clk(gclk));
	jdff dff_B_K6ApCmot7_1(.din(w_dff_B_BKCZKVgF8_1),.dout(w_dff_B_K6ApCmot7_1),.clk(gclk));
	jdff dff_B_CIxcN1lw0_1(.din(w_dff_B_K6ApCmot7_1),.dout(w_dff_B_CIxcN1lw0_1),.clk(gclk));
	jdff dff_B_XCbllKuC4_1(.din(w_dff_B_CIxcN1lw0_1),.dout(w_dff_B_XCbllKuC4_1),.clk(gclk));
	jdff dff_B_iMNuduJf2_1(.din(w_dff_B_XCbllKuC4_1),.dout(w_dff_B_iMNuduJf2_1),.clk(gclk));
	jdff dff_B_h9sZE2aB1_1(.din(w_dff_B_iMNuduJf2_1),.dout(w_dff_B_h9sZE2aB1_1),.clk(gclk));
	jdff dff_B_u3sIVnAp9_1(.din(w_dff_B_h9sZE2aB1_1),.dout(w_dff_B_u3sIVnAp9_1),.clk(gclk));
	jdff dff_B_0GqivLDO1_1(.din(w_dff_B_u3sIVnAp9_1),.dout(w_dff_B_0GqivLDO1_1),.clk(gclk));
	jdff dff_B_JSLl1Kq75_1(.din(w_dff_B_0GqivLDO1_1),.dout(w_dff_B_JSLl1Kq75_1),.clk(gclk));
	jdff dff_B_Po7J7QsB6_1(.din(w_dff_B_JSLl1Kq75_1),.dout(w_dff_B_Po7J7QsB6_1),.clk(gclk));
	jdff dff_B_JLVVm7ep3_1(.din(w_dff_B_Po7J7QsB6_1),.dout(w_dff_B_JLVVm7ep3_1),.clk(gclk));
	jdff dff_B_AsiLObze4_1(.din(w_dff_B_JLVVm7ep3_1),.dout(w_dff_B_AsiLObze4_1),.clk(gclk));
	jdff dff_B_SIE3tkeY9_1(.din(w_dff_B_AsiLObze4_1),.dout(w_dff_B_SIE3tkeY9_1),.clk(gclk));
	jdff dff_B_1PvzNOCJ8_1(.din(w_dff_B_SIE3tkeY9_1),.dout(w_dff_B_1PvzNOCJ8_1),.clk(gclk));
	jdff dff_B_JAPcQGai3_1(.din(w_dff_B_1PvzNOCJ8_1),.dout(w_dff_B_JAPcQGai3_1),.clk(gclk));
	jdff dff_B_r2QWZnGR7_1(.din(w_dff_B_JAPcQGai3_1),.dout(w_dff_B_r2QWZnGR7_1),.clk(gclk));
	jdff dff_B_5GQWkxxL9_1(.din(w_dff_B_r2QWZnGR7_1),.dout(w_dff_B_5GQWkxxL9_1),.clk(gclk));
	jdff dff_B_Q1JYRqwz0_1(.din(w_dff_B_5GQWkxxL9_1),.dout(w_dff_B_Q1JYRqwz0_1),.clk(gclk));
	jdff dff_B_Yc7NSR7p0_1(.din(w_dff_B_Q1JYRqwz0_1),.dout(w_dff_B_Yc7NSR7p0_1),.clk(gclk));
	jdff dff_B_hK4Xk5986_1(.din(w_dff_B_Yc7NSR7p0_1),.dout(w_dff_B_hK4Xk5986_1),.clk(gclk));
	jdff dff_B_mcQ4cN8r2_1(.din(w_dff_B_hK4Xk5986_1),.dout(w_dff_B_mcQ4cN8r2_1),.clk(gclk));
	jdff dff_B_cCB9zJ452_1(.din(w_dff_B_mcQ4cN8r2_1),.dout(w_dff_B_cCB9zJ452_1),.clk(gclk));
	jdff dff_B_3fsHmRIV7_1(.din(w_dff_B_cCB9zJ452_1),.dout(w_dff_B_3fsHmRIV7_1),.clk(gclk));
	jdff dff_B_lXcbVTn96_0(.din(n1057),.dout(w_dff_B_lXcbVTn96_0),.clk(gclk));
	jdff dff_B_EuJsqeSg3_0(.din(w_dff_B_lXcbVTn96_0),.dout(w_dff_B_EuJsqeSg3_0),.clk(gclk));
	jdff dff_B_MJDckVra5_0(.din(w_dff_B_EuJsqeSg3_0),.dout(w_dff_B_MJDckVra5_0),.clk(gclk));
	jdff dff_B_fisQWwGe5_0(.din(w_dff_B_MJDckVra5_0),.dout(w_dff_B_fisQWwGe5_0),.clk(gclk));
	jdff dff_B_BQ24fjm62_0(.din(w_dff_B_fisQWwGe5_0),.dout(w_dff_B_BQ24fjm62_0),.clk(gclk));
	jdff dff_B_lu8MqvrR3_0(.din(w_dff_B_BQ24fjm62_0),.dout(w_dff_B_lu8MqvrR3_0),.clk(gclk));
	jdff dff_B_jB1zSSsy8_0(.din(w_dff_B_lu8MqvrR3_0),.dout(w_dff_B_jB1zSSsy8_0),.clk(gclk));
	jdff dff_B_UjEPFYd52_0(.din(w_dff_B_jB1zSSsy8_0),.dout(w_dff_B_UjEPFYd52_0),.clk(gclk));
	jdff dff_B_HOV4m2ek6_0(.din(w_dff_B_UjEPFYd52_0),.dout(w_dff_B_HOV4m2ek6_0),.clk(gclk));
	jdff dff_B_6CVtGBpH5_0(.din(w_dff_B_HOV4m2ek6_0),.dout(w_dff_B_6CVtGBpH5_0),.clk(gclk));
	jdff dff_B_4aEeEHUi2_0(.din(w_dff_B_6CVtGBpH5_0),.dout(w_dff_B_4aEeEHUi2_0),.clk(gclk));
	jdff dff_B_JU99LIya2_0(.din(w_dff_B_4aEeEHUi2_0),.dout(w_dff_B_JU99LIya2_0),.clk(gclk));
	jdff dff_B_zrv6oWNC5_0(.din(w_dff_B_JU99LIya2_0),.dout(w_dff_B_zrv6oWNC5_0),.clk(gclk));
	jdff dff_B_6Gb5miR04_0(.din(w_dff_B_zrv6oWNC5_0),.dout(w_dff_B_6Gb5miR04_0),.clk(gclk));
	jdff dff_B_5847u9wZ4_0(.din(w_dff_B_6Gb5miR04_0),.dout(w_dff_B_5847u9wZ4_0),.clk(gclk));
	jdff dff_B_1unM9Mx92_0(.din(w_dff_B_5847u9wZ4_0),.dout(w_dff_B_1unM9Mx92_0),.clk(gclk));
	jdff dff_B_iOepQaZo4_0(.din(w_dff_B_1unM9Mx92_0),.dout(w_dff_B_iOepQaZo4_0),.clk(gclk));
	jdff dff_B_rEz9W7s84_0(.din(w_dff_B_iOepQaZo4_0),.dout(w_dff_B_rEz9W7s84_0),.clk(gclk));
	jdff dff_B_uN2cxeDa8_0(.din(w_dff_B_rEz9W7s84_0),.dout(w_dff_B_uN2cxeDa8_0),.clk(gclk));
	jdff dff_B_sctwvjzm9_0(.din(w_dff_B_uN2cxeDa8_0),.dout(w_dff_B_sctwvjzm9_0),.clk(gclk));
	jdff dff_B_adZ2zJHA6_0(.din(w_dff_B_sctwvjzm9_0),.dout(w_dff_B_adZ2zJHA6_0),.clk(gclk));
	jdff dff_B_OqUCJmYU8_0(.din(w_dff_B_adZ2zJHA6_0),.dout(w_dff_B_OqUCJmYU8_0),.clk(gclk));
	jdff dff_B_BX3hv6YD1_0(.din(w_dff_B_OqUCJmYU8_0),.dout(w_dff_B_BX3hv6YD1_0),.clk(gclk));
	jdff dff_B_m449Yf9y4_0(.din(w_dff_B_BX3hv6YD1_0),.dout(w_dff_B_m449Yf9y4_0),.clk(gclk));
	jdff dff_B_8EmH85VL8_0(.din(w_dff_B_m449Yf9y4_0),.dout(w_dff_B_8EmH85VL8_0),.clk(gclk));
	jdff dff_B_3uZFVLjP4_0(.din(w_dff_B_8EmH85VL8_0),.dout(w_dff_B_3uZFVLjP4_0),.clk(gclk));
	jdff dff_B_k3wenEl10_0(.din(w_dff_B_3uZFVLjP4_0),.dout(w_dff_B_k3wenEl10_0),.clk(gclk));
	jdff dff_B_v0QZ1dRM0_0(.din(w_dff_B_k3wenEl10_0),.dout(w_dff_B_v0QZ1dRM0_0),.clk(gclk));
	jdff dff_B_U6EboWYB7_0(.din(w_dff_B_v0QZ1dRM0_0),.dout(w_dff_B_U6EboWYB7_0),.clk(gclk));
	jdff dff_B_XJ4iQiS00_0(.din(w_dff_B_U6EboWYB7_0),.dout(w_dff_B_XJ4iQiS00_0),.clk(gclk));
	jdff dff_B_TkPSQJkp3_0(.din(w_dff_B_XJ4iQiS00_0),.dout(w_dff_B_TkPSQJkp3_0),.clk(gclk));
	jdff dff_B_jtbekEci6_0(.din(w_dff_B_TkPSQJkp3_0),.dout(w_dff_B_jtbekEci6_0),.clk(gclk));
	jdff dff_B_i71EgrhA0_0(.din(w_dff_B_jtbekEci6_0),.dout(w_dff_B_i71EgrhA0_0),.clk(gclk));
	jdff dff_B_C9pjuqWt5_0(.din(w_dff_B_i71EgrhA0_0),.dout(w_dff_B_C9pjuqWt5_0),.clk(gclk));
	jdff dff_B_dbes4qhe8_0(.din(w_dff_B_C9pjuqWt5_0),.dout(w_dff_B_dbes4qhe8_0),.clk(gclk));
	jdff dff_B_aMUB5w0v3_0(.din(w_dff_B_dbes4qhe8_0),.dout(w_dff_B_aMUB5w0v3_0),.clk(gclk));
	jdff dff_B_oWn261va5_0(.din(w_dff_B_aMUB5w0v3_0),.dout(w_dff_B_oWn261va5_0),.clk(gclk));
	jdff dff_B_sgTcgaU81_0(.din(w_dff_B_oWn261va5_0),.dout(w_dff_B_sgTcgaU81_0),.clk(gclk));
	jdff dff_B_77tqyWvs1_0(.din(w_dff_B_sgTcgaU81_0),.dout(w_dff_B_77tqyWvs1_0),.clk(gclk));
	jdff dff_B_6APz98kU2_0(.din(w_dff_B_77tqyWvs1_0),.dout(w_dff_B_6APz98kU2_0),.clk(gclk));
	jdff dff_B_TNhIk7Ih1_0(.din(w_dff_B_6APz98kU2_0),.dout(w_dff_B_TNhIk7Ih1_0),.clk(gclk));
	jdff dff_B_cU0C33If0_0(.din(w_dff_B_TNhIk7Ih1_0),.dout(w_dff_B_cU0C33If0_0),.clk(gclk));
	jdff dff_B_yJYmNmdh6_0(.din(w_dff_B_cU0C33If0_0),.dout(w_dff_B_yJYmNmdh6_0),.clk(gclk));
	jdff dff_B_iBtXgot99_0(.din(w_dff_B_yJYmNmdh6_0),.dout(w_dff_B_iBtXgot99_0),.clk(gclk));
	jdff dff_B_u5Mo357n1_0(.din(w_dff_B_iBtXgot99_0),.dout(w_dff_B_u5Mo357n1_0),.clk(gclk));
	jdff dff_B_4DzhqyBu8_0(.din(w_dff_B_u5Mo357n1_0),.dout(w_dff_B_4DzhqyBu8_0),.clk(gclk));
	jdff dff_B_WVUnn1F30_0(.din(w_dff_B_4DzhqyBu8_0),.dout(w_dff_B_WVUnn1F30_0),.clk(gclk));
	jdff dff_B_lprqYsYz7_0(.din(w_dff_B_WVUnn1F30_0),.dout(w_dff_B_lprqYsYz7_0),.clk(gclk));
	jdff dff_B_hl4FJUbS7_0(.din(w_dff_B_lprqYsYz7_0),.dout(w_dff_B_hl4FJUbS7_0),.clk(gclk));
	jdff dff_B_9A3Ssd8G5_0(.din(w_dff_B_hl4FJUbS7_0),.dout(w_dff_B_9A3Ssd8G5_0),.clk(gclk));
	jdff dff_B_G9RerJcH4_0(.din(w_dff_B_9A3Ssd8G5_0),.dout(w_dff_B_G9RerJcH4_0),.clk(gclk));
	jdff dff_B_pLT6T9RD8_0(.din(w_dff_B_G9RerJcH4_0),.dout(w_dff_B_pLT6T9RD8_0),.clk(gclk));
	jdff dff_B_PYAqlhWT4_0(.din(w_dff_B_pLT6T9RD8_0),.dout(w_dff_B_PYAqlhWT4_0),.clk(gclk));
	jdff dff_B_QemTcCs89_0(.din(w_dff_B_PYAqlhWT4_0),.dout(w_dff_B_QemTcCs89_0),.clk(gclk));
	jdff dff_B_3rWWJz0e4_0(.din(w_dff_B_QemTcCs89_0),.dout(w_dff_B_3rWWJz0e4_0),.clk(gclk));
	jdff dff_B_sVnjoQA17_0(.din(w_dff_B_3rWWJz0e4_0),.dout(w_dff_B_sVnjoQA17_0),.clk(gclk));
	jdff dff_B_Ofwh46kp5_0(.din(w_dff_B_sVnjoQA17_0),.dout(w_dff_B_Ofwh46kp5_0),.clk(gclk));
	jdff dff_B_hXscZl9E6_0(.din(w_dff_B_Ofwh46kp5_0),.dout(w_dff_B_hXscZl9E6_0),.clk(gclk));
	jdff dff_B_jWCIsWrH5_0(.din(w_dff_B_hXscZl9E6_0),.dout(w_dff_B_jWCIsWrH5_0),.clk(gclk));
	jdff dff_B_YoOEgNyD2_0(.din(w_dff_B_jWCIsWrH5_0),.dout(w_dff_B_YoOEgNyD2_0),.clk(gclk));
	jdff dff_B_56Jk0nau2_0(.din(w_dff_B_YoOEgNyD2_0),.dout(w_dff_B_56Jk0nau2_0),.clk(gclk));
	jdff dff_B_i0LZErHj4_0(.din(w_dff_B_56Jk0nau2_0),.dout(w_dff_B_i0LZErHj4_0),.clk(gclk));
	jdff dff_B_PFUkBZh20_0(.din(w_dff_B_i0LZErHj4_0),.dout(w_dff_B_PFUkBZh20_0),.clk(gclk));
	jdff dff_B_WEzCsKLz3_0(.din(w_dff_B_PFUkBZh20_0),.dout(w_dff_B_WEzCsKLz3_0),.clk(gclk));
	jdff dff_B_QvVvh4vt2_0(.din(w_dff_B_WEzCsKLz3_0),.dout(w_dff_B_QvVvh4vt2_0),.clk(gclk));
	jdff dff_B_dRo1ao7J4_0(.din(w_dff_B_QvVvh4vt2_0),.dout(w_dff_B_dRo1ao7J4_0),.clk(gclk));
	jdff dff_B_3x7bGVQX6_0(.din(w_dff_B_dRo1ao7J4_0),.dout(w_dff_B_3x7bGVQX6_0),.clk(gclk));
	jdff dff_B_GN6mD94b7_0(.din(w_dff_B_3x7bGVQX6_0),.dout(w_dff_B_GN6mD94b7_0),.clk(gclk));
	jdff dff_B_JrVCeRGC2_0(.din(w_dff_B_GN6mD94b7_0),.dout(w_dff_B_JrVCeRGC2_0),.clk(gclk));
	jdff dff_B_s3qJXBc55_0(.din(w_dff_B_JrVCeRGC2_0),.dout(w_dff_B_s3qJXBc55_0),.clk(gclk));
	jdff dff_B_jjGFx3J51_0(.din(w_dff_B_s3qJXBc55_0),.dout(w_dff_B_jjGFx3J51_0),.clk(gclk));
	jdff dff_B_D5UzCQQy8_0(.din(w_dff_B_jjGFx3J51_0),.dout(w_dff_B_D5UzCQQy8_0),.clk(gclk));
	jdff dff_B_tCqMjmsc2_0(.din(w_dff_B_D5UzCQQy8_0),.dout(w_dff_B_tCqMjmsc2_0),.clk(gclk));
	jdff dff_B_WKO7QTfx5_0(.din(w_dff_B_tCqMjmsc2_0),.dout(w_dff_B_WKO7QTfx5_0),.clk(gclk));
	jdff dff_B_p2rxYZOF2_0(.din(w_dff_B_WKO7QTfx5_0),.dout(w_dff_B_p2rxYZOF2_0),.clk(gclk));
	jdff dff_B_dHDv6ACA9_0(.din(w_dff_B_p2rxYZOF2_0),.dout(w_dff_B_dHDv6ACA9_0),.clk(gclk));
	jdff dff_B_rXzd1AYa1_0(.din(w_dff_B_dHDv6ACA9_0),.dout(w_dff_B_rXzd1AYa1_0),.clk(gclk));
	jdff dff_B_OkYKvnMa5_0(.din(w_dff_B_rXzd1AYa1_0),.dout(w_dff_B_OkYKvnMa5_0),.clk(gclk));
	jdff dff_B_6dTMppZA8_0(.din(w_dff_B_OkYKvnMa5_0),.dout(w_dff_B_6dTMppZA8_0),.clk(gclk));
	jdff dff_B_AOGUaZLi2_0(.din(w_dff_B_6dTMppZA8_0),.dout(w_dff_B_AOGUaZLi2_0),.clk(gclk));
	jdff dff_B_ApRG4ieU7_0(.din(w_dff_B_AOGUaZLi2_0),.dout(w_dff_B_ApRG4ieU7_0),.clk(gclk));
	jdff dff_B_Phgmjnkl1_0(.din(w_dff_B_ApRG4ieU7_0),.dout(w_dff_B_Phgmjnkl1_0),.clk(gclk));
	jdff dff_B_OL8cJkMh9_0(.din(w_dff_B_Phgmjnkl1_0),.dout(w_dff_B_OL8cJkMh9_0),.clk(gclk));
	jdff dff_B_z2bLtqbT5_0(.din(w_dff_B_OL8cJkMh9_0),.dout(w_dff_B_z2bLtqbT5_0),.clk(gclk));
	jdff dff_B_ALr5Fe5X0_0(.din(w_dff_B_z2bLtqbT5_0),.dout(w_dff_B_ALr5Fe5X0_0),.clk(gclk));
	jdff dff_B_ClUh65WD4_0(.din(w_dff_B_ALr5Fe5X0_0),.dout(w_dff_B_ClUh65WD4_0),.clk(gclk));
	jdff dff_B_M2iqKTpG7_0(.din(w_dff_B_ClUh65WD4_0),.dout(w_dff_B_M2iqKTpG7_0),.clk(gclk));
	jdff dff_B_UpJ9WE8l1_0(.din(w_dff_B_M2iqKTpG7_0),.dout(w_dff_B_UpJ9WE8l1_0),.clk(gclk));
	jdff dff_B_lnFB99Bj8_0(.din(w_dff_B_UpJ9WE8l1_0),.dout(w_dff_B_lnFB99Bj8_0),.clk(gclk));
	jdff dff_B_VAiZdZvZ6_0(.din(w_dff_B_lnFB99Bj8_0),.dout(w_dff_B_VAiZdZvZ6_0),.clk(gclk));
	jdff dff_B_KgQSo1s25_0(.din(w_dff_B_VAiZdZvZ6_0),.dout(w_dff_B_KgQSo1s25_0),.clk(gclk));
	jdff dff_B_kJ8if1Rz8_0(.din(w_dff_B_KgQSo1s25_0),.dout(w_dff_B_kJ8if1Rz8_0),.clk(gclk));
	jdff dff_B_aevcQyYO9_0(.din(w_dff_B_kJ8if1Rz8_0),.dout(w_dff_B_aevcQyYO9_0),.clk(gclk));
	jdff dff_B_HkGrW22G5_0(.din(w_dff_B_aevcQyYO9_0),.dout(w_dff_B_HkGrW22G5_0),.clk(gclk));
	jdff dff_B_cPtHhfw96_0(.din(w_dff_B_HkGrW22G5_0),.dout(w_dff_B_cPtHhfw96_0),.clk(gclk));
	jdff dff_B_xMjn9can3_0(.din(w_dff_B_cPtHhfw96_0),.dout(w_dff_B_xMjn9can3_0),.clk(gclk));
	jdff dff_B_qT5hyHnX6_0(.din(w_dff_B_xMjn9can3_0),.dout(w_dff_B_qT5hyHnX6_0),.clk(gclk));
	jdff dff_B_1ivdly6U4_0(.din(w_dff_B_qT5hyHnX6_0),.dout(w_dff_B_1ivdly6U4_0),.clk(gclk));
	jdff dff_B_MlZiuXDQ4_0(.din(w_dff_B_1ivdly6U4_0),.dout(w_dff_B_MlZiuXDQ4_0),.clk(gclk));
	jdff dff_B_waMMDDVc1_0(.din(w_dff_B_MlZiuXDQ4_0),.dout(w_dff_B_waMMDDVc1_0),.clk(gclk));
	jdff dff_B_2CHPNr9c3_0(.din(w_dff_B_waMMDDVc1_0),.dout(w_dff_B_2CHPNr9c3_0),.clk(gclk));
	jdff dff_B_KuGm4Giw7_0(.din(w_dff_B_2CHPNr9c3_0),.dout(w_dff_B_KuGm4Giw7_0),.clk(gclk));
	jdff dff_B_7eOg1sdf3_0(.din(w_dff_B_KuGm4Giw7_0),.dout(w_dff_B_7eOg1sdf3_0),.clk(gclk));
	jdff dff_B_1e0svXtD7_0(.din(w_dff_B_7eOg1sdf3_0),.dout(w_dff_B_1e0svXtD7_0),.clk(gclk));
	jdff dff_B_zqxBeI1X0_0(.din(w_dff_B_1e0svXtD7_0),.dout(w_dff_B_zqxBeI1X0_0),.clk(gclk));
	jdff dff_B_fcgveMbB5_0(.din(w_dff_B_zqxBeI1X0_0),.dout(w_dff_B_fcgveMbB5_0),.clk(gclk));
	jdff dff_B_vHQ6kjWz2_0(.din(w_dff_B_fcgveMbB5_0),.dout(w_dff_B_vHQ6kjWz2_0),.clk(gclk));
	jdff dff_B_phBEkl3m2_0(.din(w_dff_B_vHQ6kjWz2_0),.dout(w_dff_B_phBEkl3m2_0),.clk(gclk));
	jdff dff_B_8wUH5XTf9_0(.din(w_dff_B_phBEkl3m2_0),.dout(w_dff_B_8wUH5XTf9_0),.clk(gclk));
	jdff dff_B_aUAVFcQw1_0(.din(w_dff_B_8wUH5XTf9_0),.dout(w_dff_B_aUAVFcQw1_0),.clk(gclk));
	jdff dff_B_ncmA4MoC6_0(.din(w_dff_B_aUAVFcQw1_0),.dout(w_dff_B_ncmA4MoC6_0),.clk(gclk));
	jdff dff_B_9kk8s8Kj0_0(.din(w_dff_B_ncmA4MoC6_0),.dout(w_dff_B_9kk8s8Kj0_0),.clk(gclk));
	jdff dff_B_f5fJqnrM7_1(.din(n1050),.dout(w_dff_B_f5fJqnrM7_1),.clk(gclk));
	jdff dff_B_SCRBDtFc7_1(.din(w_dff_B_f5fJqnrM7_1),.dout(w_dff_B_SCRBDtFc7_1),.clk(gclk));
	jdff dff_B_kFZcFra90_1(.din(w_dff_B_SCRBDtFc7_1),.dout(w_dff_B_kFZcFra90_1),.clk(gclk));
	jdff dff_B_z9Ief7Ks5_1(.din(w_dff_B_kFZcFra90_1),.dout(w_dff_B_z9Ief7Ks5_1),.clk(gclk));
	jdff dff_B_3ahmI1Xs7_1(.din(w_dff_B_z9Ief7Ks5_1),.dout(w_dff_B_3ahmI1Xs7_1),.clk(gclk));
	jdff dff_B_5AiS494R3_1(.din(w_dff_B_3ahmI1Xs7_1),.dout(w_dff_B_5AiS494R3_1),.clk(gclk));
	jdff dff_B_3WgcX6Ds9_1(.din(w_dff_B_5AiS494R3_1),.dout(w_dff_B_3WgcX6Ds9_1),.clk(gclk));
	jdff dff_B_0NYHveAO2_1(.din(w_dff_B_3WgcX6Ds9_1),.dout(w_dff_B_0NYHveAO2_1),.clk(gclk));
	jdff dff_B_MNNzQLw34_1(.din(w_dff_B_0NYHveAO2_1),.dout(w_dff_B_MNNzQLw34_1),.clk(gclk));
	jdff dff_B_wuIGaYfu8_1(.din(w_dff_B_MNNzQLw34_1),.dout(w_dff_B_wuIGaYfu8_1),.clk(gclk));
	jdff dff_B_ZP15QZ0T1_1(.din(w_dff_B_wuIGaYfu8_1),.dout(w_dff_B_ZP15QZ0T1_1),.clk(gclk));
	jdff dff_B_WTNqxCAK8_1(.din(w_dff_B_ZP15QZ0T1_1),.dout(w_dff_B_WTNqxCAK8_1),.clk(gclk));
	jdff dff_B_x243EKgh1_1(.din(w_dff_B_WTNqxCAK8_1),.dout(w_dff_B_x243EKgh1_1),.clk(gclk));
	jdff dff_B_HbOt34VG0_1(.din(w_dff_B_x243EKgh1_1),.dout(w_dff_B_HbOt34VG0_1),.clk(gclk));
	jdff dff_B_Yn3RuMFN6_1(.din(w_dff_B_HbOt34VG0_1),.dout(w_dff_B_Yn3RuMFN6_1),.clk(gclk));
	jdff dff_B_87KBbj4Y4_1(.din(w_dff_B_Yn3RuMFN6_1),.dout(w_dff_B_87KBbj4Y4_1),.clk(gclk));
	jdff dff_B_4GRhYBde0_1(.din(w_dff_B_87KBbj4Y4_1),.dout(w_dff_B_4GRhYBde0_1),.clk(gclk));
	jdff dff_B_iw1OlsIB4_1(.din(w_dff_B_4GRhYBde0_1),.dout(w_dff_B_iw1OlsIB4_1),.clk(gclk));
	jdff dff_B_p8x0bEBn2_1(.din(w_dff_B_iw1OlsIB4_1),.dout(w_dff_B_p8x0bEBn2_1),.clk(gclk));
	jdff dff_B_O8akJU065_1(.din(w_dff_B_p8x0bEBn2_1),.dout(w_dff_B_O8akJU065_1),.clk(gclk));
	jdff dff_B_xIEFSa847_1(.din(w_dff_B_O8akJU065_1),.dout(w_dff_B_xIEFSa847_1),.clk(gclk));
	jdff dff_B_pXrq6MKO9_1(.din(w_dff_B_xIEFSa847_1),.dout(w_dff_B_pXrq6MKO9_1),.clk(gclk));
	jdff dff_B_xzS58Tau8_1(.din(w_dff_B_pXrq6MKO9_1),.dout(w_dff_B_xzS58Tau8_1),.clk(gclk));
	jdff dff_B_BCZ9PQjd4_1(.din(w_dff_B_xzS58Tau8_1),.dout(w_dff_B_BCZ9PQjd4_1),.clk(gclk));
	jdff dff_B_booaxSNR1_1(.din(w_dff_B_BCZ9PQjd4_1),.dout(w_dff_B_booaxSNR1_1),.clk(gclk));
	jdff dff_B_D1ghgW416_1(.din(w_dff_B_booaxSNR1_1),.dout(w_dff_B_D1ghgW416_1),.clk(gclk));
	jdff dff_B_I0RR89VS4_1(.din(w_dff_B_D1ghgW416_1),.dout(w_dff_B_I0RR89VS4_1),.clk(gclk));
	jdff dff_B_Syn8FOEL2_1(.din(w_dff_B_I0RR89VS4_1),.dout(w_dff_B_Syn8FOEL2_1),.clk(gclk));
	jdff dff_B_tQKZaWqY5_1(.din(w_dff_B_Syn8FOEL2_1),.dout(w_dff_B_tQKZaWqY5_1),.clk(gclk));
	jdff dff_B_KRNn8g490_1(.din(w_dff_B_tQKZaWqY5_1),.dout(w_dff_B_KRNn8g490_1),.clk(gclk));
	jdff dff_B_n4Cih7Cs0_1(.din(w_dff_B_KRNn8g490_1),.dout(w_dff_B_n4Cih7Cs0_1),.clk(gclk));
	jdff dff_B_V8is0NG60_1(.din(w_dff_B_n4Cih7Cs0_1),.dout(w_dff_B_V8is0NG60_1),.clk(gclk));
	jdff dff_B_uCXvTn7W7_1(.din(w_dff_B_V8is0NG60_1),.dout(w_dff_B_uCXvTn7W7_1),.clk(gclk));
	jdff dff_B_DfgfrNC04_1(.din(w_dff_B_uCXvTn7W7_1),.dout(w_dff_B_DfgfrNC04_1),.clk(gclk));
	jdff dff_B_PoDMF17E9_1(.din(w_dff_B_DfgfrNC04_1),.dout(w_dff_B_PoDMF17E9_1),.clk(gclk));
	jdff dff_B_GvWs4D6b5_1(.din(w_dff_B_PoDMF17E9_1),.dout(w_dff_B_GvWs4D6b5_1),.clk(gclk));
	jdff dff_B_jt6GZ1SQ9_1(.din(w_dff_B_GvWs4D6b5_1),.dout(w_dff_B_jt6GZ1SQ9_1),.clk(gclk));
	jdff dff_B_VEjB5MWe7_1(.din(w_dff_B_jt6GZ1SQ9_1),.dout(w_dff_B_VEjB5MWe7_1),.clk(gclk));
	jdff dff_B_JNWa2Hc12_1(.din(w_dff_B_VEjB5MWe7_1),.dout(w_dff_B_JNWa2Hc12_1),.clk(gclk));
	jdff dff_B_YedQTxBc1_1(.din(w_dff_B_JNWa2Hc12_1),.dout(w_dff_B_YedQTxBc1_1),.clk(gclk));
	jdff dff_B_MWVEk7Yy2_1(.din(w_dff_B_YedQTxBc1_1),.dout(w_dff_B_MWVEk7Yy2_1),.clk(gclk));
	jdff dff_B_SGVrIX835_1(.din(w_dff_B_MWVEk7Yy2_1),.dout(w_dff_B_SGVrIX835_1),.clk(gclk));
	jdff dff_B_iViIFdnS5_1(.din(w_dff_B_SGVrIX835_1),.dout(w_dff_B_iViIFdnS5_1),.clk(gclk));
	jdff dff_B_s0cNhQew7_1(.din(w_dff_B_iViIFdnS5_1),.dout(w_dff_B_s0cNhQew7_1),.clk(gclk));
	jdff dff_B_c9Bs7ZZT3_1(.din(w_dff_B_s0cNhQew7_1),.dout(w_dff_B_c9Bs7ZZT3_1),.clk(gclk));
	jdff dff_B_wbRhDBm88_1(.din(w_dff_B_c9Bs7ZZT3_1),.dout(w_dff_B_wbRhDBm88_1),.clk(gclk));
	jdff dff_B_9iNe9YHu5_1(.din(w_dff_B_wbRhDBm88_1),.dout(w_dff_B_9iNe9YHu5_1),.clk(gclk));
	jdff dff_B_AjXH0r3u6_1(.din(w_dff_B_9iNe9YHu5_1),.dout(w_dff_B_AjXH0r3u6_1),.clk(gclk));
	jdff dff_B_thVnRWrT7_1(.din(w_dff_B_AjXH0r3u6_1),.dout(w_dff_B_thVnRWrT7_1),.clk(gclk));
	jdff dff_B_0PTJ0m2x9_1(.din(w_dff_B_thVnRWrT7_1),.dout(w_dff_B_0PTJ0m2x9_1),.clk(gclk));
	jdff dff_B_x67HYtzZ6_1(.din(w_dff_B_0PTJ0m2x9_1),.dout(w_dff_B_x67HYtzZ6_1),.clk(gclk));
	jdff dff_B_Wyg9oLko4_1(.din(w_dff_B_x67HYtzZ6_1),.dout(w_dff_B_Wyg9oLko4_1),.clk(gclk));
	jdff dff_B_m7XQnY6f9_1(.din(w_dff_B_Wyg9oLko4_1),.dout(w_dff_B_m7XQnY6f9_1),.clk(gclk));
	jdff dff_B_86GG1ANT4_1(.din(w_dff_B_m7XQnY6f9_1),.dout(w_dff_B_86GG1ANT4_1),.clk(gclk));
	jdff dff_B_fn7ngN5V4_1(.din(w_dff_B_86GG1ANT4_1),.dout(w_dff_B_fn7ngN5V4_1),.clk(gclk));
	jdff dff_B_0NQxYXRW8_1(.din(w_dff_B_fn7ngN5V4_1),.dout(w_dff_B_0NQxYXRW8_1),.clk(gclk));
	jdff dff_B_dJdFIWHo0_1(.din(w_dff_B_0NQxYXRW8_1),.dout(w_dff_B_dJdFIWHo0_1),.clk(gclk));
	jdff dff_B_z9XltW5J7_1(.din(w_dff_B_dJdFIWHo0_1),.dout(w_dff_B_z9XltW5J7_1),.clk(gclk));
	jdff dff_B_3mqeqZlv1_1(.din(w_dff_B_z9XltW5J7_1),.dout(w_dff_B_3mqeqZlv1_1),.clk(gclk));
	jdff dff_B_0ZoUOAI12_1(.din(w_dff_B_3mqeqZlv1_1),.dout(w_dff_B_0ZoUOAI12_1),.clk(gclk));
	jdff dff_B_VsP0cSah0_1(.din(w_dff_B_0ZoUOAI12_1),.dout(w_dff_B_VsP0cSah0_1),.clk(gclk));
	jdff dff_B_JcEcZDWL8_1(.din(w_dff_B_VsP0cSah0_1),.dout(w_dff_B_JcEcZDWL8_1),.clk(gclk));
	jdff dff_B_krdChQNe4_1(.din(w_dff_B_JcEcZDWL8_1),.dout(w_dff_B_krdChQNe4_1),.clk(gclk));
	jdff dff_B_MZqqAY5K4_1(.din(w_dff_B_krdChQNe4_1),.dout(w_dff_B_MZqqAY5K4_1),.clk(gclk));
	jdff dff_B_iOZ3gROo8_1(.din(w_dff_B_MZqqAY5K4_1),.dout(w_dff_B_iOZ3gROo8_1),.clk(gclk));
	jdff dff_B_92w27m5X0_1(.din(w_dff_B_iOZ3gROo8_1),.dout(w_dff_B_92w27m5X0_1),.clk(gclk));
	jdff dff_B_ZglMHgYd9_1(.din(w_dff_B_92w27m5X0_1),.dout(w_dff_B_ZglMHgYd9_1),.clk(gclk));
	jdff dff_B_PbFPI6Fe5_1(.din(w_dff_B_ZglMHgYd9_1),.dout(w_dff_B_PbFPI6Fe5_1),.clk(gclk));
	jdff dff_B_jchvVAJs1_1(.din(w_dff_B_PbFPI6Fe5_1),.dout(w_dff_B_jchvVAJs1_1),.clk(gclk));
	jdff dff_B_1DlG3P9Z6_1(.din(w_dff_B_jchvVAJs1_1),.dout(w_dff_B_1DlG3P9Z6_1),.clk(gclk));
	jdff dff_B_dNz23Tyv9_1(.din(w_dff_B_1DlG3P9Z6_1),.dout(w_dff_B_dNz23Tyv9_1),.clk(gclk));
	jdff dff_B_E7DbAjSu7_1(.din(w_dff_B_dNz23Tyv9_1),.dout(w_dff_B_E7DbAjSu7_1),.clk(gclk));
	jdff dff_B_eHpZEKlY6_1(.din(w_dff_B_E7DbAjSu7_1),.dout(w_dff_B_eHpZEKlY6_1),.clk(gclk));
	jdff dff_B_Qj8FgEmd8_1(.din(w_dff_B_eHpZEKlY6_1),.dout(w_dff_B_Qj8FgEmd8_1),.clk(gclk));
	jdff dff_B_XnaP1RXz3_1(.din(w_dff_B_Qj8FgEmd8_1),.dout(w_dff_B_XnaP1RXz3_1),.clk(gclk));
	jdff dff_B_Jucbebss1_1(.din(w_dff_B_XnaP1RXz3_1),.dout(w_dff_B_Jucbebss1_1),.clk(gclk));
	jdff dff_B_EYBMdIFj3_1(.din(w_dff_B_Jucbebss1_1),.dout(w_dff_B_EYBMdIFj3_1),.clk(gclk));
	jdff dff_B_gwICwd4J7_1(.din(w_dff_B_EYBMdIFj3_1),.dout(w_dff_B_gwICwd4J7_1),.clk(gclk));
	jdff dff_B_hEZ8aKD22_1(.din(w_dff_B_gwICwd4J7_1),.dout(w_dff_B_hEZ8aKD22_1),.clk(gclk));
	jdff dff_B_68lFFIXZ4_1(.din(w_dff_B_hEZ8aKD22_1),.dout(w_dff_B_68lFFIXZ4_1),.clk(gclk));
	jdff dff_B_w4VXy8Sb4_1(.din(w_dff_B_68lFFIXZ4_1),.dout(w_dff_B_w4VXy8Sb4_1),.clk(gclk));
	jdff dff_B_ny3alXd71_1(.din(w_dff_B_w4VXy8Sb4_1),.dout(w_dff_B_ny3alXd71_1),.clk(gclk));
	jdff dff_B_MSi1KQ8d1_1(.din(w_dff_B_ny3alXd71_1),.dout(w_dff_B_MSi1KQ8d1_1),.clk(gclk));
	jdff dff_B_HIsATejX5_1(.din(w_dff_B_MSi1KQ8d1_1),.dout(w_dff_B_HIsATejX5_1),.clk(gclk));
	jdff dff_B_EFcE9LzN3_1(.din(w_dff_B_HIsATejX5_1),.dout(w_dff_B_EFcE9LzN3_1),.clk(gclk));
	jdff dff_B_r09dneTc2_1(.din(w_dff_B_EFcE9LzN3_1),.dout(w_dff_B_r09dneTc2_1),.clk(gclk));
	jdff dff_B_oOjE5vBU7_1(.din(w_dff_B_r09dneTc2_1),.dout(w_dff_B_oOjE5vBU7_1),.clk(gclk));
	jdff dff_B_SVsaNuYL0_1(.din(w_dff_B_oOjE5vBU7_1),.dout(w_dff_B_SVsaNuYL0_1),.clk(gclk));
	jdff dff_B_QUH1PpSS8_1(.din(w_dff_B_SVsaNuYL0_1),.dout(w_dff_B_QUH1PpSS8_1),.clk(gclk));
	jdff dff_B_bMwO5Ksz5_1(.din(w_dff_B_QUH1PpSS8_1),.dout(w_dff_B_bMwO5Ksz5_1),.clk(gclk));
	jdff dff_B_FatS89pc5_1(.din(w_dff_B_bMwO5Ksz5_1),.dout(w_dff_B_FatS89pc5_1),.clk(gclk));
	jdff dff_B_GbeDqxmI8_1(.din(w_dff_B_FatS89pc5_1),.dout(w_dff_B_GbeDqxmI8_1),.clk(gclk));
	jdff dff_B_NOPoR7ZS0_1(.din(w_dff_B_GbeDqxmI8_1),.dout(w_dff_B_NOPoR7ZS0_1),.clk(gclk));
	jdff dff_B_rgwx18Bc2_1(.din(w_dff_B_NOPoR7ZS0_1),.dout(w_dff_B_rgwx18Bc2_1),.clk(gclk));
	jdff dff_B_mEZrt6z78_1(.din(w_dff_B_rgwx18Bc2_1),.dout(w_dff_B_mEZrt6z78_1),.clk(gclk));
	jdff dff_B_PgCb1xBM1_1(.din(w_dff_B_mEZrt6z78_1),.dout(w_dff_B_PgCb1xBM1_1),.clk(gclk));
	jdff dff_B_gGE28DBO2_1(.din(w_dff_B_PgCb1xBM1_1),.dout(w_dff_B_gGE28DBO2_1),.clk(gclk));
	jdff dff_B_9xckHE418_1(.din(w_dff_B_gGE28DBO2_1),.dout(w_dff_B_9xckHE418_1),.clk(gclk));
	jdff dff_B_LHB3u8c70_1(.din(w_dff_B_9xckHE418_1),.dout(w_dff_B_LHB3u8c70_1),.clk(gclk));
	jdff dff_B_DZ6NZwNS8_1(.din(w_dff_B_LHB3u8c70_1),.dout(w_dff_B_DZ6NZwNS8_1),.clk(gclk));
	jdff dff_B_PMS6C3Ib7_1(.din(w_dff_B_DZ6NZwNS8_1),.dout(w_dff_B_PMS6C3Ib7_1),.clk(gclk));
	jdff dff_B_Y81h77nn0_1(.din(w_dff_B_PMS6C3Ib7_1),.dout(w_dff_B_Y81h77nn0_1),.clk(gclk));
	jdff dff_B_YKDPraiS0_1(.din(w_dff_B_Y81h77nn0_1),.dout(w_dff_B_YKDPraiS0_1),.clk(gclk));
	jdff dff_B_dI7R08Xx1_1(.din(w_dff_B_YKDPraiS0_1),.dout(w_dff_B_dI7R08Xx1_1),.clk(gclk));
	jdff dff_B_TNs070wt2_1(.din(w_dff_B_dI7R08Xx1_1),.dout(w_dff_B_TNs070wt2_1),.clk(gclk));
	jdff dff_B_9kifPkEd3_1(.din(w_dff_B_TNs070wt2_1),.dout(w_dff_B_9kifPkEd3_1),.clk(gclk));
	jdff dff_B_Ss2Uaxdz6_1(.din(w_dff_B_9kifPkEd3_1),.dout(w_dff_B_Ss2Uaxdz6_1),.clk(gclk));
	jdff dff_B_vm75blfX0_1(.din(w_dff_B_Ss2Uaxdz6_1),.dout(w_dff_B_vm75blfX0_1),.clk(gclk));
	jdff dff_B_2X6D9LyI9_1(.din(w_dff_B_vm75blfX0_1),.dout(w_dff_B_2X6D9LyI9_1),.clk(gclk));
	jdff dff_B_3ncbrnNb2_1(.din(w_dff_B_2X6D9LyI9_1),.dout(w_dff_B_3ncbrnNb2_1),.clk(gclk));
	jdff dff_B_7nEsIUQP7_1(.din(w_dff_B_3ncbrnNb2_1),.dout(w_dff_B_7nEsIUQP7_1),.clk(gclk));
	jdff dff_B_vh99L45W1_0(.din(n1051),.dout(w_dff_B_vh99L45W1_0),.clk(gclk));
	jdff dff_B_WpPMkpzG4_0(.din(w_dff_B_vh99L45W1_0),.dout(w_dff_B_WpPMkpzG4_0),.clk(gclk));
	jdff dff_B_Q6ZTjjX75_0(.din(w_dff_B_WpPMkpzG4_0),.dout(w_dff_B_Q6ZTjjX75_0),.clk(gclk));
	jdff dff_B_xKamv6vY8_0(.din(w_dff_B_Q6ZTjjX75_0),.dout(w_dff_B_xKamv6vY8_0),.clk(gclk));
	jdff dff_B_VCua7QkI4_0(.din(w_dff_B_xKamv6vY8_0),.dout(w_dff_B_VCua7QkI4_0),.clk(gclk));
	jdff dff_B_oxsb2J787_0(.din(w_dff_B_VCua7QkI4_0),.dout(w_dff_B_oxsb2J787_0),.clk(gclk));
	jdff dff_B_9u38LOqB5_0(.din(w_dff_B_oxsb2J787_0),.dout(w_dff_B_9u38LOqB5_0),.clk(gclk));
	jdff dff_B_loVxnU1V7_0(.din(w_dff_B_9u38LOqB5_0),.dout(w_dff_B_loVxnU1V7_0),.clk(gclk));
	jdff dff_B_scLkIwhk8_0(.din(w_dff_B_loVxnU1V7_0),.dout(w_dff_B_scLkIwhk8_0),.clk(gclk));
	jdff dff_B_18gcbKV37_0(.din(w_dff_B_scLkIwhk8_0),.dout(w_dff_B_18gcbKV37_0),.clk(gclk));
	jdff dff_B_jBeGjqSL4_0(.din(w_dff_B_18gcbKV37_0),.dout(w_dff_B_jBeGjqSL4_0),.clk(gclk));
	jdff dff_B_LucZaYKp2_0(.din(w_dff_B_jBeGjqSL4_0),.dout(w_dff_B_LucZaYKp2_0),.clk(gclk));
	jdff dff_B_f1DNbYTn6_0(.din(w_dff_B_LucZaYKp2_0),.dout(w_dff_B_f1DNbYTn6_0),.clk(gclk));
	jdff dff_B_DjVneDZu7_0(.din(w_dff_B_f1DNbYTn6_0),.dout(w_dff_B_DjVneDZu7_0),.clk(gclk));
	jdff dff_B_HRpiISse9_0(.din(w_dff_B_DjVneDZu7_0),.dout(w_dff_B_HRpiISse9_0),.clk(gclk));
	jdff dff_B_DsmGcOrD9_0(.din(w_dff_B_HRpiISse9_0),.dout(w_dff_B_DsmGcOrD9_0),.clk(gclk));
	jdff dff_B_gnlDjTcb3_0(.din(w_dff_B_DsmGcOrD9_0),.dout(w_dff_B_gnlDjTcb3_0),.clk(gclk));
	jdff dff_B_Ns3pgPzD7_0(.din(w_dff_B_gnlDjTcb3_0),.dout(w_dff_B_Ns3pgPzD7_0),.clk(gclk));
	jdff dff_B_oMCrHf1M1_0(.din(w_dff_B_Ns3pgPzD7_0),.dout(w_dff_B_oMCrHf1M1_0),.clk(gclk));
	jdff dff_B_WaEEoS817_0(.din(w_dff_B_oMCrHf1M1_0),.dout(w_dff_B_WaEEoS817_0),.clk(gclk));
	jdff dff_B_JJ8F5yyf2_0(.din(w_dff_B_WaEEoS817_0),.dout(w_dff_B_JJ8F5yyf2_0),.clk(gclk));
	jdff dff_B_8pAQ3Lj87_0(.din(w_dff_B_JJ8F5yyf2_0),.dout(w_dff_B_8pAQ3Lj87_0),.clk(gclk));
	jdff dff_B_atqK1YFV5_0(.din(w_dff_B_8pAQ3Lj87_0),.dout(w_dff_B_atqK1YFV5_0),.clk(gclk));
	jdff dff_B_jzaHvS473_0(.din(w_dff_B_atqK1YFV5_0),.dout(w_dff_B_jzaHvS473_0),.clk(gclk));
	jdff dff_B_Mr5QEqgj0_0(.din(w_dff_B_jzaHvS473_0),.dout(w_dff_B_Mr5QEqgj0_0),.clk(gclk));
	jdff dff_B_fR3Luis86_0(.din(w_dff_B_Mr5QEqgj0_0),.dout(w_dff_B_fR3Luis86_0),.clk(gclk));
	jdff dff_B_XbWQcGBV3_0(.din(w_dff_B_fR3Luis86_0),.dout(w_dff_B_XbWQcGBV3_0),.clk(gclk));
	jdff dff_B_hfM7cqph0_0(.din(w_dff_B_XbWQcGBV3_0),.dout(w_dff_B_hfM7cqph0_0),.clk(gclk));
	jdff dff_B_303QQDhd6_0(.din(w_dff_B_hfM7cqph0_0),.dout(w_dff_B_303QQDhd6_0),.clk(gclk));
	jdff dff_B_RCfuaQTD0_0(.din(w_dff_B_303QQDhd6_0),.dout(w_dff_B_RCfuaQTD0_0),.clk(gclk));
	jdff dff_B_Kt9M91KE3_0(.din(w_dff_B_RCfuaQTD0_0),.dout(w_dff_B_Kt9M91KE3_0),.clk(gclk));
	jdff dff_B_KbOef6La6_0(.din(w_dff_B_Kt9M91KE3_0),.dout(w_dff_B_KbOef6La6_0),.clk(gclk));
	jdff dff_B_hLPLZt4l5_0(.din(w_dff_B_KbOef6La6_0),.dout(w_dff_B_hLPLZt4l5_0),.clk(gclk));
	jdff dff_B_AhxYsQDU0_0(.din(w_dff_B_hLPLZt4l5_0),.dout(w_dff_B_AhxYsQDU0_0),.clk(gclk));
	jdff dff_B_Gg644Uby4_0(.din(w_dff_B_AhxYsQDU0_0),.dout(w_dff_B_Gg644Uby4_0),.clk(gclk));
	jdff dff_B_3Bnn5R344_0(.din(w_dff_B_Gg644Uby4_0),.dout(w_dff_B_3Bnn5R344_0),.clk(gclk));
	jdff dff_B_CqDmdEoC8_0(.din(w_dff_B_3Bnn5R344_0),.dout(w_dff_B_CqDmdEoC8_0),.clk(gclk));
	jdff dff_B_QFhFRcxg6_0(.din(w_dff_B_CqDmdEoC8_0),.dout(w_dff_B_QFhFRcxg6_0),.clk(gclk));
	jdff dff_B_AC1xFoOV4_0(.din(w_dff_B_QFhFRcxg6_0),.dout(w_dff_B_AC1xFoOV4_0),.clk(gclk));
	jdff dff_B_o8P8HGCg4_0(.din(w_dff_B_AC1xFoOV4_0),.dout(w_dff_B_o8P8HGCg4_0),.clk(gclk));
	jdff dff_B_tCCy3xBw1_0(.din(w_dff_B_o8P8HGCg4_0),.dout(w_dff_B_tCCy3xBw1_0),.clk(gclk));
	jdff dff_B_2uK9qrsP1_0(.din(w_dff_B_tCCy3xBw1_0),.dout(w_dff_B_2uK9qrsP1_0),.clk(gclk));
	jdff dff_B_Zu7Qzsol6_0(.din(w_dff_B_2uK9qrsP1_0),.dout(w_dff_B_Zu7Qzsol6_0),.clk(gclk));
	jdff dff_B_LuA8ccpT0_0(.din(w_dff_B_Zu7Qzsol6_0),.dout(w_dff_B_LuA8ccpT0_0),.clk(gclk));
	jdff dff_B_LXIS0KMU6_0(.din(w_dff_B_LuA8ccpT0_0),.dout(w_dff_B_LXIS0KMU6_0),.clk(gclk));
	jdff dff_B_nudrdhfk0_0(.din(w_dff_B_LXIS0KMU6_0),.dout(w_dff_B_nudrdhfk0_0),.clk(gclk));
	jdff dff_B_qaIlPDop6_0(.din(w_dff_B_nudrdhfk0_0),.dout(w_dff_B_qaIlPDop6_0),.clk(gclk));
	jdff dff_B_hzPq7EEo2_0(.din(w_dff_B_qaIlPDop6_0),.dout(w_dff_B_hzPq7EEo2_0),.clk(gclk));
	jdff dff_B_61XcsiEZ2_0(.din(w_dff_B_hzPq7EEo2_0),.dout(w_dff_B_61XcsiEZ2_0),.clk(gclk));
	jdff dff_B_hWMclC1a1_0(.din(w_dff_B_61XcsiEZ2_0),.dout(w_dff_B_hWMclC1a1_0),.clk(gclk));
	jdff dff_B_dPHn03oe7_0(.din(w_dff_B_hWMclC1a1_0),.dout(w_dff_B_dPHn03oe7_0),.clk(gclk));
	jdff dff_B_aTFnL8Uf6_0(.din(w_dff_B_dPHn03oe7_0),.dout(w_dff_B_aTFnL8Uf6_0),.clk(gclk));
	jdff dff_B_l0d8bZ0v1_0(.din(w_dff_B_aTFnL8Uf6_0),.dout(w_dff_B_l0d8bZ0v1_0),.clk(gclk));
	jdff dff_B_HufA5ZQ70_0(.din(w_dff_B_l0d8bZ0v1_0),.dout(w_dff_B_HufA5ZQ70_0),.clk(gclk));
	jdff dff_B_KVVOJQLQ0_0(.din(w_dff_B_HufA5ZQ70_0),.dout(w_dff_B_KVVOJQLQ0_0),.clk(gclk));
	jdff dff_B_bgNzMwST0_0(.din(w_dff_B_KVVOJQLQ0_0),.dout(w_dff_B_bgNzMwST0_0),.clk(gclk));
	jdff dff_B_SlPhwksZ4_0(.din(w_dff_B_bgNzMwST0_0),.dout(w_dff_B_SlPhwksZ4_0),.clk(gclk));
	jdff dff_B_tQrdhgjC0_0(.din(w_dff_B_SlPhwksZ4_0),.dout(w_dff_B_tQrdhgjC0_0),.clk(gclk));
	jdff dff_B_kynfNtjN7_0(.din(w_dff_B_tQrdhgjC0_0),.dout(w_dff_B_kynfNtjN7_0),.clk(gclk));
	jdff dff_B_Y2yw4CJS2_0(.din(w_dff_B_kynfNtjN7_0),.dout(w_dff_B_Y2yw4CJS2_0),.clk(gclk));
	jdff dff_B_DlBbqP5E9_0(.din(w_dff_B_Y2yw4CJS2_0),.dout(w_dff_B_DlBbqP5E9_0),.clk(gclk));
	jdff dff_B_Twf2Fwju5_0(.din(w_dff_B_DlBbqP5E9_0),.dout(w_dff_B_Twf2Fwju5_0),.clk(gclk));
	jdff dff_B_aQaGiu9v3_0(.din(w_dff_B_Twf2Fwju5_0),.dout(w_dff_B_aQaGiu9v3_0),.clk(gclk));
	jdff dff_B_LyVO3kP23_0(.din(w_dff_B_aQaGiu9v3_0),.dout(w_dff_B_LyVO3kP23_0),.clk(gclk));
	jdff dff_B_3fAnSOOd2_0(.din(w_dff_B_LyVO3kP23_0),.dout(w_dff_B_3fAnSOOd2_0),.clk(gclk));
	jdff dff_B_i9OJ2SyL0_0(.din(w_dff_B_3fAnSOOd2_0),.dout(w_dff_B_i9OJ2SyL0_0),.clk(gclk));
	jdff dff_B_eMBNXdNB4_0(.din(w_dff_B_i9OJ2SyL0_0),.dout(w_dff_B_eMBNXdNB4_0),.clk(gclk));
	jdff dff_B_HtrNzdA12_0(.din(w_dff_B_eMBNXdNB4_0),.dout(w_dff_B_HtrNzdA12_0),.clk(gclk));
	jdff dff_B_8k0y6odc7_0(.din(w_dff_B_HtrNzdA12_0),.dout(w_dff_B_8k0y6odc7_0),.clk(gclk));
	jdff dff_B_zzKyXlL40_0(.din(w_dff_B_8k0y6odc7_0),.dout(w_dff_B_zzKyXlL40_0),.clk(gclk));
	jdff dff_B_FqdQTw0W7_0(.din(w_dff_B_zzKyXlL40_0),.dout(w_dff_B_FqdQTw0W7_0),.clk(gclk));
	jdff dff_B_WpwrAOeV6_0(.din(w_dff_B_FqdQTw0W7_0),.dout(w_dff_B_WpwrAOeV6_0),.clk(gclk));
	jdff dff_B_51kRVBih6_0(.din(w_dff_B_WpwrAOeV6_0),.dout(w_dff_B_51kRVBih6_0),.clk(gclk));
	jdff dff_B_cVlwItkV7_0(.din(w_dff_B_51kRVBih6_0),.dout(w_dff_B_cVlwItkV7_0),.clk(gclk));
	jdff dff_B_p7WDw7xv5_0(.din(w_dff_B_cVlwItkV7_0),.dout(w_dff_B_p7WDw7xv5_0),.clk(gclk));
	jdff dff_B_Zjihcsk99_0(.din(w_dff_B_p7WDw7xv5_0),.dout(w_dff_B_Zjihcsk99_0),.clk(gclk));
	jdff dff_B_6C0fUjTS9_0(.din(w_dff_B_Zjihcsk99_0),.dout(w_dff_B_6C0fUjTS9_0),.clk(gclk));
	jdff dff_B_PZt9ZuhX2_0(.din(w_dff_B_6C0fUjTS9_0),.dout(w_dff_B_PZt9ZuhX2_0),.clk(gclk));
	jdff dff_B_l9IeCJRH7_0(.din(w_dff_B_PZt9ZuhX2_0),.dout(w_dff_B_l9IeCJRH7_0),.clk(gclk));
	jdff dff_B_LO9LHHVb9_0(.din(w_dff_B_l9IeCJRH7_0),.dout(w_dff_B_LO9LHHVb9_0),.clk(gclk));
	jdff dff_B_LDV9GZol4_0(.din(w_dff_B_LO9LHHVb9_0),.dout(w_dff_B_LDV9GZol4_0),.clk(gclk));
	jdff dff_B_5NpUfDCB0_0(.din(w_dff_B_LDV9GZol4_0),.dout(w_dff_B_5NpUfDCB0_0),.clk(gclk));
	jdff dff_B_VmNsO4Go8_0(.din(w_dff_B_5NpUfDCB0_0),.dout(w_dff_B_VmNsO4Go8_0),.clk(gclk));
	jdff dff_B_MYjzijZW4_0(.din(w_dff_B_VmNsO4Go8_0),.dout(w_dff_B_MYjzijZW4_0),.clk(gclk));
	jdff dff_B_SMQciwVq1_0(.din(w_dff_B_MYjzijZW4_0),.dout(w_dff_B_SMQciwVq1_0),.clk(gclk));
	jdff dff_B_ix9eixGn3_0(.din(w_dff_B_SMQciwVq1_0),.dout(w_dff_B_ix9eixGn3_0),.clk(gclk));
	jdff dff_B_JY5qLTsg5_0(.din(w_dff_B_ix9eixGn3_0),.dout(w_dff_B_JY5qLTsg5_0),.clk(gclk));
	jdff dff_B_kGbyK0P85_0(.din(w_dff_B_JY5qLTsg5_0),.dout(w_dff_B_kGbyK0P85_0),.clk(gclk));
	jdff dff_B_VSIalSkS8_0(.din(w_dff_B_kGbyK0P85_0),.dout(w_dff_B_VSIalSkS8_0),.clk(gclk));
	jdff dff_B_zzr6kFSZ2_0(.din(w_dff_B_VSIalSkS8_0),.dout(w_dff_B_zzr6kFSZ2_0),.clk(gclk));
	jdff dff_B_iwC1qx737_0(.din(w_dff_B_zzr6kFSZ2_0),.dout(w_dff_B_iwC1qx737_0),.clk(gclk));
	jdff dff_B_LGOGR9YC7_0(.din(w_dff_B_iwC1qx737_0),.dout(w_dff_B_LGOGR9YC7_0),.clk(gclk));
	jdff dff_B_YpLf8Nod4_0(.din(w_dff_B_LGOGR9YC7_0),.dout(w_dff_B_YpLf8Nod4_0),.clk(gclk));
	jdff dff_B_au9UPdnR0_0(.din(w_dff_B_YpLf8Nod4_0),.dout(w_dff_B_au9UPdnR0_0),.clk(gclk));
	jdff dff_B_g94g8swf6_0(.din(w_dff_B_au9UPdnR0_0),.dout(w_dff_B_g94g8swf6_0),.clk(gclk));
	jdff dff_B_D1UWS14P5_0(.din(w_dff_B_g94g8swf6_0),.dout(w_dff_B_D1UWS14P5_0),.clk(gclk));
	jdff dff_B_XmXDk5Sm5_0(.din(w_dff_B_D1UWS14P5_0),.dout(w_dff_B_XmXDk5Sm5_0),.clk(gclk));
	jdff dff_B_oXxfIAPA4_0(.din(w_dff_B_XmXDk5Sm5_0),.dout(w_dff_B_oXxfIAPA4_0),.clk(gclk));
	jdff dff_B_zEaB8Ke58_0(.din(w_dff_B_oXxfIAPA4_0),.dout(w_dff_B_zEaB8Ke58_0),.clk(gclk));
	jdff dff_B_oDifmN1a4_0(.din(w_dff_B_zEaB8Ke58_0),.dout(w_dff_B_oDifmN1a4_0),.clk(gclk));
	jdff dff_B_DvpOnxyT4_0(.din(w_dff_B_oDifmN1a4_0),.dout(w_dff_B_DvpOnxyT4_0),.clk(gclk));
	jdff dff_B_2Q35UFnP7_0(.din(w_dff_B_DvpOnxyT4_0),.dout(w_dff_B_2Q35UFnP7_0),.clk(gclk));
	jdff dff_B_MODqHYDS0_0(.din(w_dff_B_2Q35UFnP7_0),.dout(w_dff_B_MODqHYDS0_0),.clk(gclk));
	jdff dff_B_aGYC2kHH9_0(.din(w_dff_B_MODqHYDS0_0),.dout(w_dff_B_aGYC2kHH9_0),.clk(gclk));
	jdff dff_B_eNX3bVES5_0(.din(w_dff_B_aGYC2kHH9_0),.dout(w_dff_B_eNX3bVES5_0),.clk(gclk));
	jdff dff_B_t3PLhM7D0_0(.din(w_dff_B_eNX3bVES5_0),.dout(w_dff_B_t3PLhM7D0_0),.clk(gclk));
	jdff dff_B_6luBvCat5_0(.din(w_dff_B_t3PLhM7D0_0),.dout(w_dff_B_6luBvCat5_0),.clk(gclk));
	jdff dff_B_iK4jWOFR2_0(.din(w_dff_B_6luBvCat5_0),.dout(w_dff_B_iK4jWOFR2_0),.clk(gclk));
	jdff dff_B_uw84qvIf3_0(.din(w_dff_B_iK4jWOFR2_0),.dout(w_dff_B_uw84qvIf3_0),.clk(gclk));
	jdff dff_B_vOcnNdYY1_0(.din(w_dff_B_uw84qvIf3_0),.dout(w_dff_B_vOcnNdYY1_0),.clk(gclk));
	jdff dff_B_JR5SiCzG0_0(.din(w_dff_B_vOcnNdYY1_0),.dout(w_dff_B_JR5SiCzG0_0),.clk(gclk));
	jdff dff_B_TNJgKzWo1_1(.din(n1044),.dout(w_dff_B_TNJgKzWo1_1),.clk(gclk));
	jdff dff_B_lBCSnp2r7_1(.din(w_dff_B_TNJgKzWo1_1),.dout(w_dff_B_lBCSnp2r7_1),.clk(gclk));
	jdff dff_B_AVtLB6jr6_1(.din(w_dff_B_lBCSnp2r7_1),.dout(w_dff_B_AVtLB6jr6_1),.clk(gclk));
	jdff dff_B_24zzqBRI7_1(.din(w_dff_B_AVtLB6jr6_1),.dout(w_dff_B_24zzqBRI7_1),.clk(gclk));
	jdff dff_B_x00mff6S6_1(.din(w_dff_B_24zzqBRI7_1),.dout(w_dff_B_x00mff6S6_1),.clk(gclk));
	jdff dff_B_CDoGWpv02_1(.din(w_dff_B_x00mff6S6_1),.dout(w_dff_B_CDoGWpv02_1),.clk(gclk));
	jdff dff_B_VGwfrrk02_1(.din(w_dff_B_CDoGWpv02_1),.dout(w_dff_B_VGwfrrk02_1),.clk(gclk));
	jdff dff_B_R7azb7Nd0_1(.din(w_dff_B_VGwfrrk02_1),.dout(w_dff_B_R7azb7Nd0_1),.clk(gclk));
	jdff dff_B_v3RRxXsr0_1(.din(w_dff_B_R7azb7Nd0_1),.dout(w_dff_B_v3RRxXsr0_1),.clk(gclk));
	jdff dff_B_sFTrb7JH8_1(.din(w_dff_B_v3RRxXsr0_1),.dout(w_dff_B_sFTrb7JH8_1),.clk(gclk));
	jdff dff_B_JXW2zXQv5_1(.din(w_dff_B_sFTrb7JH8_1),.dout(w_dff_B_JXW2zXQv5_1),.clk(gclk));
	jdff dff_B_qLZvhUXn6_1(.din(w_dff_B_JXW2zXQv5_1),.dout(w_dff_B_qLZvhUXn6_1),.clk(gclk));
	jdff dff_B_Zs7x17fS0_1(.din(w_dff_B_qLZvhUXn6_1),.dout(w_dff_B_Zs7x17fS0_1),.clk(gclk));
	jdff dff_B_htye1RPi7_1(.din(w_dff_B_Zs7x17fS0_1),.dout(w_dff_B_htye1RPi7_1),.clk(gclk));
	jdff dff_B_uveo5U1G9_1(.din(w_dff_B_htye1RPi7_1),.dout(w_dff_B_uveo5U1G9_1),.clk(gclk));
	jdff dff_B_FC3OSfkT6_1(.din(w_dff_B_uveo5U1G9_1),.dout(w_dff_B_FC3OSfkT6_1),.clk(gclk));
	jdff dff_B_URjIChGw1_1(.din(w_dff_B_FC3OSfkT6_1),.dout(w_dff_B_URjIChGw1_1),.clk(gclk));
	jdff dff_B_cilZ3TtY0_1(.din(w_dff_B_URjIChGw1_1),.dout(w_dff_B_cilZ3TtY0_1),.clk(gclk));
	jdff dff_B_P8JUk6yn2_1(.din(w_dff_B_cilZ3TtY0_1),.dout(w_dff_B_P8JUk6yn2_1),.clk(gclk));
	jdff dff_B_sY810B3m1_1(.din(w_dff_B_P8JUk6yn2_1),.dout(w_dff_B_sY810B3m1_1),.clk(gclk));
	jdff dff_B_yfXeADdj6_1(.din(w_dff_B_sY810B3m1_1),.dout(w_dff_B_yfXeADdj6_1),.clk(gclk));
	jdff dff_B_AUyAgJEw7_1(.din(w_dff_B_yfXeADdj6_1),.dout(w_dff_B_AUyAgJEw7_1),.clk(gclk));
	jdff dff_B_oYwKGmbN0_1(.din(w_dff_B_AUyAgJEw7_1),.dout(w_dff_B_oYwKGmbN0_1),.clk(gclk));
	jdff dff_B_WNN78y1p2_1(.din(w_dff_B_oYwKGmbN0_1),.dout(w_dff_B_WNN78y1p2_1),.clk(gclk));
	jdff dff_B_BmZiL57t3_1(.din(w_dff_B_WNN78y1p2_1),.dout(w_dff_B_BmZiL57t3_1),.clk(gclk));
	jdff dff_B_l01DRcmO0_1(.din(w_dff_B_BmZiL57t3_1),.dout(w_dff_B_l01DRcmO0_1),.clk(gclk));
	jdff dff_B_IIxIsKNe0_1(.din(w_dff_B_l01DRcmO0_1),.dout(w_dff_B_IIxIsKNe0_1),.clk(gclk));
	jdff dff_B_0EvjvlxC6_1(.din(w_dff_B_IIxIsKNe0_1),.dout(w_dff_B_0EvjvlxC6_1),.clk(gclk));
	jdff dff_B_d0vS4m3V9_1(.din(w_dff_B_0EvjvlxC6_1),.dout(w_dff_B_d0vS4m3V9_1),.clk(gclk));
	jdff dff_B_ZUldIZr71_1(.din(w_dff_B_d0vS4m3V9_1),.dout(w_dff_B_ZUldIZr71_1),.clk(gclk));
	jdff dff_B_cV71bmen7_1(.din(w_dff_B_ZUldIZr71_1),.dout(w_dff_B_cV71bmen7_1),.clk(gclk));
	jdff dff_B_zWCE6COk1_1(.din(w_dff_B_cV71bmen7_1),.dout(w_dff_B_zWCE6COk1_1),.clk(gclk));
	jdff dff_B_YgtXdsHb7_1(.din(w_dff_B_zWCE6COk1_1),.dout(w_dff_B_YgtXdsHb7_1),.clk(gclk));
	jdff dff_B_iRSEWnqw4_1(.din(w_dff_B_YgtXdsHb7_1),.dout(w_dff_B_iRSEWnqw4_1),.clk(gclk));
	jdff dff_B_e1hi6Rn85_1(.din(w_dff_B_iRSEWnqw4_1),.dout(w_dff_B_e1hi6Rn85_1),.clk(gclk));
	jdff dff_B_3NjjINVj8_1(.din(w_dff_B_e1hi6Rn85_1),.dout(w_dff_B_3NjjINVj8_1),.clk(gclk));
	jdff dff_B_RAtNW0Gg1_1(.din(w_dff_B_3NjjINVj8_1),.dout(w_dff_B_RAtNW0Gg1_1),.clk(gclk));
	jdff dff_B_AqJAn9bb1_1(.din(w_dff_B_RAtNW0Gg1_1),.dout(w_dff_B_AqJAn9bb1_1),.clk(gclk));
	jdff dff_B_gZsuQJOZ9_1(.din(w_dff_B_AqJAn9bb1_1),.dout(w_dff_B_gZsuQJOZ9_1),.clk(gclk));
	jdff dff_B_7qyUS5Wd2_1(.din(w_dff_B_gZsuQJOZ9_1),.dout(w_dff_B_7qyUS5Wd2_1),.clk(gclk));
	jdff dff_B_ACuUdNia4_1(.din(w_dff_B_7qyUS5Wd2_1),.dout(w_dff_B_ACuUdNia4_1),.clk(gclk));
	jdff dff_B_X5gl6zrp8_1(.din(w_dff_B_ACuUdNia4_1),.dout(w_dff_B_X5gl6zrp8_1),.clk(gclk));
	jdff dff_B_9o42I44L6_1(.din(w_dff_B_X5gl6zrp8_1),.dout(w_dff_B_9o42I44L6_1),.clk(gclk));
	jdff dff_B_5mx11BE19_1(.din(w_dff_B_9o42I44L6_1),.dout(w_dff_B_5mx11BE19_1),.clk(gclk));
	jdff dff_B_iMrH0NZ31_1(.din(w_dff_B_5mx11BE19_1),.dout(w_dff_B_iMrH0NZ31_1),.clk(gclk));
	jdff dff_B_78QfnOWx4_1(.din(w_dff_B_iMrH0NZ31_1),.dout(w_dff_B_78QfnOWx4_1),.clk(gclk));
	jdff dff_B_iJowQtKq0_1(.din(w_dff_B_78QfnOWx4_1),.dout(w_dff_B_iJowQtKq0_1),.clk(gclk));
	jdff dff_B_cf3m5jsR2_1(.din(w_dff_B_iJowQtKq0_1),.dout(w_dff_B_cf3m5jsR2_1),.clk(gclk));
	jdff dff_B_uSgMIlFd1_1(.din(w_dff_B_cf3m5jsR2_1),.dout(w_dff_B_uSgMIlFd1_1),.clk(gclk));
	jdff dff_B_czIanC4b1_1(.din(w_dff_B_uSgMIlFd1_1),.dout(w_dff_B_czIanC4b1_1),.clk(gclk));
	jdff dff_B_0SsKP0wG1_1(.din(w_dff_B_czIanC4b1_1),.dout(w_dff_B_0SsKP0wG1_1),.clk(gclk));
	jdff dff_B_kMOcvVJd2_1(.din(w_dff_B_0SsKP0wG1_1),.dout(w_dff_B_kMOcvVJd2_1),.clk(gclk));
	jdff dff_B_AryzQLz15_1(.din(w_dff_B_kMOcvVJd2_1),.dout(w_dff_B_AryzQLz15_1),.clk(gclk));
	jdff dff_B_DQxIC9Z15_1(.din(w_dff_B_AryzQLz15_1),.dout(w_dff_B_DQxIC9Z15_1),.clk(gclk));
	jdff dff_B_bOKXOzTI4_1(.din(w_dff_B_DQxIC9Z15_1),.dout(w_dff_B_bOKXOzTI4_1),.clk(gclk));
	jdff dff_B_PJynUqyP3_1(.din(w_dff_B_bOKXOzTI4_1),.dout(w_dff_B_PJynUqyP3_1),.clk(gclk));
	jdff dff_B_BXe3PbWw8_1(.din(w_dff_B_PJynUqyP3_1),.dout(w_dff_B_BXe3PbWw8_1),.clk(gclk));
	jdff dff_B_gIFHpA6r4_1(.din(w_dff_B_BXe3PbWw8_1),.dout(w_dff_B_gIFHpA6r4_1),.clk(gclk));
	jdff dff_B_l9MmpgVJ6_1(.din(w_dff_B_gIFHpA6r4_1),.dout(w_dff_B_l9MmpgVJ6_1),.clk(gclk));
	jdff dff_B_BSPTMW9T6_1(.din(w_dff_B_l9MmpgVJ6_1),.dout(w_dff_B_BSPTMW9T6_1),.clk(gclk));
	jdff dff_B_z6XbKa2O2_1(.din(w_dff_B_BSPTMW9T6_1),.dout(w_dff_B_z6XbKa2O2_1),.clk(gclk));
	jdff dff_B_zMf20qIv4_1(.din(w_dff_B_z6XbKa2O2_1),.dout(w_dff_B_zMf20qIv4_1),.clk(gclk));
	jdff dff_B_lESTFKZ39_1(.din(w_dff_B_zMf20qIv4_1),.dout(w_dff_B_lESTFKZ39_1),.clk(gclk));
	jdff dff_B_a72zZHwv7_1(.din(w_dff_B_lESTFKZ39_1),.dout(w_dff_B_a72zZHwv7_1),.clk(gclk));
	jdff dff_B_fvfuyOux9_1(.din(w_dff_B_a72zZHwv7_1),.dout(w_dff_B_fvfuyOux9_1),.clk(gclk));
	jdff dff_B_laBtyieW9_1(.din(w_dff_B_fvfuyOux9_1),.dout(w_dff_B_laBtyieW9_1),.clk(gclk));
	jdff dff_B_tfNxG1O59_1(.din(w_dff_B_laBtyieW9_1),.dout(w_dff_B_tfNxG1O59_1),.clk(gclk));
	jdff dff_B_xSu9ZqGL9_1(.din(w_dff_B_tfNxG1O59_1),.dout(w_dff_B_xSu9ZqGL9_1),.clk(gclk));
	jdff dff_B_byiIojBQ1_1(.din(w_dff_B_xSu9ZqGL9_1),.dout(w_dff_B_byiIojBQ1_1),.clk(gclk));
	jdff dff_B_TcMM18NK4_1(.din(w_dff_B_byiIojBQ1_1),.dout(w_dff_B_TcMM18NK4_1),.clk(gclk));
	jdff dff_B_iYUPolPE7_1(.din(w_dff_B_TcMM18NK4_1),.dout(w_dff_B_iYUPolPE7_1),.clk(gclk));
	jdff dff_B_gYVM8Glb9_1(.din(w_dff_B_iYUPolPE7_1),.dout(w_dff_B_gYVM8Glb9_1),.clk(gclk));
	jdff dff_B_Sfr4aSJK3_1(.din(w_dff_B_gYVM8Glb9_1),.dout(w_dff_B_Sfr4aSJK3_1),.clk(gclk));
	jdff dff_B_VCcD85Xm0_1(.din(w_dff_B_Sfr4aSJK3_1),.dout(w_dff_B_VCcD85Xm0_1),.clk(gclk));
	jdff dff_B_dsvKWkqG3_1(.din(w_dff_B_VCcD85Xm0_1),.dout(w_dff_B_dsvKWkqG3_1),.clk(gclk));
	jdff dff_B_LKHs9SzN2_1(.din(w_dff_B_dsvKWkqG3_1),.dout(w_dff_B_LKHs9SzN2_1),.clk(gclk));
	jdff dff_B_EHMgFfpX0_1(.din(w_dff_B_LKHs9SzN2_1),.dout(w_dff_B_EHMgFfpX0_1),.clk(gclk));
	jdff dff_B_NN6hkRKp7_1(.din(w_dff_B_EHMgFfpX0_1),.dout(w_dff_B_NN6hkRKp7_1),.clk(gclk));
	jdff dff_B_8Z3PMryr0_1(.din(w_dff_B_NN6hkRKp7_1),.dout(w_dff_B_8Z3PMryr0_1),.clk(gclk));
	jdff dff_B_MWsgv9wk2_1(.din(w_dff_B_8Z3PMryr0_1),.dout(w_dff_B_MWsgv9wk2_1),.clk(gclk));
	jdff dff_B_6XyXBagH2_1(.din(w_dff_B_MWsgv9wk2_1),.dout(w_dff_B_6XyXBagH2_1),.clk(gclk));
	jdff dff_B_9IMyFUuV7_1(.din(w_dff_B_6XyXBagH2_1),.dout(w_dff_B_9IMyFUuV7_1),.clk(gclk));
	jdff dff_B_Ybge9p9p6_1(.din(w_dff_B_9IMyFUuV7_1),.dout(w_dff_B_Ybge9p9p6_1),.clk(gclk));
	jdff dff_B_BZ0kkJPv2_1(.din(w_dff_B_Ybge9p9p6_1),.dout(w_dff_B_BZ0kkJPv2_1),.clk(gclk));
	jdff dff_B_3aSt7qKB5_1(.din(w_dff_B_BZ0kkJPv2_1),.dout(w_dff_B_3aSt7qKB5_1),.clk(gclk));
	jdff dff_B_8D7NpUrs5_1(.din(w_dff_B_3aSt7qKB5_1),.dout(w_dff_B_8D7NpUrs5_1),.clk(gclk));
	jdff dff_B_1U6ocUSr9_1(.din(w_dff_B_8D7NpUrs5_1),.dout(w_dff_B_1U6ocUSr9_1),.clk(gclk));
	jdff dff_B_MZcbJ2FL9_1(.din(w_dff_B_1U6ocUSr9_1),.dout(w_dff_B_MZcbJ2FL9_1),.clk(gclk));
	jdff dff_B_ZbzCUrij7_1(.din(w_dff_B_MZcbJ2FL9_1),.dout(w_dff_B_ZbzCUrij7_1),.clk(gclk));
	jdff dff_B_Iy6YBLzm9_1(.din(w_dff_B_ZbzCUrij7_1),.dout(w_dff_B_Iy6YBLzm9_1),.clk(gclk));
	jdff dff_B_zo0eN7VF1_1(.din(w_dff_B_Iy6YBLzm9_1),.dout(w_dff_B_zo0eN7VF1_1),.clk(gclk));
	jdff dff_B_LetsnoQ83_1(.din(w_dff_B_zo0eN7VF1_1),.dout(w_dff_B_LetsnoQ83_1),.clk(gclk));
	jdff dff_B_QMtwEum80_1(.din(w_dff_B_LetsnoQ83_1),.dout(w_dff_B_QMtwEum80_1),.clk(gclk));
	jdff dff_B_XOHB2wXJ3_1(.din(w_dff_B_QMtwEum80_1),.dout(w_dff_B_XOHB2wXJ3_1),.clk(gclk));
	jdff dff_B_M33UaZg95_1(.din(w_dff_B_XOHB2wXJ3_1),.dout(w_dff_B_M33UaZg95_1),.clk(gclk));
	jdff dff_B_8nKa2SG72_1(.din(w_dff_B_M33UaZg95_1),.dout(w_dff_B_8nKa2SG72_1),.clk(gclk));
	jdff dff_B_6ys3D0sJ8_1(.din(w_dff_B_8nKa2SG72_1),.dout(w_dff_B_6ys3D0sJ8_1),.clk(gclk));
	jdff dff_B_o0TBXR9R3_1(.din(w_dff_B_6ys3D0sJ8_1),.dout(w_dff_B_o0TBXR9R3_1),.clk(gclk));
	jdff dff_B_p2oBQjh34_1(.din(w_dff_B_o0TBXR9R3_1),.dout(w_dff_B_p2oBQjh34_1),.clk(gclk));
	jdff dff_B_9abC3eYk2_1(.din(w_dff_B_p2oBQjh34_1),.dout(w_dff_B_9abC3eYk2_1),.clk(gclk));
	jdff dff_B_DV8yiukN4_1(.din(w_dff_B_9abC3eYk2_1),.dout(w_dff_B_DV8yiukN4_1),.clk(gclk));
	jdff dff_B_vUmolh8w9_1(.din(w_dff_B_DV8yiukN4_1),.dout(w_dff_B_vUmolh8w9_1),.clk(gclk));
	jdff dff_B_7DHWEMMT2_1(.din(w_dff_B_vUmolh8w9_1),.dout(w_dff_B_7DHWEMMT2_1),.clk(gclk));
	jdff dff_B_FMeYhrLy9_1(.din(w_dff_B_7DHWEMMT2_1),.dout(w_dff_B_FMeYhrLy9_1),.clk(gclk));
	jdff dff_B_V0ivtjd62_1(.din(w_dff_B_FMeYhrLy9_1),.dout(w_dff_B_V0ivtjd62_1),.clk(gclk));
	jdff dff_B_H8tSLsLj6_1(.din(w_dff_B_V0ivtjd62_1),.dout(w_dff_B_H8tSLsLj6_1),.clk(gclk));
	jdff dff_B_Vf5hwBZA4_1(.din(w_dff_B_H8tSLsLj6_1),.dout(w_dff_B_Vf5hwBZA4_1),.clk(gclk));
	jdff dff_B_ZTG1a3co6_1(.din(w_dff_B_Vf5hwBZA4_1),.dout(w_dff_B_ZTG1a3co6_1),.clk(gclk));
	jdff dff_B_3DnFUkNN0_1(.din(w_dff_B_ZTG1a3co6_1),.dout(w_dff_B_3DnFUkNN0_1),.clk(gclk));
	jdff dff_B_sX8cRBX78_1(.din(w_dff_B_3DnFUkNN0_1),.dout(w_dff_B_sX8cRBX78_1),.clk(gclk));
	jdff dff_B_eijfc5pg6_0(.din(n1045),.dout(w_dff_B_eijfc5pg6_0),.clk(gclk));
	jdff dff_B_Kki71dkq6_0(.din(w_dff_B_eijfc5pg6_0),.dout(w_dff_B_Kki71dkq6_0),.clk(gclk));
	jdff dff_B_8tQuyefM2_0(.din(w_dff_B_Kki71dkq6_0),.dout(w_dff_B_8tQuyefM2_0),.clk(gclk));
	jdff dff_B_FaedtkvH6_0(.din(w_dff_B_8tQuyefM2_0),.dout(w_dff_B_FaedtkvH6_0),.clk(gclk));
	jdff dff_B_kpbLbBbY0_0(.din(w_dff_B_FaedtkvH6_0),.dout(w_dff_B_kpbLbBbY0_0),.clk(gclk));
	jdff dff_B_wPp5KZpI7_0(.din(w_dff_B_kpbLbBbY0_0),.dout(w_dff_B_wPp5KZpI7_0),.clk(gclk));
	jdff dff_B_1bxbF8on2_0(.din(w_dff_B_wPp5KZpI7_0),.dout(w_dff_B_1bxbF8on2_0),.clk(gclk));
	jdff dff_B_vSXwfNEF7_0(.din(w_dff_B_1bxbF8on2_0),.dout(w_dff_B_vSXwfNEF7_0),.clk(gclk));
	jdff dff_B_eijOniyI3_0(.din(w_dff_B_vSXwfNEF7_0),.dout(w_dff_B_eijOniyI3_0),.clk(gclk));
	jdff dff_B_nV3SEymu4_0(.din(w_dff_B_eijOniyI3_0),.dout(w_dff_B_nV3SEymu4_0),.clk(gclk));
	jdff dff_B_8kv3raGy9_0(.din(w_dff_B_nV3SEymu4_0),.dout(w_dff_B_8kv3raGy9_0),.clk(gclk));
	jdff dff_B_eV68pfbm2_0(.din(w_dff_B_8kv3raGy9_0),.dout(w_dff_B_eV68pfbm2_0),.clk(gclk));
	jdff dff_B_100189Eh1_0(.din(w_dff_B_eV68pfbm2_0),.dout(w_dff_B_100189Eh1_0),.clk(gclk));
	jdff dff_B_OX60F6sO5_0(.din(w_dff_B_100189Eh1_0),.dout(w_dff_B_OX60F6sO5_0),.clk(gclk));
	jdff dff_B_2ZhW6l159_0(.din(w_dff_B_OX60F6sO5_0),.dout(w_dff_B_2ZhW6l159_0),.clk(gclk));
	jdff dff_B_ZxPYZXRq7_0(.din(w_dff_B_2ZhW6l159_0),.dout(w_dff_B_ZxPYZXRq7_0),.clk(gclk));
	jdff dff_B_2hpBib9f8_0(.din(w_dff_B_ZxPYZXRq7_0),.dout(w_dff_B_2hpBib9f8_0),.clk(gclk));
	jdff dff_B_wh6eX9fk6_0(.din(w_dff_B_2hpBib9f8_0),.dout(w_dff_B_wh6eX9fk6_0),.clk(gclk));
	jdff dff_B_rKbtq0A12_0(.din(w_dff_B_wh6eX9fk6_0),.dout(w_dff_B_rKbtq0A12_0),.clk(gclk));
	jdff dff_B_uYH3qtOg1_0(.din(w_dff_B_rKbtq0A12_0),.dout(w_dff_B_uYH3qtOg1_0),.clk(gclk));
	jdff dff_B_2yYLkmNq7_0(.din(w_dff_B_uYH3qtOg1_0),.dout(w_dff_B_2yYLkmNq7_0),.clk(gclk));
	jdff dff_B_31P7kpkf3_0(.din(w_dff_B_2yYLkmNq7_0),.dout(w_dff_B_31P7kpkf3_0),.clk(gclk));
	jdff dff_B_KnAeTAsA9_0(.din(w_dff_B_31P7kpkf3_0),.dout(w_dff_B_KnAeTAsA9_0),.clk(gclk));
	jdff dff_B_rrOkmwmw6_0(.din(w_dff_B_KnAeTAsA9_0),.dout(w_dff_B_rrOkmwmw6_0),.clk(gclk));
	jdff dff_B_1mOsWA3e8_0(.din(w_dff_B_rrOkmwmw6_0),.dout(w_dff_B_1mOsWA3e8_0),.clk(gclk));
	jdff dff_B_vNc2k22x5_0(.din(w_dff_B_1mOsWA3e8_0),.dout(w_dff_B_vNc2k22x5_0),.clk(gclk));
	jdff dff_B_H9jodjJU9_0(.din(w_dff_B_vNc2k22x5_0),.dout(w_dff_B_H9jodjJU9_0),.clk(gclk));
	jdff dff_B_MuNVOHU85_0(.din(w_dff_B_H9jodjJU9_0),.dout(w_dff_B_MuNVOHU85_0),.clk(gclk));
	jdff dff_B_bS1gtJIQ2_0(.din(w_dff_B_MuNVOHU85_0),.dout(w_dff_B_bS1gtJIQ2_0),.clk(gclk));
	jdff dff_B_Fy5hxjQG2_0(.din(w_dff_B_bS1gtJIQ2_0),.dout(w_dff_B_Fy5hxjQG2_0),.clk(gclk));
	jdff dff_B_ESI79r7D6_0(.din(w_dff_B_Fy5hxjQG2_0),.dout(w_dff_B_ESI79r7D6_0),.clk(gclk));
	jdff dff_B_pN7FLYz65_0(.din(w_dff_B_ESI79r7D6_0),.dout(w_dff_B_pN7FLYz65_0),.clk(gclk));
	jdff dff_B_aRPsBVvL0_0(.din(w_dff_B_pN7FLYz65_0),.dout(w_dff_B_aRPsBVvL0_0),.clk(gclk));
	jdff dff_B_x117IfYm2_0(.din(w_dff_B_aRPsBVvL0_0),.dout(w_dff_B_x117IfYm2_0),.clk(gclk));
	jdff dff_B_ayDpPYeB9_0(.din(w_dff_B_x117IfYm2_0),.dout(w_dff_B_ayDpPYeB9_0),.clk(gclk));
	jdff dff_B_8c211PYI1_0(.din(w_dff_B_ayDpPYeB9_0),.dout(w_dff_B_8c211PYI1_0),.clk(gclk));
	jdff dff_B_JurUsh7g3_0(.din(w_dff_B_8c211PYI1_0),.dout(w_dff_B_JurUsh7g3_0),.clk(gclk));
	jdff dff_B_Ny1UPnCN7_0(.din(w_dff_B_JurUsh7g3_0),.dout(w_dff_B_Ny1UPnCN7_0),.clk(gclk));
	jdff dff_B_jb4Whx431_0(.din(w_dff_B_Ny1UPnCN7_0),.dout(w_dff_B_jb4Whx431_0),.clk(gclk));
	jdff dff_B_JdekCFq97_0(.din(w_dff_B_jb4Whx431_0),.dout(w_dff_B_JdekCFq97_0),.clk(gclk));
	jdff dff_B_bCh4qLeT5_0(.din(w_dff_B_JdekCFq97_0),.dout(w_dff_B_bCh4qLeT5_0),.clk(gclk));
	jdff dff_B_larob4IN7_0(.din(w_dff_B_bCh4qLeT5_0),.dout(w_dff_B_larob4IN7_0),.clk(gclk));
	jdff dff_B_59UCg4tp4_0(.din(w_dff_B_larob4IN7_0),.dout(w_dff_B_59UCg4tp4_0),.clk(gclk));
	jdff dff_B_zWSRUSon2_0(.din(w_dff_B_59UCg4tp4_0),.dout(w_dff_B_zWSRUSon2_0),.clk(gclk));
	jdff dff_B_VmeH1jGz6_0(.din(w_dff_B_zWSRUSon2_0),.dout(w_dff_B_VmeH1jGz6_0),.clk(gclk));
	jdff dff_B_0U550N7F1_0(.din(w_dff_B_VmeH1jGz6_0),.dout(w_dff_B_0U550N7F1_0),.clk(gclk));
	jdff dff_B_ukIxxz0y6_0(.din(w_dff_B_0U550N7F1_0),.dout(w_dff_B_ukIxxz0y6_0),.clk(gclk));
	jdff dff_B_0t9lsczO6_0(.din(w_dff_B_ukIxxz0y6_0),.dout(w_dff_B_0t9lsczO6_0),.clk(gclk));
	jdff dff_B_hrQNrluM5_0(.din(w_dff_B_0t9lsczO6_0),.dout(w_dff_B_hrQNrluM5_0),.clk(gclk));
	jdff dff_B_Uai1f90i2_0(.din(w_dff_B_hrQNrluM5_0),.dout(w_dff_B_Uai1f90i2_0),.clk(gclk));
	jdff dff_B_STa2ezN83_0(.din(w_dff_B_Uai1f90i2_0),.dout(w_dff_B_STa2ezN83_0),.clk(gclk));
	jdff dff_B_Ldlh7Pm86_0(.din(w_dff_B_STa2ezN83_0),.dout(w_dff_B_Ldlh7Pm86_0),.clk(gclk));
	jdff dff_B_ERu4tLOb4_0(.din(w_dff_B_Ldlh7Pm86_0),.dout(w_dff_B_ERu4tLOb4_0),.clk(gclk));
	jdff dff_B_RiBaRBtP4_0(.din(w_dff_B_ERu4tLOb4_0),.dout(w_dff_B_RiBaRBtP4_0),.clk(gclk));
	jdff dff_B_GW4R7AIJ5_0(.din(w_dff_B_RiBaRBtP4_0),.dout(w_dff_B_GW4R7AIJ5_0),.clk(gclk));
	jdff dff_B_uPnO5vJ01_0(.din(w_dff_B_GW4R7AIJ5_0),.dout(w_dff_B_uPnO5vJ01_0),.clk(gclk));
	jdff dff_B_TzLWDAsc6_0(.din(w_dff_B_uPnO5vJ01_0),.dout(w_dff_B_TzLWDAsc6_0),.clk(gclk));
	jdff dff_B_3H9T2crH9_0(.din(w_dff_B_TzLWDAsc6_0),.dout(w_dff_B_3H9T2crH9_0),.clk(gclk));
	jdff dff_B_IBPXt5Ow0_0(.din(w_dff_B_3H9T2crH9_0),.dout(w_dff_B_IBPXt5Ow0_0),.clk(gclk));
	jdff dff_B_4hqYCYAG7_0(.din(w_dff_B_IBPXt5Ow0_0),.dout(w_dff_B_4hqYCYAG7_0),.clk(gclk));
	jdff dff_B_BH0Ge5NT6_0(.din(w_dff_B_4hqYCYAG7_0),.dout(w_dff_B_BH0Ge5NT6_0),.clk(gclk));
	jdff dff_B_2daF8TP68_0(.din(w_dff_B_BH0Ge5NT6_0),.dout(w_dff_B_2daF8TP68_0),.clk(gclk));
	jdff dff_B_o39NmiNr7_0(.din(w_dff_B_2daF8TP68_0),.dout(w_dff_B_o39NmiNr7_0),.clk(gclk));
	jdff dff_B_sF22bwQT7_0(.din(w_dff_B_o39NmiNr7_0),.dout(w_dff_B_sF22bwQT7_0),.clk(gclk));
	jdff dff_B_Ph1O0jJO8_0(.din(w_dff_B_sF22bwQT7_0),.dout(w_dff_B_Ph1O0jJO8_0),.clk(gclk));
	jdff dff_B_mis7YoWy3_0(.din(w_dff_B_Ph1O0jJO8_0),.dout(w_dff_B_mis7YoWy3_0),.clk(gclk));
	jdff dff_B_SMG1l1Rg5_0(.din(w_dff_B_mis7YoWy3_0),.dout(w_dff_B_SMG1l1Rg5_0),.clk(gclk));
	jdff dff_B_BFBtnrUY2_0(.din(w_dff_B_SMG1l1Rg5_0),.dout(w_dff_B_BFBtnrUY2_0),.clk(gclk));
	jdff dff_B_T2qhl3b43_0(.din(w_dff_B_BFBtnrUY2_0),.dout(w_dff_B_T2qhl3b43_0),.clk(gclk));
	jdff dff_B_819bPhog1_0(.din(w_dff_B_T2qhl3b43_0),.dout(w_dff_B_819bPhog1_0),.clk(gclk));
	jdff dff_B_CyGo6Nfs8_0(.din(w_dff_B_819bPhog1_0),.dout(w_dff_B_CyGo6Nfs8_0),.clk(gclk));
	jdff dff_B_JIafjria0_0(.din(w_dff_B_CyGo6Nfs8_0),.dout(w_dff_B_JIafjria0_0),.clk(gclk));
	jdff dff_B_YHutGRmb3_0(.din(w_dff_B_JIafjria0_0),.dout(w_dff_B_YHutGRmb3_0),.clk(gclk));
	jdff dff_B_OInsV6VW0_0(.din(w_dff_B_YHutGRmb3_0),.dout(w_dff_B_OInsV6VW0_0),.clk(gclk));
	jdff dff_B_WjXlSdFp5_0(.din(w_dff_B_OInsV6VW0_0),.dout(w_dff_B_WjXlSdFp5_0),.clk(gclk));
	jdff dff_B_hCeTkbMk3_0(.din(w_dff_B_WjXlSdFp5_0),.dout(w_dff_B_hCeTkbMk3_0),.clk(gclk));
	jdff dff_B_WNUB00xy9_0(.din(w_dff_B_hCeTkbMk3_0),.dout(w_dff_B_WNUB00xy9_0),.clk(gclk));
	jdff dff_B_SZ4VXvos9_0(.din(w_dff_B_WNUB00xy9_0),.dout(w_dff_B_SZ4VXvos9_0),.clk(gclk));
	jdff dff_B_yzzc5q2Q3_0(.din(w_dff_B_SZ4VXvos9_0),.dout(w_dff_B_yzzc5q2Q3_0),.clk(gclk));
	jdff dff_B_pkRr9Hfb7_0(.din(w_dff_B_yzzc5q2Q3_0),.dout(w_dff_B_pkRr9Hfb7_0),.clk(gclk));
	jdff dff_B_O7jpM7Rg7_0(.din(w_dff_B_pkRr9Hfb7_0),.dout(w_dff_B_O7jpM7Rg7_0),.clk(gclk));
	jdff dff_B_vL7lzYGD0_0(.din(w_dff_B_O7jpM7Rg7_0),.dout(w_dff_B_vL7lzYGD0_0),.clk(gclk));
	jdff dff_B_YkZUb3pQ5_0(.din(w_dff_B_vL7lzYGD0_0),.dout(w_dff_B_YkZUb3pQ5_0),.clk(gclk));
	jdff dff_B_2qwDEWHw7_0(.din(w_dff_B_YkZUb3pQ5_0),.dout(w_dff_B_2qwDEWHw7_0),.clk(gclk));
	jdff dff_B_7WIssvmJ4_0(.din(w_dff_B_2qwDEWHw7_0),.dout(w_dff_B_7WIssvmJ4_0),.clk(gclk));
	jdff dff_B_Mal5DAro1_0(.din(w_dff_B_7WIssvmJ4_0),.dout(w_dff_B_Mal5DAro1_0),.clk(gclk));
	jdff dff_B_qycH0BtL6_0(.din(w_dff_B_Mal5DAro1_0),.dout(w_dff_B_qycH0BtL6_0),.clk(gclk));
	jdff dff_B_RKNvS5rk7_0(.din(w_dff_B_qycH0BtL6_0),.dout(w_dff_B_RKNvS5rk7_0),.clk(gclk));
	jdff dff_B_dtoruauM9_0(.din(w_dff_B_RKNvS5rk7_0),.dout(w_dff_B_dtoruauM9_0),.clk(gclk));
	jdff dff_B_UqsaClGw3_0(.din(w_dff_B_dtoruauM9_0),.dout(w_dff_B_UqsaClGw3_0),.clk(gclk));
	jdff dff_B_j79nUqGF6_0(.din(w_dff_B_UqsaClGw3_0),.dout(w_dff_B_j79nUqGF6_0),.clk(gclk));
	jdff dff_B_RMfEebmb3_0(.din(w_dff_B_j79nUqGF6_0),.dout(w_dff_B_RMfEebmb3_0),.clk(gclk));
	jdff dff_B_y1FZ4rqb3_0(.din(w_dff_B_RMfEebmb3_0),.dout(w_dff_B_y1FZ4rqb3_0),.clk(gclk));
	jdff dff_B_CVQQtmVk9_0(.din(w_dff_B_y1FZ4rqb3_0),.dout(w_dff_B_CVQQtmVk9_0),.clk(gclk));
	jdff dff_B_l6CIO8uO6_0(.din(w_dff_B_CVQQtmVk9_0),.dout(w_dff_B_l6CIO8uO6_0),.clk(gclk));
	jdff dff_B_a8iR5bg72_0(.din(w_dff_B_l6CIO8uO6_0),.dout(w_dff_B_a8iR5bg72_0),.clk(gclk));
	jdff dff_B_smNCzs7c0_0(.din(w_dff_B_a8iR5bg72_0),.dout(w_dff_B_smNCzs7c0_0),.clk(gclk));
	jdff dff_B_IBJgy6V73_0(.din(w_dff_B_smNCzs7c0_0),.dout(w_dff_B_IBJgy6V73_0),.clk(gclk));
	jdff dff_B_N68b2DFq4_0(.din(w_dff_B_IBJgy6V73_0),.dout(w_dff_B_N68b2DFq4_0),.clk(gclk));
	jdff dff_B_euMyhzMj6_0(.din(w_dff_B_N68b2DFq4_0),.dout(w_dff_B_euMyhzMj6_0),.clk(gclk));
	jdff dff_B_0jmMO6n58_0(.din(w_dff_B_euMyhzMj6_0),.dout(w_dff_B_0jmMO6n58_0),.clk(gclk));
	jdff dff_B_WF6q6UMt6_0(.din(w_dff_B_0jmMO6n58_0),.dout(w_dff_B_WF6q6UMt6_0),.clk(gclk));
	jdff dff_B_L9nTN4eZ4_0(.din(w_dff_B_WF6q6UMt6_0),.dout(w_dff_B_L9nTN4eZ4_0),.clk(gclk));
	jdff dff_B_IrRSRxVR0_0(.din(w_dff_B_L9nTN4eZ4_0),.dout(w_dff_B_IrRSRxVR0_0),.clk(gclk));
	jdff dff_B_GpeT42fu3_0(.din(w_dff_B_IrRSRxVR0_0),.dout(w_dff_B_GpeT42fu3_0),.clk(gclk));
	jdff dff_B_wmA091ne9_0(.din(w_dff_B_GpeT42fu3_0),.dout(w_dff_B_wmA091ne9_0),.clk(gclk));
	jdff dff_B_fs04zcVl2_0(.din(w_dff_B_wmA091ne9_0),.dout(w_dff_B_fs04zcVl2_0),.clk(gclk));
	jdff dff_B_3duPMmKT4_0(.din(w_dff_B_fs04zcVl2_0),.dout(w_dff_B_3duPMmKT4_0),.clk(gclk));
	jdff dff_B_0ST06S6Z7_0(.din(w_dff_B_3duPMmKT4_0),.dout(w_dff_B_0ST06S6Z7_0),.clk(gclk));
	jdff dff_B_gYw3T9cY7_0(.din(w_dff_B_0ST06S6Z7_0),.dout(w_dff_B_gYw3T9cY7_0),.clk(gclk));
	jdff dff_B_GdXnogvr7_1(.din(n1038),.dout(w_dff_B_GdXnogvr7_1),.clk(gclk));
	jdff dff_B_XQwIbR8p4_1(.din(w_dff_B_GdXnogvr7_1),.dout(w_dff_B_XQwIbR8p4_1),.clk(gclk));
	jdff dff_B_XRW2itrt9_1(.din(w_dff_B_XQwIbR8p4_1),.dout(w_dff_B_XRW2itrt9_1),.clk(gclk));
	jdff dff_B_W5fOSvQ24_1(.din(w_dff_B_XRW2itrt9_1),.dout(w_dff_B_W5fOSvQ24_1),.clk(gclk));
	jdff dff_B_cIPUVuF94_1(.din(w_dff_B_W5fOSvQ24_1),.dout(w_dff_B_cIPUVuF94_1),.clk(gclk));
	jdff dff_B_7XdPC3LR4_1(.din(w_dff_B_cIPUVuF94_1),.dout(w_dff_B_7XdPC3LR4_1),.clk(gclk));
	jdff dff_B_5T81fUaD8_1(.din(w_dff_B_7XdPC3LR4_1),.dout(w_dff_B_5T81fUaD8_1),.clk(gclk));
	jdff dff_B_8bQZlJOO0_1(.din(w_dff_B_5T81fUaD8_1),.dout(w_dff_B_8bQZlJOO0_1),.clk(gclk));
	jdff dff_B_XqgXzWwt8_1(.din(w_dff_B_8bQZlJOO0_1),.dout(w_dff_B_XqgXzWwt8_1),.clk(gclk));
	jdff dff_B_oftdZZa24_1(.din(w_dff_B_XqgXzWwt8_1),.dout(w_dff_B_oftdZZa24_1),.clk(gclk));
	jdff dff_B_tT9aN8G51_1(.din(w_dff_B_oftdZZa24_1),.dout(w_dff_B_tT9aN8G51_1),.clk(gclk));
	jdff dff_B_40NbgsGD4_1(.din(w_dff_B_tT9aN8G51_1),.dout(w_dff_B_40NbgsGD4_1),.clk(gclk));
	jdff dff_B_rvr7EOT11_1(.din(w_dff_B_40NbgsGD4_1),.dout(w_dff_B_rvr7EOT11_1),.clk(gclk));
	jdff dff_B_aKGcBlSp4_1(.din(w_dff_B_rvr7EOT11_1),.dout(w_dff_B_aKGcBlSp4_1),.clk(gclk));
	jdff dff_B_vcQiqavX5_1(.din(w_dff_B_aKGcBlSp4_1),.dout(w_dff_B_vcQiqavX5_1),.clk(gclk));
	jdff dff_B_mDKkOzfl8_1(.din(w_dff_B_vcQiqavX5_1),.dout(w_dff_B_mDKkOzfl8_1),.clk(gclk));
	jdff dff_B_qaB5zHrA2_1(.din(w_dff_B_mDKkOzfl8_1),.dout(w_dff_B_qaB5zHrA2_1),.clk(gclk));
	jdff dff_B_Jya1gP1o4_1(.din(w_dff_B_qaB5zHrA2_1),.dout(w_dff_B_Jya1gP1o4_1),.clk(gclk));
	jdff dff_B_OlbHQIYo5_1(.din(w_dff_B_Jya1gP1o4_1),.dout(w_dff_B_OlbHQIYo5_1),.clk(gclk));
	jdff dff_B_DvvFtIW32_1(.din(w_dff_B_OlbHQIYo5_1),.dout(w_dff_B_DvvFtIW32_1),.clk(gclk));
	jdff dff_B_WGVbmZp47_1(.din(w_dff_B_DvvFtIW32_1),.dout(w_dff_B_WGVbmZp47_1),.clk(gclk));
	jdff dff_B_Fpv9YHTV0_1(.din(w_dff_B_WGVbmZp47_1),.dout(w_dff_B_Fpv9YHTV0_1),.clk(gclk));
	jdff dff_B_6d2eINSq6_1(.din(w_dff_B_Fpv9YHTV0_1),.dout(w_dff_B_6d2eINSq6_1),.clk(gclk));
	jdff dff_B_aKp1oa0J7_1(.din(w_dff_B_6d2eINSq6_1),.dout(w_dff_B_aKp1oa0J7_1),.clk(gclk));
	jdff dff_B_0tMQlvNh4_1(.din(w_dff_B_aKp1oa0J7_1),.dout(w_dff_B_0tMQlvNh4_1),.clk(gclk));
	jdff dff_B_Ac7jinqw7_1(.din(w_dff_B_0tMQlvNh4_1),.dout(w_dff_B_Ac7jinqw7_1),.clk(gclk));
	jdff dff_B_VmsNyaTt1_1(.din(w_dff_B_Ac7jinqw7_1),.dout(w_dff_B_VmsNyaTt1_1),.clk(gclk));
	jdff dff_B_HGFYq3Nj1_1(.din(w_dff_B_VmsNyaTt1_1),.dout(w_dff_B_HGFYq3Nj1_1),.clk(gclk));
	jdff dff_B_LUdSKeJ88_1(.din(w_dff_B_HGFYq3Nj1_1),.dout(w_dff_B_LUdSKeJ88_1),.clk(gclk));
	jdff dff_B_7L2Keg130_1(.din(w_dff_B_LUdSKeJ88_1),.dout(w_dff_B_7L2Keg130_1),.clk(gclk));
	jdff dff_B_kLnz6kAV0_1(.din(w_dff_B_7L2Keg130_1),.dout(w_dff_B_kLnz6kAV0_1),.clk(gclk));
	jdff dff_B_yOOvbO6P0_1(.din(w_dff_B_kLnz6kAV0_1),.dout(w_dff_B_yOOvbO6P0_1),.clk(gclk));
	jdff dff_B_PbUxpgOp0_1(.din(w_dff_B_yOOvbO6P0_1),.dout(w_dff_B_PbUxpgOp0_1),.clk(gclk));
	jdff dff_B_VBS6iIeL7_1(.din(w_dff_B_PbUxpgOp0_1),.dout(w_dff_B_VBS6iIeL7_1),.clk(gclk));
	jdff dff_B_U0YrBBnK6_1(.din(w_dff_B_VBS6iIeL7_1),.dout(w_dff_B_U0YrBBnK6_1),.clk(gclk));
	jdff dff_B_nE5ZQDb68_1(.din(w_dff_B_U0YrBBnK6_1),.dout(w_dff_B_nE5ZQDb68_1),.clk(gclk));
	jdff dff_B_9gi2erYH8_1(.din(w_dff_B_nE5ZQDb68_1),.dout(w_dff_B_9gi2erYH8_1),.clk(gclk));
	jdff dff_B_70vy9pFs4_1(.din(w_dff_B_9gi2erYH8_1),.dout(w_dff_B_70vy9pFs4_1),.clk(gclk));
	jdff dff_B_YLQZl8bD2_1(.din(w_dff_B_70vy9pFs4_1),.dout(w_dff_B_YLQZl8bD2_1),.clk(gclk));
	jdff dff_B_DrxjVXPS8_1(.din(w_dff_B_YLQZl8bD2_1),.dout(w_dff_B_DrxjVXPS8_1),.clk(gclk));
	jdff dff_B_gicHjYTq4_1(.din(w_dff_B_DrxjVXPS8_1),.dout(w_dff_B_gicHjYTq4_1),.clk(gclk));
	jdff dff_B_IC5KiwpU8_1(.din(w_dff_B_gicHjYTq4_1),.dout(w_dff_B_IC5KiwpU8_1),.clk(gclk));
	jdff dff_B_LCAQhOok8_1(.din(w_dff_B_IC5KiwpU8_1),.dout(w_dff_B_LCAQhOok8_1),.clk(gclk));
	jdff dff_B_Lcdse3FY4_1(.din(w_dff_B_LCAQhOok8_1),.dout(w_dff_B_Lcdse3FY4_1),.clk(gclk));
	jdff dff_B_BEtKi7yH2_1(.din(w_dff_B_Lcdse3FY4_1),.dout(w_dff_B_BEtKi7yH2_1),.clk(gclk));
	jdff dff_B_20XgnWZD6_1(.din(w_dff_B_BEtKi7yH2_1),.dout(w_dff_B_20XgnWZD6_1),.clk(gclk));
	jdff dff_B_7tWUc2sC8_1(.din(w_dff_B_20XgnWZD6_1),.dout(w_dff_B_7tWUc2sC8_1),.clk(gclk));
	jdff dff_B_MbLVCZ504_1(.din(w_dff_B_7tWUc2sC8_1),.dout(w_dff_B_MbLVCZ504_1),.clk(gclk));
	jdff dff_B_sj3oHv8P8_1(.din(w_dff_B_MbLVCZ504_1),.dout(w_dff_B_sj3oHv8P8_1),.clk(gclk));
	jdff dff_B_1SWLi7Mg2_1(.din(w_dff_B_sj3oHv8P8_1),.dout(w_dff_B_1SWLi7Mg2_1),.clk(gclk));
	jdff dff_B_BynzUjIH6_1(.din(w_dff_B_1SWLi7Mg2_1),.dout(w_dff_B_BynzUjIH6_1),.clk(gclk));
	jdff dff_B_lWhhEMYP5_1(.din(w_dff_B_BynzUjIH6_1),.dout(w_dff_B_lWhhEMYP5_1),.clk(gclk));
	jdff dff_B_RebZUSRG0_1(.din(w_dff_B_lWhhEMYP5_1),.dout(w_dff_B_RebZUSRG0_1),.clk(gclk));
	jdff dff_B_dEw66dmo6_1(.din(w_dff_B_RebZUSRG0_1),.dout(w_dff_B_dEw66dmo6_1),.clk(gclk));
	jdff dff_B_08QWJ17r5_1(.din(w_dff_B_dEw66dmo6_1),.dout(w_dff_B_08QWJ17r5_1),.clk(gclk));
	jdff dff_B_e10YDfn47_1(.din(w_dff_B_08QWJ17r5_1),.dout(w_dff_B_e10YDfn47_1),.clk(gclk));
	jdff dff_B_WWg7wf7O1_1(.din(w_dff_B_e10YDfn47_1),.dout(w_dff_B_WWg7wf7O1_1),.clk(gclk));
	jdff dff_B_7u2dcfEg9_1(.din(w_dff_B_WWg7wf7O1_1),.dout(w_dff_B_7u2dcfEg9_1),.clk(gclk));
	jdff dff_B_5lpFBKTS5_1(.din(w_dff_B_7u2dcfEg9_1),.dout(w_dff_B_5lpFBKTS5_1),.clk(gclk));
	jdff dff_B_YdZFmXL88_1(.din(w_dff_B_5lpFBKTS5_1),.dout(w_dff_B_YdZFmXL88_1),.clk(gclk));
	jdff dff_B_JfFWg1iW5_1(.din(w_dff_B_YdZFmXL88_1),.dout(w_dff_B_JfFWg1iW5_1),.clk(gclk));
	jdff dff_B_Uk3Po1dr8_1(.din(w_dff_B_JfFWg1iW5_1),.dout(w_dff_B_Uk3Po1dr8_1),.clk(gclk));
	jdff dff_B_8Mb32oqK2_1(.din(w_dff_B_Uk3Po1dr8_1),.dout(w_dff_B_8Mb32oqK2_1),.clk(gclk));
	jdff dff_B_0Wk9LVZs3_1(.din(w_dff_B_8Mb32oqK2_1),.dout(w_dff_B_0Wk9LVZs3_1),.clk(gclk));
	jdff dff_B_wuCGhu0J9_1(.din(w_dff_B_0Wk9LVZs3_1),.dout(w_dff_B_wuCGhu0J9_1),.clk(gclk));
	jdff dff_B_QHXnIcX82_1(.din(w_dff_B_wuCGhu0J9_1),.dout(w_dff_B_QHXnIcX82_1),.clk(gclk));
	jdff dff_B_z7rfscAq7_1(.din(w_dff_B_QHXnIcX82_1),.dout(w_dff_B_z7rfscAq7_1),.clk(gclk));
	jdff dff_B_Uq6s8GXI7_1(.din(w_dff_B_z7rfscAq7_1),.dout(w_dff_B_Uq6s8GXI7_1),.clk(gclk));
	jdff dff_B_gbo5BqUI5_1(.din(w_dff_B_Uq6s8GXI7_1),.dout(w_dff_B_gbo5BqUI5_1),.clk(gclk));
	jdff dff_B_ecgcdOhE0_1(.din(w_dff_B_gbo5BqUI5_1),.dout(w_dff_B_ecgcdOhE0_1),.clk(gclk));
	jdff dff_B_ijMlERTJ4_1(.din(w_dff_B_ecgcdOhE0_1),.dout(w_dff_B_ijMlERTJ4_1),.clk(gclk));
	jdff dff_B_ipn2A3FN3_1(.din(w_dff_B_ijMlERTJ4_1),.dout(w_dff_B_ipn2A3FN3_1),.clk(gclk));
	jdff dff_B_Wb3hR7mj1_1(.din(w_dff_B_ipn2A3FN3_1),.dout(w_dff_B_Wb3hR7mj1_1),.clk(gclk));
	jdff dff_B_LnGiy3TB1_1(.din(w_dff_B_Wb3hR7mj1_1),.dout(w_dff_B_LnGiy3TB1_1),.clk(gclk));
	jdff dff_B_eLaz2e8v5_1(.din(w_dff_B_LnGiy3TB1_1),.dout(w_dff_B_eLaz2e8v5_1),.clk(gclk));
	jdff dff_B_WCavkgzK5_1(.din(w_dff_B_eLaz2e8v5_1),.dout(w_dff_B_WCavkgzK5_1),.clk(gclk));
	jdff dff_B_PvztYaNT4_1(.din(w_dff_B_WCavkgzK5_1),.dout(w_dff_B_PvztYaNT4_1),.clk(gclk));
	jdff dff_B_0jZGnh2v2_1(.din(w_dff_B_PvztYaNT4_1),.dout(w_dff_B_0jZGnh2v2_1),.clk(gclk));
	jdff dff_B_EGczUprh7_1(.din(w_dff_B_0jZGnh2v2_1),.dout(w_dff_B_EGczUprh7_1),.clk(gclk));
	jdff dff_B_6Lyd6ATI7_1(.din(w_dff_B_EGczUprh7_1),.dout(w_dff_B_6Lyd6ATI7_1),.clk(gclk));
	jdff dff_B_MQg2O00O6_1(.din(w_dff_B_6Lyd6ATI7_1),.dout(w_dff_B_MQg2O00O6_1),.clk(gclk));
	jdff dff_B_vQT0tWoq5_1(.din(w_dff_B_MQg2O00O6_1),.dout(w_dff_B_vQT0tWoq5_1),.clk(gclk));
	jdff dff_B_l3qwcyBC1_1(.din(w_dff_B_vQT0tWoq5_1),.dout(w_dff_B_l3qwcyBC1_1),.clk(gclk));
	jdff dff_B_CRG8t1ah8_1(.din(w_dff_B_l3qwcyBC1_1),.dout(w_dff_B_CRG8t1ah8_1),.clk(gclk));
	jdff dff_B_LNlJZs1C4_1(.din(w_dff_B_CRG8t1ah8_1),.dout(w_dff_B_LNlJZs1C4_1),.clk(gclk));
	jdff dff_B_IWux2oHZ9_1(.din(w_dff_B_LNlJZs1C4_1),.dout(w_dff_B_IWux2oHZ9_1),.clk(gclk));
	jdff dff_B_hxw07n0o8_1(.din(w_dff_B_IWux2oHZ9_1),.dout(w_dff_B_hxw07n0o8_1),.clk(gclk));
	jdff dff_B_Jx6ohcKw2_1(.din(w_dff_B_hxw07n0o8_1),.dout(w_dff_B_Jx6ohcKw2_1),.clk(gclk));
	jdff dff_B_pldm7iwc9_1(.din(w_dff_B_Jx6ohcKw2_1),.dout(w_dff_B_pldm7iwc9_1),.clk(gclk));
	jdff dff_B_Ey1Bv6j82_1(.din(w_dff_B_pldm7iwc9_1),.dout(w_dff_B_Ey1Bv6j82_1),.clk(gclk));
	jdff dff_B_V78sD6Ie7_1(.din(w_dff_B_Ey1Bv6j82_1),.dout(w_dff_B_V78sD6Ie7_1),.clk(gclk));
	jdff dff_B_rj64pd9j9_1(.din(w_dff_B_V78sD6Ie7_1),.dout(w_dff_B_rj64pd9j9_1),.clk(gclk));
	jdff dff_B_amElfdG16_1(.din(w_dff_B_rj64pd9j9_1),.dout(w_dff_B_amElfdG16_1),.clk(gclk));
	jdff dff_B_lH6RBAX57_1(.din(w_dff_B_amElfdG16_1),.dout(w_dff_B_lH6RBAX57_1),.clk(gclk));
	jdff dff_B_cxCprxkp4_1(.din(w_dff_B_lH6RBAX57_1),.dout(w_dff_B_cxCprxkp4_1),.clk(gclk));
	jdff dff_B_eBYFtK4C2_1(.din(w_dff_B_cxCprxkp4_1),.dout(w_dff_B_eBYFtK4C2_1),.clk(gclk));
	jdff dff_B_oq2MWXEb3_1(.din(w_dff_B_eBYFtK4C2_1),.dout(w_dff_B_oq2MWXEb3_1),.clk(gclk));
	jdff dff_B_ievQsVz30_1(.din(w_dff_B_oq2MWXEb3_1),.dout(w_dff_B_ievQsVz30_1),.clk(gclk));
	jdff dff_B_EMh02utm5_1(.din(w_dff_B_ievQsVz30_1),.dout(w_dff_B_EMh02utm5_1),.clk(gclk));
	jdff dff_B_1N4e48Hr0_1(.din(w_dff_B_EMh02utm5_1),.dout(w_dff_B_1N4e48Hr0_1),.clk(gclk));
	jdff dff_B_2rj0tbAx3_1(.din(w_dff_B_1N4e48Hr0_1),.dout(w_dff_B_2rj0tbAx3_1),.clk(gclk));
	jdff dff_B_3cLY4mMu9_1(.din(w_dff_B_2rj0tbAx3_1),.dout(w_dff_B_3cLY4mMu9_1),.clk(gclk));
	jdff dff_B_lPQkhTh67_1(.din(w_dff_B_3cLY4mMu9_1),.dout(w_dff_B_lPQkhTh67_1),.clk(gclk));
	jdff dff_B_vzwRcvaQ5_1(.din(w_dff_B_lPQkhTh67_1),.dout(w_dff_B_vzwRcvaQ5_1),.clk(gclk));
	jdff dff_B_47jZaQhx6_1(.din(w_dff_B_vzwRcvaQ5_1),.dout(w_dff_B_47jZaQhx6_1),.clk(gclk));
	jdff dff_B_KQtw1Zjg3_1(.din(w_dff_B_47jZaQhx6_1),.dout(w_dff_B_KQtw1Zjg3_1),.clk(gclk));
	jdff dff_B_ji1m2Zy14_1(.din(w_dff_B_KQtw1Zjg3_1),.dout(w_dff_B_ji1m2Zy14_1),.clk(gclk));
	jdff dff_B_Zeu5QyPt7_1(.din(w_dff_B_ji1m2Zy14_1),.dout(w_dff_B_Zeu5QyPt7_1),.clk(gclk));
	jdff dff_B_mscM20U91_1(.din(w_dff_B_Zeu5QyPt7_1),.dout(w_dff_B_mscM20U91_1),.clk(gclk));
	jdff dff_B_OjgH8gAT8_0(.din(n1039),.dout(w_dff_B_OjgH8gAT8_0),.clk(gclk));
	jdff dff_B_TQ78zH5j3_0(.din(w_dff_B_OjgH8gAT8_0),.dout(w_dff_B_TQ78zH5j3_0),.clk(gclk));
	jdff dff_B_K24HpLYV1_0(.din(w_dff_B_TQ78zH5j3_0),.dout(w_dff_B_K24HpLYV1_0),.clk(gclk));
	jdff dff_B_R63ClVW62_0(.din(w_dff_B_K24HpLYV1_0),.dout(w_dff_B_R63ClVW62_0),.clk(gclk));
	jdff dff_B_ELKXiSbI5_0(.din(w_dff_B_R63ClVW62_0),.dout(w_dff_B_ELKXiSbI5_0),.clk(gclk));
	jdff dff_B_GTop6alx5_0(.din(w_dff_B_ELKXiSbI5_0),.dout(w_dff_B_GTop6alx5_0),.clk(gclk));
	jdff dff_B_isnod7H93_0(.din(w_dff_B_GTop6alx5_0),.dout(w_dff_B_isnod7H93_0),.clk(gclk));
	jdff dff_B_hYN94gql4_0(.din(w_dff_B_isnod7H93_0),.dout(w_dff_B_hYN94gql4_0),.clk(gclk));
	jdff dff_B_TYDkehFz3_0(.din(w_dff_B_hYN94gql4_0),.dout(w_dff_B_TYDkehFz3_0),.clk(gclk));
	jdff dff_B_1R1iEFKn7_0(.din(w_dff_B_TYDkehFz3_0),.dout(w_dff_B_1R1iEFKn7_0),.clk(gclk));
	jdff dff_B_hc0wCGcQ3_0(.din(w_dff_B_1R1iEFKn7_0),.dout(w_dff_B_hc0wCGcQ3_0),.clk(gclk));
	jdff dff_B_0kox4D0f8_0(.din(w_dff_B_hc0wCGcQ3_0),.dout(w_dff_B_0kox4D0f8_0),.clk(gclk));
	jdff dff_B_fSunZdvb8_0(.din(w_dff_B_0kox4D0f8_0),.dout(w_dff_B_fSunZdvb8_0),.clk(gclk));
	jdff dff_B_br6IXRvj1_0(.din(w_dff_B_fSunZdvb8_0),.dout(w_dff_B_br6IXRvj1_0),.clk(gclk));
	jdff dff_B_s0DMGbSC6_0(.din(w_dff_B_br6IXRvj1_0),.dout(w_dff_B_s0DMGbSC6_0),.clk(gclk));
	jdff dff_B_9lKQl8VW9_0(.din(w_dff_B_s0DMGbSC6_0),.dout(w_dff_B_9lKQl8VW9_0),.clk(gclk));
	jdff dff_B_yke4QKy12_0(.din(w_dff_B_9lKQl8VW9_0),.dout(w_dff_B_yke4QKy12_0),.clk(gclk));
	jdff dff_B_aah6ulmI7_0(.din(w_dff_B_yke4QKy12_0),.dout(w_dff_B_aah6ulmI7_0),.clk(gclk));
	jdff dff_B_04M2D68W8_0(.din(w_dff_B_aah6ulmI7_0),.dout(w_dff_B_04M2D68W8_0),.clk(gclk));
	jdff dff_B_rZvBXlim7_0(.din(w_dff_B_04M2D68W8_0),.dout(w_dff_B_rZvBXlim7_0),.clk(gclk));
	jdff dff_B_zD41bNiG7_0(.din(w_dff_B_rZvBXlim7_0),.dout(w_dff_B_zD41bNiG7_0),.clk(gclk));
	jdff dff_B_lkQPnXny1_0(.din(w_dff_B_zD41bNiG7_0),.dout(w_dff_B_lkQPnXny1_0),.clk(gclk));
	jdff dff_B_AMlU3bff0_0(.din(w_dff_B_lkQPnXny1_0),.dout(w_dff_B_AMlU3bff0_0),.clk(gclk));
	jdff dff_B_ih9AxHTJ2_0(.din(w_dff_B_AMlU3bff0_0),.dout(w_dff_B_ih9AxHTJ2_0),.clk(gclk));
	jdff dff_B_xvhPIzqt6_0(.din(w_dff_B_ih9AxHTJ2_0),.dout(w_dff_B_xvhPIzqt6_0),.clk(gclk));
	jdff dff_B_Uchh0Bas0_0(.din(w_dff_B_xvhPIzqt6_0),.dout(w_dff_B_Uchh0Bas0_0),.clk(gclk));
	jdff dff_B_PEgbaQ6E7_0(.din(w_dff_B_Uchh0Bas0_0),.dout(w_dff_B_PEgbaQ6E7_0),.clk(gclk));
	jdff dff_B_K10P0fQr3_0(.din(w_dff_B_PEgbaQ6E7_0),.dout(w_dff_B_K10P0fQr3_0),.clk(gclk));
	jdff dff_B_P15aDoTu2_0(.din(w_dff_B_K10P0fQr3_0),.dout(w_dff_B_P15aDoTu2_0),.clk(gclk));
	jdff dff_B_SCaMJe4u7_0(.din(w_dff_B_P15aDoTu2_0),.dout(w_dff_B_SCaMJe4u7_0),.clk(gclk));
	jdff dff_B_Nd7Fues73_0(.din(w_dff_B_SCaMJe4u7_0),.dout(w_dff_B_Nd7Fues73_0),.clk(gclk));
	jdff dff_B_Z1ueymbs7_0(.din(w_dff_B_Nd7Fues73_0),.dout(w_dff_B_Z1ueymbs7_0),.clk(gclk));
	jdff dff_B_nuJkUSOm2_0(.din(w_dff_B_Z1ueymbs7_0),.dout(w_dff_B_nuJkUSOm2_0),.clk(gclk));
	jdff dff_B_XaRpYCAd6_0(.din(w_dff_B_nuJkUSOm2_0),.dout(w_dff_B_XaRpYCAd6_0),.clk(gclk));
	jdff dff_B_6Df0zqfJ4_0(.din(w_dff_B_XaRpYCAd6_0),.dout(w_dff_B_6Df0zqfJ4_0),.clk(gclk));
	jdff dff_B_dtFngcJS1_0(.din(w_dff_B_6Df0zqfJ4_0),.dout(w_dff_B_dtFngcJS1_0),.clk(gclk));
	jdff dff_B_dCvPrrXy3_0(.din(w_dff_B_dtFngcJS1_0),.dout(w_dff_B_dCvPrrXy3_0),.clk(gclk));
	jdff dff_B_ihgSkygg2_0(.din(w_dff_B_dCvPrrXy3_0),.dout(w_dff_B_ihgSkygg2_0),.clk(gclk));
	jdff dff_B_DwdcsoqK5_0(.din(w_dff_B_ihgSkygg2_0),.dout(w_dff_B_DwdcsoqK5_0),.clk(gclk));
	jdff dff_B_vZ2dBD3F2_0(.din(w_dff_B_DwdcsoqK5_0),.dout(w_dff_B_vZ2dBD3F2_0),.clk(gclk));
	jdff dff_B_ALJcwdXU8_0(.din(w_dff_B_vZ2dBD3F2_0),.dout(w_dff_B_ALJcwdXU8_0),.clk(gclk));
	jdff dff_B_h4lfzINb3_0(.din(w_dff_B_ALJcwdXU8_0),.dout(w_dff_B_h4lfzINb3_0),.clk(gclk));
	jdff dff_B_uVu2H0jH1_0(.din(w_dff_B_h4lfzINb3_0),.dout(w_dff_B_uVu2H0jH1_0),.clk(gclk));
	jdff dff_B_oK6EAMFd5_0(.din(w_dff_B_uVu2H0jH1_0),.dout(w_dff_B_oK6EAMFd5_0),.clk(gclk));
	jdff dff_B_szAD2Rne6_0(.din(w_dff_B_oK6EAMFd5_0),.dout(w_dff_B_szAD2Rne6_0),.clk(gclk));
	jdff dff_B_V8BeWNtC3_0(.din(w_dff_B_szAD2Rne6_0),.dout(w_dff_B_V8BeWNtC3_0),.clk(gclk));
	jdff dff_B_pgydElYJ8_0(.din(w_dff_B_V8BeWNtC3_0),.dout(w_dff_B_pgydElYJ8_0),.clk(gclk));
	jdff dff_B_LDp9m6jh6_0(.din(w_dff_B_pgydElYJ8_0),.dout(w_dff_B_LDp9m6jh6_0),.clk(gclk));
	jdff dff_B_253hTXaZ8_0(.din(w_dff_B_LDp9m6jh6_0),.dout(w_dff_B_253hTXaZ8_0),.clk(gclk));
	jdff dff_B_shgoIpAe2_0(.din(w_dff_B_253hTXaZ8_0),.dout(w_dff_B_shgoIpAe2_0),.clk(gclk));
	jdff dff_B_JjU0kbAT0_0(.din(w_dff_B_shgoIpAe2_0),.dout(w_dff_B_JjU0kbAT0_0),.clk(gclk));
	jdff dff_B_Nyf1tyS72_0(.din(w_dff_B_JjU0kbAT0_0),.dout(w_dff_B_Nyf1tyS72_0),.clk(gclk));
	jdff dff_B_EVOVZtAd7_0(.din(w_dff_B_Nyf1tyS72_0),.dout(w_dff_B_EVOVZtAd7_0),.clk(gclk));
	jdff dff_B_lSezfx319_0(.din(w_dff_B_EVOVZtAd7_0),.dout(w_dff_B_lSezfx319_0),.clk(gclk));
	jdff dff_B_EeTvjZ833_0(.din(w_dff_B_lSezfx319_0),.dout(w_dff_B_EeTvjZ833_0),.clk(gclk));
	jdff dff_B_E1nOEVE68_0(.din(w_dff_B_EeTvjZ833_0),.dout(w_dff_B_E1nOEVE68_0),.clk(gclk));
	jdff dff_B_1mmysII87_0(.din(w_dff_B_E1nOEVE68_0),.dout(w_dff_B_1mmysII87_0),.clk(gclk));
	jdff dff_B_Z1nAeDqs7_0(.din(w_dff_B_1mmysII87_0),.dout(w_dff_B_Z1nAeDqs7_0),.clk(gclk));
	jdff dff_B_jiqGkYTx0_0(.din(w_dff_B_Z1nAeDqs7_0),.dout(w_dff_B_jiqGkYTx0_0),.clk(gclk));
	jdff dff_B_QXsj9D0E1_0(.din(w_dff_B_jiqGkYTx0_0),.dout(w_dff_B_QXsj9D0E1_0),.clk(gclk));
	jdff dff_B_NLb17XNZ9_0(.din(w_dff_B_QXsj9D0E1_0),.dout(w_dff_B_NLb17XNZ9_0),.clk(gclk));
	jdff dff_B_6IIpGqTX5_0(.din(w_dff_B_NLb17XNZ9_0),.dout(w_dff_B_6IIpGqTX5_0),.clk(gclk));
	jdff dff_B_0vwFyDdw3_0(.din(w_dff_B_6IIpGqTX5_0),.dout(w_dff_B_0vwFyDdw3_0),.clk(gclk));
	jdff dff_B_NkBj7BcQ2_0(.din(w_dff_B_0vwFyDdw3_0),.dout(w_dff_B_NkBj7BcQ2_0),.clk(gclk));
	jdff dff_B_DZerjOCU2_0(.din(w_dff_B_NkBj7BcQ2_0),.dout(w_dff_B_DZerjOCU2_0),.clk(gclk));
	jdff dff_B_uKsc8miY8_0(.din(w_dff_B_DZerjOCU2_0),.dout(w_dff_B_uKsc8miY8_0),.clk(gclk));
	jdff dff_B_jZYYgkKq1_0(.din(w_dff_B_uKsc8miY8_0),.dout(w_dff_B_jZYYgkKq1_0),.clk(gclk));
	jdff dff_B_H8ickXxF7_0(.din(w_dff_B_jZYYgkKq1_0),.dout(w_dff_B_H8ickXxF7_0),.clk(gclk));
	jdff dff_B_A8pRry767_0(.din(w_dff_B_H8ickXxF7_0),.dout(w_dff_B_A8pRry767_0),.clk(gclk));
	jdff dff_B_GWmOgk2V0_0(.din(w_dff_B_A8pRry767_0),.dout(w_dff_B_GWmOgk2V0_0),.clk(gclk));
	jdff dff_B_rnm3cO2Q2_0(.din(w_dff_B_GWmOgk2V0_0),.dout(w_dff_B_rnm3cO2Q2_0),.clk(gclk));
	jdff dff_B_0eO1sDOQ9_0(.din(w_dff_B_rnm3cO2Q2_0),.dout(w_dff_B_0eO1sDOQ9_0),.clk(gclk));
	jdff dff_B_Arb0ROCA4_0(.din(w_dff_B_0eO1sDOQ9_0),.dout(w_dff_B_Arb0ROCA4_0),.clk(gclk));
	jdff dff_B_hETQgg9q5_0(.din(w_dff_B_Arb0ROCA4_0),.dout(w_dff_B_hETQgg9q5_0),.clk(gclk));
	jdff dff_B_bbwbSTyP8_0(.din(w_dff_B_hETQgg9q5_0),.dout(w_dff_B_bbwbSTyP8_0),.clk(gclk));
	jdff dff_B_X6Gir7cf1_0(.din(w_dff_B_bbwbSTyP8_0),.dout(w_dff_B_X6Gir7cf1_0),.clk(gclk));
	jdff dff_B_L7CtLO6o6_0(.din(w_dff_B_X6Gir7cf1_0),.dout(w_dff_B_L7CtLO6o6_0),.clk(gclk));
	jdff dff_B_K2JIZ6ZI1_0(.din(w_dff_B_L7CtLO6o6_0),.dout(w_dff_B_K2JIZ6ZI1_0),.clk(gclk));
	jdff dff_B_uMd8AryD2_0(.din(w_dff_B_K2JIZ6ZI1_0),.dout(w_dff_B_uMd8AryD2_0),.clk(gclk));
	jdff dff_B_GrNRIarL1_0(.din(w_dff_B_uMd8AryD2_0),.dout(w_dff_B_GrNRIarL1_0),.clk(gclk));
	jdff dff_B_5Rpe5MKA3_0(.din(w_dff_B_GrNRIarL1_0),.dout(w_dff_B_5Rpe5MKA3_0),.clk(gclk));
	jdff dff_B_25jn3B9A7_0(.din(w_dff_B_5Rpe5MKA3_0),.dout(w_dff_B_25jn3B9A7_0),.clk(gclk));
	jdff dff_B_P9VzfJ9J9_0(.din(w_dff_B_25jn3B9A7_0),.dout(w_dff_B_P9VzfJ9J9_0),.clk(gclk));
	jdff dff_B_KN53MaCM1_0(.din(w_dff_B_P9VzfJ9J9_0),.dout(w_dff_B_KN53MaCM1_0),.clk(gclk));
	jdff dff_B_2XawnBzw4_0(.din(w_dff_B_KN53MaCM1_0),.dout(w_dff_B_2XawnBzw4_0),.clk(gclk));
	jdff dff_B_k9FJG9Do2_0(.din(w_dff_B_2XawnBzw4_0),.dout(w_dff_B_k9FJG9Do2_0),.clk(gclk));
	jdff dff_B_TArSJXeg5_0(.din(w_dff_B_k9FJG9Do2_0),.dout(w_dff_B_TArSJXeg5_0),.clk(gclk));
	jdff dff_B_qY3vTnCq5_0(.din(w_dff_B_TArSJXeg5_0),.dout(w_dff_B_qY3vTnCq5_0),.clk(gclk));
	jdff dff_B_toHFjzK43_0(.din(w_dff_B_qY3vTnCq5_0),.dout(w_dff_B_toHFjzK43_0),.clk(gclk));
	jdff dff_B_UtQbRfGY3_0(.din(w_dff_B_toHFjzK43_0),.dout(w_dff_B_UtQbRfGY3_0),.clk(gclk));
	jdff dff_B_qnPVfik00_0(.din(w_dff_B_UtQbRfGY3_0),.dout(w_dff_B_qnPVfik00_0),.clk(gclk));
	jdff dff_B_ZGFz7tMl6_0(.din(w_dff_B_qnPVfik00_0),.dout(w_dff_B_ZGFz7tMl6_0),.clk(gclk));
	jdff dff_B_Ml1jO7Ic0_0(.din(w_dff_B_ZGFz7tMl6_0),.dout(w_dff_B_Ml1jO7Ic0_0),.clk(gclk));
	jdff dff_B_QRC27lcQ5_0(.din(w_dff_B_Ml1jO7Ic0_0),.dout(w_dff_B_QRC27lcQ5_0),.clk(gclk));
	jdff dff_B_FJ4WNLA39_0(.din(w_dff_B_QRC27lcQ5_0),.dout(w_dff_B_FJ4WNLA39_0),.clk(gclk));
	jdff dff_B_Lbc52OQP8_0(.din(w_dff_B_FJ4WNLA39_0),.dout(w_dff_B_Lbc52OQP8_0),.clk(gclk));
	jdff dff_B_Y5afw0ZB8_0(.din(w_dff_B_Lbc52OQP8_0),.dout(w_dff_B_Y5afw0ZB8_0),.clk(gclk));
	jdff dff_B_LpU5trMT0_0(.din(w_dff_B_Y5afw0ZB8_0),.dout(w_dff_B_LpU5trMT0_0),.clk(gclk));
	jdff dff_B_eRQIpvKz8_0(.din(w_dff_B_LpU5trMT0_0),.dout(w_dff_B_eRQIpvKz8_0),.clk(gclk));
	jdff dff_B_0Z7hCwz47_0(.din(w_dff_B_eRQIpvKz8_0),.dout(w_dff_B_0Z7hCwz47_0),.clk(gclk));
	jdff dff_B_o4Svj9Vj3_0(.din(w_dff_B_0Z7hCwz47_0),.dout(w_dff_B_o4Svj9Vj3_0),.clk(gclk));
	jdff dff_B_HIERyfhj0_0(.din(w_dff_B_o4Svj9Vj3_0),.dout(w_dff_B_HIERyfhj0_0),.clk(gclk));
	jdff dff_B_s6bl0pUF6_0(.din(w_dff_B_HIERyfhj0_0),.dout(w_dff_B_s6bl0pUF6_0),.clk(gclk));
	jdff dff_B_BbZnq9aI1_0(.din(w_dff_B_s6bl0pUF6_0),.dout(w_dff_B_BbZnq9aI1_0),.clk(gclk));
	jdff dff_B_AVz3ik2a7_0(.din(w_dff_B_BbZnq9aI1_0),.dout(w_dff_B_AVz3ik2a7_0),.clk(gclk));
	jdff dff_B_6W81Yg0D1_0(.din(w_dff_B_AVz3ik2a7_0),.dout(w_dff_B_6W81Yg0D1_0),.clk(gclk));
	jdff dff_B_LJocUySI0_0(.din(w_dff_B_6W81Yg0D1_0),.dout(w_dff_B_LJocUySI0_0),.clk(gclk));
	jdff dff_B_CZKMbq7t9_0(.din(w_dff_B_LJocUySI0_0),.dout(w_dff_B_CZKMbq7t9_0),.clk(gclk));
	jdff dff_B_C9QaqcpL4_0(.din(w_dff_B_CZKMbq7t9_0),.dout(w_dff_B_C9QaqcpL4_0),.clk(gclk));
	jdff dff_B_bFVN0Qed9_1(.din(n1032),.dout(w_dff_B_bFVN0Qed9_1),.clk(gclk));
	jdff dff_B_HSBDnd5v7_1(.din(w_dff_B_bFVN0Qed9_1),.dout(w_dff_B_HSBDnd5v7_1),.clk(gclk));
	jdff dff_B_gWDft5LV8_1(.din(w_dff_B_HSBDnd5v7_1),.dout(w_dff_B_gWDft5LV8_1),.clk(gclk));
	jdff dff_B_KN7UEH1d6_1(.din(w_dff_B_gWDft5LV8_1),.dout(w_dff_B_KN7UEH1d6_1),.clk(gclk));
	jdff dff_B_IoYVsFeU4_1(.din(w_dff_B_KN7UEH1d6_1),.dout(w_dff_B_IoYVsFeU4_1),.clk(gclk));
	jdff dff_B_Ko52s5Hi0_1(.din(w_dff_B_IoYVsFeU4_1),.dout(w_dff_B_Ko52s5Hi0_1),.clk(gclk));
	jdff dff_B_wXNFg8NA9_1(.din(w_dff_B_Ko52s5Hi0_1),.dout(w_dff_B_wXNFg8NA9_1),.clk(gclk));
	jdff dff_B_cAPzcAbI6_1(.din(w_dff_B_wXNFg8NA9_1),.dout(w_dff_B_cAPzcAbI6_1),.clk(gclk));
	jdff dff_B_HyxNk1rF9_1(.din(w_dff_B_cAPzcAbI6_1),.dout(w_dff_B_HyxNk1rF9_1),.clk(gclk));
	jdff dff_B_leZFrgEh6_1(.din(w_dff_B_HyxNk1rF9_1),.dout(w_dff_B_leZFrgEh6_1),.clk(gclk));
	jdff dff_B_DN4pplCX5_1(.din(w_dff_B_leZFrgEh6_1),.dout(w_dff_B_DN4pplCX5_1),.clk(gclk));
	jdff dff_B_xXPd4XLS3_1(.din(w_dff_B_DN4pplCX5_1),.dout(w_dff_B_xXPd4XLS3_1),.clk(gclk));
	jdff dff_B_pY5DrhnD9_1(.din(w_dff_B_xXPd4XLS3_1),.dout(w_dff_B_pY5DrhnD9_1),.clk(gclk));
	jdff dff_B_ntVByL6G6_1(.din(w_dff_B_pY5DrhnD9_1),.dout(w_dff_B_ntVByL6G6_1),.clk(gclk));
	jdff dff_B_3RDIIUFW3_1(.din(w_dff_B_ntVByL6G6_1),.dout(w_dff_B_3RDIIUFW3_1),.clk(gclk));
	jdff dff_B_jtTKa6VD9_1(.din(w_dff_B_3RDIIUFW3_1),.dout(w_dff_B_jtTKa6VD9_1),.clk(gclk));
	jdff dff_B_nhs8tYnY3_1(.din(w_dff_B_jtTKa6VD9_1),.dout(w_dff_B_nhs8tYnY3_1),.clk(gclk));
	jdff dff_B_vZ7nAznE0_1(.din(w_dff_B_nhs8tYnY3_1),.dout(w_dff_B_vZ7nAznE0_1),.clk(gclk));
	jdff dff_B_kY1zTx6Z7_1(.din(w_dff_B_vZ7nAznE0_1),.dout(w_dff_B_kY1zTx6Z7_1),.clk(gclk));
	jdff dff_B_jWKVX2Bb9_1(.din(w_dff_B_kY1zTx6Z7_1),.dout(w_dff_B_jWKVX2Bb9_1),.clk(gclk));
	jdff dff_B_Pm851Ymt1_1(.din(w_dff_B_jWKVX2Bb9_1),.dout(w_dff_B_Pm851Ymt1_1),.clk(gclk));
	jdff dff_B_k3WSiMb69_1(.din(w_dff_B_Pm851Ymt1_1),.dout(w_dff_B_k3WSiMb69_1),.clk(gclk));
	jdff dff_B_z7az5cOA5_1(.din(w_dff_B_k3WSiMb69_1),.dout(w_dff_B_z7az5cOA5_1),.clk(gclk));
	jdff dff_B_9jCkwasi9_1(.din(w_dff_B_z7az5cOA5_1),.dout(w_dff_B_9jCkwasi9_1),.clk(gclk));
	jdff dff_B_8SKuRgD08_1(.din(w_dff_B_9jCkwasi9_1),.dout(w_dff_B_8SKuRgD08_1),.clk(gclk));
	jdff dff_B_WQO8gDls8_1(.din(w_dff_B_8SKuRgD08_1),.dout(w_dff_B_WQO8gDls8_1),.clk(gclk));
	jdff dff_B_LGoYdaZg6_1(.din(w_dff_B_WQO8gDls8_1),.dout(w_dff_B_LGoYdaZg6_1),.clk(gclk));
	jdff dff_B_AbSDOs336_1(.din(w_dff_B_LGoYdaZg6_1),.dout(w_dff_B_AbSDOs336_1),.clk(gclk));
	jdff dff_B_osv36UEq6_1(.din(w_dff_B_AbSDOs336_1),.dout(w_dff_B_osv36UEq6_1),.clk(gclk));
	jdff dff_B_4SZA163P8_1(.din(w_dff_B_osv36UEq6_1),.dout(w_dff_B_4SZA163P8_1),.clk(gclk));
	jdff dff_B_UesKWUS14_1(.din(w_dff_B_4SZA163P8_1),.dout(w_dff_B_UesKWUS14_1),.clk(gclk));
	jdff dff_B_gNPo2dzH8_1(.din(w_dff_B_UesKWUS14_1),.dout(w_dff_B_gNPo2dzH8_1),.clk(gclk));
	jdff dff_B_ODqNautq3_1(.din(w_dff_B_gNPo2dzH8_1),.dout(w_dff_B_ODqNautq3_1),.clk(gclk));
	jdff dff_B_jgcXi6pZ7_1(.din(w_dff_B_ODqNautq3_1),.dout(w_dff_B_jgcXi6pZ7_1),.clk(gclk));
	jdff dff_B_IXx4TcSe3_1(.din(w_dff_B_jgcXi6pZ7_1),.dout(w_dff_B_IXx4TcSe3_1),.clk(gclk));
	jdff dff_B_Ur0U9lGf8_1(.din(w_dff_B_IXx4TcSe3_1),.dout(w_dff_B_Ur0U9lGf8_1),.clk(gclk));
	jdff dff_B_L0XYUffd4_1(.din(w_dff_B_Ur0U9lGf8_1),.dout(w_dff_B_L0XYUffd4_1),.clk(gclk));
	jdff dff_B_Tlk9GDzm3_1(.din(w_dff_B_L0XYUffd4_1),.dout(w_dff_B_Tlk9GDzm3_1),.clk(gclk));
	jdff dff_B_cJvfzVON1_1(.din(w_dff_B_Tlk9GDzm3_1),.dout(w_dff_B_cJvfzVON1_1),.clk(gclk));
	jdff dff_B_k4Z7XCDJ6_1(.din(w_dff_B_cJvfzVON1_1),.dout(w_dff_B_k4Z7XCDJ6_1),.clk(gclk));
	jdff dff_B_vv4ZDUyh9_1(.din(w_dff_B_k4Z7XCDJ6_1),.dout(w_dff_B_vv4ZDUyh9_1),.clk(gclk));
	jdff dff_B_8iqiTTzx3_1(.din(w_dff_B_vv4ZDUyh9_1),.dout(w_dff_B_8iqiTTzx3_1),.clk(gclk));
	jdff dff_B_QP7WfLZS6_1(.din(w_dff_B_8iqiTTzx3_1),.dout(w_dff_B_QP7WfLZS6_1),.clk(gclk));
	jdff dff_B_3IwECteJ0_1(.din(w_dff_B_QP7WfLZS6_1),.dout(w_dff_B_3IwECteJ0_1),.clk(gclk));
	jdff dff_B_ZxEmBrr27_1(.din(w_dff_B_3IwECteJ0_1),.dout(w_dff_B_ZxEmBrr27_1),.clk(gclk));
	jdff dff_B_YaaUE8zO1_1(.din(w_dff_B_ZxEmBrr27_1),.dout(w_dff_B_YaaUE8zO1_1),.clk(gclk));
	jdff dff_B_hYH7VbdA0_1(.din(w_dff_B_YaaUE8zO1_1),.dout(w_dff_B_hYH7VbdA0_1),.clk(gclk));
	jdff dff_B_5x7Mp2Lx7_1(.din(w_dff_B_hYH7VbdA0_1),.dout(w_dff_B_5x7Mp2Lx7_1),.clk(gclk));
	jdff dff_B_H83HnVeM9_1(.din(w_dff_B_5x7Mp2Lx7_1),.dout(w_dff_B_H83HnVeM9_1),.clk(gclk));
	jdff dff_B_VDg9BtRN8_1(.din(w_dff_B_H83HnVeM9_1),.dout(w_dff_B_VDg9BtRN8_1),.clk(gclk));
	jdff dff_B_5D26V9wt3_1(.din(w_dff_B_VDg9BtRN8_1),.dout(w_dff_B_5D26V9wt3_1),.clk(gclk));
	jdff dff_B_r9KLOEtj1_1(.din(w_dff_B_5D26V9wt3_1),.dout(w_dff_B_r9KLOEtj1_1),.clk(gclk));
	jdff dff_B_94rmknWS0_1(.din(w_dff_B_r9KLOEtj1_1),.dout(w_dff_B_94rmknWS0_1),.clk(gclk));
	jdff dff_B_LF4wsQji1_1(.din(w_dff_B_94rmknWS0_1),.dout(w_dff_B_LF4wsQji1_1),.clk(gclk));
	jdff dff_B_5IofoIbI0_1(.din(w_dff_B_LF4wsQji1_1),.dout(w_dff_B_5IofoIbI0_1),.clk(gclk));
	jdff dff_B_wwyyc6zB6_1(.din(w_dff_B_5IofoIbI0_1),.dout(w_dff_B_wwyyc6zB6_1),.clk(gclk));
	jdff dff_B_5sj9XZwc7_1(.din(w_dff_B_wwyyc6zB6_1),.dout(w_dff_B_5sj9XZwc7_1),.clk(gclk));
	jdff dff_B_yOAEe7IH2_1(.din(w_dff_B_5sj9XZwc7_1),.dout(w_dff_B_yOAEe7IH2_1),.clk(gclk));
	jdff dff_B_IHkCUzU34_1(.din(w_dff_B_yOAEe7IH2_1),.dout(w_dff_B_IHkCUzU34_1),.clk(gclk));
	jdff dff_B_XaAe5UmA1_1(.din(w_dff_B_IHkCUzU34_1),.dout(w_dff_B_XaAe5UmA1_1),.clk(gclk));
	jdff dff_B_cBESAYhG1_1(.din(w_dff_B_XaAe5UmA1_1),.dout(w_dff_B_cBESAYhG1_1),.clk(gclk));
	jdff dff_B_JceMSJ8I2_1(.din(w_dff_B_cBESAYhG1_1),.dout(w_dff_B_JceMSJ8I2_1),.clk(gclk));
	jdff dff_B_1zQC9HOu0_1(.din(w_dff_B_JceMSJ8I2_1),.dout(w_dff_B_1zQC9HOu0_1),.clk(gclk));
	jdff dff_B_gv1fmmBW4_1(.din(w_dff_B_1zQC9HOu0_1),.dout(w_dff_B_gv1fmmBW4_1),.clk(gclk));
	jdff dff_B_5IyfkmIV0_1(.din(w_dff_B_gv1fmmBW4_1),.dout(w_dff_B_5IyfkmIV0_1),.clk(gclk));
	jdff dff_B_hDpjD3FY8_1(.din(w_dff_B_5IyfkmIV0_1),.dout(w_dff_B_hDpjD3FY8_1),.clk(gclk));
	jdff dff_B_taonE3Hk0_1(.din(w_dff_B_hDpjD3FY8_1),.dout(w_dff_B_taonE3Hk0_1),.clk(gclk));
	jdff dff_B_P747L8WS5_1(.din(w_dff_B_taonE3Hk0_1),.dout(w_dff_B_P747L8WS5_1),.clk(gclk));
	jdff dff_B_LciAk2zr4_1(.din(w_dff_B_P747L8WS5_1),.dout(w_dff_B_LciAk2zr4_1),.clk(gclk));
	jdff dff_B_tMB6SiXu4_1(.din(w_dff_B_LciAk2zr4_1),.dout(w_dff_B_tMB6SiXu4_1),.clk(gclk));
	jdff dff_B_Qf773v530_1(.din(w_dff_B_tMB6SiXu4_1),.dout(w_dff_B_Qf773v530_1),.clk(gclk));
	jdff dff_B_HtvzNgK15_1(.din(w_dff_B_Qf773v530_1),.dout(w_dff_B_HtvzNgK15_1),.clk(gclk));
	jdff dff_B_uIqRUHnO5_1(.din(w_dff_B_HtvzNgK15_1),.dout(w_dff_B_uIqRUHnO5_1),.clk(gclk));
	jdff dff_B_uTzEIOu43_1(.din(w_dff_B_uIqRUHnO5_1),.dout(w_dff_B_uTzEIOu43_1),.clk(gclk));
	jdff dff_B_zpmvfynv2_1(.din(w_dff_B_uTzEIOu43_1),.dout(w_dff_B_zpmvfynv2_1),.clk(gclk));
	jdff dff_B_QSY34u1X5_1(.din(w_dff_B_zpmvfynv2_1),.dout(w_dff_B_QSY34u1X5_1),.clk(gclk));
	jdff dff_B_JGl9DQes3_1(.din(w_dff_B_QSY34u1X5_1),.dout(w_dff_B_JGl9DQes3_1),.clk(gclk));
	jdff dff_B_uQaNhLDe6_1(.din(w_dff_B_JGl9DQes3_1),.dout(w_dff_B_uQaNhLDe6_1),.clk(gclk));
	jdff dff_B_YISJmDUl2_1(.din(w_dff_B_uQaNhLDe6_1),.dout(w_dff_B_YISJmDUl2_1),.clk(gclk));
	jdff dff_B_qZMmcBxe9_1(.din(w_dff_B_YISJmDUl2_1),.dout(w_dff_B_qZMmcBxe9_1),.clk(gclk));
	jdff dff_B_xgwmgfx24_1(.din(w_dff_B_qZMmcBxe9_1),.dout(w_dff_B_xgwmgfx24_1),.clk(gclk));
	jdff dff_B_ymgcPYnU6_1(.din(w_dff_B_xgwmgfx24_1),.dout(w_dff_B_ymgcPYnU6_1),.clk(gclk));
	jdff dff_B_Ne01avRW2_1(.din(w_dff_B_ymgcPYnU6_1),.dout(w_dff_B_Ne01avRW2_1),.clk(gclk));
	jdff dff_B_oH1sQqBu3_1(.din(w_dff_B_Ne01avRW2_1),.dout(w_dff_B_oH1sQqBu3_1),.clk(gclk));
	jdff dff_B_ImXwsVgn7_1(.din(w_dff_B_oH1sQqBu3_1),.dout(w_dff_B_ImXwsVgn7_1),.clk(gclk));
	jdff dff_B_5QWsOaar3_1(.din(w_dff_B_ImXwsVgn7_1),.dout(w_dff_B_5QWsOaar3_1),.clk(gclk));
	jdff dff_B_8zszqGh32_1(.din(w_dff_B_5QWsOaar3_1),.dout(w_dff_B_8zszqGh32_1),.clk(gclk));
	jdff dff_B_d0QARxKa6_1(.din(w_dff_B_8zszqGh32_1),.dout(w_dff_B_d0QARxKa6_1),.clk(gclk));
	jdff dff_B_ZOjvBBCA8_1(.din(w_dff_B_d0QARxKa6_1),.dout(w_dff_B_ZOjvBBCA8_1),.clk(gclk));
	jdff dff_B_tAY6tdAr0_1(.din(w_dff_B_ZOjvBBCA8_1),.dout(w_dff_B_tAY6tdAr0_1),.clk(gclk));
	jdff dff_B_ss4fYgPG1_1(.din(w_dff_B_tAY6tdAr0_1),.dout(w_dff_B_ss4fYgPG1_1),.clk(gclk));
	jdff dff_B_PJbZVXZ39_1(.din(w_dff_B_ss4fYgPG1_1),.dout(w_dff_B_PJbZVXZ39_1),.clk(gclk));
	jdff dff_B_UaA2q3QW0_1(.din(w_dff_B_PJbZVXZ39_1),.dout(w_dff_B_UaA2q3QW0_1),.clk(gclk));
	jdff dff_B_zXuXbAg94_1(.din(w_dff_B_UaA2q3QW0_1),.dout(w_dff_B_zXuXbAg94_1),.clk(gclk));
	jdff dff_B_kg0aVgPW1_1(.din(w_dff_B_zXuXbAg94_1),.dout(w_dff_B_kg0aVgPW1_1),.clk(gclk));
	jdff dff_B_qXDo8E5j9_1(.din(w_dff_B_kg0aVgPW1_1),.dout(w_dff_B_qXDo8E5j9_1),.clk(gclk));
	jdff dff_B_FvOkDus66_1(.din(w_dff_B_qXDo8E5j9_1),.dout(w_dff_B_FvOkDus66_1),.clk(gclk));
	jdff dff_B_ORaioyxN3_1(.din(w_dff_B_FvOkDus66_1),.dout(w_dff_B_ORaioyxN3_1),.clk(gclk));
	jdff dff_B_ENSVAwRI7_1(.din(w_dff_B_ORaioyxN3_1),.dout(w_dff_B_ENSVAwRI7_1),.clk(gclk));
	jdff dff_B_ZjnuHFbu0_1(.din(w_dff_B_ENSVAwRI7_1),.dout(w_dff_B_ZjnuHFbu0_1),.clk(gclk));
	jdff dff_B_2rSl9HV12_1(.din(w_dff_B_ZjnuHFbu0_1),.dout(w_dff_B_2rSl9HV12_1),.clk(gclk));
	jdff dff_B_yqZitFZj4_1(.din(w_dff_B_2rSl9HV12_1),.dout(w_dff_B_yqZitFZj4_1),.clk(gclk));
	jdff dff_B_ANVA01PR5_1(.din(w_dff_B_yqZitFZj4_1),.dout(w_dff_B_ANVA01PR5_1),.clk(gclk));
	jdff dff_B_gvgNoTLP7_1(.din(w_dff_B_ANVA01PR5_1),.dout(w_dff_B_gvgNoTLP7_1),.clk(gclk));
	jdff dff_B_nwX3XGbn2_1(.din(w_dff_B_gvgNoTLP7_1),.dout(w_dff_B_nwX3XGbn2_1),.clk(gclk));
	jdff dff_B_JdwvomK95_1(.din(w_dff_B_nwX3XGbn2_1),.dout(w_dff_B_JdwvomK95_1),.clk(gclk));
	jdff dff_B_D1eNItdK8_1(.din(w_dff_B_JdwvomK95_1),.dout(w_dff_B_D1eNItdK8_1),.clk(gclk));
	jdff dff_B_BMacVM8n4_1(.din(w_dff_B_D1eNItdK8_1),.dout(w_dff_B_BMacVM8n4_1),.clk(gclk));
	jdff dff_B_8deQ3RaC2_0(.din(n1033),.dout(w_dff_B_8deQ3RaC2_0),.clk(gclk));
	jdff dff_B_LZL8vLaM7_0(.din(w_dff_B_8deQ3RaC2_0),.dout(w_dff_B_LZL8vLaM7_0),.clk(gclk));
	jdff dff_B_zCoLkU1W2_0(.din(w_dff_B_LZL8vLaM7_0),.dout(w_dff_B_zCoLkU1W2_0),.clk(gclk));
	jdff dff_B_Sjo7tciE3_0(.din(w_dff_B_zCoLkU1W2_0),.dout(w_dff_B_Sjo7tciE3_0),.clk(gclk));
	jdff dff_B_1TG6dtgk4_0(.din(w_dff_B_Sjo7tciE3_0),.dout(w_dff_B_1TG6dtgk4_0),.clk(gclk));
	jdff dff_B_sDs86Ikx2_0(.din(w_dff_B_1TG6dtgk4_0),.dout(w_dff_B_sDs86Ikx2_0),.clk(gclk));
	jdff dff_B_z6PUWR8z2_0(.din(w_dff_B_sDs86Ikx2_0),.dout(w_dff_B_z6PUWR8z2_0),.clk(gclk));
	jdff dff_B_slbc8sEX2_0(.din(w_dff_B_z6PUWR8z2_0),.dout(w_dff_B_slbc8sEX2_0),.clk(gclk));
	jdff dff_B_0abywTc20_0(.din(w_dff_B_slbc8sEX2_0),.dout(w_dff_B_0abywTc20_0),.clk(gclk));
	jdff dff_B_Nxc9yxPb6_0(.din(w_dff_B_0abywTc20_0),.dout(w_dff_B_Nxc9yxPb6_0),.clk(gclk));
	jdff dff_B_Tt9BHrTK8_0(.din(w_dff_B_Nxc9yxPb6_0),.dout(w_dff_B_Tt9BHrTK8_0),.clk(gclk));
	jdff dff_B_3UweyeU27_0(.din(w_dff_B_Tt9BHrTK8_0),.dout(w_dff_B_3UweyeU27_0),.clk(gclk));
	jdff dff_B_oA47j4YF9_0(.din(w_dff_B_3UweyeU27_0),.dout(w_dff_B_oA47j4YF9_0),.clk(gclk));
	jdff dff_B_xvD4s9IZ5_0(.din(w_dff_B_oA47j4YF9_0),.dout(w_dff_B_xvD4s9IZ5_0),.clk(gclk));
	jdff dff_B_GtepwspG4_0(.din(w_dff_B_xvD4s9IZ5_0),.dout(w_dff_B_GtepwspG4_0),.clk(gclk));
	jdff dff_B_wtsmixzP9_0(.din(w_dff_B_GtepwspG4_0),.dout(w_dff_B_wtsmixzP9_0),.clk(gclk));
	jdff dff_B_xqHyY5m65_0(.din(w_dff_B_wtsmixzP9_0),.dout(w_dff_B_xqHyY5m65_0),.clk(gclk));
	jdff dff_B_CHnjgpIv6_0(.din(w_dff_B_xqHyY5m65_0),.dout(w_dff_B_CHnjgpIv6_0),.clk(gclk));
	jdff dff_B_h0Bglps86_0(.din(w_dff_B_CHnjgpIv6_0),.dout(w_dff_B_h0Bglps86_0),.clk(gclk));
	jdff dff_B_DSK2wJdV5_0(.din(w_dff_B_h0Bglps86_0),.dout(w_dff_B_DSK2wJdV5_0),.clk(gclk));
	jdff dff_B_4DyduRFv9_0(.din(w_dff_B_DSK2wJdV5_0),.dout(w_dff_B_4DyduRFv9_0),.clk(gclk));
	jdff dff_B_5ZiI9uBl4_0(.din(w_dff_B_4DyduRFv9_0),.dout(w_dff_B_5ZiI9uBl4_0),.clk(gclk));
	jdff dff_B_2QQkHLUC3_0(.din(w_dff_B_5ZiI9uBl4_0),.dout(w_dff_B_2QQkHLUC3_0),.clk(gclk));
	jdff dff_B_kVDEMbO49_0(.din(w_dff_B_2QQkHLUC3_0),.dout(w_dff_B_kVDEMbO49_0),.clk(gclk));
	jdff dff_B_pNVNweeH6_0(.din(w_dff_B_kVDEMbO49_0),.dout(w_dff_B_pNVNweeH6_0),.clk(gclk));
	jdff dff_B_crShAWPu0_0(.din(w_dff_B_pNVNweeH6_0),.dout(w_dff_B_crShAWPu0_0),.clk(gclk));
	jdff dff_B_AFVvm6CW1_0(.din(w_dff_B_crShAWPu0_0),.dout(w_dff_B_AFVvm6CW1_0),.clk(gclk));
	jdff dff_B_NuyCH00F5_0(.din(w_dff_B_AFVvm6CW1_0),.dout(w_dff_B_NuyCH00F5_0),.clk(gclk));
	jdff dff_B_Aj2o48NQ3_0(.din(w_dff_B_NuyCH00F5_0),.dout(w_dff_B_Aj2o48NQ3_0),.clk(gclk));
	jdff dff_B_16tKTqVr7_0(.din(w_dff_B_Aj2o48NQ3_0),.dout(w_dff_B_16tKTqVr7_0),.clk(gclk));
	jdff dff_B_oB0TbDs02_0(.din(w_dff_B_16tKTqVr7_0),.dout(w_dff_B_oB0TbDs02_0),.clk(gclk));
	jdff dff_B_PlGcQ7vB6_0(.din(w_dff_B_oB0TbDs02_0),.dout(w_dff_B_PlGcQ7vB6_0),.clk(gclk));
	jdff dff_B_aNbozymt3_0(.din(w_dff_B_PlGcQ7vB6_0),.dout(w_dff_B_aNbozymt3_0),.clk(gclk));
	jdff dff_B_vPiBtOGQ3_0(.din(w_dff_B_aNbozymt3_0),.dout(w_dff_B_vPiBtOGQ3_0),.clk(gclk));
	jdff dff_B_kLl3hZl09_0(.din(w_dff_B_vPiBtOGQ3_0),.dout(w_dff_B_kLl3hZl09_0),.clk(gclk));
	jdff dff_B_3mgr8RtU0_0(.din(w_dff_B_kLl3hZl09_0),.dout(w_dff_B_3mgr8RtU0_0),.clk(gclk));
	jdff dff_B_iva8plW76_0(.din(w_dff_B_3mgr8RtU0_0),.dout(w_dff_B_iva8plW76_0),.clk(gclk));
	jdff dff_B_KC5tcFuK8_0(.din(w_dff_B_iva8plW76_0),.dout(w_dff_B_KC5tcFuK8_0),.clk(gclk));
	jdff dff_B_7jJfqrHH6_0(.din(w_dff_B_KC5tcFuK8_0),.dout(w_dff_B_7jJfqrHH6_0),.clk(gclk));
	jdff dff_B_fHA6wVgn7_0(.din(w_dff_B_7jJfqrHH6_0),.dout(w_dff_B_fHA6wVgn7_0),.clk(gclk));
	jdff dff_B_yj70ytnF2_0(.din(w_dff_B_fHA6wVgn7_0),.dout(w_dff_B_yj70ytnF2_0),.clk(gclk));
	jdff dff_B_rVhPHQmC7_0(.din(w_dff_B_yj70ytnF2_0),.dout(w_dff_B_rVhPHQmC7_0),.clk(gclk));
	jdff dff_B_Kh6NGusd7_0(.din(w_dff_B_rVhPHQmC7_0),.dout(w_dff_B_Kh6NGusd7_0),.clk(gclk));
	jdff dff_B_7kj2tfp01_0(.din(w_dff_B_Kh6NGusd7_0),.dout(w_dff_B_7kj2tfp01_0),.clk(gclk));
	jdff dff_B_AyE07pT04_0(.din(w_dff_B_7kj2tfp01_0),.dout(w_dff_B_AyE07pT04_0),.clk(gclk));
	jdff dff_B_dvzjfVSt7_0(.din(w_dff_B_AyE07pT04_0),.dout(w_dff_B_dvzjfVSt7_0),.clk(gclk));
	jdff dff_B_CDxmYxKr7_0(.din(w_dff_B_dvzjfVSt7_0),.dout(w_dff_B_CDxmYxKr7_0),.clk(gclk));
	jdff dff_B_XS4DU9tw4_0(.din(w_dff_B_CDxmYxKr7_0),.dout(w_dff_B_XS4DU9tw4_0),.clk(gclk));
	jdff dff_B_2bF4EF9Z5_0(.din(w_dff_B_XS4DU9tw4_0),.dout(w_dff_B_2bF4EF9Z5_0),.clk(gclk));
	jdff dff_B_a5K1c3Bo8_0(.din(w_dff_B_2bF4EF9Z5_0),.dout(w_dff_B_a5K1c3Bo8_0),.clk(gclk));
	jdff dff_B_53qxiWqd2_0(.din(w_dff_B_a5K1c3Bo8_0),.dout(w_dff_B_53qxiWqd2_0),.clk(gclk));
	jdff dff_B_U8Cra25v2_0(.din(w_dff_B_53qxiWqd2_0),.dout(w_dff_B_U8Cra25v2_0),.clk(gclk));
	jdff dff_B_goAZPxvf2_0(.din(w_dff_B_U8Cra25v2_0),.dout(w_dff_B_goAZPxvf2_0),.clk(gclk));
	jdff dff_B_9jiy1SYX1_0(.din(w_dff_B_goAZPxvf2_0),.dout(w_dff_B_9jiy1SYX1_0),.clk(gclk));
	jdff dff_B_HkdNSkfs4_0(.din(w_dff_B_9jiy1SYX1_0),.dout(w_dff_B_HkdNSkfs4_0),.clk(gclk));
	jdff dff_B_HZ9we5PL3_0(.din(w_dff_B_HkdNSkfs4_0),.dout(w_dff_B_HZ9we5PL3_0),.clk(gclk));
	jdff dff_B_fRQ8TtFq2_0(.din(w_dff_B_HZ9we5PL3_0),.dout(w_dff_B_fRQ8TtFq2_0),.clk(gclk));
	jdff dff_B_CSKFWIas1_0(.din(w_dff_B_fRQ8TtFq2_0),.dout(w_dff_B_CSKFWIas1_0),.clk(gclk));
	jdff dff_B_hbmTbEWi8_0(.din(w_dff_B_CSKFWIas1_0),.dout(w_dff_B_hbmTbEWi8_0),.clk(gclk));
	jdff dff_B_XeCv7cN38_0(.din(w_dff_B_hbmTbEWi8_0),.dout(w_dff_B_XeCv7cN38_0),.clk(gclk));
	jdff dff_B_O85L9Tk05_0(.din(w_dff_B_XeCv7cN38_0),.dout(w_dff_B_O85L9Tk05_0),.clk(gclk));
	jdff dff_B_PUUBZXtq3_0(.din(w_dff_B_O85L9Tk05_0),.dout(w_dff_B_PUUBZXtq3_0),.clk(gclk));
	jdff dff_B_Z6CSjm9I1_0(.din(w_dff_B_PUUBZXtq3_0),.dout(w_dff_B_Z6CSjm9I1_0),.clk(gclk));
	jdff dff_B_KpPV1p3s6_0(.din(w_dff_B_Z6CSjm9I1_0),.dout(w_dff_B_KpPV1p3s6_0),.clk(gclk));
	jdff dff_B_0XYGvi6T6_0(.din(w_dff_B_KpPV1p3s6_0),.dout(w_dff_B_0XYGvi6T6_0),.clk(gclk));
	jdff dff_B_zecfbCZG9_0(.din(w_dff_B_0XYGvi6T6_0),.dout(w_dff_B_zecfbCZG9_0),.clk(gclk));
	jdff dff_B_MSyEWdwW9_0(.din(w_dff_B_zecfbCZG9_0),.dout(w_dff_B_MSyEWdwW9_0),.clk(gclk));
	jdff dff_B_zFxI68wS8_0(.din(w_dff_B_MSyEWdwW9_0),.dout(w_dff_B_zFxI68wS8_0),.clk(gclk));
	jdff dff_B_xayqS21i1_0(.din(w_dff_B_zFxI68wS8_0),.dout(w_dff_B_xayqS21i1_0),.clk(gclk));
	jdff dff_B_vtoGmsN28_0(.din(w_dff_B_xayqS21i1_0),.dout(w_dff_B_vtoGmsN28_0),.clk(gclk));
	jdff dff_B_g513HMU55_0(.din(w_dff_B_vtoGmsN28_0),.dout(w_dff_B_g513HMU55_0),.clk(gclk));
	jdff dff_B_3ZnT0QOE9_0(.din(w_dff_B_g513HMU55_0),.dout(w_dff_B_3ZnT0QOE9_0),.clk(gclk));
	jdff dff_B_e61vckDh0_0(.din(w_dff_B_3ZnT0QOE9_0),.dout(w_dff_B_e61vckDh0_0),.clk(gclk));
	jdff dff_B_aiVXdiAC4_0(.din(w_dff_B_e61vckDh0_0),.dout(w_dff_B_aiVXdiAC4_0),.clk(gclk));
	jdff dff_B_7hFEtFMA2_0(.din(w_dff_B_aiVXdiAC4_0),.dout(w_dff_B_7hFEtFMA2_0),.clk(gclk));
	jdff dff_B_Ym1v7XJ56_0(.din(w_dff_B_7hFEtFMA2_0),.dout(w_dff_B_Ym1v7XJ56_0),.clk(gclk));
	jdff dff_B_wySjj1zN5_0(.din(w_dff_B_Ym1v7XJ56_0),.dout(w_dff_B_wySjj1zN5_0),.clk(gclk));
	jdff dff_B_Hdu3tnUH8_0(.din(w_dff_B_wySjj1zN5_0),.dout(w_dff_B_Hdu3tnUH8_0),.clk(gclk));
	jdff dff_B_H3Xc0WrE1_0(.din(w_dff_B_Hdu3tnUH8_0),.dout(w_dff_B_H3Xc0WrE1_0),.clk(gclk));
	jdff dff_B_KLDaTWHJ2_0(.din(w_dff_B_H3Xc0WrE1_0),.dout(w_dff_B_KLDaTWHJ2_0),.clk(gclk));
	jdff dff_B_YEwlDs3x4_0(.din(w_dff_B_KLDaTWHJ2_0),.dout(w_dff_B_YEwlDs3x4_0),.clk(gclk));
	jdff dff_B_nmLBtDhF4_0(.din(w_dff_B_YEwlDs3x4_0),.dout(w_dff_B_nmLBtDhF4_0),.clk(gclk));
	jdff dff_B_M91nXk6g2_0(.din(w_dff_B_nmLBtDhF4_0),.dout(w_dff_B_M91nXk6g2_0),.clk(gclk));
	jdff dff_B_QiLGjchY4_0(.din(w_dff_B_M91nXk6g2_0),.dout(w_dff_B_QiLGjchY4_0),.clk(gclk));
	jdff dff_B_c15dFlmW2_0(.din(w_dff_B_QiLGjchY4_0),.dout(w_dff_B_c15dFlmW2_0),.clk(gclk));
	jdff dff_B_Re2vektU1_0(.din(w_dff_B_c15dFlmW2_0),.dout(w_dff_B_Re2vektU1_0),.clk(gclk));
	jdff dff_B_taHjV3hZ3_0(.din(w_dff_B_Re2vektU1_0),.dout(w_dff_B_taHjV3hZ3_0),.clk(gclk));
	jdff dff_B_ZjJR6ow80_0(.din(w_dff_B_taHjV3hZ3_0),.dout(w_dff_B_ZjJR6ow80_0),.clk(gclk));
	jdff dff_B_wkcVbRyr8_0(.din(w_dff_B_ZjJR6ow80_0),.dout(w_dff_B_wkcVbRyr8_0),.clk(gclk));
	jdff dff_B_cIvUoP7m0_0(.din(w_dff_B_wkcVbRyr8_0),.dout(w_dff_B_cIvUoP7m0_0),.clk(gclk));
	jdff dff_B_w7N7Xmkr3_0(.din(w_dff_B_cIvUoP7m0_0),.dout(w_dff_B_w7N7Xmkr3_0),.clk(gclk));
	jdff dff_B_NlewqK2G4_0(.din(w_dff_B_w7N7Xmkr3_0),.dout(w_dff_B_NlewqK2G4_0),.clk(gclk));
	jdff dff_B_0bBG0e9p3_0(.din(w_dff_B_NlewqK2G4_0),.dout(w_dff_B_0bBG0e9p3_0),.clk(gclk));
	jdff dff_B_FgaDW4t81_0(.din(w_dff_B_0bBG0e9p3_0),.dout(w_dff_B_FgaDW4t81_0),.clk(gclk));
	jdff dff_B_spk9uJHE8_0(.din(w_dff_B_FgaDW4t81_0),.dout(w_dff_B_spk9uJHE8_0),.clk(gclk));
	jdff dff_B_hxXzLpOP1_0(.din(w_dff_B_spk9uJHE8_0),.dout(w_dff_B_hxXzLpOP1_0),.clk(gclk));
	jdff dff_B_cIoKiF850_0(.din(w_dff_B_hxXzLpOP1_0),.dout(w_dff_B_cIoKiF850_0),.clk(gclk));
	jdff dff_B_l2or20CR9_0(.din(w_dff_B_cIoKiF850_0),.dout(w_dff_B_l2or20CR9_0),.clk(gclk));
	jdff dff_B_zvXq4FAs6_0(.din(w_dff_B_l2or20CR9_0),.dout(w_dff_B_zvXq4FAs6_0),.clk(gclk));
	jdff dff_B_v6DhjobE1_0(.din(w_dff_B_zvXq4FAs6_0),.dout(w_dff_B_v6DhjobE1_0),.clk(gclk));
	jdff dff_B_6QK2jsIT8_0(.din(w_dff_B_v6DhjobE1_0),.dout(w_dff_B_6QK2jsIT8_0),.clk(gclk));
	jdff dff_B_Tt7TPj6N2_0(.din(w_dff_B_6QK2jsIT8_0),.dout(w_dff_B_Tt7TPj6N2_0),.clk(gclk));
	jdff dff_B_a35uhzbZ9_0(.din(w_dff_B_Tt7TPj6N2_0),.dout(w_dff_B_a35uhzbZ9_0),.clk(gclk));
	jdff dff_B_4c2yPfRT6_0(.din(w_dff_B_a35uhzbZ9_0),.dout(w_dff_B_4c2yPfRT6_0),.clk(gclk));
	jdff dff_B_G9smq10s2_0(.din(w_dff_B_4c2yPfRT6_0),.dout(w_dff_B_G9smq10s2_0),.clk(gclk));
	jdff dff_B_cJVNtqKO5_0(.din(w_dff_B_G9smq10s2_0),.dout(w_dff_B_cJVNtqKO5_0),.clk(gclk));
	jdff dff_B_bJrEKCoO4_0(.din(w_dff_B_cJVNtqKO5_0),.dout(w_dff_B_bJrEKCoO4_0),.clk(gclk));
	jdff dff_B_ISqqPwDn9_0(.din(w_dff_B_bJrEKCoO4_0),.dout(w_dff_B_ISqqPwDn9_0),.clk(gclk));
	jdff dff_B_sNp6ShSz7_1(.din(n1026),.dout(w_dff_B_sNp6ShSz7_1),.clk(gclk));
	jdff dff_B_kJFprg0r5_1(.din(w_dff_B_sNp6ShSz7_1),.dout(w_dff_B_kJFprg0r5_1),.clk(gclk));
	jdff dff_B_dINkKPxx1_1(.din(w_dff_B_kJFprg0r5_1),.dout(w_dff_B_dINkKPxx1_1),.clk(gclk));
	jdff dff_B_W2v9cfAu0_1(.din(w_dff_B_dINkKPxx1_1),.dout(w_dff_B_W2v9cfAu0_1),.clk(gclk));
	jdff dff_B_DUGQt5qn9_1(.din(w_dff_B_W2v9cfAu0_1),.dout(w_dff_B_DUGQt5qn9_1),.clk(gclk));
	jdff dff_B_73CLID8z0_1(.din(w_dff_B_DUGQt5qn9_1),.dout(w_dff_B_73CLID8z0_1),.clk(gclk));
	jdff dff_B_oRCSPhpP4_1(.din(w_dff_B_73CLID8z0_1),.dout(w_dff_B_oRCSPhpP4_1),.clk(gclk));
	jdff dff_B_ZlMj3kR61_1(.din(w_dff_B_oRCSPhpP4_1),.dout(w_dff_B_ZlMj3kR61_1),.clk(gclk));
	jdff dff_B_KX2LgwsS9_1(.din(w_dff_B_ZlMj3kR61_1),.dout(w_dff_B_KX2LgwsS9_1),.clk(gclk));
	jdff dff_B_vuUqtOWm6_1(.din(w_dff_B_KX2LgwsS9_1),.dout(w_dff_B_vuUqtOWm6_1),.clk(gclk));
	jdff dff_B_Auwu0XXj6_1(.din(w_dff_B_vuUqtOWm6_1),.dout(w_dff_B_Auwu0XXj6_1),.clk(gclk));
	jdff dff_B_KB4ZfdLj2_1(.din(w_dff_B_Auwu0XXj6_1),.dout(w_dff_B_KB4ZfdLj2_1),.clk(gclk));
	jdff dff_B_HngxO0Uj0_1(.din(w_dff_B_KB4ZfdLj2_1),.dout(w_dff_B_HngxO0Uj0_1),.clk(gclk));
	jdff dff_B_2rAo27ek3_1(.din(w_dff_B_HngxO0Uj0_1),.dout(w_dff_B_2rAo27ek3_1),.clk(gclk));
	jdff dff_B_1yuMyIff2_1(.din(w_dff_B_2rAo27ek3_1),.dout(w_dff_B_1yuMyIff2_1),.clk(gclk));
	jdff dff_B_bwOPwuYv2_1(.din(w_dff_B_1yuMyIff2_1),.dout(w_dff_B_bwOPwuYv2_1),.clk(gclk));
	jdff dff_B_MTk4h14h7_1(.din(w_dff_B_bwOPwuYv2_1),.dout(w_dff_B_MTk4h14h7_1),.clk(gclk));
	jdff dff_B_d7WeVBrS5_1(.din(w_dff_B_MTk4h14h7_1),.dout(w_dff_B_d7WeVBrS5_1),.clk(gclk));
	jdff dff_B_FrWhF4Cz9_1(.din(w_dff_B_d7WeVBrS5_1),.dout(w_dff_B_FrWhF4Cz9_1),.clk(gclk));
	jdff dff_B_hJUC7WUN2_1(.din(w_dff_B_FrWhF4Cz9_1),.dout(w_dff_B_hJUC7WUN2_1),.clk(gclk));
	jdff dff_B_CxKcba1o0_1(.din(w_dff_B_hJUC7WUN2_1),.dout(w_dff_B_CxKcba1o0_1),.clk(gclk));
	jdff dff_B_6vUiK6130_1(.din(w_dff_B_CxKcba1o0_1),.dout(w_dff_B_6vUiK6130_1),.clk(gclk));
	jdff dff_B_mjDMx4ul9_1(.din(w_dff_B_6vUiK6130_1),.dout(w_dff_B_mjDMx4ul9_1),.clk(gclk));
	jdff dff_B_tYKbNTyW2_1(.din(w_dff_B_mjDMx4ul9_1),.dout(w_dff_B_tYKbNTyW2_1),.clk(gclk));
	jdff dff_B_A3wnPson6_1(.din(w_dff_B_tYKbNTyW2_1),.dout(w_dff_B_A3wnPson6_1),.clk(gclk));
	jdff dff_B_j9Jg9zDH3_1(.din(w_dff_B_A3wnPson6_1),.dout(w_dff_B_j9Jg9zDH3_1),.clk(gclk));
	jdff dff_B_QYaEuE2X5_1(.din(w_dff_B_j9Jg9zDH3_1),.dout(w_dff_B_QYaEuE2X5_1),.clk(gclk));
	jdff dff_B_tJoPPfBW7_1(.din(w_dff_B_QYaEuE2X5_1),.dout(w_dff_B_tJoPPfBW7_1),.clk(gclk));
	jdff dff_B_BcfQLpAq2_1(.din(w_dff_B_tJoPPfBW7_1),.dout(w_dff_B_BcfQLpAq2_1),.clk(gclk));
	jdff dff_B_fGdEvZyL9_1(.din(w_dff_B_BcfQLpAq2_1),.dout(w_dff_B_fGdEvZyL9_1),.clk(gclk));
	jdff dff_B_lt2uSuFn2_1(.din(w_dff_B_fGdEvZyL9_1),.dout(w_dff_B_lt2uSuFn2_1),.clk(gclk));
	jdff dff_B_eOwKKlvL6_1(.din(w_dff_B_lt2uSuFn2_1),.dout(w_dff_B_eOwKKlvL6_1),.clk(gclk));
	jdff dff_B_Kb5eZCR04_1(.din(w_dff_B_eOwKKlvL6_1),.dout(w_dff_B_Kb5eZCR04_1),.clk(gclk));
	jdff dff_B_HmmRyGwv2_1(.din(w_dff_B_Kb5eZCR04_1),.dout(w_dff_B_HmmRyGwv2_1),.clk(gclk));
	jdff dff_B_9gwTku3U3_1(.din(w_dff_B_HmmRyGwv2_1),.dout(w_dff_B_9gwTku3U3_1),.clk(gclk));
	jdff dff_B_Ob6jiuSn0_1(.din(w_dff_B_9gwTku3U3_1),.dout(w_dff_B_Ob6jiuSn0_1),.clk(gclk));
	jdff dff_B_8HEUaogz5_1(.din(w_dff_B_Ob6jiuSn0_1),.dout(w_dff_B_8HEUaogz5_1),.clk(gclk));
	jdff dff_B_Ii1lU8fb6_1(.din(w_dff_B_8HEUaogz5_1),.dout(w_dff_B_Ii1lU8fb6_1),.clk(gclk));
	jdff dff_B_DtZdYFLU3_1(.din(w_dff_B_Ii1lU8fb6_1),.dout(w_dff_B_DtZdYFLU3_1),.clk(gclk));
	jdff dff_B_AFAxx7y61_1(.din(w_dff_B_DtZdYFLU3_1),.dout(w_dff_B_AFAxx7y61_1),.clk(gclk));
	jdff dff_B_6sH0kz1P9_1(.din(w_dff_B_AFAxx7y61_1),.dout(w_dff_B_6sH0kz1P9_1),.clk(gclk));
	jdff dff_B_ljYpIwnb2_1(.din(w_dff_B_6sH0kz1P9_1),.dout(w_dff_B_ljYpIwnb2_1),.clk(gclk));
	jdff dff_B_AFjh8EhR3_1(.din(w_dff_B_ljYpIwnb2_1),.dout(w_dff_B_AFjh8EhR3_1),.clk(gclk));
	jdff dff_B_OMRA4bCC0_1(.din(w_dff_B_AFjh8EhR3_1),.dout(w_dff_B_OMRA4bCC0_1),.clk(gclk));
	jdff dff_B_GVnabYUt7_1(.din(w_dff_B_OMRA4bCC0_1),.dout(w_dff_B_GVnabYUt7_1),.clk(gclk));
	jdff dff_B_Xl68Rniz2_1(.din(w_dff_B_GVnabYUt7_1),.dout(w_dff_B_Xl68Rniz2_1),.clk(gclk));
	jdff dff_B_3zNbge5I6_1(.din(w_dff_B_Xl68Rniz2_1),.dout(w_dff_B_3zNbge5I6_1),.clk(gclk));
	jdff dff_B_5mWCnpXf3_1(.din(w_dff_B_3zNbge5I6_1),.dout(w_dff_B_5mWCnpXf3_1),.clk(gclk));
	jdff dff_B_80a8rMpB4_1(.din(w_dff_B_5mWCnpXf3_1),.dout(w_dff_B_80a8rMpB4_1),.clk(gclk));
	jdff dff_B_LcBIPVk52_1(.din(w_dff_B_80a8rMpB4_1),.dout(w_dff_B_LcBIPVk52_1),.clk(gclk));
	jdff dff_B_wkt9KDvl9_1(.din(w_dff_B_LcBIPVk52_1),.dout(w_dff_B_wkt9KDvl9_1),.clk(gclk));
	jdff dff_B_eXYZBust9_1(.din(w_dff_B_wkt9KDvl9_1),.dout(w_dff_B_eXYZBust9_1),.clk(gclk));
	jdff dff_B_UtRC0vIv2_1(.din(w_dff_B_eXYZBust9_1),.dout(w_dff_B_UtRC0vIv2_1),.clk(gclk));
	jdff dff_B_eSV6K7Yu5_1(.din(w_dff_B_UtRC0vIv2_1),.dout(w_dff_B_eSV6K7Yu5_1),.clk(gclk));
	jdff dff_B_XHpJ1g3i7_1(.din(w_dff_B_eSV6K7Yu5_1),.dout(w_dff_B_XHpJ1g3i7_1),.clk(gclk));
	jdff dff_B_tMf2eBS41_1(.din(w_dff_B_XHpJ1g3i7_1),.dout(w_dff_B_tMf2eBS41_1),.clk(gclk));
	jdff dff_B_sRPbSVa98_1(.din(w_dff_B_tMf2eBS41_1),.dout(w_dff_B_sRPbSVa98_1),.clk(gclk));
	jdff dff_B_Cv2hXfG22_1(.din(w_dff_B_sRPbSVa98_1),.dout(w_dff_B_Cv2hXfG22_1),.clk(gclk));
	jdff dff_B_0jGqNUTS9_1(.din(w_dff_B_Cv2hXfG22_1),.dout(w_dff_B_0jGqNUTS9_1),.clk(gclk));
	jdff dff_B_XmiSzfrw1_1(.din(w_dff_B_0jGqNUTS9_1),.dout(w_dff_B_XmiSzfrw1_1),.clk(gclk));
	jdff dff_B_jDHWSs2W6_1(.din(w_dff_B_XmiSzfrw1_1),.dout(w_dff_B_jDHWSs2W6_1),.clk(gclk));
	jdff dff_B_1GmN4tGU8_1(.din(w_dff_B_jDHWSs2W6_1),.dout(w_dff_B_1GmN4tGU8_1),.clk(gclk));
	jdff dff_B_Dc44K48P5_1(.din(w_dff_B_1GmN4tGU8_1),.dout(w_dff_B_Dc44K48P5_1),.clk(gclk));
	jdff dff_B_LCACFbPS9_1(.din(w_dff_B_Dc44K48P5_1),.dout(w_dff_B_LCACFbPS9_1),.clk(gclk));
	jdff dff_B_r6Eb3GYB8_1(.din(w_dff_B_LCACFbPS9_1),.dout(w_dff_B_r6Eb3GYB8_1),.clk(gclk));
	jdff dff_B_exURoR631_1(.din(w_dff_B_r6Eb3GYB8_1),.dout(w_dff_B_exURoR631_1),.clk(gclk));
	jdff dff_B_6sERNQHn1_1(.din(w_dff_B_exURoR631_1),.dout(w_dff_B_6sERNQHn1_1),.clk(gclk));
	jdff dff_B_DwNa9UBF4_1(.din(w_dff_B_6sERNQHn1_1),.dout(w_dff_B_DwNa9UBF4_1),.clk(gclk));
	jdff dff_B_Fv0wd9zd4_1(.din(w_dff_B_DwNa9UBF4_1),.dout(w_dff_B_Fv0wd9zd4_1),.clk(gclk));
	jdff dff_B_frV9Zoog4_1(.din(w_dff_B_Fv0wd9zd4_1),.dout(w_dff_B_frV9Zoog4_1),.clk(gclk));
	jdff dff_B_mUuqq02s2_1(.din(w_dff_B_frV9Zoog4_1),.dout(w_dff_B_mUuqq02s2_1),.clk(gclk));
	jdff dff_B_2Kp7A3SX6_1(.din(w_dff_B_mUuqq02s2_1),.dout(w_dff_B_2Kp7A3SX6_1),.clk(gclk));
	jdff dff_B_p73HMTjL8_1(.din(w_dff_B_2Kp7A3SX6_1),.dout(w_dff_B_p73HMTjL8_1),.clk(gclk));
	jdff dff_B_2AFVpd2l3_1(.din(w_dff_B_p73HMTjL8_1),.dout(w_dff_B_2AFVpd2l3_1),.clk(gclk));
	jdff dff_B_KJa3pqMR3_1(.din(w_dff_B_2AFVpd2l3_1),.dout(w_dff_B_KJa3pqMR3_1),.clk(gclk));
	jdff dff_B_T5YsAIWP2_1(.din(w_dff_B_KJa3pqMR3_1),.dout(w_dff_B_T5YsAIWP2_1),.clk(gclk));
	jdff dff_B_jzbrsWDm2_1(.din(w_dff_B_T5YsAIWP2_1),.dout(w_dff_B_jzbrsWDm2_1),.clk(gclk));
	jdff dff_B_GMzh451l4_1(.din(w_dff_B_jzbrsWDm2_1),.dout(w_dff_B_GMzh451l4_1),.clk(gclk));
	jdff dff_B_ycIpniEc3_1(.din(w_dff_B_GMzh451l4_1),.dout(w_dff_B_ycIpniEc3_1),.clk(gclk));
	jdff dff_B_cZ3tMkVU1_1(.din(w_dff_B_ycIpniEc3_1),.dout(w_dff_B_cZ3tMkVU1_1),.clk(gclk));
	jdff dff_B_0W3BNHKB2_1(.din(w_dff_B_cZ3tMkVU1_1),.dout(w_dff_B_0W3BNHKB2_1),.clk(gclk));
	jdff dff_B_D9zm9QL63_1(.din(w_dff_B_0W3BNHKB2_1),.dout(w_dff_B_D9zm9QL63_1),.clk(gclk));
	jdff dff_B_RjxutSIJ3_1(.din(w_dff_B_D9zm9QL63_1),.dout(w_dff_B_RjxutSIJ3_1),.clk(gclk));
	jdff dff_B_LehWGyme1_1(.din(w_dff_B_RjxutSIJ3_1),.dout(w_dff_B_LehWGyme1_1),.clk(gclk));
	jdff dff_B_IzGGpkGF4_1(.din(w_dff_B_LehWGyme1_1),.dout(w_dff_B_IzGGpkGF4_1),.clk(gclk));
	jdff dff_B_hG9jjS9b1_1(.din(w_dff_B_IzGGpkGF4_1),.dout(w_dff_B_hG9jjS9b1_1),.clk(gclk));
	jdff dff_B_Rb3hY0CN6_1(.din(w_dff_B_hG9jjS9b1_1),.dout(w_dff_B_Rb3hY0CN6_1),.clk(gclk));
	jdff dff_B_c9CPLuWJ3_1(.din(w_dff_B_Rb3hY0CN6_1),.dout(w_dff_B_c9CPLuWJ3_1),.clk(gclk));
	jdff dff_B_PHTDjAR21_1(.din(w_dff_B_c9CPLuWJ3_1),.dout(w_dff_B_PHTDjAR21_1),.clk(gclk));
	jdff dff_B_OK4Cbq2N3_1(.din(w_dff_B_PHTDjAR21_1),.dout(w_dff_B_OK4Cbq2N3_1),.clk(gclk));
	jdff dff_B_SCKtyKSI8_1(.din(w_dff_B_OK4Cbq2N3_1),.dout(w_dff_B_SCKtyKSI8_1),.clk(gclk));
	jdff dff_B_XJeY6c0D5_1(.din(w_dff_B_SCKtyKSI8_1),.dout(w_dff_B_XJeY6c0D5_1),.clk(gclk));
	jdff dff_B_SHLLeqqr4_1(.din(w_dff_B_XJeY6c0D5_1),.dout(w_dff_B_SHLLeqqr4_1),.clk(gclk));
	jdff dff_B_uP8GFxyD6_1(.din(w_dff_B_SHLLeqqr4_1),.dout(w_dff_B_uP8GFxyD6_1),.clk(gclk));
	jdff dff_B_iijEBp3U2_1(.din(w_dff_B_uP8GFxyD6_1),.dout(w_dff_B_iijEBp3U2_1),.clk(gclk));
	jdff dff_B_sTOnEMhS8_1(.din(w_dff_B_iijEBp3U2_1),.dout(w_dff_B_sTOnEMhS8_1),.clk(gclk));
	jdff dff_B_GblG97w47_1(.din(w_dff_B_sTOnEMhS8_1),.dout(w_dff_B_GblG97w47_1),.clk(gclk));
	jdff dff_B_A36wNVHx6_1(.din(w_dff_B_GblG97w47_1),.dout(w_dff_B_A36wNVHx6_1),.clk(gclk));
	jdff dff_B_USqdnUqB5_1(.din(w_dff_B_A36wNVHx6_1),.dout(w_dff_B_USqdnUqB5_1),.clk(gclk));
	jdff dff_B_KEVR8POg8_1(.din(w_dff_B_USqdnUqB5_1),.dout(w_dff_B_KEVR8POg8_1),.clk(gclk));
	jdff dff_B_JxTT3yEo9_1(.din(w_dff_B_KEVR8POg8_1),.dout(w_dff_B_JxTT3yEo9_1),.clk(gclk));
	jdff dff_B_MaMNWOS70_1(.din(w_dff_B_JxTT3yEo9_1),.dout(w_dff_B_MaMNWOS70_1),.clk(gclk));
	jdff dff_B_JELEf7Sw8_1(.din(w_dff_B_MaMNWOS70_1),.dout(w_dff_B_JELEf7Sw8_1),.clk(gclk));
	jdff dff_B_tHHHLE2j9_1(.din(w_dff_B_JELEf7Sw8_1),.dout(w_dff_B_tHHHLE2j9_1),.clk(gclk));
	jdff dff_B_VSuAiR5z5_1(.din(w_dff_B_tHHHLE2j9_1),.dout(w_dff_B_VSuAiR5z5_1),.clk(gclk));
	jdff dff_B_vJde0YQf8_1(.din(w_dff_B_VSuAiR5z5_1),.dout(w_dff_B_vJde0YQf8_1),.clk(gclk));
	jdff dff_B_XTpaCHU28_1(.din(w_dff_B_vJde0YQf8_1),.dout(w_dff_B_XTpaCHU28_1),.clk(gclk));
	jdff dff_B_pomrhoKX3_0(.din(n1027),.dout(w_dff_B_pomrhoKX3_0),.clk(gclk));
	jdff dff_B_baCcp0oq8_0(.din(w_dff_B_pomrhoKX3_0),.dout(w_dff_B_baCcp0oq8_0),.clk(gclk));
	jdff dff_B_XOUVEuQM9_0(.din(w_dff_B_baCcp0oq8_0),.dout(w_dff_B_XOUVEuQM9_0),.clk(gclk));
	jdff dff_B_iIRRvqXo2_0(.din(w_dff_B_XOUVEuQM9_0),.dout(w_dff_B_iIRRvqXo2_0),.clk(gclk));
	jdff dff_B_4ZDaoUx90_0(.din(w_dff_B_iIRRvqXo2_0),.dout(w_dff_B_4ZDaoUx90_0),.clk(gclk));
	jdff dff_B_uZ8VJFde1_0(.din(w_dff_B_4ZDaoUx90_0),.dout(w_dff_B_uZ8VJFde1_0),.clk(gclk));
	jdff dff_B_fFfeAyoS5_0(.din(w_dff_B_uZ8VJFde1_0),.dout(w_dff_B_fFfeAyoS5_0),.clk(gclk));
	jdff dff_B_vrRmLZtB7_0(.din(w_dff_B_fFfeAyoS5_0),.dout(w_dff_B_vrRmLZtB7_0),.clk(gclk));
	jdff dff_B_34i4JCfy4_0(.din(w_dff_B_vrRmLZtB7_0),.dout(w_dff_B_34i4JCfy4_0),.clk(gclk));
	jdff dff_B_e0H4W5wI5_0(.din(w_dff_B_34i4JCfy4_0),.dout(w_dff_B_e0H4W5wI5_0),.clk(gclk));
	jdff dff_B_MxyzzHXk8_0(.din(w_dff_B_e0H4W5wI5_0),.dout(w_dff_B_MxyzzHXk8_0),.clk(gclk));
	jdff dff_B_ID4vhbKP0_0(.din(w_dff_B_MxyzzHXk8_0),.dout(w_dff_B_ID4vhbKP0_0),.clk(gclk));
	jdff dff_B_lCi4MSn69_0(.din(w_dff_B_ID4vhbKP0_0),.dout(w_dff_B_lCi4MSn69_0),.clk(gclk));
	jdff dff_B_qJifAUfl6_0(.din(w_dff_B_lCi4MSn69_0),.dout(w_dff_B_qJifAUfl6_0),.clk(gclk));
	jdff dff_B_z8m25sLp9_0(.din(w_dff_B_qJifAUfl6_0),.dout(w_dff_B_z8m25sLp9_0),.clk(gclk));
	jdff dff_B_gxbjblo96_0(.din(w_dff_B_z8m25sLp9_0),.dout(w_dff_B_gxbjblo96_0),.clk(gclk));
	jdff dff_B_3yvVl3l50_0(.din(w_dff_B_gxbjblo96_0),.dout(w_dff_B_3yvVl3l50_0),.clk(gclk));
	jdff dff_B_QABOeMfz6_0(.din(w_dff_B_3yvVl3l50_0),.dout(w_dff_B_QABOeMfz6_0),.clk(gclk));
	jdff dff_B_YZSuemMn5_0(.din(w_dff_B_QABOeMfz6_0),.dout(w_dff_B_YZSuemMn5_0),.clk(gclk));
	jdff dff_B_omGWFeWB4_0(.din(w_dff_B_YZSuemMn5_0),.dout(w_dff_B_omGWFeWB4_0),.clk(gclk));
	jdff dff_B_CRL12axe7_0(.din(w_dff_B_omGWFeWB4_0),.dout(w_dff_B_CRL12axe7_0),.clk(gclk));
	jdff dff_B_SiufHU2S1_0(.din(w_dff_B_CRL12axe7_0),.dout(w_dff_B_SiufHU2S1_0),.clk(gclk));
	jdff dff_B_FKrAPskI5_0(.din(w_dff_B_SiufHU2S1_0),.dout(w_dff_B_FKrAPskI5_0),.clk(gclk));
	jdff dff_B_ee2L7aO76_0(.din(w_dff_B_FKrAPskI5_0),.dout(w_dff_B_ee2L7aO76_0),.clk(gclk));
	jdff dff_B_1hrnuihP5_0(.din(w_dff_B_ee2L7aO76_0),.dout(w_dff_B_1hrnuihP5_0),.clk(gclk));
	jdff dff_B_0iKcyB6a0_0(.din(w_dff_B_1hrnuihP5_0),.dout(w_dff_B_0iKcyB6a0_0),.clk(gclk));
	jdff dff_B_Me5b1PGq4_0(.din(w_dff_B_0iKcyB6a0_0),.dout(w_dff_B_Me5b1PGq4_0),.clk(gclk));
	jdff dff_B_oyEvkl4H7_0(.din(w_dff_B_Me5b1PGq4_0),.dout(w_dff_B_oyEvkl4H7_0),.clk(gclk));
	jdff dff_B_gDCeEwbQ4_0(.din(w_dff_B_oyEvkl4H7_0),.dout(w_dff_B_gDCeEwbQ4_0),.clk(gclk));
	jdff dff_B_3iU4jI8b5_0(.din(w_dff_B_gDCeEwbQ4_0),.dout(w_dff_B_3iU4jI8b5_0),.clk(gclk));
	jdff dff_B_gLWVFxL25_0(.din(w_dff_B_3iU4jI8b5_0),.dout(w_dff_B_gLWVFxL25_0),.clk(gclk));
	jdff dff_B_xZNckrrA1_0(.din(w_dff_B_gLWVFxL25_0),.dout(w_dff_B_xZNckrrA1_0),.clk(gclk));
	jdff dff_B_0BLRsOe23_0(.din(w_dff_B_xZNckrrA1_0),.dout(w_dff_B_0BLRsOe23_0),.clk(gclk));
	jdff dff_B_KcUXHiAH5_0(.din(w_dff_B_0BLRsOe23_0),.dout(w_dff_B_KcUXHiAH5_0),.clk(gclk));
	jdff dff_B_nKmcGCwL3_0(.din(w_dff_B_KcUXHiAH5_0),.dout(w_dff_B_nKmcGCwL3_0),.clk(gclk));
	jdff dff_B_hR41QYdD6_0(.din(w_dff_B_nKmcGCwL3_0),.dout(w_dff_B_hR41QYdD6_0),.clk(gclk));
	jdff dff_B_D48VAFVc8_0(.din(w_dff_B_hR41QYdD6_0),.dout(w_dff_B_D48VAFVc8_0),.clk(gclk));
	jdff dff_B_J36eJ6qG6_0(.din(w_dff_B_D48VAFVc8_0),.dout(w_dff_B_J36eJ6qG6_0),.clk(gclk));
	jdff dff_B_DpDdnZDY4_0(.din(w_dff_B_J36eJ6qG6_0),.dout(w_dff_B_DpDdnZDY4_0),.clk(gclk));
	jdff dff_B_xoxvbiiT5_0(.din(w_dff_B_DpDdnZDY4_0),.dout(w_dff_B_xoxvbiiT5_0),.clk(gclk));
	jdff dff_B_jXZa1wDf4_0(.din(w_dff_B_xoxvbiiT5_0),.dout(w_dff_B_jXZa1wDf4_0),.clk(gclk));
	jdff dff_B_SKy6bEDi4_0(.din(w_dff_B_jXZa1wDf4_0),.dout(w_dff_B_SKy6bEDi4_0),.clk(gclk));
	jdff dff_B_i2msDnMm6_0(.din(w_dff_B_SKy6bEDi4_0),.dout(w_dff_B_i2msDnMm6_0),.clk(gclk));
	jdff dff_B_QlPHvjD14_0(.din(w_dff_B_i2msDnMm6_0),.dout(w_dff_B_QlPHvjD14_0),.clk(gclk));
	jdff dff_B_WWffVfOq9_0(.din(w_dff_B_QlPHvjD14_0),.dout(w_dff_B_WWffVfOq9_0),.clk(gclk));
	jdff dff_B_gByYrllJ4_0(.din(w_dff_B_WWffVfOq9_0),.dout(w_dff_B_gByYrllJ4_0),.clk(gclk));
	jdff dff_B_SoARTfZF5_0(.din(w_dff_B_gByYrllJ4_0),.dout(w_dff_B_SoARTfZF5_0),.clk(gclk));
	jdff dff_B_CTyDAvbT0_0(.din(w_dff_B_SoARTfZF5_0),.dout(w_dff_B_CTyDAvbT0_0),.clk(gclk));
	jdff dff_B_pAICIYvP2_0(.din(w_dff_B_CTyDAvbT0_0),.dout(w_dff_B_pAICIYvP2_0),.clk(gclk));
	jdff dff_B_QDJNz9Tm3_0(.din(w_dff_B_pAICIYvP2_0),.dout(w_dff_B_QDJNz9Tm3_0),.clk(gclk));
	jdff dff_B_ztoT0opx6_0(.din(w_dff_B_QDJNz9Tm3_0),.dout(w_dff_B_ztoT0opx6_0),.clk(gclk));
	jdff dff_B_JxICGcUt9_0(.din(w_dff_B_ztoT0opx6_0),.dout(w_dff_B_JxICGcUt9_0),.clk(gclk));
	jdff dff_B_myoXOUum0_0(.din(w_dff_B_JxICGcUt9_0),.dout(w_dff_B_myoXOUum0_0),.clk(gclk));
	jdff dff_B_E5W8l5If0_0(.din(w_dff_B_myoXOUum0_0),.dout(w_dff_B_E5W8l5If0_0),.clk(gclk));
	jdff dff_B_Ft7QBMg95_0(.din(w_dff_B_E5W8l5If0_0),.dout(w_dff_B_Ft7QBMg95_0),.clk(gclk));
	jdff dff_B_qiBKn6Kg7_0(.din(w_dff_B_Ft7QBMg95_0),.dout(w_dff_B_qiBKn6Kg7_0),.clk(gclk));
	jdff dff_B_sTK66WS13_0(.din(w_dff_B_qiBKn6Kg7_0),.dout(w_dff_B_sTK66WS13_0),.clk(gclk));
	jdff dff_B_mV9AOvXr2_0(.din(w_dff_B_sTK66WS13_0),.dout(w_dff_B_mV9AOvXr2_0),.clk(gclk));
	jdff dff_B_btB1mEKx3_0(.din(w_dff_B_mV9AOvXr2_0),.dout(w_dff_B_btB1mEKx3_0),.clk(gclk));
	jdff dff_B_0wtbn10a4_0(.din(w_dff_B_btB1mEKx3_0),.dout(w_dff_B_0wtbn10a4_0),.clk(gclk));
	jdff dff_B_nxcFl2bI5_0(.din(w_dff_B_0wtbn10a4_0),.dout(w_dff_B_nxcFl2bI5_0),.clk(gclk));
	jdff dff_B_JVtan3Qz4_0(.din(w_dff_B_nxcFl2bI5_0),.dout(w_dff_B_JVtan3Qz4_0),.clk(gclk));
	jdff dff_B_IKBhzfGn2_0(.din(w_dff_B_JVtan3Qz4_0),.dout(w_dff_B_IKBhzfGn2_0),.clk(gclk));
	jdff dff_B_xBRBwFRm5_0(.din(w_dff_B_IKBhzfGn2_0),.dout(w_dff_B_xBRBwFRm5_0),.clk(gclk));
	jdff dff_B_xxfuCkD96_0(.din(w_dff_B_xBRBwFRm5_0),.dout(w_dff_B_xxfuCkD96_0),.clk(gclk));
	jdff dff_B_BNuSu2Ox9_0(.din(w_dff_B_xxfuCkD96_0),.dout(w_dff_B_BNuSu2Ox9_0),.clk(gclk));
	jdff dff_B_BUFmk3Cl2_0(.din(w_dff_B_BNuSu2Ox9_0),.dout(w_dff_B_BUFmk3Cl2_0),.clk(gclk));
	jdff dff_B_3RqGMbzc2_0(.din(w_dff_B_BUFmk3Cl2_0),.dout(w_dff_B_3RqGMbzc2_0),.clk(gclk));
	jdff dff_B_KF1K7Qfd5_0(.din(w_dff_B_3RqGMbzc2_0),.dout(w_dff_B_KF1K7Qfd5_0),.clk(gclk));
	jdff dff_B_PoVtOAqm5_0(.din(w_dff_B_KF1K7Qfd5_0),.dout(w_dff_B_PoVtOAqm5_0),.clk(gclk));
	jdff dff_B_5AHgWFZh4_0(.din(w_dff_B_PoVtOAqm5_0),.dout(w_dff_B_5AHgWFZh4_0),.clk(gclk));
	jdff dff_B_Mlpajz0y5_0(.din(w_dff_B_5AHgWFZh4_0),.dout(w_dff_B_Mlpajz0y5_0),.clk(gclk));
	jdff dff_B_sOaWQa9i1_0(.din(w_dff_B_Mlpajz0y5_0),.dout(w_dff_B_sOaWQa9i1_0),.clk(gclk));
	jdff dff_B_P5NahKIs3_0(.din(w_dff_B_sOaWQa9i1_0),.dout(w_dff_B_P5NahKIs3_0),.clk(gclk));
	jdff dff_B_jpCQUsBu6_0(.din(w_dff_B_P5NahKIs3_0),.dout(w_dff_B_jpCQUsBu6_0),.clk(gclk));
	jdff dff_B_cOIt78Ng7_0(.din(w_dff_B_jpCQUsBu6_0),.dout(w_dff_B_cOIt78Ng7_0),.clk(gclk));
	jdff dff_B_cvbQq8QU1_0(.din(w_dff_B_cOIt78Ng7_0),.dout(w_dff_B_cvbQq8QU1_0),.clk(gclk));
	jdff dff_B_rdF4XIZ41_0(.din(w_dff_B_cvbQq8QU1_0),.dout(w_dff_B_rdF4XIZ41_0),.clk(gclk));
	jdff dff_B_qrvbyXEo2_0(.din(w_dff_B_rdF4XIZ41_0),.dout(w_dff_B_qrvbyXEo2_0),.clk(gclk));
	jdff dff_B_6qNdAErD0_0(.din(w_dff_B_qrvbyXEo2_0),.dout(w_dff_B_6qNdAErD0_0),.clk(gclk));
	jdff dff_B_RjWmkJTb4_0(.din(w_dff_B_6qNdAErD0_0),.dout(w_dff_B_RjWmkJTb4_0),.clk(gclk));
	jdff dff_B_zFAUXzQW6_0(.din(w_dff_B_RjWmkJTb4_0),.dout(w_dff_B_zFAUXzQW6_0),.clk(gclk));
	jdff dff_B_YAx3gkgB4_0(.din(w_dff_B_zFAUXzQW6_0),.dout(w_dff_B_YAx3gkgB4_0),.clk(gclk));
	jdff dff_B_VbXmrZlD6_0(.din(w_dff_B_YAx3gkgB4_0),.dout(w_dff_B_VbXmrZlD6_0),.clk(gclk));
	jdff dff_B_gO0JsDvz1_0(.din(w_dff_B_VbXmrZlD6_0),.dout(w_dff_B_gO0JsDvz1_0),.clk(gclk));
	jdff dff_B_ONFmeABu9_0(.din(w_dff_B_gO0JsDvz1_0),.dout(w_dff_B_ONFmeABu9_0),.clk(gclk));
	jdff dff_B_LKNqEdxf1_0(.din(w_dff_B_ONFmeABu9_0),.dout(w_dff_B_LKNqEdxf1_0),.clk(gclk));
	jdff dff_B_aJ5CKMW35_0(.din(w_dff_B_LKNqEdxf1_0),.dout(w_dff_B_aJ5CKMW35_0),.clk(gclk));
	jdff dff_B_McxDPGt43_0(.din(w_dff_B_aJ5CKMW35_0),.dout(w_dff_B_McxDPGt43_0),.clk(gclk));
	jdff dff_B_wZAa0PfI2_0(.din(w_dff_B_McxDPGt43_0),.dout(w_dff_B_wZAa0PfI2_0),.clk(gclk));
	jdff dff_B_iuIi85S93_0(.din(w_dff_B_wZAa0PfI2_0),.dout(w_dff_B_iuIi85S93_0),.clk(gclk));
	jdff dff_B_xHnBmQFG1_0(.din(w_dff_B_iuIi85S93_0),.dout(w_dff_B_xHnBmQFG1_0),.clk(gclk));
	jdff dff_B_TWSyTdm77_0(.din(w_dff_B_xHnBmQFG1_0),.dout(w_dff_B_TWSyTdm77_0),.clk(gclk));
	jdff dff_B_sZjpofVw6_0(.din(w_dff_B_TWSyTdm77_0),.dout(w_dff_B_sZjpofVw6_0),.clk(gclk));
	jdff dff_B_NsxZKiOO6_0(.din(w_dff_B_sZjpofVw6_0),.dout(w_dff_B_NsxZKiOO6_0),.clk(gclk));
	jdff dff_B_oHPeoiAT6_0(.din(w_dff_B_NsxZKiOO6_0),.dout(w_dff_B_oHPeoiAT6_0),.clk(gclk));
	jdff dff_B_KT71PfDa5_0(.din(w_dff_B_oHPeoiAT6_0),.dout(w_dff_B_KT71PfDa5_0),.clk(gclk));
	jdff dff_B_AKO3xROQ2_0(.din(w_dff_B_KT71PfDa5_0),.dout(w_dff_B_AKO3xROQ2_0),.clk(gclk));
	jdff dff_B_Ew6PCfXS9_0(.din(w_dff_B_AKO3xROQ2_0),.dout(w_dff_B_Ew6PCfXS9_0),.clk(gclk));
	jdff dff_B_cdTRIFdt5_0(.din(w_dff_B_Ew6PCfXS9_0),.dout(w_dff_B_cdTRIFdt5_0),.clk(gclk));
	jdff dff_B_jEqqGPwr8_0(.din(w_dff_B_cdTRIFdt5_0),.dout(w_dff_B_jEqqGPwr8_0),.clk(gclk));
	jdff dff_B_DmEpAyja3_0(.din(w_dff_B_jEqqGPwr8_0),.dout(w_dff_B_DmEpAyja3_0),.clk(gclk));
	jdff dff_B_upEAL2tH7_0(.din(w_dff_B_DmEpAyja3_0),.dout(w_dff_B_upEAL2tH7_0),.clk(gclk));
	jdff dff_B_pZy9ywM63_0(.din(w_dff_B_upEAL2tH7_0),.dout(w_dff_B_pZy9ywM63_0),.clk(gclk));
	jdff dff_B_RSVqasus7_0(.din(w_dff_B_pZy9ywM63_0),.dout(w_dff_B_RSVqasus7_0),.clk(gclk));
	jdff dff_B_UcLcfnEH4_0(.din(w_dff_B_RSVqasus7_0),.dout(w_dff_B_UcLcfnEH4_0),.clk(gclk));
	jdff dff_B_rQs1ywwY3_0(.din(w_dff_B_UcLcfnEH4_0),.dout(w_dff_B_rQs1ywwY3_0),.clk(gclk));
	jdff dff_B_ziLTM7Mv0_1(.din(n1020),.dout(w_dff_B_ziLTM7Mv0_1),.clk(gclk));
	jdff dff_B_JppgMvTB2_1(.din(w_dff_B_ziLTM7Mv0_1),.dout(w_dff_B_JppgMvTB2_1),.clk(gclk));
	jdff dff_B_5zp088EI0_1(.din(w_dff_B_JppgMvTB2_1),.dout(w_dff_B_5zp088EI0_1),.clk(gclk));
	jdff dff_B_unK8V57A2_1(.din(w_dff_B_5zp088EI0_1),.dout(w_dff_B_unK8V57A2_1),.clk(gclk));
	jdff dff_B_JXqkLCk36_1(.din(w_dff_B_unK8V57A2_1),.dout(w_dff_B_JXqkLCk36_1),.clk(gclk));
	jdff dff_B_zkiwK9dx7_1(.din(w_dff_B_JXqkLCk36_1),.dout(w_dff_B_zkiwK9dx7_1),.clk(gclk));
	jdff dff_B_bVzakFPN1_1(.din(w_dff_B_zkiwK9dx7_1),.dout(w_dff_B_bVzakFPN1_1),.clk(gclk));
	jdff dff_B_rV34xDOI2_1(.din(w_dff_B_bVzakFPN1_1),.dout(w_dff_B_rV34xDOI2_1),.clk(gclk));
	jdff dff_B_HaBCZKri7_1(.din(w_dff_B_rV34xDOI2_1),.dout(w_dff_B_HaBCZKri7_1),.clk(gclk));
	jdff dff_B_uvp4uylE9_1(.din(w_dff_B_HaBCZKri7_1),.dout(w_dff_B_uvp4uylE9_1),.clk(gclk));
	jdff dff_B_uUagZVog8_1(.din(w_dff_B_uvp4uylE9_1),.dout(w_dff_B_uUagZVog8_1),.clk(gclk));
	jdff dff_B_pdrJnaYb7_1(.din(w_dff_B_uUagZVog8_1),.dout(w_dff_B_pdrJnaYb7_1),.clk(gclk));
	jdff dff_B_W7msf6WW5_1(.din(w_dff_B_pdrJnaYb7_1),.dout(w_dff_B_W7msf6WW5_1),.clk(gclk));
	jdff dff_B_wm3x5N3G3_1(.din(w_dff_B_W7msf6WW5_1),.dout(w_dff_B_wm3x5N3G3_1),.clk(gclk));
	jdff dff_B_DYvucooa8_1(.din(w_dff_B_wm3x5N3G3_1),.dout(w_dff_B_DYvucooa8_1),.clk(gclk));
	jdff dff_B_71pfdEjU0_1(.din(w_dff_B_DYvucooa8_1),.dout(w_dff_B_71pfdEjU0_1),.clk(gclk));
	jdff dff_B_j5GrO96V5_1(.din(w_dff_B_71pfdEjU0_1),.dout(w_dff_B_j5GrO96V5_1),.clk(gclk));
	jdff dff_B_Q8RSgHzH0_1(.din(w_dff_B_j5GrO96V5_1),.dout(w_dff_B_Q8RSgHzH0_1),.clk(gclk));
	jdff dff_B_qFIK46ND6_1(.din(w_dff_B_Q8RSgHzH0_1),.dout(w_dff_B_qFIK46ND6_1),.clk(gclk));
	jdff dff_B_i1GCqMrP5_1(.din(w_dff_B_qFIK46ND6_1),.dout(w_dff_B_i1GCqMrP5_1),.clk(gclk));
	jdff dff_B_quhWUEMl4_1(.din(w_dff_B_i1GCqMrP5_1),.dout(w_dff_B_quhWUEMl4_1),.clk(gclk));
	jdff dff_B_9QliUMWL2_1(.din(w_dff_B_quhWUEMl4_1),.dout(w_dff_B_9QliUMWL2_1),.clk(gclk));
	jdff dff_B_nWU6iosP7_1(.din(w_dff_B_9QliUMWL2_1),.dout(w_dff_B_nWU6iosP7_1),.clk(gclk));
	jdff dff_B_3munYuCa3_1(.din(w_dff_B_nWU6iosP7_1),.dout(w_dff_B_3munYuCa3_1),.clk(gclk));
	jdff dff_B_QMnnd6x60_1(.din(w_dff_B_3munYuCa3_1),.dout(w_dff_B_QMnnd6x60_1),.clk(gclk));
	jdff dff_B_n5KH8bNc1_1(.din(w_dff_B_QMnnd6x60_1),.dout(w_dff_B_n5KH8bNc1_1),.clk(gclk));
	jdff dff_B_2Fa5s8bH3_1(.din(w_dff_B_n5KH8bNc1_1),.dout(w_dff_B_2Fa5s8bH3_1),.clk(gclk));
	jdff dff_B_X9InJHaX0_1(.din(w_dff_B_2Fa5s8bH3_1),.dout(w_dff_B_X9InJHaX0_1),.clk(gclk));
	jdff dff_B_0mtu47He4_1(.din(w_dff_B_X9InJHaX0_1),.dout(w_dff_B_0mtu47He4_1),.clk(gclk));
	jdff dff_B_sdshQXGJ1_1(.din(w_dff_B_0mtu47He4_1),.dout(w_dff_B_sdshQXGJ1_1),.clk(gclk));
	jdff dff_B_kc1a2mbG4_1(.din(w_dff_B_sdshQXGJ1_1),.dout(w_dff_B_kc1a2mbG4_1),.clk(gclk));
	jdff dff_B_krp0yNrd0_1(.din(w_dff_B_kc1a2mbG4_1),.dout(w_dff_B_krp0yNrd0_1),.clk(gclk));
	jdff dff_B_SuZoj0JQ9_1(.din(w_dff_B_krp0yNrd0_1),.dout(w_dff_B_SuZoj0JQ9_1),.clk(gclk));
	jdff dff_B_jF7oMYoN4_1(.din(w_dff_B_SuZoj0JQ9_1),.dout(w_dff_B_jF7oMYoN4_1),.clk(gclk));
	jdff dff_B_84jn34NM7_1(.din(w_dff_B_jF7oMYoN4_1),.dout(w_dff_B_84jn34NM7_1),.clk(gclk));
	jdff dff_B_GEe2zmwU5_1(.din(w_dff_B_84jn34NM7_1),.dout(w_dff_B_GEe2zmwU5_1),.clk(gclk));
	jdff dff_B_o7y7ePYZ2_1(.din(w_dff_B_GEe2zmwU5_1),.dout(w_dff_B_o7y7ePYZ2_1),.clk(gclk));
	jdff dff_B_DmdVwadQ2_1(.din(w_dff_B_o7y7ePYZ2_1),.dout(w_dff_B_DmdVwadQ2_1),.clk(gclk));
	jdff dff_B_s0Zdac2D0_1(.din(w_dff_B_DmdVwadQ2_1),.dout(w_dff_B_s0Zdac2D0_1),.clk(gclk));
	jdff dff_B_d6Jw8NPt8_1(.din(w_dff_B_s0Zdac2D0_1),.dout(w_dff_B_d6Jw8NPt8_1),.clk(gclk));
	jdff dff_B_VJ2ycxkd5_1(.din(w_dff_B_d6Jw8NPt8_1),.dout(w_dff_B_VJ2ycxkd5_1),.clk(gclk));
	jdff dff_B_yBKYa5tC2_1(.din(w_dff_B_VJ2ycxkd5_1),.dout(w_dff_B_yBKYa5tC2_1),.clk(gclk));
	jdff dff_B_WwlNXJEA9_1(.din(w_dff_B_yBKYa5tC2_1),.dout(w_dff_B_WwlNXJEA9_1),.clk(gclk));
	jdff dff_B_VNuqwP7b9_1(.din(w_dff_B_WwlNXJEA9_1),.dout(w_dff_B_VNuqwP7b9_1),.clk(gclk));
	jdff dff_B_MDKUS8Pu5_1(.din(w_dff_B_VNuqwP7b9_1),.dout(w_dff_B_MDKUS8Pu5_1),.clk(gclk));
	jdff dff_B_O0H5SKCC9_1(.din(w_dff_B_MDKUS8Pu5_1),.dout(w_dff_B_O0H5SKCC9_1),.clk(gclk));
	jdff dff_B_XPoRxyEJ4_1(.din(w_dff_B_O0H5SKCC9_1),.dout(w_dff_B_XPoRxyEJ4_1),.clk(gclk));
	jdff dff_B_iIYXcv9I7_1(.din(w_dff_B_XPoRxyEJ4_1),.dout(w_dff_B_iIYXcv9I7_1),.clk(gclk));
	jdff dff_B_cGpMQEVd7_1(.din(w_dff_B_iIYXcv9I7_1),.dout(w_dff_B_cGpMQEVd7_1),.clk(gclk));
	jdff dff_B_A8motzwi4_1(.din(w_dff_B_cGpMQEVd7_1),.dout(w_dff_B_A8motzwi4_1),.clk(gclk));
	jdff dff_B_XSAuaGPJ8_1(.din(w_dff_B_A8motzwi4_1),.dout(w_dff_B_XSAuaGPJ8_1),.clk(gclk));
	jdff dff_B_jVEmj9RX3_1(.din(w_dff_B_XSAuaGPJ8_1),.dout(w_dff_B_jVEmj9RX3_1),.clk(gclk));
	jdff dff_B_pBRve9tm9_1(.din(w_dff_B_jVEmj9RX3_1),.dout(w_dff_B_pBRve9tm9_1),.clk(gclk));
	jdff dff_B_RW1RUIVr6_1(.din(w_dff_B_pBRve9tm9_1),.dout(w_dff_B_RW1RUIVr6_1),.clk(gclk));
	jdff dff_B_clRH3NjO5_1(.din(w_dff_B_RW1RUIVr6_1),.dout(w_dff_B_clRH3NjO5_1),.clk(gclk));
	jdff dff_B_3al7Lryt9_1(.din(w_dff_B_clRH3NjO5_1),.dout(w_dff_B_3al7Lryt9_1),.clk(gclk));
	jdff dff_B_qM4pHBPP0_1(.din(w_dff_B_3al7Lryt9_1),.dout(w_dff_B_qM4pHBPP0_1),.clk(gclk));
	jdff dff_B_3VREC1Y76_1(.din(w_dff_B_qM4pHBPP0_1),.dout(w_dff_B_3VREC1Y76_1),.clk(gclk));
	jdff dff_B_oaf5EENS7_1(.din(w_dff_B_3VREC1Y76_1),.dout(w_dff_B_oaf5EENS7_1),.clk(gclk));
	jdff dff_B_frKGwZtW4_1(.din(w_dff_B_oaf5EENS7_1),.dout(w_dff_B_frKGwZtW4_1),.clk(gclk));
	jdff dff_B_WKOv21Kw1_1(.din(w_dff_B_frKGwZtW4_1),.dout(w_dff_B_WKOv21Kw1_1),.clk(gclk));
	jdff dff_B_Mn5eYnsu7_1(.din(w_dff_B_WKOv21Kw1_1),.dout(w_dff_B_Mn5eYnsu7_1),.clk(gclk));
	jdff dff_B_rExBtcga4_1(.din(w_dff_B_Mn5eYnsu7_1),.dout(w_dff_B_rExBtcga4_1),.clk(gclk));
	jdff dff_B_8J85daFQ8_1(.din(w_dff_B_rExBtcga4_1),.dout(w_dff_B_8J85daFQ8_1),.clk(gclk));
	jdff dff_B_ygfmDo1b7_1(.din(w_dff_B_8J85daFQ8_1),.dout(w_dff_B_ygfmDo1b7_1),.clk(gclk));
	jdff dff_B_KvnvNw4R9_1(.din(w_dff_B_ygfmDo1b7_1),.dout(w_dff_B_KvnvNw4R9_1),.clk(gclk));
	jdff dff_B_7QLk3Ih44_1(.din(w_dff_B_KvnvNw4R9_1),.dout(w_dff_B_7QLk3Ih44_1),.clk(gclk));
	jdff dff_B_FZMpEpWQ3_1(.din(w_dff_B_7QLk3Ih44_1),.dout(w_dff_B_FZMpEpWQ3_1),.clk(gclk));
	jdff dff_B_DSFliSsu4_1(.din(w_dff_B_FZMpEpWQ3_1),.dout(w_dff_B_DSFliSsu4_1),.clk(gclk));
	jdff dff_B_878ETSX64_1(.din(w_dff_B_DSFliSsu4_1),.dout(w_dff_B_878ETSX64_1),.clk(gclk));
	jdff dff_B_J93ErqUJ7_1(.din(w_dff_B_878ETSX64_1),.dout(w_dff_B_J93ErqUJ7_1),.clk(gclk));
	jdff dff_B_NC08NBCG9_1(.din(w_dff_B_J93ErqUJ7_1),.dout(w_dff_B_NC08NBCG9_1),.clk(gclk));
	jdff dff_B_uGapLXyd4_1(.din(w_dff_B_NC08NBCG9_1),.dout(w_dff_B_uGapLXyd4_1),.clk(gclk));
	jdff dff_B_dVujtNXs2_1(.din(w_dff_B_uGapLXyd4_1),.dout(w_dff_B_dVujtNXs2_1),.clk(gclk));
	jdff dff_B_1MsgKfBg1_1(.din(w_dff_B_dVujtNXs2_1),.dout(w_dff_B_1MsgKfBg1_1),.clk(gclk));
	jdff dff_B_LFvfSxTj5_1(.din(w_dff_B_1MsgKfBg1_1),.dout(w_dff_B_LFvfSxTj5_1),.clk(gclk));
	jdff dff_B_0IluKIdd7_1(.din(w_dff_B_LFvfSxTj5_1),.dout(w_dff_B_0IluKIdd7_1),.clk(gclk));
	jdff dff_B_U1BsWREF0_1(.din(w_dff_B_0IluKIdd7_1),.dout(w_dff_B_U1BsWREF0_1),.clk(gclk));
	jdff dff_B_0fLTMB6u3_1(.din(w_dff_B_U1BsWREF0_1),.dout(w_dff_B_0fLTMB6u3_1),.clk(gclk));
	jdff dff_B_DbXPuAl33_1(.din(w_dff_B_0fLTMB6u3_1),.dout(w_dff_B_DbXPuAl33_1),.clk(gclk));
	jdff dff_B_cXuSid1T2_1(.din(w_dff_B_DbXPuAl33_1),.dout(w_dff_B_cXuSid1T2_1),.clk(gclk));
	jdff dff_B_OvgwmrmJ3_1(.din(w_dff_B_cXuSid1T2_1),.dout(w_dff_B_OvgwmrmJ3_1),.clk(gclk));
	jdff dff_B_aRnlNRVT0_1(.din(w_dff_B_OvgwmrmJ3_1),.dout(w_dff_B_aRnlNRVT0_1),.clk(gclk));
	jdff dff_B_dhbKDunM6_1(.din(w_dff_B_aRnlNRVT0_1),.dout(w_dff_B_dhbKDunM6_1),.clk(gclk));
	jdff dff_B_IuWdFmHJ7_1(.din(w_dff_B_dhbKDunM6_1),.dout(w_dff_B_IuWdFmHJ7_1),.clk(gclk));
	jdff dff_B_AlI43VYf3_1(.din(w_dff_B_IuWdFmHJ7_1),.dout(w_dff_B_AlI43VYf3_1),.clk(gclk));
	jdff dff_B_fQDL9vth7_1(.din(w_dff_B_AlI43VYf3_1),.dout(w_dff_B_fQDL9vth7_1),.clk(gclk));
	jdff dff_B_TDh6r4uK3_1(.din(w_dff_B_fQDL9vth7_1),.dout(w_dff_B_TDh6r4uK3_1),.clk(gclk));
	jdff dff_B_ANVQHhKt8_1(.din(w_dff_B_TDh6r4uK3_1),.dout(w_dff_B_ANVQHhKt8_1),.clk(gclk));
	jdff dff_B_lodUgsRh3_1(.din(w_dff_B_ANVQHhKt8_1),.dout(w_dff_B_lodUgsRh3_1),.clk(gclk));
	jdff dff_B_1ynOt1R01_1(.din(w_dff_B_lodUgsRh3_1),.dout(w_dff_B_1ynOt1R01_1),.clk(gclk));
	jdff dff_B_RF6UXE7p6_1(.din(w_dff_B_1ynOt1R01_1),.dout(w_dff_B_RF6UXE7p6_1),.clk(gclk));
	jdff dff_B_h0Ac4r5T2_1(.din(w_dff_B_RF6UXE7p6_1),.dout(w_dff_B_h0Ac4r5T2_1),.clk(gclk));
	jdff dff_B_YJVK6OyD2_1(.din(w_dff_B_h0Ac4r5T2_1),.dout(w_dff_B_YJVK6OyD2_1),.clk(gclk));
	jdff dff_B_ib1jukmZ7_1(.din(w_dff_B_YJVK6OyD2_1),.dout(w_dff_B_ib1jukmZ7_1),.clk(gclk));
	jdff dff_B_p1guUylt9_1(.din(w_dff_B_ib1jukmZ7_1),.dout(w_dff_B_p1guUylt9_1),.clk(gclk));
	jdff dff_B_yREBVfuC2_1(.din(w_dff_B_p1guUylt9_1),.dout(w_dff_B_yREBVfuC2_1),.clk(gclk));
	jdff dff_B_bE3hAoWJ1_1(.din(w_dff_B_yREBVfuC2_1),.dout(w_dff_B_bE3hAoWJ1_1),.clk(gclk));
	jdff dff_B_fMz32HQt4_1(.din(w_dff_B_bE3hAoWJ1_1),.dout(w_dff_B_fMz32HQt4_1),.clk(gclk));
	jdff dff_B_DhLmN5zo3_1(.din(w_dff_B_fMz32HQt4_1),.dout(w_dff_B_DhLmN5zo3_1),.clk(gclk));
	jdff dff_B_2F0z03f70_1(.din(w_dff_B_DhLmN5zo3_1),.dout(w_dff_B_2F0z03f70_1),.clk(gclk));
	jdff dff_B_JP2X0w3b5_1(.din(w_dff_B_2F0z03f70_1),.dout(w_dff_B_JP2X0w3b5_1),.clk(gclk));
	jdff dff_B_X4nabGQI4_1(.din(w_dff_B_JP2X0w3b5_1),.dout(w_dff_B_X4nabGQI4_1),.clk(gclk));
	jdff dff_B_9FOoyu9q4_1(.din(w_dff_B_X4nabGQI4_1),.dout(w_dff_B_9FOoyu9q4_1),.clk(gclk));
	jdff dff_B_r6CCakIW7_1(.din(w_dff_B_9FOoyu9q4_1),.dout(w_dff_B_r6CCakIW7_1),.clk(gclk));
	jdff dff_B_P8u9UvcR2_1(.din(w_dff_B_r6CCakIW7_1),.dout(w_dff_B_P8u9UvcR2_1),.clk(gclk));
	jdff dff_B_29wQ6VC00_0(.din(n1021),.dout(w_dff_B_29wQ6VC00_0),.clk(gclk));
	jdff dff_B_95cyNm3X7_0(.din(w_dff_B_29wQ6VC00_0),.dout(w_dff_B_95cyNm3X7_0),.clk(gclk));
	jdff dff_B_0pkdsav03_0(.din(w_dff_B_95cyNm3X7_0),.dout(w_dff_B_0pkdsav03_0),.clk(gclk));
	jdff dff_B_VpEujyx84_0(.din(w_dff_B_0pkdsav03_0),.dout(w_dff_B_VpEujyx84_0),.clk(gclk));
	jdff dff_B_DcU3epRh2_0(.din(w_dff_B_VpEujyx84_0),.dout(w_dff_B_DcU3epRh2_0),.clk(gclk));
	jdff dff_B_3psZYbWh2_0(.din(w_dff_B_DcU3epRh2_0),.dout(w_dff_B_3psZYbWh2_0),.clk(gclk));
	jdff dff_B_mekTVtDp1_0(.din(w_dff_B_3psZYbWh2_0),.dout(w_dff_B_mekTVtDp1_0),.clk(gclk));
	jdff dff_B_AFdrrYpY1_0(.din(w_dff_B_mekTVtDp1_0),.dout(w_dff_B_AFdrrYpY1_0),.clk(gclk));
	jdff dff_B_YlpETyDe2_0(.din(w_dff_B_AFdrrYpY1_0),.dout(w_dff_B_YlpETyDe2_0),.clk(gclk));
	jdff dff_B_LtoigXS11_0(.din(w_dff_B_YlpETyDe2_0),.dout(w_dff_B_LtoigXS11_0),.clk(gclk));
	jdff dff_B_lnAMYQyf8_0(.din(w_dff_B_LtoigXS11_0),.dout(w_dff_B_lnAMYQyf8_0),.clk(gclk));
	jdff dff_B_gOMiQl1u6_0(.din(w_dff_B_lnAMYQyf8_0),.dout(w_dff_B_gOMiQl1u6_0),.clk(gclk));
	jdff dff_B_LS5sbzif0_0(.din(w_dff_B_gOMiQl1u6_0),.dout(w_dff_B_LS5sbzif0_0),.clk(gclk));
	jdff dff_B_i6BHeBTb2_0(.din(w_dff_B_LS5sbzif0_0),.dout(w_dff_B_i6BHeBTb2_0),.clk(gclk));
	jdff dff_B_mIN3d78w1_0(.din(w_dff_B_i6BHeBTb2_0),.dout(w_dff_B_mIN3d78w1_0),.clk(gclk));
	jdff dff_B_Ye3TTZcF1_0(.din(w_dff_B_mIN3d78w1_0),.dout(w_dff_B_Ye3TTZcF1_0),.clk(gclk));
	jdff dff_B_UHk4d3Nb3_0(.din(w_dff_B_Ye3TTZcF1_0),.dout(w_dff_B_UHk4d3Nb3_0),.clk(gclk));
	jdff dff_B_ipLikkw02_0(.din(w_dff_B_UHk4d3Nb3_0),.dout(w_dff_B_ipLikkw02_0),.clk(gclk));
	jdff dff_B_2WoFnMBh7_0(.din(w_dff_B_ipLikkw02_0),.dout(w_dff_B_2WoFnMBh7_0),.clk(gclk));
	jdff dff_B_QGd9Swlp7_0(.din(w_dff_B_2WoFnMBh7_0),.dout(w_dff_B_QGd9Swlp7_0),.clk(gclk));
	jdff dff_B_Wu4FZKd05_0(.din(w_dff_B_QGd9Swlp7_0),.dout(w_dff_B_Wu4FZKd05_0),.clk(gclk));
	jdff dff_B_Vmrp97804_0(.din(w_dff_B_Wu4FZKd05_0),.dout(w_dff_B_Vmrp97804_0),.clk(gclk));
	jdff dff_B_s9xnr6Pe2_0(.din(w_dff_B_Vmrp97804_0),.dout(w_dff_B_s9xnr6Pe2_0),.clk(gclk));
	jdff dff_B_dyBrehPs0_0(.din(w_dff_B_s9xnr6Pe2_0),.dout(w_dff_B_dyBrehPs0_0),.clk(gclk));
	jdff dff_B_yR7n3T0A8_0(.din(w_dff_B_dyBrehPs0_0),.dout(w_dff_B_yR7n3T0A8_0),.clk(gclk));
	jdff dff_B_zdOnvQdf9_0(.din(w_dff_B_yR7n3T0A8_0),.dout(w_dff_B_zdOnvQdf9_0),.clk(gclk));
	jdff dff_B_HJGwPcYa6_0(.din(w_dff_B_zdOnvQdf9_0),.dout(w_dff_B_HJGwPcYa6_0),.clk(gclk));
	jdff dff_B_aWjKBzaV0_0(.din(w_dff_B_HJGwPcYa6_0),.dout(w_dff_B_aWjKBzaV0_0),.clk(gclk));
	jdff dff_B_N3vJtnMD5_0(.din(w_dff_B_aWjKBzaV0_0),.dout(w_dff_B_N3vJtnMD5_0),.clk(gclk));
	jdff dff_B_jXdoLGA43_0(.din(w_dff_B_N3vJtnMD5_0),.dout(w_dff_B_jXdoLGA43_0),.clk(gclk));
	jdff dff_B_rTapqOOZ4_0(.din(w_dff_B_jXdoLGA43_0),.dout(w_dff_B_rTapqOOZ4_0),.clk(gclk));
	jdff dff_B_IearAhPt4_0(.din(w_dff_B_rTapqOOZ4_0),.dout(w_dff_B_IearAhPt4_0),.clk(gclk));
	jdff dff_B_ac09Q1978_0(.din(w_dff_B_IearAhPt4_0),.dout(w_dff_B_ac09Q1978_0),.clk(gclk));
	jdff dff_B_SbLJRpJj8_0(.din(w_dff_B_ac09Q1978_0),.dout(w_dff_B_SbLJRpJj8_0),.clk(gclk));
	jdff dff_B_aTemLyWC2_0(.din(w_dff_B_SbLJRpJj8_0),.dout(w_dff_B_aTemLyWC2_0),.clk(gclk));
	jdff dff_B_dm1uwraT0_0(.din(w_dff_B_aTemLyWC2_0),.dout(w_dff_B_dm1uwraT0_0),.clk(gclk));
	jdff dff_B_a33z0QD25_0(.din(w_dff_B_dm1uwraT0_0),.dout(w_dff_B_a33z0QD25_0),.clk(gclk));
	jdff dff_B_cmh8g24U9_0(.din(w_dff_B_a33z0QD25_0),.dout(w_dff_B_cmh8g24U9_0),.clk(gclk));
	jdff dff_B_378AIIW14_0(.din(w_dff_B_cmh8g24U9_0),.dout(w_dff_B_378AIIW14_0),.clk(gclk));
	jdff dff_B_qo1I6EWH6_0(.din(w_dff_B_378AIIW14_0),.dout(w_dff_B_qo1I6EWH6_0),.clk(gclk));
	jdff dff_B_pmlBNUhK6_0(.din(w_dff_B_qo1I6EWH6_0),.dout(w_dff_B_pmlBNUhK6_0),.clk(gclk));
	jdff dff_B_DKcVkPuE7_0(.din(w_dff_B_pmlBNUhK6_0),.dout(w_dff_B_DKcVkPuE7_0),.clk(gclk));
	jdff dff_B_EFQSQSk04_0(.din(w_dff_B_DKcVkPuE7_0),.dout(w_dff_B_EFQSQSk04_0),.clk(gclk));
	jdff dff_B_J6XpONsp2_0(.din(w_dff_B_EFQSQSk04_0),.dout(w_dff_B_J6XpONsp2_0),.clk(gclk));
	jdff dff_B_ucZBbHJ59_0(.din(w_dff_B_J6XpONsp2_0),.dout(w_dff_B_ucZBbHJ59_0),.clk(gclk));
	jdff dff_B_HnAuSiv57_0(.din(w_dff_B_ucZBbHJ59_0),.dout(w_dff_B_HnAuSiv57_0),.clk(gclk));
	jdff dff_B_8QqAeA4W4_0(.din(w_dff_B_HnAuSiv57_0),.dout(w_dff_B_8QqAeA4W4_0),.clk(gclk));
	jdff dff_B_zDbyTkJw2_0(.din(w_dff_B_8QqAeA4W4_0),.dout(w_dff_B_zDbyTkJw2_0),.clk(gclk));
	jdff dff_B_HXOPrIN76_0(.din(w_dff_B_zDbyTkJw2_0),.dout(w_dff_B_HXOPrIN76_0),.clk(gclk));
	jdff dff_B_bblFn69R8_0(.din(w_dff_B_HXOPrIN76_0),.dout(w_dff_B_bblFn69R8_0),.clk(gclk));
	jdff dff_B_wpTdDqGr0_0(.din(w_dff_B_bblFn69R8_0),.dout(w_dff_B_wpTdDqGr0_0),.clk(gclk));
	jdff dff_B_GxbX4Cab4_0(.din(w_dff_B_wpTdDqGr0_0),.dout(w_dff_B_GxbX4Cab4_0),.clk(gclk));
	jdff dff_B_VTwEPMHl6_0(.din(w_dff_B_GxbX4Cab4_0),.dout(w_dff_B_VTwEPMHl6_0),.clk(gclk));
	jdff dff_B_gctUakBU0_0(.din(w_dff_B_VTwEPMHl6_0),.dout(w_dff_B_gctUakBU0_0),.clk(gclk));
	jdff dff_B_AgrqmcjW6_0(.din(w_dff_B_gctUakBU0_0),.dout(w_dff_B_AgrqmcjW6_0),.clk(gclk));
	jdff dff_B_tyPWyxTl2_0(.din(w_dff_B_AgrqmcjW6_0),.dout(w_dff_B_tyPWyxTl2_0),.clk(gclk));
	jdff dff_B_syhUo1cF2_0(.din(w_dff_B_tyPWyxTl2_0),.dout(w_dff_B_syhUo1cF2_0),.clk(gclk));
	jdff dff_B_HPMSueB41_0(.din(w_dff_B_syhUo1cF2_0),.dout(w_dff_B_HPMSueB41_0),.clk(gclk));
	jdff dff_B_eNs7Ry896_0(.din(w_dff_B_HPMSueB41_0),.dout(w_dff_B_eNs7Ry896_0),.clk(gclk));
	jdff dff_B_j4lf7bYQ0_0(.din(w_dff_B_eNs7Ry896_0),.dout(w_dff_B_j4lf7bYQ0_0),.clk(gclk));
	jdff dff_B_ycY1IlSU3_0(.din(w_dff_B_j4lf7bYQ0_0),.dout(w_dff_B_ycY1IlSU3_0),.clk(gclk));
	jdff dff_B_FS5rStR61_0(.din(w_dff_B_ycY1IlSU3_0),.dout(w_dff_B_FS5rStR61_0),.clk(gclk));
	jdff dff_B_hBpdjPmG0_0(.din(w_dff_B_FS5rStR61_0),.dout(w_dff_B_hBpdjPmG0_0),.clk(gclk));
	jdff dff_B_hrLVEVHK7_0(.din(w_dff_B_hBpdjPmG0_0),.dout(w_dff_B_hrLVEVHK7_0),.clk(gclk));
	jdff dff_B_nSITv95n9_0(.din(w_dff_B_hrLVEVHK7_0),.dout(w_dff_B_nSITv95n9_0),.clk(gclk));
	jdff dff_B_8CZYt4qo7_0(.din(w_dff_B_nSITv95n9_0),.dout(w_dff_B_8CZYt4qo7_0),.clk(gclk));
	jdff dff_B_at2HwvLi3_0(.din(w_dff_B_8CZYt4qo7_0),.dout(w_dff_B_at2HwvLi3_0),.clk(gclk));
	jdff dff_B_9ygDQVEG6_0(.din(w_dff_B_at2HwvLi3_0),.dout(w_dff_B_9ygDQVEG6_0),.clk(gclk));
	jdff dff_B_fZS1BtOV9_0(.din(w_dff_B_9ygDQVEG6_0),.dout(w_dff_B_fZS1BtOV9_0),.clk(gclk));
	jdff dff_B_xELxgy789_0(.din(w_dff_B_fZS1BtOV9_0),.dout(w_dff_B_xELxgy789_0),.clk(gclk));
	jdff dff_B_U09uoXR96_0(.din(w_dff_B_xELxgy789_0),.dout(w_dff_B_U09uoXR96_0),.clk(gclk));
	jdff dff_B_ccBwl2gZ4_0(.din(w_dff_B_U09uoXR96_0),.dout(w_dff_B_ccBwl2gZ4_0),.clk(gclk));
	jdff dff_B_ayx3pwgB2_0(.din(w_dff_B_ccBwl2gZ4_0),.dout(w_dff_B_ayx3pwgB2_0),.clk(gclk));
	jdff dff_B_YzWvd2OB0_0(.din(w_dff_B_ayx3pwgB2_0),.dout(w_dff_B_YzWvd2OB0_0),.clk(gclk));
	jdff dff_B_9famPQo49_0(.din(w_dff_B_YzWvd2OB0_0),.dout(w_dff_B_9famPQo49_0),.clk(gclk));
	jdff dff_B_5lZb1mgG9_0(.din(w_dff_B_9famPQo49_0),.dout(w_dff_B_5lZb1mgG9_0),.clk(gclk));
	jdff dff_B_stvrphk09_0(.din(w_dff_B_5lZb1mgG9_0),.dout(w_dff_B_stvrphk09_0),.clk(gclk));
	jdff dff_B_17cXq4X46_0(.din(w_dff_B_stvrphk09_0),.dout(w_dff_B_17cXq4X46_0),.clk(gclk));
	jdff dff_B_7vIoF1Qc0_0(.din(w_dff_B_17cXq4X46_0),.dout(w_dff_B_7vIoF1Qc0_0),.clk(gclk));
	jdff dff_B_PknXh2HB1_0(.din(w_dff_B_7vIoF1Qc0_0),.dout(w_dff_B_PknXh2HB1_0),.clk(gclk));
	jdff dff_B_mVbVs9gG9_0(.din(w_dff_B_PknXh2HB1_0),.dout(w_dff_B_mVbVs9gG9_0),.clk(gclk));
	jdff dff_B_05A0b1yf0_0(.din(w_dff_B_mVbVs9gG9_0),.dout(w_dff_B_05A0b1yf0_0),.clk(gclk));
	jdff dff_B_GW1rbx2z6_0(.din(w_dff_B_05A0b1yf0_0),.dout(w_dff_B_GW1rbx2z6_0),.clk(gclk));
	jdff dff_B_fAmRyzbQ8_0(.din(w_dff_B_GW1rbx2z6_0),.dout(w_dff_B_fAmRyzbQ8_0),.clk(gclk));
	jdff dff_B_OWtdytaD9_0(.din(w_dff_B_fAmRyzbQ8_0),.dout(w_dff_B_OWtdytaD9_0),.clk(gclk));
	jdff dff_B_FuTTeeuX1_0(.din(w_dff_B_OWtdytaD9_0),.dout(w_dff_B_FuTTeeuX1_0),.clk(gclk));
	jdff dff_B_JFml0BBk6_0(.din(w_dff_B_FuTTeeuX1_0),.dout(w_dff_B_JFml0BBk6_0),.clk(gclk));
	jdff dff_B_Q8dQkKOd8_0(.din(w_dff_B_JFml0BBk6_0),.dout(w_dff_B_Q8dQkKOd8_0),.clk(gclk));
	jdff dff_B_OKNTs6kD0_0(.din(w_dff_B_Q8dQkKOd8_0),.dout(w_dff_B_OKNTs6kD0_0),.clk(gclk));
	jdff dff_B_frAbasL66_0(.din(w_dff_B_OKNTs6kD0_0),.dout(w_dff_B_frAbasL66_0),.clk(gclk));
	jdff dff_B_cX2qw0Z04_0(.din(w_dff_B_frAbasL66_0),.dout(w_dff_B_cX2qw0Z04_0),.clk(gclk));
	jdff dff_B_tlsd6gJ52_0(.din(w_dff_B_cX2qw0Z04_0),.dout(w_dff_B_tlsd6gJ52_0),.clk(gclk));
	jdff dff_B_9jvOhias7_0(.din(w_dff_B_tlsd6gJ52_0),.dout(w_dff_B_9jvOhias7_0),.clk(gclk));
	jdff dff_B_CDenmHyS5_0(.din(w_dff_B_9jvOhias7_0),.dout(w_dff_B_CDenmHyS5_0),.clk(gclk));
	jdff dff_B_wNaBnSyQ9_0(.din(w_dff_B_CDenmHyS5_0),.dout(w_dff_B_wNaBnSyQ9_0),.clk(gclk));
	jdff dff_B_Dw3ibZ2E1_0(.din(w_dff_B_wNaBnSyQ9_0),.dout(w_dff_B_Dw3ibZ2E1_0),.clk(gclk));
	jdff dff_B_ztDSc3fz3_0(.din(w_dff_B_Dw3ibZ2E1_0),.dout(w_dff_B_ztDSc3fz3_0),.clk(gclk));
	jdff dff_B_GNKytxFO3_0(.din(w_dff_B_ztDSc3fz3_0),.dout(w_dff_B_GNKytxFO3_0),.clk(gclk));
	jdff dff_B_AUYca1hl2_0(.din(w_dff_B_GNKytxFO3_0),.dout(w_dff_B_AUYca1hl2_0),.clk(gclk));
	jdff dff_B_WifhNf3n2_0(.din(w_dff_B_AUYca1hl2_0),.dout(w_dff_B_WifhNf3n2_0),.clk(gclk));
	jdff dff_B_8t38Yj9U5_0(.din(w_dff_B_WifhNf3n2_0),.dout(w_dff_B_8t38Yj9U5_0),.clk(gclk));
	jdff dff_B_whkEqGju9_0(.din(w_dff_B_8t38Yj9U5_0),.dout(w_dff_B_whkEqGju9_0),.clk(gclk));
	jdff dff_B_1m4hZpYQ7_0(.din(w_dff_B_whkEqGju9_0),.dout(w_dff_B_1m4hZpYQ7_0),.clk(gclk));
	jdff dff_B_r0fBw0CL6_0(.din(w_dff_B_1m4hZpYQ7_0),.dout(w_dff_B_r0fBw0CL6_0),.clk(gclk));
	jdff dff_B_dFlcaupd5_0(.din(w_dff_B_r0fBw0CL6_0),.dout(w_dff_B_dFlcaupd5_0),.clk(gclk));
	jdff dff_B_OmEewm5z6_0(.din(w_dff_B_dFlcaupd5_0),.dout(w_dff_B_OmEewm5z6_0),.clk(gclk));
	jdff dff_B_JUUjm9XO7_1(.din(n1014),.dout(w_dff_B_JUUjm9XO7_1),.clk(gclk));
	jdff dff_B_ugGZOQGc4_1(.din(w_dff_B_JUUjm9XO7_1),.dout(w_dff_B_ugGZOQGc4_1),.clk(gclk));
	jdff dff_B_aaS0NVKT3_1(.din(w_dff_B_ugGZOQGc4_1),.dout(w_dff_B_aaS0NVKT3_1),.clk(gclk));
	jdff dff_B_Mag5RAyv4_1(.din(w_dff_B_aaS0NVKT3_1),.dout(w_dff_B_Mag5RAyv4_1),.clk(gclk));
	jdff dff_B_nvlWEInm8_1(.din(w_dff_B_Mag5RAyv4_1),.dout(w_dff_B_nvlWEInm8_1),.clk(gclk));
	jdff dff_B_PyDChZAP3_1(.din(w_dff_B_nvlWEInm8_1),.dout(w_dff_B_PyDChZAP3_1),.clk(gclk));
	jdff dff_B_bTtMVvBi8_1(.din(w_dff_B_PyDChZAP3_1),.dout(w_dff_B_bTtMVvBi8_1),.clk(gclk));
	jdff dff_B_6ipDwSkz7_1(.din(w_dff_B_bTtMVvBi8_1),.dout(w_dff_B_6ipDwSkz7_1),.clk(gclk));
	jdff dff_B_fvOamn8j9_1(.din(w_dff_B_6ipDwSkz7_1),.dout(w_dff_B_fvOamn8j9_1),.clk(gclk));
	jdff dff_B_W2BfAWBI3_1(.din(w_dff_B_fvOamn8j9_1),.dout(w_dff_B_W2BfAWBI3_1),.clk(gclk));
	jdff dff_B_ZDPbW5Ud3_1(.din(w_dff_B_W2BfAWBI3_1),.dout(w_dff_B_ZDPbW5Ud3_1),.clk(gclk));
	jdff dff_B_66A2Y7jx4_1(.din(w_dff_B_ZDPbW5Ud3_1),.dout(w_dff_B_66A2Y7jx4_1),.clk(gclk));
	jdff dff_B_rv9Pg3UY2_1(.din(w_dff_B_66A2Y7jx4_1),.dout(w_dff_B_rv9Pg3UY2_1),.clk(gclk));
	jdff dff_B_9EsukJjn0_1(.din(w_dff_B_rv9Pg3UY2_1),.dout(w_dff_B_9EsukJjn0_1),.clk(gclk));
	jdff dff_B_4NZxd1G13_1(.din(w_dff_B_9EsukJjn0_1),.dout(w_dff_B_4NZxd1G13_1),.clk(gclk));
	jdff dff_B_9ILGoqVG4_1(.din(w_dff_B_4NZxd1G13_1),.dout(w_dff_B_9ILGoqVG4_1),.clk(gclk));
	jdff dff_B_mKx1xcwS8_1(.din(w_dff_B_9ILGoqVG4_1),.dout(w_dff_B_mKx1xcwS8_1),.clk(gclk));
	jdff dff_B_XG1AWsmw1_1(.din(w_dff_B_mKx1xcwS8_1),.dout(w_dff_B_XG1AWsmw1_1),.clk(gclk));
	jdff dff_B_AXlW9Mng1_1(.din(w_dff_B_XG1AWsmw1_1),.dout(w_dff_B_AXlW9Mng1_1),.clk(gclk));
	jdff dff_B_0DBCNyFy1_1(.din(w_dff_B_AXlW9Mng1_1),.dout(w_dff_B_0DBCNyFy1_1),.clk(gclk));
	jdff dff_B_pbbm2fMz0_1(.din(w_dff_B_0DBCNyFy1_1),.dout(w_dff_B_pbbm2fMz0_1),.clk(gclk));
	jdff dff_B_5WUfzSRl8_1(.din(w_dff_B_pbbm2fMz0_1),.dout(w_dff_B_5WUfzSRl8_1),.clk(gclk));
	jdff dff_B_Ajc4k1FC6_1(.din(w_dff_B_5WUfzSRl8_1),.dout(w_dff_B_Ajc4k1FC6_1),.clk(gclk));
	jdff dff_B_NMq6UkGZ4_1(.din(w_dff_B_Ajc4k1FC6_1),.dout(w_dff_B_NMq6UkGZ4_1),.clk(gclk));
	jdff dff_B_ruVKIaDw4_1(.din(w_dff_B_NMq6UkGZ4_1),.dout(w_dff_B_ruVKIaDw4_1),.clk(gclk));
	jdff dff_B_tmlXTsKA8_1(.din(w_dff_B_ruVKIaDw4_1),.dout(w_dff_B_tmlXTsKA8_1),.clk(gclk));
	jdff dff_B_zEGyTuKT3_1(.din(w_dff_B_tmlXTsKA8_1),.dout(w_dff_B_zEGyTuKT3_1),.clk(gclk));
	jdff dff_B_k3xLNKhO6_1(.din(w_dff_B_zEGyTuKT3_1),.dout(w_dff_B_k3xLNKhO6_1),.clk(gclk));
	jdff dff_B_5zoKq7im8_1(.din(w_dff_B_k3xLNKhO6_1),.dout(w_dff_B_5zoKq7im8_1),.clk(gclk));
	jdff dff_B_K0pL3mhG2_1(.din(w_dff_B_5zoKq7im8_1),.dout(w_dff_B_K0pL3mhG2_1),.clk(gclk));
	jdff dff_B_1Hy5iJpa9_1(.din(w_dff_B_K0pL3mhG2_1),.dout(w_dff_B_1Hy5iJpa9_1),.clk(gclk));
	jdff dff_B_rf3tRyeL7_1(.din(w_dff_B_1Hy5iJpa9_1),.dout(w_dff_B_rf3tRyeL7_1),.clk(gclk));
	jdff dff_B_JJx3DrRV3_1(.din(w_dff_B_rf3tRyeL7_1),.dout(w_dff_B_JJx3DrRV3_1),.clk(gclk));
	jdff dff_B_hFXxEyka4_1(.din(w_dff_B_JJx3DrRV3_1),.dout(w_dff_B_hFXxEyka4_1),.clk(gclk));
	jdff dff_B_qLlHQfSq7_1(.din(w_dff_B_hFXxEyka4_1),.dout(w_dff_B_qLlHQfSq7_1),.clk(gclk));
	jdff dff_B_BLywJjcP4_1(.din(w_dff_B_qLlHQfSq7_1),.dout(w_dff_B_BLywJjcP4_1),.clk(gclk));
	jdff dff_B_g31FVAto9_1(.din(w_dff_B_BLywJjcP4_1),.dout(w_dff_B_g31FVAto9_1),.clk(gclk));
	jdff dff_B_KKO4CKx77_1(.din(w_dff_B_g31FVAto9_1),.dout(w_dff_B_KKO4CKx77_1),.clk(gclk));
	jdff dff_B_n9wBg8Et9_1(.din(w_dff_B_KKO4CKx77_1),.dout(w_dff_B_n9wBg8Et9_1),.clk(gclk));
	jdff dff_B_SIJUhVml3_1(.din(w_dff_B_n9wBg8Et9_1),.dout(w_dff_B_SIJUhVml3_1),.clk(gclk));
	jdff dff_B_YjRPGwob9_1(.din(w_dff_B_SIJUhVml3_1),.dout(w_dff_B_YjRPGwob9_1),.clk(gclk));
	jdff dff_B_tdYXr8Ue5_1(.din(w_dff_B_YjRPGwob9_1),.dout(w_dff_B_tdYXr8Ue5_1),.clk(gclk));
	jdff dff_B_2z6Xm6jk5_1(.din(w_dff_B_tdYXr8Ue5_1),.dout(w_dff_B_2z6Xm6jk5_1),.clk(gclk));
	jdff dff_B_g8eVitQw0_1(.din(w_dff_B_2z6Xm6jk5_1),.dout(w_dff_B_g8eVitQw0_1),.clk(gclk));
	jdff dff_B_vTYPfvl81_1(.din(w_dff_B_g8eVitQw0_1),.dout(w_dff_B_vTYPfvl81_1),.clk(gclk));
	jdff dff_B_UhU2nAds0_1(.din(w_dff_B_vTYPfvl81_1),.dout(w_dff_B_UhU2nAds0_1),.clk(gclk));
	jdff dff_B_zUPJRTCT3_1(.din(w_dff_B_UhU2nAds0_1),.dout(w_dff_B_zUPJRTCT3_1),.clk(gclk));
	jdff dff_B_jBODE7sf7_1(.din(w_dff_B_zUPJRTCT3_1),.dout(w_dff_B_jBODE7sf7_1),.clk(gclk));
	jdff dff_B_mvsYVhxU3_1(.din(w_dff_B_jBODE7sf7_1),.dout(w_dff_B_mvsYVhxU3_1),.clk(gclk));
	jdff dff_B_VewwZZgh6_1(.din(w_dff_B_mvsYVhxU3_1),.dout(w_dff_B_VewwZZgh6_1),.clk(gclk));
	jdff dff_B_tdA69xAC3_1(.din(w_dff_B_VewwZZgh6_1),.dout(w_dff_B_tdA69xAC3_1),.clk(gclk));
	jdff dff_B_TLG4aLnL8_1(.din(w_dff_B_tdA69xAC3_1),.dout(w_dff_B_TLG4aLnL8_1),.clk(gclk));
	jdff dff_B_kdqW6lY40_1(.din(w_dff_B_TLG4aLnL8_1),.dout(w_dff_B_kdqW6lY40_1),.clk(gclk));
	jdff dff_B_tqVtFNve8_1(.din(w_dff_B_kdqW6lY40_1),.dout(w_dff_B_tqVtFNve8_1),.clk(gclk));
	jdff dff_B_Rw87Cy3u6_1(.din(w_dff_B_tqVtFNve8_1),.dout(w_dff_B_Rw87Cy3u6_1),.clk(gclk));
	jdff dff_B_xRC3sDTn0_1(.din(w_dff_B_Rw87Cy3u6_1),.dout(w_dff_B_xRC3sDTn0_1),.clk(gclk));
	jdff dff_B_SqEdrAAx5_1(.din(w_dff_B_xRC3sDTn0_1),.dout(w_dff_B_SqEdrAAx5_1),.clk(gclk));
	jdff dff_B_m3C534ZW5_1(.din(w_dff_B_SqEdrAAx5_1),.dout(w_dff_B_m3C534ZW5_1),.clk(gclk));
	jdff dff_B_ewtK5mJ97_1(.din(w_dff_B_m3C534ZW5_1),.dout(w_dff_B_ewtK5mJ97_1),.clk(gclk));
	jdff dff_B_2GYbysjL2_1(.din(w_dff_B_ewtK5mJ97_1),.dout(w_dff_B_2GYbysjL2_1),.clk(gclk));
	jdff dff_B_uJXetQbI6_1(.din(w_dff_B_2GYbysjL2_1),.dout(w_dff_B_uJXetQbI6_1),.clk(gclk));
	jdff dff_B_5p2Uwr378_1(.din(w_dff_B_uJXetQbI6_1),.dout(w_dff_B_5p2Uwr378_1),.clk(gclk));
	jdff dff_B_hSYqCOIf6_1(.din(w_dff_B_5p2Uwr378_1),.dout(w_dff_B_hSYqCOIf6_1),.clk(gclk));
	jdff dff_B_pdGh6DDR5_1(.din(w_dff_B_hSYqCOIf6_1),.dout(w_dff_B_pdGh6DDR5_1),.clk(gclk));
	jdff dff_B_FU5WNjug3_1(.din(w_dff_B_pdGh6DDR5_1),.dout(w_dff_B_FU5WNjug3_1),.clk(gclk));
	jdff dff_B_KeLjHwOo0_1(.din(w_dff_B_FU5WNjug3_1),.dout(w_dff_B_KeLjHwOo0_1),.clk(gclk));
	jdff dff_B_E7WElCnm2_1(.din(w_dff_B_KeLjHwOo0_1),.dout(w_dff_B_E7WElCnm2_1),.clk(gclk));
	jdff dff_B_iG6VsE8q8_1(.din(w_dff_B_E7WElCnm2_1),.dout(w_dff_B_iG6VsE8q8_1),.clk(gclk));
	jdff dff_B_ttvzSkoR7_1(.din(w_dff_B_iG6VsE8q8_1),.dout(w_dff_B_ttvzSkoR7_1),.clk(gclk));
	jdff dff_B_yIVzYWdx2_1(.din(w_dff_B_ttvzSkoR7_1),.dout(w_dff_B_yIVzYWdx2_1),.clk(gclk));
	jdff dff_B_iX6WM2vv0_1(.din(w_dff_B_yIVzYWdx2_1),.dout(w_dff_B_iX6WM2vv0_1),.clk(gclk));
	jdff dff_B_k2zSO25V4_1(.din(w_dff_B_iX6WM2vv0_1),.dout(w_dff_B_k2zSO25V4_1),.clk(gclk));
	jdff dff_B_kQ2MLCEU3_1(.din(w_dff_B_k2zSO25V4_1),.dout(w_dff_B_kQ2MLCEU3_1),.clk(gclk));
	jdff dff_B_vaP66fZx3_1(.din(w_dff_B_kQ2MLCEU3_1),.dout(w_dff_B_vaP66fZx3_1),.clk(gclk));
	jdff dff_B_rXWxyiOV1_1(.din(w_dff_B_vaP66fZx3_1),.dout(w_dff_B_rXWxyiOV1_1),.clk(gclk));
	jdff dff_B_UcXmYYVp5_1(.din(w_dff_B_rXWxyiOV1_1),.dout(w_dff_B_UcXmYYVp5_1),.clk(gclk));
	jdff dff_B_fRNd6gK80_1(.din(w_dff_B_UcXmYYVp5_1),.dout(w_dff_B_fRNd6gK80_1),.clk(gclk));
	jdff dff_B_knJcnDia6_1(.din(w_dff_B_fRNd6gK80_1),.dout(w_dff_B_knJcnDia6_1),.clk(gclk));
	jdff dff_B_cBgUkfGc0_1(.din(w_dff_B_knJcnDia6_1),.dout(w_dff_B_cBgUkfGc0_1),.clk(gclk));
	jdff dff_B_GlqGkDHz4_1(.din(w_dff_B_cBgUkfGc0_1),.dout(w_dff_B_GlqGkDHz4_1),.clk(gclk));
	jdff dff_B_3Kd18oPV1_1(.din(w_dff_B_GlqGkDHz4_1),.dout(w_dff_B_3Kd18oPV1_1),.clk(gclk));
	jdff dff_B_cJyLxk779_1(.din(w_dff_B_3Kd18oPV1_1),.dout(w_dff_B_cJyLxk779_1),.clk(gclk));
	jdff dff_B_8IXRVP938_1(.din(w_dff_B_cJyLxk779_1),.dout(w_dff_B_8IXRVP938_1),.clk(gclk));
	jdff dff_B_83sdgtFi5_1(.din(w_dff_B_8IXRVP938_1),.dout(w_dff_B_83sdgtFi5_1),.clk(gclk));
	jdff dff_B_2mSg8kJD8_1(.din(w_dff_B_83sdgtFi5_1),.dout(w_dff_B_2mSg8kJD8_1),.clk(gclk));
	jdff dff_B_ItvNy3gS8_1(.din(w_dff_B_2mSg8kJD8_1),.dout(w_dff_B_ItvNy3gS8_1),.clk(gclk));
	jdff dff_B_zLaIRpRP6_1(.din(w_dff_B_ItvNy3gS8_1),.dout(w_dff_B_zLaIRpRP6_1),.clk(gclk));
	jdff dff_B_RZjEuioS1_1(.din(w_dff_B_zLaIRpRP6_1),.dout(w_dff_B_RZjEuioS1_1),.clk(gclk));
	jdff dff_B_58PEEVGP1_1(.din(w_dff_B_RZjEuioS1_1),.dout(w_dff_B_58PEEVGP1_1),.clk(gclk));
	jdff dff_B_cVjkXz2t7_1(.din(w_dff_B_58PEEVGP1_1),.dout(w_dff_B_cVjkXz2t7_1),.clk(gclk));
	jdff dff_B_dyNkmlfy8_1(.din(w_dff_B_cVjkXz2t7_1),.dout(w_dff_B_dyNkmlfy8_1),.clk(gclk));
	jdff dff_B_3oPKDMJ41_1(.din(w_dff_B_dyNkmlfy8_1),.dout(w_dff_B_3oPKDMJ41_1),.clk(gclk));
	jdff dff_B_cj7yehJr8_1(.din(w_dff_B_3oPKDMJ41_1),.dout(w_dff_B_cj7yehJr8_1),.clk(gclk));
	jdff dff_B_NHEvEhQa4_1(.din(w_dff_B_cj7yehJr8_1),.dout(w_dff_B_NHEvEhQa4_1),.clk(gclk));
	jdff dff_B_72IqebV26_1(.din(w_dff_B_NHEvEhQa4_1),.dout(w_dff_B_72IqebV26_1),.clk(gclk));
	jdff dff_B_ETzYWIxJ7_1(.din(w_dff_B_72IqebV26_1),.dout(w_dff_B_ETzYWIxJ7_1),.clk(gclk));
	jdff dff_B_BErVn2rC2_1(.din(w_dff_B_ETzYWIxJ7_1),.dout(w_dff_B_BErVn2rC2_1),.clk(gclk));
	jdff dff_B_LQNZ0gjG7_1(.din(w_dff_B_BErVn2rC2_1),.dout(w_dff_B_LQNZ0gjG7_1),.clk(gclk));
	jdff dff_B_bLOwMUpj1_1(.din(w_dff_B_LQNZ0gjG7_1),.dout(w_dff_B_bLOwMUpj1_1),.clk(gclk));
	jdff dff_B_c7EIYxgT3_1(.din(w_dff_B_bLOwMUpj1_1),.dout(w_dff_B_c7EIYxgT3_1),.clk(gclk));
	jdff dff_B_R7FpmBCw1_1(.din(w_dff_B_c7EIYxgT3_1),.dout(w_dff_B_R7FpmBCw1_1),.clk(gclk));
	jdff dff_B_3dT33HA32_1(.din(w_dff_B_R7FpmBCw1_1),.dout(w_dff_B_3dT33HA32_1),.clk(gclk));
	jdff dff_B_w0HbWKII0_1(.din(w_dff_B_3dT33HA32_1),.dout(w_dff_B_w0HbWKII0_1),.clk(gclk));
	jdff dff_B_r6KoXOnJ3_1(.din(w_dff_B_w0HbWKII0_1),.dout(w_dff_B_r6KoXOnJ3_1),.clk(gclk));
	jdff dff_B_opUbMGB49_1(.din(w_dff_B_r6KoXOnJ3_1),.dout(w_dff_B_opUbMGB49_1),.clk(gclk));
	jdff dff_B_sopoYNE76_0(.din(n1015),.dout(w_dff_B_sopoYNE76_0),.clk(gclk));
	jdff dff_B_0eGGHMlu3_0(.din(w_dff_B_sopoYNE76_0),.dout(w_dff_B_0eGGHMlu3_0),.clk(gclk));
	jdff dff_B_ZR57yI1Z8_0(.din(w_dff_B_0eGGHMlu3_0),.dout(w_dff_B_ZR57yI1Z8_0),.clk(gclk));
	jdff dff_B_gm6BWLov8_0(.din(w_dff_B_ZR57yI1Z8_0),.dout(w_dff_B_gm6BWLov8_0),.clk(gclk));
	jdff dff_B_4pl9aWMf4_0(.din(w_dff_B_gm6BWLov8_0),.dout(w_dff_B_4pl9aWMf4_0),.clk(gclk));
	jdff dff_B_leq9d4qL3_0(.din(w_dff_B_4pl9aWMf4_0),.dout(w_dff_B_leq9d4qL3_0),.clk(gclk));
	jdff dff_B_duTWINYO1_0(.din(w_dff_B_leq9d4qL3_0),.dout(w_dff_B_duTWINYO1_0),.clk(gclk));
	jdff dff_B_vB43oCBE1_0(.din(w_dff_B_duTWINYO1_0),.dout(w_dff_B_vB43oCBE1_0),.clk(gclk));
	jdff dff_B_MatlSzIi3_0(.din(w_dff_B_vB43oCBE1_0),.dout(w_dff_B_MatlSzIi3_0),.clk(gclk));
	jdff dff_B_iclNGsXo1_0(.din(w_dff_B_MatlSzIi3_0),.dout(w_dff_B_iclNGsXo1_0),.clk(gclk));
	jdff dff_B_aomv0Fqh8_0(.din(w_dff_B_iclNGsXo1_0),.dout(w_dff_B_aomv0Fqh8_0),.clk(gclk));
	jdff dff_B_fRw8MDn73_0(.din(w_dff_B_aomv0Fqh8_0),.dout(w_dff_B_fRw8MDn73_0),.clk(gclk));
	jdff dff_B_wsODJM8E6_0(.din(w_dff_B_fRw8MDn73_0),.dout(w_dff_B_wsODJM8E6_0),.clk(gclk));
	jdff dff_B_zcawso2S7_0(.din(w_dff_B_wsODJM8E6_0),.dout(w_dff_B_zcawso2S7_0),.clk(gclk));
	jdff dff_B_nNxa7va32_0(.din(w_dff_B_zcawso2S7_0),.dout(w_dff_B_nNxa7va32_0),.clk(gclk));
	jdff dff_B_JXSP59g56_0(.din(w_dff_B_nNxa7va32_0),.dout(w_dff_B_JXSP59g56_0),.clk(gclk));
	jdff dff_B_zr89SJry3_0(.din(w_dff_B_JXSP59g56_0),.dout(w_dff_B_zr89SJry3_0),.clk(gclk));
	jdff dff_B_anzB9ocb7_0(.din(w_dff_B_zr89SJry3_0),.dout(w_dff_B_anzB9ocb7_0),.clk(gclk));
	jdff dff_B_0Ha5SysI8_0(.din(w_dff_B_anzB9ocb7_0),.dout(w_dff_B_0Ha5SysI8_0),.clk(gclk));
	jdff dff_B_lai9bFW44_0(.din(w_dff_B_0Ha5SysI8_0),.dout(w_dff_B_lai9bFW44_0),.clk(gclk));
	jdff dff_B_Bcn4AlFl6_0(.din(w_dff_B_lai9bFW44_0),.dout(w_dff_B_Bcn4AlFl6_0),.clk(gclk));
	jdff dff_B_qFwM2U1V6_0(.din(w_dff_B_Bcn4AlFl6_0),.dout(w_dff_B_qFwM2U1V6_0),.clk(gclk));
	jdff dff_B_1KrcOf3k7_0(.din(w_dff_B_qFwM2U1V6_0),.dout(w_dff_B_1KrcOf3k7_0),.clk(gclk));
	jdff dff_B_ubAMaq8Q2_0(.din(w_dff_B_1KrcOf3k7_0),.dout(w_dff_B_ubAMaq8Q2_0),.clk(gclk));
	jdff dff_B_QmfOAmNk3_0(.din(w_dff_B_ubAMaq8Q2_0),.dout(w_dff_B_QmfOAmNk3_0),.clk(gclk));
	jdff dff_B_LdaOF7WW8_0(.din(w_dff_B_QmfOAmNk3_0),.dout(w_dff_B_LdaOF7WW8_0),.clk(gclk));
	jdff dff_B_nGiKIEOw8_0(.din(w_dff_B_LdaOF7WW8_0),.dout(w_dff_B_nGiKIEOw8_0),.clk(gclk));
	jdff dff_B_NjEYtfRS3_0(.din(w_dff_B_nGiKIEOw8_0),.dout(w_dff_B_NjEYtfRS3_0),.clk(gclk));
	jdff dff_B_s7NG6gVf6_0(.din(w_dff_B_NjEYtfRS3_0),.dout(w_dff_B_s7NG6gVf6_0),.clk(gclk));
	jdff dff_B_joyQhANH8_0(.din(w_dff_B_s7NG6gVf6_0),.dout(w_dff_B_joyQhANH8_0),.clk(gclk));
	jdff dff_B_MlBXG8Bf0_0(.din(w_dff_B_joyQhANH8_0),.dout(w_dff_B_MlBXG8Bf0_0),.clk(gclk));
	jdff dff_B_sALFBYPA4_0(.din(w_dff_B_MlBXG8Bf0_0),.dout(w_dff_B_sALFBYPA4_0),.clk(gclk));
	jdff dff_B_4l5xCi2h6_0(.din(w_dff_B_sALFBYPA4_0),.dout(w_dff_B_4l5xCi2h6_0),.clk(gclk));
	jdff dff_B_E4ajtg692_0(.din(w_dff_B_4l5xCi2h6_0),.dout(w_dff_B_E4ajtg692_0),.clk(gclk));
	jdff dff_B_Mv7yniZq2_0(.din(w_dff_B_E4ajtg692_0),.dout(w_dff_B_Mv7yniZq2_0),.clk(gclk));
	jdff dff_B_4hxiN5Og8_0(.din(w_dff_B_Mv7yniZq2_0),.dout(w_dff_B_4hxiN5Og8_0),.clk(gclk));
	jdff dff_B_Odmd7uzu3_0(.din(w_dff_B_4hxiN5Og8_0),.dout(w_dff_B_Odmd7uzu3_0),.clk(gclk));
	jdff dff_B_YLWAYSjY3_0(.din(w_dff_B_Odmd7uzu3_0),.dout(w_dff_B_YLWAYSjY3_0),.clk(gclk));
	jdff dff_B_sRipMn8T2_0(.din(w_dff_B_YLWAYSjY3_0),.dout(w_dff_B_sRipMn8T2_0),.clk(gclk));
	jdff dff_B_vg4Gf6lg3_0(.din(w_dff_B_sRipMn8T2_0),.dout(w_dff_B_vg4Gf6lg3_0),.clk(gclk));
	jdff dff_B_k3pfXuHF7_0(.din(w_dff_B_vg4Gf6lg3_0),.dout(w_dff_B_k3pfXuHF7_0),.clk(gclk));
	jdff dff_B_eXGVUCuG5_0(.din(w_dff_B_k3pfXuHF7_0),.dout(w_dff_B_eXGVUCuG5_0),.clk(gclk));
	jdff dff_B_33YCekoC2_0(.din(w_dff_B_eXGVUCuG5_0),.dout(w_dff_B_33YCekoC2_0),.clk(gclk));
	jdff dff_B_87DN9wnS0_0(.din(w_dff_B_33YCekoC2_0),.dout(w_dff_B_87DN9wnS0_0),.clk(gclk));
	jdff dff_B_0baUcS5p7_0(.din(w_dff_B_87DN9wnS0_0),.dout(w_dff_B_0baUcS5p7_0),.clk(gclk));
	jdff dff_B_0nZm7Sdy8_0(.din(w_dff_B_0baUcS5p7_0),.dout(w_dff_B_0nZm7Sdy8_0),.clk(gclk));
	jdff dff_B_mk7sEWke6_0(.din(w_dff_B_0nZm7Sdy8_0),.dout(w_dff_B_mk7sEWke6_0),.clk(gclk));
	jdff dff_B_fIYAB21S1_0(.din(w_dff_B_mk7sEWke6_0),.dout(w_dff_B_fIYAB21S1_0),.clk(gclk));
	jdff dff_B_nD5jHmAZ0_0(.din(w_dff_B_fIYAB21S1_0),.dout(w_dff_B_nD5jHmAZ0_0),.clk(gclk));
	jdff dff_B_u3xd9PFr8_0(.din(w_dff_B_nD5jHmAZ0_0),.dout(w_dff_B_u3xd9PFr8_0),.clk(gclk));
	jdff dff_B_lH8XCHC72_0(.din(w_dff_B_u3xd9PFr8_0),.dout(w_dff_B_lH8XCHC72_0),.clk(gclk));
	jdff dff_B_DbuqCntg1_0(.din(w_dff_B_lH8XCHC72_0),.dout(w_dff_B_DbuqCntg1_0),.clk(gclk));
	jdff dff_B_3OlBQqIe5_0(.din(w_dff_B_DbuqCntg1_0),.dout(w_dff_B_3OlBQqIe5_0),.clk(gclk));
	jdff dff_B_QjbMqjXH9_0(.din(w_dff_B_3OlBQqIe5_0),.dout(w_dff_B_QjbMqjXH9_0),.clk(gclk));
	jdff dff_B_WMDwby1R5_0(.din(w_dff_B_QjbMqjXH9_0),.dout(w_dff_B_WMDwby1R5_0),.clk(gclk));
	jdff dff_B_Mfct0s1v0_0(.din(w_dff_B_WMDwby1R5_0),.dout(w_dff_B_Mfct0s1v0_0),.clk(gclk));
	jdff dff_B_6DT5gzTT1_0(.din(w_dff_B_Mfct0s1v0_0),.dout(w_dff_B_6DT5gzTT1_0),.clk(gclk));
	jdff dff_B_L4UskE3C7_0(.din(w_dff_B_6DT5gzTT1_0),.dout(w_dff_B_L4UskE3C7_0),.clk(gclk));
	jdff dff_B_bp8t7ZE46_0(.din(w_dff_B_L4UskE3C7_0),.dout(w_dff_B_bp8t7ZE46_0),.clk(gclk));
	jdff dff_B_17eGOwd79_0(.din(w_dff_B_bp8t7ZE46_0),.dout(w_dff_B_17eGOwd79_0),.clk(gclk));
	jdff dff_B_Kmw9BlMH2_0(.din(w_dff_B_17eGOwd79_0),.dout(w_dff_B_Kmw9BlMH2_0),.clk(gclk));
	jdff dff_B_aLWfetc56_0(.din(w_dff_B_Kmw9BlMH2_0),.dout(w_dff_B_aLWfetc56_0),.clk(gclk));
	jdff dff_B_A0xtEKIQ1_0(.din(w_dff_B_aLWfetc56_0),.dout(w_dff_B_A0xtEKIQ1_0),.clk(gclk));
	jdff dff_B_b5VN4p2H0_0(.din(w_dff_B_A0xtEKIQ1_0),.dout(w_dff_B_b5VN4p2H0_0),.clk(gclk));
	jdff dff_B_B2RodtiT9_0(.din(w_dff_B_b5VN4p2H0_0),.dout(w_dff_B_B2RodtiT9_0),.clk(gclk));
	jdff dff_B_l0O7bCit6_0(.din(w_dff_B_B2RodtiT9_0),.dout(w_dff_B_l0O7bCit6_0),.clk(gclk));
	jdff dff_B_fzHBgx1X3_0(.din(w_dff_B_l0O7bCit6_0),.dout(w_dff_B_fzHBgx1X3_0),.clk(gclk));
	jdff dff_B_u8OwdW1U7_0(.din(w_dff_B_fzHBgx1X3_0),.dout(w_dff_B_u8OwdW1U7_0),.clk(gclk));
	jdff dff_B_l6H5NuBV9_0(.din(w_dff_B_u8OwdW1U7_0),.dout(w_dff_B_l6H5NuBV9_0),.clk(gclk));
	jdff dff_B_bJFMvIC76_0(.din(w_dff_B_l6H5NuBV9_0),.dout(w_dff_B_bJFMvIC76_0),.clk(gclk));
	jdff dff_B_4r81DgCj2_0(.din(w_dff_B_bJFMvIC76_0),.dout(w_dff_B_4r81DgCj2_0),.clk(gclk));
	jdff dff_B_eZdSR4q52_0(.din(w_dff_B_4r81DgCj2_0),.dout(w_dff_B_eZdSR4q52_0),.clk(gclk));
	jdff dff_B_6Js46pfn6_0(.din(w_dff_B_eZdSR4q52_0),.dout(w_dff_B_6Js46pfn6_0),.clk(gclk));
	jdff dff_B_QVqjuezl8_0(.din(w_dff_B_6Js46pfn6_0),.dout(w_dff_B_QVqjuezl8_0),.clk(gclk));
	jdff dff_B_2qPGzj4G6_0(.din(w_dff_B_QVqjuezl8_0),.dout(w_dff_B_2qPGzj4G6_0),.clk(gclk));
	jdff dff_B_8yTE7N012_0(.din(w_dff_B_2qPGzj4G6_0),.dout(w_dff_B_8yTE7N012_0),.clk(gclk));
	jdff dff_B_n41vpbyU5_0(.din(w_dff_B_8yTE7N012_0),.dout(w_dff_B_n41vpbyU5_0),.clk(gclk));
	jdff dff_B_jKZdXvcN2_0(.din(w_dff_B_n41vpbyU5_0),.dout(w_dff_B_jKZdXvcN2_0),.clk(gclk));
	jdff dff_B_us1IIPa28_0(.din(w_dff_B_jKZdXvcN2_0),.dout(w_dff_B_us1IIPa28_0),.clk(gclk));
	jdff dff_B_HgbC4rMv0_0(.din(w_dff_B_us1IIPa28_0),.dout(w_dff_B_HgbC4rMv0_0),.clk(gclk));
	jdff dff_B_y5QRl9T57_0(.din(w_dff_B_HgbC4rMv0_0),.dout(w_dff_B_y5QRl9T57_0),.clk(gclk));
	jdff dff_B_xWkFxl7Y9_0(.din(w_dff_B_y5QRl9T57_0),.dout(w_dff_B_xWkFxl7Y9_0),.clk(gclk));
	jdff dff_B_J3Ebs7Pn4_0(.din(w_dff_B_xWkFxl7Y9_0),.dout(w_dff_B_J3Ebs7Pn4_0),.clk(gclk));
	jdff dff_B_ZW4dlhnT8_0(.din(w_dff_B_J3Ebs7Pn4_0),.dout(w_dff_B_ZW4dlhnT8_0),.clk(gclk));
	jdff dff_B_jR8AcVOh7_0(.din(w_dff_B_ZW4dlhnT8_0),.dout(w_dff_B_jR8AcVOh7_0),.clk(gclk));
	jdff dff_B_sKchNxYA3_0(.din(w_dff_B_jR8AcVOh7_0),.dout(w_dff_B_sKchNxYA3_0),.clk(gclk));
	jdff dff_B_RpgGaSTt0_0(.din(w_dff_B_sKchNxYA3_0),.dout(w_dff_B_RpgGaSTt0_0),.clk(gclk));
	jdff dff_B_Xd3u2lNs0_0(.din(w_dff_B_RpgGaSTt0_0),.dout(w_dff_B_Xd3u2lNs0_0),.clk(gclk));
	jdff dff_B_Ix4QkzFX5_0(.din(w_dff_B_Xd3u2lNs0_0),.dout(w_dff_B_Ix4QkzFX5_0),.clk(gclk));
	jdff dff_B_YRvKzS0T1_0(.din(w_dff_B_Ix4QkzFX5_0),.dout(w_dff_B_YRvKzS0T1_0),.clk(gclk));
	jdff dff_B_CtZzvZcf9_0(.din(w_dff_B_YRvKzS0T1_0),.dout(w_dff_B_CtZzvZcf9_0),.clk(gclk));
	jdff dff_B_IOd6Jlkx8_0(.din(w_dff_B_CtZzvZcf9_0),.dout(w_dff_B_IOd6Jlkx8_0),.clk(gclk));
	jdff dff_B_z8sCIKSH0_0(.din(w_dff_B_IOd6Jlkx8_0),.dout(w_dff_B_z8sCIKSH0_0),.clk(gclk));
	jdff dff_B_Dp7MEQVe0_0(.din(w_dff_B_z8sCIKSH0_0),.dout(w_dff_B_Dp7MEQVe0_0),.clk(gclk));
	jdff dff_B_hf9tfxjv8_0(.din(w_dff_B_Dp7MEQVe0_0),.dout(w_dff_B_hf9tfxjv8_0),.clk(gclk));
	jdff dff_B_VwSvjwLC5_0(.din(w_dff_B_hf9tfxjv8_0),.dout(w_dff_B_VwSvjwLC5_0),.clk(gclk));
	jdff dff_B_A13X0RKi1_0(.din(w_dff_B_VwSvjwLC5_0),.dout(w_dff_B_A13X0RKi1_0),.clk(gclk));
	jdff dff_B_69jdkr2X4_0(.din(w_dff_B_A13X0RKi1_0),.dout(w_dff_B_69jdkr2X4_0),.clk(gclk));
	jdff dff_B_rOPpMwfn2_0(.din(w_dff_B_69jdkr2X4_0),.dout(w_dff_B_rOPpMwfn2_0),.clk(gclk));
	jdff dff_B_m3eUTp5i8_0(.din(w_dff_B_rOPpMwfn2_0),.dout(w_dff_B_m3eUTp5i8_0),.clk(gclk));
	jdff dff_B_KHpBvGl34_0(.din(w_dff_B_m3eUTp5i8_0),.dout(w_dff_B_KHpBvGl34_0),.clk(gclk));
	jdff dff_B_fE6COzPy2_0(.din(w_dff_B_KHpBvGl34_0),.dout(w_dff_B_fE6COzPy2_0),.clk(gclk));
	jdff dff_B_BsF4gmAC7_0(.din(w_dff_B_fE6COzPy2_0),.dout(w_dff_B_BsF4gmAC7_0),.clk(gclk));
	jdff dff_B_NEKHiB8j6_0(.din(w_dff_B_BsF4gmAC7_0),.dout(w_dff_B_NEKHiB8j6_0),.clk(gclk));
	jdff dff_B_IzQy6DU01_0(.din(w_dff_B_NEKHiB8j6_0),.dout(w_dff_B_IzQy6DU01_0),.clk(gclk));
	jdff dff_B_HJ6lVrTb0_1(.din(n1008),.dout(w_dff_B_HJ6lVrTb0_1),.clk(gclk));
	jdff dff_B_HkwNynPJ9_1(.din(w_dff_B_HJ6lVrTb0_1),.dout(w_dff_B_HkwNynPJ9_1),.clk(gclk));
	jdff dff_B_a6fYzwqM7_1(.din(w_dff_B_HkwNynPJ9_1),.dout(w_dff_B_a6fYzwqM7_1),.clk(gclk));
	jdff dff_B_W8m1CUOh6_1(.din(w_dff_B_a6fYzwqM7_1),.dout(w_dff_B_W8m1CUOh6_1),.clk(gclk));
	jdff dff_B_ZcbKwOBE0_1(.din(w_dff_B_W8m1CUOh6_1),.dout(w_dff_B_ZcbKwOBE0_1),.clk(gclk));
	jdff dff_B_xkLvKH0P2_1(.din(w_dff_B_ZcbKwOBE0_1),.dout(w_dff_B_xkLvKH0P2_1),.clk(gclk));
	jdff dff_B_5uwaqEZk0_1(.din(w_dff_B_xkLvKH0P2_1),.dout(w_dff_B_5uwaqEZk0_1),.clk(gclk));
	jdff dff_B_GrGmLSE58_1(.din(w_dff_B_5uwaqEZk0_1),.dout(w_dff_B_GrGmLSE58_1),.clk(gclk));
	jdff dff_B_JYWOJZGU1_1(.din(w_dff_B_GrGmLSE58_1),.dout(w_dff_B_JYWOJZGU1_1),.clk(gclk));
	jdff dff_B_gLcofKyE3_1(.din(w_dff_B_JYWOJZGU1_1),.dout(w_dff_B_gLcofKyE3_1),.clk(gclk));
	jdff dff_B_Eim1cGsx4_1(.din(w_dff_B_gLcofKyE3_1),.dout(w_dff_B_Eim1cGsx4_1),.clk(gclk));
	jdff dff_B_Y5O0ij5F6_1(.din(w_dff_B_Eim1cGsx4_1),.dout(w_dff_B_Y5O0ij5F6_1),.clk(gclk));
	jdff dff_B_ofxVtgf67_1(.din(w_dff_B_Y5O0ij5F6_1),.dout(w_dff_B_ofxVtgf67_1),.clk(gclk));
	jdff dff_B_7diVCkaV2_1(.din(w_dff_B_ofxVtgf67_1),.dout(w_dff_B_7diVCkaV2_1),.clk(gclk));
	jdff dff_B_pMh7tMWD6_1(.din(w_dff_B_7diVCkaV2_1),.dout(w_dff_B_pMh7tMWD6_1),.clk(gclk));
	jdff dff_B_fmQNbMFh3_1(.din(w_dff_B_pMh7tMWD6_1),.dout(w_dff_B_fmQNbMFh3_1),.clk(gclk));
	jdff dff_B_2q9IsWxb7_1(.din(w_dff_B_fmQNbMFh3_1),.dout(w_dff_B_2q9IsWxb7_1),.clk(gclk));
	jdff dff_B_RACxajck2_1(.din(w_dff_B_2q9IsWxb7_1),.dout(w_dff_B_RACxajck2_1),.clk(gclk));
	jdff dff_B_aA4nJKB04_1(.din(w_dff_B_RACxajck2_1),.dout(w_dff_B_aA4nJKB04_1),.clk(gclk));
	jdff dff_B_HFsZEE1F0_1(.din(w_dff_B_aA4nJKB04_1),.dout(w_dff_B_HFsZEE1F0_1),.clk(gclk));
	jdff dff_B_GXQsBL7t1_1(.din(w_dff_B_HFsZEE1F0_1),.dout(w_dff_B_GXQsBL7t1_1),.clk(gclk));
	jdff dff_B_UHuE8k1I4_1(.din(w_dff_B_GXQsBL7t1_1),.dout(w_dff_B_UHuE8k1I4_1),.clk(gclk));
	jdff dff_B_THM0uF6f7_1(.din(w_dff_B_UHuE8k1I4_1),.dout(w_dff_B_THM0uF6f7_1),.clk(gclk));
	jdff dff_B_PGzZk2nL0_1(.din(w_dff_B_THM0uF6f7_1),.dout(w_dff_B_PGzZk2nL0_1),.clk(gclk));
	jdff dff_B_0PKHyQ317_1(.din(w_dff_B_PGzZk2nL0_1),.dout(w_dff_B_0PKHyQ317_1),.clk(gclk));
	jdff dff_B_KR5q2HIy6_1(.din(w_dff_B_0PKHyQ317_1),.dout(w_dff_B_KR5q2HIy6_1),.clk(gclk));
	jdff dff_B_RydqBP1p9_1(.din(w_dff_B_KR5q2HIy6_1),.dout(w_dff_B_RydqBP1p9_1),.clk(gclk));
	jdff dff_B_Y22SUoGK6_1(.din(w_dff_B_RydqBP1p9_1),.dout(w_dff_B_Y22SUoGK6_1),.clk(gclk));
	jdff dff_B_yHwmgnXE8_1(.din(w_dff_B_Y22SUoGK6_1),.dout(w_dff_B_yHwmgnXE8_1),.clk(gclk));
	jdff dff_B_G2gFgPUO7_1(.din(w_dff_B_yHwmgnXE8_1),.dout(w_dff_B_G2gFgPUO7_1),.clk(gclk));
	jdff dff_B_8dit25wa2_1(.din(w_dff_B_G2gFgPUO7_1),.dout(w_dff_B_8dit25wa2_1),.clk(gclk));
	jdff dff_B_90FidDOm4_1(.din(w_dff_B_8dit25wa2_1),.dout(w_dff_B_90FidDOm4_1),.clk(gclk));
	jdff dff_B_NUURd4pn0_1(.din(w_dff_B_90FidDOm4_1),.dout(w_dff_B_NUURd4pn0_1),.clk(gclk));
	jdff dff_B_u5sGMKrC3_1(.din(w_dff_B_NUURd4pn0_1),.dout(w_dff_B_u5sGMKrC3_1),.clk(gclk));
	jdff dff_B_kdSgblys0_1(.din(w_dff_B_u5sGMKrC3_1),.dout(w_dff_B_kdSgblys0_1),.clk(gclk));
	jdff dff_B_08D9uipu3_1(.din(w_dff_B_kdSgblys0_1),.dout(w_dff_B_08D9uipu3_1),.clk(gclk));
	jdff dff_B_N8AFf5hJ8_1(.din(w_dff_B_08D9uipu3_1),.dout(w_dff_B_N8AFf5hJ8_1),.clk(gclk));
	jdff dff_B_pvAnsIew8_1(.din(w_dff_B_N8AFf5hJ8_1),.dout(w_dff_B_pvAnsIew8_1),.clk(gclk));
	jdff dff_B_iZzPuJhS9_1(.din(w_dff_B_pvAnsIew8_1),.dout(w_dff_B_iZzPuJhS9_1),.clk(gclk));
	jdff dff_B_SKauuycG8_1(.din(w_dff_B_iZzPuJhS9_1),.dout(w_dff_B_SKauuycG8_1),.clk(gclk));
	jdff dff_B_0rekuKli1_1(.din(w_dff_B_SKauuycG8_1),.dout(w_dff_B_0rekuKli1_1),.clk(gclk));
	jdff dff_B_OTPE3UwP1_1(.din(w_dff_B_0rekuKli1_1),.dout(w_dff_B_OTPE3UwP1_1),.clk(gclk));
	jdff dff_B_BwG9m3In4_1(.din(w_dff_B_OTPE3UwP1_1),.dout(w_dff_B_BwG9m3In4_1),.clk(gclk));
	jdff dff_B_DTH32o8H2_1(.din(w_dff_B_BwG9m3In4_1),.dout(w_dff_B_DTH32o8H2_1),.clk(gclk));
	jdff dff_B_SKS1RfRB5_1(.din(w_dff_B_DTH32o8H2_1),.dout(w_dff_B_SKS1RfRB5_1),.clk(gclk));
	jdff dff_B_rtdb7BK05_1(.din(w_dff_B_SKS1RfRB5_1),.dout(w_dff_B_rtdb7BK05_1),.clk(gclk));
	jdff dff_B_YTvAxG3Q3_1(.din(w_dff_B_rtdb7BK05_1),.dout(w_dff_B_YTvAxG3Q3_1),.clk(gclk));
	jdff dff_B_J7rm1AFB5_1(.din(w_dff_B_YTvAxG3Q3_1),.dout(w_dff_B_J7rm1AFB5_1),.clk(gclk));
	jdff dff_B_f6BytXrQ8_1(.din(w_dff_B_J7rm1AFB5_1),.dout(w_dff_B_f6BytXrQ8_1),.clk(gclk));
	jdff dff_B_y0Lqhrfb8_1(.din(w_dff_B_f6BytXrQ8_1),.dout(w_dff_B_y0Lqhrfb8_1),.clk(gclk));
	jdff dff_B_djeOODWI7_1(.din(w_dff_B_y0Lqhrfb8_1),.dout(w_dff_B_djeOODWI7_1),.clk(gclk));
	jdff dff_B_uliD3X7z1_1(.din(w_dff_B_djeOODWI7_1),.dout(w_dff_B_uliD3X7z1_1),.clk(gclk));
	jdff dff_B_vbnuL4pR8_1(.din(w_dff_B_uliD3X7z1_1),.dout(w_dff_B_vbnuL4pR8_1),.clk(gclk));
	jdff dff_B_atxwU3iB6_1(.din(w_dff_B_vbnuL4pR8_1),.dout(w_dff_B_atxwU3iB6_1),.clk(gclk));
	jdff dff_B_v2jjmF4A6_1(.din(w_dff_B_atxwU3iB6_1),.dout(w_dff_B_v2jjmF4A6_1),.clk(gclk));
	jdff dff_B_wDE1PLUR8_1(.din(w_dff_B_v2jjmF4A6_1),.dout(w_dff_B_wDE1PLUR8_1),.clk(gclk));
	jdff dff_B_3H8ZsqCZ7_1(.din(w_dff_B_wDE1PLUR8_1),.dout(w_dff_B_3H8ZsqCZ7_1),.clk(gclk));
	jdff dff_B_YXFcmwWs9_1(.din(w_dff_B_3H8ZsqCZ7_1),.dout(w_dff_B_YXFcmwWs9_1),.clk(gclk));
	jdff dff_B_LHKzxVsH5_1(.din(w_dff_B_YXFcmwWs9_1),.dout(w_dff_B_LHKzxVsH5_1),.clk(gclk));
	jdff dff_B_9sC2MBoT7_1(.din(w_dff_B_LHKzxVsH5_1),.dout(w_dff_B_9sC2MBoT7_1),.clk(gclk));
	jdff dff_B_jt4JEY7O0_1(.din(w_dff_B_9sC2MBoT7_1),.dout(w_dff_B_jt4JEY7O0_1),.clk(gclk));
	jdff dff_B_Rr9mJgn85_1(.din(w_dff_B_jt4JEY7O0_1),.dout(w_dff_B_Rr9mJgn85_1),.clk(gclk));
	jdff dff_B_MJ99dW0b5_1(.din(w_dff_B_Rr9mJgn85_1),.dout(w_dff_B_MJ99dW0b5_1),.clk(gclk));
	jdff dff_B_CeGqMrfq0_1(.din(w_dff_B_MJ99dW0b5_1),.dout(w_dff_B_CeGqMrfq0_1),.clk(gclk));
	jdff dff_B_gU7WsBuK3_1(.din(w_dff_B_CeGqMrfq0_1),.dout(w_dff_B_gU7WsBuK3_1),.clk(gclk));
	jdff dff_B_J15nntqZ7_1(.din(w_dff_B_gU7WsBuK3_1),.dout(w_dff_B_J15nntqZ7_1),.clk(gclk));
	jdff dff_B_WM8n7qpW1_1(.din(w_dff_B_J15nntqZ7_1),.dout(w_dff_B_WM8n7qpW1_1),.clk(gclk));
	jdff dff_B_3e0YboH48_1(.din(w_dff_B_WM8n7qpW1_1),.dout(w_dff_B_3e0YboH48_1),.clk(gclk));
	jdff dff_B_ocQ8UxSp3_1(.din(w_dff_B_3e0YboH48_1),.dout(w_dff_B_ocQ8UxSp3_1),.clk(gclk));
	jdff dff_B_BfuFaR1d6_1(.din(w_dff_B_ocQ8UxSp3_1),.dout(w_dff_B_BfuFaR1d6_1),.clk(gclk));
	jdff dff_B_07ZFZeeX9_1(.din(w_dff_B_BfuFaR1d6_1),.dout(w_dff_B_07ZFZeeX9_1),.clk(gclk));
	jdff dff_B_qvImErpT1_1(.din(w_dff_B_07ZFZeeX9_1),.dout(w_dff_B_qvImErpT1_1),.clk(gclk));
	jdff dff_B_Q3Hnkmqj8_1(.din(w_dff_B_qvImErpT1_1),.dout(w_dff_B_Q3Hnkmqj8_1),.clk(gclk));
	jdff dff_B_dBKNN4PM7_1(.din(w_dff_B_Q3Hnkmqj8_1),.dout(w_dff_B_dBKNN4PM7_1),.clk(gclk));
	jdff dff_B_SsCfeRrd7_1(.din(w_dff_B_dBKNN4PM7_1),.dout(w_dff_B_SsCfeRrd7_1),.clk(gclk));
	jdff dff_B_beMOGVr14_1(.din(w_dff_B_SsCfeRrd7_1),.dout(w_dff_B_beMOGVr14_1),.clk(gclk));
	jdff dff_B_yAAegxo65_1(.din(w_dff_B_beMOGVr14_1),.dout(w_dff_B_yAAegxo65_1),.clk(gclk));
	jdff dff_B_Wq0Zzxw80_1(.din(w_dff_B_yAAegxo65_1),.dout(w_dff_B_Wq0Zzxw80_1),.clk(gclk));
	jdff dff_B_O2Ynz6V51_1(.din(w_dff_B_Wq0Zzxw80_1),.dout(w_dff_B_O2Ynz6V51_1),.clk(gclk));
	jdff dff_B_IfGIIln55_1(.din(w_dff_B_O2Ynz6V51_1),.dout(w_dff_B_IfGIIln55_1),.clk(gclk));
	jdff dff_B_jOvVRSwm4_1(.din(w_dff_B_IfGIIln55_1),.dout(w_dff_B_jOvVRSwm4_1),.clk(gclk));
	jdff dff_B_uSbS7F3I1_1(.din(w_dff_B_jOvVRSwm4_1),.dout(w_dff_B_uSbS7F3I1_1),.clk(gclk));
	jdff dff_B_fWQu58r08_1(.din(w_dff_B_uSbS7F3I1_1),.dout(w_dff_B_fWQu58r08_1),.clk(gclk));
	jdff dff_B_5UACoK6j5_1(.din(w_dff_B_fWQu58r08_1),.dout(w_dff_B_5UACoK6j5_1),.clk(gclk));
	jdff dff_B_8GVe9j025_1(.din(w_dff_B_5UACoK6j5_1),.dout(w_dff_B_8GVe9j025_1),.clk(gclk));
	jdff dff_B_ngKcFJy79_1(.din(w_dff_B_8GVe9j025_1),.dout(w_dff_B_ngKcFJy79_1),.clk(gclk));
	jdff dff_B_jZBtkeVy6_1(.din(w_dff_B_ngKcFJy79_1),.dout(w_dff_B_jZBtkeVy6_1),.clk(gclk));
	jdff dff_B_at6GQTXv8_1(.din(w_dff_B_jZBtkeVy6_1),.dout(w_dff_B_at6GQTXv8_1),.clk(gclk));
	jdff dff_B_dHtBVGU23_1(.din(w_dff_B_at6GQTXv8_1),.dout(w_dff_B_dHtBVGU23_1),.clk(gclk));
	jdff dff_B_KT2elHrl6_1(.din(w_dff_B_dHtBVGU23_1),.dout(w_dff_B_KT2elHrl6_1),.clk(gclk));
	jdff dff_B_t8xirMW40_1(.din(w_dff_B_KT2elHrl6_1),.dout(w_dff_B_t8xirMW40_1),.clk(gclk));
	jdff dff_B_8urqMdUE3_1(.din(w_dff_B_t8xirMW40_1),.dout(w_dff_B_8urqMdUE3_1),.clk(gclk));
	jdff dff_B_U53R5WUf2_1(.din(w_dff_B_8urqMdUE3_1),.dout(w_dff_B_U53R5WUf2_1),.clk(gclk));
	jdff dff_B_8l0aIOKA3_1(.din(w_dff_B_U53R5WUf2_1),.dout(w_dff_B_8l0aIOKA3_1),.clk(gclk));
	jdff dff_B_zTD1JsW25_1(.din(w_dff_B_8l0aIOKA3_1),.dout(w_dff_B_zTD1JsW25_1),.clk(gclk));
	jdff dff_B_kN8FSfJV4_1(.din(w_dff_B_zTD1JsW25_1),.dout(w_dff_B_kN8FSfJV4_1),.clk(gclk));
	jdff dff_B_dO9uMtjr9_1(.din(w_dff_B_kN8FSfJV4_1),.dout(w_dff_B_dO9uMtjr9_1),.clk(gclk));
	jdff dff_B_E1yN1Em58_1(.din(w_dff_B_dO9uMtjr9_1),.dout(w_dff_B_E1yN1Em58_1),.clk(gclk));
	jdff dff_B_joxinVQu3_1(.din(w_dff_B_E1yN1Em58_1),.dout(w_dff_B_joxinVQu3_1),.clk(gclk));
	jdff dff_B_mvlqfd8N7_1(.din(w_dff_B_joxinVQu3_1),.dout(w_dff_B_mvlqfd8N7_1),.clk(gclk));
	jdff dff_B_OBSvF7gD7_1(.din(w_dff_B_mvlqfd8N7_1),.dout(w_dff_B_OBSvF7gD7_1),.clk(gclk));
	jdff dff_B_GAkGCBbr8_1(.din(w_dff_B_OBSvF7gD7_1),.dout(w_dff_B_GAkGCBbr8_1),.clk(gclk));
	jdff dff_B_LVI8cSBi3_1(.din(w_dff_B_GAkGCBbr8_1),.dout(w_dff_B_LVI8cSBi3_1),.clk(gclk));
	jdff dff_B_8BuCOaXp1_1(.din(w_dff_B_LVI8cSBi3_1),.dout(w_dff_B_8BuCOaXp1_1),.clk(gclk));
	jdff dff_B_LI1muG7X8_0(.din(n1009),.dout(w_dff_B_LI1muG7X8_0),.clk(gclk));
	jdff dff_B_egmYcb4j8_0(.din(w_dff_B_LI1muG7X8_0),.dout(w_dff_B_egmYcb4j8_0),.clk(gclk));
	jdff dff_B_HfoUMNU27_0(.din(w_dff_B_egmYcb4j8_0),.dout(w_dff_B_HfoUMNU27_0),.clk(gclk));
	jdff dff_B_leG3NFcU0_0(.din(w_dff_B_HfoUMNU27_0),.dout(w_dff_B_leG3NFcU0_0),.clk(gclk));
	jdff dff_B_eoOSUF5U2_0(.din(w_dff_B_leG3NFcU0_0),.dout(w_dff_B_eoOSUF5U2_0),.clk(gclk));
	jdff dff_B_qCOw17NJ7_0(.din(w_dff_B_eoOSUF5U2_0),.dout(w_dff_B_qCOw17NJ7_0),.clk(gclk));
	jdff dff_B_8qF4oLp59_0(.din(w_dff_B_qCOw17NJ7_0),.dout(w_dff_B_8qF4oLp59_0),.clk(gclk));
	jdff dff_B_sxL51aso2_0(.din(w_dff_B_8qF4oLp59_0),.dout(w_dff_B_sxL51aso2_0),.clk(gclk));
	jdff dff_B_7JLICGiQ1_0(.din(w_dff_B_sxL51aso2_0),.dout(w_dff_B_7JLICGiQ1_0),.clk(gclk));
	jdff dff_B_ZkmMBWjr2_0(.din(w_dff_B_7JLICGiQ1_0),.dout(w_dff_B_ZkmMBWjr2_0),.clk(gclk));
	jdff dff_B_b77E3YUu2_0(.din(w_dff_B_ZkmMBWjr2_0),.dout(w_dff_B_b77E3YUu2_0),.clk(gclk));
	jdff dff_B_Dhb34zyI0_0(.din(w_dff_B_b77E3YUu2_0),.dout(w_dff_B_Dhb34zyI0_0),.clk(gclk));
	jdff dff_B_Hjcx7EUi8_0(.din(w_dff_B_Dhb34zyI0_0),.dout(w_dff_B_Hjcx7EUi8_0),.clk(gclk));
	jdff dff_B_8N8u9eN09_0(.din(w_dff_B_Hjcx7EUi8_0),.dout(w_dff_B_8N8u9eN09_0),.clk(gclk));
	jdff dff_B_sI6GdHPP9_0(.din(w_dff_B_8N8u9eN09_0),.dout(w_dff_B_sI6GdHPP9_0),.clk(gclk));
	jdff dff_B_ZnyUfvvH2_0(.din(w_dff_B_sI6GdHPP9_0),.dout(w_dff_B_ZnyUfvvH2_0),.clk(gclk));
	jdff dff_B_AFG806F59_0(.din(w_dff_B_ZnyUfvvH2_0),.dout(w_dff_B_AFG806F59_0),.clk(gclk));
	jdff dff_B_XEjjwvcA2_0(.din(w_dff_B_AFG806F59_0),.dout(w_dff_B_XEjjwvcA2_0),.clk(gclk));
	jdff dff_B_iWd2cdY69_0(.din(w_dff_B_XEjjwvcA2_0),.dout(w_dff_B_iWd2cdY69_0),.clk(gclk));
	jdff dff_B_HWk4etxo7_0(.din(w_dff_B_iWd2cdY69_0),.dout(w_dff_B_HWk4etxo7_0),.clk(gclk));
	jdff dff_B_fghiXM9g4_0(.din(w_dff_B_HWk4etxo7_0),.dout(w_dff_B_fghiXM9g4_0),.clk(gclk));
	jdff dff_B_D4NjwCDp5_0(.din(w_dff_B_fghiXM9g4_0),.dout(w_dff_B_D4NjwCDp5_0),.clk(gclk));
	jdff dff_B_muBPgzAl6_0(.din(w_dff_B_D4NjwCDp5_0),.dout(w_dff_B_muBPgzAl6_0),.clk(gclk));
	jdff dff_B_n9eQtlS83_0(.din(w_dff_B_muBPgzAl6_0),.dout(w_dff_B_n9eQtlS83_0),.clk(gclk));
	jdff dff_B_3OjDPwgO6_0(.din(w_dff_B_n9eQtlS83_0),.dout(w_dff_B_3OjDPwgO6_0),.clk(gclk));
	jdff dff_B_EjSBSspc0_0(.din(w_dff_B_3OjDPwgO6_0),.dout(w_dff_B_EjSBSspc0_0),.clk(gclk));
	jdff dff_B_4mltlmjF4_0(.din(w_dff_B_EjSBSspc0_0),.dout(w_dff_B_4mltlmjF4_0),.clk(gclk));
	jdff dff_B_IWj7SB838_0(.din(w_dff_B_4mltlmjF4_0),.dout(w_dff_B_IWj7SB838_0),.clk(gclk));
	jdff dff_B_r5X8XCsD4_0(.din(w_dff_B_IWj7SB838_0),.dout(w_dff_B_r5X8XCsD4_0),.clk(gclk));
	jdff dff_B_q9kbxnmm7_0(.din(w_dff_B_r5X8XCsD4_0),.dout(w_dff_B_q9kbxnmm7_0),.clk(gclk));
	jdff dff_B_DefmhDpX7_0(.din(w_dff_B_q9kbxnmm7_0),.dout(w_dff_B_DefmhDpX7_0),.clk(gclk));
	jdff dff_B_eVJhgeTY2_0(.din(w_dff_B_DefmhDpX7_0),.dout(w_dff_B_eVJhgeTY2_0),.clk(gclk));
	jdff dff_B_fsDrF0vM9_0(.din(w_dff_B_eVJhgeTY2_0),.dout(w_dff_B_fsDrF0vM9_0),.clk(gclk));
	jdff dff_B_0tQLHKNs6_0(.din(w_dff_B_fsDrF0vM9_0),.dout(w_dff_B_0tQLHKNs6_0),.clk(gclk));
	jdff dff_B_63DrpowM4_0(.din(w_dff_B_0tQLHKNs6_0),.dout(w_dff_B_63DrpowM4_0),.clk(gclk));
	jdff dff_B_YF2Zahn03_0(.din(w_dff_B_63DrpowM4_0),.dout(w_dff_B_YF2Zahn03_0),.clk(gclk));
	jdff dff_B_Ey5PKPlS0_0(.din(w_dff_B_YF2Zahn03_0),.dout(w_dff_B_Ey5PKPlS0_0),.clk(gclk));
	jdff dff_B_3oz5WrYv2_0(.din(w_dff_B_Ey5PKPlS0_0),.dout(w_dff_B_3oz5WrYv2_0),.clk(gclk));
	jdff dff_B_op98yKlS5_0(.din(w_dff_B_3oz5WrYv2_0),.dout(w_dff_B_op98yKlS5_0),.clk(gclk));
	jdff dff_B_mcsgzguU6_0(.din(w_dff_B_op98yKlS5_0),.dout(w_dff_B_mcsgzguU6_0),.clk(gclk));
	jdff dff_B_tLYShEHZ0_0(.din(w_dff_B_mcsgzguU6_0),.dout(w_dff_B_tLYShEHZ0_0),.clk(gclk));
	jdff dff_B_6S6tvjRH1_0(.din(w_dff_B_tLYShEHZ0_0),.dout(w_dff_B_6S6tvjRH1_0),.clk(gclk));
	jdff dff_B_jplVcPNJ0_0(.din(w_dff_B_6S6tvjRH1_0),.dout(w_dff_B_jplVcPNJ0_0),.clk(gclk));
	jdff dff_B_Qhxplqxv4_0(.din(w_dff_B_jplVcPNJ0_0),.dout(w_dff_B_Qhxplqxv4_0),.clk(gclk));
	jdff dff_B_9RVKo98I3_0(.din(w_dff_B_Qhxplqxv4_0),.dout(w_dff_B_9RVKo98I3_0),.clk(gclk));
	jdff dff_B_IpDIJSNC8_0(.din(w_dff_B_9RVKo98I3_0),.dout(w_dff_B_IpDIJSNC8_0),.clk(gclk));
	jdff dff_B_fNMQA6Vj7_0(.din(w_dff_B_IpDIJSNC8_0),.dout(w_dff_B_fNMQA6Vj7_0),.clk(gclk));
	jdff dff_B_7S6qvp1Z9_0(.din(w_dff_B_fNMQA6Vj7_0),.dout(w_dff_B_7S6qvp1Z9_0),.clk(gclk));
	jdff dff_B_3IngINET2_0(.din(w_dff_B_7S6qvp1Z9_0),.dout(w_dff_B_3IngINET2_0),.clk(gclk));
	jdff dff_B_qecdS1VE6_0(.din(w_dff_B_3IngINET2_0),.dout(w_dff_B_qecdS1VE6_0),.clk(gclk));
	jdff dff_B_pXJIDVD74_0(.din(w_dff_B_qecdS1VE6_0),.dout(w_dff_B_pXJIDVD74_0),.clk(gclk));
	jdff dff_B_LeWZ4lhu7_0(.din(w_dff_B_pXJIDVD74_0),.dout(w_dff_B_LeWZ4lhu7_0),.clk(gclk));
	jdff dff_B_Rr7I6YOX2_0(.din(w_dff_B_LeWZ4lhu7_0),.dout(w_dff_B_Rr7I6YOX2_0),.clk(gclk));
	jdff dff_B_dIapvW9Q9_0(.din(w_dff_B_Rr7I6YOX2_0),.dout(w_dff_B_dIapvW9Q9_0),.clk(gclk));
	jdff dff_B_UBSKpJyw0_0(.din(w_dff_B_dIapvW9Q9_0),.dout(w_dff_B_UBSKpJyw0_0),.clk(gclk));
	jdff dff_B_nZt4nX8L4_0(.din(w_dff_B_UBSKpJyw0_0),.dout(w_dff_B_nZt4nX8L4_0),.clk(gclk));
	jdff dff_B_K5UkPmBo3_0(.din(w_dff_B_nZt4nX8L4_0),.dout(w_dff_B_K5UkPmBo3_0),.clk(gclk));
	jdff dff_B_11k69KHb6_0(.din(w_dff_B_K5UkPmBo3_0),.dout(w_dff_B_11k69KHb6_0),.clk(gclk));
	jdff dff_B_YWR2y9KU3_0(.din(w_dff_B_11k69KHb6_0),.dout(w_dff_B_YWR2y9KU3_0),.clk(gclk));
	jdff dff_B_3gak01wb9_0(.din(w_dff_B_YWR2y9KU3_0),.dout(w_dff_B_3gak01wb9_0),.clk(gclk));
	jdff dff_B_m7ehzTDk3_0(.din(w_dff_B_3gak01wb9_0),.dout(w_dff_B_m7ehzTDk3_0),.clk(gclk));
	jdff dff_B_NEgDjvWA6_0(.din(w_dff_B_m7ehzTDk3_0),.dout(w_dff_B_NEgDjvWA6_0),.clk(gclk));
	jdff dff_B_ffiE4x1C0_0(.din(w_dff_B_NEgDjvWA6_0),.dout(w_dff_B_ffiE4x1C0_0),.clk(gclk));
	jdff dff_B_r4Lt7h438_0(.din(w_dff_B_ffiE4x1C0_0),.dout(w_dff_B_r4Lt7h438_0),.clk(gclk));
	jdff dff_B_ycii6xhC3_0(.din(w_dff_B_r4Lt7h438_0),.dout(w_dff_B_ycii6xhC3_0),.clk(gclk));
	jdff dff_B_m9B9t76Q1_0(.din(w_dff_B_ycii6xhC3_0),.dout(w_dff_B_m9B9t76Q1_0),.clk(gclk));
	jdff dff_B_EhxT2tTV8_0(.din(w_dff_B_m9B9t76Q1_0),.dout(w_dff_B_EhxT2tTV8_0),.clk(gclk));
	jdff dff_B_oXh7r5bD6_0(.din(w_dff_B_EhxT2tTV8_0),.dout(w_dff_B_oXh7r5bD6_0),.clk(gclk));
	jdff dff_B_QNMF3iAj8_0(.din(w_dff_B_oXh7r5bD6_0),.dout(w_dff_B_QNMF3iAj8_0),.clk(gclk));
	jdff dff_B_xzEZGPjV0_0(.din(w_dff_B_QNMF3iAj8_0),.dout(w_dff_B_xzEZGPjV0_0),.clk(gclk));
	jdff dff_B_VeDMNrz93_0(.din(w_dff_B_xzEZGPjV0_0),.dout(w_dff_B_VeDMNrz93_0),.clk(gclk));
	jdff dff_B_N9e2qZxf6_0(.din(w_dff_B_VeDMNrz93_0),.dout(w_dff_B_N9e2qZxf6_0),.clk(gclk));
	jdff dff_B_UJ4GEoou0_0(.din(w_dff_B_N9e2qZxf6_0),.dout(w_dff_B_UJ4GEoou0_0),.clk(gclk));
	jdff dff_B_EwpETrgg3_0(.din(w_dff_B_UJ4GEoou0_0),.dout(w_dff_B_EwpETrgg3_0),.clk(gclk));
	jdff dff_B_X3WEBxMB5_0(.din(w_dff_B_EwpETrgg3_0),.dout(w_dff_B_X3WEBxMB5_0),.clk(gclk));
	jdff dff_B_zZOEJAJj1_0(.din(w_dff_B_X3WEBxMB5_0),.dout(w_dff_B_zZOEJAJj1_0),.clk(gclk));
	jdff dff_B_cTcYrSu97_0(.din(w_dff_B_zZOEJAJj1_0),.dout(w_dff_B_cTcYrSu97_0),.clk(gclk));
	jdff dff_B_S9bhGfzF2_0(.din(w_dff_B_cTcYrSu97_0),.dout(w_dff_B_S9bhGfzF2_0),.clk(gclk));
	jdff dff_B_aYcVxeT15_0(.din(w_dff_B_S9bhGfzF2_0),.dout(w_dff_B_aYcVxeT15_0),.clk(gclk));
	jdff dff_B_ap8LFJF55_0(.din(w_dff_B_aYcVxeT15_0),.dout(w_dff_B_ap8LFJF55_0),.clk(gclk));
	jdff dff_B_LgZlzfhn2_0(.din(w_dff_B_ap8LFJF55_0),.dout(w_dff_B_LgZlzfhn2_0),.clk(gclk));
	jdff dff_B_1CkPniOb4_0(.din(w_dff_B_LgZlzfhn2_0),.dout(w_dff_B_1CkPniOb4_0),.clk(gclk));
	jdff dff_B_EE51UNaF4_0(.din(w_dff_B_1CkPniOb4_0),.dout(w_dff_B_EE51UNaF4_0),.clk(gclk));
	jdff dff_B_NdNDA36K1_0(.din(w_dff_B_EE51UNaF4_0),.dout(w_dff_B_NdNDA36K1_0),.clk(gclk));
	jdff dff_B_pwtiHkDR5_0(.din(w_dff_B_NdNDA36K1_0),.dout(w_dff_B_pwtiHkDR5_0),.clk(gclk));
	jdff dff_B_A0JEfiZv9_0(.din(w_dff_B_pwtiHkDR5_0),.dout(w_dff_B_A0JEfiZv9_0),.clk(gclk));
	jdff dff_B_cTLRItGK3_0(.din(w_dff_B_A0JEfiZv9_0),.dout(w_dff_B_cTLRItGK3_0),.clk(gclk));
	jdff dff_B_Z75AlfVW4_0(.din(w_dff_B_cTLRItGK3_0),.dout(w_dff_B_Z75AlfVW4_0),.clk(gclk));
	jdff dff_B_SRJLofgB3_0(.din(w_dff_B_Z75AlfVW4_0),.dout(w_dff_B_SRJLofgB3_0),.clk(gclk));
	jdff dff_B_aW6HM6pg6_0(.din(w_dff_B_SRJLofgB3_0),.dout(w_dff_B_aW6HM6pg6_0),.clk(gclk));
	jdff dff_B_l5e3fs230_0(.din(w_dff_B_aW6HM6pg6_0),.dout(w_dff_B_l5e3fs230_0),.clk(gclk));
	jdff dff_B_WK19l0Xf4_0(.din(w_dff_B_l5e3fs230_0),.dout(w_dff_B_WK19l0Xf4_0),.clk(gclk));
	jdff dff_B_SdlSwMMp4_0(.din(w_dff_B_WK19l0Xf4_0),.dout(w_dff_B_SdlSwMMp4_0),.clk(gclk));
	jdff dff_B_zHS1dsAy1_0(.din(w_dff_B_SdlSwMMp4_0),.dout(w_dff_B_zHS1dsAy1_0),.clk(gclk));
	jdff dff_B_ODRF0p9l2_0(.din(w_dff_B_zHS1dsAy1_0),.dout(w_dff_B_ODRF0p9l2_0),.clk(gclk));
	jdff dff_B_dDPTvBqu6_0(.din(w_dff_B_ODRF0p9l2_0),.dout(w_dff_B_dDPTvBqu6_0),.clk(gclk));
	jdff dff_B_ZhfzBMLk8_0(.din(w_dff_B_dDPTvBqu6_0),.dout(w_dff_B_ZhfzBMLk8_0),.clk(gclk));
	jdff dff_B_NwPrT38H6_0(.din(w_dff_B_ZhfzBMLk8_0),.dout(w_dff_B_NwPrT38H6_0),.clk(gclk));
	jdff dff_B_s6THB9RY5_0(.din(w_dff_B_NwPrT38H6_0),.dout(w_dff_B_s6THB9RY5_0),.clk(gclk));
	jdff dff_B_uYhXifJN1_0(.din(w_dff_B_s6THB9RY5_0),.dout(w_dff_B_uYhXifJN1_0),.clk(gclk));
	jdff dff_B_Rd53p9bN8_0(.din(w_dff_B_uYhXifJN1_0),.dout(w_dff_B_Rd53p9bN8_0),.clk(gclk));
	jdff dff_B_GpMM8Ys45_0(.din(w_dff_B_Rd53p9bN8_0),.dout(w_dff_B_GpMM8Ys45_0),.clk(gclk));
	jdff dff_B_GLfXb2JO5_0(.din(w_dff_B_GpMM8Ys45_0),.dout(w_dff_B_GLfXb2JO5_0),.clk(gclk));
	jdff dff_B_lEwdgnFZ1_0(.din(w_dff_B_GLfXb2JO5_0),.dout(w_dff_B_lEwdgnFZ1_0),.clk(gclk));
	jdff dff_B_fMaqATnV1_1(.din(n1002),.dout(w_dff_B_fMaqATnV1_1),.clk(gclk));
	jdff dff_B_LczZ2fgD9_1(.din(w_dff_B_fMaqATnV1_1),.dout(w_dff_B_LczZ2fgD9_1),.clk(gclk));
	jdff dff_B_gLfPJs2k8_1(.din(w_dff_B_LczZ2fgD9_1),.dout(w_dff_B_gLfPJs2k8_1),.clk(gclk));
	jdff dff_B_z5jm6e2X4_1(.din(w_dff_B_gLfPJs2k8_1),.dout(w_dff_B_z5jm6e2X4_1),.clk(gclk));
	jdff dff_B_wLqXc8Eh1_1(.din(w_dff_B_z5jm6e2X4_1),.dout(w_dff_B_wLqXc8Eh1_1),.clk(gclk));
	jdff dff_B_SIIPbB0c8_1(.din(w_dff_B_wLqXc8Eh1_1),.dout(w_dff_B_SIIPbB0c8_1),.clk(gclk));
	jdff dff_B_4AM10sF09_1(.din(w_dff_B_SIIPbB0c8_1),.dout(w_dff_B_4AM10sF09_1),.clk(gclk));
	jdff dff_B_pd3vKY0h6_1(.din(w_dff_B_4AM10sF09_1),.dout(w_dff_B_pd3vKY0h6_1),.clk(gclk));
	jdff dff_B_0zMj7xj78_1(.din(w_dff_B_pd3vKY0h6_1),.dout(w_dff_B_0zMj7xj78_1),.clk(gclk));
	jdff dff_B_GMOIlGUD1_1(.din(w_dff_B_0zMj7xj78_1),.dout(w_dff_B_GMOIlGUD1_1),.clk(gclk));
	jdff dff_B_Ywh1KOHj5_1(.din(w_dff_B_GMOIlGUD1_1),.dout(w_dff_B_Ywh1KOHj5_1),.clk(gclk));
	jdff dff_B_b8Wb6kc55_1(.din(w_dff_B_Ywh1KOHj5_1),.dout(w_dff_B_b8Wb6kc55_1),.clk(gclk));
	jdff dff_B_Xr7aWDK08_1(.din(w_dff_B_b8Wb6kc55_1),.dout(w_dff_B_Xr7aWDK08_1),.clk(gclk));
	jdff dff_B_7DXUnPAy7_1(.din(w_dff_B_Xr7aWDK08_1),.dout(w_dff_B_7DXUnPAy7_1),.clk(gclk));
	jdff dff_B_LGzYi79Y5_1(.din(w_dff_B_7DXUnPAy7_1),.dout(w_dff_B_LGzYi79Y5_1),.clk(gclk));
	jdff dff_B_WM1q6cKc9_1(.din(w_dff_B_LGzYi79Y5_1),.dout(w_dff_B_WM1q6cKc9_1),.clk(gclk));
	jdff dff_B_FLPkBcsF3_1(.din(w_dff_B_WM1q6cKc9_1),.dout(w_dff_B_FLPkBcsF3_1),.clk(gclk));
	jdff dff_B_i6NWirmn7_1(.din(w_dff_B_FLPkBcsF3_1),.dout(w_dff_B_i6NWirmn7_1),.clk(gclk));
	jdff dff_B_Iw7HvS4c2_1(.din(w_dff_B_i6NWirmn7_1),.dout(w_dff_B_Iw7HvS4c2_1),.clk(gclk));
	jdff dff_B_RCjBSv8K1_1(.din(w_dff_B_Iw7HvS4c2_1),.dout(w_dff_B_RCjBSv8K1_1),.clk(gclk));
	jdff dff_B_OD2pNKbW2_1(.din(w_dff_B_RCjBSv8K1_1),.dout(w_dff_B_OD2pNKbW2_1),.clk(gclk));
	jdff dff_B_5TNBViO54_1(.din(w_dff_B_OD2pNKbW2_1),.dout(w_dff_B_5TNBViO54_1),.clk(gclk));
	jdff dff_B_QWOOMs9C9_1(.din(w_dff_B_5TNBViO54_1),.dout(w_dff_B_QWOOMs9C9_1),.clk(gclk));
	jdff dff_B_ztaprmkK6_1(.din(w_dff_B_QWOOMs9C9_1),.dout(w_dff_B_ztaprmkK6_1),.clk(gclk));
	jdff dff_B_SEkV0cOO8_1(.din(w_dff_B_ztaprmkK6_1),.dout(w_dff_B_SEkV0cOO8_1),.clk(gclk));
	jdff dff_B_LabkkwI49_1(.din(w_dff_B_SEkV0cOO8_1),.dout(w_dff_B_LabkkwI49_1),.clk(gclk));
	jdff dff_B_swE72mfm0_1(.din(w_dff_B_LabkkwI49_1),.dout(w_dff_B_swE72mfm0_1),.clk(gclk));
	jdff dff_B_N2aQWDGN4_1(.din(w_dff_B_swE72mfm0_1),.dout(w_dff_B_N2aQWDGN4_1),.clk(gclk));
	jdff dff_B_IRWKwa7E2_1(.din(w_dff_B_N2aQWDGN4_1),.dout(w_dff_B_IRWKwa7E2_1),.clk(gclk));
	jdff dff_B_Bl3593RG5_1(.din(w_dff_B_IRWKwa7E2_1),.dout(w_dff_B_Bl3593RG5_1),.clk(gclk));
	jdff dff_B_ExjWkram7_1(.din(w_dff_B_Bl3593RG5_1),.dout(w_dff_B_ExjWkram7_1),.clk(gclk));
	jdff dff_B_da6W8suy0_1(.din(w_dff_B_ExjWkram7_1),.dout(w_dff_B_da6W8suy0_1),.clk(gclk));
	jdff dff_B_337b6h9I7_1(.din(w_dff_B_da6W8suy0_1),.dout(w_dff_B_337b6h9I7_1),.clk(gclk));
	jdff dff_B_YlBZKN7q4_1(.din(w_dff_B_337b6h9I7_1),.dout(w_dff_B_YlBZKN7q4_1),.clk(gclk));
	jdff dff_B_r02HyutI4_1(.din(w_dff_B_YlBZKN7q4_1),.dout(w_dff_B_r02HyutI4_1),.clk(gclk));
	jdff dff_B_0wmaVvbr9_1(.din(w_dff_B_r02HyutI4_1),.dout(w_dff_B_0wmaVvbr9_1),.clk(gclk));
	jdff dff_B_J2tPZ8I21_1(.din(w_dff_B_0wmaVvbr9_1),.dout(w_dff_B_J2tPZ8I21_1),.clk(gclk));
	jdff dff_B_RvfKmCGE5_1(.din(w_dff_B_J2tPZ8I21_1),.dout(w_dff_B_RvfKmCGE5_1),.clk(gclk));
	jdff dff_B_iT8shnqG8_1(.din(w_dff_B_RvfKmCGE5_1),.dout(w_dff_B_iT8shnqG8_1),.clk(gclk));
	jdff dff_B_elOvhyhE2_1(.din(w_dff_B_iT8shnqG8_1),.dout(w_dff_B_elOvhyhE2_1),.clk(gclk));
	jdff dff_B_0OAcjmcj5_1(.din(w_dff_B_elOvhyhE2_1),.dout(w_dff_B_0OAcjmcj5_1),.clk(gclk));
	jdff dff_B_DB2vbbvL0_1(.din(w_dff_B_0OAcjmcj5_1),.dout(w_dff_B_DB2vbbvL0_1),.clk(gclk));
	jdff dff_B_crSU5yex0_1(.din(w_dff_B_DB2vbbvL0_1),.dout(w_dff_B_crSU5yex0_1),.clk(gclk));
	jdff dff_B_BNfHpmXF5_1(.din(w_dff_B_crSU5yex0_1),.dout(w_dff_B_BNfHpmXF5_1),.clk(gclk));
	jdff dff_B_SAf1DYnP0_1(.din(w_dff_B_BNfHpmXF5_1),.dout(w_dff_B_SAf1DYnP0_1),.clk(gclk));
	jdff dff_B_PdDpRUEt9_1(.din(w_dff_B_SAf1DYnP0_1),.dout(w_dff_B_PdDpRUEt9_1),.clk(gclk));
	jdff dff_B_PzdBbhbu4_1(.din(w_dff_B_PdDpRUEt9_1),.dout(w_dff_B_PzdBbhbu4_1),.clk(gclk));
	jdff dff_B_23cEm7iu6_1(.din(w_dff_B_PzdBbhbu4_1),.dout(w_dff_B_23cEm7iu6_1),.clk(gclk));
	jdff dff_B_dfyFE99p5_1(.din(w_dff_B_23cEm7iu6_1),.dout(w_dff_B_dfyFE99p5_1),.clk(gclk));
	jdff dff_B_wnOzjbsO2_1(.din(w_dff_B_dfyFE99p5_1),.dout(w_dff_B_wnOzjbsO2_1),.clk(gclk));
	jdff dff_B_x64VKMPF9_1(.din(w_dff_B_wnOzjbsO2_1),.dout(w_dff_B_x64VKMPF9_1),.clk(gclk));
	jdff dff_B_WGIs6CrK3_1(.din(w_dff_B_x64VKMPF9_1),.dout(w_dff_B_WGIs6CrK3_1),.clk(gclk));
	jdff dff_B_NDHVr71m4_1(.din(w_dff_B_WGIs6CrK3_1),.dout(w_dff_B_NDHVr71m4_1),.clk(gclk));
	jdff dff_B_jU6j1S9I3_1(.din(w_dff_B_NDHVr71m4_1),.dout(w_dff_B_jU6j1S9I3_1),.clk(gclk));
	jdff dff_B_bBW133xo7_1(.din(w_dff_B_jU6j1S9I3_1),.dout(w_dff_B_bBW133xo7_1),.clk(gclk));
	jdff dff_B_j1gTpmQG3_1(.din(w_dff_B_bBW133xo7_1),.dout(w_dff_B_j1gTpmQG3_1),.clk(gclk));
	jdff dff_B_nu4wcaFe2_1(.din(w_dff_B_j1gTpmQG3_1),.dout(w_dff_B_nu4wcaFe2_1),.clk(gclk));
	jdff dff_B_d5ww5trd6_1(.din(w_dff_B_nu4wcaFe2_1),.dout(w_dff_B_d5ww5trd6_1),.clk(gclk));
	jdff dff_B_vxSjOymS8_1(.din(w_dff_B_d5ww5trd6_1),.dout(w_dff_B_vxSjOymS8_1),.clk(gclk));
	jdff dff_B_BLHDNoIe6_1(.din(w_dff_B_vxSjOymS8_1),.dout(w_dff_B_BLHDNoIe6_1),.clk(gclk));
	jdff dff_B_JjtDlUbO9_1(.din(w_dff_B_BLHDNoIe6_1),.dout(w_dff_B_JjtDlUbO9_1),.clk(gclk));
	jdff dff_B_caypdeIr4_1(.din(w_dff_B_JjtDlUbO9_1),.dout(w_dff_B_caypdeIr4_1),.clk(gclk));
	jdff dff_B_UcCUvmwO2_1(.din(w_dff_B_caypdeIr4_1),.dout(w_dff_B_UcCUvmwO2_1),.clk(gclk));
	jdff dff_B_VjqQEqSk0_1(.din(w_dff_B_UcCUvmwO2_1),.dout(w_dff_B_VjqQEqSk0_1),.clk(gclk));
	jdff dff_B_Z0I00MCQ1_1(.din(w_dff_B_VjqQEqSk0_1),.dout(w_dff_B_Z0I00MCQ1_1),.clk(gclk));
	jdff dff_B_CINVDIGM1_1(.din(w_dff_B_Z0I00MCQ1_1),.dout(w_dff_B_CINVDIGM1_1),.clk(gclk));
	jdff dff_B_caZpxfEV1_1(.din(w_dff_B_CINVDIGM1_1),.dout(w_dff_B_caZpxfEV1_1),.clk(gclk));
	jdff dff_B_xhE3hfVr6_1(.din(w_dff_B_caZpxfEV1_1),.dout(w_dff_B_xhE3hfVr6_1),.clk(gclk));
	jdff dff_B_DdifxwCM3_1(.din(w_dff_B_xhE3hfVr6_1),.dout(w_dff_B_DdifxwCM3_1),.clk(gclk));
	jdff dff_B_FI4q1Rkk4_1(.din(w_dff_B_DdifxwCM3_1),.dout(w_dff_B_FI4q1Rkk4_1),.clk(gclk));
	jdff dff_B_hkOWJ4OF2_1(.din(w_dff_B_FI4q1Rkk4_1),.dout(w_dff_B_hkOWJ4OF2_1),.clk(gclk));
	jdff dff_B_vLWd5O6c7_1(.din(w_dff_B_hkOWJ4OF2_1),.dout(w_dff_B_vLWd5O6c7_1),.clk(gclk));
	jdff dff_B_NZd7Lg3u7_1(.din(w_dff_B_vLWd5O6c7_1),.dout(w_dff_B_NZd7Lg3u7_1),.clk(gclk));
	jdff dff_B_0Jq5KK763_1(.din(w_dff_B_NZd7Lg3u7_1),.dout(w_dff_B_0Jq5KK763_1),.clk(gclk));
	jdff dff_B_CSNzOrFa7_1(.din(w_dff_B_0Jq5KK763_1),.dout(w_dff_B_CSNzOrFa7_1),.clk(gclk));
	jdff dff_B_aOAiC69s0_1(.din(w_dff_B_CSNzOrFa7_1),.dout(w_dff_B_aOAiC69s0_1),.clk(gclk));
	jdff dff_B_8cz2WsSi6_1(.din(w_dff_B_aOAiC69s0_1),.dout(w_dff_B_8cz2WsSi6_1),.clk(gclk));
	jdff dff_B_vNNqIT0k0_1(.din(w_dff_B_8cz2WsSi6_1),.dout(w_dff_B_vNNqIT0k0_1),.clk(gclk));
	jdff dff_B_am6QIwSN5_1(.din(w_dff_B_vNNqIT0k0_1),.dout(w_dff_B_am6QIwSN5_1),.clk(gclk));
	jdff dff_B_D7UeQCsY6_1(.din(w_dff_B_am6QIwSN5_1),.dout(w_dff_B_D7UeQCsY6_1),.clk(gclk));
	jdff dff_B_WcqaJ2jn3_1(.din(w_dff_B_D7UeQCsY6_1),.dout(w_dff_B_WcqaJ2jn3_1),.clk(gclk));
	jdff dff_B_it3M0FVM2_1(.din(w_dff_B_WcqaJ2jn3_1),.dout(w_dff_B_it3M0FVM2_1),.clk(gclk));
	jdff dff_B_SsrF3jtx4_1(.din(w_dff_B_it3M0FVM2_1),.dout(w_dff_B_SsrF3jtx4_1),.clk(gclk));
	jdff dff_B_5rekw1lX6_1(.din(w_dff_B_SsrF3jtx4_1),.dout(w_dff_B_5rekw1lX6_1),.clk(gclk));
	jdff dff_B_enA95C2F9_1(.din(w_dff_B_5rekw1lX6_1),.dout(w_dff_B_enA95C2F9_1),.clk(gclk));
	jdff dff_B_0LDZx56T0_1(.din(w_dff_B_enA95C2F9_1),.dout(w_dff_B_0LDZx56T0_1),.clk(gclk));
	jdff dff_B_LYGoZoG09_1(.din(w_dff_B_0LDZx56T0_1),.dout(w_dff_B_LYGoZoG09_1),.clk(gclk));
	jdff dff_B_2PWh1po04_1(.din(w_dff_B_LYGoZoG09_1),.dout(w_dff_B_2PWh1po04_1),.clk(gclk));
	jdff dff_B_3VfNJbtd4_1(.din(w_dff_B_2PWh1po04_1),.dout(w_dff_B_3VfNJbtd4_1),.clk(gclk));
	jdff dff_B_U3MKcYr33_1(.din(w_dff_B_3VfNJbtd4_1),.dout(w_dff_B_U3MKcYr33_1),.clk(gclk));
	jdff dff_B_JZl7bUXj2_1(.din(w_dff_B_U3MKcYr33_1),.dout(w_dff_B_JZl7bUXj2_1),.clk(gclk));
	jdff dff_B_EtMzor9e5_1(.din(w_dff_B_JZl7bUXj2_1),.dout(w_dff_B_EtMzor9e5_1),.clk(gclk));
	jdff dff_B_09753Men2_1(.din(w_dff_B_EtMzor9e5_1),.dout(w_dff_B_09753Men2_1),.clk(gclk));
	jdff dff_B_SRo4UDe63_1(.din(w_dff_B_09753Men2_1),.dout(w_dff_B_SRo4UDe63_1),.clk(gclk));
	jdff dff_B_TdRn8OID0_1(.din(w_dff_B_SRo4UDe63_1),.dout(w_dff_B_TdRn8OID0_1),.clk(gclk));
	jdff dff_B_9r3EyRnt9_1(.din(w_dff_B_TdRn8OID0_1),.dout(w_dff_B_9r3EyRnt9_1),.clk(gclk));
	jdff dff_B_RV449SGC0_1(.din(w_dff_B_9r3EyRnt9_1),.dout(w_dff_B_RV449SGC0_1),.clk(gclk));
	jdff dff_B_TrlzIL7K6_1(.din(w_dff_B_RV449SGC0_1),.dout(w_dff_B_TrlzIL7K6_1),.clk(gclk));
	jdff dff_B_Rv29iDqX4_1(.din(w_dff_B_TrlzIL7K6_1),.dout(w_dff_B_Rv29iDqX4_1),.clk(gclk));
	jdff dff_B_EY4FzuFX5_1(.din(w_dff_B_Rv29iDqX4_1),.dout(w_dff_B_EY4FzuFX5_1),.clk(gclk));
	jdff dff_B_TtaQ10hk0_1(.din(w_dff_B_EY4FzuFX5_1),.dout(w_dff_B_TtaQ10hk0_1),.clk(gclk));
	jdff dff_B_ndlMbPLS5_1(.din(w_dff_B_TtaQ10hk0_1),.dout(w_dff_B_ndlMbPLS5_1),.clk(gclk));
	jdff dff_B_GI8cjqgr1_1(.din(w_dff_B_ndlMbPLS5_1),.dout(w_dff_B_GI8cjqgr1_1),.clk(gclk));
	jdff dff_B_e6lz4nSd7_0(.din(n1003),.dout(w_dff_B_e6lz4nSd7_0),.clk(gclk));
	jdff dff_B_QP1HIkg01_0(.din(w_dff_B_e6lz4nSd7_0),.dout(w_dff_B_QP1HIkg01_0),.clk(gclk));
	jdff dff_B_ej58O5Cg7_0(.din(w_dff_B_QP1HIkg01_0),.dout(w_dff_B_ej58O5Cg7_0),.clk(gclk));
	jdff dff_B_c1OS9FIc1_0(.din(w_dff_B_ej58O5Cg7_0),.dout(w_dff_B_c1OS9FIc1_0),.clk(gclk));
	jdff dff_B_UxUQjaGq6_0(.din(w_dff_B_c1OS9FIc1_0),.dout(w_dff_B_UxUQjaGq6_0),.clk(gclk));
	jdff dff_B_3IGJFiRl8_0(.din(w_dff_B_UxUQjaGq6_0),.dout(w_dff_B_3IGJFiRl8_0),.clk(gclk));
	jdff dff_B_BYw3f24c1_0(.din(w_dff_B_3IGJFiRl8_0),.dout(w_dff_B_BYw3f24c1_0),.clk(gclk));
	jdff dff_B_GCMdQVue7_0(.din(w_dff_B_BYw3f24c1_0),.dout(w_dff_B_GCMdQVue7_0),.clk(gclk));
	jdff dff_B_joe4ZUSL2_0(.din(w_dff_B_GCMdQVue7_0),.dout(w_dff_B_joe4ZUSL2_0),.clk(gclk));
	jdff dff_B_WhWE3lOn2_0(.din(w_dff_B_joe4ZUSL2_0),.dout(w_dff_B_WhWE3lOn2_0),.clk(gclk));
	jdff dff_B_XHUCO0FG0_0(.din(w_dff_B_WhWE3lOn2_0),.dout(w_dff_B_XHUCO0FG0_0),.clk(gclk));
	jdff dff_B_QN1rs2GM8_0(.din(w_dff_B_XHUCO0FG0_0),.dout(w_dff_B_QN1rs2GM8_0),.clk(gclk));
	jdff dff_B_6zu9grEN8_0(.din(w_dff_B_QN1rs2GM8_0),.dout(w_dff_B_6zu9grEN8_0),.clk(gclk));
	jdff dff_B_A8dbrEFY8_0(.din(w_dff_B_6zu9grEN8_0),.dout(w_dff_B_A8dbrEFY8_0),.clk(gclk));
	jdff dff_B_75cvf8bH4_0(.din(w_dff_B_A8dbrEFY8_0),.dout(w_dff_B_75cvf8bH4_0),.clk(gclk));
	jdff dff_B_cKKOVBjd7_0(.din(w_dff_B_75cvf8bH4_0),.dout(w_dff_B_cKKOVBjd7_0),.clk(gclk));
	jdff dff_B_qtYDwSyy0_0(.din(w_dff_B_cKKOVBjd7_0),.dout(w_dff_B_qtYDwSyy0_0),.clk(gclk));
	jdff dff_B_YVmHd4Qa5_0(.din(w_dff_B_qtYDwSyy0_0),.dout(w_dff_B_YVmHd4Qa5_0),.clk(gclk));
	jdff dff_B_uzPZcTdB4_0(.din(w_dff_B_YVmHd4Qa5_0),.dout(w_dff_B_uzPZcTdB4_0),.clk(gclk));
	jdff dff_B_LrDCyk2e9_0(.din(w_dff_B_uzPZcTdB4_0),.dout(w_dff_B_LrDCyk2e9_0),.clk(gclk));
	jdff dff_B_22TBqFiZ7_0(.din(w_dff_B_LrDCyk2e9_0),.dout(w_dff_B_22TBqFiZ7_0),.clk(gclk));
	jdff dff_B_uOgljo4N5_0(.din(w_dff_B_22TBqFiZ7_0),.dout(w_dff_B_uOgljo4N5_0),.clk(gclk));
	jdff dff_B_YmNN57yQ9_0(.din(w_dff_B_uOgljo4N5_0),.dout(w_dff_B_YmNN57yQ9_0),.clk(gclk));
	jdff dff_B_Q2Omy1N32_0(.din(w_dff_B_YmNN57yQ9_0),.dout(w_dff_B_Q2Omy1N32_0),.clk(gclk));
	jdff dff_B_p3PFj3k72_0(.din(w_dff_B_Q2Omy1N32_0),.dout(w_dff_B_p3PFj3k72_0),.clk(gclk));
	jdff dff_B_xnokRXv86_0(.din(w_dff_B_p3PFj3k72_0),.dout(w_dff_B_xnokRXv86_0),.clk(gclk));
	jdff dff_B_Vo3ZFT8P1_0(.din(w_dff_B_xnokRXv86_0),.dout(w_dff_B_Vo3ZFT8P1_0),.clk(gclk));
	jdff dff_B_XSpMbBMq5_0(.din(w_dff_B_Vo3ZFT8P1_0),.dout(w_dff_B_XSpMbBMq5_0),.clk(gclk));
	jdff dff_B_eSd5pEHh6_0(.din(w_dff_B_XSpMbBMq5_0),.dout(w_dff_B_eSd5pEHh6_0),.clk(gclk));
	jdff dff_B_qiRjCs3g2_0(.din(w_dff_B_eSd5pEHh6_0),.dout(w_dff_B_qiRjCs3g2_0),.clk(gclk));
	jdff dff_B_M9DkvZxp0_0(.din(w_dff_B_qiRjCs3g2_0),.dout(w_dff_B_M9DkvZxp0_0),.clk(gclk));
	jdff dff_B_W4DMuDQH8_0(.din(w_dff_B_M9DkvZxp0_0),.dout(w_dff_B_W4DMuDQH8_0),.clk(gclk));
	jdff dff_B_2bo03jgs9_0(.din(w_dff_B_W4DMuDQH8_0),.dout(w_dff_B_2bo03jgs9_0),.clk(gclk));
	jdff dff_B_WLNjEQDx7_0(.din(w_dff_B_2bo03jgs9_0),.dout(w_dff_B_WLNjEQDx7_0),.clk(gclk));
	jdff dff_B_I4SY4MPK0_0(.din(w_dff_B_WLNjEQDx7_0),.dout(w_dff_B_I4SY4MPK0_0),.clk(gclk));
	jdff dff_B_fJliKFbw1_0(.din(w_dff_B_I4SY4MPK0_0),.dout(w_dff_B_fJliKFbw1_0),.clk(gclk));
	jdff dff_B_MisHAYvD7_0(.din(w_dff_B_fJliKFbw1_0),.dout(w_dff_B_MisHAYvD7_0),.clk(gclk));
	jdff dff_B_Pa2q46Wb6_0(.din(w_dff_B_MisHAYvD7_0),.dout(w_dff_B_Pa2q46Wb6_0),.clk(gclk));
	jdff dff_B_OMLl9mby1_0(.din(w_dff_B_Pa2q46Wb6_0),.dout(w_dff_B_OMLl9mby1_0),.clk(gclk));
	jdff dff_B_ezRSevQT2_0(.din(w_dff_B_OMLl9mby1_0),.dout(w_dff_B_ezRSevQT2_0),.clk(gclk));
	jdff dff_B_iJCBvH4N1_0(.din(w_dff_B_ezRSevQT2_0),.dout(w_dff_B_iJCBvH4N1_0),.clk(gclk));
	jdff dff_B_hzOjO8wT3_0(.din(w_dff_B_iJCBvH4N1_0),.dout(w_dff_B_hzOjO8wT3_0),.clk(gclk));
	jdff dff_B_vZED4JAN8_0(.din(w_dff_B_hzOjO8wT3_0),.dout(w_dff_B_vZED4JAN8_0),.clk(gclk));
	jdff dff_B_BpALgirx8_0(.din(w_dff_B_vZED4JAN8_0),.dout(w_dff_B_BpALgirx8_0),.clk(gclk));
	jdff dff_B_eKWoX3Js4_0(.din(w_dff_B_BpALgirx8_0),.dout(w_dff_B_eKWoX3Js4_0),.clk(gclk));
	jdff dff_B_oxXNSdov8_0(.din(w_dff_B_eKWoX3Js4_0),.dout(w_dff_B_oxXNSdov8_0),.clk(gclk));
	jdff dff_B_L5epyQPQ9_0(.din(w_dff_B_oxXNSdov8_0),.dout(w_dff_B_L5epyQPQ9_0),.clk(gclk));
	jdff dff_B_QOkAJBUi8_0(.din(w_dff_B_L5epyQPQ9_0),.dout(w_dff_B_QOkAJBUi8_0),.clk(gclk));
	jdff dff_B_VmPocXDV2_0(.din(w_dff_B_QOkAJBUi8_0),.dout(w_dff_B_VmPocXDV2_0),.clk(gclk));
	jdff dff_B_CSBB6bv62_0(.din(w_dff_B_VmPocXDV2_0),.dout(w_dff_B_CSBB6bv62_0),.clk(gclk));
	jdff dff_B_1yL7wUaL1_0(.din(w_dff_B_CSBB6bv62_0),.dout(w_dff_B_1yL7wUaL1_0),.clk(gclk));
	jdff dff_B_v3NoQaqj4_0(.din(w_dff_B_1yL7wUaL1_0),.dout(w_dff_B_v3NoQaqj4_0),.clk(gclk));
	jdff dff_B_YZYvtNtZ8_0(.din(w_dff_B_v3NoQaqj4_0),.dout(w_dff_B_YZYvtNtZ8_0),.clk(gclk));
	jdff dff_B_ePVZN5wl8_0(.din(w_dff_B_YZYvtNtZ8_0),.dout(w_dff_B_ePVZN5wl8_0),.clk(gclk));
	jdff dff_B_kLgxzR3X1_0(.din(w_dff_B_ePVZN5wl8_0),.dout(w_dff_B_kLgxzR3X1_0),.clk(gclk));
	jdff dff_B_xGpjraOR2_0(.din(w_dff_B_kLgxzR3X1_0),.dout(w_dff_B_xGpjraOR2_0),.clk(gclk));
	jdff dff_B_iXyjUXoo0_0(.din(w_dff_B_xGpjraOR2_0),.dout(w_dff_B_iXyjUXoo0_0),.clk(gclk));
	jdff dff_B_fmJptW6U6_0(.din(w_dff_B_iXyjUXoo0_0),.dout(w_dff_B_fmJptW6U6_0),.clk(gclk));
	jdff dff_B_e2nzqi1Y5_0(.din(w_dff_B_fmJptW6U6_0),.dout(w_dff_B_e2nzqi1Y5_0),.clk(gclk));
	jdff dff_B_TakbssWp7_0(.din(w_dff_B_e2nzqi1Y5_0),.dout(w_dff_B_TakbssWp7_0),.clk(gclk));
	jdff dff_B_zW8bEz0W9_0(.din(w_dff_B_TakbssWp7_0),.dout(w_dff_B_zW8bEz0W9_0),.clk(gclk));
	jdff dff_B_vOcimzpI5_0(.din(w_dff_B_zW8bEz0W9_0),.dout(w_dff_B_vOcimzpI5_0),.clk(gclk));
	jdff dff_B_ra5hyIxk1_0(.din(w_dff_B_vOcimzpI5_0),.dout(w_dff_B_ra5hyIxk1_0),.clk(gclk));
	jdff dff_B_j9rX7nar7_0(.din(w_dff_B_ra5hyIxk1_0),.dout(w_dff_B_j9rX7nar7_0),.clk(gclk));
	jdff dff_B_ii5VuVHj2_0(.din(w_dff_B_j9rX7nar7_0),.dout(w_dff_B_ii5VuVHj2_0),.clk(gclk));
	jdff dff_B_KvW3IjMc5_0(.din(w_dff_B_ii5VuVHj2_0),.dout(w_dff_B_KvW3IjMc5_0),.clk(gclk));
	jdff dff_B_ILjjkCgc1_0(.din(w_dff_B_KvW3IjMc5_0),.dout(w_dff_B_ILjjkCgc1_0),.clk(gclk));
	jdff dff_B_OSjB8WzJ2_0(.din(w_dff_B_ILjjkCgc1_0),.dout(w_dff_B_OSjB8WzJ2_0),.clk(gclk));
	jdff dff_B_FSfjnVL29_0(.din(w_dff_B_OSjB8WzJ2_0),.dout(w_dff_B_FSfjnVL29_0),.clk(gclk));
	jdff dff_B_EkDOfp9y1_0(.din(w_dff_B_FSfjnVL29_0),.dout(w_dff_B_EkDOfp9y1_0),.clk(gclk));
	jdff dff_B_Iiumm3eR9_0(.din(w_dff_B_EkDOfp9y1_0),.dout(w_dff_B_Iiumm3eR9_0),.clk(gclk));
	jdff dff_B_z4Gd4soa7_0(.din(w_dff_B_Iiumm3eR9_0),.dout(w_dff_B_z4Gd4soa7_0),.clk(gclk));
	jdff dff_B_BKECVXw49_0(.din(w_dff_B_z4Gd4soa7_0),.dout(w_dff_B_BKECVXw49_0),.clk(gclk));
	jdff dff_B_6I1gYRnV6_0(.din(w_dff_B_BKECVXw49_0),.dout(w_dff_B_6I1gYRnV6_0),.clk(gclk));
	jdff dff_B_yhQaCsgT9_0(.din(w_dff_B_6I1gYRnV6_0),.dout(w_dff_B_yhQaCsgT9_0),.clk(gclk));
	jdff dff_B_T3heKXXc3_0(.din(w_dff_B_yhQaCsgT9_0),.dout(w_dff_B_T3heKXXc3_0),.clk(gclk));
	jdff dff_B_VAsiJoMd5_0(.din(w_dff_B_T3heKXXc3_0),.dout(w_dff_B_VAsiJoMd5_0),.clk(gclk));
	jdff dff_B_18tnDX7V4_0(.din(w_dff_B_VAsiJoMd5_0),.dout(w_dff_B_18tnDX7V4_0),.clk(gclk));
	jdff dff_B_MtOzHtfH3_0(.din(w_dff_B_18tnDX7V4_0),.dout(w_dff_B_MtOzHtfH3_0),.clk(gclk));
	jdff dff_B_QprVbgpW7_0(.din(w_dff_B_MtOzHtfH3_0),.dout(w_dff_B_QprVbgpW7_0),.clk(gclk));
	jdff dff_B_P2XHdSjZ6_0(.din(w_dff_B_QprVbgpW7_0),.dout(w_dff_B_P2XHdSjZ6_0),.clk(gclk));
	jdff dff_B_kRXfaSXs7_0(.din(w_dff_B_P2XHdSjZ6_0),.dout(w_dff_B_kRXfaSXs7_0),.clk(gclk));
	jdff dff_B_eAO4Gal12_0(.din(w_dff_B_kRXfaSXs7_0),.dout(w_dff_B_eAO4Gal12_0),.clk(gclk));
	jdff dff_B_ZsIhPlMI7_0(.din(w_dff_B_eAO4Gal12_0),.dout(w_dff_B_ZsIhPlMI7_0),.clk(gclk));
	jdff dff_B_Pj30zCB80_0(.din(w_dff_B_ZsIhPlMI7_0),.dout(w_dff_B_Pj30zCB80_0),.clk(gclk));
	jdff dff_B_AZ6NrpXW4_0(.din(w_dff_B_Pj30zCB80_0),.dout(w_dff_B_AZ6NrpXW4_0),.clk(gclk));
	jdff dff_B_6Lf2J6yg9_0(.din(w_dff_B_AZ6NrpXW4_0),.dout(w_dff_B_6Lf2J6yg9_0),.clk(gclk));
	jdff dff_B_DcjTsauK2_0(.din(w_dff_B_6Lf2J6yg9_0),.dout(w_dff_B_DcjTsauK2_0),.clk(gclk));
	jdff dff_B_rjautiqH2_0(.din(w_dff_B_DcjTsauK2_0),.dout(w_dff_B_rjautiqH2_0),.clk(gclk));
	jdff dff_B_jnCsBWIj1_0(.din(w_dff_B_rjautiqH2_0),.dout(w_dff_B_jnCsBWIj1_0),.clk(gclk));
	jdff dff_B_aGNge5uQ5_0(.din(w_dff_B_jnCsBWIj1_0),.dout(w_dff_B_aGNge5uQ5_0),.clk(gclk));
	jdff dff_B_RDjbSkuj4_0(.din(w_dff_B_aGNge5uQ5_0),.dout(w_dff_B_RDjbSkuj4_0),.clk(gclk));
	jdff dff_B_MpVggaHh6_0(.din(w_dff_B_RDjbSkuj4_0),.dout(w_dff_B_MpVggaHh6_0),.clk(gclk));
	jdff dff_B_4Ys50if07_0(.din(w_dff_B_MpVggaHh6_0),.dout(w_dff_B_4Ys50if07_0),.clk(gclk));
	jdff dff_B_i1o0bDT82_0(.din(w_dff_B_4Ys50if07_0),.dout(w_dff_B_i1o0bDT82_0),.clk(gclk));
	jdff dff_B_YniSy8aB5_0(.din(w_dff_B_i1o0bDT82_0),.dout(w_dff_B_YniSy8aB5_0),.clk(gclk));
	jdff dff_B_lck7UEvD2_0(.din(w_dff_B_YniSy8aB5_0),.dout(w_dff_B_lck7UEvD2_0),.clk(gclk));
	jdff dff_B_VU70DES38_0(.din(w_dff_B_lck7UEvD2_0),.dout(w_dff_B_VU70DES38_0),.clk(gclk));
	jdff dff_B_X0285ssm4_0(.din(w_dff_B_VU70DES38_0),.dout(w_dff_B_X0285ssm4_0),.clk(gclk));
	jdff dff_B_ms0rmQyj3_0(.din(w_dff_B_X0285ssm4_0),.dout(w_dff_B_ms0rmQyj3_0),.clk(gclk));
	jdff dff_B_CyFTqv8S8_0(.din(w_dff_B_ms0rmQyj3_0),.dout(w_dff_B_CyFTqv8S8_0),.clk(gclk));
	jdff dff_B_ap8PWfKR3_0(.din(w_dff_B_CyFTqv8S8_0),.dout(w_dff_B_ap8PWfKR3_0),.clk(gclk));
	jdff dff_B_ISBRX9kG4_0(.din(w_dff_B_ap8PWfKR3_0),.dout(w_dff_B_ISBRX9kG4_0),.clk(gclk));
	jdff dff_B_Uc08YVKY5_1(.din(n996),.dout(w_dff_B_Uc08YVKY5_1),.clk(gclk));
	jdff dff_B_JNr4uM3S9_1(.din(w_dff_B_Uc08YVKY5_1),.dout(w_dff_B_JNr4uM3S9_1),.clk(gclk));
	jdff dff_B_9h76yTlC5_1(.din(w_dff_B_JNr4uM3S9_1),.dout(w_dff_B_9h76yTlC5_1),.clk(gclk));
	jdff dff_B_Y0ZwGY1U7_1(.din(w_dff_B_9h76yTlC5_1),.dout(w_dff_B_Y0ZwGY1U7_1),.clk(gclk));
	jdff dff_B_Jlfr7Qml8_1(.din(w_dff_B_Y0ZwGY1U7_1),.dout(w_dff_B_Jlfr7Qml8_1),.clk(gclk));
	jdff dff_B_gM9vXp6G5_1(.din(w_dff_B_Jlfr7Qml8_1),.dout(w_dff_B_gM9vXp6G5_1),.clk(gclk));
	jdff dff_B_kRwJcoUK7_1(.din(w_dff_B_gM9vXp6G5_1),.dout(w_dff_B_kRwJcoUK7_1),.clk(gclk));
	jdff dff_B_u1EZgqHf5_1(.din(w_dff_B_kRwJcoUK7_1),.dout(w_dff_B_u1EZgqHf5_1),.clk(gclk));
	jdff dff_B_ushofyMb6_1(.din(w_dff_B_u1EZgqHf5_1),.dout(w_dff_B_ushofyMb6_1),.clk(gclk));
	jdff dff_B_rpfBrktU3_1(.din(w_dff_B_ushofyMb6_1),.dout(w_dff_B_rpfBrktU3_1),.clk(gclk));
	jdff dff_B_w8AP4Hsl0_1(.din(w_dff_B_rpfBrktU3_1),.dout(w_dff_B_w8AP4Hsl0_1),.clk(gclk));
	jdff dff_B_Ktjdo2Ns7_1(.din(w_dff_B_w8AP4Hsl0_1),.dout(w_dff_B_Ktjdo2Ns7_1),.clk(gclk));
	jdff dff_B_9Pr1Z7lQ3_1(.din(w_dff_B_Ktjdo2Ns7_1),.dout(w_dff_B_9Pr1Z7lQ3_1),.clk(gclk));
	jdff dff_B_KnE6zQED7_1(.din(w_dff_B_9Pr1Z7lQ3_1),.dout(w_dff_B_KnE6zQED7_1),.clk(gclk));
	jdff dff_B_3waKnxTt1_1(.din(w_dff_B_KnE6zQED7_1),.dout(w_dff_B_3waKnxTt1_1),.clk(gclk));
	jdff dff_B_DA1DP4Xd1_1(.din(w_dff_B_3waKnxTt1_1),.dout(w_dff_B_DA1DP4Xd1_1),.clk(gclk));
	jdff dff_B_MWTz8cpq3_1(.din(w_dff_B_DA1DP4Xd1_1),.dout(w_dff_B_MWTz8cpq3_1),.clk(gclk));
	jdff dff_B_eiujRRXT5_1(.din(w_dff_B_MWTz8cpq3_1),.dout(w_dff_B_eiujRRXT5_1),.clk(gclk));
	jdff dff_B_nhnZyIlb3_1(.din(w_dff_B_eiujRRXT5_1),.dout(w_dff_B_nhnZyIlb3_1),.clk(gclk));
	jdff dff_B_PKKnjG4f4_1(.din(w_dff_B_nhnZyIlb3_1),.dout(w_dff_B_PKKnjG4f4_1),.clk(gclk));
	jdff dff_B_QIQrqbdL7_1(.din(w_dff_B_PKKnjG4f4_1),.dout(w_dff_B_QIQrqbdL7_1),.clk(gclk));
	jdff dff_B_F0X5ybIW2_1(.din(w_dff_B_QIQrqbdL7_1),.dout(w_dff_B_F0X5ybIW2_1),.clk(gclk));
	jdff dff_B_nVXWQ8082_1(.din(w_dff_B_F0X5ybIW2_1),.dout(w_dff_B_nVXWQ8082_1),.clk(gclk));
	jdff dff_B_I7uVEbnw8_1(.din(w_dff_B_nVXWQ8082_1),.dout(w_dff_B_I7uVEbnw8_1),.clk(gclk));
	jdff dff_B_ER6QXdeH7_1(.din(w_dff_B_I7uVEbnw8_1),.dout(w_dff_B_ER6QXdeH7_1),.clk(gclk));
	jdff dff_B_SqcqtdqA5_1(.din(w_dff_B_ER6QXdeH7_1),.dout(w_dff_B_SqcqtdqA5_1),.clk(gclk));
	jdff dff_B_iaPnzZ829_1(.din(w_dff_B_SqcqtdqA5_1),.dout(w_dff_B_iaPnzZ829_1),.clk(gclk));
	jdff dff_B_J5R3M07j5_1(.din(w_dff_B_iaPnzZ829_1),.dout(w_dff_B_J5R3M07j5_1),.clk(gclk));
	jdff dff_B_8n1HrsKJ1_1(.din(w_dff_B_J5R3M07j5_1),.dout(w_dff_B_8n1HrsKJ1_1),.clk(gclk));
	jdff dff_B_AtOdfwoZ3_1(.din(w_dff_B_8n1HrsKJ1_1),.dout(w_dff_B_AtOdfwoZ3_1),.clk(gclk));
	jdff dff_B_mVlI4WCx0_1(.din(w_dff_B_AtOdfwoZ3_1),.dout(w_dff_B_mVlI4WCx0_1),.clk(gclk));
	jdff dff_B_GvCzs7de9_1(.din(w_dff_B_mVlI4WCx0_1),.dout(w_dff_B_GvCzs7de9_1),.clk(gclk));
	jdff dff_B_xpU7rWtj2_1(.din(w_dff_B_GvCzs7de9_1),.dout(w_dff_B_xpU7rWtj2_1),.clk(gclk));
	jdff dff_B_7ZeUikwx8_1(.din(w_dff_B_xpU7rWtj2_1),.dout(w_dff_B_7ZeUikwx8_1),.clk(gclk));
	jdff dff_B_HlQd3npy0_1(.din(w_dff_B_7ZeUikwx8_1),.dout(w_dff_B_HlQd3npy0_1),.clk(gclk));
	jdff dff_B_timINsCF3_1(.din(w_dff_B_HlQd3npy0_1),.dout(w_dff_B_timINsCF3_1),.clk(gclk));
	jdff dff_B_DXrU1c7V2_1(.din(w_dff_B_timINsCF3_1),.dout(w_dff_B_DXrU1c7V2_1),.clk(gclk));
	jdff dff_B_GeIx1So29_1(.din(w_dff_B_DXrU1c7V2_1),.dout(w_dff_B_GeIx1So29_1),.clk(gclk));
	jdff dff_B_hdMRwFTk8_1(.din(w_dff_B_GeIx1So29_1),.dout(w_dff_B_hdMRwFTk8_1),.clk(gclk));
	jdff dff_B_3fpwr5H99_1(.din(w_dff_B_hdMRwFTk8_1),.dout(w_dff_B_3fpwr5H99_1),.clk(gclk));
	jdff dff_B_V8LVNEXd4_1(.din(w_dff_B_3fpwr5H99_1),.dout(w_dff_B_V8LVNEXd4_1),.clk(gclk));
	jdff dff_B_nsx127bK8_1(.din(w_dff_B_V8LVNEXd4_1),.dout(w_dff_B_nsx127bK8_1),.clk(gclk));
	jdff dff_B_uJq1wClp0_1(.din(w_dff_B_nsx127bK8_1),.dout(w_dff_B_uJq1wClp0_1),.clk(gclk));
	jdff dff_B_z0YzCurh0_1(.din(w_dff_B_uJq1wClp0_1),.dout(w_dff_B_z0YzCurh0_1),.clk(gclk));
	jdff dff_B_qGAIjcRr7_1(.din(w_dff_B_z0YzCurh0_1),.dout(w_dff_B_qGAIjcRr7_1),.clk(gclk));
	jdff dff_B_xPHGV7GV4_1(.din(w_dff_B_qGAIjcRr7_1),.dout(w_dff_B_xPHGV7GV4_1),.clk(gclk));
	jdff dff_B_DUlgI1nE0_1(.din(w_dff_B_xPHGV7GV4_1),.dout(w_dff_B_DUlgI1nE0_1),.clk(gclk));
	jdff dff_B_wa9rmqy67_1(.din(w_dff_B_DUlgI1nE0_1),.dout(w_dff_B_wa9rmqy67_1),.clk(gclk));
	jdff dff_B_DqfPtgYI7_1(.din(w_dff_B_wa9rmqy67_1),.dout(w_dff_B_DqfPtgYI7_1),.clk(gclk));
	jdff dff_B_YK0ZpN1t9_1(.din(w_dff_B_DqfPtgYI7_1),.dout(w_dff_B_YK0ZpN1t9_1),.clk(gclk));
	jdff dff_B_w6EAt5FU2_1(.din(w_dff_B_YK0ZpN1t9_1),.dout(w_dff_B_w6EAt5FU2_1),.clk(gclk));
	jdff dff_B_QzbbztSb7_1(.din(w_dff_B_w6EAt5FU2_1),.dout(w_dff_B_QzbbztSb7_1),.clk(gclk));
	jdff dff_B_AT81xLg10_1(.din(w_dff_B_QzbbztSb7_1),.dout(w_dff_B_AT81xLg10_1),.clk(gclk));
	jdff dff_B_9MNWekpF7_1(.din(w_dff_B_AT81xLg10_1),.dout(w_dff_B_9MNWekpF7_1),.clk(gclk));
	jdff dff_B_FS5iXezl4_1(.din(w_dff_B_9MNWekpF7_1),.dout(w_dff_B_FS5iXezl4_1),.clk(gclk));
	jdff dff_B_k6rbrxsV2_1(.din(w_dff_B_FS5iXezl4_1),.dout(w_dff_B_k6rbrxsV2_1),.clk(gclk));
	jdff dff_B_YFAysJ3K5_1(.din(w_dff_B_k6rbrxsV2_1),.dout(w_dff_B_YFAysJ3K5_1),.clk(gclk));
	jdff dff_B_YHznMhmx8_1(.din(w_dff_B_YFAysJ3K5_1),.dout(w_dff_B_YHznMhmx8_1),.clk(gclk));
	jdff dff_B_E5LZrr773_1(.din(w_dff_B_YHznMhmx8_1),.dout(w_dff_B_E5LZrr773_1),.clk(gclk));
	jdff dff_B_8XugjQEe6_1(.din(w_dff_B_E5LZrr773_1),.dout(w_dff_B_8XugjQEe6_1),.clk(gclk));
	jdff dff_B_YGeeYzEU1_1(.din(w_dff_B_8XugjQEe6_1),.dout(w_dff_B_YGeeYzEU1_1),.clk(gclk));
	jdff dff_B_f02OrG1J2_1(.din(w_dff_B_YGeeYzEU1_1),.dout(w_dff_B_f02OrG1J2_1),.clk(gclk));
	jdff dff_B_hr9zR0DI5_1(.din(w_dff_B_f02OrG1J2_1),.dout(w_dff_B_hr9zR0DI5_1),.clk(gclk));
	jdff dff_B_O2uIn6pg7_1(.din(w_dff_B_hr9zR0DI5_1),.dout(w_dff_B_O2uIn6pg7_1),.clk(gclk));
	jdff dff_B_Sl5BtnIU1_1(.din(w_dff_B_O2uIn6pg7_1),.dout(w_dff_B_Sl5BtnIU1_1),.clk(gclk));
	jdff dff_B_ntE6AoX12_1(.din(w_dff_B_Sl5BtnIU1_1),.dout(w_dff_B_ntE6AoX12_1),.clk(gclk));
	jdff dff_B_anVdO9Di7_1(.din(w_dff_B_ntE6AoX12_1),.dout(w_dff_B_anVdO9Di7_1),.clk(gclk));
	jdff dff_B_KtpZAMZl6_1(.din(w_dff_B_anVdO9Di7_1),.dout(w_dff_B_KtpZAMZl6_1),.clk(gclk));
	jdff dff_B_PQoiDZgy6_1(.din(w_dff_B_KtpZAMZl6_1),.dout(w_dff_B_PQoiDZgy6_1),.clk(gclk));
	jdff dff_B_2hYxQ0tg1_1(.din(w_dff_B_PQoiDZgy6_1),.dout(w_dff_B_2hYxQ0tg1_1),.clk(gclk));
	jdff dff_B_31yiIhMV2_1(.din(w_dff_B_2hYxQ0tg1_1),.dout(w_dff_B_31yiIhMV2_1),.clk(gclk));
	jdff dff_B_c0EmdxH57_1(.din(w_dff_B_31yiIhMV2_1),.dout(w_dff_B_c0EmdxH57_1),.clk(gclk));
	jdff dff_B_vptXheoI2_1(.din(w_dff_B_c0EmdxH57_1),.dout(w_dff_B_vptXheoI2_1),.clk(gclk));
	jdff dff_B_nXwVgPLW3_1(.din(w_dff_B_vptXheoI2_1),.dout(w_dff_B_nXwVgPLW3_1),.clk(gclk));
	jdff dff_B_JuDNfIgZ0_1(.din(w_dff_B_nXwVgPLW3_1),.dout(w_dff_B_JuDNfIgZ0_1),.clk(gclk));
	jdff dff_B_ozJvyKhd1_1(.din(w_dff_B_JuDNfIgZ0_1),.dout(w_dff_B_ozJvyKhd1_1),.clk(gclk));
	jdff dff_B_nqLzc8YF2_1(.din(w_dff_B_ozJvyKhd1_1),.dout(w_dff_B_nqLzc8YF2_1),.clk(gclk));
	jdff dff_B_VftNLq0q5_1(.din(w_dff_B_nqLzc8YF2_1),.dout(w_dff_B_VftNLq0q5_1),.clk(gclk));
	jdff dff_B_4wMeMZnu6_1(.din(w_dff_B_VftNLq0q5_1),.dout(w_dff_B_4wMeMZnu6_1),.clk(gclk));
	jdff dff_B_KKWyLyDV6_1(.din(w_dff_B_4wMeMZnu6_1),.dout(w_dff_B_KKWyLyDV6_1),.clk(gclk));
	jdff dff_B_R8iTdVWC7_1(.din(w_dff_B_KKWyLyDV6_1),.dout(w_dff_B_R8iTdVWC7_1),.clk(gclk));
	jdff dff_B_S0zR8KcJ7_1(.din(w_dff_B_R8iTdVWC7_1),.dout(w_dff_B_S0zR8KcJ7_1),.clk(gclk));
	jdff dff_B_UBVTSTPL7_1(.din(w_dff_B_S0zR8KcJ7_1),.dout(w_dff_B_UBVTSTPL7_1),.clk(gclk));
	jdff dff_B_8YY9fMqH0_1(.din(w_dff_B_UBVTSTPL7_1),.dout(w_dff_B_8YY9fMqH0_1),.clk(gclk));
	jdff dff_B_0oEdJGk36_1(.din(w_dff_B_8YY9fMqH0_1),.dout(w_dff_B_0oEdJGk36_1),.clk(gclk));
	jdff dff_B_o4qTf8jB5_1(.din(w_dff_B_0oEdJGk36_1),.dout(w_dff_B_o4qTf8jB5_1),.clk(gclk));
	jdff dff_B_MPDSEuom9_1(.din(w_dff_B_o4qTf8jB5_1),.dout(w_dff_B_MPDSEuom9_1),.clk(gclk));
	jdff dff_B_c8ylioBm9_1(.din(w_dff_B_MPDSEuom9_1),.dout(w_dff_B_c8ylioBm9_1),.clk(gclk));
	jdff dff_B_nWFNcPuy9_1(.din(w_dff_B_c8ylioBm9_1),.dout(w_dff_B_nWFNcPuy9_1),.clk(gclk));
	jdff dff_B_0SwTFmC67_1(.din(w_dff_B_nWFNcPuy9_1),.dout(w_dff_B_0SwTFmC67_1),.clk(gclk));
	jdff dff_B_CeOU4EFo6_1(.din(w_dff_B_0SwTFmC67_1),.dout(w_dff_B_CeOU4EFo6_1),.clk(gclk));
	jdff dff_B_UY8LQKXX4_1(.din(w_dff_B_CeOU4EFo6_1),.dout(w_dff_B_UY8LQKXX4_1),.clk(gclk));
	jdff dff_B_fno0KeT45_1(.din(w_dff_B_UY8LQKXX4_1),.dout(w_dff_B_fno0KeT45_1),.clk(gclk));
	jdff dff_B_JlRKt4Hh9_1(.din(w_dff_B_fno0KeT45_1),.dout(w_dff_B_JlRKt4Hh9_1),.clk(gclk));
	jdff dff_B_v3VyVP3u6_1(.din(w_dff_B_JlRKt4Hh9_1),.dout(w_dff_B_v3VyVP3u6_1),.clk(gclk));
	jdff dff_B_0VnddscN1_1(.din(w_dff_B_v3VyVP3u6_1),.dout(w_dff_B_0VnddscN1_1),.clk(gclk));
	jdff dff_B_YQVrJRo68_1(.din(w_dff_B_0VnddscN1_1),.dout(w_dff_B_YQVrJRo68_1),.clk(gclk));
	jdff dff_B_MQ8eRaQ16_1(.din(w_dff_B_YQVrJRo68_1),.dout(w_dff_B_MQ8eRaQ16_1),.clk(gclk));
	jdff dff_B_Q2hFncA24_1(.din(w_dff_B_MQ8eRaQ16_1),.dout(w_dff_B_Q2hFncA24_1),.clk(gclk));
	jdff dff_B_90HziY8o0_1(.din(w_dff_B_Q2hFncA24_1),.dout(w_dff_B_90HziY8o0_1),.clk(gclk));
	jdff dff_B_R7LC8kK87_1(.din(w_dff_B_90HziY8o0_1),.dout(w_dff_B_R7LC8kK87_1),.clk(gclk));
	jdff dff_B_CTOAbFb57_1(.din(w_dff_B_R7LC8kK87_1),.dout(w_dff_B_CTOAbFb57_1),.clk(gclk));
	jdff dff_B_2DMqRswL7_0(.din(n997),.dout(w_dff_B_2DMqRswL7_0),.clk(gclk));
	jdff dff_B_xBuCHRR42_0(.din(w_dff_B_2DMqRswL7_0),.dout(w_dff_B_xBuCHRR42_0),.clk(gclk));
	jdff dff_B_XKbh560A8_0(.din(w_dff_B_xBuCHRR42_0),.dout(w_dff_B_XKbh560A8_0),.clk(gclk));
	jdff dff_B_lKBUYmLM9_0(.din(w_dff_B_XKbh560A8_0),.dout(w_dff_B_lKBUYmLM9_0),.clk(gclk));
	jdff dff_B_ScFiBwxj0_0(.din(w_dff_B_lKBUYmLM9_0),.dout(w_dff_B_ScFiBwxj0_0),.clk(gclk));
	jdff dff_B_YcTdU1gp2_0(.din(w_dff_B_ScFiBwxj0_0),.dout(w_dff_B_YcTdU1gp2_0),.clk(gclk));
	jdff dff_B_GJAjsNRd6_0(.din(w_dff_B_YcTdU1gp2_0),.dout(w_dff_B_GJAjsNRd6_0),.clk(gclk));
	jdff dff_B_MfxeiVbI4_0(.din(w_dff_B_GJAjsNRd6_0),.dout(w_dff_B_MfxeiVbI4_0),.clk(gclk));
	jdff dff_B_QcEt8eNG0_0(.din(w_dff_B_MfxeiVbI4_0),.dout(w_dff_B_QcEt8eNG0_0),.clk(gclk));
	jdff dff_B_7x8H3DV25_0(.din(w_dff_B_QcEt8eNG0_0),.dout(w_dff_B_7x8H3DV25_0),.clk(gclk));
	jdff dff_B_aekMSfWk4_0(.din(w_dff_B_7x8H3DV25_0),.dout(w_dff_B_aekMSfWk4_0),.clk(gclk));
	jdff dff_B_KXjnSbXn0_0(.din(w_dff_B_aekMSfWk4_0),.dout(w_dff_B_KXjnSbXn0_0),.clk(gclk));
	jdff dff_B_J1nJZVwh3_0(.din(w_dff_B_KXjnSbXn0_0),.dout(w_dff_B_J1nJZVwh3_0),.clk(gclk));
	jdff dff_B_qHR0xegx2_0(.din(w_dff_B_J1nJZVwh3_0),.dout(w_dff_B_qHR0xegx2_0),.clk(gclk));
	jdff dff_B_bOy7XOuS1_0(.din(w_dff_B_qHR0xegx2_0),.dout(w_dff_B_bOy7XOuS1_0),.clk(gclk));
	jdff dff_B_ypOF11ny7_0(.din(w_dff_B_bOy7XOuS1_0),.dout(w_dff_B_ypOF11ny7_0),.clk(gclk));
	jdff dff_B_mxDxIay68_0(.din(w_dff_B_ypOF11ny7_0),.dout(w_dff_B_mxDxIay68_0),.clk(gclk));
	jdff dff_B_OOC2jVv87_0(.din(w_dff_B_mxDxIay68_0),.dout(w_dff_B_OOC2jVv87_0),.clk(gclk));
	jdff dff_B_Cy9UViWe1_0(.din(w_dff_B_OOC2jVv87_0),.dout(w_dff_B_Cy9UViWe1_0),.clk(gclk));
	jdff dff_B_MrbGNQYL7_0(.din(w_dff_B_Cy9UViWe1_0),.dout(w_dff_B_MrbGNQYL7_0),.clk(gclk));
	jdff dff_B_BWYUbXs32_0(.din(w_dff_B_MrbGNQYL7_0),.dout(w_dff_B_BWYUbXs32_0),.clk(gclk));
	jdff dff_B_cGcQ3dir2_0(.din(w_dff_B_BWYUbXs32_0),.dout(w_dff_B_cGcQ3dir2_0),.clk(gclk));
	jdff dff_B_IjwtMq1Q2_0(.din(w_dff_B_cGcQ3dir2_0),.dout(w_dff_B_IjwtMq1Q2_0),.clk(gclk));
	jdff dff_B_YrkQIZLi8_0(.din(w_dff_B_IjwtMq1Q2_0),.dout(w_dff_B_YrkQIZLi8_0),.clk(gclk));
	jdff dff_B_83JO0qDw7_0(.din(w_dff_B_YrkQIZLi8_0),.dout(w_dff_B_83JO0qDw7_0),.clk(gclk));
	jdff dff_B_u4zdLjIr7_0(.din(w_dff_B_83JO0qDw7_0),.dout(w_dff_B_u4zdLjIr7_0),.clk(gclk));
	jdff dff_B_OvoTV3iT5_0(.din(w_dff_B_u4zdLjIr7_0),.dout(w_dff_B_OvoTV3iT5_0),.clk(gclk));
	jdff dff_B_AKxmYToU0_0(.din(w_dff_B_OvoTV3iT5_0),.dout(w_dff_B_AKxmYToU0_0),.clk(gclk));
	jdff dff_B_rB8X50qJ6_0(.din(w_dff_B_AKxmYToU0_0),.dout(w_dff_B_rB8X50qJ6_0),.clk(gclk));
	jdff dff_B_Xxzgxo4c9_0(.din(w_dff_B_rB8X50qJ6_0),.dout(w_dff_B_Xxzgxo4c9_0),.clk(gclk));
	jdff dff_B_SxquOrW65_0(.din(w_dff_B_Xxzgxo4c9_0),.dout(w_dff_B_SxquOrW65_0),.clk(gclk));
	jdff dff_B_KZGxgImK6_0(.din(w_dff_B_SxquOrW65_0),.dout(w_dff_B_KZGxgImK6_0),.clk(gclk));
	jdff dff_B_PJp2lxaC5_0(.din(w_dff_B_KZGxgImK6_0),.dout(w_dff_B_PJp2lxaC5_0),.clk(gclk));
	jdff dff_B_ChAtkDs68_0(.din(w_dff_B_PJp2lxaC5_0),.dout(w_dff_B_ChAtkDs68_0),.clk(gclk));
	jdff dff_B_nZxjo0XW2_0(.din(w_dff_B_ChAtkDs68_0),.dout(w_dff_B_nZxjo0XW2_0),.clk(gclk));
	jdff dff_B_5nBc7xwK0_0(.din(w_dff_B_nZxjo0XW2_0),.dout(w_dff_B_5nBc7xwK0_0),.clk(gclk));
	jdff dff_B_Xv7jY3EZ5_0(.din(w_dff_B_5nBc7xwK0_0),.dout(w_dff_B_Xv7jY3EZ5_0),.clk(gclk));
	jdff dff_B_THzs32C03_0(.din(w_dff_B_Xv7jY3EZ5_0),.dout(w_dff_B_THzs32C03_0),.clk(gclk));
	jdff dff_B_I7MFPJDM5_0(.din(w_dff_B_THzs32C03_0),.dout(w_dff_B_I7MFPJDM5_0),.clk(gclk));
	jdff dff_B_2Cn5U2F45_0(.din(w_dff_B_I7MFPJDM5_0),.dout(w_dff_B_2Cn5U2F45_0),.clk(gclk));
	jdff dff_B_lLJQocVo0_0(.din(w_dff_B_2Cn5U2F45_0),.dout(w_dff_B_lLJQocVo0_0),.clk(gclk));
	jdff dff_B_H3HluzHI1_0(.din(w_dff_B_lLJQocVo0_0),.dout(w_dff_B_H3HluzHI1_0),.clk(gclk));
	jdff dff_B_Oe8ll1Ws8_0(.din(w_dff_B_H3HluzHI1_0),.dout(w_dff_B_Oe8ll1Ws8_0),.clk(gclk));
	jdff dff_B_FnJBjWar1_0(.din(w_dff_B_Oe8ll1Ws8_0),.dout(w_dff_B_FnJBjWar1_0),.clk(gclk));
	jdff dff_B_G0qZVe1L0_0(.din(w_dff_B_FnJBjWar1_0),.dout(w_dff_B_G0qZVe1L0_0),.clk(gclk));
	jdff dff_B_bZvfMu5U8_0(.din(w_dff_B_G0qZVe1L0_0),.dout(w_dff_B_bZvfMu5U8_0),.clk(gclk));
	jdff dff_B_VFHLz0Y14_0(.din(w_dff_B_bZvfMu5U8_0),.dout(w_dff_B_VFHLz0Y14_0),.clk(gclk));
	jdff dff_B_cMimULRD4_0(.din(w_dff_B_VFHLz0Y14_0),.dout(w_dff_B_cMimULRD4_0),.clk(gclk));
	jdff dff_B_jtKpkOcZ6_0(.din(w_dff_B_cMimULRD4_0),.dout(w_dff_B_jtKpkOcZ6_0),.clk(gclk));
	jdff dff_B_IztNoIMf2_0(.din(w_dff_B_jtKpkOcZ6_0),.dout(w_dff_B_IztNoIMf2_0),.clk(gclk));
	jdff dff_B_K3mqoUfs1_0(.din(w_dff_B_IztNoIMf2_0),.dout(w_dff_B_K3mqoUfs1_0),.clk(gclk));
	jdff dff_B_fsw5iKBs5_0(.din(w_dff_B_K3mqoUfs1_0),.dout(w_dff_B_fsw5iKBs5_0),.clk(gclk));
	jdff dff_B_MZQyXlyG3_0(.din(w_dff_B_fsw5iKBs5_0),.dout(w_dff_B_MZQyXlyG3_0),.clk(gclk));
	jdff dff_B_NlwdAv251_0(.din(w_dff_B_MZQyXlyG3_0),.dout(w_dff_B_NlwdAv251_0),.clk(gclk));
	jdff dff_B_4qZsYSHs0_0(.din(w_dff_B_NlwdAv251_0),.dout(w_dff_B_4qZsYSHs0_0),.clk(gclk));
	jdff dff_B_lhi9bC4H7_0(.din(w_dff_B_4qZsYSHs0_0),.dout(w_dff_B_lhi9bC4H7_0),.clk(gclk));
	jdff dff_B_VD3Wc7S56_0(.din(w_dff_B_lhi9bC4H7_0),.dout(w_dff_B_VD3Wc7S56_0),.clk(gclk));
	jdff dff_B_JVLbNvhS5_0(.din(w_dff_B_VD3Wc7S56_0),.dout(w_dff_B_JVLbNvhS5_0),.clk(gclk));
	jdff dff_B_I1RSLtRl2_0(.din(w_dff_B_JVLbNvhS5_0),.dout(w_dff_B_I1RSLtRl2_0),.clk(gclk));
	jdff dff_B_jiebWjNd1_0(.din(w_dff_B_I1RSLtRl2_0),.dout(w_dff_B_jiebWjNd1_0),.clk(gclk));
	jdff dff_B_ZjkdADfx0_0(.din(w_dff_B_jiebWjNd1_0),.dout(w_dff_B_ZjkdADfx0_0),.clk(gclk));
	jdff dff_B_FfLSB3rV3_0(.din(w_dff_B_ZjkdADfx0_0),.dout(w_dff_B_FfLSB3rV3_0),.clk(gclk));
	jdff dff_B_JUguTPI86_0(.din(w_dff_B_FfLSB3rV3_0),.dout(w_dff_B_JUguTPI86_0),.clk(gclk));
	jdff dff_B_PcIGDrxO4_0(.din(w_dff_B_JUguTPI86_0),.dout(w_dff_B_PcIGDrxO4_0),.clk(gclk));
	jdff dff_B_BDNe8ZEZ7_0(.din(w_dff_B_PcIGDrxO4_0),.dout(w_dff_B_BDNe8ZEZ7_0),.clk(gclk));
	jdff dff_B_KH5FZZGx9_0(.din(w_dff_B_BDNe8ZEZ7_0),.dout(w_dff_B_KH5FZZGx9_0),.clk(gclk));
	jdff dff_B_5DURdh370_0(.din(w_dff_B_KH5FZZGx9_0),.dout(w_dff_B_5DURdh370_0),.clk(gclk));
	jdff dff_B_q4K6CRfJ5_0(.din(w_dff_B_5DURdh370_0),.dout(w_dff_B_q4K6CRfJ5_0),.clk(gclk));
	jdff dff_B_vXlbygkA6_0(.din(w_dff_B_q4K6CRfJ5_0),.dout(w_dff_B_vXlbygkA6_0),.clk(gclk));
	jdff dff_B_VGTIDXsV5_0(.din(w_dff_B_vXlbygkA6_0),.dout(w_dff_B_VGTIDXsV5_0),.clk(gclk));
	jdff dff_B_XXOZJK8q0_0(.din(w_dff_B_VGTIDXsV5_0),.dout(w_dff_B_XXOZJK8q0_0),.clk(gclk));
	jdff dff_B_aaQvUOy22_0(.din(w_dff_B_XXOZJK8q0_0),.dout(w_dff_B_aaQvUOy22_0),.clk(gclk));
	jdff dff_B_WpE5i4M96_0(.din(w_dff_B_aaQvUOy22_0),.dout(w_dff_B_WpE5i4M96_0),.clk(gclk));
	jdff dff_B_8qzNuaiB0_0(.din(w_dff_B_WpE5i4M96_0),.dout(w_dff_B_8qzNuaiB0_0),.clk(gclk));
	jdff dff_B_zJ6k3pij6_0(.din(w_dff_B_8qzNuaiB0_0),.dout(w_dff_B_zJ6k3pij6_0),.clk(gclk));
	jdff dff_B_tNMA2gKW9_0(.din(w_dff_B_zJ6k3pij6_0),.dout(w_dff_B_tNMA2gKW9_0),.clk(gclk));
	jdff dff_B_UcgRjmm15_0(.din(w_dff_B_tNMA2gKW9_0),.dout(w_dff_B_UcgRjmm15_0),.clk(gclk));
	jdff dff_B_FdCSyEd02_0(.din(w_dff_B_UcgRjmm15_0),.dout(w_dff_B_FdCSyEd02_0),.clk(gclk));
	jdff dff_B_AXYDZMNB2_0(.din(w_dff_B_FdCSyEd02_0),.dout(w_dff_B_AXYDZMNB2_0),.clk(gclk));
	jdff dff_B_z1wmerGy6_0(.din(w_dff_B_AXYDZMNB2_0),.dout(w_dff_B_z1wmerGy6_0),.clk(gclk));
	jdff dff_B_MdDCbMdU2_0(.din(w_dff_B_z1wmerGy6_0),.dout(w_dff_B_MdDCbMdU2_0),.clk(gclk));
	jdff dff_B_qpSaXMca4_0(.din(w_dff_B_MdDCbMdU2_0),.dout(w_dff_B_qpSaXMca4_0),.clk(gclk));
	jdff dff_B_FIpSm2XP9_0(.din(w_dff_B_qpSaXMca4_0),.dout(w_dff_B_FIpSm2XP9_0),.clk(gclk));
	jdff dff_B_BAYi9v7u5_0(.din(w_dff_B_FIpSm2XP9_0),.dout(w_dff_B_BAYi9v7u5_0),.clk(gclk));
	jdff dff_B_Uz99iBGr7_0(.din(w_dff_B_BAYi9v7u5_0),.dout(w_dff_B_Uz99iBGr7_0),.clk(gclk));
	jdff dff_B_SaRDTlUT9_0(.din(w_dff_B_Uz99iBGr7_0),.dout(w_dff_B_SaRDTlUT9_0),.clk(gclk));
	jdff dff_B_aKphVdIy6_0(.din(w_dff_B_SaRDTlUT9_0),.dout(w_dff_B_aKphVdIy6_0),.clk(gclk));
	jdff dff_B_VGjpTU1u9_0(.din(w_dff_B_aKphVdIy6_0),.dout(w_dff_B_VGjpTU1u9_0),.clk(gclk));
	jdff dff_B_E2S8nRC23_0(.din(w_dff_B_VGjpTU1u9_0),.dout(w_dff_B_E2S8nRC23_0),.clk(gclk));
	jdff dff_B_x0fgemQS2_0(.din(w_dff_B_E2S8nRC23_0),.dout(w_dff_B_x0fgemQS2_0),.clk(gclk));
	jdff dff_B_fi93cS7e7_0(.din(w_dff_B_x0fgemQS2_0),.dout(w_dff_B_fi93cS7e7_0),.clk(gclk));
	jdff dff_B_X6rYgYGA1_0(.din(w_dff_B_fi93cS7e7_0),.dout(w_dff_B_X6rYgYGA1_0),.clk(gclk));
	jdff dff_B_LFeU1zzp4_0(.din(w_dff_B_X6rYgYGA1_0),.dout(w_dff_B_LFeU1zzp4_0),.clk(gclk));
	jdff dff_B_diSNUr6c2_0(.din(w_dff_B_LFeU1zzp4_0),.dout(w_dff_B_diSNUr6c2_0),.clk(gclk));
	jdff dff_B_k0Svme9a1_0(.din(w_dff_B_diSNUr6c2_0),.dout(w_dff_B_k0Svme9a1_0),.clk(gclk));
	jdff dff_B_Gzgy1Qhg2_0(.din(w_dff_B_k0Svme9a1_0),.dout(w_dff_B_Gzgy1Qhg2_0),.clk(gclk));
	jdff dff_B_G7Zm8O1g3_0(.din(w_dff_B_Gzgy1Qhg2_0),.dout(w_dff_B_G7Zm8O1g3_0),.clk(gclk));
	jdff dff_B_iFZ3HDaO6_0(.din(w_dff_B_G7Zm8O1g3_0),.dout(w_dff_B_iFZ3HDaO6_0),.clk(gclk));
	jdff dff_B_pkVu7UHh8_0(.din(w_dff_B_iFZ3HDaO6_0),.dout(w_dff_B_pkVu7UHh8_0),.clk(gclk));
	jdff dff_B_gJWoYztq2_0(.din(w_dff_B_pkVu7UHh8_0),.dout(w_dff_B_gJWoYztq2_0),.clk(gclk));
	jdff dff_B_QphMgtJX7_0(.din(w_dff_B_gJWoYztq2_0),.dout(w_dff_B_QphMgtJX7_0),.clk(gclk));
	jdff dff_B_MNe3cJhP9_0(.din(w_dff_B_QphMgtJX7_0),.dout(w_dff_B_MNe3cJhP9_0),.clk(gclk));
	jdff dff_B_Kj5AR5fJ7_1(.din(n990),.dout(w_dff_B_Kj5AR5fJ7_1),.clk(gclk));
	jdff dff_B_oovlYFa64_1(.din(w_dff_B_Kj5AR5fJ7_1),.dout(w_dff_B_oovlYFa64_1),.clk(gclk));
	jdff dff_B_Oq3sHPJg2_1(.din(w_dff_B_oovlYFa64_1),.dout(w_dff_B_Oq3sHPJg2_1),.clk(gclk));
	jdff dff_B_xjPrILrz4_1(.din(w_dff_B_Oq3sHPJg2_1),.dout(w_dff_B_xjPrILrz4_1),.clk(gclk));
	jdff dff_B_F4lLoHk67_1(.din(w_dff_B_xjPrILrz4_1),.dout(w_dff_B_F4lLoHk67_1),.clk(gclk));
	jdff dff_B_7PrOpdYl8_1(.din(w_dff_B_F4lLoHk67_1),.dout(w_dff_B_7PrOpdYl8_1),.clk(gclk));
	jdff dff_B_wHjuVeUC1_1(.din(w_dff_B_7PrOpdYl8_1),.dout(w_dff_B_wHjuVeUC1_1),.clk(gclk));
	jdff dff_B_bRPaR6oL3_1(.din(w_dff_B_wHjuVeUC1_1),.dout(w_dff_B_bRPaR6oL3_1),.clk(gclk));
	jdff dff_B_CdFqOPkU0_1(.din(w_dff_B_bRPaR6oL3_1),.dout(w_dff_B_CdFqOPkU0_1),.clk(gclk));
	jdff dff_B_Q6drcGUE6_1(.din(w_dff_B_CdFqOPkU0_1),.dout(w_dff_B_Q6drcGUE6_1),.clk(gclk));
	jdff dff_B_JWBxPnSI7_1(.din(w_dff_B_Q6drcGUE6_1),.dout(w_dff_B_JWBxPnSI7_1),.clk(gclk));
	jdff dff_B_s9wLR4hg0_1(.din(w_dff_B_JWBxPnSI7_1),.dout(w_dff_B_s9wLR4hg0_1),.clk(gclk));
	jdff dff_B_CTnX0Qhc5_1(.din(w_dff_B_s9wLR4hg0_1),.dout(w_dff_B_CTnX0Qhc5_1),.clk(gclk));
	jdff dff_B_8iFRSUQ14_1(.din(w_dff_B_CTnX0Qhc5_1),.dout(w_dff_B_8iFRSUQ14_1),.clk(gclk));
	jdff dff_B_0gBtGdap6_1(.din(w_dff_B_8iFRSUQ14_1),.dout(w_dff_B_0gBtGdap6_1),.clk(gclk));
	jdff dff_B_15GUVvqO8_1(.din(w_dff_B_0gBtGdap6_1),.dout(w_dff_B_15GUVvqO8_1),.clk(gclk));
	jdff dff_B_zPMx39Ge7_1(.din(w_dff_B_15GUVvqO8_1),.dout(w_dff_B_zPMx39Ge7_1),.clk(gclk));
	jdff dff_B_yC50Oo7z4_1(.din(w_dff_B_zPMx39Ge7_1),.dout(w_dff_B_yC50Oo7z4_1),.clk(gclk));
	jdff dff_B_i2gZfiC96_1(.din(w_dff_B_yC50Oo7z4_1),.dout(w_dff_B_i2gZfiC96_1),.clk(gclk));
	jdff dff_B_W1GlwIdV2_1(.din(w_dff_B_i2gZfiC96_1),.dout(w_dff_B_W1GlwIdV2_1),.clk(gclk));
	jdff dff_B_GqDpNLGt6_1(.din(w_dff_B_W1GlwIdV2_1),.dout(w_dff_B_GqDpNLGt6_1),.clk(gclk));
	jdff dff_B_6jh7DCiL5_1(.din(w_dff_B_GqDpNLGt6_1),.dout(w_dff_B_6jh7DCiL5_1),.clk(gclk));
	jdff dff_B_oX0dvEqh0_1(.din(w_dff_B_6jh7DCiL5_1),.dout(w_dff_B_oX0dvEqh0_1),.clk(gclk));
	jdff dff_B_Ox9u8pFD1_1(.din(w_dff_B_oX0dvEqh0_1),.dout(w_dff_B_Ox9u8pFD1_1),.clk(gclk));
	jdff dff_B_0XUaaG3w6_1(.din(w_dff_B_Ox9u8pFD1_1),.dout(w_dff_B_0XUaaG3w6_1),.clk(gclk));
	jdff dff_B_QbeXYslI5_1(.din(w_dff_B_0XUaaG3w6_1),.dout(w_dff_B_QbeXYslI5_1),.clk(gclk));
	jdff dff_B_hdejZx0q3_1(.din(w_dff_B_QbeXYslI5_1),.dout(w_dff_B_hdejZx0q3_1),.clk(gclk));
	jdff dff_B_NsNeJRRP7_1(.din(w_dff_B_hdejZx0q3_1),.dout(w_dff_B_NsNeJRRP7_1),.clk(gclk));
	jdff dff_B_rCFS9CA73_1(.din(w_dff_B_NsNeJRRP7_1),.dout(w_dff_B_rCFS9CA73_1),.clk(gclk));
	jdff dff_B_UG2dEszc7_1(.din(w_dff_B_rCFS9CA73_1),.dout(w_dff_B_UG2dEszc7_1),.clk(gclk));
	jdff dff_B_4ekLntUr4_1(.din(w_dff_B_UG2dEszc7_1),.dout(w_dff_B_4ekLntUr4_1),.clk(gclk));
	jdff dff_B_KSbivQYk5_1(.din(w_dff_B_4ekLntUr4_1),.dout(w_dff_B_KSbivQYk5_1),.clk(gclk));
	jdff dff_B_jwm2cIUf8_1(.din(w_dff_B_KSbivQYk5_1),.dout(w_dff_B_jwm2cIUf8_1),.clk(gclk));
	jdff dff_B_wDMddMnV5_1(.din(w_dff_B_jwm2cIUf8_1),.dout(w_dff_B_wDMddMnV5_1),.clk(gclk));
	jdff dff_B_cTG46KWu8_1(.din(w_dff_B_wDMddMnV5_1),.dout(w_dff_B_cTG46KWu8_1),.clk(gclk));
	jdff dff_B_2B57DeYB5_1(.din(w_dff_B_cTG46KWu8_1),.dout(w_dff_B_2B57DeYB5_1),.clk(gclk));
	jdff dff_B_LpvxXFYX9_1(.din(w_dff_B_2B57DeYB5_1),.dout(w_dff_B_LpvxXFYX9_1),.clk(gclk));
	jdff dff_B_w4YPEJlc9_1(.din(w_dff_B_LpvxXFYX9_1),.dout(w_dff_B_w4YPEJlc9_1),.clk(gclk));
	jdff dff_B_gKUC1bO50_1(.din(w_dff_B_w4YPEJlc9_1),.dout(w_dff_B_gKUC1bO50_1),.clk(gclk));
	jdff dff_B_7nXJ67Dt8_1(.din(w_dff_B_gKUC1bO50_1),.dout(w_dff_B_7nXJ67Dt8_1),.clk(gclk));
	jdff dff_B_lfdK1lJW1_1(.din(w_dff_B_7nXJ67Dt8_1),.dout(w_dff_B_lfdK1lJW1_1),.clk(gclk));
	jdff dff_B_7L3Oi4Vy0_1(.din(w_dff_B_lfdK1lJW1_1),.dout(w_dff_B_7L3Oi4Vy0_1),.clk(gclk));
	jdff dff_B_PBi1OoMT8_1(.din(w_dff_B_7L3Oi4Vy0_1),.dout(w_dff_B_PBi1OoMT8_1),.clk(gclk));
	jdff dff_B_9auMD5uR7_1(.din(w_dff_B_PBi1OoMT8_1),.dout(w_dff_B_9auMD5uR7_1),.clk(gclk));
	jdff dff_B_eqS0iseN6_1(.din(w_dff_B_9auMD5uR7_1),.dout(w_dff_B_eqS0iseN6_1),.clk(gclk));
	jdff dff_B_Cet8uBUu6_1(.din(w_dff_B_eqS0iseN6_1),.dout(w_dff_B_Cet8uBUu6_1),.clk(gclk));
	jdff dff_B_k0F8m3NB9_1(.din(w_dff_B_Cet8uBUu6_1),.dout(w_dff_B_k0F8m3NB9_1),.clk(gclk));
	jdff dff_B_SZQUkxMM3_1(.din(w_dff_B_k0F8m3NB9_1),.dout(w_dff_B_SZQUkxMM3_1),.clk(gclk));
	jdff dff_B_v36G6yS04_1(.din(w_dff_B_SZQUkxMM3_1),.dout(w_dff_B_v36G6yS04_1),.clk(gclk));
	jdff dff_B_BkwC78Od6_1(.din(w_dff_B_v36G6yS04_1),.dout(w_dff_B_BkwC78Od6_1),.clk(gclk));
	jdff dff_B_uwb9k4xF1_1(.din(w_dff_B_BkwC78Od6_1),.dout(w_dff_B_uwb9k4xF1_1),.clk(gclk));
	jdff dff_B_nmsBbPLB4_1(.din(w_dff_B_uwb9k4xF1_1),.dout(w_dff_B_nmsBbPLB4_1),.clk(gclk));
	jdff dff_B_K8EOOJ1M7_1(.din(w_dff_B_nmsBbPLB4_1),.dout(w_dff_B_K8EOOJ1M7_1),.clk(gclk));
	jdff dff_B_5mIDOJEl0_1(.din(w_dff_B_K8EOOJ1M7_1),.dout(w_dff_B_5mIDOJEl0_1),.clk(gclk));
	jdff dff_B_ynEJA2Cc8_1(.din(w_dff_B_5mIDOJEl0_1),.dout(w_dff_B_ynEJA2Cc8_1),.clk(gclk));
	jdff dff_B_fERPU5X67_1(.din(w_dff_B_ynEJA2Cc8_1),.dout(w_dff_B_fERPU5X67_1),.clk(gclk));
	jdff dff_B_25EwPB4s3_1(.din(w_dff_B_fERPU5X67_1),.dout(w_dff_B_25EwPB4s3_1),.clk(gclk));
	jdff dff_B_9AC2eQed8_1(.din(w_dff_B_25EwPB4s3_1),.dout(w_dff_B_9AC2eQed8_1),.clk(gclk));
	jdff dff_B_wMCjXOI78_1(.din(w_dff_B_9AC2eQed8_1),.dout(w_dff_B_wMCjXOI78_1),.clk(gclk));
	jdff dff_B_M7JlE5Aj8_1(.din(w_dff_B_wMCjXOI78_1),.dout(w_dff_B_M7JlE5Aj8_1),.clk(gclk));
	jdff dff_B_vms5oa6r8_1(.din(w_dff_B_M7JlE5Aj8_1),.dout(w_dff_B_vms5oa6r8_1),.clk(gclk));
	jdff dff_B_xNZqeWOU9_1(.din(w_dff_B_vms5oa6r8_1),.dout(w_dff_B_xNZqeWOU9_1),.clk(gclk));
	jdff dff_B_TBbIDfG28_1(.din(w_dff_B_xNZqeWOU9_1),.dout(w_dff_B_TBbIDfG28_1),.clk(gclk));
	jdff dff_B_nSaVU8LB8_1(.din(w_dff_B_TBbIDfG28_1),.dout(w_dff_B_nSaVU8LB8_1),.clk(gclk));
	jdff dff_B_Li1VsOmH7_1(.din(w_dff_B_nSaVU8LB8_1),.dout(w_dff_B_Li1VsOmH7_1),.clk(gclk));
	jdff dff_B_zfahlay29_1(.din(w_dff_B_Li1VsOmH7_1),.dout(w_dff_B_zfahlay29_1),.clk(gclk));
	jdff dff_B_dUFONw517_1(.din(w_dff_B_zfahlay29_1),.dout(w_dff_B_dUFONw517_1),.clk(gclk));
	jdff dff_B_xF30TW5R7_1(.din(w_dff_B_dUFONw517_1),.dout(w_dff_B_xF30TW5R7_1),.clk(gclk));
	jdff dff_B_XTErd2bd2_1(.din(w_dff_B_xF30TW5R7_1),.dout(w_dff_B_XTErd2bd2_1),.clk(gclk));
	jdff dff_B_SKDCRRov5_1(.din(w_dff_B_XTErd2bd2_1),.dout(w_dff_B_SKDCRRov5_1),.clk(gclk));
	jdff dff_B_EufDlfqr8_1(.din(w_dff_B_SKDCRRov5_1),.dout(w_dff_B_EufDlfqr8_1),.clk(gclk));
	jdff dff_B_yc8vxl173_1(.din(w_dff_B_EufDlfqr8_1),.dout(w_dff_B_yc8vxl173_1),.clk(gclk));
	jdff dff_B_S2LNM6L52_1(.din(w_dff_B_yc8vxl173_1),.dout(w_dff_B_S2LNM6L52_1),.clk(gclk));
	jdff dff_B_TXNrvu3H2_1(.din(w_dff_B_S2LNM6L52_1),.dout(w_dff_B_TXNrvu3H2_1),.clk(gclk));
	jdff dff_B_wVkADsaW7_1(.din(w_dff_B_TXNrvu3H2_1),.dout(w_dff_B_wVkADsaW7_1),.clk(gclk));
	jdff dff_B_7pjHbMAI4_1(.din(w_dff_B_wVkADsaW7_1),.dout(w_dff_B_7pjHbMAI4_1),.clk(gclk));
	jdff dff_B_CZyv6MJn5_1(.din(w_dff_B_7pjHbMAI4_1),.dout(w_dff_B_CZyv6MJn5_1),.clk(gclk));
	jdff dff_B_RjzaxENB5_1(.din(w_dff_B_CZyv6MJn5_1),.dout(w_dff_B_RjzaxENB5_1),.clk(gclk));
	jdff dff_B_ws037e9S8_1(.din(w_dff_B_RjzaxENB5_1),.dout(w_dff_B_ws037e9S8_1),.clk(gclk));
	jdff dff_B_1RiDqpM92_1(.din(w_dff_B_ws037e9S8_1),.dout(w_dff_B_1RiDqpM92_1),.clk(gclk));
	jdff dff_B_7iulf4eM9_1(.din(w_dff_B_1RiDqpM92_1),.dout(w_dff_B_7iulf4eM9_1),.clk(gclk));
	jdff dff_B_AmMmxHSs5_1(.din(w_dff_B_7iulf4eM9_1),.dout(w_dff_B_AmMmxHSs5_1),.clk(gclk));
	jdff dff_B_L4mSRr4i5_1(.din(w_dff_B_AmMmxHSs5_1),.dout(w_dff_B_L4mSRr4i5_1),.clk(gclk));
	jdff dff_B_GDBqg1AN6_1(.din(w_dff_B_L4mSRr4i5_1),.dout(w_dff_B_GDBqg1AN6_1),.clk(gclk));
	jdff dff_B_R12BfaXI8_1(.din(w_dff_B_GDBqg1AN6_1),.dout(w_dff_B_R12BfaXI8_1),.clk(gclk));
	jdff dff_B_IuPAEgwk6_1(.din(w_dff_B_R12BfaXI8_1),.dout(w_dff_B_IuPAEgwk6_1),.clk(gclk));
	jdff dff_B_fcZduaqd0_1(.din(w_dff_B_IuPAEgwk6_1),.dout(w_dff_B_fcZduaqd0_1),.clk(gclk));
	jdff dff_B_VoNjxuvq5_1(.din(w_dff_B_fcZduaqd0_1),.dout(w_dff_B_VoNjxuvq5_1),.clk(gclk));
	jdff dff_B_wktnuJFL4_1(.din(w_dff_B_VoNjxuvq5_1),.dout(w_dff_B_wktnuJFL4_1),.clk(gclk));
	jdff dff_B_12byotXl6_1(.din(w_dff_B_wktnuJFL4_1),.dout(w_dff_B_12byotXl6_1),.clk(gclk));
	jdff dff_B_aaVNcO7N2_1(.din(w_dff_B_12byotXl6_1),.dout(w_dff_B_aaVNcO7N2_1),.clk(gclk));
	jdff dff_B_aZasClLY4_1(.din(w_dff_B_aaVNcO7N2_1),.dout(w_dff_B_aZasClLY4_1),.clk(gclk));
	jdff dff_B_qn2brB9g5_1(.din(w_dff_B_aZasClLY4_1),.dout(w_dff_B_qn2brB9g5_1),.clk(gclk));
	jdff dff_B_SiLJdpvG4_1(.din(w_dff_B_qn2brB9g5_1),.dout(w_dff_B_SiLJdpvG4_1),.clk(gclk));
	jdff dff_B_4VtBdByz4_1(.din(w_dff_B_SiLJdpvG4_1),.dout(w_dff_B_4VtBdByz4_1),.clk(gclk));
	jdff dff_B_hUe7bFZi0_1(.din(w_dff_B_4VtBdByz4_1),.dout(w_dff_B_hUe7bFZi0_1),.clk(gclk));
	jdff dff_B_Iw8yfBaD8_1(.din(w_dff_B_hUe7bFZi0_1),.dout(w_dff_B_Iw8yfBaD8_1),.clk(gclk));
	jdff dff_B_D9pND7lJ6_1(.din(w_dff_B_Iw8yfBaD8_1),.dout(w_dff_B_D9pND7lJ6_1),.clk(gclk));
	jdff dff_B_RfhM5a1Q5_1(.din(w_dff_B_D9pND7lJ6_1),.dout(w_dff_B_RfhM5a1Q5_1),.clk(gclk));
	jdff dff_B_b3qpPrCX5_1(.din(w_dff_B_RfhM5a1Q5_1),.dout(w_dff_B_b3qpPrCX5_1),.clk(gclk));
	jdff dff_B_eOrMuw528_1(.din(w_dff_B_b3qpPrCX5_1),.dout(w_dff_B_eOrMuw528_1),.clk(gclk));
	jdff dff_B_PQRirv0m1_0(.din(n991),.dout(w_dff_B_PQRirv0m1_0),.clk(gclk));
	jdff dff_B_D9gpv3kI4_0(.din(w_dff_B_PQRirv0m1_0),.dout(w_dff_B_D9gpv3kI4_0),.clk(gclk));
	jdff dff_B_4K39FXIG9_0(.din(w_dff_B_D9gpv3kI4_0),.dout(w_dff_B_4K39FXIG9_0),.clk(gclk));
	jdff dff_B_8PdTeILF8_0(.din(w_dff_B_4K39FXIG9_0),.dout(w_dff_B_8PdTeILF8_0),.clk(gclk));
	jdff dff_B_2T2924mg3_0(.din(w_dff_B_8PdTeILF8_0),.dout(w_dff_B_2T2924mg3_0),.clk(gclk));
	jdff dff_B_v4SQFyul6_0(.din(w_dff_B_2T2924mg3_0),.dout(w_dff_B_v4SQFyul6_0),.clk(gclk));
	jdff dff_B_ri0HYp239_0(.din(w_dff_B_v4SQFyul6_0),.dout(w_dff_B_ri0HYp239_0),.clk(gclk));
	jdff dff_B_1ypkeiBu2_0(.din(w_dff_B_ri0HYp239_0),.dout(w_dff_B_1ypkeiBu2_0),.clk(gclk));
	jdff dff_B_y9nRsGxj9_0(.din(w_dff_B_1ypkeiBu2_0),.dout(w_dff_B_y9nRsGxj9_0),.clk(gclk));
	jdff dff_B_TTfgeIOM0_0(.din(w_dff_B_y9nRsGxj9_0),.dout(w_dff_B_TTfgeIOM0_0),.clk(gclk));
	jdff dff_B_aHfEl3WP9_0(.din(w_dff_B_TTfgeIOM0_0),.dout(w_dff_B_aHfEl3WP9_0),.clk(gclk));
	jdff dff_B_BYKjJXzo3_0(.din(w_dff_B_aHfEl3WP9_0),.dout(w_dff_B_BYKjJXzo3_0),.clk(gclk));
	jdff dff_B_gCklSXy41_0(.din(w_dff_B_BYKjJXzo3_0),.dout(w_dff_B_gCklSXy41_0),.clk(gclk));
	jdff dff_B_7IFKvv5m7_0(.din(w_dff_B_gCklSXy41_0),.dout(w_dff_B_7IFKvv5m7_0),.clk(gclk));
	jdff dff_B_i8Xq67pF2_0(.din(w_dff_B_7IFKvv5m7_0),.dout(w_dff_B_i8Xq67pF2_0),.clk(gclk));
	jdff dff_B_FfZUezRD1_0(.din(w_dff_B_i8Xq67pF2_0),.dout(w_dff_B_FfZUezRD1_0),.clk(gclk));
	jdff dff_B_ecgCzsY40_0(.din(w_dff_B_FfZUezRD1_0),.dout(w_dff_B_ecgCzsY40_0),.clk(gclk));
	jdff dff_B_rTBFtG2P6_0(.din(w_dff_B_ecgCzsY40_0),.dout(w_dff_B_rTBFtG2P6_0),.clk(gclk));
	jdff dff_B_XDrDrEvz3_0(.din(w_dff_B_rTBFtG2P6_0),.dout(w_dff_B_XDrDrEvz3_0),.clk(gclk));
	jdff dff_B_ewOkrIJn8_0(.din(w_dff_B_XDrDrEvz3_0),.dout(w_dff_B_ewOkrIJn8_0),.clk(gclk));
	jdff dff_B_nn3scauF5_0(.din(w_dff_B_ewOkrIJn8_0),.dout(w_dff_B_nn3scauF5_0),.clk(gclk));
	jdff dff_B_dcrNNsXE3_0(.din(w_dff_B_nn3scauF5_0),.dout(w_dff_B_dcrNNsXE3_0),.clk(gclk));
	jdff dff_B_xVkHm4c43_0(.din(w_dff_B_dcrNNsXE3_0),.dout(w_dff_B_xVkHm4c43_0),.clk(gclk));
	jdff dff_B_m4vONICa3_0(.din(w_dff_B_xVkHm4c43_0),.dout(w_dff_B_m4vONICa3_0),.clk(gclk));
	jdff dff_B_lnc1Snmr9_0(.din(w_dff_B_m4vONICa3_0),.dout(w_dff_B_lnc1Snmr9_0),.clk(gclk));
	jdff dff_B_cw030unO2_0(.din(w_dff_B_lnc1Snmr9_0),.dout(w_dff_B_cw030unO2_0),.clk(gclk));
	jdff dff_B_TEO5YD8Z8_0(.din(w_dff_B_cw030unO2_0),.dout(w_dff_B_TEO5YD8Z8_0),.clk(gclk));
	jdff dff_B_LQrZYVFJ6_0(.din(w_dff_B_TEO5YD8Z8_0),.dout(w_dff_B_LQrZYVFJ6_0),.clk(gclk));
	jdff dff_B_DYhN7bMT4_0(.din(w_dff_B_LQrZYVFJ6_0),.dout(w_dff_B_DYhN7bMT4_0),.clk(gclk));
	jdff dff_B_DoVj4msS1_0(.din(w_dff_B_DYhN7bMT4_0),.dout(w_dff_B_DoVj4msS1_0),.clk(gclk));
	jdff dff_B_AN4TmMtZ1_0(.din(w_dff_B_DoVj4msS1_0),.dout(w_dff_B_AN4TmMtZ1_0),.clk(gclk));
	jdff dff_B_r1HvdoVy1_0(.din(w_dff_B_AN4TmMtZ1_0),.dout(w_dff_B_r1HvdoVy1_0),.clk(gclk));
	jdff dff_B_v8ivtiXS6_0(.din(w_dff_B_r1HvdoVy1_0),.dout(w_dff_B_v8ivtiXS6_0),.clk(gclk));
	jdff dff_B_Ng9qgkXr5_0(.din(w_dff_B_v8ivtiXS6_0),.dout(w_dff_B_Ng9qgkXr5_0),.clk(gclk));
	jdff dff_B_mCWpCiQC9_0(.din(w_dff_B_Ng9qgkXr5_0),.dout(w_dff_B_mCWpCiQC9_0),.clk(gclk));
	jdff dff_B_TVLkAODu4_0(.din(w_dff_B_mCWpCiQC9_0),.dout(w_dff_B_TVLkAODu4_0),.clk(gclk));
	jdff dff_B_gssSvAKg1_0(.din(w_dff_B_TVLkAODu4_0),.dout(w_dff_B_gssSvAKg1_0),.clk(gclk));
	jdff dff_B_Nt8AkM2W0_0(.din(w_dff_B_gssSvAKg1_0),.dout(w_dff_B_Nt8AkM2W0_0),.clk(gclk));
	jdff dff_B_uW15OETl6_0(.din(w_dff_B_Nt8AkM2W0_0),.dout(w_dff_B_uW15OETl6_0),.clk(gclk));
	jdff dff_B_OSrkWgmF6_0(.din(w_dff_B_uW15OETl6_0),.dout(w_dff_B_OSrkWgmF6_0),.clk(gclk));
	jdff dff_B_5WZOjuU90_0(.din(w_dff_B_OSrkWgmF6_0),.dout(w_dff_B_5WZOjuU90_0),.clk(gclk));
	jdff dff_B_zRNUK3wv8_0(.din(w_dff_B_5WZOjuU90_0),.dout(w_dff_B_zRNUK3wv8_0),.clk(gclk));
	jdff dff_B_rx6J8DIR6_0(.din(w_dff_B_zRNUK3wv8_0),.dout(w_dff_B_rx6J8DIR6_0),.clk(gclk));
	jdff dff_B_T5e4P5jh1_0(.din(w_dff_B_rx6J8DIR6_0),.dout(w_dff_B_T5e4P5jh1_0),.clk(gclk));
	jdff dff_B_Tw7YyZQy8_0(.din(w_dff_B_T5e4P5jh1_0),.dout(w_dff_B_Tw7YyZQy8_0),.clk(gclk));
	jdff dff_B_qzOjTNJG6_0(.din(w_dff_B_Tw7YyZQy8_0),.dout(w_dff_B_qzOjTNJG6_0),.clk(gclk));
	jdff dff_B_cIeubwr68_0(.din(w_dff_B_qzOjTNJG6_0),.dout(w_dff_B_cIeubwr68_0),.clk(gclk));
	jdff dff_B_dOMyglfL4_0(.din(w_dff_B_cIeubwr68_0),.dout(w_dff_B_dOMyglfL4_0),.clk(gclk));
	jdff dff_B_r2oqDg6g1_0(.din(w_dff_B_dOMyglfL4_0),.dout(w_dff_B_r2oqDg6g1_0),.clk(gclk));
	jdff dff_B_DP5UyGLi3_0(.din(w_dff_B_r2oqDg6g1_0),.dout(w_dff_B_DP5UyGLi3_0),.clk(gclk));
	jdff dff_B_GOXbqGGt6_0(.din(w_dff_B_DP5UyGLi3_0),.dout(w_dff_B_GOXbqGGt6_0),.clk(gclk));
	jdff dff_B_qUf7scos5_0(.din(w_dff_B_GOXbqGGt6_0),.dout(w_dff_B_qUf7scos5_0),.clk(gclk));
	jdff dff_B_hXwger6Q0_0(.din(w_dff_B_qUf7scos5_0),.dout(w_dff_B_hXwger6Q0_0),.clk(gclk));
	jdff dff_B_qaG96RCx0_0(.din(w_dff_B_hXwger6Q0_0),.dout(w_dff_B_qaG96RCx0_0),.clk(gclk));
	jdff dff_B_jR6pJF6b9_0(.din(w_dff_B_qaG96RCx0_0),.dout(w_dff_B_jR6pJF6b9_0),.clk(gclk));
	jdff dff_B_hGWJW1Oi3_0(.din(w_dff_B_jR6pJF6b9_0),.dout(w_dff_B_hGWJW1Oi3_0),.clk(gclk));
	jdff dff_B_m69YFwVh8_0(.din(w_dff_B_hGWJW1Oi3_0),.dout(w_dff_B_m69YFwVh8_0),.clk(gclk));
	jdff dff_B_XP178ACT1_0(.din(w_dff_B_m69YFwVh8_0),.dout(w_dff_B_XP178ACT1_0),.clk(gclk));
	jdff dff_B_Tyz7FRDj5_0(.din(w_dff_B_XP178ACT1_0),.dout(w_dff_B_Tyz7FRDj5_0),.clk(gclk));
	jdff dff_B_Kvp7cwzZ7_0(.din(w_dff_B_Tyz7FRDj5_0),.dout(w_dff_B_Kvp7cwzZ7_0),.clk(gclk));
	jdff dff_B_WmtFT1UX8_0(.din(w_dff_B_Kvp7cwzZ7_0),.dout(w_dff_B_WmtFT1UX8_0),.clk(gclk));
	jdff dff_B_WaZiaEi05_0(.din(w_dff_B_WmtFT1UX8_0),.dout(w_dff_B_WaZiaEi05_0),.clk(gclk));
	jdff dff_B_YcrveNHU9_0(.din(w_dff_B_WaZiaEi05_0),.dout(w_dff_B_YcrveNHU9_0),.clk(gclk));
	jdff dff_B_XzUjWw8I8_0(.din(w_dff_B_YcrveNHU9_0),.dout(w_dff_B_XzUjWw8I8_0),.clk(gclk));
	jdff dff_B_ro1gLVvR6_0(.din(w_dff_B_XzUjWw8I8_0),.dout(w_dff_B_ro1gLVvR6_0),.clk(gclk));
	jdff dff_B_4x0fcnX07_0(.din(w_dff_B_ro1gLVvR6_0),.dout(w_dff_B_4x0fcnX07_0),.clk(gclk));
	jdff dff_B_ALyepbeq7_0(.din(w_dff_B_4x0fcnX07_0),.dout(w_dff_B_ALyepbeq7_0),.clk(gclk));
	jdff dff_B_f6iUujuk5_0(.din(w_dff_B_ALyepbeq7_0),.dout(w_dff_B_f6iUujuk5_0),.clk(gclk));
	jdff dff_B_IB6jH9PE8_0(.din(w_dff_B_f6iUujuk5_0),.dout(w_dff_B_IB6jH9PE8_0),.clk(gclk));
	jdff dff_B_g88kN3uI6_0(.din(w_dff_B_IB6jH9PE8_0),.dout(w_dff_B_g88kN3uI6_0),.clk(gclk));
	jdff dff_B_D4X58SKJ5_0(.din(w_dff_B_g88kN3uI6_0),.dout(w_dff_B_D4X58SKJ5_0),.clk(gclk));
	jdff dff_B_4nhufPn46_0(.din(w_dff_B_D4X58SKJ5_0),.dout(w_dff_B_4nhufPn46_0),.clk(gclk));
	jdff dff_B_ELMaxXhd1_0(.din(w_dff_B_4nhufPn46_0),.dout(w_dff_B_ELMaxXhd1_0),.clk(gclk));
	jdff dff_B_5GHwduaf2_0(.din(w_dff_B_ELMaxXhd1_0),.dout(w_dff_B_5GHwduaf2_0),.clk(gclk));
	jdff dff_B_hycexgJs7_0(.din(w_dff_B_5GHwduaf2_0),.dout(w_dff_B_hycexgJs7_0),.clk(gclk));
	jdff dff_B_9D3h1bEM0_0(.din(w_dff_B_hycexgJs7_0),.dout(w_dff_B_9D3h1bEM0_0),.clk(gclk));
	jdff dff_B_2w9i8F3i2_0(.din(w_dff_B_9D3h1bEM0_0),.dout(w_dff_B_2w9i8F3i2_0),.clk(gclk));
	jdff dff_B_eqgPPYbX5_0(.din(w_dff_B_2w9i8F3i2_0),.dout(w_dff_B_eqgPPYbX5_0),.clk(gclk));
	jdff dff_B_G5rtZoew6_0(.din(w_dff_B_eqgPPYbX5_0),.dout(w_dff_B_G5rtZoew6_0),.clk(gclk));
	jdff dff_B_v9otEqz79_0(.din(w_dff_B_G5rtZoew6_0),.dout(w_dff_B_v9otEqz79_0),.clk(gclk));
	jdff dff_B_Fe5Cztr34_0(.din(w_dff_B_v9otEqz79_0),.dout(w_dff_B_Fe5Cztr34_0),.clk(gclk));
	jdff dff_B_HluWOPtu2_0(.din(w_dff_B_Fe5Cztr34_0),.dout(w_dff_B_HluWOPtu2_0),.clk(gclk));
	jdff dff_B_4llKQOpS1_0(.din(w_dff_B_HluWOPtu2_0),.dout(w_dff_B_4llKQOpS1_0),.clk(gclk));
	jdff dff_B_Aog8pcXj5_0(.din(w_dff_B_4llKQOpS1_0),.dout(w_dff_B_Aog8pcXj5_0),.clk(gclk));
	jdff dff_B_hSYLk0sV3_0(.din(w_dff_B_Aog8pcXj5_0),.dout(w_dff_B_hSYLk0sV3_0),.clk(gclk));
	jdff dff_B_yRRRiyKJ6_0(.din(w_dff_B_hSYLk0sV3_0),.dout(w_dff_B_yRRRiyKJ6_0),.clk(gclk));
	jdff dff_B_95jaZ1ps3_0(.din(w_dff_B_yRRRiyKJ6_0),.dout(w_dff_B_95jaZ1ps3_0),.clk(gclk));
	jdff dff_B_vU336DFM7_0(.din(w_dff_B_95jaZ1ps3_0),.dout(w_dff_B_vU336DFM7_0),.clk(gclk));
	jdff dff_B_HyPNRr7b0_0(.din(w_dff_B_vU336DFM7_0),.dout(w_dff_B_HyPNRr7b0_0),.clk(gclk));
	jdff dff_B_aK28yDJq0_0(.din(w_dff_B_HyPNRr7b0_0),.dout(w_dff_B_aK28yDJq0_0),.clk(gclk));
	jdff dff_B_RNu8fyVC8_0(.din(w_dff_B_aK28yDJq0_0),.dout(w_dff_B_RNu8fyVC8_0),.clk(gclk));
	jdff dff_B_wzn4mPF53_0(.din(w_dff_B_RNu8fyVC8_0),.dout(w_dff_B_wzn4mPF53_0),.clk(gclk));
	jdff dff_B_bFsrc20v8_0(.din(w_dff_B_wzn4mPF53_0),.dout(w_dff_B_bFsrc20v8_0),.clk(gclk));
	jdff dff_B_7jmY5U6d3_0(.din(w_dff_B_bFsrc20v8_0),.dout(w_dff_B_7jmY5U6d3_0),.clk(gclk));
	jdff dff_B_w04qloms2_0(.din(w_dff_B_7jmY5U6d3_0),.dout(w_dff_B_w04qloms2_0),.clk(gclk));
	jdff dff_B_Hdq9eNO36_0(.din(w_dff_B_w04qloms2_0),.dout(w_dff_B_Hdq9eNO36_0),.clk(gclk));
	jdff dff_B_4tDfSGdR2_0(.din(w_dff_B_Hdq9eNO36_0),.dout(w_dff_B_4tDfSGdR2_0),.clk(gclk));
	jdff dff_B_SX4kGZlS9_0(.din(w_dff_B_4tDfSGdR2_0),.dout(w_dff_B_SX4kGZlS9_0),.clk(gclk));
	jdff dff_B_wm6uFC186_0(.din(w_dff_B_SX4kGZlS9_0),.dout(w_dff_B_wm6uFC186_0),.clk(gclk));
	jdff dff_B_jse6aP2y1_0(.din(w_dff_B_wm6uFC186_0),.dout(w_dff_B_jse6aP2y1_0),.clk(gclk));
	jdff dff_B_WKYHnQ064_0(.din(w_dff_B_jse6aP2y1_0),.dout(w_dff_B_WKYHnQ064_0),.clk(gclk));
	jdff dff_B_dW3bOQsl4_1(.din(n984),.dout(w_dff_B_dW3bOQsl4_1),.clk(gclk));
	jdff dff_B_EAtwghzA5_1(.din(w_dff_B_dW3bOQsl4_1),.dout(w_dff_B_EAtwghzA5_1),.clk(gclk));
	jdff dff_B_bZUiXPwS2_1(.din(w_dff_B_EAtwghzA5_1),.dout(w_dff_B_bZUiXPwS2_1),.clk(gclk));
	jdff dff_B_tqVeCLjJ6_1(.din(w_dff_B_bZUiXPwS2_1),.dout(w_dff_B_tqVeCLjJ6_1),.clk(gclk));
	jdff dff_B_TZVevdMK9_1(.din(w_dff_B_tqVeCLjJ6_1),.dout(w_dff_B_TZVevdMK9_1),.clk(gclk));
	jdff dff_B_JSUQAoxZ4_1(.din(w_dff_B_TZVevdMK9_1),.dout(w_dff_B_JSUQAoxZ4_1),.clk(gclk));
	jdff dff_B_vzk5YVgY7_1(.din(w_dff_B_JSUQAoxZ4_1),.dout(w_dff_B_vzk5YVgY7_1),.clk(gclk));
	jdff dff_B_ahVDdP2N6_1(.din(w_dff_B_vzk5YVgY7_1),.dout(w_dff_B_ahVDdP2N6_1),.clk(gclk));
	jdff dff_B_ZxNxXE353_1(.din(w_dff_B_ahVDdP2N6_1),.dout(w_dff_B_ZxNxXE353_1),.clk(gclk));
	jdff dff_B_cd5oMpdK5_1(.din(w_dff_B_ZxNxXE353_1),.dout(w_dff_B_cd5oMpdK5_1),.clk(gclk));
	jdff dff_B_eVM8NMRf2_1(.din(w_dff_B_cd5oMpdK5_1),.dout(w_dff_B_eVM8NMRf2_1),.clk(gclk));
	jdff dff_B_ZhpnEFfF8_1(.din(w_dff_B_eVM8NMRf2_1),.dout(w_dff_B_ZhpnEFfF8_1),.clk(gclk));
	jdff dff_B_Ft4cEAzk5_1(.din(w_dff_B_ZhpnEFfF8_1),.dout(w_dff_B_Ft4cEAzk5_1),.clk(gclk));
	jdff dff_B_dHnhehqL8_1(.din(w_dff_B_Ft4cEAzk5_1),.dout(w_dff_B_dHnhehqL8_1),.clk(gclk));
	jdff dff_B_0hhvlaJU9_1(.din(w_dff_B_dHnhehqL8_1),.dout(w_dff_B_0hhvlaJU9_1),.clk(gclk));
	jdff dff_B_Z2f1xnDL8_1(.din(w_dff_B_0hhvlaJU9_1),.dout(w_dff_B_Z2f1xnDL8_1),.clk(gclk));
	jdff dff_B_ACiDnWhG9_1(.din(w_dff_B_Z2f1xnDL8_1),.dout(w_dff_B_ACiDnWhG9_1),.clk(gclk));
	jdff dff_B_H9atbfUk1_1(.din(w_dff_B_ACiDnWhG9_1),.dout(w_dff_B_H9atbfUk1_1),.clk(gclk));
	jdff dff_B_z6reGHio0_1(.din(w_dff_B_H9atbfUk1_1),.dout(w_dff_B_z6reGHio0_1),.clk(gclk));
	jdff dff_B_8prjGHfW0_1(.din(w_dff_B_z6reGHio0_1),.dout(w_dff_B_8prjGHfW0_1),.clk(gclk));
	jdff dff_B_6PZ9zAgl7_1(.din(w_dff_B_8prjGHfW0_1),.dout(w_dff_B_6PZ9zAgl7_1),.clk(gclk));
	jdff dff_B_404R34Wx4_1(.din(w_dff_B_6PZ9zAgl7_1),.dout(w_dff_B_404R34Wx4_1),.clk(gclk));
	jdff dff_B_QFVLQk999_1(.din(w_dff_B_404R34Wx4_1),.dout(w_dff_B_QFVLQk999_1),.clk(gclk));
	jdff dff_B_ZdvJztze0_1(.din(w_dff_B_QFVLQk999_1),.dout(w_dff_B_ZdvJztze0_1),.clk(gclk));
	jdff dff_B_jtUU8lLt4_1(.din(w_dff_B_ZdvJztze0_1),.dout(w_dff_B_jtUU8lLt4_1),.clk(gclk));
	jdff dff_B_ErfJELrv8_1(.din(w_dff_B_jtUU8lLt4_1),.dout(w_dff_B_ErfJELrv8_1),.clk(gclk));
	jdff dff_B_SfgdcvMN5_1(.din(w_dff_B_ErfJELrv8_1),.dout(w_dff_B_SfgdcvMN5_1),.clk(gclk));
	jdff dff_B_y6mhtZWH9_1(.din(w_dff_B_SfgdcvMN5_1),.dout(w_dff_B_y6mhtZWH9_1),.clk(gclk));
	jdff dff_B_SxZQYWiU0_1(.din(w_dff_B_y6mhtZWH9_1),.dout(w_dff_B_SxZQYWiU0_1),.clk(gclk));
	jdff dff_B_Ym66mhjs3_1(.din(w_dff_B_SxZQYWiU0_1),.dout(w_dff_B_Ym66mhjs3_1),.clk(gclk));
	jdff dff_B_zk0lrBTR9_1(.din(w_dff_B_Ym66mhjs3_1),.dout(w_dff_B_zk0lrBTR9_1),.clk(gclk));
	jdff dff_B_sBKj8tvH3_1(.din(w_dff_B_zk0lrBTR9_1),.dout(w_dff_B_sBKj8tvH3_1),.clk(gclk));
	jdff dff_B_9RGFGaUs8_1(.din(w_dff_B_sBKj8tvH3_1),.dout(w_dff_B_9RGFGaUs8_1),.clk(gclk));
	jdff dff_B_b8F8wylu8_1(.din(w_dff_B_9RGFGaUs8_1),.dout(w_dff_B_b8F8wylu8_1),.clk(gclk));
	jdff dff_B_FoGxaiXO7_1(.din(w_dff_B_b8F8wylu8_1),.dout(w_dff_B_FoGxaiXO7_1),.clk(gclk));
	jdff dff_B_htFtFf5k4_1(.din(w_dff_B_FoGxaiXO7_1),.dout(w_dff_B_htFtFf5k4_1),.clk(gclk));
	jdff dff_B_efNeOYOv9_1(.din(w_dff_B_htFtFf5k4_1),.dout(w_dff_B_efNeOYOv9_1),.clk(gclk));
	jdff dff_B_nb21rX101_1(.din(w_dff_B_efNeOYOv9_1),.dout(w_dff_B_nb21rX101_1),.clk(gclk));
	jdff dff_B_cyE9GT2i1_1(.din(w_dff_B_nb21rX101_1),.dout(w_dff_B_cyE9GT2i1_1),.clk(gclk));
	jdff dff_B_H3vbTa5N0_1(.din(w_dff_B_cyE9GT2i1_1),.dout(w_dff_B_H3vbTa5N0_1),.clk(gclk));
	jdff dff_B_0K4W2rfU6_1(.din(w_dff_B_H3vbTa5N0_1),.dout(w_dff_B_0K4W2rfU6_1),.clk(gclk));
	jdff dff_B_fU3HWTrg4_1(.din(w_dff_B_0K4W2rfU6_1),.dout(w_dff_B_fU3HWTrg4_1),.clk(gclk));
	jdff dff_B_CEJbSzhb7_1(.din(w_dff_B_fU3HWTrg4_1),.dout(w_dff_B_CEJbSzhb7_1),.clk(gclk));
	jdff dff_B_Ha899IwM9_1(.din(w_dff_B_CEJbSzhb7_1),.dout(w_dff_B_Ha899IwM9_1),.clk(gclk));
	jdff dff_B_q3iHuL7x8_1(.din(w_dff_B_Ha899IwM9_1),.dout(w_dff_B_q3iHuL7x8_1),.clk(gclk));
	jdff dff_B_rWaVp7W00_1(.din(w_dff_B_q3iHuL7x8_1),.dout(w_dff_B_rWaVp7W00_1),.clk(gclk));
	jdff dff_B_V6nJ2JND0_1(.din(w_dff_B_rWaVp7W00_1),.dout(w_dff_B_V6nJ2JND0_1),.clk(gclk));
	jdff dff_B_tKpXAavf9_1(.din(w_dff_B_V6nJ2JND0_1),.dout(w_dff_B_tKpXAavf9_1),.clk(gclk));
	jdff dff_B_W9iXaONO1_1(.din(w_dff_B_tKpXAavf9_1),.dout(w_dff_B_W9iXaONO1_1),.clk(gclk));
	jdff dff_B_dhxVqzlD7_1(.din(w_dff_B_W9iXaONO1_1),.dout(w_dff_B_dhxVqzlD7_1),.clk(gclk));
	jdff dff_B_U7TsXFN70_1(.din(w_dff_B_dhxVqzlD7_1),.dout(w_dff_B_U7TsXFN70_1),.clk(gclk));
	jdff dff_B_41vyKhgg0_1(.din(w_dff_B_U7TsXFN70_1),.dout(w_dff_B_41vyKhgg0_1),.clk(gclk));
	jdff dff_B_CGViD9Ra2_1(.din(w_dff_B_41vyKhgg0_1),.dout(w_dff_B_CGViD9Ra2_1),.clk(gclk));
	jdff dff_B_VlY5E9vk3_1(.din(w_dff_B_CGViD9Ra2_1),.dout(w_dff_B_VlY5E9vk3_1),.clk(gclk));
	jdff dff_B_PfXaZAgN8_1(.din(w_dff_B_VlY5E9vk3_1),.dout(w_dff_B_PfXaZAgN8_1),.clk(gclk));
	jdff dff_B_RHPfq9Ac8_1(.din(w_dff_B_PfXaZAgN8_1),.dout(w_dff_B_RHPfq9Ac8_1),.clk(gclk));
	jdff dff_B_PM0i3fPu5_1(.din(w_dff_B_RHPfq9Ac8_1),.dout(w_dff_B_PM0i3fPu5_1),.clk(gclk));
	jdff dff_B_qwWAUPHb8_1(.din(w_dff_B_PM0i3fPu5_1),.dout(w_dff_B_qwWAUPHb8_1),.clk(gclk));
	jdff dff_B_6ndAXiJ42_1(.din(w_dff_B_qwWAUPHb8_1),.dout(w_dff_B_6ndAXiJ42_1),.clk(gclk));
	jdff dff_B_P4W8IZrJ2_1(.din(w_dff_B_6ndAXiJ42_1),.dout(w_dff_B_P4W8IZrJ2_1),.clk(gclk));
	jdff dff_B_rtr0nblm8_1(.din(w_dff_B_P4W8IZrJ2_1),.dout(w_dff_B_rtr0nblm8_1),.clk(gclk));
	jdff dff_B_48IR0VUc0_1(.din(w_dff_B_rtr0nblm8_1),.dout(w_dff_B_48IR0VUc0_1),.clk(gclk));
	jdff dff_B_Cl5xRC565_1(.din(w_dff_B_48IR0VUc0_1),.dout(w_dff_B_Cl5xRC565_1),.clk(gclk));
	jdff dff_B_tm8WBy4I7_1(.din(w_dff_B_Cl5xRC565_1),.dout(w_dff_B_tm8WBy4I7_1),.clk(gclk));
	jdff dff_B_yFhqCxz27_1(.din(w_dff_B_tm8WBy4I7_1),.dout(w_dff_B_yFhqCxz27_1),.clk(gclk));
	jdff dff_B_Tlc9wAFJ4_1(.din(w_dff_B_yFhqCxz27_1),.dout(w_dff_B_Tlc9wAFJ4_1),.clk(gclk));
	jdff dff_B_Sc1HFL605_1(.din(w_dff_B_Tlc9wAFJ4_1),.dout(w_dff_B_Sc1HFL605_1),.clk(gclk));
	jdff dff_B_QzYujono6_1(.din(w_dff_B_Sc1HFL605_1),.dout(w_dff_B_QzYujono6_1),.clk(gclk));
	jdff dff_B_ST20qWtV2_1(.din(w_dff_B_QzYujono6_1),.dout(w_dff_B_ST20qWtV2_1),.clk(gclk));
	jdff dff_B_IMsnHKjp4_1(.din(w_dff_B_ST20qWtV2_1),.dout(w_dff_B_IMsnHKjp4_1),.clk(gclk));
	jdff dff_B_eEqRptMH7_1(.din(w_dff_B_IMsnHKjp4_1),.dout(w_dff_B_eEqRptMH7_1),.clk(gclk));
	jdff dff_B_tEtvD5pC8_1(.din(w_dff_B_eEqRptMH7_1),.dout(w_dff_B_tEtvD5pC8_1),.clk(gclk));
	jdff dff_B_PkbUtv1R1_1(.din(w_dff_B_tEtvD5pC8_1),.dout(w_dff_B_PkbUtv1R1_1),.clk(gclk));
	jdff dff_B_XQiqryRZ3_1(.din(w_dff_B_PkbUtv1R1_1),.dout(w_dff_B_XQiqryRZ3_1),.clk(gclk));
	jdff dff_B_u1hQWf5a5_1(.din(w_dff_B_XQiqryRZ3_1),.dout(w_dff_B_u1hQWf5a5_1),.clk(gclk));
	jdff dff_B_QPZUVCc46_1(.din(w_dff_B_u1hQWf5a5_1),.dout(w_dff_B_QPZUVCc46_1),.clk(gclk));
	jdff dff_B_VcIic6js6_1(.din(w_dff_B_QPZUVCc46_1),.dout(w_dff_B_VcIic6js6_1),.clk(gclk));
	jdff dff_B_ZVojjKw26_1(.din(w_dff_B_VcIic6js6_1),.dout(w_dff_B_ZVojjKw26_1),.clk(gclk));
	jdff dff_B_ZM3RHWZj3_1(.din(w_dff_B_ZVojjKw26_1),.dout(w_dff_B_ZM3RHWZj3_1),.clk(gclk));
	jdff dff_B_nMZBmZ6Y5_1(.din(w_dff_B_ZM3RHWZj3_1),.dout(w_dff_B_nMZBmZ6Y5_1),.clk(gclk));
	jdff dff_B_KxGC3tHv5_1(.din(w_dff_B_nMZBmZ6Y5_1),.dout(w_dff_B_KxGC3tHv5_1),.clk(gclk));
	jdff dff_B_46pT0eQ89_1(.din(w_dff_B_KxGC3tHv5_1),.dout(w_dff_B_46pT0eQ89_1),.clk(gclk));
	jdff dff_B_PQ9oIgaA7_1(.din(w_dff_B_46pT0eQ89_1),.dout(w_dff_B_PQ9oIgaA7_1),.clk(gclk));
	jdff dff_B_Z0StsYyh3_1(.din(w_dff_B_PQ9oIgaA7_1),.dout(w_dff_B_Z0StsYyh3_1),.clk(gclk));
	jdff dff_B_iZeFzGdY0_1(.din(w_dff_B_Z0StsYyh3_1),.dout(w_dff_B_iZeFzGdY0_1),.clk(gclk));
	jdff dff_B_eEUI45IG3_1(.din(w_dff_B_iZeFzGdY0_1),.dout(w_dff_B_eEUI45IG3_1),.clk(gclk));
	jdff dff_B_j1mj19K26_1(.din(w_dff_B_eEUI45IG3_1),.dout(w_dff_B_j1mj19K26_1),.clk(gclk));
	jdff dff_B_NIH6EfS74_1(.din(w_dff_B_j1mj19K26_1),.dout(w_dff_B_NIH6EfS74_1),.clk(gclk));
	jdff dff_B_iwPjKlG56_1(.din(w_dff_B_NIH6EfS74_1),.dout(w_dff_B_iwPjKlG56_1),.clk(gclk));
	jdff dff_B_8mtLIjRB2_1(.din(w_dff_B_iwPjKlG56_1),.dout(w_dff_B_8mtLIjRB2_1),.clk(gclk));
	jdff dff_B_aWVqOKkb0_1(.din(w_dff_B_8mtLIjRB2_1),.dout(w_dff_B_aWVqOKkb0_1),.clk(gclk));
	jdff dff_B_U5fTCsZj0_1(.din(w_dff_B_aWVqOKkb0_1),.dout(w_dff_B_U5fTCsZj0_1),.clk(gclk));
	jdff dff_B_1CDbxVMk3_1(.din(w_dff_B_U5fTCsZj0_1),.dout(w_dff_B_1CDbxVMk3_1),.clk(gclk));
	jdff dff_B_OhiKHpSY6_1(.din(w_dff_B_1CDbxVMk3_1),.dout(w_dff_B_OhiKHpSY6_1),.clk(gclk));
	jdff dff_B_pPjbgOal2_1(.din(w_dff_B_OhiKHpSY6_1),.dout(w_dff_B_pPjbgOal2_1),.clk(gclk));
	jdff dff_B_9L9tzgWz6_1(.din(w_dff_B_pPjbgOal2_1),.dout(w_dff_B_9L9tzgWz6_1),.clk(gclk));
	jdff dff_B_bHi0BR043_1(.din(w_dff_B_9L9tzgWz6_1),.dout(w_dff_B_bHi0BR043_1),.clk(gclk));
	jdff dff_B_5Nk4raz90_1(.din(w_dff_B_bHi0BR043_1),.dout(w_dff_B_5Nk4raz90_1),.clk(gclk));
	jdff dff_B_JYPc6Jnl2_1(.din(w_dff_B_5Nk4raz90_1),.dout(w_dff_B_JYPc6Jnl2_1),.clk(gclk));
	jdff dff_B_ihOKXM3G5_1(.din(w_dff_B_JYPc6Jnl2_1),.dout(w_dff_B_ihOKXM3G5_1),.clk(gclk));
	jdff dff_B_eEkl9s2m0_0(.din(n985),.dout(w_dff_B_eEkl9s2m0_0),.clk(gclk));
	jdff dff_B_D8KUBLF05_0(.din(w_dff_B_eEkl9s2m0_0),.dout(w_dff_B_D8KUBLF05_0),.clk(gclk));
	jdff dff_B_qf2xbpia8_0(.din(w_dff_B_D8KUBLF05_0),.dout(w_dff_B_qf2xbpia8_0),.clk(gclk));
	jdff dff_B_cF2Sw4nS1_0(.din(w_dff_B_qf2xbpia8_0),.dout(w_dff_B_cF2Sw4nS1_0),.clk(gclk));
	jdff dff_B_F8K1U4a32_0(.din(w_dff_B_cF2Sw4nS1_0),.dout(w_dff_B_F8K1U4a32_0),.clk(gclk));
	jdff dff_B_gzVC7ztD2_0(.din(w_dff_B_F8K1U4a32_0),.dout(w_dff_B_gzVC7ztD2_0),.clk(gclk));
	jdff dff_B_kfUrLfsQ6_0(.din(w_dff_B_gzVC7ztD2_0),.dout(w_dff_B_kfUrLfsQ6_0),.clk(gclk));
	jdff dff_B_dK0S79aT7_0(.din(w_dff_B_kfUrLfsQ6_0),.dout(w_dff_B_dK0S79aT7_0),.clk(gclk));
	jdff dff_B_x0nMv34b8_0(.din(w_dff_B_dK0S79aT7_0),.dout(w_dff_B_x0nMv34b8_0),.clk(gclk));
	jdff dff_B_eyLtVXlI7_0(.din(w_dff_B_x0nMv34b8_0),.dout(w_dff_B_eyLtVXlI7_0),.clk(gclk));
	jdff dff_B_X5hgcZze5_0(.din(w_dff_B_eyLtVXlI7_0),.dout(w_dff_B_X5hgcZze5_0),.clk(gclk));
	jdff dff_B_Pz5HTgqD6_0(.din(w_dff_B_X5hgcZze5_0),.dout(w_dff_B_Pz5HTgqD6_0),.clk(gclk));
	jdff dff_B_y4rYCSiz6_0(.din(w_dff_B_Pz5HTgqD6_0),.dout(w_dff_B_y4rYCSiz6_0),.clk(gclk));
	jdff dff_B_6ThmlYtL4_0(.din(w_dff_B_y4rYCSiz6_0),.dout(w_dff_B_6ThmlYtL4_0),.clk(gclk));
	jdff dff_B_Qt5IzyyR1_0(.din(w_dff_B_6ThmlYtL4_0),.dout(w_dff_B_Qt5IzyyR1_0),.clk(gclk));
	jdff dff_B_ObpYJLW88_0(.din(w_dff_B_Qt5IzyyR1_0),.dout(w_dff_B_ObpYJLW88_0),.clk(gclk));
	jdff dff_B_bHDtyw2h2_0(.din(w_dff_B_ObpYJLW88_0),.dout(w_dff_B_bHDtyw2h2_0),.clk(gclk));
	jdff dff_B_Rq0JrPuX7_0(.din(w_dff_B_bHDtyw2h2_0),.dout(w_dff_B_Rq0JrPuX7_0),.clk(gclk));
	jdff dff_B_F34YsqpI4_0(.din(w_dff_B_Rq0JrPuX7_0),.dout(w_dff_B_F34YsqpI4_0),.clk(gclk));
	jdff dff_B_eDZTykKZ1_0(.din(w_dff_B_F34YsqpI4_0),.dout(w_dff_B_eDZTykKZ1_0),.clk(gclk));
	jdff dff_B_x5VNB92I5_0(.din(w_dff_B_eDZTykKZ1_0),.dout(w_dff_B_x5VNB92I5_0),.clk(gclk));
	jdff dff_B_aI8VEOIL6_0(.din(w_dff_B_x5VNB92I5_0),.dout(w_dff_B_aI8VEOIL6_0),.clk(gclk));
	jdff dff_B_etFAJqn31_0(.din(w_dff_B_aI8VEOIL6_0),.dout(w_dff_B_etFAJqn31_0),.clk(gclk));
	jdff dff_B_MHIml8f18_0(.din(w_dff_B_etFAJqn31_0),.dout(w_dff_B_MHIml8f18_0),.clk(gclk));
	jdff dff_B_1atySNUl8_0(.din(w_dff_B_MHIml8f18_0),.dout(w_dff_B_1atySNUl8_0),.clk(gclk));
	jdff dff_B_FdquoYvk6_0(.din(w_dff_B_1atySNUl8_0),.dout(w_dff_B_FdquoYvk6_0),.clk(gclk));
	jdff dff_B_CFKLh3J16_0(.din(w_dff_B_FdquoYvk6_0),.dout(w_dff_B_CFKLh3J16_0),.clk(gclk));
	jdff dff_B_yENi3WCZ7_0(.din(w_dff_B_CFKLh3J16_0),.dout(w_dff_B_yENi3WCZ7_0),.clk(gclk));
	jdff dff_B_279KTDcr6_0(.din(w_dff_B_yENi3WCZ7_0),.dout(w_dff_B_279KTDcr6_0),.clk(gclk));
	jdff dff_B_ovzb43mE2_0(.din(w_dff_B_279KTDcr6_0),.dout(w_dff_B_ovzb43mE2_0),.clk(gclk));
	jdff dff_B_KWKTiTHN0_0(.din(w_dff_B_ovzb43mE2_0),.dout(w_dff_B_KWKTiTHN0_0),.clk(gclk));
	jdff dff_B_9z2B29rq6_0(.din(w_dff_B_KWKTiTHN0_0),.dout(w_dff_B_9z2B29rq6_0),.clk(gclk));
	jdff dff_B_evTDnltg1_0(.din(w_dff_B_9z2B29rq6_0),.dout(w_dff_B_evTDnltg1_0),.clk(gclk));
	jdff dff_B_rTLjHJzu6_0(.din(w_dff_B_evTDnltg1_0),.dout(w_dff_B_rTLjHJzu6_0),.clk(gclk));
	jdff dff_B_zlJc4Iql7_0(.din(w_dff_B_rTLjHJzu6_0),.dout(w_dff_B_zlJc4Iql7_0),.clk(gclk));
	jdff dff_B_BRXTv2Ar3_0(.din(w_dff_B_zlJc4Iql7_0),.dout(w_dff_B_BRXTv2Ar3_0),.clk(gclk));
	jdff dff_B_8ew50BET9_0(.din(w_dff_B_BRXTv2Ar3_0),.dout(w_dff_B_8ew50BET9_0),.clk(gclk));
	jdff dff_B_Jvy36XlD1_0(.din(w_dff_B_8ew50BET9_0),.dout(w_dff_B_Jvy36XlD1_0),.clk(gclk));
	jdff dff_B_Gzfj7Rtr1_0(.din(w_dff_B_Jvy36XlD1_0),.dout(w_dff_B_Gzfj7Rtr1_0),.clk(gclk));
	jdff dff_B_L9JCj7Nh2_0(.din(w_dff_B_Gzfj7Rtr1_0),.dout(w_dff_B_L9JCj7Nh2_0),.clk(gclk));
	jdff dff_B_DHosqy593_0(.din(w_dff_B_L9JCj7Nh2_0),.dout(w_dff_B_DHosqy593_0),.clk(gclk));
	jdff dff_B_4Vx0avMy9_0(.din(w_dff_B_DHosqy593_0),.dout(w_dff_B_4Vx0avMy9_0),.clk(gclk));
	jdff dff_B_9JBOmamy5_0(.din(w_dff_B_4Vx0avMy9_0),.dout(w_dff_B_9JBOmamy5_0),.clk(gclk));
	jdff dff_B_94Vg3t2Y5_0(.din(w_dff_B_9JBOmamy5_0),.dout(w_dff_B_94Vg3t2Y5_0),.clk(gclk));
	jdff dff_B_N0GTgjBi0_0(.din(w_dff_B_94Vg3t2Y5_0),.dout(w_dff_B_N0GTgjBi0_0),.clk(gclk));
	jdff dff_B_NAw1NFwm6_0(.din(w_dff_B_N0GTgjBi0_0),.dout(w_dff_B_NAw1NFwm6_0),.clk(gclk));
	jdff dff_B_SV7uZX0U3_0(.din(w_dff_B_NAw1NFwm6_0),.dout(w_dff_B_SV7uZX0U3_0),.clk(gclk));
	jdff dff_B_l3YsVBH02_0(.din(w_dff_B_SV7uZX0U3_0),.dout(w_dff_B_l3YsVBH02_0),.clk(gclk));
	jdff dff_B_r5fRi3ip8_0(.din(w_dff_B_l3YsVBH02_0),.dout(w_dff_B_r5fRi3ip8_0),.clk(gclk));
	jdff dff_B_ntCgpe8A0_0(.din(w_dff_B_r5fRi3ip8_0),.dout(w_dff_B_ntCgpe8A0_0),.clk(gclk));
	jdff dff_B_35GHKOE14_0(.din(w_dff_B_ntCgpe8A0_0),.dout(w_dff_B_35GHKOE14_0),.clk(gclk));
	jdff dff_B_FQSkhLyP4_0(.din(w_dff_B_35GHKOE14_0),.dout(w_dff_B_FQSkhLyP4_0),.clk(gclk));
	jdff dff_B_IvlD4qZH5_0(.din(w_dff_B_FQSkhLyP4_0),.dout(w_dff_B_IvlD4qZH5_0),.clk(gclk));
	jdff dff_B_SL43gV0Q9_0(.din(w_dff_B_IvlD4qZH5_0),.dout(w_dff_B_SL43gV0Q9_0),.clk(gclk));
	jdff dff_B_afRyoNGk8_0(.din(w_dff_B_SL43gV0Q9_0),.dout(w_dff_B_afRyoNGk8_0),.clk(gclk));
	jdff dff_B_88uefvSS1_0(.din(w_dff_B_afRyoNGk8_0),.dout(w_dff_B_88uefvSS1_0),.clk(gclk));
	jdff dff_B_kUwJ55Pl8_0(.din(w_dff_B_88uefvSS1_0),.dout(w_dff_B_kUwJ55Pl8_0),.clk(gclk));
	jdff dff_B_jyvSWpbW0_0(.din(w_dff_B_kUwJ55Pl8_0),.dout(w_dff_B_jyvSWpbW0_0),.clk(gclk));
	jdff dff_B_MHLF0uRC8_0(.din(w_dff_B_jyvSWpbW0_0),.dout(w_dff_B_MHLF0uRC8_0),.clk(gclk));
	jdff dff_B_mVgsqD6c4_0(.din(w_dff_B_MHLF0uRC8_0),.dout(w_dff_B_mVgsqD6c4_0),.clk(gclk));
	jdff dff_B_SClotsqa5_0(.din(w_dff_B_mVgsqD6c4_0),.dout(w_dff_B_SClotsqa5_0),.clk(gclk));
	jdff dff_B_LfPBmi6M8_0(.din(w_dff_B_SClotsqa5_0),.dout(w_dff_B_LfPBmi6M8_0),.clk(gclk));
	jdff dff_B_SJrdyF1v3_0(.din(w_dff_B_LfPBmi6M8_0),.dout(w_dff_B_SJrdyF1v3_0),.clk(gclk));
	jdff dff_B_X9qmn73p7_0(.din(w_dff_B_SJrdyF1v3_0),.dout(w_dff_B_X9qmn73p7_0),.clk(gclk));
	jdff dff_B_9jzDUsxY1_0(.din(w_dff_B_X9qmn73p7_0),.dout(w_dff_B_9jzDUsxY1_0),.clk(gclk));
	jdff dff_B_GRKnsCBI3_0(.din(w_dff_B_9jzDUsxY1_0),.dout(w_dff_B_GRKnsCBI3_0),.clk(gclk));
	jdff dff_B_caQ1HtKN7_0(.din(w_dff_B_GRKnsCBI3_0),.dout(w_dff_B_caQ1HtKN7_0),.clk(gclk));
	jdff dff_B_sWDZ9yAP0_0(.din(w_dff_B_caQ1HtKN7_0),.dout(w_dff_B_sWDZ9yAP0_0),.clk(gclk));
	jdff dff_B_FxuBYA3C1_0(.din(w_dff_B_sWDZ9yAP0_0),.dout(w_dff_B_FxuBYA3C1_0),.clk(gclk));
	jdff dff_B_AMLNUDZa6_0(.din(w_dff_B_FxuBYA3C1_0),.dout(w_dff_B_AMLNUDZa6_0),.clk(gclk));
	jdff dff_B_gL9ovFQ70_0(.din(w_dff_B_AMLNUDZa6_0),.dout(w_dff_B_gL9ovFQ70_0),.clk(gclk));
	jdff dff_B_v3OMlvve5_0(.din(w_dff_B_gL9ovFQ70_0),.dout(w_dff_B_v3OMlvve5_0),.clk(gclk));
	jdff dff_B_HTPqckhM9_0(.din(w_dff_B_v3OMlvve5_0),.dout(w_dff_B_HTPqckhM9_0),.clk(gclk));
	jdff dff_B_9mpvb3V42_0(.din(w_dff_B_HTPqckhM9_0),.dout(w_dff_B_9mpvb3V42_0),.clk(gclk));
	jdff dff_B_uhuyayo28_0(.din(w_dff_B_9mpvb3V42_0),.dout(w_dff_B_uhuyayo28_0),.clk(gclk));
	jdff dff_B_prU3UkQf5_0(.din(w_dff_B_uhuyayo28_0),.dout(w_dff_B_prU3UkQf5_0),.clk(gclk));
	jdff dff_B_fkAOM1JZ7_0(.din(w_dff_B_prU3UkQf5_0),.dout(w_dff_B_fkAOM1JZ7_0),.clk(gclk));
	jdff dff_B_n9KTjp973_0(.din(w_dff_B_fkAOM1JZ7_0),.dout(w_dff_B_n9KTjp973_0),.clk(gclk));
	jdff dff_B_s6T8f5YH9_0(.din(w_dff_B_n9KTjp973_0),.dout(w_dff_B_s6T8f5YH9_0),.clk(gclk));
	jdff dff_B_j09wXN7a2_0(.din(w_dff_B_s6T8f5YH9_0),.dout(w_dff_B_j09wXN7a2_0),.clk(gclk));
	jdff dff_B_vJFA0Str3_0(.din(w_dff_B_j09wXN7a2_0),.dout(w_dff_B_vJFA0Str3_0),.clk(gclk));
	jdff dff_B_MNoNaIff9_0(.din(w_dff_B_vJFA0Str3_0),.dout(w_dff_B_MNoNaIff9_0),.clk(gclk));
	jdff dff_B_sdvHJx4Z4_0(.din(w_dff_B_MNoNaIff9_0),.dout(w_dff_B_sdvHJx4Z4_0),.clk(gclk));
	jdff dff_B_DIOzZIet3_0(.din(w_dff_B_sdvHJx4Z4_0),.dout(w_dff_B_DIOzZIet3_0),.clk(gclk));
	jdff dff_B_Ly8V1W0a0_0(.din(w_dff_B_DIOzZIet3_0),.dout(w_dff_B_Ly8V1W0a0_0),.clk(gclk));
	jdff dff_B_K1JjLZHY3_0(.din(w_dff_B_Ly8V1W0a0_0),.dout(w_dff_B_K1JjLZHY3_0),.clk(gclk));
	jdff dff_B_z2W0T16R9_0(.din(w_dff_B_K1JjLZHY3_0),.dout(w_dff_B_z2W0T16R9_0),.clk(gclk));
	jdff dff_B_rAvTOp0k3_0(.din(w_dff_B_z2W0T16R9_0),.dout(w_dff_B_rAvTOp0k3_0),.clk(gclk));
	jdff dff_B_kHJmpJSC1_0(.din(w_dff_B_rAvTOp0k3_0),.dout(w_dff_B_kHJmpJSC1_0),.clk(gclk));
	jdff dff_B_tdDJgPSW1_0(.din(w_dff_B_kHJmpJSC1_0),.dout(w_dff_B_tdDJgPSW1_0),.clk(gclk));
	jdff dff_B_VVqaybmK0_0(.din(w_dff_B_tdDJgPSW1_0),.dout(w_dff_B_VVqaybmK0_0),.clk(gclk));
	jdff dff_B_hHQUy4MR1_0(.din(w_dff_B_VVqaybmK0_0),.dout(w_dff_B_hHQUy4MR1_0),.clk(gclk));
	jdff dff_B_5SgonsWr9_0(.din(w_dff_B_hHQUy4MR1_0),.dout(w_dff_B_5SgonsWr9_0),.clk(gclk));
	jdff dff_B_ut7QM3Hu0_0(.din(w_dff_B_5SgonsWr9_0),.dout(w_dff_B_ut7QM3Hu0_0),.clk(gclk));
	jdff dff_B_VHq0bp8e0_0(.din(w_dff_B_ut7QM3Hu0_0),.dout(w_dff_B_VHq0bp8e0_0),.clk(gclk));
	jdff dff_B_ACyBYY7T7_0(.din(w_dff_B_VHq0bp8e0_0),.dout(w_dff_B_ACyBYY7T7_0),.clk(gclk));
	jdff dff_B_YtryxROZ1_0(.din(w_dff_B_ACyBYY7T7_0),.dout(w_dff_B_YtryxROZ1_0),.clk(gclk));
	jdff dff_B_1a6uerT96_0(.din(w_dff_B_YtryxROZ1_0),.dout(w_dff_B_1a6uerT96_0),.clk(gclk));
	jdff dff_B_dYjiT6bc3_0(.din(w_dff_B_1a6uerT96_0),.dout(w_dff_B_dYjiT6bc3_0),.clk(gclk));
	jdff dff_B_ZBeU3nCK4_0(.din(w_dff_B_dYjiT6bc3_0),.dout(w_dff_B_ZBeU3nCK4_0),.clk(gclk));
	jdff dff_B_n82feeXJ6_1(.din(n978),.dout(w_dff_B_n82feeXJ6_1),.clk(gclk));
	jdff dff_B_WkAQ7u6W2_1(.din(w_dff_B_n82feeXJ6_1),.dout(w_dff_B_WkAQ7u6W2_1),.clk(gclk));
	jdff dff_B_Gy6kPcyJ2_1(.din(w_dff_B_WkAQ7u6W2_1),.dout(w_dff_B_Gy6kPcyJ2_1),.clk(gclk));
	jdff dff_B_0wgGlcsX2_1(.din(w_dff_B_Gy6kPcyJ2_1),.dout(w_dff_B_0wgGlcsX2_1),.clk(gclk));
	jdff dff_B_agtoXMUa0_1(.din(w_dff_B_0wgGlcsX2_1),.dout(w_dff_B_agtoXMUa0_1),.clk(gclk));
	jdff dff_B_7l8pwWSl6_1(.din(w_dff_B_agtoXMUa0_1),.dout(w_dff_B_7l8pwWSl6_1),.clk(gclk));
	jdff dff_B_tVJkpn0z3_1(.din(w_dff_B_7l8pwWSl6_1),.dout(w_dff_B_tVJkpn0z3_1),.clk(gclk));
	jdff dff_B_MfLCiWjv1_1(.din(w_dff_B_tVJkpn0z3_1),.dout(w_dff_B_MfLCiWjv1_1),.clk(gclk));
	jdff dff_B_6B6ifIgf0_1(.din(w_dff_B_MfLCiWjv1_1),.dout(w_dff_B_6B6ifIgf0_1),.clk(gclk));
	jdff dff_B_6Vvsb01V8_1(.din(w_dff_B_6B6ifIgf0_1),.dout(w_dff_B_6Vvsb01V8_1),.clk(gclk));
	jdff dff_B_JFGj1o086_1(.din(w_dff_B_6Vvsb01V8_1),.dout(w_dff_B_JFGj1o086_1),.clk(gclk));
	jdff dff_B_4kEhO6654_1(.din(w_dff_B_JFGj1o086_1),.dout(w_dff_B_4kEhO6654_1),.clk(gclk));
	jdff dff_B_gaFn8EE36_1(.din(w_dff_B_4kEhO6654_1),.dout(w_dff_B_gaFn8EE36_1),.clk(gclk));
	jdff dff_B_js56byEH9_1(.din(w_dff_B_gaFn8EE36_1),.dout(w_dff_B_js56byEH9_1),.clk(gclk));
	jdff dff_B_7FPHmqli1_1(.din(w_dff_B_js56byEH9_1),.dout(w_dff_B_7FPHmqli1_1),.clk(gclk));
	jdff dff_B_bNkFueRe3_1(.din(w_dff_B_7FPHmqli1_1),.dout(w_dff_B_bNkFueRe3_1),.clk(gclk));
	jdff dff_B_7tcyyuyz4_1(.din(w_dff_B_bNkFueRe3_1),.dout(w_dff_B_7tcyyuyz4_1),.clk(gclk));
	jdff dff_B_F14aY1DM8_1(.din(w_dff_B_7tcyyuyz4_1),.dout(w_dff_B_F14aY1DM8_1),.clk(gclk));
	jdff dff_B_vNrMpOOE0_1(.din(w_dff_B_F14aY1DM8_1),.dout(w_dff_B_vNrMpOOE0_1),.clk(gclk));
	jdff dff_B_U6VQecYl7_1(.din(w_dff_B_vNrMpOOE0_1),.dout(w_dff_B_U6VQecYl7_1),.clk(gclk));
	jdff dff_B_kVVFQFnb7_1(.din(w_dff_B_U6VQecYl7_1),.dout(w_dff_B_kVVFQFnb7_1),.clk(gclk));
	jdff dff_B_TfQjYiCO0_1(.din(w_dff_B_kVVFQFnb7_1),.dout(w_dff_B_TfQjYiCO0_1),.clk(gclk));
	jdff dff_B_FipZUJmv2_1(.din(w_dff_B_TfQjYiCO0_1),.dout(w_dff_B_FipZUJmv2_1),.clk(gclk));
	jdff dff_B_Ut6LkS6c3_1(.din(w_dff_B_FipZUJmv2_1),.dout(w_dff_B_Ut6LkS6c3_1),.clk(gclk));
	jdff dff_B_UiYvUax80_1(.din(w_dff_B_Ut6LkS6c3_1),.dout(w_dff_B_UiYvUax80_1),.clk(gclk));
	jdff dff_B_K0Lk56Wa1_1(.din(w_dff_B_UiYvUax80_1),.dout(w_dff_B_K0Lk56Wa1_1),.clk(gclk));
	jdff dff_B_Vqz7au1b1_1(.din(w_dff_B_K0Lk56Wa1_1),.dout(w_dff_B_Vqz7au1b1_1),.clk(gclk));
	jdff dff_B_C6rk0dxg7_1(.din(w_dff_B_Vqz7au1b1_1),.dout(w_dff_B_C6rk0dxg7_1),.clk(gclk));
	jdff dff_B_t9OXnGY12_1(.din(w_dff_B_C6rk0dxg7_1),.dout(w_dff_B_t9OXnGY12_1),.clk(gclk));
	jdff dff_B_0efPE6rr3_1(.din(w_dff_B_t9OXnGY12_1),.dout(w_dff_B_0efPE6rr3_1),.clk(gclk));
	jdff dff_B_HAJIT6Na0_1(.din(w_dff_B_0efPE6rr3_1),.dout(w_dff_B_HAJIT6Na0_1),.clk(gclk));
	jdff dff_B_jcnzE5Jb5_1(.din(w_dff_B_HAJIT6Na0_1),.dout(w_dff_B_jcnzE5Jb5_1),.clk(gclk));
	jdff dff_B_h02VGJpv7_1(.din(w_dff_B_jcnzE5Jb5_1),.dout(w_dff_B_h02VGJpv7_1),.clk(gclk));
	jdff dff_B_rMtvu2vC1_1(.din(w_dff_B_h02VGJpv7_1),.dout(w_dff_B_rMtvu2vC1_1),.clk(gclk));
	jdff dff_B_t1jv47dd1_1(.din(w_dff_B_rMtvu2vC1_1),.dout(w_dff_B_t1jv47dd1_1),.clk(gclk));
	jdff dff_B_X7HolBmJ8_1(.din(w_dff_B_t1jv47dd1_1),.dout(w_dff_B_X7HolBmJ8_1),.clk(gclk));
	jdff dff_B_DQgBa13G7_1(.din(w_dff_B_X7HolBmJ8_1),.dout(w_dff_B_DQgBa13G7_1),.clk(gclk));
	jdff dff_B_g5DcuphP8_1(.din(w_dff_B_DQgBa13G7_1),.dout(w_dff_B_g5DcuphP8_1),.clk(gclk));
	jdff dff_B_cwx6rjzh1_1(.din(w_dff_B_g5DcuphP8_1),.dout(w_dff_B_cwx6rjzh1_1),.clk(gclk));
	jdff dff_B_sAG6e7xv6_1(.din(w_dff_B_cwx6rjzh1_1),.dout(w_dff_B_sAG6e7xv6_1),.clk(gclk));
	jdff dff_B_n8VY4oYC7_1(.din(w_dff_B_sAG6e7xv6_1),.dout(w_dff_B_n8VY4oYC7_1),.clk(gclk));
	jdff dff_B_JnI5wO649_1(.din(w_dff_B_n8VY4oYC7_1),.dout(w_dff_B_JnI5wO649_1),.clk(gclk));
	jdff dff_B_97GSGcyp0_1(.din(w_dff_B_JnI5wO649_1),.dout(w_dff_B_97GSGcyp0_1),.clk(gclk));
	jdff dff_B_VH4azXFr3_1(.din(w_dff_B_97GSGcyp0_1),.dout(w_dff_B_VH4azXFr3_1),.clk(gclk));
	jdff dff_B_zasPMfwE5_1(.din(w_dff_B_VH4azXFr3_1),.dout(w_dff_B_zasPMfwE5_1),.clk(gclk));
	jdff dff_B_6Y1kiCmQ0_1(.din(w_dff_B_zasPMfwE5_1),.dout(w_dff_B_6Y1kiCmQ0_1),.clk(gclk));
	jdff dff_B_Uyk3Gpn20_1(.din(w_dff_B_6Y1kiCmQ0_1),.dout(w_dff_B_Uyk3Gpn20_1),.clk(gclk));
	jdff dff_B_DyElRSxN3_1(.din(w_dff_B_Uyk3Gpn20_1),.dout(w_dff_B_DyElRSxN3_1),.clk(gclk));
	jdff dff_B_2yGZeXi54_1(.din(w_dff_B_DyElRSxN3_1),.dout(w_dff_B_2yGZeXi54_1),.clk(gclk));
	jdff dff_B_615Gw5Dn4_1(.din(w_dff_B_2yGZeXi54_1),.dout(w_dff_B_615Gw5Dn4_1),.clk(gclk));
	jdff dff_B_YY4UgXBP1_1(.din(w_dff_B_615Gw5Dn4_1),.dout(w_dff_B_YY4UgXBP1_1),.clk(gclk));
	jdff dff_B_geC9abhG8_1(.din(w_dff_B_YY4UgXBP1_1),.dout(w_dff_B_geC9abhG8_1),.clk(gclk));
	jdff dff_B_wJW0CYU81_1(.din(w_dff_B_geC9abhG8_1),.dout(w_dff_B_wJW0CYU81_1),.clk(gclk));
	jdff dff_B_Hdfepvd84_1(.din(w_dff_B_wJW0CYU81_1),.dout(w_dff_B_Hdfepvd84_1),.clk(gclk));
	jdff dff_B_pRnUMcW69_1(.din(w_dff_B_Hdfepvd84_1),.dout(w_dff_B_pRnUMcW69_1),.clk(gclk));
	jdff dff_B_NzppTr7Z4_1(.din(w_dff_B_pRnUMcW69_1),.dout(w_dff_B_NzppTr7Z4_1),.clk(gclk));
	jdff dff_B_6LFlVRea8_1(.din(w_dff_B_NzppTr7Z4_1),.dout(w_dff_B_6LFlVRea8_1),.clk(gclk));
	jdff dff_B_eBTKs3XB0_1(.din(w_dff_B_6LFlVRea8_1),.dout(w_dff_B_eBTKs3XB0_1),.clk(gclk));
	jdff dff_B_oGBfP9N66_1(.din(w_dff_B_eBTKs3XB0_1),.dout(w_dff_B_oGBfP9N66_1),.clk(gclk));
	jdff dff_B_O5hCadVz8_1(.din(w_dff_B_oGBfP9N66_1),.dout(w_dff_B_O5hCadVz8_1),.clk(gclk));
	jdff dff_B_2Kb5B5Pe9_1(.din(w_dff_B_O5hCadVz8_1),.dout(w_dff_B_2Kb5B5Pe9_1),.clk(gclk));
	jdff dff_B_vbs6i2S92_1(.din(w_dff_B_2Kb5B5Pe9_1),.dout(w_dff_B_vbs6i2S92_1),.clk(gclk));
	jdff dff_B_Ci4Wnzv17_1(.din(w_dff_B_vbs6i2S92_1),.dout(w_dff_B_Ci4Wnzv17_1),.clk(gclk));
	jdff dff_B_Yxo4r10Z5_1(.din(w_dff_B_Ci4Wnzv17_1),.dout(w_dff_B_Yxo4r10Z5_1),.clk(gclk));
	jdff dff_B_F5hhH1ky1_1(.din(w_dff_B_Yxo4r10Z5_1),.dout(w_dff_B_F5hhH1ky1_1),.clk(gclk));
	jdff dff_B_ZrPO1EYw8_1(.din(w_dff_B_F5hhH1ky1_1),.dout(w_dff_B_ZrPO1EYw8_1),.clk(gclk));
	jdff dff_B_NHXs0VmM5_1(.din(w_dff_B_ZrPO1EYw8_1),.dout(w_dff_B_NHXs0VmM5_1),.clk(gclk));
	jdff dff_B_pJnEtqX11_1(.din(w_dff_B_NHXs0VmM5_1),.dout(w_dff_B_pJnEtqX11_1),.clk(gclk));
	jdff dff_B_JAiFItIv1_1(.din(w_dff_B_pJnEtqX11_1),.dout(w_dff_B_JAiFItIv1_1),.clk(gclk));
	jdff dff_B_aWURpxMI8_1(.din(w_dff_B_JAiFItIv1_1),.dout(w_dff_B_aWURpxMI8_1),.clk(gclk));
	jdff dff_B_RD3jpQJC6_1(.din(w_dff_B_aWURpxMI8_1),.dout(w_dff_B_RD3jpQJC6_1),.clk(gclk));
	jdff dff_B_fjmJSJfd4_1(.din(w_dff_B_RD3jpQJC6_1),.dout(w_dff_B_fjmJSJfd4_1),.clk(gclk));
	jdff dff_B_WSqCwYOX8_1(.din(w_dff_B_fjmJSJfd4_1),.dout(w_dff_B_WSqCwYOX8_1),.clk(gclk));
	jdff dff_B_3IJIS5TI0_1(.din(w_dff_B_WSqCwYOX8_1),.dout(w_dff_B_3IJIS5TI0_1),.clk(gclk));
	jdff dff_B_KkQQOTJO7_1(.din(w_dff_B_3IJIS5TI0_1),.dout(w_dff_B_KkQQOTJO7_1),.clk(gclk));
	jdff dff_B_yRMPGGna3_1(.din(w_dff_B_KkQQOTJO7_1),.dout(w_dff_B_yRMPGGna3_1),.clk(gclk));
	jdff dff_B_1b4SG3UD4_1(.din(w_dff_B_yRMPGGna3_1),.dout(w_dff_B_1b4SG3UD4_1),.clk(gclk));
	jdff dff_B_rjPrTpep2_1(.din(w_dff_B_1b4SG3UD4_1),.dout(w_dff_B_rjPrTpep2_1),.clk(gclk));
	jdff dff_B_v8vo6aph6_1(.din(w_dff_B_rjPrTpep2_1),.dout(w_dff_B_v8vo6aph6_1),.clk(gclk));
	jdff dff_B_GPP20TpI9_1(.din(w_dff_B_v8vo6aph6_1),.dout(w_dff_B_GPP20TpI9_1),.clk(gclk));
	jdff dff_B_DxnqTG731_1(.din(w_dff_B_GPP20TpI9_1),.dout(w_dff_B_DxnqTG731_1),.clk(gclk));
	jdff dff_B_f4A6OvnA9_1(.din(w_dff_B_DxnqTG731_1),.dout(w_dff_B_f4A6OvnA9_1),.clk(gclk));
	jdff dff_B_sXFj5RV76_1(.din(w_dff_B_f4A6OvnA9_1),.dout(w_dff_B_sXFj5RV76_1),.clk(gclk));
	jdff dff_B_t6n5teLA0_1(.din(w_dff_B_sXFj5RV76_1),.dout(w_dff_B_t6n5teLA0_1),.clk(gclk));
	jdff dff_B_eGtIiAFY6_1(.din(w_dff_B_t6n5teLA0_1),.dout(w_dff_B_eGtIiAFY6_1),.clk(gclk));
	jdff dff_B_N1GsdJ2a5_1(.din(w_dff_B_eGtIiAFY6_1),.dout(w_dff_B_N1GsdJ2a5_1),.clk(gclk));
	jdff dff_B_pkTK782F8_1(.din(w_dff_B_N1GsdJ2a5_1),.dout(w_dff_B_pkTK782F8_1),.clk(gclk));
	jdff dff_B_HmTlhb8b1_1(.din(w_dff_B_pkTK782F8_1),.dout(w_dff_B_HmTlhb8b1_1),.clk(gclk));
	jdff dff_B_gfNzXfd36_1(.din(w_dff_B_HmTlhb8b1_1),.dout(w_dff_B_gfNzXfd36_1),.clk(gclk));
	jdff dff_B_ykuba2Ed6_1(.din(w_dff_B_gfNzXfd36_1),.dout(w_dff_B_ykuba2Ed6_1),.clk(gclk));
	jdff dff_B_83jJYclD3_1(.din(w_dff_B_ykuba2Ed6_1),.dout(w_dff_B_83jJYclD3_1),.clk(gclk));
	jdff dff_B_R4vn3LvQ9_1(.din(w_dff_B_83jJYclD3_1),.dout(w_dff_B_R4vn3LvQ9_1),.clk(gclk));
	jdff dff_B_KK540xpY0_1(.din(w_dff_B_R4vn3LvQ9_1),.dout(w_dff_B_KK540xpY0_1),.clk(gclk));
	jdff dff_B_IlqIn0Sw2_1(.din(w_dff_B_KK540xpY0_1),.dout(w_dff_B_IlqIn0Sw2_1),.clk(gclk));
	jdff dff_B_q4NvRVS12_1(.din(w_dff_B_IlqIn0Sw2_1),.dout(w_dff_B_q4NvRVS12_1),.clk(gclk));
	jdff dff_B_24Tvryrg2_1(.din(w_dff_B_q4NvRVS12_1),.dout(w_dff_B_24Tvryrg2_1),.clk(gclk));
	jdff dff_B_6VIr25WK5_1(.din(w_dff_B_24Tvryrg2_1),.dout(w_dff_B_6VIr25WK5_1),.clk(gclk));
	jdff dff_B_VbfHAiNn1_1(.din(w_dff_B_6VIr25WK5_1),.dout(w_dff_B_VbfHAiNn1_1),.clk(gclk));
	jdff dff_B_miF1RlLv4_1(.din(w_dff_B_VbfHAiNn1_1),.dout(w_dff_B_miF1RlLv4_1),.clk(gclk));
	jdff dff_B_3nrQhyw92_0(.din(n979),.dout(w_dff_B_3nrQhyw92_0),.clk(gclk));
	jdff dff_B_CbbIn7De4_0(.din(w_dff_B_3nrQhyw92_0),.dout(w_dff_B_CbbIn7De4_0),.clk(gclk));
	jdff dff_B_TNhXpKTA8_0(.din(w_dff_B_CbbIn7De4_0),.dout(w_dff_B_TNhXpKTA8_0),.clk(gclk));
	jdff dff_B_XBKPienL3_0(.din(w_dff_B_TNhXpKTA8_0),.dout(w_dff_B_XBKPienL3_0),.clk(gclk));
	jdff dff_B_J4QZxdaB8_0(.din(w_dff_B_XBKPienL3_0),.dout(w_dff_B_J4QZxdaB8_0),.clk(gclk));
	jdff dff_B_VZKRyolt2_0(.din(w_dff_B_J4QZxdaB8_0),.dout(w_dff_B_VZKRyolt2_0),.clk(gclk));
	jdff dff_B_Gq4cEV8O4_0(.din(w_dff_B_VZKRyolt2_0),.dout(w_dff_B_Gq4cEV8O4_0),.clk(gclk));
	jdff dff_B_z5bhuvm83_0(.din(w_dff_B_Gq4cEV8O4_0),.dout(w_dff_B_z5bhuvm83_0),.clk(gclk));
	jdff dff_B_Cfaw5fL02_0(.din(w_dff_B_z5bhuvm83_0),.dout(w_dff_B_Cfaw5fL02_0),.clk(gclk));
	jdff dff_B_lLSfw8h66_0(.din(w_dff_B_Cfaw5fL02_0),.dout(w_dff_B_lLSfw8h66_0),.clk(gclk));
	jdff dff_B_ZPjS357q8_0(.din(w_dff_B_lLSfw8h66_0),.dout(w_dff_B_ZPjS357q8_0),.clk(gclk));
	jdff dff_B_6cCCoO4T4_0(.din(w_dff_B_ZPjS357q8_0),.dout(w_dff_B_6cCCoO4T4_0),.clk(gclk));
	jdff dff_B_51NaMtTy6_0(.din(w_dff_B_6cCCoO4T4_0),.dout(w_dff_B_51NaMtTy6_0),.clk(gclk));
	jdff dff_B_nBtYDfgE3_0(.din(w_dff_B_51NaMtTy6_0),.dout(w_dff_B_nBtYDfgE3_0),.clk(gclk));
	jdff dff_B_lrnpdaoP4_0(.din(w_dff_B_nBtYDfgE3_0),.dout(w_dff_B_lrnpdaoP4_0),.clk(gclk));
	jdff dff_B_PsZmjjBa3_0(.din(w_dff_B_lrnpdaoP4_0),.dout(w_dff_B_PsZmjjBa3_0),.clk(gclk));
	jdff dff_B_YjOEHnX96_0(.din(w_dff_B_PsZmjjBa3_0),.dout(w_dff_B_YjOEHnX96_0),.clk(gclk));
	jdff dff_B_zjCVIRYL7_0(.din(w_dff_B_YjOEHnX96_0),.dout(w_dff_B_zjCVIRYL7_0),.clk(gclk));
	jdff dff_B_LBY4wlAw6_0(.din(w_dff_B_zjCVIRYL7_0),.dout(w_dff_B_LBY4wlAw6_0),.clk(gclk));
	jdff dff_B_Zh5f54wP8_0(.din(w_dff_B_LBY4wlAw6_0),.dout(w_dff_B_Zh5f54wP8_0),.clk(gclk));
	jdff dff_B_evLOa2o75_0(.din(w_dff_B_Zh5f54wP8_0),.dout(w_dff_B_evLOa2o75_0),.clk(gclk));
	jdff dff_B_UJHFRTpn2_0(.din(w_dff_B_evLOa2o75_0),.dout(w_dff_B_UJHFRTpn2_0),.clk(gclk));
	jdff dff_B_DEjALPo85_0(.din(w_dff_B_UJHFRTpn2_0),.dout(w_dff_B_DEjALPo85_0),.clk(gclk));
	jdff dff_B_P4sEBclQ3_0(.din(w_dff_B_DEjALPo85_0),.dout(w_dff_B_P4sEBclQ3_0),.clk(gclk));
	jdff dff_B_LBIBHDpo6_0(.din(w_dff_B_P4sEBclQ3_0),.dout(w_dff_B_LBIBHDpo6_0),.clk(gclk));
	jdff dff_B_Z8GiTpec7_0(.din(w_dff_B_LBIBHDpo6_0),.dout(w_dff_B_Z8GiTpec7_0),.clk(gclk));
	jdff dff_B_4vyCtkBr9_0(.din(w_dff_B_Z8GiTpec7_0),.dout(w_dff_B_4vyCtkBr9_0),.clk(gclk));
	jdff dff_B_RVhu7ODk2_0(.din(w_dff_B_4vyCtkBr9_0),.dout(w_dff_B_RVhu7ODk2_0),.clk(gclk));
	jdff dff_B_NxIVddl43_0(.din(w_dff_B_RVhu7ODk2_0),.dout(w_dff_B_NxIVddl43_0),.clk(gclk));
	jdff dff_B_7d8uokgC2_0(.din(w_dff_B_NxIVddl43_0),.dout(w_dff_B_7d8uokgC2_0),.clk(gclk));
	jdff dff_B_13CNFcAF2_0(.din(w_dff_B_7d8uokgC2_0),.dout(w_dff_B_13CNFcAF2_0),.clk(gclk));
	jdff dff_B_PK67j5m66_0(.din(w_dff_B_13CNFcAF2_0),.dout(w_dff_B_PK67j5m66_0),.clk(gclk));
	jdff dff_B_vXvQQ8JZ8_0(.din(w_dff_B_PK67j5m66_0),.dout(w_dff_B_vXvQQ8JZ8_0),.clk(gclk));
	jdff dff_B_fEHuOur00_0(.din(w_dff_B_vXvQQ8JZ8_0),.dout(w_dff_B_fEHuOur00_0),.clk(gclk));
	jdff dff_B_pYGG8UsA7_0(.din(w_dff_B_fEHuOur00_0),.dout(w_dff_B_pYGG8UsA7_0),.clk(gclk));
	jdff dff_B_lJW7bXCv6_0(.din(w_dff_B_pYGG8UsA7_0),.dout(w_dff_B_lJW7bXCv6_0),.clk(gclk));
	jdff dff_B_AMZD781e0_0(.din(w_dff_B_lJW7bXCv6_0),.dout(w_dff_B_AMZD781e0_0),.clk(gclk));
	jdff dff_B_AzafLKOk8_0(.din(w_dff_B_AMZD781e0_0),.dout(w_dff_B_AzafLKOk8_0),.clk(gclk));
	jdff dff_B_XiEVUsl41_0(.din(w_dff_B_AzafLKOk8_0),.dout(w_dff_B_XiEVUsl41_0),.clk(gclk));
	jdff dff_B_eKyToK7j1_0(.din(w_dff_B_XiEVUsl41_0),.dout(w_dff_B_eKyToK7j1_0),.clk(gclk));
	jdff dff_B_VgmczsXf0_0(.din(w_dff_B_eKyToK7j1_0),.dout(w_dff_B_VgmczsXf0_0),.clk(gclk));
	jdff dff_B_fgcGeT7F4_0(.din(w_dff_B_VgmczsXf0_0),.dout(w_dff_B_fgcGeT7F4_0),.clk(gclk));
	jdff dff_B_yGCbEa8h2_0(.din(w_dff_B_fgcGeT7F4_0),.dout(w_dff_B_yGCbEa8h2_0),.clk(gclk));
	jdff dff_B_VGknEvuL7_0(.din(w_dff_B_yGCbEa8h2_0),.dout(w_dff_B_VGknEvuL7_0),.clk(gclk));
	jdff dff_B_wHcIpB151_0(.din(w_dff_B_VGknEvuL7_0),.dout(w_dff_B_wHcIpB151_0),.clk(gclk));
	jdff dff_B_BciolMIY8_0(.din(w_dff_B_wHcIpB151_0),.dout(w_dff_B_BciolMIY8_0),.clk(gclk));
	jdff dff_B_MmtSn4mq0_0(.din(w_dff_B_BciolMIY8_0),.dout(w_dff_B_MmtSn4mq0_0),.clk(gclk));
	jdff dff_B_dPdT549G8_0(.din(w_dff_B_MmtSn4mq0_0),.dout(w_dff_B_dPdT549G8_0),.clk(gclk));
	jdff dff_B_GxU8k5yj6_0(.din(w_dff_B_dPdT549G8_0),.dout(w_dff_B_GxU8k5yj6_0),.clk(gclk));
	jdff dff_B_aAA4G1Hu8_0(.din(w_dff_B_GxU8k5yj6_0),.dout(w_dff_B_aAA4G1Hu8_0),.clk(gclk));
	jdff dff_B_z08MuNHr2_0(.din(w_dff_B_aAA4G1Hu8_0),.dout(w_dff_B_z08MuNHr2_0),.clk(gclk));
	jdff dff_B_VrgYqoUE8_0(.din(w_dff_B_z08MuNHr2_0),.dout(w_dff_B_VrgYqoUE8_0),.clk(gclk));
	jdff dff_B_PppM4nIV6_0(.din(w_dff_B_VrgYqoUE8_0),.dout(w_dff_B_PppM4nIV6_0),.clk(gclk));
	jdff dff_B_bWRkCA5q7_0(.din(w_dff_B_PppM4nIV6_0),.dout(w_dff_B_bWRkCA5q7_0),.clk(gclk));
	jdff dff_B_Cdr4sT0g5_0(.din(w_dff_B_bWRkCA5q7_0),.dout(w_dff_B_Cdr4sT0g5_0),.clk(gclk));
	jdff dff_B_Pktez2lp6_0(.din(w_dff_B_Cdr4sT0g5_0),.dout(w_dff_B_Pktez2lp6_0),.clk(gclk));
	jdff dff_B_8blY9eG88_0(.din(w_dff_B_Pktez2lp6_0),.dout(w_dff_B_8blY9eG88_0),.clk(gclk));
	jdff dff_B_eXlQ8K6D0_0(.din(w_dff_B_8blY9eG88_0),.dout(w_dff_B_eXlQ8K6D0_0),.clk(gclk));
	jdff dff_B_NaI5Py8a7_0(.din(w_dff_B_eXlQ8K6D0_0),.dout(w_dff_B_NaI5Py8a7_0),.clk(gclk));
	jdff dff_B_AoIHz6HU1_0(.din(w_dff_B_NaI5Py8a7_0),.dout(w_dff_B_AoIHz6HU1_0),.clk(gclk));
	jdff dff_B_7e28TEzI6_0(.din(w_dff_B_AoIHz6HU1_0),.dout(w_dff_B_7e28TEzI6_0),.clk(gclk));
	jdff dff_B_6pzLgnTy5_0(.din(w_dff_B_7e28TEzI6_0),.dout(w_dff_B_6pzLgnTy5_0),.clk(gclk));
	jdff dff_B_RWrg3STi4_0(.din(w_dff_B_6pzLgnTy5_0),.dout(w_dff_B_RWrg3STi4_0),.clk(gclk));
	jdff dff_B_yFNyU4lr3_0(.din(w_dff_B_RWrg3STi4_0),.dout(w_dff_B_yFNyU4lr3_0),.clk(gclk));
	jdff dff_B_G57TeDAz0_0(.din(w_dff_B_yFNyU4lr3_0),.dout(w_dff_B_G57TeDAz0_0),.clk(gclk));
	jdff dff_B_zmQ0upcc8_0(.din(w_dff_B_G57TeDAz0_0),.dout(w_dff_B_zmQ0upcc8_0),.clk(gclk));
	jdff dff_B_2OW9FTIb4_0(.din(w_dff_B_zmQ0upcc8_0),.dout(w_dff_B_2OW9FTIb4_0),.clk(gclk));
	jdff dff_B_F8qd2xgs0_0(.din(w_dff_B_2OW9FTIb4_0),.dout(w_dff_B_F8qd2xgs0_0),.clk(gclk));
	jdff dff_B_7EkivCwc2_0(.din(w_dff_B_F8qd2xgs0_0),.dout(w_dff_B_7EkivCwc2_0),.clk(gclk));
	jdff dff_B_mI2TrU6G2_0(.din(w_dff_B_7EkivCwc2_0),.dout(w_dff_B_mI2TrU6G2_0),.clk(gclk));
	jdff dff_B_UgSyorgU1_0(.din(w_dff_B_mI2TrU6G2_0),.dout(w_dff_B_UgSyorgU1_0),.clk(gclk));
	jdff dff_B_Ib6ErwfP1_0(.din(w_dff_B_UgSyorgU1_0),.dout(w_dff_B_Ib6ErwfP1_0),.clk(gclk));
	jdff dff_B_t8JDe3iy9_0(.din(w_dff_B_Ib6ErwfP1_0),.dout(w_dff_B_t8JDe3iy9_0),.clk(gclk));
	jdff dff_B_SwrFF9Aw4_0(.din(w_dff_B_t8JDe3iy9_0),.dout(w_dff_B_SwrFF9Aw4_0),.clk(gclk));
	jdff dff_B_Vzfxnqkl2_0(.din(w_dff_B_SwrFF9Aw4_0),.dout(w_dff_B_Vzfxnqkl2_0),.clk(gclk));
	jdff dff_B_MyO7Scdb6_0(.din(w_dff_B_Vzfxnqkl2_0),.dout(w_dff_B_MyO7Scdb6_0),.clk(gclk));
	jdff dff_B_RSFQF9bE8_0(.din(w_dff_B_MyO7Scdb6_0),.dout(w_dff_B_RSFQF9bE8_0),.clk(gclk));
	jdff dff_B_WTJABp3A8_0(.din(w_dff_B_RSFQF9bE8_0),.dout(w_dff_B_WTJABp3A8_0),.clk(gclk));
	jdff dff_B_ZRJ9Tv5i7_0(.din(w_dff_B_WTJABp3A8_0),.dout(w_dff_B_ZRJ9Tv5i7_0),.clk(gclk));
	jdff dff_B_FzWP0Bfa9_0(.din(w_dff_B_ZRJ9Tv5i7_0),.dout(w_dff_B_FzWP0Bfa9_0),.clk(gclk));
	jdff dff_B_xsN5xeiE2_0(.din(w_dff_B_FzWP0Bfa9_0),.dout(w_dff_B_xsN5xeiE2_0),.clk(gclk));
	jdff dff_B_UBkYUe9l1_0(.din(w_dff_B_xsN5xeiE2_0),.dout(w_dff_B_UBkYUe9l1_0),.clk(gclk));
	jdff dff_B_cWja660D3_0(.din(w_dff_B_UBkYUe9l1_0),.dout(w_dff_B_cWja660D3_0),.clk(gclk));
	jdff dff_B_T6L9ubBb7_0(.din(w_dff_B_cWja660D3_0),.dout(w_dff_B_T6L9ubBb7_0),.clk(gclk));
	jdff dff_B_yY9hNZMB2_0(.din(w_dff_B_T6L9ubBb7_0),.dout(w_dff_B_yY9hNZMB2_0),.clk(gclk));
	jdff dff_B_KWycYczW1_0(.din(w_dff_B_yY9hNZMB2_0),.dout(w_dff_B_KWycYczW1_0),.clk(gclk));
	jdff dff_B_IHMLO9jW2_0(.din(w_dff_B_KWycYczW1_0),.dout(w_dff_B_IHMLO9jW2_0),.clk(gclk));
	jdff dff_B_rI0sIsJW4_0(.din(w_dff_B_IHMLO9jW2_0),.dout(w_dff_B_rI0sIsJW4_0),.clk(gclk));
	jdff dff_B_2dm7WGKX0_0(.din(w_dff_B_rI0sIsJW4_0),.dout(w_dff_B_2dm7WGKX0_0),.clk(gclk));
	jdff dff_B_1toynP512_0(.din(w_dff_B_2dm7WGKX0_0),.dout(w_dff_B_1toynP512_0),.clk(gclk));
	jdff dff_B_COeXabQJ7_0(.din(w_dff_B_1toynP512_0),.dout(w_dff_B_COeXabQJ7_0),.clk(gclk));
	jdff dff_B_SfJJgq0q0_0(.din(w_dff_B_COeXabQJ7_0),.dout(w_dff_B_SfJJgq0q0_0),.clk(gclk));
	jdff dff_B_PmwnDScI5_0(.din(w_dff_B_SfJJgq0q0_0),.dout(w_dff_B_PmwnDScI5_0),.clk(gclk));
	jdff dff_B_f6wAjAeX6_0(.din(w_dff_B_PmwnDScI5_0),.dout(w_dff_B_f6wAjAeX6_0),.clk(gclk));
	jdff dff_B_o5qM1l3d5_0(.din(w_dff_B_f6wAjAeX6_0),.dout(w_dff_B_o5qM1l3d5_0),.clk(gclk));
	jdff dff_B_HMy8kcEr3_0(.din(w_dff_B_o5qM1l3d5_0),.dout(w_dff_B_HMy8kcEr3_0),.clk(gclk));
	jdff dff_B_ZXdUhwdU2_0(.din(w_dff_B_HMy8kcEr3_0),.dout(w_dff_B_ZXdUhwdU2_0),.clk(gclk));
	jdff dff_B_qEjfMrsJ3_0(.din(w_dff_B_ZXdUhwdU2_0),.dout(w_dff_B_qEjfMrsJ3_0),.clk(gclk));
	jdff dff_B_wOyfHYTt8_0(.din(w_dff_B_qEjfMrsJ3_0),.dout(w_dff_B_wOyfHYTt8_0),.clk(gclk));
	jdff dff_B_Z5B1ifAp1_1(.din(n972),.dout(w_dff_B_Z5B1ifAp1_1),.clk(gclk));
	jdff dff_B_smI5au8k5_1(.din(w_dff_B_Z5B1ifAp1_1),.dout(w_dff_B_smI5au8k5_1),.clk(gclk));
	jdff dff_B_6BILCbsP8_1(.din(w_dff_B_smI5au8k5_1),.dout(w_dff_B_6BILCbsP8_1),.clk(gclk));
	jdff dff_B_dKxRMyPF3_1(.din(w_dff_B_6BILCbsP8_1),.dout(w_dff_B_dKxRMyPF3_1),.clk(gclk));
	jdff dff_B_Bfm9nvDd8_1(.din(w_dff_B_dKxRMyPF3_1),.dout(w_dff_B_Bfm9nvDd8_1),.clk(gclk));
	jdff dff_B_JFlUgZlJ2_1(.din(w_dff_B_Bfm9nvDd8_1),.dout(w_dff_B_JFlUgZlJ2_1),.clk(gclk));
	jdff dff_B_VGVnmGfa2_1(.din(w_dff_B_JFlUgZlJ2_1),.dout(w_dff_B_VGVnmGfa2_1),.clk(gclk));
	jdff dff_B_mHTX2EBj4_1(.din(w_dff_B_VGVnmGfa2_1),.dout(w_dff_B_mHTX2EBj4_1),.clk(gclk));
	jdff dff_B_2kMjsHUf0_1(.din(w_dff_B_mHTX2EBj4_1),.dout(w_dff_B_2kMjsHUf0_1),.clk(gclk));
	jdff dff_B_klBU5ysp5_1(.din(w_dff_B_2kMjsHUf0_1),.dout(w_dff_B_klBU5ysp5_1),.clk(gclk));
	jdff dff_B_NyVsTaYp6_1(.din(w_dff_B_klBU5ysp5_1),.dout(w_dff_B_NyVsTaYp6_1),.clk(gclk));
	jdff dff_B_UJoFoob13_1(.din(w_dff_B_NyVsTaYp6_1),.dout(w_dff_B_UJoFoob13_1),.clk(gclk));
	jdff dff_B_mA1B7HbN8_1(.din(w_dff_B_UJoFoob13_1),.dout(w_dff_B_mA1B7HbN8_1),.clk(gclk));
	jdff dff_B_Rlwfmm4F2_1(.din(w_dff_B_mA1B7HbN8_1),.dout(w_dff_B_Rlwfmm4F2_1),.clk(gclk));
	jdff dff_B_UIxNoNV49_1(.din(w_dff_B_Rlwfmm4F2_1),.dout(w_dff_B_UIxNoNV49_1),.clk(gclk));
	jdff dff_B_fwXK3dgO4_1(.din(w_dff_B_UIxNoNV49_1),.dout(w_dff_B_fwXK3dgO4_1),.clk(gclk));
	jdff dff_B_X8d1YTXT0_1(.din(w_dff_B_fwXK3dgO4_1),.dout(w_dff_B_X8d1YTXT0_1),.clk(gclk));
	jdff dff_B_y4DbhuP14_1(.din(w_dff_B_X8d1YTXT0_1),.dout(w_dff_B_y4DbhuP14_1),.clk(gclk));
	jdff dff_B_7ZzlPaq74_1(.din(w_dff_B_y4DbhuP14_1),.dout(w_dff_B_7ZzlPaq74_1),.clk(gclk));
	jdff dff_B_JUCpOFes5_1(.din(w_dff_B_7ZzlPaq74_1),.dout(w_dff_B_JUCpOFes5_1),.clk(gclk));
	jdff dff_B_sRnnoN4f1_1(.din(w_dff_B_JUCpOFes5_1),.dout(w_dff_B_sRnnoN4f1_1),.clk(gclk));
	jdff dff_B_UQ6ky9QJ5_1(.din(w_dff_B_sRnnoN4f1_1),.dout(w_dff_B_UQ6ky9QJ5_1),.clk(gclk));
	jdff dff_B_Hc39as0V8_1(.din(w_dff_B_UQ6ky9QJ5_1),.dout(w_dff_B_Hc39as0V8_1),.clk(gclk));
	jdff dff_B_kkQSVCxI2_1(.din(w_dff_B_Hc39as0V8_1),.dout(w_dff_B_kkQSVCxI2_1),.clk(gclk));
	jdff dff_B_tjrJW4Jp7_1(.din(w_dff_B_kkQSVCxI2_1),.dout(w_dff_B_tjrJW4Jp7_1),.clk(gclk));
	jdff dff_B_6iEMUaG30_1(.din(w_dff_B_tjrJW4Jp7_1),.dout(w_dff_B_6iEMUaG30_1),.clk(gclk));
	jdff dff_B_Dicl31VT7_1(.din(w_dff_B_6iEMUaG30_1),.dout(w_dff_B_Dicl31VT7_1),.clk(gclk));
	jdff dff_B_o9uwlSEE9_1(.din(w_dff_B_Dicl31VT7_1),.dout(w_dff_B_o9uwlSEE9_1),.clk(gclk));
	jdff dff_B_fBunnmMH4_1(.din(w_dff_B_o9uwlSEE9_1),.dout(w_dff_B_fBunnmMH4_1),.clk(gclk));
	jdff dff_B_vSdZt5K19_1(.din(w_dff_B_fBunnmMH4_1),.dout(w_dff_B_vSdZt5K19_1),.clk(gclk));
	jdff dff_B_oEcHW4UD8_1(.din(w_dff_B_vSdZt5K19_1),.dout(w_dff_B_oEcHW4UD8_1),.clk(gclk));
	jdff dff_B_hBQGymFB7_1(.din(w_dff_B_oEcHW4UD8_1),.dout(w_dff_B_hBQGymFB7_1),.clk(gclk));
	jdff dff_B_YFRf7nCJ4_1(.din(w_dff_B_hBQGymFB7_1),.dout(w_dff_B_YFRf7nCJ4_1),.clk(gclk));
	jdff dff_B_UjkGPIGk1_1(.din(w_dff_B_YFRf7nCJ4_1),.dout(w_dff_B_UjkGPIGk1_1),.clk(gclk));
	jdff dff_B_0L0OPBlx1_1(.din(w_dff_B_UjkGPIGk1_1),.dout(w_dff_B_0L0OPBlx1_1),.clk(gclk));
	jdff dff_B_dDq2mjJ57_1(.din(w_dff_B_0L0OPBlx1_1),.dout(w_dff_B_dDq2mjJ57_1),.clk(gclk));
	jdff dff_B_a33gikOx4_1(.din(w_dff_B_dDq2mjJ57_1),.dout(w_dff_B_a33gikOx4_1),.clk(gclk));
	jdff dff_B_cfv2yNw21_1(.din(w_dff_B_a33gikOx4_1),.dout(w_dff_B_cfv2yNw21_1),.clk(gclk));
	jdff dff_B_mbMDqcV79_1(.din(w_dff_B_cfv2yNw21_1),.dout(w_dff_B_mbMDqcV79_1),.clk(gclk));
	jdff dff_B_rsbBSUQk8_1(.din(w_dff_B_mbMDqcV79_1),.dout(w_dff_B_rsbBSUQk8_1),.clk(gclk));
	jdff dff_B_ArvOWERt6_1(.din(w_dff_B_rsbBSUQk8_1),.dout(w_dff_B_ArvOWERt6_1),.clk(gclk));
	jdff dff_B_GKY25DZB1_1(.din(w_dff_B_ArvOWERt6_1),.dout(w_dff_B_GKY25DZB1_1),.clk(gclk));
	jdff dff_B_P2HXyoyy1_1(.din(w_dff_B_GKY25DZB1_1),.dout(w_dff_B_P2HXyoyy1_1),.clk(gclk));
	jdff dff_B_rFmaUZyg2_1(.din(w_dff_B_P2HXyoyy1_1),.dout(w_dff_B_rFmaUZyg2_1),.clk(gclk));
	jdff dff_B_OfaP09Nb3_1(.din(w_dff_B_rFmaUZyg2_1),.dout(w_dff_B_OfaP09Nb3_1),.clk(gclk));
	jdff dff_B_5EIl57YG4_1(.din(w_dff_B_OfaP09Nb3_1),.dout(w_dff_B_5EIl57YG4_1),.clk(gclk));
	jdff dff_B_lW5Lng6G3_1(.din(w_dff_B_5EIl57YG4_1),.dout(w_dff_B_lW5Lng6G3_1),.clk(gclk));
	jdff dff_B_nJrWBbhn9_1(.din(w_dff_B_lW5Lng6G3_1),.dout(w_dff_B_nJrWBbhn9_1),.clk(gclk));
	jdff dff_B_OlKgHFTO7_1(.din(w_dff_B_nJrWBbhn9_1),.dout(w_dff_B_OlKgHFTO7_1),.clk(gclk));
	jdff dff_B_LHGOzpwD8_1(.din(w_dff_B_OlKgHFTO7_1),.dout(w_dff_B_LHGOzpwD8_1),.clk(gclk));
	jdff dff_B_6r7IHxOB7_1(.din(w_dff_B_LHGOzpwD8_1),.dout(w_dff_B_6r7IHxOB7_1),.clk(gclk));
	jdff dff_B_vyPhRNvO9_1(.din(w_dff_B_6r7IHxOB7_1),.dout(w_dff_B_vyPhRNvO9_1),.clk(gclk));
	jdff dff_B_nNk2b9Pr5_1(.din(w_dff_B_vyPhRNvO9_1),.dout(w_dff_B_nNk2b9Pr5_1),.clk(gclk));
	jdff dff_B_eZ1gYnSV0_1(.din(w_dff_B_nNk2b9Pr5_1),.dout(w_dff_B_eZ1gYnSV0_1),.clk(gclk));
	jdff dff_B_UcLdKzOT7_1(.din(w_dff_B_eZ1gYnSV0_1),.dout(w_dff_B_UcLdKzOT7_1),.clk(gclk));
	jdff dff_B_PfQFCLM56_1(.din(w_dff_B_UcLdKzOT7_1),.dout(w_dff_B_PfQFCLM56_1),.clk(gclk));
	jdff dff_B_3X21uRNw3_1(.din(w_dff_B_PfQFCLM56_1),.dout(w_dff_B_3X21uRNw3_1),.clk(gclk));
	jdff dff_B_i7oZEuPT7_1(.din(w_dff_B_3X21uRNw3_1),.dout(w_dff_B_i7oZEuPT7_1),.clk(gclk));
	jdff dff_B_jnun1KzD2_1(.din(w_dff_B_i7oZEuPT7_1),.dout(w_dff_B_jnun1KzD2_1),.clk(gclk));
	jdff dff_B_QDCFAuB92_1(.din(w_dff_B_jnun1KzD2_1),.dout(w_dff_B_QDCFAuB92_1),.clk(gclk));
	jdff dff_B_R5voHkfq6_1(.din(w_dff_B_QDCFAuB92_1),.dout(w_dff_B_R5voHkfq6_1),.clk(gclk));
	jdff dff_B_7dJi9ygn3_1(.din(w_dff_B_R5voHkfq6_1),.dout(w_dff_B_7dJi9ygn3_1),.clk(gclk));
	jdff dff_B_XV6BtSFk7_1(.din(w_dff_B_7dJi9ygn3_1),.dout(w_dff_B_XV6BtSFk7_1),.clk(gclk));
	jdff dff_B_tCpZB0Im2_1(.din(w_dff_B_XV6BtSFk7_1),.dout(w_dff_B_tCpZB0Im2_1),.clk(gclk));
	jdff dff_B_iVbImZAW4_1(.din(w_dff_B_tCpZB0Im2_1),.dout(w_dff_B_iVbImZAW4_1),.clk(gclk));
	jdff dff_B_MyOzqX2M7_1(.din(w_dff_B_iVbImZAW4_1),.dout(w_dff_B_MyOzqX2M7_1),.clk(gclk));
	jdff dff_B_hv7jnx4o7_1(.din(w_dff_B_MyOzqX2M7_1),.dout(w_dff_B_hv7jnx4o7_1),.clk(gclk));
	jdff dff_B_btcU6MIV7_1(.din(w_dff_B_hv7jnx4o7_1),.dout(w_dff_B_btcU6MIV7_1),.clk(gclk));
	jdff dff_B_d6zJbC1Z1_1(.din(w_dff_B_btcU6MIV7_1),.dout(w_dff_B_d6zJbC1Z1_1),.clk(gclk));
	jdff dff_B_P7aMs2qJ9_1(.din(w_dff_B_d6zJbC1Z1_1),.dout(w_dff_B_P7aMs2qJ9_1),.clk(gclk));
	jdff dff_B_Bd1rbLsN2_1(.din(w_dff_B_P7aMs2qJ9_1),.dout(w_dff_B_Bd1rbLsN2_1),.clk(gclk));
	jdff dff_B_0vveAfYR4_1(.din(w_dff_B_Bd1rbLsN2_1),.dout(w_dff_B_0vveAfYR4_1),.clk(gclk));
	jdff dff_B_wQrgJvMG9_1(.din(w_dff_B_0vveAfYR4_1),.dout(w_dff_B_wQrgJvMG9_1),.clk(gclk));
	jdff dff_B_jMEt6kbz1_1(.din(w_dff_B_wQrgJvMG9_1),.dout(w_dff_B_jMEt6kbz1_1),.clk(gclk));
	jdff dff_B_7DcZmRHA5_1(.din(w_dff_B_jMEt6kbz1_1),.dout(w_dff_B_7DcZmRHA5_1),.clk(gclk));
	jdff dff_B_FyB1FXnj4_1(.din(w_dff_B_7DcZmRHA5_1),.dout(w_dff_B_FyB1FXnj4_1),.clk(gclk));
	jdff dff_B_TxpvTaAI6_1(.din(w_dff_B_FyB1FXnj4_1),.dout(w_dff_B_TxpvTaAI6_1),.clk(gclk));
	jdff dff_B_EtMdV7Et3_1(.din(w_dff_B_TxpvTaAI6_1),.dout(w_dff_B_EtMdV7Et3_1),.clk(gclk));
	jdff dff_B_ddOF38Ih3_1(.din(w_dff_B_EtMdV7Et3_1),.dout(w_dff_B_ddOF38Ih3_1),.clk(gclk));
	jdff dff_B_yGYLIp2W9_1(.din(w_dff_B_ddOF38Ih3_1),.dout(w_dff_B_yGYLIp2W9_1),.clk(gclk));
	jdff dff_B_TjlEfZXk4_1(.din(w_dff_B_yGYLIp2W9_1),.dout(w_dff_B_TjlEfZXk4_1),.clk(gclk));
	jdff dff_B_l8Ja5oxY8_1(.din(w_dff_B_TjlEfZXk4_1),.dout(w_dff_B_l8Ja5oxY8_1),.clk(gclk));
	jdff dff_B_U2AwKyTz1_1(.din(w_dff_B_l8Ja5oxY8_1),.dout(w_dff_B_U2AwKyTz1_1),.clk(gclk));
	jdff dff_B_ApzrNSSa7_1(.din(w_dff_B_U2AwKyTz1_1),.dout(w_dff_B_ApzrNSSa7_1),.clk(gclk));
	jdff dff_B_kMolEM8f1_1(.din(w_dff_B_ApzrNSSa7_1),.dout(w_dff_B_kMolEM8f1_1),.clk(gclk));
	jdff dff_B_RiZp2iRJ1_1(.din(w_dff_B_kMolEM8f1_1),.dout(w_dff_B_RiZp2iRJ1_1),.clk(gclk));
	jdff dff_B_CqAEFC1Z7_1(.din(w_dff_B_RiZp2iRJ1_1),.dout(w_dff_B_CqAEFC1Z7_1),.clk(gclk));
	jdff dff_B_pYDoLRgG2_1(.din(w_dff_B_CqAEFC1Z7_1),.dout(w_dff_B_pYDoLRgG2_1),.clk(gclk));
	jdff dff_B_YezcYCFo5_1(.din(w_dff_B_pYDoLRgG2_1),.dout(w_dff_B_YezcYCFo5_1),.clk(gclk));
	jdff dff_B_fOm82p1F7_1(.din(w_dff_B_YezcYCFo5_1),.dout(w_dff_B_fOm82p1F7_1),.clk(gclk));
	jdff dff_B_Wse4aiTd1_1(.din(w_dff_B_fOm82p1F7_1),.dout(w_dff_B_Wse4aiTd1_1),.clk(gclk));
	jdff dff_B_yqELsMRu5_1(.din(w_dff_B_Wse4aiTd1_1),.dout(w_dff_B_yqELsMRu5_1),.clk(gclk));
	jdff dff_B_thnOzZPD3_1(.din(w_dff_B_yqELsMRu5_1),.dout(w_dff_B_thnOzZPD3_1),.clk(gclk));
	jdff dff_B_0hf5fLIH0_1(.din(w_dff_B_thnOzZPD3_1),.dout(w_dff_B_0hf5fLIH0_1),.clk(gclk));
	jdff dff_B_grgCfZ3C4_1(.din(w_dff_B_0hf5fLIH0_1),.dout(w_dff_B_grgCfZ3C4_1),.clk(gclk));
	jdff dff_B_TUo8Ckd70_1(.din(w_dff_B_grgCfZ3C4_1),.dout(w_dff_B_TUo8Ckd70_1),.clk(gclk));
	jdff dff_B_8mMDisi62_1(.din(w_dff_B_TUo8Ckd70_1),.dout(w_dff_B_8mMDisi62_1),.clk(gclk));
	jdff dff_B_sukvz7S18_1(.din(w_dff_B_8mMDisi62_1),.dout(w_dff_B_sukvz7S18_1),.clk(gclk));
	jdff dff_B_rUqvxiH18_0(.din(n973),.dout(w_dff_B_rUqvxiH18_0),.clk(gclk));
	jdff dff_B_Xldh1oT70_0(.din(w_dff_B_rUqvxiH18_0),.dout(w_dff_B_Xldh1oT70_0),.clk(gclk));
	jdff dff_B_o2HIcIT42_0(.din(w_dff_B_Xldh1oT70_0),.dout(w_dff_B_o2HIcIT42_0),.clk(gclk));
	jdff dff_B_6wcPQrus1_0(.din(w_dff_B_o2HIcIT42_0),.dout(w_dff_B_6wcPQrus1_0),.clk(gclk));
	jdff dff_B_VeBO6M3b3_0(.din(w_dff_B_6wcPQrus1_0),.dout(w_dff_B_VeBO6M3b3_0),.clk(gclk));
	jdff dff_B_H9JAqf418_0(.din(w_dff_B_VeBO6M3b3_0),.dout(w_dff_B_H9JAqf418_0),.clk(gclk));
	jdff dff_B_Xac74v3o8_0(.din(w_dff_B_H9JAqf418_0),.dout(w_dff_B_Xac74v3o8_0),.clk(gclk));
	jdff dff_B_i61dsSQq3_0(.din(w_dff_B_Xac74v3o8_0),.dout(w_dff_B_i61dsSQq3_0),.clk(gclk));
	jdff dff_B_5g92NNFy2_0(.din(w_dff_B_i61dsSQq3_0),.dout(w_dff_B_5g92NNFy2_0),.clk(gclk));
	jdff dff_B_HtbQ3uBa8_0(.din(w_dff_B_5g92NNFy2_0),.dout(w_dff_B_HtbQ3uBa8_0),.clk(gclk));
	jdff dff_B_P8OExxy25_0(.din(w_dff_B_HtbQ3uBa8_0),.dout(w_dff_B_P8OExxy25_0),.clk(gclk));
	jdff dff_B_fHPKsPlV9_0(.din(w_dff_B_P8OExxy25_0),.dout(w_dff_B_fHPKsPlV9_0),.clk(gclk));
	jdff dff_B_WeKWfWe80_0(.din(w_dff_B_fHPKsPlV9_0),.dout(w_dff_B_WeKWfWe80_0),.clk(gclk));
	jdff dff_B_LW4ghJrl4_0(.din(w_dff_B_WeKWfWe80_0),.dout(w_dff_B_LW4ghJrl4_0),.clk(gclk));
	jdff dff_B_LhLFQMKr0_0(.din(w_dff_B_LW4ghJrl4_0),.dout(w_dff_B_LhLFQMKr0_0),.clk(gclk));
	jdff dff_B_SJQK9jwT8_0(.din(w_dff_B_LhLFQMKr0_0),.dout(w_dff_B_SJQK9jwT8_0),.clk(gclk));
	jdff dff_B_M158QfaG4_0(.din(w_dff_B_SJQK9jwT8_0),.dout(w_dff_B_M158QfaG4_0),.clk(gclk));
	jdff dff_B_pcL1Gjfy1_0(.din(w_dff_B_M158QfaG4_0),.dout(w_dff_B_pcL1Gjfy1_0),.clk(gclk));
	jdff dff_B_kI75E0aa1_0(.din(w_dff_B_pcL1Gjfy1_0),.dout(w_dff_B_kI75E0aa1_0),.clk(gclk));
	jdff dff_B_LpKS0x3B7_0(.din(w_dff_B_kI75E0aa1_0),.dout(w_dff_B_LpKS0x3B7_0),.clk(gclk));
	jdff dff_B_uPgbB2Bz0_0(.din(w_dff_B_LpKS0x3B7_0),.dout(w_dff_B_uPgbB2Bz0_0),.clk(gclk));
	jdff dff_B_Fo9bFWL57_0(.din(w_dff_B_uPgbB2Bz0_0),.dout(w_dff_B_Fo9bFWL57_0),.clk(gclk));
	jdff dff_B_tvfTDtLb4_0(.din(w_dff_B_Fo9bFWL57_0),.dout(w_dff_B_tvfTDtLb4_0),.clk(gclk));
	jdff dff_B_nnFWtXnt4_0(.din(w_dff_B_tvfTDtLb4_0),.dout(w_dff_B_nnFWtXnt4_0),.clk(gclk));
	jdff dff_B_HMgYkUtU6_0(.din(w_dff_B_nnFWtXnt4_0),.dout(w_dff_B_HMgYkUtU6_0),.clk(gclk));
	jdff dff_B_y9doERtt2_0(.din(w_dff_B_HMgYkUtU6_0),.dout(w_dff_B_y9doERtt2_0),.clk(gclk));
	jdff dff_B_FAGuU0yQ9_0(.din(w_dff_B_y9doERtt2_0),.dout(w_dff_B_FAGuU0yQ9_0),.clk(gclk));
	jdff dff_B_H5aKfxvI6_0(.din(w_dff_B_FAGuU0yQ9_0),.dout(w_dff_B_H5aKfxvI6_0),.clk(gclk));
	jdff dff_B_Fvu5ov6C6_0(.din(w_dff_B_H5aKfxvI6_0),.dout(w_dff_B_Fvu5ov6C6_0),.clk(gclk));
	jdff dff_B_UcH42UBV5_0(.din(w_dff_B_Fvu5ov6C6_0),.dout(w_dff_B_UcH42UBV5_0),.clk(gclk));
	jdff dff_B_LB0ACfsO5_0(.din(w_dff_B_UcH42UBV5_0),.dout(w_dff_B_LB0ACfsO5_0),.clk(gclk));
	jdff dff_B_VzTEqsHa6_0(.din(w_dff_B_LB0ACfsO5_0),.dout(w_dff_B_VzTEqsHa6_0),.clk(gclk));
	jdff dff_B_Zg4NCMYi9_0(.din(w_dff_B_VzTEqsHa6_0),.dout(w_dff_B_Zg4NCMYi9_0),.clk(gclk));
	jdff dff_B_AnzSAkka4_0(.din(w_dff_B_Zg4NCMYi9_0),.dout(w_dff_B_AnzSAkka4_0),.clk(gclk));
	jdff dff_B_7GdqVjWD1_0(.din(w_dff_B_AnzSAkka4_0),.dout(w_dff_B_7GdqVjWD1_0),.clk(gclk));
	jdff dff_B_sPuPpmIu0_0(.din(w_dff_B_7GdqVjWD1_0),.dout(w_dff_B_sPuPpmIu0_0),.clk(gclk));
	jdff dff_B_pXV3OwQB5_0(.din(w_dff_B_sPuPpmIu0_0),.dout(w_dff_B_pXV3OwQB5_0),.clk(gclk));
	jdff dff_B_GGwFsP557_0(.din(w_dff_B_pXV3OwQB5_0),.dout(w_dff_B_GGwFsP557_0),.clk(gclk));
	jdff dff_B_CBJ2Dphc7_0(.din(w_dff_B_GGwFsP557_0),.dout(w_dff_B_CBJ2Dphc7_0),.clk(gclk));
	jdff dff_B_8pPbuVo30_0(.din(w_dff_B_CBJ2Dphc7_0),.dout(w_dff_B_8pPbuVo30_0),.clk(gclk));
	jdff dff_B_qNXc3wRs9_0(.din(w_dff_B_8pPbuVo30_0),.dout(w_dff_B_qNXc3wRs9_0),.clk(gclk));
	jdff dff_B_lvk3HfUk8_0(.din(w_dff_B_qNXc3wRs9_0),.dout(w_dff_B_lvk3HfUk8_0),.clk(gclk));
	jdff dff_B_uq5ctBI36_0(.din(w_dff_B_lvk3HfUk8_0),.dout(w_dff_B_uq5ctBI36_0),.clk(gclk));
	jdff dff_B_1Zi5DzAv1_0(.din(w_dff_B_uq5ctBI36_0),.dout(w_dff_B_1Zi5DzAv1_0),.clk(gclk));
	jdff dff_B_Qd6rnflo3_0(.din(w_dff_B_1Zi5DzAv1_0),.dout(w_dff_B_Qd6rnflo3_0),.clk(gclk));
	jdff dff_B_itOgf6c80_0(.din(w_dff_B_Qd6rnflo3_0),.dout(w_dff_B_itOgf6c80_0),.clk(gclk));
	jdff dff_B_l33AUiP30_0(.din(w_dff_B_itOgf6c80_0),.dout(w_dff_B_l33AUiP30_0),.clk(gclk));
	jdff dff_B_FGTJPmTo6_0(.din(w_dff_B_l33AUiP30_0),.dout(w_dff_B_FGTJPmTo6_0),.clk(gclk));
	jdff dff_B_pTSbL3mH8_0(.din(w_dff_B_FGTJPmTo6_0),.dout(w_dff_B_pTSbL3mH8_0),.clk(gclk));
	jdff dff_B_CCqJujbK5_0(.din(w_dff_B_pTSbL3mH8_0),.dout(w_dff_B_CCqJujbK5_0),.clk(gclk));
	jdff dff_B_l6N3iB2r2_0(.din(w_dff_B_CCqJujbK5_0),.dout(w_dff_B_l6N3iB2r2_0),.clk(gclk));
	jdff dff_B_AKznrzuT1_0(.din(w_dff_B_l6N3iB2r2_0),.dout(w_dff_B_AKznrzuT1_0),.clk(gclk));
	jdff dff_B_FhE4lZ2I0_0(.din(w_dff_B_AKznrzuT1_0),.dout(w_dff_B_FhE4lZ2I0_0),.clk(gclk));
	jdff dff_B_spDVAovP0_0(.din(w_dff_B_FhE4lZ2I0_0),.dout(w_dff_B_spDVAovP0_0),.clk(gclk));
	jdff dff_B_AUuyQZPs7_0(.din(w_dff_B_spDVAovP0_0),.dout(w_dff_B_AUuyQZPs7_0),.clk(gclk));
	jdff dff_B_BjrK1yoO2_0(.din(w_dff_B_AUuyQZPs7_0),.dout(w_dff_B_BjrK1yoO2_0),.clk(gclk));
	jdff dff_B_oJApgSLa1_0(.din(w_dff_B_BjrK1yoO2_0),.dout(w_dff_B_oJApgSLa1_0),.clk(gclk));
	jdff dff_B_wYkdhPUN9_0(.din(w_dff_B_oJApgSLa1_0),.dout(w_dff_B_wYkdhPUN9_0),.clk(gclk));
	jdff dff_B_HUBeeWJM7_0(.din(w_dff_B_wYkdhPUN9_0),.dout(w_dff_B_HUBeeWJM7_0),.clk(gclk));
	jdff dff_B_M9d0kA6r8_0(.din(w_dff_B_HUBeeWJM7_0),.dout(w_dff_B_M9d0kA6r8_0),.clk(gclk));
	jdff dff_B_IKCL7hOb2_0(.din(w_dff_B_M9d0kA6r8_0),.dout(w_dff_B_IKCL7hOb2_0),.clk(gclk));
	jdff dff_B_yCSblpJ54_0(.din(w_dff_B_IKCL7hOb2_0),.dout(w_dff_B_yCSblpJ54_0),.clk(gclk));
	jdff dff_B_KiYAU9YB4_0(.din(w_dff_B_yCSblpJ54_0),.dout(w_dff_B_KiYAU9YB4_0),.clk(gclk));
	jdff dff_B_DtAXHXqJ7_0(.din(w_dff_B_KiYAU9YB4_0),.dout(w_dff_B_DtAXHXqJ7_0),.clk(gclk));
	jdff dff_B_WeGVkTtR1_0(.din(w_dff_B_DtAXHXqJ7_0),.dout(w_dff_B_WeGVkTtR1_0),.clk(gclk));
	jdff dff_B_GR4eUGU35_0(.din(w_dff_B_WeGVkTtR1_0),.dout(w_dff_B_GR4eUGU35_0),.clk(gclk));
	jdff dff_B_9jjULUl33_0(.din(w_dff_B_GR4eUGU35_0),.dout(w_dff_B_9jjULUl33_0),.clk(gclk));
	jdff dff_B_LL6Z1eYE5_0(.din(w_dff_B_9jjULUl33_0),.dout(w_dff_B_LL6Z1eYE5_0),.clk(gclk));
	jdff dff_B_pRfGqLQ09_0(.din(w_dff_B_LL6Z1eYE5_0),.dout(w_dff_B_pRfGqLQ09_0),.clk(gclk));
	jdff dff_B_n1N6rYyn8_0(.din(w_dff_B_pRfGqLQ09_0),.dout(w_dff_B_n1N6rYyn8_0),.clk(gclk));
	jdff dff_B_VtPbto6B5_0(.din(w_dff_B_n1N6rYyn8_0),.dout(w_dff_B_VtPbto6B5_0),.clk(gclk));
	jdff dff_B_Kd1WDuCv8_0(.din(w_dff_B_VtPbto6B5_0),.dout(w_dff_B_Kd1WDuCv8_0),.clk(gclk));
	jdff dff_B_hWNAZ5To5_0(.din(w_dff_B_Kd1WDuCv8_0),.dout(w_dff_B_hWNAZ5To5_0),.clk(gclk));
	jdff dff_B_kq8Swrjc6_0(.din(w_dff_B_hWNAZ5To5_0),.dout(w_dff_B_kq8Swrjc6_0),.clk(gclk));
	jdff dff_B_ezraewP35_0(.din(w_dff_B_kq8Swrjc6_0),.dout(w_dff_B_ezraewP35_0),.clk(gclk));
	jdff dff_B_wOHk7AAH8_0(.din(w_dff_B_ezraewP35_0),.dout(w_dff_B_wOHk7AAH8_0),.clk(gclk));
	jdff dff_B_U8kJ5bLc9_0(.din(w_dff_B_wOHk7AAH8_0),.dout(w_dff_B_U8kJ5bLc9_0),.clk(gclk));
	jdff dff_B_kxCeRf143_0(.din(w_dff_B_U8kJ5bLc9_0),.dout(w_dff_B_kxCeRf143_0),.clk(gclk));
	jdff dff_B_0cRfT15D3_0(.din(w_dff_B_kxCeRf143_0),.dout(w_dff_B_0cRfT15D3_0),.clk(gclk));
	jdff dff_B_sBhSsg0t4_0(.din(w_dff_B_0cRfT15D3_0),.dout(w_dff_B_sBhSsg0t4_0),.clk(gclk));
	jdff dff_B_1Fyhinto4_0(.din(w_dff_B_sBhSsg0t4_0),.dout(w_dff_B_1Fyhinto4_0),.clk(gclk));
	jdff dff_B_O72zvYXv9_0(.din(w_dff_B_1Fyhinto4_0),.dout(w_dff_B_O72zvYXv9_0),.clk(gclk));
	jdff dff_B_nbRar6NA3_0(.din(w_dff_B_O72zvYXv9_0),.dout(w_dff_B_nbRar6NA3_0),.clk(gclk));
	jdff dff_B_F1EQOuCM8_0(.din(w_dff_B_nbRar6NA3_0),.dout(w_dff_B_F1EQOuCM8_0),.clk(gclk));
	jdff dff_B_oLhzaB2K7_0(.din(w_dff_B_F1EQOuCM8_0),.dout(w_dff_B_oLhzaB2K7_0),.clk(gclk));
	jdff dff_B_UzQxTQzl6_0(.din(w_dff_B_oLhzaB2K7_0),.dout(w_dff_B_UzQxTQzl6_0),.clk(gclk));
	jdff dff_B_Q4uhzlvz5_0(.din(w_dff_B_UzQxTQzl6_0),.dout(w_dff_B_Q4uhzlvz5_0),.clk(gclk));
	jdff dff_B_4ghgTtho9_0(.din(w_dff_B_Q4uhzlvz5_0),.dout(w_dff_B_4ghgTtho9_0),.clk(gclk));
	jdff dff_B_bPed92S03_0(.din(w_dff_B_4ghgTtho9_0),.dout(w_dff_B_bPed92S03_0),.clk(gclk));
	jdff dff_B_QEs5bxR17_0(.din(w_dff_B_bPed92S03_0),.dout(w_dff_B_QEs5bxR17_0),.clk(gclk));
	jdff dff_B_ClyVqHKy8_0(.din(w_dff_B_QEs5bxR17_0),.dout(w_dff_B_ClyVqHKy8_0),.clk(gclk));
	jdff dff_B_UkR6PPJC2_0(.din(w_dff_B_ClyVqHKy8_0),.dout(w_dff_B_UkR6PPJC2_0),.clk(gclk));
	jdff dff_B_AWx6xZS86_0(.din(w_dff_B_UkR6PPJC2_0),.dout(w_dff_B_AWx6xZS86_0),.clk(gclk));
	jdff dff_B_ekSGesoT8_0(.din(w_dff_B_AWx6xZS86_0),.dout(w_dff_B_ekSGesoT8_0),.clk(gclk));
	jdff dff_B_p6MYarz92_0(.din(w_dff_B_ekSGesoT8_0),.dout(w_dff_B_p6MYarz92_0),.clk(gclk));
	jdff dff_B_lsj58b6A4_0(.din(w_dff_B_p6MYarz92_0),.dout(w_dff_B_lsj58b6A4_0),.clk(gclk));
	jdff dff_B_MJq8zZki6_0(.din(w_dff_B_lsj58b6A4_0),.dout(w_dff_B_MJq8zZki6_0),.clk(gclk));
	jdff dff_B_CzElqIeo4_0(.din(w_dff_B_MJq8zZki6_0),.dout(w_dff_B_CzElqIeo4_0),.clk(gclk));
	jdff dff_B_Dbr4hHKB7_1(.din(n966),.dout(w_dff_B_Dbr4hHKB7_1),.clk(gclk));
	jdff dff_B_M1V8pSCe2_1(.din(w_dff_B_Dbr4hHKB7_1),.dout(w_dff_B_M1V8pSCe2_1),.clk(gclk));
	jdff dff_B_jt412CnA5_1(.din(w_dff_B_M1V8pSCe2_1),.dout(w_dff_B_jt412CnA5_1),.clk(gclk));
	jdff dff_B_tYMQQef54_1(.din(w_dff_B_jt412CnA5_1),.dout(w_dff_B_tYMQQef54_1),.clk(gclk));
	jdff dff_B_oTXRj5Ij4_1(.din(w_dff_B_tYMQQef54_1),.dout(w_dff_B_oTXRj5Ij4_1),.clk(gclk));
	jdff dff_B_J52uqJQr5_1(.din(w_dff_B_oTXRj5Ij4_1),.dout(w_dff_B_J52uqJQr5_1),.clk(gclk));
	jdff dff_B_AdCRbKfF8_1(.din(w_dff_B_J52uqJQr5_1),.dout(w_dff_B_AdCRbKfF8_1),.clk(gclk));
	jdff dff_B_Fh2SNVTx3_1(.din(w_dff_B_AdCRbKfF8_1),.dout(w_dff_B_Fh2SNVTx3_1),.clk(gclk));
	jdff dff_B_AfDDOqbi3_1(.din(w_dff_B_Fh2SNVTx3_1),.dout(w_dff_B_AfDDOqbi3_1),.clk(gclk));
	jdff dff_B_KumwjENN5_1(.din(w_dff_B_AfDDOqbi3_1),.dout(w_dff_B_KumwjENN5_1),.clk(gclk));
	jdff dff_B_ullppxKj1_1(.din(w_dff_B_KumwjENN5_1),.dout(w_dff_B_ullppxKj1_1),.clk(gclk));
	jdff dff_B_AXN01XtF4_1(.din(w_dff_B_ullppxKj1_1),.dout(w_dff_B_AXN01XtF4_1),.clk(gclk));
	jdff dff_B_NX2ttHWO1_1(.din(w_dff_B_AXN01XtF4_1),.dout(w_dff_B_NX2ttHWO1_1),.clk(gclk));
	jdff dff_B_06IpgZUI4_1(.din(w_dff_B_NX2ttHWO1_1),.dout(w_dff_B_06IpgZUI4_1),.clk(gclk));
	jdff dff_B_zQ5EMnhY8_1(.din(w_dff_B_06IpgZUI4_1),.dout(w_dff_B_zQ5EMnhY8_1),.clk(gclk));
	jdff dff_B_iQFTAae45_1(.din(w_dff_B_zQ5EMnhY8_1),.dout(w_dff_B_iQFTAae45_1),.clk(gclk));
	jdff dff_B_XUbB55pQ4_1(.din(w_dff_B_iQFTAae45_1),.dout(w_dff_B_XUbB55pQ4_1),.clk(gclk));
	jdff dff_B_fejEvfLA7_1(.din(w_dff_B_XUbB55pQ4_1),.dout(w_dff_B_fejEvfLA7_1),.clk(gclk));
	jdff dff_B_HxlJQza61_1(.din(w_dff_B_fejEvfLA7_1),.dout(w_dff_B_HxlJQza61_1),.clk(gclk));
	jdff dff_B_I30PErWL7_1(.din(w_dff_B_HxlJQza61_1),.dout(w_dff_B_I30PErWL7_1),.clk(gclk));
	jdff dff_B_s2I7wNWS1_1(.din(w_dff_B_I30PErWL7_1),.dout(w_dff_B_s2I7wNWS1_1),.clk(gclk));
	jdff dff_B_2GqcAZlD1_1(.din(w_dff_B_s2I7wNWS1_1),.dout(w_dff_B_2GqcAZlD1_1),.clk(gclk));
	jdff dff_B_PPIq027W4_1(.din(w_dff_B_2GqcAZlD1_1),.dout(w_dff_B_PPIq027W4_1),.clk(gclk));
	jdff dff_B_yHUIvbsh8_1(.din(w_dff_B_PPIq027W4_1),.dout(w_dff_B_yHUIvbsh8_1),.clk(gclk));
	jdff dff_B_HHagNUqw6_1(.din(w_dff_B_yHUIvbsh8_1),.dout(w_dff_B_HHagNUqw6_1),.clk(gclk));
	jdff dff_B_E88OA8zG6_1(.din(w_dff_B_HHagNUqw6_1),.dout(w_dff_B_E88OA8zG6_1),.clk(gclk));
	jdff dff_B_0MySkf4y8_1(.din(w_dff_B_E88OA8zG6_1),.dout(w_dff_B_0MySkf4y8_1),.clk(gclk));
	jdff dff_B_4DcEFcyJ8_1(.din(w_dff_B_0MySkf4y8_1),.dout(w_dff_B_4DcEFcyJ8_1),.clk(gclk));
	jdff dff_B_3nZ7x0qX0_1(.din(w_dff_B_4DcEFcyJ8_1),.dout(w_dff_B_3nZ7x0qX0_1),.clk(gclk));
	jdff dff_B_RGNbmbDh7_1(.din(w_dff_B_3nZ7x0qX0_1),.dout(w_dff_B_RGNbmbDh7_1),.clk(gclk));
	jdff dff_B_ead1Dbqk2_1(.din(w_dff_B_RGNbmbDh7_1),.dout(w_dff_B_ead1Dbqk2_1),.clk(gclk));
	jdff dff_B_dtfXQUXA3_1(.din(w_dff_B_ead1Dbqk2_1),.dout(w_dff_B_dtfXQUXA3_1),.clk(gclk));
	jdff dff_B_YcKNjoIO3_1(.din(w_dff_B_dtfXQUXA3_1),.dout(w_dff_B_YcKNjoIO3_1),.clk(gclk));
	jdff dff_B_k6ckExfr4_1(.din(w_dff_B_YcKNjoIO3_1),.dout(w_dff_B_k6ckExfr4_1),.clk(gclk));
	jdff dff_B_b02joubA6_1(.din(w_dff_B_k6ckExfr4_1),.dout(w_dff_B_b02joubA6_1),.clk(gclk));
	jdff dff_B_lFo2OMaH8_1(.din(w_dff_B_b02joubA6_1),.dout(w_dff_B_lFo2OMaH8_1),.clk(gclk));
	jdff dff_B_UcOtnxf13_1(.din(w_dff_B_lFo2OMaH8_1),.dout(w_dff_B_UcOtnxf13_1),.clk(gclk));
	jdff dff_B_6tBjxt1n6_1(.din(w_dff_B_UcOtnxf13_1),.dout(w_dff_B_6tBjxt1n6_1),.clk(gclk));
	jdff dff_B_25EGAsJT6_1(.din(w_dff_B_6tBjxt1n6_1),.dout(w_dff_B_25EGAsJT6_1),.clk(gclk));
	jdff dff_B_NNt2IY2d5_1(.din(w_dff_B_25EGAsJT6_1),.dout(w_dff_B_NNt2IY2d5_1),.clk(gclk));
	jdff dff_B_P5Ut0wK42_1(.din(w_dff_B_NNt2IY2d5_1),.dout(w_dff_B_P5Ut0wK42_1),.clk(gclk));
	jdff dff_B_eXW653uy9_1(.din(w_dff_B_P5Ut0wK42_1),.dout(w_dff_B_eXW653uy9_1),.clk(gclk));
	jdff dff_B_mmHEHHQ00_1(.din(w_dff_B_eXW653uy9_1),.dout(w_dff_B_mmHEHHQ00_1),.clk(gclk));
	jdff dff_B_X2SMlDZf2_1(.din(w_dff_B_mmHEHHQ00_1),.dout(w_dff_B_X2SMlDZf2_1),.clk(gclk));
	jdff dff_B_Gp9j5lie5_1(.din(w_dff_B_X2SMlDZf2_1),.dout(w_dff_B_Gp9j5lie5_1),.clk(gclk));
	jdff dff_B_1xe2xa2b7_1(.din(w_dff_B_Gp9j5lie5_1),.dout(w_dff_B_1xe2xa2b7_1),.clk(gclk));
	jdff dff_B_xl4ky81B8_1(.din(w_dff_B_1xe2xa2b7_1),.dout(w_dff_B_xl4ky81B8_1),.clk(gclk));
	jdff dff_B_Nf1JW0Sy8_1(.din(w_dff_B_xl4ky81B8_1),.dout(w_dff_B_Nf1JW0Sy8_1),.clk(gclk));
	jdff dff_B_N3H7juG44_1(.din(w_dff_B_Nf1JW0Sy8_1),.dout(w_dff_B_N3H7juG44_1),.clk(gclk));
	jdff dff_B_RVBQFYe26_1(.din(w_dff_B_N3H7juG44_1),.dout(w_dff_B_RVBQFYe26_1),.clk(gclk));
	jdff dff_B_SehHSgxe9_1(.din(w_dff_B_RVBQFYe26_1),.dout(w_dff_B_SehHSgxe9_1),.clk(gclk));
	jdff dff_B_q9NQ572J1_1(.din(w_dff_B_SehHSgxe9_1),.dout(w_dff_B_q9NQ572J1_1),.clk(gclk));
	jdff dff_B_WygCBZrl0_1(.din(w_dff_B_q9NQ572J1_1),.dout(w_dff_B_WygCBZrl0_1),.clk(gclk));
	jdff dff_B_iCdOZC8v7_1(.din(w_dff_B_WygCBZrl0_1),.dout(w_dff_B_iCdOZC8v7_1),.clk(gclk));
	jdff dff_B_u78A3r9W2_1(.din(w_dff_B_iCdOZC8v7_1),.dout(w_dff_B_u78A3r9W2_1),.clk(gclk));
	jdff dff_B_WRVShjn52_1(.din(w_dff_B_u78A3r9W2_1),.dout(w_dff_B_WRVShjn52_1),.clk(gclk));
	jdff dff_B_oO46UanB4_1(.din(w_dff_B_WRVShjn52_1),.dout(w_dff_B_oO46UanB4_1),.clk(gclk));
	jdff dff_B_2ET4CGcy3_1(.din(w_dff_B_oO46UanB4_1),.dout(w_dff_B_2ET4CGcy3_1),.clk(gclk));
	jdff dff_B_3WVvWm4U8_1(.din(w_dff_B_2ET4CGcy3_1),.dout(w_dff_B_3WVvWm4U8_1),.clk(gclk));
	jdff dff_B_elvslTpM4_1(.din(w_dff_B_3WVvWm4U8_1),.dout(w_dff_B_elvslTpM4_1),.clk(gclk));
	jdff dff_B_0M3DidwV5_1(.din(w_dff_B_elvslTpM4_1),.dout(w_dff_B_0M3DidwV5_1),.clk(gclk));
	jdff dff_B_OtgaCh0k0_1(.din(w_dff_B_0M3DidwV5_1),.dout(w_dff_B_OtgaCh0k0_1),.clk(gclk));
	jdff dff_B_yzn87wbr0_1(.din(w_dff_B_OtgaCh0k0_1),.dout(w_dff_B_yzn87wbr0_1),.clk(gclk));
	jdff dff_B_EtQioman0_1(.din(w_dff_B_yzn87wbr0_1),.dout(w_dff_B_EtQioman0_1),.clk(gclk));
	jdff dff_B_X4TrKgAK2_1(.din(w_dff_B_EtQioman0_1),.dout(w_dff_B_X4TrKgAK2_1),.clk(gclk));
	jdff dff_B_12GyJk4w6_1(.din(w_dff_B_X4TrKgAK2_1),.dout(w_dff_B_12GyJk4w6_1),.clk(gclk));
	jdff dff_B_1iR8VOcz6_1(.din(w_dff_B_12GyJk4w6_1),.dout(w_dff_B_1iR8VOcz6_1),.clk(gclk));
	jdff dff_B_YDgGnJyk4_1(.din(w_dff_B_1iR8VOcz6_1),.dout(w_dff_B_YDgGnJyk4_1),.clk(gclk));
	jdff dff_B_TnMoPJkA0_1(.din(w_dff_B_YDgGnJyk4_1),.dout(w_dff_B_TnMoPJkA0_1),.clk(gclk));
	jdff dff_B_RrvzXPOb5_1(.din(w_dff_B_TnMoPJkA0_1),.dout(w_dff_B_RrvzXPOb5_1),.clk(gclk));
	jdff dff_B_KdMpr6kL5_1(.din(w_dff_B_RrvzXPOb5_1),.dout(w_dff_B_KdMpr6kL5_1),.clk(gclk));
	jdff dff_B_o6atlUfx5_1(.din(w_dff_B_KdMpr6kL5_1),.dout(w_dff_B_o6atlUfx5_1),.clk(gclk));
	jdff dff_B_vA0AJS1L9_1(.din(w_dff_B_o6atlUfx5_1),.dout(w_dff_B_vA0AJS1L9_1),.clk(gclk));
	jdff dff_B_G6sJ2W8p0_1(.din(w_dff_B_vA0AJS1L9_1),.dout(w_dff_B_G6sJ2W8p0_1),.clk(gclk));
	jdff dff_B_mPQaqsW65_1(.din(w_dff_B_G6sJ2W8p0_1),.dout(w_dff_B_mPQaqsW65_1),.clk(gclk));
	jdff dff_B_0QETm1X44_1(.din(w_dff_B_mPQaqsW65_1),.dout(w_dff_B_0QETm1X44_1),.clk(gclk));
	jdff dff_B_nOrAbU4z0_1(.din(w_dff_B_0QETm1X44_1),.dout(w_dff_B_nOrAbU4z0_1),.clk(gclk));
	jdff dff_B_JgYCvPNL1_1(.din(w_dff_B_nOrAbU4z0_1),.dout(w_dff_B_JgYCvPNL1_1),.clk(gclk));
	jdff dff_B_Sb8o7SrZ3_1(.din(w_dff_B_JgYCvPNL1_1),.dout(w_dff_B_Sb8o7SrZ3_1),.clk(gclk));
	jdff dff_B_Fx8y1IPI6_1(.din(w_dff_B_Sb8o7SrZ3_1),.dout(w_dff_B_Fx8y1IPI6_1),.clk(gclk));
	jdff dff_B_BLTTxahc2_1(.din(w_dff_B_Fx8y1IPI6_1),.dout(w_dff_B_BLTTxahc2_1),.clk(gclk));
	jdff dff_B_eBj6S86y0_1(.din(w_dff_B_BLTTxahc2_1),.dout(w_dff_B_eBj6S86y0_1),.clk(gclk));
	jdff dff_B_7W2V7Ewn4_1(.din(w_dff_B_eBj6S86y0_1),.dout(w_dff_B_7W2V7Ewn4_1),.clk(gclk));
	jdff dff_B_jZPdK1kZ9_1(.din(w_dff_B_7W2V7Ewn4_1),.dout(w_dff_B_jZPdK1kZ9_1),.clk(gclk));
	jdff dff_B_NvPygvMp7_1(.din(w_dff_B_jZPdK1kZ9_1),.dout(w_dff_B_NvPygvMp7_1),.clk(gclk));
	jdff dff_B_Vor6ZZVU5_1(.din(w_dff_B_NvPygvMp7_1),.dout(w_dff_B_Vor6ZZVU5_1),.clk(gclk));
	jdff dff_B_vZsSDmqN4_1(.din(w_dff_B_Vor6ZZVU5_1),.dout(w_dff_B_vZsSDmqN4_1),.clk(gclk));
	jdff dff_B_dtYczj4u5_1(.din(w_dff_B_vZsSDmqN4_1),.dout(w_dff_B_dtYczj4u5_1),.clk(gclk));
	jdff dff_B_OcRBzI3e0_1(.din(w_dff_B_dtYczj4u5_1),.dout(w_dff_B_OcRBzI3e0_1),.clk(gclk));
	jdff dff_B_6uWEU51u0_1(.din(w_dff_B_OcRBzI3e0_1),.dout(w_dff_B_6uWEU51u0_1),.clk(gclk));
	jdff dff_B_CPLyEXKS6_1(.din(w_dff_B_6uWEU51u0_1),.dout(w_dff_B_CPLyEXKS6_1),.clk(gclk));
	jdff dff_B_Arn7DGHt6_1(.din(w_dff_B_CPLyEXKS6_1),.dout(w_dff_B_Arn7DGHt6_1),.clk(gclk));
	jdff dff_B_ZbMRvaeY4_1(.din(w_dff_B_Arn7DGHt6_1),.dout(w_dff_B_ZbMRvaeY4_1),.clk(gclk));
	jdff dff_B_Gg0qI4IW3_1(.din(w_dff_B_ZbMRvaeY4_1),.dout(w_dff_B_Gg0qI4IW3_1),.clk(gclk));
	jdff dff_B_KdYG81lr0_1(.din(w_dff_B_Gg0qI4IW3_1),.dout(w_dff_B_KdYG81lr0_1),.clk(gclk));
	jdff dff_B_DvnUCB5e3_1(.din(w_dff_B_KdYG81lr0_1),.dout(w_dff_B_DvnUCB5e3_1),.clk(gclk));
	jdff dff_B_WB80gDUQ3_1(.din(w_dff_B_DvnUCB5e3_1),.dout(w_dff_B_WB80gDUQ3_1),.clk(gclk));
	jdff dff_B_GjGh3WJu0_0(.din(n967),.dout(w_dff_B_GjGh3WJu0_0),.clk(gclk));
	jdff dff_B_87AHIjf61_0(.din(w_dff_B_GjGh3WJu0_0),.dout(w_dff_B_87AHIjf61_0),.clk(gclk));
	jdff dff_B_vha20V114_0(.din(w_dff_B_87AHIjf61_0),.dout(w_dff_B_vha20V114_0),.clk(gclk));
	jdff dff_B_IIWhL9Oy6_0(.din(w_dff_B_vha20V114_0),.dout(w_dff_B_IIWhL9Oy6_0),.clk(gclk));
	jdff dff_B_0xPVz5iZ6_0(.din(w_dff_B_IIWhL9Oy6_0),.dout(w_dff_B_0xPVz5iZ6_0),.clk(gclk));
	jdff dff_B_c73mP7TR4_0(.din(w_dff_B_0xPVz5iZ6_0),.dout(w_dff_B_c73mP7TR4_0),.clk(gclk));
	jdff dff_B_KMt2Vp601_0(.din(w_dff_B_c73mP7TR4_0),.dout(w_dff_B_KMt2Vp601_0),.clk(gclk));
	jdff dff_B_56mdr7yb8_0(.din(w_dff_B_KMt2Vp601_0),.dout(w_dff_B_56mdr7yb8_0),.clk(gclk));
	jdff dff_B_INlpUnzy1_0(.din(w_dff_B_56mdr7yb8_0),.dout(w_dff_B_INlpUnzy1_0),.clk(gclk));
	jdff dff_B_5iQ9aL7I9_0(.din(w_dff_B_INlpUnzy1_0),.dout(w_dff_B_5iQ9aL7I9_0),.clk(gclk));
	jdff dff_B_K2iAn8p76_0(.din(w_dff_B_5iQ9aL7I9_0),.dout(w_dff_B_K2iAn8p76_0),.clk(gclk));
	jdff dff_B_EHRxyDpz5_0(.din(w_dff_B_K2iAn8p76_0),.dout(w_dff_B_EHRxyDpz5_0),.clk(gclk));
	jdff dff_B_tkwPMeTL4_0(.din(w_dff_B_EHRxyDpz5_0),.dout(w_dff_B_tkwPMeTL4_0),.clk(gclk));
	jdff dff_B_k2dibsWK2_0(.din(w_dff_B_tkwPMeTL4_0),.dout(w_dff_B_k2dibsWK2_0),.clk(gclk));
	jdff dff_B_Z9ofRIyT9_0(.din(w_dff_B_k2dibsWK2_0),.dout(w_dff_B_Z9ofRIyT9_0),.clk(gclk));
	jdff dff_B_QMMpuiUz2_0(.din(w_dff_B_Z9ofRIyT9_0),.dout(w_dff_B_QMMpuiUz2_0),.clk(gclk));
	jdff dff_B_kkRvZaQa9_0(.din(w_dff_B_QMMpuiUz2_0),.dout(w_dff_B_kkRvZaQa9_0),.clk(gclk));
	jdff dff_B_RrEFziYm2_0(.din(w_dff_B_kkRvZaQa9_0),.dout(w_dff_B_RrEFziYm2_0),.clk(gclk));
	jdff dff_B_UkeEDUmI1_0(.din(w_dff_B_RrEFziYm2_0),.dout(w_dff_B_UkeEDUmI1_0),.clk(gclk));
	jdff dff_B_thld9spP1_0(.din(w_dff_B_UkeEDUmI1_0),.dout(w_dff_B_thld9spP1_0),.clk(gclk));
	jdff dff_B_5vfUe3Zu0_0(.din(w_dff_B_thld9spP1_0),.dout(w_dff_B_5vfUe3Zu0_0),.clk(gclk));
	jdff dff_B_YNbHDSyk2_0(.din(w_dff_B_5vfUe3Zu0_0),.dout(w_dff_B_YNbHDSyk2_0),.clk(gclk));
	jdff dff_B_XPehuPkM0_0(.din(w_dff_B_YNbHDSyk2_0),.dout(w_dff_B_XPehuPkM0_0),.clk(gclk));
	jdff dff_B_ZdPUWvF32_0(.din(w_dff_B_XPehuPkM0_0),.dout(w_dff_B_ZdPUWvF32_0),.clk(gclk));
	jdff dff_B_xelrXhYO3_0(.din(w_dff_B_ZdPUWvF32_0),.dout(w_dff_B_xelrXhYO3_0),.clk(gclk));
	jdff dff_B_4mo0fLKN6_0(.din(w_dff_B_xelrXhYO3_0),.dout(w_dff_B_4mo0fLKN6_0),.clk(gclk));
	jdff dff_B_JNHaoWyZ1_0(.din(w_dff_B_4mo0fLKN6_0),.dout(w_dff_B_JNHaoWyZ1_0),.clk(gclk));
	jdff dff_B_bZujMI7a4_0(.din(w_dff_B_JNHaoWyZ1_0),.dout(w_dff_B_bZujMI7a4_0),.clk(gclk));
	jdff dff_B_axWWilLA8_0(.din(w_dff_B_bZujMI7a4_0),.dout(w_dff_B_axWWilLA8_0),.clk(gclk));
	jdff dff_B_nyEmfRx03_0(.din(w_dff_B_axWWilLA8_0),.dout(w_dff_B_nyEmfRx03_0),.clk(gclk));
	jdff dff_B_xxQqm72r2_0(.din(w_dff_B_nyEmfRx03_0),.dout(w_dff_B_xxQqm72r2_0),.clk(gclk));
	jdff dff_B_sJLemPYT6_0(.din(w_dff_B_xxQqm72r2_0),.dout(w_dff_B_sJLemPYT6_0),.clk(gclk));
	jdff dff_B_7sprYiKU5_0(.din(w_dff_B_sJLemPYT6_0),.dout(w_dff_B_7sprYiKU5_0),.clk(gclk));
	jdff dff_B_e76x8MDY9_0(.din(w_dff_B_7sprYiKU5_0),.dout(w_dff_B_e76x8MDY9_0),.clk(gclk));
	jdff dff_B_KrEvJ6Em0_0(.din(w_dff_B_e76x8MDY9_0),.dout(w_dff_B_KrEvJ6Em0_0),.clk(gclk));
	jdff dff_B_9VOd76IC5_0(.din(w_dff_B_KrEvJ6Em0_0),.dout(w_dff_B_9VOd76IC5_0),.clk(gclk));
	jdff dff_B_kdcXW1Dn7_0(.din(w_dff_B_9VOd76IC5_0),.dout(w_dff_B_kdcXW1Dn7_0),.clk(gclk));
	jdff dff_B_a3CTIul14_0(.din(w_dff_B_kdcXW1Dn7_0),.dout(w_dff_B_a3CTIul14_0),.clk(gclk));
	jdff dff_B_GtMlnX143_0(.din(w_dff_B_a3CTIul14_0),.dout(w_dff_B_GtMlnX143_0),.clk(gclk));
	jdff dff_B_kF67EOkP8_0(.din(w_dff_B_GtMlnX143_0),.dout(w_dff_B_kF67EOkP8_0),.clk(gclk));
	jdff dff_B_dvgxW1fE9_0(.din(w_dff_B_kF67EOkP8_0),.dout(w_dff_B_dvgxW1fE9_0),.clk(gclk));
	jdff dff_B_fqpPdD304_0(.din(w_dff_B_dvgxW1fE9_0),.dout(w_dff_B_fqpPdD304_0),.clk(gclk));
	jdff dff_B_CAJyC8AI6_0(.din(w_dff_B_fqpPdD304_0),.dout(w_dff_B_CAJyC8AI6_0),.clk(gclk));
	jdff dff_B_NsncFfJi6_0(.din(w_dff_B_CAJyC8AI6_0),.dout(w_dff_B_NsncFfJi6_0),.clk(gclk));
	jdff dff_B_1Sn1fci71_0(.din(w_dff_B_NsncFfJi6_0),.dout(w_dff_B_1Sn1fci71_0),.clk(gclk));
	jdff dff_B_cartHQiF5_0(.din(w_dff_B_1Sn1fci71_0),.dout(w_dff_B_cartHQiF5_0),.clk(gclk));
	jdff dff_B_K7ajf5zH2_0(.din(w_dff_B_cartHQiF5_0),.dout(w_dff_B_K7ajf5zH2_0),.clk(gclk));
	jdff dff_B_9T7E4BJm4_0(.din(w_dff_B_K7ajf5zH2_0),.dout(w_dff_B_9T7E4BJm4_0),.clk(gclk));
	jdff dff_B_cBsNe0Kj1_0(.din(w_dff_B_9T7E4BJm4_0),.dout(w_dff_B_cBsNe0Kj1_0),.clk(gclk));
	jdff dff_B_EhJ4eNRk3_0(.din(w_dff_B_cBsNe0Kj1_0),.dout(w_dff_B_EhJ4eNRk3_0),.clk(gclk));
	jdff dff_B_JzYWfGWg9_0(.din(w_dff_B_EhJ4eNRk3_0),.dout(w_dff_B_JzYWfGWg9_0),.clk(gclk));
	jdff dff_B_6VMSdjb25_0(.din(w_dff_B_JzYWfGWg9_0),.dout(w_dff_B_6VMSdjb25_0),.clk(gclk));
	jdff dff_B_3pd9mDXE9_0(.din(w_dff_B_6VMSdjb25_0),.dout(w_dff_B_3pd9mDXE9_0),.clk(gclk));
	jdff dff_B_Ti5ZiTDw4_0(.din(w_dff_B_3pd9mDXE9_0),.dout(w_dff_B_Ti5ZiTDw4_0),.clk(gclk));
	jdff dff_B_Y8s4ZyLT4_0(.din(w_dff_B_Ti5ZiTDw4_0),.dout(w_dff_B_Y8s4ZyLT4_0),.clk(gclk));
	jdff dff_B_rQT0WRwO0_0(.din(w_dff_B_Y8s4ZyLT4_0),.dout(w_dff_B_rQT0WRwO0_0),.clk(gclk));
	jdff dff_B_QNrAjY2s8_0(.din(w_dff_B_rQT0WRwO0_0),.dout(w_dff_B_QNrAjY2s8_0),.clk(gclk));
	jdff dff_B_THshr7nV5_0(.din(w_dff_B_QNrAjY2s8_0),.dout(w_dff_B_THshr7nV5_0),.clk(gclk));
	jdff dff_B_q2b5Mr069_0(.din(w_dff_B_THshr7nV5_0),.dout(w_dff_B_q2b5Mr069_0),.clk(gclk));
	jdff dff_B_QcFVbgt62_0(.din(w_dff_B_q2b5Mr069_0),.dout(w_dff_B_QcFVbgt62_0),.clk(gclk));
	jdff dff_B_npoZexg99_0(.din(w_dff_B_QcFVbgt62_0),.dout(w_dff_B_npoZexg99_0),.clk(gclk));
	jdff dff_B_eyeMZbHu8_0(.din(w_dff_B_npoZexg99_0),.dout(w_dff_B_eyeMZbHu8_0),.clk(gclk));
	jdff dff_B_gpj5eUpe6_0(.din(w_dff_B_eyeMZbHu8_0),.dout(w_dff_B_gpj5eUpe6_0),.clk(gclk));
	jdff dff_B_RTy8gz0z3_0(.din(w_dff_B_gpj5eUpe6_0),.dout(w_dff_B_RTy8gz0z3_0),.clk(gclk));
	jdff dff_B_NN3NZ2ah9_0(.din(w_dff_B_RTy8gz0z3_0),.dout(w_dff_B_NN3NZ2ah9_0),.clk(gclk));
	jdff dff_B_hhjmCZRY8_0(.din(w_dff_B_NN3NZ2ah9_0),.dout(w_dff_B_hhjmCZRY8_0),.clk(gclk));
	jdff dff_B_dAOVQXDY8_0(.din(w_dff_B_hhjmCZRY8_0),.dout(w_dff_B_dAOVQXDY8_0),.clk(gclk));
	jdff dff_B_fsAZWSZI7_0(.din(w_dff_B_dAOVQXDY8_0),.dout(w_dff_B_fsAZWSZI7_0),.clk(gclk));
	jdff dff_B_M5DZCPvj6_0(.din(w_dff_B_fsAZWSZI7_0),.dout(w_dff_B_M5DZCPvj6_0),.clk(gclk));
	jdff dff_B_pdNiP3hC7_0(.din(w_dff_B_M5DZCPvj6_0),.dout(w_dff_B_pdNiP3hC7_0),.clk(gclk));
	jdff dff_B_W2REQXXw7_0(.din(w_dff_B_pdNiP3hC7_0),.dout(w_dff_B_W2REQXXw7_0),.clk(gclk));
	jdff dff_B_r47RgOHP5_0(.din(w_dff_B_W2REQXXw7_0),.dout(w_dff_B_r47RgOHP5_0),.clk(gclk));
	jdff dff_B_V7Vyc3sJ1_0(.din(w_dff_B_r47RgOHP5_0),.dout(w_dff_B_V7Vyc3sJ1_0),.clk(gclk));
	jdff dff_B_S4OLg2yr2_0(.din(w_dff_B_V7Vyc3sJ1_0),.dout(w_dff_B_S4OLg2yr2_0),.clk(gclk));
	jdff dff_B_ar8XvTH63_0(.din(w_dff_B_S4OLg2yr2_0),.dout(w_dff_B_ar8XvTH63_0),.clk(gclk));
	jdff dff_B_pJ7az45L4_0(.din(w_dff_B_ar8XvTH63_0),.dout(w_dff_B_pJ7az45L4_0),.clk(gclk));
	jdff dff_B_ag80TtA29_0(.din(w_dff_B_pJ7az45L4_0),.dout(w_dff_B_ag80TtA29_0),.clk(gclk));
	jdff dff_B_udxludNu2_0(.din(w_dff_B_ag80TtA29_0),.dout(w_dff_B_udxludNu2_0),.clk(gclk));
	jdff dff_B_c4uWKt9O0_0(.din(w_dff_B_udxludNu2_0),.dout(w_dff_B_c4uWKt9O0_0),.clk(gclk));
	jdff dff_B_d8k9JwJL6_0(.din(w_dff_B_c4uWKt9O0_0),.dout(w_dff_B_d8k9JwJL6_0),.clk(gclk));
	jdff dff_B_KQa96zfY2_0(.din(w_dff_B_d8k9JwJL6_0),.dout(w_dff_B_KQa96zfY2_0),.clk(gclk));
	jdff dff_B_HMMi7YPO4_0(.din(w_dff_B_KQa96zfY2_0),.dout(w_dff_B_HMMi7YPO4_0),.clk(gclk));
	jdff dff_B_VMDwLyZ19_0(.din(w_dff_B_HMMi7YPO4_0),.dout(w_dff_B_VMDwLyZ19_0),.clk(gclk));
	jdff dff_B_x1VH9U9f5_0(.din(w_dff_B_VMDwLyZ19_0),.dout(w_dff_B_x1VH9U9f5_0),.clk(gclk));
	jdff dff_B_e5ZhdMUD9_0(.din(w_dff_B_x1VH9U9f5_0),.dout(w_dff_B_e5ZhdMUD9_0),.clk(gclk));
	jdff dff_B_c32iPo0W0_0(.din(w_dff_B_e5ZhdMUD9_0),.dout(w_dff_B_c32iPo0W0_0),.clk(gclk));
	jdff dff_B_NvmzhQFe8_0(.din(w_dff_B_c32iPo0W0_0),.dout(w_dff_B_NvmzhQFe8_0),.clk(gclk));
	jdff dff_B_QJlmnVcJ9_0(.din(w_dff_B_NvmzhQFe8_0),.dout(w_dff_B_QJlmnVcJ9_0),.clk(gclk));
	jdff dff_B_OwnieKJd8_0(.din(w_dff_B_QJlmnVcJ9_0),.dout(w_dff_B_OwnieKJd8_0),.clk(gclk));
	jdff dff_B_fdbEgXEg2_0(.din(w_dff_B_OwnieKJd8_0),.dout(w_dff_B_fdbEgXEg2_0),.clk(gclk));
	jdff dff_B_FiNcMpAP6_0(.din(w_dff_B_fdbEgXEg2_0),.dout(w_dff_B_FiNcMpAP6_0),.clk(gclk));
	jdff dff_B_X7BNpBXy1_0(.din(w_dff_B_FiNcMpAP6_0),.dout(w_dff_B_X7BNpBXy1_0),.clk(gclk));
	jdff dff_B_DfkeKuht3_0(.din(w_dff_B_X7BNpBXy1_0),.dout(w_dff_B_DfkeKuht3_0),.clk(gclk));
	jdff dff_B_0kwJxems0_0(.din(w_dff_B_DfkeKuht3_0),.dout(w_dff_B_0kwJxems0_0),.clk(gclk));
	jdff dff_B_rO5HQhB26_0(.din(w_dff_B_0kwJxems0_0),.dout(w_dff_B_rO5HQhB26_0),.clk(gclk));
	jdff dff_B_mULJ6y7Q6_0(.din(w_dff_B_rO5HQhB26_0),.dout(w_dff_B_mULJ6y7Q6_0),.clk(gclk));
	jdff dff_B_XE2iBHU27_0(.din(w_dff_B_mULJ6y7Q6_0),.dout(w_dff_B_XE2iBHU27_0),.clk(gclk));
	jdff dff_B_X6k1QGWv0_1(.din(n960),.dout(w_dff_B_X6k1QGWv0_1),.clk(gclk));
	jdff dff_B_OhruMBzk6_1(.din(w_dff_B_X6k1QGWv0_1),.dout(w_dff_B_OhruMBzk6_1),.clk(gclk));
	jdff dff_B_gsAuGk6a3_1(.din(w_dff_B_OhruMBzk6_1),.dout(w_dff_B_gsAuGk6a3_1),.clk(gclk));
	jdff dff_B_qDbiWVZy8_1(.din(w_dff_B_gsAuGk6a3_1),.dout(w_dff_B_qDbiWVZy8_1),.clk(gclk));
	jdff dff_B_mdI0Fwlk3_1(.din(w_dff_B_qDbiWVZy8_1),.dout(w_dff_B_mdI0Fwlk3_1),.clk(gclk));
	jdff dff_B_v0aIkXA33_1(.din(w_dff_B_mdI0Fwlk3_1),.dout(w_dff_B_v0aIkXA33_1),.clk(gclk));
	jdff dff_B_eoAtNEcx1_1(.din(w_dff_B_v0aIkXA33_1),.dout(w_dff_B_eoAtNEcx1_1),.clk(gclk));
	jdff dff_B_tYpqItOU8_1(.din(w_dff_B_eoAtNEcx1_1),.dout(w_dff_B_tYpqItOU8_1),.clk(gclk));
	jdff dff_B_PgdDTKDx1_1(.din(w_dff_B_tYpqItOU8_1),.dout(w_dff_B_PgdDTKDx1_1),.clk(gclk));
	jdff dff_B_3mETEtpF9_1(.din(w_dff_B_PgdDTKDx1_1),.dout(w_dff_B_3mETEtpF9_1),.clk(gclk));
	jdff dff_B_fTJalLeC5_1(.din(w_dff_B_3mETEtpF9_1),.dout(w_dff_B_fTJalLeC5_1),.clk(gclk));
	jdff dff_B_1HEa7eRm2_1(.din(w_dff_B_fTJalLeC5_1),.dout(w_dff_B_1HEa7eRm2_1),.clk(gclk));
	jdff dff_B_hlHz8Q0g6_1(.din(w_dff_B_1HEa7eRm2_1),.dout(w_dff_B_hlHz8Q0g6_1),.clk(gclk));
	jdff dff_B_tEVcGN6p7_1(.din(w_dff_B_hlHz8Q0g6_1),.dout(w_dff_B_tEVcGN6p7_1),.clk(gclk));
	jdff dff_B_ECeAd9Bq2_1(.din(w_dff_B_tEVcGN6p7_1),.dout(w_dff_B_ECeAd9Bq2_1),.clk(gclk));
	jdff dff_B_JMLzCD4R4_1(.din(w_dff_B_ECeAd9Bq2_1),.dout(w_dff_B_JMLzCD4R4_1),.clk(gclk));
	jdff dff_B_UdIWccTE0_1(.din(w_dff_B_JMLzCD4R4_1),.dout(w_dff_B_UdIWccTE0_1),.clk(gclk));
	jdff dff_B_BpAHrHRS0_1(.din(w_dff_B_UdIWccTE0_1),.dout(w_dff_B_BpAHrHRS0_1),.clk(gclk));
	jdff dff_B_BBfgyF8V9_1(.din(w_dff_B_BpAHrHRS0_1),.dout(w_dff_B_BBfgyF8V9_1),.clk(gclk));
	jdff dff_B_tHrlVO5A4_1(.din(w_dff_B_BBfgyF8V9_1),.dout(w_dff_B_tHrlVO5A4_1),.clk(gclk));
	jdff dff_B_bdKhbPu02_1(.din(w_dff_B_tHrlVO5A4_1),.dout(w_dff_B_bdKhbPu02_1),.clk(gclk));
	jdff dff_B_ndFRSCRI2_1(.din(w_dff_B_bdKhbPu02_1),.dout(w_dff_B_ndFRSCRI2_1),.clk(gclk));
	jdff dff_B_8jsUJxoz9_1(.din(w_dff_B_ndFRSCRI2_1),.dout(w_dff_B_8jsUJxoz9_1),.clk(gclk));
	jdff dff_B_LN3jD4Wz5_1(.din(w_dff_B_8jsUJxoz9_1),.dout(w_dff_B_LN3jD4Wz5_1),.clk(gclk));
	jdff dff_B_IiLloUit1_1(.din(w_dff_B_LN3jD4Wz5_1),.dout(w_dff_B_IiLloUit1_1),.clk(gclk));
	jdff dff_B_gaRITIlM0_1(.din(w_dff_B_IiLloUit1_1),.dout(w_dff_B_gaRITIlM0_1),.clk(gclk));
	jdff dff_B_Eyru6rLW5_1(.din(w_dff_B_gaRITIlM0_1),.dout(w_dff_B_Eyru6rLW5_1),.clk(gclk));
	jdff dff_B_prMpyePJ0_1(.din(w_dff_B_Eyru6rLW5_1),.dout(w_dff_B_prMpyePJ0_1),.clk(gclk));
	jdff dff_B_M0QL4oJg0_1(.din(w_dff_B_prMpyePJ0_1),.dout(w_dff_B_M0QL4oJg0_1),.clk(gclk));
	jdff dff_B_mW5VNVn62_1(.din(w_dff_B_M0QL4oJg0_1),.dout(w_dff_B_mW5VNVn62_1),.clk(gclk));
	jdff dff_B_IYu9f9W17_1(.din(w_dff_B_mW5VNVn62_1),.dout(w_dff_B_IYu9f9W17_1),.clk(gclk));
	jdff dff_B_8aiJyBES7_1(.din(w_dff_B_IYu9f9W17_1),.dout(w_dff_B_8aiJyBES7_1),.clk(gclk));
	jdff dff_B_OvqpOZDC8_1(.din(w_dff_B_8aiJyBES7_1),.dout(w_dff_B_OvqpOZDC8_1),.clk(gclk));
	jdff dff_B_iVESutl40_1(.din(w_dff_B_OvqpOZDC8_1),.dout(w_dff_B_iVESutl40_1),.clk(gclk));
	jdff dff_B_j1Bhpc6S4_1(.din(w_dff_B_iVESutl40_1),.dout(w_dff_B_j1Bhpc6S4_1),.clk(gclk));
	jdff dff_B_sR7Zp4OF8_1(.din(w_dff_B_j1Bhpc6S4_1),.dout(w_dff_B_sR7Zp4OF8_1),.clk(gclk));
	jdff dff_B_CQ8Y6tTp1_1(.din(w_dff_B_sR7Zp4OF8_1),.dout(w_dff_B_CQ8Y6tTp1_1),.clk(gclk));
	jdff dff_B_MFws36604_1(.din(w_dff_B_CQ8Y6tTp1_1),.dout(w_dff_B_MFws36604_1),.clk(gclk));
	jdff dff_B_XtPZyC9D8_1(.din(w_dff_B_MFws36604_1),.dout(w_dff_B_XtPZyC9D8_1),.clk(gclk));
	jdff dff_B_Tmu3Mwki4_1(.din(w_dff_B_XtPZyC9D8_1),.dout(w_dff_B_Tmu3Mwki4_1),.clk(gclk));
	jdff dff_B_GC8IoMHt4_1(.din(w_dff_B_Tmu3Mwki4_1),.dout(w_dff_B_GC8IoMHt4_1),.clk(gclk));
	jdff dff_B_voBOfHj30_1(.din(w_dff_B_GC8IoMHt4_1),.dout(w_dff_B_voBOfHj30_1),.clk(gclk));
	jdff dff_B_01dYlaXF0_1(.din(w_dff_B_voBOfHj30_1),.dout(w_dff_B_01dYlaXF0_1),.clk(gclk));
	jdff dff_B_5k79iCEF9_1(.din(w_dff_B_01dYlaXF0_1),.dout(w_dff_B_5k79iCEF9_1),.clk(gclk));
	jdff dff_B_z15N4nXr3_1(.din(w_dff_B_5k79iCEF9_1),.dout(w_dff_B_z15N4nXr3_1),.clk(gclk));
	jdff dff_B_cmbJVVmN0_1(.din(w_dff_B_z15N4nXr3_1),.dout(w_dff_B_cmbJVVmN0_1),.clk(gclk));
	jdff dff_B_uVjcN9o64_1(.din(w_dff_B_cmbJVVmN0_1),.dout(w_dff_B_uVjcN9o64_1),.clk(gclk));
	jdff dff_B_C5TPksbH6_1(.din(w_dff_B_uVjcN9o64_1),.dout(w_dff_B_C5TPksbH6_1),.clk(gclk));
	jdff dff_B_itlApGNA6_1(.din(w_dff_B_C5TPksbH6_1),.dout(w_dff_B_itlApGNA6_1),.clk(gclk));
	jdff dff_B_Kv4cd13c7_1(.din(w_dff_B_itlApGNA6_1),.dout(w_dff_B_Kv4cd13c7_1),.clk(gclk));
	jdff dff_B_fEarABeZ6_1(.din(w_dff_B_Kv4cd13c7_1),.dout(w_dff_B_fEarABeZ6_1),.clk(gclk));
	jdff dff_B_kVYTvMoH9_1(.din(w_dff_B_fEarABeZ6_1),.dout(w_dff_B_kVYTvMoH9_1),.clk(gclk));
	jdff dff_B_c9ljnnf46_1(.din(w_dff_B_kVYTvMoH9_1),.dout(w_dff_B_c9ljnnf46_1),.clk(gclk));
	jdff dff_B_bIXfaSag4_1(.din(w_dff_B_c9ljnnf46_1),.dout(w_dff_B_bIXfaSag4_1),.clk(gclk));
	jdff dff_B_gUG2cZ7F5_1(.din(w_dff_B_bIXfaSag4_1),.dout(w_dff_B_gUG2cZ7F5_1),.clk(gclk));
	jdff dff_B_edydH8W29_1(.din(w_dff_B_gUG2cZ7F5_1),.dout(w_dff_B_edydH8W29_1),.clk(gclk));
	jdff dff_B_a3cgnRV14_1(.din(w_dff_B_edydH8W29_1),.dout(w_dff_B_a3cgnRV14_1),.clk(gclk));
	jdff dff_B_WA2kttRh7_1(.din(w_dff_B_a3cgnRV14_1),.dout(w_dff_B_WA2kttRh7_1),.clk(gclk));
	jdff dff_B_gSjKMQhC3_1(.din(w_dff_B_WA2kttRh7_1),.dout(w_dff_B_gSjKMQhC3_1),.clk(gclk));
	jdff dff_B_uorQ4rQZ4_1(.din(w_dff_B_gSjKMQhC3_1),.dout(w_dff_B_uorQ4rQZ4_1),.clk(gclk));
	jdff dff_B_8UMElZlA7_1(.din(w_dff_B_uorQ4rQZ4_1),.dout(w_dff_B_8UMElZlA7_1),.clk(gclk));
	jdff dff_B_JT2icPdU2_1(.din(w_dff_B_8UMElZlA7_1),.dout(w_dff_B_JT2icPdU2_1),.clk(gclk));
	jdff dff_B_jFKnzbEl5_1(.din(w_dff_B_JT2icPdU2_1),.dout(w_dff_B_jFKnzbEl5_1),.clk(gclk));
	jdff dff_B_ODhwVTrS3_1(.din(w_dff_B_jFKnzbEl5_1),.dout(w_dff_B_ODhwVTrS3_1),.clk(gclk));
	jdff dff_B_48nzjYbs5_1(.din(w_dff_B_ODhwVTrS3_1),.dout(w_dff_B_48nzjYbs5_1),.clk(gclk));
	jdff dff_B_Rsc1aUEr9_1(.din(w_dff_B_48nzjYbs5_1),.dout(w_dff_B_Rsc1aUEr9_1),.clk(gclk));
	jdff dff_B_Z7YP2Vpt9_1(.din(w_dff_B_Rsc1aUEr9_1),.dout(w_dff_B_Z7YP2Vpt9_1),.clk(gclk));
	jdff dff_B_9sDBfI0c8_1(.din(w_dff_B_Z7YP2Vpt9_1),.dout(w_dff_B_9sDBfI0c8_1),.clk(gclk));
	jdff dff_B_hiEntRbO6_1(.din(w_dff_B_9sDBfI0c8_1),.dout(w_dff_B_hiEntRbO6_1),.clk(gclk));
	jdff dff_B_1gglhluY3_1(.din(w_dff_B_hiEntRbO6_1),.dout(w_dff_B_1gglhluY3_1),.clk(gclk));
	jdff dff_B_dStCm4rp2_1(.din(w_dff_B_1gglhluY3_1),.dout(w_dff_B_dStCm4rp2_1),.clk(gclk));
	jdff dff_B_aiL9QGwt6_1(.din(w_dff_B_dStCm4rp2_1),.dout(w_dff_B_aiL9QGwt6_1),.clk(gclk));
	jdff dff_B_1Mm6isHR0_1(.din(w_dff_B_aiL9QGwt6_1),.dout(w_dff_B_1Mm6isHR0_1),.clk(gclk));
	jdff dff_B_N1y6wS8K6_1(.din(w_dff_B_1Mm6isHR0_1),.dout(w_dff_B_N1y6wS8K6_1),.clk(gclk));
	jdff dff_B_HyXTneoF4_1(.din(w_dff_B_N1y6wS8K6_1),.dout(w_dff_B_HyXTneoF4_1),.clk(gclk));
	jdff dff_B_ezmF7k1U0_1(.din(w_dff_B_HyXTneoF4_1),.dout(w_dff_B_ezmF7k1U0_1),.clk(gclk));
	jdff dff_B_t0svJczu1_1(.din(w_dff_B_ezmF7k1U0_1),.dout(w_dff_B_t0svJczu1_1),.clk(gclk));
	jdff dff_B_NGAQV2UX8_1(.din(w_dff_B_t0svJczu1_1),.dout(w_dff_B_NGAQV2UX8_1),.clk(gclk));
	jdff dff_B_etEj1QAX0_1(.din(w_dff_B_NGAQV2UX8_1),.dout(w_dff_B_etEj1QAX0_1),.clk(gclk));
	jdff dff_B_JXLDJJ4g0_1(.din(w_dff_B_etEj1QAX0_1),.dout(w_dff_B_JXLDJJ4g0_1),.clk(gclk));
	jdff dff_B_17ZWHBFQ0_1(.din(w_dff_B_JXLDJJ4g0_1),.dout(w_dff_B_17ZWHBFQ0_1),.clk(gclk));
	jdff dff_B_91IWJTxR5_1(.din(w_dff_B_17ZWHBFQ0_1),.dout(w_dff_B_91IWJTxR5_1),.clk(gclk));
	jdff dff_B_xfwwyH7Y4_1(.din(w_dff_B_91IWJTxR5_1),.dout(w_dff_B_xfwwyH7Y4_1),.clk(gclk));
	jdff dff_B_0LZhZyG82_1(.din(w_dff_B_xfwwyH7Y4_1),.dout(w_dff_B_0LZhZyG82_1),.clk(gclk));
	jdff dff_B_Tm3iqxpu1_1(.din(w_dff_B_0LZhZyG82_1),.dout(w_dff_B_Tm3iqxpu1_1),.clk(gclk));
	jdff dff_B_gNXKhCuS8_1(.din(w_dff_B_Tm3iqxpu1_1),.dout(w_dff_B_gNXKhCuS8_1),.clk(gclk));
	jdff dff_B_Ju22jkuY5_1(.din(w_dff_B_gNXKhCuS8_1),.dout(w_dff_B_Ju22jkuY5_1),.clk(gclk));
	jdff dff_B_nMUlxsrx1_1(.din(w_dff_B_Ju22jkuY5_1),.dout(w_dff_B_nMUlxsrx1_1),.clk(gclk));
	jdff dff_B_SUXm0i3Q9_1(.din(w_dff_B_nMUlxsrx1_1),.dout(w_dff_B_SUXm0i3Q9_1),.clk(gclk));
	jdff dff_B_7YGRiLKz7_1(.din(w_dff_B_SUXm0i3Q9_1),.dout(w_dff_B_7YGRiLKz7_1),.clk(gclk));
	jdff dff_B_wS9Y9S1n7_1(.din(w_dff_B_7YGRiLKz7_1),.dout(w_dff_B_wS9Y9S1n7_1),.clk(gclk));
	jdff dff_B_o6dyVh8f7_1(.din(w_dff_B_wS9Y9S1n7_1),.dout(w_dff_B_o6dyVh8f7_1),.clk(gclk));
	jdff dff_B_mGVgvzrS8_1(.din(w_dff_B_o6dyVh8f7_1),.dout(w_dff_B_mGVgvzrS8_1),.clk(gclk));
	jdff dff_B_zk07ZSL38_1(.din(w_dff_B_mGVgvzrS8_1),.dout(w_dff_B_zk07ZSL38_1),.clk(gclk));
	jdff dff_B_66FJgh837_1(.din(w_dff_B_zk07ZSL38_1),.dout(w_dff_B_66FJgh837_1),.clk(gclk));
	jdff dff_B_i16ixeFE0_1(.din(w_dff_B_66FJgh837_1),.dout(w_dff_B_i16ixeFE0_1),.clk(gclk));
	jdff dff_B_pB9ohBpz5_0(.din(n961),.dout(w_dff_B_pB9ohBpz5_0),.clk(gclk));
	jdff dff_B_qN5gVHgU3_0(.din(w_dff_B_pB9ohBpz5_0),.dout(w_dff_B_qN5gVHgU3_0),.clk(gclk));
	jdff dff_B_4t1mlIvC3_0(.din(w_dff_B_qN5gVHgU3_0),.dout(w_dff_B_4t1mlIvC3_0),.clk(gclk));
	jdff dff_B_FURDTsYV5_0(.din(w_dff_B_4t1mlIvC3_0),.dout(w_dff_B_FURDTsYV5_0),.clk(gclk));
	jdff dff_B_MBdieqMe0_0(.din(w_dff_B_FURDTsYV5_0),.dout(w_dff_B_MBdieqMe0_0),.clk(gclk));
	jdff dff_B_BfFCQTJe0_0(.din(w_dff_B_MBdieqMe0_0),.dout(w_dff_B_BfFCQTJe0_0),.clk(gclk));
	jdff dff_B_EFUNuYVk1_0(.din(w_dff_B_BfFCQTJe0_0),.dout(w_dff_B_EFUNuYVk1_0),.clk(gclk));
	jdff dff_B_yMFnqjzX7_0(.din(w_dff_B_EFUNuYVk1_0),.dout(w_dff_B_yMFnqjzX7_0),.clk(gclk));
	jdff dff_B_4T15hbcn8_0(.din(w_dff_B_yMFnqjzX7_0),.dout(w_dff_B_4T15hbcn8_0),.clk(gclk));
	jdff dff_B_AvT02vpZ9_0(.din(w_dff_B_4T15hbcn8_0),.dout(w_dff_B_AvT02vpZ9_0),.clk(gclk));
	jdff dff_B_1xIKDRRx5_0(.din(w_dff_B_AvT02vpZ9_0),.dout(w_dff_B_1xIKDRRx5_0),.clk(gclk));
	jdff dff_B_QTM9pWrH4_0(.din(w_dff_B_1xIKDRRx5_0),.dout(w_dff_B_QTM9pWrH4_0),.clk(gclk));
	jdff dff_B_IM8AeYQh7_0(.din(w_dff_B_QTM9pWrH4_0),.dout(w_dff_B_IM8AeYQh7_0),.clk(gclk));
	jdff dff_B_5owa66a82_0(.din(w_dff_B_IM8AeYQh7_0),.dout(w_dff_B_5owa66a82_0),.clk(gclk));
	jdff dff_B_m2vHSqeq3_0(.din(w_dff_B_5owa66a82_0),.dout(w_dff_B_m2vHSqeq3_0),.clk(gclk));
	jdff dff_B_UNtdUWQm7_0(.din(w_dff_B_m2vHSqeq3_0),.dout(w_dff_B_UNtdUWQm7_0),.clk(gclk));
	jdff dff_B_lIOBYjns0_0(.din(w_dff_B_UNtdUWQm7_0),.dout(w_dff_B_lIOBYjns0_0),.clk(gclk));
	jdff dff_B_2faxuY1F8_0(.din(w_dff_B_lIOBYjns0_0),.dout(w_dff_B_2faxuY1F8_0),.clk(gclk));
	jdff dff_B_PM3aSWS50_0(.din(w_dff_B_2faxuY1F8_0),.dout(w_dff_B_PM3aSWS50_0),.clk(gclk));
	jdff dff_B_Is3GgUso7_0(.din(w_dff_B_PM3aSWS50_0),.dout(w_dff_B_Is3GgUso7_0),.clk(gclk));
	jdff dff_B_4UZQvBcp9_0(.din(w_dff_B_Is3GgUso7_0),.dout(w_dff_B_4UZQvBcp9_0),.clk(gclk));
	jdff dff_B_hvYMu4RO9_0(.din(w_dff_B_4UZQvBcp9_0),.dout(w_dff_B_hvYMu4RO9_0),.clk(gclk));
	jdff dff_B_jx8JTva21_0(.din(w_dff_B_hvYMu4RO9_0),.dout(w_dff_B_jx8JTva21_0),.clk(gclk));
	jdff dff_B_h27Zusum7_0(.din(w_dff_B_jx8JTva21_0),.dout(w_dff_B_h27Zusum7_0),.clk(gclk));
	jdff dff_B_m1Zy5TGV2_0(.din(w_dff_B_h27Zusum7_0),.dout(w_dff_B_m1Zy5TGV2_0),.clk(gclk));
	jdff dff_B_ZtObcjWI4_0(.din(w_dff_B_m1Zy5TGV2_0),.dout(w_dff_B_ZtObcjWI4_0),.clk(gclk));
	jdff dff_B_5LIHS1Z84_0(.din(w_dff_B_ZtObcjWI4_0),.dout(w_dff_B_5LIHS1Z84_0),.clk(gclk));
	jdff dff_B_avFI0M5V7_0(.din(w_dff_B_5LIHS1Z84_0),.dout(w_dff_B_avFI0M5V7_0),.clk(gclk));
	jdff dff_B_9TosqZQv6_0(.din(w_dff_B_avFI0M5V7_0),.dout(w_dff_B_9TosqZQv6_0),.clk(gclk));
	jdff dff_B_dKLAarJG8_0(.din(w_dff_B_9TosqZQv6_0),.dout(w_dff_B_dKLAarJG8_0),.clk(gclk));
	jdff dff_B_IF2GADLm1_0(.din(w_dff_B_dKLAarJG8_0),.dout(w_dff_B_IF2GADLm1_0),.clk(gclk));
	jdff dff_B_7izdc4V76_0(.din(w_dff_B_IF2GADLm1_0),.dout(w_dff_B_7izdc4V76_0),.clk(gclk));
	jdff dff_B_RGkywMA92_0(.din(w_dff_B_7izdc4V76_0),.dout(w_dff_B_RGkywMA92_0),.clk(gclk));
	jdff dff_B_xjN6BYGZ6_0(.din(w_dff_B_RGkywMA92_0),.dout(w_dff_B_xjN6BYGZ6_0),.clk(gclk));
	jdff dff_B_RsrFWTXq7_0(.din(w_dff_B_xjN6BYGZ6_0),.dout(w_dff_B_RsrFWTXq7_0),.clk(gclk));
	jdff dff_B_zNMF2o3f1_0(.din(w_dff_B_RsrFWTXq7_0),.dout(w_dff_B_zNMF2o3f1_0),.clk(gclk));
	jdff dff_B_UbMj15YF7_0(.din(w_dff_B_zNMF2o3f1_0),.dout(w_dff_B_UbMj15YF7_0),.clk(gclk));
	jdff dff_B_cZ5BOPwq0_0(.din(w_dff_B_UbMj15YF7_0),.dout(w_dff_B_cZ5BOPwq0_0),.clk(gclk));
	jdff dff_B_qUsKM4NW5_0(.din(w_dff_B_cZ5BOPwq0_0),.dout(w_dff_B_qUsKM4NW5_0),.clk(gclk));
	jdff dff_B_uEIeSmiW0_0(.din(w_dff_B_qUsKM4NW5_0),.dout(w_dff_B_uEIeSmiW0_0),.clk(gclk));
	jdff dff_B_mXB4ko7Q7_0(.din(w_dff_B_uEIeSmiW0_0),.dout(w_dff_B_mXB4ko7Q7_0),.clk(gclk));
	jdff dff_B_Y5CH93RO1_0(.din(w_dff_B_mXB4ko7Q7_0),.dout(w_dff_B_Y5CH93RO1_0),.clk(gclk));
	jdff dff_B_rJlmCpRD9_0(.din(w_dff_B_Y5CH93RO1_0),.dout(w_dff_B_rJlmCpRD9_0),.clk(gclk));
	jdff dff_B_BDrkrepj7_0(.din(w_dff_B_rJlmCpRD9_0),.dout(w_dff_B_BDrkrepj7_0),.clk(gclk));
	jdff dff_B_A92dBLID0_0(.din(w_dff_B_BDrkrepj7_0),.dout(w_dff_B_A92dBLID0_0),.clk(gclk));
	jdff dff_B_Zzoca1WP0_0(.din(w_dff_B_A92dBLID0_0),.dout(w_dff_B_Zzoca1WP0_0),.clk(gclk));
	jdff dff_B_J7xGRWWQ8_0(.din(w_dff_B_Zzoca1WP0_0),.dout(w_dff_B_J7xGRWWQ8_0),.clk(gclk));
	jdff dff_B_jfthEalt2_0(.din(w_dff_B_J7xGRWWQ8_0),.dout(w_dff_B_jfthEalt2_0),.clk(gclk));
	jdff dff_B_UaJJ4Jr95_0(.din(w_dff_B_jfthEalt2_0),.dout(w_dff_B_UaJJ4Jr95_0),.clk(gclk));
	jdff dff_B_K5ygOkS13_0(.din(w_dff_B_UaJJ4Jr95_0),.dout(w_dff_B_K5ygOkS13_0),.clk(gclk));
	jdff dff_B_PN1cuHp77_0(.din(w_dff_B_K5ygOkS13_0),.dout(w_dff_B_PN1cuHp77_0),.clk(gclk));
	jdff dff_B_GejEV5Eg6_0(.din(w_dff_B_PN1cuHp77_0),.dout(w_dff_B_GejEV5Eg6_0),.clk(gclk));
	jdff dff_B_pY928UbG4_0(.din(w_dff_B_GejEV5Eg6_0),.dout(w_dff_B_pY928UbG4_0),.clk(gclk));
	jdff dff_B_vJdTy1Ut0_0(.din(w_dff_B_pY928UbG4_0),.dout(w_dff_B_vJdTy1Ut0_0),.clk(gclk));
	jdff dff_B_Yi05wNmp9_0(.din(w_dff_B_vJdTy1Ut0_0),.dout(w_dff_B_Yi05wNmp9_0),.clk(gclk));
	jdff dff_B_CJr9sUpv0_0(.din(w_dff_B_Yi05wNmp9_0),.dout(w_dff_B_CJr9sUpv0_0),.clk(gclk));
	jdff dff_B_1olkKZCp9_0(.din(w_dff_B_CJr9sUpv0_0),.dout(w_dff_B_1olkKZCp9_0),.clk(gclk));
	jdff dff_B_Yh6q8TR29_0(.din(w_dff_B_1olkKZCp9_0),.dout(w_dff_B_Yh6q8TR29_0),.clk(gclk));
	jdff dff_B_iXekFgxa6_0(.din(w_dff_B_Yh6q8TR29_0),.dout(w_dff_B_iXekFgxa6_0),.clk(gclk));
	jdff dff_B_crnV6jVU5_0(.din(w_dff_B_iXekFgxa6_0),.dout(w_dff_B_crnV6jVU5_0),.clk(gclk));
	jdff dff_B_KzHaswyh6_0(.din(w_dff_B_crnV6jVU5_0),.dout(w_dff_B_KzHaswyh6_0),.clk(gclk));
	jdff dff_B_knf8fCeI9_0(.din(w_dff_B_KzHaswyh6_0),.dout(w_dff_B_knf8fCeI9_0),.clk(gclk));
	jdff dff_B_NaGBnOLk0_0(.din(w_dff_B_knf8fCeI9_0),.dout(w_dff_B_NaGBnOLk0_0),.clk(gclk));
	jdff dff_B_jL9UKd2c2_0(.din(w_dff_B_NaGBnOLk0_0),.dout(w_dff_B_jL9UKd2c2_0),.clk(gclk));
	jdff dff_B_W3sTHeaQ4_0(.din(w_dff_B_jL9UKd2c2_0),.dout(w_dff_B_W3sTHeaQ4_0),.clk(gclk));
	jdff dff_B_smls63i15_0(.din(w_dff_B_W3sTHeaQ4_0),.dout(w_dff_B_smls63i15_0),.clk(gclk));
	jdff dff_B_rbMoLEQl6_0(.din(w_dff_B_smls63i15_0),.dout(w_dff_B_rbMoLEQl6_0),.clk(gclk));
	jdff dff_B_C6MyzLOf9_0(.din(w_dff_B_rbMoLEQl6_0),.dout(w_dff_B_C6MyzLOf9_0),.clk(gclk));
	jdff dff_B_YttT4K8E7_0(.din(w_dff_B_C6MyzLOf9_0),.dout(w_dff_B_YttT4K8E7_0),.clk(gclk));
	jdff dff_B_A8X96XcQ6_0(.din(w_dff_B_YttT4K8E7_0),.dout(w_dff_B_A8X96XcQ6_0),.clk(gclk));
	jdff dff_B_0X58FGYH0_0(.din(w_dff_B_A8X96XcQ6_0),.dout(w_dff_B_0X58FGYH0_0),.clk(gclk));
	jdff dff_B_CQz7a8gO4_0(.din(w_dff_B_0X58FGYH0_0),.dout(w_dff_B_CQz7a8gO4_0),.clk(gclk));
	jdff dff_B_zhWzqRpU0_0(.din(w_dff_B_CQz7a8gO4_0),.dout(w_dff_B_zhWzqRpU0_0),.clk(gclk));
	jdff dff_B_5sh32TL86_0(.din(w_dff_B_zhWzqRpU0_0),.dout(w_dff_B_5sh32TL86_0),.clk(gclk));
	jdff dff_B_34Xqphlm5_0(.din(w_dff_B_5sh32TL86_0),.dout(w_dff_B_34Xqphlm5_0),.clk(gclk));
	jdff dff_B_SHxPIKwg2_0(.din(w_dff_B_34Xqphlm5_0),.dout(w_dff_B_SHxPIKwg2_0),.clk(gclk));
	jdff dff_B_78ZLS5812_0(.din(w_dff_B_SHxPIKwg2_0),.dout(w_dff_B_78ZLS5812_0),.clk(gclk));
	jdff dff_B_MksQTyno0_0(.din(w_dff_B_78ZLS5812_0),.dout(w_dff_B_MksQTyno0_0),.clk(gclk));
	jdff dff_B_zdOcxGy39_0(.din(w_dff_B_MksQTyno0_0),.dout(w_dff_B_zdOcxGy39_0),.clk(gclk));
	jdff dff_B_wsW4U1dB3_0(.din(w_dff_B_zdOcxGy39_0),.dout(w_dff_B_wsW4U1dB3_0),.clk(gclk));
	jdff dff_B_w98e7xUS0_0(.din(w_dff_B_wsW4U1dB3_0),.dout(w_dff_B_w98e7xUS0_0),.clk(gclk));
	jdff dff_B_pdbfvMqH3_0(.din(w_dff_B_w98e7xUS0_0),.dout(w_dff_B_pdbfvMqH3_0),.clk(gclk));
	jdff dff_B_5cks2KkI7_0(.din(w_dff_B_pdbfvMqH3_0),.dout(w_dff_B_5cks2KkI7_0),.clk(gclk));
	jdff dff_B_7sd8C4268_0(.din(w_dff_B_5cks2KkI7_0),.dout(w_dff_B_7sd8C4268_0),.clk(gclk));
	jdff dff_B_sfEETGGb8_0(.din(w_dff_B_7sd8C4268_0),.dout(w_dff_B_sfEETGGb8_0),.clk(gclk));
	jdff dff_B_pVwxEO8f4_0(.din(w_dff_B_sfEETGGb8_0),.dout(w_dff_B_pVwxEO8f4_0),.clk(gclk));
	jdff dff_B_Ob5xSnvX8_0(.din(w_dff_B_pVwxEO8f4_0),.dout(w_dff_B_Ob5xSnvX8_0),.clk(gclk));
	jdff dff_B_9a0vFLUn0_0(.din(w_dff_B_Ob5xSnvX8_0),.dout(w_dff_B_9a0vFLUn0_0),.clk(gclk));
	jdff dff_B_S9GyfjEX9_0(.din(w_dff_B_9a0vFLUn0_0),.dout(w_dff_B_S9GyfjEX9_0),.clk(gclk));
	jdff dff_B_qiQhmBhK7_0(.din(w_dff_B_S9GyfjEX9_0),.dout(w_dff_B_qiQhmBhK7_0),.clk(gclk));
	jdff dff_B_zfZaybuE0_0(.din(w_dff_B_qiQhmBhK7_0),.dout(w_dff_B_zfZaybuE0_0),.clk(gclk));
	jdff dff_B_R8gm21p73_0(.din(w_dff_B_zfZaybuE0_0),.dout(w_dff_B_R8gm21p73_0),.clk(gclk));
	jdff dff_B_X1oxPpZf6_0(.din(w_dff_B_R8gm21p73_0),.dout(w_dff_B_X1oxPpZf6_0),.clk(gclk));
	jdff dff_B_lxbb6iv81_0(.din(w_dff_B_X1oxPpZf6_0),.dout(w_dff_B_lxbb6iv81_0),.clk(gclk));
	jdff dff_B_5r1rrR6p3_0(.din(w_dff_B_lxbb6iv81_0),.dout(w_dff_B_5r1rrR6p3_0),.clk(gclk));
	jdff dff_B_3XsPByS46_0(.din(w_dff_B_5r1rrR6p3_0),.dout(w_dff_B_3XsPByS46_0),.clk(gclk));
	jdff dff_B_5h5pEzoJ1_1(.din(n954),.dout(w_dff_B_5h5pEzoJ1_1),.clk(gclk));
	jdff dff_B_TW22cvRH5_1(.din(w_dff_B_5h5pEzoJ1_1),.dout(w_dff_B_TW22cvRH5_1),.clk(gclk));
	jdff dff_B_34SK0ARe2_1(.din(w_dff_B_TW22cvRH5_1),.dout(w_dff_B_34SK0ARe2_1),.clk(gclk));
	jdff dff_B_J7p5oi1M9_1(.din(w_dff_B_34SK0ARe2_1),.dout(w_dff_B_J7p5oi1M9_1),.clk(gclk));
	jdff dff_B_GHZwEY2s1_1(.din(w_dff_B_J7p5oi1M9_1),.dout(w_dff_B_GHZwEY2s1_1),.clk(gclk));
	jdff dff_B_g2jdiwii1_1(.din(w_dff_B_GHZwEY2s1_1),.dout(w_dff_B_g2jdiwii1_1),.clk(gclk));
	jdff dff_B_svz0r1ll2_1(.din(w_dff_B_g2jdiwii1_1),.dout(w_dff_B_svz0r1ll2_1),.clk(gclk));
	jdff dff_B_s4S94kZ96_1(.din(w_dff_B_svz0r1ll2_1),.dout(w_dff_B_s4S94kZ96_1),.clk(gclk));
	jdff dff_B_f7AWNVNL8_1(.din(w_dff_B_s4S94kZ96_1),.dout(w_dff_B_f7AWNVNL8_1),.clk(gclk));
	jdff dff_B_tfsKzCkX8_1(.din(w_dff_B_f7AWNVNL8_1),.dout(w_dff_B_tfsKzCkX8_1),.clk(gclk));
	jdff dff_B_1EsPREt61_1(.din(w_dff_B_tfsKzCkX8_1),.dout(w_dff_B_1EsPREt61_1),.clk(gclk));
	jdff dff_B_sEmo0SZx6_1(.din(w_dff_B_1EsPREt61_1),.dout(w_dff_B_sEmo0SZx6_1),.clk(gclk));
	jdff dff_B_fZEKeNit1_1(.din(w_dff_B_sEmo0SZx6_1),.dout(w_dff_B_fZEKeNit1_1),.clk(gclk));
	jdff dff_B_1xevbUJr4_1(.din(w_dff_B_fZEKeNit1_1),.dout(w_dff_B_1xevbUJr4_1),.clk(gclk));
	jdff dff_B_k0KJEXRo3_1(.din(w_dff_B_1xevbUJr4_1),.dout(w_dff_B_k0KJEXRo3_1),.clk(gclk));
	jdff dff_B_KGEILHza1_1(.din(w_dff_B_k0KJEXRo3_1),.dout(w_dff_B_KGEILHza1_1),.clk(gclk));
	jdff dff_B_FfVwj9YX7_1(.din(w_dff_B_KGEILHza1_1),.dout(w_dff_B_FfVwj9YX7_1),.clk(gclk));
	jdff dff_B_3ASk24GQ2_1(.din(w_dff_B_FfVwj9YX7_1),.dout(w_dff_B_3ASk24GQ2_1),.clk(gclk));
	jdff dff_B_NlwZVyxn1_1(.din(w_dff_B_3ASk24GQ2_1),.dout(w_dff_B_NlwZVyxn1_1),.clk(gclk));
	jdff dff_B_7pbXjwHD1_1(.din(w_dff_B_NlwZVyxn1_1),.dout(w_dff_B_7pbXjwHD1_1),.clk(gclk));
	jdff dff_B_Gg6UT4Z16_1(.din(w_dff_B_7pbXjwHD1_1),.dout(w_dff_B_Gg6UT4Z16_1),.clk(gclk));
	jdff dff_B_aa0nRbpH3_1(.din(w_dff_B_Gg6UT4Z16_1),.dout(w_dff_B_aa0nRbpH3_1),.clk(gclk));
	jdff dff_B_0InrlveO2_1(.din(w_dff_B_aa0nRbpH3_1),.dout(w_dff_B_0InrlveO2_1),.clk(gclk));
	jdff dff_B_1WjlFOcE2_1(.din(w_dff_B_0InrlveO2_1),.dout(w_dff_B_1WjlFOcE2_1),.clk(gclk));
	jdff dff_B_S8jNN0zf1_1(.din(w_dff_B_1WjlFOcE2_1),.dout(w_dff_B_S8jNN0zf1_1),.clk(gclk));
	jdff dff_B_SuZBlx139_1(.din(w_dff_B_S8jNN0zf1_1),.dout(w_dff_B_SuZBlx139_1),.clk(gclk));
	jdff dff_B_3AMKNiPJ1_1(.din(w_dff_B_SuZBlx139_1),.dout(w_dff_B_3AMKNiPJ1_1),.clk(gclk));
	jdff dff_B_jUzV742W3_1(.din(w_dff_B_3AMKNiPJ1_1),.dout(w_dff_B_jUzV742W3_1),.clk(gclk));
	jdff dff_B_FNbz4A4v3_1(.din(w_dff_B_jUzV742W3_1),.dout(w_dff_B_FNbz4A4v3_1),.clk(gclk));
	jdff dff_B_ec8KbeNC6_1(.din(w_dff_B_FNbz4A4v3_1),.dout(w_dff_B_ec8KbeNC6_1),.clk(gclk));
	jdff dff_B_LUTxwJ8h0_1(.din(w_dff_B_ec8KbeNC6_1),.dout(w_dff_B_LUTxwJ8h0_1),.clk(gclk));
	jdff dff_B_CahfPJlh5_1(.din(w_dff_B_LUTxwJ8h0_1),.dout(w_dff_B_CahfPJlh5_1),.clk(gclk));
	jdff dff_B_lx8D4W2E5_1(.din(w_dff_B_CahfPJlh5_1),.dout(w_dff_B_lx8D4W2E5_1),.clk(gclk));
	jdff dff_B_qbMiveIy7_1(.din(w_dff_B_lx8D4W2E5_1),.dout(w_dff_B_qbMiveIy7_1),.clk(gclk));
	jdff dff_B_dwX66ODU5_1(.din(w_dff_B_qbMiveIy7_1),.dout(w_dff_B_dwX66ODU5_1),.clk(gclk));
	jdff dff_B_hb4NwXxJ8_1(.din(w_dff_B_dwX66ODU5_1),.dout(w_dff_B_hb4NwXxJ8_1),.clk(gclk));
	jdff dff_B_pLZg3z3p0_1(.din(w_dff_B_hb4NwXxJ8_1),.dout(w_dff_B_pLZg3z3p0_1),.clk(gclk));
	jdff dff_B_GF7WkCUh3_1(.din(w_dff_B_pLZg3z3p0_1),.dout(w_dff_B_GF7WkCUh3_1),.clk(gclk));
	jdff dff_B_lBmk3FQv6_1(.din(w_dff_B_GF7WkCUh3_1),.dout(w_dff_B_lBmk3FQv6_1),.clk(gclk));
	jdff dff_B_rJkdbwcB7_1(.din(w_dff_B_lBmk3FQv6_1),.dout(w_dff_B_rJkdbwcB7_1),.clk(gclk));
	jdff dff_B_pjohpkrt4_1(.din(w_dff_B_rJkdbwcB7_1),.dout(w_dff_B_pjohpkrt4_1),.clk(gclk));
	jdff dff_B_iwgyciuB1_1(.din(w_dff_B_pjohpkrt4_1),.dout(w_dff_B_iwgyciuB1_1),.clk(gclk));
	jdff dff_B_GO4a9lSi5_1(.din(w_dff_B_iwgyciuB1_1),.dout(w_dff_B_GO4a9lSi5_1),.clk(gclk));
	jdff dff_B_WSA9MvCL1_1(.din(w_dff_B_GO4a9lSi5_1),.dout(w_dff_B_WSA9MvCL1_1),.clk(gclk));
	jdff dff_B_kL7HkD6D4_1(.din(w_dff_B_WSA9MvCL1_1),.dout(w_dff_B_kL7HkD6D4_1),.clk(gclk));
	jdff dff_B_EioNTpVY9_1(.din(w_dff_B_kL7HkD6D4_1),.dout(w_dff_B_EioNTpVY9_1),.clk(gclk));
	jdff dff_B_LNBmf1Xn8_1(.din(w_dff_B_EioNTpVY9_1),.dout(w_dff_B_LNBmf1Xn8_1),.clk(gclk));
	jdff dff_B_d9FZL5962_1(.din(w_dff_B_LNBmf1Xn8_1),.dout(w_dff_B_d9FZL5962_1),.clk(gclk));
	jdff dff_B_RWQrh6mq0_1(.din(w_dff_B_d9FZL5962_1),.dout(w_dff_B_RWQrh6mq0_1),.clk(gclk));
	jdff dff_B_9XaHFRwg9_1(.din(w_dff_B_RWQrh6mq0_1),.dout(w_dff_B_9XaHFRwg9_1),.clk(gclk));
	jdff dff_B_xxKQ4Ia91_1(.din(w_dff_B_9XaHFRwg9_1),.dout(w_dff_B_xxKQ4Ia91_1),.clk(gclk));
	jdff dff_B_qCh9Ijb56_1(.din(w_dff_B_xxKQ4Ia91_1),.dout(w_dff_B_qCh9Ijb56_1),.clk(gclk));
	jdff dff_B_m1QcDzfL5_1(.din(w_dff_B_qCh9Ijb56_1),.dout(w_dff_B_m1QcDzfL5_1),.clk(gclk));
	jdff dff_B_UvLUOwdL7_1(.din(w_dff_B_m1QcDzfL5_1),.dout(w_dff_B_UvLUOwdL7_1),.clk(gclk));
	jdff dff_B_af2ln9mi4_1(.din(w_dff_B_UvLUOwdL7_1),.dout(w_dff_B_af2ln9mi4_1),.clk(gclk));
	jdff dff_B_2l1X0JWa3_1(.din(w_dff_B_af2ln9mi4_1),.dout(w_dff_B_2l1X0JWa3_1),.clk(gclk));
	jdff dff_B_azVg8IOu7_1(.din(w_dff_B_2l1X0JWa3_1),.dout(w_dff_B_azVg8IOu7_1),.clk(gclk));
	jdff dff_B_h6ukKkiD4_1(.din(w_dff_B_azVg8IOu7_1),.dout(w_dff_B_h6ukKkiD4_1),.clk(gclk));
	jdff dff_B_c1aLeOMc0_1(.din(w_dff_B_h6ukKkiD4_1),.dout(w_dff_B_c1aLeOMc0_1),.clk(gclk));
	jdff dff_B_Z2zhRQzZ5_1(.din(w_dff_B_c1aLeOMc0_1),.dout(w_dff_B_Z2zhRQzZ5_1),.clk(gclk));
	jdff dff_B_Z2l5jexn7_1(.din(w_dff_B_Z2zhRQzZ5_1),.dout(w_dff_B_Z2l5jexn7_1),.clk(gclk));
	jdff dff_B_PQjUwcbL3_1(.din(w_dff_B_Z2l5jexn7_1),.dout(w_dff_B_PQjUwcbL3_1),.clk(gclk));
	jdff dff_B_K8NNNrRb2_1(.din(w_dff_B_PQjUwcbL3_1),.dout(w_dff_B_K8NNNrRb2_1),.clk(gclk));
	jdff dff_B_R3hbC0lI4_1(.din(w_dff_B_K8NNNrRb2_1),.dout(w_dff_B_R3hbC0lI4_1),.clk(gclk));
	jdff dff_B_kBZLhqis3_1(.din(w_dff_B_R3hbC0lI4_1),.dout(w_dff_B_kBZLhqis3_1),.clk(gclk));
	jdff dff_B_pBhMXUKh1_1(.din(w_dff_B_kBZLhqis3_1),.dout(w_dff_B_pBhMXUKh1_1),.clk(gclk));
	jdff dff_B_vodXbVJ26_1(.din(w_dff_B_pBhMXUKh1_1),.dout(w_dff_B_vodXbVJ26_1),.clk(gclk));
	jdff dff_B_EDTYywnX5_1(.din(w_dff_B_vodXbVJ26_1),.dout(w_dff_B_EDTYywnX5_1),.clk(gclk));
	jdff dff_B_Ci0YArzd4_1(.din(w_dff_B_EDTYywnX5_1),.dout(w_dff_B_Ci0YArzd4_1),.clk(gclk));
	jdff dff_B_4j9UoHSZ4_1(.din(w_dff_B_Ci0YArzd4_1),.dout(w_dff_B_4j9UoHSZ4_1),.clk(gclk));
	jdff dff_B_l9QuPTnE5_1(.din(w_dff_B_4j9UoHSZ4_1),.dout(w_dff_B_l9QuPTnE5_1),.clk(gclk));
	jdff dff_B_IdMkGcYU3_1(.din(w_dff_B_l9QuPTnE5_1),.dout(w_dff_B_IdMkGcYU3_1),.clk(gclk));
	jdff dff_B_oaAdyzia2_1(.din(w_dff_B_IdMkGcYU3_1),.dout(w_dff_B_oaAdyzia2_1),.clk(gclk));
	jdff dff_B_AKnU10zy5_1(.din(w_dff_B_oaAdyzia2_1),.dout(w_dff_B_AKnU10zy5_1),.clk(gclk));
	jdff dff_B_hK7GLm3G0_1(.din(w_dff_B_AKnU10zy5_1),.dout(w_dff_B_hK7GLm3G0_1),.clk(gclk));
	jdff dff_B_4EnP114U3_1(.din(w_dff_B_hK7GLm3G0_1),.dout(w_dff_B_4EnP114U3_1),.clk(gclk));
	jdff dff_B_htkj9dM24_1(.din(w_dff_B_4EnP114U3_1),.dout(w_dff_B_htkj9dM24_1),.clk(gclk));
	jdff dff_B_VuImE7Zp1_1(.din(w_dff_B_htkj9dM24_1),.dout(w_dff_B_VuImE7Zp1_1),.clk(gclk));
	jdff dff_B_V79VZpFO3_1(.din(w_dff_B_VuImE7Zp1_1),.dout(w_dff_B_V79VZpFO3_1),.clk(gclk));
	jdff dff_B_O1HARNWQ3_1(.din(w_dff_B_V79VZpFO3_1),.dout(w_dff_B_O1HARNWQ3_1),.clk(gclk));
	jdff dff_B_Z2mbYRCK4_1(.din(w_dff_B_O1HARNWQ3_1),.dout(w_dff_B_Z2mbYRCK4_1),.clk(gclk));
	jdff dff_B_aKjDdA3e7_1(.din(w_dff_B_Z2mbYRCK4_1),.dout(w_dff_B_aKjDdA3e7_1),.clk(gclk));
	jdff dff_B_e8ZoBi5d2_1(.din(w_dff_B_aKjDdA3e7_1),.dout(w_dff_B_e8ZoBi5d2_1),.clk(gclk));
	jdff dff_B_mRoO8x6R9_1(.din(w_dff_B_e8ZoBi5d2_1),.dout(w_dff_B_mRoO8x6R9_1),.clk(gclk));
	jdff dff_B_fIOfh2wh3_1(.din(w_dff_B_mRoO8x6R9_1),.dout(w_dff_B_fIOfh2wh3_1),.clk(gclk));
	jdff dff_B_kR8LnsSr2_1(.din(w_dff_B_fIOfh2wh3_1),.dout(w_dff_B_kR8LnsSr2_1),.clk(gclk));
	jdff dff_B_W13wPvvM4_1(.din(w_dff_B_kR8LnsSr2_1),.dout(w_dff_B_W13wPvvM4_1),.clk(gclk));
	jdff dff_B_HNZ5Rhd77_1(.din(w_dff_B_W13wPvvM4_1),.dout(w_dff_B_HNZ5Rhd77_1),.clk(gclk));
	jdff dff_B_AeohlU5a3_1(.din(w_dff_B_HNZ5Rhd77_1),.dout(w_dff_B_AeohlU5a3_1),.clk(gclk));
	jdff dff_B_Rugfoc3L6_1(.din(w_dff_B_AeohlU5a3_1),.dout(w_dff_B_Rugfoc3L6_1),.clk(gclk));
	jdff dff_B_FndFkS8U0_1(.din(w_dff_B_Rugfoc3L6_1),.dout(w_dff_B_FndFkS8U0_1),.clk(gclk));
	jdff dff_B_6tvLxXyI9_1(.din(w_dff_B_FndFkS8U0_1),.dout(w_dff_B_6tvLxXyI9_1),.clk(gclk));
	jdff dff_B_l2Y8TxU44_1(.din(w_dff_B_6tvLxXyI9_1),.dout(w_dff_B_l2Y8TxU44_1),.clk(gclk));
	jdff dff_B_fqdrpVbN6_1(.din(w_dff_B_l2Y8TxU44_1),.dout(w_dff_B_fqdrpVbN6_1),.clk(gclk));
	jdff dff_B_Jf6mJkjd5_1(.din(w_dff_B_fqdrpVbN6_1),.dout(w_dff_B_Jf6mJkjd5_1),.clk(gclk));
	jdff dff_B_i8hjuhlu9_0(.din(n955),.dout(w_dff_B_i8hjuhlu9_0),.clk(gclk));
	jdff dff_B_76ubyzjk6_0(.din(w_dff_B_i8hjuhlu9_0),.dout(w_dff_B_76ubyzjk6_0),.clk(gclk));
	jdff dff_B_2JUcnE6Z6_0(.din(w_dff_B_76ubyzjk6_0),.dout(w_dff_B_2JUcnE6Z6_0),.clk(gclk));
	jdff dff_B_5kkV5XQC7_0(.din(w_dff_B_2JUcnE6Z6_0),.dout(w_dff_B_5kkV5XQC7_0),.clk(gclk));
	jdff dff_B_aSytXVeC2_0(.din(w_dff_B_5kkV5XQC7_0),.dout(w_dff_B_aSytXVeC2_0),.clk(gclk));
	jdff dff_B_QJPEGd597_0(.din(w_dff_B_aSytXVeC2_0),.dout(w_dff_B_QJPEGd597_0),.clk(gclk));
	jdff dff_B_5vittjnS2_0(.din(w_dff_B_QJPEGd597_0),.dout(w_dff_B_5vittjnS2_0),.clk(gclk));
	jdff dff_B_PR9goVpm3_0(.din(w_dff_B_5vittjnS2_0),.dout(w_dff_B_PR9goVpm3_0),.clk(gclk));
	jdff dff_B_RP3oI6Nd4_0(.din(w_dff_B_PR9goVpm3_0),.dout(w_dff_B_RP3oI6Nd4_0),.clk(gclk));
	jdff dff_B_VLf54wtn9_0(.din(w_dff_B_RP3oI6Nd4_0),.dout(w_dff_B_VLf54wtn9_0),.clk(gclk));
	jdff dff_B_pzfAHvHI0_0(.din(w_dff_B_VLf54wtn9_0),.dout(w_dff_B_pzfAHvHI0_0),.clk(gclk));
	jdff dff_B_ceaM2JMS6_0(.din(w_dff_B_pzfAHvHI0_0),.dout(w_dff_B_ceaM2JMS6_0),.clk(gclk));
	jdff dff_B_hXAQVowD9_0(.din(w_dff_B_ceaM2JMS6_0),.dout(w_dff_B_hXAQVowD9_0),.clk(gclk));
	jdff dff_B_qEQVx2xH9_0(.din(w_dff_B_hXAQVowD9_0),.dout(w_dff_B_qEQVx2xH9_0),.clk(gclk));
	jdff dff_B_MuLgi9Fk0_0(.din(w_dff_B_qEQVx2xH9_0),.dout(w_dff_B_MuLgi9Fk0_0),.clk(gclk));
	jdff dff_B_xbaeqHf26_0(.din(w_dff_B_MuLgi9Fk0_0),.dout(w_dff_B_xbaeqHf26_0),.clk(gclk));
	jdff dff_B_WvpMQQrw0_0(.din(w_dff_B_xbaeqHf26_0),.dout(w_dff_B_WvpMQQrw0_0),.clk(gclk));
	jdff dff_B_NaE259Mg0_0(.din(w_dff_B_WvpMQQrw0_0),.dout(w_dff_B_NaE259Mg0_0),.clk(gclk));
	jdff dff_B_GA25x1Px6_0(.din(w_dff_B_NaE259Mg0_0),.dout(w_dff_B_GA25x1Px6_0),.clk(gclk));
	jdff dff_B_71eXY0lQ7_0(.din(w_dff_B_GA25x1Px6_0),.dout(w_dff_B_71eXY0lQ7_0),.clk(gclk));
	jdff dff_B_JbEUF7ot4_0(.din(w_dff_B_71eXY0lQ7_0),.dout(w_dff_B_JbEUF7ot4_0),.clk(gclk));
	jdff dff_B_Umb7swJJ7_0(.din(w_dff_B_JbEUF7ot4_0),.dout(w_dff_B_Umb7swJJ7_0),.clk(gclk));
	jdff dff_B_FnUuINN84_0(.din(w_dff_B_Umb7swJJ7_0),.dout(w_dff_B_FnUuINN84_0),.clk(gclk));
	jdff dff_B_Uu3FwLVp4_0(.din(w_dff_B_FnUuINN84_0),.dout(w_dff_B_Uu3FwLVp4_0),.clk(gclk));
	jdff dff_B_AHExV0Qf9_0(.din(w_dff_B_Uu3FwLVp4_0),.dout(w_dff_B_AHExV0Qf9_0),.clk(gclk));
	jdff dff_B_7VMRMB8y0_0(.din(w_dff_B_AHExV0Qf9_0),.dout(w_dff_B_7VMRMB8y0_0),.clk(gclk));
	jdff dff_B_CDaOiJ8J3_0(.din(w_dff_B_7VMRMB8y0_0),.dout(w_dff_B_CDaOiJ8J3_0),.clk(gclk));
	jdff dff_B_iXaF2lDd6_0(.din(w_dff_B_CDaOiJ8J3_0),.dout(w_dff_B_iXaF2lDd6_0),.clk(gclk));
	jdff dff_B_qtMibAbp3_0(.din(w_dff_B_iXaF2lDd6_0),.dout(w_dff_B_qtMibAbp3_0),.clk(gclk));
	jdff dff_B_xAxUj8Os9_0(.din(w_dff_B_qtMibAbp3_0),.dout(w_dff_B_xAxUj8Os9_0),.clk(gclk));
	jdff dff_B_VFQ2YYTI0_0(.din(w_dff_B_xAxUj8Os9_0),.dout(w_dff_B_VFQ2YYTI0_0),.clk(gclk));
	jdff dff_B_B1jgPaIN5_0(.din(w_dff_B_VFQ2YYTI0_0),.dout(w_dff_B_B1jgPaIN5_0),.clk(gclk));
	jdff dff_B_L5f7ZURS5_0(.din(w_dff_B_B1jgPaIN5_0),.dout(w_dff_B_L5f7ZURS5_0),.clk(gclk));
	jdff dff_B_DaGiZrT46_0(.din(w_dff_B_L5f7ZURS5_0),.dout(w_dff_B_DaGiZrT46_0),.clk(gclk));
	jdff dff_B_nJ4Ku9xO9_0(.din(w_dff_B_DaGiZrT46_0),.dout(w_dff_B_nJ4Ku9xO9_0),.clk(gclk));
	jdff dff_B_w0F39Ppm7_0(.din(w_dff_B_nJ4Ku9xO9_0),.dout(w_dff_B_w0F39Ppm7_0),.clk(gclk));
	jdff dff_B_yu8tBKAE9_0(.din(w_dff_B_w0F39Ppm7_0),.dout(w_dff_B_yu8tBKAE9_0),.clk(gclk));
	jdff dff_B_CjkOfixa4_0(.din(w_dff_B_yu8tBKAE9_0),.dout(w_dff_B_CjkOfixa4_0),.clk(gclk));
	jdff dff_B_S90VgQyU2_0(.din(w_dff_B_CjkOfixa4_0),.dout(w_dff_B_S90VgQyU2_0),.clk(gclk));
	jdff dff_B_eDsKeAmE1_0(.din(w_dff_B_S90VgQyU2_0),.dout(w_dff_B_eDsKeAmE1_0),.clk(gclk));
	jdff dff_B_haItXVPK8_0(.din(w_dff_B_eDsKeAmE1_0),.dout(w_dff_B_haItXVPK8_0),.clk(gclk));
	jdff dff_B_VgwNIEZi6_0(.din(w_dff_B_haItXVPK8_0),.dout(w_dff_B_VgwNIEZi6_0),.clk(gclk));
	jdff dff_B_ezp1duFy8_0(.din(w_dff_B_VgwNIEZi6_0),.dout(w_dff_B_ezp1duFy8_0),.clk(gclk));
	jdff dff_B_1zbwQ8W52_0(.din(w_dff_B_ezp1duFy8_0),.dout(w_dff_B_1zbwQ8W52_0),.clk(gclk));
	jdff dff_B_FWRkZ8sw0_0(.din(w_dff_B_1zbwQ8W52_0),.dout(w_dff_B_FWRkZ8sw0_0),.clk(gclk));
	jdff dff_B_6UqfWH3R3_0(.din(w_dff_B_FWRkZ8sw0_0),.dout(w_dff_B_6UqfWH3R3_0),.clk(gclk));
	jdff dff_B_6V0miGFq3_0(.din(w_dff_B_6UqfWH3R3_0),.dout(w_dff_B_6V0miGFq3_0),.clk(gclk));
	jdff dff_B_6r4CoxRh4_0(.din(w_dff_B_6V0miGFq3_0),.dout(w_dff_B_6r4CoxRh4_0),.clk(gclk));
	jdff dff_B_GwnGBeS01_0(.din(w_dff_B_6r4CoxRh4_0),.dout(w_dff_B_GwnGBeS01_0),.clk(gclk));
	jdff dff_B_lemZ41vD2_0(.din(w_dff_B_GwnGBeS01_0),.dout(w_dff_B_lemZ41vD2_0),.clk(gclk));
	jdff dff_B_SM5vYIv53_0(.din(w_dff_B_lemZ41vD2_0),.dout(w_dff_B_SM5vYIv53_0),.clk(gclk));
	jdff dff_B_iYKu0jZI7_0(.din(w_dff_B_SM5vYIv53_0),.dout(w_dff_B_iYKu0jZI7_0),.clk(gclk));
	jdff dff_B_xWCNrAXh6_0(.din(w_dff_B_iYKu0jZI7_0),.dout(w_dff_B_xWCNrAXh6_0),.clk(gclk));
	jdff dff_B_THDKSGDB9_0(.din(w_dff_B_xWCNrAXh6_0),.dout(w_dff_B_THDKSGDB9_0),.clk(gclk));
	jdff dff_B_zJsyjVAl8_0(.din(w_dff_B_THDKSGDB9_0),.dout(w_dff_B_zJsyjVAl8_0),.clk(gclk));
	jdff dff_B_UoGT25TO7_0(.din(w_dff_B_zJsyjVAl8_0),.dout(w_dff_B_UoGT25TO7_0),.clk(gclk));
	jdff dff_B_3BTz2QOv8_0(.din(w_dff_B_UoGT25TO7_0),.dout(w_dff_B_3BTz2QOv8_0),.clk(gclk));
	jdff dff_B_d8DVl0Zv9_0(.din(w_dff_B_3BTz2QOv8_0),.dout(w_dff_B_d8DVl0Zv9_0),.clk(gclk));
	jdff dff_B_ghMBkZe21_0(.din(w_dff_B_d8DVl0Zv9_0),.dout(w_dff_B_ghMBkZe21_0),.clk(gclk));
	jdff dff_B_irOuD0Bm1_0(.din(w_dff_B_ghMBkZe21_0),.dout(w_dff_B_irOuD0Bm1_0),.clk(gclk));
	jdff dff_B_lgET5Av46_0(.din(w_dff_B_irOuD0Bm1_0),.dout(w_dff_B_lgET5Av46_0),.clk(gclk));
	jdff dff_B_aK22A6Ah9_0(.din(w_dff_B_lgET5Av46_0),.dout(w_dff_B_aK22A6Ah9_0),.clk(gclk));
	jdff dff_B_xhbP446k1_0(.din(w_dff_B_aK22A6Ah9_0),.dout(w_dff_B_xhbP446k1_0),.clk(gclk));
	jdff dff_B_b8voxjEf1_0(.din(w_dff_B_xhbP446k1_0),.dout(w_dff_B_b8voxjEf1_0),.clk(gclk));
	jdff dff_B_WYhARzM81_0(.din(w_dff_B_b8voxjEf1_0),.dout(w_dff_B_WYhARzM81_0),.clk(gclk));
	jdff dff_B_kFiFUhd77_0(.din(w_dff_B_WYhARzM81_0),.dout(w_dff_B_kFiFUhd77_0),.clk(gclk));
	jdff dff_B_im71HWpd0_0(.din(w_dff_B_kFiFUhd77_0),.dout(w_dff_B_im71HWpd0_0),.clk(gclk));
	jdff dff_B_g2Gqysx42_0(.din(w_dff_B_im71HWpd0_0),.dout(w_dff_B_g2Gqysx42_0),.clk(gclk));
	jdff dff_B_cgxSuDDf5_0(.din(w_dff_B_g2Gqysx42_0),.dout(w_dff_B_cgxSuDDf5_0),.clk(gclk));
	jdff dff_B_MlQT6Hfu7_0(.din(w_dff_B_cgxSuDDf5_0),.dout(w_dff_B_MlQT6Hfu7_0),.clk(gclk));
	jdff dff_B_HjqrmXjg3_0(.din(w_dff_B_MlQT6Hfu7_0),.dout(w_dff_B_HjqrmXjg3_0),.clk(gclk));
	jdff dff_B_sGzGMXpn6_0(.din(w_dff_B_HjqrmXjg3_0),.dout(w_dff_B_sGzGMXpn6_0),.clk(gclk));
	jdff dff_B_wRIOv2bx6_0(.din(w_dff_B_sGzGMXpn6_0),.dout(w_dff_B_wRIOv2bx6_0),.clk(gclk));
	jdff dff_B_DaHKbmqu1_0(.din(w_dff_B_wRIOv2bx6_0),.dout(w_dff_B_DaHKbmqu1_0),.clk(gclk));
	jdff dff_B_x1fxOtZK0_0(.din(w_dff_B_DaHKbmqu1_0),.dout(w_dff_B_x1fxOtZK0_0),.clk(gclk));
	jdff dff_B_65OhVyop0_0(.din(w_dff_B_x1fxOtZK0_0),.dout(w_dff_B_65OhVyop0_0),.clk(gclk));
	jdff dff_B_aYKMZH9H4_0(.din(w_dff_B_65OhVyop0_0),.dout(w_dff_B_aYKMZH9H4_0),.clk(gclk));
	jdff dff_B_sW0rXPWk3_0(.din(w_dff_B_aYKMZH9H4_0),.dout(w_dff_B_sW0rXPWk3_0),.clk(gclk));
	jdff dff_B_lZ9HvCBD6_0(.din(w_dff_B_sW0rXPWk3_0),.dout(w_dff_B_lZ9HvCBD6_0),.clk(gclk));
	jdff dff_B_vkmjfrXb3_0(.din(w_dff_B_lZ9HvCBD6_0),.dout(w_dff_B_vkmjfrXb3_0),.clk(gclk));
	jdff dff_B_2xHZtOgN5_0(.din(w_dff_B_vkmjfrXb3_0),.dout(w_dff_B_2xHZtOgN5_0),.clk(gclk));
	jdff dff_B_qluoOv0f5_0(.din(w_dff_B_2xHZtOgN5_0),.dout(w_dff_B_qluoOv0f5_0),.clk(gclk));
	jdff dff_B_bQ5oZYPx1_0(.din(w_dff_B_qluoOv0f5_0),.dout(w_dff_B_bQ5oZYPx1_0),.clk(gclk));
	jdff dff_B_CSdErt2L5_0(.din(w_dff_B_bQ5oZYPx1_0),.dout(w_dff_B_CSdErt2L5_0),.clk(gclk));
	jdff dff_B_w4uv4KX34_0(.din(w_dff_B_CSdErt2L5_0),.dout(w_dff_B_w4uv4KX34_0),.clk(gclk));
	jdff dff_B_DrNNixjE3_0(.din(w_dff_B_w4uv4KX34_0),.dout(w_dff_B_DrNNixjE3_0),.clk(gclk));
	jdff dff_B_GsquZjmj7_0(.din(w_dff_B_DrNNixjE3_0),.dout(w_dff_B_GsquZjmj7_0),.clk(gclk));
	jdff dff_B_JLDbsI091_0(.din(w_dff_B_GsquZjmj7_0),.dout(w_dff_B_JLDbsI091_0),.clk(gclk));
	jdff dff_B_laECUqgj7_0(.din(w_dff_B_JLDbsI091_0),.dout(w_dff_B_laECUqgj7_0),.clk(gclk));
	jdff dff_B_h80dNyXL3_0(.din(w_dff_B_laECUqgj7_0),.dout(w_dff_B_h80dNyXL3_0),.clk(gclk));
	jdff dff_B_vfu81PqA8_0(.din(w_dff_B_h80dNyXL3_0),.dout(w_dff_B_vfu81PqA8_0),.clk(gclk));
	jdff dff_B_JqtnApUX2_0(.din(w_dff_B_vfu81PqA8_0),.dout(w_dff_B_JqtnApUX2_0),.clk(gclk));
	jdff dff_B_7QfGz7AH0_0(.din(w_dff_B_JqtnApUX2_0),.dout(w_dff_B_7QfGz7AH0_0),.clk(gclk));
	jdff dff_B_l5iuMxeB6_0(.din(w_dff_B_7QfGz7AH0_0),.dout(w_dff_B_l5iuMxeB6_0),.clk(gclk));
	jdff dff_B_gF4cW8n67_0(.din(w_dff_B_l5iuMxeB6_0),.dout(w_dff_B_gF4cW8n67_0),.clk(gclk));
	jdff dff_B_V4Id4OKl3_1(.din(n948),.dout(w_dff_B_V4Id4OKl3_1),.clk(gclk));
	jdff dff_B_FUwoILhq4_1(.din(w_dff_B_V4Id4OKl3_1),.dout(w_dff_B_FUwoILhq4_1),.clk(gclk));
	jdff dff_B_gOmB6Gj76_1(.din(w_dff_B_FUwoILhq4_1),.dout(w_dff_B_gOmB6Gj76_1),.clk(gclk));
	jdff dff_B_jqRGrULa6_1(.din(w_dff_B_gOmB6Gj76_1),.dout(w_dff_B_jqRGrULa6_1),.clk(gclk));
	jdff dff_B_W8txnoBr5_1(.din(w_dff_B_jqRGrULa6_1),.dout(w_dff_B_W8txnoBr5_1),.clk(gclk));
	jdff dff_B_ak6byy5r4_1(.din(w_dff_B_W8txnoBr5_1),.dout(w_dff_B_ak6byy5r4_1),.clk(gclk));
	jdff dff_B_PXvfUu7z8_1(.din(w_dff_B_ak6byy5r4_1),.dout(w_dff_B_PXvfUu7z8_1),.clk(gclk));
	jdff dff_B_JM3H6XI40_1(.din(w_dff_B_PXvfUu7z8_1),.dout(w_dff_B_JM3H6XI40_1),.clk(gclk));
	jdff dff_B_VVtGThzh2_1(.din(w_dff_B_JM3H6XI40_1),.dout(w_dff_B_VVtGThzh2_1),.clk(gclk));
	jdff dff_B_QDX8E3WK0_1(.din(w_dff_B_VVtGThzh2_1),.dout(w_dff_B_QDX8E3WK0_1),.clk(gclk));
	jdff dff_B_PyLaqtzv6_1(.din(w_dff_B_QDX8E3WK0_1),.dout(w_dff_B_PyLaqtzv6_1),.clk(gclk));
	jdff dff_B_D4rFeW5n7_1(.din(w_dff_B_PyLaqtzv6_1),.dout(w_dff_B_D4rFeW5n7_1),.clk(gclk));
	jdff dff_B_vtFGlBHl9_1(.din(w_dff_B_D4rFeW5n7_1),.dout(w_dff_B_vtFGlBHl9_1),.clk(gclk));
	jdff dff_B_YL9ZDojH2_1(.din(w_dff_B_vtFGlBHl9_1),.dout(w_dff_B_YL9ZDojH2_1),.clk(gclk));
	jdff dff_B_vww5tgWF5_1(.din(w_dff_B_YL9ZDojH2_1),.dout(w_dff_B_vww5tgWF5_1),.clk(gclk));
	jdff dff_B_uR5b9UZr9_1(.din(w_dff_B_vww5tgWF5_1),.dout(w_dff_B_uR5b9UZr9_1),.clk(gclk));
	jdff dff_B_nUOTufvf3_1(.din(w_dff_B_uR5b9UZr9_1),.dout(w_dff_B_nUOTufvf3_1),.clk(gclk));
	jdff dff_B_KcqX1aL82_1(.din(w_dff_B_nUOTufvf3_1),.dout(w_dff_B_KcqX1aL82_1),.clk(gclk));
	jdff dff_B_efyeNG8K8_1(.din(w_dff_B_KcqX1aL82_1),.dout(w_dff_B_efyeNG8K8_1),.clk(gclk));
	jdff dff_B_1njcdvY62_1(.din(w_dff_B_efyeNG8K8_1),.dout(w_dff_B_1njcdvY62_1),.clk(gclk));
	jdff dff_B_7eyUq7aC7_1(.din(w_dff_B_1njcdvY62_1),.dout(w_dff_B_7eyUq7aC7_1),.clk(gclk));
	jdff dff_B_ev5jeRdp2_1(.din(w_dff_B_7eyUq7aC7_1),.dout(w_dff_B_ev5jeRdp2_1),.clk(gclk));
	jdff dff_B_nOTZb0mq6_1(.din(w_dff_B_ev5jeRdp2_1),.dout(w_dff_B_nOTZb0mq6_1),.clk(gclk));
	jdff dff_B_g5AosEdZ8_1(.din(w_dff_B_nOTZb0mq6_1),.dout(w_dff_B_g5AosEdZ8_1),.clk(gclk));
	jdff dff_B_axowICWa3_1(.din(w_dff_B_g5AosEdZ8_1),.dout(w_dff_B_axowICWa3_1),.clk(gclk));
	jdff dff_B_sNAt40SC3_1(.din(w_dff_B_axowICWa3_1),.dout(w_dff_B_sNAt40SC3_1),.clk(gclk));
	jdff dff_B_K9tW33W14_1(.din(w_dff_B_sNAt40SC3_1),.dout(w_dff_B_K9tW33W14_1),.clk(gclk));
	jdff dff_B_JByQrClz1_1(.din(w_dff_B_K9tW33W14_1),.dout(w_dff_B_JByQrClz1_1),.clk(gclk));
	jdff dff_B_qxZzGxFs4_1(.din(w_dff_B_JByQrClz1_1),.dout(w_dff_B_qxZzGxFs4_1),.clk(gclk));
	jdff dff_B_dTiwJBqc5_1(.din(w_dff_B_qxZzGxFs4_1),.dout(w_dff_B_dTiwJBqc5_1),.clk(gclk));
	jdff dff_B_TYG1D1pQ0_1(.din(w_dff_B_dTiwJBqc5_1),.dout(w_dff_B_TYG1D1pQ0_1),.clk(gclk));
	jdff dff_B_Ob6aHVnN7_1(.din(w_dff_B_TYG1D1pQ0_1),.dout(w_dff_B_Ob6aHVnN7_1),.clk(gclk));
	jdff dff_B_jwyhO8Vs8_1(.din(w_dff_B_Ob6aHVnN7_1),.dout(w_dff_B_jwyhO8Vs8_1),.clk(gclk));
	jdff dff_B_7AnpxpV43_1(.din(w_dff_B_jwyhO8Vs8_1),.dout(w_dff_B_7AnpxpV43_1),.clk(gclk));
	jdff dff_B_OkSfpMsf8_1(.din(w_dff_B_7AnpxpV43_1),.dout(w_dff_B_OkSfpMsf8_1),.clk(gclk));
	jdff dff_B_WCrdtPIC6_1(.din(w_dff_B_OkSfpMsf8_1),.dout(w_dff_B_WCrdtPIC6_1),.clk(gclk));
	jdff dff_B_ElMsHhza8_1(.din(w_dff_B_WCrdtPIC6_1),.dout(w_dff_B_ElMsHhza8_1),.clk(gclk));
	jdff dff_B_RHRuAJWm6_1(.din(w_dff_B_ElMsHhza8_1),.dout(w_dff_B_RHRuAJWm6_1),.clk(gclk));
	jdff dff_B_PyBmSSVk2_1(.din(w_dff_B_RHRuAJWm6_1),.dout(w_dff_B_PyBmSSVk2_1),.clk(gclk));
	jdff dff_B_B7CZDynS5_1(.din(w_dff_B_PyBmSSVk2_1),.dout(w_dff_B_B7CZDynS5_1),.clk(gclk));
	jdff dff_B_50wj6ssY4_1(.din(w_dff_B_B7CZDynS5_1),.dout(w_dff_B_50wj6ssY4_1),.clk(gclk));
	jdff dff_B_lOZSlXPt3_1(.din(w_dff_B_50wj6ssY4_1),.dout(w_dff_B_lOZSlXPt3_1),.clk(gclk));
	jdff dff_B_ODOVFQ8H0_1(.din(w_dff_B_lOZSlXPt3_1),.dout(w_dff_B_ODOVFQ8H0_1),.clk(gclk));
	jdff dff_B_JGTGbXnm5_1(.din(w_dff_B_ODOVFQ8H0_1),.dout(w_dff_B_JGTGbXnm5_1),.clk(gclk));
	jdff dff_B_DMB2Lh6Q1_1(.din(w_dff_B_JGTGbXnm5_1),.dout(w_dff_B_DMB2Lh6Q1_1),.clk(gclk));
	jdff dff_B_dhqkdMmc0_1(.din(w_dff_B_DMB2Lh6Q1_1),.dout(w_dff_B_dhqkdMmc0_1),.clk(gclk));
	jdff dff_B_5fkAPVop7_1(.din(w_dff_B_dhqkdMmc0_1),.dout(w_dff_B_5fkAPVop7_1),.clk(gclk));
	jdff dff_B_CfX0MTeq8_1(.din(w_dff_B_5fkAPVop7_1),.dout(w_dff_B_CfX0MTeq8_1),.clk(gclk));
	jdff dff_B_f3zwWfhV4_1(.din(w_dff_B_CfX0MTeq8_1),.dout(w_dff_B_f3zwWfhV4_1),.clk(gclk));
	jdff dff_B_3WLiYBPk8_1(.din(w_dff_B_f3zwWfhV4_1),.dout(w_dff_B_3WLiYBPk8_1),.clk(gclk));
	jdff dff_B_xGimSENv5_1(.din(w_dff_B_3WLiYBPk8_1),.dout(w_dff_B_xGimSENv5_1),.clk(gclk));
	jdff dff_B_CKn9l4Kr1_1(.din(w_dff_B_xGimSENv5_1),.dout(w_dff_B_CKn9l4Kr1_1),.clk(gclk));
	jdff dff_B_9ocvr2sP9_1(.din(w_dff_B_CKn9l4Kr1_1),.dout(w_dff_B_9ocvr2sP9_1),.clk(gclk));
	jdff dff_B_O20G46hs7_1(.din(w_dff_B_9ocvr2sP9_1),.dout(w_dff_B_O20G46hs7_1),.clk(gclk));
	jdff dff_B_PoK5GwyZ2_1(.din(w_dff_B_O20G46hs7_1),.dout(w_dff_B_PoK5GwyZ2_1),.clk(gclk));
	jdff dff_B_Cv7ae5305_1(.din(w_dff_B_PoK5GwyZ2_1),.dout(w_dff_B_Cv7ae5305_1),.clk(gclk));
	jdff dff_B_mGo7EScm5_1(.din(w_dff_B_Cv7ae5305_1),.dout(w_dff_B_mGo7EScm5_1),.clk(gclk));
	jdff dff_B_lWeG9KZw3_1(.din(w_dff_B_mGo7EScm5_1),.dout(w_dff_B_lWeG9KZw3_1),.clk(gclk));
	jdff dff_B_LX5pjq8p0_1(.din(w_dff_B_lWeG9KZw3_1),.dout(w_dff_B_LX5pjq8p0_1),.clk(gclk));
	jdff dff_B_O7S507ih5_1(.din(w_dff_B_LX5pjq8p0_1),.dout(w_dff_B_O7S507ih5_1),.clk(gclk));
	jdff dff_B_YfIyJNHL8_1(.din(w_dff_B_O7S507ih5_1),.dout(w_dff_B_YfIyJNHL8_1),.clk(gclk));
	jdff dff_B_zJTwdKRq9_1(.din(w_dff_B_YfIyJNHL8_1),.dout(w_dff_B_zJTwdKRq9_1),.clk(gclk));
	jdff dff_B_m8jD3M1a0_1(.din(w_dff_B_zJTwdKRq9_1),.dout(w_dff_B_m8jD3M1a0_1),.clk(gclk));
	jdff dff_B_igDalDOA5_1(.din(w_dff_B_m8jD3M1a0_1),.dout(w_dff_B_igDalDOA5_1),.clk(gclk));
	jdff dff_B_73dKzfCz6_1(.din(w_dff_B_igDalDOA5_1),.dout(w_dff_B_73dKzfCz6_1),.clk(gclk));
	jdff dff_B_RTDxXUBi6_1(.din(w_dff_B_73dKzfCz6_1),.dout(w_dff_B_RTDxXUBi6_1),.clk(gclk));
	jdff dff_B_Gzeak3hw2_1(.din(w_dff_B_RTDxXUBi6_1),.dout(w_dff_B_Gzeak3hw2_1),.clk(gclk));
	jdff dff_B_ndxTx1pN5_1(.din(w_dff_B_Gzeak3hw2_1),.dout(w_dff_B_ndxTx1pN5_1),.clk(gclk));
	jdff dff_B_5dI8zPV48_1(.din(w_dff_B_ndxTx1pN5_1),.dout(w_dff_B_5dI8zPV48_1),.clk(gclk));
	jdff dff_B_OtzK438z1_1(.din(w_dff_B_5dI8zPV48_1),.dout(w_dff_B_OtzK438z1_1),.clk(gclk));
	jdff dff_B_UN7YaIu62_1(.din(w_dff_B_OtzK438z1_1),.dout(w_dff_B_UN7YaIu62_1),.clk(gclk));
	jdff dff_B_RwGBgBiC1_1(.din(w_dff_B_UN7YaIu62_1),.dout(w_dff_B_RwGBgBiC1_1),.clk(gclk));
	jdff dff_B_sfZVOxTI8_1(.din(w_dff_B_RwGBgBiC1_1),.dout(w_dff_B_sfZVOxTI8_1),.clk(gclk));
	jdff dff_B_q7asw41e8_1(.din(w_dff_B_sfZVOxTI8_1),.dout(w_dff_B_q7asw41e8_1),.clk(gclk));
	jdff dff_B_lrD7kicI6_1(.din(w_dff_B_q7asw41e8_1),.dout(w_dff_B_lrD7kicI6_1),.clk(gclk));
	jdff dff_B_7dA3H1dG9_1(.din(w_dff_B_lrD7kicI6_1),.dout(w_dff_B_7dA3H1dG9_1),.clk(gclk));
	jdff dff_B_MBBr2bSI5_1(.din(w_dff_B_7dA3H1dG9_1),.dout(w_dff_B_MBBr2bSI5_1),.clk(gclk));
	jdff dff_B_taRdgtTr3_1(.din(w_dff_B_MBBr2bSI5_1),.dout(w_dff_B_taRdgtTr3_1),.clk(gclk));
	jdff dff_B_SDLOufBX6_1(.din(w_dff_B_taRdgtTr3_1),.dout(w_dff_B_SDLOufBX6_1),.clk(gclk));
	jdff dff_B_TIWcSlAI4_1(.din(w_dff_B_SDLOufBX6_1),.dout(w_dff_B_TIWcSlAI4_1),.clk(gclk));
	jdff dff_B_dEodIcwZ0_1(.din(w_dff_B_TIWcSlAI4_1),.dout(w_dff_B_dEodIcwZ0_1),.clk(gclk));
	jdff dff_B_yGIVbhBp8_1(.din(w_dff_B_dEodIcwZ0_1),.dout(w_dff_B_yGIVbhBp8_1),.clk(gclk));
	jdff dff_B_pW7hpMga7_1(.din(w_dff_B_yGIVbhBp8_1),.dout(w_dff_B_pW7hpMga7_1),.clk(gclk));
	jdff dff_B_07A6QlD61_1(.din(w_dff_B_pW7hpMga7_1),.dout(w_dff_B_07A6QlD61_1),.clk(gclk));
	jdff dff_B_1SKjaigN2_1(.din(w_dff_B_07A6QlD61_1),.dout(w_dff_B_1SKjaigN2_1),.clk(gclk));
	jdff dff_B_vpwAAi2W0_1(.din(w_dff_B_1SKjaigN2_1),.dout(w_dff_B_vpwAAi2W0_1),.clk(gclk));
	jdff dff_B_Vdv0FRq96_1(.din(w_dff_B_vpwAAi2W0_1),.dout(w_dff_B_Vdv0FRq96_1),.clk(gclk));
	jdff dff_B_I9OgCQ9m8_1(.din(w_dff_B_Vdv0FRq96_1),.dout(w_dff_B_I9OgCQ9m8_1),.clk(gclk));
	jdff dff_B_nSgMasaR8_1(.din(w_dff_B_I9OgCQ9m8_1),.dout(w_dff_B_nSgMasaR8_1),.clk(gclk));
	jdff dff_B_jablWl1A6_1(.din(w_dff_B_nSgMasaR8_1),.dout(w_dff_B_jablWl1A6_1),.clk(gclk));
	jdff dff_B_x0zFPHjr0_1(.din(w_dff_B_jablWl1A6_1),.dout(w_dff_B_x0zFPHjr0_1),.clk(gclk));
	jdff dff_B_HY9tid950_1(.din(w_dff_B_x0zFPHjr0_1),.dout(w_dff_B_HY9tid950_1),.clk(gclk));
	jdff dff_B_prkOEvLy1_1(.din(w_dff_B_HY9tid950_1),.dout(w_dff_B_prkOEvLy1_1),.clk(gclk));
	jdff dff_B_gjoULGb32_1(.din(w_dff_B_prkOEvLy1_1),.dout(w_dff_B_gjoULGb32_1),.clk(gclk));
	jdff dff_B_zIDCfSlT4_0(.din(n949),.dout(w_dff_B_zIDCfSlT4_0),.clk(gclk));
	jdff dff_B_MRH0kbpu9_0(.din(w_dff_B_zIDCfSlT4_0),.dout(w_dff_B_MRH0kbpu9_0),.clk(gclk));
	jdff dff_B_7ZV0rU0I7_0(.din(w_dff_B_MRH0kbpu9_0),.dout(w_dff_B_7ZV0rU0I7_0),.clk(gclk));
	jdff dff_B_Y1Z3YWoP0_0(.din(w_dff_B_7ZV0rU0I7_0),.dout(w_dff_B_Y1Z3YWoP0_0),.clk(gclk));
	jdff dff_B_vP4xMjMZ2_0(.din(w_dff_B_Y1Z3YWoP0_0),.dout(w_dff_B_vP4xMjMZ2_0),.clk(gclk));
	jdff dff_B_wgVcbYj93_0(.din(w_dff_B_vP4xMjMZ2_0),.dout(w_dff_B_wgVcbYj93_0),.clk(gclk));
	jdff dff_B_RedyTcYe6_0(.din(w_dff_B_wgVcbYj93_0),.dout(w_dff_B_RedyTcYe6_0),.clk(gclk));
	jdff dff_B_mqeMtM671_0(.din(w_dff_B_RedyTcYe6_0),.dout(w_dff_B_mqeMtM671_0),.clk(gclk));
	jdff dff_B_J1cb6B2A0_0(.din(w_dff_B_mqeMtM671_0),.dout(w_dff_B_J1cb6B2A0_0),.clk(gclk));
	jdff dff_B_91c1GROD5_0(.din(w_dff_B_J1cb6B2A0_0),.dout(w_dff_B_91c1GROD5_0),.clk(gclk));
	jdff dff_B_vVVEWpUC4_0(.din(w_dff_B_91c1GROD5_0),.dout(w_dff_B_vVVEWpUC4_0),.clk(gclk));
	jdff dff_B_d3JOicTv0_0(.din(w_dff_B_vVVEWpUC4_0),.dout(w_dff_B_d3JOicTv0_0),.clk(gclk));
	jdff dff_B_fQw0xfZT9_0(.din(w_dff_B_d3JOicTv0_0),.dout(w_dff_B_fQw0xfZT9_0),.clk(gclk));
	jdff dff_B_ztxYsfqY5_0(.din(w_dff_B_fQw0xfZT9_0),.dout(w_dff_B_ztxYsfqY5_0),.clk(gclk));
	jdff dff_B_5vK0gKNH0_0(.din(w_dff_B_ztxYsfqY5_0),.dout(w_dff_B_5vK0gKNH0_0),.clk(gclk));
	jdff dff_B_a46F5i661_0(.din(w_dff_B_5vK0gKNH0_0),.dout(w_dff_B_a46F5i661_0),.clk(gclk));
	jdff dff_B_VO89RzTc6_0(.din(w_dff_B_a46F5i661_0),.dout(w_dff_B_VO89RzTc6_0),.clk(gclk));
	jdff dff_B_TOZpVuYs8_0(.din(w_dff_B_VO89RzTc6_0),.dout(w_dff_B_TOZpVuYs8_0),.clk(gclk));
	jdff dff_B_tcfODsTj9_0(.din(w_dff_B_TOZpVuYs8_0),.dout(w_dff_B_tcfODsTj9_0),.clk(gclk));
	jdff dff_B_Ddb5UEzH3_0(.din(w_dff_B_tcfODsTj9_0),.dout(w_dff_B_Ddb5UEzH3_0),.clk(gclk));
	jdff dff_B_rbOTEwN20_0(.din(w_dff_B_Ddb5UEzH3_0),.dout(w_dff_B_rbOTEwN20_0),.clk(gclk));
	jdff dff_B_JuoW0pJP8_0(.din(w_dff_B_rbOTEwN20_0),.dout(w_dff_B_JuoW0pJP8_0),.clk(gclk));
	jdff dff_B_DXGRnf9x0_0(.din(w_dff_B_JuoW0pJP8_0),.dout(w_dff_B_DXGRnf9x0_0),.clk(gclk));
	jdff dff_B_QkUpHHBg5_0(.din(w_dff_B_DXGRnf9x0_0),.dout(w_dff_B_QkUpHHBg5_0),.clk(gclk));
	jdff dff_B_Ny9nz9O93_0(.din(w_dff_B_QkUpHHBg5_0),.dout(w_dff_B_Ny9nz9O93_0),.clk(gclk));
	jdff dff_B_hGEzkZkF7_0(.din(w_dff_B_Ny9nz9O93_0),.dout(w_dff_B_hGEzkZkF7_0),.clk(gclk));
	jdff dff_B_8b7OOEIj0_0(.din(w_dff_B_hGEzkZkF7_0),.dout(w_dff_B_8b7OOEIj0_0),.clk(gclk));
	jdff dff_B_Db4PHfoP2_0(.din(w_dff_B_8b7OOEIj0_0),.dout(w_dff_B_Db4PHfoP2_0),.clk(gclk));
	jdff dff_B_f6hIX16U3_0(.din(w_dff_B_Db4PHfoP2_0),.dout(w_dff_B_f6hIX16U3_0),.clk(gclk));
	jdff dff_B_WngVcNBa7_0(.din(w_dff_B_f6hIX16U3_0),.dout(w_dff_B_WngVcNBa7_0),.clk(gclk));
	jdff dff_B_It7XBfVE7_0(.din(w_dff_B_WngVcNBa7_0),.dout(w_dff_B_It7XBfVE7_0),.clk(gclk));
	jdff dff_B_vf99utdR5_0(.din(w_dff_B_It7XBfVE7_0),.dout(w_dff_B_vf99utdR5_0),.clk(gclk));
	jdff dff_B_CJ835o1m4_0(.din(w_dff_B_vf99utdR5_0),.dout(w_dff_B_CJ835o1m4_0),.clk(gclk));
	jdff dff_B_kU7BB5eZ1_0(.din(w_dff_B_CJ835o1m4_0),.dout(w_dff_B_kU7BB5eZ1_0),.clk(gclk));
	jdff dff_B_Mt64mcxQ1_0(.din(w_dff_B_kU7BB5eZ1_0),.dout(w_dff_B_Mt64mcxQ1_0),.clk(gclk));
	jdff dff_B_9tpLwi0n1_0(.din(w_dff_B_Mt64mcxQ1_0),.dout(w_dff_B_9tpLwi0n1_0),.clk(gclk));
	jdff dff_B_X769e3gl8_0(.din(w_dff_B_9tpLwi0n1_0),.dout(w_dff_B_X769e3gl8_0),.clk(gclk));
	jdff dff_B_wCynEx8b6_0(.din(w_dff_B_X769e3gl8_0),.dout(w_dff_B_wCynEx8b6_0),.clk(gclk));
	jdff dff_B_nPENxYqD9_0(.din(w_dff_B_wCynEx8b6_0),.dout(w_dff_B_nPENxYqD9_0),.clk(gclk));
	jdff dff_B_8LAVOjQi0_0(.din(w_dff_B_nPENxYqD9_0),.dout(w_dff_B_8LAVOjQi0_0),.clk(gclk));
	jdff dff_B_C4fUTGvb4_0(.din(w_dff_B_8LAVOjQi0_0),.dout(w_dff_B_C4fUTGvb4_0),.clk(gclk));
	jdff dff_B_mQJFSKgO3_0(.din(w_dff_B_C4fUTGvb4_0),.dout(w_dff_B_mQJFSKgO3_0),.clk(gclk));
	jdff dff_B_mxi2saeZ8_0(.din(w_dff_B_mQJFSKgO3_0),.dout(w_dff_B_mxi2saeZ8_0),.clk(gclk));
	jdff dff_B_dhazEBQh2_0(.din(w_dff_B_mxi2saeZ8_0),.dout(w_dff_B_dhazEBQh2_0),.clk(gclk));
	jdff dff_B_narvYCok5_0(.din(w_dff_B_dhazEBQh2_0),.dout(w_dff_B_narvYCok5_0),.clk(gclk));
	jdff dff_B_HZYWSKlb8_0(.din(w_dff_B_narvYCok5_0),.dout(w_dff_B_HZYWSKlb8_0),.clk(gclk));
	jdff dff_B_qxmaXVaL1_0(.din(w_dff_B_HZYWSKlb8_0),.dout(w_dff_B_qxmaXVaL1_0),.clk(gclk));
	jdff dff_B_exqnjkt53_0(.din(w_dff_B_qxmaXVaL1_0),.dout(w_dff_B_exqnjkt53_0),.clk(gclk));
	jdff dff_B_GMIO81oT5_0(.din(w_dff_B_exqnjkt53_0),.dout(w_dff_B_GMIO81oT5_0),.clk(gclk));
	jdff dff_B_8oGHIq6R9_0(.din(w_dff_B_GMIO81oT5_0),.dout(w_dff_B_8oGHIq6R9_0),.clk(gclk));
	jdff dff_B_JL310I535_0(.din(w_dff_B_8oGHIq6R9_0),.dout(w_dff_B_JL310I535_0),.clk(gclk));
	jdff dff_B_WNY353GA7_0(.din(w_dff_B_JL310I535_0),.dout(w_dff_B_WNY353GA7_0),.clk(gclk));
	jdff dff_B_Z8jo0LFH6_0(.din(w_dff_B_WNY353GA7_0),.dout(w_dff_B_Z8jo0LFH6_0),.clk(gclk));
	jdff dff_B_iLpQhrys9_0(.din(w_dff_B_Z8jo0LFH6_0),.dout(w_dff_B_iLpQhrys9_0),.clk(gclk));
	jdff dff_B_grDKkQ9S1_0(.din(w_dff_B_iLpQhrys9_0),.dout(w_dff_B_grDKkQ9S1_0),.clk(gclk));
	jdff dff_B_YMInR4TI5_0(.din(w_dff_B_grDKkQ9S1_0),.dout(w_dff_B_YMInR4TI5_0),.clk(gclk));
	jdff dff_B_YpBGOVyZ3_0(.din(w_dff_B_YMInR4TI5_0),.dout(w_dff_B_YpBGOVyZ3_0),.clk(gclk));
	jdff dff_B_xOTPnXLV3_0(.din(w_dff_B_YpBGOVyZ3_0),.dout(w_dff_B_xOTPnXLV3_0),.clk(gclk));
	jdff dff_B_kfb600uh7_0(.din(w_dff_B_xOTPnXLV3_0),.dout(w_dff_B_kfb600uh7_0),.clk(gclk));
	jdff dff_B_MbfewOqH4_0(.din(w_dff_B_kfb600uh7_0),.dout(w_dff_B_MbfewOqH4_0),.clk(gclk));
	jdff dff_B_EeUGYaSy1_0(.din(w_dff_B_MbfewOqH4_0),.dout(w_dff_B_EeUGYaSy1_0),.clk(gclk));
	jdff dff_B_sbNHupP22_0(.din(w_dff_B_EeUGYaSy1_0),.dout(w_dff_B_sbNHupP22_0),.clk(gclk));
	jdff dff_B_U6z1YcMv7_0(.din(w_dff_B_sbNHupP22_0),.dout(w_dff_B_U6z1YcMv7_0),.clk(gclk));
	jdff dff_B_TFRxEf5t4_0(.din(w_dff_B_U6z1YcMv7_0),.dout(w_dff_B_TFRxEf5t4_0),.clk(gclk));
	jdff dff_B_AV1Y5qNW1_0(.din(w_dff_B_TFRxEf5t4_0),.dout(w_dff_B_AV1Y5qNW1_0),.clk(gclk));
	jdff dff_B_rZ5LQRvG9_0(.din(w_dff_B_AV1Y5qNW1_0),.dout(w_dff_B_rZ5LQRvG9_0),.clk(gclk));
	jdff dff_B_W6Urze7c0_0(.din(w_dff_B_rZ5LQRvG9_0),.dout(w_dff_B_W6Urze7c0_0),.clk(gclk));
	jdff dff_B_2QpAcxgm7_0(.din(w_dff_B_W6Urze7c0_0),.dout(w_dff_B_2QpAcxgm7_0),.clk(gclk));
	jdff dff_B_ic3lSNup9_0(.din(w_dff_B_2QpAcxgm7_0),.dout(w_dff_B_ic3lSNup9_0),.clk(gclk));
	jdff dff_B_oLoM5QvQ7_0(.din(w_dff_B_ic3lSNup9_0),.dout(w_dff_B_oLoM5QvQ7_0),.clk(gclk));
	jdff dff_B_UPe20AvG6_0(.din(w_dff_B_oLoM5QvQ7_0),.dout(w_dff_B_UPe20AvG6_0),.clk(gclk));
	jdff dff_B_ifnVewRr5_0(.din(w_dff_B_UPe20AvG6_0),.dout(w_dff_B_ifnVewRr5_0),.clk(gclk));
	jdff dff_B_NPkroi0A1_0(.din(w_dff_B_ifnVewRr5_0),.dout(w_dff_B_NPkroi0A1_0),.clk(gclk));
	jdff dff_B_irbehqs29_0(.din(w_dff_B_NPkroi0A1_0),.dout(w_dff_B_irbehqs29_0),.clk(gclk));
	jdff dff_B_vZDPM6ka0_0(.din(w_dff_B_irbehqs29_0),.dout(w_dff_B_vZDPM6ka0_0),.clk(gclk));
	jdff dff_B_711Y4oqI9_0(.din(w_dff_B_vZDPM6ka0_0),.dout(w_dff_B_711Y4oqI9_0),.clk(gclk));
	jdff dff_B_j5S9OtfC6_0(.din(w_dff_B_711Y4oqI9_0),.dout(w_dff_B_j5S9OtfC6_0),.clk(gclk));
	jdff dff_B_VGSlfaPw1_0(.din(w_dff_B_j5S9OtfC6_0),.dout(w_dff_B_VGSlfaPw1_0),.clk(gclk));
	jdff dff_B_ZCImlmkd5_0(.din(w_dff_B_VGSlfaPw1_0),.dout(w_dff_B_ZCImlmkd5_0),.clk(gclk));
	jdff dff_B_eJoBJKN96_0(.din(w_dff_B_ZCImlmkd5_0),.dout(w_dff_B_eJoBJKN96_0),.clk(gclk));
	jdff dff_B_jbulfgBo7_0(.din(w_dff_B_eJoBJKN96_0),.dout(w_dff_B_jbulfgBo7_0),.clk(gclk));
	jdff dff_B_TFUZBVYt3_0(.din(w_dff_B_jbulfgBo7_0),.dout(w_dff_B_TFUZBVYt3_0),.clk(gclk));
	jdff dff_B_cbkSIbUg6_0(.din(w_dff_B_TFUZBVYt3_0),.dout(w_dff_B_cbkSIbUg6_0),.clk(gclk));
	jdff dff_B_N8TKDq7N2_0(.din(w_dff_B_cbkSIbUg6_0),.dout(w_dff_B_N8TKDq7N2_0),.clk(gclk));
	jdff dff_B_5R023Dvz3_0(.din(w_dff_B_N8TKDq7N2_0),.dout(w_dff_B_5R023Dvz3_0),.clk(gclk));
	jdff dff_B_Z81DTIDr7_0(.din(w_dff_B_5R023Dvz3_0),.dout(w_dff_B_Z81DTIDr7_0),.clk(gclk));
	jdff dff_B_EF3hGMje8_0(.din(w_dff_B_Z81DTIDr7_0),.dout(w_dff_B_EF3hGMje8_0),.clk(gclk));
	jdff dff_B_CuIHmZcq4_0(.din(w_dff_B_EF3hGMje8_0),.dout(w_dff_B_CuIHmZcq4_0),.clk(gclk));
	jdff dff_B_Qd2FPUwi0_0(.din(w_dff_B_CuIHmZcq4_0),.dout(w_dff_B_Qd2FPUwi0_0),.clk(gclk));
	jdff dff_B_q3n5TzjL9_0(.din(w_dff_B_Qd2FPUwi0_0),.dout(w_dff_B_q3n5TzjL9_0),.clk(gclk));
	jdff dff_B_YuvgbGU55_0(.din(w_dff_B_q3n5TzjL9_0),.dout(w_dff_B_YuvgbGU55_0),.clk(gclk));
	jdff dff_B_bzPWadtA9_0(.din(w_dff_B_YuvgbGU55_0),.dout(w_dff_B_bzPWadtA9_0),.clk(gclk));
	jdff dff_B_G4FiTUOn2_0(.din(w_dff_B_bzPWadtA9_0),.dout(w_dff_B_G4FiTUOn2_0),.clk(gclk));
	jdff dff_B_Tlk8jcgs4_0(.din(w_dff_B_G4FiTUOn2_0),.dout(w_dff_B_Tlk8jcgs4_0),.clk(gclk));
	jdff dff_B_NIPgnmvE5_1(.din(n942),.dout(w_dff_B_NIPgnmvE5_1),.clk(gclk));
	jdff dff_B_GNazyr6z7_1(.din(w_dff_B_NIPgnmvE5_1),.dout(w_dff_B_GNazyr6z7_1),.clk(gclk));
	jdff dff_B_SRafIkTg8_1(.din(w_dff_B_GNazyr6z7_1),.dout(w_dff_B_SRafIkTg8_1),.clk(gclk));
	jdff dff_B_jfyKVKxb6_1(.din(w_dff_B_SRafIkTg8_1),.dout(w_dff_B_jfyKVKxb6_1),.clk(gclk));
	jdff dff_B_Gqoq2WRY9_1(.din(w_dff_B_jfyKVKxb6_1),.dout(w_dff_B_Gqoq2WRY9_1),.clk(gclk));
	jdff dff_B_hOjwb8ou8_1(.din(w_dff_B_Gqoq2WRY9_1),.dout(w_dff_B_hOjwb8ou8_1),.clk(gclk));
	jdff dff_B_nmnt5xcc6_1(.din(w_dff_B_hOjwb8ou8_1),.dout(w_dff_B_nmnt5xcc6_1),.clk(gclk));
	jdff dff_B_qfNir07L8_1(.din(w_dff_B_nmnt5xcc6_1),.dout(w_dff_B_qfNir07L8_1),.clk(gclk));
	jdff dff_B_tjXsTbGM0_1(.din(w_dff_B_qfNir07L8_1),.dout(w_dff_B_tjXsTbGM0_1),.clk(gclk));
	jdff dff_B_yThbUDN74_1(.din(w_dff_B_tjXsTbGM0_1),.dout(w_dff_B_yThbUDN74_1),.clk(gclk));
	jdff dff_B_i8uCCkZj0_1(.din(w_dff_B_yThbUDN74_1),.dout(w_dff_B_i8uCCkZj0_1),.clk(gclk));
	jdff dff_B_jc9rBImC3_1(.din(w_dff_B_i8uCCkZj0_1),.dout(w_dff_B_jc9rBImC3_1),.clk(gclk));
	jdff dff_B_sQd0kZYn2_1(.din(w_dff_B_jc9rBImC3_1),.dout(w_dff_B_sQd0kZYn2_1),.clk(gclk));
	jdff dff_B_qfWNX0J09_1(.din(w_dff_B_sQd0kZYn2_1),.dout(w_dff_B_qfWNX0J09_1),.clk(gclk));
	jdff dff_B_GWYui08G5_1(.din(w_dff_B_qfWNX0J09_1),.dout(w_dff_B_GWYui08G5_1),.clk(gclk));
	jdff dff_B_8HrnCfnF9_1(.din(w_dff_B_GWYui08G5_1),.dout(w_dff_B_8HrnCfnF9_1),.clk(gclk));
	jdff dff_B_9Psa5Rir3_1(.din(w_dff_B_8HrnCfnF9_1),.dout(w_dff_B_9Psa5Rir3_1),.clk(gclk));
	jdff dff_B_0pvI4qSP4_1(.din(w_dff_B_9Psa5Rir3_1),.dout(w_dff_B_0pvI4qSP4_1),.clk(gclk));
	jdff dff_B_8NRA4ImH2_1(.din(w_dff_B_0pvI4qSP4_1),.dout(w_dff_B_8NRA4ImH2_1),.clk(gclk));
	jdff dff_B_K3liEBnP7_1(.din(w_dff_B_8NRA4ImH2_1),.dout(w_dff_B_K3liEBnP7_1),.clk(gclk));
	jdff dff_B_CaDbtZGg6_1(.din(w_dff_B_K3liEBnP7_1),.dout(w_dff_B_CaDbtZGg6_1),.clk(gclk));
	jdff dff_B_LWQCpjxd2_1(.din(w_dff_B_CaDbtZGg6_1),.dout(w_dff_B_LWQCpjxd2_1),.clk(gclk));
	jdff dff_B_ZP2U6ziC1_1(.din(w_dff_B_LWQCpjxd2_1),.dout(w_dff_B_ZP2U6ziC1_1),.clk(gclk));
	jdff dff_B_6dO1q6LA8_1(.din(w_dff_B_ZP2U6ziC1_1),.dout(w_dff_B_6dO1q6LA8_1),.clk(gclk));
	jdff dff_B_3UhEkn1c9_1(.din(w_dff_B_6dO1q6LA8_1),.dout(w_dff_B_3UhEkn1c9_1),.clk(gclk));
	jdff dff_B_aqhEYIpX5_1(.din(w_dff_B_3UhEkn1c9_1),.dout(w_dff_B_aqhEYIpX5_1),.clk(gclk));
	jdff dff_B_TUtVtCGX2_1(.din(w_dff_B_aqhEYIpX5_1),.dout(w_dff_B_TUtVtCGX2_1),.clk(gclk));
	jdff dff_B_8f0LtSgp4_1(.din(w_dff_B_TUtVtCGX2_1),.dout(w_dff_B_8f0LtSgp4_1),.clk(gclk));
	jdff dff_B_aSMH59jL4_1(.din(w_dff_B_8f0LtSgp4_1),.dout(w_dff_B_aSMH59jL4_1),.clk(gclk));
	jdff dff_B_ihorJH7F9_1(.din(w_dff_B_aSMH59jL4_1),.dout(w_dff_B_ihorJH7F9_1),.clk(gclk));
	jdff dff_B_uJabjRPI5_1(.din(w_dff_B_ihorJH7F9_1),.dout(w_dff_B_uJabjRPI5_1),.clk(gclk));
	jdff dff_B_prlyCjJM6_1(.din(w_dff_B_uJabjRPI5_1),.dout(w_dff_B_prlyCjJM6_1),.clk(gclk));
	jdff dff_B_xqfmdQEK4_1(.din(w_dff_B_prlyCjJM6_1),.dout(w_dff_B_xqfmdQEK4_1),.clk(gclk));
	jdff dff_B_UTUw33b70_1(.din(w_dff_B_xqfmdQEK4_1),.dout(w_dff_B_UTUw33b70_1),.clk(gclk));
	jdff dff_B_YuVuYVtA3_1(.din(w_dff_B_UTUw33b70_1),.dout(w_dff_B_YuVuYVtA3_1),.clk(gclk));
	jdff dff_B_y3eYixxI9_1(.din(w_dff_B_YuVuYVtA3_1),.dout(w_dff_B_y3eYixxI9_1),.clk(gclk));
	jdff dff_B_4Z6DRA540_1(.din(w_dff_B_y3eYixxI9_1),.dout(w_dff_B_4Z6DRA540_1),.clk(gclk));
	jdff dff_B_4bmZvCzy4_1(.din(w_dff_B_4Z6DRA540_1),.dout(w_dff_B_4bmZvCzy4_1),.clk(gclk));
	jdff dff_B_4hvkd2lt9_1(.din(w_dff_B_4bmZvCzy4_1),.dout(w_dff_B_4hvkd2lt9_1),.clk(gclk));
	jdff dff_B_Agmltuqy7_1(.din(w_dff_B_4hvkd2lt9_1),.dout(w_dff_B_Agmltuqy7_1),.clk(gclk));
	jdff dff_B_02laE88z8_1(.din(w_dff_B_Agmltuqy7_1),.dout(w_dff_B_02laE88z8_1),.clk(gclk));
	jdff dff_B_VZAiEAtY7_1(.din(w_dff_B_02laE88z8_1),.dout(w_dff_B_VZAiEAtY7_1),.clk(gclk));
	jdff dff_B_U9UiiICj9_1(.din(w_dff_B_VZAiEAtY7_1),.dout(w_dff_B_U9UiiICj9_1),.clk(gclk));
	jdff dff_B_mhImDYsm1_1(.din(w_dff_B_U9UiiICj9_1),.dout(w_dff_B_mhImDYsm1_1),.clk(gclk));
	jdff dff_B_vkZSsfgU6_1(.din(w_dff_B_mhImDYsm1_1),.dout(w_dff_B_vkZSsfgU6_1),.clk(gclk));
	jdff dff_B_UzAKZNwJ9_1(.din(w_dff_B_vkZSsfgU6_1),.dout(w_dff_B_UzAKZNwJ9_1),.clk(gclk));
	jdff dff_B_M0O8gISK1_1(.din(w_dff_B_UzAKZNwJ9_1),.dout(w_dff_B_M0O8gISK1_1),.clk(gclk));
	jdff dff_B_URlhlWey0_1(.din(w_dff_B_M0O8gISK1_1),.dout(w_dff_B_URlhlWey0_1),.clk(gclk));
	jdff dff_B_uUawEShs2_1(.din(w_dff_B_URlhlWey0_1),.dout(w_dff_B_uUawEShs2_1),.clk(gclk));
	jdff dff_B_lRsGibNx9_1(.din(w_dff_B_uUawEShs2_1),.dout(w_dff_B_lRsGibNx9_1),.clk(gclk));
	jdff dff_B_EVhfsF6W8_1(.din(w_dff_B_lRsGibNx9_1),.dout(w_dff_B_EVhfsF6W8_1),.clk(gclk));
	jdff dff_B_aE2G8XQ32_1(.din(w_dff_B_EVhfsF6W8_1),.dout(w_dff_B_aE2G8XQ32_1),.clk(gclk));
	jdff dff_B_QTu7zUnH1_1(.din(w_dff_B_aE2G8XQ32_1),.dout(w_dff_B_QTu7zUnH1_1),.clk(gclk));
	jdff dff_B_evK6g61U2_1(.din(w_dff_B_QTu7zUnH1_1),.dout(w_dff_B_evK6g61U2_1),.clk(gclk));
	jdff dff_B_F1YmhZjp0_1(.din(w_dff_B_evK6g61U2_1),.dout(w_dff_B_F1YmhZjp0_1),.clk(gclk));
	jdff dff_B_BJPIFfZJ7_1(.din(w_dff_B_F1YmhZjp0_1),.dout(w_dff_B_BJPIFfZJ7_1),.clk(gclk));
	jdff dff_B_v4m9yThQ1_1(.din(w_dff_B_BJPIFfZJ7_1),.dout(w_dff_B_v4m9yThQ1_1),.clk(gclk));
	jdff dff_B_1Rcas2YK4_1(.din(w_dff_B_v4m9yThQ1_1),.dout(w_dff_B_1Rcas2YK4_1),.clk(gclk));
	jdff dff_B_hU198oK02_1(.din(w_dff_B_1Rcas2YK4_1),.dout(w_dff_B_hU198oK02_1),.clk(gclk));
	jdff dff_B_YRXOFSQW0_1(.din(w_dff_B_hU198oK02_1),.dout(w_dff_B_YRXOFSQW0_1),.clk(gclk));
	jdff dff_B_OsRxHc9o2_1(.din(w_dff_B_YRXOFSQW0_1),.dout(w_dff_B_OsRxHc9o2_1),.clk(gclk));
	jdff dff_B_HyBK42dg7_1(.din(w_dff_B_OsRxHc9o2_1),.dout(w_dff_B_HyBK42dg7_1),.clk(gclk));
	jdff dff_B_RfcIotNc5_1(.din(w_dff_B_HyBK42dg7_1),.dout(w_dff_B_RfcIotNc5_1),.clk(gclk));
	jdff dff_B_11nXivdv5_1(.din(w_dff_B_RfcIotNc5_1),.dout(w_dff_B_11nXivdv5_1),.clk(gclk));
	jdff dff_B_p8GAccRn6_1(.din(w_dff_B_11nXivdv5_1),.dout(w_dff_B_p8GAccRn6_1),.clk(gclk));
	jdff dff_B_NKa6mCVm3_1(.din(w_dff_B_p8GAccRn6_1),.dout(w_dff_B_NKa6mCVm3_1),.clk(gclk));
	jdff dff_B_qKm0c2PR6_1(.din(w_dff_B_NKa6mCVm3_1),.dout(w_dff_B_qKm0c2PR6_1),.clk(gclk));
	jdff dff_B_QqTC3GqG1_1(.din(w_dff_B_qKm0c2PR6_1),.dout(w_dff_B_QqTC3GqG1_1),.clk(gclk));
	jdff dff_B_d67I1yEw2_1(.din(w_dff_B_QqTC3GqG1_1),.dout(w_dff_B_d67I1yEw2_1),.clk(gclk));
	jdff dff_B_Yvz8a1Zj4_1(.din(w_dff_B_d67I1yEw2_1),.dout(w_dff_B_Yvz8a1Zj4_1),.clk(gclk));
	jdff dff_B_DTmqrhI77_1(.din(w_dff_B_Yvz8a1Zj4_1),.dout(w_dff_B_DTmqrhI77_1),.clk(gclk));
	jdff dff_B_YTMw8jbj6_1(.din(w_dff_B_DTmqrhI77_1),.dout(w_dff_B_YTMw8jbj6_1),.clk(gclk));
	jdff dff_B_ntFNMbjf3_1(.din(w_dff_B_YTMw8jbj6_1),.dout(w_dff_B_ntFNMbjf3_1),.clk(gclk));
	jdff dff_B_G2p7C0LJ4_1(.din(w_dff_B_ntFNMbjf3_1),.dout(w_dff_B_G2p7C0LJ4_1),.clk(gclk));
	jdff dff_B_kkYTFtPX6_1(.din(w_dff_B_G2p7C0LJ4_1),.dout(w_dff_B_kkYTFtPX6_1),.clk(gclk));
	jdff dff_B_nyE2hOSS6_1(.din(w_dff_B_kkYTFtPX6_1),.dout(w_dff_B_nyE2hOSS6_1),.clk(gclk));
	jdff dff_B_fFWDEjXN2_1(.din(w_dff_B_nyE2hOSS6_1),.dout(w_dff_B_fFWDEjXN2_1),.clk(gclk));
	jdff dff_B_H7D2VEHU0_1(.din(w_dff_B_fFWDEjXN2_1),.dout(w_dff_B_H7D2VEHU0_1),.clk(gclk));
	jdff dff_B_zyLsYVRs4_1(.din(w_dff_B_H7D2VEHU0_1),.dout(w_dff_B_zyLsYVRs4_1),.clk(gclk));
	jdff dff_B_ZPxGnCnY7_1(.din(w_dff_B_zyLsYVRs4_1),.dout(w_dff_B_ZPxGnCnY7_1),.clk(gclk));
	jdff dff_B_W0U7m01G1_1(.din(w_dff_B_ZPxGnCnY7_1),.dout(w_dff_B_W0U7m01G1_1),.clk(gclk));
	jdff dff_B_PUzwXvxc8_1(.din(w_dff_B_W0U7m01G1_1),.dout(w_dff_B_PUzwXvxc8_1),.clk(gclk));
	jdff dff_B_6PVqFGWO6_1(.din(w_dff_B_PUzwXvxc8_1),.dout(w_dff_B_6PVqFGWO6_1),.clk(gclk));
	jdff dff_B_DIuDIFah8_1(.din(w_dff_B_6PVqFGWO6_1),.dout(w_dff_B_DIuDIFah8_1),.clk(gclk));
	jdff dff_B_f3Wh9rEy8_1(.din(w_dff_B_DIuDIFah8_1),.dout(w_dff_B_f3Wh9rEy8_1),.clk(gclk));
	jdff dff_B_ouW4klhi7_1(.din(w_dff_B_f3Wh9rEy8_1),.dout(w_dff_B_ouW4klhi7_1),.clk(gclk));
	jdff dff_B_5JJMuoK85_1(.din(w_dff_B_ouW4klhi7_1),.dout(w_dff_B_5JJMuoK85_1),.clk(gclk));
	jdff dff_B_5xbvey3D3_1(.din(w_dff_B_5JJMuoK85_1),.dout(w_dff_B_5xbvey3D3_1),.clk(gclk));
	jdff dff_B_DqZ3krW32_1(.din(w_dff_B_5xbvey3D3_1),.dout(w_dff_B_DqZ3krW32_1),.clk(gclk));
	jdff dff_B_uLIT2wYr9_1(.din(w_dff_B_DqZ3krW32_1),.dout(w_dff_B_uLIT2wYr9_1),.clk(gclk));
	jdff dff_B_CdufCjmh8_1(.din(w_dff_B_uLIT2wYr9_1),.dout(w_dff_B_CdufCjmh8_1),.clk(gclk));
	jdff dff_B_MLhHLfZ69_1(.din(w_dff_B_CdufCjmh8_1),.dout(w_dff_B_MLhHLfZ69_1),.clk(gclk));
	jdff dff_B_qRRscppg1_1(.din(w_dff_B_MLhHLfZ69_1),.dout(w_dff_B_qRRscppg1_1),.clk(gclk));
	jdff dff_B_lu0jKwhg7_0(.din(n943),.dout(w_dff_B_lu0jKwhg7_0),.clk(gclk));
	jdff dff_B_LMG6sXCp5_0(.din(w_dff_B_lu0jKwhg7_0),.dout(w_dff_B_LMG6sXCp5_0),.clk(gclk));
	jdff dff_B_jQimGCcU4_0(.din(w_dff_B_LMG6sXCp5_0),.dout(w_dff_B_jQimGCcU4_0),.clk(gclk));
	jdff dff_B_UGbJwrK80_0(.din(w_dff_B_jQimGCcU4_0),.dout(w_dff_B_UGbJwrK80_0),.clk(gclk));
	jdff dff_B_JbfWrsew3_0(.din(w_dff_B_UGbJwrK80_0),.dout(w_dff_B_JbfWrsew3_0),.clk(gclk));
	jdff dff_B_vvLnYKPt0_0(.din(w_dff_B_JbfWrsew3_0),.dout(w_dff_B_vvLnYKPt0_0),.clk(gclk));
	jdff dff_B_SX9cjsYO7_0(.din(w_dff_B_vvLnYKPt0_0),.dout(w_dff_B_SX9cjsYO7_0),.clk(gclk));
	jdff dff_B_a7zfLXLZ1_0(.din(w_dff_B_SX9cjsYO7_0),.dout(w_dff_B_a7zfLXLZ1_0),.clk(gclk));
	jdff dff_B_0RKhL6QD0_0(.din(w_dff_B_a7zfLXLZ1_0),.dout(w_dff_B_0RKhL6QD0_0),.clk(gclk));
	jdff dff_B_PYQyE1yt0_0(.din(w_dff_B_0RKhL6QD0_0),.dout(w_dff_B_PYQyE1yt0_0),.clk(gclk));
	jdff dff_B_TjxINM5T6_0(.din(w_dff_B_PYQyE1yt0_0),.dout(w_dff_B_TjxINM5T6_0),.clk(gclk));
	jdff dff_B_LaGT85EI4_0(.din(w_dff_B_TjxINM5T6_0),.dout(w_dff_B_LaGT85EI4_0),.clk(gclk));
	jdff dff_B_98401wJs5_0(.din(w_dff_B_LaGT85EI4_0),.dout(w_dff_B_98401wJs5_0),.clk(gclk));
	jdff dff_B_7H3l43WF2_0(.din(w_dff_B_98401wJs5_0),.dout(w_dff_B_7H3l43WF2_0),.clk(gclk));
	jdff dff_B_KkNAJwhW1_0(.din(w_dff_B_7H3l43WF2_0),.dout(w_dff_B_KkNAJwhW1_0),.clk(gclk));
	jdff dff_B_kMbZVk0N2_0(.din(w_dff_B_KkNAJwhW1_0),.dout(w_dff_B_kMbZVk0N2_0),.clk(gclk));
	jdff dff_B_uhlipbo12_0(.din(w_dff_B_kMbZVk0N2_0),.dout(w_dff_B_uhlipbo12_0),.clk(gclk));
	jdff dff_B_eU1ZMQl38_0(.din(w_dff_B_uhlipbo12_0),.dout(w_dff_B_eU1ZMQl38_0),.clk(gclk));
	jdff dff_B_FYgBgGkM1_0(.din(w_dff_B_eU1ZMQl38_0),.dout(w_dff_B_FYgBgGkM1_0),.clk(gclk));
	jdff dff_B_tdaCUUCh3_0(.din(w_dff_B_FYgBgGkM1_0),.dout(w_dff_B_tdaCUUCh3_0),.clk(gclk));
	jdff dff_B_zjaA3UCz9_0(.din(w_dff_B_tdaCUUCh3_0),.dout(w_dff_B_zjaA3UCz9_0),.clk(gclk));
	jdff dff_B_j9zhAkxk0_0(.din(w_dff_B_zjaA3UCz9_0),.dout(w_dff_B_j9zhAkxk0_0),.clk(gclk));
	jdff dff_B_bjGQrSQw3_0(.din(w_dff_B_j9zhAkxk0_0),.dout(w_dff_B_bjGQrSQw3_0),.clk(gclk));
	jdff dff_B_zKR3BpMY3_0(.din(w_dff_B_bjGQrSQw3_0),.dout(w_dff_B_zKR3BpMY3_0),.clk(gclk));
	jdff dff_B_Fsv1XcOM9_0(.din(w_dff_B_zKR3BpMY3_0),.dout(w_dff_B_Fsv1XcOM9_0),.clk(gclk));
	jdff dff_B_eP80DWHN1_0(.din(w_dff_B_Fsv1XcOM9_0),.dout(w_dff_B_eP80DWHN1_0),.clk(gclk));
	jdff dff_B_uMTO6AbD9_0(.din(w_dff_B_eP80DWHN1_0),.dout(w_dff_B_uMTO6AbD9_0),.clk(gclk));
	jdff dff_B_LqzZ19jE2_0(.din(w_dff_B_uMTO6AbD9_0),.dout(w_dff_B_LqzZ19jE2_0),.clk(gclk));
	jdff dff_B_FoXkDSWr9_0(.din(w_dff_B_LqzZ19jE2_0),.dout(w_dff_B_FoXkDSWr9_0),.clk(gclk));
	jdff dff_B_ewDUfnrO5_0(.din(w_dff_B_FoXkDSWr9_0),.dout(w_dff_B_ewDUfnrO5_0),.clk(gclk));
	jdff dff_B_bYYMEXXA5_0(.din(w_dff_B_ewDUfnrO5_0),.dout(w_dff_B_bYYMEXXA5_0),.clk(gclk));
	jdff dff_B_swqyUwyx9_0(.din(w_dff_B_bYYMEXXA5_0),.dout(w_dff_B_swqyUwyx9_0),.clk(gclk));
	jdff dff_B_4L96TeJJ7_0(.din(w_dff_B_swqyUwyx9_0),.dout(w_dff_B_4L96TeJJ7_0),.clk(gclk));
	jdff dff_B_XowcDu7J3_0(.din(w_dff_B_4L96TeJJ7_0),.dout(w_dff_B_XowcDu7J3_0),.clk(gclk));
	jdff dff_B_ZdD6P1kc7_0(.din(w_dff_B_XowcDu7J3_0),.dout(w_dff_B_ZdD6P1kc7_0),.clk(gclk));
	jdff dff_B_n4T3GGwq1_0(.din(w_dff_B_ZdD6P1kc7_0),.dout(w_dff_B_n4T3GGwq1_0),.clk(gclk));
	jdff dff_B_Q1ZtM9W36_0(.din(w_dff_B_n4T3GGwq1_0),.dout(w_dff_B_Q1ZtM9W36_0),.clk(gclk));
	jdff dff_B_yD4ZP8Ky7_0(.din(w_dff_B_Q1ZtM9W36_0),.dout(w_dff_B_yD4ZP8Ky7_0),.clk(gclk));
	jdff dff_B_JFMKQI0n4_0(.din(w_dff_B_yD4ZP8Ky7_0),.dout(w_dff_B_JFMKQI0n4_0),.clk(gclk));
	jdff dff_B_BXXTbmW67_0(.din(w_dff_B_JFMKQI0n4_0),.dout(w_dff_B_BXXTbmW67_0),.clk(gclk));
	jdff dff_B_9OzdXUnA5_0(.din(w_dff_B_BXXTbmW67_0),.dout(w_dff_B_9OzdXUnA5_0),.clk(gclk));
	jdff dff_B_6ClUdtnQ0_0(.din(w_dff_B_9OzdXUnA5_0),.dout(w_dff_B_6ClUdtnQ0_0),.clk(gclk));
	jdff dff_B_8AQy0azS0_0(.din(w_dff_B_6ClUdtnQ0_0),.dout(w_dff_B_8AQy0azS0_0),.clk(gclk));
	jdff dff_B_yYGzIpmp6_0(.din(w_dff_B_8AQy0azS0_0),.dout(w_dff_B_yYGzIpmp6_0),.clk(gclk));
	jdff dff_B_eIOcBpCL5_0(.din(w_dff_B_yYGzIpmp6_0),.dout(w_dff_B_eIOcBpCL5_0),.clk(gclk));
	jdff dff_B_soHxIGkn1_0(.din(w_dff_B_eIOcBpCL5_0),.dout(w_dff_B_soHxIGkn1_0),.clk(gclk));
	jdff dff_B_Zj7Agyuo8_0(.din(w_dff_B_soHxIGkn1_0),.dout(w_dff_B_Zj7Agyuo8_0),.clk(gclk));
	jdff dff_B_GUERlje50_0(.din(w_dff_B_Zj7Agyuo8_0),.dout(w_dff_B_GUERlje50_0),.clk(gclk));
	jdff dff_B_bLc4jksm0_0(.din(w_dff_B_GUERlje50_0),.dout(w_dff_B_bLc4jksm0_0),.clk(gclk));
	jdff dff_B_DHPiFWKz8_0(.din(w_dff_B_bLc4jksm0_0),.dout(w_dff_B_DHPiFWKz8_0),.clk(gclk));
	jdff dff_B_V8YMXhhG4_0(.din(w_dff_B_DHPiFWKz8_0),.dout(w_dff_B_V8YMXhhG4_0),.clk(gclk));
	jdff dff_B_0tOAmo6v5_0(.din(w_dff_B_V8YMXhhG4_0),.dout(w_dff_B_0tOAmo6v5_0),.clk(gclk));
	jdff dff_B_mXHFyDR38_0(.din(w_dff_B_0tOAmo6v5_0),.dout(w_dff_B_mXHFyDR38_0),.clk(gclk));
	jdff dff_B_3DUEDxSV2_0(.din(w_dff_B_mXHFyDR38_0),.dout(w_dff_B_3DUEDxSV2_0),.clk(gclk));
	jdff dff_B_CFDZZqPX4_0(.din(w_dff_B_3DUEDxSV2_0),.dout(w_dff_B_CFDZZqPX4_0),.clk(gclk));
	jdff dff_B_iUZnEXYf3_0(.din(w_dff_B_CFDZZqPX4_0),.dout(w_dff_B_iUZnEXYf3_0),.clk(gclk));
	jdff dff_B_6XQagl4x4_0(.din(w_dff_B_iUZnEXYf3_0),.dout(w_dff_B_6XQagl4x4_0),.clk(gclk));
	jdff dff_B_045SAdZ08_0(.din(w_dff_B_6XQagl4x4_0),.dout(w_dff_B_045SAdZ08_0),.clk(gclk));
	jdff dff_B_6iOHQxq56_0(.din(w_dff_B_045SAdZ08_0),.dout(w_dff_B_6iOHQxq56_0),.clk(gclk));
	jdff dff_B_ZlnGgaU10_0(.din(w_dff_B_6iOHQxq56_0),.dout(w_dff_B_ZlnGgaU10_0),.clk(gclk));
	jdff dff_B_7SNsgknd4_0(.din(w_dff_B_ZlnGgaU10_0),.dout(w_dff_B_7SNsgknd4_0),.clk(gclk));
	jdff dff_B_UkjGFXeC6_0(.din(w_dff_B_7SNsgknd4_0),.dout(w_dff_B_UkjGFXeC6_0),.clk(gclk));
	jdff dff_B_ZM99NR263_0(.din(w_dff_B_UkjGFXeC6_0),.dout(w_dff_B_ZM99NR263_0),.clk(gclk));
	jdff dff_B_giyBhSGG8_0(.din(w_dff_B_ZM99NR263_0),.dout(w_dff_B_giyBhSGG8_0),.clk(gclk));
	jdff dff_B_bC88Rmr72_0(.din(w_dff_B_giyBhSGG8_0),.dout(w_dff_B_bC88Rmr72_0),.clk(gclk));
	jdff dff_B_BFiisW189_0(.din(w_dff_B_bC88Rmr72_0),.dout(w_dff_B_BFiisW189_0),.clk(gclk));
	jdff dff_B_6e7R4Sh14_0(.din(w_dff_B_BFiisW189_0),.dout(w_dff_B_6e7R4Sh14_0),.clk(gclk));
	jdff dff_B_WbJF2mNq0_0(.din(w_dff_B_6e7R4Sh14_0),.dout(w_dff_B_WbJF2mNq0_0),.clk(gclk));
	jdff dff_B_Pd1XC5Qu7_0(.din(w_dff_B_WbJF2mNq0_0),.dout(w_dff_B_Pd1XC5Qu7_0),.clk(gclk));
	jdff dff_B_eyJLCFYt9_0(.din(w_dff_B_Pd1XC5Qu7_0),.dout(w_dff_B_eyJLCFYt9_0),.clk(gclk));
	jdff dff_B_FKDsgxv23_0(.din(w_dff_B_eyJLCFYt9_0),.dout(w_dff_B_FKDsgxv23_0),.clk(gclk));
	jdff dff_B_n4YjFBQ69_0(.din(w_dff_B_FKDsgxv23_0),.dout(w_dff_B_n4YjFBQ69_0),.clk(gclk));
	jdff dff_B_qbF6fOU16_0(.din(w_dff_B_n4YjFBQ69_0),.dout(w_dff_B_qbF6fOU16_0),.clk(gclk));
	jdff dff_B_tcBIdS1F9_0(.din(w_dff_B_qbF6fOU16_0),.dout(w_dff_B_tcBIdS1F9_0),.clk(gclk));
	jdff dff_B_5yv60ErV3_0(.din(w_dff_B_tcBIdS1F9_0),.dout(w_dff_B_5yv60ErV3_0),.clk(gclk));
	jdff dff_B_PV6UTCN74_0(.din(w_dff_B_5yv60ErV3_0),.dout(w_dff_B_PV6UTCN74_0),.clk(gclk));
	jdff dff_B_DN0IvlKQ2_0(.din(w_dff_B_PV6UTCN74_0),.dout(w_dff_B_DN0IvlKQ2_0),.clk(gclk));
	jdff dff_B_4JQHIIHQ9_0(.din(w_dff_B_DN0IvlKQ2_0),.dout(w_dff_B_4JQHIIHQ9_0),.clk(gclk));
	jdff dff_B_VlFtOg230_0(.din(w_dff_B_4JQHIIHQ9_0),.dout(w_dff_B_VlFtOg230_0),.clk(gclk));
	jdff dff_B_iRaeLmCR6_0(.din(w_dff_B_VlFtOg230_0),.dout(w_dff_B_iRaeLmCR6_0),.clk(gclk));
	jdff dff_B_pS5Sx5fS8_0(.din(w_dff_B_iRaeLmCR6_0),.dout(w_dff_B_pS5Sx5fS8_0),.clk(gclk));
	jdff dff_B_LHsiC0Jf1_0(.din(w_dff_B_pS5Sx5fS8_0),.dout(w_dff_B_LHsiC0Jf1_0),.clk(gclk));
	jdff dff_B_5madsnMo3_0(.din(w_dff_B_LHsiC0Jf1_0),.dout(w_dff_B_5madsnMo3_0),.clk(gclk));
	jdff dff_B_208MumJ28_0(.din(w_dff_B_5madsnMo3_0),.dout(w_dff_B_208MumJ28_0),.clk(gclk));
	jdff dff_B_XvplUUQN7_0(.din(w_dff_B_208MumJ28_0),.dout(w_dff_B_XvplUUQN7_0),.clk(gclk));
	jdff dff_B_d2zxyvRn8_0(.din(w_dff_B_XvplUUQN7_0),.dout(w_dff_B_d2zxyvRn8_0),.clk(gclk));
	jdff dff_B_Vs4X5a7l1_0(.din(w_dff_B_d2zxyvRn8_0),.dout(w_dff_B_Vs4X5a7l1_0),.clk(gclk));
	jdff dff_B_dEEZRkyX6_0(.din(w_dff_B_Vs4X5a7l1_0),.dout(w_dff_B_dEEZRkyX6_0),.clk(gclk));
	jdff dff_B_5OC06DAu9_0(.din(w_dff_B_dEEZRkyX6_0),.dout(w_dff_B_5OC06DAu9_0),.clk(gclk));
	jdff dff_B_RAmAeZvY4_0(.din(w_dff_B_5OC06DAu9_0),.dout(w_dff_B_RAmAeZvY4_0),.clk(gclk));
	jdff dff_B_gBxUcg4g0_0(.din(w_dff_B_RAmAeZvY4_0),.dout(w_dff_B_gBxUcg4g0_0),.clk(gclk));
	jdff dff_B_ikZRNFc48_0(.din(w_dff_B_gBxUcg4g0_0),.dout(w_dff_B_ikZRNFc48_0),.clk(gclk));
	jdff dff_B_Z53VFgFh4_0(.din(w_dff_B_ikZRNFc48_0),.dout(w_dff_B_Z53VFgFh4_0),.clk(gclk));
	jdff dff_B_gJdq2iFW4_1(.din(n936),.dout(w_dff_B_gJdq2iFW4_1),.clk(gclk));
	jdff dff_B_kxp8UXUu7_1(.din(w_dff_B_gJdq2iFW4_1),.dout(w_dff_B_kxp8UXUu7_1),.clk(gclk));
	jdff dff_B_Y8AS3hzT7_1(.din(w_dff_B_kxp8UXUu7_1),.dout(w_dff_B_Y8AS3hzT7_1),.clk(gclk));
	jdff dff_B_rYUKApbL1_1(.din(w_dff_B_Y8AS3hzT7_1),.dout(w_dff_B_rYUKApbL1_1),.clk(gclk));
	jdff dff_B_1D6fcqmm4_1(.din(w_dff_B_rYUKApbL1_1),.dout(w_dff_B_1D6fcqmm4_1),.clk(gclk));
	jdff dff_B_XTDzDp7s6_1(.din(w_dff_B_1D6fcqmm4_1),.dout(w_dff_B_XTDzDp7s6_1),.clk(gclk));
	jdff dff_B_o8HThdOc9_1(.din(w_dff_B_XTDzDp7s6_1),.dout(w_dff_B_o8HThdOc9_1),.clk(gclk));
	jdff dff_B_BVLnBUKQ7_1(.din(w_dff_B_o8HThdOc9_1),.dout(w_dff_B_BVLnBUKQ7_1),.clk(gclk));
	jdff dff_B_Q72bFlLb5_1(.din(w_dff_B_BVLnBUKQ7_1),.dout(w_dff_B_Q72bFlLb5_1),.clk(gclk));
	jdff dff_B_7w8HJnUw1_1(.din(w_dff_B_Q72bFlLb5_1),.dout(w_dff_B_7w8HJnUw1_1),.clk(gclk));
	jdff dff_B_Earm1Lbh5_1(.din(w_dff_B_7w8HJnUw1_1),.dout(w_dff_B_Earm1Lbh5_1),.clk(gclk));
	jdff dff_B_AQCtyrYs0_1(.din(w_dff_B_Earm1Lbh5_1),.dout(w_dff_B_AQCtyrYs0_1),.clk(gclk));
	jdff dff_B_XLPQlUWJ3_1(.din(w_dff_B_AQCtyrYs0_1),.dout(w_dff_B_XLPQlUWJ3_1),.clk(gclk));
	jdff dff_B_a40VwrMN9_1(.din(w_dff_B_XLPQlUWJ3_1),.dout(w_dff_B_a40VwrMN9_1),.clk(gclk));
	jdff dff_B_OXHbIwbY8_1(.din(w_dff_B_a40VwrMN9_1),.dout(w_dff_B_OXHbIwbY8_1),.clk(gclk));
	jdff dff_B_nClTPOUA0_1(.din(w_dff_B_OXHbIwbY8_1),.dout(w_dff_B_nClTPOUA0_1),.clk(gclk));
	jdff dff_B_x0WGYBFI3_1(.din(w_dff_B_nClTPOUA0_1),.dout(w_dff_B_x0WGYBFI3_1),.clk(gclk));
	jdff dff_B_l0Mk3j9i2_1(.din(w_dff_B_x0WGYBFI3_1),.dout(w_dff_B_l0Mk3j9i2_1),.clk(gclk));
	jdff dff_B_oTfozGIW0_1(.din(w_dff_B_l0Mk3j9i2_1),.dout(w_dff_B_oTfozGIW0_1),.clk(gclk));
	jdff dff_B_WWOZ8LHr2_1(.din(w_dff_B_oTfozGIW0_1),.dout(w_dff_B_WWOZ8LHr2_1),.clk(gclk));
	jdff dff_B_z7ZTOhm55_1(.din(w_dff_B_WWOZ8LHr2_1),.dout(w_dff_B_z7ZTOhm55_1),.clk(gclk));
	jdff dff_B_yQOybGYQ3_1(.din(w_dff_B_z7ZTOhm55_1),.dout(w_dff_B_yQOybGYQ3_1),.clk(gclk));
	jdff dff_B_AkQFHqJJ2_1(.din(w_dff_B_yQOybGYQ3_1),.dout(w_dff_B_AkQFHqJJ2_1),.clk(gclk));
	jdff dff_B_nN68PjVC6_1(.din(w_dff_B_AkQFHqJJ2_1),.dout(w_dff_B_nN68PjVC6_1),.clk(gclk));
	jdff dff_B_2kpzQNDz3_1(.din(w_dff_B_nN68PjVC6_1),.dout(w_dff_B_2kpzQNDz3_1),.clk(gclk));
	jdff dff_B_Juay2Nov4_1(.din(w_dff_B_2kpzQNDz3_1),.dout(w_dff_B_Juay2Nov4_1),.clk(gclk));
	jdff dff_B_FXvrNmQ59_1(.din(w_dff_B_Juay2Nov4_1),.dout(w_dff_B_FXvrNmQ59_1),.clk(gclk));
	jdff dff_B_VBUE0oDI6_1(.din(w_dff_B_FXvrNmQ59_1),.dout(w_dff_B_VBUE0oDI6_1),.clk(gclk));
	jdff dff_B_fqREJ3yI4_1(.din(w_dff_B_VBUE0oDI6_1),.dout(w_dff_B_fqREJ3yI4_1),.clk(gclk));
	jdff dff_B_p4o6w6TL1_1(.din(w_dff_B_fqREJ3yI4_1),.dout(w_dff_B_p4o6w6TL1_1),.clk(gclk));
	jdff dff_B_umbdZvZk2_1(.din(w_dff_B_p4o6w6TL1_1),.dout(w_dff_B_umbdZvZk2_1),.clk(gclk));
	jdff dff_B_T0G0K86w9_1(.din(w_dff_B_umbdZvZk2_1),.dout(w_dff_B_T0G0K86w9_1),.clk(gclk));
	jdff dff_B_gjYt8e504_1(.din(w_dff_B_T0G0K86w9_1),.dout(w_dff_B_gjYt8e504_1),.clk(gclk));
	jdff dff_B_WxshiquB5_1(.din(w_dff_B_gjYt8e504_1),.dout(w_dff_B_WxshiquB5_1),.clk(gclk));
	jdff dff_B_pvL3FjqO3_1(.din(w_dff_B_WxshiquB5_1),.dout(w_dff_B_pvL3FjqO3_1),.clk(gclk));
	jdff dff_B_Oo9lCkc38_1(.din(w_dff_B_pvL3FjqO3_1),.dout(w_dff_B_Oo9lCkc38_1),.clk(gclk));
	jdff dff_B_LqZkMe9J7_1(.din(w_dff_B_Oo9lCkc38_1),.dout(w_dff_B_LqZkMe9J7_1),.clk(gclk));
	jdff dff_B_bdmcPQ3E0_1(.din(w_dff_B_LqZkMe9J7_1),.dout(w_dff_B_bdmcPQ3E0_1),.clk(gclk));
	jdff dff_B_UKYfU18j8_1(.din(w_dff_B_bdmcPQ3E0_1),.dout(w_dff_B_UKYfU18j8_1),.clk(gclk));
	jdff dff_B_xgvNeYYX7_1(.din(w_dff_B_UKYfU18j8_1),.dout(w_dff_B_xgvNeYYX7_1),.clk(gclk));
	jdff dff_B_pf5bLrZd2_1(.din(w_dff_B_xgvNeYYX7_1),.dout(w_dff_B_pf5bLrZd2_1),.clk(gclk));
	jdff dff_B_2qVzltxa0_1(.din(w_dff_B_pf5bLrZd2_1),.dout(w_dff_B_2qVzltxa0_1),.clk(gclk));
	jdff dff_B_iXjBJbqQ0_1(.din(w_dff_B_2qVzltxa0_1),.dout(w_dff_B_iXjBJbqQ0_1),.clk(gclk));
	jdff dff_B_GQOHcUtf8_1(.din(w_dff_B_iXjBJbqQ0_1),.dout(w_dff_B_GQOHcUtf8_1),.clk(gclk));
	jdff dff_B_G6aCvdQ98_1(.din(w_dff_B_GQOHcUtf8_1),.dout(w_dff_B_G6aCvdQ98_1),.clk(gclk));
	jdff dff_B_VQFU9dlP5_1(.din(w_dff_B_G6aCvdQ98_1),.dout(w_dff_B_VQFU9dlP5_1),.clk(gclk));
	jdff dff_B_HGr7RPbD3_1(.din(w_dff_B_VQFU9dlP5_1),.dout(w_dff_B_HGr7RPbD3_1),.clk(gclk));
	jdff dff_B_dDCKUA7p7_1(.din(w_dff_B_HGr7RPbD3_1),.dout(w_dff_B_dDCKUA7p7_1),.clk(gclk));
	jdff dff_B_Q4Trv6Kx3_1(.din(w_dff_B_dDCKUA7p7_1),.dout(w_dff_B_Q4Trv6Kx3_1),.clk(gclk));
	jdff dff_B_Ky9FZmxw7_1(.din(w_dff_B_Q4Trv6Kx3_1),.dout(w_dff_B_Ky9FZmxw7_1),.clk(gclk));
	jdff dff_B_kp9m1rdh1_1(.din(w_dff_B_Ky9FZmxw7_1),.dout(w_dff_B_kp9m1rdh1_1),.clk(gclk));
	jdff dff_B_dNsFh5629_1(.din(w_dff_B_kp9m1rdh1_1),.dout(w_dff_B_dNsFh5629_1),.clk(gclk));
	jdff dff_B_CMXQOyfh5_1(.din(w_dff_B_dNsFh5629_1),.dout(w_dff_B_CMXQOyfh5_1),.clk(gclk));
	jdff dff_B_g0dV1RIx1_1(.din(w_dff_B_CMXQOyfh5_1),.dout(w_dff_B_g0dV1RIx1_1),.clk(gclk));
	jdff dff_B_SLZO7cTh8_1(.din(w_dff_B_g0dV1RIx1_1),.dout(w_dff_B_SLZO7cTh8_1),.clk(gclk));
	jdff dff_B_v30Q16nc3_1(.din(w_dff_B_SLZO7cTh8_1),.dout(w_dff_B_v30Q16nc3_1),.clk(gclk));
	jdff dff_B_sFRDUQyu4_1(.din(w_dff_B_v30Q16nc3_1),.dout(w_dff_B_sFRDUQyu4_1),.clk(gclk));
	jdff dff_B_c3qqaAIE7_1(.din(w_dff_B_sFRDUQyu4_1),.dout(w_dff_B_c3qqaAIE7_1),.clk(gclk));
	jdff dff_B_1Z84bdlj8_1(.din(w_dff_B_c3qqaAIE7_1),.dout(w_dff_B_1Z84bdlj8_1),.clk(gclk));
	jdff dff_B_HeBMupr65_1(.din(w_dff_B_1Z84bdlj8_1),.dout(w_dff_B_HeBMupr65_1),.clk(gclk));
	jdff dff_B_ZtZW9Vkp9_1(.din(w_dff_B_HeBMupr65_1),.dout(w_dff_B_ZtZW9Vkp9_1),.clk(gclk));
	jdff dff_B_bTWyxHBG4_1(.din(w_dff_B_ZtZW9Vkp9_1),.dout(w_dff_B_bTWyxHBG4_1),.clk(gclk));
	jdff dff_B_JSjapsW71_1(.din(w_dff_B_bTWyxHBG4_1),.dout(w_dff_B_JSjapsW71_1),.clk(gclk));
	jdff dff_B_modIlHbJ9_1(.din(w_dff_B_JSjapsW71_1),.dout(w_dff_B_modIlHbJ9_1),.clk(gclk));
	jdff dff_B_ju0FS38I7_1(.din(w_dff_B_modIlHbJ9_1),.dout(w_dff_B_ju0FS38I7_1),.clk(gclk));
	jdff dff_B_SR7yMiT46_1(.din(w_dff_B_ju0FS38I7_1),.dout(w_dff_B_SR7yMiT46_1),.clk(gclk));
	jdff dff_B_qPlGZ4Op4_1(.din(w_dff_B_SR7yMiT46_1),.dout(w_dff_B_qPlGZ4Op4_1),.clk(gclk));
	jdff dff_B_zgHESNBO2_1(.din(w_dff_B_qPlGZ4Op4_1),.dout(w_dff_B_zgHESNBO2_1),.clk(gclk));
	jdff dff_B_6MyFkASg8_1(.din(w_dff_B_zgHESNBO2_1),.dout(w_dff_B_6MyFkASg8_1),.clk(gclk));
	jdff dff_B_1jpzhTsR7_1(.din(w_dff_B_6MyFkASg8_1),.dout(w_dff_B_1jpzhTsR7_1),.clk(gclk));
	jdff dff_B_f17KTT2q2_1(.din(w_dff_B_1jpzhTsR7_1),.dout(w_dff_B_f17KTT2q2_1),.clk(gclk));
	jdff dff_B_thw9dMyV7_1(.din(w_dff_B_f17KTT2q2_1),.dout(w_dff_B_thw9dMyV7_1),.clk(gclk));
	jdff dff_B_7tDgPT6H2_1(.din(w_dff_B_thw9dMyV7_1),.dout(w_dff_B_7tDgPT6H2_1),.clk(gclk));
	jdff dff_B_XM37YRli8_1(.din(w_dff_B_7tDgPT6H2_1),.dout(w_dff_B_XM37YRli8_1),.clk(gclk));
	jdff dff_B_AL8Jhazv9_1(.din(w_dff_B_XM37YRli8_1),.dout(w_dff_B_AL8Jhazv9_1),.clk(gclk));
	jdff dff_B_aHVoLH9V4_1(.din(w_dff_B_AL8Jhazv9_1),.dout(w_dff_B_aHVoLH9V4_1),.clk(gclk));
	jdff dff_B_PCRJhqxl5_1(.din(w_dff_B_aHVoLH9V4_1),.dout(w_dff_B_PCRJhqxl5_1),.clk(gclk));
	jdff dff_B_6Zi3mZRg6_1(.din(w_dff_B_PCRJhqxl5_1),.dout(w_dff_B_6Zi3mZRg6_1),.clk(gclk));
	jdff dff_B_5p6VndcG9_1(.din(w_dff_B_6Zi3mZRg6_1),.dout(w_dff_B_5p6VndcG9_1),.clk(gclk));
	jdff dff_B_hK8IBF6Z7_1(.din(w_dff_B_5p6VndcG9_1),.dout(w_dff_B_hK8IBF6Z7_1),.clk(gclk));
	jdff dff_B_xBgQUeLM5_1(.din(w_dff_B_hK8IBF6Z7_1),.dout(w_dff_B_xBgQUeLM5_1),.clk(gclk));
	jdff dff_B_pUYlLAwu1_1(.din(w_dff_B_xBgQUeLM5_1),.dout(w_dff_B_pUYlLAwu1_1),.clk(gclk));
	jdff dff_B_riFVKxaT3_1(.din(w_dff_B_pUYlLAwu1_1),.dout(w_dff_B_riFVKxaT3_1),.clk(gclk));
	jdff dff_B_CAxX5keN2_1(.din(w_dff_B_riFVKxaT3_1),.dout(w_dff_B_CAxX5keN2_1),.clk(gclk));
	jdff dff_B_hT9uO1Sj6_1(.din(w_dff_B_CAxX5keN2_1),.dout(w_dff_B_hT9uO1Sj6_1),.clk(gclk));
	jdff dff_B_2XG7dEL79_1(.din(w_dff_B_hT9uO1Sj6_1),.dout(w_dff_B_2XG7dEL79_1),.clk(gclk));
	jdff dff_B_aRJdYECd0_1(.din(w_dff_B_2XG7dEL79_1),.dout(w_dff_B_aRJdYECd0_1),.clk(gclk));
	jdff dff_B_Q8vzqKRK2_1(.din(w_dff_B_aRJdYECd0_1),.dout(w_dff_B_Q8vzqKRK2_1),.clk(gclk));
	jdff dff_B_NJXi8wR85_1(.din(w_dff_B_Q8vzqKRK2_1),.dout(w_dff_B_NJXi8wR85_1),.clk(gclk));
	jdff dff_B_HmwWwxAw6_1(.din(w_dff_B_NJXi8wR85_1),.dout(w_dff_B_HmwWwxAw6_1),.clk(gclk));
	jdff dff_B_ATTpfHUD2_1(.din(w_dff_B_HmwWwxAw6_1),.dout(w_dff_B_ATTpfHUD2_1),.clk(gclk));
	jdff dff_B_Vnmk2IHa8_1(.din(w_dff_B_ATTpfHUD2_1),.dout(w_dff_B_Vnmk2IHa8_1),.clk(gclk));
	jdff dff_B_lM2dOOfg6_0(.din(n937),.dout(w_dff_B_lM2dOOfg6_0),.clk(gclk));
	jdff dff_B_UVBbWmA94_0(.din(w_dff_B_lM2dOOfg6_0),.dout(w_dff_B_UVBbWmA94_0),.clk(gclk));
	jdff dff_B_O5EZFslc0_0(.din(w_dff_B_UVBbWmA94_0),.dout(w_dff_B_O5EZFslc0_0),.clk(gclk));
	jdff dff_B_wpQvMyOr8_0(.din(w_dff_B_O5EZFslc0_0),.dout(w_dff_B_wpQvMyOr8_0),.clk(gclk));
	jdff dff_B_ffZKLTDW9_0(.din(w_dff_B_wpQvMyOr8_0),.dout(w_dff_B_ffZKLTDW9_0),.clk(gclk));
	jdff dff_B_AtwWn1ak4_0(.din(w_dff_B_ffZKLTDW9_0),.dout(w_dff_B_AtwWn1ak4_0),.clk(gclk));
	jdff dff_B_JFXGJ8Q57_0(.din(w_dff_B_AtwWn1ak4_0),.dout(w_dff_B_JFXGJ8Q57_0),.clk(gclk));
	jdff dff_B_cM0XTWPi0_0(.din(w_dff_B_JFXGJ8Q57_0),.dout(w_dff_B_cM0XTWPi0_0),.clk(gclk));
	jdff dff_B_gBbmHKQx9_0(.din(w_dff_B_cM0XTWPi0_0),.dout(w_dff_B_gBbmHKQx9_0),.clk(gclk));
	jdff dff_B_8wkIgPVT6_0(.din(w_dff_B_gBbmHKQx9_0),.dout(w_dff_B_8wkIgPVT6_0),.clk(gclk));
	jdff dff_B_7IbJrvUK8_0(.din(w_dff_B_8wkIgPVT6_0),.dout(w_dff_B_7IbJrvUK8_0),.clk(gclk));
	jdff dff_B_ZFjcT3Mm6_0(.din(w_dff_B_7IbJrvUK8_0),.dout(w_dff_B_ZFjcT3Mm6_0),.clk(gclk));
	jdff dff_B_vyqccrap3_0(.din(w_dff_B_ZFjcT3Mm6_0),.dout(w_dff_B_vyqccrap3_0),.clk(gclk));
	jdff dff_B_wBEh1cYs8_0(.din(w_dff_B_vyqccrap3_0),.dout(w_dff_B_wBEh1cYs8_0),.clk(gclk));
	jdff dff_B_LEvP48ZI4_0(.din(w_dff_B_wBEh1cYs8_0),.dout(w_dff_B_LEvP48ZI4_0),.clk(gclk));
	jdff dff_B_O7o0v4391_0(.din(w_dff_B_LEvP48ZI4_0),.dout(w_dff_B_O7o0v4391_0),.clk(gclk));
	jdff dff_B_Vu0dGa9d7_0(.din(w_dff_B_O7o0v4391_0),.dout(w_dff_B_Vu0dGa9d7_0),.clk(gclk));
	jdff dff_B_ScmTPTjs2_0(.din(w_dff_B_Vu0dGa9d7_0),.dout(w_dff_B_ScmTPTjs2_0),.clk(gclk));
	jdff dff_B_CSPiqqkT7_0(.din(w_dff_B_ScmTPTjs2_0),.dout(w_dff_B_CSPiqqkT7_0),.clk(gclk));
	jdff dff_B_DAvgV9gY4_0(.din(w_dff_B_CSPiqqkT7_0),.dout(w_dff_B_DAvgV9gY4_0),.clk(gclk));
	jdff dff_B_dbwZnmVb1_0(.din(w_dff_B_DAvgV9gY4_0),.dout(w_dff_B_dbwZnmVb1_0),.clk(gclk));
	jdff dff_B_b4oSywtt6_0(.din(w_dff_B_dbwZnmVb1_0),.dout(w_dff_B_b4oSywtt6_0),.clk(gclk));
	jdff dff_B_heADqEni1_0(.din(w_dff_B_b4oSywtt6_0),.dout(w_dff_B_heADqEni1_0),.clk(gclk));
	jdff dff_B_jaJEzduF5_0(.din(w_dff_B_heADqEni1_0),.dout(w_dff_B_jaJEzduF5_0),.clk(gclk));
	jdff dff_B_ZI4LEGYH2_0(.din(w_dff_B_jaJEzduF5_0),.dout(w_dff_B_ZI4LEGYH2_0),.clk(gclk));
	jdff dff_B_yYDFQRsZ7_0(.din(w_dff_B_ZI4LEGYH2_0),.dout(w_dff_B_yYDFQRsZ7_0),.clk(gclk));
	jdff dff_B_goIIgDJs7_0(.din(w_dff_B_yYDFQRsZ7_0),.dout(w_dff_B_goIIgDJs7_0),.clk(gclk));
	jdff dff_B_wydOFzRy6_0(.din(w_dff_B_goIIgDJs7_0),.dout(w_dff_B_wydOFzRy6_0),.clk(gclk));
	jdff dff_B_eWJ5OrwX9_0(.din(w_dff_B_wydOFzRy6_0),.dout(w_dff_B_eWJ5OrwX9_0),.clk(gclk));
	jdff dff_B_dg6eiWIh2_0(.din(w_dff_B_eWJ5OrwX9_0),.dout(w_dff_B_dg6eiWIh2_0),.clk(gclk));
	jdff dff_B_WOH5FebT2_0(.din(w_dff_B_dg6eiWIh2_0),.dout(w_dff_B_WOH5FebT2_0),.clk(gclk));
	jdff dff_B_SuOwa5ZY2_0(.din(w_dff_B_WOH5FebT2_0),.dout(w_dff_B_SuOwa5ZY2_0),.clk(gclk));
	jdff dff_B_ztuftAGP7_0(.din(w_dff_B_SuOwa5ZY2_0),.dout(w_dff_B_ztuftAGP7_0),.clk(gclk));
	jdff dff_B_jWwmd1iH4_0(.din(w_dff_B_ztuftAGP7_0),.dout(w_dff_B_jWwmd1iH4_0),.clk(gclk));
	jdff dff_B_qrkXPVzr1_0(.din(w_dff_B_jWwmd1iH4_0),.dout(w_dff_B_qrkXPVzr1_0),.clk(gclk));
	jdff dff_B_NeygJGxY4_0(.din(w_dff_B_qrkXPVzr1_0),.dout(w_dff_B_NeygJGxY4_0),.clk(gclk));
	jdff dff_B_5mlTtPy62_0(.din(w_dff_B_NeygJGxY4_0),.dout(w_dff_B_5mlTtPy62_0),.clk(gclk));
	jdff dff_B_SgFXI4tH1_0(.din(w_dff_B_5mlTtPy62_0),.dout(w_dff_B_SgFXI4tH1_0),.clk(gclk));
	jdff dff_B_9xBA2FgC8_0(.din(w_dff_B_SgFXI4tH1_0),.dout(w_dff_B_9xBA2FgC8_0),.clk(gclk));
	jdff dff_B_Pn8DZBJI7_0(.din(w_dff_B_9xBA2FgC8_0),.dout(w_dff_B_Pn8DZBJI7_0),.clk(gclk));
	jdff dff_B_6BNrlVVG6_0(.din(w_dff_B_Pn8DZBJI7_0),.dout(w_dff_B_6BNrlVVG6_0),.clk(gclk));
	jdff dff_B_mSbK4Cra5_0(.din(w_dff_B_6BNrlVVG6_0),.dout(w_dff_B_mSbK4Cra5_0),.clk(gclk));
	jdff dff_B_DTSA04BY1_0(.din(w_dff_B_mSbK4Cra5_0),.dout(w_dff_B_DTSA04BY1_0),.clk(gclk));
	jdff dff_B_BB6gZxnl4_0(.din(w_dff_B_DTSA04BY1_0),.dout(w_dff_B_BB6gZxnl4_0),.clk(gclk));
	jdff dff_B_mU06QV8i2_0(.din(w_dff_B_BB6gZxnl4_0),.dout(w_dff_B_mU06QV8i2_0),.clk(gclk));
	jdff dff_B_ZZPsf6WI2_0(.din(w_dff_B_mU06QV8i2_0),.dout(w_dff_B_ZZPsf6WI2_0),.clk(gclk));
	jdff dff_B_e1xU3K620_0(.din(w_dff_B_ZZPsf6WI2_0),.dout(w_dff_B_e1xU3K620_0),.clk(gclk));
	jdff dff_B_vsYwFBOP4_0(.din(w_dff_B_e1xU3K620_0),.dout(w_dff_B_vsYwFBOP4_0),.clk(gclk));
	jdff dff_B_AQzJivG39_0(.din(w_dff_B_vsYwFBOP4_0),.dout(w_dff_B_AQzJivG39_0),.clk(gclk));
	jdff dff_B_B26oeoLo6_0(.din(w_dff_B_AQzJivG39_0),.dout(w_dff_B_B26oeoLo6_0),.clk(gclk));
	jdff dff_B_TLcpQ3IQ1_0(.din(w_dff_B_B26oeoLo6_0),.dout(w_dff_B_TLcpQ3IQ1_0),.clk(gclk));
	jdff dff_B_MGPMoaRv0_0(.din(w_dff_B_TLcpQ3IQ1_0),.dout(w_dff_B_MGPMoaRv0_0),.clk(gclk));
	jdff dff_B_wuhFgHP11_0(.din(w_dff_B_MGPMoaRv0_0),.dout(w_dff_B_wuhFgHP11_0),.clk(gclk));
	jdff dff_B_vYUpdkdO0_0(.din(w_dff_B_wuhFgHP11_0),.dout(w_dff_B_vYUpdkdO0_0),.clk(gclk));
	jdff dff_B_sbK29lDI3_0(.din(w_dff_B_vYUpdkdO0_0),.dout(w_dff_B_sbK29lDI3_0),.clk(gclk));
	jdff dff_B_GH1p1qcc2_0(.din(w_dff_B_sbK29lDI3_0),.dout(w_dff_B_GH1p1qcc2_0),.clk(gclk));
	jdff dff_B_SNATx7hZ5_0(.din(w_dff_B_GH1p1qcc2_0),.dout(w_dff_B_SNATx7hZ5_0),.clk(gclk));
	jdff dff_B_Sx5BBdHK2_0(.din(w_dff_B_SNATx7hZ5_0),.dout(w_dff_B_Sx5BBdHK2_0),.clk(gclk));
	jdff dff_B_uKMBZZ7b1_0(.din(w_dff_B_Sx5BBdHK2_0),.dout(w_dff_B_uKMBZZ7b1_0),.clk(gclk));
	jdff dff_B_B2AAVMVs9_0(.din(w_dff_B_uKMBZZ7b1_0),.dout(w_dff_B_B2AAVMVs9_0),.clk(gclk));
	jdff dff_B_T3LNFtu92_0(.din(w_dff_B_B2AAVMVs9_0),.dout(w_dff_B_T3LNFtu92_0),.clk(gclk));
	jdff dff_B_x2ILHnnz5_0(.din(w_dff_B_T3LNFtu92_0),.dout(w_dff_B_x2ILHnnz5_0),.clk(gclk));
	jdff dff_B_x9qszdhL8_0(.din(w_dff_B_x2ILHnnz5_0),.dout(w_dff_B_x9qszdhL8_0),.clk(gclk));
	jdff dff_B_UftfQlIV1_0(.din(w_dff_B_x9qszdhL8_0),.dout(w_dff_B_UftfQlIV1_0),.clk(gclk));
	jdff dff_B_vz3zVUZd8_0(.din(w_dff_B_UftfQlIV1_0),.dout(w_dff_B_vz3zVUZd8_0),.clk(gclk));
	jdff dff_B_fmk6QcDA9_0(.din(w_dff_B_vz3zVUZd8_0),.dout(w_dff_B_fmk6QcDA9_0),.clk(gclk));
	jdff dff_B_cJOc17Dj2_0(.din(w_dff_B_fmk6QcDA9_0),.dout(w_dff_B_cJOc17Dj2_0),.clk(gclk));
	jdff dff_B_lzFljsCR2_0(.din(w_dff_B_cJOc17Dj2_0),.dout(w_dff_B_lzFljsCR2_0),.clk(gclk));
	jdff dff_B_PtfeqFIx3_0(.din(w_dff_B_lzFljsCR2_0),.dout(w_dff_B_PtfeqFIx3_0),.clk(gclk));
	jdff dff_B_yep4vL4G0_0(.din(w_dff_B_PtfeqFIx3_0),.dout(w_dff_B_yep4vL4G0_0),.clk(gclk));
	jdff dff_B_NheNfkYk8_0(.din(w_dff_B_yep4vL4G0_0),.dout(w_dff_B_NheNfkYk8_0),.clk(gclk));
	jdff dff_B_UebbZUQr0_0(.din(w_dff_B_NheNfkYk8_0),.dout(w_dff_B_UebbZUQr0_0),.clk(gclk));
	jdff dff_B_br2B6fth1_0(.din(w_dff_B_UebbZUQr0_0),.dout(w_dff_B_br2B6fth1_0),.clk(gclk));
	jdff dff_B_syA4iOfo1_0(.din(w_dff_B_br2B6fth1_0),.dout(w_dff_B_syA4iOfo1_0),.clk(gclk));
	jdff dff_B_QJiujBaq8_0(.din(w_dff_B_syA4iOfo1_0),.dout(w_dff_B_QJiujBaq8_0),.clk(gclk));
	jdff dff_B_2FUlOjPf6_0(.din(w_dff_B_QJiujBaq8_0),.dout(w_dff_B_2FUlOjPf6_0),.clk(gclk));
	jdff dff_B_VBqk8ThL3_0(.din(w_dff_B_2FUlOjPf6_0),.dout(w_dff_B_VBqk8ThL3_0),.clk(gclk));
	jdff dff_B_TncV616K6_0(.din(w_dff_B_VBqk8ThL3_0),.dout(w_dff_B_TncV616K6_0),.clk(gclk));
	jdff dff_B_c5JrsnKV6_0(.din(w_dff_B_TncV616K6_0),.dout(w_dff_B_c5JrsnKV6_0),.clk(gclk));
	jdff dff_B_RbbPDLYO1_0(.din(w_dff_B_c5JrsnKV6_0),.dout(w_dff_B_RbbPDLYO1_0),.clk(gclk));
	jdff dff_B_kOGm8zEs9_0(.din(w_dff_B_RbbPDLYO1_0),.dout(w_dff_B_kOGm8zEs9_0),.clk(gclk));
	jdff dff_B_KBgZBmGc5_0(.din(w_dff_B_kOGm8zEs9_0),.dout(w_dff_B_KBgZBmGc5_0),.clk(gclk));
	jdff dff_B_ZtxR5PI36_0(.din(w_dff_B_KBgZBmGc5_0),.dout(w_dff_B_ZtxR5PI36_0),.clk(gclk));
	jdff dff_B_l6ocIsuX2_0(.din(w_dff_B_ZtxR5PI36_0),.dout(w_dff_B_l6ocIsuX2_0),.clk(gclk));
	jdff dff_B_eMlvmWyc5_0(.din(w_dff_B_l6ocIsuX2_0),.dout(w_dff_B_eMlvmWyc5_0),.clk(gclk));
	jdff dff_B_waAhaXlM4_0(.din(w_dff_B_eMlvmWyc5_0),.dout(w_dff_B_waAhaXlM4_0),.clk(gclk));
	jdff dff_B_yIo0sQNo8_0(.din(w_dff_B_waAhaXlM4_0),.dout(w_dff_B_yIo0sQNo8_0),.clk(gclk));
	jdff dff_B_Tjg5JjoQ5_0(.din(w_dff_B_yIo0sQNo8_0),.dout(w_dff_B_Tjg5JjoQ5_0),.clk(gclk));
	jdff dff_B_c3Num61Z6_0(.din(w_dff_B_Tjg5JjoQ5_0),.dout(w_dff_B_c3Num61Z6_0),.clk(gclk));
	jdff dff_B_RiUHyLMr8_0(.din(w_dff_B_c3Num61Z6_0),.dout(w_dff_B_RiUHyLMr8_0),.clk(gclk));
	jdff dff_B_t57R8BJk5_0(.din(w_dff_B_RiUHyLMr8_0),.dout(w_dff_B_t57R8BJk5_0),.clk(gclk));
	jdff dff_B_2tpIruTy5_0(.din(w_dff_B_t57R8BJk5_0),.dout(w_dff_B_2tpIruTy5_0),.clk(gclk));
	jdff dff_B_ZQKKpnKS0_1(.din(n930),.dout(w_dff_B_ZQKKpnKS0_1),.clk(gclk));
	jdff dff_B_hyvVoXDq5_1(.din(w_dff_B_ZQKKpnKS0_1),.dout(w_dff_B_hyvVoXDq5_1),.clk(gclk));
	jdff dff_B_2rlWrmKE8_1(.din(w_dff_B_hyvVoXDq5_1),.dout(w_dff_B_2rlWrmKE8_1),.clk(gclk));
	jdff dff_B_b77XAnMR0_1(.din(w_dff_B_2rlWrmKE8_1),.dout(w_dff_B_b77XAnMR0_1),.clk(gclk));
	jdff dff_B_XTx48BFZ6_1(.din(w_dff_B_b77XAnMR0_1),.dout(w_dff_B_XTx48BFZ6_1),.clk(gclk));
	jdff dff_B_qdXgJKKH5_1(.din(w_dff_B_XTx48BFZ6_1),.dout(w_dff_B_qdXgJKKH5_1),.clk(gclk));
	jdff dff_B_OeO1Wmeq0_1(.din(w_dff_B_qdXgJKKH5_1),.dout(w_dff_B_OeO1Wmeq0_1),.clk(gclk));
	jdff dff_B_TZxNTdXT0_1(.din(w_dff_B_OeO1Wmeq0_1),.dout(w_dff_B_TZxNTdXT0_1),.clk(gclk));
	jdff dff_B_i6woalFV3_1(.din(w_dff_B_TZxNTdXT0_1),.dout(w_dff_B_i6woalFV3_1),.clk(gclk));
	jdff dff_B_WQiHXRey7_1(.din(w_dff_B_i6woalFV3_1),.dout(w_dff_B_WQiHXRey7_1),.clk(gclk));
	jdff dff_B_eKpshZld5_1(.din(w_dff_B_WQiHXRey7_1),.dout(w_dff_B_eKpshZld5_1),.clk(gclk));
	jdff dff_B_rBhIkbGK4_1(.din(w_dff_B_eKpshZld5_1),.dout(w_dff_B_rBhIkbGK4_1),.clk(gclk));
	jdff dff_B_5AcocSIw2_1(.din(w_dff_B_rBhIkbGK4_1),.dout(w_dff_B_5AcocSIw2_1),.clk(gclk));
	jdff dff_B_upL5tNg77_1(.din(w_dff_B_5AcocSIw2_1),.dout(w_dff_B_upL5tNg77_1),.clk(gclk));
	jdff dff_B_hAwyS8Ed9_1(.din(w_dff_B_upL5tNg77_1),.dout(w_dff_B_hAwyS8Ed9_1),.clk(gclk));
	jdff dff_B_hMCqLxTx9_1(.din(w_dff_B_hAwyS8Ed9_1),.dout(w_dff_B_hMCqLxTx9_1),.clk(gclk));
	jdff dff_B_ABREldef9_1(.din(w_dff_B_hMCqLxTx9_1),.dout(w_dff_B_ABREldef9_1),.clk(gclk));
	jdff dff_B_Za16KxHz1_1(.din(w_dff_B_ABREldef9_1),.dout(w_dff_B_Za16KxHz1_1),.clk(gclk));
	jdff dff_B_g9BEGyV38_1(.din(w_dff_B_Za16KxHz1_1),.dout(w_dff_B_g9BEGyV38_1),.clk(gclk));
	jdff dff_B_q2dsZIkH5_1(.din(w_dff_B_g9BEGyV38_1),.dout(w_dff_B_q2dsZIkH5_1),.clk(gclk));
	jdff dff_B_HCkqZFVx7_1(.din(w_dff_B_q2dsZIkH5_1),.dout(w_dff_B_HCkqZFVx7_1),.clk(gclk));
	jdff dff_B_wuh39z5h0_1(.din(w_dff_B_HCkqZFVx7_1),.dout(w_dff_B_wuh39z5h0_1),.clk(gclk));
	jdff dff_B_KZVJ1Uil1_1(.din(w_dff_B_wuh39z5h0_1),.dout(w_dff_B_KZVJ1Uil1_1),.clk(gclk));
	jdff dff_B_BWpVNCCC2_1(.din(w_dff_B_KZVJ1Uil1_1),.dout(w_dff_B_BWpVNCCC2_1),.clk(gclk));
	jdff dff_B_DKdYYBA96_1(.din(w_dff_B_BWpVNCCC2_1),.dout(w_dff_B_DKdYYBA96_1),.clk(gclk));
	jdff dff_B_qwEHv9v82_1(.din(w_dff_B_DKdYYBA96_1),.dout(w_dff_B_qwEHv9v82_1),.clk(gclk));
	jdff dff_B_kTqFJaj26_1(.din(w_dff_B_qwEHv9v82_1),.dout(w_dff_B_kTqFJaj26_1),.clk(gclk));
	jdff dff_B_NOLA7Ut27_1(.din(w_dff_B_kTqFJaj26_1),.dout(w_dff_B_NOLA7Ut27_1),.clk(gclk));
	jdff dff_B_fsJEECv94_1(.din(w_dff_B_NOLA7Ut27_1),.dout(w_dff_B_fsJEECv94_1),.clk(gclk));
	jdff dff_B_LuYGpeAY1_1(.din(w_dff_B_fsJEECv94_1),.dout(w_dff_B_LuYGpeAY1_1),.clk(gclk));
	jdff dff_B_le184tYM0_1(.din(w_dff_B_LuYGpeAY1_1),.dout(w_dff_B_le184tYM0_1),.clk(gclk));
	jdff dff_B_T9eTpHAR9_1(.din(w_dff_B_le184tYM0_1),.dout(w_dff_B_T9eTpHAR9_1),.clk(gclk));
	jdff dff_B_uH14Dbid2_1(.din(w_dff_B_T9eTpHAR9_1),.dout(w_dff_B_uH14Dbid2_1),.clk(gclk));
	jdff dff_B_2Lkym8bN9_1(.din(w_dff_B_uH14Dbid2_1),.dout(w_dff_B_2Lkym8bN9_1),.clk(gclk));
	jdff dff_B_a9kFii4x0_1(.din(w_dff_B_2Lkym8bN9_1),.dout(w_dff_B_a9kFii4x0_1),.clk(gclk));
	jdff dff_B_lmmnAsfP6_1(.din(w_dff_B_a9kFii4x0_1),.dout(w_dff_B_lmmnAsfP6_1),.clk(gclk));
	jdff dff_B_EnxXsfQC6_1(.din(w_dff_B_lmmnAsfP6_1),.dout(w_dff_B_EnxXsfQC6_1),.clk(gclk));
	jdff dff_B_RVIrtoho8_1(.din(w_dff_B_EnxXsfQC6_1),.dout(w_dff_B_RVIrtoho8_1),.clk(gclk));
	jdff dff_B_V8mjDS7W3_1(.din(w_dff_B_RVIrtoho8_1),.dout(w_dff_B_V8mjDS7W3_1),.clk(gclk));
	jdff dff_B_jnQNt3aD2_1(.din(w_dff_B_V8mjDS7W3_1),.dout(w_dff_B_jnQNt3aD2_1),.clk(gclk));
	jdff dff_B_7gg0bx6b0_1(.din(w_dff_B_jnQNt3aD2_1),.dout(w_dff_B_7gg0bx6b0_1),.clk(gclk));
	jdff dff_B_JY0KhHLO8_1(.din(w_dff_B_7gg0bx6b0_1),.dout(w_dff_B_JY0KhHLO8_1),.clk(gclk));
	jdff dff_B_iLXZ0D6q2_1(.din(w_dff_B_JY0KhHLO8_1),.dout(w_dff_B_iLXZ0D6q2_1),.clk(gclk));
	jdff dff_B_FsLwiPBW3_1(.din(w_dff_B_iLXZ0D6q2_1),.dout(w_dff_B_FsLwiPBW3_1),.clk(gclk));
	jdff dff_B_loGaXOrq4_1(.din(w_dff_B_FsLwiPBW3_1),.dout(w_dff_B_loGaXOrq4_1),.clk(gclk));
	jdff dff_B_5aBw9nLi5_1(.din(w_dff_B_loGaXOrq4_1),.dout(w_dff_B_5aBw9nLi5_1),.clk(gclk));
	jdff dff_B_mZpK3axG0_1(.din(w_dff_B_5aBw9nLi5_1),.dout(w_dff_B_mZpK3axG0_1),.clk(gclk));
	jdff dff_B_XyRs4s4z3_1(.din(w_dff_B_mZpK3axG0_1),.dout(w_dff_B_XyRs4s4z3_1),.clk(gclk));
	jdff dff_B_ACmCXSDy4_1(.din(w_dff_B_XyRs4s4z3_1),.dout(w_dff_B_ACmCXSDy4_1),.clk(gclk));
	jdff dff_B_GJh7p58r5_1(.din(w_dff_B_ACmCXSDy4_1),.dout(w_dff_B_GJh7p58r5_1),.clk(gclk));
	jdff dff_B_2frT5aZ90_1(.din(w_dff_B_GJh7p58r5_1),.dout(w_dff_B_2frT5aZ90_1),.clk(gclk));
	jdff dff_B_KzN9yxYq6_1(.din(w_dff_B_2frT5aZ90_1),.dout(w_dff_B_KzN9yxYq6_1),.clk(gclk));
	jdff dff_B_AJZCYnvk9_1(.din(w_dff_B_KzN9yxYq6_1),.dout(w_dff_B_AJZCYnvk9_1),.clk(gclk));
	jdff dff_B_DbsOHvFM7_1(.din(w_dff_B_AJZCYnvk9_1),.dout(w_dff_B_DbsOHvFM7_1),.clk(gclk));
	jdff dff_B_BP6jGezL7_1(.din(w_dff_B_DbsOHvFM7_1),.dout(w_dff_B_BP6jGezL7_1),.clk(gclk));
	jdff dff_B_VamXzUl30_1(.din(w_dff_B_BP6jGezL7_1),.dout(w_dff_B_VamXzUl30_1),.clk(gclk));
	jdff dff_B_AWRB28MV2_1(.din(w_dff_B_VamXzUl30_1),.dout(w_dff_B_AWRB28MV2_1),.clk(gclk));
	jdff dff_B_5AjSqHfD8_1(.din(w_dff_B_AWRB28MV2_1),.dout(w_dff_B_5AjSqHfD8_1),.clk(gclk));
	jdff dff_B_9dV47HvI6_1(.din(w_dff_B_5AjSqHfD8_1),.dout(w_dff_B_9dV47HvI6_1),.clk(gclk));
	jdff dff_B_bOBWRJGc1_1(.din(w_dff_B_9dV47HvI6_1),.dout(w_dff_B_bOBWRJGc1_1),.clk(gclk));
	jdff dff_B_Mvp7oTsm1_1(.din(w_dff_B_bOBWRJGc1_1),.dout(w_dff_B_Mvp7oTsm1_1),.clk(gclk));
	jdff dff_B_bZJSGiR79_1(.din(w_dff_B_Mvp7oTsm1_1),.dout(w_dff_B_bZJSGiR79_1),.clk(gclk));
	jdff dff_B_Pfl3HMCX3_1(.din(w_dff_B_bZJSGiR79_1),.dout(w_dff_B_Pfl3HMCX3_1),.clk(gclk));
	jdff dff_B_UiKAMvgk0_1(.din(w_dff_B_Pfl3HMCX3_1),.dout(w_dff_B_UiKAMvgk0_1),.clk(gclk));
	jdff dff_B_dIa7nWvw1_1(.din(w_dff_B_UiKAMvgk0_1),.dout(w_dff_B_dIa7nWvw1_1),.clk(gclk));
	jdff dff_B_IG3ckOWe8_1(.din(w_dff_B_dIa7nWvw1_1),.dout(w_dff_B_IG3ckOWe8_1),.clk(gclk));
	jdff dff_B_8nE5qFnE0_1(.din(w_dff_B_IG3ckOWe8_1),.dout(w_dff_B_8nE5qFnE0_1),.clk(gclk));
	jdff dff_B_HL2xPlH74_1(.din(w_dff_B_8nE5qFnE0_1),.dout(w_dff_B_HL2xPlH74_1),.clk(gclk));
	jdff dff_B_mcEoyKTN6_1(.din(w_dff_B_HL2xPlH74_1),.dout(w_dff_B_mcEoyKTN6_1),.clk(gclk));
	jdff dff_B_oXFS6tjS9_1(.din(w_dff_B_mcEoyKTN6_1),.dout(w_dff_B_oXFS6tjS9_1),.clk(gclk));
	jdff dff_B_3Mi9Gsdu5_1(.din(w_dff_B_oXFS6tjS9_1),.dout(w_dff_B_3Mi9Gsdu5_1),.clk(gclk));
	jdff dff_B_ELejFTVp7_1(.din(w_dff_B_3Mi9Gsdu5_1),.dout(w_dff_B_ELejFTVp7_1),.clk(gclk));
	jdff dff_B_sn5Wp6Fr4_1(.din(w_dff_B_ELejFTVp7_1),.dout(w_dff_B_sn5Wp6Fr4_1),.clk(gclk));
	jdff dff_B_j8SCVz7e6_1(.din(w_dff_B_sn5Wp6Fr4_1),.dout(w_dff_B_j8SCVz7e6_1),.clk(gclk));
	jdff dff_B_VUiFq6jH9_1(.din(w_dff_B_j8SCVz7e6_1),.dout(w_dff_B_VUiFq6jH9_1),.clk(gclk));
	jdff dff_B_IxpQ1gpW4_1(.din(w_dff_B_VUiFq6jH9_1),.dout(w_dff_B_IxpQ1gpW4_1),.clk(gclk));
	jdff dff_B_MP9moO1H6_1(.din(w_dff_B_IxpQ1gpW4_1),.dout(w_dff_B_MP9moO1H6_1),.clk(gclk));
	jdff dff_B_CMYRLp6X7_1(.din(w_dff_B_MP9moO1H6_1),.dout(w_dff_B_CMYRLp6X7_1),.clk(gclk));
	jdff dff_B_uNurphcp6_1(.din(w_dff_B_CMYRLp6X7_1),.dout(w_dff_B_uNurphcp6_1),.clk(gclk));
	jdff dff_B_XktcUBUX7_1(.din(w_dff_B_uNurphcp6_1),.dout(w_dff_B_XktcUBUX7_1),.clk(gclk));
	jdff dff_B_iN8WgXyO6_1(.din(w_dff_B_XktcUBUX7_1),.dout(w_dff_B_iN8WgXyO6_1),.clk(gclk));
	jdff dff_B_3XjSxaxE6_1(.din(w_dff_B_iN8WgXyO6_1),.dout(w_dff_B_3XjSxaxE6_1),.clk(gclk));
	jdff dff_B_MlD79jp26_1(.din(w_dff_B_3XjSxaxE6_1),.dout(w_dff_B_MlD79jp26_1),.clk(gclk));
	jdff dff_B_bA6E01ro1_1(.din(w_dff_B_MlD79jp26_1),.dout(w_dff_B_bA6E01ro1_1),.clk(gclk));
	jdff dff_B_J5bPjCEh8_1(.din(w_dff_B_bA6E01ro1_1),.dout(w_dff_B_J5bPjCEh8_1),.clk(gclk));
	jdff dff_B_PKpGVWci4_1(.din(w_dff_B_J5bPjCEh8_1),.dout(w_dff_B_PKpGVWci4_1),.clk(gclk));
	jdff dff_B_b4Yyg7Wb8_1(.din(w_dff_B_PKpGVWci4_1),.dout(w_dff_B_b4Yyg7Wb8_1),.clk(gclk));
	jdff dff_B_y35aUNqV9_1(.din(w_dff_B_b4Yyg7Wb8_1),.dout(w_dff_B_y35aUNqV9_1),.clk(gclk));
	jdff dff_B_8Kymw5863_1(.din(w_dff_B_y35aUNqV9_1),.dout(w_dff_B_8Kymw5863_1),.clk(gclk));
	jdff dff_B_YvcDHCUq5_1(.din(w_dff_B_8Kymw5863_1),.dout(w_dff_B_YvcDHCUq5_1),.clk(gclk));
	jdff dff_B_eoY4eUdu5_1(.din(w_dff_B_YvcDHCUq5_1),.dout(w_dff_B_eoY4eUdu5_1),.clk(gclk));
	jdff dff_B_r6oiuFx05_0(.din(n931),.dout(w_dff_B_r6oiuFx05_0),.clk(gclk));
	jdff dff_B_2bawyn1r8_0(.din(w_dff_B_r6oiuFx05_0),.dout(w_dff_B_2bawyn1r8_0),.clk(gclk));
	jdff dff_B_ziqfpptT1_0(.din(w_dff_B_2bawyn1r8_0),.dout(w_dff_B_ziqfpptT1_0),.clk(gclk));
	jdff dff_B_37JprzNU9_0(.din(w_dff_B_ziqfpptT1_0),.dout(w_dff_B_37JprzNU9_0),.clk(gclk));
	jdff dff_B_akUv6lz74_0(.din(w_dff_B_37JprzNU9_0),.dout(w_dff_B_akUv6lz74_0),.clk(gclk));
	jdff dff_B_OGMDRS3F7_0(.din(w_dff_B_akUv6lz74_0),.dout(w_dff_B_OGMDRS3F7_0),.clk(gclk));
	jdff dff_B_UnjYyCk78_0(.din(w_dff_B_OGMDRS3F7_0),.dout(w_dff_B_UnjYyCk78_0),.clk(gclk));
	jdff dff_B_nhdnsPRK0_0(.din(w_dff_B_UnjYyCk78_0),.dout(w_dff_B_nhdnsPRK0_0),.clk(gclk));
	jdff dff_B_HQE5uNHq0_0(.din(w_dff_B_nhdnsPRK0_0),.dout(w_dff_B_HQE5uNHq0_0),.clk(gclk));
	jdff dff_B_HHmdn0UE9_0(.din(w_dff_B_HQE5uNHq0_0),.dout(w_dff_B_HHmdn0UE9_0),.clk(gclk));
	jdff dff_B_V6tFQHXl8_0(.din(w_dff_B_HHmdn0UE9_0),.dout(w_dff_B_V6tFQHXl8_0),.clk(gclk));
	jdff dff_B_nXVvsL5x3_0(.din(w_dff_B_V6tFQHXl8_0),.dout(w_dff_B_nXVvsL5x3_0),.clk(gclk));
	jdff dff_B_1wvDl6qs8_0(.din(w_dff_B_nXVvsL5x3_0),.dout(w_dff_B_1wvDl6qs8_0),.clk(gclk));
	jdff dff_B_ravbEzCR9_0(.din(w_dff_B_1wvDl6qs8_0),.dout(w_dff_B_ravbEzCR9_0),.clk(gclk));
	jdff dff_B_8KhRWNQ71_0(.din(w_dff_B_ravbEzCR9_0),.dout(w_dff_B_8KhRWNQ71_0),.clk(gclk));
	jdff dff_B_cyzAh48f6_0(.din(w_dff_B_8KhRWNQ71_0),.dout(w_dff_B_cyzAh48f6_0),.clk(gclk));
	jdff dff_B_s5e8FSEN1_0(.din(w_dff_B_cyzAh48f6_0),.dout(w_dff_B_s5e8FSEN1_0),.clk(gclk));
	jdff dff_B_mK1nylq38_0(.din(w_dff_B_s5e8FSEN1_0),.dout(w_dff_B_mK1nylq38_0),.clk(gclk));
	jdff dff_B_Um5pdJSm4_0(.din(w_dff_B_mK1nylq38_0),.dout(w_dff_B_Um5pdJSm4_0),.clk(gclk));
	jdff dff_B_oZzS8cBA7_0(.din(w_dff_B_Um5pdJSm4_0),.dout(w_dff_B_oZzS8cBA7_0),.clk(gclk));
	jdff dff_B_Rsw4HFE22_0(.din(w_dff_B_oZzS8cBA7_0),.dout(w_dff_B_Rsw4HFE22_0),.clk(gclk));
	jdff dff_B_FUtx1SPN0_0(.din(w_dff_B_Rsw4HFE22_0),.dout(w_dff_B_FUtx1SPN0_0),.clk(gclk));
	jdff dff_B_FJrcUHrM5_0(.din(w_dff_B_FUtx1SPN0_0),.dout(w_dff_B_FJrcUHrM5_0),.clk(gclk));
	jdff dff_B_qVH48R986_0(.din(w_dff_B_FJrcUHrM5_0),.dout(w_dff_B_qVH48R986_0),.clk(gclk));
	jdff dff_B_VKbE30s90_0(.din(w_dff_B_qVH48R986_0),.dout(w_dff_B_VKbE30s90_0),.clk(gclk));
	jdff dff_B_otbRIaFe2_0(.din(w_dff_B_VKbE30s90_0),.dout(w_dff_B_otbRIaFe2_0),.clk(gclk));
	jdff dff_B_oSXLY6E07_0(.din(w_dff_B_otbRIaFe2_0),.dout(w_dff_B_oSXLY6E07_0),.clk(gclk));
	jdff dff_B_XEENkSAO6_0(.din(w_dff_B_oSXLY6E07_0),.dout(w_dff_B_XEENkSAO6_0),.clk(gclk));
	jdff dff_B_9avH78Dr5_0(.din(w_dff_B_XEENkSAO6_0),.dout(w_dff_B_9avH78Dr5_0),.clk(gclk));
	jdff dff_B_SwwZKrUg8_0(.din(w_dff_B_9avH78Dr5_0),.dout(w_dff_B_SwwZKrUg8_0),.clk(gclk));
	jdff dff_B_Dzixfz0g7_0(.din(w_dff_B_SwwZKrUg8_0),.dout(w_dff_B_Dzixfz0g7_0),.clk(gclk));
	jdff dff_B_jYBkZqFp1_0(.din(w_dff_B_Dzixfz0g7_0),.dout(w_dff_B_jYBkZqFp1_0),.clk(gclk));
	jdff dff_B_DHIPo0I45_0(.din(w_dff_B_jYBkZqFp1_0),.dout(w_dff_B_DHIPo0I45_0),.clk(gclk));
	jdff dff_B_wx8zFKNI8_0(.din(w_dff_B_DHIPo0I45_0),.dout(w_dff_B_wx8zFKNI8_0),.clk(gclk));
	jdff dff_B_PmlhirSB8_0(.din(w_dff_B_wx8zFKNI8_0),.dout(w_dff_B_PmlhirSB8_0),.clk(gclk));
	jdff dff_B_6RWenhc93_0(.din(w_dff_B_PmlhirSB8_0),.dout(w_dff_B_6RWenhc93_0),.clk(gclk));
	jdff dff_B_mzqpiX8W6_0(.din(w_dff_B_6RWenhc93_0),.dout(w_dff_B_mzqpiX8W6_0),.clk(gclk));
	jdff dff_B_PjwitYUW4_0(.din(w_dff_B_mzqpiX8W6_0),.dout(w_dff_B_PjwitYUW4_0),.clk(gclk));
	jdff dff_B_nYfbVR5P4_0(.din(w_dff_B_PjwitYUW4_0),.dout(w_dff_B_nYfbVR5P4_0),.clk(gclk));
	jdff dff_B_ud0NlXKT4_0(.din(w_dff_B_nYfbVR5P4_0),.dout(w_dff_B_ud0NlXKT4_0),.clk(gclk));
	jdff dff_B_hR6qfRFe9_0(.din(w_dff_B_ud0NlXKT4_0),.dout(w_dff_B_hR6qfRFe9_0),.clk(gclk));
	jdff dff_B_ojaHAo0n5_0(.din(w_dff_B_hR6qfRFe9_0),.dout(w_dff_B_ojaHAo0n5_0),.clk(gclk));
	jdff dff_B_iIXUgi9K5_0(.din(w_dff_B_ojaHAo0n5_0),.dout(w_dff_B_iIXUgi9K5_0),.clk(gclk));
	jdff dff_B_RQfKjI439_0(.din(w_dff_B_iIXUgi9K5_0),.dout(w_dff_B_RQfKjI439_0),.clk(gclk));
	jdff dff_B_a8ZPmP1q9_0(.din(w_dff_B_RQfKjI439_0),.dout(w_dff_B_a8ZPmP1q9_0),.clk(gclk));
	jdff dff_B_7zFFgnua2_0(.din(w_dff_B_a8ZPmP1q9_0),.dout(w_dff_B_7zFFgnua2_0),.clk(gclk));
	jdff dff_B_7gxoReoM7_0(.din(w_dff_B_7zFFgnua2_0),.dout(w_dff_B_7gxoReoM7_0),.clk(gclk));
	jdff dff_B_8cXdFcyZ5_0(.din(w_dff_B_7gxoReoM7_0),.dout(w_dff_B_8cXdFcyZ5_0),.clk(gclk));
	jdff dff_B_oaQ0FsZ10_0(.din(w_dff_B_8cXdFcyZ5_0),.dout(w_dff_B_oaQ0FsZ10_0),.clk(gclk));
	jdff dff_B_oZvnS2510_0(.din(w_dff_B_oaQ0FsZ10_0),.dout(w_dff_B_oZvnS2510_0),.clk(gclk));
	jdff dff_B_EXC8SVu56_0(.din(w_dff_B_oZvnS2510_0),.dout(w_dff_B_EXC8SVu56_0),.clk(gclk));
	jdff dff_B_2PcolzLq4_0(.din(w_dff_B_EXC8SVu56_0),.dout(w_dff_B_2PcolzLq4_0),.clk(gclk));
	jdff dff_B_LDhGuWmx4_0(.din(w_dff_B_2PcolzLq4_0),.dout(w_dff_B_LDhGuWmx4_0),.clk(gclk));
	jdff dff_B_M4qapaot3_0(.din(w_dff_B_LDhGuWmx4_0),.dout(w_dff_B_M4qapaot3_0),.clk(gclk));
	jdff dff_B_pCRKaWQa6_0(.din(w_dff_B_M4qapaot3_0),.dout(w_dff_B_pCRKaWQa6_0),.clk(gclk));
	jdff dff_B_QD9euuLG9_0(.din(w_dff_B_pCRKaWQa6_0),.dout(w_dff_B_QD9euuLG9_0),.clk(gclk));
	jdff dff_B_a88WwJJP7_0(.din(w_dff_B_QD9euuLG9_0),.dout(w_dff_B_a88WwJJP7_0),.clk(gclk));
	jdff dff_B_9iyKrfid3_0(.din(w_dff_B_a88WwJJP7_0),.dout(w_dff_B_9iyKrfid3_0),.clk(gclk));
	jdff dff_B_4HyRwzR37_0(.din(w_dff_B_9iyKrfid3_0),.dout(w_dff_B_4HyRwzR37_0),.clk(gclk));
	jdff dff_B_EaD88TUA8_0(.din(w_dff_B_4HyRwzR37_0),.dout(w_dff_B_EaD88TUA8_0),.clk(gclk));
	jdff dff_B_r4dh04yK0_0(.din(w_dff_B_EaD88TUA8_0),.dout(w_dff_B_r4dh04yK0_0),.clk(gclk));
	jdff dff_B_wqR3NJMA7_0(.din(w_dff_B_r4dh04yK0_0),.dout(w_dff_B_wqR3NJMA7_0),.clk(gclk));
	jdff dff_B_Qnjbbc5T4_0(.din(w_dff_B_wqR3NJMA7_0),.dout(w_dff_B_Qnjbbc5T4_0),.clk(gclk));
	jdff dff_B_C0f42nzF8_0(.din(w_dff_B_Qnjbbc5T4_0),.dout(w_dff_B_C0f42nzF8_0),.clk(gclk));
	jdff dff_B_lo9QwvLM4_0(.din(w_dff_B_C0f42nzF8_0),.dout(w_dff_B_lo9QwvLM4_0),.clk(gclk));
	jdff dff_B_vTH0mWKG9_0(.din(w_dff_B_lo9QwvLM4_0),.dout(w_dff_B_vTH0mWKG9_0),.clk(gclk));
	jdff dff_B_Kt6wot8k7_0(.din(w_dff_B_vTH0mWKG9_0),.dout(w_dff_B_Kt6wot8k7_0),.clk(gclk));
	jdff dff_B_epyffjIx6_0(.din(w_dff_B_Kt6wot8k7_0),.dout(w_dff_B_epyffjIx6_0),.clk(gclk));
	jdff dff_B_wm3QBzfu2_0(.din(w_dff_B_epyffjIx6_0),.dout(w_dff_B_wm3QBzfu2_0),.clk(gclk));
	jdff dff_B_umGt7O0q9_0(.din(w_dff_B_wm3QBzfu2_0),.dout(w_dff_B_umGt7O0q9_0),.clk(gclk));
	jdff dff_B_UngqZoyv3_0(.din(w_dff_B_umGt7O0q9_0),.dout(w_dff_B_UngqZoyv3_0),.clk(gclk));
	jdff dff_B_l87SoIcI6_0(.din(w_dff_B_UngqZoyv3_0),.dout(w_dff_B_l87SoIcI6_0),.clk(gclk));
	jdff dff_B_oVjMHjQe7_0(.din(w_dff_B_l87SoIcI6_0),.dout(w_dff_B_oVjMHjQe7_0),.clk(gclk));
	jdff dff_B_63sWTRei1_0(.din(w_dff_B_oVjMHjQe7_0),.dout(w_dff_B_63sWTRei1_0),.clk(gclk));
	jdff dff_B_SkGqrsQ32_0(.din(w_dff_B_63sWTRei1_0),.dout(w_dff_B_SkGqrsQ32_0),.clk(gclk));
	jdff dff_B_1f1zlaui2_0(.din(w_dff_B_SkGqrsQ32_0),.dout(w_dff_B_1f1zlaui2_0),.clk(gclk));
	jdff dff_B_VhcQO4xz5_0(.din(w_dff_B_1f1zlaui2_0),.dout(w_dff_B_VhcQO4xz5_0),.clk(gclk));
	jdff dff_B_XpQCptHj0_0(.din(w_dff_B_VhcQO4xz5_0),.dout(w_dff_B_XpQCptHj0_0),.clk(gclk));
	jdff dff_B_UCouXUMV6_0(.din(w_dff_B_XpQCptHj0_0),.dout(w_dff_B_UCouXUMV6_0),.clk(gclk));
	jdff dff_B_dpDwdH1y6_0(.din(w_dff_B_UCouXUMV6_0),.dout(w_dff_B_dpDwdH1y6_0),.clk(gclk));
	jdff dff_B_nOwIypRd1_0(.din(w_dff_B_dpDwdH1y6_0),.dout(w_dff_B_nOwIypRd1_0),.clk(gclk));
	jdff dff_B_2ACqmBer0_0(.din(w_dff_B_nOwIypRd1_0),.dout(w_dff_B_2ACqmBer0_0),.clk(gclk));
	jdff dff_B_sLkbvnto5_0(.din(w_dff_B_2ACqmBer0_0),.dout(w_dff_B_sLkbvnto5_0),.clk(gclk));
	jdff dff_B_0fb6EK129_0(.din(w_dff_B_sLkbvnto5_0),.dout(w_dff_B_0fb6EK129_0),.clk(gclk));
	jdff dff_B_LJfbNuao1_0(.din(w_dff_B_0fb6EK129_0),.dout(w_dff_B_LJfbNuao1_0),.clk(gclk));
	jdff dff_B_QaEH5rye9_0(.din(w_dff_B_LJfbNuao1_0),.dout(w_dff_B_QaEH5rye9_0),.clk(gclk));
	jdff dff_B_aldOUR2M3_0(.din(w_dff_B_QaEH5rye9_0),.dout(w_dff_B_aldOUR2M3_0),.clk(gclk));
	jdff dff_B_E5Shiag94_0(.din(w_dff_B_aldOUR2M3_0),.dout(w_dff_B_E5Shiag94_0),.clk(gclk));
	jdff dff_B_iHxN2qeg1_0(.din(w_dff_B_E5Shiag94_0),.dout(w_dff_B_iHxN2qeg1_0),.clk(gclk));
	jdff dff_B_uiXlNlYP1_0(.din(w_dff_B_iHxN2qeg1_0),.dout(w_dff_B_uiXlNlYP1_0),.clk(gclk));
	jdff dff_B_yQ9eGirj0_0(.din(w_dff_B_uiXlNlYP1_0),.dout(w_dff_B_yQ9eGirj0_0),.clk(gclk));
	jdff dff_B_se6uw62Z3_1(.din(n924),.dout(w_dff_B_se6uw62Z3_1),.clk(gclk));
	jdff dff_B_YDFTS4SQ8_1(.din(w_dff_B_se6uw62Z3_1),.dout(w_dff_B_YDFTS4SQ8_1),.clk(gclk));
	jdff dff_B_cpUYpy5L2_1(.din(w_dff_B_YDFTS4SQ8_1),.dout(w_dff_B_cpUYpy5L2_1),.clk(gclk));
	jdff dff_B_At484BH01_1(.din(w_dff_B_cpUYpy5L2_1),.dout(w_dff_B_At484BH01_1),.clk(gclk));
	jdff dff_B_TwSipUUb6_1(.din(w_dff_B_At484BH01_1),.dout(w_dff_B_TwSipUUb6_1),.clk(gclk));
	jdff dff_B_442PVjyk4_1(.din(w_dff_B_TwSipUUb6_1),.dout(w_dff_B_442PVjyk4_1),.clk(gclk));
	jdff dff_B_VeLr0Mw59_1(.din(w_dff_B_442PVjyk4_1),.dout(w_dff_B_VeLr0Mw59_1),.clk(gclk));
	jdff dff_B_LxYosw3b0_1(.din(w_dff_B_VeLr0Mw59_1),.dout(w_dff_B_LxYosw3b0_1),.clk(gclk));
	jdff dff_B_fiyfH08J3_1(.din(w_dff_B_LxYosw3b0_1),.dout(w_dff_B_fiyfH08J3_1),.clk(gclk));
	jdff dff_B_pg9ajxEX1_1(.din(w_dff_B_fiyfH08J3_1),.dout(w_dff_B_pg9ajxEX1_1),.clk(gclk));
	jdff dff_B_BHOL2XNv4_1(.din(w_dff_B_pg9ajxEX1_1),.dout(w_dff_B_BHOL2XNv4_1),.clk(gclk));
	jdff dff_B_Dnw9AESR8_1(.din(w_dff_B_BHOL2XNv4_1),.dout(w_dff_B_Dnw9AESR8_1),.clk(gclk));
	jdff dff_B_vuaxBBiN0_1(.din(w_dff_B_Dnw9AESR8_1),.dout(w_dff_B_vuaxBBiN0_1),.clk(gclk));
	jdff dff_B_fm1ljZqU0_1(.din(w_dff_B_vuaxBBiN0_1),.dout(w_dff_B_fm1ljZqU0_1),.clk(gclk));
	jdff dff_B_Pi1MUNvl8_1(.din(w_dff_B_fm1ljZqU0_1),.dout(w_dff_B_Pi1MUNvl8_1),.clk(gclk));
	jdff dff_B_xiWacX7r8_1(.din(w_dff_B_Pi1MUNvl8_1),.dout(w_dff_B_xiWacX7r8_1),.clk(gclk));
	jdff dff_B_ZmshhO0M4_1(.din(w_dff_B_xiWacX7r8_1),.dout(w_dff_B_ZmshhO0M4_1),.clk(gclk));
	jdff dff_B_2RM2zhVA6_1(.din(w_dff_B_ZmshhO0M4_1),.dout(w_dff_B_2RM2zhVA6_1),.clk(gclk));
	jdff dff_B_aadhiS0u7_1(.din(w_dff_B_2RM2zhVA6_1),.dout(w_dff_B_aadhiS0u7_1),.clk(gclk));
	jdff dff_B_ODs7ZHdc9_1(.din(w_dff_B_aadhiS0u7_1),.dout(w_dff_B_ODs7ZHdc9_1),.clk(gclk));
	jdff dff_B_uuTht2yX7_1(.din(w_dff_B_ODs7ZHdc9_1),.dout(w_dff_B_uuTht2yX7_1),.clk(gclk));
	jdff dff_B_8PNwltkp0_1(.din(w_dff_B_uuTht2yX7_1),.dout(w_dff_B_8PNwltkp0_1),.clk(gclk));
	jdff dff_B_UagfwMXB8_1(.din(w_dff_B_8PNwltkp0_1),.dout(w_dff_B_UagfwMXB8_1),.clk(gclk));
	jdff dff_B_N9UWKVbL3_1(.din(w_dff_B_UagfwMXB8_1),.dout(w_dff_B_N9UWKVbL3_1),.clk(gclk));
	jdff dff_B_UenmgPv27_1(.din(w_dff_B_N9UWKVbL3_1),.dout(w_dff_B_UenmgPv27_1),.clk(gclk));
	jdff dff_B_l8eCAZ7q8_1(.din(w_dff_B_UenmgPv27_1),.dout(w_dff_B_l8eCAZ7q8_1),.clk(gclk));
	jdff dff_B_e4SZfojh6_1(.din(w_dff_B_l8eCAZ7q8_1),.dout(w_dff_B_e4SZfojh6_1),.clk(gclk));
	jdff dff_B_MahyBmm61_1(.din(w_dff_B_e4SZfojh6_1),.dout(w_dff_B_MahyBmm61_1),.clk(gclk));
	jdff dff_B_poG3bfMf7_1(.din(w_dff_B_MahyBmm61_1),.dout(w_dff_B_poG3bfMf7_1),.clk(gclk));
	jdff dff_B_hXyV80Eh8_1(.din(w_dff_B_poG3bfMf7_1),.dout(w_dff_B_hXyV80Eh8_1),.clk(gclk));
	jdff dff_B_96Y8Y0Xn7_1(.din(w_dff_B_hXyV80Eh8_1),.dout(w_dff_B_96Y8Y0Xn7_1),.clk(gclk));
	jdff dff_B_u8LgfXdD4_1(.din(w_dff_B_96Y8Y0Xn7_1),.dout(w_dff_B_u8LgfXdD4_1),.clk(gclk));
	jdff dff_B_YZrnAZso7_1(.din(w_dff_B_u8LgfXdD4_1),.dout(w_dff_B_YZrnAZso7_1),.clk(gclk));
	jdff dff_B_6q36HsiP7_1(.din(w_dff_B_YZrnAZso7_1),.dout(w_dff_B_6q36HsiP7_1),.clk(gclk));
	jdff dff_B_gfBpOPU05_1(.din(w_dff_B_6q36HsiP7_1),.dout(w_dff_B_gfBpOPU05_1),.clk(gclk));
	jdff dff_B_ayQVFRgc6_1(.din(w_dff_B_gfBpOPU05_1),.dout(w_dff_B_ayQVFRgc6_1),.clk(gclk));
	jdff dff_B_D7Bq0hXG9_1(.din(w_dff_B_ayQVFRgc6_1),.dout(w_dff_B_D7Bq0hXG9_1),.clk(gclk));
	jdff dff_B_RAqRx4YC3_1(.din(w_dff_B_D7Bq0hXG9_1),.dout(w_dff_B_RAqRx4YC3_1),.clk(gclk));
	jdff dff_B_rrTAiO973_1(.din(w_dff_B_RAqRx4YC3_1),.dout(w_dff_B_rrTAiO973_1),.clk(gclk));
	jdff dff_B_PdmRQyhx4_1(.din(w_dff_B_rrTAiO973_1),.dout(w_dff_B_PdmRQyhx4_1),.clk(gclk));
	jdff dff_B_jlTdkK9s5_1(.din(w_dff_B_PdmRQyhx4_1),.dout(w_dff_B_jlTdkK9s5_1),.clk(gclk));
	jdff dff_B_q6r7xMLt3_1(.din(w_dff_B_jlTdkK9s5_1),.dout(w_dff_B_q6r7xMLt3_1),.clk(gclk));
	jdff dff_B_v7cnN4s29_1(.din(w_dff_B_q6r7xMLt3_1),.dout(w_dff_B_v7cnN4s29_1),.clk(gclk));
	jdff dff_B_SX529mAj1_1(.din(w_dff_B_v7cnN4s29_1),.dout(w_dff_B_SX529mAj1_1),.clk(gclk));
	jdff dff_B_girElLVg7_1(.din(w_dff_B_SX529mAj1_1),.dout(w_dff_B_girElLVg7_1),.clk(gclk));
	jdff dff_B_4016CAJ11_1(.din(w_dff_B_girElLVg7_1),.dout(w_dff_B_4016CAJ11_1),.clk(gclk));
	jdff dff_B_cMLBt9kp1_1(.din(w_dff_B_4016CAJ11_1),.dout(w_dff_B_cMLBt9kp1_1),.clk(gclk));
	jdff dff_B_uLTtgTGu2_1(.din(w_dff_B_cMLBt9kp1_1),.dout(w_dff_B_uLTtgTGu2_1),.clk(gclk));
	jdff dff_B_zF8Wz0fX8_1(.din(w_dff_B_uLTtgTGu2_1),.dout(w_dff_B_zF8Wz0fX8_1),.clk(gclk));
	jdff dff_B_DzR02vbf7_1(.din(w_dff_B_zF8Wz0fX8_1),.dout(w_dff_B_DzR02vbf7_1),.clk(gclk));
	jdff dff_B_EsGhCumm9_1(.din(w_dff_B_DzR02vbf7_1),.dout(w_dff_B_EsGhCumm9_1),.clk(gclk));
	jdff dff_B_tyTJrobg6_1(.din(w_dff_B_EsGhCumm9_1),.dout(w_dff_B_tyTJrobg6_1),.clk(gclk));
	jdff dff_B_xZ1dsy4Y4_1(.din(w_dff_B_tyTJrobg6_1),.dout(w_dff_B_xZ1dsy4Y4_1),.clk(gclk));
	jdff dff_B_0rzug1X50_1(.din(w_dff_B_xZ1dsy4Y4_1),.dout(w_dff_B_0rzug1X50_1),.clk(gclk));
	jdff dff_B_9yUdXD7Q0_1(.din(w_dff_B_0rzug1X50_1),.dout(w_dff_B_9yUdXD7Q0_1),.clk(gclk));
	jdff dff_B_P6ZBZUna8_1(.din(w_dff_B_9yUdXD7Q0_1),.dout(w_dff_B_P6ZBZUna8_1),.clk(gclk));
	jdff dff_B_ehxFBoAy6_1(.din(w_dff_B_P6ZBZUna8_1),.dout(w_dff_B_ehxFBoAy6_1),.clk(gclk));
	jdff dff_B_O6uoHPkp0_1(.din(w_dff_B_ehxFBoAy6_1),.dout(w_dff_B_O6uoHPkp0_1),.clk(gclk));
	jdff dff_B_KXCWaXlA1_1(.din(w_dff_B_O6uoHPkp0_1),.dout(w_dff_B_KXCWaXlA1_1),.clk(gclk));
	jdff dff_B_h5SArAYA8_1(.din(w_dff_B_KXCWaXlA1_1),.dout(w_dff_B_h5SArAYA8_1),.clk(gclk));
	jdff dff_B_67xymoO71_1(.din(w_dff_B_h5SArAYA8_1),.dout(w_dff_B_67xymoO71_1),.clk(gclk));
	jdff dff_B_fhEPmXiH3_1(.din(w_dff_B_67xymoO71_1),.dout(w_dff_B_fhEPmXiH3_1),.clk(gclk));
	jdff dff_B_dTsEZXC33_1(.din(w_dff_B_fhEPmXiH3_1),.dout(w_dff_B_dTsEZXC33_1),.clk(gclk));
	jdff dff_B_yogbt60R8_1(.din(w_dff_B_dTsEZXC33_1),.dout(w_dff_B_yogbt60R8_1),.clk(gclk));
	jdff dff_B_9EkWQFFq8_1(.din(w_dff_B_yogbt60R8_1),.dout(w_dff_B_9EkWQFFq8_1),.clk(gclk));
	jdff dff_B_gAaNQ4jQ3_1(.din(w_dff_B_9EkWQFFq8_1),.dout(w_dff_B_gAaNQ4jQ3_1),.clk(gclk));
	jdff dff_B_Ab1nIuMG4_1(.din(w_dff_B_gAaNQ4jQ3_1),.dout(w_dff_B_Ab1nIuMG4_1),.clk(gclk));
	jdff dff_B_xfIxl0zk7_1(.din(w_dff_B_Ab1nIuMG4_1),.dout(w_dff_B_xfIxl0zk7_1),.clk(gclk));
	jdff dff_B_T7EngNF43_1(.din(w_dff_B_xfIxl0zk7_1),.dout(w_dff_B_T7EngNF43_1),.clk(gclk));
	jdff dff_B_Z4x5vGIF6_1(.din(w_dff_B_T7EngNF43_1),.dout(w_dff_B_Z4x5vGIF6_1),.clk(gclk));
	jdff dff_B_mSYnoF7c0_1(.din(w_dff_B_Z4x5vGIF6_1),.dout(w_dff_B_mSYnoF7c0_1),.clk(gclk));
	jdff dff_B_eMqWX1mv4_1(.din(w_dff_B_mSYnoF7c0_1),.dout(w_dff_B_eMqWX1mv4_1),.clk(gclk));
	jdff dff_B_2j8yGB2t7_1(.din(w_dff_B_eMqWX1mv4_1),.dout(w_dff_B_2j8yGB2t7_1),.clk(gclk));
	jdff dff_B_oBGuM9CJ9_1(.din(w_dff_B_2j8yGB2t7_1),.dout(w_dff_B_oBGuM9CJ9_1),.clk(gclk));
	jdff dff_B_xjNVOoN11_1(.din(w_dff_B_oBGuM9CJ9_1),.dout(w_dff_B_xjNVOoN11_1),.clk(gclk));
	jdff dff_B_V0t9D08C8_1(.din(w_dff_B_xjNVOoN11_1),.dout(w_dff_B_V0t9D08C8_1),.clk(gclk));
	jdff dff_B_u67vymPe9_1(.din(w_dff_B_V0t9D08C8_1),.dout(w_dff_B_u67vymPe9_1),.clk(gclk));
	jdff dff_B_uEGT0HKF9_1(.din(w_dff_B_u67vymPe9_1),.dout(w_dff_B_uEGT0HKF9_1),.clk(gclk));
	jdff dff_B_bwbXM5zf9_1(.din(w_dff_B_uEGT0HKF9_1),.dout(w_dff_B_bwbXM5zf9_1),.clk(gclk));
	jdff dff_B_vPk5cKqa5_1(.din(w_dff_B_bwbXM5zf9_1),.dout(w_dff_B_vPk5cKqa5_1),.clk(gclk));
	jdff dff_B_ENDknJRO4_1(.din(w_dff_B_vPk5cKqa5_1),.dout(w_dff_B_ENDknJRO4_1),.clk(gclk));
	jdff dff_B_AoiiewfB8_1(.din(w_dff_B_ENDknJRO4_1),.dout(w_dff_B_AoiiewfB8_1),.clk(gclk));
	jdff dff_B_aXE0BQV53_1(.din(w_dff_B_AoiiewfB8_1),.dout(w_dff_B_aXE0BQV53_1),.clk(gclk));
	jdff dff_B_rhDmmGVz7_1(.din(w_dff_B_aXE0BQV53_1),.dout(w_dff_B_rhDmmGVz7_1),.clk(gclk));
	jdff dff_B_9Ny2l7y05_1(.din(w_dff_B_rhDmmGVz7_1),.dout(w_dff_B_9Ny2l7y05_1),.clk(gclk));
	jdff dff_B_MR3g1Rmd9_1(.din(w_dff_B_9Ny2l7y05_1),.dout(w_dff_B_MR3g1Rmd9_1),.clk(gclk));
	jdff dff_B_GJxbffZN1_1(.din(w_dff_B_MR3g1Rmd9_1),.dout(w_dff_B_GJxbffZN1_1),.clk(gclk));
	jdff dff_B_VrVeXKav6_1(.din(w_dff_B_GJxbffZN1_1),.dout(w_dff_B_VrVeXKav6_1),.clk(gclk));
	jdff dff_B_QhDgwt0p3_1(.din(w_dff_B_VrVeXKav6_1),.dout(w_dff_B_QhDgwt0p3_1),.clk(gclk));
	jdff dff_B_8T9xx6qV1_1(.din(w_dff_B_QhDgwt0p3_1),.dout(w_dff_B_8T9xx6qV1_1),.clk(gclk));
	jdff dff_B_9TIwEGfL8_0(.din(n925),.dout(w_dff_B_9TIwEGfL8_0),.clk(gclk));
	jdff dff_B_sIteoKyL8_0(.din(w_dff_B_9TIwEGfL8_0),.dout(w_dff_B_sIteoKyL8_0),.clk(gclk));
	jdff dff_B_00Epb6yB9_0(.din(w_dff_B_sIteoKyL8_0),.dout(w_dff_B_00Epb6yB9_0),.clk(gclk));
	jdff dff_B_tk6ZurhK2_0(.din(w_dff_B_00Epb6yB9_0),.dout(w_dff_B_tk6ZurhK2_0),.clk(gclk));
	jdff dff_B_TDPGJW6W9_0(.din(w_dff_B_tk6ZurhK2_0),.dout(w_dff_B_TDPGJW6W9_0),.clk(gclk));
	jdff dff_B_r0bZlsZ27_0(.din(w_dff_B_TDPGJW6W9_0),.dout(w_dff_B_r0bZlsZ27_0),.clk(gclk));
	jdff dff_B_P55q99eh7_0(.din(w_dff_B_r0bZlsZ27_0),.dout(w_dff_B_P55q99eh7_0),.clk(gclk));
	jdff dff_B_qOMxUOQB0_0(.din(w_dff_B_P55q99eh7_0),.dout(w_dff_B_qOMxUOQB0_0),.clk(gclk));
	jdff dff_B_GA7N7gGi1_0(.din(w_dff_B_qOMxUOQB0_0),.dout(w_dff_B_GA7N7gGi1_0),.clk(gclk));
	jdff dff_B_KM0OfOSB7_0(.din(w_dff_B_GA7N7gGi1_0),.dout(w_dff_B_KM0OfOSB7_0),.clk(gclk));
	jdff dff_B_63mw0JeE4_0(.din(w_dff_B_KM0OfOSB7_0),.dout(w_dff_B_63mw0JeE4_0),.clk(gclk));
	jdff dff_B_CeIS1ebV3_0(.din(w_dff_B_63mw0JeE4_0),.dout(w_dff_B_CeIS1ebV3_0),.clk(gclk));
	jdff dff_B_ZuLkiFml4_0(.din(w_dff_B_CeIS1ebV3_0),.dout(w_dff_B_ZuLkiFml4_0),.clk(gclk));
	jdff dff_B_CUCnWHdZ8_0(.din(w_dff_B_ZuLkiFml4_0),.dout(w_dff_B_CUCnWHdZ8_0),.clk(gclk));
	jdff dff_B_UImQlz6O0_0(.din(w_dff_B_CUCnWHdZ8_0),.dout(w_dff_B_UImQlz6O0_0),.clk(gclk));
	jdff dff_B_RnKs8BBT4_0(.din(w_dff_B_UImQlz6O0_0),.dout(w_dff_B_RnKs8BBT4_0),.clk(gclk));
	jdff dff_B_XrGY9wZF1_0(.din(w_dff_B_RnKs8BBT4_0),.dout(w_dff_B_XrGY9wZF1_0),.clk(gclk));
	jdff dff_B_D7Gg0IyA5_0(.din(w_dff_B_XrGY9wZF1_0),.dout(w_dff_B_D7Gg0IyA5_0),.clk(gclk));
	jdff dff_B_RyOQ2TAX1_0(.din(w_dff_B_D7Gg0IyA5_0),.dout(w_dff_B_RyOQ2TAX1_0),.clk(gclk));
	jdff dff_B_Ud0Mwmln4_0(.din(w_dff_B_RyOQ2TAX1_0),.dout(w_dff_B_Ud0Mwmln4_0),.clk(gclk));
	jdff dff_B_Qi56saku0_0(.din(w_dff_B_Ud0Mwmln4_0),.dout(w_dff_B_Qi56saku0_0),.clk(gclk));
	jdff dff_B_dM2qqaU35_0(.din(w_dff_B_Qi56saku0_0),.dout(w_dff_B_dM2qqaU35_0),.clk(gclk));
	jdff dff_B_cW5EmClX9_0(.din(w_dff_B_dM2qqaU35_0),.dout(w_dff_B_cW5EmClX9_0),.clk(gclk));
	jdff dff_B_jn3TTuLa2_0(.din(w_dff_B_cW5EmClX9_0),.dout(w_dff_B_jn3TTuLa2_0),.clk(gclk));
	jdff dff_B_ME6W3FR53_0(.din(w_dff_B_jn3TTuLa2_0),.dout(w_dff_B_ME6W3FR53_0),.clk(gclk));
	jdff dff_B_fGtxDOeT3_0(.din(w_dff_B_ME6W3FR53_0),.dout(w_dff_B_fGtxDOeT3_0),.clk(gclk));
	jdff dff_B_Yl4aPK3S6_0(.din(w_dff_B_fGtxDOeT3_0),.dout(w_dff_B_Yl4aPK3S6_0),.clk(gclk));
	jdff dff_B_LQGJATPE7_0(.din(w_dff_B_Yl4aPK3S6_0),.dout(w_dff_B_LQGJATPE7_0),.clk(gclk));
	jdff dff_B_zgYswCqo8_0(.din(w_dff_B_LQGJATPE7_0),.dout(w_dff_B_zgYswCqo8_0),.clk(gclk));
	jdff dff_B_qJVr2lAM9_0(.din(w_dff_B_zgYswCqo8_0),.dout(w_dff_B_qJVr2lAM9_0),.clk(gclk));
	jdff dff_B_iKbkbYNq5_0(.din(w_dff_B_qJVr2lAM9_0),.dout(w_dff_B_iKbkbYNq5_0),.clk(gclk));
	jdff dff_B_wbbMIOMZ0_0(.din(w_dff_B_iKbkbYNq5_0),.dout(w_dff_B_wbbMIOMZ0_0),.clk(gclk));
	jdff dff_B_qK2JSXFx0_0(.din(w_dff_B_wbbMIOMZ0_0),.dout(w_dff_B_qK2JSXFx0_0),.clk(gclk));
	jdff dff_B_0ENvKeQX2_0(.din(w_dff_B_qK2JSXFx0_0),.dout(w_dff_B_0ENvKeQX2_0),.clk(gclk));
	jdff dff_B_2nv5Y9tz5_0(.din(w_dff_B_0ENvKeQX2_0),.dout(w_dff_B_2nv5Y9tz5_0),.clk(gclk));
	jdff dff_B_NwWtRiby8_0(.din(w_dff_B_2nv5Y9tz5_0),.dout(w_dff_B_NwWtRiby8_0),.clk(gclk));
	jdff dff_B_8f9lUmVY2_0(.din(w_dff_B_NwWtRiby8_0),.dout(w_dff_B_8f9lUmVY2_0),.clk(gclk));
	jdff dff_B_MOJaemYw3_0(.din(w_dff_B_8f9lUmVY2_0),.dout(w_dff_B_MOJaemYw3_0),.clk(gclk));
	jdff dff_B_ubiPk2dv7_0(.din(w_dff_B_MOJaemYw3_0),.dout(w_dff_B_ubiPk2dv7_0),.clk(gclk));
	jdff dff_B_4Ah5fmIz1_0(.din(w_dff_B_ubiPk2dv7_0),.dout(w_dff_B_4Ah5fmIz1_0),.clk(gclk));
	jdff dff_B_eo5i8lER0_0(.din(w_dff_B_4Ah5fmIz1_0),.dout(w_dff_B_eo5i8lER0_0),.clk(gclk));
	jdff dff_B_fSBLeV4Y6_0(.din(w_dff_B_eo5i8lER0_0),.dout(w_dff_B_fSBLeV4Y6_0),.clk(gclk));
	jdff dff_B_8FG9T9k87_0(.din(w_dff_B_fSBLeV4Y6_0),.dout(w_dff_B_8FG9T9k87_0),.clk(gclk));
	jdff dff_B_RLiXS2969_0(.din(w_dff_B_8FG9T9k87_0),.dout(w_dff_B_RLiXS2969_0),.clk(gclk));
	jdff dff_B_MnNLDbuF8_0(.din(w_dff_B_RLiXS2969_0),.dout(w_dff_B_MnNLDbuF8_0),.clk(gclk));
	jdff dff_B_oKEFgqO73_0(.din(w_dff_B_MnNLDbuF8_0),.dout(w_dff_B_oKEFgqO73_0),.clk(gclk));
	jdff dff_B_cbwPiUJS3_0(.din(w_dff_B_oKEFgqO73_0),.dout(w_dff_B_cbwPiUJS3_0),.clk(gclk));
	jdff dff_B_1eid7WdF0_0(.din(w_dff_B_cbwPiUJS3_0),.dout(w_dff_B_1eid7WdF0_0),.clk(gclk));
	jdff dff_B_CytOpRm93_0(.din(w_dff_B_1eid7WdF0_0),.dout(w_dff_B_CytOpRm93_0),.clk(gclk));
	jdff dff_B_A5aCXa3M9_0(.din(w_dff_B_CytOpRm93_0),.dout(w_dff_B_A5aCXa3M9_0),.clk(gclk));
	jdff dff_B_Sr9ARhcy1_0(.din(w_dff_B_A5aCXa3M9_0),.dout(w_dff_B_Sr9ARhcy1_0),.clk(gclk));
	jdff dff_B_O2MXcG8D1_0(.din(w_dff_B_Sr9ARhcy1_0),.dout(w_dff_B_O2MXcG8D1_0),.clk(gclk));
	jdff dff_B_fw0AaPIr8_0(.din(w_dff_B_O2MXcG8D1_0),.dout(w_dff_B_fw0AaPIr8_0),.clk(gclk));
	jdff dff_B_8DxRkOeI1_0(.din(w_dff_B_fw0AaPIr8_0),.dout(w_dff_B_8DxRkOeI1_0),.clk(gclk));
	jdff dff_B_ChaCEjcx6_0(.din(w_dff_B_8DxRkOeI1_0),.dout(w_dff_B_ChaCEjcx6_0),.clk(gclk));
	jdff dff_B_LE7h1kVx6_0(.din(w_dff_B_ChaCEjcx6_0),.dout(w_dff_B_LE7h1kVx6_0),.clk(gclk));
	jdff dff_B_SR7lmSk17_0(.din(w_dff_B_LE7h1kVx6_0),.dout(w_dff_B_SR7lmSk17_0),.clk(gclk));
	jdff dff_B_upYOXlrG2_0(.din(w_dff_B_SR7lmSk17_0),.dout(w_dff_B_upYOXlrG2_0),.clk(gclk));
	jdff dff_B_ETyYKwbI8_0(.din(w_dff_B_upYOXlrG2_0),.dout(w_dff_B_ETyYKwbI8_0),.clk(gclk));
	jdff dff_B_A3JkxCNg8_0(.din(w_dff_B_ETyYKwbI8_0),.dout(w_dff_B_A3JkxCNg8_0),.clk(gclk));
	jdff dff_B_3sgCRIyf1_0(.din(w_dff_B_A3JkxCNg8_0),.dout(w_dff_B_3sgCRIyf1_0),.clk(gclk));
	jdff dff_B_SjXgULOd1_0(.din(w_dff_B_3sgCRIyf1_0),.dout(w_dff_B_SjXgULOd1_0),.clk(gclk));
	jdff dff_B_Mqk47ZQl3_0(.din(w_dff_B_SjXgULOd1_0),.dout(w_dff_B_Mqk47ZQl3_0),.clk(gclk));
	jdff dff_B_39aR6EaX5_0(.din(w_dff_B_Mqk47ZQl3_0),.dout(w_dff_B_39aR6EaX5_0),.clk(gclk));
	jdff dff_B_ZNXax4Ux1_0(.din(w_dff_B_39aR6EaX5_0),.dout(w_dff_B_ZNXax4Ux1_0),.clk(gclk));
	jdff dff_B_lL0rgrqc6_0(.din(w_dff_B_ZNXax4Ux1_0),.dout(w_dff_B_lL0rgrqc6_0),.clk(gclk));
	jdff dff_B_zWHxyE0u6_0(.din(w_dff_B_lL0rgrqc6_0),.dout(w_dff_B_zWHxyE0u6_0),.clk(gclk));
	jdff dff_B_azEX5QrN2_0(.din(w_dff_B_zWHxyE0u6_0),.dout(w_dff_B_azEX5QrN2_0),.clk(gclk));
	jdff dff_B_39Hqd9fk9_0(.din(w_dff_B_azEX5QrN2_0),.dout(w_dff_B_39Hqd9fk9_0),.clk(gclk));
	jdff dff_B_cYGe8lOB3_0(.din(w_dff_B_39Hqd9fk9_0),.dout(w_dff_B_cYGe8lOB3_0),.clk(gclk));
	jdff dff_B_XzuFU1fd3_0(.din(w_dff_B_cYGe8lOB3_0),.dout(w_dff_B_XzuFU1fd3_0),.clk(gclk));
	jdff dff_B_GVEkaWq78_0(.din(w_dff_B_XzuFU1fd3_0),.dout(w_dff_B_GVEkaWq78_0),.clk(gclk));
	jdff dff_B_SPYaZBIt9_0(.din(w_dff_B_GVEkaWq78_0),.dout(w_dff_B_SPYaZBIt9_0),.clk(gclk));
	jdff dff_B_IKK8GyuH4_0(.din(w_dff_B_SPYaZBIt9_0),.dout(w_dff_B_IKK8GyuH4_0),.clk(gclk));
	jdff dff_B_WPAHE3mh3_0(.din(w_dff_B_IKK8GyuH4_0),.dout(w_dff_B_WPAHE3mh3_0),.clk(gclk));
	jdff dff_B_nIdPCuCc6_0(.din(w_dff_B_WPAHE3mh3_0),.dout(w_dff_B_nIdPCuCc6_0),.clk(gclk));
	jdff dff_B_LyL1bnj37_0(.din(w_dff_B_nIdPCuCc6_0),.dout(w_dff_B_LyL1bnj37_0),.clk(gclk));
	jdff dff_B_r3MtVTUV4_0(.din(w_dff_B_LyL1bnj37_0),.dout(w_dff_B_r3MtVTUV4_0),.clk(gclk));
	jdff dff_B_49A45O3U7_0(.din(w_dff_B_r3MtVTUV4_0),.dout(w_dff_B_49A45O3U7_0),.clk(gclk));
	jdff dff_B_SPYIYyVM1_0(.din(w_dff_B_49A45O3U7_0),.dout(w_dff_B_SPYIYyVM1_0),.clk(gclk));
	jdff dff_B_3ITYnHvH3_0(.din(w_dff_B_SPYIYyVM1_0),.dout(w_dff_B_3ITYnHvH3_0),.clk(gclk));
	jdff dff_B_JIjQ7XFx8_0(.din(w_dff_B_3ITYnHvH3_0),.dout(w_dff_B_JIjQ7XFx8_0),.clk(gclk));
	jdff dff_B_xJ5r5Fbi2_0(.din(w_dff_B_JIjQ7XFx8_0),.dout(w_dff_B_xJ5r5Fbi2_0),.clk(gclk));
	jdff dff_B_uVjbqEq83_0(.din(w_dff_B_xJ5r5Fbi2_0),.dout(w_dff_B_uVjbqEq83_0),.clk(gclk));
	jdff dff_B_tDjI2Xgg9_0(.din(w_dff_B_uVjbqEq83_0),.dout(w_dff_B_tDjI2Xgg9_0),.clk(gclk));
	jdff dff_B_PDwlWK5J4_0(.din(w_dff_B_tDjI2Xgg9_0),.dout(w_dff_B_PDwlWK5J4_0),.clk(gclk));
	jdff dff_B_jxrQ0aod0_0(.din(w_dff_B_PDwlWK5J4_0),.dout(w_dff_B_jxrQ0aod0_0),.clk(gclk));
	jdff dff_B_zzWVvkcD6_0(.din(w_dff_B_jxrQ0aod0_0),.dout(w_dff_B_zzWVvkcD6_0),.clk(gclk));
	jdff dff_B_dh0e9h5F0_0(.din(w_dff_B_zzWVvkcD6_0),.dout(w_dff_B_dh0e9h5F0_0),.clk(gclk));
	jdff dff_B_wsbERzgk2_0(.din(w_dff_B_dh0e9h5F0_0),.dout(w_dff_B_wsbERzgk2_0),.clk(gclk));
	jdff dff_B_rKDKmjhn1_1(.din(n918),.dout(w_dff_B_rKDKmjhn1_1),.clk(gclk));
	jdff dff_B_er6DPLDV9_1(.din(w_dff_B_rKDKmjhn1_1),.dout(w_dff_B_er6DPLDV9_1),.clk(gclk));
	jdff dff_B_ODFTmzQx6_1(.din(w_dff_B_er6DPLDV9_1),.dout(w_dff_B_ODFTmzQx6_1),.clk(gclk));
	jdff dff_B_cdw8X4H16_1(.din(w_dff_B_ODFTmzQx6_1),.dout(w_dff_B_cdw8X4H16_1),.clk(gclk));
	jdff dff_B_mD0hgiOU4_1(.din(w_dff_B_cdw8X4H16_1),.dout(w_dff_B_mD0hgiOU4_1),.clk(gclk));
	jdff dff_B_XLPWQ5T59_1(.din(w_dff_B_mD0hgiOU4_1),.dout(w_dff_B_XLPWQ5T59_1),.clk(gclk));
	jdff dff_B_mHQpz9YE1_1(.din(w_dff_B_XLPWQ5T59_1),.dout(w_dff_B_mHQpz9YE1_1),.clk(gclk));
	jdff dff_B_KyEJI5Bt8_1(.din(w_dff_B_mHQpz9YE1_1),.dout(w_dff_B_KyEJI5Bt8_1),.clk(gclk));
	jdff dff_B_wq03rv2k6_1(.din(w_dff_B_KyEJI5Bt8_1),.dout(w_dff_B_wq03rv2k6_1),.clk(gclk));
	jdff dff_B_aiNAYzaR4_1(.din(w_dff_B_wq03rv2k6_1),.dout(w_dff_B_aiNAYzaR4_1),.clk(gclk));
	jdff dff_B_bx2HPkwq1_1(.din(w_dff_B_aiNAYzaR4_1),.dout(w_dff_B_bx2HPkwq1_1),.clk(gclk));
	jdff dff_B_6zDt640a2_1(.din(w_dff_B_bx2HPkwq1_1),.dout(w_dff_B_6zDt640a2_1),.clk(gclk));
	jdff dff_B_XxjHxdxX5_1(.din(w_dff_B_6zDt640a2_1),.dout(w_dff_B_XxjHxdxX5_1),.clk(gclk));
	jdff dff_B_XxhCUhdQ1_1(.din(w_dff_B_XxjHxdxX5_1),.dout(w_dff_B_XxhCUhdQ1_1),.clk(gclk));
	jdff dff_B_Zc7zOHuv6_1(.din(w_dff_B_XxhCUhdQ1_1),.dout(w_dff_B_Zc7zOHuv6_1),.clk(gclk));
	jdff dff_B_o8Akz7Mt5_1(.din(w_dff_B_Zc7zOHuv6_1),.dout(w_dff_B_o8Akz7Mt5_1),.clk(gclk));
	jdff dff_B_QEHvMTz34_1(.din(w_dff_B_o8Akz7Mt5_1),.dout(w_dff_B_QEHvMTz34_1),.clk(gclk));
	jdff dff_B_JsxK5gxm1_1(.din(w_dff_B_QEHvMTz34_1),.dout(w_dff_B_JsxK5gxm1_1),.clk(gclk));
	jdff dff_B_CQRFALly7_1(.din(w_dff_B_JsxK5gxm1_1),.dout(w_dff_B_CQRFALly7_1),.clk(gclk));
	jdff dff_B_Uf6KxqXy3_1(.din(w_dff_B_CQRFALly7_1),.dout(w_dff_B_Uf6KxqXy3_1),.clk(gclk));
	jdff dff_B_nl9xqzwR2_1(.din(w_dff_B_Uf6KxqXy3_1),.dout(w_dff_B_nl9xqzwR2_1),.clk(gclk));
	jdff dff_B_jPPhEZsJ2_1(.din(w_dff_B_nl9xqzwR2_1),.dout(w_dff_B_jPPhEZsJ2_1),.clk(gclk));
	jdff dff_B_FiU7s8qO1_1(.din(w_dff_B_jPPhEZsJ2_1),.dout(w_dff_B_FiU7s8qO1_1),.clk(gclk));
	jdff dff_B_kNypXD1Q4_1(.din(w_dff_B_FiU7s8qO1_1),.dout(w_dff_B_kNypXD1Q4_1),.clk(gclk));
	jdff dff_B_0RkdU8Dk8_1(.din(w_dff_B_kNypXD1Q4_1),.dout(w_dff_B_0RkdU8Dk8_1),.clk(gclk));
	jdff dff_B_EZSTBJhw7_1(.din(w_dff_B_0RkdU8Dk8_1),.dout(w_dff_B_EZSTBJhw7_1),.clk(gclk));
	jdff dff_B_tsV3vvCx4_1(.din(w_dff_B_EZSTBJhw7_1),.dout(w_dff_B_tsV3vvCx4_1),.clk(gclk));
	jdff dff_B_zL04EztH8_1(.din(w_dff_B_tsV3vvCx4_1),.dout(w_dff_B_zL04EztH8_1),.clk(gclk));
	jdff dff_B_bnYS9BIZ0_1(.din(w_dff_B_zL04EztH8_1),.dout(w_dff_B_bnYS9BIZ0_1),.clk(gclk));
	jdff dff_B_0HmWMjm60_1(.din(w_dff_B_bnYS9BIZ0_1),.dout(w_dff_B_0HmWMjm60_1),.clk(gclk));
	jdff dff_B_7cLCiQrE9_1(.din(w_dff_B_0HmWMjm60_1),.dout(w_dff_B_7cLCiQrE9_1),.clk(gclk));
	jdff dff_B_a43D8jlE0_1(.din(w_dff_B_7cLCiQrE9_1),.dout(w_dff_B_a43D8jlE0_1),.clk(gclk));
	jdff dff_B_ClCzBaz86_1(.din(w_dff_B_a43D8jlE0_1),.dout(w_dff_B_ClCzBaz86_1),.clk(gclk));
	jdff dff_B_H59AaPml8_1(.din(w_dff_B_ClCzBaz86_1),.dout(w_dff_B_H59AaPml8_1),.clk(gclk));
	jdff dff_B_zGXCVR4D2_1(.din(w_dff_B_H59AaPml8_1),.dout(w_dff_B_zGXCVR4D2_1),.clk(gclk));
	jdff dff_B_yowb84Xb8_1(.din(w_dff_B_zGXCVR4D2_1),.dout(w_dff_B_yowb84Xb8_1),.clk(gclk));
	jdff dff_B_bkDWcV3o3_1(.din(w_dff_B_yowb84Xb8_1),.dout(w_dff_B_bkDWcV3o3_1),.clk(gclk));
	jdff dff_B_VLrIIkL24_1(.din(w_dff_B_bkDWcV3o3_1),.dout(w_dff_B_VLrIIkL24_1),.clk(gclk));
	jdff dff_B_HuOV8PjD9_1(.din(w_dff_B_VLrIIkL24_1),.dout(w_dff_B_HuOV8PjD9_1),.clk(gclk));
	jdff dff_B_8dftSuwz0_1(.din(w_dff_B_HuOV8PjD9_1),.dout(w_dff_B_8dftSuwz0_1),.clk(gclk));
	jdff dff_B_SSKgH0KB3_1(.din(w_dff_B_8dftSuwz0_1),.dout(w_dff_B_SSKgH0KB3_1),.clk(gclk));
	jdff dff_B_JMRYtb9y7_1(.din(w_dff_B_SSKgH0KB3_1),.dout(w_dff_B_JMRYtb9y7_1),.clk(gclk));
	jdff dff_B_NEnxLnDV7_1(.din(w_dff_B_JMRYtb9y7_1),.dout(w_dff_B_NEnxLnDV7_1),.clk(gclk));
	jdff dff_B_amkxZG7q1_1(.din(w_dff_B_NEnxLnDV7_1),.dout(w_dff_B_amkxZG7q1_1),.clk(gclk));
	jdff dff_B_3HSDIFXS2_1(.din(w_dff_B_amkxZG7q1_1),.dout(w_dff_B_3HSDIFXS2_1),.clk(gclk));
	jdff dff_B_9wVIedni4_1(.din(w_dff_B_3HSDIFXS2_1),.dout(w_dff_B_9wVIedni4_1),.clk(gclk));
	jdff dff_B_ZSRuF6jb7_1(.din(w_dff_B_9wVIedni4_1),.dout(w_dff_B_ZSRuF6jb7_1),.clk(gclk));
	jdff dff_B_US6vRUHY0_1(.din(w_dff_B_ZSRuF6jb7_1),.dout(w_dff_B_US6vRUHY0_1),.clk(gclk));
	jdff dff_B_RzfUZ08N9_1(.din(w_dff_B_US6vRUHY0_1),.dout(w_dff_B_RzfUZ08N9_1),.clk(gclk));
	jdff dff_B_S7D9ZjUa7_1(.din(w_dff_B_RzfUZ08N9_1),.dout(w_dff_B_S7D9ZjUa7_1),.clk(gclk));
	jdff dff_B_V1bKtOVA2_1(.din(w_dff_B_S7D9ZjUa7_1),.dout(w_dff_B_V1bKtOVA2_1),.clk(gclk));
	jdff dff_B_ltlyL98u1_1(.din(w_dff_B_V1bKtOVA2_1),.dout(w_dff_B_ltlyL98u1_1),.clk(gclk));
	jdff dff_B_GiMVxJ3q9_1(.din(w_dff_B_ltlyL98u1_1),.dout(w_dff_B_GiMVxJ3q9_1),.clk(gclk));
	jdff dff_B_fKLzQruU2_1(.din(w_dff_B_GiMVxJ3q9_1),.dout(w_dff_B_fKLzQruU2_1),.clk(gclk));
	jdff dff_B_IMDbmNky4_1(.din(w_dff_B_fKLzQruU2_1),.dout(w_dff_B_IMDbmNky4_1),.clk(gclk));
	jdff dff_B_2YRG67FH6_1(.din(w_dff_B_IMDbmNky4_1),.dout(w_dff_B_2YRG67FH6_1),.clk(gclk));
	jdff dff_B_YM06LLsm5_1(.din(w_dff_B_2YRG67FH6_1),.dout(w_dff_B_YM06LLsm5_1),.clk(gclk));
	jdff dff_B_3e0Nst5O6_1(.din(w_dff_B_YM06LLsm5_1),.dout(w_dff_B_3e0Nst5O6_1),.clk(gclk));
	jdff dff_B_MBWRp3Ey3_1(.din(w_dff_B_3e0Nst5O6_1),.dout(w_dff_B_MBWRp3Ey3_1),.clk(gclk));
	jdff dff_B_PLdqrGPO2_1(.din(w_dff_B_MBWRp3Ey3_1),.dout(w_dff_B_PLdqrGPO2_1),.clk(gclk));
	jdff dff_B_BLqyRjBX1_1(.din(w_dff_B_PLdqrGPO2_1),.dout(w_dff_B_BLqyRjBX1_1),.clk(gclk));
	jdff dff_B_DKc8bUBK8_1(.din(w_dff_B_BLqyRjBX1_1),.dout(w_dff_B_DKc8bUBK8_1),.clk(gclk));
	jdff dff_B_GAlLQwWb0_1(.din(w_dff_B_DKc8bUBK8_1),.dout(w_dff_B_GAlLQwWb0_1),.clk(gclk));
	jdff dff_B_pwXVKTPS2_1(.din(w_dff_B_GAlLQwWb0_1),.dout(w_dff_B_pwXVKTPS2_1),.clk(gclk));
	jdff dff_B_2YBe1GuN5_1(.din(w_dff_B_pwXVKTPS2_1),.dout(w_dff_B_2YBe1GuN5_1),.clk(gclk));
	jdff dff_B_ieOnnjQB6_1(.din(w_dff_B_2YBe1GuN5_1),.dout(w_dff_B_ieOnnjQB6_1),.clk(gclk));
	jdff dff_B_ScSKBDkm6_1(.din(w_dff_B_ieOnnjQB6_1),.dout(w_dff_B_ScSKBDkm6_1),.clk(gclk));
	jdff dff_B_tr7FRnQa7_1(.din(w_dff_B_ScSKBDkm6_1),.dout(w_dff_B_tr7FRnQa7_1),.clk(gclk));
	jdff dff_B_bWrAbkGA7_1(.din(w_dff_B_tr7FRnQa7_1),.dout(w_dff_B_bWrAbkGA7_1),.clk(gclk));
	jdff dff_B_gohdcBDQ3_1(.din(w_dff_B_bWrAbkGA7_1),.dout(w_dff_B_gohdcBDQ3_1),.clk(gclk));
	jdff dff_B_Dql4hhBu7_1(.din(w_dff_B_gohdcBDQ3_1),.dout(w_dff_B_Dql4hhBu7_1),.clk(gclk));
	jdff dff_B_WVh3pUMT9_1(.din(w_dff_B_Dql4hhBu7_1),.dout(w_dff_B_WVh3pUMT9_1),.clk(gclk));
	jdff dff_B_WKXVA4Ld0_1(.din(w_dff_B_WVh3pUMT9_1),.dout(w_dff_B_WKXVA4Ld0_1),.clk(gclk));
	jdff dff_B_k2AYrc4j4_1(.din(w_dff_B_WKXVA4Ld0_1),.dout(w_dff_B_k2AYrc4j4_1),.clk(gclk));
	jdff dff_B_AdKJ3Hcc8_1(.din(w_dff_B_k2AYrc4j4_1),.dout(w_dff_B_AdKJ3Hcc8_1),.clk(gclk));
	jdff dff_B_jcSfwrUx9_1(.din(w_dff_B_AdKJ3Hcc8_1),.dout(w_dff_B_jcSfwrUx9_1),.clk(gclk));
	jdff dff_B_csSKlNFX4_1(.din(w_dff_B_jcSfwrUx9_1),.dout(w_dff_B_csSKlNFX4_1),.clk(gclk));
	jdff dff_B_ar2mZ5eW9_1(.din(w_dff_B_csSKlNFX4_1),.dout(w_dff_B_ar2mZ5eW9_1),.clk(gclk));
	jdff dff_B_6iVhIGeW4_1(.din(w_dff_B_ar2mZ5eW9_1),.dout(w_dff_B_6iVhIGeW4_1),.clk(gclk));
	jdff dff_B_404uCMXz1_1(.din(w_dff_B_6iVhIGeW4_1),.dout(w_dff_B_404uCMXz1_1),.clk(gclk));
	jdff dff_B_kYuYXyIp6_1(.din(w_dff_B_404uCMXz1_1),.dout(w_dff_B_kYuYXyIp6_1),.clk(gclk));
	jdff dff_B_k7t0G1JG8_1(.din(w_dff_B_kYuYXyIp6_1),.dout(w_dff_B_k7t0G1JG8_1),.clk(gclk));
	jdff dff_B_qxFNxcRM7_1(.din(w_dff_B_k7t0G1JG8_1),.dout(w_dff_B_qxFNxcRM7_1),.clk(gclk));
	jdff dff_B_FpTQl5Wl9_1(.din(w_dff_B_qxFNxcRM7_1),.dout(w_dff_B_FpTQl5Wl9_1),.clk(gclk));
	jdff dff_B_flJCG5ug4_1(.din(w_dff_B_FpTQl5Wl9_1),.dout(w_dff_B_flJCG5ug4_1),.clk(gclk));
	jdff dff_B_aOkUFpOL7_1(.din(w_dff_B_flJCG5ug4_1),.dout(w_dff_B_aOkUFpOL7_1),.clk(gclk));
	jdff dff_B_OLNO1eLj9_1(.din(w_dff_B_aOkUFpOL7_1),.dout(w_dff_B_OLNO1eLj9_1),.clk(gclk));
	jdff dff_B_AVhDbNiO2_1(.din(w_dff_B_OLNO1eLj9_1),.dout(w_dff_B_AVhDbNiO2_1),.clk(gclk));
	jdff dff_B_fXOzDmTA4_1(.din(w_dff_B_AVhDbNiO2_1),.dout(w_dff_B_fXOzDmTA4_1),.clk(gclk));
	jdff dff_B_CWY8rxXl1_0(.din(n919),.dout(w_dff_B_CWY8rxXl1_0),.clk(gclk));
	jdff dff_B_Ny70iVOY9_0(.din(w_dff_B_CWY8rxXl1_0),.dout(w_dff_B_Ny70iVOY9_0),.clk(gclk));
	jdff dff_B_Q9H4HAL91_0(.din(w_dff_B_Ny70iVOY9_0),.dout(w_dff_B_Q9H4HAL91_0),.clk(gclk));
	jdff dff_B_30UWpCw58_0(.din(w_dff_B_Q9H4HAL91_0),.dout(w_dff_B_30UWpCw58_0),.clk(gclk));
	jdff dff_B_omDmp2vB0_0(.din(w_dff_B_30UWpCw58_0),.dout(w_dff_B_omDmp2vB0_0),.clk(gclk));
	jdff dff_B_LGRf6koU9_0(.din(w_dff_B_omDmp2vB0_0),.dout(w_dff_B_LGRf6koU9_0),.clk(gclk));
	jdff dff_B_vwZCHmW48_0(.din(w_dff_B_LGRf6koU9_0),.dout(w_dff_B_vwZCHmW48_0),.clk(gclk));
	jdff dff_B_af6AY2XI5_0(.din(w_dff_B_vwZCHmW48_0),.dout(w_dff_B_af6AY2XI5_0),.clk(gclk));
	jdff dff_B_zDJTeMAT6_0(.din(w_dff_B_af6AY2XI5_0),.dout(w_dff_B_zDJTeMAT6_0),.clk(gclk));
	jdff dff_B_oifYlsDu9_0(.din(w_dff_B_zDJTeMAT6_0),.dout(w_dff_B_oifYlsDu9_0),.clk(gclk));
	jdff dff_B_zSKEdXgu0_0(.din(w_dff_B_oifYlsDu9_0),.dout(w_dff_B_zSKEdXgu0_0),.clk(gclk));
	jdff dff_B_FLTnRCvU1_0(.din(w_dff_B_zSKEdXgu0_0),.dout(w_dff_B_FLTnRCvU1_0),.clk(gclk));
	jdff dff_B_EWjKqhVF3_0(.din(w_dff_B_FLTnRCvU1_0),.dout(w_dff_B_EWjKqhVF3_0),.clk(gclk));
	jdff dff_B_uEblP9m40_0(.din(w_dff_B_EWjKqhVF3_0),.dout(w_dff_B_uEblP9m40_0),.clk(gclk));
	jdff dff_B_vLSkXsNv3_0(.din(w_dff_B_uEblP9m40_0),.dout(w_dff_B_vLSkXsNv3_0),.clk(gclk));
	jdff dff_B_0WWw44gL1_0(.din(w_dff_B_vLSkXsNv3_0),.dout(w_dff_B_0WWw44gL1_0),.clk(gclk));
	jdff dff_B_cT684YBL8_0(.din(w_dff_B_0WWw44gL1_0),.dout(w_dff_B_cT684YBL8_0),.clk(gclk));
	jdff dff_B_2iu8I3dq9_0(.din(w_dff_B_cT684YBL8_0),.dout(w_dff_B_2iu8I3dq9_0),.clk(gclk));
	jdff dff_B_n8Z6Ey0N6_0(.din(w_dff_B_2iu8I3dq9_0),.dout(w_dff_B_n8Z6Ey0N6_0),.clk(gclk));
	jdff dff_B_8kuPXEBp8_0(.din(w_dff_B_n8Z6Ey0N6_0),.dout(w_dff_B_8kuPXEBp8_0),.clk(gclk));
	jdff dff_B_n25xiboc3_0(.din(w_dff_B_8kuPXEBp8_0),.dout(w_dff_B_n25xiboc3_0),.clk(gclk));
	jdff dff_B_DM63jPwM4_0(.din(w_dff_B_n25xiboc3_0),.dout(w_dff_B_DM63jPwM4_0),.clk(gclk));
	jdff dff_B_q4Bj0sIl0_0(.din(w_dff_B_DM63jPwM4_0),.dout(w_dff_B_q4Bj0sIl0_0),.clk(gclk));
	jdff dff_B_I0hi6NFe2_0(.din(w_dff_B_q4Bj0sIl0_0),.dout(w_dff_B_I0hi6NFe2_0),.clk(gclk));
	jdff dff_B_EtL3VBlb5_0(.din(w_dff_B_I0hi6NFe2_0),.dout(w_dff_B_EtL3VBlb5_0),.clk(gclk));
	jdff dff_B_FSx0JAlp5_0(.din(w_dff_B_EtL3VBlb5_0),.dout(w_dff_B_FSx0JAlp5_0),.clk(gclk));
	jdff dff_B_x1PaXvSn0_0(.din(w_dff_B_FSx0JAlp5_0),.dout(w_dff_B_x1PaXvSn0_0),.clk(gclk));
	jdff dff_B_rMpptube3_0(.din(w_dff_B_x1PaXvSn0_0),.dout(w_dff_B_rMpptube3_0),.clk(gclk));
	jdff dff_B_4LXFm2cM8_0(.din(w_dff_B_rMpptube3_0),.dout(w_dff_B_4LXFm2cM8_0),.clk(gclk));
	jdff dff_B_MEdwn9WO6_0(.din(w_dff_B_4LXFm2cM8_0),.dout(w_dff_B_MEdwn9WO6_0),.clk(gclk));
	jdff dff_B_YZA7a6bx2_0(.din(w_dff_B_MEdwn9WO6_0),.dout(w_dff_B_YZA7a6bx2_0),.clk(gclk));
	jdff dff_B_pGg2c7GD7_0(.din(w_dff_B_YZA7a6bx2_0),.dout(w_dff_B_pGg2c7GD7_0),.clk(gclk));
	jdff dff_B_eCMr5V4a0_0(.din(w_dff_B_pGg2c7GD7_0),.dout(w_dff_B_eCMr5V4a0_0),.clk(gclk));
	jdff dff_B_3PDhePEA7_0(.din(w_dff_B_eCMr5V4a0_0),.dout(w_dff_B_3PDhePEA7_0),.clk(gclk));
	jdff dff_B_YjJH8gE13_0(.din(w_dff_B_3PDhePEA7_0),.dout(w_dff_B_YjJH8gE13_0),.clk(gclk));
	jdff dff_B_DtD70DHb6_0(.din(w_dff_B_YjJH8gE13_0),.dout(w_dff_B_DtD70DHb6_0),.clk(gclk));
	jdff dff_B_JPIFBaPW5_0(.din(w_dff_B_DtD70DHb6_0),.dout(w_dff_B_JPIFBaPW5_0),.clk(gclk));
	jdff dff_B_fC8vDLJp1_0(.din(w_dff_B_JPIFBaPW5_0),.dout(w_dff_B_fC8vDLJp1_0),.clk(gclk));
	jdff dff_B_R3uBh1WE3_0(.din(w_dff_B_fC8vDLJp1_0),.dout(w_dff_B_R3uBh1WE3_0),.clk(gclk));
	jdff dff_B_xX63uc1T8_0(.din(w_dff_B_R3uBh1WE3_0),.dout(w_dff_B_xX63uc1T8_0),.clk(gclk));
	jdff dff_B_IBGy8Mal3_0(.din(w_dff_B_xX63uc1T8_0),.dout(w_dff_B_IBGy8Mal3_0),.clk(gclk));
	jdff dff_B_CRlFtMDL1_0(.din(w_dff_B_IBGy8Mal3_0),.dout(w_dff_B_CRlFtMDL1_0),.clk(gclk));
	jdff dff_B_fhayUEiM1_0(.din(w_dff_B_CRlFtMDL1_0),.dout(w_dff_B_fhayUEiM1_0),.clk(gclk));
	jdff dff_B_CTT2RzvP6_0(.din(w_dff_B_fhayUEiM1_0),.dout(w_dff_B_CTT2RzvP6_0),.clk(gclk));
	jdff dff_B_GNpGWrch2_0(.din(w_dff_B_CTT2RzvP6_0),.dout(w_dff_B_GNpGWrch2_0),.clk(gclk));
	jdff dff_B_79o3CK3J5_0(.din(w_dff_B_GNpGWrch2_0),.dout(w_dff_B_79o3CK3J5_0),.clk(gclk));
	jdff dff_B_wJccEvqV2_0(.din(w_dff_B_79o3CK3J5_0),.dout(w_dff_B_wJccEvqV2_0),.clk(gclk));
	jdff dff_B_qZc6Kva81_0(.din(w_dff_B_wJccEvqV2_0),.dout(w_dff_B_qZc6Kva81_0),.clk(gclk));
	jdff dff_B_58n5S6Og6_0(.din(w_dff_B_qZc6Kva81_0),.dout(w_dff_B_58n5S6Og6_0),.clk(gclk));
	jdff dff_B_gbbwywZx9_0(.din(w_dff_B_58n5S6Og6_0),.dout(w_dff_B_gbbwywZx9_0),.clk(gclk));
	jdff dff_B_DBQAm4B07_0(.din(w_dff_B_gbbwywZx9_0),.dout(w_dff_B_DBQAm4B07_0),.clk(gclk));
	jdff dff_B_M1BI0gGk2_0(.din(w_dff_B_DBQAm4B07_0),.dout(w_dff_B_M1BI0gGk2_0),.clk(gclk));
	jdff dff_B_2qmu4oG88_0(.din(w_dff_B_M1BI0gGk2_0),.dout(w_dff_B_2qmu4oG88_0),.clk(gclk));
	jdff dff_B_FT5BDjny3_0(.din(w_dff_B_2qmu4oG88_0),.dout(w_dff_B_FT5BDjny3_0),.clk(gclk));
	jdff dff_B_Q9hu3h5h6_0(.din(w_dff_B_FT5BDjny3_0),.dout(w_dff_B_Q9hu3h5h6_0),.clk(gclk));
	jdff dff_B_MVyVtx7U7_0(.din(w_dff_B_Q9hu3h5h6_0),.dout(w_dff_B_MVyVtx7U7_0),.clk(gclk));
	jdff dff_B_ksW94IBm2_0(.din(w_dff_B_MVyVtx7U7_0),.dout(w_dff_B_ksW94IBm2_0),.clk(gclk));
	jdff dff_B_edURTfez4_0(.din(w_dff_B_ksW94IBm2_0),.dout(w_dff_B_edURTfez4_0),.clk(gclk));
	jdff dff_B_moy20kW28_0(.din(w_dff_B_edURTfez4_0),.dout(w_dff_B_moy20kW28_0),.clk(gclk));
	jdff dff_B_AES7Vx9z9_0(.din(w_dff_B_moy20kW28_0),.dout(w_dff_B_AES7Vx9z9_0),.clk(gclk));
	jdff dff_B_wTLA7ySI6_0(.din(w_dff_B_AES7Vx9z9_0),.dout(w_dff_B_wTLA7ySI6_0),.clk(gclk));
	jdff dff_B_KKmk6h587_0(.din(w_dff_B_wTLA7ySI6_0),.dout(w_dff_B_KKmk6h587_0),.clk(gclk));
	jdff dff_B_mUBHhjhV0_0(.din(w_dff_B_KKmk6h587_0),.dout(w_dff_B_mUBHhjhV0_0),.clk(gclk));
	jdff dff_B_6t2YTT5n9_0(.din(w_dff_B_mUBHhjhV0_0),.dout(w_dff_B_6t2YTT5n9_0),.clk(gclk));
	jdff dff_B_iyju2Npd6_0(.din(w_dff_B_6t2YTT5n9_0),.dout(w_dff_B_iyju2Npd6_0),.clk(gclk));
	jdff dff_B_MbGZNfAM5_0(.din(w_dff_B_iyju2Npd6_0),.dout(w_dff_B_MbGZNfAM5_0),.clk(gclk));
	jdff dff_B_n0UEG5tt1_0(.din(w_dff_B_MbGZNfAM5_0),.dout(w_dff_B_n0UEG5tt1_0),.clk(gclk));
	jdff dff_B_gf76WM7O6_0(.din(w_dff_B_n0UEG5tt1_0),.dout(w_dff_B_gf76WM7O6_0),.clk(gclk));
	jdff dff_B_BUsnqW3l9_0(.din(w_dff_B_gf76WM7O6_0),.dout(w_dff_B_BUsnqW3l9_0),.clk(gclk));
	jdff dff_B_O49HHtdK9_0(.din(w_dff_B_BUsnqW3l9_0),.dout(w_dff_B_O49HHtdK9_0),.clk(gclk));
	jdff dff_B_U0LAbCxi3_0(.din(w_dff_B_O49HHtdK9_0),.dout(w_dff_B_U0LAbCxi3_0),.clk(gclk));
	jdff dff_B_tmd08aPY9_0(.din(w_dff_B_U0LAbCxi3_0),.dout(w_dff_B_tmd08aPY9_0),.clk(gclk));
	jdff dff_B_gLwQOAJk1_0(.din(w_dff_B_tmd08aPY9_0),.dout(w_dff_B_gLwQOAJk1_0),.clk(gclk));
	jdff dff_B_ouLHRigy8_0(.din(w_dff_B_gLwQOAJk1_0),.dout(w_dff_B_ouLHRigy8_0),.clk(gclk));
	jdff dff_B_tPkjOYBy4_0(.din(w_dff_B_ouLHRigy8_0),.dout(w_dff_B_tPkjOYBy4_0),.clk(gclk));
	jdff dff_B_vILfiHHU9_0(.din(w_dff_B_tPkjOYBy4_0),.dout(w_dff_B_vILfiHHU9_0),.clk(gclk));
	jdff dff_B_R2PnrNGY4_0(.din(w_dff_B_vILfiHHU9_0),.dout(w_dff_B_R2PnrNGY4_0),.clk(gclk));
	jdff dff_B_FqO1L7OJ6_0(.din(w_dff_B_R2PnrNGY4_0),.dout(w_dff_B_FqO1L7OJ6_0),.clk(gclk));
	jdff dff_B_wyKOe8zS5_0(.din(w_dff_B_FqO1L7OJ6_0),.dout(w_dff_B_wyKOe8zS5_0),.clk(gclk));
	jdff dff_B_ufcbxOSq4_0(.din(w_dff_B_wyKOe8zS5_0),.dout(w_dff_B_ufcbxOSq4_0),.clk(gclk));
	jdff dff_B_D7GKjPWf6_0(.din(w_dff_B_ufcbxOSq4_0),.dout(w_dff_B_D7GKjPWf6_0),.clk(gclk));
	jdff dff_B_sD6exW0m0_0(.din(w_dff_B_D7GKjPWf6_0),.dout(w_dff_B_sD6exW0m0_0),.clk(gclk));
	jdff dff_B_MoMNsD464_0(.din(w_dff_B_sD6exW0m0_0),.dout(w_dff_B_MoMNsD464_0),.clk(gclk));
	jdff dff_B_a01Bcux69_0(.din(w_dff_B_MoMNsD464_0),.dout(w_dff_B_a01Bcux69_0),.clk(gclk));
	jdff dff_B_HWHgsry20_0(.din(w_dff_B_a01Bcux69_0),.dout(w_dff_B_HWHgsry20_0),.clk(gclk));
	jdff dff_B_QsNjBccf5_0(.din(w_dff_B_HWHgsry20_0),.dout(w_dff_B_QsNjBccf5_0),.clk(gclk));
	jdff dff_B_TgKETz5Q9_0(.din(w_dff_B_QsNjBccf5_0),.dout(w_dff_B_TgKETz5Q9_0),.clk(gclk));
	jdff dff_B_JZOXfO6O4_0(.din(w_dff_B_TgKETz5Q9_0),.dout(w_dff_B_JZOXfO6O4_0),.clk(gclk));
	jdff dff_B_AOA64WTK7_0(.din(w_dff_B_JZOXfO6O4_0),.dout(w_dff_B_AOA64WTK7_0),.clk(gclk));
	jdff dff_B_UPtvfWU60_1(.din(n912),.dout(w_dff_B_UPtvfWU60_1),.clk(gclk));
	jdff dff_B_UuOGWOQp9_1(.din(w_dff_B_UPtvfWU60_1),.dout(w_dff_B_UuOGWOQp9_1),.clk(gclk));
	jdff dff_B_yMt3zrPz8_1(.din(w_dff_B_UuOGWOQp9_1),.dout(w_dff_B_yMt3zrPz8_1),.clk(gclk));
	jdff dff_B_8P3Gnk313_1(.din(w_dff_B_yMt3zrPz8_1),.dout(w_dff_B_8P3Gnk313_1),.clk(gclk));
	jdff dff_B_LYUouN115_1(.din(w_dff_B_8P3Gnk313_1),.dout(w_dff_B_LYUouN115_1),.clk(gclk));
	jdff dff_B_h0DfzFCB3_1(.din(w_dff_B_LYUouN115_1),.dout(w_dff_B_h0DfzFCB3_1),.clk(gclk));
	jdff dff_B_knu0rVNO2_1(.din(w_dff_B_h0DfzFCB3_1),.dout(w_dff_B_knu0rVNO2_1),.clk(gclk));
	jdff dff_B_CZDWk2PV0_1(.din(w_dff_B_knu0rVNO2_1),.dout(w_dff_B_CZDWk2PV0_1),.clk(gclk));
	jdff dff_B_EA5nR9F51_1(.din(w_dff_B_CZDWk2PV0_1),.dout(w_dff_B_EA5nR9F51_1),.clk(gclk));
	jdff dff_B_duyFeznp0_1(.din(w_dff_B_EA5nR9F51_1),.dout(w_dff_B_duyFeznp0_1),.clk(gclk));
	jdff dff_B_TcBiiXrJ3_1(.din(w_dff_B_duyFeznp0_1),.dout(w_dff_B_TcBiiXrJ3_1),.clk(gclk));
	jdff dff_B_uLSGMLcW8_1(.din(w_dff_B_TcBiiXrJ3_1),.dout(w_dff_B_uLSGMLcW8_1),.clk(gclk));
	jdff dff_B_v0TSw7JI3_1(.din(w_dff_B_uLSGMLcW8_1),.dout(w_dff_B_v0TSw7JI3_1),.clk(gclk));
	jdff dff_B_4t17URdi6_1(.din(w_dff_B_v0TSw7JI3_1),.dout(w_dff_B_4t17URdi6_1),.clk(gclk));
	jdff dff_B_vE3UuXuF7_1(.din(w_dff_B_4t17URdi6_1),.dout(w_dff_B_vE3UuXuF7_1),.clk(gclk));
	jdff dff_B_R5k7A6RI9_1(.din(w_dff_B_vE3UuXuF7_1),.dout(w_dff_B_R5k7A6RI9_1),.clk(gclk));
	jdff dff_B_WlfhKH3U5_1(.din(w_dff_B_R5k7A6RI9_1),.dout(w_dff_B_WlfhKH3U5_1),.clk(gclk));
	jdff dff_B_cI3IDdS14_1(.din(w_dff_B_WlfhKH3U5_1),.dout(w_dff_B_cI3IDdS14_1),.clk(gclk));
	jdff dff_B_aeAVzOg09_1(.din(w_dff_B_cI3IDdS14_1),.dout(w_dff_B_aeAVzOg09_1),.clk(gclk));
	jdff dff_B_cFj5Rkyd6_1(.din(w_dff_B_aeAVzOg09_1),.dout(w_dff_B_cFj5Rkyd6_1),.clk(gclk));
	jdff dff_B_qTb8J63n7_1(.din(w_dff_B_cFj5Rkyd6_1),.dout(w_dff_B_qTb8J63n7_1),.clk(gclk));
	jdff dff_B_uOx7elwQ2_1(.din(w_dff_B_qTb8J63n7_1),.dout(w_dff_B_uOx7elwQ2_1),.clk(gclk));
	jdff dff_B_JSZ2VZWM4_1(.din(w_dff_B_uOx7elwQ2_1),.dout(w_dff_B_JSZ2VZWM4_1),.clk(gclk));
	jdff dff_B_F7FYp8q85_1(.din(w_dff_B_JSZ2VZWM4_1),.dout(w_dff_B_F7FYp8q85_1),.clk(gclk));
	jdff dff_B_V1ZQmTS75_1(.din(w_dff_B_F7FYp8q85_1),.dout(w_dff_B_V1ZQmTS75_1),.clk(gclk));
	jdff dff_B_g8Zm9LJX0_1(.din(w_dff_B_V1ZQmTS75_1),.dout(w_dff_B_g8Zm9LJX0_1),.clk(gclk));
	jdff dff_B_iufyHvuQ4_1(.din(w_dff_B_g8Zm9LJX0_1),.dout(w_dff_B_iufyHvuQ4_1),.clk(gclk));
	jdff dff_B_Wa2XdwjX7_1(.din(w_dff_B_iufyHvuQ4_1),.dout(w_dff_B_Wa2XdwjX7_1),.clk(gclk));
	jdff dff_B_K6xUvzdL9_1(.din(w_dff_B_Wa2XdwjX7_1),.dout(w_dff_B_K6xUvzdL9_1),.clk(gclk));
	jdff dff_B_OgvBeiFM7_1(.din(w_dff_B_K6xUvzdL9_1),.dout(w_dff_B_OgvBeiFM7_1),.clk(gclk));
	jdff dff_B_sLV6BVkR5_1(.din(w_dff_B_OgvBeiFM7_1),.dout(w_dff_B_sLV6BVkR5_1),.clk(gclk));
	jdff dff_B_Ej2EvRIy2_1(.din(w_dff_B_sLV6BVkR5_1),.dout(w_dff_B_Ej2EvRIy2_1),.clk(gclk));
	jdff dff_B_HGsJMk7P0_1(.din(w_dff_B_Ej2EvRIy2_1),.dout(w_dff_B_HGsJMk7P0_1),.clk(gclk));
	jdff dff_B_gjfCaYEd9_1(.din(w_dff_B_HGsJMk7P0_1),.dout(w_dff_B_gjfCaYEd9_1),.clk(gclk));
	jdff dff_B_urQqdP6W4_1(.din(w_dff_B_gjfCaYEd9_1),.dout(w_dff_B_urQqdP6W4_1),.clk(gclk));
	jdff dff_B_rd9rnUmv2_1(.din(w_dff_B_urQqdP6W4_1),.dout(w_dff_B_rd9rnUmv2_1),.clk(gclk));
	jdff dff_B_7zEgOf3D5_1(.din(w_dff_B_rd9rnUmv2_1),.dout(w_dff_B_7zEgOf3D5_1),.clk(gclk));
	jdff dff_B_R4kYRWuP0_1(.din(w_dff_B_7zEgOf3D5_1),.dout(w_dff_B_R4kYRWuP0_1),.clk(gclk));
	jdff dff_B_7yUVFmDn0_1(.din(w_dff_B_R4kYRWuP0_1),.dout(w_dff_B_7yUVFmDn0_1),.clk(gclk));
	jdff dff_B_WUXOmaGF5_1(.din(w_dff_B_7yUVFmDn0_1),.dout(w_dff_B_WUXOmaGF5_1),.clk(gclk));
	jdff dff_B_AyXoPT2q4_1(.din(w_dff_B_WUXOmaGF5_1),.dout(w_dff_B_AyXoPT2q4_1),.clk(gclk));
	jdff dff_B_yoITZG6x9_1(.din(w_dff_B_AyXoPT2q4_1),.dout(w_dff_B_yoITZG6x9_1),.clk(gclk));
	jdff dff_B_j8H2qCDz2_1(.din(w_dff_B_yoITZG6x9_1),.dout(w_dff_B_j8H2qCDz2_1),.clk(gclk));
	jdff dff_B_cxJ5m42a9_1(.din(w_dff_B_j8H2qCDz2_1),.dout(w_dff_B_cxJ5m42a9_1),.clk(gclk));
	jdff dff_B_3kJ06I5f3_1(.din(w_dff_B_cxJ5m42a9_1),.dout(w_dff_B_3kJ06I5f3_1),.clk(gclk));
	jdff dff_B_7G3xDoNL0_1(.din(w_dff_B_3kJ06I5f3_1),.dout(w_dff_B_7G3xDoNL0_1),.clk(gclk));
	jdff dff_B_kdItoFeT0_1(.din(w_dff_B_7G3xDoNL0_1),.dout(w_dff_B_kdItoFeT0_1),.clk(gclk));
	jdff dff_B_qPjCYXlb9_1(.din(w_dff_B_kdItoFeT0_1),.dout(w_dff_B_qPjCYXlb9_1),.clk(gclk));
	jdff dff_B_KjKFHHGJ3_1(.din(w_dff_B_qPjCYXlb9_1),.dout(w_dff_B_KjKFHHGJ3_1),.clk(gclk));
	jdff dff_B_4H8rZfp22_1(.din(w_dff_B_KjKFHHGJ3_1),.dout(w_dff_B_4H8rZfp22_1),.clk(gclk));
	jdff dff_B_I6ZHTxQ72_1(.din(w_dff_B_4H8rZfp22_1),.dout(w_dff_B_I6ZHTxQ72_1),.clk(gclk));
	jdff dff_B_mAIZ0iRx5_1(.din(w_dff_B_I6ZHTxQ72_1),.dout(w_dff_B_mAIZ0iRx5_1),.clk(gclk));
	jdff dff_B_N671BKDk2_1(.din(w_dff_B_mAIZ0iRx5_1),.dout(w_dff_B_N671BKDk2_1),.clk(gclk));
	jdff dff_B_zoxs8NpC1_1(.din(w_dff_B_N671BKDk2_1),.dout(w_dff_B_zoxs8NpC1_1),.clk(gclk));
	jdff dff_B_Q8WXGUNJ9_1(.din(w_dff_B_zoxs8NpC1_1),.dout(w_dff_B_Q8WXGUNJ9_1),.clk(gclk));
	jdff dff_B_Eq45sx0L3_1(.din(w_dff_B_Q8WXGUNJ9_1),.dout(w_dff_B_Eq45sx0L3_1),.clk(gclk));
	jdff dff_B_pYASwdi28_1(.din(w_dff_B_Eq45sx0L3_1),.dout(w_dff_B_pYASwdi28_1),.clk(gclk));
	jdff dff_B_tMOh0O4u2_1(.din(w_dff_B_pYASwdi28_1),.dout(w_dff_B_tMOh0O4u2_1),.clk(gclk));
	jdff dff_B_0roOkXH24_1(.din(w_dff_B_tMOh0O4u2_1),.dout(w_dff_B_0roOkXH24_1),.clk(gclk));
	jdff dff_B_MH69ShYO8_1(.din(w_dff_B_0roOkXH24_1),.dout(w_dff_B_MH69ShYO8_1),.clk(gclk));
	jdff dff_B_vSiNR5eF4_1(.din(w_dff_B_MH69ShYO8_1),.dout(w_dff_B_vSiNR5eF4_1),.clk(gclk));
	jdff dff_B_YPeD6d7k1_1(.din(w_dff_B_vSiNR5eF4_1),.dout(w_dff_B_YPeD6d7k1_1),.clk(gclk));
	jdff dff_B_fHsyco9E6_1(.din(w_dff_B_YPeD6d7k1_1),.dout(w_dff_B_fHsyco9E6_1),.clk(gclk));
	jdff dff_B_CnWOAJ7q1_1(.din(w_dff_B_fHsyco9E6_1),.dout(w_dff_B_CnWOAJ7q1_1),.clk(gclk));
	jdff dff_B_Mxv6c0mD9_1(.din(w_dff_B_CnWOAJ7q1_1),.dout(w_dff_B_Mxv6c0mD9_1),.clk(gclk));
	jdff dff_B_yAllGcT59_1(.din(w_dff_B_Mxv6c0mD9_1),.dout(w_dff_B_yAllGcT59_1),.clk(gclk));
	jdff dff_B_qWiGnwCm2_1(.din(w_dff_B_yAllGcT59_1),.dout(w_dff_B_qWiGnwCm2_1),.clk(gclk));
	jdff dff_B_iZqOtCPt9_1(.din(w_dff_B_qWiGnwCm2_1),.dout(w_dff_B_iZqOtCPt9_1),.clk(gclk));
	jdff dff_B_BBhfh24u9_1(.din(w_dff_B_iZqOtCPt9_1),.dout(w_dff_B_BBhfh24u9_1),.clk(gclk));
	jdff dff_B_rI29TUNV0_1(.din(w_dff_B_BBhfh24u9_1),.dout(w_dff_B_rI29TUNV0_1),.clk(gclk));
	jdff dff_B_4zmlxP5B9_1(.din(w_dff_B_rI29TUNV0_1),.dout(w_dff_B_4zmlxP5B9_1),.clk(gclk));
	jdff dff_B_9BlZBOlK0_1(.din(w_dff_B_4zmlxP5B9_1),.dout(w_dff_B_9BlZBOlK0_1),.clk(gclk));
	jdff dff_B_dGbXgqSD7_1(.din(w_dff_B_9BlZBOlK0_1),.dout(w_dff_B_dGbXgqSD7_1),.clk(gclk));
	jdff dff_B_vfag6Alh2_1(.din(w_dff_B_dGbXgqSD7_1),.dout(w_dff_B_vfag6Alh2_1),.clk(gclk));
	jdff dff_B_viRKEOL81_1(.din(w_dff_B_vfag6Alh2_1),.dout(w_dff_B_viRKEOL81_1),.clk(gclk));
	jdff dff_B_GwWNSl3K4_1(.din(w_dff_B_viRKEOL81_1),.dout(w_dff_B_GwWNSl3K4_1),.clk(gclk));
	jdff dff_B_mmGaHJCF4_1(.din(w_dff_B_GwWNSl3K4_1),.dout(w_dff_B_mmGaHJCF4_1),.clk(gclk));
	jdff dff_B_EuDKPksJ8_1(.din(w_dff_B_mmGaHJCF4_1),.dout(w_dff_B_EuDKPksJ8_1),.clk(gclk));
	jdff dff_B_vJdIGQTd9_1(.din(w_dff_B_EuDKPksJ8_1),.dout(w_dff_B_vJdIGQTd9_1),.clk(gclk));
	jdff dff_B_6Q20xzzj1_1(.din(w_dff_B_vJdIGQTd9_1),.dout(w_dff_B_6Q20xzzj1_1),.clk(gclk));
	jdff dff_B_z6lZE8jM0_1(.din(w_dff_B_6Q20xzzj1_1),.dout(w_dff_B_z6lZE8jM0_1),.clk(gclk));
	jdff dff_B_JzzNGpKQ4_1(.din(w_dff_B_z6lZE8jM0_1),.dout(w_dff_B_JzzNGpKQ4_1),.clk(gclk));
	jdff dff_B_EoiDjHmx8_1(.din(w_dff_B_JzzNGpKQ4_1),.dout(w_dff_B_EoiDjHmx8_1),.clk(gclk));
	jdff dff_B_aYMo1f8Q1_1(.din(w_dff_B_EoiDjHmx8_1),.dout(w_dff_B_aYMo1f8Q1_1),.clk(gclk));
	jdff dff_B_9wosPKm44_1(.din(w_dff_B_aYMo1f8Q1_1),.dout(w_dff_B_9wosPKm44_1),.clk(gclk));
	jdff dff_B_cAUCsaW39_1(.din(w_dff_B_9wosPKm44_1),.dout(w_dff_B_cAUCsaW39_1),.clk(gclk));
	jdff dff_B_TPpqxXKK1_1(.din(w_dff_B_cAUCsaW39_1),.dout(w_dff_B_TPpqxXKK1_1),.clk(gclk));
	jdff dff_B_brSNaHyt4_1(.din(w_dff_B_TPpqxXKK1_1),.dout(w_dff_B_brSNaHyt4_1),.clk(gclk));
	jdff dff_B_gj9BSaQ32_0(.din(n913),.dout(w_dff_B_gj9BSaQ32_0),.clk(gclk));
	jdff dff_B_zScffpru6_0(.din(w_dff_B_gj9BSaQ32_0),.dout(w_dff_B_zScffpru6_0),.clk(gclk));
	jdff dff_B_eRTzEZpJ6_0(.din(w_dff_B_zScffpru6_0),.dout(w_dff_B_eRTzEZpJ6_0),.clk(gclk));
	jdff dff_B_01rWgdmJ3_0(.din(w_dff_B_eRTzEZpJ6_0),.dout(w_dff_B_01rWgdmJ3_0),.clk(gclk));
	jdff dff_B_QuU0yevI8_0(.din(w_dff_B_01rWgdmJ3_0),.dout(w_dff_B_QuU0yevI8_0),.clk(gclk));
	jdff dff_B_WuP55TXA7_0(.din(w_dff_B_QuU0yevI8_0),.dout(w_dff_B_WuP55TXA7_0),.clk(gclk));
	jdff dff_B_zn9j9xCW5_0(.din(w_dff_B_WuP55TXA7_0),.dout(w_dff_B_zn9j9xCW5_0),.clk(gclk));
	jdff dff_B_wqVOPVUm3_0(.din(w_dff_B_zn9j9xCW5_0),.dout(w_dff_B_wqVOPVUm3_0),.clk(gclk));
	jdff dff_B_dN4gfwnQ8_0(.din(w_dff_B_wqVOPVUm3_0),.dout(w_dff_B_dN4gfwnQ8_0),.clk(gclk));
	jdff dff_B_RenkfMsc9_0(.din(w_dff_B_dN4gfwnQ8_0),.dout(w_dff_B_RenkfMsc9_0),.clk(gclk));
	jdff dff_B_cqGmaX3E7_0(.din(w_dff_B_RenkfMsc9_0),.dout(w_dff_B_cqGmaX3E7_0),.clk(gclk));
	jdff dff_B_PtwmYSdd5_0(.din(w_dff_B_cqGmaX3E7_0),.dout(w_dff_B_PtwmYSdd5_0),.clk(gclk));
	jdff dff_B_WuZw9MOB7_0(.din(w_dff_B_PtwmYSdd5_0),.dout(w_dff_B_WuZw9MOB7_0),.clk(gclk));
	jdff dff_B_IXVE1zvs5_0(.din(w_dff_B_WuZw9MOB7_0),.dout(w_dff_B_IXVE1zvs5_0),.clk(gclk));
	jdff dff_B_fimdODgY4_0(.din(w_dff_B_IXVE1zvs5_0),.dout(w_dff_B_fimdODgY4_0),.clk(gclk));
	jdff dff_B_O4nudeKV7_0(.din(w_dff_B_fimdODgY4_0),.dout(w_dff_B_O4nudeKV7_0),.clk(gclk));
	jdff dff_B_HjBxPVmu6_0(.din(w_dff_B_O4nudeKV7_0),.dout(w_dff_B_HjBxPVmu6_0),.clk(gclk));
	jdff dff_B_QNx5d1kF9_0(.din(w_dff_B_HjBxPVmu6_0),.dout(w_dff_B_QNx5d1kF9_0),.clk(gclk));
	jdff dff_B_u8AICUb41_0(.din(w_dff_B_QNx5d1kF9_0),.dout(w_dff_B_u8AICUb41_0),.clk(gclk));
	jdff dff_B_Nw9h7WSn4_0(.din(w_dff_B_u8AICUb41_0),.dout(w_dff_B_Nw9h7WSn4_0),.clk(gclk));
	jdff dff_B_WFLAkxCm6_0(.din(w_dff_B_Nw9h7WSn4_0),.dout(w_dff_B_WFLAkxCm6_0),.clk(gclk));
	jdff dff_B_dIO8Od0q6_0(.din(w_dff_B_WFLAkxCm6_0),.dout(w_dff_B_dIO8Od0q6_0),.clk(gclk));
	jdff dff_B_OnURPUhk5_0(.din(w_dff_B_dIO8Od0q6_0),.dout(w_dff_B_OnURPUhk5_0),.clk(gclk));
	jdff dff_B_1fbtBmKS0_0(.din(w_dff_B_OnURPUhk5_0),.dout(w_dff_B_1fbtBmKS0_0),.clk(gclk));
	jdff dff_B_wX4S2dqZ2_0(.din(w_dff_B_1fbtBmKS0_0),.dout(w_dff_B_wX4S2dqZ2_0),.clk(gclk));
	jdff dff_B_weSLLnbF3_0(.din(w_dff_B_wX4S2dqZ2_0),.dout(w_dff_B_weSLLnbF3_0),.clk(gclk));
	jdff dff_B_hEbhc98o2_0(.din(w_dff_B_weSLLnbF3_0),.dout(w_dff_B_hEbhc98o2_0),.clk(gclk));
	jdff dff_B_O5FKdVO75_0(.din(w_dff_B_hEbhc98o2_0),.dout(w_dff_B_O5FKdVO75_0),.clk(gclk));
	jdff dff_B_lwZGOtEz8_0(.din(w_dff_B_O5FKdVO75_0),.dout(w_dff_B_lwZGOtEz8_0),.clk(gclk));
	jdff dff_B_j8v2niyu4_0(.din(w_dff_B_lwZGOtEz8_0),.dout(w_dff_B_j8v2niyu4_0),.clk(gclk));
	jdff dff_B_Cgw5QtpC0_0(.din(w_dff_B_j8v2niyu4_0),.dout(w_dff_B_Cgw5QtpC0_0),.clk(gclk));
	jdff dff_B_2b8Jtanv8_0(.din(w_dff_B_Cgw5QtpC0_0),.dout(w_dff_B_2b8Jtanv8_0),.clk(gclk));
	jdff dff_B_kBRfDvoP4_0(.din(w_dff_B_2b8Jtanv8_0),.dout(w_dff_B_kBRfDvoP4_0),.clk(gclk));
	jdff dff_B_Nw7jXWAZ9_0(.din(w_dff_B_kBRfDvoP4_0),.dout(w_dff_B_Nw7jXWAZ9_0),.clk(gclk));
	jdff dff_B_Mf0LqrWX5_0(.din(w_dff_B_Nw7jXWAZ9_0),.dout(w_dff_B_Mf0LqrWX5_0),.clk(gclk));
	jdff dff_B_qyZixoqC9_0(.din(w_dff_B_Mf0LqrWX5_0),.dout(w_dff_B_qyZixoqC9_0),.clk(gclk));
	jdff dff_B_aiZLZEq63_0(.din(w_dff_B_qyZixoqC9_0),.dout(w_dff_B_aiZLZEq63_0),.clk(gclk));
	jdff dff_B_1AaDvqDm1_0(.din(w_dff_B_aiZLZEq63_0),.dout(w_dff_B_1AaDvqDm1_0),.clk(gclk));
	jdff dff_B_gH7gHrNK6_0(.din(w_dff_B_1AaDvqDm1_0),.dout(w_dff_B_gH7gHrNK6_0),.clk(gclk));
	jdff dff_B_EIVlY7Gq6_0(.din(w_dff_B_gH7gHrNK6_0),.dout(w_dff_B_EIVlY7Gq6_0),.clk(gclk));
	jdff dff_B_hAg9ZTMY9_0(.din(w_dff_B_EIVlY7Gq6_0),.dout(w_dff_B_hAg9ZTMY9_0),.clk(gclk));
	jdff dff_B_fiBGJqbq1_0(.din(w_dff_B_hAg9ZTMY9_0),.dout(w_dff_B_fiBGJqbq1_0),.clk(gclk));
	jdff dff_B_ZGRaC1kQ2_0(.din(w_dff_B_fiBGJqbq1_0),.dout(w_dff_B_ZGRaC1kQ2_0),.clk(gclk));
	jdff dff_B_eNxLlYtU5_0(.din(w_dff_B_ZGRaC1kQ2_0),.dout(w_dff_B_eNxLlYtU5_0),.clk(gclk));
	jdff dff_B_oNVlvjEm9_0(.din(w_dff_B_eNxLlYtU5_0),.dout(w_dff_B_oNVlvjEm9_0),.clk(gclk));
	jdff dff_B_ypipYVnK0_0(.din(w_dff_B_oNVlvjEm9_0),.dout(w_dff_B_ypipYVnK0_0),.clk(gclk));
	jdff dff_B_G3wt2Ihy5_0(.din(w_dff_B_ypipYVnK0_0),.dout(w_dff_B_G3wt2Ihy5_0),.clk(gclk));
	jdff dff_B_LbuN2S981_0(.din(w_dff_B_G3wt2Ihy5_0),.dout(w_dff_B_LbuN2S981_0),.clk(gclk));
	jdff dff_B_TW3FMs1W4_0(.din(w_dff_B_LbuN2S981_0),.dout(w_dff_B_TW3FMs1W4_0),.clk(gclk));
	jdff dff_B_qKGSCiFM8_0(.din(w_dff_B_TW3FMs1W4_0),.dout(w_dff_B_qKGSCiFM8_0),.clk(gclk));
	jdff dff_B_0Sd2KXnC8_0(.din(w_dff_B_qKGSCiFM8_0),.dout(w_dff_B_0Sd2KXnC8_0),.clk(gclk));
	jdff dff_B_QNWKoSPe6_0(.din(w_dff_B_0Sd2KXnC8_0),.dout(w_dff_B_QNWKoSPe6_0),.clk(gclk));
	jdff dff_B_xLmYmdXH5_0(.din(w_dff_B_QNWKoSPe6_0),.dout(w_dff_B_xLmYmdXH5_0),.clk(gclk));
	jdff dff_B_hYBJVPYE0_0(.din(w_dff_B_xLmYmdXH5_0),.dout(w_dff_B_hYBJVPYE0_0),.clk(gclk));
	jdff dff_B_XMqHatDK8_0(.din(w_dff_B_hYBJVPYE0_0),.dout(w_dff_B_XMqHatDK8_0),.clk(gclk));
	jdff dff_B_f5WRGiSU7_0(.din(w_dff_B_XMqHatDK8_0),.dout(w_dff_B_f5WRGiSU7_0),.clk(gclk));
	jdff dff_B_YBjguptx0_0(.din(w_dff_B_f5WRGiSU7_0),.dout(w_dff_B_YBjguptx0_0),.clk(gclk));
	jdff dff_B_cFs0iOoL4_0(.din(w_dff_B_YBjguptx0_0),.dout(w_dff_B_cFs0iOoL4_0),.clk(gclk));
	jdff dff_B_kzJ4k9HD4_0(.din(w_dff_B_cFs0iOoL4_0),.dout(w_dff_B_kzJ4k9HD4_0),.clk(gclk));
	jdff dff_B_vHReqyac4_0(.din(w_dff_B_kzJ4k9HD4_0),.dout(w_dff_B_vHReqyac4_0),.clk(gclk));
	jdff dff_B_lXj30V6V2_0(.din(w_dff_B_vHReqyac4_0),.dout(w_dff_B_lXj30V6V2_0),.clk(gclk));
	jdff dff_B_Yr3uBJhz8_0(.din(w_dff_B_lXj30V6V2_0),.dout(w_dff_B_Yr3uBJhz8_0),.clk(gclk));
	jdff dff_B_P8fyoIaN1_0(.din(w_dff_B_Yr3uBJhz8_0),.dout(w_dff_B_P8fyoIaN1_0),.clk(gclk));
	jdff dff_B_ooeeHe1Z9_0(.din(w_dff_B_P8fyoIaN1_0),.dout(w_dff_B_ooeeHe1Z9_0),.clk(gclk));
	jdff dff_B_1qN8zhd62_0(.din(w_dff_B_ooeeHe1Z9_0),.dout(w_dff_B_1qN8zhd62_0),.clk(gclk));
	jdff dff_B_q8WGGNTC8_0(.din(w_dff_B_1qN8zhd62_0),.dout(w_dff_B_q8WGGNTC8_0),.clk(gclk));
	jdff dff_B_Ofpdrk672_0(.din(w_dff_B_q8WGGNTC8_0),.dout(w_dff_B_Ofpdrk672_0),.clk(gclk));
	jdff dff_B_dmE7wIib9_0(.din(w_dff_B_Ofpdrk672_0),.dout(w_dff_B_dmE7wIib9_0),.clk(gclk));
	jdff dff_B_WCARSoGH8_0(.din(w_dff_B_dmE7wIib9_0),.dout(w_dff_B_WCARSoGH8_0),.clk(gclk));
	jdff dff_B_RMTzlVVX2_0(.din(w_dff_B_WCARSoGH8_0),.dout(w_dff_B_RMTzlVVX2_0),.clk(gclk));
	jdff dff_B_gPiENw7M9_0(.din(w_dff_B_RMTzlVVX2_0),.dout(w_dff_B_gPiENw7M9_0),.clk(gclk));
	jdff dff_B_cx2KtWNM1_0(.din(w_dff_B_gPiENw7M9_0),.dout(w_dff_B_cx2KtWNM1_0),.clk(gclk));
	jdff dff_B_jgNPEzhL6_0(.din(w_dff_B_cx2KtWNM1_0),.dout(w_dff_B_jgNPEzhL6_0),.clk(gclk));
	jdff dff_B_vyv3QZRw0_0(.din(w_dff_B_jgNPEzhL6_0),.dout(w_dff_B_vyv3QZRw0_0),.clk(gclk));
	jdff dff_B_ATufaRAT8_0(.din(w_dff_B_vyv3QZRw0_0),.dout(w_dff_B_ATufaRAT8_0),.clk(gclk));
	jdff dff_B_RMFUD2fO6_0(.din(w_dff_B_ATufaRAT8_0),.dout(w_dff_B_RMFUD2fO6_0),.clk(gclk));
	jdff dff_B_IGVwytqN2_0(.din(w_dff_B_RMFUD2fO6_0),.dout(w_dff_B_IGVwytqN2_0),.clk(gclk));
	jdff dff_B_VkCKYLEW6_0(.din(w_dff_B_IGVwytqN2_0),.dout(w_dff_B_VkCKYLEW6_0),.clk(gclk));
	jdff dff_B_p465ngL27_0(.din(w_dff_B_VkCKYLEW6_0),.dout(w_dff_B_p465ngL27_0),.clk(gclk));
	jdff dff_B_44xOJOdM7_0(.din(w_dff_B_p465ngL27_0),.dout(w_dff_B_44xOJOdM7_0),.clk(gclk));
	jdff dff_B_UGl0cc1T6_0(.din(w_dff_B_44xOJOdM7_0),.dout(w_dff_B_UGl0cc1T6_0),.clk(gclk));
	jdff dff_B_fBiDhWsS6_0(.din(w_dff_B_UGl0cc1T6_0),.dout(w_dff_B_fBiDhWsS6_0),.clk(gclk));
	jdff dff_B_w8lFOCaz9_0(.din(w_dff_B_fBiDhWsS6_0),.dout(w_dff_B_w8lFOCaz9_0),.clk(gclk));
	jdff dff_B_fKUl863m0_0(.din(w_dff_B_w8lFOCaz9_0),.dout(w_dff_B_fKUl863m0_0),.clk(gclk));
	jdff dff_B_UYLDZLJM4_0(.din(w_dff_B_fKUl863m0_0),.dout(w_dff_B_UYLDZLJM4_0),.clk(gclk));
	jdff dff_B_WTuT0sRw7_0(.din(w_dff_B_UYLDZLJM4_0),.dout(w_dff_B_WTuT0sRw7_0),.clk(gclk));
	jdff dff_B_D1pBStHq0_0(.din(w_dff_B_WTuT0sRw7_0),.dout(w_dff_B_D1pBStHq0_0),.clk(gclk));
	jdff dff_B_N7vmbMkQ0_0(.din(w_dff_B_D1pBStHq0_0),.dout(w_dff_B_N7vmbMkQ0_0),.clk(gclk));
	jdff dff_B_3nxITtqi1_1(.din(n906),.dout(w_dff_B_3nxITtqi1_1),.clk(gclk));
	jdff dff_B_OY2rNriK2_1(.din(w_dff_B_3nxITtqi1_1),.dout(w_dff_B_OY2rNriK2_1),.clk(gclk));
	jdff dff_B_KxDJtCsC5_1(.din(w_dff_B_OY2rNriK2_1),.dout(w_dff_B_KxDJtCsC5_1),.clk(gclk));
	jdff dff_B_MRznJZ2V8_1(.din(w_dff_B_KxDJtCsC5_1),.dout(w_dff_B_MRznJZ2V8_1),.clk(gclk));
	jdff dff_B_6hJao4te2_1(.din(w_dff_B_MRznJZ2V8_1),.dout(w_dff_B_6hJao4te2_1),.clk(gclk));
	jdff dff_B_aNDxRmSo2_1(.din(w_dff_B_6hJao4te2_1),.dout(w_dff_B_aNDxRmSo2_1),.clk(gclk));
	jdff dff_B_9mDzCuTh4_1(.din(w_dff_B_aNDxRmSo2_1),.dout(w_dff_B_9mDzCuTh4_1),.clk(gclk));
	jdff dff_B_TkGFrCbe0_1(.din(w_dff_B_9mDzCuTh4_1),.dout(w_dff_B_TkGFrCbe0_1),.clk(gclk));
	jdff dff_B_MvI5NZum1_1(.din(w_dff_B_TkGFrCbe0_1),.dout(w_dff_B_MvI5NZum1_1),.clk(gclk));
	jdff dff_B_OvDfYURa0_1(.din(w_dff_B_MvI5NZum1_1),.dout(w_dff_B_OvDfYURa0_1),.clk(gclk));
	jdff dff_B_seEix5eN4_1(.din(w_dff_B_OvDfYURa0_1),.dout(w_dff_B_seEix5eN4_1),.clk(gclk));
	jdff dff_B_YGK7MZPn7_1(.din(w_dff_B_seEix5eN4_1),.dout(w_dff_B_YGK7MZPn7_1),.clk(gclk));
	jdff dff_B_YMcqpjlG1_1(.din(w_dff_B_YGK7MZPn7_1),.dout(w_dff_B_YMcqpjlG1_1),.clk(gclk));
	jdff dff_B_oR5AoGfk2_1(.din(w_dff_B_YMcqpjlG1_1),.dout(w_dff_B_oR5AoGfk2_1),.clk(gclk));
	jdff dff_B_M2eZ4DfO4_1(.din(w_dff_B_oR5AoGfk2_1),.dout(w_dff_B_M2eZ4DfO4_1),.clk(gclk));
	jdff dff_B_UJmA2lav7_1(.din(w_dff_B_M2eZ4DfO4_1),.dout(w_dff_B_UJmA2lav7_1),.clk(gclk));
	jdff dff_B_hfkTVK7o6_1(.din(w_dff_B_UJmA2lav7_1),.dout(w_dff_B_hfkTVK7o6_1),.clk(gclk));
	jdff dff_B_EIInKr7E9_1(.din(w_dff_B_hfkTVK7o6_1),.dout(w_dff_B_EIInKr7E9_1),.clk(gclk));
	jdff dff_B_b9XhOSpz8_1(.din(w_dff_B_EIInKr7E9_1),.dout(w_dff_B_b9XhOSpz8_1),.clk(gclk));
	jdff dff_B_i8DE75Ze0_1(.din(w_dff_B_b9XhOSpz8_1),.dout(w_dff_B_i8DE75Ze0_1),.clk(gclk));
	jdff dff_B_etvdKZ7e5_1(.din(w_dff_B_i8DE75Ze0_1),.dout(w_dff_B_etvdKZ7e5_1),.clk(gclk));
	jdff dff_B_xT6XSek77_1(.din(w_dff_B_etvdKZ7e5_1),.dout(w_dff_B_xT6XSek77_1),.clk(gclk));
	jdff dff_B_N8ze5nwB4_1(.din(w_dff_B_xT6XSek77_1),.dout(w_dff_B_N8ze5nwB4_1),.clk(gclk));
	jdff dff_B_2fPf9uIc4_1(.din(w_dff_B_N8ze5nwB4_1),.dout(w_dff_B_2fPf9uIc4_1),.clk(gclk));
	jdff dff_B_pWiraKkQ6_1(.din(w_dff_B_2fPf9uIc4_1),.dout(w_dff_B_pWiraKkQ6_1),.clk(gclk));
	jdff dff_B_hxGFuNEE1_1(.din(w_dff_B_pWiraKkQ6_1),.dout(w_dff_B_hxGFuNEE1_1),.clk(gclk));
	jdff dff_B_9uXZVZ7o6_1(.din(w_dff_B_hxGFuNEE1_1),.dout(w_dff_B_9uXZVZ7o6_1),.clk(gclk));
	jdff dff_B_2n8yYbkH4_1(.din(w_dff_B_9uXZVZ7o6_1),.dout(w_dff_B_2n8yYbkH4_1),.clk(gclk));
	jdff dff_B_qGvwWjX74_1(.din(w_dff_B_2n8yYbkH4_1),.dout(w_dff_B_qGvwWjX74_1),.clk(gclk));
	jdff dff_B_570ADOlS3_1(.din(w_dff_B_qGvwWjX74_1),.dout(w_dff_B_570ADOlS3_1),.clk(gclk));
	jdff dff_B_fGGrn6YP6_1(.din(w_dff_B_570ADOlS3_1),.dout(w_dff_B_fGGrn6YP6_1),.clk(gclk));
	jdff dff_B_JhhTo1ZE2_1(.din(w_dff_B_fGGrn6YP6_1),.dout(w_dff_B_JhhTo1ZE2_1),.clk(gclk));
	jdff dff_B_g5NZvvAt8_1(.din(w_dff_B_JhhTo1ZE2_1),.dout(w_dff_B_g5NZvvAt8_1),.clk(gclk));
	jdff dff_B_LaGgbmqZ2_1(.din(w_dff_B_g5NZvvAt8_1),.dout(w_dff_B_LaGgbmqZ2_1),.clk(gclk));
	jdff dff_B_PAlhKosg6_1(.din(w_dff_B_LaGgbmqZ2_1),.dout(w_dff_B_PAlhKosg6_1),.clk(gclk));
	jdff dff_B_gyA1OFlq0_1(.din(w_dff_B_PAlhKosg6_1),.dout(w_dff_B_gyA1OFlq0_1),.clk(gclk));
	jdff dff_B_ovgXJbXd2_1(.din(w_dff_B_gyA1OFlq0_1),.dout(w_dff_B_ovgXJbXd2_1),.clk(gclk));
	jdff dff_B_A5e2ravW8_1(.din(w_dff_B_ovgXJbXd2_1),.dout(w_dff_B_A5e2ravW8_1),.clk(gclk));
	jdff dff_B_6Q0caIYh0_1(.din(w_dff_B_A5e2ravW8_1),.dout(w_dff_B_6Q0caIYh0_1),.clk(gclk));
	jdff dff_B_TJLpKMo57_1(.din(w_dff_B_6Q0caIYh0_1),.dout(w_dff_B_TJLpKMo57_1),.clk(gclk));
	jdff dff_B_Iwu02DDs8_1(.din(w_dff_B_TJLpKMo57_1),.dout(w_dff_B_Iwu02DDs8_1),.clk(gclk));
	jdff dff_B_sskXV6pq5_1(.din(w_dff_B_Iwu02DDs8_1),.dout(w_dff_B_sskXV6pq5_1),.clk(gclk));
	jdff dff_B_RixVdW8j2_1(.din(w_dff_B_sskXV6pq5_1),.dout(w_dff_B_RixVdW8j2_1),.clk(gclk));
	jdff dff_B_CDB3Pimm3_1(.din(w_dff_B_RixVdW8j2_1),.dout(w_dff_B_CDB3Pimm3_1),.clk(gclk));
	jdff dff_B_TsnxBlJj6_1(.din(w_dff_B_CDB3Pimm3_1),.dout(w_dff_B_TsnxBlJj6_1),.clk(gclk));
	jdff dff_B_gnt9diSQ7_1(.din(w_dff_B_TsnxBlJj6_1),.dout(w_dff_B_gnt9diSQ7_1),.clk(gclk));
	jdff dff_B_ahDyzhe43_1(.din(w_dff_B_gnt9diSQ7_1),.dout(w_dff_B_ahDyzhe43_1),.clk(gclk));
	jdff dff_B_fl9kYm1H7_1(.din(w_dff_B_ahDyzhe43_1),.dout(w_dff_B_fl9kYm1H7_1),.clk(gclk));
	jdff dff_B_KySJAlVy8_1(.din(w_dff_B_fl9kYm1H7_1),.dout(w_dff_B_KySJAlVy8_1),.clk(gclk));
	jdff dff_B_kGAcvuc99_1(.din(w_dff_B_KySJAlVy8_1),.dout(w_dff_B_kGAcvuc99_1),.clk(gclk));
	jdff dff_B_IBE3bsOk7_1(.din(w_dff_B_kGAcvuc99_1),.dout(w_dff_B_IBE3bsOk7_1),.clk(gclk));
	jdff dff_B_U3epGkXT2_1(.din(w_dff_B_IBE3bsOk7_1),.dout(w_dff_B_U3epGkXT2_1),.clk(gclk));
	jdff dff_B_K1CLJtb48_1(.din(w_dff_B_U3epGkXT2_1),.dout(w_dff_B_K1CLJtb48_1),.clk(gclk));
	jdff dff_B_Rqg5JfTZ5_1(.din(w_dff_B_K1CLJtb48_1),.dout(w_dff_B_Rqg5JfTZ5_1),.clk(gclk));
	jdff dff_B_1hafOUpw8_1(.din(w_dff_B_Rqg5JfTZ5_1),.dout(w_dff_B_1hafOUpw8_1),.clk(gclk));
	jdff dff_B_kc0k9wSE7_1(.din(w_dff_B_1hafOUpw8_1),.dout(w_dff_B_kc0k9wSE7_1),.clk(gclk));
	jdff dff_B_vtFiJc4h0_1(.din(w_dff_B_kc0k9wSE7_1),.dout(w_dff_B_vtFiJc4h0_1),.clk(gclk));
	jdff dff_B_tEBBFEtC9_1(.din(w_dff_B_vtFiJc4h0_1),.dout(w_dff_B_tEBBFEtC9_1),.clk(gclk));
	jdff dff_B_0nZBMp6Y4_1(.din(w_dff_B_tEBBFEtC9_1),.dout(w_dff_B_0nZBMp6Y4_1),.clk(gclk));
	jdff dff_B_zJ7KyBYy5_1(.din(w_dff_B_0nZBMp6Y4_1),.dout(w_dff_B_zJ7KyBYy5_1),.clk(gclk));
	jdff dff_B_gsENW5VE5_1(.din(w_dff_B_zJ7KyBYy5_1),.dout(w_dff_B_gsENW5VE5_1),.clk(gclk));
	jdff dff_B_z2nQMeJU1_1(.din(w_dff_B_gsENW5VE5_1),.dout(w_dff_B_z2nQMeJU1_1),.clk(gclk));
	jdff dff_B_ccxG0Q207_1(.din(w_dff_B_z2nQMeJU1_1),.dout(w_dff_B_ccxG0Q207_1),.clk(gclk));
	jdff dff_B_o24hhAGX8_1(.din(w_dff_B_ccxG0Q207_1),.dout(w_dff_B_o24hhAGX8_1),.clk(gclk));
	jdff dff_B_NYlA2kK67_1(.din(w_dff_B_o24hhAGX8_1),.dout(w_dff_B_NYlA2kK67_1),.clk(gclk));
	jdff dff_B_z2U4Prsj6_1(.din(w_dff_B_NYlA2kK67_1),.dout(w_dff_B_z2U4Prsj6_1),.clk(gclk));
	jdff dff_B_y6G2xfc01_1(.din(w_dff_B_z2U4Prsj6_1),.dout(w_dff_B_y6G2xfc01_1),.clk(gclk));
	jdff dff_B_CAzTvFjT7_1(.din(w_dff_B_y6G2xfc01_1),.dout(w_dff_B_CAzTvFjT7_1),.clk(gclk));
	jdff dff_B_HZtwRYYs1_1(.din(w_dff_B_CAzTvFjT7_1),.dout(w_dff_B_HZtwRYYs1_1),.clk(gclk));
	jdff dff_B_2wOj47B74_1(.din(w_dff_B_HZtwRYYs1_1),.dout(w_dff_B_2wOj47B74_1),.clk(gclk));
	jdff dff_B_3Sqezcf91_1(.din(w_dff_B_2wOj47B74_1),.dout(w_dff_B_3Sqezcf91_1),.clk(gclk));
	jdff dff_B_4jvZRNPu1_1(.din(w_dff_B_3Sqezcf91_1),.dout(w_dff_B_4jvZRNPu1_1),.clk(gclk));
	jdff dff_B_zNbb8qII5_1(.din(w_dff_B_4jvZRNPu1_1),.dout(w_dff_B_zNbb8qII5_1),.clk(gclk));
	jdff dff_B_6ySqU7NU6_1(.din(w_dff_B_zNbb8qII5_1),.dout(w_dff_B_6ySqU7NU6_1),.clk(gclk));
	jdff dff_B_4sa4L1va5_1(.din(w_dff_B_6ySqU7NU6_1),.dout(w_dff_B_4sa4L1va5_1),.clk(gclk));
	jdff dff_B_bVK9UKFi6_1(.din(w_dff_B_4sa4L1va5_1),.dout(w_dff_B_bVK9UKFi6_1),.clk(gclk));
	jdff dff_B_mLXAfc796_1(.din(w_dff_B_bVK9UKFi6_1),.dout(w_dff_B_mLXAfc796_1),.clk(gclk));
	jdff dff_B_TRjy6evf4_1(.din(w_dff_B_mLXAfc796_1),.dout(w_dff_B_TRjy6evf4_1),.clk(gclk));
	jdff dff_B_QDBbrq6c2_1(.din(w_dff_B_TRjy6evf4_1),.dout(w_dff_B_QDBbrq6c2_1),.clk(gclk));
	jdff dff_B_fvWpofjd2_1(.din(w_dff_B_QDBbrq6c2_1),.dout(w_dff_B_fvWpofjd2_1),.clk(gclk));
	jdff dff_B_pM9LgozB4_1(.din(w_dff_B_fvWpofjd2_1),.dout(w_dff_B_pM9LgozB4_1),.clk(gclk));
	jdff dff_B_LswJxzVi3_1(.din(w_dff_B_pM9LgozB4_1),.dout(w_dff_B_LswJxzVi3_1),.clk(gclk));
	jdff dff_B_KBOyUbQG1_1(.din(w_dff_B_LswJxzVi3_1),.dout(w_dff_B_KBOyUbQG1_1),.clk(gclk));
	jdff dff_B_axP6W0ux6_1(.din(w_dff_B_KBOyUbQG1_1),.dout(w_dff_B_axP6W0ux6_1),.clk(gclk));
	jdff dff_B_1eQjlJ7B5_1(.din(w_dff_B_axP6W0ux6_1),.dout(w_dff_B_1eQjlJ7B5_1),.clk(gclk));
	jdff dff_B_LPntHGIh3_1(.din(w_dff_B_1eQjlJ7B5_1),.dout(w_dff_B_LPntHGIh3_1),.clk(gclk));
	jdff dff_B_utDSKdr27_1(.din(w_dff_B_LPntHGIh3_1),.dout(w_dff_B_utDSKdr27_1),.clk(gclk));
	jdff dff_B_9OfuBhph8_0(.din(n907),.dout(w_dff_B_9OfuBhph8_0),.clk(gclk));
	jdff dff_B_fSvMGx083_0(.din(w_dff_B_9OfuBhph8_0),.dout(w_dff_B_fSvMGx083_0),.clk(gclk));
	jdff dff_B_PbQQjmcP1_0(.din(w_dff_B_fSvMGx083_0),.dout(w_dff_B_PbQQjmcP1_0),.clk(gclk));
	jdff dff_B_UmIzH0ra0_0(.din(w_dff_B_PbQQjmcP1_0),.dout(w_dff_B_UmIzH0ra0_0),.clk(gclk));
	jdff dff_B_2EOuS1kW7_0(.din(w_dff_B_UmIzH0ra0_0),.dout(w_dff_B_2EOuS1kW7_0),.clk(gclk));
	jdff dff_B_HJjDZQ491_0(.din(w_dff_B_2EOuS1kW7_0),.dout(w_dff_B_HJjDZQ491_0),.clk(gclk));
	jdff dff_B_FsIxBUry9_0(.din(w_dff_B_HJjDZQ491_0),.dout(w_dff_B_FsIxBUry9_0),.clk(gclk));
	jdff dff_B_QdOryrZ81_0(.din(w_dff_B_FsIxBUry9_0),.dout(w_dff_B_QdOryrZ81_0),.clk(gclk));
	jdff dff_B_qDO5vPBl7_0(.din(w_dff_B_QdOryrZ81_0),.dout(w_dff_B_qDO5vPBl7_0),.clk(gclk));
	jdff dff_B_tszjXaEA4_0(.din(w_dff_B_qDO5vPBl7_0),.dout(w_dff_B_tszjXaEA4_0),.clk(gclk));
	jdff dff_B_wlJRwORz2_0(.din(w_dff_B_tszjXaEA4_0),.dout(w_dff_B_wlJRwORz2_0),.clk(gclk));
	jdff dff_B_SK5LwVko8_0(.din(w_dff_B_wlJRwORz2_0),.dout(w_dff_B_SK5LwVko8_0),.clk(gclk));
	jdff dff_B_YeYxrDAV9_0(.din(w_dff_B_SK5LwVko8_0),.dout(w_dff_B_YeYxrDAV9_0),.clk(gclk));
	jdff dff_B_5Qp7hdX02_0(.din(w_dff_B_YeYxrDAV9_0),.dout(w_dff_B_5Qp7hdX02_0),.clk(gclk));
	jdff dff_B_8ICqi3Ox9_0(.din(w_dff_B_5Qp7hdX02_0),.dout(w_dff_B_8ICqi3Ox9_0),.clk(gclk));
	jdff dff_B_vyJ9grxt2_0(.din(w_dff_B_8ICqi3Ox9_0),.dout(w_dff_B_vyJ9grxt2_0),.clk(gclk));
	jdff dff_B_bfs9zKE79_0(.din(w_dff_B_vyJ9grxt2_0),.dout(w_dff_B_bfs9zKE79_0),.clk(gclk));
	jdff dff_B_bxdeaFXv6_0(.din(w_dff_B_bfs9zKE79_0),.dout(w_dff_B_bxdeaFXv6_0),.clk(gclk));
	jdff dff_B_QsY6qUnX4_0(.din(w_dff_B_bxdeaFXv6_0),.dout(w_dff_B_QsY6qUnX4_0),.clk(gclk));
	jdff dff_B_j59beE0U8_0(.din(w_dff_B_QsY6qUnX4_0),.dout(w_dff_B_j59beE0U8_0),.clk(gclk));
	jdff dff_B_z0hlPxAr6_0(.din(w_dff_B_j59beE0U8_0),.dout(w_dff_B_z0hlPxAr6_0),.clk(gclk));
	jdff dff_B_4tL7UEOV2_0(.din(w_dff_B_z0hlPxAr6_0),.dout(w_dff_B_4tL7UEOV2_0),.clk(gclk));
	jdff dff_B_1dkoGQx85_0(.din(w_dff_B_4tL7UEOV2_0),.dout(w_dff_B_1dkoGQx85_0),.clk(gclk));
	jdff dff_B_lm0gTiO35_0(.din(w_dff_B_1dkoGQx85_0),.dout(w_dff_B_lm0gTiO35_0),.clk(gclk));
	jdff dff_B_srwZ13vA8_0(.din(w_dff_B_lm0gTiO35_0),.dout(w_dff_B_srwZ13vA8_0),.clk(gclk));
	jdff dff_B_T9q9rx4k3_0(.din(w_dff_B_srwZ13vA8_0),.dout(w_dff_B_T9q9rx4k3_0),.clk(gclk));
	jdff dff_B_S07tiac19_0(.din(w_dff_B_T9q9rx4k3_0),.dout(w_dff_B_S07tiac19_0),.clk(gclk));
	jdff dff_B_xUgD5UNb5_0(.din(w_dff_B_S07tiac19_0),.dout(w_dff_B_xUgD5UNb5_0),.clk(gclk));
	jdff dff_B_A6fW8pRB0_0(.din(w_dff_B_xUgD5UNb5_0),.dout(w_dff_B_A6fW8pRB0_0),.clk(gclk));
	jdff dff_B_crgzXCqM1_0(.din(w_dff_B_A6fW8pRB0_0),.dout(w_dff_B_crgzXCqM1_0),.clk(gclk));
	jdff dff_B_aIqpclKv9_0(.din(w_dff_B_crgzXCqM1_0),.dout(w_dff_B_aIqpclKv9_0),.clk(gclk));
	jdff dff_B_rYpOO1Mu6_0(.din(w_dff_B_aIqpclKv9_0),.dout(w_dff_B_rYpOO1Mu6_0),.clk(gclk));
	jdff dff_B_vm8WZ0yM2_0(.din(w_dff_B_rYpOO1Mu6_0),.dout(w_dff_B_vm8WZ0yM2_0),.clk(gclk));
	jdff dff_B_L3hDfd8S0_0(.din(w_dff_B_vm8WZ0yM2_0),.dout(w_dff_B_L3hDfd8S0_0),.clk(gclk));
	jdff dff_B_wMRyWpiD0_0(.din(w_dff_B_L3hDfd8S0_0),.dout(w_dff_B_wMRyWpiD0_0),.clk(gclk));
	jdff dff_B_Vf80f1Lw3_0(.din(w_dff_B_wMRyWpiD0_0),.dout(w_dff_B_Vf80f1Lw3_0),.clk(gclk));
	jdff dff_B_zraub0fj5_0(.din(w_dff_B_Vf80f1Lw3_0),.dout(w_dff_B_zraub0fj5_0),.clk(gclk));
	jdff dff_B_uY4V9vDI4_0(.din(w_dff_B_zraub0fj5_0),.dout(w_dff_B_uY4V9vDI4_0),.clk(gclk));
	jdff dff_B_hPLKAhbe9_0(.din(w_dff_B_uY4V9vDI4_0),.dout(w_dff_B_hPLKAhbe9_0),.clk(gclk));
	jdff dff_B_XeI2PEdj6_0(.din(w_dff_B_hPLKAhbe9_0),.dout(w_dff_B_XeI2PEdj6_0),.clk(gclk));
	jdff dff_B_byRcTbez4_0(.din(w_dff_B_XeI2PEdj6_0),.dout(w_dff_B_byRcTbez4_0),.clk(gclk));
	jdff dff_B_aUxFGFSR6_0(.din(w_dff_B_byRcTbez4_0),.dout(w_dff_B_aUxFGFSR6_0),.clk(gclk));
	jdff dff_B_GONssTcG3_0(.din(w_dff_B_aUxFGFSR6_0),.dout(w_dff_B_GONssTcG3_0),.clk(gclk));
	jdff dff_B_hZS5ek4N0_0(.din(w_dff_B_GONssTcG3_0),.dout(w_dff_B_hZS5ek4N0_0),.clk(gclk));
	jdff dff_B_mYEE4hLh4_0(.din(w_dff_B_hZS5ek4N0_0),.dout(w_dff_B_mYEE4hLh4_0),.clk(gclk));
	jdff dff_B_utaoV4oG5_0(.din(w_dff_B_mYEE4hLh4_0),.dout(w_dff_B_utaoV4oG5_0),.clk(gclk));
	jdff dff_B_l9AqLoT11_0(.din(w_dff_B_utaoV4oG5_0),.dout(w_dff_B_l9AqLoT11_0),.clk(gclk));
	jdff dff_B_uexlpWaD7_0(.din(w_dff_B_l9AqLoT11_0),.dout(w_dff_B_uexlpWaD7_0),.clk(gclk));
	jdff dff_B_3UwJZ2Us6_0(.din(w_dff_B_uexlpWaD7_0),.dout(w_dff_B_3UwJZ2Us6_0),.clk(gclk));
	jdff dff_B_ph05CXZ16_0(.din(w_dff_B_3UwJZ2Us6_0),.dout(w_dff_B_ph05CXZ16_0),.clk(gclk));
	jdff dff_B_CW0eQWU43_0(.din(w_dff_B_ph05CXZ16_0),.dout(w_dff_B_CW0eQWU43_0),.clk(gclk));
	jdff dff_B_SmHGQilD7_0(.din(w_dff_B_CW0eQWU43_0),.dout(w_dff_B_SmHGQilD7_0),.clk(gclk));
	jdff dff_B_Rzn23w105_0(.din(w_dff_B_SmHGQilD7_0),.dout(w_dff_B_Rzn23w105_0),.clk(gclk));
	jdff dff_B_QnCJ3FFM2_0(.din(w_dff_B_Rzn23w105_0),.dout(w_dff_B_QnCJ3FFM2_0),.clk(gclk));
	jdff dff_B_egwZnSYa0_0(.din(w_dff_B_QnCJ3FFM2_0),.dout(w_dff_B_egwZnSYa0_0),.clk(gclk));
	jdff dff_B_0yDvGr9g3_0(.din(w_dff_B_egwZnSYa0_0),.dout(w_dff_B_0yDvGr9g3_0),.clk(gclk));
	jdff dff_B_0598e1ao2_0(.din(w_dff_B_0yDvGr9g3_0),.dout(w_dff_B_0598e1ao2_0),.clk(gclk));
	jdff dff_B_QSoSxXWZ6_0(.din(w_dff_B_0598e1ao2_0),.dout(w_dff_B_QSoSxXWZ6_0),.clk(gclk));
	jdff dff_B_VdjDn69y3_0(.din(w_dff_B_QSoSxXWZ6_0),.dout(w_dff_B_VdjDn69y3_0),.clk(gclk));
	jdff dff_B_fTT29wPF9_0(.din(w_dff_B_VdjDn69y3_0),.dout(w_dff_B_fTT29wPF9_0),.clk(gclk));
	jdff dff_B_zxfVbPlO8_0(.din(w_dff_B_fTT29wPF9_0),.dout(w_dff_B_zxfVbPlO8_0),.clk(gclk));
	jdff dff_B_TA34UdTz7_0(.din(w_dff_B_zxfVbPlO8_0),.dout(w_dff_B_TA34UdTz7_0),.clk(gclk));
	jdff dff_B_MoN52Izk1_0(.din(w_dff_B_TA34UdTz7_0),.dout(w_dff_B_MoN52Izk1_0),.clk(gclk));
	jdff dff_B_Sor7zlqY9_0(.din(w_dff_B_MoN52Izk1_0),.dout(w_dff_B_Sor7zlqY9_0),.clk(gclk));
	jdff dff_B_ZANXWw0N6_0(.din(w_dff_B_Sor7zlqY9_0),.dout(w_dff_B_ZANXWw0N6_0),.clk(gclk));
	jdff dff_B_qkDf3kKX9_0(.din(w_dff_B_ZANXWw0N6_0),.dout(w_dff_B_qkDf3kKX9_0),.clk(gclk));
	jdff dff_B_b1Qaza8E9_0(.din(w_dff_B_qkDf3kKX9_0),.dout(w_dff_B_b1Qaza8E9_0),.clk(gclk));
	jdff dff_B_cpmt8CvA4_0(.din(w_dff_B_b1Qaza8E9_0),.dout(w_dff_B_cpmt8CvA4_0),.clk(gclk));
	jdff dff_B_SHVva91F4_0(.din(w_dff_B_cpmt8CvA4_0),.dout(w_dff_B_SHVva91F4_0),.clk(gclk));
	jdff dff_B_r6PKqLfI1_0(.din(w_dff_B_SHVva91F4_0),.dout(w_dff_B_r6PKqLfI1_0),.clk(gclk));
	jdff dff_B_AAvzp0KW5_0(.din(w_dff_B_r6PKqLfI1_0),.dout(w_dff_B_AAvzp0KW5_0),.clk(gclk));
	jdff dff_B_p3uAXoKr8_0(.din(w_dff_B_AAvzp0KW5_0),.dout(w_dff_B_p3uAXoKr8_0),.clk(gclk));
	jdff dff_B_WmF1feBH6_0(.din(w_dff_B_p3uAXoKr8_0),.dout(w_dff_B_WmF1feBH6_0),.clk(gclk));
	jdff dff_B_gIrCgn8u6_0(.din(w_dff_B_WmF1feBH6_0),.dout(w_dff_B_gIrCgn8u6_0),.clk(gclk));
	jdff dff_B_SwLUpiyP0_0(.din(w_dff_B_gIrCgn8u6_0),.dout(w_dff_B_SwLUpiyP0_0),.clk(gclk));
	jdff dff_B_XHHSkZBs7_0(.din(w_dff_B_SwLUpiyP0_0),.dout(w_dff_B_XHHSkZBs7_0),.clk(gclk));
	jdff dff_B_ZmfgwsEv4_0(.din(w_dff_B_XHHSkZBs7_0),.dout(w_dff_B_ZmfgwsEv4_0),.clk(gclk));
	jdff dff_B_fJU91JOB5_0(.din(w_dff_B_ZmfgwsEv4_0),.dout(w_dff_B_fJU91JOB5_0),.clk(gclk));
	jdff dff_B_SK2pSLPr2_0(.din(w_dff_B_fJU91JOB5_0),.dout(w_dff_B_SK2pSLPr2_0),.clk(gclk));
	jdff dff_B_KSDyklnh5_0(.din(w_dff_B_SK2pSLPr2_0),.dout(w_dff_B_KSDyklnh5_0),.clk(gclk));
	jdff dff_B_AfyInHg87_0(.din(w_dff_B_KSDyklnh5_0),.dout(w_dff_B_AfyInHg87_0),.clk(gclk));
	jdff dff_B_bIh4yIkm9_0(.din(w_dff_B_AfyInHg87_0),.dout(w_dff_B_bIh4yIkm9_0),.clk(gclk));
	jdff dff_B_bD2ZHqTj2_0(.din(w_dff_B_bIh4yIkm9_0),.dout(w_dff_B_bD2ZHqTj2_0),.clk(gclk));
	jdff dff_B_hc8SK1Fi3_0(.din(w_dff_B_bD2ZHqTj2_0),.dout(w_dff_B_hc8SK1Fi3_0),.clk(gclk));
	jdff dff_B_PPPR0yO03_0(.din(w_dff_B_hc8SK1Fi3_0),.dout(w_dff_B_PPPR0yO03_0),.clk(gclk));
	jdff dff_B_NxxGUlsv8_0(.din(w_dff_B_PPPR0yO03_0),.dout(w_dff_B_NxxGUlsv8_0),.clk(gclk));
	jdff dff_B_dfcAYDfk0_0(.din(w_dff_B_NxxGUlsv8_0),.dout(w_dff_B_dfcAYDfk0_0),.clk(gclk));
	jdff dff_B_qcSVTYBt6_1(.din(n900),.dout(w_dff_B_qcSVTYBt6_1),.clk(gclk));
	jdff dff_B_kCUZfYTp3_1(.din(w_dff_B_qcSVTYBt6_1),.dout(w_dff_B_kCUZfYTp3_1),.clk(gclk));
	jdff dff_B_l9JmYZuV0_1(.din(w_dff_B_kCUZfYTp3_1),.dout(w_dff_B_l9JmYZuV0_1),.clk(gclk));
	jdff dff_B_MUTLEILN0_1(.din(w_dff_B_l9JmYZuV0_1),.dout(w_dff_B_MUTLEILN0_1),.clk(gclk));
	jdff dff_B_t1DlIuwm4_1(.din(w_dff_B_MUTLEILN0_1),.dout(w_dff_B_t1DlIuwm4_1),.clk(gclk));
	jdff dff_B_MDmwKUKd8_1(.din(w_dff_B_t1DlIuwm4_1),.dout(w_dff_B_MDmwKUKd8_1),.clk(gclk));
	jdff dff_B_ggdNpTeq7_1(.din(w_dff_B_MDmwKUKd8_1),.dout(w_dff_B_ggdNpTeq7_1),.clk(gclk));
	jdff dff_B_Sl6ehuhW1_1(.din(w_dff_B_ggdNpTeq7_1),.dout(w_dff_B_Sl6ehuhW1_1),.clk(gclk));
	jdff dff_B_L2g6XaFm5_1(.din(w_dff_B_Sl6ehuhW1_1),.dout(w_dff_B_L2g6XaFm5_1),.clk(gclk));
	jdff dff_B_IX9sPtvr1_1(.din(w_dff_B_L2g6XaFm5_1),.dout(w_dff_B_IX9sPtvr1_1),.clk(gclk));
	jdff dff_B_faNiQ44i5_1(.din(w_dff_B_IX9sPtvr1_1),.dout(w_dff_B_faNiQ44i5_1),.clk(gclk));
	jdff dff_B_5teCjQA89_1(.din(w_dff_B_faNiQ44i5_1),.dout(w_dff_B_5teCjQA89_1),.clk(gclk));
	jdff dff_B_pHMIlqKv2_1(.din(w_dff_B_5teCjQA89_1),.dout(w_dff_B_pHMIlqKv2_1),.clk(gclk));
	jdff dff_B_0WXk4iqa7_1(.din(w_dff_B_pHMIlqKv2_1),.dout(w_dff_B_0WXk4iqa7_1),.clk(gclk));
	jdff dff_B_BU8p5kxc3_1(.din(w_dff_B_0WXk4iqa7_1),.dout(w_dff_B_BU8p5kxc3_1),.clk(gclk));
	jdff dff_B_KwNJ0nR89_1(.din(w_dff_B_BU8p5kxc3_1),.dout(w_dff_B_KwNJ0nR89_1),.clk(gclk));
	jdff dff_B_HD1v7Uex0_1(.din(w_dff_B_KwNJ0nR89_1),.dout(w_dff_B_HD1v7Uex0_1),.clk(gclk));
	jdff dff_B_1XKQHulc3_1(.din(w_dff_B_HD1v7Uex0_1),.dout(w_dff_B_1XKQHulc3_1),.clk(gclk));
	jdff dff_B_uYRl3mGy6_1(.din(w_dff_B_1XKQHulc3_1),.dout(w_dff_B_uYRl3mGy6_1),.clk(gclk));
	jdff dff_B_O7LXoTaD2_1(.din(w_dff_B_uYRl3mGy6_1),.dout(w_dff_B_O7LXoTaD2_1),.clk(gclk));
	jdff dff_B_H1ESkHXW7_1(.din(w_dff_B_O7LXoTaD2_1),.dout(w_dff_B_H1ESkHXW7_1),.clk(gclk));
	jdff dff_B_NN6KyhtX9_1(.din(w_dff_B_H1ESkHXW7_1),.dout(w_dff_B_NN6KyhtX9_1),.clk(gclk));
	jdff dff_B_Pd2Ycupa4_1(.din(w_dff_B_NN6KyhtX9_1),.dout(w_dff_B_Pd2Ycupa4_1),.clk(gclk));
	jdff dff_B_03GxbXdr8_1(.din(w_dff_B_Pd2Ycupa4_1),.dout(w_dff_B_03GxbXdr8_1),.clk(gclk));
	jdff dff_B_MaSD429G4_1(.din(w_dff_B_03GxbXdr8_1),.dout(w_dff_B_MaSD429G4_1),.clk(gclk));
	jdff dff_B_DRNPArfw6_1(.din(w_dff_B_MaSD429G4_1),.dout(w_dff_B_DRNPArfw6_1),.clk(gclk));
	jdff dff_B_wVgaMNmO0_1(.din(w_dff_B_DRNPArfw6_1),.dout(w_dff_B_wVgaMNmO0_1),.clk(gclk));
	jdff dff_B_CNG9TtUj2_1(.din(w_dff_B_wVgaMNmO0_1),.dout(w_dff_B_CNG9TtUj2_1),.clk(gclk));
	jdff dff_B_fDJqvT1B2_1(.din(w_dff_B_CNG9TtUj2_1),.dout(w_dff_B_fDJqvT1B2_1),.clk(gclk));
	jdff dff_B_0UytVQ538_1(.din(w_dff_B_fDJqvT1B2_1),.dout(w_dff_B_0UytVQ538_1),.clk(gclk));
	jdff dff_B_1Zi6cly41_1(.din(w_dff_B_0UytVQ538_1),.dout(w_dff_B_1Zi6cly41_1),.clk(gclk));
	jdff dff_B_ZfrVhfV95_1(.din(w_dff_B_1Zi6cly41_1),.dout(w_dff_B_ZfrVhfV95_1),.clk(gclk));
	jdff dff_B_FKubNhMB5_1(.din(w_dff_B_ZfrVhfV95_1),.dout(w_dff_B_FKubNhMB5_1),.clk(gclk));
	jdff dff_B_il7oxq9A9_1(.din(w_dff_B_FKubNhMB5_1),.dout(w_dff_B_il7oxq9A9_1),.clk(gclk));
	jdff dff_B_r4gNjLID6_1(.din(w_dff_B_il7oxq9A9_1),.dout(w_dff_B_r4gNjLID6_1),.clk(gclk));
	jdff dff_B_gBvwLckV9_1(.din(w_dff_B_r4gNjLID6_1),.dout(w_dff_B_gBvwLckV9_1),.clk(gclk));
	jdff dff_B_KAgHEonp2_1(.din(w_dff_B_gBvwLckV9_1),.dout(w_dff_B_KAgHEonp2_1),.clk(gclk));
	jdff dff_B_NWOYjdxL1_1(.din(w_dff_B_KAgHEonp2_1),.dout(w_dff_B_NWOYjdxL1_1),.clk(gclk));
	jdff dff_B_w5kPSTO77_1(.din(w_dff_B_NWOYjdxL1_1),.dout(w_dff_B_w5kPSTO77_1),.clk(gclk));
	jdff dff_B_mBurp2Wg1_1(.din(w_dff_B_w5kPSTO77_1),.dout(w_dff_B_mBurp2Wg1_1),.clk(gclk));
	jdff dff_B_8ikH037v5_1(.din(w_dff_B_mBurp2Wg1_1),.dout(w_dff_B_8ikH037v5_1),.clk(gclk));
	jdff dff_B_Jc5yxD6j4_1(.din(w_dff_B_8ikH037v5_1),.dout(w_dff_B_Jc5yxD6j4_1),.clk(gclk));
	jdff dff_B_RIpNZff03_1(.din(w_dff_B_Jc5yxD6j4_1),.dout(w_dff_B_RIpNZff03_1),.clk(gclk));
	jdff dff_B_D6Qr4FjS6_1(.din(w_dff_B_RIpNZff03_1),.dout(w_dff_B_D6Qr4FjS6_1),.clk(gclk));
	jdff dff_B_hatumkC54_1(.din(w_dff_B_D6Qr4FjS6_1),.dout(w_dff_B_hatumkC54_1),.clk(gclk));
	jdff dff_B_xvc7aVNj9_1(.din(w_dff_B_hatumkC54_1),.dout(w_dff_B_xvc7aVNj9_1),.clk(gclk));
	jdff dff_B_dJmtbbsb4_1(.din(w_dff_B_xvc7aVNj9_1),.dout(w_dff_B_dJmtbbsb4_1),.clk(gclk));
	jdff dff_B_fH8U0KNH8_1(.din(w_dff_B_dJmtbbsb4_1),.dout(w_dff_B_fH8U0KNH8_1),.clk(gclk));
	jdff dff_B_DVfUTmGv6_1(.din(w_dff_B_fH8U0KNH8_1),.dout(w_dff_B_DVfUTmGv6_1),.clk(gclk));
	jdff dff_B_wkFIHAjd8_1(.din(w_dff_B_DVfUTmGv6_1),.dout(w_dff_B_wkFIHAjd8_1),.clk(gclk));
	jdff dff_B_eQUQcj2A8_1(.din(w_dff_B_wkFIHAjd8_1),.dout(w_dff_B_eQUQcj2A8_1),.clk(gclk));
	jdff dff_B_5mEazVqq0_1(.din(w_dff_B_eQUQcj2A8_1),.dout(w_dff_B_5mEazVqq0_1),.clk(gclk));
	jdff dff_B_z8quFIX49_1(.din(w_dff_B_5mEazVqq0_1),.dout(w_dff_B_z8quFIX49_1),.clk(gclk));
	jdff dff_B_5ehHha4I4_1(.din(w_dff_B_z8quFIX49_1),.dout(w_dff_B_5ehHha4I4_1),.clk(gclk));
	jdff dff_B_B7sZWNWV2_1(.din(w_dff_B_5ehHha4I4_1),.dout(w_dff_B_B7sZWNWV2_1),.clk(gclk));
	jdff dff_B_1R8BjQso5_1(.din(w_dff_B_B7sZWNWV2_1),.dout(w_dff_B_1R8BjQso5_1),.clk(gclk));
	jdff dff_B_4aMiubAG9_1(.din(w_dff_B_1R8BjQso5_1),.dout(w_dff_B_4aMiubAG9_1),.clk(gclk));
	jdff dff_B_El0fXTge8_1(.din(w_dff_B_4aMiubAG9_1),.dout(w_dff_B_El0fXTge8_1),.clk(gclk));
	jdff dff_B_RtkevHbs4_1(.din(w_dff_B_El0fXTge8_1),.dout(w_dff_B_RtkevHbs4_1),.clk(gclk));
	jdff dff_B_eagTtNFW7_1(.din(w_dff_B_RtkevHbs4_1),.dout(w_dff_B_eagTtNFW7_1),.clk(gclk));
	jdff dff_B_HnY2EmTT9_1(.din(w_dff_B_eagTtNFW7_1),.dout(w_dff_B_HnY2EmTT9_1),.clk(gclk));
	jdff dff_B_yibIVmkH0_1(.din(w_dff_B_HnY2EmTT9_1),.dout(w_dff_B_yibIVmkH0_1),.clk(gclk));
	jdff dff_B_DMfWNayZ1_1(.din(w_dff_B_yibIVmkH0_1),.dout(w_dff_B_DMfWNayZ1_1),.clk(gclk));
	jdff dff_B_AdMQCjDj7_1(.din(w_dff_B_DMfWNayZ1_1),.dout(w_dff_B_AdMQCjDj7_1),.clk(gclk));
	jdff dff_B_VE2qHRlP4_1(.din(w_dff_B_AdMQCjDj7_1),.dout(w_dff_B_VE2qHRlP4_1),.clk(gclk));
	jdff dff_B_5PgKb5Di1_1(.din(w_dff_B_VE2qHRlP4_1),.dout(w_dff_B_5PgKb5Di1_1),.clk(gclk));
	jdff dff_B_kJwU9FMJ3_1(.din(w_dff_B_5PgKb5Di1_1),.dout(w_dff_B_kJwU9FMJ3_1),.clk(gclk));
	jdff dff_B_WCDyewqD5_1(.din(w_dff_B_kJwU9FMJ3_1),.dout(w_dff_B_WCDyewqD5_1),.clk(gclk));
	jdff dff_B_Rsfv1YQS6_1(.din(w_dff_B_WCDyewqD5_1),.dout(w_dff_B_Rsfv1YQS6_1),.clk(gclk));
	jdff dff_B_20oLA5Fu7_1(.din(w_dff_B_Rsfv1YQS6_1),.dout(w_dff_B_20oLA5Fu7_1),.clk(gclk));
	jdff dff_B_NEh4Ars43_1(.din(w_dff_B_20oLA5Fu7_1),.dout(w_dff_B_NEh4Ars43_1),.clk(gclk));
	jdff dff_B_MuZtmzvI0_1(.din(w_dff_B_NEh4Ars43_1),.dout(w_dff_B_MuZtmzvI0_1),.clk(gclk));
	jdff dff_B_VqP7gHLh7_1(.din(w_dff_B_MuZtmzvI0_1),.dout(w_dff_B_VqP7gHLh7_1),.clk(gclk));
	jdff dff_B_EXarQuNl8_1(.din(w_dff_B_VqP7gHLh7_1),.dout(w_dff_B_EXarQuNl8_1),.clk(gclk));
	jdff dff_B_SYtHEa4P5_1(.din(w_dff_B_EXarQuNl8_1),.dout(w_dff_B_SYtHEa4P5_1),.clk(gclk));
	jdff dff_B_fmhA17n98_1(.din(w_dff_B_SYtHEa4P5_1),.dout(w_dff_B_fmhA17n98_1),.clk(gclk));
	jdff dff_B_yhtsF8Sz7_1(.din(w_dff_B_fmhA17n98_1),.dout(w_dff_B_yhtsF8Sz7_1),.clk(gclk));
	jdff dff_B_Cn2hHtih0_1(.din(w_dff_B_yhtsF8Sz7_1),.dout(w_dff_B_Cn2hHtih0_1),.clk(gclk));
	jdff dff_B_8xIVSn6b0_1(.din(w_dff_B_Cn2hHtih0_1),.dout(w_dff_B_8xIVSn6b0_1),.clk(gclk));
	jdff dff_B_toIxr72N6_1(.din(w_dff_B_8xIVSn6b0_1),.dout(w_dff_B_toIxr72N6_1),.clk(gclk));
	jdff dff_B_BFLvQCNi1_1(.din(w_dff_B_toIxr72N6_1),.dout(w_dff_B_BFLvQCNi1_1),.clk(gclk));
	jdff dff_B_zlMrmKcm4_1(.din(w_dff_B_BFLvQCNi1_1),.dout(w_dff_B_zlMrmKcm4_1),.clk(gclk));
	jdff dff_B_cO5bJQqp0_1(.din(w_dff_B_zlMrmKcm4_1),.dout(w_dff_B_cO5bJQqp0_1),.clk(gclk));
	jdff dff_B_phmxwEJS6_1(.din(w_dff_B_cO5bJQqp0_1),.dout(w_dff_B_phmxwEJS6_1),.clk(gclk));
	jdff dff_B_cCTExRmf2_1(.din(w_dff_B_phmxwEJS6_1),.dout(w_dff_B_cCTExRmf2_1),.clk(gclk));
	jdff dff_B_epsTtTK93_1(.din(w_dff_B_cCTExRmf2_1),.dout(w_dff_B_epsTtTK93_1),.clk(gclk));
	jdff dff_B_lJKhvoH82_0(.din(n901),.dout(w_dff_B_lJKhvoH82_0),.clk(gclk));
	jdff dff_B_tYJqsr5I9_0(.din(w_dff_B_lJKhvoH82_0),.dout(w_dff_B_tYJqsr5I9_0),.clk(gclk));
	jdff dff_B_Z3Z7ZH8q4_0(.din(w_dff_B_tYJqsr5I9_0),.dout(w_dff_B_Z3Z7ZH8q4_0),.clk(gclk));
	jdff dff_B_RGMB55Qg6_0(.din(w_dff_B_Z3Z7ZH8q4_0),.dout(w_dff_B_RGMB55Qg6_0),.clk(gclk));
	jdff dff_B_DpLshpnH9_0(.din(w_dff_B_RGMB55Qg6_0),.dout(w_dff_B_DpLshpnH9_0),.clk(gclk));
	jdff dff_B_UT2eOLfP0_0(.din(w_dff_B_DpLshpnH9_0),.dout(w_dff_B_UT2eOLfP0_0),.clk(gclk));
	jdff dff_B_rhzop9Wj6_0(.din(w_dff_B_UT2eOLfP0_0),.dout(w_dff_B_rhzop9Wj6_0),.clk(gclk));
	jdff dff_B_8Lx8gHrN0_0(.din(w_dff_B_rhzop9Wj6_0),.dout(w_dff_B_8Lx8gHrN0_0),.clk(gclk));
	jdff dff_B_3cAwkOm45_0(.din(w_dff_B_8Lx8gHrN0_0),.dout(w_dff_B_3cAwkOm45_0),.clk(gclk));
	jdff dff_B_HNHTCCXO0_0(.din(w_dff_B_3cAwkOm45_0),.dout(w_dff_B_HNHTCCXO0_0),.clk(gclk));
	jdff dff_B_F8LxUllA6_0(.din(w_dff_B_HNHTCCXO0_0),.dout(w_dff_B_F8LxUllA6_0),.clk(gclk));
	jdff dff_B_rX82UoT69_0(.din(w_dff_B_F8LxUllA6_0),.dout(w_dff_B_rX82UoT69_0),.clk(gclk));
	jdff dff_B_Ak7edaud8_0(.din(w_dff_B_rX82UoT69_0),.dout(w_dff_B_Ak7edaud8_0),.clk(gclk));
	jdff dff_B_RCebTlL39_0(.din(w_dff_B_Ak7edaud8_0),.dout(w_dff_B_RCebTlL39_0),.clk(gclk));
	jdff dff_B_59V0tLYw0_0(.din(w_dff_B_RCebTlL39_0),.dout(w_dff_B_59V0tLYw0_0),.clk(gclk));
	jdff dff_B_D3UdOmYb1_0(.din(w_dff_B_59V0tLYw0_0),.dout(w_dff_B_D3UdOmYb1_0),.clk(gclk));
	jdff dff_B_xxoqTyml6_0(.din(w_dff_B_D3UdOmYb1_0),.dout(w_dff_B_xxoqTyml6_0),.clk(gclk));
	jdff dff_B_BMkInMR34_0(.din(w_dff_B_xxoqTyml6_0),.dout(w_dff_B_BMkInMR34_0),.clk(gclk));
	jdff dff_B_xc42WZ2K7_0(.din(w_dff_B_BMkInMR34_0),.dout(w_dff_B_xc42WZ2K7_0),.clk(gclk));
	jdff dff_B_3u70UCbM7_0(.din(w_dff_B_xc42WZ2K7_0),.dout(w_dff_B_3u70UCbM7_0),.clk(gclk));
	jdff dff_B_qcnVjCEA7_0(.din(w_dff_B_3u70UCbM7_0),.dout(w_dff_B_qcnVjCEA7_0),.clk(gclk));
	jdff dff_B_3t1jWBqX8_0(.din(w_dff_B_qcnVjCEA7_0),.dout(w_dff_B_3t1jWBqX8_0),.clk(gclk));
	jdff dff_B_3sEaB4hb2_0(.din(w_dff_B_3t1jWBqX8_0),.dout(w_dff_B_3sEaB4hb2_0),.clk(gclk));
	jdff dff_B_bOJPNF9p3_0(.din(w_dff_B_3sEaB4hb2_0),.dout(w_dff_B_bOJPNF9p3_0),.clk(gclk));
	jdff dff_B_LSbV7o3T6_0(.din(w_dff_B_bOJPNF9p3_0),.dout(w_dff_B_LSbV7o3T6_0),.clk(gclk));
	jdff dff_B_0gVHR0mp2_0(.din(w_dff_B_LSbV7o3T6_0),.dout(w_dff_B_0gVHR0mp2_0),.clk(gclk));
	jdff dff_B_CcVqdpX83_0(.din(w_dff_B_0gVHR0mp2_0),.dout(w_dff_B_CcVqdpX83_0),.clk(gclk));
	jdff dff_B_HhYHRB5A6_0(.din(w_dff_B_CcVqdpX83_0),.dout(w_dff_B_HhYHRB5A6_0),.clk(gclk));
	jdff dff_B_xdK0AGMy6_0(.din(w_dff_B_HhYHRB5A6_0),.dout(w_dff_B_xdK0AGMy6_0),.clk(gclk));
	jdff dff_B_mNqA4OR71_0(.din(w_dff_B_xdK0AGMy6_0),.dout(w_dff_B_mNqA4OR71_0),.clk(gclk));
	jdff dff_B_DuajkWtH8_0(.din(w_dff_B_mNqA4OR71_0),.dout(w_dff_B_DuajkWtH8_0),.clk(gclk));
	jdff dff_B_yiRRm0pg0_0(.din(w_dff_B_DuajkWtH8_0),.dout(w_dff_B_yiRRm0pg0_0),.clk(gclk));
	jdff dff_B_dquNXKj92_0(.din(w_dff_B_yiRRm0pg0_0),.dout(w_dff_B_dquNXKj92_0),.clk(gclk));
	jdff dff_B_MY61xwSR8_0(.din(w_dff_B_dquNXKj92_0),.dout(w_dff_B_MY61xwSR8_0),.clk(gclk));
	jdff dff_B_OqlVEJAF1_0(.din(w_dff_B_MY61xwSR8_0),.dout(w_dff_B_OqlVEJAF1_0),.clk(gclk));
	jdff dff_B_Z3LdAn8U1_0(.din(w_dff_B_OqlVEJAF1_0),.dout(w_dff_B_Z3LdAn8U1_0),.clk(gclk));
	jdff dff_B_4WiDP0Jz6_0(.din(w_dff_B_Z3LdAn8U1_0),.dout(w_dff_B_4WiDP0Jz6_0),.clk(gclk));
	jdff dff_B_zNVdezlO2_0(.din(w_dff_B_4WiDP0Jz6_0),.dout(w_dff_B_zNVdezlO2_0),.clk(gclk));
	jdff dff_B_6G5koO6k8_0(.din(w_dff_B_zNVdezlO2_0),.dout(w_dff_B_6G5koO6k8_0),.clk(gclk));
	jdff dff_B_qnyw3YUh8_0(.din(w_dff_B_6G5koO6k8_0),.dout(w_dff_B_qnyw3YUh8_0),.clk(gclk));
	jdff dff_B_hVQt8W721_0(.din(w_dff_B_qnyw3YUh8_0),.dout(w_dff_B_hVQt8W721_0),.clk(gclk));
	jdff dff_B_h6j9IioH2_0(.din(w_dff_B_hVQt8W721_0),.dout(w_dff_B_h6j9IioH2_0),.clk(gclk));
	jdff dff_B_qpQOSbSI1_0(.din(w_dff_B_h6j9IioH2_0),.dout(w_dff_B_qpQOSbSI1_0),.clk(gclk));
	jdff dff_B_dtO7tGe90_0(.din(w_dff_B_qpQOSbSI1_0),.dout(w_dff_B_dtO7tGe90_0),.clk(gclk));
	jdff dff_B_XtxS4THl4_0(.din(w_dff_B_dtO7tGe90_0),.dout(w_dff_B_XtxS4THl4_0),.clk(gclk));
	jdff dff_B_LyroC0pO7_0(.din(w_dff_B_XtxS4THl4_0),.dout(w_dff_B_LyroC0pO7_0),.clk(gclk));
	jdff dff_B_se7GK7f21_0(.din(w_dff_B_LyroC0pO7_0),.dout(w_dff_B_se7GK7f21_0),.clk(gclk));
	jdff dff_B_DlLxr2Yu4_0(.din(w_dff_B_se7GK7f21_0),.dout(w_dff_B_DlLxr2Yu4_0),.clk(gclk));
	jdff dff_B_HD8vbn4S1_0(.din(w_dff_B_DlLxr2Yu4_0),.dout(w_dff_B_HD8vbn4S1_0),.clk(gclk));
	jdff dff_B_oDuOkmWK7_0(.din(w_dff_B_HD8vbn4S1_0),.dout(w_dff_B_oDuOkmWK7_0),.clk(gclk));
	jdff dff_B_9TE1E8X39_0(.din(w_dff_B_oDuOkmWK7_0),.dout(w_dff_B_9TE1E8X39_0),.clk(gclk));
	jdff dff_B_noti4kox8_0(.din(w_dff_B_9TE1E8X39_0),.dout(w_dff_B_noti4kox8_0),.clk(gclk));
	jdff dff_B_tdplmZdU6_0(.din(w_dff_B_noti4kox8_0),.dout(w_dff_B_tdplmZdU6_0),.clk(gclk));
	jdff dff_B_7EeOCSTE5_0(.din(w_dff_B_tdplmZdU6_0),.dout(w_dff_B_7EeOCSTE5_0),.clk(gclk));
	jdff dff_B_BzLW0QeY4_0(.din(w_dff_B_7EeOCSTE5_0),.dout(w_dff_B_BzLW0QeY4_0),.clk(gclk));
	jdff dff_B_TfodfJ7I6_0(.din(w_dff_B_BzLW0QeY4_0),.dout(w_dff_B_TfodfJ7I6_0),.clk(gclk));
	jdff dff_B_TeAOA5997_0(.din(w_dff_B_TfodfJ7I6_0),.dout(w_dff_B_TeAOA5997_0),.clk(gclk));
	jdff dff_B_O2GFG1zm8_0(.din(w_dff_B_TeAOA5997_0),.dout(w_dff_B_O2GFG1zm8_0),.clk(gclk));
	jdff dff_B_mFtGdxyv1_0(.din(w_dff_B_O2GFG1zm8_0),.dout(w_dff_B_mFtGdxyv1_0),.clk(gclk));
	jdff dff_B_wuYptM569_0(.din(w_dff_B_mFtGdxyv1_0),.dout(w_dff_B_wuYptM569_0),.clk(gclk));
	jdff dff_B_sIjMrqwr4_0(.din(w_dff_B_wuYptM569_0),.dout(w_dff_B_sIjMrqwr4_0),.clk(gclk));
	jdff dff_B_2PfwSk4k2_0(.din(w_dff_B_sIjMrqwr4_0),.dout(w_dff_B_2PfwSk4k2_0),.clk(gclk));
	jdff dff_B_Lgz7XXpd8_0(.din(w_dff_B_2PfwSk4k2_0),.dout(w_dff_B_Lgz7XXpd8_0),.clk(gclk));
	jdff dff_B_mvmbzmkD9_0(.din(w_dff_B_Lgz7XXpd8_0),.dout(w_dff_B_mvmbzmkD9_0),.clk(gclk));
	jdff dff_B_RMiPg7n25_0(.din(w_dff_B_mvmbzmkD9_0),.dout(w_dff_B_RMiPg7n25_0),.clk(gclk));
	jdff dff_B_hE5szb6K7_0(.din(w_dff_B_RMiPg7n25_0),.dout(w_dff_B_hE5szb6K7_0),.clk(gclk));
	jdff dff_B_Qvfx0zTR0_0(.din(w_dff_B_hE5szb6K7_0),.dout(w_dff_B_Qvfx0zTR0_0),.clk(gclk));
	jdff dff_B_3ElEBm7Y3_0(.din(w_dff_B_Qvfx0zTR0_0),.dout(w_dff_B_3ElEBm7Y3_0),.clk(gclk));
	jdff dff_B_sSJRl0zJ3_0(.din(w_dff_B_3ElEBm7Y3_0),.dout(w_dff_B_sSJRl0zJ3_0),.clk(gclk));
	jdff dff_B_nkWTR3151_0(.din(w_dff_B_sSJRl0zJ3_0),.dout(w_dff_B_nkWTR3151_0),.clk(gclk));
	jdff dff_B_9XRJmcUB6_0(.din(w_dff_B_nkWTR3151_0),.dout(w_dff_B_9XRJmcUB6_0),.clk(gclk));
	jdff dff_B_J2wQ01T72_0(.din(w_dff_B_9XRJmcUB6_0),.dout(w_dff_B_J2wQ01T72_0),.clk(gclk));
	jdff dff_B_weR9CNAu3_0(.din(w_dff_B_J2wQ01T72_0),.dout(w_dff_B_weR9CNAu3_0),.clk(gclk));
	jdff dff_B_81W8Bcd78_0(.din(w_dff_B_weR9CNAu3_0),.dout(w_dff_B_81W8Bcd78_0),.clk(gclk));
	jdff dff_B_WEX9TPsK2_0(.din(w_dff_B_81W8Bcd78_0),.dout(w_dff_B_WEX9TPsK2_0),.clk(gclk));
	jdff dff_B_CxjRKDCx8_0(.din(w_dff_B_WEX9TPsK2_0),.dout(w_dff_B_CxjRKDCx8_0),.clk(gclk));
	jdff dff_B_sKnetmQq7_0(.din(w_dff_B_CxjRKDCx8_0),.dout(w_dff_B_sKnetmQq7_0),.clk(gclk));
	jdff dff_B_oA16ioMu6_0(.din(w_dff_B_sKnetmQq7_0),.dout(w_dff_B_oA16ioMu6_0),.clk(gclk));
	jdff dff_B_TLmonIpi5_0(.din(w_dff_B_oA16ioMu6_0),.dout(w_dff_B_TLmonIpi5_0),.clk(gclk));
	jdff dff_B_HqjuU3ck9_0(.din(w_dff_B_TLmonIpi5_0),.dout(w_dff_B_HqjuU3ck9_0),.clk(gclk));
	jdff dff_B_jG98F9on0_0(.din(w_dff_B_HqjuU3ck9_0),.dout(w_dff_B_jG98F9on0_0),.clk(gclk));
	jdff dff_B_GwOesIIM8_0(.din(w_dff_B_jG98F9on0_0),.dout(w_dff_B_GwOesIIM8_0),.clk(gclk));
	jdff dff_B_ni1zVnKN5_0(.din(w_dff_B_GwOesIIM8_0),.dout(w_dff_B_ni1zVnKN5_0),.clk(gclk));
	jdff dff_B_xJLu7Dhv0_0(.din(w_dff_B_ni1zVnKN5_0),.dout(w_dff_B_xJLu7Dhv0_0),.clk(gclk));
	jdff dff_B_BTdgaiJE3_0(.din(w_dff_B_xJLu7Dhv0_0),.dout(w_dff_B_BTdgaiJE3_0),.clk(gclk));
	jdff dff_B_f56FFK1t6_0(.din(w_dff_B_BTdgaiJE3_0),.dout(w_dff_B_f56FFK1t6_0),.clk(gclk));
	jdff dff_B_zbQvJ6C20_1(.din(n894),.dout(w_dff_B_zbQvJ6C20_1),.clk(gclk));
	jdff dff_B_qkZKEyZM5_1(.din(w_dff_B_zbQvJ6C20_1),.dout(w_dff_B_qkZKEyZM5_1),.clk(gclk));
	jdff dff_B_j4xkmDK01_1(.din(w_dff_B_qkZKEyZM5_1),.dout(w_dff_B_j4xkmDK01_1),.clk(gclk));
	jdff dff_B_zatxTxgJ2_1(.din(w_dff_B_j4xkmDK01_1),.dout(w_dff_B_zatxTxgJ2_1),.clk(gclk));
	jdff dff_B_z23GvKJy1_1(.din(w_dff_B_zatxTxgJ2_1),.dout(w_dff_B_z23GvKJy1_1),.clk(gclk));
	jdff dff_B_FU5uW0LL5_1(.din(w_dff_B_z23GvKJy1_1),.dout(w_dff_B_FU5uW0LL5_1),.clk(gclk));
	jdff dff_B_0JOslABT7_1(.din(w_dff_B_FU5uW0LL5_1),.dout(w_dff_B_0JOslABT7_1),.clk(gclk));
	jdff dff_B_zfaeMbhO7_1(.din(w_dff_B_0JOslABT7_1),.dout(w_dff_B_zfaeMbhO7_1),.clk(gclk));
	jdff dff_B_By6RENUn8_1(.din(w_dff_B_zfaeMbhO7_1),.dout(w_dff_B_By6RENUn8_1),.clk(gclk));
	jdff dff_B_Cm0JmzQM0_1(.din(w_dff_B_By6RENUn8_1),.dout(w_dff_B_Cm0JmzQM0_1),.clk(gclk));
	jdff dff_B_MRWRJWiv5_1(.din(w_dff_B_Cm0JmzQM0_1),.dout(w_dff_B_MRWRJWiv5_1),.clk(gclk));
	jdff dff_B_bKcHDVgq7_1(.din(w_dff_B_MRWRJWiv5_1),.dout(w_dff_B_bKcHDVgq7_1),.clk(gclk));
	jdff dff_B_agEp6D0J7_1(.din(w_dff_B_bKcHDVgq7_1),.dout(w_dff_B_agEp6D0J7_1),.clk(gclk));
	jdff dff_B_yXzGxSnQ9_1(.din(w_dff_B_agEp6D0J7_1),.dout(w_dff_B_yXzGxSnQ9_1),.clk(gclk));
	jdff dff_B_27yZqm3R3_1(.din(w_dff_B_yXzGxSnQ9_1),.dout(w_dff_B_27yZqm3R3_1),.clk(gclk));
	jdff dff_B_jOX0Y95X4_1(.din(w_dff_B_27yZqm3R3_1),.dout(w_dff_B_jOX0Y95X4_1),.clk(gclk));
	jdff dff_B_JG3sCRf83_1(.din(w_dff_B_jOX0Y95X4_1),.dout(w_dff_B_JG3sCRf83_1),.clk(gclk));
	jdff dff_B_ofZCAthg4_1(.din(w_dff_B_JG3sCRf83_1),.dout(w_dff_B_ofZCAthg4_1),.clk(gclk));
	jdff dff_B_Wlj5ZjIk6_1(.din(w_dff_B_ofZCAthg4_1),.dout(w_dff_B_Wlj5ZjIk6_1),.clk(gclk));
	jdff dff_B_Ct3kltv05_1(.din(w_dff_B_Wlj5ZjIk6_1),.dout(w_dff_B_Ct3kltv05_1),.clk(gclk));
	jdff dff_B_lp7XH4td4_1(.din(w_dff_B_Ct3kltv05_1),.dout(w_dff_B_lp7XH4td4_1),.clk(gclk));
	jdff dff_B_t8nnAsFa4_1(.din(w_dff_B_lp7XH4td4_1),.dout(w_dff_B_t8nnAsFa4_1),.clk(gclk));
	jdff dff_B_iIHAmn9P9_1(.din(w_dff_B_t8nnAsFa4_1),.dout(w_dff_B_iIHAmn9P9_1),.clk(gclk));
	jdff dff_B_9QUtU3ri9_1(.din(w_dff_B_iIHAmn9P9_1),.dout(w_dff_B_9QUtU3ri9_1),.clk(gclk));
	jdff dff_B_JJZDMfo27_1(.din(w_dff_B_9QUtU3ri9_1),.dout(w_dff_B_JJZDMfo27_1),.clk(gclk));
	jdff dff_B_hdB5Vu0Y0_1(.din(w_dff_B_JJZDMfo27_1),.dout(w_dff_B_hdB5Vu0Y0_1),.clk(gclk));
	jdff dff_B_GCPQZIcq3_1(.din(w_dff_B_hdB5Vu0Y0_1),.dout(w_dff_B_GCPQZIcq3_1),.clk(gclk));
	jdff dff_B_aLlYiWik5_1(.din(w_dff_B_GCPQZIcq3_1),.dout(w_dff_B_aLlYiWik5_1),.clk(gclk));
	jdff dff_B_grzNRwks5_1(.din(w_dff_B_aLlYiWik5_1),.dout(w_dff_B_grzNRwks5_1),.clk(gclk));
	jdff dff_B_XYADlfYb7_1(.din(w_dff_B_grzNRwks5_1),.dout(w_dff_B_XYADlfYb7_1),.clk(gclk));
	jdff dff_B_MiP3P8gZ6_1(.din(w_dff_B_XYADlfYb7_1),.dout(w_dff_B_MiP3P8gZ6_1),.clk(gclk));
	jdff dff_B_L2NoJ0596_1(.din(w_dff_B_MiP3P8gZ6_1),.dout(w_dff_B_L2NoJ0596_1),.clk(gclk));
	jdff dff_B_8RkYEkTS8_1(.din(w_dff_B_L2NoJ0596_1),.dout(w_dff_B_8RkYEkTS8_1),.clk(gclk));
	jdff dff_B_k2IuLtRU2_1(.din(w_dff_B_8RkYEkTS8_1),.dout(w_dff_B_k2IuLtRU2_1),.clk(gclk));
	jdff dff_B_05SpV9JD0_1(.din(w_dff_B_k2IuLtRU2_1),.dout(w_dff_B_05SpV9JD0_1),.clk(gclk));
	jdff dff_B_vRPA8CpO5_1(.din(w_dff_B_05SpV9JD0_1),.dout(w_dff_B_vRPA8CpO5_1),.clk(gclk));
	jdff dff_B_Iss29SFq5_1(.din(w_dff_B_vRPA8CpO5_1),.dout(w_dff_B_Iss29SFq5_1),.clk(gclk));
	jdff dff_B_MkWsVnk81_1(.din(w_dff_B_Iss29SFq5_1),.dout(w_dff_B_MkWsVnk81_1),.clk(gclk));
	jdff dff_B_SnWspLte0_1(.din(w_dff_B_MkWsVnk81_1),.dout(w_dff_B_SnWspLte0_1),.clk(gclk));
	jdff dff_B_v7h1jybE7_1(.din(w_dff_B_SnWspLte0_1),.dout(w_dff_B_v7h1jybE7_1),.clk(gclk));
	jdff dff_B_tWfbd1wB9_1(.din(w_dff_B_v7h1jybE7_1),.dout(w_dff_B_tWfbd1wB9_1),.clk(gclk));
	jdff dff_B_uiYCYSo46_1(.din(w_dff_B_tWfbd1wB9_1),.dout(w_dff_B_uiYCYSo46_1),.clk(gclk));
	jdff dff_B_hef6HTNh4_1(.din(w_dff_B_uiYCYSo46_1),.dout(w_dff_B_hef6HTNh4_1),.clk(gclk));
	jdff dff_B_KsnqZkag3_1(.din(w_dff_B_hef6HTNh4_1),.dout(w_dff_B_KsnqZkag3_1),.clk(gclk));
	jdff dff_B_zoYKeZuQ2_1(.din(w_dff_B_KsnqZkag3_1),.dout(w_dff_B_zoYKeZuQ2_1),.clk(gclk));
	jdff dff_B_lqUlsJr93_1(.din(w_dff_B_zoYKeZuQ2_1),.dout(w_dff_B_lqUlsJr93_1),.clk(gclk));
	jdff dff_B_2qg6iKSM7_1(.din(w_dff_B_lqUlsJr93_1),.dout(w_dff_B_2qg6iKSM7_1),.clk(gclk));
	jdff dff_B_caYLUQbm4_1(.din(w_dff_B_2qg6iKSM7_1),.dout(w_dff_B_caYLUQbm4_1),.clk(gclk));
	jdff dff_B_0rqwwXhM5_1(.din(w_dff_B_caYLUQbm4_1),.dout(w_dff_B_0rqwwXhM5_1),.clk(gclk));
	jdff dff_B_xfgpOJRk4_1(.din(w_dff_B_0rqwwXhM5_1),.dout(w_dff_B_xfgpOJRk4_1),.clk(gclk));
	jdff dff_B_QrJq7BVy9_1(.din(w_dff_B_xfgpOJRk4_1),.dout(w_dff_B_QrJq7BVy9_1),.clk(gclk));
	jdff dff_B_r62YTe5a1_1(.din(w_dff_B_QrJq7BVy9_1),.dout(w_dff_B_r62YTe5a1_1),.clk(gclk));
	jdff dff_B_wXIeoSUK9_1(.din(w_dff_B_r62YTe5a1_1),.dout(w_dff_B_wXIeoSUK9_1),.clk(gclk));
	jdff dff_B_FtB8rJSI9_1(.din(w_dff_B_wXIeoSUK9_1),.dout(w_dff_B_FtB8rJSI9_1),.clk(gclk));
	jdff dff_B_889gqyHm2_1(.din(w_dff_B_FtB8rJSI9_1),.dout(w_dff_B_889gqyHm2_1),.clk(gclk));
	jdff dff_B_yRAVixMX4_1(.din(w_dff_B_889gqyHm2_1),.dout(w_dff_B_yRAVixMX4_1),.clk(gclk));
	jdff dff_B_Kv6Gql8K6_1(.din(w_dff_B_yRAVixMX4_1),.dout(w_dff_B_Kv6Gql8K6_1),.clk(gclk));
	jdff dff_B_9ongw8eY6_1(.din(w_dff_B_Kv6Gql8K6_1),.dout(w_dff_B_9ongw8eY6_1),.clk(gclk));
	jdff dff_B_VFdd7dNM6_1(.din(w_dff_B_9ongw8eY6_1),.dout(w_dff_B_VFdd7dNM6_1),.clk(gclk));
	jdff dff_B_johDkqTX1_1(.din(w_dff_B_VFdd7dNM6_1),.dout(w_dff_B_johDkqTX1_1),.clk(gclk));
	jdff dff_B_xG0IAOyf5_1(.din(w_dff_B_johDkqTX1_1),.dout(w_dff_B_xG0IAOyf5_1),.clk(gclk));
	jdff dff_B_ontINZd45_1(.din(w_dff_B_xG0IAOyf5_1),.dout(w_dff_B_ontINZd45_1),.clk(gclk));
	jdff dff_B_mponBiiv1_1(.din(w_dff_B_ontINZd45_1),.dout(w_dff_B_mponBiiv1_1),.clk(gclk));
	jdff dff_B_7oyNpD7Y9_1(.din(w_dff_B_mponBiiv1_1),.dout(w_dff_B_7oyNpD7Y9_1),.clk(gclk));
	jdff dff_B_MHFPgTmc5_1(.din(w_dff_B_7oyNpD7Y9_1),.dout(w_dff_B_MHFPgTmc5_1),.clk(gclk));
	jdff dff_B_Un8VFwHd3_1(.din(w_dff_B_MHFPgTmc5_1),.dout(w_dff_B_Un8VFwHd3_1),.clk(gclk));
	jdff dff_B_AZY4aIGL8_1(.din(w_dff_B_Un8VFwHd3_1),.dout(w_dff_B_AZY4aIGL8_1),.clk(gclk));
	jdff dff_B_hWbl4can7_1(.din(w_dff_B_AZY4aIGL8_1),.dout(w_dff_B_hWbl4can7_1),.clk(gclk));
	jdff dff_B_zTtvZ0Ge9_1(.din(w_dff_B_hWbl4can7_1),.dout(w_dff_B_zTtvZ0Ge9_1),.clk(gclk));
	jdff dff_B_HgqGc6jD2_1(.din(w_dff_B_zTtvZ0Ge9_1),.dout(w_dff_B_HgqGc6jD2_1),.clk(gclk));
	jdff dff_B_kbJGJARV1_1(.din(w_dff_B_HgqGc6jD2_1),.dout(w_dff_B_kbJGJARV1_1),.clk(gclk));
	jdff dff_B_3TvpvZzv1_1(.din(w_dff_B_kbJGJARV1_1),.dout(w_dff_B_3TvpvZzv1_1),.clk(gclk));
	jdff dff_B_q0e6NACN2_1(.din(w_dff_B_3TvpvZzv1_1),.dout(w_dff_B_q0e6NACN2_1),.clk(gclk));
	jdff dff_B_Pb5dlJDf5_1(.din(w_dff_B_q0e6NACN2_1),.dout(w_dff_B_Pb5dlJDf5_1),.clk(gclk));
	jdff dff_B_rZYql6Ih7_1(.din(w_dff_B_Pb5dlJDf5_1),.dout(w_dff_B_rZYql6Ih7_1),.clk(gclk));
	jdff dff_B_RPzSUgBZ5_1(.din(w_dff_B_rZYql6Ih7_1),.dout(w_dff_B_RPzSUgBZ5_1),.clk(gclk));
	jdff dff_B_ugtsLmQ65_1(.din(w_dff_B_RPzSUgBZ5_1),.dout(w_dff_B_ugtsLmQ65_1),.clk(gclk));
	jdff dff_B_U3ER6DbH1_1(.din(w_dff_B_ugtsLmQ65_1),.dout(w_dff_B_U3ER6DbH1_1),.clk(gclk));
	jdff dff_B_BMdQNpqJ9_1(.din(w_dff_B_U3ER6DbH1_1),.dout(w_dff_B_BMdQNpqJ9_1),.clk(gclk));
	jdff dff_B_BClkdMQc4_1(.din(w_dff_B_BMdQNpqJ9_1),.dout(w_dff_B_BClkdMQc4_1),.clk(gclk));
	jdff dff_B_gBg1UEpp0_1(.din(w_dff_B_BClkdMQc4_1),.dout(w_dff_B_gBg1UEpp0_1),.clk(gclk));
	jdff dff_B_qFVlKnSy1_1(.din(w_dff_B_gBg1UEpp0_1),.dout(w_dff_B_qFVlKnSy1_1),.clk(gclk));
	jdff dff_B_TBbi45624_1(.din(w_dff_B_qFVlKnSy1_1),.dout(w_dff_B_TBbi45624_1),.clk(gclk));
	jdff dff_B_nZFY3ZaV0_1(.din(w_dff_B_TBbi45624_1),.dout(w_dff_B_nZFY3ZaV0_1),.clk(gclk));
	jdff dff_B_8UlPWcMp1_1(.din(w_dff_B_nZFY3ZaV0_1),.dout(w_dff_B_8UlPWcMp1_1),.clk(gclk));
	jdff dff_B_3msDc8HK9_0(.din(n895),.dout(w_dff_B_3msDc8HK9_0),.clk(gclk));
	jdff dff_B_dmrV2Ji61_0(.din(w_dff_B_3msDc8HK9_0),.dout(w_dff_B_dmrV2Ji61_0),.clk(gclk));
	jdff dff_B_FdG9gOQB6_0(.din(w_dff_B_dmrV2Ji61_0),.dout(w_dff_B_FdG9gOQB6_0),.clk(gclk));
	jdff dff_B_0n35iexP7_0(.din(w_dff_B_FdG9gOQB6_0),.dout(w_dff_B_0n35iexP7_0),.clk(gclk));
	jdff dff_B_QWhhxulS7_0(.din(w_dff_B_0n35iexP7_0),.dout(w_dff_B_QWhhxulS7_0),.clk(gclk));
	jdff dff_B_EVumF80J0_0(.din(w_dff_B_QWhhxulS7_0),.dout(w_dff_B_EVumF80J0_0),.clk(gclk));
	jdff dff_B_PTML7Nqq4_0(.din(w_dff_B_EVumF80J0_0),.dout(w_dff_B_PTML7Nqq4_0),.clk(gclk));
	jdff dff_B_4esAWS705_0(.din(w_dff_B_PTML7Nqq4_0),.dout(w_dff_B_4esAWS705_0),.clk(gclk));
	jdff dff_B_lMgLuAUV7_0(.din(w_dff_B_4esAWS705_0),.dout(w_dff_B_lMgLuAUV7_0),.clk(gclk));
	jdff dff_B_UVXGxXoK5_0(.din(w_dff_B_lMgLuAUV7_0),.dout(w_dff_B_UVXGxXoK5_0),.clk(gclk));
	jdff dff_B_iBUuvlbL8_0(.din(w_dff_B_UVXGxXoK5_0),.dout(w_dff_B_iBUuvlbL8_0),.clk(gclk));
	jdff dff_B_g7anM3Pd5_0(.din(w_dff_B_iBUuvlbL8_0),.dout(w_dff_B_g7anM3Pd5_0),.clk(gclk));
	jdff dff_B_MFxd858v7_0(.din(w_dff_B_g7anM3Pd5_0),.dout(w_dff_B_MFxd858v7_0),.clk(gclk));
	jdff dff_B_k18YaPRN6_0(.din(w_dff_B_MFxd858v7_0),.dout(w_dff_B_k18YaPRN6_0),.clk(gclk));
	jdff dff_B_yFmWwlCQ8_0(.din(w_dff_B_k18YaPRN6_0),.dout(w_dff_B_yFmWwlCQ8_0),.clk(gclk));
	jdff dff_B_aRYMJqhW1_0(.din(w_dff_B_yFmWwlCQ8_0),.dout(w_dff_B_aRYMJqhW1_0),.clk(gclk));
	jdff dff_B_VZTQcXus1_0(.din(w_dff_B_aRYMJqhW1_0),.dout(w_dff_B_VZTQcXus1_0),.clk(gclk));
	jdff dff_B_QdAZzkMb6_0(.din(w_dff_B_VZTQcXus1_0),.dout(w_dff_B_QdAZzkMb6_0),.clk(gclk));
	jdff dff_B_SoPw7wRM5_0(.din(w_dff_B_QdAZzkMb6_0),.dout(w_dff_B_SoPw7wRM5_0),.clk(gclk));
	jdff dff_B_5BTjZDLb8_0(.din(w_dff_B_SoPw7wRM5_0),.dout(w_dff_B_5BTjZDLb8_0),.clk(gclk));
	jdff dff_B_FHSyB3Yj9_0(.din(w_dff_B_5BTjZDLb8_0),.dout(w_dff_B_FHSyB3Yj9_0),.clk(gclk));
	jdff dff_B_aX53TefW5_0(.din(w_dff_B_FHSyB3Yj9_0),.dout(w_dff_B_aX53TefW5_0),.clk(gclk));
	jdff dff_B_QIUiqdd55_0(.din(w_dff_B_aX53TefW5_0),.dout(w_dff_B_QIUiqdd55_0),.clk(gclk));
	jdff dff_B_qLMAomy10_0(.din(w_dff_B_QIUiqdd55_0),.dout(w_dff_B_qLMAomy10_0),.clk(gclk));
	jdff dff_B_dzJuL4r81_0(.din(w_dff_B_qLMAomy10_0),.dout(w_dff_B_dzJuL4r81_0),.clk(gclk));
	jdff dff_B_qExanZTJ3_0(.din(w_dff_B_dzJuL4r81_0),.dout(w_dff_B_qExanZTJ3_0),.clk(gclk));
	jdff dff_B_DMVlJJIf6_0(.din(w_dff_B_qExanZTJ3_0),.dout(w_dff_B_DMVlJJIf6_0),.clk(gclk));
	jdff dff_B_b6kgwMDK7_0(.din(w_dff_B_DMVlJJIf6_0),.dout(w_dff_B_b6kgwMDK7_0),.clk(gclk));
	jdff dff_B_BC2WxAwk3_0(.din(w_dff_B_b6kgwMDK7_0),.dout(w_dff_B_BC2WxAwk3_0),.clk(gclk));
	jdff dff_B_z3GeC4HW3_0(.din(w_dff_B_BC2WxAwk3_0),.dout(w_dff_B_z3GeC4HW3_0),.clk(gclk));
	jdff dff_B_ihpTs5eF0_0(.din(w_dff_B_z3GeC4HW3_0),.dout(w_dff_B_ihpTs5eF0_0),.clk(gclk));
	jdff dff_B_sETUEPwu2_0(.din(w_dff_B_ihpTs5eF0_0),.dout(w_dff_B_sETUEPwu2_0),.clk(gclk));
	jdff dff_B_4U1pC6Ie1_0(.din(w_dff_B_sETUEPwu2_0),.dout(w_dff_B_4U1pC6Ie1_0),.clk(gclk));
	jdff dff_B_RtEXnXBG7_0(.din(w_dff_B_4U1pC6Ie1_0),.dout(w_dff_B_RtEXnXBG7_0),.clk(gclk));
	jdff dff_B_udzItZ6C4_0(.din(w_dff_B_RtEXnXBG7_0),.dout(w_dff_B_udzItZ6C4_0),.clk(gclk));
	jdff dff_B_weMw1psK9_0(.din(w_dff_B_udzItZ6C4_0),.dout(w_dff_B_weMw1psK9_0),.clk(gclk));
	jdff dff_B_C2G07WEF1_0(.din(w_dff_B_weMw1psK9_0),.dout(w_dff_B_C2G07WEF1_0),.clk(gclk));
	jdff dff_B_8TRDEEBO4_0(.din(w_dff_B_C2G07WEF1_0),.dout(w_dff_B_8TRDEEBO4_0),.clk(gclk));
	jdff dff_B_QB1IXyew8_0(.din(w_dff_B_8TRDEEBO4_0),.dout(w_dff_B_QB1IXyew8_0),.clk(gclk));
	jdff dff_B_qp26auB63_0(.din(w_dff_B_QB1IXyew8_0),.dout(w_dff_B_qp26auB63_0),.clk(gclk));
	jdff dff_B_kI2dXGRk5_0(.din(w_dff_B_qp26auB63_0),.dout(w_dff_B_kI2dXGRk5_0),.clk(gclk));
	jdff dff_B_XqOtYwS99_0(.din(w_dff_B_kI2dXGRk5_0),.dout(w_dff_B_XqOtYwS99_0),.clk(gclk));
	jdff dff_B_YFmMzJDX4_0(.din(w_dff_B_XqOtYwS99_0),.dout(w_dff_B_YFmMzJDX4_0),.clk(gclk));
	jdff dff_B_puvZOHJr3_0(.din(w_dff_B_YFmMzJDX4_0),.dout(w_dff_B_puvZOHJr3_0),.clk(gclk));
	jdff dff_B_MnVza0pd2_0(.din(w_dff_B_puvZOHJr3_0),.dout(w_dff_B_MnVza0pd2_0),.clk(gclk));
	jdff dff_B_GIMAJzJL7_0(.din(w_dff_B_MnVza0pd2_0),.dout(w_dff_B_GIMAJzJL7_0),.clk(gclk));
	jdff dff_B_4exDOfFQ0_0(.din(w_dff_B_GIMAJzJL7_0),.dout(w_dff_B_4exDOfFQ0_0),.clk(gclk));
	jdff dff_B_UnNaBk9q7_0(.din(w_dff_B_4exDOfFQ0_0),.dout(w_dff_B_UnNaBk9q7_0),.clk(gclk));
	jdff dff_B_6jzhcUbu5_0(.din(w_dff_B_UnNaBk9q7_0),.dout(w_dff_B_6jzhcUbu5_0),.clk(gclk));
	jdff dff_B_eM0hB67C3_0(.din(w_dff_B_6jzhcUbu5_0),.dout(w_dff_B_eM0hB67C3_0),.clk(gclk));
	jdff dff_B_s4pMU2ic3_0(.din(w_dff_B_eM0hB67C3_0),.dout(w_dff_B_s4pMU2ic3_0),.clk(gclk));
	jdff dff_B_WV0Zihy29_0(.din(w_dff_B_s4pMU2ic3_0),.dout(w_dff_B_WV0Zihy29_0),.clk(gclk));
	jdff dff_B_A4ytXW2y6_0(.din(w_dff_B_WV0Zihy29_0),.dout(w_dff_B_A4ytXW2y6_0),.clk(gclk));
	jdff dff_B_3mDjKqEZ6_0(.din(w_dff_B_A4ytXW2y6_0),.dout(w_dff_B_3mDjKqEZ6_0),.clk(gclk));
	jdff dff_B_bf2FZPon1_0(.din(w_dff_B_3mDjKqEZ6_0),.dout(w_dff_B_bf2FZPon1_0),.clk(gclk));
	jdff dff_B_xJBqJB2M5_0(.din(w_dff_B_bf2FZPon1_0),.dout(w_dff_B_xJBqJB2M5_0),.clk(gclk));
	jdff dff_B_ZZU372l87_0(.din(w_dff_B_xJBqJB2M5_0),.dout(w_dff_B_ZZU372l87_0),.clk(gclk));
	jdff dff_B_F0kdrYZa2_0(.din(w_dff_B_ZZU372l87_0),.dout(w_dff_B_F0kdrYZa2_0),.clk(gclk));
	jdff dff_B_UiJ1EqSr9_0(.din(w_dff_B_F0kdrYZa2_0),.dout(w_dff_B_UiJ1EqSr9_0),.clk(gclk));
	jdff dff_B_uWwRSsrZ1_0(.din(w_dff_B_UiJ1EqSr9_0),.dout(w_dff_B_uWwRSsrZ1_0),.clk(gclk));
	jdff dff_B_haQDWQAZ6_0(.din(w_dff_B_uWwRSsrZ1_0),.dout(w_dff_B_haQDWQAZ6_0),.clk(gclk));
	jdff dff_B_SwhZn6SF5_0(.din(w_dff_B_haQDWQAZ6_0),.dout(w_dff_B_SwhZn6SF5_0),.clk(gclk));
	jdff dff_B_wezeHtDL5_0(.din(w_dff_B_SwhZn6SF5_0),.dout(w_dff_B_wezeHtDL5_0),.clk(gclk));
	jdff dff_B_RBTvXJq86_0(.din(w_dff_B_wezeHtDL5_0),.dout(w_dff_B_RBTvXJq86_0),.clk(gclk));
	jdff dff_B_mSny4DcO2_0(.din(w_dff_B_RBTvXJq86_0),.dout(w_dff_B_mSny4DcO2_0),.clk(gclk));
	jdff dff_B_KtRvRu983_0(.din(w_dff_B_mSny4DcO2_0),.dout(w_dff_B_KtRvRu983_0),.clk(gclk));
	jdff dff_B_TFZFbgvc4_0(.din(w_dff_B_KtRvRu983_0),.dout(w_dff_B_TFZFbgvc4_0),.clk(gclk));
	jdff dff_B_H4O1GOiU3_0(.din(w_dff_B_TFZFbgvc4_0),.dout(w_dff_B_H4O1GOiU3_0),.clk(gclk));
	jdff dff_B_VSQ0QRtf2_0(.din(w_dff_B_H4O1GOiU3_0),.dout(w_dff_B_VSQ0QRtf2_0),.clk(gclk));
	jdff dff_B_TuVIazGH6_0(.din(w_dff_B_VSQ0QRtf2_0),.dout(w_dff_B_TuVIazGH6_0),.clk(gclk));
	jdff dff_B_nB4Z9b8r8_0(.din(w_dff_B_TuVIazGH6_0),.dout(w_dff_B_nB4Z9b8r8_0),.clk(gclk));
	jdff dff_B_qTBND50X4_0(.din(w_dff_B_nB4Z9b8r8_0),.dout(w_dff_B_qTBND50X4_0),.clk(gclk));
	jdff dff_B_DoYeaq9e6_0(.din(w_dff_B_qTBND50X4_0),.dout(w_dff_B_DoYeaq9e6_0),.clk(gclk));
	jdff dff_B_ijtOPvtT0_0(.din(w_dff_B_DoYeaq9e6_0),.dout(w_dff_B_ijtOPvtT0_0),.clk(gclk));
	jdff dff_B_YUpIWiZ31_0(.din(w_dff_B_ijtOPvtT0_0),.dout(w_dff_B_YUpIWiZ31_0),.clk(gclk));
	jdff dff_B_s266H8zw3_0(.din(w_dff_B_YUpIWiZ31_0),.dout(w_dff_B_s266H8zw3_0),.clk(gclk));
	jdff dff_B_D3oVOrNU8_0(.din(w_dff_B_s266H8zw3_0),.dout(w_dff_B_D3oVOrNU8_0),.clk(gclk));
	jdff dff_B_7aN59Uv71_0(.din(w_dff_B_D3oVOrNU8_0),.dout(w_dff_B_7aN59Uv71_0),.clk(gclk));
	jdff dff_B_uSN6thyP8_0(.din(w_dff_B_7aN59Uv71_0),.dout(w_dff_B_uSN6thyP8_0),.clk(gclk));
	jdff dff_B_ldrRvn527_0(.din(w_dff_B_uSN6thyP8_0),.dout(w_dff_B_ldrRvn527_0),.clk(gclk));
	jdff dff_B_eHTTBcll6_0(.din(w_dff_B_ldrRvn527_0),.dout(w_dff_B_eHTTBcll6_0),.clk(gclk));
	jdff dff_B_vdCbUMJ06_0(.din(w_dff_B_eHTTBcll6_0),.dout(w_dff_B_vdCbUMJ06_0),.clk(gclk));
	jdff dff_B_HvHUCB9z8_0(.din(w_dff_B_vdCbUMJ06_0),.dout(w_dff_B_HvHUCB9z8_0),.clk(gclk));
	jdff dff_B_Sx2NmIou8_0(.din(w_dff_B_HvHUCB9z8_0),.dout(w_dff_B_Sx2NmIou8_0),.clk(gclk));
	jdff dff_B_LbDxoEnS2_0(.din(w_dff_B_Sx2NmIou8_0),.dout(w_dff_B_LbDxoEnS2_0),.clk(gclk));
	jdff dff_B_GKtRYPrW2_1(.din(n888),.dout(w_dff_B_GKtRYPrW2_1),.clk(gclk));
	jdff dff_B_3F1aMPwX3_1(.din(w_dff_B_GKtRYPrW2_1),.dout(w_dff_B_3F1aMPwX3_1),.clk(gclk));
	jdff dff_B_7ipyUibD1_1(.din(w_dff_B_3F1aMPwX3_1),.dout(w_dff_B_7ipyUibD1_1),.clk(gclk));
	jdff dff_B_3Z4uc6Es6_1(.din(w_dff_B_7ipyUibD1_1),.dout(w_dff_B_3Z4uc6Es6_1),.clk(gclk));
	jdff dff_B_RprIe1Dt1_1(.din(w_dff_B_3Z4uc6Es6_1),.dout(w_dff_B_RprIe1Dt1_1),.clk(gclk));
	jdff dff_B_rjLJBud54_1(.din(w_dff_B_RprIe1Dt1_1),.dout(w_dff_B_rjLJBud54_1),.clk(gclk));
	jdff dff_B_8fv1Bf5S2_1(.din(w_dff_B_rjLJBud54_1),.dout(w_dff_B_8fv1Bf5S2_1),.clk(gclk));
	jdff dff_B_ZrPlNy286_1(.din(w_dff_B_8fv1Bf5S2_1),.dout(w_dff_B_ZrPlNy286_1),.clk(gclk));
	jdff dff_B_9W4sielV8_1(.din(w_dff_B_ZrPlNy286_1),.dout(w_dff_B_9W4sielV8_1),.clk(gclk));
	jdff dff_B_Kt2JAZpY6_1(.din(w_dff_B_9W4sielV8_1),.dout(w_dff_B_Kt2JAZpY6_1),.clk(gclk));
	jdff dff_B_HCpcGmzM1_1(.din(w_dff_B_Kt2JAZpY6_1),.dout(w_dff_B_HCpcGmzM1_1),.clk(gclk));
	jdff dff_B_cx7bQocO7_1(.din(w_dff_B_HCpcGmzM1_1),.dout(w_dff_B_cx7bQocO7_1),.clk(gclk));
	jdff dff_B_EhfcKy846_1(.din(w_dff_B_cx7bQocO7_1),.dout(w_dff_B_EhfcKy846_1),.clk(gclk));
	jdff dff_B_tphxZSMk1_1(.din(w_dff_B_EhfcKy846_1),.dout(w_dff_B_tphxZSMk1_1),.clk(gclk));
	jdff dff_B_Ndad2jbe8_1(.din(w_dff_B_tphxZSMk1_1),.dout(w_dff_B_Ndad2jbe8_1),.clk(gclk));
	jdff dff_B_hS1wXzlv5_1(.din(w_dff_B_Ndad2jbe8_1),.dout(w_dff_B_hS1wXzlv5_1),.clk(gclk));
	jdff dff_B_jtawZMZS5_1(.din(w_dff_B_hS1wXzlv5_1),.dout(w_dff_B_jtawZMZS5_1),.clk(gclk));
	jdff dff_B_rqfDRn3X2_1(.din(w_dff_B_jtawZMZS5_1),.dout(w_dff_B_rqfDRn3X2_1),.clk(gclk));
	jdff dff_B_r6g8H71W1_1(.din(w_dff_B_rqfDRn3X2_1),.dout(w_dff_B_r6g8H71W1_1),.clk(gclk));
	jdff dff_B_sqEqgQik3_1(.din(w_dff_B_r6g8H71W1_1),.dout(w_dff_B_sqEqgQik3_1),.clk(gclk));
	jdff dff_B_Ws5szzQx2_1(.din(w_dff_B_sqEqgQik3_1),.dout(w_dff_B_Ws5szzQx2_1),.clk(gclk));
	jdff dff_B_sjsLXqOQ3_1(.din(w_dff_B_Ws5szzQx2_1),.dout(w_dff_B_sjsLXqOQ3_1),.clk(gclk));
	jdff dff_B_GmlnaTke8_1(.din(w_dff_B_sjsLXqOQ3_1),.dout(w_dff_B_GmlnaTke8_1),.clk(gclk));
	jdff dff_B_B5BYmlYS1_1(.din(w_dff_B_GmlnaTke8_1),.dout(w_dff_B_B5BYmlYS1_1),.clk(gclk));
	jdff dff_B_QKoKqY614_1(.din(w_dff_B_B5BYmlYS1_1),.dout(w_dff_B_QKoKqY614_1),.clk(gclk));
	jdff dff_B_7Chx3MfP0_1(.din(w_dff_B_QKoKqY614_1),.dout(w_dff_B_7Chx3MfP0_1),.clk(gclk));
	jdff dff_B_LGkYfDpn3_1(.din(w_dff_B_7Chx3MfP0_1),.dout(w_dff_B_LGkYfDpn3_1),.clk(gclk));
	jdff dff_B_gudizypC1_1(.din(w_dff_B_LGkYfDpn3_1),.dout(w_dff_B_gudizypC1_1),.clk(gclk));
	jdff dff_B_jHkHUqva5_1(.din(w_dff_B_gudizypC1_1),.dout(w_dff_B_jHkHUqva5_1),.clk(gclk));
	jdff dff_B_dQCzMzMy0_1(.din(w_dff_B_jHkHUqva5_1),.dout(w_dff_B_dQCzMzMy0_1),.clk(gclk));
	jdff dff_B_OF3ywdzv0_1(.din(w_dff_B_dQCzMzMy0_1),.dout(w_dff_B_OF3ywdzv0_1),.clk(gclk));
	jdff dff_B_E3TqWAjh0_1(.din(w_dff_B_OF3ywdzv0_1),.dout(w_dff_B_E3TqWAjh0_1),.clk(gclk));
	jdff dff_B_HBSvAhJa4_1(.din(w_dff_B_E3TqWAjh0_1),.dout(w_dff_B_HBSvAhJa4_1),.clk(gclk));
	jdff dff_B_itaB3R5g2_1(.din(w_dff_B_HBSvAhJa4_1),.dout(w_dff_B_itaB3R5g2_1),.clk(gclk));
	jdff dff_B_SD4QNh4g1_1(.din(w_dff_B_itaB3R5g2_1),.dout(w_dff_B_SD4QNh4g1_1),.clk(gclk));
	jdff dff_B_XvZXIE296_1(.din(w_dff_B_SD4QNh4g1_1),.dout(w_dff_B_XvZXIE296_1),.clk(gclk));
	jdff dff_B_K87zYtj92_1(.din(w_dff_B_XvZXIE296_1),.dout(w_dff_B_K87zYtj92_1),.clk(gclk));
	jdff dff_B_2qWdqTH73_1(.din(w_dff_B_K87zYtj92_1),.dout(w_dff_B_2qWdqTH73_1),.clk(gclk));
	jdff dff_B_4odDBRJw6_1(.din(w_dff_B_2qWdqTH73_1),.dout(w_dff_B_4odDBRJw6_1),.clk(gclk));
	jdff dff_B_BBh2S4Na3_1(.din(w_dff_B_4odDBRJw6_1),.dout(w_dff_B_BBh2S4Na3_1),.clk(gclk));
	jdff dff_B_cnhIEryX7_1(.din(w_dff_B_BBh2S4Na3_1),.dout(w_dff_B_cnhIEryX7_1),.clk(gclk));
	jdff dff_B_ztrWRd7J8_1(.din(w_dff_B_cnhIEryX7_1),.dout(w_dff_B_ztrWRd7J8_1),.clk(gclk));
	jdff dff_B_j39FyQzb7_1(.din(w_dff_B_ztrWRd7J8_1),.dout(w_dff_B_j39FyQzb7_1),.clk(gclk));
	jdff dff_B_eBM8205w1_1(.din(w_dff_B_j39FyQzb7_1),.dout(w_dff_B_eBM8205w1_1),.clk(gclk));
	jdff dff_B_CURzSjlm4_1(.din(w_dff_B_eBM8205w1_1),.dout(w_dff_B_CURzSjlm4_1),.clk(gclk));
	jdff dff_B_Q4VwXRyH6_1(.din(w_dff_B_CURzSjlm4_1),.dout(w_dff_B_Q4VwXRyH6_1),.clk(gclk));
	jdff dff_B_8xYdzrIY1_1(.din(w_dff_B_Q4VwXRyH6_1),.dout(w_dff_B_8xYdzrIY1_1),.clk(gclk));
	jdff dff_B_4yV7nJBP4_1(.din(w_dff_B_8xYdzrIY1_1),.dout(w_dff_B_4yV7nJBP4_1),.clk(gclk));
	jdff dff_B_l6Ltd7GT5_1(.din(w_dff_B_4yV7nJBP4_1),.dout(w_dff_B_l6Ltd7GT5_1),.clk(gclk));
	jdff dff_B_qMEhjrSU0_1(.din(w_dff_B_l6Ltd7GT5_1),.dout(w_dff_B_qMEhjrSU0_1),.clk(gclk));
	jdff dff_B_tnyo2G0o6_1(.din(w_dff_B_qMEhjrSU0_1),.dout(w_dff_B_tnyo2G0o6_1),.clk(gclk));
	jdff dff_B_u3kneydC3_1(.din(w_dff_B_tnyo2G0o6_1),.dout(w_dff_B_u3kneydC3_1),.clk(gclk));
	jdff dff_B_nj8hUOoP3_1(.din(w_dff_B_u3kneydC3_1),.dout(w_dff_B_nj8hUOoP3_1),.clk(gclk));
	jdff dff_B_S1fm64og5_1(.din(w_dff_B_nj8hUOoP3_1),.dout(w_dff_B_S1fm64og5_1),.clk(gclk));
	jdff dff_B_8e04RCjO4_1(.din(w_dff_B_S1fm64og5_1),.dout(w_dff_B_8e04RCjO4_1),.clk(gclk));
	jdff dff_B_JIUf7FBz2_1(.din(w_dff_B_8e04RCjO4_1),.dout(w_dff_B_JIUf7FBz2_1),.clk(gclk));
	jdff dff_B_5pIGDXSh9_1(.din(w_dff_B_JIUf7FBz2_1),.dout(w_dff_B_5pIGDXSh9_1),.clk(gclk));
	jdff dff_B_bu60NKrG4_1(.din(w_dff_B_5pIGDXSh9_1),.dout(w_dff_B_bu60NKrG4_1),.clk(gclk));
	jdff dff_B_97A3pkXr7_1(.din(w_dff_B_bu60NKrG4_1),.dout(w_dff_B_97A3pkXr7_1),.clk(gclk));
	jdff dff_B_tuagi6Ba0_1(.din(w_dff_B_97A3pkXr7_1),.dout(w_dff_B_tuagi6Ba0_1),.clk(gclk));
	jdff dff_B_u5SYOHUA9_1(.din(w_dff_B_tuagi6Ba0_1),.dout(w_dff_B_u5SYOHUA9_1),.clk(gclk));
	jdff dff_B_Kd09eGeT9_1(.din(w_dff_B_u5SYOHUA9_1),.dout(w_dff_B_Kd09eGeT9_1),.clk(gclk));
	jdff dff_B_UWURkiLl8_1(.din(w_dff_B_Kd09eGeT9_1),.dout(w_dff_B_UWURkiLl8_1),.clk(gclk));
	jdff dff_B_bHHS2Dnx6_1(.din(w_dff_B_UWURkiLl8_1),.dout(w_dff_B_bHHS2Dnx6_1),.clk(gclk));
	jdff dff_B_CYcAG6bC2_1(.din(w_dff_B_bHHS2Dnx6_1),.dout(w_dff_B_CYcAG6bC2_1),.clk(gclk));
	jdff dff_B_ZQ5XIhPt2_1(.din(w_dff_B_CYcAG6bC2_1),.dout(w_dff_B_ZQ5XIhPt2_1),.clk(gclk));
	jdff dff_B_9DhvbhLG9_1(.din(w_dff_B_ZQ5XIhPt2_1),.dout(w_dff_B_9DhvbhLG9_1),.clk(gclk));
	jdff dff_B_mwg3qWgc6_1(.din(w_dff_B_9DhvbhLG9_1),.dout(w_dff_B_mwg3qWgc6_1),.clk(gclk));
	jdff dff_B_Od2dIDMp2_1(.din(w_dff_B_mwg3qWgc6_1),.dout(w_dff_B_Od2dIDMp2_1),.clk(gclk));
	jdff dff_B_PY1v2Rwt9_1(.din(w_dff_B_Od2dIDMp2_1),.dout(w_dff_B_PY1v2Rwt9_1),.clk(gclk));
	jdff dff_B_vSuWtJfl2_1(.din(w_dff_B_PY1v2Rwt9_1),.dout(w_dff_B_vSuWtJfl2_1),.clk(gclk));
	jdff dff_B_MukH1qL56_1(.din(w_dff_B_vSuWtJfl2_1),.dout(w_dff_B_MukH1qL56_1),.clk(gclk));
	jdff dff_B_oC8QApYL6_1(.din(w_dff_B_MukH1qL56_1),.dout(w_dff_B_oC8QApYL6_1),.clk(gclk));
	jdff dff_B_2AeYhtpO0_1(.din(w_dff_B_oC8QApYL6_1),.dout(w_dff_B_2AeYhtpO0_1),.clk(gclk));
	jdff dff_B_nyqwvJoK4_1(.din(w_dff_B_2AeYhtpO0_1),.dout(w_dff_B_nyqwvJoK4_1),.clk(gclk));
	jdff dff_B_ysxui0172_1(.din(w_dff_B_nyqwvJoK4_1),.dout(w_dff_B_ysxui0172_1),.clk(gclk));
	jdff dff_B_LVVtV4Qm1_1(.din(w_dff_B_ysxui0172_1),.dout(w_dff_B_LVVtV4Qm1_1),.clk(gclk));
	jdff dff_B_FMVPXCWy1_1(.din(w_dff_B_LVVtV4Qm1_1),.dout(w_dff_B_FMVPXCWy1_1),.clk(gclk));
	jdff dff_B_COstpe8X7_1(.din(w_dff_B_FMVPXCWy1_1),.dout(w_dff_B_COstpe8X7_1),.clk(gclk));
	jdff dff_B_CBkZ6ETZ4_1(.din(w_dff_B_COstpe8X7_1),.dout(w_dff_B_CBkZ6ETZ4_1),.clk(gclk));
	jdff dff_B_Vbuzfyop4_1(.din(w_dff_B_CBkZ6ETZ4_1),.dout(w_dff_B_Vbuzfyop4_1),.clk(gclk));
	jdff dff_B_FjY0zC7k0_1(.din(w_dff_B_Vbuzfyop4_1),.dout(w_dff_B_FjY0zC7k0_1),.clk(gclk));
	jdff dff_B_n0qrL1M48_1(.din(w_dff_B_FjY0zC7k0_1),.dout(w_dff_B_n0qrL1M48_1),.clk(gclk));
	jdff dff_B_etx97ig43_1(.din(w_dff_B_n0qrL1M48_1),.dout(w_dff_B_etx97ig43_1),.clk(gclk));
	jdff dff_B_IS9gqbo12_0(.din(n889),.dout(w_dff_B_IS9gqbo12_0),.clk(gclk));
	jdff dff_B_9Vj3Nt8X5_0(.din(w_dff_B_IS9gqbo12_0),.dout(w_dff_B_9Vj3Nt8X5_0),.clk(gclk));
	jdff dff_B_SXu1pMQS5_0(.din(w_dff_B_9Vj3Nt8X5_0),.dout(w_dff_B_SXu1pMQS5_0),.clk(gclk));
	jdff dff_B_n3WVT6mU1_0(.din(w_dff_B_SXu1pMQS5_0),.dout(w_dff_B_n3WVT6mU1_0),.clk(gclk));
	jdff dff_B_raRSMuC74_0(.din(w_dff_B_n3WVT6mU1_0),.dout(w_dff_B_raRSMuC74_0),.clk(gclk));
	jdff dff_B_fPUHfe4T1_0(.din(w_dff_B_raRSMuC74_0),.dout(w_dff_B_fPUHfe4T1_0),.clk(gclk));
	jdff dff_B_5vzL2BVh1_0(.din(w_dff_B_fPUHfe4T1_0),.dout(w_dff_B_5vzL2BVh1_0),.clk(gclk));
	jdff dff_B_2OmAh31x7_0(.din(w_dff_B_5vzL2BVh1_0),.dout(w_dff_B_2OmAh31x7_0),.clk(gclk));
	jdff dff_B_zJ4FtWxm1_0(.din(w_dff_B_2OmAh31x7_0),.dout(w_dff_B_zJ4FtWxm1_0),.clk(gclk));
	jdff dff_B_JsgkxfMI9_0(.din(w_dff_B_zJ4FtWxm1_0),.dout(w_dff_B_JsgkxfMI9_0),.clk(gclk));
	jdff dff_B_blQQ2uMx4_0(.din(w_dff_B_JsgkxfMI9_0),.dout(w_dff_B_blQQ2uMx4_0),.clk(gclk));
	jdff dff_B_gepnvB4j8_0(.din(w_dff_B_blQQ2uMx4_0),.dout(w_dff_B_gepnvB4j8_0),.clk(gclk));
	jdff dff_B_oX5E9BmF8_0(.din(w_dff_B_gepnvB4j8_0),.dout(w_dff_B_oX5E9BmF8_0),.clk(gclk));
	jdff dff_B_HVeHePan1_0(.din(w_dff_B_oX5E9BmF8_0),.dout(w_dff_B_HVeHePan1_0),.clk(gclk));
	jdff dff_B_zHp0ZRjP8_0(.din(w_dff_B_HVeHePan1_0),.dout(w_dff_B_zHp0ZRjP8_0),.clk(gclk));
	jdff dff_B_vXtK9Mlt5_0(.din(w_dff_B_zHp0ZRjP8_0),.dout(w_dff_B_vXtK9Mlt5_0),.clk(gclk));
	jdff dff_B_h7tdAW7D8_0(.din(w_dff_B_vXtK9Mlt5_0),.dout(w_dff_B_h7tdAW7D8_0),.clk(gclk));
	jdff dff_B_Zlikh2j86_0(.din(w_dff_B_h7tdAW7D8_0),.dout(w_dff_B_Zlikh2j86_0),.clk(gclk));
	jdff dff_B_VPTpC2H45_0(.din(w_dff_B_Zlikh2j86_0),.dout(w_dff_B_VPTpC2H45_0),.clk(gclk));
	jdff dff_B_VvMr97nE3_0(.din(w_dff_B_VPTpC2H45_0),.dout(w_dff_B_VvMr97nE3_0),.clk(gclk));
	jdff dff_B_NahAC0Eo9_0(.din(w_dff_B_VvMr97nE3_0),.dout(w_dff_B_NahAC0Eo9_0),.clk(gclk));
	jdff dff_B_280qH7kL6_0(.din(w_dff_B_NahAC0Eo9_0),.dout(w_dff_B_280qH7kL6_0),.clk(gclk));
	jdff dff_B_MlKTwdTh4_0(.din(w_dff_B_280qH7kL6_0),.dout(w_dff_B_MlKTwdTh4_0),.clk(gclk));
	jdff dff_B_aGjj0Nh93_0(.din(w_dff_B_MlKTwdTh4_0),.dout(w_dff_B_aGjj0Nh93_0),.clk(gclk));
	jdff dff_B_LAOfmeim3_0(.din(w_dff_B_aGjj0Nh93_0),.dout(w_dff_B_LAOfmeim3_0),.clk(gclk));
	jdff dff_B_h0ZQAsrA1_0(.din(w_dff_B_LAOfmeim3_0),.dout(w_dff_B_h0ZQAsrA1_0),.clk(gclk));
	jdff dff_B_Rbgkyd2G8_0(.din(w_dff_B_h0ZQAsrA1_0),.dout(w_dff_B_Rbgkyd2G8_0),.clk(gclk));
	jdff dff_B_RUOWKRLc3_0(.din(w_dff_B_Rbgkyd2G8_0),.dout(w_dff_B_RUOWKRLc3_0),.clk(gclk));
	jdff dff_B_Zqy47IMD9_0(.din(w_dff_B_RUOWKRLc3_0),.dout(w_dff_B_Zqy47IMD9_0),.clk(gclk));
	jdff dff_B_Xck9EUzY8_0(.din(w_dff_B_Zqy47IMD9_0),.dout(w_dff_B_Xck9EUzY8_0),.clk(gclk));
	jdff dff_B_ypyvD6Bz4_0(.din(w_dff_B_Xck9EUzY8_0),.dout(w_dff_B_ypyvD6Bz4_0),.clk(gclk));
	jdff dff_B_HpUYi8oQ3_0(.din(w_dff_B_ypyvD6Bz4_0),.dout(w_dff_B_HpUYi8oQ3_0),.clk(gclk));
	jdff dff_B_cRZ5Imnm4_0(.din(w_dff_B_HpUYi8oQ3_0),.dout(w_dff_B_cRZ5Imnm4_0),.clk(gclk));
	jdff dff_B_mDCQl1v25_0(.din(w_dff_B_cRZ5Imnm4_0),.dout(w_dff_B_mDCQl1v25_0),.clk(gclk));
	jdff dff_B_mIiKfnyG8_0(.din(w_dff_B_mDCQl1v25_0),.dout(w_dff_B_mIiKfnyG8_0),.clk(gclk));
	jdff dff_B_lgZJCgZP1_0(.din(w_dff_B_mIiKfnyG8_0),.dout(w_dff_B_lgZJCgZP1_0),.clk(gclk));
	jdff dff_B_7ndmbS6K9_0(.din(w_dff_B_lgZJCgZP1_0),.dout(w_dff_B_7ndmbS6K9_0),.clk(gclk));
	jdff dff_B_rTCVd5N99_0(.din(w_dff_B_7ndmbS6K9_0),.dout(w_dff_B_rTCVd5N99_0),.clk(gclk));
	jdff dff_B_7E3pJjH17_0(.din(w_dff_B_rTCVd5N99_0),.dout(w_dff_B_7E3pJjH17_0),.clk(gclk));
	jdff dff_B_g6nplmB82_0(.din(w_dff_B_7E3pJjH17_0),.dout(w_dff_B_g6nplmB82_0),.clk(gclk));
	jdff dff_B_h9cRijoQ3_0(.din(w_dff_B_g6nplmB82_0),.dout(w_dff_B_h9cRijoQ3_0),.clk(gclk));
	jdff dff_B_fFVisHlT2_0(.din(w_dff_B_h9cRijoQ3_0),.dout(w_dff_B_fFVisHlT2_0),.clk(gclk));
	jdff dff_B_FIWK01KE2_0(.din(w_dff_B_fFVisHlT2_0),.dout(w_dff_B_FIWK01KE2_0),.clk(gclk));
	jdff dff_B_gs5iODbn6_0(.din(w_dff_B_FIWK01KE2_0),.dout(w_dff_B_gs5iODbn6_0),.clk(gclk));
	jdff dff_B_DMyofCCZ7_0(.din(w_dff_B_gs5iODbn6_0),.dout(w_dff_B_DMyofCCZ7_0),.clk(gclk));
	jdff dff_B_bhVr24TV4_0(.din(w_dff_B_DMyofCCZ7_0),.dout(w_dff_B_bhVr24TV4_0),.clk(gclk));
	jdff dff_B_tI6gCD1J8_0(.din(w_dff_B_bhVr24TV4_0),.dout(w_dff_B_tI6gCD1J8_0),.clk(gclk));
	jdff dff_B_Q3fAfedx4_0(.din(w_dff_B_tI6gCD1J8_0),.dout(w_dff_B_Q3fAfedx4_0),.clk(gclk));
	jdff dff_B_2hHLb52J6_0(.din(w_dff_B_Q3fAfedx4_0),.dout(w_dff_B_2hHLb52J6_0),.clk(gclk));
	jdff dff_B_UXHygEj31_0(.din(w_dff_B_2hHLb52J6_0),.dout(w_dff_B_UXHygEj31_0),.clk(gclk));
	jdff dff_B_MPWVDqaN0_0(.din(w_dff_B_UXHygEj31_0),.dout(w_dff_B_MPWVDqaN0_0),.clk(gclk));
	jdff dff_B_dwHbIRQV6_0(.din(w_dff_B_MPWVDqaN0_0),.dout(w_dff_B_dwHbIRQV6_0),.clk(gclk));
	jdff dff_B_kFtrtvSs1_0(.din(w_dff_B_dwHbIRQV6_0),.dout(w_dff_B_kFtrtvSs1_0),.clk(gclk));
	jdff dff_B_Ys4FiAHx0_0(.din(w_dff_B_kFtrtvSs1_0),.dout(w_dff_B_Ys4FiAHx0_0),.clk(gclk));
	jdff dff_B_9YrrfuX94_0(.din(w_dff_B_Ys4FiAHx0_0),.dout(w_dff_B_9YrrfuX94_0),.clk(gclk));
	jdff dff_B_5AGYM25N5_0(.din(w_dff_B_9YrrfuX94_0),.dout(w_dff_B_5AGYM25N5_0),.clk(gclk));
	jdff dff_B_qHUkpTyI3_0(.din(w_dff_B_5AGYM25N5_0),.dout(w_dff_B_qHUkpTyI3_0),.clk(gclk));
	jdff dff_B_fOUDaivR3_0(.din(w_dff_B_qHUkpTyI3_0),.dout(w_dff_B_fOUDaivR3_0),.clk(gclk));
	jdff dff_B_alYZk9ks1_0(.din(w_dff_B_fOUDaivR3_0),.dout(w_dff_B_alYZk9ks1_0),.clk(gclk));
	jdff dff_B_IO2CtH3y3_0(.din(w_dff_B_alYZk9ks1_0),.dout(w_dff_B_IO2CtH3y3_0),.clk(gclk));
	jdff dff_B_KtHIdWub0_0(.din(w_dff_B_IO2CtH3y3_0),.dout(w_dff_B_KtHIdWub0_0),.clk(gclk));
	jdff dff_B_XP0zdyAC9_0(.din(w_dff_B_KtHIdWub0_0),.dout(w_dff_B_XP0zdyAC9_0),.clk(gclk));
	jdff dff_B_zU4AQxrN6_0(.din(w_dff_B_XP0zdyAC9_0),.dout(w_dff_B_zU4AQxrN6_0),.clk(gclk));
	jdff dff_B_UcJWm4uf0_0(.din(w_dff_B_zU4AQxrN6_0),.dout(w_dff_B_UcJWm4uf0_0),.clk(gclk));
	jdff dff_B_uiSNVyjp4_0(.din(w_dff_B_UcJWm4uf0_0),.dout(w_dff_B_uiSNVyjp4_0),.clk(gclk));
	jdff dff_B_QZiYkCeo5_0(.din(w_dff_B_uiSNVyjp4_0),.dout(w_dff_B_QZiYkCeo5_0),.clk(gclk));
	jdff dff_B_V9sIaIe34_0(.din(w_dff_B_QZiYkCeo5_0),.dout(w_dff_B_V9sIaIe34_0),.clk(gclk));
	jdff dff_B_mRo9FUhG9_0(.din(w_dff_B_V9sIaIe34_0),.dout(w_dff_B_mRo9FUhG9_0),.clk(gclk));
	jdff dff_B_32yQTYIV2_0(.din(w_dff_B_mRo9FUhG9_0),.dout(w_dff_B_32yQTYIV2_0),.clk(gclk));
	jdff dff_B_50EwaRSy4_0(.din(w_dff_B_32yQTYIV2_0),.dout(w_dff_B_50EwaRSy4_0),.clk(gclk));
	jdff dff_B_ekMlRWdn7_0(.din(w_dff_B_50EwaRSy4_0),.dout(w_dff_B_ekMlRWdn7_0),.clk(gclk));
	jdff dff_B_Em4aZHXi9_0(.din(w_dff_B_ekMlRWdn7_0),.dout(w_dff_B_Em4aZHXi9_0),.clk(gclk));
	jdff dff_B_kEpVFEnH7_0(.din(w_dff_B_Em4aZHXi9_0),.dout(w_dff_B_kEpVFEnH7_0),.clk(gclk));
	jdff dff_B_YZgb51P05_0(.din(w_dff_B_kEpVFEnH7_0),.dout(w_dff_B_YZgb51P05_0),.clk(gclk));
	jdff dff_B_WxaoF8hO3_0(.din(w_dff_B_YZgb51P05_0),.dout(w_dff_B_WxaoF8hO3_0),.clk(gclk));
	jdff dff_B_44JFbs0e0_0(.din(w_dff_B_WxaoF8hO3_0),.dout(w_dff_B_44JFbs0e0_0),.clk(gclk));
	jdff dff_B_bWFses4t8_0(.din(w_dff_B_44JFbs0e0_0),.dout(w_dff_B_bWFses4t8_0),.clk(gclk));
	jdff dff_B_EVWYhNQk7_0(.din(w_dff_B_bWFses4t8_0),.dout(w_dff_B_EVWYhNQk7_0),.clk(gclk));
	jdff dff_B_fEoxjw221_0(.din(w_dff_B_EVWYhNQk7_0),.dout(w_dff_B_fEoxjw221_0),.clk(gclk));
	jdff dff_B_SJ3NDSfr7_0(.din(w_dff_B_fEoxjw221_0),.dout(w_dff_B_SJ3NDSfr7_0),.clk(gclk));
	jdff dff_B_xf81cLkS2_0(.din(w_dff_B_SJ3NDSfr7_0),.dout(w_dff_B_xf81cLkS2_0),.clk(gclk));
	jdff dff_B_NfmeXSyA9_0(.din(w_dff_B_xf81cLkS2_0),.dout(w_dff_B_NfmeXSyA9_0),.clk(gclk));
	jdff dff_B_ihb62fBO1_0(.din(w_dff_B_NfmeXSyA9_0),.dout(w_dff_B_ihb62fBO1_0),.clk(gclk));
	jdff dff_B_mRYvO6bw1_0(.din(w_dff_B_ihb62fBO1_0),.dout(w_dff_B_mRYvO6bw1_0),.clk(gclk));
	jdff dff_B_Mq8qISei8_1(.din(n882),.dout(w_dff_B_Mq8qISei8_1),.clk(gclk));
	jdff dff_B_zVwl7onX2_1(.din(w_dff_B_Mq8qISei8_1),.dout(w_dff_B_zVwl7onX2_1),.clk(gclk));
	jdff dff_B_jkhEDHER3_1(.din(w_dff_B_zVwl7onX2_1),.dout(w_dff_B_jkhEDHER3_1),.clk(gclk));
	jdff dff_B_sjCYmBud1_1(.din(w_dff_B_jkhEDHER3_1),.dout(w_dff_B_sjCYmBud1_1),.clk(gclk));
	jdff dff_B_jovfwT9y8_1(.din(w_dff_B_sjCYmBud1_1),.dout(w_dff_B_jovfwT9y8_1),.clk(gclk));
	jdff dff_B_dByslP4G1_1(.din(w_dff_B_jovfwT9y8_1),.dout(w_dff_B_dByslP4G1_1),.clk(gclk));
	jdff dff_B_TqaYnsJW8_1(.din(w_dff_B_dByslP4G1_1),.dout(w_dff_B_TqaYnsJW8_1),.clk(gclk));
	jdff dff_B_2N9Enggv5_1(.din(w_dff_B_TqaYnsJW8_1),.dout(w_dff_B_2N9Enggv5_1),.clk(gclk));
	jdff dff_B_M2l7D4P54_1(.din(w_dff_B_2N9Enggv5_1),.dout(w_dff_B_M2l7D4P54_1),.clk(gclk));
	jdff dff_B_CUaXZ9OF8_1(.din(w_dff_B_M2l7D4P54_1),.dout(w_dff_B_CUaXZ9OF8_1),.clk(gclk));
	jdff dff_B_ajq5lKV57_1(.din(w_dff_B_CUaXZ9OF8_1),.dout(w_dff_B_ajq5lKV57_1),.clk(gclk));
	jdff dff_B_0Oeh6Ivd1_1(.din(w_dff_B_ajq5lKV57_1),.dout(w_dff_B_0Oeh6Ivd1_1),.clk(gclk));
	jdff dff_B_ALDAxfQp4_1(.din(w_dff_B_0Oeh6Ivd1_1),.dout(w_dff_B_ALDAxfQp4_1),.clk(gclk));
	jdff dff_B_XujCND2b7_1(.din(w_dff_B_ALDAxfQp4_1),.dout(w_dff_B_XujCND2b7_1),.clk(gclk));
	jdff dff_B_YZ3L0UOX4_1(.din(w_dff_B_XujCND2b7_1),.dout(w_dff_B_YZ3L0UOX4_1),.clk(gclk));
	jdff dff_B_wLzp8yy96_1(.din(w_dff_B_YZ3L0UOX4_1),.dout(w_dff_B_wLzp8yy96_1),.clk(gclk));
	jdff dff_B_1W53RdhW9_1(.din(w_dff_B_wLzp8yy96_1),.dout(w_dff_B_1W53RdhW9_1),.clk(gclk));
	jdff dff_B_8sVhLcJ53_1(.din(w_dff_B_1W53RdhW9_1),.dout(w_dff_B_8sVhLcJ53_1),.clk(gclk));
	jdff dff_B_VneuQfHg2_1(.din(w_dff_B_8sVhLcJ53_1),.dout(w_dff_B_VneuQfHg2_1),.clk(gclk));
	jdff dff_B_d9oWTCcI3_1(.din(w_dff_B_VneuQfHg2_1),.dout(w_dff_B_d9oWTCcI3_1),.clk(gclk));
	jdff dff_B_Ib90Bc2V6_1(.din(w_dff_B_d9oWTCcI3_1),.dout(w_dff_B_Ib90Bc2V6_1),.clk(gclk));
	jdff dff_B_ZO7bX5aP4_1(.din(w_dff_B_Ib90Bc2V6_1),.dout(w_dff_B_ZO7bX5aP4_1),.clk(gclk));
	jdff dff_B_fy2DG2792_1(.din(w_dff_B_ZO7bX5aP4_1),.dout(w_dff_B_fy2DG2792_1),.clk(gclk));
	jdff dff_B_x9u41iBL8_1(.din(w_dff_B_fy2DG2792_1),.dout(w_dff_B_x9u41iBL8_1),.clk(gclk));
	jdff dff_B_qBqDGxo13_1(.din(w_dff_B_x9u41iBL8_1),.dout(w_dff_B_qBqDGxo13_1),.clk(gclk));
	jdff dff_B_HZUFPXbX1_1(.din(w_dff_B_qBqDGxo13_1),.dout(w_dff_B_HZUFPXbX1_1),.clk(gclk));
	jdff dff_B_piUxztbY6_1(.din(w_dff_B_HZUFPXbX1_1),.dout(w_dff_B_piUxztbY6_1),.clk(gclk));
	jdff dff_B_KTdvDgsl7_1(.din(w_dff_B_piUxztbY6_1),.dout(w_dff_B_KTdvDgsl7_1),.clk(gclk));
	jdff dff_B_0ejnl01W7_1(.din(w_dff_B_KTdvDgsl7_1),.dout(w_dff_B_0ejnl01W7_1),.clk(gclk));
	jdff dff_B_gmtA3fTG3_1(.din(w_dff_B_0ejnl01W7_1),.dout(w_dff_B_gmtA3fTG3_1),.clk(gclk));
	jdff dff_B_ZeE6vPmm5_1(.din(w_dff_B_gmtA3fTG3_1),.dout(w_dff_B_ZeE6vPmm5_1),.clk(gclk));
	jdff dff_B_pkTlWEEt6_1(.din(w_dff_B_ZeE6vPmm5_1),.dout(w_dff_B_pkTlWEEt6_1),.clk(gclk));
	jdff dff_B_K0xiAILb1_1(.din(w_dff_B_pkTlWEEt6_1),.dout(w_dff_B_K0xiAILb1_1),.clk(gclk));
	jdff dff_B_Fa6nHqKX9_1(.din(w_dff_B_K0xiAILb1_1),.dout(w_dff_B_Fa6nHqKX9_1),.clk(gclk));
	jdff dff_B_iP1Y05CH9_1(.din(w_dff_B_Fa6nHqKX9_1),.dout(w_dff_B_iP1Y05CH9_1),.clk(gclk));
	jdff dff_B_hSyM2ESL0_1(.din(w_dff_B_iP1Y05CH9_1),.dout(w_dff_B_hSyM2ESL0_1),.clk(gclk));
	jdff dff_B_SUJ9gpXS1_1(.din(w_dff_B_hSyM2ESL0_1),.dout(w_dff_B_SUJ9gpXS1_1),.clk(gclk));
	jdff dff_B_Gj7GG32j2_1(.din(w_dff_B_SUJ9gpXS1_1),.dout(w_dff_B_Gj7GG32j2_1),.clk(gclk));
	jdff dff_B_o68rxA8H6_1(.din(w_dff_B_Gj7GG32j2_1),.dout(w_dff_B_o68rxA8H6_1),.clk(gclk));
	jdff dff_B_Rr9TWc367_1(.din(w_dff_B_o68rxA8H6_1),.dout(w_dff_B_Rr9TWc367_1),.clk(gclk));
	jdff dff_B_NDxObvPn9_1(.din(w_dff_B_Rr9TWc367_1),.dout(w_dff_B_NDxObvPn9_1),.clk(gclk));
	jdff dff_B_dPqgRTiZ7_1(.din(w_dff_B_NDxObvPn9_1),.dout(w_dff_B_dPqgRTiZ7_1),.clk(gclk));
	jdff dff_B_6vK1fI4O5_1(.din(w_dff_B_dPqgRTiZ7_1),.dout(w_dff_B_6vK1fI4O5_1),.clk(gclk));
	jdff dff_B_IYn3bxHz2_1(.din(w_dff_B_6vK1fI4O5_1),.dout(w_dff_B_IYn3bxHz2_1),.clk(gclk));
	jdff dff_B_qVwDrg6t2_1(.din(w_dff_B_IYn3bxHz2_1),.dout(w_dff_B_qVwDrg6t2_1),.clk(gclk));
	jdff dff_B_ia5XpHfb1_1(.din(w_dff_B_qVwDrg6t2_1),.dout(w_dff_B_ia5XpHfb1_1),.clk(gclk));
	jdff dff_B_Q9RYIJyk5_1(.din(w_dff_B_ia5XpHfb1_1),.dout(w_dff_B_Q9RYIJyk5_1),.clk(gclk));
	jdff dff_B_zoX5ATlX5_1(.din(w_dff_B_Q9RYIJyk5_1),.dout(w_dff_B_zoX5ATlX5_1),.clk(gclk));
	jdff dff_B_wbM3uAG80_1(.din(w_dff_B_zoX5ATlX5_1),.dout(w_dff_B_wbM3uAG80_1),.clk(gclk));
	jdff dff_B_7Xdc5KDA2_1(.din(w_dff_B_wbM3uAG80_1),.dout(w_dff_B_7Xdc5KDA2_1),.clk(gclk));
	jdff dff_B_eMjTXNVt2_1(.din(w_dff_B_7Xdc5KDA2_1),.dout(w_dff_B_eMjTXNVt2_1),.clk(gclk));
	jdff dff_B_OyvQbfIX6_1(.din(w_dff_B_eMjTXNVt2_1),.dout(w_dff_B_OyvQbfIX6_1),.clk(gclk));
	jdff dff_B_LkLd7c4S5_1(.din(w_dff_B_OyvQbfIX6_1),.dout(w_dff_B_LkLd7c4S5_1),.clk(gclk));
	jdff dff_B_D1JzKo7d1_1(.din(w_dff_B_LkLd7c4S5_1),.dout(w_dff_B_D1JzKo7d1_1),.clk(gclk));
	jdff dff_B_8eNJeAIF6_1(.din(w_dff_B_D1JzKo7d1_1),.dout(w_dff_B_8eNJeAIF6_1),.clk(gclk));
	jdff dff_B_VMsSEPD41_1(.din(w_dff_B_8eNJeAIF6_1),.dout(w_dff_B_VMsSEPD41_1),.clk(gclk));
	jdff dff_B_3V3AGUMO8_1(.din(w_dff_B_VMsSEPD41_1),.dout(w_dff_B_3V3AGUMO8_1),.clk(gclk));
	jdff dff_B_n5zI5kEv0_1(.din(w_dff_B_3V3AGUMO8_1),.dout(w_dff_B_n5zI5kEv0_1),.clk(gclk));
	jdff dff_B_cOFKFadO3_1(.din(w_dff_B_n5zI5kEv0_1),.dout(w_dff_B_cOFKFadO3_1),.clk(gclk));
	jdff dff_B_PwtDI52T9_1(.din(w_dff_B_cOFKFadO3_1),.dout(w_dff_B_PwtDI52T9_1),.clk(gclk));
	jdff dff_B_09g35pyA2_1(.din(w_dff_B_PwtDI52T9_1),.dout(w_dff_B_09g35pyA2_1),.clk(gclk));
	jdff dff_B_FeR02UvE6_1(.din(w_dff_B_09g35pyA2_1),.dout(w_dff_B_FeR02UvE6_1),.clk(gclk));
	jdff dff_B_5kcb8wRv6_1(.din(w_dff_B_FeR02UvE6_1),.dout(w_dff_B_5kcb8wRv6_1),.clk(gclk));
	jdff dff_B_XLby0v3k4_1(.din(w_dff_B_5kcb8wRv6_1),.dout(w_dff_B_XLby0v3k4_1),.clk(gclk));
	jdff dff_B_YIcD3ovG5_1(.din(w_dff_B_XLby0v3k4_1),.dout(w_dff_B_YIcD3ovG5_1),.clk(gclk));
	jdff dff_B_lJ7GpQk82_1(.din(w_dff_B_YIcD3ovG5_1),.dout(w_dff_B_lJ7GpQk82_1),.clk(gclk));
	jdff dff_B_CbZ06e4w7_1(.din(w_dff_B_lJ7GpQk82_1),.dout(w_dff_B_CbZ06e4w7_1),.clk(gclk));
	jdff dff_B_g0qywdFH7_1(.din(w_dff_B_CbZ06e4w7_1),.dout(w_dff_B_g0qywdFH7_1),.clk(gclk));
	jdff dff_B_R7UTxnki4_1(.din(w_dff_B_g0qywdFH7_1),.dout(w_dff_B_R7UTxnki4_1),.clk(gclk));
	jdff dff_B_wri3YED41_1(.din(w_dff_B_R7UTxnki4_1),.dout(w_dff_B_wri3YED41_1),.clk(gclk));
	jdff dff_B_O8bczUst3_1(.din(w_dff_B_wri3YED41_1),.dout(w_dff_B_O8bczUst3_1),.clk(gclk));
	jdff dff_B_38fwY4Ln6_1(.din(w_dff_B_O8bczUst3_1),.dout(w_dff_B_38fwY4Ln6_1),.clk(gclk));
	jdff dff_B_faHhFQx39_1(.din(w_dff_B_38fwY4Ln6_1),.dout(w_dff_B_faHhFQx39_1),.clk(gclk));
	jdff dff_B_rAkmUrHa2_1(.din(w_dff_B_faHhFQx39_1),.dout(w_dff_B_rAkmUrHa2_1),.clk(gclk));
	jdff dff_B_8IY2qjMo0_1(.din(w_dff_B_rAkmUrHa2_1),.dout(w_dff_B_8IY2qjMo0_1),.clk(gclk));
	jdff dff_B_DVsHxG738_1(.din(w_dff_B_8IY2qjMo0_1),.dout(w_dff_B_DVsHxG738_1),.clk(gclk));
	jdff dff_B_Dz1BOvfe3_1(.din(w_dff_B_DVsHxG738_1),.dout(w_dff_B_Dz1BOvfe3_1),.clk(gclk));
	jdff dff_B_2OLArSu79_1(.din(w_dff_B_Dz1BOvfe3_1),.dout(w_dff_B_2OLArSu79_1),.clk(gclk));
	jdff dff_B_uvEgy2uw2_1(.din(w_dff_B_2OLArSu79_1),.dout(w_dff_B_uvEgy2uw2_1),.clk(gclk));
	jdff dff_B_gFNdgW0F4_1(.din(w_dff_B_uvEgy2uw2_1),.dout(w_dff_B_gFNdgW0F4_1),.clk(gclk));
	jdff dff_B_9iZ9wvN55_1(.din(w_dff_B_gFNdgW0F4_1),.dout(w_dff_B_9iZ9wvN55_1),.clk(gclk));
	jdff dff_B_R04kQDea7_1(.din(w_dff_B_9iZ9wvN55_1),.dout(w_dff_B_R04kQDea7_1),.clk(gclk));
	jdff dff_B_pqpOHVfn2_1(.din(w_dff_B_R04kQDea7_1),.dout(w_dff_B_pqpOHVfn2_1),.clk(gclk));
	jdff dff_B_lbx0bJ3I1_0(.din(n883),.dout(w_dff_B_lbx0bJ3I1_0),.clk(gclk));
	jdff dff_B_UgaUlG2h9_0(.din(w_dff_B_lbx0bJ3I1_0),.dout(w_dff_B_UgaUlG2h9_0),.clk(gclk));
	jdff dff_B_bgm9I2RO3_0(.din(w_dff_B_UgaUlG2h9_0),.dout(w_dff_B_bgm9I2RO3_0),.clk(gclk));
	jdff dff_B_YQcMCGIS2_0(.din(w_dff_B_bgm9I2RO3_0),.dout(w_dff_B_YQcMCGIS2_0),.clk(gclk));
	jdff dff_B_w58wDCjv1_0(.din(w_dff_B_YQcMCGIS2_0),.dout(w_dff_B_w58wDCjv1_0),.clk(gclk));
	jdff dff_B_kywKR1cJ6_0(.din(w_dff_B_w58wDCjv1_0),.dout(w_dff_B_kywKR1cJ6_0),.clk(gclk));
	jdff dff_B_ulUMzjEr8_0(.din(w_dff_B_kywKR1cJ6_0),.dout(w_dff_B_ulUMzjEr8_0),.clk(gclk));
	jdff dff_B_4ZxSj76o7_0(.din(w_dff_B_ulUMzjEr8_0),.dout(w_dff_B_4ZxSj76o7_0),.clk(gclk));
	jdff dff_B_eMYbxtrk4_0(.din(w_dff_B_4ZxSj76o7_0),.dout(w_dff_B_eMYbxtrk4_0),.clk(gclk));
	jdff dff_B_fSm2hHlu7_0(.din(w_dff_B_eMYbxtrk4_0),.dout(w_dff_B_fSm2hHlu7_0),.clk(gclk));
	jdff dff_B_yXjcUZOK0_0(.din(w_dff_B_fSm2hHlu7_0),.dout(w_dff_B_yXjcUZOK0_0),.clk(gclk));
	jdff dff_B_1zLrhq7K1_0(.din(w_dff_B_yXjcUZOK0_0),.dout(w_dff_B_1zLrhq7K1_0),.clk(gclk));
	jdff dff_B_5wjrOJs38_0(.din(w_dff_B_1zLrhq7K1_0),.dout(w_dff_B_5wjrOJs38_0),.clk(gclk));
	jdff dff_B_XMzR0ZiJ0_0(.din(w_dff_B_5wjrOJs38_0),.dout(w_dff_B_XMzR0ZiJ0_0),.clk(gclk));
	jdff dff_B_gPfC5QxC4_0(.din(w_dff_B_XMzR0ZiJ0_0),.dout(w_dff_B_gPfC5QxC4_0),.clk(gclk));
	jdff dff_B_syhuGrkJ1_0(.din(w_dff_B_gPfC5QxC4_0),.dout(w_dff_B_syhuGrkJ1_0),.clk(gclk));
	jdff dff_B_xMp1MZqg5_0(.din(w_dff_B_syhuGrkJ1_0),.dout(w_dff_B_xMp1MZqg5_0),.clk(gclk));
	jdff dff_B_5RpfC5KX3_0(.din(w_dff_B_xMp1MZqg5_0),.dout(w_dff_B_5RpfC5KX3_0),.clk(gclk));
	jdff dff_B_8mrylY1Q0_0(.din(w_dff_B_5RpfC5KX3_0),.dout(w_dff_B_8mrylY1Q0_0),.clk(gclk));
	jdff dff_B_ovHkF9IV0_0(.din(w_dff_B_8mrylY1Q0_0),.dout(w_dff_B_ovHkF9IV0_0),.clk(gclk));
	jdff dff_B_rvcFtqMG9_0(.din(w_dff_B_ovHkF9IV0_0),.dout(w_dff_B_rvcFtqMG9_0),.clk(gclk));
	jdff dff_B_2sfw3t971_0(.din(w_dff_B_rvcFtqMG9_0),.dout(w_dff_B_2sfw3t971_0),.clk(gclk));
	jdff dff_B_rlgkM11P5_0(.din(w_dff_B_2sfw3t971_0),.dout(w_dff_B_rlgkM11P5_0),.clk(gclk));
	jdff dff_B_N7gOJYOh8_0(.din(w_dff_B_rlgkM11P5_0),.dout(w_dff_B_N7gOJYOh8_0),.clk(gclk));
	jdff dff_B_Ipbu9Ot25_0(.din(w_dff_B_N7gOJYOh8_0),.dout(w_dff_B_Ipbu9Ot25_0),.clk(gclk));
	jdff dff_B_wYqg17or3_0(.din(w_dff_B_Ipbu9Ot25_0),.dout(w_dff_B_wYqg17or3_0),.clk(gclk));
	jdff dff_B_52rEqSmP5_0(.din(w_dff_B_wYqg17or3_0),.dout(w_dff_B_52rEqSmP5_0),.clk(gclk));
	jdff dff_B_Y4dLJha30_0(.din(w_dff_B_52rEqSmP5_0),.dout(w_dff_B_Y4dLJha30_0),.clk(gclk));
	jdff dff_B_1dsZkoae8_0(.din(w_dff_B_Y4dLJha30_0),.dout(w_dff_B_1dsZkoae8_0),.clk(gclk));
	jdff dff_B_TAyn4PGm2_0(.din(w_dff_B_1dsZkoae8_0),.dout(w_dff_B_TAyn4PGm2_0),.clk(gclk));
	jdff dff_B_zR8DzHqz5_0(.din(w_dff_B_TAyn4PGm2_0),.dout(w_dff_B_zR8DzHqz5_0),.clk(gclk));
	jdff dff_B_JPxwGHbe9_0(.din(w_dff_B_zR8DzHqz5_0),.dout(w_dff_B_JPxwGHbe9_0),.clk(gclk));
	jdff dff_B_F1bEbhZw3_0(.din(w_dff_B_JPxwGHbe9_0),.dout(w_dff_B_F1bEbhZw3_0),.clk(gclk));
	jdff dff_B_Ovtj5Uu34_0(.din(w_dff_B_F1bEbhZw3_0),.dout(w_dff_B_Ovtj5Uu34_0),.clk(gclk));
	jdff dff_B_mlE9rzgM9_0(.din(w_dff_B_Ovtj5Uu34_0),.dout(w_dff_B_mlE9rzgM9_0),.clk(gclk));
	jdff dff_B_F2dJ8WjC6_0(.din(w_dff_B_mlE9rzgM9_0),.dout(w_dff_B_F2dJ8WjC6_0),.clk(gclk));
	jdff dff_B_LQ3kaRtF8_0(.din(w_dff_B_F2dJ8WjC6_0),.dout(w_dff_B_LQ3kaRtF8_0),.clk(gclk));
	jdff dff_B_Qb5hRfiD2_0(.din(w_dff_B_LQ3kaRtF8_0),.dout(w_dff_B_Qb5hRfiD2_0),.clk(gclk));
	jdff dff_B_luqFBp6l0_0(.din(w_dff_B_Qb5hRfiD2_0),.dout(w_dff_B_luqFBp6l0_0),.clk(gclk));
	jdff dff_B_JSXjiCEQ0_0(.din(w_dff_B_luqFBp6l0_0),.dout(w_dff_B_JSXjiCEQ0_0),.clk(gclk));
	jdff dff_B_nyu6l83o3_0(.din(w_dff_B_JSXjiCEQ0_0),.dout(w_dff_B_nyu6l83o3_0),.clk(gclk));
	jdff dff_B_DUPsTurq4_0(.din(w_dff_B_nyu6l83o3_0),.dout(w_dff_B_DUPsTurq4_0),.clk(gclk));
	jdff dff_B_3J4ZgUEC1_0(.din(w_dff_B_DUPsTurq4_0),.dout(w_dff_B_3J4ZgUEC1_0),.clk(gclk));
	jdff dff_B_1IBbH39q0_0(.din(w_dff_B_3J4ZgUEC1_0),.dout(w_dff_B_1IBbH39q0_0),.clk(gclk));
	jdff dff_B_pn6a7Tt96_0(.din(w_dff_B_1IBbH39q0_0),.dout(w_dff_B_pn6a7Tt96_0),.clk(gclk));
	jdff dff_B_Bbq4SO8H0_0(.din(w_dff_B_pn6a7Tt96_0),.dout(w_dff_B_Bbq4SO8H0_0),.clk(gclk));
	jdff dff_B_ujHpbwvQ9_0(.din(w_dff_B_Bbq4SO8H0_0),.dout(w_dff_B_ujHpbwvQ9_0),.clk(gclk));
	jdff dff_B_TNQBdK2p8_0(.din(w_dff_B_ujHpbwvQ9_0),.dout(w_dff_B_TNQBdK2p8_0),.clk(gclk));
	jdff dff_B_UoMHYi4T2_0(.din(w_dff_B_TNQBdK2p8_0),.dout(w_dff_B_UoMHYi4T2_0),.clk(gclk));
	jdff dff_B_ZVSmNbLf7_0(.din(w_dff_B_UoMHYi4T2_0),.dout(w_dff_B_ZVSmNbLf7_0),.clk(gclk));
	jdff dff_B_49oXdpNJ2_0(.din(w_dff_B_ZVSmNbLf7_0),.dout(w_dff_B_49oXdpNJ2_0),.clk(gclk));
	jdff dff_B_nTfSG4iy3_0(.din(w_dff_B_49oXdpNJ2_0),.dout(w_dff_B_nTfSG4iy3_0),.clk(gclk));
	jdff dff_B_Oy80N22j5_0(.din(w_dff_B_nTfSG4iy3_0),.dout(w_dff_B_Oy80N22j5_0),.clk(gclk));
	jdff dff_B_CHQb8XLy8_0(.din(w_dff_B_Oy80N22j5_0),.dout(w_dff_B_CHQb8XLy8_0),.clk(gclk));
	jdff dff_B_YJkhyArE6_0(.din(w_dff_B_CHQb8XLy8_0),.dout(w_dff_B_YJkhyArE6_0),.clk(gclk));
	jdff dff_B_QAH5LVWN5_0(.din(w_dff_B_YJkhyArE6_0),.dout(w_dff_B_QAH5LVWN5_0),.clk(gclk));
	jdff dff_B_mh4uii889_0(.din(w_dff_B_QAH5LVWN5_0),.dout(w_dff_B_mh4uii889_0),.clk(gclk));
	jdff dff_B_zfdsILgT3_0(.din(w_dff_B_mh4uii889_0),.dout(w_dff_B_zfdsILgT3_0),.clk(gclk));
	jdff dff_B_SzkvICuc8_0(.din(w_dff_B_zfdsILgT3_0),.dout(w_dff_B_SzkvICuc8_0),.clk(gclk));
	jdff dff_B_uqsLirJX5_0(.din(w_dff_B_SzkvICuc8_0),.dout(w_dff_B_uqsLirJX5_0),.clk(gclk));
	jdff dff_B_uskQaVMn5_0(.din(w_dff_B_uqsLirJX5_0),.dout(w_dff_B_uskQaVMn5_0),.clk(gclk));
	jdff dff_B_BHZ6k7Y53_0(.din(w_dff_B_uskQaVMn5_0),.dout(w_dff_B_BHZ6k7Y53_0),.clk(gclk));
	jdff dff_B_XH8yS9iD4_0(.din(w_dff_B_BHZ6k7Y53_0),.dout(w_dff_B_XH8yS9iD4_0),.clk(gclk));
	jdff dff_B_R5zlN7zy5_0(.din(w_dff_B_XH8yS9iD4_0),.dout(w_dff_B_R5zlN7zy5_0),.clk(gclk));
	jdff dff_B_V8anR2zM2_0(.din(w_dff_B_R5zlN7zy5_0),.dout(w_dff_B_V8anR2zM2_0),.clk(gclk));
	jdff dff_B_ETi7pgUl8_0(.din(w_dff_B_V8anR2zM2_0),.dout(w_dff_B_ETi7pgUl8_0),.clk(gclk));
	jdff dff_B_lVz8UHwx9_0(.din(w_dff_B_ETi7pgUl8_0),.dout(w_dff_B_lVz8UHwx9_0),.clk(gclk));
	jdff dff_B_KvRRpVXS0_0(.din(w_dff_B_lVz8UHwx9_0),.dout(w_dff_B_KvRRpVXS0_0),.clk(gclk));
	jdff dff_B_wPXMR1n72_0(.din(w_dff_B_KvRRpVXS0_0),.dout(w_dff_B_wPXMR1n72_0),.clk(gclk));
	jdff dff_B_RgdBGlg80_0(.din(w_dff_B_wPXMR1n72_0),.dout(w_dff_B_RgdBGlg80_0),.clk(gclk));
	jdff dff_B_dCaPC60s2_0(.din(w_dff_B_RgdBGlg80_0),.dout(w_dff_B_dCaPC60s2_0),.clk(gclk));
	jdff dff_B_zftcPdEp8_0(.din(w_dff_B_dCaPC60s2_0),.dout(w_dff_B_zftcPdEp8_0),.clk(gclk));
	jdff dff_B_3UL5uNh81_0(.din(w_dff_B_zftcPdEp8_0),.dout(w_dff_B_3UL5uNh81_0),.clk(gclk));
	jdff dff_B_XBqXH6D92_0(.din(w_dff_B_3UL5uNh81_0),.dout(w_dff_B_XBqXH6D92_0),.clk(gclk));
	jdff dff_B_QmfgcSuP6_0(.din(w_dff_B_XBqXH6D92_0),.dout(w_dff_B_QmfgcSuP6_0),.clk(gclk));
	jdff dff_B_tNRYvELa2_0(.din(w_dff_B_QmfgcSuP6_0),.dout(w_dff_B_tNRYvELa2_0),.clk(gclk));
	jdff dff_B_QGUwBrrA3_0(.din(w_dff_B_tNRYvELa2_0),.dout(w_dff_B_QGUwBrrA3_0),.clk(gclk));
	jdff dff_B_vOhWD8ma3_0(.din(w_dff_B_QGUwBrrA3_0),.dout(w_dff_B_vOhWD8ma3_0),.clk(gclk));
	jdff dff_B_fNLVoglA7_0(.din(w_dff_B_vOhWD8ma3_0),.dout(w_dff_B_fNLVoglA7_0),.clk(gclk));
	jdff dff_B_oeLcs5Fp4_0(.din(w_dff_B_fNLVoglA7_0),.dout(w_dff_B_oeLcs5Fp4_0),.clk(gclk));
	jdff dff_B_v73dFm1n7_0(.din(w_dff_B_oeLcs5Fp4_0),.dout(w_dff_B_v73dFm1n7_0),.clk(gclk));
	jdff dff_B_AtsoBtob9_0(.din(w_dff_B_v73dFm1n7_0),.dout(w_dff_B_AtsoBtob9_0),.clk(gclk));
	jdff dff_B_XuAALr0W2_0(.din(w_dff_B_AtsoBtob9_0),.dout(w_dff_B_XuAALr0W2_0),.clk(gclk));
	jdff dff_B_Xd3qesh12_1(.din(n876),.dout(w_dff_B_Xd3qesh12_1),.clk(gclk));
	jdff dff_B_Eokc923Z1_1(.din(w_dff_B_Xd3qesh12_1),.dout(w_dff_B_Eokc923Z1_1),.clk(gclk));
	jdff dff_B_oAHzyOSn4_1(.din(w_dff_B_Eokc923Z1_1),.dout(w_dff_B_oAHzyOSn4_1),.clk(gclk));
	jdff dff_B_ICP5pvP52_1(.din(w_dff_B_oAHzyOSn4_1),.dout(w_dff_B_ICP5pvP52_1),.clk(gclk));
	jdff dff_B_QXMlNoS57_1(.din(w_dff_B_ICP5pvP52_1),.dout(w_dff_B_QXMlNoS57_1),.clk(gclk));
	jdff dff_B_HhcMAKUO9_1(.din(w_dff_B_QXMlNoS57_1),.dout(w_dff_B_HhcMAKUO9_1),.clk(gclk));
	jdff dff_B_z2dU9mrH0_1(.din(w_dff_B_HhcMAKUO9_1),.dout(w_dff_B_z2dU9mrH0_1),.clk(gclk));
	jdff dff_B_DTG1yr730_1(.din(w_dff_B_z2dU9mrH0_1),.dout(w_dff_B_DTG1yr730_1),.clk(gclk));
	jdff dff_B_kPYFWJQU5_1(.din(w_dff_B_DTG1yr730_1),.dout(w_dff_B_kPYFWJQU5_1),.clk(gclk));
	jdff dff_B_eldJobIu1_1(.din(w_dff_B_kPYFWJQU5_1),.dout(w_dff_B_eldJobIu1_1),.clk(gclk));
	jdff dff_B_seIxoZZz2_1(.din(w_dff_B_eldJobIu1_1),.dout(w_dff_B_seIxoZZz2_1),.clk(gclk));
	jdff dff_B_L1ssJrKX0_1(.din(w_dff_B_seIxoZZz2_1),.dout(w_dff_B_L1ssJrKX0_1),.clk(gclk));
	jdff dff_B_zjULwgap5_1(.din(w_dff_B_L1ssJrKX0_1),.dout(w_dff_B_zjULwgap5_1),.clk(gclk));
	jdff dff_B_1gm5Ydf39_1(.din(w_dff_B_zjULwgap5_1),.dout(w_dff_B_1gm5Ydf39_1),.clk(gclk));
	jdff dff_B_8eSX5zWY4_1(.din(w_dff_B_1gm5Ydf39_1),.dout(w_dff_B_8eSX5zWY4_1),.clk(gclk));
	jdff dff_B_DFHIWMFM8_1(.din(w_dff_B_8eSX5zWY4_1),.dout(w_dff_B_DFHIWMFM8_1),.clk(gclk));
	jdff dff_B_oXXmaJfU7_1(.din(w_dff_B_DFHIWMFM8_1),.dout(w_dff_B_oXXmaJfU7_1),.clk(gclk));
	jdff dff_B_E88Fkyhd9_1(.din(w_dff_B_oXXmaJfU7_1),.dout(w_dff_B_E88Fkyhd9_1),.clk(gclk));
	jdff dff_B_sGUqVLio2_1(.din(w_dff_B_E88Fkyhd9_1),.dout(w_dff_B_sGUqVLio2_1),.clk(gclk));
	jdff dff_B_9uUW4FKq6_1(.din(w_dff_B_sGUqVLio2_1),.dout(w_dff_B_9uUW4FKq6_1),.clk(gclk));
	jdff dff_B_cApTODzx3_1(.din(w_dff_B_9uUW4FKq6_1),.dout(w_dff_B_cApTODzx3_1),.clk(gclk));
	jdff dff_B_u9Y1Kk1M2_1(.din(w_dff_B_cApTODzx3_1),.dout(w_dff_B_u9Y1Kk1M2_1),.clk(gclk));
	jdff dff_B_yzvPv0Gf2_1(.din(w_dff_B_u9Y1Kk1M2_1),.dout(w_dff_B_yzvPv0Gf2_1),.clk(gclk));
	jdff dff_B_e277gc5k7_1(.din(w_dff_B_yzvPv0Gf2_1),.dout(w_dff_B_e277gc5k7_1),.clk(gclk));
	jdff dff_B_5yP6dijU2_1(.din(w_dff_B_e277gc5k7_1),.dout(w_dff_B_5yP6dijU2_1),.clk(gclk));
	jdff dff_B_syBHCo5S8_1(.din(w_dff_B_5yP6dijU2_1),.dout(w_dff_B_syBHCo5S8_1),.clk(gclk));
	jdff dff_B_s6tREeMO8_1(.din(w_dff_B_syBHCo5S8_1),.dout(w_dff_B_s6tREeMO8_1),.clk(gclk));
	jdff dff_B_RnLjzHSX0_1(.din(w_dff_B_s6tREeMO8_1),.dout(w_dff_B_RnLjzHSX0_1),.clk(gclk));
	jdff dff_B_eCalJcio6_1(.din(w_dff_B_RnLjzHSX0_1),.dout(w_dff_B_eCalJcio6_1),.clk(gclk));
	jdff dff_B_ksb7gZyq3_1(.din(w_dff_B_eCalJcio6_1),.dout(w_dff_B_ksb7gZyq3_1),.clk(gclk));
	jdff dff_B_9qaNjVeX6_1(.din(w_dff_B_ksb7gZyq3_1),.dout(w_dff_B_9qaNjVeX6_1),.clk(gclk));
	jdff dff_B_O8bgULBf5_1(.din(w_dff_B_9qaNjVeX6_1),.dout(w_dff_B_O8bgULBf5_1),.clk(gclk));
	jdff dff_B_qY474FcQ6_1(.din(w_dff_B_O8bgULBf5_1),.dout(w_dff_B_qY474FcQ6_1),.clk(gclk));
	jdff dff_B_CFFeTcxm3_1(.din(w_dff_B_qY474FcQ6_1),.dout(w_dff_B_CFFeTcxm3_1),.clk(gclk));
	jdff dff_B_399lFJV69_1(.din(w_dff_B_CFFeTcxm3_1),.dout(w_dff_B_399lFJV69_1),.clk(gclk));
	jdff dff_B_53UHsDp51_1(.din(w_dff_B_399lFJV69_1),.dout(w_dff_B_53UHsDp51_1),.clk(gclk));
	jdff dff_B_tYs46H4D0_1(.din(w_dff_B_53UHsDp51_1),.dout(w_dff_B_tYs46H4D0_1),.clk(gclk));
	jdff dff_B_rt75IlMh2_1(.din(w_dff_B_tYs46H4D0_1),.dout(w_dff_B_rt75IlMh2_1),.clk(gclk));
	jdff dff_B_2O0ggyf76_1(.din(w_dff_B_rt75IlMh2_1),.dout(w_dff_B_2O0ggyf76_1),.clk(gclk));
	jdff dff_B_0o1vNFXX9_1(.din(w_dff_B_2O0ggyf76_1),.dout(w_dff_B_0o1vNFXX9_1),.clk(gclk));
	jdff dff_B_5rKo3sG89_1(.din(w_dff_B_0o1vNFXX9_1),.dout(w_dff_B_5rKo3sG89_1),.clk(gclk));
	jdff dff_B_YRGyUjuk0_1(.din(w_dff_B_5rKo3sG89_1),.dout(w_dff_B_YRGyUjuk0_1),.clk(gclk));
	jdff dff_B_doE5mHOh9_1(.din(w_dff_B_YRGyUjuk0_1),.dout(w_dff_B_doE5mHOh9_1),.clk(gclk));
	jdff dff_B_fmMw772B1_1(.din(w_dff_B_doE5mHOh9_1),.dout(w_dff_B_fmMw772B1_1),.clk(gclk));
	jdff dff_B_KvZawl2d8_1(.din(w_dff_B_fmMw772B1_1),.dout(w_dff_B_KvZawl2d8_1),.clk(gclk));
	jdff dff_B_u9Yjhk0a5_1(.din(w_dff_B_KvZawl2d8_1),.dout(w_dff_B_u9Yjhk0a5_1),.clk(gclk));
	jdff dff_B_kgyJzPCJ1_1(.din(w_dff_B_u9Yjhk0a5_1),.dout(w_dff_B_kgyJzPCJ1_1),.clk(gclk));
	jdff dff_B_O1FazG0M5_1(.din(w_dff_B_kgyJzPCJ1_1),.dout(w_dff_B_O1FazG0M5_1),.clk(gclk));
	jdff dff_B_w4H1VIdU4_1(.din(w_dff_B_O1FazG0M5_1),.dout(w_dff_B_w4H1VIdU4_1),.clk(gclk));
	jdff dff_B_774dSw5z2_1(.din(w_dff_B_w4H1VIdU4_1),.dout(w_dff_B_774dSw5z2_1),.clk(gclk));
	jdff dff_B_lMaWDzSI2_1(.din(w_dff_B_774dSw5z2_1),.dout(w_dff_B_lMaWDzSI2_1),.clk(gclk));
	jdff dff_B_y6CplWrf0_1(.din(w_dff_B_lMaWDzSI2_1),.dout(w_dff_B_y6CplWrf0_1),.clk(gclk));
	jdff dff_B_bnYHiXBW9_1(.din(w_dff_B_y6CplWrf0_1),.dout(w_dff_B_bnYHiXBW9_1),.clk(gclk));
	jdff dff_B_3kQGj0Cf9_1(.din(w_dff_B_bnYHiXBW9_1),.dout(w_dff_B_3kQGj0Cf9_1),.clk(gclk));
	jdff dff_B_2WtXukM07_1(.din(w_dff_B_3kQGj0Cf9_1),.dout(w_dff_B_2WtXukM07_1),.clk(gclk));
	jdff dff_B_sSUNASYl8_1(.din(w_dff_B_2WtXukM07_1),.dout(w_dff_B_sSUNASYl8_1),.clk(gclk));
	jdff dff_B_zveSQgSV5_1(.din(w_dff_B_sSUNASYl8_1),.dout(w_dff_B_zveSQgSV5_1),.clk(gclk));
	jdff dff_B_b3HkcRC63_1(.din(w_dff_B_zveSQgSV5_1),.dout(w_dff_B_b3HkcRC63_1),.clk(gclk));
	jdff dff_B_DCuFrT1Q1_1(.din(w_dff_B_b3HkcRC63_1),.dout(w_dff_B_DCuFrT1Q1_1),.clk(gclk));
	jdff dff_B_FqulapPz9_1(.din(w_dff_B_DCuFrT1Q1_1),.dout(w_dff_B_FqulapPz9_1),.clk(gclk));
	jdff dff_B_jACIDB1M8_1(.din(w_dff_B_FqulapPz9_1),.dout(w_dff_B_jACIDB1M8_1),.clk(gclk));
	jdff dff_B_PqOy7b1u8_1(.din(w_dff_B_jACIDB1M8_1),.dout(w_dff_B_PqOy7b1u8_1),.clk(gclk));
	jdff dff_B_ef8zidSD8_1(.din(w_dff_B_PqOy7b1u8_1),.dout(w_dff_B_ef8zidSD8_1),.clk(gclk));
	jdff dff_B_ly868IGg7_1(.din(w_dff_B_ef8zidSD8_1),.dout(w_dff_B_ly868IGg7_1),.clk(gclk));
	jdff dff_B_48xh1Xbv7_1(.din(w_dff_B_ly868IGg7_1),.dout(w_dff_B_48xh1Xbv7_1),.clk(gclk));
	jdff dff_B_ENuE0Vz92_1(.din(w_dff_B_48xh1Xbv7_1),.dout(w_dff_B_ENuE0Vz92_1),.clk(gclk));
	jdff dff_B_POWywMl40_1(.din(w_dff_B_ENuE0Vz92_1),.dout(w_dff_B_POWywMl40_1),.clk(gclk));
	jdff dff_B_vImdWakB7_1(.din(w_dff_B_POWywMl40_1),.dout(w_dff_B_vImdWakB7_1),.clk(gclk));
	jdff dff_B_hx1EwlHH6_1(.din(w_dff_B_vImdWakB7_1),.dout(w_dff_B_hx1EwlHH6_1),.clk(gclk));
	jdff dff_B_rdN34DIu8_1(.din(w_dff_B_hx1EwlHH6_1),.dout(w_dff_B_rdN34DIu8_1),.clk(gclk));
	jdff dff_B_AyvGowR26_1(.din(w_dff_B_rdN34DIu8_1),.dout(w_dff_B_AyvGowR26_1),.clk(gclk));
	jdff dff_B_z7cI5L9c8_1(.din(w_dff_B_AyvGowR26_1),.dout(w_dff_B_z7cI5L9c8_1),.clk(gclk));
	jdff dff_B_25t8uufX2_1(.din(w_dff_B_z7cI5L9c8_1),.dout(w_dff_B_25t8uufX2_1),.clk(gclk));
	jdff dff_B_x7ePNm8y5_1(.din(w_dff_B_25t8uufX2_1),.dout(w_dff_B_x7ePNm8y5_1),.clk(gclk));
	jdff dff_B_aUdLdDXa1_1(.din(w_dff_B_x7ePNm8y5_1),.dout(w_dff_B_aUdLdDXa1_1),.clk(gclk));
	jdff dff_B_IjxD3l1I6_1(.din(w_dff_B_aUdLdDXa1_1),.dout(w_dff_B_IjxD3l1I6_1),.clk(gclk));
	jdff dff_B_gisVeJyT4_1(.din(w_dff_B_IjxD3l1I6_1),.dout(w_dff_B_gisVeJyT4_1),.clk(gclk));
	jdff dff_B_9oyZfYz89_1(.din(w_dff_B_gisVeJyT4_1),.dout(w_dff_B_9oyZfYz89_1),.clk(gclk));
	jdff dff_B_PTXz50yE3_1(.din(w_dff_B_9oyZfYz89_1),.dout(w_dff_B_PTXz50yE3_1),.clk(gclk));
	jdff dff_B_PkGbuQfZ3_1(.din(w_dff_B_PTXz50yE3_1),.dout(w_dff_B_PkGbuQfZ3_1),.clk(gclk));
	jdff dff_B_RuSpPh4Y8_1(.din(w_dff_B_PkGbuQfZ3_1),.dout(w_dff_B_RuSpPh4Y8_1),.clk(gclk));
	jdff dff_B_GzgJUVn93_1(.din(w_dff_B_RuSpPh4Y8_1),.dout(w_dff_B_GzgJUVn93_1),.clk(gclk));
	jdff dff_B_XcvAxMVt9_0(.din(n877),.dout(w_dff_B_XcvAxMVt9_0),.clk(gclk));
	jdff dff_B_RpVKE8vT4_0(.din(w_dff_B_XcvAxMVt9_0),.dout(w_dff_B_RpVKE8vT4_0),.clk(gclk));
	jdff dff_B_9vBSIjVw6_0(.din(w_dff_B_RpVKE8vT4_0),.dout(w_dff_B_9vBSIjVw6_0),.clk(gclk));
	jdff dff_B_NRtPG4HM1_0(.din(w_dff_B_9vBSIjVw6_0),.dout(w_dff_B_NRtPG4HM1_0),.clk(gclk));
	jdff dff_B_iTFCQodU7_0(.din(w_dff_B_NRtPG4HM1_0),.dout(w_dff_B_iTFCQodU7_0),.clk(gclk));
	jdff dff_B_eNZRrUkz9_0(.din(w_dff_B_iTFCQodU7_0),.dout(w_dff_B_eNZRrUkz9_0),.clk(gclk));
	jdff dff_B_FNGg0k8D4_0(.din(w_dff_B_eNZRrUkz9_0),.dout(w_dff_B_FNGg0k8D4_0),.clk(gclk));
	jdff dff_B_a50DlNCi9_0(.din(w_dff_B_FNGg0k8D4_0),.dout(w_dff_B_a50DlNCi9_0),.clk(gclk));
	jdff dff_B_bTonFqOW3_0(.din(w_dff_B_a50DlNCi9_0),.dout(w_dff_B_bTonFqOW3_0),.clk(gclk));
	jdff dff_B_b73D48xU6_0(.din(w_dff_B_bTonFqOW3_0),.dout(w_dff_B_b73D48xU6_0),.clk(gclk));
	jdff dff_B_wiavP2YL6_0(.din(w_dff_B_b73D48xU6_0),.dout(w_dff_B_wiavP2YL6_0),.clk(gclk));
	jdff dff_B_xDx47EjO1_0(.din(w_dff_B_wiavP2YL6_0),.dout(w_dff_B_xDx47EjO1_0),.clk(gclk));
	jdff dff_B_t4SJtfgz5_0(.din(w_dff_B_xDx47EjO1_0),.dout(w_dff_B_t4SJtfgz5_0),.clk(gclk));
	jdff dff_B_m8rltR9S8_0(.din(w_dff_B_t4SJtfgz5_0),.dout(w_dff_B_m8rltR9S8_0),.clk(gclk));
	jdff dff_B_FUZynIAS5_0(.din(w_dff_B_m8rltR9S8_0),.dout(w_dff_B_FUZynIAS5_0),.clk(gclk));
	jdff dff_B_SNJC5Cqh2_0(.din(w_dff_B_FUZynIAS5_0),.dout(w_dff_B_SNJC5Cqh2_0),.clk(gclk));
	jdff dff_B_PuTqYIrU5_0(.din(w_dff_B_SNJC5Cqh2_0),.dout(w_dff_B_PuTqYIrU5_0),.clk(gclk));
	jdff dff_B_bswICrJG7_0(.din(w_dff_B_PuTqYIrU5_0),.dout(w_dff_B_bswICrJG7_0),.clk(gclk));
	jdff dff_B_jr1mpQMw5_0(.din(w_dff_B_bswICrJG7_0),.dout(w_dff_B_jr1mpQMw5_0),.clk(gclk));
	jdff dff_B_IpenWHNU5_0(.din(w_dff_B_jr1mpQMw5_0),.dout(w_dff_B_IpenWHNU5_0),.clk(gclk));
	jdff dff_B_T7qsEW3G4_0(.din(w_dff_B_IpenWHNU5_0),.dout(w_dff_B_T7qsEW3G4_0),.clk(gclk));
	jdff dff_B_bVuI5yqA8_0(.din(w_dff_B_T7qsEW3G4_0),.dout(w_dff_B_bVuI5yqA8_0),.clk(gclk));
	jdff dff_B_xJ3iZ2ii1_0(.din(w_dff_B_bVuI5yqA8_0),.dout(w_dff_B_xJ3iZ2ii1_0),.clk(gclk));
	jdff dff_B_rusifKPM8_0(.din(w_dff_B_xJ3iZ2ii1_0),.dout(w_dff_B_rusifKPM8_0),.clk(gclk));
	jdff dff_B_32aZPd3X6_0(.din(w_dff_B_rusifKPM8_0),.dout(w_dff_B_32aZPd3X6_0),.clk(gclk));
	jdff dff_B_L8Cgwdgs0_0(.din(w_dff_B_32aZPd3X6_0),.dout(w_dff_B_L8Cgwdgs0_0),.clk(gclk));
	jdff dff_B_6rAVLAmc7_0(.din(w_dff_B_L8Cgwdgs0_0),.dout(w_dff_B_6rAVLAmc7_0),.clk(gclk));
	jdff dff_B_yg4SBqH26_0(.din(w_dff_B_6rAVLAmc7_0),.dout(w_dff_B_yg4SBqH26_0),.clk(gclk));
	jdff dff_B_6wzUchkh8_0(.din(w_dff_B_yg4SBqH26_0),.dout(w_dff_B_6wzUchkh8_0),.clk(gclk));
	jdff dff_B_XAEVdv4h6_0(.din(w_dff_B_6wzUchkh8_0),.dout(w_dff_B_XAEVdv4h6_0),.clk(gclk));
	jdff dff_B_sseBOyvc7_0(.din(w_dff_B_XAEVdv4h6_0),.dout(w_dff_B_sseBOyvc7_0),.clk(gclk));
	jdff dff_B_GlzUnj512_0(.din(w_dff_B_sseBOyvc7_0),.dout(w_dff_B_GlzUnj512_0),.clk(gclk));
	jdff dff_B_f2oUjk3w3_0(.din(w_dff_B_GlzUnj512_0),.dout(w_dff_B_f2oUjk3w3_0),.clk(gclk));
	jdff dff_B_2zzWnXtA3_0(.din(w_dff_B_f2oUjk3w3_0),.dout(w_dff_B_2zzWnXtA3_0),.clk(gclk));
	jdff dff_B_T2vaAMqJ2_0(.din(w_dff_B_2zzWnXtA3_0),.dout(w_dff_B_T2vaAMqJ2_0),.clk(gclk));
	jdff dff_B_dYNyFugB3_0(.din(w_dff_B_T2vaAMqJ2_0),.dout(w_dff_B_dYNyFugB3_0),.clk(gclk));
	jdff dff_B_XxUQXtJi6_0(.din(w_dff_B_dYNyFugB3_0),.dout(w_dff_B_XxUQXtJi6_0),.clk(gclk));
	jdff dff_B_ptd5B7Z85_0(.din(w_dff_B_XxUQXtJi6_0),.dout(w_dff_B_ptd5B7Z85_0),.clk(gclk));
	jdff dff_B_49ppE5Yu2_0(.din(w_dff_B_ptd5B7Z85_0),.dout(w_dff_B_49ppE5Yu2_0),.clk(gclk));
	jdff dff_B_EIqH16tS9_0(.din(w_dff_B_49ppE5Yu2_0),.dout(w_dff_B_EIqH16tS9_0),.clk(gclk));
	jdff dff_B_s72BTiyB5_0(.din(w_dff_B_EIqH16tS9_0),.dout(w_dff_B_s72BTiyB5_0),.clk(gclk));
	jdff dff_B_IULCqqVL5_0(.din(w_dff_B_s72BTiyB5_0),.dout(w_dff_B_IULCqqVL5_0),.clk(gclk));
	jdff dff_B_OPCZ2pQK8_0(.din(w_dff_B_IULCqqVL5_0),.dout(w_dff_B_OPCZ2pQK8_0),.clk(gclk));
	jdff dff_B_ttK48AQt5_0(.din(w_dff_B_OPCZ2pQK8_0),.dout(w_dff_B_ttK48AQt5_0),.clk(gclk));
	jdff dff_B_yUjJGqob2_0(.din(w_dff_B_ttK48AQt5_0),.dout(w_dff_B_yUjJGqob2_0),.clk(gclk));
	jdff dff_B_a3fZ0Rio8_0(.din(w_dff_B_yUjJGqob2_0),.dout(w_dff_B_a3fZ0Rio8_0),.clk(gclk));
	jdff dff_B_3GhrjSsy0_0(.din(w_dff_B_a3fZ0Rio8_0),.dout(w_dff_B_3GhrjSsy0_0),.clk(gclk));
	jdff dff_B_3i1rE0Li9_0(.din(w_dff_B_3GhrjSsy0_0),.dout(w_dff_B_3i1rE0Li9_0),.clk(gclk));
	jdff dff_B_iz6Tp54D5_0(.din(w_dff_B_3i1rE0Li9_0),.dout(w_dff_B_iz6Tp54D5_0),.clk(gclk));
	jdff dff_B_eDt15EWn3_0(.din(w_dff_B_iz6Tp54D5_0),.dout(w_dff_B_eDt15EWn3_0),.clk(gclk));
	jdff dff_B_QNakKLW77_0(.din(w_dff_B_eDt15EWn3_0),.dout(w_dff_B_QNakKLW77_0),.clk(gclk));
	jdff dff_B_HDVIR3J11_0(.din(w_dff_B_QNakKLW77_0),.dout(w_dff_B_HDVIR3J11_0),.clk(gclk));
	jdff dff_B_UCeS1BTq5_0(.din(w_dff_B_HDVIR3J11_0),.dout(w_dff_B_UCeS1BTq5_0),.clk(gclk));
	jdff dff_B_1GCpW4xq1_0(.din(w_dff_B_UCeS1BTq5_0),.dout(w_dff_B_1GCpW4xq1_0),.clk(gclk));
	jdff dff_B_SCkx9vpA6_0(.din(w_dff_B_1GCpW4xq1_0),.dout(w_dff_B_SCkx9vpA6_0),.clk(gclk));
	jdff dff_B_sUS44pZR7_0(.din(w_dff_B_SCkx9vpA6_0),.dout(w_dff_B_sUS44pZR7_0),.clk(gclk));
	jdff dff_B_Jz3Hz0aB0_0(.din(w_dff_B_sUS44pZR7_0),.dout(w_dff_B_Jz3Hz0aB0_0),.clk(gclk));
	jdff dff_B_HPb3SAhM2_0(.din(w_dff_B_Jz3Hz0aB0_0),.dout(w_dff_B_HPb3SAhM2_0),.clk(gclk));
	jdff dff_B_GCwkzC5l9_0(.din(w_dff_B_HPb3SAhM2_0),.dout(w_dff_B_GCwkzC5l9_0),.clk(gclk));
	jdff dff_B_SSiLXWJO5_0(.din(w_dff_B_GCwkzC5l9_0),.dout(w_dff_B_SSiLXWJO5_0),.clk(gclk));
	jdff dff_B_GSc3vhSl1_0(.din(w_dff_B_SSiLXWJO5_0),.dout(w_dff_B_GSc3vhSl1_0),.clk(gclk));
	jdff dff_B_SzGCLdj83_0(.din(w_dff_B_GSc3vhSl1_0),.dout(w_dff_B_SzGCLdj83_0),.clk(gclk));
	jdff dff_B_ny6XWGds6_0(.din(w_dff_B_SzGCLdj83_0),.dout(w_dff_B_ny6XWGds6_0),.clk(gclk));
	jdff dff_B_cQbPTwoj5_0(.din(w_dff_B_ny6XWGds6_0),.dout(w_dff_B_cQbPTwoj5_0),.clk(gclk));
	jdff dff_B_tKxglLIJ7_0(.din(w_dff_B_cQbPTwoj5_0),.dout(w_dff_B_tKxglLIJ7_0),.clk(gclk));
	jdff dff_B_wDB7Jm120_0(.din(w_dff_B_tKxglLIJ7_0),.dout(w_dff_B_wDB7Jm120_0),.clk(gclk));
	jdff dff_B_JpQ9tElH8_0(.din(w_dff_B_wDB7Jm120_0),.dout(w_dff_B_JpQ9tElH8_0),.clk(gclk));
	jdff dff_B_FSeBSD4l2_0(.din(w_dff_B_JpQ9tElH8_0),.dout(w_dff_B_FSeBSD4l2_0),.clk(gclk));
	jdff dff_B_m2PCLPWI8_0(.din(w_dff_B_FSeBSD4l2_0),.dout(w_dff_B_m2PCLPWI8_0),.clk(gclk));
	jdff dff_B_foavRE1o9_0(.din(w_dff_B_m2PCLPWI8_0),.dout(w_dff_B_foavRE1o9_0),.clk(gclk));
	jdff dff_B_3iAyf6st6_0(.din(w_dff_B_foavRE1o9_0),.dout(w_dff_B_3iAyf6st6_0),.clk(gclk));
	jdff dff_B_x7wKRM273_0(.din(w_dff_B_3iAyf6st6_0),.dout(w_dff_B_x7wKRM273_0),.clk(gclk));
	jdff dff_B_FYwZKf7J8_0(.din(w_dff_B_x7wKRM273_0),.dout(w_dff_B_FYwZKf7J8_0),.clk(gclk));
	jdff dff_B_VgtKyPMi1_0(.din(w_dff_B_FYwZKf7J8_0),.dout(w_dff_B_VgtKyPMi1_0),.clk(gclk));
	jdff dff_B_AL7UwVBw4_0(.din(w_dff_B_VgtKyPMi1_0),.dout(w_dff_B_AL7UwVBw4_0),.clk(gclk));
	jdff dff_B_7KeJblEc5_0(.din(w_dff_B_AL7UwVBw4_0),.dout(w_dff_B_7KeJblEc5_0),.clk(gclk));
	jdff dff_B_DPn3BabI4_0(.din(w_dff_B_7KeJblEc5_0),.dout(w_dff_B_DPn3BabI4_0),.clk(gclk));
	jdff dff_B_JmnLm2Ir4_0(.din(w_dff_B_DPn3BabI4_0),.dout(w_dff_B_JmnLm2Ir4_0),.clk(gclk));
	jdff dff_B_OZ0Y5C9I6_0(.din(w_dff_B_JmnLm2Ir4_0),.dout(w_dff_B_OZ0Y5C9I6_0),.clk(gclk));
	jdff dff_B_urhxRM5H3_0(.din(w_dff_B_OZ0Y5C9I6_0),.dout(w_dff_B_urhxRM5H3_0),.clk(gclk));
	jdff dff_B_HnA7n8nv2_0(.din(w_dff_B_urhxRM5H3_0),.dout(w_dff_B_HnA7n8nv2_0),.clk(gclk));
	jdff dff_B_kq0cFdQ24_0(.din(w_dff_B_HnA7n8nv2_0),.dout(w_dff_B_kq0cFdQ24_0),.clk(gclk));
	jdff dff_B_HGLUILcM4_1(.din(n870),.dout(w_dff_B_HGLUILcM4_1),.clk(gclk));
	jdff dff_B_FAQyOcLZ7_1(.din(w_dff_B_HGLUILcM4_1),.dout(w_dff_B_FAQyOcLZ7_1),.clk(gclk));
	jdff dff_B_ecvuUYPK7_1(.din(w_dff_B_FAQyOcLZ7_1),.dout(w_dff_B_ecvuUYPK7_1),.clk(gclk));
	jdff dff_B_rHN2QkmK2_1(.din(w_dff_B_ecvuUYPK7_1),.dout(w_dff_B_rHN2QkmK2_1),.clk(gclk));
	jdff dff_B_oSpA3vca2_1(.din(w_dff_B_rHN2QkmK2_1),.dout(w_dff_B_oSpA3vca2_1),.clk(gclk));
	jdff dff_B_5ogCHQop0_1(.din(w_dff_B_oSpA3vca2_1),.dout(w_dff_B_5ogCHQop0_1),.clk(gclk));
	jdff dff_B_LLEgP7sp0_1(.din(w_dff_B_5ogCHQop0_1),.dout(w_dff_B_LLEgP7sp0_1),.clk(gclk));
	jdff dff_B_WtEFNwD22_1(.din(w_dff_B_LLEgP7sp0_1),.dout(w_dff_B_WtEFNwD22_1),.clk(gclk));
	jdff dff_B_SdvpqJ9I0_1(.din(w_dff_B_WtEFNwD22_1),.dout(w_dff_B_SdvpqJ9I0_1),.clk(gclk));
	jdff dff_B_kmjw1zPo7_1(.din(w_dff_B_SdvpqJ9I0_1),.dout(w_dff_B_kmjw1zPo7_1),.clk(gclk));
	jdff dff_B_9tJZEBie7_1(.din(w_dff_B_kmjw1zPo7_1),.dout(w_dff_B_9tJZEBie7_1),.clk(gclk));
	jdff dff_B_ZL2b8DO29_1(.din(w_dff_B_9tJZEBie7_1),.dout(w_dff_B_ZL2b8DO29_1),.clk(gclk));
	jdff dff_B_Oytvunn13_1(.din(w_dff_B_ZL2b8DO29_1),.dout(w_dff_B_Oytvunn13_1),.clk(gclk));
	jdff dff_B_bqTIOM818_1(.din(w_dff_B_Oytvunn13_1),.dout(w_dff_B_bqTIOM818_1),.clk(gclk));
	jdff dff_B_zvgoz3Or6_1(.din(w_dff_B_bqTIOM818_1),.dout(w_dff_B_zvgoz3Or6_1),.clk(gclk));
	jdff dff_B_DjlqhmOH2_1(.din(w_dff_B_zvgoz3Or6_1),.dout(w_dff_B_DjlqhmOH2_1),.clk(gclk));
	jdff dff_B_HRPm5ceE0_1(.din(w_dff_B_DjlqhmOH2_1),.dout(w_dff_B_HRPm5ceE0_1),.clk(gclk));
	jdff dff_B_y0e9V7Le4_1(.din(w_dff_B_HRPm5ceE0_1),.dout(w_dff_B_y0e9V7Le4_1),.clk(gclk));
	jdff dff_B_D3sBofnd3_1(.din(w_dff_B_y0e9V7Le4_1),.dout(w_dff_B_D3sBofnd3_1),.clk(gclk));
	jdff dff_B_bIqpzd0J6_1(.din(w_dff_B_D3sBofnd3_1),.dout(w_dff_B_bIqpzd0J6_1),.clk(gclk));
	jdff dff_B_w46QEcus9_1(.din(w_dff_B_bIqpzd0J6_1),.dout(w_dff_B_w46QEcus9_1),.clk(gclk));
	jdff dff_B_VnurZ78S7_1(.din(w_dff_B_w46QEcus9_1),.dout(w_dff_B_VnurZ78S7_1),.clk(gclk));
	jdff dff_B_rvsf82Hy9_1(.din(w_dff_B_VnurZ78S7_1),.dout(w_dff_B_rvsf82Hy9_1),.clk(gclk));
	jdff dff_B_KCY6jKxL8_1(.din(w_dff_B_rvsf82Hy9_1),.dout(w_dff_B_KCY6jKxL8_1),.clk(gclk));
	jdff dff_B_neuIDJ094_1(.din(w_dff_B_KCY6jKxL8_1),.dout(w_dff_B_neuIDJ094_1),.clk(gclk));
	jdff dff_B_LLlnUf0X8_1(.din(w_dff_B_neuIDJ094_1),.dout(w_dff_B_LLlnUf0X8_1),.clk(gclk));
	jdff dff_B_XnIRbzHe1_1(.din(w_dff_B_LLlnUf0X8_1),.dout(w_dff_B_XnIRbzHe1_1),.clk(gclk));
	jdff dff_B_GlfsU0pY0_1(.din(w_dff_B_XnIRbzHe1_1),.dout(w_dff_B_GlfsU0pY0_1),.clk(gclk));
	jdff dff_B_HkvM7tUT2_1(.din(w_dff_B_GlfsU0pY0_1),.dout(w_dff_B_HkvM7tUT2_1),.clk(gclk));
	jdff dff_B_Jc0uU5PP2_1(.din(w_dff_B_HkvM7tUT2_1),.dout(w_dff_B_Jc0uU5PP2_1),.clk(gclk));
	jdff dff_B_t8S2V3MC4_1(.din(w_dff_B_Jc0uU5PP2_1),.dout(w_dff_B_t8S2V3MC4_1),.clk(gclk));
	jdff dff_B_aaEYDhan0_1(.din(w_dff_B_t8S2V3MC4_1),.dout(w_dff_B_aaEYDhan0_1),.clk(gclk));
	jdff dff_B_pPZqv6HN4_1(.din(w_dff_B_aaEYDhan0_1),.dout(w_dff_B_pPZqv6HN4_1),.clk(gclk));
	jdff dff_B_6Q9PEvRh8_1(.din(w_dff_B_pPZqv6HN4_1),.dout(w_dff_B_6Q9PEvRh8_1),.clk(gclk));
	jdff dff_B_zwpm3GUc5_1(.din(w_dff_B_6Q9PEvRh8_1),.dout(w_dff_B_zwpm3GUc5_1),.clk(gclk));
	jdff dff_B_uJWYmW7H4_1(.din(w_dff_B_zwpm3GUc5_1),.dout(w_dff_B_uJWYmW7H4_1),.clk(gclk));
	jdff dff_B_NZk7PCDX8_1(.din(w_dff_B_uJWYmW7H4_1),.dout(w_dff_B_NZk7PCDX8_1),.clk(gclk));
	jdff dff_B_7EzHJnX21_1(.din(w_dff_B_NZk7PCDX8_1),.dout(w_dff_B_7EzHJnX21_1),.clk(gclk));
	jdff dff_B_cqLup7jz7_1(.din(w_dff_B_7EzHJnX21_1),.dout(w_dff_B_cqLup7jz7_1),.clk(gclk));
	jdff dff_B_P6j9Uit05_1(.din(w_dff_B_cqLup7jz7_1),.dout(w_dff_B_P6j9Uit05_1),.clk(gclk));
	jdff dff_B_yjodbsVS4_1(.din(w_dff_B_P6j9Uit05_1),.dout(w_dff_B_yjodbsVS4_1),.clk(gclk));
	jdff dff_B_HJUaiY828_1(.din(w_dff_B_yjodbsVS4_1),.dout(w_dff_B_HJUaiY828_1),.clk(gclk));
	jdff dff_B_qzyPgkD27_1(.din(w_dff_B_HJUaiY828_1),.dout(w_dff_B_qzyPgkD27_1),.clk(gclk));
	jdff dff_B_X0uR2JGV6_1(.din(w_dff_B_qzyPgkD27_1),.dout(w_dff_B_X0uR2JGV6_1),.clk(gclk));
	jdff dff_B_ER3U3fqg6_1(.din(w_dff_B_X0uR2JGV6_1),.dout(w_dff_B_ER3U3fqg6_1),.clk(gclk));
	jdff dff_B_OKF48mbL2_1(.din(w_dff_B_ER3U3fqg6_1),.dout(w_dff_B_OKF48mbL2_1),.clk(gclk));
	jdff dff_B_VthZKeJx5_1(.din(w_dff_B_OKF48mbL2_1),.dout(w_dff_B_VthZKeJx5_1),.clk(gclk));
	jdff dff_B_BZMoRq1H3_1(.din(w_dff_B_VthZKeJx5_1),.dout(w_dff_B_BZMoRq1H3_1),.clk(gclk));
	jdff dff_B_1556L6KT5_1(.din(w_dff_B_BZMoRq1H3_1),.dout(w_dff_B_1556L6KT5_1),.clk(gclk));
	jdff dff_B_rg0cl9838_1(.din(w_dff_B_1556L6KT5_1),.dout(w_dff_B_rg0cl9838_1),.clk(gclk));
	jdff dff_B_Dvmvkiei3_1(.din(w_dff_B_rg0cl9838_1),.dout(w_dff_B_Dvmvkiei3_1),.clk(gclk));
	jdff dff_B_dS5eIGWr2_1(.din(w_dff_B_Dvmvkiei3_1),.dout(w_dff_B_dS5eIGWr2_1),.clk(gclk));
	jdff dff_B_G9zIIImv0_1(.din(w_dff_B_dS5eIGWr2_1),.dout(w_dff_B_G9zIIImv0_1),.clk(gclk));
	jdff dff_B_7ka1G4sx6_1(.din(w_dff_B_G9zIIImv0_1),.dout(w_dff_B_7ka1G4sx6_1),.clk(gclk));
	jdff dff_B_KWT6pzHw7_1(.din(w_dff_B_7ka1G4sx6_1),.dout(w_dff_B_KWT6pzHw7_1),.clk(gclk));
	jdff dff_B_VpeHMeY28_1(.din(w_dff_B_KWT6pzHw7_1),.dout(w_dff_B_VpeHMeY28_1),.clk(gclk));
	jdff dff_B_IXZHpsWX0_1(.din(w_dff_B_VpeHMeY28_1),.dout(w_dff_B_IXZHpsWX0_1),.clk(gclk));
	jdff dff_B_XMZThkG69_1(.din(w_dff_B_IXZHpsWX0_1),.dout(w_dff_B_XMZThkG69_1),.clk(gclk));
	jdff dff_B_OJU6tlcr3_1(.din(w_dff_B_XMZThkG69_1),.dout(w_dff_B_OJU6tlcr3_1),.clk(gclk));
	jdff dff_B_2FY1RBD26_1(.din(w_dff_B_OJU6tlcr3_1),.dout(w_dff_B_2FY1RBD26_1),.clk(gclk));
	jdff dff_B_XUKOerNr6_1(.din(w_dff_B_2FY1RBD26_1),.dout(w_dff_B_XUKOerNr6_1),.clk(gclk));
	jdff dff_B_cSjM4ZjR3_1(.din(w_dff_B_XUKOerNr6_1),.dout(w_dff_B_cSjM4ZjR3_1),.clk(gclk));
	jdff dff_B_xiwPHwZO0_1(.din(w_dff_B_cSjM4ZjR3_1),.dout(w_dff_B_xiwPHwZO0_1),.clk(gclk));
	jdff dff_B_rmy2HHye7_1(.din(w_dff_B_xiwPHwZO0_1),.dout(w_dff_B_rmy2HHye7_1),.clk(gclk));
	jdff dff_B_4A1CkX5B4_1(.din(w_dff_B_rmy2HHye7_1),.dout(w_dff_B_4A1CkX5B4_1),.clk(gclk));
	jdff dff_B_vbbWAHtj0_1(.din(w_dff_B_4A1CkX5B4_1),.dout(w_dff_B_vbbWAHtj0_1),.clk(gclk));
	jdff dff_B_smF1nojO0_1(.din(w_dff_B_vbbWAHtj0_1),.dout(w_dff_B_smF1nojO0_1),.clk(gclk));
	jdff dff_B_57FFLbto4_1(.din(w_dff_B_smF1nojO0_1),.dout(w_dff_B_57FFLbto4_1),.clk(gclk));
	jdff dff_B_C2Y1m1Yv7_1(.din(w_dff_B_57FFLbto4_1),.dout(w_dff_B_C2Y1m1Yv7_1),.clk(gclk));
	jdff dff_B_wtrTuE9s1_1(.din(w_dff_B_C2Y1m1Yv7_1),.dout(w_dff_B_wtrTuE9s1_1),.clk(gclk));
	jdff dff_B_7V0Zc7gS5_1(.din(w_dff_B_wtrTuE9s1_1),.dout(w_dff_B_7V0Zc7gS5_1),.clk(gclk));
	jdff dff_B_fRWjVBnI8_1(.din(w_dff_B_7V0Zc7gS5_1),.dout(w_dff_B_fRWjVBnI8_1),.clk(gclk));
	jdff dff_B_svFv9JXO5_1(.din(w_dff_B_fRWjVBnI8_1),.dout(w_dff_B_svFv9JXO5_1),.clk(gclk));
	jdff dff_B_UIKRhfJj1_1(.din(w_dff_B_svFv9JXO5_1),.dout(w_dff_B_UIKRhfJj1_1),.clk(gclk));
	jdff dff_B_lfWYUkE89_1(.din(w_dff_B_UIKRhfJj1_1),.dout(w_dff_B_lfWYUkE89_1),.clk(gclk));
	jdff dff_B_jz0eAxfA5_1(.din(w_dff_B_lfWYUkE89_1),.dout(w_dff_B_jz0eAxfA5_1),.clk(gclk));
	jdff dff_B_p5Y4LAwZ6_1(.din(w_dff_B_jz0eAxfA5_1),.dout(w_dff_B_p5Y4LAwZ6_1),.clk(gclk));
	jdff dff_B_4ZXn5FRc7_1(.din(w_dff_B_p5Y4LAwZ6_1),.dout(w_dff_B_4ZXn5FRc7_1),.clk(gclk));
	jdff dff_B_fNWVTgnR3_1(.din(w_dff_B_4ZXn5FRc7_1),.dout(w_dff_B_fNWVTgnR3_1),.clk(gclk));
	jdff dff_B_yXHeBq5g7_1(.din(w_dff_B_fNWVTgnR3_1),.dout(w_dff_B_yXHeBq5g7_1),.clk(gclk));
	jdff dff_B_tvjawTBP1_1(.din(w_dff_B_yXHeBq5g7_1),.dout(w_dff_B_tvjawTBP1_1),.clk(gclk));
	jdff dff_B_G5qkCL0X7_0(.din(n871),.dout(w_dff_B_G5qkCL0X7_0),.clk(gclk));
	jdff dff_B_W0Qjtbz47_0(.din(w_dff_B_G5qkCL0X7_0),.dout(w_dff_B_W0Qjtbz47_0),.clk(gclk));
	jdff dff_B_FrTXzQKt6_0(.din(w_dff_B_W0Qjtbz47_0),.dout(w_dff_B_FrTXzQKt6_0),.clk(gclk));
	jdff dff_B_85UZipWH4_0(.din(w_dff_B_FrTXzQKt6_0),.dout(w_dff_B_85UZipWH4_0),.clk(gclk));
	jdff dff_B_Qwhn3Ko87_0(.din(w_dff_B_85UZipWH4_0),.dout(w_dff_B_Qwhn3Ko87_0),.clk(gclk));
	jdff dff_B_cKlewMrP2_0(.din(w_dff_B_Qwhn3Ko87_0),.dout(w_dff_B_cKlewMrP2_0),.clk(gclk));
	jdff dff_B_LjzyfdRH7_0(.din(w_dff_B_cKlewMrP2_0),.dout(w_dff_B_LjzyfdRH7_0),.clk(gclk));
	jdff dff_B_ZXyzgNCw8_0(.din(w_dff_B_LjzyfdRH7_0),.dout(w_dff_B_ZXyzgNCw8_0),.clk(gclk));
	jdff dff_B_6uLSzrLn5_0(.din(w_dff_B_ZXyzgNCw8_0),.dout(w_dff_B_6uLSzrLn5_0),.clk(gclk));
	jdff dff_B_Sr54sdTA5_0(.din(w_dff_B_6uLSzrLn5_0),.dout(w_dff_B_Sr54sdTA5_0),.clk(gclk));
	jdff dff_B_AyMcy5ei3_0(.din(w_dff_B_Sr54sdTA5_0),.dout(w_dff_B_AyMcy5ei3_0),.clk(gclk));
	jdff dff_B_JLvX7JJU4_0(.din(w_dff_B_AyMcy5ei3_0),.dout(w_dff_B_JLvX7JJU4_0),.clk(gclk));
	jdff dff_B_bBz64bGA2_0(.din(w_dff_B_JLvX7JJU4_0),.dout(w_dff_B_bBz64bGA2_0),.clk(gclk));
	jdff dff_B_pKhh7Bse3_0(.din(w_dff_B_bBz64bGA2_0),.dout(w_dff_B_pKhh7Bse3_0),.clk(gclk));
	jdff dff_B_QMFevvUf8_0(.din(w_dff_B_pKhh7Bse3_0),.dout(w_dff_B_QMFevvUf8_0),.clk(gclk));
	jdff dff_B_ixUx4s6R0_0(.din(w_dff_B_QMFevvUf8_0),.dout(w_dff_B_ixUx4s6R0_0),.clk(gclk));
	jdff dff_B_e4ioJ66S3_0(.din(w_dff_B_ixUx4s6R0_0),.dout(w_dff_B_e4ioJ66S3_0),.clk(gclk));
	jdff dff_B_mcwjGYuR6_0(.din(w_dff_B_e4ioJ66S3_0),.dout(w_dff_B_mcwjGYuR6_0),.clk(gclk));
	jdff dff_B_W2uRE0Cp8_0(.din(w_dff_B_mcwjGYuR6_0),.dout(w_dff_B_W2uRE0Cp8_0),.clk(gclk));
	jdff dff_B_e3df2hCj1_0(.din(w_dff_B_W2uRE0Cp8_0),.dout(w_dff_B_e3df2hCj1_0),.clk(gclk));
	jdff dff_B_WWMhl39V7_0(.din(w_dff_B_e3df2hCj1_0),.dout(w_dff_B_WWMhl39V7_0),.clk(gclk));
	jdff dff_B_KuPQB4Se4_0(.din(w_dff_B_WWMhl39V7_0),.dout(w_dff_B_KuPQB4Se4_0),.clk(gclk));
	jdff dff_B_cCXIpIxk5_0(.din(w_dff_B_KuPQB4Se4_0),.dout(w_dff_B_cCXIpIxk5_0),.clk(gclk));
	jdff dff_B_j3AMZp8F3_0(.din(w_dff_B_cCXIpIxk5_0),.dout(w_dff_B_j3AMZp8F3_0),.clk(gclk));
	jdff dff_B_Qy23gWSG3_0(.din(w_dff_B_j3AMZp8F3_0),.dout(w_dff_B_Qy23gWSG3_0),.clk(gclk));
	jdff dff_B_8ZKhRNLZ9_0(.din(w_dff_B_Qy23gWSG3_0),.dout(w_dff_B_8ZKhRNLZ9_0),.clk(gclk));
	jdff dff_B_2IFjmLoA3_0(.din(w_dff_B_8ZKhRNLZ9_0),.dout(w_dff_B_2IFjmLoA3_0),.clk(gclk));
	jdff dff_B_HWP9ru513_0(.din(w_dff_B_2IFjmLoA3_0),.dout(w_dff_B_HWP9ru513_0),.clk(gclk));
	jdff dff_B_0CdQbKA81_0(.din(w_dff_B_HWP9ru513_0),.dout(w_dff_B_0CdQbKA81_0),.clk(gclk));
	jdff dff_B_tHPKEO575_0(.din(w_dff_B_0CdQbKA81_0),.dout(w_dff_B_tHPKEO575_0),.clk(gclk));
	jdff dff_B_snBOq5kJ0_0(.din(w_dff_B_tHPKEO575_0),.dout(w_dff_B_snBOq5kJ0_0),.clk(gclk));
	jdff dff_B_oTZTnS232_0(.din(w_dff_B_snBOq5kJ0_0),.dout(w_dff_B_oTZTnS232_0),.clk(gclk));
	jdff dff_B_lAezKzTq6_0(.din(w_dff_B_oTZTnS232_0),.dout(w_dff_B_lAezKzTq6_0),.clk(gclk));
	jdff dff_B_pQvZFp9X9_0(.din(w_dff_B_lAezKzTq6_0),.dout(w_dff_B_pQvZFp9X9_0),.clk(gclk));
	jdff dff_B_yqLXZtf07_0(.din(w_dff_B_pQvZFp9X9_0),.dout(w_dff_B_yqLXZtf07_0),.clk(gclk));
	jdff dff_B_fhzR3x2f4_0(.din(w_dff_B_yqLXZtf07_0),.dout(w_dff_B_fhzR3x2f4_0),.clk(gclk));
	jdff dff_B_PZZ92WMf6_0(.din(w_dff_B_fhzR3x2f4_0),.dout(w_dff_B_PZZ92WMf6_0),.clk(gclk));
	jdff dff_B_xV5VhJBE8_0(.din(w_dff_B_PZZ92WMf6_0),.dout(w_dff_B_xV5VhJBE8_0),.clk(gclk));
	jdff dff_B_udSN2HBo6_0(.din(w_dff_B_xV5VhJBE8_0),.dout(w_dff_B_udSN2HBo6_0),.clk(gclk));
	jdff dff_B_UznRq11J3_0(.din(w_dff_B_udSN2HBo6_0),.dout(w_dff_B_UznRq11J3_0),.clk(gclk));
	jdff dff_B_UwRvC1K20_0(.din(w_dff_B_UznRq11J3_0),.dout(w_dff_B_UwRvC1K20_0),.clk(gclk));
	jdff dff_B_E6zqEYfG2_0(.din(w_dff_B_UwRvC1K20_0),.dout(w_dff_B_E6zqEYfG2_0),.clk(gclk));
	jdff dff_B_vAcTpdOW4_0(.din(w_dff_B_E6zqEYfG2_0),.dout(w_dff_B_vAcTpdOW4_0),.clk(gclk));
	jdff dff_B_pdYnTYPI3_0(.din(w_dff_B_vAcTpdOW4_0),.dout(w_dff_B_pdYnTYPI3_0),.clk(gclk));
	jdff dff_B_4NhGbutW7_0(.din(w_dff_B_pdYnTYPI3_0),.dout(w_dff_B_4NhGbutW7_0),.clk(gclk));
	jdff dff_B_xKT1u53Y9_0(.din(w_dff_B_4NhGbutW7_0),.dout(w_dff_B_xKT1u53Y9_0),.clk(gclk));
	jdff dff_B_bgmYoS3D8_0(.din(w_dff_B_xKT1u53Y9_0),.dout(w_dff_B_bgmYoS3D8_0),.clk(gclk));
	jdff dff_B_K9nWt2Yx3_0(.din(w_dff_B_bgmYoS3D8_0),.dout(w_dff_B_K9nWt2Yx3_0),.clk(gclk));
	jdff dff_B_zzyP0Zp78_0(.din(w_dff_B_K9nWt2Yx3_0),.dout(w_dff_B_zzyP0Zp78_0),.clk(gclk));
	jdff dff_B_Izliwfpz0_0(.din(w_dff_B_zzyP0Zp78_0),.dout(w_dff_B_Izliwfpz0_0),.clk(gclk));
	jdff dff_B_s2TekWhD5_0(.din(w_dff_B_Izliwfpz0_0),.dout(w_dff_B_s2TekWhD5_0),.clk(gclk));
	jdff dff_B_zucnam1y8_0(.din(w_dff_B_s2TekWhD5_0),.dout(w_dff_B_zucnam1y8_0),.clk(gclk));
	jdff dff_B_7zs0lD3d3_0(.din(w_dff_B_zucnam1y8_0),.dout(w_dff_B_7zs0lD3d3_0),.clk(gclk));
	jdff dff_B_fU7zMoX06_0(.din(w_dff_B_7zs0lD3d3_0),.dout(w_dff_B_fU7zMoX06_0),.clk(gclk));
	jdff dff_B_ql6LDvXf6_0(.din(w_dff_B_fU7zMoX06_0),.dout(w_dff_B_ql6LDvXf6_0),.clk(gclk));
	jdff dff_B_G3bu3MRX2_0(.din(w_dff_B_ql6LDvXf6_0),.dout(w_dff_B_G3bu3MRX2_0),.clk(gclk));
	jdff dff_B_VCVnfmzm3_0(.din(w_dff_B_G3bu3MRX2_0),.dout(w_dff_B_VCVnfmzm3_0),.clk(gclk));
	jdff dff_B_TPK0c9xf2_0(.din(w_dff_B_VCVnfmzm3_0),.dout(w_dff_B_TPK0c9xf2_0),.clk(gclk));
	jdff dff_B_nlsQP6292_0(.din(w_dff_B_TPK0c9xf2_0),.dout(w_dff_B_nlsQP6292_0),.clk(gclk));
	jdff dff_B_WAmrd0AY3_0(.din(w_dff_B_nlsQP6292_0),.dout(w_dff_B_WAmrd0AY3_0),.clk(gclk));
	jdff dff_B_vVMEnPU32_0(.din(w_dff_B_WAmrd0AY3_0),.dout(w_dff_B_vVMEnPU32_0),.clk(gclk));
	jdff dff_B_xQkZ1Kwc9_0(.din(w_dff_B_vVMEnPU32_0),.dout(w_dff_B_xQkZ1Kwc9_0),.clk(gclk));
	jdff dff_B_CnnuCVmE3_0(.din(w_dff_B_xQkZ1Kwc9_0),.dout(w_dff_B_CnnuCVmE3_0),.clk(gclk));
	jdff dff_B_bCsX3cDJ5_0(.din(w_dff_B_CnnuCVmE3_0),.dout(w_dff_B_bCsX3cDJ5_0),.clk(gclk));
	jdff dff_B_41grjv8w0_0(.din(w_dff_B_bCsX3cDJ5_0),.dout(w_dff_B_41grjv8w0_0),.clk(gclk));
	jdff dff_B_cudNGoO26_0(.din(w_dff_B_41grjv8w0_0),.dout(w_dff_B_cudNGoO26_0),.clk(gclk));
	jdff dff_B_chimribU5_0(.din(w_dff_B_cudNGoO26_0),.dout(w_dff_B_chimribU5_0),.clk(gclk));
	jdff dff_B_UHzd7LdG8_0(.din(w_dff_B_chimribU5_0),.dout(w_dff_B_UHzd7LdG8_0),.clk(gclk));
	jdff dff_B_3wWRXdiY2_0(.din(w_dff_B_UHzd7LdG8_0),.dout(w_dff_B_3wWRXdiY2_0),.clk(gclk));
	jdff dff_B_xbj2Qh1V4_0(.din(w_dff_B_3wWRXdiY2_0),.dout(w_dff_B_xbj2Qh1V4_0),.clk(gclk));
	jdff dff_B_UnoDeeOr7_0(.din(w_dff_B_xbj2Qh1V4_0),.dout(w_dff_B_UnoDeeOr7_0),.clk(gclk));
	jdff dff_B_tCwpCsJa9_0(.din(w_dff_B_UnoDeeOr7_0),.dout(w_dff_B_tCwpCsJa9_0),.clk(gclk));
	jdff dff_B_pCwSTHxS9_0(.din(w_dff_B_tCwpCsJa9_0),.dout(w_dff_B_pCwSTHxS9_0),.clk(gclk));
	jdff dff_B_Tfa6iLBB6_0(.din(w_dff_B_pCwSTHxS9_0),.dout(w_dff_B_Tfa6iLBB6_0),.clk(gclk));
	jdff dff_B_JCmdtD7q6_0(.din(w_dff_B_Tfa6iLBB6_0),.dout(w_dff_B_JCmdtD7q6_0),.clk(gclk));
	jdff dff_B_FIzmcAae6_0(.din(w_dff_B_JCmdtD7q6_0),.dout(w_dff_B_FIzmcAae6_0),.clk(gclk));
	jdff dff_B_WYMQiob36_0(.din(w_dff_B_FIzmcAae6_0),.dout(w_dff_B_WYMQiob36_0),.clk(gclk));
	jdff dff_B_anDCubS42_0(.din(w_dff_B_WYMQiob36_0),.dout(w_dff_B_anDCubS42_0),.clk(gclk));
	jdff dff_B_PygIc9OI4_0(.din(w_dff_B_anDCubS42_0),.dout(w_dff_B_PygIc9OI4_0),.clk(gclk));
	jdff dff_B_nSy1uQnu2_0(.din(w_dff_B_PygIc9OI4_0),.dout(w_dff_B_nSy1uQnu2_0),.clk(gclk));
	jdff dff_B_JvDs4JAs1_0(.din(w_dff_B_nSy1uQnu2_0),.dout(w_dff_B_JvDs4JAs1_0),.clk(gclk));
	jdff dff_B_1fNWwNfy0_1(.din(n864),.dout(w_dff_B_1fNWwNfy0_1),.clk(gclk));
	jdff dff_B_0hMFpWJF4_1(.din(w_dff_B_1fNWwNfy0_1),.dout(w_dff_B_0hMFpWJF4_1),.clk(gclk));
	jdff dff_B_ohVW7VIx3_1(.din(w_dff_B_0hMFpWJF4_1),.dout(w_dff_B_ohVW7VIx3_1),.clk(gclk));
	jdff dff_B_bojFVHxi6_1(.din(w_dff_B_ohVW7VIx3_1),.dout(w_dff_B_bojFVHxi6_1),.clk(gclk));
	jdff dff_B_U1RRFvWX4_1(.din(w_dff_B_bojFVHxi6_1),.dout(w_dff_B_U1RRFvWX4_1),.clk(gclk));
	jdff dff_B_k6RWaLjO8_1(.din(w_dff_B_U1RRFvWX4_1),.dout(w_dff_B_k6RWaLjO8_1),.clk(gclk));
	jdff dff_B_kwOVKXfA7_1(.din(w_dff_B_k6RWaLjO8_1),.dout(w_dff_B_kwOVKXfA7_1),.clk(gclk));
	jdff dff_B_5UzRbjzr2_1(.din(w_dff_B_kwOVKXfA7_1),.dout(w_dff_B_5UzRbjzr2_1),.clk(gclk));
	jdff dff_B_FODG8SnM9_1(.din(w_dff_B_5UzRbjzr2_1),.dout(w_dff_B_FODG8SnM9_1),.clk(gclk));
	jdff dff_B_e6TUD5kF7_1(.din(w_dff_B_FODG8SnM9_1),.dout(w_dff_B_e6TUD5kF7_1),.clk(gclk));
	jdff dff_B_3ahSLU0f5_1(.din(w_dff_B_e6TUD5kF7_1),.dout(w_dff_B_3ahSLU0f5_1),.clk(gclk));
	jdff dff_B_GIKKA03y8_1(.din(w_dff_B_3ahSLU0f5_1),.dout(w_dff_B_GIKKA03y8_1),.clk(gclk));
	jdff dff_B_SS6WDjzM5_1(.din(w_dff_B_GIKKA03y8_1),.dout(w_dff_B_SS6WDjzM5_1),.clk(gclk));
	jdff dff_B_cWw19qAf3_1(.din(w_dff_B_SS6WDjzM5_1),.dout(w_dff_B_cWw19qAf3_1),.clk(gclk));
	jdff dff_B_BFNjEJig8_1(.din(w_dff_B_cWw19qAf3_1),.dout(w_dff_B_BFNjEJig8_1),.clk(gclk));
	jdff dff_B_Kjp1X3wj4_1(.din(w_dff_B_BFNjEJig8_1),.dout(w_dff_B_Kjp1X3wj4_1),.clk(gclk));
	jdff dff_B_yxCjC1Eo5_1(.din(w_dff_B_Kjp1X3wj4_1),.dout(w_dff_B_yxCjC1Eo5_1),.clk(gclk));
	jdff dff_B_SeajZeG01_1(.din(w_dff_B_yxCjC1Eo5_1),.dout(w_dff_B_SeajZeG01_1),.clk(gclk));
	jdff dff_B_1brRFTAQ7_1(.din(w_dff_B_SeajZeG01_1),.dout(w_dff_B_1brRFTAQ7_1),.clk(gclk));
	jdff dff_B_jVBvabbt5_1(.din(w_dff_B_1brRFTAQ7_1),.dout(w_dff_B_jVBvabbt5_1),.clk(gclk));
	jdff dff_B_1ZYustJz1_1(.din(w_dff_B_jVBvabbt5_1),.dout(w_dff_B_1ZYustJz1_1),.clk(gclk));
	jdff dff_B_YVdG32KG6_1(.din(w_dff_B_1ZYustJz1_1),.dout(w_dff_B_YVdG32KG6_1),.clk(gclk));
	jdff dff_B_P6WDcFKN9_1(.din(w_dff_B_YVdG32KG6_1),.dout(w_dff_B_P6WDcFKN9_1),.clk(gclk));
	jdff dff_B_IGqHtOAZ5_1(.din(w_dff_B_P6WDcFKN9_1),.dout(w_dff_B_IGqHtOAZ5_1),.clk(gclk));
	jdff dff_B_oCAn17SR0_1(.din(w_dff_B_IGqHtOAZ5_1),.dout(w_dff_B_oCAn17SR0_1),.clk(gclk));
	jdff dff_B_KXbAAbK76_1(.din(w_dff_B_oCAn17SR0_1),.dout(w_dff_B_KXbAAbK76_1),.clk(gclk));
	jdff dff_B_pwEezPyR0_1(.din(w_dff_B_KXbAAbK76_1),.dout(w_dff_B_pwEezPyR0_1),.clk(gclk));
	jdff dff_B_A5znvr275_1(.din(w_dff_B_pwEezPyR0_1),.dout(w_dff_B_A5znvr275_1),.clk(gclk));
	jdff dff_B_VXehlGKy3_1(.din(w_dff_B_A5znvr275_1),.dout(w_dff_B_VXehlGKy3_1),.clk(gclk));
	jdff dff_B_EdIecont7_1(.din(w_dff_B_VXehlGKy3_1),.dout(w_dff_B_EdIecont7_1),.clk(gclk));
	jdff dff_B_tx1DN6rz5_1(.din(w_dff_B_EdIecont7_1),.dout(w_dff_B_tx1DN6rz5_1),.clk(gclk));
	jdff dff_B_fnIfyBF51_1(.din(w_dff_B_tx1DN6rz5_1),.dout(w_dff_B_fnIfyBF51_1),.clk(gclk));
	jdff dff_B_bAT882n93_1(.din(w_dff_B_fnIfyBF51_1),.dout(w_dff_B_bAT882n93_1),.clk(gclk));
	jdff dff_B_OhRJB9ro3_1(.din(w_dff_B_bAT882n93_1),.dout(w_dff_B_OhRJB9ro3_1),.clk(gclk));
	jdff dff_B_cZfPFW8I5_1(.din(w_dff_B_OhRJB9ro3_1),.dout(w_dff_B_cZfPFW8I5_1),.clk(gclk));
	jdff dff_B_DQG9O0KZ1_1(.din(w_dff_B_cZfPFW8I5_1),.dout(w_dff_B_DQG9O0KZ1_1),.clk(gclk));
	jdff dff_B_pRpKWNyO9_1(.din(w_dff_B_DQG9O0KZ1_1),.dout(w_dff_B_pRpKWNyO9_1),.clk(gclk));
	jdff dff_B_aWFkOS0o6_1(.din(w_dff_B_pRpKWNyO9_1),.dout(w_dff_B_aWFkOS0o6_1),.clk(gclk));
	jdff dff_B_dRiK9Ukz0_1(.din(w_dff_B_aWFkOS0o6_1),.dout(w_dff_B_dRiK9Ukz0_1),.clk(gclk));
	jdff dff_B_cduITGCM4_1(.din(w_dff_B_dRiK9Ukz0_1),.dout(w_dff_B_cduITGCM4_1),.clk(gclk));
	jdff dff_B_gqbX7jdF0_1(.din(w_dff_B_cduITGCM4_1),.dout(w_dff_B_gqbX7jdF0_1),.clk(gclk));
	jdff dff_B_hFQT1YAU5_1(.din(w_dff_B_gqbX7jdF0_1),.dout(w_dff_B_hFQT1YAU5_1),.clk(gclk));
	jdff dff_B_hkJ3ShXI0_1(.din(w_dff_B_hFQT1YAU5_1),.dout(w_dff_B_hkJ3ShXI0_1),.clk(gclk));
	jdff dff_B_5vb6oOpc8_1(.din(w_dff_B_hkJ3ShXI0_1),.dout(w_dff_B_5vb6oOpc8_1),.clk(gclk));
	jdff dff_B_nZg0GdcQ2_1(.din(w_dff_B_5vb6oOpc8_1),.dout(w_dff_B_nZg0GdcQ2_1),.clk(gclk));
	jdff dff_B_EFlFV7KA5_1(.din(w_dff_B_nZg0GdcQ2_1),.dout(w_dff_B_EFlFV7KA5_1),.clk(gclk));
	jdff dff_B_FSmo0P7R4_1(.din(w_dff_B_EFlFV7KA5_1),.dout(w_dff_B_FSmo0P7R4_1),.clk(gclk));
	jdff dff_B_3J7wgZMo8_1(.din(w_dff_B_FSmo0P7R4_1),.dout(w_dff_B_3J7wgZMo8_1),.clk(gclk));
	jdff dff_B_sYvKG95B8_1(.din(w_dff_B_3J7wgZMo8_1),.dout(w_dff_B_sYvKG95B8_1),.clk(gclk));
	jdff dff_B_YJaQeKRC6_1(.din(w_dff_B_sYvKG95B8_1),.dout(w_dff_B_YJaQeKRC6_1),.clk(gclk));
	jdff dff_B_ZxSgdjvF3_1(.din(w_dff_B_YJaQeKRC6_1),.dout(w_dff_B_ZxSgdjvF3_1),.clk(gclk));
	jdff dff_B_eLDVdvK05_1(.din(w_dff_B_ZxSgdjvF3_1),.dout(w_dff_B_eLDVdvK05_1),.clk(gclk));
	jdff dff_B_leSJa8mv3_1(.din(w_dff_B_eLDVdvK05_1),.dout(w_dff_B_leSJa8mv3_1),.clk(gclk));
	jdff dff_B_emB1c9tb6_1(.din(w_dff_B_leSJa8mv3_1),.dout(w_dff_B_emB1c9tb6_1),.clk(gclk));
	jdff dff_B_ovrDLKBA1_1(.din(w_dff_B_emB1c9tb6_1),.dout(w_dff_B_ovrDLKBA1_1),.clk(gclk));
	jdff dff_B_CSf3cnQF3_1(.din(w_dff_B_ovrDLKBA1_1),.dout(w_dff_B_CSf3cnQF3_1),.clk(gclk));
	jdff dff_B_qWbXoKNO7_1(.din(w_dff_B_CSf3cnQF3_1),.dout(w_dff_B_qWbXoKNO7_1),.clk(gclk));
	jdff dff_B_ODxQMLDb6_1(.din(w_dff_B_qWbXoKNO7_1),.dout(w_dff_B_ODxQMLDb6_1),.clk(gclk));
	jdff dff_B_ZwTNwGA55_1(.din(w_dff_B_ODxQMLDb6_1),.dout(w_dff_B_ZwTNwGA55_1),.clk(gclk));
	jdff dff_B_R3xUGviu9_1(.din(w_dff_B_ZwTNwGA55_1),.dout(w_dff_B_R3xUGviu9_1),.clk(gclk));
	jdff dff_B_EN1NQcku8_1(.din(w_dff_B_R3xUGviu9_1),.dout(w_dff_B_EN1NQcku8_1),.clk(gclk));
	jdff dff_B_1LGb7X9i6_1(.din(w_dff_B_EN1NQcku8_1),.dout(w_dff_B_1LGb7X9i6_1),.clk(gclk));
	jdff dff_B_y4Vxv6FO7_1(.din(w_dff_B_1LGb7X9i6_1),.dout(w_dff_B_y4Vxv6FO7_1),.clk(gclk));
	jdff dff_B_csX0uRYy5_1(.din(w_dff_B_y4Vxv6FO7_1),.dout(w_dff_B_csX0uRYy5_1),.clk(gclk));
	jdff dff_B_mFe7Unt29_1(.din(w_dff_B_csX0uRYy5_1),.dout(w_dff_B_mFe7Unt29_1),.clk(gclk));
	jdff dff_B_WAZikE3v7_1(.din(w_dff_B_mFe7Unt29_1),.dout(w_dff_B_WAZikE3v7_1),.clk(gclk));
	jdff dff_B_8tIQy2SM3_1(.din(w_dff_B_WAZikE3v7_1),.dout(w_dff_B_8tIQy2SM3_1),.clk(gclk));
	jdff dff_B_1S442Ar52_1(.din(w_dff_B_8tIQy2SM3_1),.dout(w_dff_B_1S442Ar52_1),.clk(gclk));
	jdff dff_B_aj23fqra7_1(.din(w_dff_B_1S442Ar52_1),.dout(w_dff_B_aj23fqra7_1),.clk(gclk));
	jdff dff_B_8SQNheKS0_1(.din(w_dff_B_aj23fqra7_1),.dout(w_dff_B_8SQNheKS0_1),.clk(gclk));
	jdff dff_B_nviS5O506_1(.din(w_dff_B_8SQNheKS0_1),.dout(w_dff_B_nviS5O506_1),.clk(gclk));
	jdff dff_B_eIl5V82O6_1(.din(w_dff_B_nviS5O506_1),.dout(w_dff_B_eIl5V82O6_1),.clk(gclk));
	jdff dff_B_3pOx5mzZ5_1(.din(w_dff_B_eIl5V82O6_1),.dout(w_dff_B_3pOx5mzZ5_1),.clk(gclk));
	jdff dff_B_w3vnM6zc0_1(.din(w_dff_B_3pOx5mzZ5_1),.dout(w_dff_B_w3vnM6zc0_1),.clk(gclk));
	jdff dff_B_5SuKWVLd3_1(.din(w_dff_B_w3vnM6zc0_1),.dout(w_dff_B_5SuKWVLd3_1),.clk(gclk));
	jdff dff_B_PDF1HE6X2_1(.din(w_dff_B_5SuKWVLd3_1),.dout(w_dff_B_PDF1HE6X2_1),.clk(gclk));
	jdff dff_B_xD6nLRAA9_1(.din(w_dff_B_PDF1HE6X2_1),.dout(w_dff_B_xD6nLRAA9_1),.clk(gclk));
	jdff dff_B_5Zwwjfqu1_1(.din(w_dff_B_xD6nLRAA9_1),.dout(w_dff_B_5Zwwjfqu1_1),.clk(gclk));
	jdff dff_B_nRpberWk8_1(.din(w_dff_B_5Zwwjfqu1_1),.dout(w_dff_B_nRpberWk8_1),.clk(gclk));
	jdff dff_B_e84DdMJl5_1(.din(w_dff_B_nRpberWk8_1),.dout(w_dff_B_e84DdMJl5_1),.clk(gclk));
	jdff dff_B_LA8nUIhW1_0(.din(n865),.dout(w_dff_B_LA8nUIhW1_0),.clk(gclk));
	jdff dff_B_UlwaVDyo4_0(.din(w_dff_B_LA8nUIhW1_0),.dout(w_dff_B_UlwaVDyo4_0),.clk(gclk));
	jdff dff_B_WsGbYJHm5_0(.din(w_dff_B_UlwaVDyo4_0),.dout(w_dff_B_WsGbYJHm5_0),.clk(gclk));
	jdff dff_B_joZJAjTz7_0(.din(w_dff_B_WsGbYJHm5_0),.dout(w_dff_B_joZJAjTz7_0),.clk(gclk));
	jdff dff_B_bGHwirTb0_0(.din(w_dff_B_joZJAjTz7_0),.dout(w_dff_B_bGHwirTb0_0),.clk(gclk));
	jdff dff_B_sjPjaM7I3_0(.din(w_dff_B_bGHwirTb0_0),.dout(w_dff_B_sjPjaM7I3_0),.clk(gclk));
	jdff dff_B_uA4c2xIE5_0(.din(w_dff_B_sjPjaM7I3_0),.dout(w_dff_B_uA4c2xIE5_0),.clk(gclk));
	jdff dff_B_5EoqFvgV4_0(.din(w_dff_B_uA4c2xIE5_0),.dout(w_dff_B_5EoqFvgV4_0),.clk(gclk));
	jdff dff_B_ohalHl3I7_0(.din(w_dff_B_5EoqFvgV4_0),.dout(w_dff_B_ohalHl3I7_0),.clk(gclk));
	jdff dff_B_VuRCtj7r9_0(.din(w_dff_B_ohalHl3I7_0),.dout(w_dff_B_VuRCtj7r9_0),.clk(gclk));
	jdff dff_B_93txWX9V4_0(.din(w_dff_B_VuRCtj7r9_0),.dout(w_dff_B_93txWX9V4_0),.clk(gclk));
	jdff dff_B_fjicCr5Z6_0(.din(w_dff_B_93txWX9V4_0),.dout(w_dff_B_fjicCr5Z6_0),.clk(gclk));
	jdff dff_B_mGafTpnt9_0(.din(w_dff_B_fjicCr5Z6_0),.dout(w_dff_B_mGafTpnt9_0),.clk(gclk));
	jdff dff_B_hOdSlX2K2_0(.din(w_dff_B_mGafTpnt9_0),.dout(w_dff_B_hOdSlX2K2_0),.clk(gclk));
	jdff dff_B_BusYKFN71_0(.din(w_dff_B_hOdSlX2K2_0),.dout(w_dff_B_BusYKFN71_0),.clk(gclk));
	jdff dff_B_yJ07B1S13_0(.din(w_dff_B_BusYKFN71_0),.dout(w_dff_B_yJ07B1S13_0),.clk(gclk));
	jdff dff_B_07V96llp4_0(.din(w_dff_B_yJ07B1S13_0),.dout(w_dff_B_07V96llp4_0),.clk(gclk));
	jdff dff_B_hjFWNCWA7_0(.din(w_dff_B_07V96llp4_0),.dout(w_dff_B_hjFWNCWA7_0),.clk(gclk));
	jdff dff_B_SOpCPN7r2_0(.din(w_dff_B_hjFWNCWA7_0),.dout(w_dff_B_SOpCPN7r2_0),.clk(gclk));
	jdff dff_B_FTtsVcvj6_0(.din(w_dff_B_SOpCPN7r2_0),.dout(w_dff_B_FTtsVcvj6_0),.clk(gclk));
	jdff dff_B_EtWZMNfG2_0(.din(w_dff_B_FTtsVcvj6_0),.dout(w_dff_B_EtWZMNfG2_0),.clk(gclk));
	jdff dff_B_L677Jlfv4_0(.din(w_dff_B_EtWZMNfG2_0),.dout(w_dff_B_L677Jlfv4_0),.clk(gclk));
	jdff dff_B_sZfXbixm5_0(.din(w_dff_B_L677Jlfv4_0),.dout(w_dff_B_sZfXbixm5_0),.clk(gclk));
	jdff dff_B_IPzOYziY9_0(.din(w_dff_B_sZfXbixm5_0),.dout(w_dff_B_IPzOYziY9_0),.clk(gclk));
	jdff dff_B_1XvA1Jmo0_0(.din(w_dff_B_IPzOYziY9_0),.dout(w_dff_B_1XvA1Jmo0_0),.clk(gclk));
	jdff dff_B_9gBZcg8H3_0(.din(w_dff_B_1XvA1Jmo0_0),.dout(w_dff_B_9gBZcg8H3_0),.clk(gclk));
	jdff dff_B_12hH4dGZ5_0(.din(w_dff_B_9gBZcg8H3_0),.dout(w_dff_B_12hH4dGZ5_0),.clk(gclk));
	jdff dff_B_7LbisSyT2_0(.din(w_dff_B_12hH4dGZ5_0),.dout(w_dff_B_7LbisSyT2_0),.clk(gclk));
	jdff dff_B_mtPh5xJ10_0(.din(w_dff_B_7LbisSyT2_0),.dout(w_dff_B_mtPh5xJ10_0),.clk(gclk));
	jdff dff_B_FPDXdtsm1_0(.din(w_dff_B_mtPh5xJ10_0),.dout(w_dff_B_FPDXdtsm1_0),.clk(gclk));
	jdff dff_B_07N54mPD2_0(.din(w_dff_B_FPDXdtsm1_0),.dout(w_dff_B_07N54mPD2_0),.clk(gclk));
	jdff dff_B_gJ0yOhSL0_0(.din(w_dff_B_07N54mPD2_0),.dout(w_dff_B_gJ0yOhSL0_0),.clk(gclk));
	jdff dff_B_R6xK6GA07_0(.din(w_dff_B_gJ0yOhSL0_0),.dout(w_dff_B_R6xK6GA07_0),.clk(gclk));
	jdff dff_B_Nz9McD6Q8_0(.din(w_dff_B_R6xK6GA07_0),.dout(w_dff_B_Nz9McD6Q8_0),.clk(gclk));
	jdff dff_B_tsPwY25c3_0(.din(w_dff_B_Nz9McD6Q8_0),.dout(w_dff_B_tsPwY25c3_0),.clk(gclk));
	jdff dff_B_Sa3VBwqB5_0(.din(w_dff_B_tsPwY25c3_0),.dout(w_dff_B_Sa3VBwqB5_0),.clk(gclk));
	jdff dff_B_QPv0mvlg0_0(.din(w_dff_B_Sa3VBwqB5_0),.dout(w_dff_B_QPv0mvlg0_0),.clk(gclk));
	jdff dff_B_eO1IIRFA4_0(.din(w_dff_B_QPv0mvlg0_0),.dout(w_dff_B_eO1IIRFA4_0),.clk(gclk));
	jdff dff_B_S1UjzQh42_0(.din(w_dff_B_eO1IIRFA4_0),.dout(w_dff_B_S1UjzQh42_0),.clk(gclk));
	jdff dff_B_N5ROz9rz6_0(.din(w_dff_B_S1UjzQh42_0),.dout(w_dff_B_N5ROz9rz6_0),.clk(gclk));
	jdff dff_B_eFnN80HK4_0(.din(w_dff_B_N5ROz9rz6_0),.dout(w_dff_B_eFnN80HK4_0),.clk(gclk));
	jdff dff_B_O5e8Amcy6_0(.din(w_dff_B_eFnN80HK4_0),.dout(w_dff_B_O5e8Amcy6_0),.clk(gclk));
	jdff dff_B_VD38JG0M7_0(.din(w_dff_B_O5e8Amcy6_0),.dout(w_dff_B_VD38JG0M7_0),.clk(gclk));
	jdff dff_B_mEcvTa2v6_0(.din(w_dff_B_VD38JG0M7_0),.dout(w_dff_B_mEcvTa2v6_0),.clk(gclk));
	jdff dff_B_MvVy2GtC7_0(.din(w_dff_B_mEcvTa2v6_0),.dout(w_dff_B_MvVy2GtC7_0),.clk(gclk));
	jdff dff_B_BMZ9kfZd3_0(.din(w_dff_B_MvVy2GtC7_0),.dout(w_dff_B_BMZ9kfZd3_0),.clk(gclk));
	jdff dff_B_EISWj2oM1_0(.din(w_dff_B_BMZ9kfZd3_0),.dout(w_dff_B_EISWj2oM1_0),.clk(gclk));
	jdff dff_B_BzdIBGA48_0(.din(w_dff_B_EISWj2oM1_0),.dout(w_dff_B_BzdIBGA48_0),.clk(gclk));
	jdff dff_B_iSM6W20w8_0(.din(w_dff_B_BzdIBGA48_0),.dout(w_dff_B_iSM6W20w8_0),.clk(gclk));
	jdff dff_B_sogyuxOg0_0(.din(w_dff_B_iSM6W20w8_0),.dout(w_dff_B_sogyuxOg0_0),.clk(gclk));
	jdff dff_B_VE8BkZXE0_0(.din(w_dff_B_sogyuxOg0_0),.dout(w_dff_B_VE8BkZXE0_0),.clk(gclk));
	jdff dff_B_cpt6ZdiB9_0(.din(w_dff_B_VE8BkZXE0_0),.dout(w_dff_B_cpt6ZdiB9_0),.clk(gclk));
	jdff dff_B_8Ywpla247_0(.din(w_dff_B_cpt6ZdiB9_0),.dout(w_dff_B_8Ywpla247_0),.clk(gclk));
	jdff dff_B_CHNqhXo22_0(.din(w_dff_B_8Ywpla247_0),.dout(w_dff_B_CHNqhXo22_0),.clk(gclk));
	jdff dff_B_DsBOklLR6_0(.din(w_dff_B_CHNqhXo22_0),.dout(w_dff_B_DsBOklLR6_0),.clk(gclk));
	jdff dff_B_fVhNd03m0_0(.din(w_dff_B_DsBOklLR6_0),.dout(w_dff_B_fVhNd03m0_0),.clk(gclk));
	jdff dff_B_inBtQ2Fh1_0(.din(w_dff_B_fVhNd03m0_0),.dout(w_dff_B_inBtQ2Fh1_0),.clk(gclk));
	jdff dff_B_LvRMYlsV7_0(.din(w_dff_B_inBtQ2Fh1_0),.dout(w_dff_B_LvRMYlsV7_0),.clk(gclk));
	jdff dff_B_mWZPlMUn1_0(.din(w_dff_B_LvRMYlsV7_0),.dout(w_dff_B_mWZPlMUn1_0),.clk(gclk));
	jdff dff_B_FG0yEm768_0(.din(w_dff_B_mWZPlMUn1_0),.dout(w_dff_B_FG0yEm768_0),.clk(gclk));
	jdff dff_B_Wgklik3i7_0(.din(w_dff_B_FG0yEm768_0),.dout(w_dff_B_Wgklik3i7_0),.clk(gclk));
	jdff dff_B_e4ZRLmT65_0(.din(w_dff_B_Wgklik3i7_0),.dout(w_dff_B_e4ZRLmT65_0),.clk(gclk));
	jdff dff_B_uc4EemAt8_0(.din(w_dff_B_e4ZRLmT65_0),.dout(w_dff_B_uc4EemAt8_0),.clk(gclk));
	jdff dff_B_v62cHd8i6_0(.din(w_dff_B_uc4EemAt8_0),.dout(w_dff_B_v62cHd8i6_0),.clk(gclk));
	jdff dff_B_8bZh3vep5_0(.din(w_dff_B_v62cHd8i6_0),.dout(w_dff_B_8bZh3vep5_0),.clk(gclk));
	jdff dff_B_IN6Z1lU39_0(.din(w_dff_B_8bZh3vep5_0),.dout(w_dff_B_IN6Z1lU39_0),.clk(gclk));
	jdff dff_B_xO2ENmm82_0(.din(w_dff_B_IN6Z1lU39_0),.dout(w_dff_B_xO2ENmm82_0),.clk(gclk));
	jdff dff_B_bc4YtK6Z7_0(.din(w_dff_B_xO2ENmm82_0),.dout(w_dff_B_bc4YtK6Z7_0),.clk(gclk));
	jdff dff_B_YhHx2WQc0_0(.din(w_dff_B_bc4YtK6Z7_0),.dout(w_dff_B_YhHx2WQc0_0),.clk(gclk));
	jdff dff_B_JSwaYugR5_0(.din(w_dff_B_YhHx2WQc0_0),.dout(w_dff_B_JSwaYugR5_0),.clk(gclk));
	jdff dff_B_XRyY7pT98_0(.din(w_dff_B_JSwaYugR5_0),.dout(w_dff_B_XRyY7pT98_0),.clk(gclk));
	jdff dff_B_sKB8gmvT8_0(.din(w_dff_B_XRyY7pT98_0),.dout(w_dff_B_sKB8gmvT8_0),.clk(gclk));
	jdff dff_B_VaegOeAt7_0(.din(w_dff_B_sKB8gmvT8_0),.dout(w_dff_B_VaegOeAt7_0),.clk(gclk));
	jdff dff_B_gXkYNe7n9_0(.din(w_dff_B_VaegOeAt7_0),.dout(w_dff_B_gXkYNe7n9_0),.clk(gclk));
	jdff dff_B_pW8kc4Be2_0(.din(w_dff_B_gXkYNe7n9_0),.dout(w_dff_B_pW8kc4Be2_0),.clk(gclk));
	jdff dff_B_tnRPek717_0(.din(w_dff_B_pW8kc4Be2_0),.dout(w_dff_B_tnRPek717_0),.clk(gclk));
	jdff dff_B_ysmONgPT3_0(.din(w_dff_B_tnRPek717_0),.dout(w_dff_B_ysmONgPT3_0),.clk(gclk));
	jdff dff_B_o5w7wT8k3_0(.din(w_dff_B_ysmONgPT3_0),.dout(w_dff_B_o5w7wT8k3_0),.clk(gclk));
	jdff dff_B_HgzYxPhY9_0(.din(w_dff_B_o5w7wT8k3_0),.dout(w_dff_B_HgzYxPhY9_0),.clk(gclk));
	jdff dff_B_MhnprG8l9_0(.din(w_dff_B_HgzYxPhY9_0),.dout(w_dff_B_MhnprG8l9_0),.clk(gclk));
	jdff dff_B_qceRoBmQ1_1(.din(n858),.dout(w_dff_B_qceRoBmQ1_1),.clk(gclk));
	jdff dff_B_nuicdX2j0_1(.din(w_dff_B_qceRoBmQ1_1),.dout(w_dff_B_nuicdX2j0_1),.clk(gclk));
	jdff dff_B_KhD2OBuk3_1(.din(w_dff_B_nuicdX2j0_1),.dout(w_dff_B_KhD2OBuk3_1),.clk(gclk));
	jdff dff_B_4JJj7Ghw4_1(.din(w_dff_B_KhD2OBuk3_1),.dout(w_dff_B_4JJj7Ghw4_1),.clk(gclk));
	jdff dff_B_QHMVQmaQ1_1(.din(w_dff_B_4JJj7Ghw4_1),.dout(w_dff_B_QHMVQmaQ1_1),.clk(gclk));
	jdff dff_B_706k3QG64_1(.din(w_dff_B_QHMVQmaQ1_1),.dout(w_dff_B_706k3QG64_1),.clk(gclk));
	jdff dff_B_i0ZmiZkZ5_1(.din(w_dff_B_706k3QG64_1),.dout(w_dff_B_i0ZmiZkZ5_1),.clk(gclk));
	jdff dff_B_RWCUxv5t6_1(.din(w_dff_B_i0ZmiZkZ5_1),.dout(w_dff_B_RWCUxv5t6_1),.clk(gclk));
	jdff dff_B_7B9YVItL2_1(.din(w_dff_B_RWCUxv5t6_1),.dout(w_dff_B_7B9YVItL2_1),.clk(gclk));
	jdff dff_B_oO4vhS9F3_1(.din(w_dff_B_7B9YVItL2_1),.dout(w_dff_B_oO4vhS9F3_1),.clk(gclk));
	jdff dff_B_uEi0WiuB0_1(.din(w_dff_B_oO4vhS9F3_1),.dout(w_dff_B_uEi0WiuB0_1),.clk(gclk));
	jdff dff_B_abEnW9Zc4_1(.din(w_dff_B_uEi0WiuB0_1),.dout(w_dff_B_abEnW9Zc4_1),.clk(gclk));
	jdff dff_B_UzQodXDE8_1(.din(w_dff_B_abEnW9Zc4_1),.dout(w_dff_B_UzQodXDE8_1),.clk(gclk));
	jdff dff_B_zPdKUbsG2_1(.din(w_dff_B_UzQodXDE8_1),.dout(w_dff_B_zPdKUbsG2_1),.clk(gclk));
	jdff dff_B_CYJARK1g6_1(.din(w_dff_B_zPdKUbsG2_1),.dout(w_dff_B_CYJARK1g6_1),.clk(gclk));
	jdff dff_B_Oii4CUX08_1(.din(w_dff_B_CYJARK1g6_1),.dout(w_dff_B_Oii4CUX08_1),.clk(gclk));
	jdff dff_B_hF4uKHVr3_1(.din(w_dff_B_Oii4CUX08_1),.dout(w_dff_B_hF4uKHVr3_1),.clk(gclk));
	jdff dff_B_lOMYp8Kt3_1(.din(w_dff_B_hF4uKHVr3_1),.dout(w_dff_B_lOMYp8Kt3_1),.clk(gclk));
	jdff dff_B_2ahuWX887_1(.din(w_dff_B_lOMYp8Kt3_1),.dout(w_dff_B_2ahuWX887_1),.clk(gclk));
	jdff dff_B_JMGiE6G57_1(.din(w_dff_B_2ahuWX887_1),.dout(w_dff_B_JMGiE6G57_1),.clk(gclk));
	jdff dff_B_TDtMm0XF1_1(.din(w_dff_B_JMGiE6G57_1),.dout(w_dff_B_TDtMm0XF1_1),.clk(gclk));
	jdff dff_B_UWnr3xXR6_1(.din(w_dff_B_TDtMm0XF1_1),.dout(w_dff_B_UWnr3xXR6_1),.clk(gclk));
	jdff dff_B_lFTYaQDp8_1(.din(w_dff_B_UWnr3xXR6_1),.dout(w_dff_B_lFTYaQDp8_1),.clk(gclk));
	jdff dff_B_L7kOx4Gv5_1(.din(w_dff_B_lFTYaQDp8_1),.dout(w_dff_B_L7kOx4Gv5_1),.clk(gclk));
	jdff dff_B_sAWqPKB59_1(.din(w_dff_B_L7kOx4Gv5_1),.dout(w_dff_B_sAWqPKB59_1),.clk(gclk));
	jdff dff_B_VzLpQoOw6_1(.din(w_dff_B_sAWqPKB59_1),.dout(w_dff_B_VzLpQoOw6_1),.clk(gclk));
	jdff dff_B_rhEZciPG6_1(.din(w_dff_B_VzLpQoOw6_1),.dout(w_dff_B_rhEZciPG6_1),.clk(gclk));
	jdff dff_B_fVOMApE95_1(.din(w_dff_B_rhEZciPG6_1),.dout(w_dff_B_fVOMApE95_1),.clk(gclk));
	jdff dff_B_jgMf64ZO3_1(.din(w_dff_B_fVOMApE95_1),.dout(w_dff_B_jgMf64ZO3_1),.clk(gclk));
	jdff dff_B_FjREz1Ko1_1(.din(w_dff_B_jgMf64ZO3_1),.dout(w_dff_B_FjREz1Ko1_1),.clk(gclk));
	jdff dff_B_RWsC1hqg3_1(.din(w_dff_B_FjREz1Ko1_1),.dout(w_dff_B_RWsC1hqg3_1),.clk(gclk));
	jdff dff_B_YcC5qUWt7_1(.din(w_dff_B_RWsC1hqg3_1),.dout(w_dff_B_YcC5qUWt7_1),.clk(gclk));
	jdff dff_B_OjJcsPVX5_1(.din(w_dff_B_YcC5qUWt7_1),.dout(w_dff_B_OjJcsPVX5_1),.clk(gclk));
	jdff dff_B_rddN5v7d1_1(.din(w_dff_B_OjJcsPVX5_1),.dout(w_dff_B_rddN5v7d1_1),.clk(gclk));
	jdff dff_B_0VDSB8Kz6_1(.din(w_dff_B_rddN5v7d1_1),.dout(w_dff_B_0VDSB8Kz6_1),.clk(gclk));
	jdff dff_B_n7bb6j482_1(.din(w_dff_B_0VDSB8Kz6_1),.dout(w_dff_B_n7bb6j482_1),.clk(gclk));
	jdff dff_B_27vDazFn0_1(.din(w_dff_B_n7bb6j482_1),.dout(w_dff_B_27vDazFn0_1),.clk(gclk));
	jdff dff_B_cgp6ZmvE8_1(.din(w_dff_B_27vDazFn0_1),.dout(w_dff_B_cgp6ZmvE8_1),.clk(gclk));
	jdff dff_B_PcwTg4Nf8_1(.din(w_dff_B_cgp6ZmvE8_1),.dout(w_dff_B_PcwTg4Nf8_1),.clk(gclk));
	jdff dff_B_q5rNOSs75_1(.din(w_dff_B_PcwTg4Nf8_1),.dout(w_dff_B_q5rNOSs75_1),.clk(gclk));
	jdff dff_B_yFqsHu4m0_1(.din(w_dff_B_q5rNOSs75_1),.dout(w_dff_B_yFqsHu4m0_1),.clk(gclk));
	jdff dff_B_QYl9RcJo7_1(.din(w_dff_B_yFqsHu4m0_1),.dout(w_dff_B_QYl9RcJo7_1),.clk(gclk));
	jdff dff_B_zwRJYAip8_1(.din(w_dff_B_QYl9RcJo7_1),.dout(w_dff_B_zwRJYAip8_1),.clk(gclk));
	jdff dff_B_cB6U3jUe6_1(.din(w_dff_B_zwRJYAip8_1),.dout(w_dff_B_cB6U3jUe6_1),.clk(gclk));
	jdff dff_B_CWf4T7Q14_1(.din(w_dff_B_cB6U3jUe6_1),.dout(w_dff_B_CWf4T7Q14_1),.clk(gclk));
	jdff dff_B_YXNjCd5l2_1(.din(w_dff_B_CWf4T7Q14_1),.dout(w_dff_B_YXNjCd5l2_1),.clk(gclk));
	jdff dff_B_I7mOOrUk8_1(.din(w_dff_B_YXNjCd5l2_1),.dout(w_dff_B_I7mOOrUk8_1),.clk(gclk));
	jdff dff_B_xWYdAhSV0_1(.din(w_dff_B_I7mOOrUk8_1),.dout(w_dff_B_xWYdAhSV0_1),.clk(gclk));
	jdff dff_B_LWVgbbQf8_1(.din(w_dff_B_xWYdAhSV0_1),.dout(w_dff_B_LWVgbbQf8_1),.clk(gclk));
	jdff dff_B_ro2YST8v1_1(.din(w_dff_B_LWVgbbQf8_1),.dout(w_dff_B_ro2YST8v1_1),.clk(gclk));
	jdff dff_B_LYP36CjP9_1(.din(w_dff_B_ro2YST8v1_1),.dout(w_dff_B_LYP36CjP9_1),.clk(gclk));
	jdff dff_B_FWGwVdIL3_1(.din(w_dff_B_LYP36CjP9_1),.dout(w_dff_B_FWGwVdIL3_1),.clk(gclk));
	jdff dff_B_SZmvxS565_1(.din(w_dff_B_FWGwVdIL3_1),.dout(w_dff_B_SZmvxS565_1),.clk(gclk));
	jdff dff_B_osRZc0eC4_1(.din(w_dff_B_SZmvxS565_1),.dout(w_dff_B_osRZc0eC4_1),.clk(gclk));
	jdff dff_B_UIZFMvfW9_1(.din(w_dff_B_osRZc0eC4_1),.dout(w_dff_B_UIZFMvfW9_1),.clk(gclk));
	jdff dff_B_YcXqJC6S0_1(.din(w_dff_B_UIZFMvfW9_1),.dout(w_dff_B_YcXqJC6S0_1),.clk(gclk));
	jdff dff_B_w7HSpxz76_1(.din(w_dff_B_YcXqJC6S0_1),.dout(w_dff_B_w7HSpxz76_1),.clk(gclk));
	jdff dff_B_a33IaeeV4_1(.din(w_dff_B_w7HSpxz76_1),.dout(w_dff_B_a33IaeeV4_1),.clk(gclk));
	jdff dff_B_kVzCrytA1_1(.din(w_dff_B_a33IaeeV4_1),.dout(w_dff_B_kVzCrytA1_1),.clk(gclk));
	jdff dff_B_8PC2PrYQ7_1(.din(w_dff_B_kVzCrytA1_1),.dout(w_dff_B_8PC2PrYQ7_1),.clk(gclk));
	jdff dff_B_hA6Esfvs9_1(.din(w_dff_B_8PC2PrYQ7_1),.dout(w_dff_B_hA6Esfvs9_1),.clk(gclk));
	jdff dff_B_tUvVXCne1_1(.din(w_dff_B_hA6Esfvs9_1),.dout(w_dff_B_tUvVXCne1_1),.clk(gclk));
	jdff dff_B_n8NVf91s7_1(.din(w_dff_B_tUvVXCne1_1),.dout(w_dff_B_n8NVf91s7_1),.clk(gclk));
	jdff dff_B_7dc5sPpq5_1(.din(w_dff_B_n8NVf91s7_1),.dout(w_dff_B_7dc5sPpq5_1),.clk(gclk));
	jdff dff_B_ELIHhym96_1(.din(w_dff_B_7dc5sPpq5_1),.dout(w_dff_B_ELIHhym96_1),.clk(gclk));
	jdff dff_B_VFbNHcqM6_1(.din(w_dff_B_ELIHhym96_1),.dout(w_dff_B_VFbNHcqM6_1),.clk(gclk));
	jdff dff_B_xIwOwtEl0_1(.din(w_dff_B_VFbNHcqM6_1),.dout(w_dff_B_xIwOwtEl0_1),.clk(gclk));
	jdff dff_B_KFRsv0e36_1(.din(w_dff_B_xIwOwtEl0_1),.dout(w_dff_B_KFRsv0e36_1),.clk(gclk));
	jdff dff_B_WErrMpK48_1(.din(w_dff_B_KFRsv0e36_1),.dout(w_dff_B_WErrMpK48_1),.clk(gclk));
	jdff dff_B_IY6u5P0P2_1(.din(w_dff_B_WErrMpK48_1),.dout(w_dff_B_IY6u5P0P2_1),.clk(gclk));
	jdff dff_B_T8tVNFsk9_1(.din(w_dff_B_IY6u5P0P2_1),.dout(w_dff_B_T8tVNFsk9_1),.clk(gclk));
	jdff dff_B_HGObvQ0B4_1(.din(w_dff_B_T8tVNFsk9_1),.dout(w_dff_B_HGObvQ0B4_1),.clk(gclk));
	jdff dff_B_WmVuxury4_1(.din(w_dff_B_HGObvQ0B4_1),.dout(w_dff_B_WmVuxury4_1),.clk(gclk));
	jdff dff_B_rrrI6D1L4_1(.din(w_dff_B_WmVuxury4_1),.dout(w_dff_B_rrrI6D1L4_1),.clk(gclk));
	jdff dff_B_kWY03dVN0_1(.din(w_dff_B_rrrI6D1L4_1),.dout(w_dff_B_kWY03dVN0_1),.clk(gclk));
	jdff dff_B_qABRW3tr6_1(.din(w_dff_B_kWY03dVN0_1),.dout(w_dff_B_qABRW3tr6_1),.clk(gclk));
	jdff dff_B_RYu0Dyl48_1(.din(w_dff_B_qABRW3tr6_1),.dout(w_dff_B_RYu0Dyl48_1),.clk(gclk));
	jdff dff_B_HNvMBpKf9_1(.din(w_dff_B_RYu0Dyl48_1),.dout(w_dff_B_HNvMBpKf9_1),.clk(gclk));
	jdff dff_B_sIPXzDkp4_1(.din(w_dff_B_HNvMBpKf9_1),.dout(w_dff_B_sIPXzDkp4_1),.clk(gclk));
	jdff dff_B_C0HHHzh75_0(.din(n859),.dout(w_dff_B_C0HHHzh75_0),.clk(gclk));
	jdff dff_B_0unVWWyq5_0(.din(w_dff_B_C0HHHzh75_0),.dout(w_dff_B_0unVWWyq5_0),.clk(gclk));
	jdff dff_B_DYKWDjoX2_0(.din(w_dff_B_0unVWWyq5_0),.dout(w_dff_B_DYKWDjoX2_0),.clk(gclk));
	jdff dff_B_IYubbnKR7_0(.din(w_dff_B_DYKWDjoX2_0),.dout(w_dff_B_IYubbnKR7_0),.clk(gclk));
	jdff dff_B_QQk97jog6_0(.din(w_dff_B_IYubbnKR7_0),.dout(w_dff_B_QQk97jog6_0),.clk(gclk));
	jdff dff_B_01JquW444_0(.din(w_dff_B_QQk97jog6_0),.dout(w_dff_B_01JquW444_0),.clk(gclk));
	jdff dff_B_bJg4TdHi2_0(.din(w_dff_B_01JquW444_0),.dout(w_dff_B_bJg4TdHi2_0),.clk(gclk));
	jdff dff_B_qIRSSsbt1_0(.din(w_dff_B_bJg4TdHi2_0),.dout(w_dff_B_qIRSSsbt1_0),.clk(gclk));
	jdff dff_B_ahFmu9QF6_0(.din(w_dff_B_qIRSSsbt1_0),.dout(w_dff_B_ahFmu9QF6_0),.clk(gclk));
	jdff dff_B_ldvR4YwX7_0(.din(w_dff_B_ahFmu9QF6_0),.dout(w_dff_B_ldvR4YwX7_0),.clk(gclk));
	jdff dff_B_tn0WhfQ49_0(.din(w_dff_B_ldvR4YwX7_0),.dout(w_dff_B_tn0WhfQ49_0),.clk(gclk));
	jdff dff_B_aIbwPofl7_0(.din(w_dff_B_tn0WhfQ49_0),.dout(w_dff_B_aIbwPofl7_0),.clk(gclk));
	jdff dff_B_gDq3y9cm1_0(.din(w_dff_B_aIbwPofl7_0),.dout(w_dff_B_gDq3y9cm1_0),.clk(gclk));
	jdff dff_B_jh7p3t3W0_0(.din(w_dff_B_gDq3y9cm1_0),.dout(w_dff_B_jh7p3t3W0_0),.clk(gclk));
	jdff dff_B_Azk00dkJ0_0(.din(w_dff_B_jh7p3t3W0_0),.dout(w_dff_B_Azk00dkJ0_0),.clk(gclk));
	jdff dff_B_GkE1YKNl1_0(.din(w_dff_B_Azk00dkJ0_0),.dout(w_dff_B_GkE1YKNl1_0),.clk(gclk));
	jdff dff_B_DRBOY5cU8_0(.din(w_dff_B_GkE1YKNl1_0),.dout(w_dff_B_DRBOY5cU8_0),.clk(gclk));
	jdff dff_B_YyZ3OxUL0_0(.din(w_dff_B_DRBOY5cU8_0),.dout(w_dff_B_YyZ3OxUL0_0),.clk(gclk));
	jdff dff_B_qSezP5MA4_0(.din(w_dff_B_YyZ3OxUL0_0),.dout(w_dff_B_qSezP5MA4_0),.clk(gclk));
	jdff dff_B_EwXafume2_0(.din(w_dff_B_qSezP5MA4_0),.dout(w_dff_B_EwXafume2_0),.clk(gclk));
	jdff dff_B_SidiTEaW2_0(.din(w_dff_B_EwXafume2_0),.dout(w_dff_B_SidiTEaW2_0),.clk(gclk));
	jdff dff_B_WI4iuNYk9_0(.din(w_dff_B_SidiTEaW2_0),.dout(w_dff_B_WI4iuNYk9_0),.clk(gclk));
	jdff dff_B_gC1FqZfa3_0(.din(w_dff_B_WI4iuNYk9_0),.dout(w_dff_B_gC1FqZfa3_0),.clk(gclk));
	jdff dff_B_5dywQ92U5_0(.din(w_dff_B_gC1FqZfa3_0),.dout(w_dff_B_5dywQ92U5_0),.clk(gclk));
	jdff dff_B_Y9gyQyNF6_0(.din(w_dff_B_5dywQ92U5_0),.dout(w_dff_B_Y9gyQyNF6_0),.clk(gclk));
	jdff dff_B_RBi06g3M8_0(.din(w_dff_B_Y9gyQyNF6_0),.dout(w_dff_B_RBi06g3M8_0),.clk(gclk));
	jdff dff_B_xYbX8bbr1_0(.din(w_dff_B_RBi06g3M8_0),.dout(w_dff_B_xYbX8bbr1_0),.clk(gclk));
	jdff dff_B_WImmKUQa0_0(.din(w_dff_B_xYbX8bbr1_0),.dout(w_dff_B_WImmKUQa0_0),.clk(gclk));
	jdff dff_B_i13Vv1PM3_0(.din(w_dff_B_WImmKUQa0_0),.dout(w_dff_B_i13Vv1PM3_0),.clk(gclk));
	jdff dff_B_k4qQKCLj6_0(.din(w_dff_B_i13Vv1PM3_0),.dout(w_dff_B_k4qQKCLj6_0),.clk(gclk));
	jdff dff_B_Yd0LhWEN2_0(.din(w_dff_B_k4qQKCLj6_0),.dout(w_dff_B_Yd0LhWEN2_0),.clk(gclk));
	jdff dff_B_Eej5KYxV4_0(.din(w_dff_B_Yd0LhWEN2_0),.dout(w_dff_B_Eej5KYxV4_0),.clk(gclk));
	jdff dff_B_wgeHFxXT0_0(.din(w_dff_B_Eej5KYxV4_0),.dout(w_dff_B_wgeHFxXT0_0),.clk(gclk));
	jdff dff_B_LKW7eHky4_0(.din(w_dff_B_wgeHFxXT0_0),.dout(w_dff_B_LKW7eHky4_0),.clk(gclk));
	jdff dff_B_lLoufkls1_0(.din(w_dff_B_LKW7eHky4_0),.dout(w_dff_B_lLoufkls1_0),.clk(gclk));
	jdff dff_B_4rSgmUun2_0(.din(w_dff_B_lLoufkls1_0),.dout(w_dff_B_4rSgmUun2_0),.clk(gclk));
	jdff dff_B_cfoVcOpw7_0(.din(w_dff_B_4rSgmUun2_0),.dout(w_dff_B_cfoVcOpw7_0),.clk(gclk));
	jdff dff_B_2xrE3NSH1_0(.din(w_dff_B_cfoVcOpw7_0),.dout(w_dff_B_2xrE3NSH1_0),.clk(gclk));
	jdff dff_B_CcYX6sPK8_0(.din(w_dff_B_2xrE3NSH1_0),.dout(w_dff_B_CcYX6sPK8_0),.clk(gclk));
	jdff dff_B_Jwr9ud9u8_0(.din(w_dff_B_CcYX6sPK8_0),.dout(w_dff_B_Jwr9ud9u8_0),.clk(gclk));
	jdff dff_B_Y05VgRx63_0(.din(w_dff_B_Jwr9ud9u8_0),.dout(w_dff_B_Y05VgRx63_0),.clk(gclk));
	jdff dff_B_tv9e17wr1_0(.din(w_dff_B_Y05VgRx63_0),.dout(w_dff_B_tv9e17wr1_0),.clk(gclk));
	jdff dff_B_yjmp301p1_0(.din(w_dff_B_tv9e17wr1_0),.dout(w_dff_B_yjmp301p1_0),.clk(gclk));
	jdff dff_B_WFn3IAxy3_0(.din(w_dff_B_yjmp301p1_0),.dout(w_dff_B_WFn3IAxy3_0),.clk(gclk));
	jdff dff_B_fuOQSH5C1_0(.din(w_dff_B_WFn3IAxy3_0),.dout(w_dff_B_fuOQSH5C1_0),.clk(gclk));
	jdff dff_B_5ITfGVaQ2_0(.din(w_dff_B_fuOQSH5C1_0),.dout(w_dff_B_5ITfGVaQ2_0),.clk(gclk));
	jdff dff_B_0VD5m62i0_0(.din(w_dff_B_5ITfGVaQ2_0),.dout(w_dff_B_0VD5m62i0_0),.clk(gclk));
	jdff dff_B_not8cW135_0(.din(w_dff_B_0VD5m62i0_0),.dout(w_dff_B_not8cW135_0),.clk(gclk));
	jdff dff_B_9jvl69mj8_0(.din(w_dff_B_not8cW135_0),.dout(w_dff_B_9jvl69mj8_0),.clk(gclk));
	jdff dff_B_4TrvZjcd5_0(.din(w_dff_B_9jvl69mj8_0),.dout(w_dff_B_4TrvZjcd5_0),.clk(gclk));
	jdff dff_B_FSKLiabn8_0(.din(w_dff_B_4TrvZjcd5_0),.dout(w_dff_B_FSKLiabn8_0),.clk(gclk));
	jdff dff_B_qb8zBmN64_0(.din(w_dff_B_FSKLiabn8_0),.dout(w_dff_B_qb8zBmN64_0),.clk(gclk));
	jdff dff_B_isw0vxTt7_0(.din(w_dff_B_qb8zBmN64_0),.dout(w_dff_B_isw0vxTt7_0),.clk(gclk));
	jdff dff_B_4AHxuAkV4_0(.din(w_dff_B_isw0vxTt7_0),.dout(w_dff_B_4AHxuAkV4_0),.clk(gclk));
	jdff dff_B_SH38UfqO5_0(.din(w_dff_B_4AHxuAkV4_0),.dout(w_dff_B_SH38UfqO5_0),.clk(gclk));
	jdff dff_B_ezIRKy3t8_0(.din(w_dff_B_SH38UfqO5_0),.dout(w_dff_B_ezIRKy3t8_0),.clk(gclk));
	jdff dff_B_OCQCRQcb0_0(.din(w_dff_B_ezIRKy3t8_0),.dout(w_dff_B_OCQCRQcb0_0),.clk(gclk));
	jdff dff_B_05Kch9JF6_0(.din(w_dff_B_OCQCRQcb0_0),.dout(w_dff_B_05Kch9JF6_0),.clk(gclk));
	jdff dff_B_XO7Wi3Gt8_0(.din(w_dff_B_05Kch9JF6_0),.dout(w_dff_B_XO7Wi3Gt8_0),.clk(gclk));
	jdff dff_B_dOPWldWu1_0(.din(w_dff_B_XO7Wi3Gt8_0),.dout(w_dff_B_dOPWldWu1_0),.clk(gclk));
	jdff dff_B_u0CkkhaS3_0(.din(w_dff_B_dOPWldWu1_0),.dout(w_dff_B_u0CkkhaS3_0),.clk(gclk));
	jdff dff_B_SWGrBkMc8_0(.din(w_dff_B_u0CkkhaS3_0),.dout(w_dff_B_SWGrBkMc8_0),.clk(gclk));
	jdff dff_B_Y4tj5F2l3_0(.din(w_dff_B_SWGrBkMc8_0),.dout(w_dff_B_Y4tj5F2l3_0),.clk(gclk));
	jdff dff_B_AVhl6SGa2_0(.din(w_dff_B_Y4tj5F2l3_0),.dout(w_dff_B_AVhl6SGa2_0),.clk(gclk));
	jdff dff_B_k68Mwf0C2_0(.din(w_dff_B_AVhl6SGa2_0),.dout(w_dff_B_k68Mwf0C2_0),.clk(gclk));
	jdff dff_B_gUV6Cqb07_0(.din(w_dff_B_k68Mwf0C2_0),.dout(w_dff_B_gUV6Cqb07_0),.clk(gclk));
	jdff dff_B_uJ8bQSmx0_0(.din(w_dff_B_gUV6Cqb07_0),.dout(w_dff_B_uJ8bQSmx0_0),.clk(gclk));
	jdff dff_B_EnIhzMOw3_0(.din(w_dff_B_uJ8bQSmx0_0),.dout(w_dff_B_EnIhzMOw3_0),.clk(gclk));
	jdff dff_B_qNCpt48b4_0(.din(w_dff_B_EnIhzMOw3_0),.dout(w_dff_B_qNCpt48b4_0),.clk(gclk));
	jdff dff_B_YQu8q8eu7_0(.din(w_dff_B_qNCpt48b4_0),.dout(w_dff_B_YQu8q8eu7_0),.clk(gclk));
	jdff dff_B_QQoj9x9n2_0(.din(w_dff_B_YQu8q8eu7_0),.dout(w_dff_B_QQoj9x9n2_0),.clk(gclk));
	jdff dff_B_hccerYTj0_0(.din(w_dff_B_QQoj9x9n2_0),.dout(w_dff_B_hccerYTj0_0),.clk(gclk));
	jdff dff_B_cAvIqjhH2_0(.din(w_dff_B_hccerYTj0_0),.dout(w_dff_B_cAvIqjhH2_0),.clk(gclk));
	jdff dff_B_lvBtN87r4_0(.din(w_dff_B_cAvIqjhH2_0),.dout(w_dff_B_lvBtN87r4_0),.clk(gclk));
	jdff dff_B_N9aWi0P60_0(.din(w_dff_B_lvBtN87r4_0),.dout(w_dff_B_N9aWi0P60_0),.clk(gclk));
	jdff dff_B_srqhhSHi4_0(.din(w_dff_B_N9aWi0P60_0),.dout(w_dff_B_srqhhSHi4_0),.clk(gclk));
	jdff dff_B_nqBuXuO03_0(.din(w_dff_B_srqhhSHi4_0),.dout(w_dff_B_nqBuXuO03_0),.clk(gclk));
	jdff dff_B_8VOKdXdQ9_0(.din(w_dff_B_nqBuXuO03_0),.dout(w_dff_B_8VOKdXdQ9_0),.clk(gclk));
	jdff dff_B_OkjULAnL9_0(.din(w_dff_B_8VOKdXdQ9_0),.dout(w_dff_B_OkjULAnL9_0),.clk(gclk));
	jdff dff_B_9NJgM24b5_1(.din(n852),.dout(w_dff_B_9NJgM24b5_1),.clk(gclk));
	jdff dff_B_Ee89ZGrN4_1(.din(w_dff_B_9NJgM24b5_1),.dout(w_dff_B_Ee89ZGrN4_1),.clk(gclk));
	jdff dff_B_ZF42x9ts0_1(.din(w_dff_B_Ee89ZGrN4_1),.dout(w_dff_B_ZF42x9ts0_1),.clk(gclk));
	jdff dff_B_QjswzR6b7_1(.din(w_dff_B_ZF42x9ts0_1),.dout(w_dff_B_QjswzR6b7_1),.clk(gclk));
	jdff dff_B_Louy74bJ1_1(.din(w_dff_B_QjswzR6b7_1),.dout(w_dff_B_Louy74bJ1_1),.clk(gclk));
	jdff dff_B_KSXvOQt49_1(.din(w_dff_B_Louy74bJ1_1),.dout(w_dff_B_KSXvOQt49_1),.clk(gclk));
	jdff dff_B_vWIbbuSJ2_1(.din(w_dff_B_KSXvOQt49_1),.dout(w_dff_B_vWIbbuSJ2_1),.clk(gclk));
	jdff dff_B_FenRkLh27_1(.din(w_dff_B_vWIbbuSJ2_1),.dout(w_dff_B_FenRkLh27_1),.clk(gclk));
	jdff dff_B_26b3Zlqq7_1(.din(w_dff_B_FenRkLh27_1),.dout(w_dff_B_26b3Zlqq7_1),.clk(gclk));
	jdff dff_B_Muweay6I7_1(.din(w_dff_B_26b3Zlqq7_1),.dout(w_dff_B_Muweay6I7_1),.clk(gclk));
	jdff dff_B_CMWFYgjn0_1(.din(w_dff_B_Muweay6I7_1),.dout(w_dff_B_CMWFYgjn0_1),.clk(gclk));
	jdff dff_B_j8KqCyKQ6_1(.din(w_dff_B_CMWFYgjn0_1),.dout(w_dff_B_j8KqCyKQ6_1),.clk(gclk));
	jdff dff_B_sT0Hmm989_1(.din(w_dff_B_j8KqCyKQ6_1),.dout(w_dff_B_sT0Hmm989_1),.clk(gclk));
	jdff dff_B_tozgOeZS8_1(.din(w_dff_B_sT0Hmm989_1),.dout(w_dff_B_tozgOeZS8_1),.clk(gclk));
	jdff dff_B_Y7x8ms9G3_1(.din(w_dff_B_tozgOeZS8_1),.dout(w_dff_B_Y7x8ms9G3_1),.clk(gclk));
	jdff dff_B_bsT20mAX8_1(.din(w_dff_B_Y7x8ms9G3_1),.dout(w_dff_B_bsT20mAX8_1),.clk(gclk));
	jdff dff_B_tINAJHrN2_1(.din(w_dff_B_bsT20mAX8_1),.dout(w_dff_B_tINAJHrN2_1),.clk(gclk));
	jdff dff_B_zjO5cdOm8_1(.din(w_dff_B_tINAJHrN2_1),.dout(w_dff_B_zjO5cdOm8_1),.clk(gclk));
	jdff dff_B_4DUWaUx61_1(.din(w_dff_B_zjO5cdOm8_1),.dout(w_dff_B_4DUWaUx61_1),.clk(gclk));
	jdff dff_B_Ol3ZBT5B5_1(.din(w_dff_B_4DUWaUx61_1),.dout(w_dff_B_Ol3ZBT5B5_1),.clk(gclk));
	jdff dff_B_A1uC9sbx9_1(.din(w_dff_B_Ol3ZBT5B5_1),.dout(w_dff_B_A1uC9sbx9_1),.clk(gclk));
	jdff dff_B_pwMQRzIi0_1(.din(w_dff_B_A1uC9sbx9_1),.dout(w_dff_B_pwMQRzIi0_1),.clk(gclk));
	jdff dff_B_mjZS1bgC8_1(.din(w_dff_B_pwMQRzIi0_1),.dout(w_dff_B_mjZS1bgC8_1),.clk(gclk));
	jdff dff_B_ysFgUrBC8_1(.din(w_dff_B_mjZS1bgC8_1),.dout(w_dff_B_ysFgUrBC8_1),.clk(gclk));
	jdff dff_B_co0ctbka3_1(.din(w_dff_B_ysFgUrBC8_1),.dout(w_dff_B_co0ctbka3_1),.clk(gclk));
	jdff dff_B_iS99qmpY0_1(.din(w_dff_B_co0ctbka3_1),.dout(w_dff_B_iS99qmpY0_1),.clk(gclk));
	jdff dff_B_9VmRnF7I2_1(.din(w_dff_B_iS99qmpY0_1),.dout(w_dff_B_9VmRnF7I2_1),.clk(gclk));
	jdff dff_B_t4eQxJZH6_1(.din(w_dff_B_9VmRnF7I2_1),.dout(w_dff_B_t4eQxJZH6_1),.clk(gclk));
	jdff dff_B_XwUgOE3E5_1(.din(w_dff_B_t4eQxJZH6_1),.dout(w_dff_B_XwUgOE3E5_1),.clk(gclk));
	jdff dff_B_Nm5IPIl41_1(.din(w_dff_B_XwUgOE3E5_1),.dout(w_dff_B_Nm5IPIl41_1),.clk(gclk));
	jdff dff_B_JaKKb2p29_1(.din(w_dff_B_Nm5IPIl41_1),.dout(w_dff_B_JaKKb2p29_1),.clk(gclk));
	jdff dff_B_ICBZ6n092_1(.din(w_dff_B_JaKKb2p29_1),.dout(w_dff_B_ICBZ6n092_1),.clk(gclk));
	jdff dff_B_oo2OxxsJ1_1(.din(w_dff_B_ICBZ6n092_1),.dout(w_dff_B_oo2OxxsJ1_1),.clk(gclk));
	jdff dff_B_tTj9umva9_1(.din(w_dff_B_oo2OxxsJ1_1),.dout(w_dff_B_tTj9umva9_1),.clk(gclk));
	jdff dff_B_Wy7hGWI61_1(.din(w_dff_B_tTj9umva9_1),.dout(w_dff_B_Wy7hGWI61_1),.clk(gclk));
	jdff dff_B_IQJhi7uQ9_1(.din(w_dff_B_Wy7hGWI61_1),.dout(w_dff_B_IQJhi7uQ9_1),.clk(gclk));
	jdff dff_B_qhye2kpX3_1(.din(w_dff_B_IQJhi7uQ9_1),.dout(w_dff_B_qhye2kpX3_1),.clk(gclk));
	jdff dff_B_cVDBCvHa0_1(.din(w_dff_B_qhye2kpX3_1),.dout(w_dff_B_cVDBCvHa0_1),.clk(gclk));
	jdff dff_B_hcdN6NNH1_1(.din(w_dff_B_cVDBCvHa0_1),.dout(w_dff_B_hcdN6NNH1_1),.clk(gclk));
	jdff dff_B_52ms6wAm9_1(.din(w_dff_B_hcdN6NNH1_1),.dout(w_dff_B_52ms6wAm9_1),.clk(gclk));
	jdff dff_B_e8cBAJ450_1(.din(w_dff_B_52ms6wAm9_1),.dout(w_dff_B_e8cBAJ450_1),.clk(gclk));
	jdff dff_B_BFddvJTE7_1(.din(w_dff_B_e8cBAJ450_1),.dout(w_dff_B_BFddvJTE7_1),.clk(gclk));
	jdff dff_B_FsUz8bED2_1(.din(w_dff_B_BFddvJTE7_1),.dout(w_dff_B_FsUz8bED2_1),.clk(gclk));
	jdff dff_B_F7zOgjsA2_1(.din(w_dff_B_FsUz8bED2_1),.dout(w_dff_B_F7zOgjsA2_1),.clk(gclk));
	jdff dff_B_ed99a9fb5_1(.din(w_dff_B_F7zOgjsA2_1),.dout(w_dff_B_ed99a9fb5_1),.clk(gclk));
	jdff dff_B_901DdbOZ7_1(.din(w_dff_B_ed99a9fb5_1),.dout(w_dff_B_901DdbOZ7_1),.clk(gclk));
	jdff dff_B_NcAKWOW76_1(.din(w_dff_B_901DdbOZ7_1),.dout(w_dff_B_NcAKWOW76_1),.clk(gclk));
	jdff dff_B_45zR5xGK2_1(.din(w_dff_B_NcAKWOW76_1),.dout(w_dff_B_45zR5xGK2_1),.clk(gclk));
	jdff dff_B_O7c4UxYo3_1(.din(w_dff_B_45zR5xGK2_1),.dout(w_dff_B_O7c4UxYo3_1),.clk(gclk));
	jdff dff_B_v0LDFqJ10_1(.din(w_dff_B_O7c4UxYo3_1),.dout(w_dff_B_v0LDFqJ10_1),.clk(gclk));
	jdff dff_B_VHa9mYIA3_1(.din(w_dff_B_v0LDFqJ10_1),.dout(w_dff_B_VHa9mYIA3_1),.clk(gclk));
	jdff dff_B_ktlZVb6b6_1(.din(w_dff_B_VHa9mYIA3_1),.dout(w_dff_B_ktlZVb6b6_1),.clk(gclk));
	jdff dff_B_CGC6woTF7_1(.din(w_dff_B_ktlZVb6b6_1),.dout(w_dff_B_CGC6woTF7_1),.clk(gclk));
	jdff dff_B_40M3lrbG9_1(.din(w_dff_B_CGC6woTF7_1),.dout(w_dff_B_40M3lrbG9_1),.clk(gclk));
	jdff dff_B_EJ4RaDyY2_1(.din(w_dff_B_40M3lrbG9_1),.dout(w_dff_B_EJ4RaDyY2_1),.clk(gclk));
	jdff dff_B_PRIf5Z2A2_1(.din(w_dff_B_EJ4RaDyY2_1),.dout(w_dff_B_PRIf5Z2A2_1),.clk(gclk));
	jdff dff_B_qCgnp5tw7_1(.din(w_dff_B_PRIf5Z2A2_1),.dout(w_dff_B_qCgnp5tw7_1),.clk(gclk));
	jdff dff_B_2WZarVJq6_1(.din(w_dff_B_qCgnp5tw7_1),.dout(w_dff_B_2WZarVJq6_1),.clk(gclk));
	jdff dff_B_Lg6v5lBM4_1(.din(w_dff_B_2WZarVJq6_1),.dout(w_dff_B_Lg6v5lBM4_1),.clk(gclk));
	jdff dff_B_s43XP0Le3_1(.din(w_dff_B_Lg6v5lBM4_1),.dout(w_dff_B_s43XP0Le3_1),.clk(gclk));
	jdff dff_B_wfRhvxgL3_1(.din(w_dff_B_s43XP0Le3_1),.dout(w_dff_B_wfRhvxgL3_1),.clk(gclk));
	jdff dff_B_TndS5KXC9_1(.din(w_dff_B_wfRhvxgL3_1),.dout(w_dff_B_TndS5KXC9_1),.clk(gclk));
	jdff dff_B_r8PlXZlq0_1(.din(w_dff_B_TndS5KXC9_1),.dout(w_dff_B_r8PlXZlq0_1),.clk(gclk));
	jdff dff_B_UuuzylPH3_1(.din(w_dff_B_r8PlXZlq0_1),.dout(w_dff_B_UuuzylPH3_1),.clk(gclk));
	jdff dff_B_zftX87tM0_1(.din(w_dff_B_UuuzylPH3_1),.dout(w_dff_B_zftX87tM0_1),.clk(gclk));
	jdff dff_B_bbA0ckeX8_1(.din(w_dff_B_zftX87tM0_1),.dout(w_dff_B_bbA0ckeX8_1),.clk(gclk));
	jdff dff_B_HlBBpU5P9_1(.din(w_dff_B_bbA0ckeX8_1),.dout(w_dff_B_HlBBpU5P9_1),.clk(gclk));
	jdff dff_B_jfFDA3w71_1(.din(w_dff_B_HlBBpU5P9_1),.dout(w_dff_B_jfFDA3w71_1),.clk(gclk));
	jdff dff_B_15P4j7GD1_1(.din(w_dff_B_jfFDA3w71_1),.dout(w_dff_B_15P4j7GD1_1),.clk(gclk));
	jdff dff_B_u8RZ4i7D2_1(.din(w_dff_B_15P4j7GD1_1),.dout(w_dff_B_u8RZ4i7D2_1),.clk(gclk));
	jdff dff_B_jtXBEZHH1_1(.din(w_dff_B_u8RZ4i7D2_1),.dout(w_dff_B_jtXBEZHH1_1),.clk(gclk));
	jdff dff_B_rg7QbqaU7_1(.din(w_dff_B_jtXBEZHH1_1),.dout(w_dff_B_rg7QbqaU7_1),.clk(gclk));
	jdff dff_B_kAeLitOl4_1(.din(w_dff_B_rg7QbqaU7_1),.dout(w_dff_B_kAeLitOl4_1),.clk(gclk));
	jdff dff_B_TejR0zQI9_1(.din(w_dff_B_kAeLitOl4_1),.dout(w_dff_B_TejR0zQI9_1),.clk(gclk));
	jdff dff_B_xdTQ0fQL4_1(.din(w_dff_B_TejR0zQI9_1),.dout(w_dff_B_xdTQ0fQL4_1),.clk(gclk));
	jdff dff_B_CQwcGSaj4_1(.din(w_dff_B_xdTQ0fQL4_1),.dout(w_dff_B_CQwcGSaj4_1),.clk(gclk));
	jdff dff_B_Amfob1qH1_1(.din(w_dff_B_CQwcGSaj4_1),.dout(w_dff_B_Amfob1qH1_1),.clk(gclk));
	jdff dff_B_PPpQ5mdn1_1(.din(w_dff_B_Amfob1qH1_1),.dout(w_dff_B_PPpQ5mdn1_1),.clk(gclk));
	jdff dff_B_AKYzejYo5_0(.din(n853),.dout(w_dff_B_AKYzejYo5_0),.clk(gclk));
	jdff dff_B_7IDtgNJk7_0(.din(w_dff_B_AKYzejYo5_0),.dout(w_dff_B_7IDtgNJk7_0),.clk(gclk));
	jdff dff_B_8HrLto0e2_0(.din(w_dff_B_7IDtgNJk7_0),.dout(w_dff_B_8HrLto0e2_0),.clk(gclk));
	jdff dff_B_JpX2n4bg1_0(.din(w_dff_B_8HrLto0e2_0),.dout(w_dff_B_JpX2n4bg1_0),.clk(gclk));
	jdff dff_B_IaEbr7209_0(.din(w_dff_B_JpX2n4bg1_0),.dout(w_dff_B_IaEbr7209_0),.clk(gclk));
	jdff dff_B_nSyI0P9w4_0(.din(w_dff_B_IaEbr7209_0),.dout(w_dff_B_nSyI0P9w4_0),.clk(gclk));
	jdff dff_B_vrUairEN8_0(.din(w_dff_B_nSyI0P9w4_0),.dout(w_dff_B_vrUairEN8_0),.clk(gclk));
	jdff dff_B_wcO3udsH0_0(.din(w_dff_B_vrUairEN8_0),.dout(w_dff_B_wcO3udsH0_0),.clk(gclk));
	jdff dff_B_QMIJgd9Z3_0(.din(w_dff_B_wcO3udsH0_0),.dout(w_dff_B_QMIJgd9Z3_0),.clk(gclk));
	jdff dff_B_olCUdMbx8_0(.din(w_dff_B_QMIJgd9Z3_0),.dout(w_dff_B_olCUdMbx8_0),.clk(gclk));
	jdff dff_B_vOpYVEes8_0(.din(w_dff_B_olCUdMbx8_0),.dout(w_dff_B_vOpYVEes8_0),.clk(gclk));
	jdff dff_B_Mj2dEgYd3_0(.din(w_dff_B_vOpYVEes8_0),.dout(w_dff_B_Mj2dEgYd3_0),.clk(gclk));
	jdff dff_B_ZdScPvL71_0(.din(w_dff_B_Mj2dEgYd3_0),.dout(w_dff_B_ZdScPvL71_0),.clk(gclk));
	jdff dff_B_mtYlnKgr1_0(.din(w_dff_B_ZdScPvL71_0),.dout(w_dff_B_mtYlnKgr1_0),.clk(gclk));
	jdff dff_B_eMSlw0Pt4_0(.din(w_dff_B_mtYlnKgr1_0),.dout(w_dff_B_eMSlw0Pt4_0),.clk(gclk));
	jdff dff_B_MaRdwAHT1_0(.din(w_dff_B_eMSlw0Pt4_0),.dout(w_dff_B_MaRdwAHT1_0),.clk(gclk));
	jdff dff_B_ZmpmK7St6_0(.din(w_dff_B_MaRdwAHT1_0),.dout(w_dff_B_ZmpmK7St6_0),.clk(gclk));
	jdff dff_B_VaDQCl2Y8_0(.din(w_dff_B_ZmpmK7St6_0),.dout(w_dff_B_VaDQCl2Y8_0),.clk(gclk));
	jdff dff_B_KvghZkei9_0(.din(w_dff_B_VaDQCl2Y8_0),.dout(w_dff_B_KvghZkei9_0),.clk(gclk));
	jdff dff_B_gi1vx5sq4_0(.din(w_dff_B_KvghZkei9_0),.dout(w_dff_B_gi1vx5sq4_0),.clk(gclk));
	jdff dff_B_7EnuHvxh9_0(.din(w_dff_B_gi1vx5sq4_0),.dout(w_dff_B_7EnuHvxh9_0),.clk(gclk));
	jdff dff_B_qwhUHJDk8_0(.din(w_dff_B_7EnuHvxh9_0),.dout(w_dff_B_qwhUHJDk8_0),.clk(gclk));
	jdff dff_B_xpLm7AOd1_0(.din(w_dff_B_qwhUHJDk8_0),.dout(w_dff_B_xpLm7AOd1_0),.clk(gclk));
	jdff dff_B_37slPqMN9_0(.din(w_dff_B_xpLm7AOd1_0),.dout(w_dff_B_37slPqMN9_0),.clk(gclk));
	jdff dff_B_gtWRKnly7_0(.din(w_dff_B_37slPqMN9_0),.dout(w_dff_B_gtWRKnly7_0),.clk(gclk));
	jdff dff_B_gECJYpll1_0(.din(w_dff_B_gtWRKnly7_0),.dout(w_dff_B_gECJYpll1_0),.clk(gclk));
	jdff dff_B_I4muCoFR5_0(.din(w_dff_B_gECJYpll1_0),.dout(w_dff_B_I4muCoFR5_0),.clk(gclk));
	jdff dff_B_3Vo90gVp6_0(.din(w_dff_B_I4muCoFR5_0),.dout(w_dff_B_3Vo90gVp6_0),.clk(gclk));
	jdff dff_B_J97ykhr25_0(.din(w_dff_B_3Vo90gVp6_0),.dout(w_dff_B_J97ykhr25_0),.clk(gclk));
	jdff dff_B_lhCECIPs9_0(.din(w_dff_B_J97ykhr25_0),.dout(w_dff_B_lhCECIPs9_0),.clk(gclk));
	jdff dff_B_Af5AdqYE5_0(.din(w_dff_B_lhCECIPs9_0),.dout(w_dff_B_Af5AdqYE5_0),.clk(gclk));
	jdff dff_B_p88eS73Q0_0(.din(w_dff_B_Af5AdqYE5_0),.dout(w_dff_B_p88eS73Q0_0),.clk(gclk));
	jdff dff_B_H7hjs9Kc4_0(.din(w_dff_B_p88eS73Q0_0),.dout(w_dff_B_H7hjs9Kc4_0),.clk(gclk));
	jdff dff_B_gkb9CDrm3_0(.din(w_dff_B_H7hjs9Kc4_0),.dout(w_dff_B_gkb9CDrm3_0),.clk(gclk));
	jdff dff_B_aIyQQONY1_0(.din(w_dff_B_gkb9CDrm3_0),.dout(w_dff_B_aIyQQONY1_0),.clk(gclk));
	jdff dff_B_HrQm4c5a8_0(.din(w_dff_B_aIyQQONY1_0),.dout(w_dff_B_HrQm4c5a8_0),.clk(gclk));
	jdff dff_B_wvS1Pqwl2_0(.din(w_dff_B_HrQm4c5a8_0),.dout(w_dff_B_wvS1Pqwl2_0),.clk(gclk));
	jdff dff_B_oYJAh0cj9_0(.din(w_dff_B_wvS1Pqwl2_0),.dout(w_dff_B_oYJAh0cj9_0),.clk(gclk));
	jdff dff_B_gDE3kUwP1_0(.din(w_dff_B_oYJAh0cj9_0),.dout(w_dff_B_gDE3kUwP1_0),.clk(gclk));
	jdff dff_B_IpocvKzj5_0(.din(w_dff_B_gDE3kUwP1_0),.dout(w_dff_B_IpocvKzj5_0),.clk(gclk));
	jdff dff_B_hMYQshit6_0(.din(w_dff_B_IpocvKzj5_0),.dout(w_dff_B_hMYQshit6_0),.clk(gclk));
	jdff dff_B_vvfUGRbh0_0(.din(w_dff_B_hMYQshit6_0),.dout(w_dff_B_vvfUGRbh0_0),.clk(gclk));
	jdff dff_B_stdu2BJX2_0(.din(w_dff_B_vvfUGRbh0_0),.dout(w_dff_B_stdu2BJX2_0),.clk(gclk));
	jdff dff_B_4rpeBBVQ0_0(.din(w_dff_B_stdu2BJX2_0),.dout(w_dff_B_4rpeBBVQ0_0),.clk(gclk));
	jdff dff_B_hEZrfaVQ7_0(.din(w_dff_B_4rpeBBVQ0_0),.dout(w_dff_B_hEZrfaVQ7_0),.clk(gclk));
	jdff dff_B_dk8Gjgog4_0(.din(w_dff_B_hEZrfaVQ7_0),.dout(w_dff_B_dk8Gjgog4_0),.clk(gclk));
	jdff dff_B_i2eCqOGc5_0(.din(w_dff_B_dk8Gjgog4_0),.dout(w_dff_B_i2eCqOGc5_0),.clk(gclk));
	jdff dff_B_BolPvYss6_0(.din(w_dff_B_i2eCqOGc5_0),.dout(w_dff_B_BolPvYss6_0),.clk(gclk));
	jdff dff_B_uoqHmwnq3_0(.din(w_dff_B_BolPvYss6_0),.dout(w_dff_B_uoqHmwnq3_0),.clk(gclk));
	jdff dff_B_iMLRkoUN5_0(.din(w_dff_B_uoqHmwnq3_0),.dout(w_dff_B_iMLRkoUN5_0),.clk(gclk));
	jdff dff_B_QIBLQZZa0_0(.din(w_dff_B_iMLRkoUN5_0),.dout(w_dff_B_QIBLQZZa0_0),.clk(gclk));
	jdff dff_B_bFJKcIP87_0(.din(w_dff_B_QIBLQZZa0_0),.dout(w_dff_B_bFJKcIP87_0),.clk(gclk));
	jdff dff_B_lhZFRcmq9_0(.din(w_dff_B_bFJKcIP87_0),.dout(w_dff_B_lhZFRcmq9_0),.clk(gclk));
	jdff dff_B_z6rvqgCH2_0(.din(w_dff_B_lhZFRcmq9_0),.dout(w_dff_B_z6rvqgCH2_0),.clk(gclk));
	jdff dff_B_oQcsgDTN6_0(.din(w_dff_B_z6rvqgCH2_0),.dout(w_dff_B_oQcsgDTN6_0),.clk(gclk));
	jdff dff_B_qPjFxPqP6_0(.din(w_dff_B_oQcsgDTN6_0),.dout(w_dff_B_qPjFxPqP6_0),.clk(gclk));
	jdff dff_B_cfFdhhoE2_0(.din(w_dff_B_qPjFxPqP6_0),.dout(w_dff_B_cfFdhhoE2_0),.clk(gclk));
	jdff dff_B_18yjfYTz5_0(.din(w_dff_B_cfFdhhoE2_0),.dout(w_dff_B_18yjfYTz5_0),.clk(gclk));
	jdff dff_B_jsRJJOYz8_0(.din(w_dff_B_18yjfYTz5_0),.dout(w_dff_B_jsRJJOYz8_0),.clk(gclk));
	jdff dff_B_5xgLIorn9_0(.din(w_dff_B_jsRJJOYz8_0),.dout(w_dff_B_5xgLIorn9_0),.clk(gclk));
	jdff dff_B_mmH7ljqM2_0(.din(w_dff_B_5xgLIorn9_0),.dout(w_dff_B_mmH7ljqM2_0),.clk(gclk));
	jdff dff_B_qA1OOnNy6_0(.din(w_dff_B_mmH7ljqM2_0),.dout(w_dff_B_qA1OOnNy6_0),.clk(gclk));
	jdff dff_B_QcxskTGc8_0(.din(w_dff_B_qA1OOnNy6_0),.dout(w_dff_B_QcxskTGc8_0),.clk(gclk));
	jdff dff_B_MPlmTR1w1_0(.din(w_dff_B_QcxskTGc8_0),.dout(w_dff_B_MPlmTR1w1_0),.clk(gclk));
	jdff dff_B_seD2LrPD7_0(.din(w_dff_B_MPlmTR1w1_0),.dout(w_dff_B_seD2LrPD7_0),.clk(gclk));
	jdff dff_B_2s0OEdS27_0(.din(w_dff_B_seD2LrPD7_0),.dout(w_dff_B_2s0OEdS27_0),.clk(gclk));
	jdff dff_B_4OOlJfPb9_0(.din(w_dff_B_2s0OEdS27_0),.dout(w_dff_B_4OOlJfPb9_0),.clk(gclk));
	jdff dff_B_sE3eZfIE4_0(.din(w_dff_B_4OOlJfPb9_0),.dout(w_dff_B_sE3eZfIE4_0),.clk(gclk));
	jdff dff_B_whJyrNNb9_0(.din(w_dff_B_sE3eZfIE4_0),.dout(w_dff_B_whJyrNNb9_0),.clk(gclk));
	jdff dff_B_fgDz39rj3_0(.din(w_dff_B_whJyrNNb9_0),.dout(w_dff_B_fgDz39rj3_0),.clk(gclk));
	jdff dff_B_c5MKNbQr9_0(.din(w_dff_B_fgDz39rj3_0),.dout(w_dff_B_c5MKNbQr9_0),.clk(gclk));
	jdff dff_B_1dUNJKul3_0(.din(w_dff_B_c5MKNbQr9_0),.dout(w_dff_B_1dUNJKul3_0),.clk(gclk));
	jdff dff_B_vSJ6okrh6_0(.din(w_dff_B_1dUNJKul3_0),.dout(w_dff_B_vSJ6okrh6_0),.clk(gclk));
	jdff dff_B_7HOhPr9F3_0(.din(w_dff_B_vSJ6okrh6_0),.dout(w_dff_B_7HOhPr9F3_0),.clk(gclk));
	jdff dff_B_eDTMfV4R7_0(.din(w_dff_B_7HOhPr9F3_0),.dout(w_dff_B_eDTMfV4R7_0),.clk(gclk));
	jdff dff_B_7OfKxHUE9_0(.din(w_dff_B_eDTMfV4R7_0),.dout(w_dff_B_7OfKxHUE9_0),.clk(gclk));
	jdff dff_B_OAi2xSZU9_0(.din(w_dff_B_7OfKxHUE9_0),.dout(w_dff_B_OAi2xSZU9_0),.clk(gclk));
	jdff dff_B_nx8MnoHd2_0(.din(w_dff_B_OAi2xSZU9_0),.dout(w_dff_B_nx8MnoHd2_0),.clk(gclk));
	jdff dff_B_lCknWwrj8_1(.din(n846),.dout(w_dff_B_lCknWwrj8_1),.clk(gclk));
	jdff dff_B_xZsUVpB96_1(.din(w_dff_B_lCknWwrj8_1),.dout(w_dff_B_xZsUVpB96_1),.clk(gclk));
	jdff dff_B_OdyCepR85_1(.din(w_dff_B_xZsUVpB96_1),.dout(w_dff_B_OdyCepR85_1),.clk(gclk));
	jdff dff_B_TdQA974I2_1(.din(w_dff_B_OdyCepR85_1),.dout(w_dff_B_TdQA974I2_1),.clk(gclk));
	jdff dff_B_1OLK7WvQ2_1(.din(w_dff_B_TdQA974I2_1),.dout(w_dff_B_1OLK7WvQ2_1),.clk(gclk));
	jdff dff_B_QRCLJIzF2_1(.din(w_dff_B_1OLK7WvQ2_1),.dout(w_dff_B_QRCLJIzF2_1),.clk(gclk));
	jdff dff_B_zgky6dEv8_1(.din(w_dff_B_QRCLJIzF2_1),.dout(w_dff_B_zgky6dEv8_1),.clk(gclk));
	jdff dff_B_FGEnxrmt2_1(.din(w_dff_B_zgky6dEv8_1),.dout(w_dff_B_FGEnxrmt2_1),.clk(gclk));
	jdff dff_B_iHU1lMPN3_1(.din(w_dff_B_FGEnxrmt2_1),.dout(w_dff_B_iHU1lMPN3_1),.clk(gclk));
	jdff dff_B_JdgEoIGi3_1(.din(w_dff_B_iHU1lMPN3_1),.dout(w_dff_B_JdgEoIGi3_1),.clk(gclk));
	jdff dff_B_vbCn5soC4_1(.din(w_dff_B_JdgEoIGi3_1),.dout(w_dff_B_vbCn5soC4_1),.clk(gclk));
	jdff dff_B_pwwNt5c28_1(.din(w_dff_B_vbCn5soC4_1),.dout(w_dff_B_pwwNt5c28_1),.clk(gclk));
	jdff dff_B_ROq1uc8L7_1(.din(w_dff_B_pwwNt5c28_1),.dout(w_dff_B_ROq1uc8L7_1),.clk(gclk));
	jdff dff_B_MurowAlE7_1(.din(w_dff_B_ROq1uc8L7_1),.dout(w_dff_B_MurowAlE7_1),.clk(gclk));
	jdff dff_B_6XfR9vIt1_1(.din(w_dff_B_MurowAlE7_1),.dout(w_dff_B_6XfR9vIt1_1),.clk(gclk));
	jdff dff_B_WXvnlxJT5_1(.din(w_dff_B_6XfR9vIt1_1),.dout(w_dff_B_WXvnlxJT5_1),.clk(gclk));
	jdff dff_B_yaRblRQ46_1(.din(w_dff_B_WXvnlxJT5_1),.dout(w_dff_B_yaRblRQ46_1),.clk(gclk));
	jdff dff_B_DIohpfQV5_1(.din(w_dff_B_yaRblRQ46_1),.dout(w_dff_B_DIohpfQV5_1),.clk(gclk));
	jdff dff_B_YvKgTTZQ7_1(.din(w_dff_B_DIohpfQV5_1),.dout(w_dff_B_YvKgTTZQ7_1),.clk(gclk));
	jdff dff_B_kG1QNLdi9_1(.din(w_dff_B_YvKgTTZQ7_1),.dout(w_dff_B_kG1QNLdi9_1),.clk(gclk));
	jdff dff_B_sXuXqJmA8_1(.din(w_dff_B_kG1QNLdi9_1),.dout(w_dff_B_sXuXqJmA8_1),.clk(gclk));
	jdff dff_B_iNq0GzVs2_1(.din(w_dff_B_sXuXqJmA8_1),.dout(w_dff_B_iNq0GzVs2_1),.clk(gclk));
	jdff dff_B_fXK9lR2Q4_1(.din(w_dff_B_iNq0GzVs2_1),.dout(w_dff_B_fXK9lR2Q4_1),.clk(gclk));
	jdff dff_B_LvndWEaJ3_1(.din(w_dff_B_fXK9lR2Q4_1),.dout(w_dff_B_LvndWEaJ3_1),.clk(gclk));
	jdff dff_B_H74PVpH53_1(.din(w_dff_B_LvndWEaJ3_1),.dout(w_dff_B_H74PVpH53_1),.clk(gclk));
	jdff dff_B_8qyhmj779_1(.din(w_dff_B_H74PVpH53_1),.dout(w_dff_B_8qyhmj779_1),.clk(gclk));
	jdff dff_B_LlZHsgZg7_1(.din(w_dff_B_8qyhmj779_1),.dout(w_dff_B_LlZHsgZg7_1),.clk(gclk));
	jdff dff_B_vnR7Vhd15_1(.din(w_dff_B_LlZHsgZg7_1),.dout(w_dff_B_vnR7Vhd15_1),.clk(gclk));
	jdff dff_B_hJS2rmOb2_1(.din(w_dff_B_vnR7Vhd15_1),.dout(w_dff_B_hJS2rmOb2_1),.clk(gclk));
	jdff dff_B_lPCprq4y1_1(.din(w_dff_B_hJS2rmOb2_1),.dout(w_dff_B_lPCprq4y1_1),.clk(gclk));
	jdff dff_B_JwWZkULi6_1(.din(w_dff_B_lPCprq4y1_1),.dout(w_dff_B_JwWZkULi6_1),.clk(gclk));
	jdff dff_B_T1QzJsnp7_1(.din(w_dff_B_JwWZkULi6_1),.dout(w_dff_B_T1QzJsnp7_1),.clk(gclk));
	jdff dff_B_yuMrqQsK6_1(.din(w_dff_B_T1QzJsnp7_1),.dout(w_dff_B_yuMrqQsK6_1),.clk(gclk));
	jdff dff_B_hFX3SBAr1_1(.din(w_dff_B_yuMrqQsK6_1),.dout(w_dff_B_hFX3SBAr1_1),.clk(gclk));
	jdff dff_B_VvxhphEV2_1(.din(w_dff_B_hFX3SBAr1_1),.dout(w_dff_B_VvxhphEV2_1),.clk(gclk));
	jdff dff_B_KP6iEftl2_1(.din(w_dff_B_VvxhphEV2_1),.dout(w_dff_B_KP6iEftl2_1),.clk(gclk));
	jdff dff_B_wHB3vvVW5_1(.din(w_dff_B_KP6iEftl2_1),.dout(w_dff_B_wHB3vvVW5_1),.clk(gclk));
	jdff dff_B_bQ9tjdIx0_1(.din(w_dff_B_wHB3vvVW5_1),.dout(w_dff_B_bQ9tjdIx0_1),.clk(gclk));
	jdff dff_B_rXxfZgr74_1(.din(w_dff_B_bQ9tjdIx0_1),.dout(w_dff_B_rXxfZgr74_1),.clk(gclk));
	jdff dff_B_0l0nvwRK1_1(.din(w_dff_B_rXxfZgr74_1),.dout(w_dff_B_0l0nvwRK1_1),.clk(gclk));
	jdff dff_B_knOUVsni5_1(.din(w_dff_B_0l0nvwRK1_1),.dout(w_dff_B_knOUVsni5_1),.clk(gclk));
	jdff dff_B_ANDRZreF6_1(.din(w_dff_B_knOUVsni5_1),.dout(w_dff_B_ANDRZreF6_1),.clk(gclk));
	jdff dff_B_it1pg5m83_1(.din(w_dff_B_ANDRZreF6_1),.dout(w_dff_B_it1pg5m83_1),.clk(gclk));
	jdff dff_B_T6y7wXMy3_1(.din(w_dff_B_it1pg5m83_1),.dout(w_dff_B_T6y7wXMy3_1),.clk(gclk));
	jdff dff_B_eUYgLd0Z4_1(.din(w_dff_B_T6y7wXMy3_1),.dout(w_dff_B_eUYgLd0Z4_1),.clk(gclk));
	jdff dff_B_Q01jJjEK7_1(.din(w_dff_B_eUYgLd0Z4_1),.dout(w_dff_B_Q01jJjEK7_1),.clk(gclk));
	jdff dff_B_jI1RE9so4_1(.din(w_dff_B_Q01jJjEK7_1),.dout(w_dff_B_jI1RE9so4_1),.clk(gclk));
	jdff dff_B_uQNoylBf7_1(.din(w_dff_B_jI1RE9so4_1),.dout(w_dff_B_uQNoylBf7_1),.clk(gclk));
	jdff dff_B_i6FkjAbK9_1(.din(w_dff_B_uQNoylBf7_1),.dout(w_dff_B_i6FkjAbK9_1),.clk(gclk));
	jdff dff_B_jKzmRNqQ0_1(.din(w_dff_B_i6FkjAbK9_1),.dout(w_dff_B_jKzmRNqQ0_1),.clk(gclk));
	jdff dff_B_4FQAICTw7_1(.din(w_dff_B_jKzmRNqQ0_1),.dout(w_dff_B_4FQAICTw7_1),.clk(gclk));
	jdff dff_B_nYL3Nx2S9_1(.din(w_dff_B_4FQAICTw7_1),.dout(w_dff_B_nYL3Nx2S9_1),.clk(gclk));
	jdff dff_B_WENE3vIV8_1(.din(w_dff_B_nYL3Nx2S9_1),.dout(w_dff_B_WENE3vIV8_1),.clk(gclk));
	jdff dff_B_qxrqIai26_1(.din(w_dff_B_WENE3vIV8_1),.dout(w_dff_B_qxrqIai26_1),.clk(gclk));
	jdff dff_B_EffnkreD7_1(.din(w_dff_B_qxrqIai26_1),.dout(w_dff_B_EffnkreD7_1),.clk(gclk));
	jdff dff_B_QNB56xWq6_1(.din(w_dff_B_EffnkreD7_1),.dout(w_dff_B_QNB56xWq6_1),.clk(gclk));
	jdff dff_B_r5AYdCqd9_1(.din(w_dff_B_QNB56xWq6_1),.dout(w_dff_B_r5AYdCqd9_1),.clk(gclk));
	jdff dff_B_2YAzXdR91_1(.din(w_dff_B_r5AYdCqd9_1),.dout(w_dff_B_2YAzXdR91_1),.clk(gclk));
	jdff dff_B_cMVQaYHH7_1(.din(w_dff_B_2YAzXdR91_1),.dout(w_dff_B_cMVQaYHH7_1),.clk(gclk));
	jdff dff_B_Qyq5nCpg1_1(.din(w_dff_B_cMVQaYHH7_1),.dout(w_dff_B_Qyq5nCpg1_1),.clk(gclk));
	jdff dff_B_3sp0g04m1_1(.din(w_dff_B_Qyq5nCpg1_1),.dout(w_dff_B_3sp0g04m1_1),.clk(gclk));
	jdff dff_B_tpDNhVmN3_1(.din(w_dff_B_3sp0g04m1_1),.dout(w_dff_B_tpDNhVmN3_1),.clk(gclk));
	jdff dff_B_WYLn8ZGZ6_1(.din(w_dff_B_tpDNhVmN3_1),.dout(w_dff_B_WYLn8ZGZ6_1),.clk(gclk));
	jdff dff_B_GYHJmo1p7_1(.din(w_dff_B_WYLn8ZGZ6_1),.dout(w_dff_B_GYHJmo1p7_1),.clk(gclk));
	jdff dff_B_BDprvJWN4_1(.din(w_dff_B_GYHJmo1p7_1),.dout(w_dff_B_BDprvJWN4_1),.clk(gclk));
	jdff dff_B_o8C8aFx62_1(.din(w_dff_B_BDprvJWN4_1),.dout(w_dff_B_o8C8aFx62_1),.clk(gclk));
	jdff dff_B_gYgMndHP4_1(.din(w_dff_B_o8C8aFx62_1),.dout(w_dff_B_gYgMndHP4_1),.clk(gclk));
	jdff dff_B_2iKCVqqj6_1(.din(w_dff_B_gYgMndHP4_1),.dout(w_dff_B_2iKCVqqj6_1),.clk(gclk));
	jdff dff_B_IDPg7c2D3_1(.din(w_dff_B_2iKCVqqj6_1),.dout(w_dff_B_IDPg7c2D3_1),.clk(gclk));
	jdff dff_B_UrHN7OS58_1(.din(w_dff_B_IDPg7c2D3_1),.dout(w_dff_B_UrHN7OS58_1),.clk(gclk));
	jdff dff_B_tKxokccA5_1(.din(w_dff_B_UrHN7OS58_1),.dout(w_dff_B_tKxokccA5_1),.clk(gclk));
	jdff dff_B_9jxuSUNa7_1(.din(w_dff_B_tKxokccA5_1),.dout(w_dff_B_9jxuSUNa7_1),.clk(gclk));
	jdff dff_B_GCQ35GD83_1(.din(w_dff_B_9jxuSUNa7_1),.dout(w_dff_B_GCQ35GD83_1),.clk(gclk));
	jdff dff_B_EBMD30yN5_1(.din(w_dff_B_GCQ35GD83_1),.dout(w_dff_B_EBMD30yN5_1),.clk(gclk));
	jdff dff_B_oI973qly7_1(.din(w_dff_B_EBMD30yN5_1),.dout(w_dff_B_oI973qly7_1),.clk(gclk));
	jdff dff_B_jqQA2aqk2_1(.din(w_dff_B_oI973qly7_1),.dout(w_dff_B_jqQA2aqk2_1),.clk(gclk));
	jdff dff_B_HA2BJTtt9_1(.din(w_dff_B_jqQA2aqk2_1),.dout(w_dff_B_HA2BJTtt9_1),.clk(gclk));
	jdff dff_B_8pR5AibF7_0(.din(n847),.dout(w_dff_B_8pR5AibF7_0),.clk(gclk));
	jdff dff_B_PTgSigU62_0(.din(w_dff_B_8pR5AibF7_0),.dout(w_dff_B_PTgSigU62_0),.clk(gclk));
	jdff dff_B_XbVtRYNq9_0(.din(w_dff_B_PTgSigU62_0),.dout(w_dff_B_XbVtRYNq9_0),.clk(gclk));
	jdff dff_B_Rt1ZJNqG2_0(.din(w_dff_B_XbVtRYNq9_0),.dout(w_dff_B_Rt1ZJNqG2_0),.clk(gclk));
	jdff dff_B_vbS1gE4f5_0(.din(w_dff_B_Rt1ZJNqG2_0),.dout(w_dff_B_vbS1gE4f5_0),.clk(gclk));
	jdff dff_B_ezEXvfl51_0(.din(w_dff_B_vbS1gE4f5_0),.dout(w_dff_B_ezEXvfl51_0),.clk(gclk));
	jdff dff_B_d37Hi4Od5_0(.din(w_dff_B_ezEXvfl51_0),.dout(w_dff_B_d37Hi4Od5_0),.clk(gclk));
	jdff dff_B_IO1WzdKW2_0(.din(w_dff_B_d37Hi4Od5_0),.dout(w_dff_B_IO1WzdKW2_0),.clk(gclk));
	jdff dff_B_SEyXEGbi5_0(.din(w_dff_B_IO1WzdKW2_0),.dout(w_dff_B_SEyXEGbi5_0),.clk(gclk));
	jdff dff_B_888l08rT3_0(.din(w_dff_B_SEyXEGbi5_0),.dout(w_dff_B_888l08rT3_0),.clk(gclk));
	jdff dff_B_1irBXwd25_0(.din(w_dff_B_888l08rT3_0),.dout(w_dff_B_1irBXwd25_0),.clk(gclk));
	jdff dff_B_Lvej4ssC6_0(.din(w_dff_B_1irBXwd25_0),.dout(w_dff_B_Lvej4ssC6_0),.clk(gclk));
	jdff dff_B_j8jljDa79_0(.din(w_dff_B_Lvej4ssC6_0),.dout(w_dff_B_j8jljDa79_0),.clk(gclk));
	jdff dff_B_3RhFFOSC6_0(.din(w_dff_B_j8jljDa79_0),.dout(w_dff_B_3RhFFOSC6_0),.clk(gclk));
	jdff dff_B_4JDAeqte3_0(.din(w_dff_B_3RhFFOSC6_0),.dout(w_dff_B_4JDAeqte3_0),.clk(gclk));
	jdff dff_B_iWkEtxVz3_0(.din(w_dff_B_4JDAeqte3_0),.dout(w_dff_B_iWkEtxVz3_0),.clk(gclk));
	jdff dff_B_yaX44PMA7_0(.din(w_dff_B_iWkEtxVz3_0),.dout(w_dff_B_yaX44PMA7_0),.clk(gclk));
	jdff dff_B_k3pIdAEr1_0(.din(w_dff_B_yaX44PMA7_0),.dout(w_dff_B_k3pIdAEr1_0),.clk(gclk));
	jdff dff_B_LD2sgsV22_0(.din(w_dff_B_k3pIdAEr1_0),.dout(w_dff_B_LD2sgsV22_0),.clk(gclk));
	jdff dff_B_ufiDitnS4_0(.din(w_dff_B_LD2sgsV22_0),.dout(w_dff_B_ufiDitnS4_0),.clk(gclk));
	jdff dff_B_OhJ9YZ951_0(.din(w_dff_B_ufiDitnS4_0),.dout(w_dff_B_OhJ9YZ951_0),.clk(gclk));
	jdff dff_B_74CaXz5Z5_0(.din(w_dff_B_OhJ9YZ951_0),.dout(w_dff_B_74CaXz5Z5_0),.clk(gclk));
	jdff dff_B_DOQQAgLu4_0(.din(w_dff_B_74CaXz5Z5_0),.dout(w_dff_B_DOQQAgLu4_0),.clk(gclk));
	jdff dff_B_dsp8lnif5_0(.din(w_dff_B_DOQQAgLu4_0),.dout(w_dff_B_dsp8lnif5_0),.clk(gclk));
	jdff dff_B_aAp71gpb7_0(.din(w_dff_B_dsp8lnif5_0),.dout(w_dff_B_aAp71gpb7_0),.clk(gclk));
	jdff dff_B_T0LA9Nw03_0(.din(w_dff_B_aAp71gpb7_0),.dout(w_dff_B_T0LA9Nw03_0),.clk(gclk));
	jdff dff_B_10nzDHj67_0(.din(w_dff_B_T0LA9Nw03_0),.dout(w_dff_B_10nzDHj67_0),.clk(gclk));
	jdff dff_B_DahEASI98_0(.din(w_dff_B_10nzDHj67_0),.dout(w_dff_B_DahEASI98_0),.clk(gclk));
	jdff dff_B_C5OsTMEn8_0(.din(w_dff_B_DahEASI98_0),.dout(w_dff_B_C5OsTMEn8_0),.clk(gclk));
	jdff dff_B_bLvUkQ5E1_0(.din(w_dff_B_C5OsTMEn8_0),.dout(w_dff_B_bLvUkQ5E1_0),.clk(gclk));
	jdff dff_B_afsvWgQ33_0(.din(w_dff_B_bLvUkQ5E1_0),.dout(w_dff_B_afsvWgQ33_0),.clk(gclk));
	jdff dff_B_KXhgsZnd3_0(.din(w_dff_B_afsvWgQ33_0),.dout(w_dff_B_KXhgsZnd3_0),.clk(gclk));
	jdff dff_B_x37VCLaJ0_0(.din(w_dff_B_KXhgsZnd3_0),.dout(w_dff_B_x37VCLaJ0_0),.clk(gclk));
	jdff dff_B_fjmfZY1A0_0(.din(w_dff_B_x37VCLaJ0_0),.dout(w_dff_B_fjmfZY1A0_0),.clk(gclk));
	jdff dff_B_In4uh2SE9_0(.din(w_dff_B_fjmfZY1A0_0),.dout(w_dff_B_In4uh2SE9_0),.clk(gclk));
	jdff dff_B_fH5HQvAi4_0(.din(w_dff_B_In4uh2SE9_0),.dout(w_dff_B_fH5HQvAi4_0),.clk(gclk));
	jdff dff_B_dVSyXFwA2_0(.din(w_dff_B_fH5HQvAi4_0),.dout(w_dff_B_dVSyXFwA2_0),.clk(gclk));
	jdff dff_B_F18WAuQ17_0(.din(w_dff_B_dVSyXFwA2_0),.dout(w_dff_B_F18WAuQ17_0),.clk(gclk));
	jdff dff_B_RxYBCtvV6_0(.din(w_dff_B_F18WAuQ17_0),.dout(w_dff_B_RxYBCtvV6_0),.clk(gclk));
	jdff dff_B_DeLRJMnl2_0(.din(w_dff_B_RxYBCtvV6_0),.dout(w_dff_B_DeLRJMnl2_0),.clk(gclk));
	jdff dff_B_BaBZuiMe0_0(.din(w_dff_B_DeLRJMnl2_0),.dout(w_dff_B_BaBZuiMe0_0),.clk(gclk));
	jdff dff_B_zFfxEav43_0(.din(w_dff_B_BaBZuiMe0_0),.dout(w_dff_B_zFfxEav43_0),.clk(gclk));
	jdff dff_B_cKbfnsVF5_0(.din(w_dff_B_zFfxEav43_0),.dout(w_dff_B_cKbfnsVF5_0),.clk(gclk));
	jdff dff_B_QoErXhUF6_0(.din(w_dff_B_cKbfnsVF5_0),.dout(w_dff_B_QoErXhUF6_0),.clk(gclk));
	jdff dff_B_ab9VWgkK0_0(.din(w_dff_B_QoErXhUF6_0),.dout(w_dff_B_ab9VWgkK0_0),.clk(gclk));
	jdff dff_B_3NTnxzKy3_0(.din(w_dff_B_ab9VWgkK0_0),.dout(w_dff_B_3NTnxzKy3_0),.clk(gclk));
	jdff dff_B_lMaiTyyr7_0(.din(w_dff_B_3NTnxzKy3_0),.dout(w_dff_B_lMaiTyyr7_0),.clk(gclk));
	jdff dff_B_tRYKaLhl0_0(.din(w_dff_B_lMaiTyyr7_0),.dout(w_dff_B_tRYKaLhl0_0),.clk(gclk));
	jdff dff_B_XIlI9xkP5_0(.din(w_dff_B_tRYKaLhl0_0),.dout(w_dff_B_XIlI9xkP5_0),.clk(gclk));
	jdff dff_B_RSF77Hhi8_0(.din(w_dff_B_XIlI9xkP5_0),.dout(w_dff_B_RSF77Hhi8_0),.clk(gclk));
	jdff dff_B_jqJrSM7f2_0(.din(w_dff_B_RSF77Hhi8_0),.dout(w_dff_B_jqJrSM7f2_0),.clk(gclk));
	jdff dff_B_MRsiVjKc1_0(.din(w_dff_B_jqJrSM7f2_0),.dout(w_dff_B_MRsiVjKc1_0),.clk(gclk));
	jdff dff_B_ZXbgPzE16_0(.din(w_dff_B_MRsiVjKc1_0),.dout(w_dff_B_ZXbgPzE16_0),.clk(gclk));
	jdff dff_B_odyB82xQ8_0(.din(w_dff_B_ZXbgPzE16_0),.dout(w_dff_B_odyB82xQ8_0),.clk(gclk));
	jdff dff_B_Jm9rZfzg2_0(.din(w_dff_B_odyB82xQ8_0),.dout(w_dff_B_Jm9rZfzg2_0),.clk(gclk));
	jdff dff_B_E3fYC9Lc7_0(.din(w_dff_B_Jm9rZfzg2_0),.dout(w_dff_B_E3fYC9Lc7_0),.clk(gclk));
	jdff dff_B_OZmjox1e6_0(.din(w_dff_B_E3fYC9Lc7_0),.dout(w_dff_B_OZmjox1e6_0),.clk(gclk));
	jdff dff_B_0DRsR5bf0_0(.din(w_dff_B_OZmjox1e6_0),.dout(w_dff_B_0DRsR5bf0_0),.clk(gclk));
	jdff dff_B_ktgXCOXu0_0(.din(w_dff_B_0DRsR5bf0_0),.dout(w_dff_B_ktgXCOXu0_0),.clk(gclk));
	jdff dff_B_IbSg46bX1_0(.din(w_dff_B_ktgXCOXu0_0),.dout(w_dff_B_IbSg46bX1_0),.clk(gclk));
	jdff dff_B_QBBQkVIG8_0(.din(w_dff_B_IbSg46bX1_0),.dout(w_dff_B_QBBQkVIG8_0),.clk(gclk));
	jdff dff_B_J6L1RD5k0_0(.din(w_dff_B_QBBQkVIG8_0),.dout(w_dff_B_J6L1RD5k0_0),.clk(gclk));
	jdff dff_B_uzcBvMxk0_0(.din(w_dff_B_J6L1RD5k0_0),.dout(w_dff_B_uzcBvMxk0_0),.clk(gclk));
	jdff dff_B_JKpHx7LD2_0(.din(w_dff_B_uzcBvMxk0_0),.dout(w_dff_B_JKpHx7LD2_0),.clk(gclk));
	jdff dff_B_ma2r9Cls1_0(.din(w_dff_B_JKpHx7LD2_0),.dout(w_dff_B_ma2r9Cls1_0),.clk(gclk));
	jdff dff_B_kgpuzd063_0(.din(w_dff_B_ma2r9Cls1_0),.dout(w_dff_B_kgpuzd063_0),.clk(gclk));
	jdff dff_B_h483iYpH0_0(.din(w_dff_B_kgpuzd063_0),.dout(w_dff_B_h483iYpH0_0),.clk(gclk));
	jdff dff_B_LDmWxb6H9_0(.din(w_dff_B_h483iYpH0_0),.dout(w_dff_B_LDmWxb6H9_0),.clk(gclk));
	jdff dff_B_sZwG3PZS6_0(.din(w_dff_B_LDmWxb6H9_0),.dout(w_dff_B_sZwG3PZS6_0),.clk(gclk));
	jdff dff_B_K19q3U5j0_0(.din(w_dff_B_sZwG3PZS6_0),.dout(w_dff_B_K19q3U5j0_0),.clk(gclk));
	jdff dff_B_SfYFSYlY8_0(.din(w_dff_B_K19q3U5j0_0),.dout(w_dff_B_SfYFSYlY8_0),.clk(gclk));
	jdff dff_B_0At1ML9x5_0(.din(w_dff_B_SfYFSYlY8_0),.dout(w_dff_B_0At1ML9x5_0),.clk(gclk));
	jdff dff_B_4vR1Fg8b0_0(.din(w_dff_B_0At1ML9x5_0),.dout(w_dff_B_4vR1Fg8b0_0),.clk(gclk));
	jdff dff_B_y4cCk3QS7_0(.din(w_dff_B_4vR1Fg8b0_0),.dout(w_dff_B_y4cCk3QS7_0),.clk(gclk));
	jdff dff_B_kjQazQ2J0_0(.din(w_dff_B_y4cCk3QS7_0),.dout(w_dff_B_kjQazQ2J0_0),.clk(gclk));
	jdff dff_B_tFfMyx684_0(.din(w_dff_B_kjQazQ2J0_0),.dout(w_dff_B_tFfMyx684_0),.clk(gclk));
	jdff dff_B_tkkHea3i0_0(.din(w_dff_B_tFfMyx684_0),.dout(w_dff_B_tkkHea3i0_0),.clk(gclk));
	jdff dff_B_vWkwsoob5_1(.din(n840),.dout(w_dff_B_vWkwsoob5_1),.clk(gclk));
	jdff dff_B_kHKmM3Us2_1(.din(w_dff_B_vWkwsoob5_1),.dout(w_dff_B_kHKmM3Us2_1),.clk(gclk));
	jdff dff_B_QuhYpKCW9_1(.din(w_dff_B_kHKmM3Us2_1),.dout(w_dff_B_QuhYpKCW9_1),.clk(gclk));
	jdff dff_B_LALH7kbx2_1(.din(w_dff_B_QuhYpKCW9_1),.dout(w_dff_B_LALH7kbx2_1),.clk(gclk));
	jdff dff_B_M6b94v5q0_1(.din(w_dff_B_LALH7kbx2_1),.dout(w_dff_B_M6b94v5q0_1),.clk(gclk));
	jdff dff_B_dIFwdDTK5_1(.din(w_dff_B_M6b94v5q0_1),.dout(w_dff_B_dIFwdDTK5_1),.clk(gclk));
	jdff dff_B_cyp5PYob1_1(.din(w_dff_B_dIFwdDTK5_1),.dout(w_dff_B_cyp5PYob1_1),.clk(gclk));
	jdff dff_B_AC1l9Bnu7_1(.din(w_dff_B_cyp5PYob1_1),.dout(w_dff_B_AC1l9Bnu7_1),.clk(gclk));
	jdff dff_B_UNxvzmta7_1(.din(w_dff_B_AC1l9Bnu7_1),.dout(w_dff_B_UNxvzmta7_1),.clk(gclk));
	jdff dff_B_dwMsz9xw0_1(.din(w_dff_B_UNxvzmta7_1),.dout(w_dff_B_dwMsz9xw0_1),.clk(gclk));
	jdff dff_B_pX2UXhnk6_1(.din(w_dff_B_dwMsz9xw0_1),.dout(w_dff_B_pX2UXhnk6_1),.clk(gclk));
	jdff dff_B_pzGV0cx13_1(.din(w_dff_B_pX2UXhnk6_1),.dout(w_dff_B_pzGV0cx13_1),.clk(gclk));
	jdff dff_B_Tr32mQqt8_1(.din(w_dff_B_pzGV0cx13_1),.dout(w_dff_B_Tr32mQqt8_1),.clk(gclk));
	jdff dff_B_Qzrdw8Sa6_1(.din(w_dff_B_Tr32mQqt8_1),.dout(w_dff_B_Qzrdw8Sa6_1),.clk(gclk));
	jdff dff_B_PdTKADZr3_1(.din(w_dff_B_Qzrdw8Sa6_1),.dout(w_dff_B_PdTKADZr3_1),.clk(gclk));
	jdff dff_B_gM71vmhI7_1(.din(w_dff_B_PdTKADZr3_1),.dout(w_dff_B_gM71vmhI7_1),.clk(gclk));
	jdff dff_B_Rhwm3rHQ4_1(.din(w_dff_B_gM71vmhI7_1),.dout(w_dff_B_Rhwm3rHQ4_1),.clk(gclk));
	jdff dff_B_OWsBmfZN5_1(.din(w_dff_B_Rhwm3rHQ4_1),.dout(w_dff_B_OWsBmfZN5_1),.clk(gclk));
	jdff dff_B_iD3D3xJB5_1(.din(w_dff_B_OWsBmfZN5_1),.dout(w_dff_B_iD3D3xJB5_1),.clk(gclk));
	jdff dff_B_ThbPfWDJ1_1(.din(w_dff_B_iD3D3xJB5_1),.dout(w_dff_B_ThbPfWDJ1_1),.clk(gclk));
	jdff dff_B_UKXhGR6F1_1(.din(w_dff_B_ThbPfWDJ1_1),.dout(w_dff_B_UKXhGR6F1_1),.clk(gclk));
	jdff dff_B_5kQ52v5b1_1(.din(w_dff_B_UKXhGR6F1_1),.dout(w_dff_B_5kQ52v5b1_1),.clk(gclk));
	jdff dff_B_PenMa5rR3_1(.din(w_dff_B_5kQ52v5b1_1),.dout(w_dff_B_PenMa5rR3_1),.clk(gclk));
	jdff dff_B_t7zXDa3p1_1(.din(w_dff_B_PenMa5rR3_1),.dout(w_dff_B_t7zXDa3p1_1),.clk(gclk));
	jdff dff_B_u732Smtf0_1(.din(w_dff_B_t7zXDa3p1_1),.dout(w_dff_B_u732Smtf0_1),.clk(gclk));
	jdff dff_B_td6gkA3P9_1(.din(w_dff_B_u732Smtf0_1),.dout(w_dff_B_td6gkA3P9_1),.clk(gclk));
	jdff dff_B_URAlXzOj5_1(.din(w_dff_B_td6gkA3P9_1),.dout(w_dff_B_URAlXzOj5_1),.clk(gclk));
	jdff dff_B_wLs0cD850_1(.din(w_dff_B_URAlXzOj5_1),.dout(w_dff_B_wLs0cD850_1),.clk(gclk));
	jdff dff_B_EcA06yZa4_1(.din(w_dff_B_wLs0cD850_1),.dout(w_dff_B_EcA06yZa4_1),.clk(gclk));
	jdff dff_B_Dsiq8tRm8_1(.din(w_dff_B_EcA06yZa4_1),.dout(w_dff_B_Dsiq8tRm8_1),.clk(gclk));
	jdff dff_B_5RzThljG4_1(.din(w_dff_B_Dsiq8tRm8_1),.dout(w_dff_B_5RzThljG4_1),.clk(gclk));
	jdff dff_B_iD28wjrw3_1(.din(w_dff_B_5RzThljG4_1),.dout(w_dff_B_iD28wjrw3_1),.clk(gclk));
	jdff dff_B_nt5ccctD4_1(.din(w_dff_B_iD28wjrw3_1),.dout(w_dff_B_nt5ccctD4_1),.clk(gclk));
	jdff dff_B_bWOW1rZQ6_1(.din(w_dff_B_nt5ccctD4_1),.dout(w_dff_B_bWOW1rZQ6_1),.clk(gclk));
	jdff dff_B_9Vz53FNo6_1(.din(w_dff_B_bWOW1rZQ6_1),.dout(w_dff_B_9Vz53FNo6_1),.clk(gclk));
	jdff dff_B_TFANf9cN6_1(.din(w_dff_B_9Vz53FNo6_1),.dout(w_dff_B_TFANf9cN6_1),.clk(gclk));
	jdff dff_B_74ruwPTI7_1(.din(w_dff_B_TFANf9cN6_1),.dout(w_dff_B_74ruwPTI7_1),.clk(gclk));
	jdff dff_B_8UFPFhdU6_1(.din(w_dff_B_74ruwPTI7_1),.dout(w_dff_B_8UFPFhdU6_1),.clk(gclk));
	jdff dff_B_qVFtB9gW4_1(.din(w_dff_B_8UFPFhdU6_1),.dout(w_dff_B_qVFtB9gW4_1),.clk(gclk));
	jdff dff_B_E8ov80fE0_1(.din(w_dff_B_qVFtB9gW4_1),.dout(w_dff_B_E8ov80fE0_1),.clk(gclk));
	jdff dff_B_saiEfAmf8_1(.din(w_dff_B_E8ov80fE0_1),.dout(w_dff_B_saiEfAmf8_1),.clk(gclk));
	jdff dff_B_yVTKt6Cz2_1(.din(w_dff_B_saiEfAmf8_1),.dout(w_dff_B_yVTKt6Cz2_1),.clk(gclk));
	jdff dff_B_YLArECpI4_1(.din(w_dff_B_yVTKt6Cz2_1),.dout(w_dff_B_YLArECpI4_1),.clk(gclk));
	jdff dff_B_dmi9TOxo7_1(.din(w_dff_B_YLArECpI4_1),.dout(w_dff_B_dmi9TOxo7_1),.clk(gclk));
	jdff dff_B_W2j8eTxx6_1(.din(w_dff_B_dmi9TOxo7_1),.dout(w_dff_B_W2j8eTxx6_1),.clk(gclk));
	jdff dff_B_XB4D5V0k0_1(.din(w_dff_B_W2j8eTxx6_1),.dout(w_dff_B_XB4D5V0k0_1),.clk(gclk));
	jdff dff_B_1ir5ZE9B3_1(.din(w_dff_B_XB4D5V0k0_1),.dout(w_dff_B_1ir5ZE9B3_1),.clk(gclk));
	jdff dff_B_8fEKguUf5_1(.din(w_dff_B_1ir5ZE9B3_1),.dout(w_dff_B_8fEKguUf5_1),.clk(gclk));
	jdff dff_B_Q2SbXHbd3_1(.din(w_dff_B_8fEKguUf5_1),.dout(w_dff_B_Q2SbXHbd3_1),.clk(gclk));
	jdff dff_B_jMQM2M6y5_1(.din(w_dff_B_Q2SbXHbd3_1),.dout(w_dff_B_jMQM2M6y5_1),.clk(gclk));
	jdff dff_B_nzRnGZpe3_1(.din(w_dff_B_jMQM2M6y5_1),.dout(w_dff_B_nzRnGZpe3_1),.clk(gclk));
	jdff dff_B_ReEGW0oi9_1(.din(w_dff_B_nzRnGZpe3_1),.dout(w_dff_B_ReEGW0oi9_1),.clk(gclk));
	jdff dff_B_K5gh1g9W8_1(.din(w_dff_B_ReEGW0oi9_1),.dout(w_dff_B_K5gh1g9W8_1),.clk(gclk));
	jdff dff_B_vgk24bdc8_1(.din(w_dff_B_K5gh1g9W8_1),.dout(w_dff_B_vgk24bdc8_1),.clk(gclk));
	jdff dff_B_i4rzaCrW7_1(.din(w_dff_B_vgk24bdc8_1),.dout(w_dff_B_i4rzaCrW7_1),.clk(gclk));
	jdff dff_B_NdjYAE8v1_1(.din(w_dff_B_i4rzaCrW7_1),.dout(w_dff_B_NdjYAE8v1_1),.clk(gclk));
	jdff dff_B_hqtRGZx85_1(.din(w_dff_B_NdjYAE8v1_1),.dout(w_dff_B_hqtRGZx85_1),.clk(gclk));
	jdff dff_B_jpfjsvFt6_1(.din(w_dff_B_hqtRGZx85_1),.dout(w_dff_B_jpfjsvFt6_1),.clk(gclk));
	jdff dff_B_aypb6kBz2_1(.din(w_dff_B_jpfjsvFt6_1),.dout(w_dff_B_aypb6kBz2_1),.clk(gclk));
	jdff dff_B_PkxuWRtq7_1(.din(w_dff_B_aypb6kBz2_1),.dout(w_dff_B_PkxuWRtq7_1),.clk(gclk));
	jdff dff_B_c8JM0jut5_1(.din(w_dff_B_PkxuWRtq7_1),.dout(w_dff_B_c8JM0jut5_1),.clk(gclk));
	jdff dff_B_PBpMSWtP2_1(.din(w_dff_B_c8JM0jut5_1),.dout(w_dff_B_PBpMSWtP2_1),.clk(gclk));
	jdff dff_B_AmIYtOuT1_1(.din(w_dff_B_PBpMSWtP2_1),.dout(w_dff_B_AmIYtOuT1_1),.clk(gclk));
	jdff dff_B_dI38pliI1_1(.din(w_dff_B_AmIYtOuT1_1),.dout(w_dff_B_dI38pliI1_1),.clk(gclk));
	jdff dff_B_EayRjbrE3_1(.din(w_dff_B_dI38pliI1_1),.dout(w_dff_B_EayRjbrE3_1),.clk(gclk));
	jdff dff_B_RWW4oKsi1_1(.din(w_dff_B_EayRjbrE3_1),.dout(w_dff_B_RWW4oKsi1_1),.clk(gclk));
	jdff dff_B_cDBqrpOP5_1(.din(w_dff_B_RWW4oKsi1_1),.dout(w_dff_B_cDBqrpOP5_1),.clk(gclk));
	jdff dff_B_D8ukmdFy4_1(.din(w_dff_B_cDBqrpOP5_1),.dout(w_dff_B_D8ukmdFy4_1),.clk(gclk));
	jdff dff_B_W8Vmw1lW3_1(.din(w_dff_B_D8ukmdFy4_1),.dout(w_dff_B_W8Vmw1lW3_1),.clk(gclk));
	jdff dff_B_JlLdtDBr9_1(.din(w_dff_B_W8Vmw1lW3_1),.dout(w_dff_B_JlLdtDBr9_1),.clk(gclk));
	jdff dff_B_GyjGYEKW3_1(.din(w_dff_B_JlLdtDBr9_1),.dout(w_dff_B_GyjGYEKW3_1),.clk(gclk));
	jdff dff_B_SSsgMMn53_1(.din(w_dff_B_GyjGYEKW3_1),.dout(w_dff_B_SSsgMMn53_1),.clk(gclk));
	jdff dff_B_1BfijTHY6_1(.din(w_dff_B_SSsgMMn53_1),.dout(w_dff_B_1BfijTHY6_1),.clk(gclk));
	jdff dff_B_B2QvJI0J3_1(.din(w_dff_B_1BfijTHY6_1),.dout(w_dff_B_B2QvJI0J3_1),.clk(gclk));
	jdff dff_B_7CxKjaeA3_1(.din(w_dff_B_B2QvJI0J3_1),.dout(w_dff_B_7CxKjaeA3_1),.clk(gclk));
	jdff dff_B_NwsfVLEn3_1(.din(w_dff_B_7CxKjaeA3_1),.dout(w_dff_B_NwsfVLEn3_1),.clk(gclk));
	jdff dff_B_xhrH6Nm59_0(.din(n841),.dout(w_dff_B_xhrH6Nm59_0),.clk(gclk));
	jdff dff_B_IIVCRSfT9_0(.din(w_dff_B_xhrH6Nm59_0),.dout(w_dff_B_IIVCRSfT9_0),.clk(gclk));
	jdff dff_B_Vz75Hc9N1_0(.din(w_dff_B_IIVCRSfT9_0),.dout(w_dff_B_Vz75Hc9N1_0),.clk(gclk));
	jdff dff_B_ryUncve94_0(.din(w_dff_B_Vz75Hc9N1_0),.dout(w_dff_B_ryUncve94_0),.clk(gclk));
	jdff dff_B_fzwsv5Ng7_0(.din(w_dff_B_ryUncve94_0),.dout(w_dff_B_fzwsv5Ng7_0),.clk(gclk));
	jdff dff_B_02ur9dbA6_0(.din(w_dff_B_fzwsv5Ng7_0),.dout(w_dff_B_02ur9dbA6_0),.clk(gclk));
	jdff dff_B_Ukbytt5a0_0(.din(w_dff_B_02ur9dbA6_0),.dout(w_dff_B_Ukbytt5a0_0),.clk(gclk));
	jdff dff_B_upfwbd9v5_0(.din(w_dff_B_Ukbytt5a0_0),.dout(w_dff_B_upfwbd9v5_0),.clk(gclk));
	jdff dff_B_jVU0m9z81_0(.din(w_dff_B_upfwbd9v5_0),.dout(w_dff_B_jVU0m9z81_0),.clk(gclk));
	jdff dff_B_m6jinLyX8_0(.din(w_dff_B_jVU0m9z81_0),.dout(w_dff_B_m6jinLyX8_0),.clk(gclk));
	jdff dff_B_q3f2w4hW9_0(.din(w_dff_B_m6jinLyX8_0),.dout(w_dff_B_q3f2w4hW9_0),.clk(gclk));
	jdff dff_B_EelgDfDz9_0(.din(w_dff_B_q3f2w4hW9_0),.dout(w_dff_B_EelgDfDz9_0),.clk(gclk));
	jdff dff_B_YWDRUUir3_0(.din(w_dff_B_EelgDfDz9_0),.dout(w_dff_B_YWDRUUir3_0),.clk(gclk));
	jdff dff_B_2jGsQFbT9_0(.din(w_dff_B_YWDRUUir3_0),.dout(w_dff_B_2jGsQFbT9_0),.clk(gclk));
	jdff dff_B_FFxz1r686_0(.din(w_dff_B_2jGsQFbT9_0),.dout(w_dff_B_FFxz1r686_0),.clk(gclk));
	jdff dff_B_LjfOJKfn9_0(.din(w_dff_B_FFxz1r686_0),.dout(w_dff_B_LjfOJKfn9_0),.clk(gclk));
	jdff dff_B_bhF2X3nJ8_0(.din(w_dff_B_LjfOJKfn9_0),.dout(w_dff_B_bhF2X3nJ8_0),.clk(gclk));
	jdff dff_B_q78C42SI4_0(.din(w_dff_B_bhF2X3nJ8_0),.dout(w_dff_B_q78C42SI4_0),.clk(gclk));
	jdff dff_B_ZTfgykT46_0(.din(w_dff_B_q78C42SI4_0),.dout(w_dff_B_ZTfgykT46_0),.clk(gclk));
	jdff dff_B_MFr8crzT2_0(.din(w_dff_B_ZTfgykT46_0),.dout(w_dff_B_MFr8crzT2_0),.clk(gclk));
	jdff dff_B_C5Pddw0X6_0(.din(w_dff_B_MFr8crzT2_0),.dout(w_dff_B_C5Pddw0X6_0),.clk(gclk));
	jdff dff_B_Qw0Yx3lN7_0(.din(w_dff_B_C5Pddw0X6_0),.dout(w_dff_B_Qw0Yx3lN7_0),.clk(gclk));
	jdff dff_B_yZ4UumJW5_0(.din(w_dff_B_Qw0Yx3lN7_0),.dout(w_dff_B_yZ4UumJW5_0),.clk(gclk));
	jdff dff_B_t9XNvqfh7_0(.din(w_dff_B_yZ4UumJW5_0),.dout(w_dff_B_t9XNvqfh7_0),.clk(gclk));
	jdff dff_B_Naen5Ig93_0(.din(w_dff_B_t9XNvqfh7_0),.dout(w_dff_B_Naen5Ig93_0),.clk(gclk));
	jdff dff_B_iJ5WC9Jq0_0(.din(w_dff_B_Naen5Ig93_0),.dout(w_dff_B_iJ5WC9Jq0_0),.clk(gclk));
	jdff dff_B_SLGAKHsB9_0(.din(w_dff_B_iJ5WC9Jq0_0),.dout(w_dff_B_SLGAKHsB9_0),.clk(gclk));
	jdff dff_B_6Ays6BV72_0(.din(w_dff_B_SLGAKHsB9_0),.dout(w_dff_B_6Ays6BV72_0),.clk(gclk));
	jdff dff_B_h98fre8B9_0(.din(w_dff_B_6Ays6BV72_0),.dout(w_dff_B_h98fre8B9_0),.clk(gclk));
	jdff dff_B_M0PymkID7_0(.din(w_dff_B_h98fre8B9_0),.dout(w_dff_B_M0PymkID7_0),.clk(gclk));
	jdff dff_B_8VV1FZOi7_0(.din(w_dff_B_M0PymkID7_0),.dout(w_dff_B_8VV1FZOi7_0),.clk(gclk));
	jdff dff_B_npTNlMOa8_0(.din(w_dff_B_8VV1FZOi7_0),.dout(w_dff_B_npTNlMOa8_0),.clk(gclk));
	jdff dff_B_cUMyGulG0_0(.din(w_dff_B_npTNlMOa8_0),.dout(w_dff_B_cUMyGulG0_0),.clk(gclk));
	jdff dff_B_o8G2JyCb5_0(.din(w_dff_B_cUMyGulG0_0),.dout(w_dff_B_o8G2JyCb5_0),.clk(gclk));
	jdff dff_B_myRu39ur8_0(.din(w_dff_B_o8G2JyCb5_0),.dout(w_dff_B_myRu39ur8_0),.clk(gclk));
	jdff dff_B_xZA5tJ8K2_0(.din(w_dff_B_myRu39ur8_0),.dout(w_dff_B_xZA5tJ8K2_0),.clk(gclk));
	jdff dff_B_61J9Poug7_0(.din(w_dff_B_xZA5tJ8K2_0),.dout(w_dff_B_61J9Poug7_0),.clk(gclk));
	jdff dff_B_2baMkR5X5_0(.din(w_dff_B_61J9Poug7_0),.dout(w_dff_B_2baMkR5X5_0),.clk(gclk));
	jdff dff_B_SshvMVj89_0(.din(w_dff_B_2baMkR5X5_0),.dout(w_dff_B_SshvMVj89_0),.clk(gclk));
	jdff dff_B_X2z7ayJJ8_0(.din(w_dff_B_SshvMVj89_0),.dout(w_dff_B_X2z7ayJJ8_0),.clk(gclk));
	jdff dff_B_Yg0dPY2j1_0(.din(w_dff_B_X2z7ayJJ8_0),.dout(w_dff_B_Yg0dPY2j1_0),.clk(gclk));
	jdff dff_B_2G52tnv12_0(.din(w_dff_B_Yg0dPY2j1_0),.dout(w_dff_B_2G52tnv12_0),.clk(gclk));
	jdff dff_B_0hAfMPkm1_0(.din(w_dff_B_2G52tnv12_0),.dout(w_dff_B_0hAfMPkm1_0),.clk(gclk));
	jdff dff_B_rD9euaHI7_0(.din(w_dff_B_0hAfMPkm1_0),.dout(w_dff_B_rD9euaHI7_0),.clk(gclk));
	jdff dff_B_hEsduBhp0_0(.din(w_dff_B_rD9euaHI7_0),.dout(w_dff_B_hEsduBhp0_0),.clk(gclk));
	jdff dff_B_V7sCtpSY6_0(.din(w_dff_B_hEsduBhp0_0),.dout(w_dff_B_V7sCtpSY6_0),.clk(gclk));
	jdff dff_B_qOv9yfU77_0(.din(w_dff_B_V7sCtpSY6_0),.dout(w_dff_B_qOv9yfU77_0),.clk(gclk));
	jdff dff_B_PoNosoNN3_0(.din(w_dff_B_qOv9yfU77_0),.dout(w_dff_B_PoNosoNN3_0),.clk(gclk));
	jdff dff_B_lIBmC1Rw9_0(.din(w_dff_B_PoNosoNN3_0),.dout(w_dff_B_lIBmC1Rw9_0),.clk(gclk));
	jdff dff_B_t16Darf14_0(.din(w_dff_B_lIBmC1Rw9_0),.dout(w_dff_B_t16Darf14_0),.clk(gclk));
	jdff dff_B_0han21e32_0(.din(w_dff_B_t16Darf14_0),.dout(w_dff_B_0han21e32_0),.clk(gclk));
	jdff dff_B_q0Txbzls2_0(.din(w_dff_B_0han21e32_0),.dout(w_dff_B_q0Txbzls2_0),.clk(gclk));
	jdff dff_B_bd2CmCoH1_0(.din(w_dff_B_q0Txbzls2_0),.dout(w_dff_B_bd2CmCoH1_0),.clk(gclk));
	jdff dff_B_DFh0NfmB0_0(.din(w_dff_B_bd2CmCoH1_0),.dout(w_dff_B_DFh0NfmB0_0),.clk(gclk));
	jdff dff_B_0ACsdpkW0_0(.din(w_dff_B_DFh0NfmB0_0),.dout(w_dff_B_0ACsdpkW0_0),.clk(gclk));
	jdff dff_B_OSkzEPVq1_0(.din(w_dff_B_0ACsdpkW0_0),.dout(w_dff_B_OSkzEPVq1_0),.clk(gclk));
	jdff dff_B_IGcDcHAI4_0(.din(w_dff_B_OSkzEPVq1_0),.dout(w_dff_B_IGcDcHAI4_0),.clk(gclk));
	jdff dff_B_IhMaCvDh6_0(.din(w_dff_B_IGcDcHAI4_0),.dout(w_dff_B_IhMaCvDh6_0),.clk(gclk));
	jdff dff_B_dySYdNLk3_0(.din(w_dff_B_IhMaCvDh6_0),.dout(w_dff_B_dySYdNLk3_0),.clk(gclk));
	jdff dff_B_q5toYGPF8_0(.din(w_dff_B_dySYdNLk3_0),.dout(w_dff_B_q5toYGPF8_0),.clk(gclk));
	jdff dff_B_gaqWYEvY9_0(.din(w_dff_B_q5toYGPF8_0),.dout(w_dff_B_gaqWYEvY9_0),.clk(gclk));
	jdff dff_B_WE0qIHoN2_0(.din(w_dff_B_gaqWYEvY9_0),.dout(w_dff_B_WE0qIHoN2_0),.clk(gclk));
	jdff dff_B_X4w4jAka2_0(.din(w_dff_B_WE0qIHoN2_0),.dout(w_dff_B_X4w4jAka2_0),.clk(gclk));
	jdff dff_B_0r5nbhGq5_0(.din(w_dff_B_X4w4jAka2_0),.dout(w_dff_B_0r5nbhGq5_0),.clk(gclk));
	jdff dff_B_en0bcXGN9_0(.din(w_dff_B_0r5nbhGq5_0),.dout(w_dff_B_en0bcXGN9_0),.clk(gclk));
	jdff dff_B_F4xZ3c6h7_0(.din(w_dff_B_en0bcXGN9_0),.dout(w_dff_B_F4xZ3c6h7_0),.clk(gclk));
	jdff dff_B_ViVPGS8l2_0(.din(w_dff_B_F4xZ3c6h7_0),.dout(w_dff_B_ViVPGS8l2_0),.clk(gclk));
	jdff dff_B_l0Yf07rA0_0(.din(w_dff_B_ViVPGS8l2_0),.dout(w_dff_B_l0Yf07rA0_0),.clk(gclk));
	jdff dff_B_B5LtcFVG6_0(.din(w_dff_B_l0Yf07rA0_0),.dout(w_dff_B_B5LtcFVG6_0),.clk(gclk));
	jdff dff_B_vRbftr4M2_0(.din(w_dff_B_B5LtcFVG6_0),.dout(w_dff_B_vRbftr4M2_0),.clk(gclk));
	jdff dff_B_pC7rqyHu3_0(.din(w_dff_B_vRbftr4M2_0),.dout(w_dff_B_pC7rqyHu3_0),.clk(gclk));
	jdff dff_B_hlndAAMl5_0(.din(w_dff_B_pC7rqyHu3_0),.dout(w_dff_B_hlndAAMl5_0),.clk(gclk));
	jdff dff_B_qozOIvyD4_0(.din(w_dff_B_hlndAAMl5_0),.dout(w_dff_B_qozOIvyD4_0),.clk(gclk));
	jdff dff_B_XAE10I893_0(.din(w_dff_B_qozOIvyD4_0),.dout(w_dff_B_XAE10I893_0),.clk(gclk));
	jdff dff_B_SeDS6H6O2_0(.din(w_dff_B_XAE10I893_0),.dout(w_dff_B_SeDS6H6O2_0),.clk(gclk));
	jdff dff_B_ogHkkQPV9_0(.din(w_dff_B_SeDS6H6O2_0),.dout(w_dff_B_ogHkkQPV9_0),.clk(gclk));
	jdff dff_B_fHBzS1Qj2_1(.din(n834),.dout(w_dff_B_fHBzS1Qj2_1),.clk(gclk));
	jdff dff_B_GRopQDNe2_1(.din(w_dff_B_fHBzS1Qj2_1),.dout(w_dff_B_GRopQDNe2_1),.clk(gclk));
	jdff dff_B_mHqdaL8S5_1(.din(w_dff_B_GRopQDNe2_1),.dout(w_dff_B_mHqdaL8S5_1),.clk(gclk));
	jdff dff_B_NkKEE4hf8_1(.din(w_dff_B_mHqdaL8S5_1),.dout(w_dff_B_NkKEE4hf8_1),.clk(gclk));
	jdff dff_B_5HJd2Ywu1_1(.din(w_dff_B_NkKEE4hf8_1),.dout(w_dff_B_5HJd2Ywu1_1),.clk(gclk));
	jdff dff_B_0V7iFQOI8_1(.din(w_dff_B_5HJd2Ywu1_1),.dout(w_dff_B_0V7iFQOI8_1),.clk(gclk));
	jdff dff_B_yzYSvzCT6_1(.din(w_dff_B_0V7iFQOI8_1),.dout(w_dff_B_yzYSvzCT6_1),.clk(gclk));
	jdff dff_B_J5V2NcVn0_1(.din(w_dff_B_yzYSvzCT6_1),.dout(w_dff_B_J5V2NcVn0_1),.clk(gclk));
	jdff dff_B_iG1sVmlX9_1(.din(w_dff_B_J5V2NcVn0_1),.dout(w_dff_B_iG1sVmlX9_1),.clk(gclk));
	jdff dff_B_aaq4mC4U7_1(.din(w_dff_B_iG1sVmlX9_1),.dout(w_dff_B_aaq4mC4U7_1),.clk(gclk));
	jdff dff_B_Pz9yoNB81_1(.din(w_dff_B_aaq4mC4U7_1),.dout(w_dff_B_Pz9yoNB81_1),.clk(gclk));
	jdff dff_B_5htoz7wO1_1(.din(w_dff_B_Pz9yoNB81_1),.dout(w_dff_B_5htoz7wO1_1),.clk(gclk));
	jdff dff_B_IMRkCq3l5_1(.din(w_dff_B_5htoz7wO1_1),.dout(w_dff_B_IMRkCq3l5_1),.clk(gclk));
	jdff dff_B_jfHSZsx56_1(.din(w_dff_B_IMRkCq3l5_1),.dout(w_dff_B_jfHSZsx56_1),.clk(gclk));
	jdff dff_B_SqclJWp48_1(.din(w_dff_B_jfHSZsx56_1),.dout(w_dff_B_SqclJWp48_1),.clk(gclk));
	jdff dff_B_keN5G0ag7_1(.din(w_dff_B_SqclJWp48_1),.dout(w_dff_B_keN5G0ag7_1),.clk(gclk));
	jdff dff_B_pEHqStHt6_1(.din(w_dff_B_keN5G0ag7_1),.dout(w_dff_B_pEHqStHt6_1),.clk(gclk));
	jdff dff_B_Fpis1flx9_1(.din(w_dff_B_pEHqStHt6_1),.dout(w_dff_B_Fpis1flx9_1),.clk(gclk));
	jdff dff_B_ENUDrgFV6_1(.din(w_dff_B_Fpis1flx9_1),.dout(w_dff_B_ENUDrgFV6_1),.clk(gclk));
	jdff dff_B_QiucTPP74_1(.din(w_dff_B_ENUDrgFV6_1),.dout(w_dff_B_QiucTPP74_1),.clk(gclk));
	jdff dff_B_0bzNuzCC6_1(.din(w_dff_B_QiucTPP74_1),.dout(w_dff_B_0bzNuzCC6_1),.clk(gclk));
	jdff dff_B_WKWUERgi6_1(.din(w_dff_B_0bzNuzCC6_1),.dout(w_dff_B_WKWUERgi6_1),.clk(gclk));
	jdff dff_B_CE07WeNE8_1(.din(w_dff_B_WKWUERgi6_1),.dout(w_dff_B_CE07WeNE8_1),.clk(gclk));
	jdff dff_B_6Gxr33yF0_1(.din(w_dff_B_CE07WeNE8_1),.dout(w_dff_B_6Gxr33yF0_1),.clk(gclk));
	jdff dff_B_smrgTVRZ0_1(.din(w_dff_B_6Gxr33yF0_1),.dout(w_dff_B_smrgTVRZ0_1),.clk(gclk));
	jdff dff_B_HKmPsPlD7_1(.din(w_dff_B_smrgTVRZ0_1),.dout(w_dff_B_HKmPsPlD7_1),.clk(gclk));
	jdff dff_B_w4gle9Fi8_1(.din(w_dff_B_HKmPsPlD7_1),.dout(w_dff_B_w4gle9Fi8_1),.clk(gclk));
	jdff dff_B_0l6Fwr7h9_1(.din(w_dff_B_w4gle9Fi8_1),.dout(w_dff_B_0l6Fwr7h9_1),.clk(gclk));
	jdff dff_B_yX8FJu2R6_1(.din(w_dff_B_0l6Fwr7h9_1),.dout(w_dff_B_yX8FJu2R6_1),.clk(gclk));
	jdff dff_B_rfFExPzG2_1(.din(w_dff_B_yX8FJu2R6_1),.dout(w_dff_B_rfFExPzG2_1),.clk(gclk));
	jdff dff_B_mVKGQXKT0_1(.din(w_dff_B_rfFExPzG2_1),.dout(w_dff_B_mVKGQXKT0_1),.clk(gclk));
	jdff dff_B_wRfypqQU9_1(.din(w_dff_B_mVKGQXKT0_1),.dout(w_dff_B_wRfypqQU9_1),.clk(gclk));
	jdff dff_B_FFaY4lUK9_1(.din(w_dff_B_wRfypqQU9_1),.dout(w_dff_B_FFaY4lUK9_1),.clk(gclk));
	jdff dff_B_iTYtuHjh7_1(.din(w_dff_B_FFaY4lUK9_1),.dout(w_dff_B_iTYtuHjh7_1),.clk(gclk));
	jdff dff_B_A6BE0GtO2_1(.din(w_dff_B_iTYtuHjh7_1),.dout(w_dff_B_A6BE0GtO2_1),.clk(gclk));
	jdff dff_B_cJyNYkpL9_1(.din(w_dff_B_A6BE0GtO2_1),.dout(w_dff_B_cJyNYkpL9_1),.clk(gclk));
	jdff dff_B_vTdJpKuB7_1(.din(w_dff_B_cJyNYkpL9_1),.dout(w_dff_B_vTdJpKuB7_1),.clk(gclk));
	jdff dff_B_SBVp6tmq7_1(.din(w_dff_B_vTdJpKuB7_1),.dout(w_dff_B_SBVp6tmq7_1),.clk(gclk));
	jdff dff_B_XIgoaezm7_1(.din(w_dff_B_SBVp6tmq7_1),.dout(w_dff_B_XIgoaezm7_1),.clk(gclk));
	jdff dff_B_fgqZTn0Y2_1(.din(w_dff_B_XIgoaezm7_1),.dout(w_dff_B_fgqZTn0Y2_1),.clk(gclk));
	jdff dff_B_dBGCToTY4_1(.din(w_dff_B_fgqZTn0Y2_1),.dout(w_dff_B_dBGCToTY4_1),.clk(gclk));
	jdff dff_B_f1na4EFN5_1(.din(w_dff_B_dBGCToTY4_1),.dout(w_dff_B_f1na4EFN5_1),.clk(gclk));
	jdff dff_B_5RN1rz7j2_1(.din(w_dff_B_f1na4EFN5_1),.dout(w_dff_B_5RN1rz7j2_1),.clk(gclk));
	jdff dff_B_KL748LSw3_1(.din(w_dff_B_5RN1rz7j2_1),.dout(w_dff_B_KL748LSw3_1),.clk(gclk));
	jdff dff_B_LVEgZ2y84_1(.din(w_dff_B_KL748LSw3_1),.dout(w_dff_B_LVEgZ2y84_1),.clk(gclk));
	jdff dff_B_Pz0C8YGX5_1(.din(w_dff_B_LVEgZ2y84_1),.dout(w_dff_B_Pz0C8YGX5_1),.clk(gclk));
	jdff dff_B_fIIhbOo01_1(.din(w_dff_B_Pz0C8YGX5_1),.dout(w_dff_B_fIIhbOo01_1),.clk(gclk));
	jdff dff_B_AgVwI4mG7_1(.din(w_dff_B_fIIhbOo01_1),.dout(w_dff_B_AgVwI4mG7_1),.clk(gclk));
	jdff dff_B_gb5X35pF6_1(.din(w_dff_B_AgVwI4mG7_1),.dout(w_dff_B_gb5X35pF6_1),.clk(gclk));
	jdff dff_B_lTF4DvuM2_1(.din(w_dff_B_gb5X35pF6_1),.dout(w_dff_B_lTF4DvuM2_1),.clk(gclk));
	jdff dff_B_fpQBtV6F4_1(.din(w_dff_B_lTF4DvuM2_1),.dout(w_dff_B_fpQBtV6F4_1),.clk(gclk));
	jdff dff_B_cXx7hrRE8_1(.din(w_dff_B_fpQBtV6F4_1),.dout(w_dff_B_cXx7hrRE8_1),.clk(gclk));
	jdff dff_B_yU8IOQd13_1(.din(w_dff_B_cXx7hrRE8_1),.dout(w_dff_B_yU8IOQd13_1),.clk(gclk));
	jdff dff_B_EBuIYaZv1_1(.din(w_dff_B_yU8IOQd13_1),.dout(w_dff_B_EBuIYaZv1_1),.clk(gclk));
	jdff dff_B_NhG75iV78_1(.din(w_dff_B_EBuIYaZv1_1),.dout(w_dff_B_NhG75iV78_1),.clk(gclk));
	jdff dff_B_P1xugy5g5_1(.din(w_dff_B_NhG75iV78_1),.dout(w_dff_B_P1xugy5g5_1),.clk(gclk));
	jdff dff_B_qJKTQRMG5_1(.din(w_dff_B_P1xugy5g5_1),.dout(w_dff_B_qJKTQRMG5_1),.clk(gclk));
	jdff dff_B_HSAtnPCm9_1(.din(w_dff_B_qJKTQRMG5_1),.dout(w_dff_B_HSAtnPCm9_1),.clk(gclk));
	jdff dff_B_2OI6n3n12_1(.din(w_dff_B_HSAtnPCm9_1),.dout(w_dff_B_2OI6n3n12_1),.clk(gclk));
	jdff dff_B_HNtekZpL1_1(.din(w_dff_B_2OI6n3n12_1),.dout(w_dff_B_HNtekZpL1_1),.clk(gclk));
	jdff dff_B_reYtGFKb0_1(.din(w_dff_B_HNtekZpL1_1),.dout(w_dff_B_reYtGFKb0_1),.clk(gclk));
	jdff dff_B_RlHvAOD07_1(.din(w_dff_B_reYtGFKb0_1),.dout(w_dff_B_RlHvAOD07_1),.clk(gclk));
	jdff dff_B_sPPHuCiZ6_1(.din(w_dff_B_RlHvAOD07_1),.dout(w_dff_B_sPPHuCiZ6_1),.clk(gclk));
	jdff dff_B_FazavZOt9_1(.din(w_dff_B_sPPHuCiZ6_1),.dout(w_dff_B_FazavZOt9_1),.clk(gclk));
	jdff dff_B_JtloA87w9_1(.din(w_dff_B_FazavZOt9_1),.dout(w_dff_B_JtloA87w9_1),.clk(gclk));
	jdff dff_B_XMzLTVwp1_1(.din(w_dff_B_JtloA87w9_1),.dout(w_dff_B_XMzLTVwp1_1),.clk(gclk));
	jdff dff_B_e0QxKCJC7_1(.din(w_dff_B_XMzLTVwp1_1),.dout(w_dff_B_e0QxKCJC7_1),.clk(gclk));
	jdff dff_B_fYxI2bvJ1_1(.din(w_dff_B_e0QxKCJC7_1),.dout(w_dff_B_fYxI2bvJ1_1),.clk(gclk));
	jdff dff_B_29qVH3sF3_1(.din(w_dff_B_fYxI2bvJ1_1),.dout(w_dff_B_29qVH3sF3_1),.clk(gclk));
	jdff dff_B_yDHr625w2_1(.din(w_dff_B_29qVH3sF3_1),.dout(w_dff_B_yDHr625w2_1),.clk(gclk));
	jdff dff_B_2nt6yQUH0_1(.din(w_dff_B_yDHr625w2_1),.dout(w_dff_B_2nt6yQUH0_1),.clk(gclk));
	jdff dff_B_BMA8R8kp0_1(.din(w_dff_B_2nt6yQUH0_1),.dout(w_dff_B_BMA8R8kp0_1),.clk(gclk));
	jdff dff_B_CWvGASmY1_1(.din(w_dff_B_BMA8R8kp0_1),.dout(w_dff_B_CWvGASmY1_1),.clk(gclk));
	jdff dff_B_zXeAHdLL5_1(.din(w_dff_B_CWvGASmY1_1),.dout(w_dff_B_zXeAHdLL5_1),.clk(gclk));
	jdff dff_B_iCcYTe8i1_1(.din(w_dff_B_zXeAHdLL5_1),.dout(w_dff_B_iCcYTe8i1_1),.clk(gclk));
	jdff dff_B_KKQakevS5_0(.din(n835),.dout(w_dff_B_KKQakevS5_0),.clk(gclk));
	jdff dff_B_IhDGF9wD5_0(.din(w_dff_B_KKQakevS5_0),.dout(w_dff_B_IhDGF9wD5_0),.clk(gclk));
	jdff dff_B_4RNSSUwD7_0(.din(w_dff_B_IhDGF9wD5_0),.dout(w_dff_B_4RNSSUwD7_0),.clk(gclk));
	jdff dff_B_pJYJVPvG1_0(.din(w_dff_B_4RNSSUwD7_0),.dout(w_dff_B_pJYJVPvG1_0),.clk(gclk));
	jdff dff_B_MeZqI1Vs8_0(.din(w_dff_B_pJYJVPvG1_0),.dout(w_dff_B_MeZqI1Vs8_0),.clk(gclk));
	jdff dff_B_NUmgf4hR3_0(.din(w_dff_B_MeZqI1Vs8_0),.dout(w_dff_B_NUmgf4hR3_0),.clk(gclk));
	jdff dff_B_NaEsykuF6_0(.din(w_dff_B_NUmgf4hR3_0),.dout(w_dff_B_NaEsykuF6_0),.clk(gclk));
	jdff dff_B_djV25LEY0_0(.din(w_dff_B_NaEsykuF6_0),.dout(w_dff_B_djV25LEY0_0),.clk(gclk));
	jdff dff_B_5Ye4GQGV8_0(.din(w_dff_B_djV25LEY0_0),.dout(w_dff_B_5Ye4GQGV8_0),.clk(gclk));
	jdff dff_B_S1Ux8Jpl1_0(.din(w_dff_B_5Ye4GQGV8_0),.dout(w_dff_B_S1Ux8Jpl1_0),.clk(gclk));
	jdff dff_B_BuJDb4Zd8_0(.din(w_dff_B_S1Ux8Jpl1_0),.dout(w_dff_B_BuJDb4Zd8_0),.clk(gclk));
	jdff dff_B_vyYoU76S7_0(.din(w_dff_B_BuJDb4Zd8_0),.dout(w_dff_B_vyYoU76S7_0),.clk(gclk));
	jdff dff_B_j4eDO0iq0_0(.din(w_dff_B_vyYoU76S7_0),.dout(w_dff_B_j4eDO0iq0_0),.clk(gclk));
	jdff dff_B_vzYntVQH4_0(.din(w_dff_B_j4eDO0iq0_0),.dout(w_dff_B_vzYntVQH4_0),.clk(gclk));
	jdff dff_B_DhLw4Sf48_0(.din(w_dff_B_vzYntVQH4_0),.dout(w_dff_B_DhLw4Sf48_0),.clk(gclk));
	jdff dff_B_kRnq9FQR5_0(.din(w_dff_B_DhLw4Sf48_0),.dout(w_dff_B_kRnq9FQR5_0),.clk(gclk));
	jdff dff_B_Clh0ZgdA4_0(.din(w_dff_B_kRnq9FQR5_0),.dout(w_dff_B_Clh0ZgdA4_0),.clk(gclk));
	jdff dff_B_s7LPLWVc3_0(.din(w_dff_B_Clh0ZgdA4_0),.dout(w_dff_B_s7LPLWVc3_0),.clk(gclk));
	jdff dff_B_HUEhu5CO6_0(.din(w_dff_B_s7LPLWVc3_0),.dout(w_dff_B_HUEhu5CO6_0),.clk(gclk));
	jdff dff_B_4ABZhlbX6_0(.din(w_dff_B_HUEhu5CO6_0),.dout(w_dff_B_4ABZhlbX6_0),.clk(gclk));
	jdff dff_B_t4q3b0OU9_0(.din(w_dff_B_4ABZhlbX6_0),.dout(w_dff_B_t4q3b0OU9_0),.clk(gclk));
	jdff dff_B_l9eIGpDQ4_0(.din(w_dff_B_t4q3b0OU9_0),.dout(w_dff_B_l9eIGpDQ4_0),.clk(gclk));
	jdff dff_B_I20CSoCB9_0(.din(w_dff_B_l9eIGpDQ4_0),.dout(w_dff_B_I20CSoCB9_0),.clk(gclk));
	jdff dff_B_w5YhRXmd8_0(.din(w_dff_B_I20CSoCB9_0),.dout(w_dff_B_w5YhRXmd8_0),.clk(gclk));
	jdff dff_B_en541yeg8_0(.din(w_dff_B_w5YhRXmd8_0),.dout(w_dff_B_en541yeg8_0),.clk(gclk));
	jdff dff_B_wdo74DPK9_0(.din(w_dff_B_en541yeg8_0),.dout(w_dff_B_wdo74DPK9_0),.clk(gclk));
	jdff dff_B_KQ7vyMZB6_0(.din(w_dff_B_wdo74DPK9_0),.dout(w_dff_B_KQ7vyMZB6_0),.clk(gclk));
	jdff dff_B_QqJtAtlP6_0(.din(w_dff_B_KQ7vyMZB6_0),.dout(w_dff_B_QqJtAtlP6_0),.clk(gclk));
	jdff dff_B_HpDSNcJq8_0(.din(w_dff_B_QqJtAtlP6_0),.dout(w_dff_B_HpDSNcJq8_0),.clk(gclk));
	jdff dff_B_nhUFAeSf1_0(.din(w_dff_B_HpDSNcJq8_0),.dout(w_dff_B_nhUFAeSf1_0),.clk(gclk));
	jdff dff_B_Lrerls4A4_0(.din(w_dff_B_nhUFAeSf1_0),.dout(w_dff_B_Lrerls4A4_0),.clk(gclk));
	jdff dff_B_yL4zEJyM6_0(.din(w_dff_B_Lrerls4A4_0),.dout(w_dff_B_yL4zEJyM6_0),.clk(gclk));
	jdff dff_B_YUfHx6So4_0(.din(w_dff_B_yL4zEJyM6_0),.dout(w_dff_B_YUfHx6So4_0),.clk(gclk));
	jdff dff_B_co16vS2v1_0(.din(w_dff_B_YUfHx6So4_0),.dout(w_dff_B_co16vS2v1_0),.clk(gclk));
	jdff dff_B_eJ5ImPck9_0(.din(w_dff_B_co16vS2v1_0),.dout(w_dff_B_eJ5ImPck9_0),.clk(gclk));
	jdff dff_B_GvsBcK7a3_0(.din(w_dff_B_eJ5ImPck9_0),.dout(w_dff_B_GvsBcK7a3_0),.clk(gclk));
	jdff dff_B_DDvavwnA4_0(.din(w_dff_B_GvsBcK7a3_0),.dout(w_dff_B_DDvavwnA4_0),.clk(gclk));
	jdff dff_B_XG1tvJuA4_0(.din(w_dff_B_DDvavwnA4_0),.dout(w_dff_B_XG1tvJuA4_0),.clk(gclk));
	jdff dff_B_i4gwd2VF1_0(.din(w_dff_B_XG1tvJuA4_0),.dout(w_dff_B_i4gwd2VF1_0),.clk(gclk));
	jdff dff_B_OOAWPb6Z3_0(.din(w_dff_B_i4gwd2VF1_0),.dout(w_dff_B_OOAWPb6Z3_0),.clk(gclk));
	jdff dff_B_Df0fWIFc7_0(.din(w_dff_B_OOAWPb6Z3_0),.dout(w_dff_B_Df0fWIFc7_0),.clk(gclk));
	jdff dff_B_hHnVT1au1_0(.din(w_dff_B_Df0fWIFc7_0),.dout(w_dff_B_hHnVT1au1_0),.clk(gclk));
	jdff dff_B_gGPz1dSO0_0(.din(w_dff_B_hHnVT1au1_0),.dout(w_dff_B_gGPz1dSO0_0),.clk(gclk));
	jdff dff_B_kQFMvZhe5_0(.din(w_dff_B_gGPz1dSO0_0),.dout(w_dff_B_kQFMvZhe5_0),.clk(gclk));
	jdff dff_B_bUueOIPZ0_0(.din(w_dff_B_kQFMvZhe5_0),.dout(w_dff_B_bUueOIPZ0_0),.clk(gclk));
	jdff dff_B_PfqZblfI4_0(.din(w_dff_B_bUueOIPZ0_0),.dout(w_dff_B_PfqZblfI4_0),.clk(gclk));
	jdff dff_B_J0s7zKTJ6_0(.din(w_dff_B_PfqZblfI4_0),.dout(w_dff_B_J0s7zKTJ6_0),.clk(gclk));
	jdff dff_B_lmfqUDMB1_0(.din(w_dff_B_J0s7zKTJ6_0),.dout(w_dff_B_lmfqUDMB1_0),.clk(gclk));
	jdff dff_B_LVKqfL9B0_0(.din(w_dff_B_lmfqUDMB1_0),.dout(w_dff_B_LVKqfL9B0_0),.clk(gclk));
	jdff dff_B_q7Ocs7Ei2_0(.din(w_dff_B_LVKqfL9B0_0),.dout(w_dff_B_q7Ocs7Ei2_0),.clk(gclk));
	jdff dff_B_kW0hc2Fd0_0(.din(w_dff_B_q7Ocs7Ei2_0),.dout(w_dff_B_kW0hc2Fd0_0),.clk(gclk));
	jdff dff_B_kOk8aa1D3_0(.din(w_dff_B_kW0hc2Fd0_0),.dout(w_dff_B_kOk8aa1D3_0),.clk(gclk));
	jdff dff_B_4Mppnres1_0(.din(w_dff_B_kOk8aa1D3_0),.dout(w_dff_B_4Mppnres1_0),.clk(gclk));
	jdff dff_B_u23GWRg08_0(.din(w_dff_B_4Mppnres1_0),.dout(w_dff_B_u23GWRg08_0),.clk(gclk));
	jdff dff_B_JQaMCbOl3_0(.din(w_dff_B_u23GWRg08_0),.dout(w_dff_B_JQaMCbOl3_0),.clk(gclk));
	jdff dff_B_tzwRobKE2_0(.din(w_dff_B_JQaMCbOl3_0),.dout(w_dff_B_tzwRobKE2_0),.clk(gclk));
	jdff dff_B_6GPTC3jI3_0(.din(w_dff_B_tzwRobKE2_0),.dout(w_dff_B_6GPTC3jI3_0),.clk(gclk));
	jdff dff_B_0A23CzIg8_0(.din(w_dff_B_6GPTC3jI3_0),.dout(w_dff_B_0A23CzIg8_0),.clk(gclk));
	jdff dff_B_1gHyfTLa9_0(.din(w_dff_B_0A23CzIg8_0),.dout(w_dff_B_1gHyfTLa9_0),.clk(gclk));
	jdff dff_B_VBw2aKEP2_0(.din(w_dff_B_1gHyfTLa9_0),.dout(w_dff_B_VBw2aKEP2_0),.clk(gclk));
	jdff dff_B_DttoBILE6_0(.din(w_dff_B_VBw2aKEP2_0),.dout(w_dff_B_DttoBILE6_0),.clk(gclk));
	jdff dff_B_Qop7ZEK13_0(.din(w_dff_B_DttoBILE6_0),.dout(w_dff_B_Qop7ZEK13_0),.clk(gclk));
	jdff dff_B_Sd9TXsMA3_0(.din(w_dff_B_Qop7ZEK13_0),.dout(w_dff_B_Sd9TXsMA3_0),.clk(gclk));
	jdff dff_B_nXZZwd4K5_0(.din(w_dff_B_Sd9TXsMA3_0),.dout(w_dff_B_nXZZwd4K5_0),.clk(gclk));
	jdff dff_B_NmUpZhn23_0(.din(w_dff_B_nXZZwd4K5_0),.dout(w_dff_B_NmUpZhn23_0),.clk(gclk));
	jdff dff_B_YO3I10x21_0(.din(w_dff_B_NmUpZhn23_0),.dout(w_dff_B_YO3I10x21_0),.clk(gclk));
	jdff dff_B_uLZagXrY4_0(.din(w_dff_B_YO3I10x21_0),.dout(w_dff_B_uLZagXrY4_0),.clk(gclk));
	jdff dff_B_0adFijnY2_0(.din(w_dff_B_uLZagXrY4_0),.dout(w_dff_B_0adFijnY2_0),.clk(gclk));
	jdff dff_B_OPUjSWhz6_0(.din(w_dff_B_0adFijnY2_0),.dout(w_dff_B_OPUjSWhz6_0),.clk(gclk));
	jdff dff_B_vBjknD2k1_0(.din(w_dff_B_OPUjSWhz6_0),.dout(w_dff_B_vBjknD2k1_0),.clk(gclk));
	jdff dff_B_Ze6FlNRD1_0(.din(w_dff_B_vBjknD2k1_0),.dout(w_dff_B_Ze6FlNRD1_0),.clk(gclk));
	jdff dff_B_ZGHgKduP7_0(.din(w_dff_B_Ze6FlNRD1_0),.dout(w_dff_B_ZGHgKduP7_0),.clk(gclk));
	jdff dff_B_6xRazE0Z0_0(.din(w_dff_B_ZGHgKduP7_0),.dout(w_dff_B_6xRazE0Z0_0),.clk(gclk));
	jdff dff_B_1LX0OJy92_0(.din(w_dff_B_6xRazE0Z0_0),.dout(w_dff_B_1LX0OJy92_0),.clk(gclk));
	jdff dff_B_eQj5PWyb8_0(.din(w_dff_B_1LX0OJy92_0),.dout(w_dff_B_eQj5PWyb8_0),.clk(gclk));
	jdff dff_B_fzcQWGjQ1_1(.din(n828),.dout(w_dff_B_fzcQWGjQ1_1),.clk(gclk));
	jdff dff_B_iWqqy8Ef0_1(.din(w_dff_B_fzcQWGjQ1_1),.dout(w_dff_B_iWqqy8Ef0_1),.clk(gclk));
	jdff dff_B_9Av6yP9T3_1(.din(w_dff_B_iWqqy8Ef0_1),.dout(w_dff_B_9Av6yP9T3_1),.clk(gclk));
	jdff dff_B_YXx2SfdY1_1(.din(w_dff_B_9Av6yP9T3_1),.dout(w_dff_B_YXx2SfdY1_1),.clk(gclk));
	jdff dff_B_oIYmjxts5_1(.din(w_dff_B_YXx2SfdY1_1),.dout(w_dff_B_oIYmjxts5_1),.clk(gclk));
	jdff dff_B_p8yNM6qJ2_1(.din(w_dff_B_oIYmjxts5_1),.dout(w_dff_B_p8yNM6qJ2_1),.clk(gclk));
	jdff dff_B_FCCUOyOc5_1(.din(w_dff_B_p8yNM6qJ2_1),.dout(w_dff_B_FCCUOyOc5_1),.clk(gclk));
	jdff dff_B_QT1NzXQi2_1(.din(w_dff_B_FCCUOyOc5_1),.dout(w_dff_B_QT1NzXQi2_1),.clk(gclk));
	jdff dff_B_U8HTmwp55_1(.din(w_dff_B_QT1NzXQi2_1),.dout(w_dff_B_U8HTmwp55_1),.clk(gclk));
	jdff dff_B_FUmWtdDH4_1(.din(w_dff_B_U8HTmwp55_1),.dout(w_dff_B_FUmWtdDH4_1),.clk(gclk));
	jdff dff_B_MEOVQKAS1_1(.din(w_dff_B_FUmWtdDH4_1),.dout(w_dff_B_MEOVQKAS1_1),.clk(gclk));
	jdff dff_B_UdPpq5NB9_1(.din(w_dff_B_MEOVQKAS1_1),.dout(w_dff_B_UdPpq5NB9_1),.clk(gclk));
	jdff dff_B_Mhc9hgNk9_1(.din(w_dff_B_UdPpq5NB9_1),.dout(w_dff_B_Mhc9hgNk9_1),.clk(gclk));
	jdff dff_B_Qapas9H97_1(.din(w_dff_B_Mhc9hgNk9_1),.dout(w_dff_B_Qapas9H97_1),.clk(gclk));
	jdff dff_B_eLBOgaF59_1(.din(w_dff_B_Qapas9H97_1),.dout(w_dff_B_eLBOgaF59_1),.clk(gclk));
	jdff dff_B_MoASXsnZ0_1(.din(w_dff_B_eLBOgaF59_1),.dout(w_dff_B_MoASXsnZ0_1),.clk(gclk));
	jdff dff_B_5jhs2Gql9_1(.din(w_dff_B_MoASXsnZ0_1),.dout(w_dff_B_5jhs2Gql9_1),.clk(gclk));
	jdff dff_B_rHroq8Um7_1(.din(w_dff_B_5jhs2Gql9_1),.dout(w_dff_B_rHroq8Um7_1),.clk(gclk));
	jdff dff_B_hM0BHclV2_1(.din(w_dff_B_rHroq8Um7_1),.dout(w_dff_B_hM0BHclV2_1),.clk(gclk));
	jdff dff_B_XIoaE5mR7_1(.din(w_dff_B_hM0BHclV2_1),.dout(w_dff_B_XIoaE5mR7_1),.clk(gclk));
	jdff dff_B_5orr76Oy5_1(.din(w_dff_B_XIoaE5mR7_1),.dout(w_dff_B_5orr76Oy5_1),.clk(gclk));
	jdff dff_B_MBvwhF022_1(.din(w_dff_B_5orr76Oy5_1),.dout(w_dff_B_MBvwhF022_1),.clk(gclk));
	jdff dff_B_1ZAhBf8L2_1(.din(w_dff_B_MBvwhF022_1),.dout(w_dff_B_1ZAhBf8L2_1),.clk(gclk));
	jdff dff_B_on9oBKIb0_1(.din(w_dff_B_1ZAhBf8L2_1),.dout(w_dff_B_on9oBKIb0_1),.clk(gclk));
	jdff dff_B_nuwwpKgZ5_1(.din(w_dff_B_on9oBKIb0_1),.dout(w_dff_B_nuwwpKgZ5_1),.clk(gclk));
	jdff dff_B_Ce1x3yho2_1(.din(w_dff_B_nuwwpKgZ5_1),.dout(w_dff_B_Ce1x3yho2_1),.clk(gclk));
	jdff dff_B_DhjtPnGr8_1(.din(w_dff_B_Ce1x3yho2_1),.dout(w_dff_B_DhjtPnGr8_1),.clk(gclk));
	jdff dff_B_2oCfYTSA5_1(.din(w_dff_B_DhjtPnGr8_1),.dout(w_dff_B_2oCfYTSA5_1),.clk(gclk));
	jdff dff_B_Xm2qg5Nn8_1(.din(w_dff_B_2oCfYTSA5_1),.dout(w_dff_B_Xm2qg5Nn8_1),.clk(gclk));
	jdff dff_B_CAmA70hQ5_1(.din(w_dff_B_Xm2qg5Nn8_1),.dout(w_dff_B_CAmA70hQ5_1),.clk(gclk));
	jdff dff_B_Ql0RvhiW8_1(.din(w_dff_B_CAmA70hQ5_1),.dout(w_dff_B_Ql0RvhiW8_1),.clk(gclk));
	jdff dff_B_UD7L9CII8_1(.din(w_dff_B_Ql0RvhiW8_1),.dout(w_dff_B_UD7L9CII8_1),.clk(gclk));
	jdff dff_B_CpsaaURa7_1(.din(w_dff_B_UD7L9CII8_1),.dout(w_dff_B_CpsaaURa7_1),.clk(gclk));
	jdff dff_B_VSOnUax70_1(.din(w_dff_B_CpsaaURa7_1),.dout(w_dff_B_VSOnUax70_1),.clk(gclk));
	jdff dff_B_bTZjxV3X9_1(.din(w_dff_B_VSOnUax70_1),.dout(w_dff_B_bTZjxV3X9_1),.clk(gclk));
	jdff dff_B_m9XojbnU1_1(.din(w_dff_B_bTZjxV3X9_1),.dout(w_dff_B_m9XojbnU1_1),.clk(gclk));
	jdff dff_B_ec05QcVN4_1(.din(w_dff_B_m9XojbnU1_1),.dout(w_dff_B_ec05QcVN4_1),.clk(gclk));
	jdff dff_B_UWWylQYY9_1(.din(w_dff_B_ec05QcVN4_1),.dout(w_dff_B_UWWylQYY9_1),.clk(gclk));
	jdff dff_B_UBv1pgTI6_1(.din(w_dff_B_UWWylQYY9_1),.dout(w_dff_B_UBv1pgTI6_1),.clk(gclk));
	jdff dff_B_93kHH1z81_1(.din(w_dff_B_UBv1pgTI6_1),.dout(w_dff_B_93kHH1z81_1),.clk(gclk));
	jdff dff_B_vh4YDzLy3_1(.din(w_dff_B_93kHH1z81_1),.dout(w_dff_B_vh4YDzLy3_1),.clk(gclk));
	jdff dff_B_ngm6uAAi4_1(.din(w_dff_B_vh4YDzLy3_1),.dout(w_dff_B_ngm6uAAi4_1),.clk(gclk));
	jdff dff_B_0H8Cm9Ip6_1(.din(w_dff_B_ngm6uAAi4_1),.dout(w_dff_B_0H8Cm9Ip6_1),.clk(gclk));
	jdff dff_B_li0ODhpa9_1(.din(w_dff_B_0H8Cm9Ip6_1),.dout(w_dff_B_li0ODhpa9_1),.clk(gclk));
	jdff dff_B_ICpyKWgS1_1(.din(w_dff_B_li0ODhpa9_1),.dout(w_dff_B_ICpyKWgS1_1),.clk(gclk));
	jdff dff_B_POTFi3md5_1(.din(w_dff_B_ICpyKWgS1_1),.dout(w_dff_B_POTFi3md5_1),.clk(gclk));
	jdff dff_B_pXRCJx5B8_1(.din(w_dff_B_POTFi3md5_1),.dout(w_dff_B_pXRCJx5B8_1),.clk(gclk));
	jdff dff_B_g56UXDze6_1(.din(w_dff_B_pXRCJx5B8_1),.dout(w_dff_B_g56UXDze6_1),.clk(gclk));
	jdff dff_B_0Gx8e77j0_1(.din(w_dff_B_g56UXDze6_1),.dout(w_dff_B_0Gx8e77j0_1),.clk(gclk));
	jdff dff_B_JWiXsLj33_1(.din(w_dff_B_0Gx8e77j0_1),.dout(w_dff_B_JWiXsLj33_1),.clk(gclk));
	jdff dff_B_HdJm9LvW7_1(.din(w_dff_B_JWiXsLj33_1),.dout(w_dff_B_HdJm9LvW7_1),.clk(gclk));
	jdff dff_B_WiI54ckC1_1(.din(w_dff_B_HdJm9LvW7_1),.dout(w_dff_B_WiI54ckC1_1),.clk(gclk));
	jdff dff_B_WTtqsecn6_1(.din(w_dff_B_WiI54ckC1_1),.dout(w_dff_B_WTtqsecn6_1),.clk(gclk));
	jdff dff_B_idsXCX3d9_1(.din(w_dff_B_WTtqsecn6_1),.dout(w_dff_B_idsXCX3d9_1),.clk(gclk));
	jdff dff_B_y2F4RiEV4_1(.din(w_dff_B_idsXCX3d9_1),.dout(w_dff_B_y2F4RiEV4_1),.clk(gclk));
	jdff dff_B_11Vt3sBK0_1(.din(w_dff_B_y2F4RiEV4_1),.dout(w_dff_B_11Vt3sBK0_1),.clk(gclk));
	jdff dff_B_wM9oTRtT9_1(.din(w_dff_B_11Vt3sBK0_1),.dout(w_dff_B_wM9oTRtT9_1),.clk(gclk));
	jdff dff_B_aaiF4Yzg2_1(.din(w_dff_B_wM9oTRtT9_1),.dout(w_dff_B_aaiF4Yzg2_1),.clk(gclk));
	jdff dff_B_WJdfKBfg4_1(.din(w_dff_B_aaiF4Yzg2_1),.dout(w_dff_B_WJdfKBfg4_1),.clk(gclk));
	jdff dff_B_cwwrwLCm6_1(.din(w_dff_B_WJdfKBfg4_1),.dout(w_dff_B_cwwrwLCm6_1),.clk(gclk));
	jdff dff_B_Y6qNhR5p3_1(.din(w_dff_B_cwwrwLCm6_1),.dout(w_dff_B_Y6qNhR5p3_1),.clk(gclk));
	jdff dff_B_sUdhBr9E5_1(.din(w_dff_B_Y6qNhR5p3_1),.dout(w_dff_B_sUdhBr9E5_1),.clk(gclk));
	jdff dff_B_cA5cZ6907_1(.din(w_dff_B_sUdhBr9E5_1),.dout(w_dff_B_cA5cZ6907_1),.clk(gclk));
	jdff dff_B_b9BLn1h61_1(.din(w_dff_B_cA5cZ6907_1),.dout(w_dff_B_b9BLn1h61_1),.clk(gclk));
	jdff dff_B_hnEdSN8A2_1(.din(w_dff_B_b9BLn1h61_1),.dout(w_dff_B_hnEdSN8A2_1),.clk(gclk));
	jdff dff_B_W7FVO3aG1_1(.din(w_dff_B_hnEdSN8A2_1),.dout(w_dff_B_W7FVO3aG1_1),.clk(gclk));
	jdff dff_B_9cvDDs469_1(.din(w_dff_B_W7FVO3aG1_1),.dout(w_dff_B_9cvDDs469_1),.clk(gclk));
	jdff dff_B_2K7tkW5v1_1(.din(w_dff_B_9cvDDs469_1),.dout(w_dff_B_2K7tkW5v1_1),.clk(gclk));
	jdff dff_B_pbgoh5Qd8_1(.din(w_dff_B_2K7tkW5v1_1),.dout(w_dff_B_pbgoh5Qd8_1),.clk(gclk));
	jdff dff_B_rBwhVI587_1(.din(w_dff_B_pbgoh5Qd8_1),.dout(w_dff_B_rBwhVI587_1),.clk(gclk));
	jdff dff_B_cVeA81v10_1(.din(w_dff_B_rBwhVI587_1),.dout(w_dff_B_cVeA81v10_1),.clk(gclk));
	jdff dff_B_c4AgP0Gh0_1(.din(w_dff_B_cVeA81v10_1),.dout(w_dff_B_c4AgP0Gh0_1),.clk(gclk));
	jdff dff_B_h5ChKpm86_1(.din(w_dff_B_c4AgP0Gh0_1),.dout(w_dff_B_h5ChKpm86_1),.clk(gclk));
	jdff dff_B_yknhl01q3_1(.din(w_dff_B_h5ChKpm86_1),.dout(w_dff_B_yknhl01q3_1),.clk(gclk));
	jdff dff_B_NXdUOz5k1_0(.din(n829),.dout(w_dff_B_NXdUOz5k1_0),.clk(gclk));
	jdff dff_B_rvLNVcuE6_0(.din(w_dff_B_NXdUOz5k1_0),.dout(w_dff_B_rvLNVcuE6_0),.clk(gclk));
	jdff dff_B_gHuqydpu1_0(.din(w_dff_B_rvLNVcuE6_0),.dout(w_dff_B_gHuqydpu1_0),.clk(gclk));
	jdff dff_B_Womz66i84_0(.din(w_dff_B_gHuqydpu1_0),.dout(w_dff_B_Womz66i84_0),.clk(gclk));
	jdff dff_B_AyNzqpIh4_0(.din(w_dff_B_Womz66i84_0),.dout(w_dff_B_AyNzqpIh4_0),.clk(gclk));
	jdff dff_B_AXGHcgiM1_0(.din(w_dff_B_AyNzqpIh4_0),.dout(w_dff_B_AXGHcgiM1_0),.clk(gclk));
	jdff dff_B_OLgFLNcu7_0(.din(w_dff_B_AXGHcgiM1_0),.dout(w_dff_B_OLgFLNcu7_0),.clk(gclk));
	jdff dff_B_fGmBEd840_0(.din(w_dff_B_OLgFLNcu7_0),.dout(w_dff_B_fGmBEd840_0),.clk(gclk));
	jdff dff_B_LAE4i4Nd7_0(.din(w_dff_B_fGmBEd840_0),.dout(w_dff_B_LAE4i4Nd7_0),.clk(gclk));
	jdff dff_B_5nYvM20E9_0(.din(w_dff_B_LAE4i4Nd7_0),.dout(w_dff_B_5nYvM20E9_0),.clk(gclk));
	jdff dff_B_FLISnqZ31_0(.din(w_dff_B_5nYvM20E9_0),.dout(w_dff_B_FLISnqZ31_0),.clk(gclk));
	jdff dff_B_kgskhX5U8_0(.din(w_dff_B_FLISnqZ31_0),.dout(w_dff_B_kgskhX5U8_0),.clk(gclk));
	jdff dff_B_pseM8KBi5_0(.din(w_dff_B_kgskhX5U8_0),.dout(w_dff_B_pseM8KBi5_0),.clk(gclk));
	jdff dff_B_NCZ3iCjn1_0(.din(w_dff_B_pseM8KBi5_0),.dout(w_dff_B_NCZ3iCjn1_0),.clk(gclk));
	jdff dff_B_yfd8K9kw0_0(.din(w_dff_B_NCZ3iCjn1_0),.dout(w_dff_B_yfd8K9kw0_0),.clk(gclk));
	jdff dff_B_soHwuBmQ0_0(.din(w_dff_B_yfd8K9kw0_0),.dout(w_dff_B_soHwuBmQ0_0),.clk(gclk));
	jdff dff_B_ttlUcDMf3_0(.din(w_dff_B_soHwuBmQ0_0),.dout(w_dff_B_ttlUcDMf3_0),.clk(gclk));
	jdff dff_B_wDJ7CNjL7_0(.din(w_dff_B_ttlUcDMf3_0),.dout(w_dff_B_wDJ7CNjL7_0),.clk(gclk));
	jdff dff_B_DBH5LdSb4_0(.din(w_dff_B_wDJ7CNjL7_0),.dout(w_dff_B_DBH5LdSb4_0),.clk(gclk));
	jdff dff_B_aSbcZRhu5_0(.din(w_dff_B_DBH5LdSb4_0),.dout(w_dff_B_aSbcZRhu5_0),.clk(gclk));
	jdff dff_B_BU8ADFap7_0(.din(w_dff_B_aSbcZRhu5_0),.dout(w_dff_B_BU8ADFap7_0),.clk(gclk));
	jdff dff_B_2QBwY8623_0(.din(w_dff_B_BU8ADFap7_0),.dout(w_dff_B_2QBwY8623_0),.clk(gclk));
	jdff dff_B_NMCoNdre5_0(.din(w_dff_B_2QBwY8623_0),.dout(w_dff_B_NMCoNdre5_0),.clk(gclk));
	jdff dff_B_4JlLuIGm7_0(.din(w_dff_B_NMCoNdre5_0),.dout(w_dff_B_4JlLuIGm7_0),.clk(gclk));
	jdff dff_B_7k2r6Ht79_0(.din(w_dff_B_4JlLuIGm7_0),.dout(w_dff_B_7k2r6Ht79_0),.clk(gclk));
	jdff dff_B_kuLBzDew0_0(.din(w_dff_B_7k2r6Ht79_0),.dout(w_dff_B_kuLBzDew0_0),.clk(gclk));
	jdff dff_B_VbRP7utx1_0(.din(w_dff_B_kuLBzDew0_0),.dout(w_dff_B_VbRP7utx1_0),.clk(gclk));
	jdff dff_B_BgjkTimB9_0(.din(w_dff_B_VbRP7utx1_0),.dout(w_dff_B_BgjkTimB9_0),.clk(gclk));
	jdff dff_B_pOWyAVL76_0(.din(w_dff_B_BgjkTimB9_0),.dout(w_dff_B_pOWyAVL76_0),.clk(gclk));
	jdff dff_B_txbNW4CK3_0(.din(w_dff_B_pOWyAVL76_0),.dout(w_dff_B_txbNW4CK3_0),.clk(gclk));
	jdff dff_B_8YcG4hoe3_0(.din(w_dff_B_txbNW4CK3_0),.dout(w_dff_B_8YcG4hoe3_0),.clk(gclk));
	jdff dff_B_VHsc707M3_0(.din(w_dff_B_8YcG4hoe3_0),.dout(w_dff_B_VHsc707M3_0),.clk(gclk));
	jdff dff_B_FoqpMuCn2_0(.din(w_dff_B_VHsc707M3_0),.dout(w_dff_B_FoqpMuCn2_0),.clk(gclk));
	jdff dff_B_MOUfJ2bf1_0(.din(w_dff_B_FoqpMuCn2_0),.dout(w_dff_B_MOUfJ2bf1_0),.clk(gclk));
	jdff dff_B_zKYMz6YK5_0(.din(w_dff_B_MOUfJ2bf1_0),.dout(w_dff_B_zKYMz6YK5_0),.clk(gclk));
	jdff dff_B_W1CSDG8t9_0(.din(w_dff_B_zKYMz6YK5_0),.dout(w_dff_B_W1CSDG8t9_0),.clk(gclk));
	jdff dff_B_lkMNodfX8_0(.din(w_dff_B_W1CSDG8t9_0),.dout(w_dff_B_lkMNodfX8_0),.clk(gclk));
	jdff dff_B_DeuUb19m8_0(.din(w_dff_B_lkMNodfX8_0),.dout(w_dff_B_DeuUb19m8_0),.clk(gclk));
	jdff dff_B_2T2l4kmR7_0(.din(w_dff_B_DeuUb19m8_0),.dout(w_dff_B_2T2l4kmR7_0),.clk(gclk));
	jdff dff_B_vildeu6e0_0(.din(w_dff_B_2T2l4kmR7_0),.dout(w_dff_B_vildeu6e0_0),.clk(gclk));
	jdff dff_B_CG00E0vw7_0(.din(w_dff_B_vildeu6e0_0),.dout(w_dff_B_CG00E0vw7_0),.clk(gclk));
	jdff dff_B_ApCQjulg9_0(.din(w_dff_B_CG00E0vw7_0),.dout(w_dff_B_ApCQjulg9_0),.clk(gclk));
	jdff dff_B_74o4HdjE8_0(.din(w_dff_B_ApCQjulg9_0),.dout(w_dff_B_74o4HdjE8_0),.clk(gclk));
	jdff dff_B_zDCkAEWQ3_0(.din(w_dff_B_74o4HdjE8_0),.dout(w_dff_B_zDCkAEWQ3_0),.clk(gclk));
	jdff dff_B_fK4nLh8r9_0(.din(w_dff_B_zDCkAEWQ3_0),.dout(w_dff_B_fK4nLh8r9_0),.clk(gclk));
	jdff dff_B_3fBo5HpL0_0(.din(w_dff_B_fK4nLh8r9_0),.dout(w_dff_B_3fBo5HpL0_0),.clk(gclk));
	jdff dff_B_FKZmoGFT1_0(.din(w_dff_B_3fBo5HpL0_0),.dout(w_dff_B_FKZmoGFT1_0),.clk(gclk));
	jdff dff_B_UShcwkED6_0(.din(w_dff_B_FKZmoGFT1_0),.dout(w_dff_B_UShcwkED6_0),.clk(gclk));
	jdff dff_B_4PUDOwNs3_0(.din(w_dff_B_UShcwkED6_0),.dout(w_dff_B_4PUDOwNs3_0),.clk(gclk));
	jdff dff_B_9Fa55XcT1_0(.din(w_dff_B_4PUDOwNs3_0),.dout(w_dff_B_9Fa55XcT1_0),.clk(gclk));
	jdff dff_B_sLTfuto52_0(.din(w_dff_B_9Fa55XcT1_0),.dout(w_dff_B_sLTfuto52_0),.clk(gclk));
	jdff dff_B_etjT0UeA0_0(.din(w_dff_B_sLTfuto52_0),.dout(w_dff_B_etjT0UeA0_0),.clk(gclk));
	jdff dff_B_nr2Yngns4_0(.din(w_dff_B_etjT0UeA0_0),.dout(w_dff_B_nr2Yngns4_0),.clk(gclk));
	jdff dff_B_ttamoL4V1_0(.din(w_dff_B_nr2Yngns4_0),.dout(w_dff_B_ttamoL4V1_0),.clk(gclk));
	jdff dff_B_40zbkknR9_0(.din(w_dff_B_ttamoL4V1_0),.dout(w_dff_B_40zbkknR9_0),.clk(gclk));
	jdff dff_B_0WwOXIgK8_0(.din(w_dff_B_40zbkknR9_0),.dout(w_dff_B_0WwOXIgK8_0),.clk(gclk));
	jdff dff_B_VKAWpe2X1_0(.din(w_dff_B_0WwOXIgK8_0),.dout(w_dff_B_VKAWpe2X1_0),.clk(gclk));
	jdff dff_B_uSx5Ur0E4_0(.din(w_dff_B_VKAWpe2X1_0),.dout(w_dff_B_uSx5Ur0E4_0),.clk(gclk));
	jdff dff_B_JDqwaRfV9_0(.din(w_dff_B_uSx5Ur0E4_0),.dout(w_dff_B_JDqwaRfV9_0),.clk(gclk));
	jdff dff_B_mo9r74Aw1_0(.din(w_dff_B_JDqwaRfV9_0),.dout(w_dff_B_mo9r74Aw1_0),.clk(gclk));
	jdff dff_B_J9W8VrJi2_0(.din(w_dff_B_mo9r74Aw1_0),.dout(w_dff_B_J9W8VrJi2_0),.clk(gclk));
	jdff dff_B_w1JhITiY6_0(.din(w_dff_B_J9W8VrJi2_0),.dout(w_dff_B_w1JhITiY6_0),.clk(gclk));
	jdff dff_B_3YhGHSeV9_0(.din(w_dff_B_w1JhITiY6_0),.dout(w_dff_B_3YhGHSeV9_0),.clk(gclk));
	jdff dff_B_T9IyBr3I4_0(.din(w_dff_B_3YhGHSeV9_0),.dout(w_dff_B_T9IyBr3I4_0),.clk(gclk));
	jdff dff_B_DRhjfae82_0(.din(w_dff_B_T9IyBr3I4_0),.dout(w_dff_B_DRhjfae82_0),.clk(gclk));
	jdff dff_B_G75xdA971_0(.din(w_dff_B_DRhjfae82_0),.dout(w_dff_B_G75xdA971_0),.clk(gclk));
	jdff dff_B_ZcdO2RPK4_0(.din(w_dff_B_G75xdA971_0),.dout(w_dff_B_ZcdO2RPK4_0),.clk(gclk));
	jdff dff_B_E2sDRwcC4_0(.din(w_dff_B_ZcdO2RPK4_0),.dout(w_dff_B_E2sDRwcC4_0),.clk(gclk));
	jdff dff_B_vnDJJop06_0(.din(w_dff_B_E2sDRwcC4_0),.dout(w_dff_B_vnDJJop06_0),.clk(gclk));
	jdff dff_B_6K4WLKcr8_0(.din(w_dff_B_vnDJJop06_0),.dout(w_dff_B_6K4WLKcr8_0),.clk(gclk));
	jdff dff_B_3n7DBwv68_0(.din(w_dff_B_6K4WLKcr8_0),.dout(w_dff_B_3n7DBwv68_0),.clk(gclk));
	jdff dff_B_7Ak4wJe99_0(.din(w_dff_B_3n7DBwv68_0),.dout(w_dff_B_7Ak4wJe99_0),.clk(gclk));
	jdff dff_B_PLV9oANz4_0(.din(w_dff_B_7Ak4wJe99_0),.dout(w_dff_B_PLV9oANz4_0),.clk(gclk));
	jdff dff_B_zTdSogfq8_0(.din(w_dff_B_PLV9oANz4_0),.dout(w_dff_B_zTdSogfq8_0),.clk(gclk));
	jdff dff_B_P1a241067_1(.din(n822),.dout(w_dff_B_P1a241067_1),.clk(gclk));
	jdff dff_B_WBtJ2fqY2_1(.din(w_dff_B_P1a241067_1),.dout(w_dff_B_WBtJ2fqY2_1),.clk(gclk));
	jdff dff_B_9jD9mowu5_1(.din(w_dff_B_WBtJ2fqY2_1),.dout(w_dff_B_9jD9mowu5_1),.clk(gclk));
	jdff dff_B_0fmoSMOy1_1(.din(w_dff_B_9jD9mowu5_1),.dout(w_dff_B_0fmoSMOy1_1),.clk(gclk));
	jdff dff_B_VTyKecC02_1(.din(w_dff_B_0fmoSMOy1_1),.dout(w_dff_B_VTyKecC02_1),.clk(gclk));
	jdff dff_B_4C4bnUWE3_1(.din(w_dff_B_VTyKecC02_1),.dout(w_dff_B_4C4bnUWE3_1),.clk(gclk));
	jdff dff_B_SKBPGTCL9_1(.din(w_dff_B_4C4bnUWE3_1),.dout(w_dff_B_SKBPGTCL9_1),.clk(gclk));
	jdff dff_B_OvVv21AE5_1(.din(w_dff_B_SKBPGTCL9_1),.dout(w_dff_B_OvVv21AE5_1),.clk(gclk));
	jdff dff_B_k11z6bDt0_1(.din(w_dff_B_OvVv21AE5_1),.dout(w_dff_B_k11z6bDt0_1),.clk(gclk));
	jdff dff_B_OQ1vd6TP3_1(.din(w_dff_B_k11z6bDt0_1),.dout(w_dff_B_OQ1vd6TP3_1),.clk(gclk));
	jdff dff_B_9Uxuewrh6_1(.din(w_dff_B_OQ1vd6TP3_1),.dout(w_dff_B_9Uxuewrh6_1),.clk(gclk));
	jdff dff_B_UQpsdQPT1_1(.din(w_dff_B_9Uxuewrh6_1),.dout(w_dff_B_UQpsdQPT1_1),.clk(gclk));
	jdff dff_B_3NH9F9hi3_1(.din(w_dff_B_UQpsdQPT1_1),.dout(w_dff_B_3NH9F9hi3_1),.clk(gclk));
	jdff dff_B_XDXpJEb01_1(.din(w_dff_B_3NH9F9hi3_1),.dout(w_dff_B_XDXpJEb01_1),.clk(gclk));
	jdff dff_B_G1DgOKdE8_1(.din(w_dff_B_XDXpJEb01_1),.dout(w_dff_B_G1DgOKdE8_1),.clk(gclk));
	jdff dff_B_pwewoXo13_1(.din(w_dff_B_G1DgOKdE8_1),.dout(w_dff_B_pwewoXo13_1),.clk(gclk));
	jdff dff_B_pAjrQGmh3_1(.din(w_dff_B_pwewoXo13_1),.dout(w_dff_B_pAjrQGmh3_1),.clk(gclk));
	jdff dff_B_Aw8S6JcH2_1(.din(w_dff_B_pAjrQGmh3_1),.dout(w_dff_B_Aw8S6JcH2_1),.clk(gclk));
	jdff dff_B_CKKMrjSH4_1(.din(w_dff_B_Aw8S6JcH2_1),.dout(w_dff_B_CKKMrjSH4_1),.clk(gclk));
	jdff dff_B_OiZm2VEm8_1(.din(w_dff_B_CKKMrjSH4_1),.dout(w_dff_B_OiZm2VEm8_1),.clk(gclk));
	jdff dff_B_A3iCMKUs1_1(.din(w_dff_B_OiZm2VEm8_1),.dout(w_dff_B_A3iCMKUs1_1),.clk(gclk));
	jdff dff_B_10It760G9_1(.din(w_dff_B_A3iCMKUs1_1),.dout(w_dff_B_10It760G9_1),.clk(gclk));
	jdff dff_B_DX4UyAc42_1(.din(w_dff_B_10It760G9_1),.dout(w_dff_B_DX4UyAc42_1),.clk(gclk));
	jdff dff_B_lU8vVODj6_1(.din(w_dff_B_DX4UyAc42_1),.dout(w_dff_B_lU8vVODj6_1),.clk(gclk));
	jdff dff_B_H2pjsWzT9_1(.din(w_dff_B_lU8vVODj6_1),.dout(w_dff_B_H2pjsWzT9_1),.clk(gclk));
	jdff dff_B_AcJPtQK80_1(.din(w_dff_B_H2pjsWzT9_1),.dout(w_dff_B_AcJPtQK80_1),.clk(gclk));
	jdff dff_B_bNtDkg091_1(.din(w_dff_B_AcJPtQK80_1),.dout(w_dff_B_bNtDkg091_1),.clk(gclk));
	jdff dff_B_YpFb5RHt5_1(.din(w_dff_B_bNtDkg091_1),.dout(w_dff_B_YpFb5RHt5_1),.clk(gclk));
	jdff dff_B_MwbFFXpn5_1(.din(w_dff_B_YpFb5RHt5_1),.dout(w_dff_B_MwbFFXpn5_1),.clk(gclk));
	jdff dff_B_MGixn9EF7_1(.din(w_dff_B_MwbFFXpn5_1),.dout(w_dff_B_MGixn9EF7_1),.clk(gclk));
	jdff dff_B_CrK3a6ka5_1(.din(w_dff_B_MGixn9EF7_1),.dout(w_dff_B_CrK3a6ka5_1),.clk(gclk));
	jdff dff_B_fADA8nPu2_1(.din(w_dff_B_CrK3a6ka5_1),.dout(w_dff_B_fADA8nPu2_1),.clk(gclk));
	jdff dff_B_iDDLOMSv5_1(.din(w_dff_B_fADA8nPu2_1),.dout(w_dff_B_iDDLOMSv5_1),.clk(gclk));
	jdff dff_B_bupoSeDY8_1(.din(w_dff_B_iDDLOMSv5_1),.dout(w_dff_B_bupoSeDY8_1),.clk(gclk));
	jdff dff_B_E9pOElhA6_1(.din(w_dff_B_bupoSeDY8_1),.dout(w_dff_B_E9pOElhA6_1),.clk(gclk));
	jdff dff_B_VPlwSNKi2_1(.din(w_dff_B_E9pOElhA6_1),.dout(w_dff_B_VPlwSNKi2_1),.clk(gclk));
	jdff dff_B_9UZzjdqH8_1(.din(w_dff_B_VPlwSNKi2_1),.dout(w_dff_B_9UZzjdqH8_1),.clk(gclk));
	jdff dff_B_N1eUPrLV7_1(.din(w_dff_B_9UZzjdqH8_1),.dout(w_dff_B_N1eUPrLV7_1),.clk(gclk));
	jdff dff_B_fXdK2AGn0_1(.din(w_dff_B_N1eUPrLV7_1),.dout(w_dff_B_fXdK2AGn0_1),.clk(gclk));
	jdff dff_B_mErZx3rd6_1(.din(w_dff_B_fXdK2AGn0_1),.dout(w_dff_B_mErZx3rd6_1),.clk(gclk));
	jdff dff_B_pe0G3Tzl6_1(.din(w_dff_B_mErZx3rd6_1),.dout(w_dff_B_pe0G3Tzl6_1),.clk(gclk));
	jdff dff_B_80W7Q4dK1_1(.din(w_dff_B_pe0G3Tzl6_1),.dout(w_dff_B_80W7Q4dK1_1),.clk(gclk));
	jdff dff_B_kE4D6ikc6_1(.din(w_dff_B_80W7Q4dK1_1),.dout(w_dff_B_kE4D6ikc6_1),.clk(gclk));
	jdff dff_B_NZR66vAv1_1(.din(w_dff_B_kE4D6ikc6_1),.dout(w_dff_B_NZR66vAv1_1),.clk(gclk));
	jdff dff_B_i7grhFx50_1(.din(w_dff_B_NZR66vAv1_1),.dout(w_dff_B_i7grhFx50_1),.clk(gclk));
	jdff dff_B_41zHWW3w6_1(.din(w_dff_B_i7grhFx50_1),.dout(w_dff_B_41zHWW3w6_1),.clk(gclk));
	jdff dff_B_7bi29k8c5_1(.din(w_dff_B_41zHWW3w6_1),.dout(w_dff_B_7bi29k8c5_1),.clk(gclk));
	jdff dff_B_LpPMhu5y7_1(.din(w_dff_B_7bi29k8c5_1),.dout(w_dff_B_LpPMhu5y7_1),.clk(gclk));
	jdff dff_B_0zcTE1Bs3_1(.din(w_dff_B_LpPMhu5y7_1),.dout(w_dff_B_0zcTE1Bs3_1),.clk(gclk));
	jdff dff_B_0qLLWQmH0_1(.din(w_dff_B_0zcTE1Bs3_1),.dout(w_dff_B_0qLLWQmH0_1),.clk(gclk));
	jdff dff_B_kSOBHOgB4_1(.din(w_dff_B_0qLLWQmH0_1),.dout(w_dff_B_kSOBHOgB4_1),.clk(gclk));
	jdff dff_B_GejgVfJ74_1(.din(w_dff_B_kSOBHOgB4_1),.dout(w_dff_B_GejgVfJ74_1),.clk(gclk));
	jdff dff_B_Jl2NPXL00_1(.din(w_dff_B_GejgVfJ74_1),.dout(w_dff_B_Jl2NPXL00_1),.clk(gclk));
	jdff dff_B_2lcY77pa2_1(.din(w_dff_B_Jl2NPXL00_1),.dout(w_dff_B_2lcY77pa2_1),.clk(gclk));
	jdff dff_B_8L5gM2XY0_1(.din(w_dff_B_2lcY77pa2_1),.dout(w_dff_B_8L5gM2XY0_1),.clk(gclk));
	jdff dff_B_3ktVkiK66_1(.din(w_dff_B_8L5gM2XY0_1),.dout(w_dff_B_3ktVkiK66_1),.clk(gclk));
	jdff dff_B_a3npL29q4_1(.din(w_dff_B_3ktVkiK66_1),.dout(w_dff_B_a3npL29q4_1),.clk(gclk));
	jdff dff_B_IWrQNUuz6_1(.din(w_dff_B_a3npL29q4_1),.dout(w_dff_B_IWrQNUuz6_1),.clk(gclk));
	jdff dff_B_aZkSvajn3_1(.din(w_dff_B_IWrQNUuz6_1),.dout(w_dff_B_aZkSvajn3_1),.clk(gclk));
	jdff dff_B_l8u35DY66_1(.din(w_dff_B_aZkSvajn3_1),.dout(w_dff_B_l8u35DY66_1),.clk(gclk));
	jdff dff_B_8igXaLMG6_1(.din(w_dff_B_l8u35DY66_1),.dout(w_dff_B_8igXaLMG6_1),.clk(gclk));
	jdff dff_B_JrGG7lIa6_1(.din(w_dff_B_8igXaLMG6_1),.dout(w_dff_B_JrGG7lIa6_1),.clk(gclk));
	jdff dff_B_JnJbw1BE6_1(.din(w_dff_B_JrGG7lIa6_1),.dout(w_dff_B_JnJbw1BE6_1),.clk(gclk));
	jdff dff_B_ZOZbBxey3_1(.din(w_dff_B_JnJbw1BE6_1),.dout(w_dff_B_ZOZbBxey3_1),.clk(gclk));
	jdff dff_B_jXTzPP9m4_1(.din(w_dff_B_ZOZbBxey3_1),.dout(w_dff_B_jXTzPP9m4_1),.clk(gclk));
	jdff dff_B_NoabEJFQ3_1(.din(w_dff_B_jXTzPP9m4_1),.dout(w_dff_B_NoabEJFQ3_1),.clk(gclk));
	jdff dff_B_LoQRTAu85_1(.din(w_dff_B_NoabEJFQ3_1),.dout(w_dff_B_LoQRTAu85_1),.clk(gclk));
	jdff dff_B_btPsXjUD0_1(.din(w_dff_B_LoQRTAu85_1),.dout(w_dff_B_btPsXjUD0_1),.clk(gclk));
	jdff dff_B_NQmElksK9_1(.din(w_dff_B_btPsXjUD0_1),.dout(w_dff_B_NQmElksK9_1),.clk(gclk));
	jdff dff_B_Gv8tLM9X0_1(.din(w_dff_B_NQmElksK9_1),.dout(w_dff_B_Gv8tLM9X0_1),.clk(gclk));
	jdff dff_B_3omyXlQ26_1(.din(w_dff_B_Gv8tLM9X0_1),.dout(w_dff_B_3omyXlQ26_1),.clk(gclk));
	jdff dff_B_LnUCF9vy8_1(.din(w_dff_B_3omyXlQ26_1),.dout(w_dff_B_LnUCF9vy8_1),.clk(gclk));
	jdff dff_B_yBmv7bjw0_1(.din(w_dff_B_LnUCF9vy8_1),.dout(w_dff_B_yBmv7bjw0_1),.clk(gclk));
	jdff dff_B_RAHituV56_0(.din(n823),.dout(w_dff_B_RAHituV56_0),.clk(gclk));
	jdff dff_B_aA9MMUZg1_0(.din(w_dff_B_RAHituV56_0),.dout(w_dff_B_aA9MMUZg1_0),.clk(gclk));
	jdff dff_B_MiQYWdBZ7_0(.din(w_dff_B_aA9MMUZg1_0),.dout(w_dff_B_MiQYWdBZ7_0),.clk(gclk));
	jdff dff_B_ZEsAe6eD3_0(.din(w_dff_B_MiQYWdBZ7_0),.dout(w_dff_B_ZEsAe6eD3_0),.clk(gclk));
	jdff dff_B_i6VhmQwu4_0(.din(w_dff_B_ZEsAe6eD3_0),.dout(w_dff_B_i6VhmQwu4_0),.clk(gclk));
	jdff dff_B_L3ynKQpL0_0(.din(w_dff_B_i6VhmQwu4_0),.dout(w_dff_B_L3ynKQpL0_0),.clk(gclk));
	jdff dff_B_S3mZmyAG0_0(.din(w_dff_B_L3ynKQpL0_0),.dout(w_dff_B_S3mZmyAG0_0),.clk(gclk));
	jdff dff_B_ZYTmjL1Y3_0(.din(w_dff_B_S3mZmyAG0_0),.dout(w_dff_B_ZYTmjL1Y3_0),.clk(gclk));
	jdff dff_B_VOoMSUSD9_0(.din(w_dff_B_ZYTmjL1Y3_0),.dout(w_dff_B_VOoMSUSD9_0),.clk(gclk));
	jdff dff_B_zFqCZzvi4_0(.din(w_dff_B_VOoMSUSD9_0),.dout(w_dff_B_zFqCZzvi4_0),.clk(gclk));
	jdff dff_B_uSlPX1qB3_0(.din(w_dff_B_zFqCZzvi4_0),.dout(w_dff_B_uSlPX1qB3_0),.clk(gclk));
	jdff dff_B_VlSZki5Q5_0(.din(w_dff_B_uSlPX1qB3_0),.dout(w_dff_B_VlSZki5Q5_0),.clk(gclk));
	jdff dff_B_6IxXXMo99_0(.din(w_dff_B_VlSZki5Q5_0),.dout(w_dff_B_6IxXXMo99_0),.clk(gclk));
	jdff dff_B_tS0SPITA0_0(.din(w_dff_B_6IxXXMo99_0),.dout(w_dff_B_tS0SPITA0_0),.clk(gclk));
	jdff dff_B_dLKL2beP3_0(.din(w_dff_B_tS0SPITA0_0),.dout(w_dff_B_dLKL2beP3_0),.clk(gclk));
	jdff dff_B_0GqKqaxd3_0(.din(w_dff_B_dLKL2beP3_0),.dout(w_dff_B_0GqKqaxd3_0),.clk(gclk));
	jdff dff_B_x9E4GK9J7_0(.din(w_dff_B_0GqKqaxd3_0),.dout(w_dff_B_x9E4GK9J7_0),.clk(gclk));
	jdff dff_B_H8rbAbgZ0_0(.din(w_dff_B_x9E4GK9J7_0),.dout(w_dff_B_H8rbAbgZ0_0),.clk(gclk));
	jdff dff_B_eAxQyGb48_0(.din(w_dff_B_H8rbAbgZ0_0),.dout(w_dff_B_eAxQyGb48_0),.clk(gclk));
	jdff dff_B_DOSvCxMA8_0(.din(w_dff_B_eAxQyGb48_0),.dout(w_dff_B_DOSvCxMA8_0),.clk(gclk));
	jdff dff_B_nZ7TMs2t3_0(.din(w_dff_B_DOSvCxMA8_0),.dout(w_dff_B_nZ7TMs2t3_0),.clk(gclk));
	jdff dff_B_Q4jb6NL63_0(.din(w_dff_B_nZ7TMs2t3_0),.dout(w_dff_B_Q4jb6NL63_0),.clk(gclk));
	jdff dff_B_Rrqr1Uj90_0(.din(w_dff_B_Q4jb6NL63_0),.dout(w_dff_B_Rrqr1Uj90_0),.clk(gclk));
	jdff dff_B_mfjnUpzA1_0(.din(w_dff_B_Rrqr1Uj90_0),.dout(w_dff_B_mfjnUpzA1_0),.clk(gclk));
	jdff dff_B_jRAkfUvh2_0(.din(w_dff_B_mfjnUpzA1_0),.dout(w_dff_B_jRAkfUvh2_0),.clk(gclk));
	jdff dff_B_OZJFt1Jz9_0(.din(w_dff_B_jRAkfUvh2_0),.dout(w_dff_B_OZJFt1Jz9_0),.clk(gclk));
	jdff dff_B_oYk5U38s2_0(.din(w_dff_B_OZJFt1Jz9_0),.dout(w_dff_B_oYk5U38s2_0),.clk(gclk));
	jdff dff_B_HWRZgDLW4_0(.din(w_dff_B_oYk5U38s2_0),.dout(w_dff_B_HWRZgDLW4_0),.clk(gclk));
	jdff dff_B_MlqYv43V0_0(.din(w_dff_B_HWRZgDLW4_0),.dout(w_dff_B_MlqYv43V0_0),.clk(gclk));
	jdff dff_B_5ej493qt9_0(.din(w_dff_B_MlqYv43V0_0),.dout(w_dff_B_5ej493qt9_0),.clk(gclk));
	jdff dff_B_NqJiMSj51_0(.din(w_dff_B_5ej493qt9_0),.dout(w_dff_B_NqJiMSj51_0),.clk(gclk));
	jdff dff_B_87PaAeXd0_0(.din(w_dff_B_NqJiMSj51_0),.dout(w_dff_B_87PaAeXd0_0),.clk(gclk));
	jdff dff_B_pruRAMB99_0(.din(w_dff_B_87PaAeXd0_0),.dout(w_dff_B_pruRAMB99_0),.clk(gclk));
	jdff dff_B_1MNEhZdI5_0(.din(w_dff_B_pruRAMB99_0),.dout(w_dff_B_1MNEhZdI5_0),.clk(gclk));
	jdff dff_B_IpnBBlcW6_0(.din(w_dff_B_1MNEhZdI5_0),.dout(w_dff_B_IpnBBlcW6_0),.clk(gclk));
	jdff dff_B_hiA6z7NU1_0(.din(w_dff_B_IpnBBlcW6_0),.dout(w_dff_B_hiA6z7NU1_0),.clk(gclk));
	jdff dff_B_QzJp9Tl70_0(.din(w_dff_B_hiA6z7NU1_0),.dout(w_dff_B_QzJp9Tl70_0),.clk(gclk));
	jdff dff_B_7O96u6dz3_0(.din(w_dff_B_QzJp9Tl70_0),.dout(w_dff_B_7O96u6dz3_0),.clk(gclk));
	jdff dff_B_6dwmHMj61_0(.din(w_dff_B_7O96u6dz3_0),.dout(w_dff_B_6dwmHMj61_0),.clk(gclk));
	jdff dff_B_lsEPhBgi2_0(.din(w_dff_B_6dwmHMj61_0),.dout(w_dff_B_lsEPhBgi2_0),.clk(gclk));
	jdff dff_B_0qBd94Ap8_0(.din(w_dff_B_lsEPhBgi2_0),.dout(w_dff_B_0qBd94Ap8_0),.clk(gclk));
	jdff dff_B_fEVehGMh4_0(.din(w_dff_B_0qBd94Ap8_0),.dout(w_dff_B_fEVehGMh4_0),.clk(gclk));
	jdff dff_B_DSndmckA4_0(.din(w_dff_B_fEVehGMh4_0),.dout(w_dff_B_DSndmckA4_0),.clk(gclk));
	jdff dff_B_2ogHnr3U7_0(.din(w_dff_B_DSndmckA4_0),.dout(w_dff_B_2ogHnr3U7_0),.clk(gclk));
	jdff dff_B_qrPuhFOX2_0(.din(w_dff_B_2ogHnr3U7_0),.dout(w_dff_B_qrPuhFOX2_0),.clk(gclk));
	jdff dff_B_su8gd8sq2_0(.din(w_dff_B_qrPuhFOX2_0),.dout(w_dff_B_su8gd8sq2_0),.clk(gclk));
	jdff dff_B_KbhraIE22_0(.din(w_dff_B_su8gd8sq2_0),.dout(w_dff_B_KbhraIE22_0),.clk(gclk));
	jdff dff_B_iKk4QUEi2_0(.din(w_dff_B_KbhraIE22_0),.dout(w_dff_B_iKk4QUEi2_0),.clk(gclk));
	jdff dff_B_zyjU2V6i8_0(.din(w_dff_B_iKk4QUEi2_0),.dout(w_dff_B_zyjU2V6i8_0),.clk(gclk));
	jdff dff_B_dlmvgXlg2_0(.din(w_dff_B_zyjU2V6i8_0),.dout(w_dff_B_dlmvgXlg2_0),.clk(gclk));
	jdff dff_B_VNb5ncHS1_0(.din(w_dff_B_dlmvgXlg2_0),.dout(w_dff_B_VNb5ncHS1_0),.clk(gclk));
	jdff dff_B_KfjkTy7X0_0(.din(w_dff_B_VNb5ncHS1_0),.dout(w_dff_B_KfjkTy7X0_0),.clk(gclk));
	jdff dff_B_Bb9Mwo246_0(.din(w_dff_B_KfjkTy7X0_0),.dout(w_dff_B_Bb9Mwo246_0),.clk(gclk));
	jdff dff_B_YnB2EQJc4_0(.din(w_dff_B_Bb9Mwo246_0),.dout(w_dff_B_YnB2EQJc4_0),.clk(gclk));
	jdff dff_B_qpnWWWUU5_0(.din(w_dff_B_YnB2EQJc4_0),.dout(w_dff_B_qpnWWWUU5_0),.clk(gclk));
	jdff dff_B_FgWrSpTH5_0(.din(w_dff_B_qpnWWWUU5_0),.dout(w_dff_B_FgWrSpTH5_0),.clk(gclk));
	jdff dff_B_BYDiHvZm4_0(.din(w_dff_B_FgWrSpTH5_0),.dout(w_dff_B_BYDiHvZm4_0),.clk(gclk));
	jdff dff_B_Do5MkOoQ6_0(.din(w_dff_B_BYDiHvZm4_0),.dout(w_dff_B_Do5MkOoQ6_0),.clk(gclk));
	jdff dff_B_yrz9v0t61_0(.din(w_dff_B_Do5MkOoQ6_0),.dout(w_dff_B_yrz9v0t61_0),.clk(gclk));
	jdff dff_B_5z3U7XQD0_0(.din(w_dff_B_yrz9v0t61_0),.dout(w_dff_B_5z3U7XQD0_0),.clk(gclk));
	jdff dff_B_3XnMhdo41_0(.din(w_dff_B_5z3U7XQD0_0),.dout(w_dff_B_3XnMhdo41_0),.clk(gclk));
	jdff dff_B_eBPAsBAR6_0(.din(w_dff_B_3XnMhdo41_0),.dout(w_dff_B_eBPAsBAR6_0),.clk(gclk));
	jdff dff_B_IZUlk9BH6_0(.din(w_dff_B_eBPAsBAR6_0),.dout(w_dff_B_IZUlk9BH6_0),.clk(gclk));
	jdff dff_B_dxMJb1gP3_0(.din(w_dff_B_IZUlk9BH6_0),.dout(w_dff_B_dxMJb1gP3_0),.clk(gclk));
	jdff dff_B_vPvwatj83_0(.din(w_dff_B_dxMJb1gP3_0),.dout(w_dff_B_vPvwatj83_0),.clk(gclk));
	jdff dff_B_wRo5T9ko6_0(.din(w_dff_B_vPvwatj83_0),.dout(w_dff_B_wRo5T9ko6_0),.clk(gclk));
	jdff dff_B_Zc2pNYTa5_0(.din(w_dff_B_wRo5T9ko6_0),.dout(w_dff_B_Zc2pNYTa5_0),.clk(gclk));
	jdff dff_B_lpghyYVv7_0(.din(w_dff_B_Zc2pNYTa5_0),.dout(w_dff_B_lpghyYVv7_0),.clk(gclk));
	jdff dff_B_2Hi23M2r2_0(.din(w_dff_B_lpghyYVv7_0),.dout(w_dff_B_2Hi23M2r2_0),.clk(gclk));
	jdff dff_B_PZz4M9hI3_0(.din(w_dff_B_2Hi23M2r2_0),.dout(w_dff_B_PZz4M9hI3_0),.clk(gclk));
	jdff dff_B_Y9Cdh24Z6_0(.din(w_dff_B_PZz4M9hI3_0),.dout(w_dff_B_Y9Cdh24Z6_0),.clk(gclk));
	jdff dff_B_BODBuvVB6_0(.din(w_dff_B_Y9Cdh24Z6_0),.dout(w_dff_B_BODBuvVB6_0),.clk(gclk));
	jdff dff_B_rKut0M2W1_0(.din(w_dff_B_BODBuvVB6_0),.dout(w_dff_B_rKut0M2W1_0),.clk(gclk));
	jdff dff_B_b4HSidhS9_1(.din(n816),.dout(w_dff_B_b4HSidhS9_1),.clk(gclk));
	jdff dff_B_GrqHro6J9_1(.din(w_dff_B_b4HSidhS9_1),.dout(w_dff_B_GrqHro6J9_1),.clk(gclk));
	jdff dff_B_QwqtT17P6_1(.din(w_dff_B_GrqHro6J9_1),.dout(w_dff_B_QwqtT17P6_1),.clk(gclk));
	jdff dff_B_SvqzD8iR4_1(.din(w_dff_B_QwqtT17P6_1),.dout(w_dff_B_SvqzD8iR4_1),.clk(gclk));
	jdff dff_B_5N730P6n1_1(.din(w_dff_B_SvqzD8iR4_1),.dout(w_dff_B_5N730P6n1_1),.clk(gclk));
	jdff dff_B_PN4JjQXV6_1(.din(w_dff_B_5N730P6n1_1),.dout(w_dff_B_PN4JjQXV6_1),.clk(gclk));
	jdff dff_B_xvcyzseX9_1(.din(w_dff_B_PN4JjQXV6_1),.dout(w_dff_B_xvcyzseX9_1),.clk(gclk));
	jdff dff_B_SmHblLy75_1(.din(w_dff_B_xvcyzseX9_1),.dout(w_dff_B_SmHblLy75_1),.clk(gclk));
	jdff dff_B_T5smbZTS3_1(.din(w_dff_B_SmHblLy75_1),.dout(w_dff_B_T5smbZTS3_1),.clk(gclk));
	jdff dff_B_GACa4STw2_1(.din(w_dff_B_T5smbZTS3_1),.dout(w_dff_B_GACa4STw2_1),.clk(gclk));
	jdff dff_B_M4lhjITy5_1(.din(w_dff_B_GACa4STw2_1),.dout(w_dff_B_M4lhjITy5_1),.clk(gclk));
	jdff dff_B_PRzfMe5g1_1(.din(w_dff_B_M4lhjITy5_1),.dout(w_dff_B_PRzfMe5g1_1),.clk(gclk));
	jdff dff_B_5OcTVZmz6_1(.din(w_dff_B_PRzfMe5g1_1),.dout(w_dff_B_5OcTVZmz6_1),.clk(gclk));
	jdff dff_B_1g5NA4Bn0_1(.din(w_dff_B_5OcTVZmz6_1),.dout(w_dff_B_1g5NA4Bn0_1),.clk(gclk));
	jdff dff_B_AtgLpfYf0_1(.din(w_dff_B_1g5NA4Bn0_1),.dout(w_dff_B_AtgLpfYf0_1),.clk(gclk));
	jdff dff_B_pl2Jfj7l2_1(.din(w_dff_B_AtgLpfYf0_1),.dout(w_dff_B_pl2Jfj7l2_1),.clk(gclk));
	jdff dff_B_l2TMvDHP2_1(.din(w_dff_B_pl2Jfj7l2_1),.dout(w_dff_B_l2TMvDHP2_1),.clk(gclk));
	jdff dff_B_6MYnmPOk8_1(.din(w_dff_B_l2TMvDHP2_1),.dout(w_dff_B_6MYnmPOk8_1),.clk(gclk));
	jdff dff_B_7up5ZRKX0_1(.din(w_dff_B_6MYnmPOk8_1),.dout(w_dff_B_7up5ZRKX0_1),.clk(gclk));
	jdff dff_B_WkErKG0L6_1(.din(w_dff_B_7up5ZRKX0_1),.dout(w_dff_B_WkErKG0L6_1),.clk(gclk));
	jdff dff_B_mun8BVp62_1(.din(w_dff_B_WkErKG0L6_1),.dout(w_dff_B_mun8BVp62_1),.clk(gclk));
	jdff dff_B_epqHRWpi1_1(.din(w_dff_B_mun8BVp62_1),.dout(w_dff_B_epqHRWpi1_1),.clk(gclk));
	jdff dff_B_Oy2Vne6r4_1(.din(w_dff_B_epqHRWpi1_1),.dout(w_dff_B_Oy2Vne6r4_1),.clk(gclk));
	jdff dff_B_2Y9W4CfV7_1(.din(w_dff_B_Oy2Vne6r4_1),.dout(w_dff_B_2Y9W4CfV7_1),.clk(gclk));
	jdff dff_B_NNLff3Lt3_1(.din(w_dff_B_2Y9W4CfV7_1),.dout(w_dff_B_NNLff3Lt3_1),.clk(gclk));
	jdff dff_B_K686eWDB7_1(.din(w_dff_B_NNLff3Lt3_1),.dout(w_dff_B_K686eWDB7_1),.clk(gclk));
	jdff dff_B_r7aCH8wM3_1(.din(w_dff_B_K686eWDB7_1),.dout(w_dff_B_r7aCH8wM3_1),.clk(gclk));
	jdff dff_B_zSS8ZzN40_1(.din(w_dff_B_r7aCH8wM3_1),.dout(w_dff_B_zSS8ZzN40_1),.clk(gclk));
	jdff dff_B_9LHZBG0E0_1(.din(w_dff_B_zSS8ZzN40_1),.dout(w_dff_B_9LHZBG0E0_1),.clk(gclk));
	jdff dff_B_xk1N7SbQ3_1(.din(w_dff_B_9LHZBG0E0_1),.dout(w_dff_B_xk1N7SbQ3_1),.clk(gclk));
	jdff dff_B_tcFwzUeZ0_1(.din(w_dff_B_xk1N7SbQ3_1),.dout(w_dff_B_tcFwzUeZ0_1),.clk(gclk));
	jdff dff_B_cJsWbnMT9_1(.din(w_dff_B_tcFwzUeZ0_1),.dout(w_dff_B_cJsWbnMT9_1),.clk(gclk));
	jdff dff_B_cpxgLhzs4_1(.din(w_dff_B_cJsWbnMT9_1),.dout(w_dff_B_cpxgLhzs4_1),.clk(gclk));
	jdff dff_B_PNSolVS35_1(.din(w_dff_B_cpxgLhzs4_1),.dout(w_dff_B_PNSolVS35_1),.clk(gclk));
	jdff dff_B_KTV7JitT7_1(.din(w_dff_B_PNSolVS35_1),.dout(w_dff_B_KTV7JitT7_1),.clk(gclk));
	jdff dff_B_S5kF8oyp1_1(.din(w_dff_B_KTV7JitT7_1),.dout(w_dff_B_S5kF8oyp1_1),.clk(gclk));
	jdff dff_B_4eOrq1hD2_1(.din(w_dff_B_S5kF8oyp1_1),.dout(w_dff_B_4eOrq1hD2_1),.clk(gclk));
	jdff dff_B_jYEZptSz4_1(.din(w_dff_B_4eOrq1hD2_1),.dout(w_dff_B_jYEZptSz4_1),.clk(gclk));
	jdff dff_B_84AFV4wZ4_1(.din(w_dff_B_jYEZptSz4_1),.dout(w_dff_B_84AFV4wZ4_1),.clk(gclk));
	jdff dff_B_SbOqHVtP9_1(.din(w_dff_B_84AFV4wZ4_1),.dout(w_dff_B_SbOqHVtP9_1),.clk(gclk));
	jdff dff_B_PihnK1wM7_1(.din(w_dff_B_SbOqHVtP9_1),.dout(w_dff_B_PihnK1wM7_1),.clk(gclk));
	jdff dff_B_pC7Qi3dg8_1(.din(w_dff_B_PihnK1wM7_1),.dout(w_dff_B_pC7Qi3dg8_1),.clk(gclk));
	jdff dff_B_kFReKYZS6_1(.din(w_dff_B_pC7Qi3dg8_1),.dout(w_dff_B_kFReKYZS6_1),.clk(gclk));
	jdff dff_B_HgL6vTZ53_1(.din(w_dff_B_kFReKYZS6_1),.dout(w_dff_B_HgL6vTZ53_1),.clk(gclk));
	jdff dff_B_M6R53h0c2_1(.din(w_dff_B_HgL6vTZ53_1),.dout(w_dff_B_M6R53h0c2_1),.clk(gclk));
	jdff dff_B_jVlFUBsW6_1(.din(w_dff_B_M6R53h0c2_1),.dout(w_dff_B_jVlFUBsW6_1),.clk(gclk));
	jdff dff_B_o9X0LLj41_1(.din(w_dff_B_jVlFUBsW6_1),.dout(w_dff_B_o9X0LLj41_1),.clk(gclk));
	jdff dff_B_ydGaxygF9_1(.din(w_dff_B_o9X0LLj41_1),.dout(w_dff_B_ydGaxygF9_1),.clk(gclk));
	jdff dff_B_pvG1Bkes5_1(.din(w_dff_B_ydGaxygF9_1),.dout(w_dff_B_pvG1Bkes5_1),.clk(gclk));
	jdff dff_B_zJdmmRxx5_1(.din(w_dff_B_pvG1Bkes5_1),.dout(w_dff_B_zJdmmRxx5_1),.clk(gclk));
	jdff dff_B_hZMGqjXs4_1(.din(w_dff_B_zJdmmRxx5_1),.dout(w_dff_B_hZMGqjXs4_1),.clk(gclk));
	jdff dff_B_pM2AWCf15_1(.din(w_dff_B_hZMGqjXs4_1),.dout(w_dff_B_pM2AWCf15_1),.clk(gclk));
	jdff dff_B_BWm5S38Q9_1(.din(w_dff_B_pM2AWCf15_1),.dout(w_dff_B_BWm5S38Q9_1),.clk(gclk));
	jdff dff_B_pJmzltft3_1(.din(w_dff_B_BWm5S38Q9_1),.dout(w_dff_B_pJmzltft3_1),.clk(gclk));
	jdff dff_B_aH3rfv8h8_1(.din(w_dff_B_pJmzltft3_1),.dout(w_dff_B_aH3rfv8h8_1),.clk(gclk));
	jdff dff_B_TK7dTSFu2_1(.din(w_dff_B_aH3rfv8h8_1),.dout(w_dff_B_TK7dTSFu2_1),.clk(gclk));
	jdff dff_B_apqCesxp5_1(.din(w_dff_B_TK7dTSFu2_1),.dout(w_dff_B_apqCesxp5_1),.clk(gclk));
	jdff dff_B_fTtlmO4F2_1(.din(w_dff_B_apqCesxp5_1),.dout(w_dff_B_fTtlmO4F2_1),.clk(gclk));
	jdff dff_B_9JdUVkl86_1(.din(w_dff_B_fTtlmO4F2_1),.dout(w_dff_B_9JdUVkl86_1),.clk(gclk));
	jdff dff_B_gfWeo0Ef7_1(.din(w_dff_B_9JdUVkl86_1),.dout(w_dff_B_gfWeo0Ef7_1),.clk(gclk));
	jdff dff_B_B2rUbfEZ7_1(.din(w_dff_B_gfWeo0Ef7_1),.dout(w_dff_B_B2rUbfEZ7_1),.clk(gclk));
	jdff dff_B_A6hKXfm65_1(.din(w_dff_B_B2rUbfEZ7_1),.dout(w_dff_B_A6hKXfm65_1),.clk(gclk));
	jdff dff_B_rgd4q4JO6_1(.din(w_dff_B_A6hKXfm65_1),.dout(w_dff_B_rgd4q4JO6_1),.clk(gclk));
	jdff dff_B_qTTQQUpr0_1(.din(w_dff_B_rgd4q4JO6_1),.dout(w_dff_B_qTTQQUpr0_1),.clk(gclk));
	jdff dff_B_ATxwmUt31_1(.din(w_dff_B_qTTQQUpr0_1),.dout(w_dff_B_ATxwmUt31_1),.clk(gclk));
	jdff dff_B_HaKLKpFt1_1(.din(w_dff_B_ATxwmUt31_1),.dout(w_dff_B_HaKLKpFt1_1),.clk(gclk));
	jdff dff_B_GYiACixA2_1(.din(w_dff_B_HaKLKpFt1_1),.dout(w_dff_B_GYiACixA2_1),.clk(gclk));
	jdff dff_B_O8vQytY30_1(.din(w_dff_B_GYiACixA2_1),.dout(w_dff_B_O8vQytY30_1),.clk(gclk));
	jdff dff_B_qARWhyZh9_1(.din(w_dff_B_O8vQytY30_1),.dout(w_dff_B_qARWhyZh9_1),.clk(gclk));
	jdff dff_B_XT4w1tQi0_1(.din(w_dff_B_qARWhyZh9_1),.dout(w_dff_B_XT4w1tQi0_1),.clk(gclk));
	jdff dff_B_nAL383XY7_1(.din(w_dff_B_XT4w1tQi0_1),.dout(w_dff_B_nAL383XY7_1),.clk(gclk));
	jdff dff_B_CmLHlizM1_1(.din(w_dff_B_nAL383XY7_1),.dout(w_dff_B_CmLHlizM1_1),.clk(gclk));
	jdff dff_B_GFyTLlSL7_0(.din(n817),.dout(w_dff_B_GFyTLlSL7_0),.clk(gclk));
	jdff dff_B_PxTmtekB1_0(.din(w_dff_B_GFyTLlSL7_0),.dout(w_dff_B_PxTmtekB1_0),.clk(gclk));
	jdff dff_B_QHM1ATau8_0(.din(w_dff_B_PxTmtekB1_0),.dout(w_dff_B_QHM1ATau8_0),.clk(gclk));
	jdff dff_B_dRDueS452_0(.din(w_dff_B_QHM1ATau8_0),.dout(w_dff_B_dRDueS452_0),.clk(gclk));
	jdff dff_B_AH6aannt7_0(.din(w_dff_B_dRDueS452_0),.dout(w_dff_B_AH6aannt7_0),.clk(gclk));
	jdff dff_B_3rV3KiuU9_0(.din(w_dff_B_AH6aannt7_0),.dout(w_dff_B_3rV3KiuU9_0),.clk(gclk));
	jdff dff_B_9YAuWKnM3_0(.din(w_dff_B_3rV3KiuU9_0),.dout(w_dff_B_9YAuWKnM3_0),.clk(gclk));
	jdff dff_B_ssRh6omy8_0(.din(w_dff_B_9YAuWKnM3_0),.dout(w_dff_B_ssRh6omy8_0),.clk(gclk));
	jdff dff_B_B8JeIfJd8_0(.din(w_dff_B_ssRh6omy8_0),.dout(w_dff_B_B8JeIfJd8_0),.clk(gclk));
	jdff dff_B_cjHgWY2H3_0(.din(w_dff_B_B8JeIfJd8_0),.dout(w_dff_B_cjHgWY2H3_0),.clk(gclk));
	jdff dff_B_ywvVU7Mf4_0(.din(w_dff_B_cjHgWY2H3_0),.dout(w_dff_B_ywvVU7Mf4_0),.clk(gclk));
	jdff dff_B_BwVmR7SR8_0(.din(w_dff_B_ywvVU7Mf4_0),.dout(w_dff_B_BwVmR7SR8_0),.clk(gclk));
	jdff dff_B_nfUXkAuU9_0(.din(w_dff_B_BwVmR7SR8_0),.dout(w_dff_B_nfUXkAuU9_0),.clk(gclk));
	jdff dff_B_NQ3hdSku8_0(.din(w_dff_B_nfUXkAuU9_0),.dout(w_dff_B_NQ3hdSku8_0),.clk(gclk));
	jdff dff_B_DBcCHZp04_0(.din(w_dff_B_NQ3hdSku8_0),.dout(w_dff_B_DBcCHZp04_0),.clk(gclk));
	jdff dff_B_n4cvWEd38_0(.din(w_dff_B_DBcCHZp04_0),.dout(w_dff_B_n4cvWEd38_0),.clk(gclk));
	jdff dff_B_b02EVVu31_0(.din(w_dff_B_n4cvWEd38_0),.dout(w_dff_B_b02EVVu31_0),.clk(gclk));
	jdff dff_B_tmeqqpIg0_0(.din(w_dff_B_b02EVVu31_0),.dout(w_dff_B_tmeqqpIg0_0),.clk(gclk));
	jdff dff_B_aaBQF0Cn8_0(.din(w_dff_B_tmeqqpIg0_0),.dout(w_dff_B_aaBQF0Cn8_0),.clk(gclk));
	jdff dff_B_Fk1cmqpc9_0(.din(w_dff_B_aaBQF0Cn8_0),.dout(w_dff_B_Fk1cmqpc9_0),.clk(gclk));
	jdff dff_B_jAcp4NRB0_0(.din(w_dff_B_Fk1cmqpc9_0),.dout(w_dff_B_jAcp4NRB0_0),.clk(gclk));
	jdff dff_B_z424nFrH6_0(.din(w_dff_B_jAcp4NRB0_0),.dout(w_dff_B_z424nFrH6_0),.clk(gclk));
	jdff dff_B_5gWowZOH2_0(.din(w_dff_B_z424nFrH6_0),.dout(w_dff_B_5gWowZOH2_0),.clk(gclk));
	jdff dff_B_5n6abP317_0(.din(w_dff_B_5gWowZOH2_0),.dout(w_dff_B_5n6abP317_0),.clk(gclk));
	jdff dff_B_4AL1rcrm0_0(.din(w_dff_B_5n6abP317_0),.dout(w_dff_B_4AL1rcrm0_0),.clk(gclk));
	jdff dff_B_NxJ7c8hl3_0(.din(w_dff_B_4AL1rcrm0_0),.dout(w_dff_B_NxJ7c8hl3_0),.clk(gclk));
	jdff dff_B_YUV4qxrB6_0(.din(w_dff_B_NxJ7c8hl3_0),.dout(w_dff_B_YUV4qxrB6_0),.clk(gclk));
	jdff dff_B_WBcw1FaZ6_0(.din(w_dff_B_YUV4qxrB6_0),.dout(w_dff_B_WBcw1FaZ6_0),.clk(gclk));
	jdff dff_B_Y40OrlF30_0(.din(w_dff_B_WBcw1FaZ6_0),.dout(w_dff_B_Y40OrlF30_0),.clk(gclk));
	jdff dff_B_n08nwpdU0_0(.din(w_dff_B_Y40OrlF30_0),.dout(w_dff_B_n08nwpdU0_0),.clk(gclk));
	jdff dff_B_zVLiVMKA8_0(.din(w_dff_B_n08nwpdU0_0),.dout(w_dff_B_zVLiVMKA8_0),.clk(gclk));
	jdff dff_B_ddsPfdrH4_0(.din(w_dff_B_zVLiVMKA8_0),.dout(w_dff_B_ddsPfdrH4_0),.clk(gclk));
	jdff dff_B_nK1cSWgf8_0(.din(w_dff_B_ddsPfdrH4_0),.dout(w_dff_B_nK1cSWgf8_0),.clk(gclk));
	jdff dff_B_zhO5B4ZN8_0(.din(w_dff_B_nK1cSWgf8_0),.dout(w_dff_B_zhO5B4ZN8_0),.clk(gclk));
	jdff dff_B_GLenQ7nM6_0(.din(w_dff_B_zhO5B4ZN8_0),.dout(w_dff_B_GLenQ7nM6_0),.clk(gclk));
	jdff dff_B_rURqX3Tj8_0(.din(w_dff_B_GLenQ7nM6_0),.dout(w_dff_B_rURqX3Tj8_0),.clk(gclk));
	jdff dff_B_DvVKpehl2_0(.din(w_dff_B_rURqX3Tj8_0),.dout(w_dff_B_DvVKpehl2_0),.clk(gclk));
	jdff dff_B_WVedm75X3_0(.din(w_dff_B_DvVKpehl2_0),.dout(w_dff_B_WVedm75X3_0),.clk(gclk));
	jdff dff_B_zkc0RCJ48_0(.din(w_dff_B_WVedm75X3_0),.dout(w_dff_B_zkc0RCJ48_0),.clk(gclk));
	jdff dff_B_etj6C3jq1_0(.din(w_dff_B_zkc0RCJ48_0),.dout(w_dff_B_etj6C3jq1_0),.clk(gclk));
	jdff dff_B_pow9Xqhp8_0(.din(w_dff_B_etj6C3jq1_0),.dout(w_dff_B_pow9Xqhp8_0),.clk(gclk));
	jdff dff_B_IM238BUL5_0(.din(w_dff_B_pow9Xqhp8_0),.dout(w_dff_B_IM238BUL5_0),.clk(gclk));
	jdff dff_B_BvDFv2aE3_0(.din(w_dff_B_IM238BUL5_0),.dout(w_dff_B_BvDFv2aE3_0),.clk(gclk));
	jdff dff_B_goKe2PLj9_0(.din(w_dff_B_BvDFv2aE3_0),.dout(w_dff_B_goKe2PLj9_0),.clk(gclk));
	jdff dff_B_GtVZ4Owg1_0(.din(w_dff_B_goKe2PLj9_0),.dout(w_dff_B_GtVZ4Owg1_0),.clk(gclk));
	jdff dff_B_bB84obzN0_0(.din(w_dff_B_GtVZ4Owg1_0),.dout(w_dff_B_bB84obzN0_0),.clk(gclk));
	jdff dff_B_TVpGm1bL0_0(.din(w_dff_B_bB84obzN0_0),.dout(w_dff_B_TVpGm1bL0_0),.clk(gclk));
	jdff dff_B_iGMFxjY16_0(.din(w_dff_B_TVpGm1bL0_0),.dout(w_dff_B_iGMFxjY16_0),.clk(gclk));
	jdff dff_B_HftuvI6x5_0(.din(w_dff_B_iGMFxjY16_0),.dout(w_dff_B_HftuvI6x5_0),.clk(gclk));
	jdff dff_B_6KgP9fnU4_0(.din(w_dff_B_HftuvI6x5_0),.dout(w_dff_B_6KgP9fnU4_0),.clk(gclk));
	jdff dff_B_n1c7whd10_0(.din(w_dff_B_6KgP9fnU4_0),.dout(w_dff_B_n1c7whd10_0),.clk(gclk));
	jdff dff_B_utgJJrcv4_0(.din(w_dff_B_n1c7whd10_0),.dout(w_dff_B_utgJJrcv4_0),.clk(gclk));
	jdff dff_B_pSIxGsn99_0(.din(w_dff_B_utgJJrcv4_0),.dout(w_dff_B_pSIxGsn99_0),.clk(gclk));
	jdff dff_B_ZbWtIy7L5_0(.din(w_dff_B_pSIxGsn99_0),.dout(w_dff_B_ZbWtIy7L5_0),.clk(gclk));
	jdff dff_B_Z3Qc2kDf4_0(.din(w_dff_B_ZbWtIy7L5_0),.dout(w_dff_B_Z3Qc2kDf4_0),.clk(gclk));
	jdff dff_B_L1VMpWZE9_0(.din(w_dff_B_Z3Qc2kDf4_0),.dout(w_dff_B_L1VMpWZE9_0),.clk(gclk));
	jdff dff_B_sTh5CHzI9_0(.din(w_dff_B_L1VMpWZE9_0),.dout(w_dff_B_sTh5CHzI9_0),.clk(gclk));
	jdff dff_B_cf2HexZ64_0(.din(w_dff_B_sTh5CHzI9_0),.dout(w_dff_B_cf2HexZ64_0),.clk(gclk));
	jdff dff_B_qgPPnmKV3_0(.din(w_dff_B_cf2HexZ64_0),.dout(w_dff_B_qgPPnmKV3_0),.clk(gclk));
	jdff dff_B_JKcuVPDt2_0(.din(w_dff_B_qgPPnmKV3_0),.dout(w_dff_B_JKcuVPDt2_0),.clk(gclk));
	jdff dff_B_k51KdTd10_0(.din(w_dff_B_JKcuVPDt2_0),.dout(w_dff_B_k51KdTd10_0),.clk(gclk));
	jdff dff_B_mdfpRZoz6_0(.din(w_dff_B_k51KdTd10_0),.dout(w_dff_B_mdfpRZoz6_0),.clk(gclk));
	jdff dff_B_hwjwXKxG5_0(.din(w_dff_B_mdfpRZoz6_0),.dout(w_dff_B_hwjwXKxG5_0),.clk(gclk));
	jdff dff_B_duZOeWpI5_0(.din(w_dff_B_hwjwXKxG5_0),.dout(w_dff_B_duZOeWpI5_0),.clk(gclk));
	jdff dff_B_HAoUd2zw6_0(.din(w_dff_B_duZOeWpI5_0),.dout(w_dff_B_HAoUd2zw6_0),.clk(gclk));
	jdff dff_B_chVpCn8l2_0(.din(w_dff_B_HAoUd2zw6_0),.dout(w_dff_B_chVpCn8l2_0),.clk(gclk));
	jdff dff_B_KZNYSLRT7_0(.din(w_dff_B_chVpCn8l2_0),.dout(w_dff_B_KZNYSLRT7_0),.clk(gclk));
	jdff dff_B_vLichBWZ1_0(.din(w_dff_B_KZNYSLRT7_0),.dout(w_dff_B_vLichBWZ1_0),.clk(gclk));
	jdff dff_B_xgV7aKI32_0(.din(w_dff_B_vLichBWZ1_0),.dout(w_dff_B_xgV7aKI32_0),.clk(gclk));
	jdff dff_B_ukBXUbxV1_0(.din(w_dff_B_xgV7aKI32_0),.dout(w_dff_B_ukBXUbxV1_0),.clk(gclk));
	jdff dff_B_XnXEUs236_0(.din(w_dff_B_ukBXUbxV1_0),.dout(w_dff_B_XnXEUs236_0),.clk(gclk));
	jdff dff_B_FLEVHsvk5_0(.din(w_dff_B_XnXEUs236_0),.dout(w_dff_B_FLEVHsvk5_0),.clk(gclk));
	jdff dff_B_Fn07mpj66_1(.din(n810),.dout(w_dff_B_Fn07mpj66_1),.clk(gclk));
	jdff dff_B_CPMG4O5U9_1(.din(w_dff_B_Fn07mpj66_1),.dout(w_dff_B_CPMG4O5U9_1),.clk(gclk));
	jdff dff_B_SZoP2WA16_1(.din(w_dff_B_CPMG4O5U9_1),.dout(w_dff_B_SZoP2WA16_1),.clk(gclk));
	jdff dff_B_21kpJTjy4_1(.din(w_dff_B_SZoP2WA16_1),.dout(w_dff_B_21kpJTjy4_1),.clk(gclk));
	jdff dff_B_sREIaAun7_1(.din(w_dff_B_21kpJTjy4_1),.dout(w_dff_B_sREIaAun7_1),.clk(gclk));
	jdff dff_B_rHsmr3kF0_1(.din(w_dff_B_sREIaAun7_1),.dout(w_dff_B_rHsmr3kF0_1),.clk(gclk));
	jdff dff_B_iJqtsLo26_1(.din(w_dff_B_rHsmr3kF0_1),.dout(w_dff_B_iJqtsLo26_1),.clk(gclk));
	jdff dff_B_ofuibS3N9_1(.din(w_dff_B_iJqtsLo26_1),.dout(w_dff_B_ofuibS3N9_1),.clk(gclk));
	jdff dff_B_dWbTqyrF3_1(.din(w_dff_B_ofuibS3N9_1),.dout(w_dff_B_dWbTqyrF3_1),.clk(gclk));
	jdff dff_B_5ycJ3PHi8_1(.din(w_dff_B_dWbTqyrF3_1),.dout(w_dff_B_5ycJ3PHi8_1),.clk(gclk));
	jdff dff_B_23mOysOv2_1(.din(w_dff_B_5ycJ3PHi8_1),.dout(w_dff_B_23mOysOv2_1),.clk(gclk));
	jdff dff_B_wt0vfdau2_1(.din(w_dff_B_23mOysOv2_1),.dout(w_dff_B_wt0vfdau2_1),.clk(gclk));
	jdff dff_B_5Gfz4Cbu7_1(.din(w_dff_B_wt0vfdau2_1),.dout(w_dff_B_5Gfz4Cbu7_1),.clk(gclk));
	jdff dff_B_0z0OIQZK0_1(.din(w_dff_B_5Gfz4Cbu7_1),.dout(w_dff_B_0z0OIQZK0_1),.clk(gclk));
	jdff dff_B_Qucn0uoQ0_1(.din(w_dff_B_0z0OIQZK0_1),.dout(w_dff_B_Qucn0uoQ0_1),.clk(gclk));
	jdff dff_B_u2B7voVP8_1(.din(w_dff_B_Qucn0uoQ0_1),.dout(w_dff_B_u2B7voVP8_1),.clk(gclk));
	jdff dff_B_OsrTxzBq6_1(.din(w_dff_B_u2B7voVP8_1),.dout(w_dff_B_OsrTxzBq6_1),.clk(gclk));
	jdff dff_B_D08ZMa047_1(.din(w_dff_B_OsrTxzBq6_1),.dout(w_dff_B_D08ZMa047_1),.clk(gclk));
	jdff dff_B_evWj6xiq4_1(.din(w_dff_B_D08ZMa047_1),.dout(w_dff_B_evWj6xiq4_1),.clk(gclk));
	jdff dff_B_J40iZ6Ho9_1(.din(w_dff_B_evWj6xiq4_1),.dout(w_dff_B_J40iZ6Ho9_1),.clk(gclk));
	jdff dff_B_nWKsqVu08_1(.din(w_dff_B_J40iZ6Ho9_1),.dout(w_dff_B_nWKsqVu08_1),.clk(gclk));
	jdff dff_B_viNll7tx8_1(.din(w_dff_B_nWKsqVu08_1),.dout(w_dff_B_viNll7tx8_1),.clk(gclk));
	jdff dff_B_qGJVV4M45_1(.din(w_dff_B_viNll7tx8_1),.dout(w_dff_B_qGJVV4M45_1),.clk(gclk));
	jdff dff_B_HkIhst496_1(.din(w_dff_B_qGJVV4M45_1),.dout(w_dff_B_HkIhst496_1),.clk(gclk));
	jdff dff_B_VZq9cFdL7_1(.din(w_dff_B_HkIhst496_1),.dout(w_dff_B_VZq9cFdL7_1),.clk(gclk));
	jdff dff_B_ounaAOLQ4_1(.din(w_dff_B_VZq9cFdL7_1),.dout(w_dff_B_ounaAOLQ4_1),.clk(gclk));
	jdff dff_B_2duDj88d2_1(.din(w_dff_B_ounaAOLQ4_1),.dout(w_dff_B_2duDj88d2_1),.clk(gclk));
	jdff dff_B_XGy4m2J89_1(.din(w_dff_B_2duDj88d2_1),.dout(w_dff_B_XGy4m2J89_1),.clk(gclk));
	jdff dff_B_s29Eg6PN9_1(.din(w_dff_B_XGy4m2J89_1),.dout(w_dff_B_s29Eg6PN9_1),.clk(gclk));
	jdff dff_B_NmxiH5lS5_1(.din(w_dff_B_s29Eg6PN9_1),.dout(w_dff_B_NmxiH5lS5_1),.clk(gclk));
	jdff dff_B_nBGMMrt79_1(.din(w_dff_B_NmxiH5lS5_1),.dout(w_dff_B_nBGMMrt79_1),.clk(gclk));
	jdff dff_B_NjWXLlhu1_1(.din(w_dff_B_nBGMMrt79_1),.dout(w_dff_B_NjWXLlhu1_1),.clk(gclk));
	jdff dff_B_QJaX1yLt5_1(.din(w_dff_B_NjWXLlhu1_1),.dout(w_dff_B_QJaX1yLt5_1),.clk(gclk));
	jdff dff_B_1nZXS5tk2_1(.din(w_dff_B_QJaX1yLt5_1),.dout(w_dff_B_1nZXS5tk2_1),.clk(gclk));
	jdff dff_B_HgjxWLeM9_1(.din(w_dff_B_1nZXS5tk2_1),.dout(w_dff_B_HgjxWLeM9_1),.clk(gclk));
	jdff dff_B_QzBSIu435_1(.din(w_dff_B_HgjxWLeM9_1),.dout(w_dff_B_QzBSIu435_1),.clk(gclk));
	jdff dff_B_NBZzaYUS9_1(.din(w_dff_B_QzBSIu435_1),.dout(w_dff_B_NBZzaYUS9_1),.clk(gclk));
	jdff dff_B_GqbdVfgC8_1(.din(w_dff_B_NBZzaYUS9_1),.dout(w_dff_B_GqbdVfgC8_1),.clk(gclk));
	jdff dff_B_erHLbXQL4_1(.din(w_dff_B_GqbdVfgC8_1),.dout(w_dff_B_erHLbXQL4_1),.clk(gclk));
	jdff dff_B_eUUKJn3q6_1(.din(w_dff_B_erHLbXQL4_1),.dout(w_dff_B_eUUKJn3q6_1),.clk(gclk));
	jdff dff_B_H1ytEKT36_1(.din(w_dff_B_eUUKJn3q6_1),.dout(w_dff_B_H1ytEKT36_1),.clk(gclk));
	jdff dff_B_GGB3ALZY0_1(.din(w_dff_B_H1ytEKT36_1),.dout(w_dff_B_GGB3ALZY0_1),.clk(gclk));
	jdff dff_B_JAfcG5719_1(.din(w_dff_B_GGB3ALZY0_1),.dout(w_dff_B_JAfcG5719_1),.clk(gclk));
	jdff dff_B_Mxvq50P53_1(.din(w_dff_B_JAfcG5719_1),.dout(w_dff_B_Mxvq50P53_1),.clk(gclk));
	jdff dff_B_lVh7q02f0_1(.din(w_dff_B_Mxvq50P53_1),.dout(w_dff_B_lVh7q02f0_1),.clk(gclk));
	jdff dff_B_yJxWgjrK7_1(.din(w_dff_B_lVh7q02f0_1),.dout(w_dff_B_yJxWgjrK7_1),.clk(gclk));
	jdff dff_B_7bj5zypn6_1(.din(w_dff_B_yJxWgjrK7_1),.dout(w_dff_B_7bj5zypn6_1),.clk(gclk));
	jdff dff_B_bWnn7mRa7_1(.din(w_dff_B_7bj5zypn6_1),.dout(w_dff_B_bWnn7mRa7_1),.clk(gclk));
	jdff dff_B_YFgZ2xtI1_1(.din(w_dff_B_bWnn7mRa7_1),.dout(w_dff_B_YFgZ2xtI1_1),.clk(gclk));
	jdff dff_B_2q3ifhJd6_1(.din(w_dff_B_YFgZ2xtI1_1),.dout(w_dff_B_2q3ifhJd6_1),.clk(gclk));
	jdff dff_B_br2dRU665_1(.din(w_dff_B_2q3ifhJd6_1),.dout(w_dff_B_br2dRU665_1),.clk(gclk));
	jdff dff_B_jcF9v2hz5_1(.din(w_dff_B_br2dRU665_1),.dout(w_dff_B_jcF9v2hz5_1),.clk(gclk));
	jdff dff_B_mNc6PFXQ0_1(.din(w_dff_B_jcF9v2hz5_1),.dout(w_dff_B_mNc6PFXQ0_1),.clk(gclk));
	jdff dff_B_nFYobDWW9_1(.din(w_dff_B_mNc6PFXQ0_1),.dout(w_dff_B_nFYobDWW9_1),.clk(gclk));
	jdff dff_B_AmehRiI93_1(.din(w_dff_B_nFYobDWW9_1),.dout(w_dff_B_AmehRiI93_1),.clk(gclk));
	jdff dff_B_YCHQ6EdZ0_1(.din(w_dff_B_AmehRiI93_1),.dout(w_dff_B_YCHQ6EdZ0_1),.clk(gclk));
	jdff dff_B_n1SoDHzL9_1(.din(w_dff_B_YCHQ6EdZ0_1),.dout(w_dff_B_n1SoDHzL9_1),.clk(gclk));
	jdff dff_B_DLIX49hN9_1(.din(w_dff_B_n1SoDHzL9_1),.dout(w_dff_B_DLIX49hN9_1),.clk(gclk));
	jdff dff_B_k8xOooFM4_1(.din(w_dff_B_DLIX49hN9_1),.dout(w_dff_B_k8xOooFM4_1),.clk(gclk));
	jdff dff_B_XwnUYPgR2_1(.din(w_dff_B_k8xOooFM4_1),.dout(w_dff_B_XwnUYPgR2_1),.clk(gclk));
	jdff dff_B_3UQkUfI68_1(.din(w_dff_B_XwnUYPgR2_1),.dout(w_dff_B_3UQkUfI68_1),.clk(gclk));
	jdff dff_B_POirTfb49_1(.din(w_dff_B_3UQkUfI68_1),.dout(w_dff_B_POirTfb49_1),.clk(gclk));
	jdff dff_B_Jm5xqbpj7_1(.din(w_dff_B_POirTfb49_1),.dout(w_dff_B_Jm5xqbpj7_1),.clk(gclk));
	jdff dff_B_sgnaPnVx9_1(.din(w_dff_B_Jm5xqbpj7_1),.dout(w_dff_B_sgnaPnVx9_1),.clk(gclk));
	jdff dff_B_zxY0mHzY3_1(.din(w_dff_B_sgnaPnVx9_1),.dout(w_dff_B_zxY0mHzY3_1),.clk(gclk));
	jdff dff_B_iWu0Xn025_1(.din(w_dff_B_zxY0mHzY3_1),.dout(w_dff_B_iWu0Xn025_1),.clk(gclk));
	jdff dff_B_VGUWiZmZ8_1(.din(w_dff_B_iWu0Xn025_1),.dout(w_dff_B_VGUWiZmZ8_1),.clk(gclk));
	jdff dff_B_w3E6nsfT5_1(.din(w_dff_B_VGUWiZmZ8_1),.dout(w_dff_B_w3E6nsfT5_1),.clk(gclk));
	jdff dff_B_5nh3WXtJ0_1(.din(w_dff_B_w3E6nsfT5_1),.dout(w_dff_B_5nh3WXtJ0_1),.clk(gclk));
	jdff dff_B_VkNunJB06_1(.din(w_dff_B_5nh3WXtJ0_1),.dout(w_dff_B_VkNunJB06_1),.clk(gclk));
	jdff dff_B_2xeLz8H77_1(.din(w_dff_B_VkNunJB06_1),.dout(w_dff_B_2xeLz8H77_1),.clk(gclk));
	jdff dff_B_nvl1DsuF6_0(.din(n811),.dout(w_dff_B_nvl1DsuF6_0),.clk(gclk));
	jdff dff_B_UxUSEnrq9_0(.din(w_dff_B_nvl1DsuF6_0),.dout(w_dff_B_UxUSEnrq9_0),.clk(gclk));
	jdff dff_B_qk7OKlME8_0(.din(w_dff_B_UxUSEnrq9_0),.dout(w_dff_B_qk7OKlME8_0),.clk(gclk));
	jdff dff_B_ljzoi7Gx0_0(.din(w_dff_B_qk7OKlME8_0),.dout(w_dff_B_ljzoi7Gx0_0),.clk(gclk));
	jdff dff_B_GyxbHnTi1_0(.din(w_dff_B_ljzoi7Gx0_0),.dout(w_dff_B_GyxbHnTi1_0),.clk(gclk));
	jdff dff_B_RF2xT56F1_0(.din(w_dff_B_GyxbHnTi1_0),.dout(w_dff_B_RF2xT56F1_0),.clk(gclk));
	jdff dff_B_qtiZPLq51_0(.din(w_dff_B_RF2xT56F1_0),.dout(w_dff_B_qtiZPLq51_0),.clk(gclk));
	jdff dff_B_poDzi82x6_0(.din(w_dff_B_qtiZPLq51_0),.dout(w_dff_B_poDzi82x6_0),.clk(gclk));
	jdff dff_B_F7jtAGL09_0(.din(w_dff_B_poDzi82x6_0),.dout(w_dff_B_F7jtAGL09_0),.clk(gclk));
	jdff dff_B_u5nVXoww7_0(.din(w_dff_B_F7jtAGL09_0),.dout(w_dff_B_u5nVXoww7_0),.clk(gclk));
	jdff dff_B_TT9lRUQV8_0(.din(w_dff_B_u5nVXoww7_0),.dout(w_dff_B_TT9lRUQV8_0),.clk(gclk));
	jdff dff_B_xUbNhu9M1_0(.din(w_dff_B_TT9lRUQV8_0),.dout(w_dff_B_xUbNhu9M1_0),.clk(gclk));
	jdff dff_B_TjgeKRwY9_0(.din(w_dff_B_xUbNhu9M1_0),.dout(w_dff_B_TjgeKRwY9_0),.clk(gclk));
	jdff dff_B_k8kRByqR6_0(.din(w_dff_B_TjgeKRwY9_0),.dout(w_dff_B_k8kRByqR6_0),.clk(gclk));
	jdff dff_B_tnZDjq6y5_0(.din(w_dff_B_k8kRByqR6_0),.dout(w_dff_B_tnZDjq6y5_0),.clk(gclk));
	jdff dff_B_rCJs1lad9_0(.din(w_dff_B_tnZDjq6y5_0),.dout(w_dff_B_rCJs1lad9_0),.clk(gclk));
	jdff dff_B_PoxsRFmk6_0(.din(w_dff_B_rCJs1lad9_0),.dout(w_dff_B_PoxsRFmk6_0),.clk(gclk));
	jdff dff_B_dd5hwphR4_0(.din(w_dff_B_PoxsRFmk6_0),.dout(w_dff_B_dd5hwphR4_0),.clk(gclk));
	jdff dff_B_CNylEeYP7_0(.din(w_dff_B_dd5hwphR4_0),.dout(w_dff_B_CNylEeYP7_0),.clk(gclk));
	jdff dff_B_At2ilMbM0_0(.din(w_dff_B_CNylEeYP7_0),.dout(w_dff_B_At2ilMbM0_0),.clk(gclk));
	jdff dff_B_Jd4F5Olk6_0(.din(w_dff_B_At2ilMbM0_0),.dout(w_dff_B_Jd4F5Olk6_0),.clk(gclk));
	jdff dff_B_4QhqIe667_0(.din(w_dff_B_Jd4F5Olk6_0),.dout(w_dff_B_4QhqIe667_0),.clk(gclk));
	jdff dff_B_i9pUHtxJ6_0(.din(w_dff_B_4QhqIe667_0),.dout(w_dff_B_i9pUHtxJ6_0),.clk(gclk));
	jdff dff_B_uRen2yrE3_0(.din(w_dff_B_i9pUHtxJ6_0),.dout(w_dff_B_uRen2yrE3_0),.clk(gclk));
	jdff dff_B_vafBg3Vk3_0(.din(w_dff_B_uRen2yrE3_0),.dout(w_dff_B_vafBg3Vk3_0),.clk(gclk));
	jdff dff_B_xuIisjlp4_0(.din(w_dff_B_vafBg3Vk3_0),.dout(w_dff_B_xuIisjlp4_0),.clk(gclk));
	jdff dff_B_eWLD32ma0_0(.din(w_dff_B_xuIisjlp4_0),.dout(w_dff_B_eWLD32ma0_0),.clk(gclk));
	jdff dff_B_SNQz7Q316_0(.din(w_dff_B_eWLD32ma0_0),.dout(w_dff_B_SNQz7Q316_0),.clk(gclk));
	jdff dff_B_GsUAQ68U8_0(.din(w_dff_B_SNQz7Q316_0),.dout(w_dff_B_GsUAQ68U8_0),.clk(gclk));
	jdff dff_B_RSaTXRfz7_0(.din(w_dff_B_GsUAQ68U8_0),.dout(w_dff_B_RSaTXRfz7_0),.clk(gclk));
	jdff dff_B_USp6mICs2_0(.din(w_dff_B_RSaTXRfz7_0),.dout(w_dff_B_USp6mICs2_0),.clk(gclk));
	jdff dff_B_4ExvazqS9_0(.din(w_dff_B_USp6mICs2_0),.dout(w_dff_B_4ExvazqS9_0),.clk(gclk));
	jdff dff_B_Jd1gpXR12_0(.din(w_dff_B_4ExvazqS9_0),.dout(w_dff_B_Jd1gpXR12_0),.clk(gclk));
	jdff dff_B_5M7EyEsQ4_0(.din(w_dff_B_Jd1gpXR12_0),.dout(w_dff_B_5M7EyEsQ4_0),.clk(gclk));
	jdff dff_B_IcM4Ep1U6_0(.din(w_dff_B_5M7EyEsQ4_0),.dout(w_dff_B_IcM4Ep1U6_0),.clk(gclk));
	jdff dff_B_I4kbpMhW8_0(.din(w_dff_B_IcM4Ep1U6_0),.dout(w_dff_B_I4kbpMhW8_0),.clk(gclk));
	jdff dff_B_S3z89LHJ1_0(.din(w_dff_B_I4kbpMhW8_0),.dout(w_dff_B_S3z89LHJ1_0),.clk(gclk));
	jdff dff_B_XLnaXlOQ9_0(.din(w_dff_B_S3z89LHJ1_0),.dout(w_dff_B_XLnaXlOQ9_0),.clk(gclk));
	jdff dff_B_h5fbgJQb2_0(.din(w_dff_B_XLnaXlOQ9_0),.dout(w_dff_B_h5fbgJQb2_0),.clk(gclk));
	jdff dff_B_4HukJdoK4_0(.din(w_dff_B_h5fbgJQb2_0),.dout(w_dff_B_4HukJdoK4_0),.clk(gclk));
	jdff dff_B_5IG5ManI3_0(.din(w_dff_B_4HukJdoK4_0),.dout(w_dff_B_5IG5ManI3_0),.clk(gclk));
	jdff dff_B_rkLa2H1l3_0(.din(w_dff_B_5IG5ManI3_0),.dout(w_dff_B_rkLa2H1l3_0),.clk(gclk));
	jdff dff_B_ZEcAbrYv0_0(.din(w_dff_B_rkLa2H1l3_0),.dout(w_dff_B_ZEcAbrYv0_0),.clk(gclk));
	jdff dff_B_2E1Auvo42_0(.din(w_dff_B_ZEcAbrYv0_0),.dout(w_dff_B_2E1Auvo42_0),.clk(gclk));
	jdff dff_B_3isJtvCp9_0(.din(w_dff_B_2E1Auvo42_0),.dout(w_dff_B_3isJtvCp9_0),.clk(gclk));
	jdff dff_B_rW8HDDwB0_0(.din(w_dff_B_3isJtvCp9_0),.dout(w_dff_B_rW8HDDwB0_0),.clk(gclk));
	jdff dff_B_rM39nGdq6_0(.din(w_dff_B_rW8HDDwB0_0),.dout(w_dff_B_rM39nGdq6_0),.clk(gclk));
	jdff dff_B_0wB66zH80_0(.din(w_dff_B_rM39nGdq6_0),.dout(w_dff_B_0wB66zH80_0),.clk(gclk));
	jdff dff_B_oFUvSo5u3_0(.din(w_dff_B_0wB66zH80_0),.dout(w_dff_B_oFUvSo5u3_0),.clk(gclk));
	jdff dff_B_NOZCM0cf2_0(.din(w_dff_B_oFUvSo5u3_0),.dout(w_dff_B_NOZCM0cf2_0),.clk(gclk));
	jdff dff_B_x0K9wlQz2_0(.din(w_dff_B_NOZCM0cf2_0),.dout(w_dff_B_x0K9wlQz2_0),.clk(gclk));
	jdff dff_B_NhC7MEUy1_0(.din(w_dff_B_x0K9wlQz2_0),.dout(w_dff_B_NhC7MEUy1_0),.clk(gclk));
	jdff dff_B_vRFCuuG98_0(.din(w_dff_B_NhC7MEUy1_0),.dout(w_dff_B_vRFCuuG98_0),.clk(gclk));
	jdff dff_B_UzQOeXxz6_0(.din(w_dff_B_vRFCuuG98_0),.dout(w_dff_B_UzQOeXxz6_0),.clk(gclk));
	jdff dff_B_uuGrenYI4_0(.din(w_dff_B_UzQOeXxz6_0),.dout(w_dff_B_uuGrenYI4_0),.clk(gclk));
	jdff dff_B_HfD8uDU70_0(.din(w_dff_B_uuGrenYI4_0),.dout(w_dff_B_HfD8uDU70_0),.clk(gclk));
	jdff dff_B_hfjeN3Wx6_0(.din(w_dff_B_HfD8uDU70_0),.dout(w_dff_B_hfjeN3Wx6_0),.clk(gclk));
	jdff dff_B_ECUwhUDy0_0(.din(w_dff_B_hfjeN3Wx6_0),.dout(w_dff_B_ECUwhUDy0_0),.clk(gclk));
	jdff dff_B_fU2RXRtI8_0(.din(w_dff_B_ECUwhUDy0_0),.dout(w_dff_B_fU2RXRtI8_0),.clk(gclk));
	jdff dff_B_CbEXAH8a8_0(.din(w_dff_B_fU2RXRtI8_0),.dout(w_dff_B_CbEXAH8a8_0),.clk(gclk));
	jdff dff_B_iR9EAUy26_0(.din(w_dff_B_CbEXAH8a8_0),.dout(w_dff_B_iR9EAUy26_0),.clk(gclk));
	jdff dff_B_Le0kiDce0_0(.din(w_dff_B_iR9EAUy26_0),.dout(w_dff_B_Le0kiDce0_0),.clk(gclk));
	jdff dff_B_7QGzODXK6_0(.din(w_dff_B_Le0kiDce0_0),.dout(w_dff_B_7QGzODXK6_0),.clk(gclk));
	jdff dff_B_fRDxdxij7_0(.din(w_dff_B_7QGzODXK6_0),.dout(w_dff_B_fRDxdxij7_0),.clk(gclk));
	jdff dff_B_c4Pa7EKc0_0(.din(w_dff_B_fRDxdxij7_0),.dout(w_dff_B_c4Pa7EKc0_0),.clk(gclk));
	jdff dff_B_nQwA0zln9_0(.din(w_dff_B_c4Pa7EKc0_0),.dout(w_dff_B_nQwA0zln9_0),.clk(gclk));
	jdff dff_B_LmJdCNY68_0(.din(w_dff_B_nQwA0zln9_0),.dout(w_dff_B_LmJdCNY68_0),.clk(gclk));
	jdff dff_B_hgg32NFA5_0(.din(w_dff_B_LmJdCNY68_0),.dout(w_dff_B_hgg32NFA5_0),.clk(gclk));
	jdff dff_B_m9LK9m683_0(.din(w_dff_B_hgg32NFA5_0),.dout(w_dff_B_m9LK9m683_0),.clk(gclk));
	jdff dff_B_FuCsEnzB2_0(.din(w_dff_B_m9LK9m683_0),.dout(w_dff_B_FuCsEnzB2_0),.clk(gclk));
	jdff dff_B_opoKmvzR0_0(.din(w_dff_B_FuCsEnzB2_0),.dout(w_dff_B_opoKmvzR0_0),.clk(gclk));
	jdff dff_B_fPtnV4ne1_1(.din(n804),.dout(w_dff_B_fPtnV4ne1_1),.clk(gclk));
	jdff dff_B_u5KB2iBC0_1(.din(w_dff_B_fPtnV4ne1_1),.dout(w_dff_B_u5KB2iBC0_1),.clk(gclk));
	jdff dff_B_jdWkOwwN7_1(.din(w_dff_B_u5KB2iBC0_1),.dout(w_dff_B_jdWkOwwN7_1),.clk(gclk));
	jdff dff_B_uwYk1ykc6_1(.din(w_dff_B_jdWkOwwN7_1),.dout(w_dff_B_uwYk1ykc6_1),.clk(gclk));
	jdff dff_B_SiluVxBi9_1(.din(w_dff_B_uwYk1ykc6_1),.dout(w_dff_B_SiluVxBi9_1),.clk(gclk));
	jdff dff_B_VAACcGSx5_1(.din(w_dff_B_SiluVxBi9_1),.dout(w_dff_B_VAACcGSx5_1),.clk(gclk));
	jdff dff_B_h3w4uTr13_1(.din(w_dff_B_VAACcGSx5_1),.dout(w_dff_B_h3w4uTr13_1),.clk(gclk));
	jdff dff_B_39zBnsb43_1(.din(w_dff_B_h3w4uTr13_1),.dout(w_dff_B_39zBnsb43_1),.clk(gclk));
	jdff dff_B_aZtWOlo36_1(.din(w_dff_B_39zBnsb43_1),.dout(w_dff_B_aZtWOlo36_1),.clk(gclk));
	jdff dff_B_A1Dsif1O2_1(.din(w_dff_B_aZtWOlo36_1),.dout(w_dff_B_A1Dsif1O2_1),.clk(gclk));
	jdff dff_B_UNfAREHO0_1(.din(w_dff_B_A1Dsif1O2_1),.dout(w_dff_B_UNfAREHO0_1),.clk(gclk));
	jdff dff_B_Sgz1soDP7_1(.din(w_dff_B_UNfAREHO0_1),.dout(w_dff_B_Sgz1soDP7_1),.clk(gclk));
	jdff dff_B_2JK0dxAD0_1(.din(w_dff_B_Sgz1soDP7_1),.dout(w_dff_B_2JK0dxAD0_1),.clk(gclk));
	jdff dff_B_iFw6OVHl8_1(.din(w_dff_B_2JK0dxAD0_1),.dout(w_dff_B_iFw6OVHl8_1),.clk(gclk));
	jdff dff_B_RjclR5278_1(.din(w_dff_B_iFw6OVHl8_1),.dout(w_dff_B_RjclR5278_1),.clk(gclk));
	jdff dff_B_6uAudWPB3_1(.din(w_dff_B_RjclR5278_1),.dout(w_dff_B_6uAudWPB3_1),.clk(gclk));
	jdff dff_B_plIOSQUf0_1(.din(w_dff_B_6uAudWPB3_1),.dout(w_dff_B_plIOSQUf0_1),.clk(gclk));
	jdff dff_B_jKEPCnNX6_1(.din(w_dff_B_plIOSQUf0_1),.dout(w_dff_B_jKEPCnNX6_1),.clk(gclk));
	jdff dff_B_YVaQyCet2_1(.din(w_dff_B_jKEPCnNX6_1),.dout(w_dff_B_YVaQyCet2_1),.clk(gclk));
	jdff dff_B_iz4QeOnO6_1(.din(w_dff_B_YVaQyCet2_1),.dout(w_dff_B_iz4QeOnO6_1),.clk(gclk));
	jdff dff_B_rFPliHwR7_1(.din(w_dff_B_iz4QeOnO6_1),.dout(w_dff_B_rFPliHwR7_1),.clk(gclk));
	jdff dff_B_awJCPDGO5_1(.din(w_dff_B_rFPliHwR7_1),.dout(w_dff_B_awJCPDGO5_1),.clk(gclk));
	jdff dff_B_2C25k7Jb7_1(.din(w_dff_B_awJCPDGO5_1),.dout(w_dff_B_2C25k7Jb7_1),.clk(gclk));
	jdff dff_B_rVS7Kz5u7_1(.din(w_dff_B_2C25k7Jb7_1),.dout(w_dff_B_rVS7Kz5u7_1),.clk(gclk));
	jdff dff_B_trc6snZY1_1(.din(w_dff_B_rVS7Kz5u7_1),.dout(w_dff_B_trc6snZY1_1),.clk(gclk));
	jdff dff_B_eQjwPyqC5_1(.din(w_dff_B_trc6snZY1_1),.dout(w_dff_B_eQjwPyqC5_1),.clk(gclk));
	jdff dff_B_jP9xQUtG5_1(.din(w_dff_B_eQjwPyqC5_1),.dout(w_dff_B_jP9xQUtG5_1),.clk(gclk));
	jdff dff_B_jqdsOLBy4_1(.din(w_dff_B_jP9xQUtG5_1),.dout(w_dff_B_jqdsOLBy4_1),.clk(gclk));
	jdff dff_B_9wvJyR1H1_1(.din(w_dff_B_jqdsOLBy4_1),.dout(w_dff_B_9wvJyR1H1_1),.clk(gclk));
	jdff dff_B_5tdoIqmD1_1(.din(w_dff_B_9wvJyR1H1_1),.dout(w_dff_B_5tdoIqmD1_1),.clk(gclk));
	jdff dff_B_1McRnk3w4_1(.din(w_dff_B_5tdoIqmD1_1),.dout(w_dff_B_1McRnk3w4_1),.clk(gclk));
	jdff dff_B_NuFG2oGH1_1(.din(w_dff_B_1McRnk3w4_1),.dout(w_dff_B_NuFG2oGH1_1),.clk(gclk));
	jdff dff_B_0NdLb2sr3_1(.din(w_dff_B_NuFG2oGH1_1),.dout(w_dff_B_0NdLb2sr3_1),.clk(gclk));
	jdff dff_B_EdpR58VJ4_1(.din(w_dff_B_0NdLb2sr3_1),.dout(w_dff_B_EdpR58VJ4_1),.clk(gclk));
	jdff dff_B_vCoVINpe7_1(.din(w_dff_B_EdpR58VJ4_1),.dout(w_dff_B_vCoVINpe7_1),.clk(gclk));
	jdff dff_B_q3H8vo2M7_1(.din(w_dff_B_vCoVINpe7_1),.dout(w_dff_B_q3H8vo2M7_1),.clk(gclk));
	jdff dff_B_gU6I6iIH9_1(.din(w_dff_B_q3H8vo2M7_1),.dout(w_dff_B_gU6I6iIH9_1),.clk(gclk));
	jdff dff_B_X8rZibmw1_1(.din(w_dff_B_gU6I6iIH9_1),.dout(w_dff_B_X8rZibmw1_1),.clk(gclk));
	jdff dff_B_8BSjqyq00_1(.din(w_dff_B_X8rZibmw1_1),.dout(w_dff_B_8BSjqyq00_1),.clk(gclk));
	jdff dff_B_MZKGPgIk0_1(.din(w_dff_B_8BSjqyq00_1),.dout(w_dff_B_MZKGPgIk0_1),.clk(gclk));
	jdff dff_B_vfoBeLG48_1(.din(w_dff_B_MZKGPgIk0_1),.dout(w_dff_B_vfoBeLG48_1),.clk(gclk));
	jdff dff_B_pxtXzr5M9_1(.din(w_dff_B_vfoBeLG48_1),.dout(w_dff_B_pxtXzr5M9_1),.clk(gclk));
	jdff dff_B_akxC9Onn9_1(.din(w_dff_B_pxtXzr5M9_1),.dout(w_dff_B_akxC9Onn9_1),.clk(gclk));
	jdff dff_B_kAmT2Wwo3_1(.din(w_dff_B_akxC9Onn9_1),.dout(w_dff_B_kAmT2Wwo3_1),.clk(gclk));
	jdff dff_B_x9OiuhUO1_1(.din(w_dff_B_kAmT2Wwo3_1),.dout(w_dff_B_x9OiuhUO1_1),.clk(gclk));
	jdff dff_B_sDbcG5VX0_1(.din(w_dff_B_x9OiuhUO1_1),.dout(w_dff_B_sDbcG5VX0_1),.clk(gclk));
	jdff dff_B_ohXgzFRg6_1(.din(w_dff_B_sDbcG5VX0_1),.dout(w_dff_B_ohXgzFRg6_1),.clk(gclk));
	jdff dff_B_tuFLE2z73_1(.din(w_dff_B_ohXgzFRg6_1),.dout(w_dff_B_tuFLE2z73_1),.clk(gclk));
	jdff dff_B_a8Wm1DCm6_1(.din(w_dff_B_tuFLE2z73_1),.dout(w_dff_B_a8Wm1DCm6_1),.clk(gclk));
	jdff dff_B_nTMYM4Ce6_1(.din(w_dff_B_a8Wm1DCm6_1),.dout(w_dff_B_nTMYM4Ce6_1),.clk(gclk));
	jdff dff_B_1Zj5aoxT5_1(.din(w_dff_B_nTMYM4Ce6_1),.dout(w_dff_B_1Zj5aoxT5_1),.clk(gclk));
	jdff dff_B_khpJAC276_1(.din(w_dff_B_1Zj5aoxT5_1),.dout(w_dff_B_khpJAC276_1),.clk(gclk));
	jdff dff_B_5h2KiXqU1_1(.din(w_dff_B_khpJAC276_1),.dout(w_dff_B_5h2KiXqU1_1),.clk(gclk));
	jdff dff_B_3OZt11gE3_1(.din(w_dff_B_5h2KiXqU1_1),.dout(w_dff_B_3OZt11gE3_1),.clk(gclk));
	jdff dff_B_Z14jyo114_1(.din(w_dff_B_3OZt11gE3_1),.dout(w_dff_B_Z14jyo114_1),.clk(gclk));
	jdff dff_B_vIyHb3Mq2_1(.din(w_dff_B_Z14jyo114_1),.dout(w_dff_B_vIyHb3Mq2_1),.clk(gclk));
	jdff dff_B_aCtDj9Ow4_1(.din(w_dff_B_vIyHb3Mq2_1),.dout(w_dff_B_aCtDj9Ow4_1),.clk(gclk));
	jdff dff_B_mR77MZ8I0_1(.din(w_dff_B_aCtDj9Ow4_1),.dout(w_dff_B_mR77MZ8I0_1),.clk(gclk));
	jdff dff_B_DBZVxHnp3_1(.din(w_dff_B_mR77MZ8I0_1),.dout(w_dff_B_DBZVxHnp3_1),.clk(gclk));
	jdff dff_B_AhsGIHbx2_1(.din(w_dff_B_DBZVxHnp3_1),.dout(w_dff_B_AhsGIHbx2_1),.clk(gclk));
	jdff dff_B_yhVf4j9i5_1(.din(w_dff_B_AhsGIHbx2_1),.dout(w_dff_B_yhVf4j9i5_1),.clk(gclk));
	jdff dff_B_u2csuEJ05_1(.din(w_dff_B_yhVf4j9i5_1),.dout(w_dff_B_u2csuEJ05_1),.clk(gclk));
	jdff dff_B_qgLzhbVe3_1(.din(w_dff_B_u2csuEJ05_1),.dout(w_dff_B_qgLzhbVe3_1),.clk(gclk));
	jdff dff_B_QWLTNVuz7_1(.din(w_dff_B_qgLzhbVe3_1),.dout(w_dff_B_QWLTNVuz7_1),.clk(gclk));
	jdff dff_B_Nn3e0hev5_1(.din(w_dff_B_QWLTNVuz7_1),.dout(w_dff_B_Nn3e0hev5_1),.clk(gclk));
	jdff dff_B_aCH4LLod8_1(.din(w_dff_B_Nn3e0hev5_1),.dout(w_dff_B_aCH4LLod8_1),.clk(gclk));
	jdff dff_B_shoRslMY0_1(.din(w_dff_B_aCH4LLod8_1),.dout(w_dff_B_shoRslMY0_1),.clk(gclk));
	jdff dff_B_uXXOUjCv2_1(.din(w_dff_B_shoRslMY0_1),.dout(w_dff_B_uXXOUjCv2_1),.clk(gclk));
	jdff dff_B_9VcyI3r83_1(.din(w_dff_B_uXXOUjCv2_1),.dout(w_dff_B_9VcyI3r83_1),.clk(gclk));
	jdff dff_B_pVF4M0wG0_1(.din(w_dff_B_9VcyI3r83_1),.dout(w_dff_B_pVF4M0wG0_1),.clk(gclk));
	jdff dff_B_5Ni2CrgP5_0(.din(n805),.dout(w_dff_B_5Ni2CrgP5_0),.clk(gclk));
	jdff dff_B_FSDDnmCR6_0(.din(w_dff_B_5Ni2CrgP5_0),.dout(w_dff_B_FSDDnmCR6_0),.clk(gclk));
	jdff dff_B_UM8lSR7m2_0(.din(w_dff_B_FSDDnmCR6_0),.dout(w_dff_B_UM8lSR7m2_0),.clk(gclk));
	jdff dff_B_D21i3gug7_0(.din(w_dff_B_UM8lSR7m2_0),.dout(w_dff_B_D21i3gug7_0),.clk(gclk));
	jdff dff_B_9ObiCvZv1_0(.din(w_dff_B_D21i3gug7_0),.dout(w_dff_B_9ObiCvZv1_0),.clk(gclk));
	jdff dff_B_Lm0XaGbR3_0(.din(w_dff_B_9ObiCvZv1_0),.dout(w_dff_B_Lm0XaGbR3_0),.clk(gclk));
	jdff dff_B_2YMpziwZ3_0(.din(w_dff_B_Lm0XaGbR3_0),.dout(w_dff_B_2YMpziwZ3_0),.clk(gclk));
	jdff dff_B_C44ROdL24_0(.din(w_dff_B_2YMpziwZ3_0),.dout(w_dff_B_C44ROdL24_0),.clk(gclk));
	jdff dff_B_TabcxDqg2_0(.din(w_dff_B_C44ROdL24_0),.dout(w_dff_B_TabcxDqg2_0),.clk(gclk));
	jdff dff_B_h2KZ6CGk5_0(.din(w_dff_B_TabcxDqg2_0),.dout(w_dff_B_h2KZ6CGk5_0),.clk(gclk));
	jdff dff_B_sAvbZ5hM3_0(.din(w_dff_B_h2KZ6CGk5_0),.dout(w_dff_B_sAvbZ5hM3_0),.clk(gclk));
	jdff dff_B_quVmLe8D7_0(.din(w_dff_B_sAvbZ5hM3_0),.dout(w_dff_B_quVmLe8D7_0),.clk(gclk));
	jdff dff_B_vdaOlCqG6_0(.din(w_dff_B_quVmLe8D7_0),.dout(w_dff_B_vdaOlCqG6_0),.clk(gclk));
	jdff dff_B_yQqVSCO33_0(.din(w_dff_B_vdaOlCqG6_0),.dout(w_dff_B_yQqVSCO33_0),.clk(gclk));
	jdff dff_B_eH7kOKHS9_0(.din(w_dff_B_yQqVSCO33_0),.dout(w_dff_B_eH7kOKHS9_0),.clk(gclk));
	jdff dff_B_FLRfAfIX1_0(.din(w_dff_B_eH7kOKHS9_0),.dout(w_dff_B_FLRfAfIX1_0),.clk(gclk));
	jdff dff_B_kGFRuOZH4_0(.din(w_dff_B_FLRfAfIX1_0),.dout(w_dff_B_kGFRuOZH4_0),.clk(gclk));
	jdff dff_B_eXcRlOOD7_0(.din(w_dff_B_kGFRuOZH4_0),.dout(w_dff_B_eXcRlOOD7_0),.clk(gclk));
	jdff dff_B_TaQKXIL92_0(.din(w_dff_B_eXcRlOOD7_0),.dout(w_dff_B_TaQKXIL92_0),.clk(gclk));
	jdff dff_B_7sHwa8Mc9_0(.din(w_dff_B_TaQKXIL92_0),.dout(w_dff_B_7sHwa8Mc9_0),.clk(gclk));
	jdff dff_B_zO5Y0dJj3_0(.din(w_dff_B_7sHwa8Mc9_0),.dout(w_dff_B_zO5Y0dJj3_0),.clk(gclk));
	jdff dff_B_FUHHROpm6_0(.din(w_dff_B_zO5Y0dJj3_0),.dout(w_dff_B_FUHHROpm6_0),.clk(gclk));
	jdff dff_B_hg6yJ2KZ4_0(.din(w_dff_B_FUHHROpm6_0),.dout(w_dff_B_hg6yJ2KZ4_0),.clk(gclk));
	jdff dff_B_3U56scaO3_0(.din(w_dff_B_hg6yJ2KZ4_0),.dout(w_dff_B_3U56scaO3_0),.clk(gclk));
	jdff dff_B_0IdauRGb0_0(.din(w_dff_B_3U56scaO3_0),.dout(w_dff_B_0IdauRGb0_0),.clk(gclk));
	jdff dff_B_6E5XANT57_0(.din(w_dff_B_0IdauRGb0_0),.dout(w_dff_B_6E5XANT57_0),.clk(gclk));
	jdff dff_B_0LwHkpT39_0(.din(w_dff_B_6E5XANT57_0),.dout(w_dff_B_0LwHkpT39_0),.clk(gclk));
	jdff dff_B_W5LqX5Ho0_0(.din(w_dff_B_0LwHkpT39_0),.dout(w_dff_B_W5LqX5Ho0_0),.clk(gclk));
	jdff dff_B_GB0jboq45_0(.din(w_dff_B_W5LqX5Ho0_0),.dout(w_dff_B_GB0jboq45_0),.clk(gclk));
	jdff dff_B_RfGtvzon1_0(.din(w_dff_B_GB0jboq45_0),.dout(w_dff_B_RfGtvzon1_0),.clk(gclk));
	jdff dff_B_vA3eJbty0_0(.din(w_dff_B_RfGtvzon1_0),.dout(w_dff_B_vA3eJbty0_0),.clk(gclk));
	jdff dff_B_fMkP9Uic2_0(.din(w_dff_B_vA3eJbty0_0),.dout(w_dff_B_fMkP9Uic2_0),.clk(gclk));
	jdff dff_B_hyPuF6Ow8_0(.din(w_dff_B_fMkP9Uic2_0),.dout(w_dff_B_hyPuF6Ow8_0),.clk(gclk));
	jdff dff_B_RIhNgZz05_0(.din(w_dff_B_hyPuF6Ow8_0),.dout(w_dff_B_RIhNgZz05_0),.clk(gclk));
	jdff dff_B_EKHbUWMj5_0(.din(w_dff_B_RIhNgZz05_0),.dout(w_dff_B_EKHbUWMj5_0),.clk(gclk));
	jdff dff_B_geDmSBno5_0(.din(w_dff_B_EKHbUWMj5_0),.dout(w_dff_B_geDmSBno5_0),.clk(gclk));
	jdff dff_B_OriJUwel6_0(.din(w_dff_B_geDmSBno5_0),.dout(w_dff_B_OriJUwel6_0),.clk(gclk));
	jdff dff_B_xgMQCIlB4_0(.din(w_dff_B_OriJUwel6_0),.dout(w_dff_B_xgMQCIlB4_0),.clk(gclk));
	jdff dff_B_zsbImneq4_0(.din(w_dff_B_xgMQCIlB4_0),.dout(w_dff_B_zsbImneq4_0),.clk(gclk));
	jdff dff_B_sk0oR1Kf4_0(.din(w_dff_B_zsbImneq4_0),.dout(w_dff_B_sk0oR1Kf4_0),.clk(gclk));
	jdff dff_B_q3RSenw00_0(.din(w_dff_B_sk0oR1Kf4_0),.dout(w_dff_B_q3RSenw00_0),.clk(gclk));
	jdff dff_B_Tx9pgges0_0(.din(w_dff_B_q3RSenw00_0),.dout(w_dff_B_Tx9pgges0_0),.clk(gclk));
	jdff dff_B_1PuhqfBk1_0(.din(w_dff_B_Tx9pgges0_0),.dout(w_dff_B_1PuhqfBk1_0),.clk(gclk));
	jdff dff_B_S3oheR1K1_0(.din(w_dff_B_1PuhqfBk1_0),.dout(w_dff_B_S3oheR1K1_0),.clk(gclk));
	jdff dff_B_lxh7nCk79_0(.din(w_dff_B_S3oheR1K1_0),.dout(w_dff_B_lxh7nCk79_0),.clk(gclk));
	jdff dff_B_T7cWo3xx4_0(.din(w_dff_B_lxh7nCk79_0),.dout(w_dff_B_T7cWo3xx4_0),.clk(gclk));
	jdff dff_B_7GSxoU2g5_0(.din(w_dff_B_T7cWo3xx4_0),.dout(w_dff_B_7GSxoU2g5_0),.clk(gclk));
	jdff dff_B_zHi0uYkY5_0(.din(w_dff_B_7GSxoU2g5_0),.dout(w_dff_B_zHi0uYkY5_0),.clk(gclk));
	jdff dff_B_eGWX7n3w8_0(.din(w_dff_B_zHi0uYkY5_0),.dout(w_dff_B_eGWX7n3w8_0),.clk(gclk));
	jdff dff_B_h0nfvhi62_0(.din(w_dff_B_eGWX7n3w8_0),.dout(w_dff_B_h0nfvhi62_0),.clk(gclk));
	jdff dff_B_vFEo9h5K5_0(.din(w_dff_B_h0nfvhi62_0),.dout(w_dff_B_vFEo9h5K5_0),.clk(gclk));
	jdff dff_B_0SoYbOul9_0(.din(w_dff_B_vFEo9h5K5_0),.dout(w_dff_B_0SoYbOul9_0),.clk(gclk));
	jdff dff_B_mpidmNvA2_0(.din(w_dff_B_0SoYbOul9_0),.dout(w_dff_B_mpidmNvA2_0),.clk(gclk));
	jdff dff_B_1MmgSsZ66_0(.din(w_dff_B_mpidmNvA2_0),.dout(w_dff_B_1MmgSsZ66_0),.clk(gclk));
	jdff dff_B_3azS8yEz2_0(.din(w_dff_B_1MmgSsZ66_0),.dout(w_dff_B_3azS8yEz2_0),.clk(gclk));
	jdff dff_B_dYF03m3J8_0(.din(w_dff_B_3azS8yEz2_0),.dout(w_dff_B_dYF03m3J8_0),.clk(gclk));
	jdff dff_B_7wkog4mP8_0(.din(w_dff_B_dYF03m3J8_0),.dout(w_dff_B_7wkog4mP8_0),.clk(gclk));
	jdff dff_B_mOWiLkdh4_0(.din(w_dff_B_7wkog4mP8_0),.dout(w_dff_B_mOWiLkdh4_0),.clk(gclk));
	jdff dff_B_6AcOMnso4_0(.din(w_dff_B_mOWiLkdh4_0),.dout(w_dff_B_6AcOMnso4_0),.clk(gclk));
	jdff dff_B_OTTj2QL28_0(.din(w_dff_B_6AcOMnso4_0),.dout(w_dff_B_OTTj2QL28_0),.clk(gclk));
	jdff dff_B_VYksLNI65_0(.din(w_dff_B_OTTj2QL28_0),.dout(w_dff_B_VYksLNI65_0),.clk(gclk));
	jdff dff_B_Z8NxScdf1_0(.din(w_dff_B_VYksLNI65_0),.dout(w_dff_B_Z8NxScdf1_0),.clk(gclk));
	jdff dff_B_3ldWa6gA5_0(.din(w_dff_B_Z8NxScdf1_0),.dout(w_dff_B_3ldWa6gA5_0),.clk(gclk));
	jdff dff_B_C0O7QFSI4_0(.din(w_dff_B_3ldWa6gA5_0),.dout(w_dff_B_C0O7QFSI4_0),.clk(gclk));
	jdff dff_B_wSLYOuqJ4_0(.din(w_dff_B_C0O7QFSI4_0),.dout(w_dff_B_wSLYOuqJ4_0),.clk(gclk));
	jdff dff_B_JrId8InE1_0(.din(w_dff_B_wSLYOuqJ4_0),.dout(w_dff_B_JrId8InE1_0),.clk(gclk));
	jdff dff_B_7K3aF9Vz9_0(.din(w_dff_B_JrId8InE1_0),.dout(w_dff_B_7K3aF9Vz9_0),.clk(gclk));
	jdff dff_B_5f4GkgB66_0(.din(w_dff_B_7K3aF9Vz9_0),.dout(w_dff_B_5f4GkgB66_0),.clk(gclk));
	jdff dff_B_1ntz2iTa3_0(.din(w_dff_B_5f4GkgB66_0),.dout(w_dff_B_1ntz2iTa3_0),.clk(gclk));
	jdff dff_B_ok8xe67Q0_0(.din(w_dff_B_1ntz2iTa3_0),.dout(w_dff_B_ok8xe67Q0_0),.clk(gclk));
	jdff dff_B_ptW8XoVC7_1(.din(n798),.dout(w_dff_B_ptW8XoVC7_1),.clk(gclk));
	jdff dff_B_3pJQMJoW5_1(.din(w_dff_B_ptW8XoVC7_1),.dout(w_dff_B_3pJQMJoW5_1),.clk(gclk));
	jdff dff_B_cekGFxVL7_1(.din(w_dff_B_3pJQMJoW5_1),.dout(w_dff_B_cekGFxVL7_1),.clk(gclk));
	jdff dff_B_ixlxO9H45_1(.din(w_dff_B_cekGFxVL7_1),.dout(w_dff_B_ixlxO9H45_1),.clk(gclk));
	jdff dff_B_dA0IOJR33_1(.din(w_dff_B_ixlxO9H45_1),.dout(w_dff_B_dA0IOJR33_1),.clk(gclk));
	jdff dff_B_FlMMIyM59_1(.din(w_dff_B_dA0IOJR33_1),.dout(w_dff_B_FlMMIyM59_1),.clk(gclk));
	jdff dff_B_Jxka773Z0_1(.din(w_dff_B_FlMMIyM59_1),.dout(w_dff_B_Jxka773Z0_1),.clk(gclk));
	jdff dff_B_rdR2pFcl4_1(.din(w_dff_B_Jxka773Z0_1),.dout(w_dff_B_rdR2pFcl4_1),.clk(gclk));
	jdff dff_B_DTbs7MKm6_1(.din(w_dff_B_rdR2pFcl4_1),.dout(w_dff_B_DTbs7MKm6_1),.clk(gclk));
	jdff dff_B_XPvgE4Qs9_1(.din(w_dff_B_DTbs7MKm6_1),.dout(w_dff_B_XPvgE4Qs9_1),.clk(gclk));
	jdff dff_B_jz8Re5ZI2_1(.din(w_dff_B_XPvgE4Qs9_1),.dout(w_dff_B_jz8Re5ZI2_1),.clk(gclk));
	jdff dff_B_zJlMaynd1_1(.din(w_dff_B_jz8Re5ZI2_1),.dout(w_dff_B_zJlMaynd1_1),.clk(gclk));
	jdff dff_B_KqMN3XV17_1(.din(w_dff_B_zJlMaynd1_1),.dout(w_dff_B_KqMN3XV17_1),.clk(gclk));
	jdff dff_B_h1jjEvu12_1(.din(w_dff_B_KqMN3XV17_1),.dout(w_dff_B_h1jjEvu12_1),.clk(gclk));
	jdff dff_B_nmVmKBVL3_1(.din(w_dff_B_h1jjEvu12_1),.dout(w_dff_B_nmVmKBVL3_1),.clk(gclk));
	jdff dff_B_QTPcrAO08_1(.din(w_dff_B_nmVmKBVL3_1),.dout(w_dff_B_QTPcrAO08_1),.clk(gclk));
	jdff dff_B_KuOuFnyX7_1(.din(w_dff_B_QTPcrAO08_1),.dout(w_dff_B_KuOuFnyX7_1),.clk(gclk));
	jdff dff_B_MFUfr5Qa6_1(.din(w_dff_B_KuOuFnyX7_1),.dout(w_dff_B_MFUfr5Qa6_1),.clk(gclk));
	jdff dff_B_8qzSMwtE9_1(.din(w_dff_B_MFUfr5Qa6_1),.dout(w_dff_B_8qzSMwtE9_1),.clk(gclk));
	jdff dff_B_mxmjQZhX3_1(.din(w_dff_B_8qzSMwtE9_1),.dout(w_dff_B_mxmjQZhX3_1),.clk(gclk));
	jdff dff_B_nOE1QFe26_1(.din(w_dff_B_mxmjQZhX3_1),.dout(w_dff_B_nOE1QFe26_1),.clk(gclk));
	jdff dff_B_0YsZnwW28_1(.din(w_dff_B_nOE1QFe26_1),.dout(w_dff_B_0YsZnwW28_1),.clk(gclk));
	jdff dff_B_gfXIpjCS2_1(.din(w_dff_B_0YsZnwW28_1),.dout(w_dff_B_gfXIpjCS2_1),.clk(gclk));
	jdff dff_B_6Yu3s5tv7_1(.din(w_dff_B_gfXIpjCS2_1),.dout(w_dff_B_6Yu3s5tv7_1),.clk(gclk));
	jdff dff_B_8DQWRRrg3_1(.din(w_dff_B_6Yu3s5tv7_1),.dout(w_dff_B_8DQWRRrg3_1),.clk(gclk));
	jdff dff_B_D82Loipc7_1(.din(w_dff_B_8DQWRRrg3_1),.dout(w_dff_B_D82Loipc7_1),.clk(gclk));
	jdff dff_B_8r3015HU7_1(.din(w_dff_B_D82Loipc7_1),.dout(w_dff_B_8r3015HU7_1),.clk(gclk));
	jdff dff_B_JtQLUTeL5_1(.din(w_dff_B_8r3015HU7_1),.dout(w_dff_B_JtQLUTeL5_1),.clk(gclk));
	jdff dff_B_8Cr0TDEK8_1(.din(w_dff_B_JtQLUTeL5_1),.dout(w_dff_B_8Cr0TDEK8_1),.clk(gclk));
	jdff dff_B_delF4Zas1_1(.din(w_dff_B_8Cr0TDEK8_1),.dout(w_dff_B_delF4Zas1_1),.clk(gclk));
	jdff dff_B_tbdtF29X5_1(.din(w_dff_B_delF4Zas1_1),.dout(w_dff_B_tbdtF29X5_1),.clk(gclk));
	jdff dff_B_shH6qQGn7_1(.din(w_dff_B_tbdtF29X5_1),.dout(w_dff_B_shH6qQGn7_1),.clk(gclk));
	jdff dff_B_RpVWgE2a6_1(.din(w_dff_B_shH6qQGn7_1),.dout(w_dff_B_RpVWgE2a6_1),.clk(gclk));
	jdff dff_B_hZ079ath5_1(.din(w_dff_B_RpVWgE2a6_1),.dout(w_dff_B_hZ079ath5_1),.clk(gclk));
	jdff dff_B_6VVkpMPZ1_1(.din(w_dff_B_hZ079ath5_1),.dout(w_dff_B_6VVkpMPZ1_1),.clk(gclk));
	jdff dff_B_hFiHPxHv8_1(.din(w_dff_B_6VVkpMPZ1_1),.dout(w_dff_B_hFiHPxHv8_1),.clk(gclk));
	jdff dff_B_faYWkUvB7_1(.din(w_dff_B_hFiHPxHv8_1),.dout(w_dff_B_faYWkUvB7_1),.clk(gclk));
	jdff dff_B_ncU3zyj54_1(.din(w_dff_B_faYWkUvB7_1),.dout(w_dff_B_ncU3zyj54_1),.clk(gclk));
	jdff dff_B_b47Ey68k6_1(.din(w_dff_B_ncU3zyj54_1),.dout(w_dff_B_b47Ey68k6_1),.clk(gclk));
	jdff dff_B_04oEdqq83_1(.din(w_dff_B_b47Ey68k6_1),.dout(w_dff_B_04oEdqq83_1),.clk(gclk));
	jdff dff_B_sYoD3wKb8_1(.din(w_dff_B_04oEdqq83_1),.dout(w_dff_B_sYoD3wKb8_1),.clk(gclk));
	jdff dff_B_U3ijMOQ21_1(.din(w_dff_B_sYoD3wKb8_1),.dout(w_dff_B_U3ijMOQ21_1),.clk(gclk));
	jdff dff_B_xuERZg8e0_1(.din(w_dff_B_U3ijMOQ21_1),.dout(w_dff_B_xuERZg8e0_1),.clk(gclk));
	jdff dff_B_C0aIYlpK2_1(.din(w_dff_B_xuERZg8e0_1),.dout(w_dff_B_C0aIYlpK2_1),.clk(gclk));
	jdff dff_B_AUKxi8sQ2_1(.din(w_dff_B_C0aIYlpK2_1),.dout(w_dff_B_AUKxi8sQ2_1),.clk(gclk));
	jdff dff_B_MkIcXSec5_1(.din(w_dff_B_AUKxi8sQ2_1),.dout(w_dff_B_MkIcXSec5_1),.clk(gclk));
	jdff dff_B_hLk0iwCI2_1(.din(w_dff_B_MkIcXSec5_1),.dout(w_dff_B_hLk0iwCI2_1),.clk(gclk));
	jdff dff_B_kAZSBhwF8_1(.din(w_dff_B_hLk0iwCI2_1),.dout(w_dff_B_kAZSBhwF8_1),.clk(gclk));
	jdff dff_B_car6Iadq0_1(.din(w_dff_B_kAZSBhwF8_1),.dout(w_dff_B_car6Iadq0_1),.clk(gclk));
	jdff dff_B_JQLYd7Gz9_1(.din(w_dff_B_car6Iadq0_1),.dout(w_dff_B_JQLYd7Gz9_1),.clk(gclk));
	jdff dff_B_6TxBxlq59_1(.din(w_dff_B_JQLYd7Gz9_1),.dout(w_dff_B_6TxBxlq59_1),.clk(gclk));
	jdff dff_B_8j8EdYPm6_1(.din(w_dff_B_6TxBxlq59_1),.dout(w_dff_B_8j8EdYPm6_1),.clk(gclk));
	jdff dff_B_eTmHU9F74_1(.din(w_dff_B_8j8EdYPm6_1),.dout(w_dff_B_eTmHU9F74_1),.clk(gclk));
	jdff dff_B_vdi7sNWe8_1(.din(w_dff_B_eTmHU9F74_1),.dout(w_dff_B_vdi7sNWe8_1),.clk(gclk));
	jdff dff_B_UVST5Psl6_1(.din(w_dff_B_vdi7sNWe8_1),.dout(w_dff_B_UVST5Psl6_1),.clk(gclk));
	jdff dff_B_sV5OFSWG8_1(.din(w_dff_B_UVST5Psl6_1),.dout(w_dff_B_sV5OFSWG8_1),.clk(gclk));
	jdff dff_B_TnQ11QdE6_1(.din(w_dff_B_sV5OFSWG8_1),.dout(w_dff_B_TnQ11QdE6_1),.clk(gclk));
	jdff dff_B_r7INjLgL2_1(.din(w_dff_B_TnQ11QdE6_1),.dout(w_dff_B_r7INjLgL2_1),.clk(gclk));
	jdff dff_B_Vf8B4GpP1_1(.din(w_dff_B_r7INjLgL2_1),.dout(w_dff_B_Vf8B4GpP1_1),.clk(gclk));
	jdff dff_B_hvlMPTQU4_1(.din(w_dff_B_Vf8B4GpP1_1),.dout(w_dff_B_hvlMPTQU4_1),.clk(gclk));
	jdff dff_B_o8Q9QmFf8_1(.din(w_dff_B_hvlMPTQU4_1),.dout(w_dff_B_o8Q9QmFf8_1),.clk(gclk));
	jdff dff_B_VyhL9ZbR7_1(.din(w_dff_B_o8Q9QmFf8_1),.dout(w_dff_B_VyhL9ZbR7_1),.clk(gclk));
	jdff dff_B_Vx6SkBpy5_1(.din(w_dff_B_VyhL9ZbR7_1),.dout(w_dff_B_Vx6SkBpy5_1),.clk(gclk));
	jdff dff_B_V3roUK6J2_1(.din(w_dff_B_Vx6SkBpy5_1),.dout(w_dff_B_V3roUK6J2_1),.clk(gclk));
	jdff dff_B_j0hqHtfN0_1(.din(w_dff_B_V3roUK6J2_1),.dout(w_dff_B_j0hqHtfN0_1),.clk(gclk));
	jdff dff_B_79PLedoF0_1(.din(w_dff_B_j0hqHtfN0_1),.dout(w_dff_B_79PLedoF0_1),.clk(gclk));
	jdff dff_B_IYp0UUHq6_1(.din(w_dff_B_79PLedoF0_1),.dout(w_dff_B_IYp0UUHq6_1),.clk(gclk));
	jdff dff_B_kANsNCpt4_1(.din(w_dff_B_IYp0UUHq6_1),.dout(w_dff_B_kANsNCpt4_1),.clk(gclk));
	jdff dff_B_7PPvMfFA7_1(.din(w_dff_B_kANsNCpt4_1),.dout(w_dff_B_7PPvMfFA7_1),.clk(gclk));
	jdff dff_B_I6WIoN6h9_0(.din(n799),.dout(w_dff_B_I6WIoN6h9_0),.clk(gclk));
	jdff dff_B_v20YfTkz6_0(.din(w_dff_B_I6WIoN6h9_0),.dout(w_dff_B_v20YfTkz6_0),.clk(gclk));
	jdff dff_B_PfraoEG97_0(.din(w_dff_B_v20YfTkz6_0),.dout(w_dff_B_PfraoEG97_0),.clk(gclk));
	jdff dff_B_imbyAO0c0_0(.din(w_dff_B_PfraoEG97_0),.dout(w_dff_B_imbyAO0c0_0),.clk(gclk));
	jdff dff_B_W1o7TQaN3_0(.din(w_dff_B_imbyAO0c0_0),.dout(w_dff_B_W1o7TQaN3_0),.clk(gclk));
	jdff dff_B_okqyDaim1_0(.din(w_dff_B_W1o7TQaN3_0),.dout(w_dff_B_okqyDaim1_0),.clk(gclk));
	jdff dff_B_OfCh70Dx4_0(.din(w_dff_B_okqyDaim1_0),.dout(w_dff_B_OfCh70Dx4_0),.clk(gclk));
	jdff dff_B_u4IfrlRY8_0(.din(w_dff_B_OfCh70Dx4_0),.dout(w_dff_B_u4IfrlRY8_0),.clk(gclk));
	jdff dff_B_tu2SQGoP4_0(.din(w_dff_B_u4IfrlRY8_0),.dout(w_dff_B_tu2SQGoP4_0),.clk(gclk));
	jdff dff_B_V96De1zx0_0(.din(w_dff_B_tu2SQGoP4_0),.dout(w_dff_B_V96De1zx0_0),.clk(gclk));
	jdff dff_B_6rRrfUwT2_0(.din(w_dff_B_V96De1zx0_0),.dout(w_dff_B_6rRrfUwT2_0),.clk(gclk));
	jdff dff_B_gleQx6wI2_0(.din(w_dff_B_6rRrfUwT2_0),.dout(w_dff_B_gleQx6wI2_0),.clk(gclk));
	jdff dff_B_qf9QqL4M3_0(.din(w_dff_B_gleQx6wI2_0),.dout(w_dff_B_qf9QqL4M3_0),.clk(gclk));
	jdff dff_B_mmjojyzO8_0(.din(w_dff_B_qf9QqL4M3_0),.dout(w_dff_B_mmjojyzO8_0),.clk(gclk));
	jdff dff_B_PUgkccG65_0(.din(w_dff_B_mmjojyzO8_0),.dout(w_dff_B_PUgkccG65_0),.clk(gclk));
	jdff dff_B_bzzPzEFh1_0(.din(w_dff_B_PUgkccG65_0),.dout(w_dff_B_bzzPzEFh1_0),.clk(gclk));
	jdff dff_B_LY3rvpL17_0(.din(w_dff_B_bzzPzEFh1_0),.dout(w_dff_B_LY3rvpL17_0),.clk(gclk));
	jdff dff_B_zQxkMZYt4_0(.din(w_dff_B_LY3rvpL17_0),.dout(w_dff_B_zQxkMZYt4_0),.clk(gclk));
	jdff dff_B_vtTpJuU04_0(.din(w_dff_B_zQxkMZYt4_0),.dout(w_dff_B_vtTpJuU04_0),.clk(gclk));
	jdff dff_B_AcgPGI5J9_0(.din(w_dff_B_vtTpJuU04_0),.dout(w_dff_B_AcgPGI5J9_0),.clk(gclk));
	jdff dff_B_3ISiST9S4_0(.din(w_dff_B_AcgPGI5J9_0),.dout(w_dff_B_3ISiST9S4_0),.clk(gclk));
	jdff dff_B_Hny5F13O7_0(.din(w_dff_B_3ISiST9S4_0),.dout(w_dff_B_Hny5F13O7_0),.clk(gclk));
	jdff dff_B_KoMGABHe1_0(.din(w_dff_B_Hny5F13O7_0),.dout(w_dff_B_KoMGABHe1_0),.clk(gclk));
	jdff dff_B_AYmvd9PC9_0(.din(w_dff_B_KoMGABHe1_0),.dout(w_dff_B_AYmvd9PC9_0),.clk(gclk));
	jdff dff_B_VTqx7xA56_0(.din(w_dff_B_AYmvd9PC9_0),.dout(w_dff_B_VTqx7xA56_0),.clk(gclk));
	jdff dff_B_jFSt2hhA9_0(.din(w_dff_B_VTqx7xA56_0),.dout(w_dff_B_jFSt2hhA9_0),.clk(gclk));
	jdff dff_B_2ElLLR002_0(.din(w_dff_B_jFSt2hhA9_0),.dout(w_dff_B_2ElLLR002_0),.clk(gclk));
	jdff dff_B_VBmHLkhk4_0(.din(w_dff_B_2ElLLR002_0),.dout(w_dff_B_VBmHLkhk4_0),.clk(gclk));
	jdff dff_B_uu8e0X9u2_0(.din(w_dff_B_VBmHLkhk4_0),.dout(w_dff_B_uu8e0X9u2_0),.clk(gclk));
	jdff dff_B_rxm1CEDV3_0(.din(w_dff_B_uu8e0X9u2_0),.dout(w_dff_B_rxm1CEDV3_0),.clk(gclk));
	jdff dff_B_POCj02fA0_0(.din(w_dff_B_rxm1CEDV3_0),.dout(w_dff_B_POCj02fA0_0),.clk(gclk));
	jdff dff_B_QZmL1ut17_0(.din(w_dff_B_POCj02fA0_0),.dout(w_dff_B_QZmL1ut17_0),.clk(gclk));
	jdff dff_B_is1RNg5Z7_0(.din(w_dff_B_QZmL1ut17_0),.dout(w_dff_B_is1RNg5Z7_0),.clk(gclk));
	jdff dff_B_F448UmfK5_0(.din(w_dff_B_is1RNg5Z7_0),.dout(w_dff_B_F448UmfK5_0),.clk(gclk));
	jdff dff_B_dYvtZ8Df4_0(.din(w_dff_B_F448UmfK5_0),.dout(w_dff_B_dYvtZ8Df4_0),.clk(gclk));
	jdff dff_B_Jlo8iZXm1_0(.din(w_dff_B_dYvtZ8Df4_0),.dout(w_dff_B_Jlo8iZXm1_0),.clk(gclk));
	jdff dff_B_1lD11DCz5_0(.din(w_dff_B_Jlo8iZXm1_0),.dout(w_dff_B_1lD11DCz5_0),.clk(gclk));
	jdff dff_B_X7lFK10V4_0(.din(w_dff_B_1lD11DCz5_0),.dout(w_dff_B_X7lFK10V4_0),.clk(gclk));
	jdff dff_B_ByIfzr0X7_0(.din(w_dff_B_X7lFK10V4_0),.dout(w_dff_B_ByIfzr0X7_0),.clk(gclk));
	jdff dff_B_IM7RNfKI9_0(.din(w_dff_B_ByIfzr0X7_0),.dout(w_dff_B_IM7RNfKI9_0),.clk(gclk));
	jdff dff_B_l25djXMi1_0(.din(w_dff_B_IM7RNfKI9_0),.dout(w_dff_B_l25djXMi1_0),.clk(gclk));
	jdff dff_B_NtXcXJe15_0(.din(w_dff_B_l25djXMi1_0),.dout(w_dff_B_NtXcXJe15_0),.clk(gclk));
	jdff dff_B_7tdbdGb58_0(.din(w_dff_B_NtXcXJe15_0),.dout(w_dff_B_7tdbdGb58_0),.clk(gclk));
	jdff dff_B_b3nx18Dx2_0(.din(w_dff_B_7tdbdGb58_0),.dout(w_dff_B_b3nx18Dx2_0),.clk(gclk));
	jdff dff_B_wSys2fMt6_0(.din(w_dff_B_b3nx18Dx2_0),.dout(w_dff_B_wSys2fMt6_0),.clk(gclk));
	jdff dff_B_RQiFxszD5_0(.din(w_dff_B_wSys2fMt6_0),.dout(w_dff_B_RQiFxszD5_0),.clk(gclk));
	jdff dff_B_TJy3hCGi0_0(.din(w_dff_B_RQiFxszD5_0),.dout(w_dff_B_TJy3hCGi0_0),.clk(gclk));
	jdff dff_B_QAVTeGs81_0(.din(w_dff_B_TJy3hCGi0_0),.dout(w_dff_B_QAVTeGs81_0),.clk(gclk));
	jdff dff_B_SHZTPkSY3_0(.din(w_dff_B_QAVTeGs81_0),.dout(w_dff_B_SHZTPkSY3_0),.clk(gclk));
	jdff dff_B_BVceaEl17_0(.din(w_dff_B_SHZTPkSY3_0),.dout(w_dff_B_BVceaEl17_0),.clk(gclk));
	jdff dff_B_oEZnnk893_0(.din(w_dff_B_BVceaEl17_0),.dout(w_dff_B_oEZnnk893_0),.clk(gclk));
	jdff dff_B_g2qzq5Uk0_0(.din(w_dff_B_oEZnnk893_0),.dout(w_dff_B_g2qzq5Uk0_0),.clk(gclk));
	jdff dff_B_pZ0wTiXF3_0(.din(w_dff_B_g2qzq5Uk0_0),.dout(w_dff_B_pZ0wTiXF3_0),.clk(gclk));
	jdff dff_B_pRlFmw680_0(.din(w_dff_B_pZ0wTiXF3_0),.dout(w_dff_B_pRlFmw680_0),.clk(gclk));
	jdff dff_B_PrE4Y01E3_0(.din(w_dff_B_pRlFmw680_0),.dout(w_dff_B_PrE4Y01E3_0),.clk(gclk));
	jdff dff_B_UPycdJTr5_0(.din(w_dff_B_PrE4Y01E3_0),.dout(w_dff_B_UPycdJTr5_0),.clk(gclk));
	jdff dff_B_REgZMpD55_0(.din(w_dff_B_UPycdJTr5_0),.dout(w_dff_B_REgZMpD55_0),.clk(gclk));
	jdff dff_B_kvaykdB33_0(.din(w_dff_B_REgZMpD55_0),.dout(w_dff_B_kvaykdB33_0),.clk(gclk));
	jdff dff_B_l5TD8cJi8_0(.din(w_dff_B_kvaykdB33_0),.dout(w_dff_B_l5TD8cJi8_0),.clk(gclk));
	jdff dff_B_bKY8m1741_0(.din(w_dff_B_l5TD8cJi8_0),.dout(w_dff_B_bKY8m1741_0),.clk(gclk));
	jdff dff_B_He72oM2c0_0(.din(w_dff_B_bKY8m1741_0),.dout(w_dff_B_He72oM2c0_0),.clk(gclk));
	jdff dff_B_1Nni3J8A7_0(.din(w_dff_B_He72oM2c0_0),.dout(w_dff_B_1Nni3J8A7_0),.clk(gclk));
	jdff dff_B_FQYrsurh4_0(.din(w_dff_B_1Nni3J8A7_0),.dout(w_dff_B_FQYrsurh4_0),.clk(gclk));
	jdff dff_B_IKOjdOM87_0(.din(w_dff_B_FQYrsurh4_0),.dout(w_dff_B_IKOjdOM87_0),.clk(gclk));
	jdff dff_B_paRCc5t83_0(.din(w_dff_B_IKOjdOM87_0),.dout(w_dff_B_paRCc5t83_0),.clk(gclk));
	jdff dff_B_RQgA9OTF1_0(.din(w_dff_B_paRCc5t83_0),.dout(w_dff_B_RQgA9OTF1_0),.clk(gclk));
	jdff dff_B_LscnLPzu1_0(.din(w_dff_B_RQgA9OTF1_0),.dout(w_dff_B_LscnLPzu1_0),.clk(gclk));
	jdff dff_B_ZVOHQZK42_0(.din(w_dff_B_LscnLPzu1_0),.dout(w_dff_B_ZVOHQZK42_0),.clk(gclk));
	jdff dff_B_iAHi3cHM6_0(.din(w_dff_B_ZVOHQZK42_0),.dout(w_dff_B_iAHi3cHM6_0),.clk(gclk));
	jdff dff_B_ccPsAbWf9_1(.din(n792),.dout(w_dff_B_ccPsAbWf9_1),.clk(gclk));
	jdff dff_B_dmbCAVom9_1(.din(w_dff_B_ccPsAbWf9_1),.dout(w_dff_B_dmbCAVom9_1),.clk(gclk));
	jdff dff_B_MgeQSUbk5_1(.din(w_dff_B_dmbCAVom9_1),.dout(w_dff_B_MgeQSUbk5_1),.clk(gclk));
	jdff dff_B_0DkQeKzB3_1(.din(w_dff_B_MgeQSUbk5_1),.dout(w_dff_B_0DkQeKzB3_1),.clk(gclk));
	jdff dff_B_24do6nwZ7_1(.din(w_dff_B_0DkQeKzB3_1),.dout(w_dff_B_24do6nwZ7_1),.clk(gclk));
	jdff dff_B_5CsvRKcR9_1(.din(w_dff_B_24do6nwZ7_1),.dout(w_dff_B_5CsvRKcR9_1),.clk(gclk));
	jdff dff_B_BwLXSL496_1(.din(w_dff_B_5CsvRKcR9_1),.dout(w_dff_B_BwLXSL496_1),.clk(gclk));
	jdff dff_B_X5SdyCPi4_1(.din(w_dff_B_BwLXSL496_1),.dout(w_dff_B_X5SdyCPi4_1),.clk(gclk));
	jdff dff_B_pBcaSdze7_1(.din(w_dff_B_X5SdyCPi4_1),.dout(w_dff_B_pBcaSdze7_1),.clk(gclk));
	jdff dff_B_oF7TpXhf2_1(.din(w_dff_B_pBcaSdze7_1),.dout(w_dff_B_oF7TpXhf2_1),.clk(gclk));
	jdff dff_B_0Jb9fXQB2_1(.din(w_dff_B_oF7TpXhf2_1),.dout(w_dff_B_0Jb9fXQB2_1),.clk(gclk));
	jdff dff_B_uMDf2A0X9_1(.din(w_dff_B_0Jb9fXQB2_1),.dout(w_dff_B_uMDf2A0X9_1),.clk(gclk));
	jdff dff_B_TgXIkbVz9_1(.din(w_dff_B_uMDf2A0X9_1),.dout(w_dff_B_TgXIkbVz9_1),.clk(gclk));
	jdff dff_B_bn0PNVvC9_1(.din(w_dff_B_TgXIkbVz9_1),.dout(w_dff_B_bn0PNVvC9_1),.clk(gclk));
	jdff dff_B_Rs4oPUVF0_1(.din(w_dff_B_bn0PNVvC9_1),.dout(w_dff_B_Rs4oPUVF0_1),.clk(gclk));
	jdff dff_B_FgAafpcG0_1(.din(w_dff_B_Rs4oPUVF0_1),.dout(w_dff_B_FgAafpcG0_1),.clk(gclk));
	jdff dff_B_UwaFiXc28_1(.din(w_dff_B_FgAafpcG0_1),.dout(w_dff_B_UwaFiXc28_1),.clk(gclk));
	jdff dff_B_gm5GmJDo1_1(.din(w_dff_B_UwaFiXc28_1),.dout(w_dff_B_gm5GmJDo1_1),.clk(gclk));
	jdff dff_B_bF6joxCt6_1(.din(w_dff_B_gm5GmJDo1_1),.dout(w_dff_B_bF6joxCt6_1),.clk(gclk));
	jdff dff_B_P5K6vhlN1_1(.din(w_dff_B_bF6joxCt6_1),.dout(w_dff_B_P5K6vhlN1_1),.clk(gclk));
	jdff dff_B_7ry2rKjK0_1(.din(w_dff_B_P5K6vhlN1_1),.dout(w_dff_B_7ry2rKjK0_1),.clk(gclk));
	jdff dff_B_lMzls0By5_1(.din(w_dff_B_7ry2rKjK0_1),.dout(w_dff_B_lMzls0By5_1),.clk(gclk));
	jdff dff_B_qtCAoueu8_1(.din(w_dff_B_lMzls0By5_1),.dout(w_dff_B_qtCAoueu8_1),.clk(gclk));
	jdff dff_B_nyelgwX72_1(.din(w_dff_B_qtCAoueu8_1),.dout(w_dff_B_nyelgwX72_1),.clk(gclk));
	jdff dff_B_RU54vTfO6_1(.din(w_dff_B_nyelgwX72_1),.dout(w_dff_B_RU54vTfO6_1),.clk(gclk));
	jdff dff_B_dhGlGXz38_1(.din(w_dff_B_RU54vTfO6_1),.dout(w_dff_B_dhGlGXz38_1),.clk(gclk));
	jdff dff_B_TJvcmoAJ6_1(.din(w_dff_B_dhGlGXz38_1),.dout(w_dff_B_TJvcmoAJ6_1),.clk(gclk));
	jdff dff_B_VGuaFH3C4_1(.din(w_dff_B_TJvcmoAJ6_1),.dout(w_dff_B_VGuaFH3C4_1),.clk(gclk));
	jdff dff_B_bCdNpNb82_1(.din(w_dff_B_VGuaFH3C4_1),.dout(w_dff_B_bCdNpNb82_1),.clk(gclk));
	jdff dff_B_cd4ZdLXE0_1(.din(w_dff_B_bCdNpNb82_1),.dout(w_dff_B_cd4ZdLXE0_1),.clk(gclk));
	jdff dff_B_gCWmVbHO2_1(.din(w_dff_B_cd4ZdLXE0_1),.dout(w_dff_B_gCWmVbHO2_1),.clk(gclk));
	jdff dff_B_uIH1LtwR0_1(.din(w_dff_B_gCWmVbHO2_1),.dout(w_dff_B_uIH1LtwR0_1),.clk(gclk));
	jdff dff_B_aBLe5VPw2_1(.din(w_dff_B_uIH1LtwR0_1),.dout(w_dff_B_aBLe5VPw2_1),.clk(gclk));
	jdff dff_B_Mew2iMBG1_1(.din(w_dff_B_aBLe5VPw2_1),.dout(w_dff_B_Mew2iMBG1_1),.clk(gclk));
	jdff dff_B_B1HOIyvz8_1(.din(w_dff_B_Mew2iMBG1_1),.dout(w_dff_B_B1HOIyvz8_1),.clk(gclk));
	jdff dff_B_x7a7HDjW2_1(.din(w_dff_B_B1HOIyvz8_1),.dout(w_dff_B_x7a7HDjW2_1),.clk(gclk));
	jdff dff_B_MVEgX4ZT6_1(.din(w_dff_B_x7a7HDjW2_1),.dout(w_dff_B_MVEgX4ZT6_1),.clk(gclk));
	jdff dff_B_X6gl0TC57_1(.din(w_dff_B_MVEgX4ZT6_1),.dout(w_dff_B_X6gl0TC57_1),.clk(gclk));
	jdff dff_B_RnXb8XwF7_1(.din(w_dff_B_X6gl0TC57_1),.dout(w_dff_B_RnXb8XwF7_1),.clk(gclk));
	jdff dff_B_WdejpLEj2_1(.din(w_dff_B_RnXb8XwF7_1),.dout(w_dff_B_WdejpLEj2_1),.clk(gclk));
	jdff dff_B_tGg6C0Gf2_1(.din(w_dff_B_WdejpLEj2_1),.dout(w_dff_B_tGg6C0Gf2_1),.clk(gclk));
	jdff dff_B_bYaLPosM8_1(.din(w_dff_B_tGg6C0Gf2_1),.dout(w_dff_B_bYaLPosM8_1),.clk(gclk));
	jdff dff_B_96qtvItC4_1(.din(w_dff_B_bYaLPosM8_1),.dout(w_dff_B_96qtvItC4_1),.clk(gclk));
	jdff dff_B_1DzZ794W0_1(.din(w_dff_B_96qtvItC4_1),.dout(w_dff_B_1DzZ794W0_1),.clk(gclk));
	jdff dff_B_V0YdEzAl6_1(.din(w_dff_B_1DzZ794W0_1),.dout(w_dff_B_V0YdEzAl6_1),.clk(gclk));
	jdff dff_B_u9Iyaxzs1_1(.din(w_dff_B_V0YdEzAl6_1),.dout(w_dff_B_u9Iyaxzs1_1),.clk(gclk));
	jdff dff_B_10iTyhZc8_1(.din(w_dff_B_u9Iyaxzs1_1),.dout(w_dff_B_10iTyhZc8_1),.clk(gclk));
	jdff dff_B_jQCpIzdn1_1(.din(w_dff_B_10iTyhZc8_1),.dout(w_dff_B_jQCpIzdn1_1),.clk(gclk));
	jdff dff_B_Y7qClh7w5_1(.din(w_dff_B_jQCpIzdn1_1),.dout(w_dff_B_Y7qClh7w5_1),.clk(gclk));
	jdff dff_B_Jl6hGn6p0_1(.din(w_dff_B_Y7qClh7w5_1),.dout(w_dff_B_Jl6hGn6p0_1),.clk(gclk));
	jdff dff_B_rXbfx66U8_1(.din(w_dff_B_Jl6hGn6p0_1),.dout(w_dff_B_rXbfx66U8_1),.clk(gclk));
	jdff dff_B_pnOqBFsZ5_1(.din(w_dff_B_rXbfx66U8_1),.dout(w_dff_B_pnOqBFsZ5_1),.clk(gclk));
	jdff dff_B_PfcHVto03_1(.din(w_dff_B_pnOqBFsZ5_1),.dout(w_dff_B_PfcHVto03_1),.clk(gclk));
	jdff dff_B_R5prVtWR3_1(.din(w_dff_B_PfcHVto03_1),.dout(w_dff_B_R5prVtWR3_1),.clk(gclk));
	jdff dff_B_g0FnvyOO0_1(.din(w_dff_B_R5prVtWR3_1),.dout(w_dff_B_g0FnvyOO0_1),.clk(gclk));
	jdff dff_B_X5WDxEki9_1(.din(w_dff_B_g0FnvyOO0_1),.dout(w_dff_B_X5WDxEki9_1),.clk(gclk));
	jdff dff_B_6rFnZItM8_1(.din(w_dff_B_X5WDxEki9_1),.dout(w_dff_B_6rFnZItM8_1),.clk(gclk));
	jdff dff_B_rVcEjktx8_1(.din(w_dff_B_6rFnZItM8_1),.dout(w_dff_B_rVcEjktx8_1),.clk(gclk));
	jdff dff_B_bZcmDoP90_1(.din(w_dff_B_rVcEjktx8_1),.dout(w_dff_B_bZcmDoP90_1),.clk(gclk));
	jdff dff_B_9yJEvkvp4_1(.din(w_dff_B_bZcmDoP90_1),.dout(w_dff_B_9yJEvkvp4_1),.clk(gclk));
	jdff dff_B_kbGi0tiY5_1(.din(w_dff_B_9yJEvkvp4_1),.dout(w_dff_B_kbGi0tiY5_1),.clk(gclk));
	jdff dff_B_qIt9bu6a7_1(.din(w_dff_B_kbGi0tiY5_1),.dout(w_dff_B_qIt9bu6a7_1),.clk(gclk));
	jdff dff_B_W5g0AisX0_1(.din(w_dff_B_qIt9bu6a7_1),.dout(w_dff_B_W5g0AisX0_1),.clk(gclk));
	jdff dff_B_uccJS0r33_1(.din(w_dff_B_W5g0AisX0_1),.dout(w_dff_B_uccJS0r33_1),.clk(gclk));
	jdff dff_B_zZI2lwkB3_1(.din(w_dff_B_uccJS0r33_1),.dout(w_dff_B_zZI2lwkB3_1),.clk(gclk));
	jdff dff_B_Q2rwYFRl1_1(.din(w_dff_B_zZI2lwkB3_1),.dout(w_dff_B_Q2rwYFRl1_1),.clk(gclk));
	jdff dff_B_uEErvOl90_1(.din(w_dff_B_Q2rwYFRl1_1),.dout(w_dff_B_uEErvOl90_1),.clk(gclk));
	jdff dff_B_qVRyJbno5_1(.din(w_dff_B_uEErvOl90_1),.dout(w_dff_B_qVRyJbno5_1),.clk(gclk));
	jdff dff_B_Z7Sirpij6_0(.din(n793),.dout(w_dff_B_Z7Sirpij6_0),.clk(gclk));
	jdff dff_B_Xt0IZgU98_0(.din(w_dff_B_Z7Sirpij6_0),.dout(w_dff_B_Xt0IZgU98_0),.clk(gclk));
	jdff dff_B_SscclUei3_0(.din(w_dff_B_Xt0IZgU98_0),.dout(w_dff_B_SscclUei3_0),.clk(gclk));
	jdff dff_B_06Ha8EZo0_0(.din(w_dff_B_SscclUei3_0),.dout(w_dff_B_06Ha8EZo0_0),.clk(gclk));
	jdff dff_B_rW9Os9Be3_0(.din(w_dff_B_06Ha8EZo0_0),.dout(w_dff_B_rW9Os9Be3_0),.clk(gclk));
	jdff dff_B_aLTFwZJy5_0(.din(w_dff_B_rW9Os9Be3_0),.dout(w_dff_B_aLTFwZJy5_0),.clk(gclk));
	jdff dff_B_tNkFvcdR8_0(.din(w_dff_B_aLTFwZJy5_0),.dout(w_dff_B_tNkFvcdR8_0),.clk(gclk));
	jdff dff_B_tcxaZwbW0_0(.din(w_dff_B_tNkFvcdR8_0),.dout(w_dff_B_tcxaZwbW0_0),.clk(gclk));
	jdff dff_B_Q4pd3c0U9_0(.din(w_dff_B_tcxaZwbW0_0),.dout(w_dff_B_Q4pd3c0U9_0),.clk(gclk));
	jdff dff_B_aEOuJAQW1_0(.din(w_dff_B_Q4pd3c0U9_0),.dout(w_dff_B_aEOuJAQW1_0),.clk(gclk));
	jdff dff_B_sXlyN3LW9_0(.din(w_dff_B_aEOuJAQW1_0),.dout(w_dff_B_sXlyN3LW9_0),.clk(gclk));
	jdff dff_B_ysnb1nD20_0(.din(w_dff_B_sXlyN3LW9_0),.dout(w_dff_B_ysnb1nD20_0),.clk(gclk));
	jdff dff_B_ZDo2W9112_0(.din(w_dff_B_ysnb1nD20_0),.dout(w_dff_B_ZDo2W9112_0),.clk(gclk));
	jdff dff_B_pH8Al40V3_0(.din(w_dff_B_ZDo2W9112_0),.dout(w_dff_B_pH8Al40V3_0),.clk(gclk));
	jdff dff_B_h3AyDBmA5_0(.din(w_dff_B_pH8Al40V3_0),.dout(w_dff_B_h3AyDBmA5_0),.clk(gclk));
	jdff dff_B_BTcpYFCC2_0(.din(w_dff_B_h3AyDBmA5_0),.dout(w_dff_B_BTcpYFCC2_0),.clk(gclk));
	jdff dff_B_2TLyYWgn4_0(.din(w_dff_B_BTcpYFCC2_0),.dout(w_dff_B_2TLyYWgn4_0),.clk(gclk));
	jdff dff_B_1PXVEvfi7_0(.din(w_dff_B_2TLyYWgn4_0),.dout(w_dff_B_1PXVEvfi7_0),.clk(gclk));
	jdff dff_B_j9uYYPGg2_0(.din(w_dff_B_1PXVEvfi7_0),.dout(w_dff_B_j9uYYPGg2_0),.clk(gclk));
	jdff dff_B_FMkCthkR8_0(.din(w_dff_B_j9uYYPGg2_0),.dout(w_dff_B_FMkCthkR8_0),.clk(gclk));
	jdff dff_B_OzMDdI7f5_0(.din(w_dff_B_FMkCthkR8_0),.dout(w_dff_B_OzMDdI7f5_0),.clk(gclk));
	jdff dff_B_B3Qfqtdn6_0(.din(w_dff_B_OzMDdI7f5_0),.dout(w_dff_B_B3Qfqtdn6_0),.clk(gclk));
	jdff dff_B_azkTL9Ge3_0(.din(w_dff_B_B3Qfqtdn6_0),.dout(w_dff_B_azkTL9Ge3_0),.clk(gclk));
	jdff dff_B_167uqdjx2_0(.din(w_dff_B_azkTL9Ge3_0),.dout(w_dff_B_167uqdjx2_0),.clk(gclk));
	jdff dff_B_pbofjOQ73_0(.din(w_dff_B_167uqdjx2_0),.dout(w_dff_B_pbofjOQ73_0),.clk(gclk));
	jdff dff_B_WBFFFfyu5_0(.din(w_dff_B_pbofjOQ73_0),.dout(w_dff_B_WBFFFfyu5_0),.clk(gclk));
	jdff dff_B_lSLEwKtG5_0(.din(w_dff_B_WBFFFfyu5_0),.dout(w_dff_B_lSLEwKtG5_0),.clk(gclk));
	jdff dff_B_in8KpmEK3_0(.din(w_dff_B_lSLEwKtG5_0),.dout(w_dff_B_in8KpmEK3_0),.clk(gclk));
	jdff dff_B_lpWVG82G3_0(.din(w_dff_B_in8KpmEK3_0),.dout(w_dff_B_lpWVG82G3_0),.clk(gclk));
	jdff dff_B_196kHsNn6_0(.din(w_dff_B_lpWVG82G3_0),.dout(w_dff_B_196kHsNn6_0),.clk(gclk));
	jdff dff_B_DaWn44x37_0(.din(w_dff_B_196kHsNn6_0),.dout(w_dff_B_DaWn44x37_0),.clk(gclk));
	jdff dff_B_ixTnrwlj0_0(.din(w_dff_B_DaWn44x37_0),.dout(w_dff_B_ixTnrwlj0_0),.clk(gclk));
	jdff dff_B_TZ6t1DcZ9_0(.din(w_dff_B_ixTnrwlj0_0),.dout(w_dff_B_TZ6t1DcZ9_0),.clk(gclk));
	jdff dff_B_73Eyf9sN5_0(.din(w_dff_B_TZ6t1DcZ9_0),.dout(w_dff_B_73Eyf9sN5_0),.clk(gclk));
	jdff dff_B_JUgVaWZe5_0(.din(w_dff_B_73Eyf9sN5_0),.dout(w_dff_B_JUgVaWZe5_0),.clk(gclk));
	jdff dff_B_HQt7KFSI4_0(.din(w_dff_B_JUgVaWZe5_0),.dout(w_dff_B_HQt7KFSI4_0),.clk(gclk));
	jdff dff_B_nljmBTFz4_0(.din(w_dff_B_HQt7KFSI4_0),.dout(w_dff_B_nljmBTFz4_0),.clk(gclk));
	jdff dff_B_XUqcbzYd3_0(.din(w_dff_B_nljmBTFz4_0),.dout(w_dff_B_XUqcbzYd3_0),.clk(gclk));
	jdff dff_B_qEBXuOTc1_0(.din(w_dff_B_XUqcbzYd3_0),.dout(w_dff_B_qEBXuOTc1_0),.clk(gclk));
	jdff dff_B_0IUP9tQc4_0(.din(w_dff_B_qEBXuOTc1_0),.dout(w_dff_B_0IUP9tQc4_0),.clk(gclk));
	jdff dff_B_1N6TIWUA9_0(.din(w_dff_B_0IUP9tQc4_0),.dout(w_dff_B_1N6TIWUA9_0),.clk(gclk));
	jdff dff_B_NqEojNv73_0(.din(w_dff_B_1N6TIWUA9_0),.dout(w_dff_B_NqEojNv73_0),.clk(gclk));
	jdff dff_B_dZXrFEHE3_0(.din(w_dff_B_NqEojNv73_0),.dout(w_dff_B_dZXrFEHE3_0),.clk(gclk));
	jdff dff_B_fquEqgDn0_0(.din(w_dff_B_dZXrFEHE3_0),.dout(w_dff_B_fquEqgDn0_0),.clk(gclk));
	jdff dff_B_NipIEUO12_0(.din(w_dff_B_fquEqgDn0_0),.dout(w_dff_B_NipIEUO12_0),.clk(gclk));
	jdff dff_B_H2nginmZ3_0(.din(w_dff_B_NipIEUO12_0),.dout(w_dff_B_H2nginmZ3_0),.clk(gclk));
	jdff dff_B_zNukDOmz4_0(.din(w_dff_B_H2nginmZ3_0),.dout(w_dff_B_zNukDOmz4_0),.clk(gclk));
	jdff dff_B_OcdQusVV4_0(.din(w_dff_B_zNukDOmz4_0),.dout(w_dff_B_OcdQusVV4_0),.clk(gclk));
	jdff dff_B_Z3I96UfL8_0(.din(w_dff_B_OcdQusVV4_0),.dout(w_dff_B_Z3I96UfL8_0),.clk(gclk));
	jdff dff_B_GR16x9f84_0(.din(w_dff_B_Z3I96UfL8_0),.dout(w_dff_B_GR16x9f84_0),.clk(gclk));
	jdff dff_B_YWVEAJNb3_0(.din(w_dff_B_GR16x9f84_0),.dout(w_dff_B_YWVEAJNb3_0),.clk(gclk));
	jdff dff_B_DTwAlIz35_0(.din(w_dff_B_YWVEAJNb3_0),.dout(w_dff_B_DTwAlIz35_0),.clk(gclk));
	jdff dff_B_pESVZrL72_0(.din(w_dff_B_DTwAlIz35_0),.dout(w_dff_B_pESVZrL72_0),.clk(gclk));
	jdff dff_B_oIGVC5e15_0(.din(w_dff_B_pESVZrL72_0),.dout(w_dff_B_oIGVC5e15_0),.clk(gclk));
	jdff dff_B_z9VmCxm43_0(.din(w_dff_B_oIGVC5e15_0),.dout(w_dff_B_z9VmCxm43_0),.clk(gclk));
	jdff dff_B_nAAcQ5dS9_0(.din(w_dff_B_z9VmCxm43_0),.dout(w_dff_B_nAAcQ5dS9_0),.clk(gclk));
	jdff dff_B_qBEN5rIH6_0(.din(w_dff_B_nAAcQ5dS9_0),.dout(w_dff_B_qBEN5rIH6_0),.clk(gclk));
	jdff dff_B_LdGie02W9_0(.din(w_dff_B_qBEN5rIH6_0),.dout(w_dff_B_LdGie02W9_0),.clk(gclk));
	jdff dff_B_q6hamDKF4_0(.din(w_dff_B_LdGie02W9_0),.dout(w_dff_B_q6hamDKF4_0),.clk(gclk));
	jdff dff_B_EWIV7aT86_0(.din(w_dff_B_q6hamDKF4_0),.dout(w_dff_B_EWIV7aT86_0),.clk(gclk));
	jdff dff_B_XgdVLFX05_0(.din(w_dff_B_EWIV7aT86_0),.dout(w_dff_B_XgdVLFX05_0),.clk(gclk));
	jdff dff_B_da93tegn2_0(.din(w_dff_B_XgdVLFX05_0),.dout(w_dff_B_da93tegn2_0),.clk(gclk));
	jdff dff_B_oTCFVaiB9_0(.din(w_dff_B_da93tegn2_0),.dout(w_dff_B_oTCFVaiB9_0),.clk(gclk));
	jdff dff_B_yN0uHUf27_0(.din(w_dff_B_oTCFVaiB9_0),.dout(w_dff_B_yN0uHUf27_0),.clk(gclk));
	jdff dff_B_Ql5QI0JW4_0(.din(w_dff_B_yN0uHUf27_0),.dout(w_dff_B_Ql5QI0JW4_0),.clk(gclk));
	jdff dff_B_4WKBwRrS5_0(.din(w_dff_B_Ql5QI0JW4_0),.dout(w_dff_B_4WKBwRrS5_0),.clk(gclk));
	jdff dff_B_jLpXYLo19_0(.din(w_dff_B_4WKBwRrS5_0),.dout(w_dff_B_jLpXYLo19_0),.clk(gclk));
	jdff dff_B_2OXQnYqp2_0(.din(w_dff_B_jLpXYLo19_0),.dout(w_dff_B_2OXQnYqp2_0),.clk(gclk));
	jdff dff_B_GYLbdOCX1_1(.din(n786),.dout(w_dff_B_GYLbdOCX1_1),.clk(gclk));
	jdff dff_B_XTMiRIhg6_1(.din(w_dff_B_GYLbdOCX1_1),.dout(w_dff_B_XTMiRIhg6_1),.clk(gclk));
	jdff dff_B_fca62qz78_1(.din(w_dff_B_XTMiRIhg6_1),.dout(w_dff_B_fca62qz78_1),.clk(gclk));
	jdff dff_B_CA96vvcK6_1(.din(w_dff_B_fca62qz78_1),.dout(w_dff_B_CA96vvcK6_1),.clk(gclk));
	jdff dff_B_AxC8Bn919_1(.din(w_dff_B_CA96vvcK6_1),.dout(w_dff_B_AxC8Bn919_1),.clk(gclk));
	jdff dff_B_VnGEQUVf8_1(.din(w_dff_B_AxC8Bn919_1),.dout(w_dff_B_VnGEQUVf8_1),.clk(gclk));
	jdff dff_B_gz805dBu9_1(.din(w_dff_B_VnGEQUVf8_1),.dout(w_dff_B_gz805dBu9_1),.clk(gclk));
	jdff dff_B_OYSgM1FI7_1(.din(w_dff_B_gz805dBu9_1),.dout(w_dff_B_OYSgM1FI7_1),.clk(gclk));
	jdff dff_B_kVgENUOB3_1(.din(w_dff_B_OYSgM1FI7_1),.dout(w_dff_B_kVgENUOB3_1),.clk(gclk));
	jdff dff_B_a5FLGmfM2_1(.din(w_dff_B_kVgENUOB3_1),.dout(w_dff_B_a5FLGmfM2_1),.clk(gclk));
	jdff dff_B_pudAD3l09_1(.din(w_dff_B_a5FLGmfM2_1),.dout(w_dff_B_pudAD3l09_1),.clk(gclk));
	jdff dff_B_Ry7mGxoA4_1(.din(w_dff_B_pudAD3l09_1),.dout(w_dff_B_Ry7mGxoA4_1),.clk(gclk));
	jdff dff_B_ayRfBUuD5_1(.din(w_dff_B_Ry7mGxoA4_1),.dout(w_dff_B_ayRfBUuD5_1),.clk(gclk));
	jdff dff_B_8TdiQmeR0_1(.din(w_dff_B_ayRfBUuD5_1),.dout(w_dff_B_8TdiQmeR0_1),.clk(gclk));
	jdff dff_B_15tzuv726_1(.din(w_dff_B_8TdiQmeR0_1),.dout(w_dff_B_15tzuv726_1),.clk(gclk));
	jdff dff_B_a4rhMODF8_1(.din(w_dff_B_15tzuv726_1),.dout(w_dff_B_a4rhMODF8_1),.clk(gclk));
	jdff dff_B_h5kncKbx2_1(.din(w_dff_B_a4rhMODF8_1),.dout(w_dff_B_h5kncKbx2_1),.clk(gclk));
	jdff dff_B_c7UWHLAU3_1(.din(w_dff_B_h5kncKbx2_1),.dout(w_dff_B_c7UWHLAU3_1),.clk(gclk));
	jdff dff_B_vK6RYFCF5_1(.din(w_dff_B_c7UWHLAU3_1),.dout(w_dff_B_vK6RYFCF5_1),.clk(gclk));
	jdff dff_B_dV7qbMGB7_1(.din(w_dff_B_vK6RYFCF5_1),.dout(w_dff_B_dV7qbMGB7_1),.clk(gclk));
	jdff dff_B_nIhwms0s2_1(.din(w_dff_B_dV7qbMGB7_1),.dout(w_dff_B_nIhwms0s2_1),.clk(gclk));
	jdff dff_B_5xgyrkik8_1(.din(w_dff_B_nIhwms0s2_1),.dout(w_dff_B_5xgyrkik8_1),.clk(gclk));
	jdff dff_B_kXpfZHYh6_1(.din(w_dff_B_5xgyrkik8_1),.dout(w_dff_B_kXpfZHYh6_1),.clk(gclk));
	jdff dff_B_P4D5bdzx3_1(.din(w_dff_B_kXpfZHYh6_1),.dout(w_dff_B_P4D5bdzx3_1),.clk(gclk));
	jdff dff_B_nbDHKJqV7_1(.din(w_dff_B_P4D5bdzx3_1),.dout(w_dff_B_nbDHKJqV7_1),.clk(gclk));
	jdff dff_B_VBapY2Xc5_1(.din(w_dff_B_nbDHKJqV7_1),.dout(w_dff_B_VBapY2Xc5_1),.clk(gclk));
	jdff dff_B_m3ahZ0hv3_1(.din(w_dff_B_VBapY2Xc5_1),.dout(w_dff_B_m3ahZ0hv3_1),.clk(gclk));
	jdff dff_B_npLZaldD7_1(.din(w_dff_B_m3ahZ0hv3_1),.dout(w_dff_B_npLZaldD7_1),.clk(gclk));
	jdff dff_B_rY1AjtU16_1(.din(w_dff_B_npLZaldD7_1),.dout(w_dff_B_rY1AjtU16_1),.clk(gclk));
	jdff dff_B_OB3r4e8T6_1(.din(w_dff_B_rY1AjtU16_1),.dout(w_dff_B_OB3r4e8T6_1),.clk(gclk));
	jdff dff_B_3EkqwtWF6_1(.din(w_dff_B_OB3r4e8T6_1),.dout(w_dff_B_3EkqwtWF6_1),.clk(gclk));
	jdff dff_B_FlCYy9XC2_1(.din(w_dff_B_3EkqwtWF6_1),.dout(w_dff_B_FlCYy9XC2_1),.clk(gclk));
	jdff dff_B_7WQkiWTC5_1(.din(w_dff_B_FlCYy9XC2_1),.dout(w_dff_B_7WQkiWTC5_1),.clk(gclk));
	jdff dff_B_ekxYldbM2_1(.din(w_dff_B_7WQkiWTC5_1),.dout(w_dff_B_ekxYldbM2_1),.clk(gclk));
	jdff dff_B_4nrSJw3b6_1(.din(w_dff_B_ekxYldbM2_1),.dout(w_dff_B_4nrSJw3b6_1),.clk(gclk));
	jdff dff_B_eSczoEVk3_1(.din(w_dff_B_4nrSJw3b6_1),.dout(w_dff_B_eSczoEVk3_1),.clk(gclk));
	jdff dff_B_VfiN7Kqr7_1(.din(w_dff_B_eSczoEVk3_1),.dout(w_dff_B_VfiN7Kqr7_1),.clk(gclk));
	jdff dff_B_yDWaDszt7_1(.din(w_dff_B_VfiN7Kqr7_1),.dout(w_dff_B_yDWaDszt7_1),.clk(gclk));
	jdff dff_B_KV7PT3no8_1(.din(w_dff_B_yDWaDszt7_1),.dout(w_dff_B_KV7PT3no8_1),.clk(gclk));
	jdff dff_B_Mamc8fYB6_1(.din(w_dff_B_KV7PT3no8_1),.dout(w_dff_B_Mamc8fYB6_1),.clk(gclk));
	jdff dff_B_R7fWHnxx9_1(.din(w_dff_B_Mamc8fYB6_1),.dout(w_dff_B_R7fWHnxx9_1),.clk(gclk));
	jdff dff_B_ebdebRnl0_1(.din(w_dff_B_R7fWHnxx9_1),.dout(w_dff_B_ebdebRnl0_1),.clk(gclk));
	jdff dff_B_IMkukUns7_1(.din(w_dff_B_ebdebRnl0_1),.dout(w_dff_B_IMkukUns7_1),.clk(gclk));
	jdff dff_B_BHFm5u7A9_1(.din(w_dff_B_IMkukUns7_1),.dout(w_dff_B_BHFm5u7A9_1),.clk(gclk));
	jdff dff_B_Fh8EvCGF5_1(.din(w_dff_B_BHFm5u7A9_1),.dout(w_dff_B_Fh8EvCGF5_1),.clk(gclk));
	jdff dff_B_aSirw5ni6_1(.din(w_dff_B_Fh8EvCGF5_1),.dout(w_dff_B_aSirw5ni6_1),.clk(gclk));
	jdff dff_B_MckXILbF5_1(.din(w_dff_B_aSirw5ni6_1),.dout(w_dff_B_MckXILbF5_1),.clk(gclk));
	jdff dff_B_7b54I00q0_1(.din(w_dff_B_MckXILbF5_1),.dout(w_dff_B_7b54I00q0_1),.clk(gclk));
	jdff dff_B_ew2uIHn05_1(.din(w_dff_B_7b54I00q0_1),.dout(w_dff_B_ew2uIHn05_1),.clk(gclk));
	jdff dff_B_E9YuMPL53_1(.din(w_dff_B_ew2uIHn05_1),.dout(w_dff_B_E9YuMPL53_1),.clk(gclk));
	jdff dff_B_JlnpJguO9_1(.din(w_dff_B_E9YuMPL53_1),.dout(w_dff_B_JlnpJguO9_1),.clk(gclk));
	jdff dff_B_t6xqW9AH7_1(.din(w_dff_B_JlnpJguO9_1),.dout(w_dff_B_t6xqW9AH7_1),.clk(gclk));
	jdff dff_B_GUvPEhZy4_1(.din(w_dff_B_t6xqW9AH7_1),.dout(w_dff_B_GUvPEhZy4_1),.clk(gclk));
	jdff dff_B_fKPjesXu7_1(.din(w_dff_B_GUvPEhZy4_1),.dout(w_dff_B_fKPjesXu7_1),.clk(gclk));
	jdff dff_B_QqPNInrF5_1(.din(w_dff_B_fKPjesXu7_1),.dout(w_dff_B_QqPNInrF5_1),.clk(gclk));
	jdff dff_B_9BafUZ3m2_1(.din(w_dff_B_QqPNInrF5_1),.dout(w_dff_B_9BafUZ3m2_1),.clk(gclk));
	jdff dff_B_r4FeSYkW5_1(.din(w_dff_B_9BafUZ3m2_1),.dout(w_dff_B_r4FeSYkW5_1),.clk(gclk));
	jdff dff_B_qqW4rb7h8_1(.din(w_dff_B_r4FeSYkW5_1),.dout(w_dff_B_qqW4rb7h8_1),.clk(gclk));
	jdff dff_B_bd0Chshm7_1(.din(w_dff_B_qqW4rb7h8_1),.dout(w_dff_B_bd0Chshm7_1),.clk(gclk));
	jdff dff_B_YNTY3V7G0_1(.din(w_dff_B_bd0Chshm7_1),.dout(w_dff_B_YNTY3V7G0_1),.clk(gclk));
	jdff dff_B_bFmVn5FG1_1(.din(w_dff_B_YNTY3V7G0_1),.dout(w_dff_B_bFmVn5FG1_1),.clk(gclk));
	jdff dff_B_mfpjVyzb5_1(.din(w_dff_B_bFmVn5FG1_1),.dout(w_dff_B_mfpjVyzb5_1),.clk(gclk));
	jdff dff_B_Hqpq0lHO1_1(.din(w_dff_B_mfpjVyzb5_1),.dout(w_dff_B_Hqpq0lHO1_1),.clk(gclk));
	jdff dff_B_q8PTZoPo1_1(.din(w_dff_B_Hqpq0lHO1_1),.dout(w_dff_B_q8PTZoPo1_1),.clk(gclk));
	jdff dff_B_webqAdQe2_1(.din(w_dff_B_q8PTZoPo1_1),.dout(w_dff_B_webqAdQe2_1),.clk(gclk));
	jdff dff_B_xE1QwoiX4_1(.din(w_dff_B_webqAdQe2_1),.dout(w_dff_B_xE1QwoiX4_1),.clk(gclk));
	jdff dff_B_cSmyQJfw1_1(.din(w_dff_B_xE1QwoiX4_1),.dout(w_dff_B_cSmyQJfw1_1),.clk(gclk));
	jdff dff_B_2kuov4Ma5_0(.din(n787),.dout(w_dff_B_2kuov4Ma5_0),.clk(gclk));
	jdff dff_B_hgcS7yAr1_0(.din(w_dff_B_2kuov4Ma5_0),.dout(w_dff_B_hgcS7yAr1_0),.clk(gclk));
	jdff dff_B_VFTWXQwn3_0(.din(w_dff_B_hgcS7yAr1_0),.dout(w_dff_B_VFTWXQwn3_0),.clk(gclk));
	jdff dff_B_IyIOkS585_0(.din(w_dff_B_VFTWXQwn3_0),.dout(w_dff_B_IyIOkS585_0),.clk(gclk));
	jdff dff_B_J5TPWZ5A2_0(.din(w_dff_B_IyIOkS585_0),.dout(w_dff_B_J5TPWZ5A2_0),.clk(gclk));
	jdff dff_B_xpa1SDpE3_0(.din(w_dff_B_J5TPWZ5A2_0),.dout(w_dff_B_xpa1SDpE3_0),.clk(gclk));
	jdff dff_B_MEZD3l295_0(.din(w_dff_B_xpa1SDpE3_0),.dout(w_dff_B_MEZD3l295_0),.clk(gclk));
	jdff dff_B_pMjUpsoh0_0(.din(w_dff_B_MEZD3l295_0),.dout(w_dff_B_pMjUpsoh0_0),.clk(gclk));
	jdff dff_B_eCCIluiV0_0(.din(w_dff_B_pMjUpsoh0_0),.dout(w_dff_B_eCCIluiV0_0),.clk(gclk));
	jdff dff_B_JcJcVjnT0_0(.din(w_dff_B_eCCIluiV0_0),.dout(w_dff_B_JcJcVjnT0_0),.clk(gclk));
	jdff dff_B_Y3F6E1Cv9_0(.din(w_dff_B_JcJcVjnT0_0),.dout(w_dff_B_Y3F6E1Cv9_0),.clk(gclk));
	jdff dff_B_aUYGUOPZ0_0(.din(w_dff_B_Y3F6E1Cv9_0),.dout(w_dff_B_aUYGUOPZ0_0),.clk(gclk));
	jdff dff_B_tmivuLWk9_0(.din(w_dff_B_aUYGUOPZ0_0),.dout(w_dff_B_tmivuLWk9_0),.clk(gclk));
	jdff dff_B_JHQmj32y2_0(.din(w_dff_B_tmivuLWk9_0),.dout(w_dff_B_JHQmj32y2_0),.clk(gclk));
	jdff dff_B_x6STL4N87_0(.din(w_dff_B_JHQmj32y2_0),.dout(w_dff_B_x6STL4N87_0),.clk(gclk));
	jdff dff_B_f79Gd9jy3_0(.din(w_dff_B_x6STL4N87_0),.dout(w_dff_B_f79Gd9jy3_0),.clk(gclk));
	jdff dff_B_nT9Ppg2E5_0(.din(w_dff_B_f79Gd9jy3_0),.dout(w_dff_B_nT9Ppg2E5_0),.clk(gclk));
	jdff dff_B_g4wSRRW03_0(.din(w_dff_B_nT9Ppg2E5_0),.dout(w_dff_B_g4wSRRW03_0),.clk(gclk));
	jdff dff_B_vcQEEfC96_0(.din(w_dff_B_g4wSRRW03_0),.dout(w_dff_B_vcQEEfC96_0),.clk(gclk));
	jdff dff_B_X1PT3bfU4_0(.din(w_dff_B_vcQEEfC96_0),.dout(w_dff_B_X1PT3bfU4_0),.clk(gclk));
	jdff dff_B_zOmvvbsf7_0(.din(w_dff_B_X1PT3bfU4_0),.dout(w_dff_B_zOmvvbsf7_0),.clk(gclk));
	jdff dff_B_pa1ivYoB2_0(.din(w_dff_B_zOmvvbsf7_0),.dout(w_dff_B_pa1ivYoB2_0),.clk(gclk));
	jdff dff_B_gNrW1Hqd8_0(.din(w_dff_B_pa1ivYoB2_0),.dout(w_dff_B_gNrW1Hqd8_0),.clk(gclk));
	jdff dff_B_VCz6KMAP0_0(.din(w_dff_B_gNrW1Hqd8_0),.dout(w_dff_B_VCz6KMAP0_0),.clk(gclk));
	jdff dff_B_LIMABhSd5_0(.din(w_dff_B_VCz6KMAP0_0),.dout(w_dff_B_LIMABhSd5_0),.clk(gclk));
	jdff dff_B_vzyPKbW73_0(.din(w_dff_B_LIMABhSd5_0),.dout(w_dff_B_vzyPKbW73_0),.clk(gclk));
	jdff dff_B_imAPqwS29_0(.din(w_dff_B_vzyPKbW73_0),.dout(w_dff_B_imAPqwS29_0),.clk(gclk));
	jdff dff_B_bNVQeznS5_0(.din(w_dff_B_imAPqwS29_0),.dout(w_dff_B_bNVQeznS5_0),.clk(gclk));
	jdff dff_B_LXjMrRfl1_0(.din(w_dff_B_bNVQeznS5_0),.dout(w_dff_B_LXjMrRfl1_0),.clk(gclk));
	jdff dff_B_4GDqU3Y27_0(.din(w_dff_B_LXjMrRfl1_0),.dout(w_dff_B_4GDqU3Y27_0),.clk(gclk));
	jdff dff_B_L6Md8L6y4_0(.din(w_dff_B_4GDqU3Y27_0),.dout(w_dff_B_L6Md8L6y4_0),.clk(gclk));
	jdff dff_B_1JB8yVNP5_0(.din(w_dff_B_L6Md8L6y4_0),.dout(w_dff_B_1JB8yVNP5_0),.clk(gclk));
	jdff dff_B_gj84PKrv2_0(.din(w_dff_B_1JB8yVNP5_0),.dout(w_dff_B_gj84PKrv2_0),.clk(gclk));
	jdff dff_B_WTAsiURZ6_0(.din(w_dff_B_gj84PKrv2_0),.dout(w_dff_B_WTAsiURZ6_0),.clk(gclk));
	jdff dff_B_GqDHW8ku9_0(.din(w_dff_B_WTAsiURZ6_0),.dout(w_dff_B_GqDHW8ku9_0),.clk(gclk));
	jdff dff_B_arDvEw2o7_0(.din(w_dff_B_GqDHW8ku9_0),.dout(w_dff_B_arDvEw2o7_0),.clk(gclk));
	jdff dff_B_9O6ALU7A7_0(.din(w_dff_B_arDvEw2o7_0),.dout(w_dff_B_9O6ALU7A7_0),.clk(gclk));
	jdff dff_B_AyMsjAM11_0(.din(w_dff_B_9O6ALU7A7_0),.dout(w_dff_B_AyMsjAM11_0),.clk(gclk));
	jdff dff_B_kSiyrEyt6_0(.din(w_dff_B_AyMsjAM11_0),.dout(w_dff_B_kSiyrEyt6_0),.clk(gclk));
	jdff dff_B_nYpzzvIZ5_0(.din(w_dff_B_kSiyrEyt6_0),.dout(w_dff_B_nYpzzvIZ5_0),.clk(gclk));
	jdff dff_B_BTwfQMWg4_0(.din(w_dff_B_nYpzzvIZ5_0),.dout(w_dff_B_BTwfQMWg4_0),.clk(gclk));
	jdff dff_B_HcS9eDNk2_0(.din(w_dff_B_BTwfQMWg4_0),.dout(w_dff_B_HcS9eDNk2_0),.clk(gclk));
	jdff dff_B_bfB4mSgk7_0(.din(w_dff_B_HcS9eDNk2_0),.dout(w_dff_B_bfB4mSgk7_0),.clk(gclk));
	jdff dff_B_zqzTntQx4_0(.din(w_dff_B_bfB4mSgk7_0),.dout(w_dff_B_zqzTntQx4_0),.clk(gclk));
	jdff dff_B_BPyDJHz75_0(.din(w_dff_B_zqzTntQx4_0),.dout(w_dff_B_BPyDJHz75_0),.clk(gclk));
	jdff dff_B_Zy20p5QQ9_0(.din(w_dff_B_BPyDJHz75_0),.dout(w_dff_B_Zy20p5QQ9_0),.clk(gclk));
	jdff dff_B_78wEVBwe5_0(.din(w_dff_B_Zy20p5QQ9_0),.dout(w_dff_B_78wEVBwe5_0),.clk(gclk));
	jdff dff_B_olI84OtP1_0(.din(w_dff_B_78wEVBwe5_0),.dout(w_dff_B_olI84OtP1_0),.clk(gclk));
	jdff dff_B_mAjfHW8s2_0(.din(w_dff_B_olI84OtP1_0),.dout(w_dff_B_mAjfHW8s2_0),.clk(gclk));
	jdff dff_B_IJube8Tl3_0(.din(w_dff_B_mAjfHW8s2_0),.dout(w_dff_B_IJube8Tl3_0),.clk(gclk));
	jdff dff_B_bLRExcag1_0(.din(w_dff_B_IJube8Tl3_0),.dout(w_dff_B_bLRExcag1_0),.clk(gclk));
	jdff dff_B_otck3mYW7_0(.din(w_dff_B_bLRExcag1_0),.dout(w_dff_B_otck3mYW7_0),.clk(gclk));
	jdff dff_B_OW0lfqG68_0(.din(w_dff_B_otck3mYW7_0),.dout(w_dff_B_OW0lfqG68_0),.clk(gclk));
	jdff dff_B_KLDZkxPv9_0(.din(w_dff_B_OW0lfqG68_0),.dout(w_dff_B_KLDZkxPv9_0),.clk(gclk));
	jdff dff_B_0ioHCZkX2_0(.din(w_dff_B_KLDZkxPv9_0),.dout(w_dff_B_0ioHCZkX2_0),.clk(gclk));
	jdff dff_B_8wWhhm1t0_0(.din(w_dff_B_0ioHCZkX2_0),.dout(w_dff_B_8wWhhm1t0_0),.clk(gclk));
	jdff dff_B_Ye7Ynpi14_0(.din(w_dff_B_8wWhhm1t0_0),.dout(w_dff_B_Ye7Ynpi14_0),.clk(gclk));
	jdff dff_B_4OiEwAw81_0(.din(w_dff_B_Ye7Ynpi14_0),.dout(w_dff_B_4OiEwAw81_0),.clk(gclk));
	jdff dff_B_tCwxgcz61_0(.din(w_dff_B_4OiEwAw81_0),.dout(w_dff_B_tCwxgcz61_0),.clk(gclk));
	jdff dff_B_n8ypLifR2_0(.din(w_dff_B_tCwxgcz61_0),.dout(w_dff_B_n8ypLifR2_0),.clk(gclk));
	jdff dff_B_9f3vnqCZ2_0(.din(w_dff_B_n8ypLifR2_0),.dout(w_dff_B_9f3vnqCZ2_0),.clk(gclk));
	jdff dff_B_q22xhbRt6_0(.din(w_dff_B_9f3vnqCZ2_0),.dout(w_dff_B_q22xhbRt6_0),.clk(gclk));
	jdff dff_B_8bx1wEvl6_0(.din(w_dff_B_q22xhbRt6_0),.dout(w_dff_B_8bx1wEvl6_0),.clk(gclk));
	jdff dff_B_Ok9Fv8JV6_0(.din(w_dff_B_8bx1wEvl6_0),.dout(w_dff_B_Ok9Fv8JV6_0),.clk(gclk));
	jdff dff_B_SAdbhHjd5_0(.din(w_dff_B_Ok9Fv8JV6_0),.dout(w_dff_B_SAdbhHjd5_0),.clk(gclk));
	jdff dff_B_K3XBmhG19_0(.din(w_dff_B_SAdbhHjd5_0),.dout(w_dff_B_K3XBmhG19_0),.clk(gclk));
	jdff dff_B_bDbh5nUT3_0(.din(w_dff_B_K3XBmhG19_0),.dout(w_dff_B_bDbh5nUT3_0),.clk(gclk));
	jdff dff_B_56bX8R0X1_1(.din(n780),.dout(w_dff_B_56bX8R0X1_1),.clk(gclk));
	jdff dff_B_J1VBtjpb7_1(.din(w_dff_B_56bX8R0X1_1),.dout(w_dff_B_J1VBtjpb7_1),.clk(gclk));
	jdff dff_B_kT8blCOC1_1(.din(w_dff_B_J1VBtjpb7_1),.dout(w_dff_B_kT8blCOC1_1),.clk(gclk));
	jdff dff_B_TSzDlOlD2_1(.din(w_dff_B_kT8blCOC1_1),.dout(w_dff_B_TSzDlOlD2_1),.clk(gclk));
	jdff dff_B_mONv6dmT2_1(.din(w_dff_B_TSzDlOlD2_1),.dout(w_dff_B_mONv6dmT2_1),.clk(gclk));
	jdff dff_B_zpmgjFJA0_1(.din(w_dff_B_mONv6dmT2_1),.dout(w_dff_B_zpmgjFJA0_1),.clk(gclk));
	jdff dff_B_tOzNchBf7_1(.din(w_dff_B_zpmgjFJA0_1),.dout(w_dff_B_tOzNchBf7_1),.clk(gclk));
	jdff dff_B_McKFDm483_1(.din(w_dff_B_tOzNchBf7_1),.dout(w_dff_B_McKFDm483_1),.clk(gclk));
	jdff dff_B_kN4zv8fZ9_1(.din(w_dff_B_McKFDm483_1),.dout(w_dff_B_kN4zv8fZ9_1),.clk(gclk));
	jdff dff_B_lkp6yAJk8_1(.din(w_dff_B_kN4zv8fZ9_1),.dout(w_dff_B_lkp6yAJk8_1),.clk(gclk));
	jdff dff_B_Kx9gPkVX2_1(.din(w_dff_B_lkp6yAJk8_1),.dout(w_dff_B_Kx9gPkVX2_1),.clk(gclk));
	jdff dff_B_knTFINpX0_1(.din(w_dff_B_Kx9gPkVX2_1),.dout(w_dff_B_knTFINpX0_1),.clk(gclk));
	jdff dff_B_BdKWTzfq3_1(.din(w_dff_B_knTFINpX0_1),.dout(w_dff_B_BdKWTzfq3_1),.clk(gclk));
	jdff dff_B_ue7wsvFG8_1(.din(w_dff_B_BdKWTzfq3_1),.dout(w_dff_B_ue7wsvFG8_1),.clk(gclk));
	jdff dff_B_9ZMM5I1P3_1(.din(w_dff_B_ue7wsvFG8_1),.dout(w_dff_B_9ZMM5I1P3_1),.clk(gclk));
	jdff dff_B_Btqj4csN3_1(.din(w_dff_B_9ZMM5I1P3_1),.dout(w_dff_B_Btqj4csN3_1),.clk(gclk));
	jdff dff_B_FuXT22V75_1(.din(w_dff_B_Btqj4csN3_1),.dout(w_dff_B_FuXT22V75_1),.clk(gclk));
	jdff dff_B_9XYUF4Y51_1(.din(w_dff_B_FuXT22V75_1),.dout(w_dff_B_9XYUF4Y51_1),.clk(gclk));
	jdff dff_B_7fcbPlL34_1(.din(w_dff_B_9XYUF4Y51_1),.dout(w_dff_B_7fcbPlL34_1),.clk(gclk));
	jdff dff_B_KbrJpvMN9_1(.din(w_dff_B_7fcbPlL34_1),.dout(w_dff_B_KbrJpvMN9_1),.clk(gclk));
	jdff dff_B_wHeGzfyO0_1(.din(w_dff_B_KbrJpvMN9_1),.dout(w_dff_B_wHeGzfyO0_1),.clk(gclk));
	jdff dff_B_rbCrlYIc2_1(.din(w_dff_B_wHeGzfyO0_1),.dout(w_dff_B_rbCrlYIc2_1),.clk(gclk));
	jdff dff_B_XlYlYdku0_1(.din(w_dff_B_rbCrlYIc2_1),.dout(w_dff_B_XlYlYdku0_1),.clk(gclk));
	jdff dff_B_LU0eBLHF4_1(.din(w_dff_B_XlYlYdku0_1),.dout(w_dff_B_LU0eBLHF4_1),.clk(gclk));
	jdff dff_B_9KSkMU2o8_1(.din(w_dff_B_LU0eBLHF4_1),.dout(w_dff_B_9KSkMU2o8_1),.clk(gclk));
	jdff dff_B_wt0LdzhI8_1(.din(w_dff_B_9KSkMU2o8_1),.dout(w_dff_B_wt0LdzhI8_1),.clk(gclk));
	jdff dff_B_G8hwBcFe3_1(.din(w_dff_B_wt0LdzhI8_1),.dout(w_dff_B_G8hwBcFe3_1),.clk(gclk));
	jdff dff_B_Berkjg9t1_1(.din(w_dff_B_G8hwBcFe3_1),.dout(w_dff_B_Berkjg9t1_1),.clk(gclk));
	jdff dff_B_7Rl9qeDe3_1(.din(w_dff_B_Berkjg9t1_1),.dout(w_dff_B_7Rl9qeDe3_1),.clk(gclk));
	jdff dff_B_EuE4d9l20_1(.din(w_dff_B_7Rl9qeDe3_1),.dout(w_dff_B_EuE4d9l20_1),.clk(gclk));
	jdff dff_B_NYdYAMfg2_1(.din(w_dff_B_EuE4d9l20_1),.dout(w_dff_B_NYdYAMfg2_1),.clk(gclk));
	jdff dff_B_SJoVikYW5_1(.din(w_dff_B_NYdYAMfg2_1),.dout(w_dff_B_SJoVikYW5_1),.clk(gclk));
	jdff dff_B_q6GBacby4_1(.din(w_dff_B_SJoVikYW5_1),.dout(w_dff_B_q6GBacby4_1),.clk(gclk));
	jdff dff_B_JrXM8Gur7_1(.din(w_dff_B_q6GBacby4_1),.dout(w_dff_B_JrXM8Gur7_1),.clk(gclk));
	jdff dff_B_srMCdosz4_1(.din(w_dff_B_JrXM8Gur7_1),.dout(w_dff_B_srMCdosz4_1),.clk(gclk));
	jdff dff_B_4hKse7bY4_1(.din(w_dff_B_srMCdosz4_1),.dout(w_dff_B_4hKse7bY4_1),.clk(gclk));
	jdff dff_B_TFs6LkqF2_1(.din(w_dff_B_4hKse7bY4_1),.dout(w_dff_B_TFs6LkqF2_1),.clk(gclk));
	jdff dff_B_go67H1jV6_1(.din(w_dff_B_TFs6LkqF2_1),.dout(w_dff_B_go67H1jV6_1),.clk(gclk));
	jdff dff_B_c3DWREm90_1(.din(w_dff_B_go67H1jV6_1),.dout(w_dff_B_c3DWREm90_1),.clk(gclk));
	jdff dff_B_wcaO8rLs8_1(.din(w_dff_B_c3DWREm90_1),.dout(w_dff_B_wcaO8rLs8_1),.clk(gclk));
	jdff dff_B_Goglo8i51_1(.din(w_dff_B_wcaO8rLs8_1),.dout(w_dff_B_Goglo8i51_1),.clk(gclk));
	jdff dff_B_gxgFigMS6_1(.din(w_dff_B_Goglo8i51_1),.dout(w_dff_B_gxgFigMS6_1),.clk(gclk));
	jdff dff_B_1MknRRtB0_1(.din(w_dff_B_gxgFigMS6_1),.dout(w_dff_B_1MknRRtB0_1),.clk(gclk));
	jdff dff_B_FYp2ifzv6_1(.din(w_dff_B_1MknRRtB0_1),.dout(w_dff_B_FYp2ifzv6_1),.clk(gclk));
	jdff dff_B_tBEhIhY80_1(.din(w_dff_B_FYp2ifzv6_1),.dout(w_dff_B_tBEhIhY80_1),.clk(gclk));
	jdff dff_B_URwioq5W9_1(.din(w_dff_B_tBEhIhY80_1),.dout(w_dff_B_URwioq5W9_1),.clk(gclk));
	jdff dff_B_rH3K16z08_1(.din(w_dff_B_URwioq5W9_1),.dout(w_dff_B_rH3K16z08_1),.clk(gclk));
	jdff dff_B_Z4XxR2Vj7_1(.din(w_dff_B_rH3K16z08_1),.dout(w_dff_B_Z4XxR2Vj7_1),.clk(gclk));
	jdff dff_B_POg0RIHh7_1(.din(w_dff_B_Z4XxR2Vj7_1),.dout(w_dff_B_POg0RIHh7_1),.clk(gclk));
	jdff dff_B_pB6jNztE3_1(.din(w_dff_B_POg0RIHh7_1),.dout(w_dff_B_pB6jNztE3_1),.clk(gclk));
	jdff dff_B_gAWATq4q7_1(.din(w_dff_B_pB6jNztE3_1),.dout(w_dff_B_gAWATq4q7_1),.clk(gclk));
	jdff dff_B_zmDSTPOg8_1(.din(w_dff_B_gAWATq4q7_1),.dout(w_dff_B_zmDSTPOg8_1),.clk(gclk));
	jdff dff_B_7HZk2J4Z2_1(.din(w_dff_B_zmDSTPOg8_1),.dout(w_dff_B_7HZk2J4Z2_1),.clk(gclk));
	jdff dff_B_x19aOJ4G4_1(.din(w_dff_B_7HZk2J4Z2_1),.dout(w_dff_B_x19aOJ4G4_1),.clk(gclk));
	jdff dff_B_7YOlw7Rq5_1(.din(w_dff_B_x19aOJ4G4_1),.dout(w_dff_B_7YOlw7Rq5_1),.clk(gclk));
	jdff dff_B_rADkxrbZ0_1(.din(w_dff_B_7YOlw7Rq5_1),.dout(w_dff_B_rADkxrbZ0_1),.clk(gclk));
	jdff dff_B_xvXgV9UQ2_1(.din(w_dff_B_rADkxrbZ0_1),.dout(w_dff_B_xvXgV9UQ2_1),.clk(gclk));
	jdff dff_B_CrMqGhrX5_1(.din(w_dff_B_xvXgV9UQ2_1),.dout(w_dff_B_CrMqGhrX5_1),.clk(gclk));
	jdff dff_B_tazpeA5A9_1(.din(w_dff_B_CrMqGhrX5_1),.dout(w_dff_B_tazpeA5A9_1),.clk(gclk));
	jdff dff_B_3mG95Zq31_1(.din(w_dff_B_tazpeA5A9_1),.dout(w_dff_B_3mG95Zq31_1),.clk(gclk));
	jdff dff_B_VeAwDMtq4_1(.din(w_dff_B_3mG95Zq31_1),.dout(w_dff_B_VeAwDMtq4_1),.clk(gclk));
	jdff dff_B_qzF6vHka3_1(.din(w_dff_B_VeAwDMtq4_1),.dout(w_dff_B_qzF6vHka3_1),.clk(gclk));
	jdff dff_B_CX5qG5KJ2_1(.din(w_dff_B_qzF6vHka3_1),.dout(w_dff_B_CX5qG5KJ2_1),.clk(gclk));
	jdff dff_B_jT6bcSwr0_1(.din(w_dff_B_CX5qG5KJ2_1),.dout(w_dff_B_jT6bcSwr0_1),.clk(gclk));
	jdff dff_B_0jkwT1wb5_1(.din(w_dff_B_jT6bcSwr0_1),.dout(w_dff_B_0jkwT1wb5_1),.clk(gclk));
	jdff dff_B_SvQrjUup5_1(.din(w_dff_B_0jkwT1wb5_1),.dout(w_dff_B_SvQrjUup5_1),.clk(gclk));
	jdff dff_B_lC8L2YxA4_0(.din(n781),.dout(w_dff_B_lC8L2YxA4_0),.clk(gclk));
	jdff dff_B_UPgIhrhr4_0(.din(w_dff_B_lC8L2YxA4_0),.dout(w_dff_B_UPgIhrhr4_0),.clk(gclk));
	jdff dff_B_51ulyRTI6_0(.din(w_dff_B_UPgIhrhr4_0),.dout(w_dff_B_51ulyRTI6_0),.clk(gclk));
	jdff dff_B_IQ0VR6wP1_0(.din(w_dff_B_51ulyRTI6_0),.dout(w_dff_B_IQ0VR6wP1_0),.clk(gclk));
	jdff dff_B_ZjGJvPSI4_0(.din(w_dff_B_IQ0VR6wP1_0),.dout(w_dff_B_ZjGJvPSI4_0),.clk(gclk));
	jdff dff_B_tvqjYEwZ2_0(.din(w_dff_B_ZjGJvPSI4_0),.dout(w_dff_B_tvqjYEwZ2_0),.clk(gclk));
	jdff dff_B_Le8Canjh3_0(.din(w_dff_B_tvqjYEwZ2_0),.dout(w_dff_B_Le8Canjh3_0),.clk(gclk));
	jdff dff_B_lhdOWkJI7_0(.din(w_dff_B_Le8Canjh3_0),.dout(w_dff_B_lhdOWkJI7_0),.clk(gclk));
	jdff dff_B_sfWgnykp5_0(.din(w_dff_B_lhdOWkJI7_0),.dout(w_dff_B_sfWgnykp5_0),.clk(gclk));
	jdff dff_B_nQjRrXT37_0(.din(w_dff_B_sfWgnykp5_0),.dout(w_dff_B_nQjRrXT37_0),.clk(gclk));
	jdff dff_B_9dfk2v6l8_0(.din(w_dff_B_nQjRrXT37_0),.dout(w_dff_B_9dfk2v6l8_0),.clk(gclk));
	jdff dff_B_4Sk6MFFu2_0(.din(w_dff_B_9dfk2v6l8_0),.dout(w_dff_B_4Sk6MFFu2_0),.clk(gclk));
	jdff dff_B_0sNlxbt18_0(.din(w_dff_B_4Sk6MFFu2_0),.dout(w_dff_B_0sNlxbt18_0),.clk(gclk));
	jdff dff_B_0F3aU7Xk2_0(.din(w_dff_B_0sNlxbt18_0),.dout(w_dff_B_0F3aU7Xk2_0),.clk(gclk));
	jdff dff_B_IETck1EM7_0(.din(w_dff_B_0F3aU7Xk2_0),.dout(w_dff_B_IETck1EM7_0),.clk(gclk));
	jdff dff_B_iDnLCt3V6_0(.din(w_dff_B_IETck1EM7_0),.dout(w_dff_B_iDnLCt3V6_0),.clk(gclk));
	jdff dff_B_oT6Q1veI4_0(.din(w_dff_B_iDnLCt3V6_0),.dout(w_dff_B_oT6Q1veI4_0),.clk(gclk));
	jdff dff_B_Qddfi4658_0(.din(w_dff_B_oT6Q1veI4_0),.dout(w_dff_B_Qddfi4658_0),.clk(gclk));
	jdff dff_B_asck50dK0_0(.din(w_dff_B_Qddfi4658_0),.dout(w_dff_B_asck50dK0_0),.clk(gclk));
	jdff dff_B_xc1yyz7X4_0(.din(w_dff_B_asck50dK0_0),.dout(w_dff_B_xc1yyz7X4_0),.clk(gclk));
	jdff dff_B_4WbD3Ruu4_0(.din(w_dff_B_xc1yyz7X4_0),.dout(w_dff_B_4WbD3Ruu4_0),.clk(gclk));
	jdff dff_B_ygJPhuTH1_0(.din(w_dff_B_4WbD3Ruu4_0),.dout(w_dff_B_ygJPhuTH1_0),.clk(gclk));
	jdff dff_B_t4ihs8jP1_0(.din(w_dff_B_ygJPhuTH1_0),.dout(w_dff_B_t4ihs8jP1_0),.clk(gclk));
	jdff dff_B_OOmlmDZy0_0(.din(w_dff_B_t4ihs8jP1_0),.dout(w_dff_B_OOmlmDZy0_0),.clk(gclk));
	jdff dff_B_q3sb1ZZ37_0(.din(w_dff_B_OOmlmDZy0_0),.dout(w_dff_B_q3sb1ZZ37_0),.clk(gclk));
	jdff dff_B_fDvSImvh6_0(.din(w_dff_B_q3sb1ZZ37_0),.dout(w_dff_B_fDvSImvh6_0),.clk(gclk));
	jdff dff_B_eAv5gTy56_0(.din(w_dff_B_fDvSImvh6_0),.dout(w_dff_B_eAv5gTy56_0),.clk(gclk));
	jdff dff_B_tu1W32LA1_0(.din(w_dff_B_eAv5gTy56_0),.dout(w_dff_B_tu1W32LA1_0),.clk(gclk));
	jdff dff_B_4fpJw69N2_0(.din(w_dff_B_tu1W32LA1_0),.dout(w_dff_B_4fpJw69N2_0),.clk(gclk));
	jdff dff_B_j8top92t0_0(.din(w_dff_B_4fpJw69N2_0),.dout(w_dff_B_j8top92t0_0),.clk(gclk));
	jdff dff_B_giU7u6ow1_0(.din(w_dff_B_j8top92t0_0),.dout(w_dff_B_giU7u6ow1_0),.clk(gclk));
	jdff dff_B_ybnAhAMc9_0(.din(w_dff_B_giU7u6ow1_0),.dout(w_dff_B_ybnAhAMc9_0),.clk(gclk));
	jdff dff_B_pEIs1MsE1_0(.din(w_dff_B_ybnAhAMc9_0),.dout(w_dff_B_pEIs1MsE1_0),.clk(gclk));
	jdff dff_B_Iv4h4NTC2_0(.din(w_dff_B_pEIs1MsE1_0),.dout(w_dff_B_Iv4h4NTC2_0),.clk(gclk));
	jdff dff_B_uixhFbrS8_0(.din(w_dff_B_Iv4h4NTC2_0),.dout(w_dff_B_uixhFbrS8_0),.clk(gclk));
	jdff dff_B_VdGqVnLr0_0(.din(w_dff_B_uixhFbrS8_0),.dout(w_dff_B_VdGqVnLr0_0),.clk(gclk));
	jdff dff_B_zQLbocjZ8_0(.din(w_dff_B_VdGqVnLr0_0),.dout(w_dff_B_zQLbocjZ8_0),.clk(gclk));
	jdff dff_B_7zcYi1To6_0(.din(w_dff_B_zQLbocjZ8_0),.dout(w_dff_B_7zcYi1To6_0),.clk(gclk));
	jdff dff_B_v4lHygoC3_0(.din(w_dff_B_7zcYi1To6_0),.dout(w_dff_B_v4lHygoC3_0),.clk(gclk));
	jdff dff_B_proeNED82_0(.din(w_dff_B_v4lHygoC3_0),.dout(w_dff_B_proeNED82_0),.clk(gclk));
	jdff dff_B_Ud0vc5AS6_0(.din(w_dff_B_proeNED82_0),.dout(w_dff_B_Ud0vc5AS6_0),.clk(gclk));
	jdff dff_B_JAvHcDPl3_0(.din(w_dff_B_Ud0vc5AS6_0),.dout(w_dff_B_JAvHcDPl3_0),.clk(gclk));
	jdff dff_B_x19qJt542_0(.din(w_dff_B_JAvHcDPl3_0),.dout(w_dff_B_x19qJt542_0),.clk(gclk));
	jdff dff_B_Xo2I9Atg9_0(.din(w_dff_B_x19qJt542_0),.dout(w_dff_B_Xo2I9Atg9_0),.clk(gclk));
	jdff dff_B_dVLQmnYY3_0(.din(w_dff_B_Xo2I9Atg9_0),.dout(w_dff_B_dVLQmnYY3_0),.clk(gclk));
	jdff dff_B_AlsrzvHm5_0(.din(w_dff_B_dVLQmnYY3_0),.dout(w_dff_B_AlsrzvHm5_0),.clk(gclk));
	jdff dff_B_zVmuojRz8_0(.din(w_dff_B_AlsrzvHm5_0),.dout(w_dff_B_zVmuojRz8_0),.clk(gclk));
	jdff dff_B_gr65bRSH8_0(.din(w_dff_B_zVmuojRz8_0),.dout(w_dff_B_gr65bRSH8_0),.clk(gclk));
	jdff dff_B_Vih6pky98_0(.din(w_dff_B_gr65bRSH8_0),.dout(w_dff_B_Vih6pky98_0),.clk(gclk));
	jdff dff_B_DREh6Ggg1_0(.din(w_dff_B_Vih6pky98_0),.dout(w_dff_B_DREh6Ggg1_0),.clk(gclk));
	jdff dff_B_kVLy3ipX6_0(.din(w_dff_B_DREh6Ggg1_0),.dout(w_dff_B_kVLy3ipX6_0),.clk(gclk));
	jdff dff_B_Di5LgRRX3_0(.din(w_dff_B_kVLy3ipX6_0),.dout(w_dff_B_Di5LgRRX3_0),.clk(gclk));
	jdff dff_B_kvlNU53N1_0(.din(w_dff_B_Di5LgRRX3_0),.dout(w_dff_B_kvlNU53N1_0),.clk(gclk));
	jdff dff_B_0aMKTrjg4_0(.din(w_dff_B_kvlNU53N1_0),.dout(w_dff_B_0aMKTrjg4_0),.clk(gclk));
	jdff dff_B_yFJWLOEU1_0(.din(w_dff_B_0aMKTrjg4_0),.dout(w_dff_B_yFJWLOEU1_0),.clk(gclk));
	jdff dff_B_6ZjTiqxA7_0(.din(w_dff_B_yFJWLOEU1_0),.dout(w_dff_B_6ZjTiqxA7_0),.clk(gclk));
	jdff dff_B_JA9I5uAh1_0(.din(w_dff_B_6ZjTiqxA7_0),.dout(w_dff_B_JA9I5uAh1_0),.clk(gclk));
	jdff dff_B_Vr1dtRmG6_0(.din(w_dff_B_JA9I5uAh1_0),.dout(w_dff_B_Vr1dtRmG6_0),.clk(gclk));
	jdff dff_B_nFCXKPYZ1_0(.din(w_dff_B_Vr1dtRmG6_0),.dout(w_dff_B_nFCXKPYZ1_0),.clk(gclk));
	jdff dff_B_1TqtO5gz9_0(.din(w_dff_B_nFCXKPYZ1_0),.dout(w_dff_B_1TqtO5gz9_0),.clk(gclk));
	jdff dff_B_vwtDePh67_0(.din(w_dff_B_1TqtO5gz9_0),.dout(w_dff_B_vwtDePh67_0),.clk(gclk));
	jdff dff_B_efUGQzXU9_0(.din(w_dff_B_vwtDePh67_0),.dout(w_dff_B_efUGQzXU9_0),.clk(gclk));
	jdff dff_B_c2gXUocZ1_0(.din(w_dff_B_efUGQzXU9_0),.dout(w_dff_B_c2gXUocZ1_0),.clk(gclk));
	jdff dff_B_a7wPIu1f1_0(.din(w_dff_B_c2gXUocZ1_0),.dout(w_dff_B_a7wPIu1f1_0),.clk(gclk));
	jdff dff_B_8SgZofGF7_0(.din(w_dff_B_a7wPIu1f1_0),.dout(w_dff_B_8SgZofGF7_0),.clk(gclk));
	jdff dff_B_Mcr16eGs4_0(.din(w_dff_B_8SgZofGF7_0),.dout(w_dff_B_Mcr16eGs4_0),.clk(gclk));
	jdff dff_B_7RUTZ4zU2_1(.din(n774),.dout(w_dff_B_7RUTZ4zU2_1),.clk(gclk));
	jdff dff_B_zh4yBwlC6_1(.din(w_dff_B_7RUTZ4zU2_1),.dout(w_dff_B_zh4yBwlC6_1),.clk(gclk));
	jdff dff_B_6kluDntq0_1(.din(w_dff_B_zh4yBwlC6_1),.dout(w_dff_B_6kluDntq0_1),.clk(gclk));
	jdff dff_B_69QmJAUD5_1(.din(w_dff_B_6kluDntq0_1),.dout(w_dff_B_69QmJAUD5_1),.clk(gclk));
	jdff dff_B_eUsldsk62_1(.din(w_dff_B_69QmJAUD5_1),.dout(w_dff_B_eUsldsk62_1),.clk(gclk));
	jdff dff_B_eDqPIPgc3_1(.din(w_dff_B_eUsldsk62_1),.dout(w_dff_B_eDqPIPgc3_1),.clk(gclk));
	jdff dff_B_CKXEPosv7_1(.din(w_dff_B_eDqPIPgc3_1),.dout(w_dff_B_CKXEPosv7_1),.clk(gclk));
	jdff dff_B_g71M3N2a3_1(.din(w_dff_B_CKXEPosv7_1),.dout(w_dff_B_g71M3N2a3_1),.clk(gclk));
	jdff dff_B_ROXgn1xk4_1(.din(w_dff_B_g71M3N2a3_1),.dout(w_dff_B_ROXgn1xk4_1),.clk(gclk));
	jdff dff_B_UBk1rUiz5_1(.din(w_dff_B_ROXgn1xk4_1),.dout(w_dff_B_UBk1rUiz5_1),.clk(gclk));
	jdff dff_B_grIg65Bo8_1(.din(w_dff_B_UBk1rUiz5_1),.dout(w_dff_B_grIg65Bo8_1),.clk(gclk));
	jdff dff_B_3su8UvJ92_1(.din(w_dff_B_grIg65Bo8_1),.dout(w_dff_B_3su8UvJ92_1),.clk(gclk));
	jdff dff_B_y2O6myBI6_1(.din(w_dff_B_3su8UvJ92_1),.dout(w_dff_B_y2O6myBI6_1),.clk(gclk));
	jdff dff_B_JMfa18Nx5_1(.din(w_dff_B_y2O6myBI6_1),.dout(w_dff_B_JMfa18Nx5_1),.clk(gclk));
	jdff dff_B_d1WlfRUu6_1(.din(w_dff_B_JMfa18Nx5_1),.dout(w_dff_B_d1WlfRUu6_1),.clk(gclk));
	jdff dff_B_Bgc7zlAf7_1(.din(w_dff_B_d1WlfRUu6_1),.dout(w_dff_B_Bgc7zlAf7_1),.clk(gclk));
	jdff dff_B_tLE6cLRp7_1(.din(w_dff_B_Bgc7zlAf7_1),.dout(w_dff_B_tLE6cLRp7_1),.clk(gclk));
	jdff dff_B_CiVge8Qz6_1(.din(w_dff_B_tLE6cLRp7_1),.dout(w_dff_B_CiVge8Qz6_1),.clk(gclk));
	jdff dff_B_hjHbACXu9_1(.din(w_dff_B_CiVge8Qz6_1),.dout(w_dff_B_hjHbACXu9_1),.clk(gclk));
	jdff dff_B_iUWCiWiG5_1(.din(w_dff_B_hjHbACXu9_1),.dout(w_dff_B_iUWCiWiG5_1),.clk(gclk));
	jdff dff_B_ym415l320_1(.din(w_dff_B_iUWCiWiG5_1),.dout(w_dff_B_ym415l320_1),.clk(gclk));
	jdff dff_B_RR2qjc2W0_1(.din(w_dff_B_ym415l320_1),.dout(w_dff_B_RR2qjc2W0_1),.clk(gclk));
	jdff dff_B_G7vkg4dJ7_1(.din(w_dff_B_RR2qjc2W0_1),.dout(w_dff_B_G7vkg4dJ7_1),.clk(gclk));
	jdff dff_B_kfw8nkjS4_1(.din(w_dff_B_G7vkg4dJ7_1),.dout(w_dff_B_kfw8nkjS4_1),.clk(gclk));
	jdff dff_B_L2I1VkNL2_1(.din(w_dff_B_kfw8nkjS4_1),.dout(w_dff_B_L2I1VkNL2_1),.clk(gclk));
	jdff dff_B_pCmAb4DC9_1(.din(w_dff_B_L2I1VkNL2_1),.dout(w_dff_B_pCmAb4DC9_1),.clk(gclk));
	jdff dff_B_CkGmlYcr0_1(.din(w_dff_B_pCmAb4DC9_1),.dout(w_dff_B_CkGmlYcr0_1),.clk(gclk));
	jdff dff_B_02oPRZOV9_1(.din(w_dff_B_CkGmlYcr0_1),.dout(w_dff_B_02oPRZOV9_1),.clk(gclk));
	jdff dff_B_saTYnvjd4_1(.din(w_dff_B_02oPRZOV9_1),.dout(w_dff_B_saTYnvjd4_1),.clk(gclk));
	jdff dff_B_xSds98j35_1(.din(w_dff_B_saTYnvjd4_1),.dout(w_dff_B_xSds98j35_1),.clk(gclk));
	jdff dff_B_8G5Feubv2_1(.din(w_dff_B_xSds98j35_1),.dout(w_dff_B_8G5Feubv2_1),.clk(gclk));
	jdff dff_B_il0oKbyf7_1(.din(w_dff_B_8G5Feubv2_1),.dout(w_dff_B_il0oKbyf7_1),.clk(gclk));
	jdff dff_B_gKyPP9wD0_1(.din(w_dff_B_il0oKbyf7_1),.dout(w_dff_B_gKyPP9wD0_1),.clk(gclk));
	jdff dff_B_2tFGeIHX4_1(.din(w_dff_B_gKyPP9wD0_1),.dout(w_dff_B_2tFGeIHX4_1),.clk(gclk));
	jdff dff_B_6IZBCQvH0_1(.din(w_dff_B_2tFGeIHX4_1),.dout(w_dff_B_6IZBCQvH0_1),.clk(gclk));
	jdff dff_B_3bwl2I039_1(.din(w_dff_B_6IZBCQvH0_1),.dout(w_dff_B_3bwl2I039_1),.clk(gclk));
	jdff dff_B_0bTe5xoN7_1(.din(w_dff_B_3bwl2I039_1),.dout(w_dff_B_0bTe5xoN7_1),.clk(gclk));
	jdff dff_B_gho2VcCs6_1(.din(w_dff_B_0bTe5xoN7_1),.dout(w_dff_B_gho2VcCs6_1),.clk(gclk));
	jdff dff_B_3gaMNsXM6_1(.din(w_dff_B_gho2VcCs6_1),.dout(w_dff_B_3gaMNsXM6_1),.clk(gclk));
	jdff dff_B_BbFk8HaN1_1(.din(w_dff_B_3gaMNsXM6_1),.dout(w_dff_B_BbFk8HaN1_1),.clk(gclk));
	jdff dff_B_ffg2xW9O3_1(.din(w_dff_B_BbFk8HaN1_1),.dout(w_dff_B_ffg2xW9O3_1),.clk(gclk));
	jdff dff_B_IeNIno6q0_1(.din(w_dff_B_ffg2xW9O3_1),.dout(w_dff_B_IeNIno6q0_1),.clk(gclk));
	jdff dff_B_XBQnb87s0_1(.din(w_dff_B_IeNIno6q0_1),.dout(w_dff_B_XBQnb87s0_1),.clk(gclk));
	jdff dff_B_wgL2iy9s2_1(.din(w_dff_B_XBQnb87s0_1),.dout(w_dff_B_wgL2iy9s2_1),.clk(gclk));
	jdff dff_B_ulxkTynz5_1(.din(w_dff_B_wgL2iy9s2_1),.dout(w_dff_B_ulxkTynz5_1),.clk(gclk));
	jdff dff_B_iSyD2i7a9_1(.din(w_dff_B_ulxkTynz5_1),.dout(w_dff_B_iSyD2i7a9_1),.clk(gclk));
	jdff dff_B_zVhLE4EG2_1(.din(w_dff_B_iSyD2i7a9_1),.dout(w_dff_B_zVhLE4EG2_1),.clk(gclk));
	jdff dff_B_mFwyxYtW1_1(.din(w_dff_B_zVhLE4EG2_1),.dout(w_dff_B_mFwyxYtW1_1),.clk(gclk));
	jdff dff_B_KqXYvtun4_1(.din(w_dff_B_mFwyxYtW1_1),.dout(w_dff_B_KqXYvtun4_1),.clk(gclk));
	jdff dff_B_0zHvMaRL8_1(.din(w_dff_B_KqXYvtun4_1),.dout(w_dff_B_0zHvMaRL8_1),.clk(gclk));
	jdff dff_B_FTiAOK5M1_1(.din(w_dff_B_0zHvMaRL8_1),.dout(w_dff_B_FTiAOK5M1_1),.clk(gclk));
	jdff dff_B_k13IfzzH0_1(.din(w_dff_B_FTiAOK5M1_1),.dout(w_dff_B_k13IfzzH0_1),.clk(gclk));
	jdff dff_B_x5Xq9cFG9_1(.din(w_dff_B_k13IfzzH0_1),.dout(w_dff_B_x5Xq9cFG9_1),.clk(gclk));
	jdff dff_B_6yQkGmP23_1(.din(w_dff_B_x5Xq9cFG9_1),.dout(w_dff_B_6yQkGmP23_1),.clk(gclk));
	jdff dff_B_qzzrmTg50_1(.din(w_dff_B_6yQkGmP23_1),.dout(w_dff_B_qzzrmTg50_1),.clk(gclk));
	jdff dff_B_xMjyzten7_1(.din(w_dff_B_qzzrmTg50_1),.dout(w_dff_B_xMjyzten7_1),.clk(gclk));
	jdff dff_B_uaBMf0Ov5_1(.din(w_dff_B_xMjyzten7_1),.dout(w_dff_B_uaBMf0Ov5_1),.clk(gclk));
	jdff dff_B_rrrKqrcF5_1(.din(w_dff_B_uaBMf0Ov5_1),.dout(w_dff_B_rrrKqrcF5_1),.clk(gclk));
	jdff dff_B_JsQwJtSs2_1(.din(w_dff_B_rrrKqrcF5_1),.dout(w_dff_B_JsQwJtSs2_1),.clk(gclk));
	jdff dff_B_O21dVdx15_1(.din(w_dff_B_JsQwJtSs2_1),.dout(w_dff_B_O21dVdx15_1),.clk(gclk));
	jdff dff_B_ZideBjrU7_1(.din(w_dff_B_O21dVdx15_1),.dout(w_dff_B_ZideBjrU7_1),.clk(gclk));
	jdff dff_B_Gjyh2fKb3_1(.din(w_dff_B_ZideBjrU7_1),.dout(w_dff_B_Gjyh2fKb3_1),.clk(gclk));
	jdff dff_B_1rSLPhl06_1(.din(w_dff_B_Gjyh2fKb3_1),.dout(w_dff_B_1rSLPhl06_1),.clk(gclk));
	jdff dff_B_hKx3fuL67_1(.din(w_dff_B_1rSLPhl06_1),.dout(w_dff_B_hKx3fuL67_1),.clk(gclk));
	jdff dff_B_NsY7JH502_1(.din(w_dff_B_hKx3fuL67_1),.dout(w_dff_B_NsY7JH502_1),.clk(gclk));
	jdff dff_B_GEUzZB1m6_0(.din(n775),.dout(w_dff_B_GEUzZB1m6_0),.clk(gclk));
	jdff dff_B_EgxhAFsZ9_0(.din(w_dff_B_GEUzZB1m6_0),.dout(w_dff_B_EgxhAFsZ9_0),.clk(gclk));
	jdff dff_B_lmHDZMkk9_0(.din(w_dff_B_EgxhAFsZ9_0),.dout(w_dff_B_lmHDZMkk9_0),.clk(gclk));
	jdff dff_B_NtrhFY9P1_0(.din(w_dff_B_lmHDZMkk9_0),.dout(w_dff_B_NtrhFY9P1_0),.clk(gclk));
	jdff dff_B_Era2yddZ9_0(.din(w_dff_B_NtrhFY9P1_0),.dout(w_dff_B_Era2yddZ9_0),.clk(gclk));
	jdff dff_B_u1dbi5Aj6_0(.din(w_dff_B_Era2yddZ9_0),.dout(w_dff_B_u1dbi5Aj6_0),.clk(gclk));
	jdff dff_B_wfLV2Djz7_0(.din(w_dff_B_u1dbi5Aj6_0),.dout(w_dff_B_wfLV2Djz7_0),.clk(gclk));
	jdff dff_B_p6vknCGc5_0(.din(w_dff_B_wfLV2Djz7_0),.dout(w_dff_B_p6vknCGc5_0),.clk(gclk));
	jdff dff_B_rk60TxdO8_0(.din(w_dff_B_p6vknCGc5_0),.dout(w_dff_B_rk60TxdO8_0),.clk(gclk));
	jdff dff_B_wOTquhKX1_0(.din(w_dff_B_rk60TxdO8_0),.dout(w_dff_B_wOTquhKX1_0),.clk(gclk));
	jdff dff_B_cabrGrRQ6_0(.din(w_dff_B_wOTquhKX1_0),.dout(w_dff_B_cabrGrRQ6_0),.clk(gclk));
	jdff dff_B_172tfGOf4_0(.din(w_dff_B_cabrGrRQ6_0),.dout(w_dff_B_172tfGOf4_0),.clk(gclk));
	jdff dff_B_AA3vfSq39_0(.din(w_dff_B_172tfGOf4_0),.dout(w_dff_B_AA3vfSq39_0),.clk(gclk));
	jdff dff_B_ZVdcox9C2_0(.din(w_dff_B_AA3vfSq39_0),.dout(w_dff_B_ZVdcox9C2_0),.clk(gclk));
	jdff dff_B_cspLt6N93_0(.din(w_dff_B_ZVdcox9C2_0),.dout(w_dff_B_cspLt6N93_0),.clk(gclk));
	jdff dff_B_EDBypqyU3_0(.din(w_dff_B_cspLt6N93_0),.dout(w_dff_B_EDBypqyU3_0),.clk(gclk));
	jdff dff_B_4HkFUDsW2_0(.din(w_dff_B_EDBypqyU3_0),.dout(w_dff_B_4HkFUDsW2_0),.clk(gclk));
	jdff dff_B_RKuAUXUZ9_0(.din(w_dff_B_4HkFUDsW2_0),.dout(w_dff_B_RKuAUXUZ9_0),.clk(gclk));
	jdff dff_B_1USPPnLV9_0(.din(w_dff_B_RKuAUXUZ9_0),.dout(w_dff_B_1USPPnLV9_0),.clk(gclk));
	jdff dff_B_66L2saSR9_0(.din(w_dff_B_1USPPnLV9_0),.dout(w_dff_B_66L2saSR9_0),.clk(gclk));
	jdff dff_B_WFUGenHp2_0(.din(w_dff_B_66L2saSR9_0),.dout(w_dff_B_WFUGenHp2_0),.clk(gclk));
	jdff dff_B_uOZQLOrV2_0(.din(w_dff_B_WFUGenHp2_0),.dout(w_dff_B_uOZQLOrV2_0),.clk(gclk));
	jdff dff_B_uW1X7DZu7_0(.din(w_dff_B_uOZQLOrV2_0),.dout(w_dff_B_uW1X7DZu7_0),.clk(gclk));
	jdff dff_B_hoaUnRl34_0(.din(w_dff_B_uW1X7DZu7_0),.dout(w_dff_B_hoaUnRl34_0),.clk(gclk));
	jdff dff_B_hkM24vPM3_0(.din(w_dff_B_hoaUnRl34_0),.dout(w_dff_B_hkM24vPM3_0),.clk(gclk));
	jdff dff_B_l2EG3j3S2_0(.din(w_dff_B_hkM24vPM3_0),.dout(w_dff_B_l2EG3j3S2_0),.clk(gclk));
	jdff dff_B_CfEy3taW2_0(.din(w_dff_B_l2EG3j3S2_0),.dout(w_dff_B_CfEy3taW2_0),.clk(gclk));
	jdff dff_B_Skt9gxQk7_0(.din(w_dff_B_CfEy3taW2_0),.dout(w_dff_B_Skt9gxQk7_0),.clk(gclk));
	jdff dff_B_y8oJOJv10_0(.din(w_dff_B_Skt9gxQk7_0),.dout(w_dff_B_y8oJOJv10_0),.clk(gclk));
	jdff dff_B_Zp8rVhpO8_0(.din(w_dff_B_y8oJOJv10_0),.dout(w_dff_B_Zp8rVhpO8_0),.clk(gclk));
	jdff dff_B_sdxLvkqM2_0(.din(w_dff_B_Zp8rVhpO8_0),.dout(w_dff_B_sdxLvkqM2_0),.clk(gclk));
	jdff dff_B_dz5ojoSk0_0(.din(w_dff_B_sdxLvkqM2_0),.dout(w_dff_B_dz5ojoSk0_0),.clk(gclk));
	jdff dff_B_D09QsuvI5_0(.din(w_dff_B_dz5ojoSk0_0),.dout(w_dff_B_D09QsuvI5_0),.clk(gclk));
	jdff dff_B_vYWBSVrn3_0(.din(w_dff_B_D09QsuvI5_0),.dout(w_dff_B_vYWBSVrn3_0),.clk(gclk));
	jdff dff_B_EQZcIIy48_0(.din(w_dff_B_vYWBSVrn3_0),.dout(w_dff_B_EQZcIIy48_0),.clk(gclk));
	jdff dff_B_fPOg4O0G3_0(.din(w_dff_B_EQZcIIy48_0),.dout(w_dff_B_fPOg4O0G3_0),.clk(gclk));
	jdff dff_B_ze07Q5ma2_0(.din(w_dff_B_fPOg4O0G3_0),.dout(w_dff_B_ze07Q5ma2_0),.clk(gclk));
	jdff dff_B_0xlaqssf2_0(.din(w_dff_B_ze07Q5ma2_0),.dout(w_dff_B_0xlaqssf2_0),.clk(gclk));
	jdff dff_B_N9PkOXHb4_0(.din(w_dff_B_0xlaqssf2_0),.dout(w_dff_B_N9PkOXHb4_0),.clk(gclk));
	jdff dff_B_M94hMR660_0(.din(w_dff_B_N9PkOXHb4_0),.dout(w_dff_B_M94hMR660_0),.clk(gclk));
	jdff dff_B_W8njf6Rr0_0(.din(w_dff_B_M94hMR660_0),.dout(w_dff_B_W8njf6Rr0_0),.clk(gclk));
	jdff dff_B_VHMMMsFQ0_0(.din(w_dff_B_W8njf6Rr0_0),.dout(w_dff_B_VHMMMsFQ0_0),.clk(gclk));
	jdff dff_B_wViNcPEe6_0(.din(w_dff_B_VHMMMsFQ0_0),.dout(w_dff_B_wViNcPEe6_0),.clk(gclk));
	jdff dff_B_dmqzSnUX6_0(.din(w_dff_B_wViNcPEe6_0),.dout(w_dff_B_dmqzSnUX6_0),.clk(gclk));
	jdff dff_B_do8guoy77_0(.din(w_dff_B_dmqzSnUX6_0),.dout(w_dff_B_do8guoy77_0),.clk(gclk));
	jdff dff_B_IR1vPNZS1_0(.din(w_dff_B_do8guoy77_0),.dout(w_dff_B_IR1vPNZS1_0),.clk(gclk));
	jdff dff_B_X2HsWHIV2_0(.din(w_dff_B_IR1vPNZS1_0),.dout(w_dff_B_X2HsWHIV2_0),.clk(gclk));
	jdff dff_B_uOFHBJ8Q2_0(.din(w_dff_B_X2HsWHIV2_0),.dout(w_dff_B_uOFHBJ8Q2_0),.clk(gclk));
	jdff dff_B_G6aAfiPF9_0(.din(w_dff_B_uOFHBJ8Q2_0),.dout(w_dff_B_G6aAfiPF9_0),.clk(gclk));
	jdff dff_B_m4LbWDCE6_0(.din(w_dff_B_G6aAfiPF9_0),.dout(w_dff_B_m4LbWDCE6_0),.clk(gclk));
	jdff dff_B_wGnGLw7v7_0(.din(w_dff_B_m4LbWDCE6_0),.dout(w_dff_B_wGnGLw7v7_0),.clk(gclk));
	jdff dff_B_JEVXnVFX1_0(.din(w_dff_B_wGnGLw7v7_0),.dout(w_dff_B_JEVXnVFX1_0),.clk(gclk));
	jdff dff_B_eD2NTRBl2_0(.din(w_dff_B_JEVXnVFX1_0),.dout(w_dff_B_eD2NTRBl2_0),.clk(gclk));
	jdff dff_B_m5t01a8u0_0(.din(w_dff_B_eD2NTRBl2_0),.dout(w_dff_B_m5t01a8u0_0),.clk(gclk));
	jdff dff_B_FKoGc5pu2_0(.din(w_dff_B_m5t01a8u0_0),.dout(w_dff_B_FKoGc5pu2_0),.clk(gclk));
	jdff dff_B_cLQrrrTq9_0(.din(w_dff_B_FKoGc5pu2_0),.dout(w_dff_B_cLQrrrTq9_0),.clk(gclk));
	jdff dff_B_8OAmP6dJ4_0(.din(w_dff_B_cLQrrrTq9_0),.dout(w_dff_B_8OAmP6dJ4_0),.clk(gclk));
	jdff dff_B_JupuSsmG5_0(.din(w_dff_B_8OAmP6dJ4_0),.dout(w_dff_B_JupuSsmG5_0),.clk(gclk));
	jdff dff_B_ZYq0H2iY3_0(.din(w_dff_B_JupuSsmG5_0),.dout(w_dff_B_ZYq0H2iY3_0),.clk(gclk));
	jdff dff_B_blAMKkR16_0(.din(w_dff_B_ZYq0H2iY3_0),.dout(w_dff_B_blAMKkR16_0),.clk(gclk));
	jdff dff_B_q2LgQ0Gs2_0(.din(w_dff_B_blAMKkR16_0),.dout(w_dff_B_q2LgQ0Gs2_0),.clk(gclk));
	jdff dff_B_SEkSkBZV6_0(.din(w_dff_B_q2LgQ0Gs2_0),.dout(w_dff_B_SEkSkBZV6_0),.clk(gclk));
	jdff dff_B_GAvcsof61_0(.din(w_dff_B_SEkSkBZV6_0),.dout(w_dff_B_GAvcsof61_0),.clk(gclk));
	jdff dff_B_m8F3KBwR0_0(.din(w_dff_B_GAvcsof61_0),.dout(w_dff_B_m8F3KBwR0_0),.clk(gclk));
	jdff dff_B_CuQ7QQJA6_0(.din(w_dff_B_m8F3KBwR0_0),.dout(w_dff_B_CuQ7QQJA6_0),.clk(gclk));
	jdff dff_B_nS8rjJeB5_1(.din(n768),.dout(w_dff_B_nS8rjJeB5_1),.clk(gclk));
	jdff dff_B_VTPBg5wx6_1(.din(w_dff_B_nS8rjJeB5_1),.dout(w_dff_B_VTPBg5wx6_1),.clk(gclk));
	jdff dff_B_eBidpytV4_1(.din(w_dff_B_VTPBg5wx6_1),.dout(w_dff_B_eBidpytV4_1),.clk(gclk));
	jdff dff_B_Jj6e9lh24_1(.din(w_dff_B_eBidpytV4_1),.dout(w_dff_B_Jj6e9lh24_1),.clk(gclk));
	jdff dff_B_A7suurIY2_1(.din(w_dff_B_Jj6e9lh24_1),.dout(w_dff_B_A7suurIY2_1),.clk(gclk));
	jdff dff_B_hsOgVLe48_1(.din(w_dff_B_A7suurIY2_1),.dout(w_dff_B_hsOgVLe48_1),.clk(gclk));
	jdff dff_B_yjjAjc7x8_1(.din(w_dff_B_hsOgVLe48_1),.dout(w_dff_B_yjjAjc7x8_1),.clk(gclk));
	jdff dff_B_QpFQWZ810_1(.din(w_dff_B_yjjAjc7x8_1),.dout(w_dff_B_QpFQWZ810_1),.clk(gclk));
	jdff dff_B_nQ7HpCc60_1(.din(w_dff_B_QpFQWZ810_1),.dout(w_dff_B_nQ7HpCc60_1),.clk(gclk));
	jdff dff_B_AHIsHExp9_1(.din(w_dff_B_nQ7HpCc60_1),.dout(w_dff_B_AHIsHExp9_1),.clk(gclk));
	jdff dff_B_I3MQ57Gs4_1(.din(w_dff_B_AHIsHExp9_1),.dout(w_dff_B_I3MQ57Gs4_1),.clk(gclk));
	jdff dff_B_FH0zwPGi3_1(.din(w_dff_B_I3MQ57Gs4_1),.dout(w_dff_B_FH0zwPGi3_1),.clk(gclk));
	jdff dff_B_d78C6Lkt9_1(.din(w_dff_B_FH0zwPGi3_1),.dout(w_dff_B_d78C6Lkt9_1),.clk(gclk));
	jdff dff_B_Hz39arMe4_1(.din(w_dff_B_d78C6Lkt9_1),.dout(w_dff_B_Hz39arMe4_1),.clk(gclk));
	jdff dff_B_2toyf6gO0_1(.din(w_dff_B_Hz39arMe4_1),.dout(w_dff_B_2toyf6gO0_1),.clk(gclk));
	jdff dff_B_S4z1YssN2_1(.din(w_dff_B_2toyf6gO0_1),.dout(w_dff_B_S4z1YssN2_1),.clk(gclk));
	jdff dff_B_w668kYAL8_1(.din(w_dff_B_S4z1YssN2_1),.dout(w_dff_B_w668kYAL8_1),.clk(gclk));
	jdff dff_B_7Odta9Xs7_1(.din(w_dff_B_w668kYAL8_1),.dout(w_dff_B_7Odta9Xs7_1),.clk(gclk));
	jdff dff_B_FK8CKacm3_1(.din(w_dff_B_7Odta9Xs7_1),.dout(w_dff_B_FK8CKacm3_1),.clk(gclk));
	jdff dff_B_A6gyFyOH3_1(.din(w_dff_B_FK8CKacm3_1),.dout(w_dff_B_A6gyFyOH3_1),.clk(gclk));
	jdff dff_B_laPivbMg4_1(.din(w_dff_B_A6gyFyOH3_1),.dout(w_dff_B_laPivbMg4_1),.clk(gclk));
	jdff dff_B_vyb1i9MF2_1(.din(w_dff_B_laPivbMg4_1),.dout(w_dff_B_vyb1i9MF2_1),.clk(gclk));
	jdff dff_B_3KTwAvUB4_1(.din(w_dff_B_vyb1i9MF2_1),.dout(w_dff_B_3KTwAvUB4_1),.clk(gclk));
	jdff dff_B_zs3MaSr95_1(.din(w_dff_B_3KTwAvUB4_1),.dout(w_dff_B_zs3MaSr95_1),.clk(gclk));
	jdff dff_B_7OdJvSyP8_1(.din(w_dff_B_zs3MaSr95_1),.dout(w_dff_B_7OdJvSyP8_1),.clk(gclk));
	jdff dff_B_4jD6a6Bo2_1(.din(w_dff_B_7OdJvSyP8_1),.dout(w_dff_B_4jD6a6Bo2_1),.clk(gclk));
	jdff dff_B_iNB1kBqi3_1(.din(w_dff_B_4jD6a6Bo2_1),.dout(w_dff_B_iNB1kBqi3_1),.clk(gclk));
	jdff dff_B_IoUT6ftK3_1(.din(w_dff_B_iNB1kBqi3_1),.dout(w_dff_B_IoUT6ftK3_1),.clk(gclk));
	jdff dff_B_9TmBcy0q4_1(.din(w_dff_B_IoUT6ftK3_1),.dout(w_dff_B_9TmBcy0q4_1),.clk(gclk));
	jdff dff_B_NwqlbZuE0_1(.din(w_dff_B_9TmBcy0q4_1),.dout(w_dff_B_NwqlbZuE0_1),.clk(gclk));
	jdff dff_B_7PxXoN4N0_1(.din(w_dff_B_NwqlbZuE0_1),.dout(w_dff_B_7PxXoN4N0_1),.clk(gclk));
	jdff dff_B_spE9vrh28_1(.din(w_dff_B_7PxXoN4N0_1),.dout(w_dff_B_spE9vrh28_1),.clk(gclk));
	jdff dff_B_S176hAA30_1(.din(w_dff_B_spE9vrh28_1),.dout(w_dff_B_S176hAA30_1),.clk(gclk));
	jdff dff_B_8AQbBgk44_1(.din(w_dff_B_S176hAA30_1),.dout(w_dff_B_8AQbBgk44_1),.clk(gclk));
	jdff dff_B_kqP8Zlwi1_1(.din(w_dff_B_8AQbBgk44_1),.dout(w_dff_B_kqP8Zlwi1_1),.clk(gclk));
	jdff dff_B_63wyduLu5_1(.din(w_dff_B_kqP8Zlwi1_1),.dout(w_dff_B_63wyduLu5_1),.clk(gclk));
	jdff dff_B_tIK3KKXj6_1(.din(w_dff_B_63wyduLu5_1),.dout(w_dff_B_tIK3KKXj6_1),.clk(gclk));
	jdff dff_B_UJK6vTrf5_1(.din(w_dff_B_tIK3KKXj6_1),.dout(w_dff_B_UJK6vTrf5_1),.clk(gclk));
	jdff dff_B_2NviqDDV3_1(.din(w_dff_B_UJK6vTrf5_1),.dout(w_dff_B_2NviqDDV3_1),.clk(gclk));
	jdff dff_B_AYUOc8Gs5_1(.din(w_dff_B_2NviqDDV3_1),.dout(w_dff_B_AYUOc8Gs5_1),.clk(gclk));
	jdff dff_B_j15IcKmA1_1(.din(w_dff_B_AYUOc8Gs5_1),.dout(w_dff_B_j15IcKmA1_1),.clk(gclk));
	jdff dff_B_OhtQOzVD0_1(.din(w_dff_B_j15IcKmA1_1),.dout(w_dff_B_OhtQOzVD0_1),.clk(gclk));
	jdff dff_B_KLCzHLKu7_1(.din(w_dff_B_OhtQOzVD0_1),.dout(w_dff_B_KLCzHLKu7_1),.clk(gclk));
	jdff dff_B_MdeiuEh41_1(.din(w_dff_B_KLCzHLKu7_1),.dout(w_dff_B_MdeiuEh41_1),.clk(gclk));
	jdff dff_B_5EvCmtn50_1(.din(w_dff_B_MdeiuEh41_1),.dout(w_dff_B_5EvCmtn50_1),.clk(gclk));
	jdff dff_B_SZYbdwEX3_1(.din(w_dff_B_5EvCmtn50_1),.dout(w_dff_B_SZYbdwEX3_1),.clk(gclk));
	jdff dff_B_6oy73FDB8_1(.din(w_dff_B_SZYbdwEX3_1),.dout(w_dff_B_6oy73FDB8_1),.clk(gclk));
	jdff dff_B_REoTtRit1_1(.din(w_dff_B_6oy73FDB8_1),.dout(w_dff_B_REoTtRit1_1),.clk(gclk));
	jdff dff_B_9avp0UTU2_1(.din(w_dff_B_REoTtRit1_1),.dout(w_dff_B_9avp0UTU2_1),.clk(gclk));
	jdff dff_B_hWNOZcnz8_1(.din(w_dff_B_9avp0UTU2_1),.dout(w_dff_B_hWNOZcnz8_1),.clk(gclk));
	jdff dff_B_HEGWyX2r6_1(.din(w_dff_B_hWNOZcnz8_1),.dout(w_dff_B_HEGWyX2r6_1),.clk(gclk));
	jdff dff_B_nfwDGdAw9_1(.din(w_dff_B_HEGWyX2r6_1),.dout(w_dff_B_nfwDGdAw9_1),.clk(gclk));
	jdff dff_B_d6AQp35w2_1(.din(w_dff_B_nfwDGdAw9_1),.dout(w_dff_B_d6AQp35w2_1),.clk(gclk));
	jdff dff_B_4jLjwKaP1_1(.din(w_dff_B_d6AQp35w2_1),.dout(w_dff_B_4jLjwKaP1_1),.clk(gclk));
	jdff dff_B_H4M4vGHf9_1(.din(w_dff_B_4jLjwKaP1_1),.dout(w_dff_B_H4M4vGHf9_1),.clk(gclk));
	jdff dff_B_waGw9LyA0_1(.din(w_dff_B_H4M4vGHf9_1),.dout(w_dff_B_waGw9LyA0_1),.clk(gclk));
	jdff dff_B_2Qva7Bku8_1(.din(w_dff_B_waGw9LyA0_1),.dout(w_dff_B_2Qva7Bku8_1),.clk(gclk));
	jdff dff_B_j2zzwqhC0_1(.din(w_dff_B_2Qva7Bku8_1),.dout(w_dff_B_j2zzwqhC0_1),.clk(gclk));
	jdff dff_B_JUIiLmhv4_1(.din(w_dff_B_j2zzwqhC0_1),.dout(w_dff_B_JUIiLmhv4_1),.clk(gclk));
	jdff dff_B_dhkiUpHi9_1(.din(w_dff_B_JUIiLmhv4_1),.dout(w_dff_B_dhkiUpHi9_1),.clk(gclk));
	jdff dff_B_vuJXoeI63_1(.din(w_dff_B_dhkiUpHi9_1),.dout(w_dff_B_vuJXoeI63_1),.clk(gclk));
	jdff dff_B_JYX8rV1H7_1(.din(w_dff_B_vuJXoeI63_1),.dout(w_dff_B_JYX8rV1H7_1),.clk(gclk));
	jdff dff_B_8Wtnif2L2_1(.din(w_dff_B_JYX8rV1H7_1),.dout(w_dff_B_8Wtnif2L2_1),.clk(gclk));
	jdff dff_B_7KmGZ0V04_1(.din(w_dff_B_8Wtnif2L2_1),.dout(w_dff_B_7KmGZ0V04_1),.clk(gclk));
	jdff dff_B_8jvt49m20_0(.din(n769),.dout(w_dff_B_8jvt49m20_0),.clk(gclk));
	jdff dff_B_y8kKgoeP1_0(.din(w_dff_B_8jvt49m20_0),.dout(w_dff_B_y8kKgoeP1_0),.clk(gclk));
	jdff dff_B_0dx886Ab3_0(.din(w_dff_B_y8kKgoeP1_0),.dout(w_dff_B_0dx886Ab3_0),.clk(gclk));
	jdff dff_B_sUlcGnsL9_0(.din(w_dff_B_0dx886Ab3_0),.dout(w_dff_B_sUlcGnsL9_0),.clk(gclk));
	jdff dff_B_Wa7HuQ6Q1_0(.din(w_dff_B_sUlcGnsL9_0),.dout(w_dff_B_Wa7HuQ6Q1_0),.clk(gclk));
	jdff dff_B_ZNWjGReA2_0(.din(w_dff_B_Wa7HuQ6Q1_0),.dout(w_dff_B_ZNWjGReA2_0),.clk(gclk));
	jdff dff_B_PAZl7fDR1_0(.din(w_dff_B_ZNWjGReA2_0),.dout(w_dff_B_PAZl7fDR1_0),.clk(gclk));
	jdff dff_B_32Fn1vWW5_0(.din(w_dff_B_PAZl7fDR1_0),.dout(w_dff_B_32Fn1vWW5_0),.clk(gclk));
	jdff dff_B_uc1vmQNc3_0(.din(w_dff_B_32Fn1vWW5_0),.dout(w_dff_B_uc1vmQNc3_0),.clk(gclk));
	jdff dff_B_AQwrQfHK9_0(.din(w_dff_B_uc1vmQNc3_0),.dout(w_dff_B_AQwrQfHK9_0),.clk(gclk));
	jdff dff_B_bC5jBocF6_0(.din(w_dff_B_AQwrQfHK9_0),.dout(w_dff_B_bC5jBocF6_0),.clk(gclk));
	jdff dff_B_ci4c5CF33_0(.din(w_dff_B_bC5jBocF6_0),.dout(w_dff_B_ci4c5CF33_0),.clk(gclk));
	jdff dff_B_nuzmbeWP1_0(.din(w_dff_B_ci4c5CF33_0),.dout(w_dff_B_nuzmbeWP1_0),.clk(gclk));
	jdff dff_B_B7Hw1spn0_0(.din(w_dff_B_nuzmbeWP1_0),.dout(w_dff_B_B7Hw1spn0_0),.clk(gclk));
	jdff dff_B_mlnM6kO62_0(.din(w_dff_B_B7Hw1spn0_0),.dout(w_dff_B_mlnM6kO62_0),.clk(gclk));
	jdff dff_B_EuUOriNB7_0(.din(w_dff_B_mlnM6kO62_0),.dout(w_dff_B_EuUOriNB7_0),.clk(gclk));
	jdff dff_B_gV2aYLZu5_0(.din(w_dff_B_EuUOriNB7_0),.dout(w_dff_B_gV2aYLZu5_0),.clk(gclk));
	jdff dff_B_SzQKEmyD2_0(.din(w_dff_B_gV2aYLZu5_0),.dout(w_dff_B_SzQKEmyD2_0),.clk(gclk));
	jdff dff_B_CTKMIZTy8_0(.din(w_dff_B_SzQKEmyD2_0),.dout(w_dff_B_CTKMIZTy8_0),.clk(gclk));
	jdff dff_B_3gdFVuvg4_0(.din(w_dff_B_CTKMIZTy8_0),.dout(w_dff_B_3gdFVuvg4_0),.clk(gclk));
	jdff dff_B_cewDTCxe9_0(.din(w_dff_B_3gdFVuvg4_0),.dout(w_dff_B_cewDTCxe9_0),.clk(gclk));
	jdff dff_B_XcDV76281_0(.din(w_dff_B_cewDTCxe9_0),.dout(w_dff_B_XcDV76281_0),.clk(gclk));
	jdff dff_B_zInW8uel6_0(.din(w_dff_B_XcDV76281_0),.dout(w_dff_B_zInW8uel6_0),.clk(gclk));
	jdff dff_B_180jp84y5_0(.din(w_dff_B_zInW8uel6_0),.dout(w_dff_B_180jp84y5_0),.clk(gclk));
	jdff dff_B_i6YDqOyM0_0(.din(w_dff_B_180jp84y5_0),.dout(w_dff_B_i6YDqOyM0_0),.clk(gclk));
	jdff dff_B_pSF9T5Pf2_0(.din(w_dff_B_i6YDqOyM0_0),.dout(w_dff_B_pSF9T5Pf2_0),.clk(gclk));
	jdff dff_B_bVFiigHL8_0(.din(w_dff_B_pSF9T5Pf2_0),.dout(w_dff_B_bVFiigHL8_0),.clk(gclk));
	jdff dff_B_lHP5kb4g2_0(.din(w_dff_B_bVFiigHL8_0),.dout(w_dff_B_lHP5kb4g2_0),.clk(gclk));
	jdff dff_B_dYhXjvMW5_0(.din(w_dff_B_lHP5kb4g2_0),.dout(w_dff_B_dYhXjvMW5_0),.clk(gclk));
	jdff dff_B_zV3Bh9KR9_0(.din(w_dff_B_dYhXjvMW5_0),.dout(w_dff_B_zV3Bh9KR9_0),.clk(gclk));
	jdff dff_B_p2uARIOa3_0(.din(w_dff_B_zV3Bh9KR9_0),.dout(w_dff_B_p2uARIOa3_0),.clk(gclk));
	jdff dff_B_PYTZ8VtL4_0(.din(w_dff_B_p2uARIOa3_0),.dout(w_dff_B_PYTZ8VtL4_0),.clk(gclk));
	jdff dff_B_EGkNCrWW0_0(.din(w_dff_B_PYTZ8VtL4_0),.dout(w_dff_B_EGkNCrWW0_0),.clk(gclk));
	jdff dff_B_SV1DUznb6_0(.din(w_dff_B_EGkNCrWW0_0),.dout(w_dff_B_SV1DUznb6_0),.clk(gclk));
	jdff dff_B_OOSxOqMm7_0(.din(w_dff_B_SV1DUznb6_0),.dout(w_dff_B_OOSxOqMm7_0),.clk(gclk));
	jdff dff_B_0TrsDzSo0_0(.din(w_dff_B_OOSxOqMm7_0),.dout(w_dff_B_0TrsDzSo0_0),.clk(gclk));
	jdff dff_B_sOPMhTBd5_0(.din(w_dff_B_0TrsDzSo0_0),.dout(w_dff_B_sOPMhTBd5_0),.clk(gclk));
	jdff dff_B_qRRGCDx71_0(.din(w_dff_B_sOPMhTBd5_0),.dout(w_dff_B_qRRGCDx71_0),.clk(gclk));
	jdff dff_B_kU4aM4Ij4_0(.din(w_dff_B_qRRGCDx71_0),.dout(w_dff_B_kU4aM4Ij4_0),.clk(gclk));
	jdff dff_B_isPekpHg1_0(.din(w_dff_B_kU4aM4Ij4_0),.dout(w_dff_B_isPekpHg1_0),.clk(gclk));
	jdff dff_B_sUxngRBc5_0(.din(w_dff_B_isPekpHg1_0),.dout(w_dff_B_sUxngRBc5_0),.clk(gclk));
	jdff dff_B_mO4k8g2u9_0(.din(w_dff_B_sUxngRBc5_0),.dout(w_dff_B_mO4k8g2u9_0),.clk(gclk));
	jdff dff_B_zaxnlJSa6_0(.din(w_dff_B_mO4k8g2u9_0),.dout(w_dff_B_zaxnlJSa6_0),.clk(gclk));
	jdff dff_B_xBDjz1107_0(.din(w_dff_B_zaxnlJSa6_0),.dout(w_dff_B_xBDjz1107_0),.clk(gclk));
	jdff dff_B_WGiSRHLC9_0(.din(w_dff_B_xBDjz1107_0),.dout(w_dff_B_WGiSRHLC9_0),.clk(gclk));
	jdff dff_B_SiXnnu6K5_0(.din(w_dff_B_WGiSRHLC9_0),.dout(w_dff_B_SiXnnu6K5_0),.clk(gclk));
	jdff dff_B_aXmc2KFr1_0(.din(w_dff_B_SiXnnu6K5_0),.dout(w_dff_B_aXmc2KFr1_0),.clk(gclk));
	jdff dff_B_XQ8nriLS7_0(.din(w_dff_B_aXmc2KFr1_0),.dout(w_dff_B_XQ8nriLS7_0),.clk(gclk));
	jdff dff_B_zELcjJ1u1_0(.din(w_dff_B_XQ8nriLS7_0),.dout(w_dff_B_zELcjJ1u1_0),.clk(gclk));
	jdff dff_B_F516xxhK4_0(.din(w_dff_B_zELcjJ1u1_0),.dout(w_dff_B_F516xxhK4_0),.clk(gclk));
	jdff dff_B_LN8GzzQ85_0(.din(w_dff_B_F516xxhK4_0),.dout(w_dff_B_LN8GzzQ85_0),.clk(gclk));
	jdff dff_B_SDd9pG3g6_0(.din(w_dff_B_LN8GzzQ85_0),.dout(w_dff_B_SDd9pG3g6_0),.clk(gclk));
	jdff dff_B_n2BpADnQ6_0(.din(w_dff_B_SDd9pG3g6_0),.dout(w_dff_B_n2BpADnQ6_0),.clk(gclk));
	jdff dff_B_hYq1GgVC3_0(.din(w_dff_B_n2BpADnQ6_0),.dout(w_dff_B_hYq1GgVC3_0),.clk(gclk));
	jdff dff_B_le5p1kjZ9_0(.din(w_dff_B_hYq1GgVC3_0),.dout(w_dff_B_le5p1kjZ9_0),.clk(gclk));
	jdff dff_B_JcQE2Eb47_0(.din(w_dff_B_le5p1kjZ9_0),.dout(w_dff_B_JcQE2Eb47_0),.clk(gclk));
	jdff dff_B_G0PReR3J0_0(.din(w_dff_B_JcQE2Eb47_0),.dout(w_dff_B_G0PReR3J0_0),.clk(gclk));
	jdff dff_B_9PGRykE52_0(.din(w_dff_B_G0PReR3J0_0),.dout(w_dff_B_9PGRykE52_0),.clk(gclk));
	jdff dff_B_UEunsgaB1_0(.din(w_dff_B_9PGRykE52_0),.dout(w_dff_B_UEunsgaB1_0),.clk(gclk));
	jdff dff_B_hx8YtgrH1_0(.din(w_dff_B_UEunsgaB1_0),.dout(w_dff_B_hx8YtgrH1_0),.clk(gclk));
	jdff dff_B_KuEIbo5y0_0(.din(w_dff_B_hx8YtgrH1_0),.dout(w_dff_B_KuEIbo5y0_0),.clk(gclk));
	jdff dff_B_kits9ir32_0(.din(w_dff_B_KuEIbo5y0_0),.dout(w_dff_B_kits9ir32_0),.clk(gclk));
	jdff dff_B_4e2hgKf74_0(.din(w_dff_B_kits9ir32_0),.dout(w_dff_B_4e2hgKf74_0),.clk(gclk));
	jdff dff_B_Xj7EsTj23_0(.din(w_dff_B_4e2hgKf74_0),.dout(w_dff_B_Xj7EsTj23_0),.clk(gclk));
	jdff dff_B_7cu7BDBS8_1(.din(n762),.dout(w_dff_B_7cu7BDBS8_1),.clk(gclk));
	jdff dff_B_uDqwjLj17_1(.din(w_dff_B_7cu7BDBS8_1),.dout(w_dff_B_uDqwjLj17_1),.clk(gclk));
	jdff dff_B_4Yb516S16_1(.din(w_dff_B_uDqwjLj17_1),.dout(w_dff_B_4Yb516S16_1),.clk(gclk));
	jdff dff_B_2YcgcUE42_1(.din(w_dff_B_4Yb516S16_1),.dout(w_dff_B_2YcgcUE42_1),.clk(gclk));
	jdff dff_B_odBgWBtx6_1(.din(w_dff_B_2YcgcUE42_1),.dout(w_dff_B_odBgWBtx6_1),.clk(gclk));
	jdff dff_B_cbCgOXKC4_1(.din(w_dff_B_odBgWBtx6_1),.dout(w_dff_B_cbCgOXKC4_1),.clk(gclk));
	jdff dff_B_vhwz3dOr6_1(.din(w_dff_B_cbCgOXKC4_1),.dout(w_dff_B_vhwz3dOr6_1),.clk(gclk));
	jdff dff_B_PsA58lrt6_1(.din(w_dff_B_vhwz3dOr6_1),.dout(w_dff_B_PsA58lrt6_1),.clk(gclk));
	jdff dff_B_imCIvpUZ8_1(.din(w_dff_B_PsA58lrt6_1),.dout(w_dff_B_imCIvpUZ8_1),.clk(gclk));
	jdff dff_B_IdW1OJU97_1(.din(w_dff_B_imCIvpUZ8_1),.dout(w_dff_B_IdW1OJU97_1),.clk(gclk));
	jdff dff_B_OsfbAIuW6_1(.din(w_dff_B_IdW1OJU97_1),.dout(w_dff_B_OsfbAIuW6_1),.clk(gclk));
	jdff dff_B_z2fJUlJw0_1(.din(w_dff_B_OsfbAIuW6_1),.dout(w_dff_B_z2fJUlJw0_1),.clk(gclk));
	jdff dff_B_XCUHLsZ74_1(.din(w_dff_B_z2fJUlJw0_1),.dout(w_dff_B_XCUHLsZ74_1),.clk(gclk));
	jdff dff_B_j9NGT5YK2_1(.din(w_dff_B_XCUHLsZ74_1),.dout(w_dff_B_j9NGT5YK2_1),.clk(gclk));
	jdff dff_B_IGRL3lqn4_1(.din(w_dff_B_j9NGT5YK2_1),.dout(w_dff_B_IGRL3lqn4_1),.clk(gclk));
	jdff dff_B_vXANSm6S1_1(.din(w_dff_B_IGRL3lqn4_1),.dout(w_dff_B_vXANSm6S1_1),.clk(gclk));
	jdff dff_B_gcJo1ROv2_1(.din(w_dff_B_vXANSm6S1_1),.dout(w_dff_B_gcJo1ROv2_1),.clk(gclk));
	jdff dff_B_CjMoUz0g9_1(.din(w_dff_B_gcJo1ROv2_1),.dout(w_dff_B_CjMoUz0g9_1),.clk(gclk));
	jdff dff_B_aZ8nqmGT8_1(.din(w_dff_B_CjMoUz0g9_1),.dout(w_dff_B_aZ8nqmGT8_1),.clk(gclk));
	jdff dff_B_A7PZ9GsO1_1(.din(w_dff_B_aZ8nqmGT8_1),.dout(w_dff_B_A7PZ9GsO1_1),.clk(gclk));
	jdff dff_B_iT5MW0qn5_1(.din(w_dff_B_A7PZ9GsO1_1),.dout(w_dff_B_iT5MW0qn5_1),.clk(gclk));
	jdff dff_B_n9Ig3jhR8_1(.din(w_dff_B_iT5MW0qn5_1),.dout(w_dff_B_n9Ig3jhR8_1),.clk(gclk));
	jdff dff_B_Cu5mas7q6_1(.din(w_dff_B_n9Ig3jhR8_1),.dout(w_dff_B_Cu5mas7q6_1),.clk(gclk));
	jdff dff_B_I65WPdcW8_1(.din(w_dff_B_Cu5mas7q6_1),.dout(w_dff_B_I65WPdcW8_1),.clk(gclk));
	jdff dff_B_kFN790u39_1(.din(w_dff_B_I65WPdcW8_1),.dout(w_dff_B_kFN790u39_1),.clk(gclk));
	jdff dff_B_S5lGZ8J95_1(.din(w_dff_B_kFN790u39_1),.dout(w_dff_B_S5lGZ8J95_1),.clk(gclk));
	jdff dff_B_uIpOpjSU2_1(.din(w_dff_B_S5lGZ8J95_1),.dout(w_dff_B_uIpOpjSU2_1),.clk(gclk));
	jdff dff_B_2Isikgdt0_1(.din(w_dff_B_uIpOpjSU2_1),.dout(w_dff_B_2Isikgdt0_1),.clk(gclk));
	jdff dff_B_1uaBUYjd8_1(.din(w_dff_B_2Isikgdt0_1),.dout(w_dff_B_1uaBUYjd8_1),.clk(gclk));
	jdff dff_B_6BWM4xHe6_1(.din(w_dff_B_1uaBUYjd8_1),.dout(w_dff_B_6BWM4xHe6_1),.clk(gclk));
	jdff dff_B_D2t2dySb7_1(.din(w_dff_B_6BWM4xHe6_1),.dout(w_dff_B_D2t2dySb7_1),.clk(gclk));
	jdff dff_B_z6WYQSXk4_1(.din(w_dff_B_D2t2dySb7_1),.dout(w_dff_B_z6WYQSXk4_1),.clk(gclk));
	jdff dff_B_JWFXxkoL4_1(.din(w_dff_B_z6WYQSXk4_1),.dout(w_dff_B_JWFXxkoL4_1),.clk(gclk));
	jdff dff_B_FDYeKO5A5_1(.din(w_dff_B_JWFXxkoL4_1),.dout(w_dff_B_FDYeKO5A5_1),.clk(gclk));
	jdff dff_B_c8TtplOB7_1(.din(w_dff_B_FDYeKO5A5_1),.dout(w_dff_B_c8TtplOB7_1),.clk(gclk));
	jdff dff_B_c0MzHVnU4_1(.din(w_dff_B_c8TtplOB7_1),.dout(w_dff_B_c0MzHVnU4_1),.clk(gclk));
	jdff dff_B_TPpuQTEn7_1(.din(w_dff_B_c0MzHVnU4_1),.dout(w_dff_B_TPpuQTEn7_1),.clk(gclk));
	jdff dff_B_BVr4Ymur2_1(.din(w_dff_B_TPpuQTEn7_1),.dout(w_dff_B_BVr4Ymur2_1),.clk(gclk));
	jdff dff_B_Cx89FCXi5_1(.din(w_dff_B_BVr4Ymur2_1),.dout(w_dff_B_Cx89FCXi5_1),.clk(gclk));
	jdff dff_B_2hlkU6Dy2_1(.din(w_dff_B_Cx89FCXi5_1),.dout(w_dff_B_2hlkU6Dy2_1),.clk(gclk));
	jdff dff_B_zwqOC2Hw2_1(.din(w_dff_B_2hlkU6Dy2_1),.dout(w_dff_B_zwqOC2Hw2_1),.clk(gclk));
	jdff dff_B_wuoZo4Q99_1(.din(w_dff_B_zwqOC2Hw2_1),.dout(w_dff_B_wuoZo4Q99_1),.clk(gclk));
	jdff dff_B_m0kHz9zy9_1(.din(w_dff_B_wuoZo4Q99_1),.dout(w_dff_B_m0kHz9zy9_1),.clk(gclk));
	jdff dff_B_oZnF0VNm8_1(.din(w_dff_B_m0kHz9zy9_1),.dout(w_dff_B_oZnF0VNm8_1),.clk(gclk));
	jdff dff_B_vaqKKXb76_1(.din(w_dff_B_oZnF0VNm8_1),.dout(w_dff_B_vaqKKXb76_1),.clk(gclk));
	jdff dff_B_n1oRl45p3_1(.din(w_dff_B_vaqKKXb76_1),.dout(w_dff_B_n1oRl45p3_1),.clk(gclk));
	jdff dff_B_VMz29ONC9_1(.din(w_dff_B_n1oRl45p3_1),.dout(w_dff_B_VMz29ONC9_1),.clk(gclk));
	jdff dff_B_bx9muena6_1(.din(w_dff_B_VMz29ONC9_1),.dout(w_dff_B_bx9muena6_1),.clk(gclk));
	jdff dff_B_0UuwdQhS5_1(.din(w_dff_B_bx9muena6_1),.dout(w_dff_B_0UuwdQhS5_1),.clk(gclk));
	jdff dff_B_1imDCN9U1_1(.din(w_dff_B_0UuwdQhS5_1),.dout(w_dff_B_1imDCN9U1_1),.clk(gclk));
	jdff dff_B_l6Oug9xJ1_1(.din(w_dff_B_1imDCN9U1_1),.dout(w_dff_B_l6Oug9xJ1_1),.clk(gclk));
	jdff dff_B_4fQmefUB9_1(.din(w_dff_B_l6Oug9xJ1_1),.dout(w_dff_B_4fQmefUB9_1),.clk(gclk));
	jdff dff_B_dKIuqhRF8_1(.din(w_dff_B_4fQmefUB9_1),.dout(w_dff_B_dKIuqhRF8_1),.clk(gclk));
	jdff dff_B_saMclL7J2_1(.din(w_dff_B_dKIuqhRF8_1),.dout(w_dff_B_saMclL7J2_1),.clk(gclk));
	jdff dff_B_M5nzTvhP9_1(.din(w_dff_B_saMclL7J2_1),.dout(w_dff_B_M5nzTvhP9_1),.clk(gclk));
	jdff dff_B_bvtfSewb1_1(.din(w_dff_B_M5nzTvhP9_1),.dout(w_dff_B_bvtfSewb1_1),.clk(gclk));
	jdff dff_B_15G1G7e40_1(.din(w_dff_B_bvtfSewb1_1),.dout(w_dff_B_15G1G7e40_1),.clk(gclk));
	jdff dff_B_XMoTTNRF2_1(.din(w_dff_B_15G1G7e40_1),.dout(w_dff_B_XMoTTNRF2_1),.clk(gclk));
	jdff dff_B_QcjToezX0_1(.din(w_dff_B_XMoTTNRF2_1),.dout(w_dff_B_QcjToezX0_1),.clk(gclk));
	jdff dff_B_mXyo8GpD5_1(.din(w_dff_B_QcjToezX0_1),.dout(w_dff_B_mXyo8GpD5_1),.clk(gclk));
	jdff dff_B_oyx70XJx7_1(.din(w_dff_B_mXyo8GpD5_1),.dout(w_dff_B_oyx70XJx7_1),.clk(gclk));
	jdff dff_B_4g3ciLln4_1(.din(w_dff_B_oyx70XJx7_1),.dout(w_dff_B_4g3ciLln4_1),.clk(gclk));
	jdff dff_B_HRhAL3Ck5_1(.din(w_dff_B_4g3ciLln4_1),.dout(w_dff_B_HRhAL3Ck5_1),.clk(gclk));
	jdff dff_B_Iq5SIEBg6_0(.din(n763),.dout(w_dff_B_Iq5SIEBg6_0),.clk(gclk));
	jdff dff_B_bmrF8RiS9_0(.din(w_dff_B_Iq5SIEBg6_0),.dout(w_dff_B_bmrF8RiS9_0),.clk(gclk));
	jdff dff_B_r7MNbbqV7_0(.din(w_dff_B_bmrF8RiS9_0),.dout(w_dff_B_r7MNbbqV7_0),.clk(gclk));
	jdff dff_B_gQHgiSjD3_0(.din(w_dff_B_r7MNbbqV7_0),.dout(w_dff_B_gQHgiSjD3_0),.clk(gclk));
	jdff dff_B_qnPmHTNX8_0(.din(w_dff_B_gQHgiSjD3_0),.dout(w_dff_B_qnPmHTNX8_0),.clk(gclk));
	jdff dff_B_TAEV7iu27_0(.din(w_dff_B_qnPmHTNX8_0),.dout(w_dff_B_TAEV7iu27_0),.clk(gclk));
	jdff dff_B_SZ66MXMF7_0(.din(w_dff_B_TAEV7iu27_0),.dout(w_dff_B_SZ66MXMF7_0),.clk(gclk));
	jdff dff_B_YHjvIQoi4_0(.din(w_dff_B_SZ66MXMF7_0),.dout(w_dff_B_YHjvIQoi4_0),.clk(gclk));
	jdff dff_B_xoksyxlb4_0(.din(w_dff_B_YHjvIQoi4_0),.dout(w_dff_B_xoksyxlb4_0),.clk(gclk));
	jdff dff_B_KvxheGpT2_0(.din(w_dff_B_xoksyxlb4_0),.dout(w_dff_B_KvxheGpT2_0),.clk(gclk));
	jdff dff_B_Ea58jBqh6_0(.din(w_dff_B_KvxheGpT2_0),.dout(w_dff_B_Ea58jBqh6_0),.clk(gclk));
	jdff dff_B_4Y4zcUxE3_0(.din(w_dff_B_Ea58jBqh6_0),.dout(w_dff_B_4Y4zcUxE3_0),.clk(gclk));
	jdff dff_B_2kjiat809_0(.din(w_dff_B_4Y4zcUxE3_0),.dout(w_dff_B_2kjiat809_0),.clk(gclk));
	jdff dff_B_I780kHOK0_0(.din(w_dff_B_2kjiat809_0),.dout(w_dff_B_I780kHOK0_0),.clk(gclk));
	jdff dff_B_7Xq193pV4_0(.din(w_dff_B_I780kHOK0_0),.dout(w_dff_B_7Xq193pV4_0),.clk(gclk));
	jdff dff_B_zNDcUXjD9_0(.din(w_dff_B_7Xq193pV4_0),.dout(w_dff_B_zNDcUXjD9_0),.clk(gclk));
	jdff dff_B_ZoZt7Vke9_0(.din(w_dff_B_zNDcUXjD9_0),.dout(w_dff_B_ZoZt7Vke9_0),.clk(gclk));
	jdff dff_B_yAXdDuId3_0(.din(w_dff_B_ZoZt7Vke9_0),.dout(w_dff_B_yAXdDuId3_0),.clk(gclk));
	jdff dff_B_FNPm2xdt1_0(.din(w_dff_B_yAXdDuId3_0),.dout(w_dff_B_FNPm2xdt1_0),.clk(gclk));
	jdff dff_B_MSY8yK4a2_0(.din(w_dff_B_FNPm2xdt1_0),.dout(w_dff_B_MSY8yK4a2_0),.clk(gclk));
	jdff dff_B_UllGlyU07_0(.din(w_dff_B_MSY8yK4a2_0),.dout(w_dff_B_UllGlyU07_0),.clk(gclk));
	jdff dff_B_yHPFuprz2_0(.din(w_dff_B_UllGlyU07_0),.dout(w_dff_B_yHPFuprz2_0),.clk(gclk));
	jdff dff_B_uT4LyiFS9_0(.din(w_dff_B_yHPFuprz2_0),.dout(w_dff_B_uT4LyiFS9_0),.clk(gclk));
	jdff dff_B_i90G6ENc0_0(.din(w_dff_B_uT4LyiFS9_0),.dout(w_dff_B_i90G6ENc0_0),.clk(gclk));
	jdff dff_B_2VnWw6Lw7_0(.din(w_dff_B_i90G6ENc0_0),.dout(w_dff_B_2VnWw6Lw7_0),.clk(gclk));
	jdff dff_B_dgSVkDSR7_0(.din(w_dff_B_2VnWw6Lw7_0),.dout(w_dff_B_dgSVkDSR7_0),.clk(gclk));
	jdff dff_B_yw9Aq1s27_0(.din(w_dff_B_dgSVkDSR7_0),.dout(w_dff_B_yw9Aq1s27_0),.clk(gclk));
	jdff dff_B_xiVuwzzH4_0(.din(w_dff_B_yw9Aq1s27_0),.dout(w_dff_B_xiVuwzzH4_0),.clk(gclk));
	jdff dff_B_ZOEY9g4g0_0(.din(w_dff_B_xiVuwzzH4_0),.dout(w_dff_B_ZOEY9g4g0_0),.clk(gclk));
	jdff dff_B_8yuHZmbB1_0(.din(w_dff_B_ZOEY9g4g0_0),.dout(w_dff_B_8yuHZmbB1_0),.clk(gclk));
	jdff dff_B_D11GE3nS0_0(.din(w_dff_B_8yuHZmbB1_0),.dout(w_dff_B_D11GE3nS0_0),.clk(gclk));
	jdff dff_B_6Di2tpgr8_0(.din(w_dff_B_D11GE3nS0_0),.dout(w_dff_B_6Di2tpgr8_0),.clk(gclk));
	jdff dff_B_gfZQfCSD6_0(.din(w_dff_B_6Di2tpgr8_0),.dout(w_dff_B_gfZQfCSD6_0),.clk(gclk));
	jdff dff_B_n1wrFb1w8_0(.din(w_dff_B_gfZQfCSD6_0),.dout(w_dff_B_n1wrFb1w8_0),.clk(gclk));
	jdff dff_B_cVAJMW9Z7_0(.din(w_dff_B_n1wrFb1w8_0),.dout(w_dff_B_cVAJMW9Z7_0),.clk(gclk));
	jdff dff_B_5E48SLub1_0(.din(w_dff_B_cVAJMW9Z7_0),.dout(w_dff_B_5E48SLub1_0),.clk(gclk));
	jdff dff_B_qsyeCCur8_0(.din(w_dff_B_5E48SLub1_0),.dout(w_dff_B_qsyeCCur8_0),.clk(gclk));
	jdff dff_B_8rvzTbZY2_0(.din(w_dff_B_qsyeCCur8_0),.dout(w_dff_B_8rvzTbZY2_0),.clk(gclk));
	jdff dff_B_gGh3ub9W9_0(.din(w_dff_B_8rvzTbZY2_0),.dout(w_dff_B_gGh3ub9W9_0),.clk(gclk));
	jdff dff_B_JtWItMy44_0(.din(w_dff_B_gGh3ub9W9_0),.dout(w_dff_B_JtWItMy44_0),.clk(gclk));
	jdff dff_B_CuhD3rm99_0(.din(w_dff_B_JtWItMy44_0),.dout(w_dff_B_CuhD3rm99_0),.clk(gclk));
	jdff dff_B_tpLSu2OR1_0(.din(w_dff_B_CuhD3rm99_0),.dout(w_dff_B_tpLSu2OR1_0),.clk(gclk));
	jdff dff_B_QSQ8UDAV1_0(.din(w_dff_B_tpLSu2OR1_0),.dout(w_dff_B_QSQ8UDAV1_0),.clk(gclk));
	jdff dff_B_GrGS9iFN1_0(.din(w_dff_B_QSQ8UDAV1_0),.dout(w_dff_B_GrGS9iFN1_0),.clk(gclk));
	jdff dff_B_MU7OR6QM1_0(.din(w_dff_B_GrGS9iFN1_0),.dout(w_dff_B_MU7OR6QM1_0),.clk(gclk));
	jdff dff_B_fflddMHi4_0(.din(w_dff_B_MU7OR6QM1_0),.dout(w_dff_B_fflddMHi4_0),.clk(gclk));
	jdff dff_B_1gjHNwWc6_0(.din(w_dff_B_fflddMHi4_0),.dout(w_dff_B_1gjHNwWc6_0),.clk(gclk));
	jdff dff_B_50W7jHId4_0(.din(w_dff_B_1gjHNwWc6_0),.dout(w_dff_B_50W7jHId4_0),.clk(gclk));
	jdff dff_B_D1TrHkD97_0(.din(w_dff_B_50W7jHId4_0),.dout(w_dff_B_D1TrHkD97_0),.clk(gclk));
	jdff dff_B_RqaAzPuO6_0(.din(w_dff_B_D1TrHkD97_0),.dout(w_dff_B_RqaAzPuO6_0),.clk(gclk));
	jdff dff_B_1FnkpiRx8_0(.din(w_dff_B_RqaAzPuO6_0),.dout(w_dff_B_1FnkpiRx8_0),.clk(gclk));
	jdff dff_B_TvPafgFc4_0(.din(w_dff_B_1FnkpiRx8_0),.dout(w_dff_B_TvPafgFc4_0),.clk(gclk));
	jdff dff_B_oRv6gGLj3_0(.din(w_dff_B_TvPafgFc4_0),.dout(w_dff_B_oRv6gGLj3_0),.clk(gclk));
	jdff dff_B_FZhMXYUO1_0(.din(w_dff_B_oRv6gGLj3_0),.dout(w_dff_B_FZhMXYUO1_0),.clk(gclk));
	jdff dff_B_AvlaCdJf9_0(.din(w_dff_B_FZhMXYUO1_0),.dout(w_dff_B_AvlaCdJf9_0),.clk(gclk));
	jdff dff_B_IGcHJelU4_0(.din(w_dff_B_AvlaCdJf9_0),.dout(w_dff_B_IGcHJelU4_0),.clk(gclk));
	jdff dff_B_C1ixfA4R2_0(.din(w_dff_B_IGcHJelU4_0),.dout(w_dff_B_C1ixfA4R2_0),.clk(gclk));
	jdff dff_B_dnzUGiSt8_0(.din(w_dff_B_C1ixfA4R2_0),.dout(w_dff_B_dnzUGiSt8_0),.clk(gclk));
	jdff dff_B_6qouszEI7_0(.din(w_dff_B_dnzUGiSt8_0),.dout(w_dff_B_6qouszEI7_0),.clk(gclk));
	jdff dff_B_ouioeusH9_0(.din(w_dff_B_6qouszEI7_0),.dout(w_dff_B_ouioeusH9_0),.clk(gclk));
	jdff dff_B_er01xbRt3_0(.din(w_dff_B_ouioeusH9_0),.dout(w_dff_B_er01xbRt3_0),.clk(gclk));
	jdff dff_B_pzmkeITL1_0(.din(w_dff_B_er01xbRt3_0),.dout(w_dff_B_pzmkeITL1_0),.clk(gclk));
	jdff dff_B_J5sqkVLr6_0(.din(w_dff_B_pzmkeITL1_0),.dout(w_dff_B_J5sqkVLr6_0),.clk(gclk));
	jdff dff_B_pCM6Lm6q5_1(.din(n756),.dout(w_dff_B_pCM6Lm6q5_1),.clk(gclk));
	jdff dff_B_6g0XpZPS6_1(.din(w_dff_B_pCM6Lm6q5_1),.dout(w_dff_B_6g0XpZPS6_1),.clk(gclk));
	jdff dff_B_HIcw1Ujt6_1(.din(w_dff_B_6g0XpZPS6_1),.dout(w_dff_B_HIcw1Ujt6_1),.clk(gclk));
	jdff dff_B_JSWdv6P78_1(.din(w_dff_B_HIcw1Ujt6_1),.dout(w_dff_B_JSWdv6P78_1),.clk(gclk));
	jdff dff_B_q0KVr8gt5_1(.din(w_dff_B_JSWdv6P78_1),.dout(w_dff_B_q0KVr8gt5_1),.clk(gclk));
	jdff dff_B_FAsyEvzp0_1(.din(w_dff_B_q0KVr8gt5_1),.dout(w_dff_B_FAsyEvzp0_1),.clk(gclk));
	jdff dff_B_FJCFVEKQ8_1(.din(w_dff_B_FAsyEvzp0_1),.dout(w_dff_B_FJCFVEKQ8_1),.clk(gclk));
	jdff dff_B_4OO3EZD56_1(.din(w_dff_B_FJCFVEKQ8_1),.dout(w_dff_B_4OO3EZD56_1),.clk(gclk));
	jdff dff_B_RyX0zQpk7_1(.din(w_dff_B_4OO3EZD56_1),.dout(w_dff_B_RyX0zQpk7_1),.clk(gclk));
	jdff dff_B_zeC7bnIP2_1(.din(w_dff_B_RyX0zQpk7_1),.dout(w_dff_B_zeC7bnIP2_1),.clk(gclk));
	jdff dff_B_TnpxSOum1_1(.din(w_dff_B_zeC7bnIP2_1),.dout(w_dff_B_TnpxSOum1_1),.clk(gclk));
	jdff dff_B_M3WoWmAY6_1(.din(w_dff_B_TnpxSOum1_1),.dout(w_dff_B_M3WoWmAY6_1),.clk(gclk));
	jdff dff_B_4MO54Gg99_1(.din(w_dff_B_M3WoWmAY6_1),.dout(w_dff_B_4MO54Gg99_1),.clk(gclk));
	jdff dff_B_kJHuamjg4_1(.din(w_dff_B_4MO54Gg99_1),.dout(w_dff_B_kJHuamjg4_1),.clk(gclk));
	jdff dff_B_AZrgnmcb3_1(.din(w_dff_B_kJHuamjg4_1),.dout(w_dff_B_AZrgnmcb3_1),.clk(gclk));
	jdff dff_B_WsjUi3Z02_1(.din(w_dff_B_AZrgnmcb3_1),.dout(w_dff_B_WsjUi3Z02_1),.clk(gclk));
	jdff dff_B_wnGOngvr1_1(.din(w_dff_B_WsjUi3Z02_1),.dout(w_dff_B_wnGOngvr1_1),.clk(gclk));
	jdff dff_B_4o4fRPLS7_1(.din(w_dff_B_wnGOngvr1_1),.dout(w_dff_B_4o4fRPLS7_1),.clk(gclk));
	jdff dff_B_GffUK5y29_1(.din(w_dff_B_4o4fRPLS7_1),.dout(w_dff_B_GffUK5y29_1),.clk(gclk));
	jdff dff_B_r3xQzSi28_1(.din(w_dff_B_GffUK5y29_1),.dout(w_dff_B_r3xQzSi28_1),.clk(gclk));
	jdff dff_B_G4vRyjta4_1(.din(w_dff_B_r3xQzSi28_1),.dout(w_dff_B_G4vRyjta4_1),.clk(gclk));
	jdff dff_B_SoEiGnIc9_1(.din(w_dff_B_G4vRyjta4_1),.dout(w_dff_B_SoEiGnIc9_1),.clk(gclk));
	jdff dff_B_cSy2rZTF5_1(.din(w_dff_B_SoEiGnIc9_1),.dout(w_dff_B_cSy2rZTF5_1),.clk(gclk));
	jdff dff_B_jcpNYGoa8_1(.din(w_dff_B_cSy2rZTF5_1),.dout(w_dff_B_jcpNYGoa8_1),.clk(gclk));
	jdff dff_B_V7x0HHom5_1(.din(w_dff_B_jcpNYGoa8_1),.dout(w_dff_B_V7x0HHom5_1),.clk(gclk));
	jdff dff_B_YhIb3nKD3_1(.din(w_dff_B_V7x0HHom5_1),.dout(w_dff_B_YhIb3nKD3_1),.clk(gclk));
	jdff dff_B_BSNDtTVs0_1(.din(w_dff_B_YhIb3nKD3_1),.dout(w_dff_B_BSNDtTVs0_1),.clk(gclk));
	jdff dff_B_8fXS1JJJ3_1(.din(w_dff_B_BSNDtTVs0_1),.dout(w_dff_B_8fXS1JJJ3_1),.clk(gclk));
	jdff dff_B_bgE0axYw4_1(.din(w_dff_B_8fXS1JJJ3_1),.dout(w_dff_B_bgE0axYw4_1),.clk(gclk));
	jdff dff_B_5wZkBvJB4_1(.din(w_dff_B_bgE0axYw4_1),.dout(w_dff_B_5wZkBvJB4_1),.clk(gclk));
	jdff dff_B_TSyG6yGQ7_1(.din(w_dff_B_5wZkBvJB4_1),.dout(w_dff_B_TSyG6yGQ7_1),.clk(gclk));
	jdff dff_B_GnSoo2yZ0_1(.din(w_dff_B_TSyG6yGQ7_1),.dout(w_dff_B_GnSoo2yZ0_1),.clk(gclk));
	jdff dff_B_ApU1RraW2_1(.din(w_dff_B_GnSoo2yZ0_1),.dout(w_dff_B_ApU1RraW2_1),.clk(gclk));
	jdff dff_B_dXxRocCG3_1(.din(w_dff_B_ApU1RraW2_1),.dout(w_dff_B_dXxRocCG3_1),.clk(gclk));
	jdff dff_B_NyCSVVwW0_1(.din(w_dff_B_dXxRocCG3_1),.dout(w_dff_B_NyCSVVwW0_1),.clk(gclk));
	jdff dff_B_SkTkYTez9_1(.din(w_dff_B_NyCSVVwW0_1),.dout(w_dff_B_SkTkYTez9_1),.clk(gclk));
	jdff dff_B_ThLrF0L50_1(.din(w_dff_B_SkTkYTez9_1),.dout(w_dff_B_ThLrF0L50_1),.clk(gclk));
	jdff dff_B_EGNoTHZr6_1(.din(w_dff_B_ThLrF0L50_1),.dout(w_dff_B_EGNoTHZr6_1),.clk(gclk));
	jdff dff_B_iAAgjrVY4_1(.din(w_dff_B_EGNoTHZr6_1),.dout(w_dff_B_iAAgjrVY4_1),.clk(gclk));
	jdff dff_B_Ch9Js3uL3_1(.din(w_dff_B_iAAgjrVY4_1),.dout(w_dff_B_Ch9Js3uL3_1),.clk(gclk));
	jdff dff_B_BJJQJOLT0_1(.din(w_dff_B_Ch9Js3uL3_1),.dout(w_dff_B_BJJQJOLT0_1),.clk(gclk));
	jdff dff_B_COHzw3Zv6_1(.din(w_dff_B_BJJQJOLT0_1),.dout(w_dff_B_COHzw3Zv6_1),.clk(gclk));
	jdff dff_B_QireFWjw0_1(.din(w_dff_B_COHzw3Zv6_1),.dout(w_dff_B_QireFWjw0_1),.clk(gclk));
	jdff dff_B_iDWWtNtt6_1(.din(w_dff_B_QireFWjw0_1),.dout(w_dff_B_iDWWtNtt6_1),.clk(gclk));
	jdff dff_B_NwnT28Ys4_1(.din(w_dff_B_iDWWtNtt6_1),.dout(w_dff_B_NwnT28Ys4_1),.clk(gclk));
	jdff dff_B_8w4rU8iO1_1(.din(w_dff_B_NwnT28Ys4_1),.dout(w_dff_B_8w4rU8iO1_1),.clk(gclk));
	jdff dff_B_Nnsn6uhN7_1(.din(w_dff_B_8w4rU8iO1_1),.dout(w_dff_B_Nnsn6uhN7_1),.clk(gclk));
	jdff dff_B_sTCo5yyV6_1(.din(w_dff_B_Nnsn6uhN7_1),.dout(w_dff_B_sTCo5yyV6_1),.clk(gclk));
	jdff dff_B_JfrxKUFD2_1(.din(w_dff_B_sTCo5yyV6_1),.dout(w_dff_B_JfrxKUFD2_1),.clk(gclk));
	jdff dff_B_hFcX7sdE2_1(.din(w_dff_B_JfrxKUFD2_1),.dout(w_dff_B_hFcX7sdE2_1),.clk(gclk));
	jdff dff_B_0Eg3HpmP6_1(.din(w_dff_B_hFcX7sdE2_1),.dout(w_dff_B_0Eg3HpmP6_1),.clk(gclk));
	jdff dff_B_XiZ30F528_1(.din(w_dff_B_0Eg3HpmP6_1),.dout(w_dff_B_XiZ30F528_1),.clk(gclk));
	jdff dff_B_SkJKHoaU3_1(.din(w_dff_B_XiZ30F528_1),.dout(w_dff_B_SkJKHoaU3_1),.clk(gclk));
	jdff dff_B_vkt6hixL8_1(.din(w_dff_B_SkJKHoaU3_1),.dout(w_dff_B_vkt6hixL8_1),.clk(gclk));
	jdff dff_B_8C6yja3S5_1(.din(w_dff_B_vkt6hixL8_1),.dout(w_dff_B_8C6yja3S5_1),.clk(gclk));
	jdff dff_B_L2a0jLLv7_1(.din(w_dff_B_8C6yja3S5_1),.dout(w_dff_B_L2a0jLLv7_1),.clk(gclk));
	jdff dff_B_3DIWUwOC8_1(.din(w_dff_B_L2a0jLLv7_1),.dout(w_dff_B_3DIWUwOC8_1),.clk(gclk));
	jdff dff_B_dsiL7QO31_1(.din(w_dff_B_3DIWUwOC8_1),.dout(w_dff_B_dsiL7QO31_1),.clk(gclk));
	jdff dff_B_bZkssdEr2_1(.din(w_dff_B_dsiL7QO31_1),.dout(w_dff_B_bZkssdEr2_1),.clk(gclk));
	jdff dff_B_AoekRums7_1(.din(w_dff_B_bZkssdEr2_1),.dout(w_dff_B_AoekRums7_1),.clk(gclk));
	jdff dff_B_uPtNt3TD0_1(.din(w_dff_B_AoekRums7_1),.dout(w_dff_B_uPtNt3TD0_1),.clk(gclk));
	jdff dff_B_cMTGAhWx0_1(.din(w_dff_B_uPtNt3TD0_1),.dout(w_dff_B_cMTGAhWx0_1),.clk(gclk));
	jdff dff_B_Gb948lxH1_0(.din(n757),.dout(w_dff_B_Gb948lxH1_0),.clk(gclk));
	jdff dff_B_xCgC25rv5_0(.din(w_dff_B_Gb948lxH1_0),.dout(w_dff_B_xCgC25rv5_0),.clk(gclk));
	jdff dff_B_0T5yJljr6_0(.din(w_dff_B_xCgC25rv5_0),.dout(w_dff_B_0T5yJljr6_0),.clk(gclk));
	jdff dff_B_Cx6GdO1b6_0(.din(w_dff_B_0T5yJljr6_0),.dout(w_dff_B_Cx6GdO1b6_0),.clk(gclk));
	jdff dff_B_9FA9bqwa3_0(.din(w_dff_B_Cx6GdO1b6_0),.dout(w_dff_B_9FA9bqwa3_0),.clk(gclk));
	jdff dff_B_omhxUjMQ2_0(.din(w_dff_B_9FA9bqwa3_0),.dout(w_dff_B_omhxUjMQ2_0),.clk(gclk));
	jdff dff_B_RWbulGMU8_0(.din(w_dff_B_omhxUjMQ2_0),.dout(w_dff_B_RWbulGMU8_0),.clk(gclk));
	jdff dff_B_biOsRHvH5_0(.din(w_dff_B_RWbulGMU8_0),.dout(w_dff_B_biOsRHvH5_0),.clk(gclk));
	jdff dff_B_AajU3Poq2_0(.din(w_dff_B_biOsRHvH5_0),.dout(w_dff_B_AajU3Poq2_0),.clk(gclk));
	jdff dff_B_9k83aELm8_0(.din(w_dff_B_AajU3Poq2_0),.dout(w_dff_B_9k83aELm8_0),.clk(gclk));
	jdff dff_B_twXb4y336_0(.din(w_dff_B_9k83aELm8_0),.dout(w_dff_B_twXb4y336_0),.clk(gclk));
	jdff dff_B_nwoVfyvi7_0(.din(w_dff_B_twXb4y336_0),.dout(w_dff_B_nwoVfyvi7_0),.clk(gclk));
	jdff dff_B_oTNcbAP31_0(.din(w_dff_B_nwoVfyvi7_0),.dout(w_dff_B_oTNcbAP31_0),.clk(gclk));
	jdff dff_B_Mluztiq98_0(.din(w_dff_B_oTNcbAP31_0),.dout(w_dff_B_Mluztiq98_0),.clk(gclk));
	jdff dff_B_NkpLAXM08_0(.din(w_dff_B_Mluztiq98_0),.dout(w_dff_B_NkpLAXM08_0),.clk(gclk));
	jdff dff_B_2Oxc3Bb70_0(.din(w_dff_B_NkpLAXM08_0),.dout(w_dff_B_2Oxc3Bb70_0),.clk(gclk));
	jdff dff_B_fcvkr44d8_0(.din(w_dff_B_2Oxc3Bb70_0),.dout(w_dff_B_fcvkr44d8_0),.clk(gclk));
	jdff dff_B_GZpZuG998_0(.din(w_dff_B_fcvkr44d8_0),.dout(w_dff_B_GZpZuG998_0),.clk(gclk));
	jdff dff_B_7bd4c1KM4_0(.din(w_dff_B_GZpZuG998_0),.dout(w_dff_B_7bd4c1KM4_0),.clk(gclk));
	jdff dff_B_g3XloexJ9_0(.din(w_dff_B_7bd4c1KM4_0),.dout(w_dff_B_g3XloexJ9_0),.clk(gclk));
	jdff dff_B_zHKfXbTo6_0(.din(w_dff_B_g3XloexJ9_0),.dout(w_dff_B_zHKfXbTo6_0),.clk(gclk));
	jdff dff_B_L79zxG8M9_0(.din(w_dff_B_zHKfXbTo6_0),.dout(w_dff_B_L79zxG8M9_0),.clk(gclk));
	jdff dff_B_H7AFWyFd4_0(.din(w_dff_B_L79zxG8M9_0),.dout(w_dff_B_H7AFWyFd4_0),.clk(gclk));
	jdff dff_B_MI2VsTuJ0_0(.din(w_dff_B_H7AFWyFd4_0),.dout(w_dff_B_MI2VsTuJ0_0),.clk(gclk));
	jdff dff_B_R5A55xmn6_0(.din(w_dff_B_MI2VsTuJ0_0),.dout(w_dff_B_R5A55xmn6_0),.clk(gclk));
	jdff dff_B_bocE3cjN9_0(.din(w_dff_B_R5A55xmn6_0),.dout(w_dff_B_bocE3cjN9_0),.clk(gclk));
	jdff dff_B_3iMJ1vi79_0(.din(w_dff_B_bocE3cjN9_0),.dout(w_dff_B_3iMJ1vi79_0),.clk(gclk));
	jdff dff_B_XH7l6pFw1_0(.din(w_dff_B_3iMJ1vi79_0),.dout(w_dff_B_XH7l6pFw1_0),.clk(gclk));
	jdff dff_B_xkz7X7su9_0(.din(w_dff_B_XH7l6pFw1_0),.dout(w_dff_B_xkz7X7su9_0),.clk(gclk));
	jdff dff_B_P7Ttqsm60_0(.din(w_dff_B_xkz7X7su9_0),.dout(w_dff_B_P7Ttqsm60_0),.clk(gclk));
	jdff dff_B_r78hXM8n4_0(.din(w_dff_B_P7Ttqsm60_0),.dout(w_dff_B_r78hXM8n4_0),.clk(gclk));
	jdff dff_B_QnUHT7aa9_0(.din(w_dff_B_r78hXM8n4_0),.dout(w_dff_B_QnUHT7aa9_0),.clk(gclk));
	jdff dff_B_Aaj1fTkD9_0(.din(w_dff_B_QnUHT7aa9_0),.dout(w_dff_B_Aaj1fTkD9_0),.clk(gclk));
	jdff dff_B_NiN5AGtF5_0(.din(w_dff_B_Aaj1fTkD9_0),.dout(w_dff_B_NiN5AGtF5_0),.clk(gclk));
	jdff dff_B_wlC7SorM1_0(.din(w_dff_B_NiN5AGtF5_0),.dout(w_dff_B_wlC7SorM1_0),.clk(gclk));
	jdff dff_B_eSmT3Kxy0_0(.din(w_dff_B_wlC7SorM1_0),.dout(w_dff_B_eSmT3Kxy0_0),.clk(gclk));
	jdff dff_B_En9mGDM56_0(.din(w_dff_B_eSmT3Kxy0_0),.dout(w_dff_B_En9mGDM56_0),.clk(gclk));
	jdff dff_B_JU8Pvl128_0(.din(w_dff_B_En9mGDM56_0),.dout(w_dff_B_JU8Pvl128_0),.clk(gclk));
	jdff dff_B_qUFc0Ed45_0(.din(w_dff_B_JU8Pvl128_0),.dout(w_dff_B_qUFc0Ed45_0),.clk(gclk));
	jdff dff_B_JPN8PLhI2_0(.din(w_dff_B_qUFc0Ed45_0),.dout(w_dff_B_JPN8PLhI2_0),.clk(gclk));
	jdff dff_B_IMtlwL1c8_0(.din(w_dff_B_JPN8PLhI2_0),.dout(w_dff_B_IMtlwL1c8_0),.clk(gclk));
	jdff dff_B_U9HNst065_0(.din(w_dff_B_IMtlwL1c8_0),.dout(w_dff_B_U9HNst065_0),.clk(gclk));
	jdff dff_B_W0AM2YSI3_0(.din(w_dff_B_U9HNst065_0),.dout(w_dff_B_W0AM2YSI3_0),.clk(gclk));
	jdff dff_B_NiNbrwPS6_0(.din(w_dff_B_W0AM2YSI3_0),.dout(w_dff_B_NiNbrwPS6_0),.clk(gclk));
	jdff dff_B_qPNot8fL7_0(.din(w_dff_B_NiNbrwPS6_0),.dout(w_dff_B_qPNot8fL7_0),.clk(gclk));
	jdff dff_B_bTkhISM76_0(.din(w_dff_B_qPNot8fL7_0),.dout(w_dff_B_bTkhISM76_0),.clk(gclk));
	jdff dff_B_3zXwjCk84_0(.din(w_dff_B_bTkhISM76_0),.dout(w_dff_B_3zXwjCk84_0),.clk(gclk));
	jdff dff_B_qSeJNasX3_0(.din(w_dff_B_3zXwjCk84_0),.dout(w_dff_B_qSeJNasX3_0),.clk(gclk));
	jdff dff_B_VsC3ZK6P6_0(.din(w_dff_B_qSeJNasX3_0),.dout(w_dff_B_VsC3ZK6P6_0),.clk(gclk));
	jdff dff_B_mbanrVUj6_0(.din(w_dff_B_VsC3ZK6P6_0),.dout(w_dff_B_mbanrVUj6_0),.clk(gclk));
	jdff dff_B_mKZRQVP83_0(.din(w_dff_B_mbanrVUj6_0),.dout(w_dff_B_mKZRQVP83_0),.clk(gclk));
	jdff dff_B_ukn8lQJC0_0(.din(w_dff_B_mKZRQVP83_0),.dout(w_dff_B_ukn8lQJC0_0),.clk(gclk));
	jdff dff_B_07t8K00Q6_0(.din(w_dff_B_ukn8lQJC0_0),.dout(w_dff_B_07t8K00Q6_0),.clk(gclk));
	jdff dff_B_ln577FH27_0(.din(w_dff_B_07t8K00Q6_0),.dout(w_dff_B_ln577FH27_0),.clk(gclk));
	jdff dff_B_wAbb5i1f6_0(.din(w_dff_B_ln577FH27_0),.dout(w_dff_B_wAbb5i1f6_0),.clk(gclk));
	jdff dff_B_PggIU1MR3_0(.din(w_dff_B_wAbb5i1f6_0),.dout(w_dff_B_PggIU1MR3_0),.clk(gclk));
	jdff dff_B_csLlCdeo0_0(.din(w_dff_B_PggIU1MR3_0),.dout(w_dff_B_csLlCdeo0_0),.clk(gclk));
	jdff dff_B_1wKRBaic4_0(.din(w_dff_B_csLlCdeo0_0),.dout(w_dff_B_1wKRBaic4_0),.clk(gclk));
	jdff dff_B_A5xpSkoS7_0(.din(w_dff_B_1wKRBaic4_0),.dout(w_dff_B_A5xpSkoS7_0),.clk(gclk));
	jdff dff_B_D316AO3t0_0(.din(w_dff_B_A5xpSkoS7_0),.dout(w_dff_B_D316AO3t0_0),.clk(gclk));
	jdff dff_B_M4MGvFqE3_0(.din(w_dff_B_D316AO3t0_0),.dout(w_dff_B_M4MGvFqE3_0),.clk(gclk));
	jdff dff_B_fIXrmCN75_0(.din(w_dff_B_M4MGvFqE3_0),.dout(w_dff_B_fIXrmCN75_0),.clk(gclk));
	jdff dff_B_cJXCeA0y1_1(.din(n750),.dout(w_dff_B_cJXCeA0y1_1),.clk(gclk));
	jdff dff_B_59HshVZs5_1(.din(w_dff_B_cJXCeA0y1_1),.dout(w_dff_B_59HshVZs5_1),.clk(gclk));
	jdff dff_B_7TbwzYyW6_1(.din(w_dff_B_59HshVZs5_1),.dout(w_dff_B_7TbwzYyW6_1),.clk(gclk));
	jdff dff_B_VYJOMNCg2_1(.din(w_dff_B_7TbwzYyW6_1),.dout(w_dff_B_VYJOMNCg2_1),.clk(gclk));
	jdff dff_B_zyAYYDJ41_1(.din(w_dff_B_VYJOMNCg2_1),.dout(w_dff_B_zyAYYDJ41_1),.clk(gclk));
	jdff dff_B_KEu0eFlD6_1(.din(w_dff_B_zyAYYDJ41_1),.dout(w_dff_B_KEu0eFlD6_1),.clk(gclk));
	jdff dff_B_z3BTkWCm6_1(.din(w_dff_B_KEu0eFlD6_1),.dout(w_dff_B_z3BTkWCm6_1),.clk(gclk));
	jdff dff_B_IEYnuEbp6_1(.din(w_dff_B_z3BTkWCm6_1),.dout(w_dff_B_IEYnuEbp6_1),.clk(gclk));
	jdff dff_B_WocVIAZP4_1(.din(w_dff_B_IEYnuEbp6_1),.dout(w_dff_B_WocVIAZP4_1),.clk(gclk));
	jdff dff_B_16KqC2lq3_1(.din(w_dff_B_WocVIAZP4_1),.dout(w_dff_B_16KqC2lq3_1),.clk(gclk));
	jdff dff_B_f52Galrs2_1(.din(w_dff_B_16KqC2lq3_1),.dout(w_dff_B_f52Galrs2_1),.clk(gclk));
	jdff dff_B_79iSBHbn9_1(.din(w_dff_B_f52Galrs2_1),.dout(w_dff_B_79iSBHbn9_1),.clk(gclk));
	jdff dff_B_MREGjirp4_1(.din(w_dff_B_79iSBHbn9_1),.dout(w_dff_B_MREGjirp4_1),.clk(gclk));
	jdff dff_B_lcyCrvdg1_1(.din(w_dff_B_MREGjirp4_1),.dout(w_dff_B_lcyCrvdg1_1),.clk(gclk));
	jdff dff_B_cjHB07l78_1(.din(w_dff_B_lcyCrvdg1_1),.dout(w_dff_B_cjHB07l78_1),.clk(gclk));
	jdff dff_B_cQVTuwlt3_1(.din(w_dff_B_cjHB07l78_1),.dout(w_dff_B_cQVTuwlt3_1),.clk(gclk));
	jdff dff_B_NFXRdkBp2_1(.din(w_dff_B_cQVTuwlt3_1),.dout(w_dff_B_NFXRdkBp2_1),.clk(gclk));
	jdff dff_B_bw4tAdz56_1(.din(w_dff_B_NFXRdkBp2_1),.dout(w_dff_B_bw4tAdz56_1),.clk(gclk));
	jdff dff_B_MmC0O3Jy9_1(.din(w_dff_B_bw4tAdz56_1),.dout(w_dff_B_MmC0O3Jy9_1),.clk(gclk));
	jdff dff_B_2m4yg1en4_1(.din(w_dff_B_MmC0O3Jy9_1),.dout(w_dff_B_2m4yg1en4_1),.clk(gclk));
	jdff dff_B_b9Pjx3a21_1(.din(w_dff_B_2m4yg1en4_1),.dout(w_dff_B_b9Pjx3a21_1),.clk(gclk));
	jdff dff_B_MCwlDmhL0_1(.din(w_dff_B_b9Pjx3a21_1),.dout(w_dff_B_MCwlDmhL0_1),.clk(gclk));
	jdff dff_B_HkRpkuox2_1(.din(w_dff_B_MCwlDmhL0_1),.dout(w_dff_B_HkRpkuox2_1),.clk(gclk));
	jdff dff_B_3EPNxRK11_1(.din(w_dff_B_HkRpkuox2_1),.dout(w_dff_B_3EPNxRK11_1),.clk(gclk));
	jdff dff_B_kMm4iLo02_1(.din(w_dff_B_3EPNxRK11_1),.dout(w_dff_B_kMm4iLo02_1),.clk(gclk));
	jdff dff_B_mwm4f3jj5_1(.din(w_dff_B_kMm4iLo02_1),.dout(w_dff_B_mwm4f3jj5_1),.clk(gclk));
	jdff dff_B_2Z2DBqI25_1(.din(w_dff_B_mwm4f3jj5_1),.dout(w_dff_B_2Z2DBqI25_1),.clk(gclk));
	jdff dff_B_AMwvfgvg0_1(.din(w_dff_B_2Z2DBqI25_1),.dout(w_dff_B_AMwvfgvg0_1),.clk(gclk));
	jdff dff_B_Lm7HFJFP8_1(.din(w_dff_B_AMwvfgvg0_1),.dout(w_dff_B_Lm7HFJFP8_1),.clk(gclk));
	jdff dff_B_CocpBhrM1_1(.din(w_dff_B_Lm7HFJFP8_1),.dout(w_dff_B_CocpBhrM1_1),.clk(gclk));
	jdff dff_B_bTMeguTl4_1(.din(w_dff_B_CocpBhrM1_1),.dout(w_dff_B_bTMeguTl4_1),.clk(gclk));
	jdff dff_B_dbV42ggt3_1(.din(w_dff_B_bTMeguTl4_1),.dout(w_dff_B_dbV42ggt3_1),.clk(gclk));
	jdff dff_B_X5Nj5lhu8_1(.din(w_dff_B_dbV42ggt3_1),.dout(w_dff_B_X5Nj5lhu8_1),.clk(gclk));
	jdff dff_B_3TZnnSnD0_1(.din(w_dff_B_X5Nj5lhu8_1),.dout(w_dff_B_3TZnnSnD0_1),.clk(gclk));
	jdff dff_B_7qc1KcHe9_1(.din(w_dff_B_3TZnnSnD0_1),.dout(w_dff_B_7qc1KcHe9_1),.clk(gclk));
	jdff dff_B_gnWiF34h1_1(.din(w_dff_B_7qc1KcHe9_1),.dout(w_dff_B_gnWiF34h1_1),.clk(gclk));
	jdff dff_B_6GIRifoM8_1(.din(w_dff_B_gnWiF34h1_1),.dout(w_dff_B_6GIRifoM8_1),.clk(gclk));
	jdff dff_B_HhwQyiw53_1(.din(w_dff_B_6GIRifoM8_1),.dout(w_dff_B_HhwQyiw53_1),.clk(gclk));
	jdff dff_B_3txzdJ769_1(.din(w_dff_B_HhwQyiw53_1),.dout(w_dff_B_3txzdJ769_1),.clk(gclk));
	jdff dff_B_Vz5VF6nz6_1(.din(w_dff_B_3txzdJ769_1),.dout(w_dff_B_Vz5VF6nz6_1),.clk(gclk));
	jdff dff_B_KLbxjjcm3_1(.din(w_dff_B_Vz5VF6nz6_1),.dout(w_dff_B_KLbxjjcm3_1),.clk(gclk));
	jdff dff_B_phGo1tTR9_1(.din(w_dff_B_KLbxjjcm3_1),.dout(w_dff_B_phGo1tTR9_1),.clk(gclk));
	jdff dff_B_yTcGv9Tp8_1(.din(w_dff_B_phGo1tTR9_1),.dout(w_dff_B_yTcGv9Tp8_1),.clk(gclk));
	jdff dff_B_SShyMNgN8_1(.din(w_dff_B_yTcGv9Tp8_1),.dout(w_dff_B_SShyMNgN8_1),.clk(gclk));
	jdff dff_B_yKFOmL6P5_1(.din(w_dff_B_SShyMNgN8_1),.dout(w_dff_B_yKFOmL6P5_1),.clk(gclk));
	jdff dff_B_RkEsnCnM8_1(.din(w_dff_B_yKFOmL6P5_1),.dout(w_dff_B_RkEsnCnM8_1),.clk(gclk));
	jdff dff_B_m9lvf0eN6_1(.din(w_dff_B_RkEsnCnM8_1),.dout(w_dff_B_m9lvf0eN6_1),.clk(gclk));
	jdff dff_B_qc9FyenM2_1(.din(w_dff_B_m9lvf0eN6_1),.dout(w_dff_B_qc9FyenM2_1),.clk(gclk));
	jdff dff_B_LNX9EyJ24_1(.din(w_dff_B_qc9FyenM2_1),.dout(w_dff_B_LNX9EyJ24_1),.clk(gclk));
	jdff dff_B_wyWpdCvO3_1(.din(w_dff_B_LNX9EyJ24_1),.dout(w_dff_B_wyWpdCvO3_1),.clk(gclk));
	jdff dff_B_jmD3nOY58_1(.din(w_dff_B_wyWpdCvO3_1),.dout(w_dff_B_jmD3nOY58_1),.clk(gclk));
	jdff dff_B_bi72tpfm5_1(.din(w_dff_B_jmD3nOY58_1),.dout(w_dff_B_bi72tpfm5_1),.clk(gclk));
	jdff dff_B_bVL4ArLi6_1(.din(w_dff_B_bi72tpfm5_1),.dout(w_dff_B_bVL4ArLi6_1),.clk(gclk));
	jdff dff_B_OLHl6SlF6_1(.din(w_dff_B_bVL4ArLi6_1),.dout(w_dff_B_OLHl6SlF6_1),.clk(gclk));
	jdff dff_B_cC1TbIde8_1(.din(w_dff_B_OLHl6SlF6_1),.dout(w_dff_B_cC1TbIde8_1),.clk(gclk));
	jdff dff_B_npTdC99a0_1(.din(w_dff_B_cC1TbIde8_1),.dout(w_dff_B_npTdC99a0_1),.clk(gclk));
	jdff dff_B_BCnOsJAV2_1(.din(w_dff_B_npTdC99a0_1),.dout(w_dff_B_BCnOsJAV2_1),.clk(gclk));
	jdff dff_B_B2GyJLRl2_1(.din(w_dff_B_BCnOsJAV2_1),.dout(w_dff_B_B2GyJLRl2_1),.clk(gclk));
	jdff dff_B_zTg9Asyt2_1(.din(w_dff_B_B2GyJLRl2_1),.dout(w_dff_B_zTg9Asyt2_1),.clk(gclk));
	jdff dff_B_6HxPxKS97_1(.din(w_dff_B_zTg9Asyt2_1),.dout(w_dff_B_6HxPxKS97_1),.clk(gclk));
	jdff dff_B_uGDXx6qa1_1(.din(w_dff_B_6HxPxKS97_1),.dout(w_dff_B_uGDXx6qa1_1),.clk(gclk));
	jdff dff_B_iCIplsYd1_0(.din(n751),.dout(w_dff_B_iCIplsYd1_0),.clk(gclk));
	jdff dff_B_R032ZZRg9_0(.din(w_dff_B_iCIplsYd1_0),.dout(w_dff_B_R032ZZRg9_0),.clk(gclk));
	jdff dff_B_lIV4UJEk4_0(.din(w_dff_B_R032ZZRg9_0),.dout(w_dff_B_lIV4UJEk4_0),.clk(gclk));
	jdff dff_B_xTqWbW790_0(.din(w_dff_B_lIV4UJEk4_0),.dout(w_dff_B_xTqWbW790_0),.clk(gclk));
	jdff dff_B_ixbL4vuu8_0(.din(w_dff_B_xTqWbW790_0),.dout(w_dff_B_ixbL4vuu8_0),.clk(gclk));
	jdff dff_B_s5uNid6B0_0(.din(w_dff_B_ixbL4vuu8_0),.dout(w_dff_B_s5uNid6B0_0),.clk(gclk));
	jdff dff_B_Gx1wuIWB0_0(.din(w_dff_B_s5uNid6B0_0),.dout(w_dff_B_Gx1wuIWB0_0),.clk(gclk));
	jdff dff_B_QLhEGMfl8_0(.din(w_dff_B_Gx1wuIWB0_0),.dout(w_dff_B_QLhEGMfl8_0),.clk(gclk));
	jdff dff_B_GyKup3Yz8_0(.din(w_dff_B_QLhEGMfl8_0),.dout(w_dff_B_GyKup3Yz8_0),.clk(gclk));
	jdff dff_B_pG0Tfhxu4_0(.din(w_dff_B_GyKup3Yz8_0),.dout(w_dff_B_pG0Tfhxu4_0),.clk(gclk));
	jdff dff_B_Y0MESBHd9_0(.din(w_dff_B_pG0Tfhxu4_0),.dout(w_dff_B_Y0MESBHd9_0),.clk(gclk));
	jdff dff_B_0GCi309a2_0(.din(w_dff_B_Y0MESBHd9_0),.dout(w_dff_B_0GCi309a2_0),.clk(gclk));
	jdff dff_B_qr15E9pm1_0(.din(w_dff_B_0GCi309a2_0),.dout(w_dff_B_qr15E9pm1_0),.clk(gclk));
	jdff dff_B_SviJMRe40_0(.din(w_dff_B_qr15E9pm1_0),.dout(w_dff_B_SviJMRe40_0),.clk(gclk));
	jdff dff_B_98L6txer0_0(.din(w_dff_B_SviJMRe40_0),.dout(w_dff_B_98L6txer0_0),.clk(gclk));
	jdff dff_B_pQ67VDW02_0(.din(w_dff_B_98L6txer0_0),.dout(w_dff_B_pQ67VDW02_0),.clk(gclk));
	jdff dff_B_Riw8sEhq4_0(.din(w_dff_B_pQ67VDW02_0),.dout(w_dff_B_Riw8sEhq4_0),.clk(gclk));
	jdff dff_B_8d5uUr404_0(.din(w_dff_B_Riw8sEhq4_0),.dout(w_dff_B_8d5uUr404_0),.clk(gclk));
	jdff dff_B_2BDAb8Ld1_0(.din(w_dff_B_8d5uUr404_0),.dout(w_dff_B_2BDAb8Ld1_0),.clk(gclk));
	jdff dff_B_gaPI7QpK9_0(.din(w_dff_B_2BDAb8Ld1_0),.dout(w_dff_B_gaPI7QpK9_0),.clk(gclk));
	jdff dff_B_bckyv8fy8_0(.din(w_dff_B_gaPI7QpK9_0),.dout(w_dff_B_bckyv8fy8_0),.clk(gclk));
	jdff dff_B_z2CUQsrk8_0(.din(w_dff_B_bckyv8fy8_0),.dout(w_dff_B_z2CUQsrk8_0),.clk(gclk));
	jdff dff_B_UFE4WZqR9_0(.din(w_dff_B_z2CUQsrk8_0),.dout(w_dff_B_UFE4WZqR9_0),.clk(gclk));
	jdff dff_B_kc1zoTdG8_0(.din(w_dff_B_UFE4WZqR9_0),.dout(w_dff_B_kc1zoTdG8_0),.clk(gclk));
	jdff dff_B_Umk802Ry1_0(.din(w_dff_B_kc1zoTdG8_0),.dout(w_dff_B_Umk802Ry1_0),.clk(gclk));
	jdff dff_B_zpBsNDiN3_0(.din(w_dff_B_Umk802Ry1_0),.dout(w_dff_B_zpBsNDiN3_0),.clk(gclk));
	jdff dff_B_0jKSU1ix0_0(.din(w_dff_B_zpBsNDiN3_0),.dout(w_dff_B_0jKSU1ix0_0),.clk(gclk));
	jdff dff_B_koYusXgY5_0(.din(w_dff_B_0jKSU1ix0_0),.dout(w_dff_B_koYusXgY5_0),.clk(gclk));
	jdff dff_B_BoSNCSfl0_0(.din(w_dff_B_koYusXgY5_0),.dout(w_dff_B_BoSNCSfl0_0),.clk(gclk));
	jdff dff_B_NxkGtQvq7_0(.din(w_dff_B_BoSNCSfl0_0),.dout(w_dff_B_NxkGtQvq7_0),.clk(gclk));
	jdff dff_B_6Q9rhIwi3_0(.din(w_dff_B_NxkGtQvq7_0),.dout(w_dff_B_6Q9rhIwi3_0),.clk(gclk));
	jdff dff_B_Md306bRj5_0(.din(w_dff_B_6Q9rhIwi3_0),.dout(w_dff_B_Md306bRj5_0),.clk(gclk));
	jdff dff_B_Qbf0zgD62_0(.din(w_dff_B_Md306bRj5_0),.dout(w_dff_B_Qbf0zgD62_0),.clk(gclk));
	jdff dff_B_zvgZVG6U5_0(.din(w_dff_B_Qbf0zgD62_0),.dout(w_dff_B_zvgZVG6U5_0),.clk(gclk));
	jdff dff_B_7M3zvLsv9_0(.din(w_dff_B_zvgZVG6U5_0),.dout(w_dff_B_7M3zvLsv9_0),.clk(gclk));
	jdff dff_B_iGEiv4fl9_0(.din(w_dff_B_7M3zvLsv9_0),.dout(w_dff_B_iGEiv4fl9_0),.clk(gclk));
	jdff dff_B_bXOGno0P0_0(.din(w_dff_B_iGEiv4fl9_0),.dout(w_dff_B_bXOGno0P0_0),.clk(gclk));
	jdff dff_B_mE0JMGW64_0(.din(w_dff_B_bXOGno0P0_0),.dout(w_dff_B_mE0JMGW64_0),.clk(gclk));
	jdff dff_B_LpsdSPht5_0(.din(w_dff_B_mE0JMGW64_0),.dout(w_dff_B_LpsdSPht5_0),.clk(gclk));
	jdff dff_B_4PbJHVNJ1_0(.din(w_dff_B_LpsdSPht5_0),.dout(w_dff_B_4PbJHVNJ1_0),.clk(gclk));
	jdff dff_B_KBNebchZ7_0(.din(w_dff_B_4PbJHVNJ1_0),.dout(w_dff_B_KBNebchZ7_0),.clk(gclk));
	jdff dff_B_ymRIN3jK2_0(.din(w_dff_B_KBNebchZ7_0),.dout(w_dff_B_ymRIN3jK2_0),.clk(gclk));
	jdff dff_B_nsGtLrzT6_0(.din(w_dff_B_ymRIN3jK2_0),.dout(w_dff_B_nsGtLrzT6_0),.clk(gclk));
	jdff dff_B_eXgiMATL4_0(.din(w_dff_B_nsGtLrzT6_0),.dout(w_dff_B_eXgiMATL4_0),.clk(gclk));
	jdff dff_B_eDqZ8lPw9_0(.din(w_dff_B_eXgiMATL4_0),.dout(w_dff_B_eDqZ8lPw9_0),.clk(gclk));
	jdff dff_B_otWcS33k2_0(.din(w_dff_B_eDqZ8lPw9_0),.dout(w_dff_B_otWcS33k2_0),.clk(gclk));
	jdff dff_B_5NocYk2f2_0(.din(w_dff_B_otWcS33k2_0),.dout(w_dff_B_5NocYk2f2_0),.clk(gclk));
	jdff dff_B_BHGDl4sJ3_0(.din(w_dff_B_5NocYk2f2_0),.dout(w_dff_B_BHGDl4sJ3_0),.clk(gclk));
	jdff dff_B_0ot5iYN30_0(.din(w_dff_B_BHGDl4sJ3_0),.dout(w_dff_B_0ot5iYN30_0),.clk(gclk));
	jdff dff_B_aB7eZaWZ9_0(.din(w_dff_B_0ot5iYN30_0),.dout(w_dff_B_aB7eZaWZ9_0),.clk(gclk));
	jdff dff_B_8uCdyeHM3_0(.din(w_dff_B_aB7eZaWZ9_0),.dout(w_dff_B_8uCdyeHM3_0),.clk(gclk));
	jdff dff_B_yg1H9zqC3_0(.din(w_dff_B_8uCdyeHM3_0),.dout(w_dff_B_yg1H9zqC3_0),.clk(gclk));
	jdff dff_B_jUvToiwx6_0(.din(w_dff_B_yg1H9zqC3_0),.dout(w_dff_B_jUvToiwx6_0),.clk(gclk));
	jdff dff_B_JAIq4SKV0_0(.din(w_dff_B_jUvToiwx6_0),.dout(w_dff_B_JAIq4SKV0_0),.clk(gclk));
	jdff dff_B_CIQ32VdY8_0(.din(w_dff_B_JAIq4SKV0_0),.dout(w_dff_B_CIQ32VdY8_0),.clk(gclk));
	jdff dff_B_JYr9aXgA9_0(.din(w_dff_B_CIQ32VdY8_0),.dout(w_dff_B_JYr9aXgA9_0),.clk(gclk));
	jdff dff_B_PWDjvkGs6_0(.din(w_dff_B_JYr9aXgA9_0),.dout(w_dff_B_PWDjvkGs6_0),.clk(gclk));
	jdff dff_B_POJGLbQe0_0(.din(w_dff_B_PWDjvkGs6_0),.dout(w_dff_B_POJGLbQe0_0),.clk(gclk));
	jdff dff_B_VobqMd4O4_0(.din(w_dff_B_POJGLbQe0_0),.dout(w_dff_B_VobqMd4O4_0),.clk(gclk));
	jdff dff_B_SLEJI2E67_0(.din(w_dff_B_VobqMd4O4_0),.dout(w_dff_B_SLEJI2E67_0),.clk(gclk));
	jdff dff_B_nUECFkPE3_0(.din(w_dff_B_SLEJI2E67_0),.dout(w_dff_B_nUECFkPE3_0),.clk(gclk));
	jdff dff_B_4r2a8qYn0_1(.din(n744),.dout(w_dff_B_4r2a8qYn0_1),.clk(gclk));
	jdff dff_B_Sly2Rx7X7_1(.din(w_dff_B_4r2a8qYn0_1),.dout(w_dff_B_Sly2Rx7X7_1),.clk(gclk));
	jdff dff_B_hlydHVMl8_1(.din(w_dff_B_Sly2Rx7X7_1),.dout(w_dff_B_hlydHVMl8_1),.clk(gclk));
	jdff dff_B_yzeIPWWA1_1(.din(w_dff_B_hlydHVMl8_1),.dout(w_dff_B_yzeIPWWA1_1),.clk(gclk));
	jdff dff_B_wPodME3e2_1(.din(w_dff_B_yzeIPWWA1_1),.dout(w_dff_B_wPodME3e2_1),.clk(gclk));
	jdff dff_B_7GjLbvzm7_1(.din(w_dff_B_wPodME3e2_1),.dout(w_dff_B_7GjLbvzm7_1),.clk(gclk));
	jdff dff_B_juRmGHoY0_1(.din(w_dff_B_7GjLbvzm7_1),.dout(w_dff_B_juRmGHoY0_1),.clk(gclk));
	jdff dff_B_nDTvbOWK6_1(.din(w_dff_B_juRmGHoY0_1),.dout(w_dff_B_nDTvbOWK6_1),.clk(gclk));
	jdff dff_B_p0CKGQ2U5_1(.din(w_dff_B_nDTvbOWK6_1),.dout(w_dff_B_p0CKGQ2U5_1),.clk(gclk));
	jdff dff_B_lvVXzTXP7_1(.din(w_dff_B_p0CKGQ2U5_1),.dout(w_dff_B_lvVXzTXP7_1),.clk(gclk));
	jdff dff_B_ojAQA5Aw1_1(.din(w_dff_B_lvVXzTXP7_1),.dout(w_dff_B_ojAQA5Aw1_1),.clk(gclk));
	jdff dff_B_gDSCbj817_1(.din(w_dff_B_ojAQA5Aw1_1),.dout(w_dff_B_gDSCbj817_1),.clk(gclk));
	jdff dff_B_mbs9phc69_1(.din(w_dff_B_gDSCbj817_1),.dout(w_dff_B_mbs9phc69_1),.clk(gclk));
	jdff dff_B_I94G633r6_1(.din(w_dff_B_mbs9phc69_1),.dout(w_dff_B_I94G633r6_1),.clk(gclk));
	jdff dff_B_dnST0awd2_1(.din(w_dff_B_I94G633r6_1),.dout(w_dff_B_dnST0awd2_1),.clk(gclk));
	jdff dff_B_IZg8B82I0_1(.din(w_dff_B_dnST0awd2_1),.dout(w_dff_B_IZg8B82I0_1),.clk(gclk));
	jdff dff_B_gtrt0q9Z4_1(.din(w_dff_B_IZg8B82I0_1),.dout(w_dff_B_gtrt0q9Z4_1),.clk(gclk));
	jdff dff_B_jKTcvnDw0_1(.din(w_dff_B_gtrt0q9Z4_1),.dout(w_dff_B_jKTcvnDw0_1),.clk(gclk));
	jdff dff_B_HT2QJnO22_1(.din(w_dff_B_jKTcvnDw0_1),.dout(w_dff_B_HT2QJnO22_1),.clk(gclk));
	jdff dff_B_Ewicx5MI8_1(.din(w_dff_B_HT2QJnO22_1),.dout(w_dff_B_Ewicx5MI8_1),.clk(gclk));
	jdff dff_B_7Uusi3WG0_1(.din(w_dff_B_Ewicx5MI8_1),.dout(w_dff_B_7Uusi3WG0_1),.clk(gclk));
	jdff dff_B_Pj6balu61_1(.din(w_dff_B_7Uusi3WG0_1),.dout(w_dff_B_Pj6balu61_1),.clk(gclk));
	jdff dff_B_Su5dXGqT0_1(.din(w_dff_B_Pj6balu61_1),.dout(w_dff_B_Su5dXGqT0_1),.clk(gclk));
	jdff dff_B_1CGdUx5Y7_1(.din(w_dff_B_Su5dXGqT0_1),.dout(w_dff_B_1CGdUx5Y7_1),.clk(gclk));
	jdff dff_B_tDR81CLx2_1(.din(w_dff_B_1CGdUx5Y7_1),.dout(w_dff_B_tDR81CLx2_1),.clk(gclk));
	jdff dff_B_bs1PMIkH7_1(.din(w_dff_B_tDR81CLx2_1),.dout(w_dff_B_bs1PMIkH7_1),.clk(gclk));
	jdff dff_B_Y7OhseaZ9_1(.din(w_dff_B_bs1PMIkH7_1),.dout(w_dff_B_Y7OhseaZ9_1),.clk(gclk));
	jdff dff_B_BOeVL6ve7_1(.din(w_dff_B_Y7OhseaZ9_1),.dout(w_dff_B_BOeVL6ve7_1),.clk(gclk));
	jdff dff_B_g0tsrqBD1_1(.din(w_dff_B_BOeVL6ve7_1),.dout(w_dff_B_g0tsrqBD1_1),.clk(gclk));
	jdff dff_B_h5QnmR809_1(.din(w_dff_B_g0tsrqBD1_1),.dout(w_dff_B_h5QnmR809_1),.clk(gclk));
	jdff dff_B_xRkDJq5h9_1(.din(w_dff_B_h5QnmR809_1),.dout(w_dff_B_xRkDJq5h9_1),.clk(gclk));
	jdff dff_B_WWKSD8Cq4_1(.din(w_dff_B_xRkDJq5h9_1),.dout(w_dff_B_WWKSD8Cq4_1),.clk(gclk));
	jdff dff_B_Ig8YdTV84_1(.din(w_dff_B_WWKSD8Cq4_1),.dout(w_dff_B_Ig8YdTV84_1),.clk(gclk));
	jdff dff_B_pXHdOA077_1(.din(w_dff_B_Ig8YdTV84_1),.dout(w_dff_B_pXHdOA077_1),.clk(gclk));
	jdff dff_B_t2l5o3Ta6_1(.din(w_dff_B_pXHdOA077_1),.dout(w_dff_B_t2l5o3Ta6_1),.clk(gclk));
	jdff dff_B_boxmnPnb1_1(.din(w_dff_B_t2l5o3Ta6_1),.dout(w_dff_B_boxmnPnb1_1),.clk(gclk));
	jdff dff_B_HoysxmWq2_1(.din(w_dff_B_boxmnPnb1_1),.dout(w_dff_B_HoysxmWq2_1),.clk(gclk));
	jdff dff_B_cEPoh1h64_1(.din(w_dff_B_HoysxmWq2_1),.dout(w_dff_B_cEPoh1h64_1),.clk(gclk));
	jdff dff_B_u9DOPFVB9_1(.din(w_dff_B_cEPoh1h64_1),.dout(w_dff_B_u9DOPFVB9_1),.clk(gclk));
	jdff dff_B_JmMp7Cdw4_1(.din(w_dff_B_u9DOPFVB9_1),.dout(w_dff_B_JmMp7Cdw4_1),.clk(gclk));
	jdff dff_B_JQVCBCXc7_1(.din(w_dff_B_JmMp7Cdw4_1),.dout(w_dff_B_JQVCBCXc7_1),.clk(gclk));
	jdff dff_B_pZzBcMIm0_1(.din(w_dff_B_JQVCBCXc7_1),.dout(w_dff_B_pZzBcMIm0_1),.clk(gclk));
	jdff dff_B_l9WmSUtg4_1(.din(w_dff_B_pZzBcMIm0_1),.dout(w_dff_B_l9WmSUtg4_1),.clk(gclk));
	jdff dff_B_WgfPajVu1_1(.din(w_dff_B_l9WmSUtg4_1),.dout(w_dff_B_WgfPajVu1_1),.clk(gclk));
	jdff dff_B_mzaSY1Zu9_1(.din(w_dff_B_WgfPajVu1_1),.dout(w_dff_B_mzaSY1Zu9_1),.clk(gclk));
	jdff dff_B_OfoRcyLI7_1(.din(w_dff_B_mzaSY1Zu9_1),.dout(w_dff_B_OfoRcyLI7_1),.clk(gclk));
	jdff dff_B_9ZXlClCf9_1(.din(w_dff_B_OfoRcyLI7_1),.dout(w_dff_B_9ZXlClCf9_1),.clk(gclk));
	jdff dff_B_M4UGntXx5_1(.din(w_dff_B_9ZXlClCf9_1),.dout(w_dff_B_M4UGntXx5_1),.clk(gclk));
	jdff dff_B_LDXOTzf36_1(.din(w_dff_B_M4UGntXx5_1),.dout(w_dff_B_LDXOTzf36_1),.clk(gclk));
	jdff dff_B_yIbndY3H6_1(.din(w_dff_B_LDXOTzf36_1),.dout(w_dff_B_yIbndY3H6_1),.clk(gclk));
	jdff dff_B_A9D3q4lP5_1(.din(w_dff_B_yIbndY3H6_1),.dout(w_dff_B_A9D3q4lP5_1),.clk(gclk));
	jdff dff_B_n5TTfjRT9_1(.din(w_dff_B_A9D3q4lP5_1),.dout(w_dff_B_n5TTfjRT9_1),.clk(gclk));
	jdff dff_B_LzQpxSza9_1(.din(w_dff_B_n5TTfjRT9_1),.dout(w_dff_B_LzQpxSza9_1),.clk(gclk));
	jdff dff_B_NN0hhJfy2_1(.din(w_dff_B_LzQpxSza9_1),.dout(w_dff_B_NN0hhJfy2_1),.clk(gclk));
	jdff dff_B_AZxMxgX31_1(.din(w_dff_B_NN0hhJfy2_1),.dout(w_dff_B_AZxMxgX31_1),.clk(gclk));
	jdff dff_B_f9dMONXb3_1(.din(w_dff_B_AZxMxgX31_1),.dout(w_dff_B_f9dMONXb3_1),.clk(gclk));
	jdff dff_B_0HXGUKem9_1(.din(w_dff_B_f9dMONXb3_1),.dout(w_dff_B_0HXGUKem9_1),.clk(gclk));
	jdff dff_B_IBvWu3Eh6_1(.din(w_dff_B_0HXGUKem9_1),.dout(w_dff_B_IBvWu3Eh6_1),.clk(gclk));
	jdff dff_B_ma7LURTy0_1(.din(w_dff_B_IBvWu3Eh6_1),.dout(w_dff_B_ma7LURTy0_1),.clk(gclk));
	jdff dff_B_gZ9xFATs7_1(.din(w_dff_B_ma7LURTy0_1),.dout(w_dff_B_gZ9xFATs7_1),.clk(gclk));
	jdff dff_B_bK7ToB561_0(.din(n745),.dout(w_dff_B_bK7ToB561_0),.clk(gclk));
	jdff dff_B_vrl6EvLN9_0(.din(w_dff_B_bK7ToB561_0),.dout(w_dff_B_vrl6EvLN9_0),.clk(gclk));
	jdff dff_B_iyGeSKHv5_0(.din(w_dff_B_vrl6EvLN9_0),.dout(w_dff_B_iyGeSKHv5_0),.clk(gclk));
	jdff dff_B_wKyKD5oY3_0(.din(w_dff_B_iyGeSKHv5_0),.dout(w_dff_B_wKyKD5oY3_0),.clk(gclk));
	jdff dff_B_xh3lNg544_0(.din(w_dff_B_wKyKD5oY3_0),.dout(w_dff_B_xh3lNg544_0),.clk(gclk));
	jdff dff_B_33RCGcIN7_0(.din(w_dff_B_xh3lNg544_0),.dout(w_dff_B_33RCGcIN7_0),.clk(gclk));
	jdff dff_B_yAEvh6ME1_0(.din(w_dff_B_33RCGcIN7_0),.dout(w_dff_B_yAEvh6ME1_0),.clk(gclk));
	jdff dff_B_TqNbQJRH0_0(.din(w_dff_B_yAEvh6ME1_0),.dout(w_dff_B_TqNbQJRH0_0),.clk(gclk));
	jdff dff_B_C7RB8ZTe4_0(.din(w_dff_B_TqNbQJRH0_0),.dout(w_dff_B_C7RB8ZTe4_0),.clk(gclk));
	jdff dff_B_etSwmNbZ3_0(.din(w_dff_B_C7RB8ZTe4_0),.dout(w_dff_B_etSwmNbZ3_0),.clk(gclk));
	jdff dff_B_uZAVrlBY3_0(.din(w_dff_B_etSwmNbZ3_0),.dout(w_dff_B_uZAVrlBY3_0),.clk(gclk));
	jdff dff_B_xe8Wi7jE8_0(.din(w_dff_B_uZAVrlBY3_0),.dout(w_dff_B_xe8Wi7jE8_0),.clk(gclk));
	jdff dff_B_VOWqZwoz5_0(.din(w_dff_B_xe8Wi7jE8_0),.dout(w_dff_B_VOWqZwoz5_0),.clk(gclk));
	jdff dff_B_zESnTcPO2_0(.din(w_dff_B_VOWqZwoz5_0),.dout(w_dff_B_zESnTcPO2_0),.clk(gclk));
	jdff dff_B_OxueMZJc8_0(.din(w_dff_B_zESnTcPO2_0),.dout(w_dff_B_OxueMZJc8_0),.clk(gclk));
	jdff dff_B_pGG8WJUa9_0(.din(w_dff_B_OxueMZJc8_0),.dout(w_dff_B_pGG8WJUa9_0),.clk(gclk));
	jdff dff_B_Oq0fkz0l7_0(.din(w_dff_B_pGG8WJUa9_0),.dout(w_dff_B_Oq0fkz0l7_0),.clk(gclk));
	jdff dff_B_3RUhCgWm2_0(.din(w_dff_B_Oq0fkz0l7_0),.dout(w_dff_B_3RUhCgWm2_0),.clk(gclk));
	jdff dff_B_iKVZ2m0e4_0(.din(w_dff_B_3RUhCgWm2_0),.dout(w_dff_B_iKVZ2m0e4_0),.clk(gclk));
	jdff dff_B_HzNFQLS72_0(.din(w_dff_B_iKVZ2m0e4_0),.dout(w_dff_B_HzNFQLS72_0),.clk(gclk));
	jdff dff_B_6I4EmERV8_0(.din(w_dff_B_HzNFQLS72_0),.dout(w_dff_B_6I4EmERV8_0),.clk(gclk));
	jdff dff_B_EYevRhXP5_0(.din(w_dff_B_6I4EmERV8_0),.dout(w_dff_B_EYevRhXP5_0),.clk(gclk));
	jdff dff_B_CUAjfqae4_0(.din(w_dff_B_EYevRhXP5_0),.dout(w_dff_B_CUAjfqae4_0),.clk(gclk));
	jdff dff_B_OY5QezOA2_0(.din(w_dff_B_CUAjfqae4_0),.dout(w_dff_B_OY5QezOA2_0),.clk(gclk));
	jdff dff_B_xrVkakDe4_0(.din(w_dff_B_OY5QezOA2_0),.dout(w_dff_B_xrVkakDe4_0),.clk(gclk));
	jdff dff_B_o9dmVp507_0(.din(w_dff_B_xrVkakDe4_0),.dout(w_dff_B_o9dmVp507_0),.clk(gclk));
	jdff dff_B_bwGMiDeP9_0(.din(w_dff_B_o9dmVp507_0),.dout(w_dff_B_bwGMiDeP9_0),.clk(gclk));
	jdff dff_B_jvm9tsOV5_0(.din(w_dff_B_bwGMiDeP9_0),.dout(w_dff_B_jvm9tsOV5_0),.clk(gclk));
	jdff dff_B_AVi0ttD09_0(.din(w_dff_B_jvm9tsOV5_0),.dout(w_dff_B_AVi0ttD09_0),.clk(gclk));
	jdff dff_B_xTLU9toU0_0(.din(w_dff_B_AVi0ttD09_0),.dout(w_dff_B_xTLU9toU0_0),.clk(gclk));
	jdff dff_B_BUuWtqCV3_0(.din(w_dff_B_xTLU9toU0_0),.dout(w_dff_B_BUuWtqCV3_0),.clk(gclk));
	jdff dff_B_VO0v5epf5_0(.din(w_dff_B_BUuWtqCV3_0),.dout(w_dff_B_VO0v5epf5_0),.clk(gclk));
	jdff dff_B_oOuD9jeo5_0(.din(w_dff_B_VO0v5epf5_0),.dout(w_dff_B_oOuD9jeo5_0),.clk(gclk));
	jdff dff_B_EXleF4Sd9_0(.din(w_dff_B_oOuD9jeo5_0),.dout(w_dff_B_EXleF4Sd9_0),.clk(gclk));
	jdff dff_B_kKqLcXHM0_0(.din(w_dff_B_EXleF4Sd9_0),.dout(w_dff_B_kKqLcXHM0_0),.clk(gclk));
	jdff dff_B_zbY4bD9a6_0(.din(w_dff_B_kKqLcXHM0_0),.dout(w_dff_B_zbY4bD9a6_0),.clk(gclk));
	jdff dff_B_zQyWVxrd6_0(.din(w_dff_B_zbY4bD9a6_0),.dout(w_dff_B_zQyWVxrd6_0),.clk(gclk));
	jdff dff_B_nmKAHa1f6_0(.din(w_dff_B_zQyWVxrd6_0),.dout(w_dff_B_nmKAHa1f6_0),.clk(gclk));
	jdff dff_B_3aWDFIBf9_0(.din(w_dff_B_nmKAHa1f6_0),.dout(w_dff_B_3aWDFIBf9_0),.clk(gclk));
	jdff dff_B_IEBmjdSg9_0(.din(w_dff_B_3aWDFIBf9_0),.dout(w_dff_B_IEBmjdSg9_0),.clk(gclk));
	jdff dff_B_Bjty1Tt67_0(.din(w_dff_B_IEBmjdSg9_0),.dout(w_dff_B_Bjty1Tt67_0),.clk(gclk));
	jdff dff_B_53aklnda2_0(.din(w_dff_B_Bjty1Tt67_0),.dout(w_dff_B_53aklnda2_0),.clk(gclk));
	jdff dff_B_Bu79q6876_0(.din(w_dff_B_53aklnda2_0),.dout(w_dff_B_Bu79q6876_0),.clk(gclk));
	jdff dff_B_1yWYUlkS8_0(.din(w_dff_B_Bu79q6876_0),.dout(w_dff_B_1yWYUlkS8_0),.clk(gclk));
	jdff dff_B_0XKY71Rh7_0(.din(w_dff_B_1yWYUlkS8_0),.dout(w_dff_B_0XKY71Rh7_0),.clk(gclk));
	jdff dff_B_0XRA4b5v2_0(.din(w_dff_B_0XKY71Rh7_0),.dout(w_dff_B_0XRA4b5v2_0),.clk(gclk));
	jdff dff_B_rpPTQowr0_0(.din(w_dff_B_0XRA4b5v2_0),.dout(w_dff_B_rpPTQowr0_0),.clk(gclk));
	jdff dff_B_5TswgD3O8_0(.din(w_dff_B_rpPTQowr0_0),.dout(w_dff_B_5TswgD3O8_0),.clk(gclk));
	jdff dff_B_ckk5nHEA2_0(.din(w_dff_B_5TswgD3O8_0),.dout(w_dff_B_ckk5nHEA2_0),.clk(gclk));
	jdff dff_B_lQqTLJ0Q0_0(.din(w_dff_B_ckk5nHEA2_0),.dout(w_dff_B_lQqTLJ0Q0_0),.clk(gclk));
	jdff dff_B_yXlWp8g34_0(.din(w_dff_B_lQqTLJ0Q0_0),.dout(w_dff_B_yXlWp8g34_0),.clk(gclk));
	jdff dff_B_4J8UpfmA3_0(.din(w_dff_B_yXlWp8g34_0),.dout(w_dff_B_4J8UpfmA3_0),.clk(gclk));
	jdff dff_B_xnoGFQho2_0(.din(w_dff_B_4J8UpfmA3_0),.dout(w_dff_B_xnoGFQho2_0),.clk(gclk));
	jdff dff_B_83aPIXcz7_0(.din(w_dff_B_xnoGFQho2_0),.dout(w_dff_B_83aPIXcz7_0),.clk(gclk));
	jdff dff_B_UAS5stHz9_0(.din(w_dff_B_83aPIXcz7_0),.dout(w_dff_B_UAS5stHz9_0),.clk(gclk));
	jdff dff_B_TP3oONU42_0(.din(w_dff_B_UAS5stHz9_0),.dout(w_dff_B_TP3oONU42_0),.clk(gclk));
	jdff dff_B_iPaydoqZ6_0(.din(w_dff_B_TP3oONU42_0),.dout(w_dff_B_iPaydoqZ6_0),.clk(gclk));
	jdff dff_B_Ryv6wlV94_0(.din(w_dff_B_iPaydoqZ6_0),.dout(w_dff_B_Ryv6wlV94_0),.clk(gclk));
	jdff dff_B_i64hvzJ48_0(.din(w_dff_B_Ryv6wlV94_0),.dout(w_dff_B_i64hvzJ48_0),.clk(gclk));
	jdff dff_B_LsprbBuG0_0(.din(w_dff_B_i64hvzJ48_0),.dout(w_dff_B_LsprbBuG0_0),.clk(gclk));
	jdff dff_B_1Cx2caxz2_1(.din(n738),.dout(w_dff_B_1Cx2caxz2_1),.clk(gclk));
	jdff dff_B_vbRcEPTh3_1(.din(w_dff_B_1Cx2caxz2_1),.dout(w_dff_B_vbRcEPTh3_1),.clk(gclk));
	jdff dff_B_LvCxr4V80_1(.din(w_dff_B_vbRcEPTh3_1),.dout(w_dff_B_LvCxr4V80_1),.clk(gclk));
	jdff dff_B_z3WnlphU0_1(.din(w_dff_B_LvCxr4V80_1),.dout(w_dff_B_z3WnlphU0_1),.clk(gclk));
	jdff dff_B_mn7LwfYp9_1(.din(w_dff_B_z3WnlphU0_1),.dout(w_dff_B_mn7LwfYp9_1),.clk(gclk));
	jdff dff_B_KzmADoTA4_1(.din(w_dff_B_mn7LwfYp9_1),.dout(w_dff_B_KzmADoTA4_1),.clk(gclk));
	jdff dff_B_QODcd1RD4_1(.din(w_dff_B_KzmADoTA4_1),.dout(w_dff_B_QODcd1RD4_1),.clk(gclk));
	jdff dff_B_5L3Io06b1_1(.din(w_dff_B_QODcd1RD4_1),.dout(w_dff_B_5L3Io06b1_1),.clk(gclk));
	jdff dff_B_K7cmhTgc0_1(.din(w_dff_B_5L3Io06b1_1),.dout(w_dff_B_K7cmhTgc0_1),.clk(gclk));
	jdff dff_B_IoDvpxl32_1(.din(w_dff_B_K7cmhTgc0_1),.dout(w_dff_B_IoDvpxl32_1),.clk(gclk));
	jdff dff_B_fv4E2Fld4_1(.din(w_dff_B_IoDvpxl32_1),.dout(w_dff_B_fv4E2Fld4_1),.clk(gclk));
	jdff dff_B_sjdERbEs4_1(.din(w_dff_B_fv4E2Fld4_1),.dout(w_dff_B_sjdERbEs4_1),.clk(gclk));
	jdff dff_B_zfoIswA72_1(.din(w_dff_B_sjdERbEs4_1),.dout(w_dff_B_zfoIswA72_1),.clk(gclk));
	jdff dff_B_5l7hGFXW0_1(.din(w_dff_B_zfoIswA72_1),.dout(w_dff_B_5l7hGFXW0_1),.clk(gclk));
	jdff dff_B_bRSljdGJ7_1(.din(w_dff_B_5l7hGFXW0_1),.dout(w_dff_B_bRSljdGJ7_1),.clk(gclk));
	jdff dff_B_ZgQK24zP8_1(.din(w_dff_B_bRSljdGJ7_1),.dout(w_dff_B_ZgQK24zP8_1),.clk(gclk));
	jdff dff_B_naXpGiBI6_1(.din(w_dff_B_ZgQK24zP8_1),.dout(w_dff_B_naXpGiBI6_1),.clk(gclk));
	jdff dff_B_JMiN8GXZ6_1(.din(w_dff_B_naXpGiBI6_1),.dout(w_dff_B_JMiN8GXZ6_1),.clk(gclk));
	jdff dff_B_HUg9T4C80_1(.din(w_dff_B_JMiN8GXZ6_1),.dout(w_dff_B_HUg9T4C80_1),.clk(gclk));
	jdff dff_B_eq6ugiHg7_1(.din(w_dff_B_HUg9T4C80_1),.dout(w_dff_B_eq6ugiHg7_1),.clk(gclk));
	jdff dff_B_aPGmollr7_1(.din(w_dff_B_eq6ugiHg7_1),.dout(w_dff_B_aPGmollr7_1),.clk(gclk));
	jdff dff_B_mB9Nlvsz9_1(.din(w_dff_B_aPGmollr7_1),.dout(w_dff_B_mB9Nlvsz9_1),.clk(gclk));
	jdff dff_B_ViyzJoYs0_1(.din(w_dff_B_mB9Nlvsz9_1),.dout(w_dff_B_ViyzJoYs0_1),.clk(gclk));
	jdff dff_B_AtqpOaXn3_1(.din(w_dff_B_ViyzJoYs0_1),.dout(w_dff_B_AtqpOaXn3_1),.clk(gclk));
	jdff dff_B_FpYOZrTm9_1(.din(w_dff_B_AtqpOaXn3_1),.dout(w_dff_B_FpYOZrTm9_1),.clk(gclk));
	jdff dff_B_BHwGjug68_1(.din(w_dff_B_FpYOZrTm9_1),.dout(w_dff_B_BHwGjug68_1),.clk(gclk));
	jdff dff_B_DDfvJhH70_1(.din(w_dff_B_BHwGjug68_1),.dout(w_dff_B_DDfvJhH70_1),.clk(gclk));
	jdff dff_B_y389G3vK0_1(.din(w_dff_B_DDfvJhH70_1),.dout(w_dff_B_y389G3vK0_1),.clk(gclk));
	jdff dff_B_5FgpWpnl6_1(.din(w_dff_B_y389G3vK0_1),.dout(w_dff_B_5FgpWpnl6_1),.clk(gclk));
	jdff dff_B_U3JRfg9Z1_1(.din(w_dff_B_5FgpWpnl6_1),.dout(w_dff_B_U3JRfg9Z1_1),.clk(gclk));
	jdff dff_B_ClW58C9k4_1(.din(w_dff_B_U3JRfg9Z1_1),.dout(w_dff_B_ClW58C9k4_1),.clk(gclk));
	jdff dff_B_FK5tsFwb2_1(.din(w_dff_B_ClW58C9k4_1),.dout(w_dff_B_FK5tsFwb2_1),.clk(gclk));
	jdff dff_B_IYCZTfX03_1(.din(w_dff_B_FK5tsFwb2_1),.dout(w_dff_B_IYCZTfX03_1),.clk(gclk));
	jdff dff_B_PCAzmfHq9_1(.din(w_dff_B_IYCZTfX03_1),.dout(w_dff_B_PCAzmfHq9_1),.clk(gclk));
	jdff dff_B_wODzMxyA4_1(.din(w_dff_B_PCAzmfHq9_1),.dout(w_dff_B_wODzMxyA4_1),.clk(gclk));
	jdff dff_B_1gQkhwGp9_1(.din(w_dff_B_wODzMxyA4_1),.dout(w_dff_B_1gQkhwGp9_1),.clk(gclk));
	jdff dff_B_8Ue2Hj8O5_1(.din(w_dff_B_1gQkhwGp9_1),.dout(w_dff_B_8Ue2Hj8O5_1),.clk(gclk));
	jdff dff_B_90SkqCke5_1(.din(w_dff_B_8Ue2Hj8O5_1),.dout(w_dff_B_90SkqCke5_1),.clk(gclk));
	jdff dff_B_LaURsvA52_1(.din(w_dff_B_90SkqCke5_1),.dout(w_dff_B_LaURsvA52_1),.clk(gclk));
	jdff dff_B_K1nORJFn0_1(.din(w_dff_B_LaURsvA52_1),.dout(w_dff_B_K1nORJFn0_1),.clk(gclk));
	jdff dff_B_3LbkweKt7_1(.din(w_dff_B_K1nORJFn0_1),.dout(w_dff_B_3LbkweKt7_1),.clk(gclk));
	jdff dff_B_J0NPgAzB3_1(.din(w_dff_B_3LbkweKt7_1),.dout(w_dff_B_J0NPgAzB3_1),.clk(gclk));
	jdff dff_B_Datb44zb4_1(.din(w_dff_B_J0NPgAzB3_1),.dout(w_dff_B_Datb44zb4_1),.clk(gclk));
	jdff dff_B_0trhLKQ41_1(.din(w_dff_B_Datb44zb4_1),.dout(w_dff_B_0trhLKQ41_1),.clk(gclk));
	jdff dff_B_JhjYVBbm1_1(.din(w_dff_B_0trhLKQ41_1),.dout(w_dff_B_JhjYVBbm1_1),.clk(gclk));
	jdff dff_B_WU9ViVsG2_1(.din(w_dff_B_JhjYVBbm1_1),.dout(w_dff_B_WU9ViVsG2_1),.clk(gclk));
	jdff dff_B_sT70E6fh1_1(.din(w_dff_B_WU9ViVsG2_1),.dout(w_dff_B_sT70E6fh1_1),.clk(gclk));
	jdff dff_B_g8JdIeNz5_1(.din(w_dff_B_sT70E6fh1_1),.dout(w_dff_B_g8JdIeNz5_1),.clk(gclk));
	jdff dff_B_C8dI7RKM9_1(.din(w_dff_B_g8JdIeNz5_1),.dout(w_dff_B_C8dI7RKM9_1),.clk(gclk));
	jdff dff_B_dogrt0bY4_1(.din(w_dff_B_C8dI7RKM9_1),.dout(w_dff_B_dogrt0bY4_1),.clk(gclk));
	jdff dff_B_VAGySKC93_1(.din(w_dff_B_dogrt0bY4_1),.dout(w_dff_B_VAGySKC93_1),.clk(gclk));
	jdff dff_B_U7uE6QrZ9_1(.din(w_dff_B_VAGySKC93_1),.dout(w_dff_B_U7uE6QrZ9_1),.clk(gclk));
	jdff dff_B_9aBkHysO8_1(.din(w_dff_B_U7uE6QrZ9_1),.dout(w_dff_B_9aBkHysO8_1),.clk(gclk));
	jdff dff_B_DWyBmJIV0_1(.din(w_dff_B_9aBkHysO8_1),.dout(w_dff_B_DWyBmJIV0_1),.clk(gclk));
	jdff dff_B_ozCyyVsh4_1(.din(w_dff_B_DWyBmJIV0_1),.dout(w_dff_B_ozCyyVsh4_1),.clk(gclk));
	jdff dff_B_cI4GD7xH9_1(.din(w_dff_B_ozCyyVsh4_1),.dout(w_dff_B_cI4GD7xH9_1),.clk(gclk));
	jdff dff_B_0U4Zp4el5_1(.din(w_dff_B_cI4GD7xH9_1),.dout(w_dff_B_0U4Zp4el5_1),.clk(gclk));
	jdff dff_B_6BCzzzIk1_1(.din(w_dff_B_0U4Zp4el5_1),.dout(w_dff_B_6BCzzzIk1_1),.clk(gclk));
	jdff dff_B_NtYVoxbX5_1(.din(w_dff_B_6BCzzzIk1_1),.dout(w_dff_B_NtYVoxbX5_1),.clk(gclk));
	jdff dff_B_xMJ8Ciao7_0(.din(n739),.dout(w_dff_B_xMJ8Ciao7_0),.clk(gclk));
	jdff dff_B_vSFhHKni3_0(.din(w_dff_B_xMJ8Ciao7_0),.dout(w_dff_B_vSFhHKni3_0),.clk(gclk));
	jdff dff_B_w1imK7my9_0(.din(w_dff_B_vSFhHKni3_0),.dout(w_dff_B_w1imK7my9_0),.clk(gclk));
	jdff dff_B_pjCs8IJ28_0(.din(w_dff_B_w1imK7my9_0),.dout(w_dff_B_pjCs8IJ28_0),.clk(gclk));
	jdff dff_B_aNzkU1O32_0(.din(w_dff_B_pjCs8IJ28_0),.dout(w_dff_B_aNzkU1O32_0),.clk(gclk));
	jdff dff_B_vYZOsSVd9_0(.din(w_dff_B_aNzkU1O32_0),.dout(w_dff_B_vYZOsSVd9_0),.clk(gclk));
	jdff dff_B_DZYx8Q680_0(.din(w_dff_B_vYZOsSVd9_0),.dout(w_dff_B_DZYx8Q680_0),.clk(gclk));
	jdff dff_B_0oRIfecE9_0(.din(w_dff_B_DZYx8Q680_0),.dout(w_dff_B_0oRIfecE9_0),.clk(gclk));
	jdff dff_B_JzWFCzIV0_0(.din(w_dff_B_0oRIfecE9_0),.dout(w_dff_B_JzWFCzIV0_0),.clk(gclk));
	jdff dff_B_mltLMu050_0(.din(w_dff_B_JzWFCzIV0_0),.dout(w_dff_B_mltLMu050_0),.clk(gclk));
	jdff dff_B_ZjHoYKYX7_0(.din(w_dff_B_mltLMu050_0),.dout(w_dff_B_ZjHoYKYX7_0),.clk(gclk));
	jdff dff_B_7xxrVNAZ8_0(.din(w_dff_B_ZjHoYKYX7_0),.dout(w_dff_B_7xxrVNAZ8_0),.clk(gclk));
	jdff dff_B_f6YrUZjQ6_0(.din(w_dff_B_7xxrVNAZ8_0),.dout(w_dff_B_f6YrUZjQ6_0),.clk(gclk));
	jdff dff_B_zrv7936S3_0(.din(w_dff_B_f6YrUZjQ6_0),.dout(w_dff_B_zrv7936S3_0),.clk(gclk));
	jdff dff_B_GnqGi2xD8_0(.din(w_dff_B_zrv7936S3_0),.dout(w_dff_B_GnqGi2xD8_0),.clk(gclk));
	jdff dff_B_ubtHYmWE4_0(.din(w_dff_B_GnqGi2xD8_0),.dout(w_dff_B_ubtHYmWE4_0),.clk(gclk));
	jdff dff_B_AdTpG3142_0(.din(w_dff_B_ubtHYmWE4_0),.dout(w_dff_B_AdTpG3142_0),.clk(gclk));
	jdff dff_B_VNBffzMG2_0(.din(w_dff_B_AdTpG3142_0),.dout(w_dff_B_VNBffzMG2_0),.clk(gclk));
	jdff dff_B_NIWY21Si3_0(.din(w_dff_B_VNBffzMG2_0),.dout(w_dff_B_NIWY21Si3_0),.clk(gclk));
	jdff dff_B_tu8JMW301_0(.din(w_dff_B_NIWY21Si3_0),.dout(w_dff_B_tu8JMW301_0),.clk(gclk));
	jdff dff_B_qwIKNpJb1_0(.din(w_dff_B_tu8JMW301_0),.dout(w_dff_B_qwIKNpJb1_0),.clk(gclk));
	jdff dff_B_b68fVYw63_0(.din(w_dff_B_qwIKNpJb1_0),.dout(w_dff_B_b68fVYw63_0),.clk(gclk));
	jdff dff_B_MYI5QRP06_0(.din(w_dff_B_b68fVYw63_0),.dout(w_dff_B_MYI5QRP06_0),.clk(gclk));
	jdff dff_B_mpMpEfFL5_0(.din(w_dff_B_MYI5QRP06_0),.dout(w_dff_B_mpMpEfFL5_0),.clk(gclk));
	jdff dff_B_msFyOpjd9_0(.din(w_dff_B_mpMpEfFL5_0),.dout(w_dff_B_msFyOpjd9_0),.clk(gclk));
	jdff dff_B_kUPQ2jMn5_0(.din(w_dff_B_msFyOpjd9_0),.dout(w_dff_B_kUPQ2jMn5_0),.clk(gclk));
	jdff dff_B_bTjTUVwT6_0(.din(w_dff_B_kUPQ2jMn5_0),.dout(w_dff_B_bTjTUVwT6_0),.clk(gclk));
	jdff dff_B_WxdEABRo7_0(.din(w_dff_B_bTjTUVwT6_0),.dout(w_dff_B_WxdEABRo7_0),.clk(gclk));
	jdff dff_B_lGW2T8n41_0(.din(w_dff_B_WxdEABRo7_0),.dout(w_dff_B_lGW2T8n41_0),.clk(gclk));
	jdff dff_B_1X46zTKq0_0(.din(w_dff_B_lGW2T8n41_0),.dout(w_dff_B_1X46zTKq0_0),.clk(gclk));
	jdff dff_B_QwWCDhRA2_0(.din(w_dff_B_1X46zTKq0_0),.dout(w_dff_B_QwWCDhRA2_0),.clk(gclk));
	jdff dff_B_CdquVX552_0(.din(w_dff_B_QwWCDhRA2_0),.dout(w_dff_B_CdquVX552_0),.clk(gclk));
	jdff dff_B_wkifLEgs5_0(.din(w_dff_B_CdquVX552_0),.dout(w_dff_B_wkifLEgs5_0),.clk(gclk));
	jdff dff_B_J60MzZXP7_0(.din(w_dff_B_wkifLEgs5_0),.dout(w_dff_B_J60MzZXP7_0),.clk(gclk));
	jdff dff_B_GzHbQOhD1_0(.din(w_dff_B_J60MzZXP7_0),.dout(w_dff_B_GzHbQOhD1_0),.clk(gclk));
	jdff dff_B_tUntfrAW0_0(.din(w_dff_B_GzHbQOhD1_0),.dout(w_dff_B_tUntfrAW0_0),.clk(gclk));
	jdff dff_B_Ey4vlT174_0(.din(w_dff_B_tUntfrAW0_0),.dout(w_dff_B_Ey4vlT174_0),.clk(gclk));
	jdff dff_B_YxR7vpTH6_0(.din(w_dff_B_Ey4vlT174_0),.dout(w_dff_B_YxR7vpTH6_0),.clk(gclk));
	jdff dff_B_dpcinvtm0_0(.din(w_dff_B_YxR7vpTH6_0),.dout(w_dff_B_dpcinvtm0_0),.clk(gclk));
	jdff dff_B_K9nMNI3k6_0(.din(w_dff_B_dpcinvtm0_0),.dout(w_dff_B_K9nMNI3k6_0),.clk(gclk));
	jdff dff_B_6Pgs1x7T0_0(.din(w_dff_B_K9nMNI3k6_0),.dout(w_dff_B_6Pgs1x7T0_0),.clk(gclk));
	jdff dff_B_0b8BnNLT3_0(.din(w_dff_B_6Pgs1x7T0_0),.dout(w_dff_B_0b8BnNLT3_0),.clk(gclk));
	jdff dff_B_wqsYkcVq0_0(.din(w_dff_B_0b8BnNLT3_0),.dout(w_dff_B_wqsYkcVq0_0),.clk(gclk));
	jdff dff_B_SEL0GGUA1_0(.din(w_dff_B_wqsYkcVq0_0),.dout(w_dff_B_SEL0GGUA1_0),.clk(gclk));
	jdff dff_B_tjrxL4aE1_0(.din(w_dff_B_SEL0GGUA1_0),.dout(w_dff_B_tjrxL4aE1_0),.clk(gclk));
	jdff dff_B_UKmlommC3_0(.din(w_dff_B_tjrxL4aE1_0),.dout(w_dff_B_UKmlommC3_0),.clk(gclk));
	jdff dff_B_wVFqXuWr5_0(.din(w_dff_B_UKmlommC3_0),.dout(w_dff_B_wVFqXuWr5_0),.clk(gclk));
	jdff dff_B_UdpaqKrt7_0(.din(w_dff_B_wVFqXuWr5_0),.dout(w_dff_B_UdpaqKrt7_0),.clk(gclk));
	jdff dff_B_4gwA4mz83_0(.din(w_dff_B_UdpaqKrt7_0),.dout(w_dff_B_4gwA4mz83_0),.clk(gclk));
	jdff dff_B_vkPQatIp2_0(.din(w_dff_B_4gwA4mz83_0),.dout(w_dff_B_vkPQatIp2_0),.clk(gclk));
	jdff dff_B_LvLXhLf50_0(.din(w_dff_B_vkPQatIp2_0),.dout(w_dff_B_LvLXhLf50_0),.clk(gclk));
	jdff dff_B_9yAIr1Ce7_0(.din(w_dff_B_LvLXhLf50_0),.dout(w_dff_B_9yAIr1Ce7_0),.clk(gclk));
	jdff dff_B_iH32c2aR6_0(.din(w_dff_B_9yAIr1Ce7_0),.dout(w_dff_B_iH32c2aR6_0),.clk(gclk));
	jdff dff_B_8aJjRu5i1_0(.din(w_dff_B_iH32c2aR6_0),.dout(w_dff_B_8aJjRu5i1_0),.clk(gclk));
	jdff dff_B_FnTFnsir7_0(.din(w_dff_B_8aJjRu5i1_0),.dout(w_dff_B_FnTFnsir7_0),.clk(gclk));
	jdff dff_B_JKwARmW67_0(.din(w_dff_B_FnTFnsir7_0),.dout(w_dff_B_JKwARmW67_0),.clk(gclk));
	jdff dff_B_hxxUxdVp6_0(.din(w_dff_B_JKwARmW67_0),.dout(w_dff_B_hxxUxdVp6_0),.clk(gclk));
	jdff dff_B_LgOqTvTR3_0(.din(w_dff_B_hxxUxdVp6_0),.dout(w_dff_B_LgOqTvTR3_0),.clk(gclk));
	jdff dff_B_pQOVSYfd7_0(.din(w_dff_B_LgOqTvTR3_0),.dout(w_dff_B_pQOVSYfd7_0),.clk(gclk));
	jdff dff_B_QtN5qD899_1(.din(n732),.dout(w_dff_B_QtN5qD899_1),.clk(gclk));
	jdff dff_B_BhK3uIPd2_1(.din(w_dff_B_QtN5qD899_1),.dout(w_dff_B_BhK3uIPd2_1),.clk(gclk));
	jdff dff_B_nVyzy8dO1_1(.din(w_dff_B_BhK3uIPd2_1),.dout(w_dff_B_nVyzy8dO1_1),.clk(gclk));
	jdff dff_B_M2GbGVRc7_1(.din(w_dff_B_nVyzy8dO1_1),.dout(w_dff_B_M2GbGVRc7_1),.clk(gclk));
	jdff dff_B_rON9mXIN5_1(.din(w_dff_B_M2GbGVRc7_1),.dout(w_dff_B_rON9mXIN5_1),.clk(gclk));
	jdff dff_B_ZbMvnJ8n7_1(.din(w_dff_B_rON9mXIN5_1),.dout(w_dff_B_ZbMvnJ8n7_1),.clk(gclk));
	jdff dff_B_Ww93OQfn0_1(.din(w_dff_B_ZbMvnJ8n7_1),.dout(w_dff_B_Ww93OQfn0_1),.clk(gclk));
	jdff dff_B_Q8dcIBKq6_1(.din(w_dff_B_Ww93OQfn0_1),.dout(w_dff_B_Q8dcIBKq6_1),.clk(gclk));
	jdff dff_B_2tNelLJL8_1(.din(w_dff_B_Q8dcIBKq6_1),.dout(w_dff_B_2tNelLJL8_1),.clk(gclk));
	jdff dff_B_9oDwAZwX2_1(.din(w_dff_B_2tNelLJL8_1),.dout(w_dff_B_9oDwAZwX2_1),.clk(gclk));
	jdff dff_B_qytbBNr40_1(.din(w_dff_B_9oDwAZwX2_1),.dout(w_dff_B_qytbBNr40_1),.clk(gclk));
	jdff dff_B_DQzX6z0F2_1(.din(w_dff_B_qytbBNr40_1),.dout(w_dff_B_DQzX6z0F2_1),.clk(gclk));
	jdff dff_B_qsKPAzlQ3_1(.din(w_dff_B_DQzX6z0F2_1),.dout(w_dff_B_qsKPAzlQ3_1),.clk(gclk));
	jdff dff_B_XaqLyrZn8_1(.din(w_dff_B_qsKPAzlQ3_1),.dout(w_dff_B_XaqLyrZn8_1),.clk(gclk));
	jdff dff_B_gumfe9L20_1(.din(w_dff_B_XaqLyrZn8_1),.dout(w_dff_B_gumfe9L20_1),.clk(gclk));
	jdff dff_B_6pAGLQS84_1(.din(w_dff_B_gumfe9L20_1),.dout(w_dff_B_6pAGLQS84_1),.clk(gclk));
	jdff dff_B_jyyO2smQ6_1(.din(w_dff_B_6pAGLQS84_1),.dout(w_dff_B_jyyO2smQ6_1),.clk(gclk));
	jdff dff_B_QMgJQDr59_1(.din(w_dff_B_jyyO2smQ6_1),.dout(w_dff_B_QMgJQDr59_1),.clk(gclk));
	jdff dff_B_UkEvQpEm5_1(.din(w_dff_B_QMgJQDr59_1),.dout(w_dff_B_UkEvQpEm5_1),.clk(gclk));
	jdff dff_B_rxigErof6_1(.din(w_dff_B_UkEvQpEm5_1),.dout(w_dff_B_rxigErof6_1),.clk(gclk));
	jdff dff_B_xBO1dK357_1(.din(w_dff_B_rxigErof6_1),.dout(w_dff_B_xBO1dK357_1),.clk(gclk));
	jdff dff_B_rHaX9fF95_1(.din(w_dff_B_xBO1dK357_1),.dout(w_dff_B_rHaX9fF95_1),.clk(gclk));
	jdff dff_B_GAd2QaDS8_1(.din(w_dff_B_rHaX9fF95_1),.dout(w_dff_B_GAd2QaDS8_1),.clk(gclk));
	jdff dff_B_GclAZwzu5_1(.din(w_dff_B_GAd2QaDS8_1),.dout(w_dff_B_GclAZwzu5_1),.clk(gclk));
	jdff dff_B_7vnjpK433_1(.din(w_dff_B_GclAZwzu5_1),.dout(w_dff_B_7vnjpK433_1),.clk(gclk));
	jdff dff_B_qul3X06P7_1(.din(w_dff_B_7vnjpK433_1),.dout(w_dff_B_qul3X06P7_1),.clk(gclk));
	jdff dff_B_RwsYYg4w0_1(.din(w_dff_B_qul3X06P7_1),.dout(w_dff_B_RwsYYg4w0_1),.clk(gclk));
	jdff dff_B_PqEnw8Th4_1(.din(w_dff_B_RwsYYg4w0_1),.dout(w_dff_B_PqEnw8Th4_1),.clk(gclk));
	jdff dff_B_4hwD080H1_1(.din(w_dff_B_PqEnw8Th4_1),.dout(w_dff_B_4hwD080H1_1),.clk(gclk));
	jdff dff_B_GWk0qToj9_1(.din(w_dff_B_4hwD080H1_1),.dout(w_dff_B_GWk0qToj9_1),.clk(gclk));
	jdff dff_B_tV5ewyNb8_1(.din(w_dff_B_GWk0qToj9_1),.dout(w_dff_B_tV5ewyNb8_1),.clk(gclk));
	jdff dff_B_OFBrhHVk2_1(.din(w_dff_B_tV5ewyNb8_1),.dout(w_dff_B_OFBrhHVk2_1),.clk(gclk));
	jdff dff_B_ZPdKca7b7_1(.din(w_dff_B_OFBrhHVk2_1),.dout(w_dff_B_ZPdKca7b7_1),.clk(gclk));
	jdff dff_B_WMiaqdY48_1(.din(w_dff_B_ZPdKca7b7_1),.dout(w_dff_B_WMiaqdY48_1),.clk(gclk));
	jdff dff_B_50aNQJna7_1(.din(w_dff_B_WMiaqdY48_1),.dout(w_dff_B_50aNQJna7_1),.clk(gclk));
	jdff dff_B_YTBJ8uZ56_1(.din(w_dff_B_50aNQJna7_1),.dout(w_dff_B_YTBJ8uZ56_1),.clk(gclk));
	jdff dff_B_ZEWd1Usu6_1(.din(w_dff_B_YTBJ8uZ56_1),.dout(w_dff_B_ZEWd1Usu6_1),.clk(gclk));
	jdff dff_B_Ro5PxidI0_1(.din(w_dff_B_ZEWd1Usu6_1),.dout(w_dff_B_Ro5PxidI0_1),.clk(gclk));
	jdff dff_B_fxRK22Ws0_1(.din(w_dff_B_Ro5PxidI0_1),.dout(w_dff_B_fxRK22Ws0_1),.clk(gclk));
	jdff dff_B_ebgIrvys7_1(.din(w_dff_B_fxRK22Ws0_1),.dout(w_dff_B_ebgIrvys7_1),.clk(gclk));
	jdff dff_B_BCWSgJn99_1(.din(w_dff_B_ebgIrvys7_1),.dout(w_dff_B_BCWSgJn99_1),.clk(gclk));
	jdff dff_B_vv69iHma1_1(.din(w_dff_B_BCWSgJn99_1),.dout(w_dff_B_vv69iHma1_1),.clk(gclk));
	jdff dff_B_SpovpCDb4_1(.din(w_dff_B_vv69iHma1_1),.dout(w_dff_B_SpovpCDb4_1),.clk(gclk));
	jdff dff_B_01gwM5td1_1(.din(w_dff_B_SpovpCDb4_1),.dout(w_dff_B_01gwM5td1_1),.clk(gclk));
	jdff dff_B_3ydsrsbU9_1(.din(w_dff_B_01gwM5td1_1),.dout(w_dff_B_3ydsrsbU9_1),.clk(gclk));
	jdff dff_B_19EKRhkE9_1(.din(w_dff_B_3ydsrsbU9_1),.dout(w_dff_B_19EKRhkE9_1),.clk(gclk));
	jdff dff_B_GPuZbTUg8_1(.din(w_dff_B_19EKRhkE9_1),.dout(w_dff_B_GPuZbTUg8_1),.clk(gclk));
	jdff dff_B_KcXhrDlg6_1(.din(w_dff_B_GPuZbTUg8_1),.dout(w_dff_B_KcXhrDlg6_1),.clk(gclk));
	jdff dff_B_s7jEAdkM2_1(.din(w_dff_B_KcXhrDlg6_1),.dout(w_dff_B_s7jEAdkM2_1),.clk(gclk));
	jdff dff_B_m3mI4AfZ0_1(.din(w_dff_B_s7jEAdkM2_1),.dout(w_dff_B_m3mI4AfZ0_1),.clk(gclk));
	jdff dff_B_LhlkRvhW5_1(.din(w_dff_B_m3mI4AfZ0_1),.dout(w_dff_B_LhlkRvhW5_1),.clk(gclk));
	jdff dff_B_t3UiMecJ2_1(.din(w_dff_B_LhlkRvhW5_1),.dout(w_dff_B_t3UiMecJ2_1),.clk(gclk));
	jdff dff_B_c2MWpj7p1_1(.din(w_dff_B_t3UiMecJ2_1),.dout(w_dff_B_c2MWpj7p1_1),.clk(gclk));
	jdff dff_B_MmIq7VXG8_1(.din(w_dff_B_c2MWpj7p1_1),.dout(w_dff_B_MmIq7VXG8_1),.clk(gclk));
	jdff dff_B_92kAfPWp0_1(.din(w_dff_B_MmIq7VXG8_1),.dout(w_dff_B_92kAfPWp0_1),.clk(gclk));
	jdff dff_B_PMoP7dQt5_1(.din(w_dff_B_92kAfPWp0_1),.dout(w_dff_B_PMoP7dQt5_1),.clk(gclk));
	jdff dff_B_vdKdPBZQ8_1(.din(w_dff_B_PMoP7dQt5_1),.dout(w_dff_B_vdKdPBZQ8_1),.clk(gclk));
	jdff dff_B_WezfSukm9_1(.din(w_dff_B_vdKdPBZQ8_1),.dout(w_dff_B_WezfSukm9_1),.clk(gclk));
	jdff dff_B_3EbZKUZW6_0(.din(n733),.dout(w_dff_B_3EbZKUZW6_0),.clk(gclk));
	jdff dff_B_m5xhbG9y8_0(.din(w_dff_B_3EbZKUZW6_0),.dout(w_dff_B_m5xhbG9y8_0),.clk(gclk));
	jdff dff_B_xVRGVVqd6_0(.din(w_dff_B_m5xhbG9y8_0),.dout(w_dff_B_xVRGVVqd6_0),.clk(gclk));
	jdff dff_B_OLecySnw0_0(.din(w_dff_B_xVRGVVqd6_0),.dout(w_dff_B_OLecySnw0_0),.clk(gclk));
	jdff dff_B_RdAXibh13_0(.din(w_dff_B_OLecySnw0_0),.dout(w_dff_B_RdAXibh13_0),.clk(gclk));
	jdff dff_B_A5rMYJBz8_0(.din(w_dff_B_RdAXibh13_0),.dout(w_dff_B_A5rMYJBz8_0),.clk(gclk));
	jdff dff_B_qobfzLXL2_0(.din(w_dff_B_A5rMYJBz8_0),.dout(w_dff_B_qobfzLXL2_0),.clk(gclk));
	jdff dff_B_Nyf5Y3g61_0(.din(w_dff_B_qobfzLXL2_0),.dout(w_dff_B_Nyf5Y3g61_0),.clk(gclk));
	jdff dff_B_Hkf1kb616_0(.din(w_dff_B_Nyf5Y3g61_0),.dout(w_dff_B_Hkf1kb616_0),.clk(gclk));
	jdff dff_B_kF2fPO3l1_0(.din(w_dff_B_Hkf1kb616_0),.dout(w_dff_B_kF2fPO3l1_0),.clk(gclk));
	jdff dff_B_EvNMMVMc0_0(.din(w_dff_B_kF2fPO3l1_0),.dout(w_dff_B_EvNMMVMc0_0),.clk(gclk));
	jdff dff_B_EHP7Ju2R1_0(.din(w_dff_B_EvNMMVMc0_0),.dout(w_dff_B_EHP7Ju2R1_0),.clk(gclk));
	jdff dff_B_nov3DkHn6_0(.din(w_dff_B_EHP7Ju2R1_0),.dout(w_dff_B_nov3DkHn6_0),.clk(gclk));
	jdff dff_B_skjKwW3f6_0(.din(w_dff_B_nov3DkHn6_0),.dout(w_dff_B_skjKwW3f6_0),.clk(gclk));
	jdff dff_B_rcR9tqwC3_0(.din(w_dff_B_skjKwW3f6_0),.dout(w_dff_B_rcR9tqwC3_0),.clk(gclk));
	jdff dff_B_O1mV4QtD9_0(.din(w_dff_B_rcR9tqwC3_0),.dout(w_dff_B_O1mV4QtD9_0),.clk(gclk));
	jdff dff_B_mTyNPoAB0_0(.din(w_dff_B_O1mV4QtD9_0),.dout(w_dff_B_mTyNPoAB0_0),.clk(gclk));
	jdff dff_B_rv76iRzu1_0(.din(w_dff_B_mTyNPoAB0_0),.dout(w_dff_B_rv76iRzu1_0),.clk(gclk));
	jdff dff_B_9BhQMxDU9_0(.din(w_dff_B_rv76iRzu1_0),.dout(w_dff_B_9BhQMxDU9_0),.clk(gclk));
	jdff dff_B_E03CVzQb8_0(.din(w_dff_B_9BhQMxDU9_0),.dout(w_dff_B_E03CVzQb8_0),.clk(gclk));
	jdff dff_B_3YGaRqIu4_0(.din(w_dff_B_E03CVzQb8_0),.dout(w_dff_B_3YGaRqIu4_0),.clk(gclk));
	jdff dff_B_qOrN67cM1_0(.din(w_dff_B_3YGaRqIu4_0),.dout(w_dff_B_qOrN67cM1_0),.clk(gclk));
	jdff dff_B_ZlhKjNc12_0(.din(w_dff_B_qOrN67cM1_0),.dout(w_dff_B_ZlhKjNc12_0),.clk(gclk));
	jdff dff_B_dOn35z4Y0_0(.din(w_dff_B_ZlhKjNc12_0),.dout(w_dff_B_dOn35z4Y0_0),.clk(gclk));
	jdff dff_B_58atLflz6_0(.din(w_dff_B_dOn35z4Y0_0),.dout(w_dff_B_58atLflz6_0),.clk(gclk));
	jdff dff_B_njGhdoid9_0(.din(w_dff_B_58atLflz6_0),.dout(w_dff_B_njGhdoid9_0),.clk(gclk));
	jdff dff_B_58U6EFxH0_0(.din(w_dff_B_njGhdoid9_0),.dout(w_dff_B_58U6EFxH0_0),.clk(gclk));
	jdff dff_B_GKoaAw8s3_0(.din(w_dff_B_58U6EFxH0_0),.dout(w_dff_B_GKoaAw8s3_0),.clk(gclk));
	jdff dff_B_bAz2h1C45_0(.din(w_dff_B_GKoaAw8s3_0),.dout(w_dff_B_bAz2h1C45_0),.clk(gclk));
	jdff dff_B_UO4rzyae3_0(.din(w_dff_B_bAz2h1C45_0),.dout(w_dff_B_UO4rzyae3_0),.clk(gclk));
	jdff dff_B_095kRksM1_0(.din(w_dff_B_UO4rzyae3_0),.dout(w_dff_B_095kRksM1_0),.clk(gclk));
	jdff dff_B_lcov63Po0_0(.din(w_dff_B_095kRksM1_0),.dout(w_dff_B_lcov63Po0_0),.clk(gclk));
	jdff dff_B_V6tpfWNY7_0(.din(w_dff_B_lcov63Po0_0),.dout(w_dff_B_V6tpfWNY7_0),.clk(gclk));
	jdff dff_B_0pDBbWT35_0(.din(w_dff_B_V6tpfWNY7_0),.dout(w_dff_B_0pDBbWT35_0),.clk(gclk));
	jdff dff_B_Lm5xfr8P1_0(.din(w_dff_B_0pDBbWT35_0),.dout(w_dff_B_Lm5xfr8P1_0),.clk(gclk));
	jdff dff_B_W3tYjjy10_0(.din(w_dff_B_Lm5xfr8P1_0),.dout(w_dff_B_W3tYjjy10_0),.clk(gclk));
	jdff dff_B_6as0KEqd5_0(.din(w_dff_B_W3tYjjy10_0),.dout(w_dff_B_6as0KEqd5_0),.clk(gclk));
	jdff dff_B_6CVVIedW9_0(.din(w_dff_B_6as0KEqd5_0),.dout(w_dff_B_6CVVIedW9_0),.clk(gclk));
	jdff dff_B_cgymDpta2_0(.din(w_dff_B_6CVVIedW9_0),.dout(w_dff_B_cgymDpta2_0),.clk(gclk));
	jdff dff_B_OxTSltq28_0(.din(w_dff_B_cgymDpta2_0),.dout(w_dff_B_OxTSltq28_0),.clk(gclk));
	jdff dff_B_NYBhYppf2_0(.din(w_dff_B_OxTSltq28_0),.dout(w_dff_B_NYBhYppf2_0),.clk(gclk));
	jdff dff_B_oMx0QT8S6_0(.din(w_dff_B_NYBhYppf2_0),.dout(w_dff_B_oMx0QT8S6_0),.clk(gclk));
	jdff dff_B_84DNG2JZ9_0(.din(w_dff_B_oMx0QT8S6_0),.dout(w_dff_B_84DNG2JZ9_0),.clk(gclk));
	jdff dff_B_EWryNmyW9_0(.din(w_dff_B_84DNG2JZ9_0),.dout(w_dff_B_EWryNmyW9_0),.clk(gclk));
	jdff dff_B_arYWH0Ma9_0(.din(w_dff_B_EWryNmyW9_0),.dout(w_dff_B_arYWH0Ma9_0),.clk(gclk));
	jdff dff_B_ug4mcUrf6_0(.din(w_dff_B_arYWH0Ma9_0),.dout(w_dff_B_ug4mcUrf6_0),.clk(gclk));
	jdff dff_B_pPom2blk5_0(.din(w_dff_B_ug4mcUrf6_0),.dout(w_dff_B_pPom2blk5_0),.clk(gclk));
	jdff dff_B_8LByvSlY7_0(.din(w_dff_B_pPom2blk5_0),.dout(w_dff_B_8LByvSlY7_0),.clk(gclk));
	jdff dff_B_vxmWHeNr3_0(.din(w_dff_B_8LByvSlY7_0),.dout(w_dff_B_vxmWHeNr3_0),.clk(gclk));
	jdff dff_B_C0ENE8n84_0(.din(w_dff_B_vxmWHeNr3_0),.dout(w_dff_B_C0ENE8n84_0),.clk(gclk));
	jdff dff_B_HRkudgNT9_0(.din(w_dff_B_C0ENE8n84_0),.dout(w_dff_B_HRkudgNT9_0),.clk(gclk));
	jdff dff_B_Gcz3vLz62_0(.din(w_dff_B_HRkudgNT9_0),.dout(w_dff_B_Gcz3vLz62_0),.clk(gclk));
	jdff dff_B_EhHOQVgi4_0(.din(w_dff_B_Gcz3vLz62_0),.dout(w_dff_B_EhHOQVgi4_0),.clk(gclk));
	jdff dff_B_zJxe281o8_0(.din(w_dff_B_EhHOQVgi4_0),.dout(w_dff_B_zJxe281o8_0),.clk(gclk));
	jdff dff_B_vMQXSUN57_0(.din(w_dff_B_zJxe281o8_0),.dout(w_dff_B_vMQXSUN57_0),.clk(gclk));
	jdff dff_B_Z2LiN9iz2_0(.din(w_dff_B_vMQXSUN57_0),.dout(w_dff_B_Z2LiN9iz2_0),.clk(gclk));
	jdff dff_B_nQBMPS0x9_0(.din(w_dff_B_Z2LiN9iz2_0),.dout(w_dff_B_nQBMPS0x9_0),.clk(gclk));
	jdff dff_B_jX94jsrp1_0(.din(w_dff_B_nQBMPS0x9_0),.dout(w_dff_B_jX94jsrp1_0),.clk(gclk));
	jdff dff_B_2Fh0fFQ36_1(.din(n726),.dout(w_dff_B_2Fh0fFQ36_1),.clk(gclk));
	jdff dff_B_cna6aabl3_1(.din(w_dff_B_2Fh0fFQ36_1),.dout(w_dff_B_cna6aabl3_1),.clk(gclk));
	jdff dff_B_8pNKKJkC4_1(.din(w_dff_B_cna6aabl3_1),.dout(w_dff_B_8pNKKJkC4_1),.clk(gclk));
	jdff dff_B_IEwzXTD45_1(.din(w_dff_B_8pNKKJkC4_1),.dout(w_dff_B_IEwzXTD45_1),.clk(gclk));
	jdff dff_B_Lvyjbjhr6_1(.din(w_dff_B_IEwzXTD45_1),.dout(w_dff_B_Lvyjbjhr6_1),.clk(gclk));
	jdff dff_B_BvQqoA6l3_1(.din(w_dff_B_Lvyjbjhr6_1),.dout(w_dff_B_BvQqoA6l3_1),.clk(gclk));
	jdff dff_B_wqk3qosK7_1(.din(w_dff_B_BvQqoA6l3_1),.dout(w_dff_B_wqk3qosK7_1),.clk(gclk));
	jdff dff_B_4wpnnK5J2_1(.din(w_dff_B_wqk3qosK7_1),.dout(w_dff_B_4wpnnK5J2_1),.clk(gclk));
	jdff dff_B_3Jf4ZWm04_1(.din(w_dff_B_4wpnnK5J2_1),.dout(w_dff_B_3Jf4ZWm04_1),.clk(gclk));
	jdff dff_B_YwLuvEKI6_1(.din(w_dff_B_3Jf4ZWm04_1),.dout(w_dff_B_YwLuvEKI6_1),.clk(gclk));
	jdff dff_B_4YHJtBmE0_1(.din(w_dff_B_YwLuvEKI6_1),.dout(w_dff_B_4YHJtBmE0_1),.clk(gclk));
	jdff dff_B_Vr3CkPg10_1(.din(w_dff_B_4YHJtBmE0_1),.dout(w_dff_B_Vr3CkPg10_1),.clk(gclk));
	jdff dff_B_eUPKISmw4_1(.din(w_dff_B_Vr3CkPg10_1),.dout(w_dff_B_eUPKISmw4_1),.clk(gclk));
	jdff dff_B_jioS5rU41_1(.din(w_dff_B_eUPKISmw4_1),.dout(w_dff_B_jioS5rU41_1),.clk(gclk));
	jdff dff_B_k4Cw3Myd1_1(.din(w_dff_B_jioS5rU41_1),.dout(w_dff_B_k4Cw3Myd1_1),.clk(gclk));
	jdff dff_B_DZv0marw9_1(.din(w_dff_B_k4Cw3Myd1_1),.dout(w_dff_B_DZv0marw9_1),.clk(gclk));
	jdff dff_B_AdoR8d0i0_1(.din(w_dff_B_DZv0marw9_1),.dout(w_dff_B_AdoR8d0i0_1),.clk(gclk));
	jdff dff_B_zUmhhjUJ0_1(.din(w_dff_B_AdoR8d0i0_1),.dout(w_dff_B_zUmhhjUJ0_1),.clk(gclk));
	jdff dff_B_g0wot8bn0_1(.din(w_dff_B_zUmhhjUJ0_1),.dout(w_dff_B_g0wot8bn0_1),.clk(gclk));
	jdff dff_B_863NnPMp2_1(.din(w_dff_B_g0wot8bn0_1),.dout(w_dff_B_863NnPMp2_1),.clk(gclk));
	jdff dff_B_bwXv3Nma9_1(.din(w_dff_B_863NnPMp2_1),.dout(w_dff_B_bwXv3Nma9_1),.clk(gclk));
	jdff dff_B_POVRJj548_1(.din(w_dff_B_bwXv3Nma9_1),.dout(w_dff_B_POVRJj548_1),.clk(gclk));
	jdff dff_B_0V30eLpk9_1(.din(w_dff_B_POVRJj548_1),.dout(w_dff_B_0V30eLpk9_1),.clk(gclk));
	jdff dff_B_5gds8XUZ4_1(.din(w_dff_B_0V30eLpk9_1),.dout(w_dff_B_5gds8XUZ4_1),.clk(gclk));
	jdff dff_B_lPqfSb8b0_1(.din(w_dff_B_5gds8XUZ4_1),.dout(w_dff_B_lPqfSb8b0_1),.clk(gclk));
	jdff dff_B_fipJqsSe8_1(.din(w_dff_B_lPqfSb8b0_1),.dout(w_dff_B_fipJqsSe8_1),.clk(gclk));
	jdff dff_B_dLIrZH2K6_1(.din(w_dff_B_fipJqsSe8_1),.dout(w_dff_B_dLIrZH2K6_1),.clk(gclk));
	jdff dff_B_4Rz9h9rD4_1(.din(w_dff_B_dLIrZH2K6_1),.dout(w_dff_B_4Rz9h9rD4_1),.clk(gclk));
	jdff dff_B_S4w2GT5n6_1(.din(w_dff_B_4Rz9h9rD4_1),.dout(w_dff_B_S4w2GT5n6_1),.clk(gclk));
	jdff dff_B_eQ1qDrA86_1(.din(w_dff_B_S4w2GT5n6_1),.dout(w_dff_B_eQ1qDrA86_1),.clk(gclk));
	jdff dff_B_eiYeq4ox4_1(.din(w_dff_B_eQ1qDrA86_1),.dout(w_dff_B_eiYeq4ox4_1),.clk(gclk));
	jdff dff_B_ou0RgOdy9_1(.din(w_dff_B_eiYeq4ox4_1),.dout(w_dff_B_ou0RgOdy9_1),.clk(gclk));
	jdff dff_B_gDyc3p8b0_1(.din(w_dff_B_ou0RgOdy9_1),.dout(w_dff_B_gDyc3p8b0_1),.clk(gclk));
	jdff dff_B_Hb4m2qnY3_1(.din(w_dff_B_gDyc3p8b0_1),.dout(w_dff_B_Hb4m2qnY3_1),.clk(gclk));
	jdff dff_B_1K76nVgS4_1(.din(w_dff_B_Hb4m2qnY3_1),.dout(w_dff_B_1K76nVgS4_1),.clk(gclk));
	jdff dff_B_eoP3Yex09_1(.din(w_dff_B_1K76nVgS4_1),.dout(w_dff_B_eoP3Yex09_1),.clk(gclk));
	jdff dff_B_2Uj1LSKp3_1(.din(w_dff_B_eoP3Yex09_1),.dout(w_dff_B_2Uj1LSKp3_1),.clk(gclk));
	jdff dff_B_ghSR0Zmw4_1(.din(w_dff_B_2Uj1LSKp3_1),.dout(w_dff_B_ghSR0Zmw4_1),.clk(gclk));
	jdff dff_B_5RaPRw7l4_1(.din(w_dff_B_ghSR0Zmw4_1),.dout(w_dff_B_5RaPRw7l4_1),.clk(gclk));
	jdff dff_B_27uAV64G6_1(.din(w_dff_B_5RaPRw7l4_1),.dout(w_dff_B_27uAV64G6_1),.clk(gclk));
	jdff dff_B_JgpuGL5Q5_1(.din(w_dff_B_27uAV64G6_1),.dout(w_dff_B_JgpuGL5Q5_1),.clk(gclk));
	jdff dff_B_7N4MKayX3_1(.din(w_dff_B_JgpuGL5Q5_1),.dout(w_dff_B_7N4MKayX3_1),.clk(gclk));
	jdff dff_B_GhL8ah425_1(.din(w_dff_B_7N4MKayX3_1),.dout(w_dff_B_GhL8ah425_1),.clk(gclk));
	jdff dff_B_IGujUGsJ2_1(.din(w_dff_B_GhL8ah425_1),.dout(w_dff_B_IGujUGsJ2_1),.clk(gclk));
	jdff dff_B_gesBFxlK8_1(.din(w_dff_B_IGujUGsJ2_1),.dout(w_dff_B_gesBFxlK8_1),.clk(gclk));
	jdff dff_B_5Mzt9yVe4_1(.din(w_dff_B_gesBFxlK8_1),.dout(w_dff_B_5Mzt9yVe4_1),.clk(gclk));
	jdff dff_B_3672zwHl0_1(.din(w_dff_B_5Mzt9yVe4_1),.dout(w_dff_B_3672zwHl0_1),.clk(gclk));
	jdff dff_B_OsJ4Xwr37_1(.din(w_dff_B_3672zwHl0_1),.dout(w_dff_B_OsJ4Xwr37_1),.clk(gclk));
	jdff dff_B_MjGSkulR6_1(.din(w_dff_B_OsJ4Xwr37_1),.dout(w_dff_B_MjGSkulR6_1),.clk(gclk));
	jdff dff_B_TmOPLkar1_1(.din(w_dff_B_MjGSkulR6_1),.dout(w_dff_B_TmOPLkar1_1),.clk(gclk));
	jdff dff_B_T9xEWAhQ2_1(.din(w_dff_B_TmOPLkar1_1),.dout(w_dff_B_T9xEWAhQ2_1),.clk(gclk));
	jdff dff_B_c8fB6bqp0_1(.din(w_dff_B_T9xEWAhQ2_1),.dout(w_dff_B_c8fB6bqp0_1),.clk(gclk));
	jdff dff_B_cjFPaJhc7_1(.din(w_dff_B_c8fB6bqp0_1),.dout(w_dff_B_cjFPaJhc7_1),.clk(gclk));
	jdff dff_B_do1dJ43T8_1(.din(w_dff_B_cjFPaJhc7_1),.dout(w_dff_B_do1dJ43T8_1),.clk(gclk));
	jdff dff_B_lG5DkX6d0_1(.din(w_dff_B_do1dJ43T8_1),.dout(w_dff_B_lG5DkX6d0_1),.clk(gclk));
	jdff dff_B_Tf7WMqGk9_1(.din(w_dff_B_lG5DkX6d0_1),.dout(w_dff_B_Tf7WMqGk9_1),.clk(gclk));
	jdff dff_B_oG1alkJt9_1(.din(w_dff_B_Tf7WMqGk9_1),.dout(w_dff_B_oG1alkJt9_1),.clk(gclk));
	jdff dff_B_dBdjK4Go2_0(.din(n727),.dout(w_dff_B_dBdjK4Go2_0),.clk(gclk));
	jdff dff_B_wyPIm1UZ3_0(.din(w_dff_B_dBdjK4Go2_0),.dout(w_dff_B_wyPIm1UZ3_0),.clk(gclk));
	jdff dff_B_BjFyTSEJ1_0(.din(w_dff_B_wyPIm1UZ3_0),.dout(w_dff_B_BjFyTSEJ1_0),.clk(gclk));
	jdff dff_B_jXLLyTQO5_0(.din(w_dff_B_BjFyTSEJ1_0),.dout(w_dff_B_jXLLyTQO5_0),.clk(gclk));
	jdff dff_B_OMiCFaPv5_0(.din(w_dff_B_jXLLyTQO5_0),.dout(w_dff_B_OMiCFaPv5_0),.clk(gclk));
	jdff dff_B_OP7PK68l7_0(.din(w_dff_B_OMiCFaPv5_0),.dout(w_dff_B_OP7PK68l7_0),.clk(gclk));
	jdff dff_B_FpX1ZdTa1_0(.din(w_dff_B_OP7PK68l7_0),.dout(w_dff_B_FpX1ZdTa1_0),.clk(gclk));
	jdff dff_B_8DMekzTk8_0(.din(w_dff_B_FpX1ZdTa1_0),.dout(w_dff_B_8DMekzTk8_0),.clk(gclk));
	jdff dff_B_G4sePo7S0_0(.din(w_dff_B_8DMekzTk8_0),.dout(w_dff_B_G4sePo7S0_0),.clk(gclk));
	jdff dff_B_t8rmk72t4_0(.din(w_dff_B_G4sePo7S0_0),.dout(w_dff_B_t8rmk72t4_0),.clk(gclk));
	jdff dff_B_LlxRW8C52_0(.din(w_dff_B_t8rmk72t4_0),.dout(w_dff_B_LlxRW8C52_0),.clk(gclk));
	jdff dff_B_Ky9pUCVw5_0(.din(w_dff_B_LlxRW8C52_0),.dout(w_dff_B_Ky9pUCVw5_0),.clk(gclk));
	jdff dff_B_Oy0NuylO8_0(.din(w_dff_B_Ky9pUCVw5_0),.dout(w_dff_B_Oy0NuylO8_0),.clk(gclk));
	jdff dff_B_2noy2oTJ2_0(.din(w_dff_B_Oy0NuylO8_0),.dout(w_dff_B_2noy2oTJ2_0),.clk(gclk));
	jdff dff_B_dLBVVI7u3_0(.din(w_dff_B_2noy2oTJ2_0),.dout(w_dff_B_dLBVVI7u3_0),.clk(gclk));
	jdff dff_B_NRbQ4r6x2_0(.din(w_dff_B_dLBVVI7u3_0),.dout(w_dff_B_NRbQ4r6x2_0),.clk(gclk));
	jdff dff_B_NBvesLd92_0(.din(w_dff_B_NRbQ4r6x2_0),.dout(w_dff_B_NBvesLd92_0),.clk(gclk));
	jdff dff_B_K3H4kZND4_0(.din(w_dff_B_NBvesLd92_0),.dout(w_dff_B_K3H4kZND4_0),.clk(gclk));
	jdff dff_B_MjByZoJH9_0(.din(w_dff_B_K3H4kZND4_0),.dout(w_dff_B_MjByZoJH9_0),.clk(gclk));
	jdff dff_B_56sHsrca8_0(.din(w_dff_B_MjByZoJH9_0),.dout(w_dff_B_56sHsrca8_0),.clk(gclk));
	jdff dff_B_cwC5cs5I1_0(.din(w_dff_B_56sHsrca8_0),.dout(w_dff_B_cwC5cs5I1_0),.clk(gclk));
	jdff dff_B_g9qqL6A16_0(.din(w_dff_B_cwC5cs5I1_0),.dout(w_dff_B_g9qqL6A16_0),.clk(gclk));
	jdff dff_B_TuWm4ZfD5_0(.din(w_dff_B_g9qqL6A16_0),.dout(w_dff_B_TuWm4ZfD5_0),.clk(gclk));
	jdff dff_B_4xiv5mHj9_0(.din(w_dff_B_TuWm4ZfD5_0),.dout(w_dff_B_4xiv5mHj9_0),.clk(gclk));
	jdff dff_B_YRzchkIR9_0(.din(w_dff_B_4xiv5mHj9_0),.dout(w_dff_B_YRzchkIR9_0),.clk(gclk));
	jdff dff_B_K74nRoLS3_0(.din(w_dff_B_YRzchkIR9_0),.dout(w_dff_B_K74nRoLS3_0),.clk(gclk));
	jdff dff_B_cLWezrlL6_0(.din(w_dff_B_K74nRoLS3_0),.dout(w_dff_B_cLWezrlL6_0),.clk(gclk));
	jdff dff_B_qcSg3F8k4_0(.din(w_dff_B_cLWezrlL6_0),.dout(w_dff_B_qcSg3F8k4_0),.clk(gclk));
	jdff dff_B_3aZscX4A1_0(.din(w_dff_B_qcSg3F8k4_0),.dout(w_dff_B_3aZscX4A1_0),.clk(gclk));
	jdff dff_B_s7nhyX6k9_0(.din(w_dff_B_3aZscX4A1_0),.dout(w_dff_B_s7nhyX6k9_0),.clk(gclk));
	jdff dff_B_rTPn8nXI6_0(.din(w_dff_B_s7nhyX6k9_0),.dout(w_dff_B_rTPn8nXI6_0),.clk(gclk));
	jdff dff_B_kGnHDunW8_0(.din(w_dff_B_rTPn8nXI6_0),.dout(w_dff_B_kGnHDunW8_0),.clk(gclk));
	jdff dff_B_dQRXvK4c9_0(.din(w_dff_B_kGnHDunW8_0),.dout(w_dff_B_dQRXvK4c9_0),.clk(gclk));
	jdff dff_B_LPBJXOcQ8_0(.din(w_dff_B_dQRXvK4c9_0),.dout(w_dff_B_LPBJXOcQ8_0),.clk(gclk));
	jdff dff_B_b5AQC59K3_0(.din(w_dff_B_LPBJXOcQ8_0),.dout(w_dff_B_b5AQC59K3_0),.clk(gclk));
	jdff dff_B_dhivIDxT2_0(.din(w_dff_B_b5AQC59K3_0),.dout(w_dff_B_dhivIDxT2_0),.clk(gclk));
	jdff dff_B_6vd3IVKb2_0(.din(w_dff_B_dhivIDxT2_0),.dout(w_dff_B_6vd3IVKb2_0),.clk(gclk));
	jdff dff_B_P0g11IjR1_0(.din(w_dff_B_6vd3IVKb2_0),.dout(w_dff_B_P0g11IjR1_0),.clk(gclk));
	jdff dff_B_DGjguLL43_0(.din(w_dff_B_P0g11IjR1_0),.dout(w_dff_B_DGjguLL43_0),.clk(gclk));
	jdff dff_B_dTFCTEre2_0(.din(w_dff_B_DGjguLL43_0),.dout(w_dff_B_dTFCTEre2_0),.clk(gclk));
	jdff dff_B_ciAR4HWn8_0(.din(w_dff_B_dTFCTEre2_0),.dout(w_dff_B_ciAR4HWn8_0),.clk(gclk));
	jdff dff_B_IbE5Bi4l7_0(.din(w_dff_B_ciAR4HWn8_0),.dout(w_dff_B_IbE5Bi4l7_0),.clk(gclk));
	jdff dff_B_Q59msCFu4_0(.din(w_dff_B_IbE5Bi4l7_0),.dout(w_dff_B_Q59msCFu4_0),.clk(gclk));
	jdff dff_B_jXcU14ww5_0(.din(w_dff_B_Q59msCFu4_0),.dout(w_dff_B_jXcU14ww5_0),.clk(gclk));
	jdff dff_B_eWohGabJ7_0(.din(w_dff_B_jXcU14ww5_0),.dout(w_dff_B_eWohGabJ7_0),.clk(gclk));
	jdff dff_B_T7F6FABL1_0(.din(w_dff_B_eWohGabJ7_0),.dout(w_dff_B_T7F6FABL1_0),.clk(gclk));
	jdff dff_B_2JdPZ1OT5_0(.din(w_dff_B_T7F6FABL1_0),.dout(w_dff_B_2JdPZ1OT5_0),.clk(gclk));
	jdff dff_B_4NRa4jZy9_0(.din(w_dff_B_2JdPZ1OT5_0),.dout(w_dff_B_4NRa4jZy9_0),.clk(gclk));
	jdff dff_B_q8M4SDgg7_0(.din(w_dff_B_4NRa4jZy9_0),.dout(w_dff_B_q8M4SDgg7_0),.clk(gclk));
	jdff dff_B_NMOeFRYK4_0(.din(w_dff_B_q8M4SDgg7_0),.dout(w_dff_B_NMOeFRYK4_0),.clk(gclk));
	jdff dff_B_Ju8OmXTI0_0(.din(w_dff_B_NMOeFRYK4_0),.dout(w_dff_B_Ju8OmXTI0_0),.clk(gclk));
	jdff dff_B_Iwn6LkHQ1_0(.din(w_dff_B_Ju8OmXTI0_0),.dout(w_dff_B_Iwn6LkHQ1_0),.clk(gclk));
	jdff dff_B_pvhokLI60_0(.din(w_dff_B_Iwn6LkHQ1_0),.dout(w_dff_B_pvhokLI60_0),.clk(gclk));
	jdff dff_B_YdQR1MtD3_0(.din(w_dff_B_pvhokLI60_0),.dout(w_dff_B_YdQR1MtD3_0),.clk(gclk));
	jdff dff_B_MuFHsWWb0_0(.din(w_dff_B_YdQR1MtD3_0),.dout(w_dff_B_MuFHsWWb0_0),.clk(gclk));
	jdff dff_B_DJknTa6t8_0(.din(w_dff_B_MuFHsWWb0_0),.dout(w_dff_B_DJknTa6t8_0),.clk(gclk));
	jdff dff_B_y4LeRC6T7_0(.din(w_dff_B_DJknTa6t8_0),.dout(w_dff_B_y4LeRC6T7_0),.clk(gclk));
	jdff dff_B_GpWeFU1s5_1(.din(n720),.dout(w_dff_B_GpWeFU1s5_1),.clk(gclk));
	jdff dff_B_FgTKZoKY3_1(.din(w_dff_B_GpWeFU1s5_1),.dout(w_dff_B_FgTKZoKY3_1),.clk(gclk));
	jdff dff_B_aiiSi7yj2_1(.din(w_dff_B_FgTKZoKY3_1),.dout(w_dff_B_aiiSi7yj2_1),.clk(gclk));
	jdff dff_B_k9uGIfOT2_1(.din(w_dff_B_aiiSi7yj2_1),.dout(w_dff_B_k9uGIfOT2_1),.clk(gclk));
	jdff dff_B_VsnQUbqM6_1(.din(w_dff_B_k9uGIfOT2_1),.dout(w_dff_B_VsnQUbqM6_1),.clk(gclk));
	jdff dff_B_H86GVT4Y9_1(.din(w_dff_B_VsnQUbqM6_1),.dout(w_dff_B_H86GVT4Y9_1),.clk(gclk));
	jdff dff_B_noW4LybY3_1(.din(w_dff_B_H86GVT4Y9_1),.dout(w_dff_B_noW4LybY3_1),.clk(gclk));
	jdff dff_B_v5JRCwk38_1(.din(w_dff_B_noW4LybY3_1),.dout(w_dff_B_v5JRCwk38_1),.clk(gclk));
	jdff dff_B_WZSkCvgY7_1(.din(w_dff_B_v5JRCwk38_1),.dout(w_dff_B_WZSkCvgY7_1),.clk(gclk));
	jdff dff_B_zhg9jDwQ9_1(.din(w_dff_B_WZSkCvgY7_1),.dout(w_dff_B_zhg9jDwQ9_1),.clk(gclk));
	jdff dff_B_dI8eMT2e2_1(.din(w_dff_B_zhg9jDwQ9_1),.dout(w_dff_B_dI8eMT2e2_1),.clk(gclk));
	jdff dff_B_OOl40zg64_1(.din(w_dff_B_dI8eMT2e2_1),.dout(w_dff_B_OOl40zg64_1),.clk(gclk));
	jdff dff_B_a2jHVhPZ4_1(.din(w_dff_B_OOl40zg64_1),.dout(w_dff_B_a2jHVhPZ4_1),.clk(gclk));
	jdff dff_B_2ew70LjY4_1(.din(w_dff_B_a2jHVhPZ4_1),.dout(w_dff_B_2ew70LjY4_1),.clk(gclk));
	jdff dff_B_2QNNBvTf6_1(.din(w_dff_B_2ew70LjY4_1),.dout(w_dff_B_2QNNBvTf6_1),.clk(gclk));
	jdff dff_B_sFOQtUNk8_1(.din(w_dff_B_2QNNBvTf6_1),.dout(w_dff_B_sFOQtUNk8_1),.clk(gclk));
	jdff dff_B_87nCt9bA0_1(.din(w_dff_B_sFOQtUNk8_1),.dout(w_dff_B_87nCt9bA0_1),.clk(gclk));
	jdff dff_B_buDyeB7T7_1(.din(w_dff_B_87nCt9bA0_1),.dout(w_dff_B_buDyeB7T7_1),.clk(gclk));
	jdff dff_B_6KmE9TuB0_1(.din(w_dff_B_buDyeB7T7_1),.dout(w_dff_B_6KmE9TuB0_1),.clk(gclk));
	jdff dff_B_eVO0fgWg6_1(.din(w_dff_B_6KmE9TuB0_1),.dout(w_dff_B_eVO0fgWg6_1),.clk(gclk));
	jdff dff_B_NQZZxeGt0_1(.din(w_dff_B_eVO0fgWg6_1),.dout(w_dff_B_NQZZxeGt0_1),.clk(gclk));
	jdff dff_B_daK270jr9_1(.din(w_dff_B_NQZZxeGt0_1),.dout(w_dff_B_daK270jr9_1),.clk(gclk));
	jdff dff_B_Ehbjd6Ch0_1(.din(w_dff_B_daK270jr9_1),.dout(w_dff_B_Ehbjd6Ch0_1),.clk(gclk));
	jdff dff_B_MniuClbY7_1(.din(w_dff_B_Ehbjd6Ch0_1),.dout(w_dff_B_MniuClbY7_1),.clk(gclk));
	jdff dff_B_3uFndIfq4_1(.din(w_dff_B_MniuClbY7_1),.dout(w_dff_B_3uFndIfq4_1),.clk(gclk));
	jdff dff_B_NGaQbojq4_1(.din(w_dff_B_3uFndIfq4_1),.dout(w_dff_B_NGaQbojq4_1),.clk(gclk));
	jdff dff_B_IiwrG0eu4_1(.din(w_dff_B_NGaQbojq4_1),.dout(w_dff_B_IiwrG0eu4_1),.clk(gclk));
	jdff dff_B_v5Inhmz92_1(.din(w_dff_B_IiwrG0eu4_1),.dout(w_dff_B_v5Inhmz92_1),.clk(gclk));
	jdff dff_B_3x5CRNck3_1(.din(w_dff_B_v5Inhmz92_1),.dout(w_dff_B_3x5CRNck3_1),.clk(gclk));
	jdff dff_B_dPvXVYw16_1(.din(w_dff_B_3x5CRNck3_1),.dout(w_dff_B_dPvXVYw16_1),.clk(gclk));
	jdff dff_B_x6ouehoS0_1(.din(w_dff_B_dPvXVYw16_1),.dout(w_dff_B_x6ouehoS0_1),.clk(gclk));
	jdff dff_B_Py0FRrTG8_1(.din(w_dff_B_x6ouehoS0_1),.dout(w_dff_B_Py0FRrTG8_1),.clk(gclk));
	jdff dff_B_vZXReVgw5_1(.din(w_dff_B_Py0FRrTG8_1),.dout(w_dff_B_vZXReVgw5_1),.clk(gclk));
	jdff dff_B_T7n84AaM3_1(.din(w_dff_B_vZXReVgw5_1),.dout(w_dff_B_T7n84AaM3_1),.clk(gclk));
	jdff dff_B_vYEUeJoc9_1(.din(w_dff_B_T7n84AaM3_1),.dout(w_dff_B_vYEUeJoc9_1),.clk(gclk));
	jdff dff_B_2T110TmO9_1(.din(w_dff_B_vYEUeJoc9_1),.dout(w_dff_B_2T110TmO9_1),.clk(gclk));
	jdff dff_B_GCyTDkA14_1(.din(w_dff_B_2T110TmO9_1),.dout(w_dff_B_GCyTDkA14_1),.clk(gclk));
	jdff dff_B_sNmnjWOY1_1(.din(w_dff_B_GCyTDkA14_1),.dout(w_dff_B_sNmnjWOY1_1),.clk(gclk));
	jdff dff_B_YEnXssFw8_1(.din(w_dff_B_sNmnjWOY1_1),.dout(w_dff_B_YEnXssFw8_1),.clk(gclk));
	jdff dff_B_0iwNGo6Z5_1(.din(w_dff_B_YEnXssFw8_1),.dout(w_dff_B_0iwNGo6Z5_1),.clk(gclk));
	jdff dff_B_9V7Hm9qW8_1(.din(w_dff_B_0iwNGo6Z5_1),.dout(w_dff_B_9V7Hm9qW8_1),.clk(gclk));
	jdff dff_B_pKtxPdUH5_1(.din(w_dff_B_9V7Hm9qW8_1),.dout(w_dff_B_pKtxPdUH5_1),.clk(gclk));
	jdff dff_B_U05Knw5y5_1(.din(w_dff_B_pKtxPdUH5_1),.dout(w_dff_B_U05Knw5y5_1),.clk(gclk));
	jdff dff_B_pzI1WzRe5_1(.din(w_dff_B_U05Knw5y5_1),.dout(w_dff_B_pzI1WzRe5_1),.clk(gclk));
	jdff dff_B_98pEpBOP1_1(.din(w_dff_B_pzI1WzRe5_1),.dout(w_dff_B_98pEpBOP1_1),.clk(gclk));
	jdff dff_B_3VVTgbij2_1(.din(w_dff_B_98pEpBOP1_1),.dout(w_dff_B_3VVTgbij2_1),.clk(gclk));
	jdff dff_B_dsFFpdN42_1(.din(w_dff_B_3VVTgbij2_1),.dout(w_dff_B_dsFFpdN42_1),.clk(gclk));
	jdff dff_B_QdYTwScb1_1(.din(w_dff_B_dsFFpdN42_1),.dout(w_dff_B_QdYTwScb1_1),.clk(gclk));
	jdff dff_B_IAurgHSJ4_1(.din(w_dff_B_QdYTwScb1_1),.dout(w_dff_B_IAurgHSJ4_1),.clk(gclk));
	jdff dff_B_BgMUHX8R5_1(.din(w_dff_B_IAurgHSJ4_1),.dout(w_dff_B_BgMUHX8R5_1),.clk(gclk));
	jdff dff_B_yCjwOozj4_1(.din(w_dff_B_BgMUHX8R5_1),.dout(w_dff_B_yCjwOozj4_1),.clk(gclk));
	jdff dff_B_OQj0EPzU8_1(.din(w_dff_B_yCjwOozj4_1),.dout(w_dff_B_OQj0EPzU8_1),.clk(gclk));
	jdff dff_B_OUMAHm6x3_1(.din(w_dff_B_OQj0EPzU8_1),.dout(w_dff_B_OUMAHm6x3_1),.clk(gclk));
	jdff dff_B_CW9Chxyz6_1(.din(w_dff_B_OUMAHm6x3_1),.dout(w_dff_B_CW9Chxyz6_1),.clk(gclk));
	jdff dff_B_PhaSoyuf9_1(.din(w_dff_B_CW9Chxyz6_1),.dout(w_dff_B_PhaSoyuf9_1),.clk(gclk));
	jdff dff_B_7hG8iOrA5_1(.din(w_dff_B_PhaSoyuf9_1),.dout(w_dff_B_7hG8iOrA5_1),.clk(gclk));
	jdff dff_B_lCwjjydv0_0(.din(n721),.dout(w_dff_B_lCwjjydv0_0),.clk(gclk));
	jdff dff_B_ucmcO5Ml9_0(.din(w_dff_B_lCwjjydv0_0),.dout(w_dff_B_ucmcO5Ml9_0),.clk(gclk));
	jdff dff_B_0mLqRJyn2_0(.din(w_dff_B_ucmcO5Ml9_0),.dout(w_dff_B_0mLqRJyn2_0),.clk(gclk));
	jdff dff_B_7nWxuOlI8_0(.din(w_dff_B_0mLqRJyn2_0),.dout(w_dff_B_7nWxuOlI8_0),.clk(gclk));
	jdff dff_B_qAiuHkW09_0(.din(w_dff_B_7nWxuOlI8_0),.dout(w_dff_B_qAiuHkW09_0),.clk(gclk));
	jdff dff_B_XoioK0yV9_0(.din(w_dff_B_qAiuHkW09_0),.dout(w_dff_B_XoioK0yV9_0),.clk(gclk));
	jdff dff_B_9GQ1TgWU3_0(.din(w_dff_B_XoioK0yV9_0),.dout(w_dff_B_9GQ1TgWU3_0),.clk(gclk));
	jdff dff_B_59gJDSWg4_0(.din(w_dff_B_9GQ1TgWU3_0),.dout(w_dff_B_59gJDSWg4_0),.clk(gclk));
	jdff dff_B_Fqri8rU17_0(.din(w_dff_B_59gJDSWg4_0),.dout(w_dff_B_Fqri8rU17_0),.clk(gclk));
	jdff dff_B_fusZp0wO4_0(.din(w_dff_B_Fqri8rU17_0),.dout(w_dff_B_fusZp0wO4_0),.clk(gclk));
	jdff dff_B_qfiPzsTJ0_0(.din(w_dff_B_fusZp0wO4_0),.dout(w_dff_B_qfiPzsTJ0_0),.clk(gclk));
	jdff dff_B_1IHRjypV6_0(.din(w_dff_B_qfiPzsTJ0_0),.dout(w_dff_B_1IHRjypV6_0),.clk(gclk));
	jdff dff_B_Mt73eZIK8_0(.din(w_dff_B_1IHRjypV6_0),.dout(w_dff_B_Mt73eZIK8_0),.clk(gclk));
	jdff dff_B_L8tAwmN70_0(.din(w_dff_B_Mt73eZIK8_0),.dout(w_dff_B_L8tAwmN70_0),.clk(gclk));
	jdff dff_B_Rg5dGiZJ9_0(.din(w_dff_B_L8tAwmN70_0),.dout(w_dff_B_Rg5dGiZJ9_0),.clk(gclk));
	jdff dff_B_U09o2vKe9_0(.din(w_dff_B_Rg5dGiZJ9_0),.dout(w_dff_B_U09o2vKe9_0),.clk(gclk));
	jdff dff_B_UBub5VMl4_0(.din(w_dff_B_U09o2vKe9_0),.dout(w_dff_B_UBub5VMl4_0),.clk(gclk));
	jdff dff_B_Y5Hjnyb33_0(.din(w_dff_B_UBub5VMl4_0),.dout(w_dff_B_Y5Hjnyb33_0),.clk(gclk));
	jdff dff_B_izX1EhWs3_0(.din(w_dff_B_Y5Hjnyb33_0),.dout(w_dff_B_izX1EhWs3_0),.clk(gclk));
	jdff dff_B_GFojTKFQ4_0(.din(w_dff_B_izX1EhWs3_0),.dout(w_dff_B_GFojTKFQ4_0),.clk(gclk));
	jdff dff_B_HgByJuwt0_0(.din(w_dff_B_GFojTKFQ4_0),.dout(w_dff_B_HgByJuwt0_0),.clk(gclk));
	jdff dff_B_AAhMz0cT7_0(.din(w_dff_B_HgByJuwt0_0),.dout(w_dff_B_AAhMz0cT7_0),.clk(gclk));
	jdff dff_B_IVtehnJB2_0(.din(w_dff_B_AAhMz0cT7_0),.dout(w_dff_B_IVtehnJB2_0),.clk(gclk));
	jdff dff_B_ppAay2wQ0_0(.din(w_dff_B_IVtehnJB2_0),.dout(w_dff_B_ppAay2wQ0_0),.clk(gclk));
	jdff dff_B_fvd8OPgU6_0(.din(w_dff_B_ppAay2wQ0_0),.dout(w_dff_B_fvd8OPgU6_0),.clk(gclk));
	jdff dff_B_ud6T4sad7_0(.din(w_dff_B_fvd8OPgU6_0),.dout(w_dff_B_ud6T4sad7_0),.clk(gclk));
	jdff dff_B_R2RMJGAo2_0(.din(w_dff_B_ud6T4sad7_0),.dout(w_dff_B_R2RMJGAo2_0),.clk(gclk));
	jdff dff_B_Udu3LCzL3_0(.din(w_dff_B_R2RMJGAo2_0),.dout(w_dff_B_Udu3LCzL3_0),.clk(gclk));
	jdff dff_B_cPRnuFfU0_0(.din(w_dff_B_Udu3LCzL3_0),.dout(w_dff_B_cPRnuFfU0_0),.clk(gclk));
	jdff dff_B_VfYi89cV3_0(.din(w_dff_B_cPRnuFfU0_0),.dout(w_dff_B_VfYi89cV3_0),.clk(gclk));
	jdff dff_B_crlkUjKD0_0(.din(w_dff_B_VfYi89cV3_0),.dout(w_dff_B_crlkUjKD0_0),.clk(gclk));
	jdff dff_B_lnwW7c1Z6_0(.din(w_dff_B_crlkUjKD0_0),.dout(w_dff_B_lnwW7c1Z6_0),.clk(gclk));
	jdff dff_B_MjnPmnjI0_0(.din(w_dff_B_lnwW7c1Z6_0),.dout(w_dff_B_MjnPmnjI0_0),.clk(gclk));
	jdff dff_B_5rPxPaU28_0(.din(w_dff_B_MjnPmnjI0_0),.dout(w_dff_B_5rPxPaU28_0),.clk(gclk));
	jdff dff_B_TAYMsVAj8_0(.din(w_dff_B_5rPxPaU28_0),.dout(w_dff_B_TAYMsVAj8_0),.clk(gclk));
	jdff dff_B_m0gHZEVP0_0(.din(w_dff_B_TAYMsVAj8_0),.dout(w_dff_B_m0gHZEVP0_0),.clk(gclk));
	jdff dff_B_CHvgD6cr3_0(.din(w_dff_B_m0gHZEVP0_0),.dout(w_dff_B_CHvgD6cr3_0),.clk(gclk));
	jdff dff_B_Swy415Fb5_0(.din(w_dff_B_CHvgD6cr3_0),.dout(w_dff_B_Swy415Fb5_0),.clk(gclk));
	jdff dff_B_rS4why0S1_0(.din(w_dff_B_Swy415Fb5_0),.dout(w_dff_B_rS4why0S1_0),.clk(gclk));
	jdff dff_B_FAS5VmN86_0(.din(w_dff_B_rS4why0S1_0),.dout(w_dff_B_FAS5VmN86_0),.clk(gclk));
	jdff dff_B_8bMGc5ws7_0(.din(w_dff_B_FAS5VmN86_0),.dout(w_dff_B_8bMGc5ws7_0),.clk(gclk));
	jdff dff_B_TamJ9C3q4_0(.din(w_dff_B_8bMGc5ws7_0),.dout(w_dff_B_TamJ9C3q4_0),.clk(gclk));
	jdff dff_B_EDiQGhZA2_0(.din(w_dff_B_TamJ9C3q4_0),.dout(w_dff_B_EDiQGhZA2_0),.clk(gclk));
	jdff dff_B_tG9RCre11_0(.din(w_dff_B_EDiQGhZA2_0),.dout(w_dff_B_tG9RCre11_0),.clk(gclk));
	jdff dff_B_9HgKTcxd6_0(.din(w_dff_B_tG9RCre11_0),.dout(w_dff_B_9HgKTcxd6_0),.clk(gclk));
	jdff dff_B_jE0d3Y2q4_0(.din(w_dff_B_9HgKTcxd6_0),.dout(w_dff_B_jE0d3Y2q4_0),.clk(gclk));
	jdff dff_B_IewIwsfG9_0(.din(w_dff_B_jE0d3Y2q4_0),.dout(w_dff_B_IewIwsfG9_0),.clk(gclk));
	jdff dff_B_u20dojIx1_0(.din(w_dff_B_IewIwsfG9_0),.dout(w_dff_B_u20dojIx1_0),.clk(gclk));
	jdff dff_B_4pg06WGH8_0(.din(w_dff_B_u20dojIx1_0),.dout(w_dff_B_4pg06WGH8_0),.clk(gclk));
	jdff dff_B_3KJRWdtl7_0(.din(w_dff_B_4pg06WGH8_0),.dout(w_dff_B_3KJRWdtl7_0),.clk(gclk));
	jdff dff_B_EFceaqyR5_0(.din(w_dff_B_3KJRWdtl7_0),.dout(w_dff_B_EFceaqyR5_0),.clk(gclk));
	jdff dff_B_J9OGBn7A9_0(.din(w_dff_B_EFceaqyR5_0),.dout(w_dff_B_J9OGBn7A9_0),.clk(gclk));
	jdff dff_B_nN040jiK9_0(.din(w_dff_B_J9OGBn7A9_0),.dout(w_dff_B_nN040jiK9_0),.clk(gclk));
	jdff dff_B_tVW8F4P63_0(.din(w_dff_B_nN040jiK9_0),.dout(w_dff_B_tVW8F4P63_0),.clk(gclk));
	jdff dff_B_qRjaLalN4_0(.din(w_dff_B_tVW8F4P63_0),.dout(w_dff_B_qRjaLalN4_0),.clk(gclk));
	jdff dff_B_3PM2Wo7i4_0(.din(w_dff_B_qRjaLalN4_0),.dout(w_dff_B_3PM2Wo7i4_0),.clk(gclk));
	jdff dff_B_u3TmHQQg3_1(.din(n714),.dout(w_dff_B_u3TmHQQg3_1),.clk(gclk));
	jdff dff_B_WyI1cjee2_1(.din(w_dff_B_u3TmHQQg3_1),.dout(w_dff_B_WyI1cjee2_1),.clk(gclk));
	jdff dff_B_QwI2VE026_1(.din(w_dff_B_WyI1cjee2_1),.dout(w_dff_B_QwI2VE026_1),.clk(gclk));
	jdff dff_B_f3OOC1vX5_1(.din(w_dff_B_QwI2VE026_1),.dout(w_dff_B_f3OOC1vX5_1),.clk(gclk));
	jdff dff_B_kObOhMPQ6_1(.din(w_dff_B_f3OOC1vX5_1),.dout(w_dff_B_kObOhMPQ6_1),.clk(gclk));
	jdff dff_B_UXXiYhTZ7_1(.din(w_dff_B_kObOhMPQ6_1),.dout(w_dff_B_UXXiYhTZ7_1),.clk(gclk));
	jdff dff_B_vSzIN6NW1_1(.din(w_dff_B_UXXiYhTZ7_1),.dout(w_dff_B_vSzIN6NW1_1),.clk(gclk));
	jdff dff_B_zx7wZkaR9_1(.din(w_dff_B_vSzIN6NW1_1),.dout(w_dff_B_zx7wZkaR9_1),.clk(gclk));
	jdff dff_B_qjQmHTsH3_1(.din(w_dff_B_zx7wZkaR9_1),.dout(w_dff_B_qjQmHTsH3_1),.clk(gclk));
	jdff dff_B_gxCBoZzF0_1(.din(w_dff_B_qjQmHTsH3_1),.dout(w_dff_B_gxCBoZzF0_1),.clk(gclk));
	jdff dff_B_T1Nxxa6N3_1(.din(w_dff_B_gxCBoZzF0_1),.dout(w_dff_B_T1Nxxa6N3_1),.clk(gclk));
	jdff dff_B_aItBSbms7_1(.din(w_dff_B_T1Nxxa6N3_1),.dout(w_dff_B_aItBSbms7_1),.clk(gclk));
	jdff dff_B_m9z39zzQ9_1(.din(w_dff_B_aItBSbms7_1),.dout(w_dff_B_m9z39zzQ9_1),.clk(gclk));
	jdff dff_B_wLFJeXXi6_1(.din(w_dff_B_m9z39zzQ9_1),.dout(w_dff_B_wLFJeXXi6_1),.clk(gclk));
	jdff dff_B_98y3Vefh8_1(.din(w_dff_B_wLFJeXXi6_1),.dout(w_dff_B_98y3Vefh8_1),.clk(gclk));
	jdff dff_B_TOqFGqCT9_1(.din(w_dff_B_98y3Vefh8_1),.dout(w_dff_B_TOqFGqCT9_1),.clk(gclk));
	jdff dff_B_WWse1KpF5_1(.din(w_dff_B_TOqFGqCT9_1),.dout(w_dff_B_WWse1KpF5_1),.clk(gclk));
	jdff dff_B_QNEaobnf7_1(.din(w_dff_B_WWse1KpF5_1),.dout(w_dff_B_QNEaobnf7_1),.clk(gclk));
	jdff dff_B_mSkhTW764_1(.din(w_dff_B_QNEaobnf7_1),.dout(w_dff_B_mSkhTW764_1),.clk(gclk));
	jdff dff_B_xMWIwYl62_1(.din(w_dff_B_mSkhTW764_1),.dout(w_dff_B_xMWIwYl62_1),.clk(gclk));
	jdff dff_B_x02PzPzH6_1(.din(w_dff_B_xMWIwYl62_1),.dout(w_dff_B_x02PzPzH6_1),.clk(gclk));
	jdff dff_B_VLUkPEy28_1(.din(w_dff_B_x02PzPzH6_1),.dout(w_dff_B_VLUkPEy28_1),.clk(gclk));
	jdff dff_B_8sX3xPsl3_1(.din(w_dff_B_VLUkPEy28_1),.dout(w_dff_B_8sX3xPsl3_1),.clk(gclk));
	jdff dff_B_GBVOD50H0_1(.din(w_dff_B_8sX3xPsl3_1),.dout(w_dff_B_GBVOD50H0_1),.clk(gclk));
	jdff dff_B_jNtNys3P5_1(.din(w_dff_B_GBVOD50H0_1),.dout(w_dff_B_jNtNys3P5_1),.clk(gclk));
	jdff dff_B_OubD3WKZ2_1(.din(w_dff_B_jNtNys3P5_1),.dout(w_dff_B_OubD3WKZ2_1),.clk(gclk));
	jdff dff_B_pcaQ4YbL7_1(.din(w_dff_B_OubD3WKZ2_1),.dout(w_dff_B_pcaQ4YbL7_1),.clk(gclk));
	jdff dff_B_7Ni4p2F14_1(.din(w_dff_B_pcaQ4YbL7_1),.dout(w_dff_B_7Ni4p2F14_1),.clk(gclk));
	jdff dff_B_URUERMh85_1(.din(w_dff_B_7Ni4p2F14_1),.dout(w_dff_B_URUERMh85_1),.clk(gclk));
	jdff dff_B_KsDpCKZB3_1(.din(w_dff_B_URUERMh85_1),.dout(w_dff_B_KsDpCKZB3_1),.clk(gclk));
	jdff dff_B_xx3DzdvC8_1(.din(w_dff_B_KsDpCKZB3_1),.dout(w_dff_B_xx3DzdvC8_1),.clk(gclk));
	jdff dff_B_3vi7eenL8_1(.din(w_dff_B_xx3DzdvC8_1),.dout(w_dff_B_3vi7eenL8_1),.clk(gclk));
	jdff dff_B_xm2P1eNU0_1(.din(w_dff_B_3vi7eenL8_1),.dout(w_dff_B_xm2P1eNU0_1),.clk(gclk));
	jdff dff_B_1hSD98Bj1_1(.din(w_dff_B_xm2P1eNU0_1),.dout(w_dff_B_1hSD98Bj1_1),.clk(gclk));
	jdff dff_B_31MJ7sCG5_1(.din(w_dff_B_1hSD98Bj1_1),.dout(w_dff_B_31MJ7sCG5_1),.clk(gclk));
	jdff dff_B_qFsfFMl80_1(.din(w_dff_B_31MJ7sCG5_1),.dout(w_dff_B_qFsfFMl80_1),.clk(gclk));
	jdff dff_B_MVByffY11_1(.din(w_dff_B_qFsfFMl80_1),.dout(w_dff_B_MVByffY11_1),.clk(gclk));
	jdff dff_B_rlPV8eVZ9_1(.din(w_dff_B_MVByffY11_1),.dout(w_dff_B_rlPV8eVZ9_1),.clk(gclk));
	jdff dff_B_iVd6ZCv73_1(.din(w_dff_B_rlPV8eVZ9_1),.dout(w_dff_B_iVd6ZCv73_1),.clk(gclk));
	jdff dff_B_XQftyCr26_1(.din(w_dff_B_iVd6ZCv73_1),.dout(w_dff_B_XQftyCr26_1),.clk(gclk));
	jdff dff_B_bCEJJ1tn6_1(.din(w_dff_B_XQftyCr26_1),.dout(w_dff_B_bCEJJ1tn6_1),.clk(gclk));
	jdff dff_B_N7h1wGxT8_1(.din(w_dff_B_bCEJJ1tn6_1),.dout(w_dff_B_N7h1wGxT8_1),.clk(gclk));
	jdff dff_B_YXV3KCnD0_1(.din(w_dff_B_N7h1wGxT8_1),.dout(w_dff_B_YXV3KCnD0_1),.clk(gclk));
	jdff dff_B_W7Dg6nDB7_1(.din(w_dff_B_YXV3KCnD0_1),.dout(w_dff_B_W7Dg6nDB7_1),.clk(gclk));
	jdff dff_B_jdkH2UOj7_1(.din(w_dff_B_W7Dg6nDB7_1),.dout(w_dff_B_jdkH2UOj7_1),.clk(gclk));
	jdff dff_B_Ra4Icv467_1(.din(w_dff_B_jdkH2UOj7_1),.dout(w_dff_B_Ra4Icv467_1),.clk(gclk));
	jdff dff_B_oBUgjbJu4_1(.din(w_dff_B_Ra4Icv467_1),.dout(w_dff_B_oBUgjbJu4_1),.clk(gclk));
	jdff dff_B_5LUFVdB82_1(.din(w_dff_B_oBUgjbJu4_1),.dout(w_dff_B_5LUFVdB82_1),.clk(gclk));
	jdff dff_B_x8gIbswR4_1(.din(w_dff_B_5LUFVdB82_1),.dout(w_dff_B_x8gIbswR4_1),.clk(gclk));
	jdff dff_B_83yftHTo3_1(.din(w_dff_B_x8gIbswR4_1),.dout(w_dff_B_83yftHTo3_1),.clk(gclk));
	jdff dff_B_5pXggwZi5_1(.din(w_dff_B_83yftHTo3_1),.dout(w_dff_B_5pXggwZi5_1),.clk(gclk));
	jdff dff_B_S4ZFBNfZ5_1(.din(w_dff_B_5pXggwZi5_1),.dout(w_dff_B_S4ZFBNfZ5_1),.clk(gclk));
	jdff dff_B_Eq02vrvz2_1(.din(w_dff_B_S4ZFBNfZ5_1),.dout(w_dff_B_Eq02vrvz2_1),.clk(gclk));
	jdff dff_B_ObDGcnQU8_1(.din(w_dff_B_Eq02vrvz2_1),.dout(w_dff_B_ObDGcnQU8_1),.clk(gclk));
	jdff dff_B_2n0kw3zB1_1(.din(w_dff_B_ObDGcnQU8_1),.dout(w_dff_B_2n0kw3zB1_1),.clk(gclk));
	jdff dff_B_EsGJzq0m3_0(.din(n715),.dout(w_dff_B_EsGJzq0m3_0),.clk(gclk));
	jdff dff_B_sU19rznP3_0(.din(w_dff_B_EsGJzq0m3_0),.dout(w_dff_B_sU19rznP3_0),.clk(gclk));
	jdff dff_B_IPWvB2Wl9_0(.din(w_dff_B_sU19rznP3_0),.dout(w_dff_B_IPWvB2Wl9_0),.clk(gclk));
	jdff dff_B_6bizC6M54_0(.din(w_dff_B_IPWvB2Wl9_0),.dout(w_dff_B_6bizC6M54_0),.clk(gclk));
	jdff dff_B_sCD3mHk49_0(.din(w_dff_B_6bizC6M54_0),.dout(w_dff_B_sCD3mHk49_0),.clk(gclk));
	jdff dff_B_fhRiEnQz3_0(.din(w_dff_B_sCD3mHk49_0),.dout(w_dff_B_fhRiEnQz3_0),.clk(gclk));
	jdff dff_B_bmpbmBlk3_0(.din(w_dff_B_fhRiEnQz3_0),.dout(w_dff_B_bmpbmBlk3_0),.clk(gclk));
	jdff dff_B_9umcwsmN4_0(.din(w_dff_B_bmpbmBlk3_0),.dout(w_dff_B_9umcwsmN4_0),.clk(gclk));
	jdff dff_B_0IDKInX46_0(.din(w_dff_B_9umcwsmN4_0),.dout(w_dff_B_0IDKInX46_0),.clk(gclk));
	jdff dff_B_LA6dKFUh9_0(.din(w_dff_B_0IDKInX46_0),.dout(w_dff_B_LA6dKFUh9_0),.clk(gclk));
	jdff dff_B_uAfYTa8O8_0(.din(w_dff_B_LA6dKFUh9_0),.dout(w_dff_B_uAfYTa8O8_0),.clk(gclk));
	jdff dff_B_g6jccsU59_0(.din(w_dff_B_uAfYTa8O8_0),.dout(w_dff_B_g6jccsU59_0),.clk(gclk));
	jdff dff_B_1iButynI2_0(.din(w_dff_B_g6jccsU59_0),.dout(w_dff_B_1iButynI2_0),.clk(gclk));
	jdff dff_B_sQowIlt83_0(.din(w_dff_B_1iButynI2_0),.dout(w_dff_B_sQowIlt83_0),.clk(gclk));
	jdff dff_B_PAiQ2VbV8_0(.din(w_dff_B_sQowIlt83_0),.dout(w_dff_B_PAiQ2VbV8_0),.clk(gclk));
	jdff dff_B_jVnUIAVA9_0(.din(w_dff_B_PAiQ2VbV8_0),.dout(w_dff_B_jVnUIAVA9_0),.clk(gclk));
	jdff dff_B_cINYgPb58_0(.din(w_dff_B_jVnUIAVA9_0),.dout(w_dff_B_cINYgPb58_0),.clk(gclk));
	jdff dff_B_rDEHEZWj5_0(.din(w_dff_B_cINYgPb58_0),.dout(w_dff_B_rDEHEZWj5_0),.clk(gclk));
	jdff dff_B_6KIz9v888_0(.din(w_dff_B_rDEHEZWj5_0),.dout(w_dff_B_6KIz9v888_0),.clk(gclk));
	jdff dff_B_JOgEGpBe8_0(.din(w_dff_B_6KIz9v888_0),.dout(w_dff_B_JOgEGpBe8_0),.clk(gclk));
	jdff dff_B_cUoiqd011_0(.din(w_dff_B_JOgEGpBe8_0),.dout(w_dff_B_cUoiqd011_0),.clk(gclk));
	jdff dff_B_n5qNuo1S7_0(.din(w_dff_B_cUoiqd011_0),.dout(w_dff_B_n5qNuo1S7_0),.clk(gclk));
	jdff dff_B_RmDJbPsU9_0(.din(w_dff_B_n5qNuo1S7_0),.dout(w_dff_B_RmDJbPsU9_0),.clk(gclk));
	jdff dff_B_sa9SjKqv1_0(.din(w_dff_B_RmDJbPsU9_0),.dout(w_dff_B_sa9SjKqv1_0),.clk(gclk));
	jdff dff_B_PBFYuqlC4_0(.din(w_dff_B_sa9SjKqv1_0),.dout(w_dff_B_PBFYuqlC4_0),.clk(gclk));
	jdff dff_B_hkSqgQ6W2_0(.din(w_dff_B_PBFYuqlC4_0),.dout(w_dff_B_hkSqgQ6W2_0),.clk(gclk));
	jdff dff_B_TwtWAeLD6_0(.din(w_dff_B_hkSqgQ6W2_0),.dout(w_dff_B_TwtWAeLD6_0),.clk(gclk));
	jdff dff_B_5YaTVtET9_0(.din(w_dff_B_TwtWAeLD6_0),.dout(w_dff_B_5YaTVtET9_0),.clk(gclk));
	jdff dff_B_VftSinlm9_0(.din(w_dff_B_5YaTVtET9_0),.dout(w_dff_B_VftSinlm9_0),.clk(gclk));
	jdff dff_B_bhnbH8kj1_0(.din(w_dff_B_VftSinlm9_0),.dout(w_dff_B_bhnbH8kj1_0),.clk(gclk));
	jdff dff_B_UxywJgzz8_0(.din(w_dff_B_bhnbH8kj1_0),.dout(w_dff_B_UxywJgzz8_0),.clk(gclk));
	jdff dff_B_OtYc43D56_0(.din(w_dff_B_UxywJgzz8_0),.dout(w_dff_B_OtYc43D56_0),.clk(gclk));
	jdff dff_B_LC9d0Ljk9_0(.din(w_dff_B_OtYc43D56_0),.dout(w_dff_B_LC9d0Ljk9_0),.clk(gclk));
	jdff dff_B_gku3dSbK8_0(.din(w_dff_B_LC9d0Ljk9_0),.dout(w_dff_B_gku3dSbK8_0),.clk(gclk));
	jdff dff_B_Rbpqcn241_0(.din(w_dff_B_gku3dSbK8_0),.dout(w_dff_B_Rbpqcn241_0),.clk(gclk));
	jdff dff_B_FDtEjWJY3_0(.din(w_dff_B_Rbpqcn241_0),.dout(w_dff_B_FDtEjWJY3_0),.clk(gclk));
	jdff dff_B_QUl09qph3_0(.din(w_dff_B_FDtEjWJY3_0),.dout(w_dff_B_QUl09qph3_0),.clk(gclk));
	jdff dff_B_AaQaOd5P7_0(.din(w_dff_B_QUl09qph3_0),.dout(w_dff_B_AaQaOd5P7_0),.clk(gclk));
	jdff dff_B_ovWruR753_0(.din(w_dff_B_AaQaOd5P7_0),.dout(w_dff_B_ovWruR753_0),.clk(gclk));
	jdff dff_B_cgX8LBHo8_0(.din(w_dff_B_ovWruR753_0),.dout(w_dff_B_cgX8LBHo8_0),.clk(gclk));
	jdff dff_B_rjylf6od7_0(.din(w_dff_B_cgX8LBHo8_0),.dout(w_dff_B_rjylf6od7_0),.clk(gclk));
	jdff dff_B_Bt632EuU5_0(.din(w_dff_B_rjylf6od7_0),.dout(w_dff_B_Bt632EuU5_0),.clk(gclk));
	jdff dff_B_WMWMEPWe4_0(.din(w_dff_B_Bt632EuU5_0),.dout(w_dff_B_WMWMEPWe4_0),.clk(gclk));
	jdff dff_B_3BR8YzSM9_0(.din(w_dff_B_WMWMEPWe4_0),.dout(w_dff_B_3BR8YzSM9_0),.clk(gclk));
	jdff dff_B_dk3ZerKI6_0(.din(w_dff_B_3BR8YzSM9_0),.dout(w_dff_B_dk3ZerKI6_0),.clk(gclk));
	jdff dff_B_i6kUDe318_0(.din(w_dff_B_dk3ZerKI6_0),.dout(w_dff_B_i6kUDe318_0),.clk(gclk));
	jdff dff_B_33Nb1gZU4_0(.din(w_dff_B_i6kUDe318_0),.dout(w_dff_B_33Nb1gZU4_0),.clk(gclk));
	jdff dff_B_EA8KARRM1_0(.din(w_dff_B_33Nb1gZU4_0),.dout(w_dff_B_EA8KARRM1_0),.clk(gclk));
	jdff dff_B_vWQAAiWQ6_0(.din(w_dff_B_EA8KARRM1_0),.dout(w_dff_B_vWQAAiWQ6_0),.clk(gclk));
	jdff dff_B_WM0tBsn91_0(.din(w_dff_B_vWQAAiWQ6_0),.dout(w_dff_B_WM0tBsn91_0),.clk(gclk));
	jdff dff_B_z8rNMEFI7_0(.din(w_dff_B_WM0tBsn91_0),.dout(w_dff_B_z8rNMEFI7_0),.clk(gclk));
	jdff dff_B_W4LRAtjG4_0(.din(w_dff_B_z8rNMEFI7_0),.dout(w_dff_B_W4LRAtjG4_0),.clk(gclk));
	jdff dff_B_n2SzxAAr1_0(.din(w_dff_B_W4LRAtjG4_0),.dout(w_dff_B_n2SzxAAr1_0),.clk(gclk));
	jdff dff_B_m5ibI5Kj7_0(.din(w_dff_B_n2SzxAAr1_0),.dout(w_dff_B_m5ibI5Kj7_0),.clk(gclk));
	jdff dff_B_krSKQ8iz1_0(.din(w_dff_B_m5ibI5Kj7_0),.dout(w_dff_B_krSKQ8iz1_0),.clk(gclk));
	jdff dff_B_b5cRaWfO3_1(.din(n708),.dout(w_dff_B_b5cRaWfO3_1),.clk(gclk));
	jdff dff_B_xlaGHZpv9_1(.din(w_dff_B_b5cRaWfO3_1),.dout(w_dff_B_xlaGHZpv9_1),.clk(gclk));
	jdff dff_B_gFzSFs251_1(.din(w_dff_B_xlaGHZpv9_1),.dout(w_dff_B_gFzSFs251_1),.clk(gclk));
	jdff dff_B_RAkB4lKs8_1(.din(w_dff_B_gFzSFs251_1),.dout(w_dff_B_RAkB4lKs8_1),.clk(gclk));
	jdff dff_B_J0A4sMAg3_1(.din(w_dff_B_RAkB4lKs8_1),.dout(w_dff_B_J0A4sMAg3_1),.clk(gclk));
	jdff dff_B_qITCs0Z54_1(.din(w_dff_B_J0A4sMAg3_1),.dout(w_dff_B_qITCs0Z54_1),.clk(gclk));
	jdff dff_B_z81S9qzx5_1(.din(w_dff_B_qITCs0Z54_1),.dout(w_dff_B_z81S9qzx5_1),.clk(gclk));
	jdff dff_B_9O7j9BaX8_1(.din(w_dff_B_z81S9qzx5_1),.dout(w_dff_B_9O7j9BaX8_1),.clk(gclk));
	jdff dff_B_eBqnDMTA3_1(.din(w_dff_B_9O7j9BaX8_1),.dout(w_dff_B_eBqnDMTA3_1),.clk(gclk));
	jdff dff_B_ZS581Y7Y7_1(.din(w_dff_B_eBqnDMTA3_1),.dout(w_dff_B_ZS581Y7Y7_1),.clk(gclk));
	jdff dff_B_RNOrmn2G3_1(.din(w_dff_B_ZS581Y7Y7_1),.dout(w_dff_B_RNOrmn2G3_1),.clk(gclk));
	jdff dff_B_GWmmUahR8_1(.din(w_dff_B_RNOrmn2G3_1),.dout(w_dff_B_GWmmUahR8_1),.clk(gclk));
	jdff dff_B_5dtNx9NK9_1(.din(w_dff_B_GWmmUahR8_1),.dout(w_dff_B_5dtNx9NK9_1),.clk(gclk));
	jdff dff_B_pHCAYkUu6_1(.din(w_dff_B_5dtNx9NK9_1),.dout(w_dff_B_pHCAYkUu6_1),.clk(gclk));
	jdff dff_B_6ooHb8145_1(.din(w_dff_B_pHCAYkUu6_1),.dout(w_dff_B_6ooHb8145_1),.clk(gclk));
	jdff dff_B_6z6YJeSJ8_1(.din(w_dff_B_6ooHb8145_1),.dout(w_dff_B_6z6YJeSJ8_1),.clk(gclk));
	jdff dff_B_ZDPkAR0O8_1(.din(w_dff_B_6z6YJeSJ8_1),.dout(w_dff_B_ZDPkAR0O8_1),.clk(gclk));
	jdff dff_B_yV5BnaNt6_1(.din(w_dff_B_ZDPkAR0O8_1),.dout(w_dff_B_yV5BnaNt6_1),.clk(gclk));
	jdff dff_B_aZkUgmSp5_1(.din(w_dff_B_yV5BnaNt6_1),.dout(w_dff_B_aZkUgmSp5_1),.clk(gclk));
	jdff dff_B_iNNRgKN24_1(.din(w_dff_B_aZkUgmSp5_1),.dout(w_dff_B_iNNRgKN24_1),.clk(gclk));
	jdff dff_B_qvEcccPS0_1(.din(w_dff_B_iNNRgKN24_1),.dout(w_dff_B_qvEcccPS0_1),.clk(gclk));
	jdff dff_B_ogrzD7CN0_1(.din(w_dff_B_qvEcccPS0_1),.dout(w_dff_B_ogrzD7CN0_1),.clk(gclk));
	jdff dff_B_V7mgggxv6_1(.din(w_dff_B_ogrzD7CN0_1),.dout(w_dff_B_V7mgggxv6_1),.clk(gclk));
	jdff dff_B_0qy9Xb9k3_1(.din(w_dff_B_V7mgggxv6_1),.dout(w_dff_B_0qy9Xb9k3_1),.clk(gclk));
	jdff dff_B_hV2arTAE2_1(.din(w_dff_B_0qy9Xb9k3_1),.dout(w_dff_B_hV2arTAE2_1),.clk(gclk));
	jdff dff_B_0gg7424s5_1(.din(w_dff_B_hV2arTAE2_1),.dout(w_dff_B_0gg7424s5_1),.clk(gclk));
	jdff dff_B_cN3qZ7nT9_1(.din(w_dff_B_0gg7424s5_1),.dout(w_dff_B_cN3qZ7nT9_1),.clk(gclk));
	jdff dff_B_QmAHih4Q6_1(.din(w_dff_B_cN3qZ7nT9_1),.dout(w_dff_B_QmAHih4Q6_1),.clk(gclk));
	jdff dff_B_lNAl2PBD8_1(.din(w_dff_B_QmAHih4Q6_1),.dout(w_dff_B_lNAl2PBD8_1),.clk(gclk));
	jdff dff_B_FEOjUxHq4_1(.din(w_dff_B_lNAl2PBD8_1),.dout(w_dff_B_FEOjUxHq4_1),.clk(gclk));
	jdff dff_B_GqgF33Vm5_1(.din(w_dff_B_FEOjUxHq4_1),.dout(w_dff_B_GqgF33Vm5_1),.clk(gclk));
	jdff dff_B_dpeDIHqQ1_1(.din(w_dff_B_GqgF33Vm5_1),.dout(w_dff_B_dpeDIHqQ1_1),.clk(gclk));
	jdff dff_B_3GytPG7M5_1(.din(w_dff_B_dpeDIHqQ1_1),.dout(w_dff_B_3GytPG7M5_1),.clk(gclk));
	jdff dff_B_eYVPShpD2_1(.din(w_dff_B_3GytPG7M5_1),.dout(w_dff_B_eYVPShpD2_1),.clk(gclk));
	jdff dff_B_czpvQJoN5_1(.din(w_dff_B_eYVPShpD2_1),.dout(w_dff_B_czpvQJoN5_1),.clk(gclk));
	jdff dff_B_OwoURhs59_1(.din(w_dff_B_czpvQJoN5_1),.dout(w_dff_B_OwoURhs59_1),.clk(gclk));
	jdff dff_B_BtgBJ39c3_1(.din(w_dff_B_OwoURhs59_1),.dout(w_dff_B_BtgBJ39c3_1),.clk(gclk));
	jdff dff_B_uwsbOTxx4_1(.din(w_dff_B_BtgBJ39c3_1),.dout(w_dff_B_uwsbOTxx4_1),.clk(gclk));
	jdff dff_B_Vnojznox4_1(.din(w_dff_B_uwsbOTxx4_1),.dout(w_dff_B_Vnojznox4_1),.clk(gclk));
	jdff dff_B_ZeRwnd7x6_1(.din(w_dff_B_Vnojznox4_1),.dout(w_dff_B_ZeRwnd7x6_1),.clk(gclk));
	jdff dff_B_dtjxjMSz0_1(.din(w_dff_B_ZeRwnd7x6_1),.dout(w_dff_B_dtjxjMSz0_1),.clk(gclk));
	jdff dff_B_jTDhGBs07_1(.din(w_dff_B_dtjxjMSz0_1),.dout(w_dff_B_jTDhGBs07_1),.clk(gclk));
	jdff dff_B_PTcwSUUh3_1(.din(w_dff_B_jTDhGBs07_1),.dout(w_dff_B_PTcwSUUh3_1),.clk(gclk));
	jdff dff_B_QnUnaBCc7_1(.din(w_dff_B_PTcwSUUh3_1),.dout(w_dff_B_QnUnaBCc7_1),.clk(gclk));
	jdff dff_B_GBGM6Wqj1_1(.din(w_dff_B_QnUnaBCc7_1),.dout(w_dff_B_GBGM6Wqj1_1),.clk(gclk));
	jdff dff_B_ycVE9GKq1_1(.din(w_dff_B_GBGM6Wqj1_1),.dout(w_dff_B_ycVE9GKq1_1),.clk(gclk));
	jdff dff_B_UM3geSuB2_1(.din(w_dff_B_ycVE9GKq1_1),.dout(w_dff_B_UM3geSuB2_1),.clk(gclk));
	jdff dff_B_in75Yttl2_1(.din(w_dff_B_UM3geSuB2_1),.dout(w_dff_B_in75Yttl2_1),.clk(gclk));
	jdff dff_B_sYnq7Z1t6_1(.din(w_dff_B_in75Yttl2_1),.dout(w_dff_B_sYnq7Z1t6_1),.clk(gclk));
	jdff dff_B_G1EGA7eb7_1(.din(w_dff_B_sYnq7Z1t6_1),.dout(w_dff_B_G1EGA7eb7_1),.clk(gclk));
	jdff dff_B_9TEw2b3a3_1(.din(w_dff_B_G1EGA7eb7_1),.dout(w_dff_B_9TEw2b3a3_1),.clk(gclk));
	jdff dff_B_7gPiBWga2_1(.din(w_dff_B_9TEw2b3a3_1),.dout(w_dff_B_7gPiBWga2_1),.clk(gclk));
	jdff dff_B_Y1BbdXkY5_1(.din(w_dff_B_7gPiBWga2_1),.dout(w_dff_B_Y1BbdXkY5_1),.clk(gclk));
	jdff dff_B_o4QB8nIG6_1(.din(w_dff_B_Y1BbdXkY5_1),.dout(w_dff_B_o4QB8nIG6_1),.clk(gclk));
	jdff dff_B_qgluD6W81_0(.din(n709),.dout(w_dff_B_qgluD6W81_0),.clk(gclk));
	jdff dff_B_P3tZvSFY8_0(.din(w_dff_B_qgluD6W81_0),.dout(w_dff_B_P3tZvSFY8_0),.clk(gclk));
	jdff dff_B_cjmn3daQ8_0(.din(w_dff_B_P3tZvSFY8_0),.dout(w_dff_B_cjmn3daQ8_0),.clk(gclk));
	jdff dff_B_lkP51Fe28_0(.din(w_dff_B_cjmn3daQ8_0),.dout(w_dff_B_lkP51Fe28_0),.clk(gclk));
	jdff dff_B_RX372wIP1_0(.din(w_dff_B_lkP51Fe28_0),.dout(w_dff_B_RX372wIP1_0),.clk(gclk));
	jdff dff_B_LODRxVuP3_0(.din(w_dff_B_RX372wIP1_0),.dout(w_dff_B_LODRxVuP3_0),.clk(gclk));
	jdff dff_B_CMvbWlZI9_0(.din(w_dff_B_LODRxVuP3_0),.dout(w_dff_B_CMvbWlZI9_0),.clk(gclk));
	jdff dff_B_Qw4zpn3i3_0(.din(w_dff_B_CMvbWlZI9_0),.dout(w_dff_B_Qw4zpn3i3_0),.clk(gclk));
	jdff dff_B_XSkCxKzz4_0(.din(w_dff_B_Qw4zpn3i3_0),.dout(w_dff_B_XSkCxKzz4_0),.clk(gclk));
	jdff dff_B_kdriNoI87_0(.din(w_dff_B_XSkCxKzz4_0),.dout(w_dff_B_kdriNoI87_0),.clk(gclk));
	jdff dff_B_U6JGT3CN0_0(.din(w_dff_B_kdriNoI87_0),.dout(w_dff_B_U6JGT3CN0_0),.clk(gclk));
	jdff dff_B_AYF1fGEB5_0(.din(w_dff_B_U6JGT3CN0_0),.dout(w_dff_B_AYF1fGEB5_0),.clk(gclk));
	jdff dff_B_NsXxB5lA3_0(.din(w_dff_B_AYF1fGEB5_0),.dout(w_dff_B_NsXxB5lA3_0),.clk(gclk));
	jdff dff_B_5EflqxPj3_0(.din(w_dff_B_NsXxB5lA3_0),.dout(w_dff_B_5EflqxPj3_0),.clk(gclk));
	jdff dff_B_ltqeW4Ki0_0(.din(w_dff_B_5EflqxPj3_0),.dout(w_dff_B_ltqeW4Ki0_0),.clk(gclk));
	jdff dff_B_ktfDYClP5_0(.din(w_dff_B_ltqeW4Ki0_0),.dout(w_dff_B_ktfDYClP5_0),.clk(gclk));
	jdff dff_B_lt1VzINv0_0(.din(w_dff_B_ktfDYClP5_0),.dout(w_dff_B_lt1VzINv0_0),.clk(gclk));
	jdff dff_B_cc3jXEfG1_0(.din(w_dff_B_lt1VzINv0_0),.dout(w_dff_B_cc3jXEfG1_0),.clk(gclk));
	jdff dff_B_bzOPL8I80_0(.din(w_dff_B_cc3jXEfG1_0),.dout(w_dff_B_bzOPL8I80_0),.clk(gclk));
	jdff dff_B_qWehV0hB2_0(.din(w_dff_B_bzOPL8I80_0),.dout(w_dff_B_qWehV0hB2_0),.clk(gclk));
	jdff dff_B_xlDhjvz07_0(.din(w_dff_B_qWehV0hB2_0),.dout(w_dff_B_xlDhjvz07_0),.clk(gclk));
	jdff dff_B_pUaOUwjp9_0(.din(w_dff_B_xlDhjvz07_0),.dout(w_dff_B_pUaOUwjp9_0),.clk(gclk));
	jdff dff_B_UIwajwPo0_0(.din(w_dff_B_pUaOUwjp9_0),.dout(w_dff_B_UIwajwPo0_0),.clk(gclk));
	jdff dff_B_d0BF7Ojp6_0(.din(w_dff_B_UIwajwPo0_0),.dout(w_dff_B_d0BF7Ojp6_0),.clk(gclk));
	jdff dff_B_izH7tfVv4_0(.din(w_dff_B_d0BF7Ojp6_0),.dout(w_dff_B_izH7tfVv4_0),.clk(gclk));
	jdff dff_B_LfQudMwg9_0(.din(w_dff_B_izH7tfVv4_0),.dout(w_dff_B_LfQudMwg9_0),.clk(gclk));
	jdff dff_B_hhFLWRJV0_0(.din(w_dff_B_LfQudMwg9_0),.dout(w_dff_B_hhFLWRJV0_0),.clk(gclk));
	jdff dff_B_OXUtnckG6_0(.din(w_dff_B_hhFLWRJV0_0),.dout(w_dff_B_OXUtnckG6_0),.clk(gclk));
	jdff dff_B_eOyAxgCh7_0(.din(w_dff_B_OXUtnckG6_0),.dout(w_dff_B_eOyAxgCh7_0),.clk(gclk));
	jdff dff_B_XVCZhUN09_0(.din(w_dff_B_eOyAxgCh7_0),.dout(w_dff_B_XVCZhUN09_0),.clk(gclk));
	jdff dff_B_0v9ArSCW1_0(.din(w_dff_B_XVCZhUN09_0),.dout(w_dff_B_0v9ArSCW1_0),.clk(gclk));
	jdff dff_B_Yw3riKHO0_0(.din(w_dff_B_0v9ArSCW1_0),.dout(w_dff_B_Yw3riKHO0_0),.clk(gclk));
	jdff dff_B_OtOLNGDa9_0(.din(w_dff_B_Yw3riKHO0_0),.dout(w_dff_B_OtOLNGDa9_0),.clk(gclk));
	jdff dff_B_yYSI4l345_0(.din(w_dff_B_OtOLNGDa9_0),.dout(w_dff_B_yYSI4l345_0),.clk(gclk));
	jdff dff_B_Ax22BgcJ8_0(.din(w_dff_B_yYSI4l345_0),.dout(w_dff_B_Ax22BgcJ8_0),.clk(gclk));
	jdff dff_B_M1iRof4g1_0(.din(w_dff_B_Ax22BgcJ8_0),.dout(w_dff_B_M1iRof4g1_0),.clk(gclk));
	jdff dff_B_HqLo0pTa7_0(.din(w_dff_B_M1iRof4g1_0),.dout(w_dff_B_HqLo0pTa7_0),.clk(gclk));
	jdff dff_B_ios72luL7_0(.din(w_dff_B_HqLo0pTa7_0),.dout(w_dff_B_ios72luL7_0),.clk(gclk));
	jdff dff_B_S4FK22xX7_0(.din(w_dff_B_ios72luL7_0),.dout(w_dff_B_S4FK22xX7_0),.clk(gclk));
	jdff dff_B_KfRSqJR12_0(.din(w_dff_B_S4FK22xX7_0),.dout(w_dff_B_KfRSqJR12_0),.clk(gclk));
	jdff dff_B_4UyExW7n7_0(.din(w_dff_B_KfRSqJR12_0),.dout(w_dff_B_4UyExW7n7_0),.clk(gclk));
	jdff dff_B_eQU5zz4z1_0(.din(w_dff_B_4UyExW7n7_0),.dout(w_dff_B_eQU5zz4z1_0),.clk(gclk));
	jdff dff_B_4oDxjTBS4_0(.din(w_dff_B_eQU5zz4z1_0),.dout(w_dff_B_4oDxjTBS4_0),.clk(gclk));
	jdff dff_B_Xo416V730_0(.din(w_dff_B_4oDxjTBS4_0),.dout(w_dff_B_Xo416V730_0),.clk(gclk));
	jdff dff_B_Vqvyy7Tn2_0(.din(w_dff_B_Xo416V730_0),.dout(w_dff_B_Vqvyy7Tn2_0),.clk(gclk));
	jdff dff_B_4xJChCV04_0(.din(w_dff_B_Vqvyy7Tn2_0),.dout(w_dff_B_4xJChCV04_0),.clk(gclk));
	jdff dff_B_Oi3s39gH7_0(.din(w_dff_B_4xJChCV04_0),.dout(w_dff_B_Oi3s39gH7_0),.clk(gclk));
	jdff dff_B_pIXfFVxd7_0(.din(w_dff_B_Oi3s39gH7_0),.dout(w_dff_B_pIXfFVxd7_0),.clk(gclk));
	jdff dff_B_ie4FZ6xV3_0(.din(w_dff_B_pIXfFVxd7_0),.dout(w_dff_B_ie4FZ6xV3_0),.clk(gclk));
	jdff dff_B_LJi9gYe52_0(.din(w_dff_B_ie4FZ6xV3_0),.dout(w_dff_B_LJi9gYe52_0),.clk(gclk));
	jdff dff_B_UPmU200N5_0(.din(w_dff_B_LJi9gYe52_0),.dout(w_dff_B_UPmU200N5_0),.clk(gclk));
	jdff dff_B_5KI7Y7LT5_0(.din(w_dff_B_UPmU200N5_0),.dout(w_dff_B_5KI7Y7LT5_0),.clk(gclk));
	jdff dff_B_f3oqTQmX3_0(.din(w_dff_B_5KI7Y7LT5_0),.dout(w_dff_B_f3oqTQmX3_0),.clk(gclk));
	jdff dff_B_PGiiN9Zt6_0(.din(w_dff_B_f3oqTQmX3_0),.dout(w_dff_B_PGiiN9Zt6_0),.clk(gclk));
	jdff dff_B_3NitMkSn5_1(.din(n702),.dout(w_dff_B_3NitMkSn5_1),.clk(gclk));
	jdff dff_B_TD2Z713j1_1(.din(w_dff_B_3NitMkSn5_1),.dout(w_dff_B_TD2Z713j1_1),.clk(gclk));
	jdff dff_B_fP6arkUA1_1(.din(w_dff_B_TD2Z713j1_1),.dout(w_dff_B_fP6arkUA1_1),.clk(gclk));
	jdff dff_B_5hibjoB12_1(.din(w_dff_B_fP6arkUA1_1),.dout(w_dff_B_5hibjoB12_1),.clk(gclk));
	jdff dff_B_SBj1vHub8_1(.din(w_dff_B_5hibjoB12_1),.dout(w_dff_B_SBj1vHub8_1),.clk(gclk));
	jdff dff_B_zbKmpZxD4_1(.din(w_dff_B_SBj1vHub8_1),.dout(w_dff_B_zbKmpZxD4_1),.clk(gclk));
	jdff dff_B_lqY1FCXF4_1(.din(w_dff_B_zbKmpZxD4_1),.dout(w_dff_B_lqY1FCXF4_1),.clk(gclk));
	jdff dff_B_dM9s1a8J8_1(.din(w_dff_B_lqY1FCXF4_1),.dout(w_dff_B_dM9s1a8J8_1),.clk(gclk));
	jdff dff_B_LM3SgKNk9_1(.din(w_dff_B_dM9s1a8J8_1),.dout(w_dff_B_LM3SgKNk9_1),.clk(gclk));
	jdff dff_B_SDopu2EN1_1(.din(w_dff_B_LM3SgKNk9_1),.dout(w_dff_B_SDopu2EN1_1),.clk(gclk));
	jdff dff_B_N4MNZalv6_1(.din(w_dff_B_SDopu2EN1_1),.dout(w_dff_B_N4MNZalv6_1),.clk(gclk));
	jdff dff_B_YiirUJhj9_1(.din(w_dff_B_N4MNZalv6_1),.dout(w_dff_B_YiirUJhj9_1),.clk(gclk));
	jdff dff_B_OwSdZTxt6_1(.din(w_dff_B_YiirUJhj9_1),.dout(w_dff_B_OwSdZTxt6_1),.clk(gclk));
	jdff dff_B_2VqZHS2R7_1(.din(w_dff_B_OwSdZTxt6_1),.dout(w_dff_B_2VqZHS2R7_1),.clk(gclk));
	jdff dff_B_XHsRDCG96_1(.din(w_dff_B_2VqZHS2R7_1),.dout(w_dff_B_XHsRDCG96_1),.clk(gclk));
	jdff dff_B_6q7Z3Cw30_1(.din(w_dff_B_XHsRDCG96_1),.dout(w_dff_B_6q7Z3Cw30_1),.clk(gclk));
	jdff dff_B_EkEgcoTD9_1(.din(w_dff_B_6q7Z3Cw30_1),.dout(w_dff_B_EkEgcoTD9_1),.clk(gclk));
	jdff dff_B_hXtkLu3D3_1(.din(w_dff_B_EkEgcoTD9_1),.dout(w_dff_B_hXtkLu3D3_1),.clk(gclk));
	jdff dff_B_ZcVTmXbd9_1(.din(w_dff_B_hXtkLu3D3_1),.dout(w_dff_B_ZcVTmXbd9_1),.clk(gclk));
	jdff dff_B_A1XMNnPh8_1(.din(w_dff_B_ZcVTmXbd9_1),.dout(w_dff_B_A1XMNnPh8_1),.clk(gclk));
	jdff dff_B_WI4lMTSO2_1(.din(w_dff_B_A1XMNnPh8_1),.dout(w_dff_B_WI4lMTSO2_1),.clk(gclk));
	jdff dff_B_tREcRG0L5_1(.din(w_dff_B_WI4lMTSO2_1),.dout(w_dff_B_tREcRG0L5_1),.clk(gclk));
	jdff dff_B_U0HNQjfI9_1(.din(w_dff_B_tREcRG0L5_1),.dout(w_dff_B_U0HNQjfI9_1),.clk(gclk));
	jdff dff_B_mG0IVshm0_1(.din(w_dff_B_U0HNQjfI9_1),.dout(w_dff_B_mG0IVshm0_1),.clk(gclk));
	jdff dff_B_t6azt6QS3_1(.din(w_dff_B_mG0IVshm0_1),.dout(w_dff_B_t6azt6QS3_1),.clk(gclk));
	jdff dff_B_dRas7cl43_1(.din(w_dff_B_t6azt6QS3_1),.dout(w_dff_B_dRas7cl43_1),.clk(gclk));
	jdff dff_B_J8Lii8eP9_1(.din(w_dff_B_dRas7cl43_1),.dout(w_dff_B_J8Lii8eP9_1),.clk(gclk));
	jdff dff_B_Lvmat3IV1_1(.din(w_dff_B_J8Lii8eP9_1),.dout(w_dff_B_Lvmat3IV1_1),.clk(gclk));
	jdff dff_B_cIoF13n37_1(.din(w_dff_B_Lvmat3IV1_1),.dout(w_dff_B_cIoF13n37_1),.clk(gclk));
	jdff dff_B_WXyncf266_1(.din(w_dff_B_cIoF13n37_1),.dout(w_dff_B_WXyncf266_1),.clk(gclk));
	jdff dff_B_SbnysYY39_1(.din(w_dff_B_WXyncf266_1),.dout(w_dff_B_SbnysYY39_1),.clk(gclk));
	jdff dff_B_mB3fUMUv3_1(.din(w_dff_B_SbnysYY39_1),.dout(w_dff_B_mB3fUMUv3_1),.clk(gclk));
	jdff dff_B_NFX3FAcm5_1(.din(w_dff_B_mB3fUMUv3_1),.dout(w_dff_B_NFX3FAcm5_1),.clk(gclk));
	jdff dff_B_34KXOmbo1_1(.din(w_dff_B_NFX3FAcm5_1),.dout(w_dff_B_34KXOmbo1_1),.clk(gclk));
	jdff dff_B_gntJ5zFW8_1(.din(w_dff_B_34KXOmbo1_1),.dout(w_dff_B_gntJ5zFW8_1),.clk(gclk));
	jdff dff_B_Fd5aVKKW5_1(.din(w_dff_B_gntJ5zFW8_1),.dout(w_dff_B_Fd5aVKKW5_1),.clk(gclk));
	jdff dff_B_V1Fzn0Hz3_1(.din(w_dff_B_Fd5aVKKW5_1),.dout(w_dff_B_V1Fzn0Hz3_1),.clk(gclk));
	jdff dff_B_SHzVeHZz1_1(.din(w_dff_B_V1Fzn0Hz3_1),.dout(w_dff_B_SHzVeHZz1_1),.clk(gclk));
	jdff dff_B_ABl7DXHU3_1(.din(w_dff_B_SHzVeHZz1_1),.dout(w_dff_B_ABl7DXHU3_1),.clk(gclk));
	jdff dff_B_Oa0XLna62_1(.din(w_dff_B_ABl7DXHU3_1),.dout(w_dff_B_Oa0XLna62_1),.clk(gclk));
	jdff dff_B_NSKaInd08_1(.din(w_dff_B_Oa0XLna62_1),.dout(w_dff_B_NSKaInd08_1),.clk(gclk));
	jdff dff_B_jrGGJek59_1(.din(w_dff_B_NSKaInd08_1),.dout(w_dff_B_jrGGJek59_1),.clk(gclk));
	jdff dff_B_mD9wOaOj6_1(.din(w_dff_B_jrGGJek59_1),.dout(w_dff_B_mD9wOaOj6_1),.clk(gclk));
	jdff dff_B_XdEyA1PA6_1(.din(w_dff_B_mD9wOaOj6_1),.dout(w_dff_B_XdEyA1PA6_1),.clk(gclk));
	jdff dff_B_GUKttWlt3_1(.din(w_dff_B_XdEyA1PA6_1),.dout(w_dff_B_GUKttWlt3_1),.clk(gclk));
	jdff dff_B_7TkwSu6j1_1(.din(w_dff_B_GUKttWlt3_1),.dout(w_dff_B_7TkwSu6j1_1),.clk(gclk));
	jdff dff_B_MC81BYoT1_1(.din(w_dff_B_7TkwSu6j1_1),.dout(w_dff_B_MC81BYoT1_1),.clk(gclk));
	jdff dff_B_pOxdbK7F9_1(.din(w_dff_B_MC81BYoT1_1),.dout(w_dff_B_pOxdbK7F9_1),.clk(gclk));
	jdff dff_B_SGlrsFHN7_1(.din(w_dff_B_pOxdbK7F9_1),.dout(w_dff_B_SGlrsFHN7_1),.clk(gclk));
	jdff dff_B_BwevHhOt9_1(.din(w_dff_B_SGlrsFHN7_1),.dout(w_dff_B_BwevHhOt9_1),.clk(gclk));
	jdff dff_B_aeNYWdBC5_1(.din(w_dff_B_BwevHhOt9_1),.dout(w_dff_B_aeNYWdBC5_1),.clk(gclk));
	jdff dff_B_ASGowOXa9_1(.din(w_dff_B_aeNYWdBC5_1),.dout(w_dff_B_ASGowOXa9_1),.clk(gclk));
	jdff dff_B_NmBOBsht4_1(.din(w_dff_B_ASGowOXa9_1),.dout(w_dff_B_NmBOBsht4_1),.clk(gclk));
	jdff dff_B_LZiz5Mk84_0(.din(n703),.dout(w_dff_B_LZiz5Mk84_0),.clk(gclk));
	jdff dff_B_Cg7oUIvo6_0(.din(w_dff_B_LZiz5Mk84_0),.dout(w_dff_B_Cg7oUIvo6_0),.clk(gclk));
	jdff dff_B_qmpjg2xX3_0(.din(w_dff_B_Cg7oUIvo6_0),.dout(w_dff_B_qmpjg2xX3_0),.clk(gclk));
	jdff dff_B_8MeaT4Re8_0(.din(w_dff_B_qmpjg2xX3_0),.dout(w_dff_B_8MeaT4Re8_0),.clk(gclk));
	jdff dff_B_rU1WovaH5_0(.din(w_dff_B_8MeaT4Re8_0),.dout(w_dff_B_rU1WovaH5_0),.clk(gclk));
	jdff dff_B_cCDqW4AS3_0(.din(w_dff_B_rU1WovaH5_0),.dout(w_dff_B_cCDqW4AS3_0),.clk(gclk));
	jdff dff_B_bSODKpen8_0(.din(w_dff_B_cCDqW4AS3_0),.dout(w_dff_B_bSODKpen8_0),.clk(gclk));
	jdff dff_B_59KfPeM54_0(.din(w_dff_B_bSODKpen8_0),.dout(w_dff_B_59KfPeM54_0),.clk(gclk));
	jdff dff_B_CQIrmEjv0_0(.din(w_dff_B_59KfPeM54_0),.dout(w_dff_B_CQIrmEjv0_0),.clk(gclk));
	jdff dff_B_M5z9CxST4_0(.din(w_dff_B_CQIrmEjv0_0),.dout(w_dff_B_M5z9CxST4_0),.clk(gclk));
	jdff dff_B_uOUHpAvM3_0(.din(w_dff_B_M5z9CxST4_0),.dout(w_dff_B_uOUHpAvM3_0),.clk(gclk));
	jdff dff_B_tFlWG7Wd3_0(.din(w_dff_B_uOUHpAvM3_0),.dout(w_dff_B_tFlWG7Wd3_0),.clk(gclk));
	jdff dff_B_s4OlzC849_0(.din(w_dff_B_tFlWG7Wd3_0),.dout(w_dff_B_s4OlzC849_0),.clk(gclk));
	jdff dff_B_jogyRlTu0_0(.din(w_dff_B_s4OlzC849_0),.dout(w_dff_B_jogyRlTu0_0),.clk(gclk));
	jdff dff_B_8KxzbwZY6_0(.din(w_dff_B_jogyRlTu0_0),.dout(w_dff_B_8KxzbwZY6_0),.clk(gclk));
	jdff dff_B_KZvx0bmv9_0(.din(w_dff_B_8KxzbwZY6_0),.dout(w_dff_B_KZvx0bmv9_0),.clk(gclk));
	jdff dff_B_ENkhQy1m6_0(.din(w_dff_B_KZvx0bmv9_0),.dout(w_dff_B_ENkhQy1m6_0),.clk(gclk));
	jdff dff_B_Q8vIP5FK5_0(.din(w_dff_B_ENkhQy1m6_0),.dout(w_dff_B_Q8vIP5FK5_0),.clk(gclk));
	jdff dff_B_wvrTyQXF7_0(.din(w_dff_B_Q8vIP5FK5_0),.dout(w_dff_B_wvrTyQXF7_0),.clk(gclk));
	jdff dff_B_qIg12tJV1_0(.din(w_dff_B_wvrTyQXF7_0),.dout(w_dff_B_qIg12tJV1_0),.clk(gclk));
	jdff dff_B_4R10EknX2_0(.din(w_dff_B_qIg12tJV1_0),.dout(w_dff_B_4R10EknX2_0),.clk(gclk));
	jdff dff_B_x6m6PfM41_0(.din(w_dff_B_4R10EknX2_0),.dout(w_dff_B_x6m6PfM41_0),.clk(gclk));
	jdff dff_B_IuGJVSDc4_0(.din(w_dff_B_x6m6PfM41_0),.dout(w_dff_B_IuGJVSDc4_0),.clk(gclk));
	jdff dff_B_EaB2OiFS9_0(.din(w_dff_B_IuGJVSDc4_0),.dout(w_dff_B_EaB2OiFS9_0),.clk(gclk));
	jdff dff_B_7tLK8jSy8_0(.din(w_dff_B_EaB2OiFS9_0),.dout(w_dff_B_7tLK8jSy8_0),.clk(gclk));
	jdff dff_B_abJ5S8bA8_0(.din(w_dff_B_7tLK8jSy8_0),.dout(w_dff_B_abJ5S8bA8_0),.clk(gclk));
	jdff dff_B_wyHXDwFz2_0(.din(w_dff_B_abJ5S8bA8_0),.dout(w_dff_B_wyHXDwFz2_0),.clk(gclk));
	jdff dff_B_nqfoKhld4_0(.din(w_dff_B_wyHXDwFz2_0),.dout(w_dff_B_nqfoKhld4_0),.clk(gclk));
	jdff dff_B_UeIP226U6_0(.din(w_dff_B_nqfoKhld4_0),.dout(w_dff_B_UeIP226U6_0),.clk(gclk));
	jdff dff_B_hMQyWIQ96_0(.din(w_dff_B_UeIP226U6_0),.dout(w_dff_B_hMQyWIQ96_0),.clk(gclk));
	jdff dff_B_rY8jcPou3_0(.din(w_dff_B_hMQyWIQ96_0),.dout(w_dff_B_rY8jcPou3_0),.clk(gclk));
	jdff dff_B_77ox5Eyr9_0(.din(w_dff_B_rY8jcPou3_0),.dout(w_dff_B_77ox5Eyr9_0),.clk(gclk));
	jdff dff_B_ARztImsF2_0(.din(w_dff_B_77ox5Eyr9_0),.dout(w_dff_B_ARztImsF2_0),.clk(gclk));
	jdff dff_B_9Ieo69JZ3_0(.din(w_dff_B_ARztImsF2_0),.dout(w_dff_B_9Ieo69JZ3_0),.clk(gclk));
	jdff dff_B_yaH6cuNL9_0(.din(w_dff_B_9Ieo69JZ3_0),.dout(w_dff_B_yaH6cuNL9_0),.clk(gclk));
	jdff dff_B_P9wUUOL93_0(.din(w_dff_B_yaH6cuNL9_0),.dout(w_dff_B_P9wUUOL93_0),.clk(gclk));
	jdff dff_B_cDXCglxj5_0(.din(w_dff_B_P9wUUOL93_0),.dout(w_dff_B_cDXCglxj5_0),.clk(gclk));
	jdff dff_B_OiBhCLLK5_0(.din(w_dff_B_cDXCglxj5_0),.dout(w_dff_B_OiBhCLLK5_0),.clk(gclk));
	jdff dff_B_PmXYMJ4Q5_0(.din(w_dff_B_OiBhCLLK5_0),.dout(w_dff_B_PmXYMJ4Q5_0),.clk(gclk));
	jdff dff_B_J8TpZcJc0_0(.din(w_dff_B_PmXYMJ4Q5_0),.dout(w_dff_B_J8TpZcJc0_0),.clk(gclk));
	jdff dff_B_cA507CoC5_0(.din(w_dff_B_J8TpZcJc0_0),.dout(w_dff_B_cA507CoC5_0),.clk(gclk));
	jdff dff_B_XjlxePQq2_0(.din(w_dff_B_cA507CoC5_0),.dout(w_dff_B_XjlxePQq2_0),.clk(gclk));
	jdff dff_B_KdPouap28_0(.din(w_dff_B_XjlxePQq2_0),.dout(w_dff_B_KdPouap28_0),.clk(gclk));
	jdff dff_B_caKrQ1o24_0(.din(w_dff_B_KdPouap28_0),.dout(w_dff_B_caKrQ1o24_0),.clk(gclk));
	jdff dff_B_fiSm5DT83_0(.din(w_dff_B_caKrQ1o24_0),.dout(w_dff_B_fiSm5DT83_0),.clk(gclk));
	jdff dff_B_uocp1eZa9_0(.din(w_dff_B_fiSm5DT83_0),.dout(w_dff_B_uocp1eZa9_0),.clk(gclk));
	jdff dff_B_tlaMApI32_0(.din(w_dff_B_uocp1eZa9_0),.dout(w_dff_B_tlaMApI32_0),.clk(gclk));
	jdff dff_B_yFCLzRZ81_0(.din(w_dff_B_tlaMApI32_0),.dout(w_dff_B_yFCLzRZ81_0),.clk(gclk));
	jdff dff_B_hNPlTbA14_0(.din(w_dff_B_yFCLzRZ81_0),.dout(w_dff_B_hNPlTbA14_0),.clk(gclk));
	jdff dff_B_fy7XqznP4_0(.din(w_dff_B_hNPlTbA14_0),.dout(w_dff_B_fy7XqznP4_0),.clk(gclk));
	jdff dff_B_OOSx4D8S7_0(.din(w_dff_B_fy7XqznP4_0),.dout(w_dff_B_OOSx4D8S7_0),.clk(gclk));
	jdff dff_B_YAYWLjIP7_0(.din(w_dff_B_OOSx4D8S7_0),.dout(w_dff_B_YAYWLjIP7_0),.clk(gclk));
	jdff dff_B_PKOhVjuX2_0(.din(w_dff_B_YAYWLjIP7_0),.dout(w_dff_B_PKOhVjuX2_0),.clk(gclk));
	jdff dff_B_UaRV9XiG9_1(.din(n696),.dout(w_dff_B_UaRV9XiG9_1),.clk(gclk));
	jdff dff_B_ai6QQYtD2_1(.din(w_dff_B_UaRV9XiG9_1),.dout(w_dff_B_ai6QQYtD2_1),.clk(gclk));
	jdff dff_B_6ulGzJuO0_1(.din(w_dff_B_ai6QQYtD2_1),.dout(w_dff_B_6ulGzJuO0_1),.clk(gclk));
	jdff dff_B_Yh8x01by5_1(.din(w_dff_B_6ulGzJuO0_1),.dout(w_dff_B_Yh8x01by5_1),.clk(gclk));
	jdff dff_B_cZz7PcrI2_1(.din(w_dff_B_Yh8x01by5_1),.dout(w_dff_B_cZz7PcrI2_1),.clk(gclk));
	jdff dff_B_HXraKzYR1_1(.din(w_dff_B_cZz7PcrI2_1),.dout(w_dff_B_HXraKzYR1_1),.clk(gclk));
	jdff dff_B_hDoW6Imj0_1(.din(w_dff_B_HXraKzYR1_1),.dout(w_dff_B_hDoW6Imj0_1),.clk(gclk));
	jdff dff_B_9BhmjCQ98_1(.din(w_dff_B_hDoW6Imj0_1),.dout(w_dff_B_9BhmjCQ98_1),.clk(gclk));
	jdff dff_B_z1A0BqMQ0_1(.din(w_dff_B_9BhmjCQ98_1),.dout(w_dff_B_z1A0BqMQ0_1),.clk(gclk));
	jdff dff_B_cQw5Ygzh8_1(.din(w_dff_B_z1A0BqMQ0_1),.dout(w_dff_B_cQw5Ygzh8_1),.clk(gclk));
	jdff dff_B_geHnPb5o1_1(.din(w_dff_B_cQw5Ygzh8_1),.dout(w_dff_B_geHnPb5o1_1),.clk(gclk));
	jdff dff_B_rL0o6L9n1_1(.din(w_dff_B_geHnPb5o1_1),.dout(w_dff_B_rL0o6L9n1_1),.clk(gclk));
	jdff dff_B_fGXVZiE07_1(.din(w_dff_B_rL0o6L9n1_1),.dout(w_dff_B_fGXVZiE07_1),.clk(gclk));
	jdff dff_B_r5eIxA1C1_1(.din(w_dff_B_fGXVZiE07_1),.dout(w_dff_B_r5eIxA1C1_1),.clk(gclk));
	jdff dff_B_5Zr7A37h7_1(.din(w_dff_B_r5eIxA1C1_1),.dout(w_dff_B_5Zr7A37h7_1),.clk(gclk));
	jdff dff_B_8YGySTQb1_1(.din(w_dff_B_5Zr7A37h7_1),.dout(w_dff_B_8YGySTQb1_1),.clk(gclk));
	jdff dff_B_qkQiWXg85_1(.din(w_dff_B_8YGySTQb1_1),.dout(w_dff_B_qkQiWXg85_1),.clk(gclk));
	jdff dff_B_Lnf1Vxmy8_1(.din(w_dff_B_qkQiWXg85_1),.dout(w_dff_B_Lnf1Vxmy8_1),.clk(gclk));
	jdff dff_B_gNg2Bj4n7_1(.din(w_dff_B_Lnf1Vxmy8_1),.dout(w_dff_B_gNg2Bj4n7_1),.clk(gclk));
	jdff dff_B_F5BkbjlA0_1(.din(w_dff_B_gNg2Bj4n7_1),.dout(w_dff_B_F5BkbjlA0_1),.clk(gclk));
	jdff dff_B_nSSjuBxj0_1(.din(w_dff_B_F5BkbjlA0_1),.dout(w_dff_B_nSSjuBxj0_1),.clk(gclk));
	jdff dff_B_jRNSO7Ad9_1(.din(w_dff_B_nSSjuBxj0_1),.dout(w_dff_B_jRNSO7Ad9_1),.clk(gclk));
	jdff dff_B_CfZtREaj7_1(.din(w_dff_B_jRNSO7Ad9_1),.dout(w_dff_B_CfZtREaj7_1),.clk(gclk));
	jdff dff_B_pcNBA27f6_1(.din(w_dff_B_CfZtREaj7_1),.dout(w_dff_B_pcNBA27f6_1),.clk(gclk));
	jdff dff_B_YjQIUFxD7_1(.din(w_dff_B_pcNBA27f6_1),.dout(w_dff_B_YjQIUFxD7_1),.clk(gclk));
	jdff dff_B_elgCwbZ71_1(.din(w_dff_B_YjQIUFxD7_1),.dout(w_dff_B_elgCwbZ71_1),.clk(gclk));
	jdff dff_B_nOIukjqm0_1(.din(w_dff_B_elgCwbZ71_1),.dout(w_dff_B_nOIukjqm0_1),.clk(gclk));
	jdff dff_B_vSQHOlay9_1(.din(w_dff_B_nOIukjqm0_1),.dout(w_dff_B_vSQHOlay9_1),.clk(gclk));
	jdff dff_B_HagQRFEJ2_1(.din(w_dff_B_vSQHOlay9_1),.dout(w_dff_B_HagQRFEJ2_1),.clk(gclk));
	jdff dff_B_moWyMS6c6_1(.din(w_dff_B_HagQRFEJ2_1),.dout(w_dff_B_moWyMS6c6_1),.clk(gclk));
	jdff dff_B_FgbhDgid5_1(.din(w_dff_B_moWyMS6c6_1),.dout(w_dff_B_FgbhDgid5_1),.clk(gclk));
	jdff dff_B_YnndI7fC7_1(.din(w_dff_B_FgbhDgid5_1),.dout(w_dff_B_YnndI7fC7_1),.clk(gclk));
	jdff dff_B_8AjHEswg3_1(.din(w_dff_B_YnndI7fC7_1),.dout(w_dff_B_8AjHEswg3_1),.clk(gclk));
	jdff dff_B_omF8WcBY1_1(.din(w_dff_B_8AjHEswg3_1),.dout(w_dff_B_omF8WcBY1_1),.clk(gclk));
	jdff dff_B_4cQ0tuWt0_1(.din(w_dff_B_omF8WcBY1_1),.dout(w_dff_B_4cQ0tuWt0_1),.clk(gclk));
	jdff dff_B_y9xgnwPd1_1(.din(w_dff_B_4cQ0tuWt0_1),.dout(w_dff_B_y9xgnwPd1_1),.clk(gclk));
	jdff dff_B_Ssa1m4iN3_1(.din(w_dff_B_y9xgnwPd1_1),.dout(w_dff_B_Ssa1m4iN3_1),.clk(gclk));
	jdff dff_B_JRrVcOLQ0_1(.din(w_dff_B_Ssa1m4iN3_1),.dout(w_dff_B_JRrVcOLQ0_1),.clk(gclk));
	jdff dff_B_ym9V9iZV0_1(.din(w_dff_B_JRrVcOLQ0_1),.dout(w_dff_B_ym9V9iZV0_1),.clk(gclk));
	jdff dff_B_vQyt8eDB7_1(.din(w_dff_B_ym9V9iZV0_1),.dout(w_dff_B_vQyt8eDB7_1),.clk(gclk));
	jdff dff_B_CWijj2xq6_1(.din(w_dff_B_vQyt8eDB7_1),.dout(w_dff_B_CWijj2xq6_1),.clk(gclk));
	jdff dff_B_sYfMa7sh8_1(.din(w_dff_B_CWijj2xq6_1),.dout(w_dff_B_sYfMa7sh8_1),.clk(gclk));
	jdff dff_B_zYeuVKsX5_1(.din(w_dff_B_sYfMa7sh8_1),.dout(w_dff_B_zYeuVKsX5_1),.clk(gclk));
	jdff dff_B_0qKHwpwa0_1(.din(w_dff_B_zYeuVKsX5_1),.dout(w_dff_B_0qKHwpwa0_1),.clk(gclk));
	jdff dff_B_LrrV8GhS1_1(.din(w_dff_B_0qKHwpwa0_1),.dout(w_dff_B_LrrV8GhS1_1),.clk(gclk));
	jdff dff_B_YxQft1Qn7_1(.din(w_dff_B_LrrV8GhS1_1),.dout(w_dff_B_YxQft1Qn7_1),.clk(gclk));
	jdff dff_B_GUSPqldz7_1(.din(w_dff_B_YxQft1Qn7_1),.dout(w_dff_B_GUSPqldz7_1),.clk(gclk));
	jdff dff_B_tHHP3yKU1_1(.din(w_dff_B_GUSPqldz7_1),.dout(w_dff_B_tHHP3yKU1_1),.clk(gclk));
	jdff dff_B_hlgryvHg4_1(.din(w_dff_B_tHHP3yKU1_1),.dout(w_dff_B_hlgryvHg4_1),.clk(gclk));
	jdff dff_B_4o7gxzqN8_1(.din(w_dff_B_hlgryvHg4_1),.dout(w_dff_B_4o7gxzqN8_1),.clk(gclk));
	jdff dff_B_cluyeuU07_1(.din(w_dff_B_4o7gxzqN8_1),.dout(w_dff_B_cluyeuU07_1),.clk(gclk));
	jdff dff_B_79nILaoK7_1(.din(w_dff_B_cluyeuU07_1),.dout(w_dff_B_79nILaoK7_1),.clk(gclk));
	jdff dff_B_pGUbVjsV3_0(.din(n697),.dout(w_dff_B_pGUbVjsV3_0),.clk(gclk));
	jdff dff_B_d3rqFy5D5_0(.din(w_dff_B_pGUbVjsV3_0),.dout(w_dff_B_d3rqFy5D5_0),.clk(gclk));
	jdff dff_B_BNdNpxkY9_0(.din(w_dff_B_d3rqFy5D5_0),.dout(w_dff_B_BNdNpxkY9_0),.clk(gclk));
	jdff dff_B_Jeo6SBNY1_0(.din(w_dff_B_BNdNpxkY9_0),.dout(w_dff_B_Jeo6SBNY1_0),.clk(gclk));
	jdff dff_B_kOYnA20F5_0(.din(w_dff_B_Jeo6SBNY1_0),.dout(w_dff_B_kOYnA20F5_0),.clk(gclk));
	jdff dff_B_rGvnW9783_0(.din(w_dff_B_kOYnA20F5_0),.dout(w_dff_B_rGvnW9783_0),.clk(gclk));
	jdff dff_B_kOfgVrCm8_0(.din(w_dff_B_rGvnW9783_0),.dout(w_dff_B_kOfgVrCm8_0),.clk(gclk));
	jdff dff_B_4vEHYa0W6_0(.din(w_dff_B_kOfgVrCm8_0),.dout(w_dff_B_4vEHYa0W6_0),.clk(gclk));
	jdff dff_B_1OLEl31J2_0(.din(w_dff_B_4vEHYa0W6_0),.dout(w_dff_B_1OLEl31J2_0),.clk(gclk));
	jdff dff_B_bnqNQYyD9_0(.din(w_dff_B_1OLEl31J2_0),.dout(w_dff_B_bnqNQYyD9_0),.clk(gclk));
	jdff dff_B_yI2g0aOB6_0(.din(w_dff_B_bnqNQYyD9_0),.dout(w_dff_B_yI2g0aOB6_0),.clk(gclk));
	jdff dff_B_8q1AVIyY0_0(.din(w_dff_B_yI2g0aOB6_0),.dout(w_dff_B_8q1AVIyY0_0),.clk(gclk));
	jdff dff_B_9uoMbIDX1_0(.din(w_dff_B_8q1AVIyY0_0),.dout(w_dff_B_9uoMbIDX1_0),.clk(gclk));
	jdff dff_B_90ENeEdu6_0(.din(w_dff_B_9uoMbIDX1_0),.dout(w_dff_B_90ENeEdu6_0),.clk(gclk));
	jdff dff_B_wTcAe09v7_0(.din(w_dff_B_90ENeEdu6_0),.dout(w_dff_B_wTcAe09v7_0),.clk(gclk));
	jdff dff_B_PxMenEEx5_0(.din(w_dff_B_wTcAe09v7_0),.dout(w_dff_B_PxMenEEx5_0),.clk(gclk));
	jdff dff_B_KAVa2u9w1_0(.din(w_dff_B_PxMenEEx5_0),.dout(w_dff_B_KAVa2u9w1_0),.clk(gclk));
	jdff dff_B_NZpfTpyH8_0(.din(w_dff_B_KAVa2u9w1_0),.dout(w_dff_B_NZpfTpyH8_0),.clk(gclk));
	jdff dff_B_1e1mwxTc2_0(.din(w_dff_B_NZpfTpyH8_0),.dout(w_dff_B_1e1mwxTc2_0),.clk(gclk));
	jdff dff_B_LBSYbJPY9_0(.din(w_dff_B_1e1mwxTc2_0),.dout(w_dff_B_LBSYbJPY9_0),.clk(gclk));
	jdff dff_B_FL3l4UmT4_0(.din(w_dff_B_LBSYbJPY9_0),.dout(w_dff_B_FL3l4UmT4_0),.clk(gclk));
	jdff dff_B_egqqIj7F9_0(.din(w_dff_B_FL3l4UmT4_0),.dout(w_dff_B_egqqIj7F9_0),.clk(gclk));
	jdff dff_B_uGfySTqf5_0(.din(w_dff_B_egqqIj7F9_0),.dout(w_dff_B_uGfySTqf5_0),.clk(gclk));
	jdff dff_B_FBFGkjD36_0(.din(w_dff_B_uGfySTqf5_0),.dout(w_dff_B_FBFGkjD36_0),.clk(gclk));
	jdff dff_B_9bywbQDE0_0(.din(w_dff_B_FBFGkjD36_0),.dout(w_dff_B_9bywbQDE0_0),.clk(gclk));
	jdff dff_B_p0RUlMGR9_0(.din(w_dff_B_9bywbQDE0_0),.dout(w_dff_B_p0RUlMGR9_0),.clk(gclk));
	jdff dff_B_NvXMLp5e8_0(.din(w_dff_B_p0RUlMGR9_0),.dout(w_dff_B_NvXMLp5e8_0),.clk(gclk));
	jdff dff_B_cIy6U2Dg3_0(.din(w_dff_B_NvXMLp5e8_0),.dout(w_dff_B_cIy6U2Dg3_0),.clk(gclk));
	jdff dff_B_RpSPZDMK5_0(.din(w_dff_B_cIy6U2Dg3_0),.dout(w_dff_B_RpSPZDMK5_0),.clk(gclk));
	jdff dff_B_cpjiHNqP9_0(.din(w_dff_B_RpSPZDMK5_0),.dout(w_dff_B_cpjiHNqP9_0),.clk(gclk));
	jdff dff_B_bo1EpKJ08_0(.din(w_dff_B_cpjiHNqP9_0),.dout(w_dff_B_bo1EpKJ08_0),.clk(gclk));
	jdff dff_B_0Jjtd9Ny6_0(.din(w_dff_B_bo1EpKJ08_0),.dout(w_dff_B_0Jjtd9Ny6_0),.clk(gclk));
	jdff dff_B_NRRVuZBu9_0(.din(w_dff_B_0Jjtd9Ny6_0),.dout(w_dff_B_NRRVuZBu9_0),.clk(gclk));
	jdff dff_B_9inLRKhL5_0(.din(w_dff_B_NRRVuZBu9_0),.dout(w_dff_B_9inLRKhL5_0),.clk(gclk));
	jdff dff_B_10rHqYex3_0(.din(w_dff_B_9inLRKhL5_0),.dout(w_dff_B_10rHqYex3_0),.clk(gclk));
	jdff dff_B_oQ31CafH6_0(.din(w_dff_B_10rHqYex3_0),.dout(w_dff_B_oQ31CafH6_0),.clk(gclk));
	jdff dff_B_psv2ZGRp5_0(.din(w_dff_B_oQ31CafH6_0),.dout(w_dff_B_psv2ZGRp5_0),.clk(gclk));
	jdff dff_B_S5DVYHzT2_0(.din(w_dff_B_psv2ZGRp5_0),.dout(w_dff_B_S5DVYHzT2_0),.clk(gclk));
	jdff dff_B_nHiGZgZ04_0(.din(w_dff_B_S5DVYHzT2_0),.dout(w_dff_B_nHiGZgZ04_0),.clk(gclk));
	jdff dff_B_XF69njg37_0(.din(w_dff_B_nHiGZgZ04_0),.dout(w_dff_B_XF69njg37_0),.clk(gclk));
	jdff dff_B_vnNfoRqy5_0(.din(w_dff_B_XF69njg37_0),.dout(w_dff_B_vnNfoRqy5_0),.clk(gclk));
	jdff dff_B_6job68c48_0(.din(w_dff_B_vnNfoRqy5_0),.dout(w_dff_B_6job68c48_0),.clk(gclk));
	jdff dff_B_ZvxRwRnz6_0(.din(w_dff_B_6job68c48_0),.dout(w_dff_B_ZvxRwRnz6_0),.clk(gclk));
	jdff dff_B_ODhguznM4_0(.din(w_dff_B_ZvxRwRnz6_0),.dout(w_dff_B_ODhguznM4_0),.clk(gclk));
	jdff dff_B_il1gIN9f0_0(.din(w_dff_B_ODhguznM4_0),.dout(w_dff_B_il1gIN9f0_0),.clk(gclk));
	jdff dff_B_BD0PLByC2_0(.din(w_dff_B_il1gIN9f0_0),.dout(w_dff_B_BD0PLByC2_0),.clk(gclk));
	jdff dff_B_NjlY0O9g5_0(.din(w_dff_B_BD0PLByC2_0),.dout(w_dff_B_NjlY0O9g5_0),.clk(gclk));
	jdff dff_B_VEx44Apl7_0(.din(w_dff_B_NjlY0O9g5_0),.dout(w_dff_B_VEx44Apl7_0),.clk(gclk));
	jdff dff_B_DeHnzkIw8_0(.din(w_dff_B_VEx44Apl7_0),.dout(w_dff_B_DeHnzkIw8_0),.clk(gclk));
	jdff dff_B_OJQ39A6f8_0(.din(w_dff_B_DeHnzkIw8_0),.dout(w_dff_B_OJQ39A6f8_0),.clk(gclk));
	jdff dff_B_YTJNs6OE9_0(.din(w_dff_B_OJQ39A6f8_0),.dout(w_dff_B_YTJNs6OE9_0),.clk(gclk));
	jdff dff_B_YyW5ipZv0_0(.din(w_dff_B_YTJNs6OE9_0),.dout(w_dff_B_YyW5ipZv0_0),.clk(gclk));
	jdff dff_B_bQJvc0Ve4_1(.din(n690),.dout(w_dff_B_bQJvc0Ve4_1),.clk(gclk));
	jdff dff_B_zpqlmqQV7_1(.din(w_dff_B_bQJvc0Ve4_1),.dout(w_dff_B_zpqlmqQV7_1),.clk(gclk));
	jdff dff_B_rXaYLGdB1_1(.din(w_dff_B_zpqlmqQV7_1),.dout(w_dff_B_rXaYLGdB1_1),.clk(gclk));
	jdff dff_B_tDQKSBf49_1(.din(w_dff_B_rXaYLGdB1_1),.dout(w_dff_B_tDQKSBf49_1),.clk(gclk));
	jdff dff_B_ZgIzSM0g2_1(.din(w_dff_B_tDQKSBf49_1),.dout(w_dff_B_ZgIzSM0g2_1),.clk(gclk));
	jdff dff_B_EzlASfqV0_1(.din(w_dff_B_ZgIzSM0g2_1),.dout(w_dff_B_EzlASfqV0_1),.clk(gclk));
	jdff dff_B_zOtsgs4y5_1(.din(w_dff_B_EzlASfqV0_1),.dout(w_dff_B_zOtsgs4y5_1),.clk(gclk));
	jdff dff_B_3HiJEepv8_1(.din(w_dff_B_zOtsgs4y5_1),.dout(w_dff_B_3HiJEepv8_1),.clk(gclk));
	jdff dff_B_mH5nxX8w0_1(.din(w_dff_B_3HiJEepv8_1),.dout(w_dff_B_mH5nxX8w0_1),.clk(gclk));
	jdff dff_B_yXRxkrjl3_1(.din(w_dff_B_mH5nxX8w0_1),.dout(w_dff_B_yXRxkrjl3_1),.clk(gclk));
	jdff dff_B_EsEpf7x14_1(.din(w_dff_B_yXRxkrjl3_1),.dout(w_dff_B_EsEpf7x14_1),.clk(gclk));
	jdff dff_B_ePEQmxLZ0_1(.din(w_dff_B_EsEpf7x14_1),.dout(w_dff_B_ePEQmxLZ0_1),.clk(gclk));
	jdff dff_B_cwlunOWY5_1(.din(w_dff_B_ePEQmxLZ0_1),.dout(w_dff_B_cwlunOWY5_1),.clk(gclk));
	jdff dff_B_2raQsTBN5_1(.din(w_dff_B_cwlunOWY5_1),.dout(w_dff_B_2raQsTBN5_1),.clk(gclk));
	jdff dff_B_VtKk39hK5_1(.din(w_dff_B_2raQsTBN5_1),.dout(w_dff_B_VtKk39hK5_1),.clk(gclk));
	jdff dff_B_GDcWeBkl4_1(.din(w_dff_B_VtKk39hK5_1),.dout(w_dff_B_GDcWeBkl4_1),.clk(gclk));
	jdff dff_B_0nDkNwCJ9_1(.din(w_dff_B_GDcWeBkl4_1),.dout(w_dff_B_0nDkNwCJ9_1),.clk(gclk));
	jdff dff_B_xQaQhewD5_1(.din(w_dff_B_0nDkNwCJ9_1),.dout(w_dff_B_xQaQhewD5_1),.clk(gclk));
	jdff dff_B_NwSl4ljJ9_1(.din(w_dff_B_xQaQhewD5_1),.dout(w_dff_B_NwSl4ljJ9_1),.clk(gclk));
	jdff dff_B_fzFNLoXH8_1(.din(w_dff_B_NwSl4ljJ9_1),.dout(w_dff_B_fzFNLoXH8_1),.clk(gclk));
	jdff dff_B_THQVFNnC3_1(.din(w_dff_B_fzFNLoXH8_1),.dout(w_dff_B_THQVFNnC3_1),.clk(gclk));
	jdff dff_B_BVvyncLx5_1(.din(w_dff_B_THQVFNnC3_1),.dout(w_dff_B_BVvyncLx5_1),.clk(gclk));
	jdff dff_B_oBdoHUk20_1(.din(w_dff_B_BVvyncLx5_1),.dout(w_dff_B_oBdoHUk20_1),.clk(gclk));
	jdff dff_B_77BlTrmI7_1(.din(w_dff_B_oBdoHUk20_1),.dout(w_dff_B_77BlTrmI7_1),.clk(gclk));
	jdff dff_B_Akj4xQoO2_1(.din(w_dff_B_77BlTrmI7_1),.dout(w_dff_B_Akj4xQoO2_1),.clk(gclk));
	jdff dff_B_F63teBN88_1(.din(w_dff_B_Akj4xQoO2_1),.dout(w_dff_B_F63teBN88_1),.clk(gclk));
	jdff dff_B_I2cJFXtg8_1(.din(w_dff_B_F63teBN88_1),.dout(w_dff_B_I2cJFXtg8_1),.clk(gclk));
	jdff dff_B_1cEWMqRE4_1(.din(w_dff_B_I2cJFXtg8_1),.dout(w_dff_B_1cEWMqRE4_1),.clk(gclk));
	jdff dff_B_okmk8ej78_1(.din(w_dff_B_1cEWMqRE4_1),.dout(w_dff_B_okmk8ej78_1),.clk(gclk));
	jdff dff_B_kkLOaFPG5_1(.din(w_dff_B_okmk8ej78_1),.dout(w_dff_B_kkLOaFPG5_1),.clk(gclk));
	jdff dff_B_EjC2iTcd4_1(.din(w_dff_B_kkLOaFPG5_1),.dout(w_dff_B_EjC2iTcd4_1),.clk(gclk));
	jdff dff_B_vHvRE9FN1_1(.din(w_dff_B_EjC2iTcd4_1),.dout(w_dff_B_vHvRE9FN1_1),.clk(gclk));
	jdff dff_B_BI742HCc7_1(.din(w_dff_B_vHvRE9FN1_1),.dout(w_dff_B_BI742HCc7_1),.clk(gclk));
	jdff dff_B_MqfxA0Lp3_1(.din(w_dff_B_BI742HCc7_1),.dout(w_dff_B_MqfxA0Lp3_1),.clk(gclk));
	jdff dff_B_Nn016g5K1_1(.din(w_dff_B_MqfxA0Lp3_1),.dout(w_dff_B_Nn016g5K1_1),.clk(gclk));
	jdff dff_B_nfwkgyr70_1(.din(w_dff_B_Nn016g5K1_1),.dout(w_dff_B_nfwkgyr70_1),.clk(gclk));
	jdff dff_B_HYC4HdS17_1(.din(w_dff_B_nfwkgyr70_1),.dout(w_dff_B_HYC4HdS17_1),.clk(gclk));
	jdff dff_B_4Y4qqm3i7_1(.din(w_dff_B_HYC4HdS17_1),.dout(w_dff_B_4Y4qqm3i7_1),.clk(gclk));
	jdff dff_B_CozIy5H87_1(.din(w_dff_B_4Y4qqm3i7_1),.dout(w_dff_B_CozIy5H87_1),.clk(gclk));
	jdff dff_B_06amHgLg0_1(.din(w_dff_B_CozIy5H87_1),.dout(w_dff_B_06amHgLg0_1),.clk(gclk));
	jdff dff_B_dlS9G38y9_1(.din(w_dff_B_06amHgLg0_1),.dout(w_dff_B_dlS9G38y9_1),.clk(gclk));
	jdff dff_B_eCym5FEC1_1(.din(w_dff_B_dlS9G38y9_1),.dout(w_dff_B_eCym5FEC1_1),.clk(gclk));
	jdff dff_B_rmWpV3nV5_1(.din(w_dff_B_eCym5FEC1_1),.dout(w_dff_B_rmWpV3nV5_1),.clk(gclk));
	jdff dff_B_fTEJk2RJ7_1(.din(w_dff_B_rmWpV3nV5_1),.dout(w_dff_B_fTEJk2RJ7_1),.clk(gclk));
	jdff dff_B_YmAS7Fvg3_1(.din(w_dff_B_fTEJk2RJ7_1),.dout(w_dff_B_YmAS7Fvg3_1),.clk(gclk));
	jdff dff_B_ypTX0I4J3_1(.din(w_dff_B_YmAS7Fvg3_1),.dout(w_dff_B_ypTX0I4J3_1),.clk(gclk));
	jdff dff_B_VLimmRyo2_1(.din(w_dff_B_ypTX0I4J3_1),.dout(w_dff_B_VLimmRyo2_1),.clk(gclk));
	jdff dff_B_OmDnhRHM5_1(.din(w_dff_B_VLimmRyo2_1),.dout(w_dff_B_OmDnhRHM5_1),.clk(gclk));
	jdff dff_B_ALskcCGj8_1(.din(w_dff_B_OmDnhRHM5_1),.dout(w_dff_B_ALskcCGj8_1),.clk(gclk));
	jdff dff_B_qfGrphfe9_1(.din(w_dff_B_ALskcCGj8_1),.dout(w_dff_B_qfGrphfe9_1),.clk(gclk));
	jdff dff_B_YvJN65Kw3_1(.din(w_dff_B_qfGrphfe9_1),.dout(w_dff_B_YvJN65Kw3_1),.clk(gclk));
	jdff dff_B_M2Z2Zpi32_0(.din(n691),.dout(w_dff_B_M2Z2Zpi32_0),.clk(gclk));
	jdff dff_B_9BNZtYOb1_0(.din(w_dff_B_M2Z2Zpi32_0),.dout(w_dff_B_9BNZtYOb1_0),.clk(gclk));
	jdff dff_B_urkHJcp67_0(.din(w_dff_B_9BNZtYOb1_0),.dout(w_dff_B_urkHJcp67_0),.clk(gclk));
	jdff dff_B_HYUQAbQz0_0(.din(w_dff_B_urkHJcp67_0),.dout(w_dff_B_HYUQAbQz0_0),.clk(gclk));
	jdff dff_B_6dR6rfDE6_0(.din(w_dff_B_HYUQAbQz0_0),.dout(w_dff_B_6dR6rfDE6_0),.clk(gclk));
	jdff dff_B_NdN26ESU3_0(.din(w_dff_B_6dR6rfDE6_0),.dout(w_dff_B_NdN26ESU3_0),.clk(gclk));
	jdff dff_B_bcAtTlFa1_0(.din(w_dff_B_NdN26ESU3_0),.dout(w_dff_B_bcAtTlFa1_0),.clk(gclk));
	jdff dff_B_cjyUP6Kr0_0(.din(w_dff_B_bcAtTlFa1_0),.dout(w_dff_B_cjyUP6Kr0_0),.clk(gclk));
	jdff dff_B_3AjLE3qU1_0(.din(w_dff_B_cjyUP6Kr0_0),.dout(w_dff_B_3AjLE3qU1_0),.clk(gclk));
	jdff dff_B_QfEyjW9I7_0(.din(w_dff_B_3AjLE3qU1_0),.dout(w_dff_B_QfEyjW9I7_0),.clk(gclk));
	jdff dff_B_I8jMhcO03_0(.din(w_dff_B_QfEyjW9I7_0),.dout(w_dff_B_I8jMhcO03_0),.clk(gclk));
	jdff dff_B_k7RHcAAU8_0(.din(w_dff_B_I8jMhcO03_0),.dout(w_dff_B_k7RHcAAU8_0),.clk(gclk));
	jdff dff_B_FAE4LRK28_0(.din(w_dff_B_k7RHcAAU8_0),.dout(w_dff_B_FAE4LRK28_0),.clk(gclk));
	jdff dff_B_Tsy8CsY51_0(.din(w_dff_B_FAE4LRK28_0),.dout(w_dff_B_Tsy8CsY51_0),.clk(gclk));
	jdff dff_B_qzVPgNDZ8_0(.din(w_dff_B_Tsy8CsY51_0),.dout(w_dff_B_qzVPgNDZ8_0),.clk(gclk));
	jdff dff_B_Gezd239A1_0(.din(w_dff_B_qzVPgNDZ8_0),.dout(w_dff_B_Gezd239A1_0),.clk(gclk));
	jdff dff_B_nyhxF0bx7_0(.din(w_dff_B_Gezd239A1_0),.dout(w_dff_B_nyhxF0bx7_0),.clk(gclk));
	jdff dff_B_d24qscAP0_0(.din(w_dff_B_nyhxF0bx7_0),.dout(w_dff_B_d24qscAP0_0),.clk(gclk));
	jdff dff_B_DDGoja6p3_0(.din(w_dff_B_d24qscAP0_0),.dout(w_dff_B_DDGoja6p3_0),.clk(gclk));
	jdff dff_B_HLsuJNa15_0(.din(w_dff_B_DDGoja6p3_0),.dout(w_dff_B_HLsuJNa15_0),.clk(gclk));
	jdff dff_B_sTveYXAB5_0(.din(w_dff_B_HLsuJNa15_0),.dout(w_dff_B_sTveYXAB5_0),.clk(gclk));
	jdff dff_B_HidMJlhl6_0(.din(w_dff_B_sTveYXAB5_0),.dout(w_dff_B_HidMJlhl6_0),.clk(gclk));
	jdff dff_B_ls5QBqFE3_0(.din(w_dff_B_HidMJlhl6_0),.dout(w_dff_B_ls5QBqFE3_0),.clk(gclk));
	jdff dff_B_RJOXyWdE1_0(.din(w_dff_B_ls5QBqFE3_0),.dout(w_dff_B_RJOXyWdE1_0),.clk(gclk));
	jdff dff_B_GPTPpF4S8_0(.din(w_dff_B_RJOXyWdE1_0),.dout(w_dff_B_GPTPpF4S8_0),.clk(gclk));
	jdff dff_B_jnx3XdYU8_0(.din(w_dff_B_GPTPpF4S8_0),.dout(w_dff_B_jnx3XdYU8_0),.clk(gclk));
	jdff dff_B_pD6aRnsO7_0(.din(w_dff_B_jnx3XdYU8_0),.dout(w_dff_B_pD6aRnsO7_0),.clk(gclk));
	jdff dff_B_U3E4HFq46_0(.din(w_dff_B_pD6aRnsO7_0),.dout(w_dff_B_U3E4HFq46_0),.clk(gclk));
	jdff dff_B_lyp4tZrL0_0(.din(w_dff_B_U3E4HFq46_0),.dout(w_dff_B_lyp4tZrL0_0),.clk(gclk));
	jdff dff_B_9hDLQRiJ7_0(.din(w_dff_B_lyp4tZrL0_0),.dout(w_dff_B_9hDLQRiJ7_0),.clk(gclk));
	jdff dff_B_HoUpFYSE5_0(.din(w_dff_B_9hDLQRiJ7_0),.dout(w_dff_B_HoUpFYSE5_0),.clk(gclk));
	jdff dff_B_TvI30jHQ4_0(.din(w_dff_B_HoUpFYSE5_0),.dout(w_dff_B_TvI30jHQ4_0),.clk(gclk));
	jdff dff_B_5V8MuIts4_0(.din(w_dff_B_TvI30jHQ4_0),.dout(w_dff_B_5V8MuIts4_0),.clk(gclk));
	jdff dff_B_G1HHMFcq3_0(.din(w_dff_B_5V8MuIts4_0),.dout(w_dff_B_G1HHMFcq3_0),.clk(gclk));
	jdff dff_B_KGGzbHOG1_0(.din(w_dff_B_G1HHMFcq3_0),.dout(w_dff_B_KGGzbHOG1_0),.clk(gclk));
	jdff dff_B_3F0HRwKR7_0(.din(w_dff_B_KGGzbHOG1_0),.dout(w_dff_B_3F0HRwKR7_0),.clk(gclk));
	jdff dff_B_UfRH370V6_0(.din(w_dff_B_3F0HRwKR7_0),.dout(w_dff_B_UfRH370V6_0),.clk(gclk));
	jdff dff_B_p0lZTIYI2_0(.din(w_dff_B_UfRH370V6_0),.dout(w_dff_B_p0lZTIYI2_0),.clk(gclk));
	jdff dff_B_6Sp6LpxQ3_0(.din(w_dff_B_p0lZTIYI2_0),.dout(w_dff_B_6Sp6LpxQ3_0),.clk(gclk));
	jdff dff_B_mYyvAyXV9_0(.din(w_dff_B_6Sp6LpxQ3_0),.dout(w_dff_B_mYyvAyXV9_0),.clk(gclk));
	jdff dff_B_qPvW9PJ80_0(.din(w_dff_B_mYyvAyXV9_0),.dout(w_dff_B_qPvW9PJ80_0),.clk(gclk));
	jdff dff_B_a5RrtU5Q3_0(.din(w_dff_B_qPvW9PJ80_0),.dout(w_dff_B_a5RrtU5Q3_0),.clk(gclk));
	jdff dff_B_Tcb12aoD3_0(.din(w_dff_B_a5RrtU5Q3_0),.dout(w_dff_B_Tcb12aoD3_0),.clk(gclk));
	jdff dff_B_JIoB9FaU8_0(.din(w_dff_B_Tcb12aoD3_0),.dout(w_dff_B_JIoB9FaU8_0),.clk(gclk));
	jdff dff_B_6YMK5mcd7_0(.din(w_dff_B_JIoB9FaU8_0),.dout(w_dff_B_6YMK5mcd7_0),.clk(gclk));
	jdff dff_B_K2CBbsIh3_0(.din(w_dff_B_6YMK5mcd7_0),.dout(w_dff_B_K2CBbsIh3_0),.clk(gclk));
	jdff dff_B_nDNyBPl96_0(.din(w_dff_B_K2CBbsIh3_0),.dout(w_dff_B_nDNyBPl96_0),.clk(gclk));
	jdff dff_B_K3fYR1rs1_0(.din(w_dff_B_nDNyBPl96_0),.dout(w_dff_B_K3fYR1rs1_0),.clk(gclk));
	jdff dff_B_4RgPXNwX4_0(.din(w_dff_B_K3fYR1rs1_0),.dout(w_dff_B_4RgPXNwX4_0),.clk(gclk));
	jdff dff_B_zD5kcOtr8_0(.din(w_dff_B_4RgPXNwX4_0),.dout(w_dff_B_zD5kcOtr8_0),.clk(gclk));
	jdff dff_B_pJXXJjmH2_0(.din(w_dff_B_zD5kcOtr8_0),.dout(w_dff_B_pJXXJjmH2_0),.clk(gclk));
	jdff dff_B_Bn0ayf4l4_1(.din(n684),.dout(w_dff_B_Bn0ayf4l4_1),.clk(gclk));
	jdff dff_B_OPBHspa78_1(.din(w_dff_B_Bn0ayf4l4_1),.dout(w_dff_B_OPBHspa78_1),.clk(gclk));
	jdff dff_B_bUr2KpR36_1(.din(w_dff_B_OPBHspa78_1),.dout(w_dff_B_bUr2KpR36_1),.clk(gclk));
	jdff dff_B_wcblMY8k6_1(.din(w_dff_B_bUr2KpR36_1),.dout(w_dff_B_wcblMY8k6_1),.clk(gclk));
	jdff dff_B_icjOWe594_1(.din(w_dff_B_wcblMY8k6_1),.dout(w_dff_B_icjOWe594_1),.clk(gclk));
	jdff dff_B_gZfppW2h5_1(.din(w_dff_B_icjOWe594_1),.dout(w_dff_B_gZfppW2h5_1),.clk(gclk));
	jdff dff_B_si1WYAmm3_1(.din(w_dff_B_gZfppW2h5_1),.dout(w_dff_B_si1WYAmm3_1),.clk(gclk));
	jdff dff_B_zm2c9Z7N0_1(.din(w_dff_B_si1WYAmm3_1),.dout(w_dff_B_zm2c9Z7N0_1),.clk(gclk));
	jdff dff_B_72KwYpSV6_1(.din(w_dff_B_zm2c9Z7N0_1),.dout(w_dff_B_72KwYpSV6_1),.clk(gclk));
	jdff dff_B_8NxQKTM29_1(.din(w_dff_B_72KwYpSV6_1),.dout(w_dff_B_8NxQKTM29_1),.clk(gclk));
	jdff dff_B_d5auuZ082_1(.din(w_dff_B_8NxQKTM29_1),.dout(w_dff_B_d5auuZ082_1),.clk(gclk));
	jdff dff_B_zUOcucZ45_1(.din(w_dff_B_d5auuZ082_1),.dout(w_dff_B_zUOcucZ45_1),.clk(gclk));
	jdff dff_B_9Doe7fob0_1(.din(w_dff_B_zUOcucZ45_1),.dout(w_dff_B_9Doe7fob0_1),.clk(gclk));
	jdff dff_B_IItQNjhK6_1(.din(w_dff_B_9Doe7fob0_1),.dout(w_dff_B_IItQNjhK6_1),.clk(gclk));
	jdff dff_B_JjFlQL1Y5_1(.din(w_dff_B_IItQNjhK6_1),.dout(w_dff_B_JjFlQL1Y5_1),.clk(gclk));
	jdff dff_B_CNa3mE9S8_1(.din(w_dff_B_JjFlQL1Y5_1),.dout(w_dff_B_CNa3mE9S8_1),.clk(gclk));
	jdff dff_B_CTxuITsz9_1(.din(w_dff_B_CNa3mE9S8_1),.dout(w_dff_B_CTxuITsz9_1),.clk(gclk));
	jdff dff_B_AiRXKI9w3_1(.din(w_dff_B_CTxuITsz9_1),.dout(w_dff_B_AiRXKI9w3_1),.clk(gclk));
	jdff dff_B_5UzYnNcM5_1(.din(w_dff_B_AiRXKI9w3_1),.dout(w_dff_B_5UzYnNcM5_1),.clk(gclk));
	jdff dff_B_UKfwHjPq0_1(.din(w_dff_B_5UzYnNcM5_1),.dout(w_dff_B_UKfwHjPq0_1),.clk(gclk));
	jdff dff_B_me5Mvwh82_1(.din(w_dff_B_UKfwHjPq0_1),.dout(w_dff_B_me5Mvwh82_1),.clk(gclk));
	jdff dff_B_C7YKzlWL4_1(.din(w_dff_B_me5Mvwh82_1),.dout(w_dff_B_C7YKzlWL4_1),.clk(gclk));
	jdff dff_B_SiCu6AZd6_1(.din(w_dff_B_C7YKzlWL4_1),.dout(w_dff_B_SiCu6AZd6_1),.clk(gclk));
	jdff dff_B_1f6dY7SB4_1(.din(w_dff_B_SiCu6AZd6_1),.dout(w_dff_B_1f6dY7SB4_1),.clk(gclk));
	jdff dff_B_cBkaatC65_1(.din(w_dff_B_1f6dY7SB4_1),.dout(w_dff_B_cBkaatC65_1),.clk(gclk));
	jdff dff_B_Py9Fyv2e4_1(.din(w_dff_B_cBkaatC65_1),.dout(w_dff_B_Py9Fyv2e4_1),.clk(gclk));
	jdff dff_B_XR1rBt5N7_1(.din(w_dff_B_Py9Fyv2e4_1),.dout(w_dff_B_XR1rBt5N7_1),.clk(gclk));
	jdff dff_B_TUCQCzOL1_1(.din(w_dff_B_XR1rBt5N7_1),.dout(w_dff_B_TUCQCzOL1_1),.clk(gclk));
	jdff dff_B_b9Fa4T0N5_1(.din(w_dff_B_TUCQCzOL1_1),.dout(w_dff_B_b9Fa4T0N5_1),.clk(gclk));
	jdff dff_B_dLhp6r1k5_1(.din(w_dff_B_b9Fa4T0N5_1),.dout(w_dff_B_dLhp6r1k5_1),.clk(gclk));
	jdff dff_B_KesjSdmP3_1(.din(w_dff_B_dLhp6r1k5_1),.dout(w_dff_B_KesjSdmP3_1),.clk(gclk));
	jdff dff_B_y5dEn2zu7_1(.din(w_dff_B_KesjSdmP3_1),.dout(w_dff_B_y5dEn2zu7_1),.clk(gclk));
	jdff dff_B_U8JxLU4j7_1(.din(w_dff_B_y5dEn2zu7_1),.dout(w_dff_B_U8JxLU4j7_1),.clk(gclk));
	jdff dff_B_rDJUI1sC4_1(.din(w_dff_B_U8JxLU4j7_1),.dout(w_dff_B_rDJUI1sC4_1),.clk(gclk));
	jdff dff_B_Xk4bNTa88_1(.din(w_dff_B_rDJUI1sC4_1),.dout(w_dff_B_Xk4bNTa88_1),.clk(gclk));
	jdff dff_B_n4Po8Bdw4_1(.din(w_dff_B_Xk4bNTa88_1),.dout(w_dff_B_n4Po8Bdw4_1),.clk(gclk));
	jdff dff_B_srHselSA2_1(.din(w_dff_B_n4Po8Bdw4_1),.dout(w_dff_B_srHselSA2_1),.clk(gclk));
	jdff dff_B_OdB1l3Ip0_1(.din(w_dff_B_srHselSA2_1),.dout(w_dff_B_OdB1l3Ip0_1),.clk(gclk));
	jdff dff_B_wF9PpH6P0_1(.din(w_dff_B_OdB1l3Ip0_1),.dout(w_dff_B_wF9PpH6P0_1),.clk(gclk));
	jdff dff_B_923Ba2Vi2_1(.din(w_dff_B_wF9PpH6P0_1),.dout(w_dff_B_923Ba2Vi2_1),.clk(gclk));
	jdff dff_B_t9LnWkL38_1(.din(w_dff_B_923Ba2Vi2_1),.dout(w_dff_B_t9LnWkL38_1),.clk(gclk));
	jdff dff_B_R1frhqzv4_1(.din(w_dff_B_t9LnWkL38_1),.dout(w_dff_B_R1frhqzv4_1),.clk(gclk));
	jdff dff_B_XTZGcLFe9_1(.din(w_dff_B_R1frhqzv4_1),.dout(w_dff_B_XTZGcLFe9_1),.clk(gclk));
	jdff dff_B_2bzqm8vX8_1(.din(w_dff_B_XTZGcLFe9_1),.dout(w_dff_B_2bzqm8vX8_1),.clk(gclk));
	jdff dff_B_giOac33U5_1(.din(w_dff_B_2bzqm8vX8_1),.dout(w_dff_B_giOac33U5_1),.clk(gclk));
	jdff dff_B_juqi6SO07_1(.din(w_dff_B_giOac33U5_1),.dout(w_dff_B_juqi6SO07_1),.clk(gclk));
	jdff dff_B_bkVmEFIp3_1(.din(w_dff_B_juqi6SO07_1),.dout(w_dff_B_bkVmEFIp3_1),.clk(gclk));
	jdff dff_B_NpUfs0ua2_1(.din(w_dff_B_bkVmEFIp3_1),.dout(w_dff_B_NpUfs0ua2_1),.clk(gclk));
	jdff dff_B_j6Xz2bdg7_1(.din(w_dff_B_NpUfs0ua2_1),.dout(w_dff_B_j6Xz2bdg7_1),.clk(gclk));
	jdff dff_B_YfcGYVQq4_1(.din(w_dff_B_j6Xz2bdg7_1),.dout(w_dff_B_YfcGYVQq4_1),.clk(gclk));
	jdff dff_B_o8lKl7m83_0(.din(n685),.dout(w_dff_B_o8lKl7m83_0),.clk(gclk));
	jdff dff_B_m9OuHavv5_0(.din(w_dff_B_o8lKl7m83_0),.dout(w_dff_B_m9OuHavv5_0),.clk(gclk));
	jdff dff_B_gNsFavlC5_0(.din(w_dff_B_m9OuHavv5_0),.dout(w_dff_B_gNsFavlC5_0),.clk(gclk));
	jdff dff_B_GNFIWxiW6_0(.din(w_dff_B_gNsFavlC5_0),.dout(w_dff_B_GNFIWxiW6_0),.clk(gclk));
	jdff dff_B_yztwk1Wg8_0(.din(w_dff_B_GNFIWxiW6_0),.dout(w_dff_B_yztwk1Wg8_0),.clk(gclk));
	jdff dff_B_J5gNqZO42_0(.din(w_dff_B_yztwk1Wg8_0),.dout(w_dff_B_J5gNqZO42_0),.clk(gclk));
	jdff dff_B_jecSgOEO2_0(.din(w_dff_B_J5gNqZO42_0),.dout(w_dff_B_jecSgOEO2_0),.clk(gclk));
	jdff dff_B_nAMmXpDe1_0(.din(w_dff_B_jecSgOEO2_0),.dout(w_dff_B_nAMmXpDe1_0),.clk(gclk));
	jdff dff_B_2CGPr0jL7_0(.din(w_dff_B_nAMmXpDe1_0),.dout(w_dff_B_2CGPr0jL7_0),.clk(gclk));
	jdff dff_B_C8aTMibt1_0(.din(w_dff_B_2CGPr0jL7_0),.dout(w_dff_B_C8aTMibt1_0),.clk(gclk));
	jdff dff_B_oEasvFXR1_0(.din(w_dff_B_C8aTMibt1_0),.dout(w_dff_B_oEasvFXR1_0),.clk(gclk));
	jdff dff_B_jX7N9V0l2_0(.din(w_dff_B_oEasvFXR1_0),.dout(w_dff_B_jX7N9V0l2_0),.clk(gclk));
	jdff dff_B_nhHmOG3l9_0(.din(w_dff_B_jX7N9V0l2_0),.dout(w_dff_B_nhHmOG3l9_0),.clk(gclk));
	jdff dff_B_2zfAyqfA1_0(.din(w_dff_B_nhHmOG3l9_0),.dout(w_dff_B_2zfAyqfA1_0),.clk(gclk));
	jdff dff_B_79j2RWhB7_0(.din(w_dff_B_2zfAyqfA1_0),.dout(w_dff_B_79j2RWhB7_0),.clk(gclk));
	jdff dff_B_Mipow4lI7_0(.din(w_dff_B_79j2RWhB7_0),.dout(w_dff_B_Mipow4lI7_0),.clk(gclk));
	jdff dff_B_tgjkLOLF0_0(.din(w_dff_B_Mipow4lI7_0),.dout(w_dff_B_tgjkLOLF0_0),.clk(gclk));
	jdff dff_B_M8j2y6Gb9_0(.din(w_dff_B_tgjkLOLF0_0),.dout(w_dff_B_M8j2y6Gb9_0),.clk(gclk));
	jdff dff_B_GcV2SYhj9_0(.din(w_dff_B_M8j2y6Gb9_0),.dout(w_dff_B_GcV2SYhj9_0),.clk(gclk));
	jdff dff_B_3wIQeuvn5_0(.din(w_dff_B_GcV2SYhj9_0),.dout(w_dff_B_3wIQeuvn5_0),.clk(gclk));
	jdff dff_B_6PdG8ZXr7_0(.din(w_dff_B_3wIQeuvn5_0),.dout(w_dff_B_6PdG8ZXr7_0),.clk(gclk));
	jdff dff_B_nSRU9s8V7_0(.din(w_dff_B_6PdG8ZXr7_0),.dout(w_dff_B_nSRU9s8V7_0),.clk(gclk));
	jdff dff_B_XQuVQhQs3_0(.din(w_dff_B_nSRU9s8V7_0),.dout(w_dff_B_XQuVQhQs3_0),.clk(gclk));
	jdff dff_B_0ZJBcOC74_0(.din(w_dff_B_XQuVQhQs3_0),.dout(w_dff_B_0ZJBcOC74_0),.clk(gclk));
	jdff dff_B_lTAhuV0P1_0(.din(w_dff_B_0ZJBcOC74_0),.dout(w_dff_B_lTAhuV0P1_0),.clk(gclk));
	jdff dff_B_iZTbxxbL3_0(.din(w_dff_B_lTAhuV0P1_0),.dout(w_dff_B_iZTbxxbL3_0),.clk(gclk));
	jdff dff_B_xNYiCHiy4_0(.din(w_dff_B_iZTbxxbL3_0),.dout(w_dff_B_xNYiCHiy4_0),.clk(gclk));
	jdff dff_B_ZdkeEZqT4_0(.din(w_dff_B_xNYiCHiy4_0),.dout(w_dff_B_ZdkeEZqT4_0),.clk(gclk));
	jdff dff_B_6wYHZRJa3_0(.din(w_dff_B_ZdkeEZqT4_0),.dout(w_dff_B_6wYHZRJa3_0),.clk(gclk));
	jdff dff_B_nLpqIPr92_0(.din(w_dff_B_6wYHZRJa3_0),.dout(w_dff_B_nLpqIPr92_0),.clk(gclk));
	jdff dff_B_rypsM0rh5_0(.din(w_dff_B_nLpqIPr92_0),.dout(w_dff_B_rypsM0rh5_0),.clk(gclk));
	jdff dff_B_oJrbA7549_0(.din(w_dff_B_rypsM0rh5_0),.dout(w_dff_B_oJrbA7549_0),.clk(gclk));
	jdff dff_B_2MgsdNv10_0(.din(w_dff_B_oJrbA7549_0),.dout(w_dff_B_2MgsdNv10_0),.clk(gclk));
	jdff dff_B_nvUQFevb7_0(.din(w_dff_B_2MgsdNv10_0),.dout(w_dff_B_nvUQFevb7_0),.clk(gclk));
	jdff dff_B_Qz2Aludt3_0(.din(w_dff_B_nvUQFevb7_0),.dout(w_dff_B_Qz2Aludt3_0),.clk(gclk));
	jdff dff_B_aFt5mB8r1_0(.din(w_dff_B_Qz2Aludt3_0),.dout(w_dff_B_aFt5mB8r1_0),.clk(gclk));
	jdff dff_B_nCJQ1OO02_0(.din(w_dff_B_aFt5mB8r1_0),.dout(w_dff_B_nCJQ1OO02_0),.clk(gclk));
	jdff dff_B_GOrBIJIZ5_0(.din(w_dff_B_nCJQ1OO02_0),.dout(w_dff_B_GOrBIJIZ5_0),.clk(gclk));
	jdff dff_B_HWXM8W3R5_0(.din(w_dff_B_GOrBIJIZ5_0),.dout(w_dff_B_HWXM8W3R5_0),.clk(gclk));
	jdff dff_B_0HvLrBnk7_0(.din(w_dff_B_HWXM8W3R5_0),.dout(w_dff_B_0HvLrBnk7_0),.clk(gclk));
	jdff dff_B_wMph96Ty8_0(.din(w_dff_B_0HvLrBnk7_0),.dout(w_dff_B_wMph96Ty8_0),.clk(gclk));
	jdff dff_B_Bf7cOeaZ6_0(.din(w_dff_B_wMph96Ty8_0),.dout(w_dff_B_Bf7cOeaZ6_0),.clk(gclk));
	jdff dff_B_tVxHdxMC3_0(.din(w_dff_B_Bf7cOeaZ6_0),.dout(w_dff_B_tVxHdxMC3_0),.clk(gclk));
	jdff dff_B_cCv8HaBD0_0(.din(w_dff_B_tVxHdxMC3_0),.dout(w_dff_B_cCv8HaBD0_0),.clk(gclk));
	jdff dff_B_0Tpg07rk5_0(.din(w_dff_B_cCv8HaBD0_0),.dout(w_dff_B_0Tpg07rk5_0),.clk(gclk));
	jdff dff_B_bKzotIXb8_0(.din(w_dff_B_0Tpg07rk5_0),.dout(w_dff_B_bKzotIXb8_0),.clk(gclk));
	jdff dff_B_QTJk9WmN1_0(.din(w_dff_B_bKzotIXb8_0),.dout(w_dff_B_QTJk9WmN1_0),.clk(gclk));
	jdff dff_B_XUO0cnc56_0(.din(w_dff_B_QTJk9WmN1_0),.dout(w_dff_B_XUO0cnc56_0),.clk(gclk));
	jdff dff_B_zAV1WpsN2_0(.din(w_dff_B_XUO0cnc56_0),.dout(w_dff_B_zAV1WpsN2_0),.clk(gclk));
	jdff dff_B_puRmXWhG3_0(.din(w_dff_B_zAV1WpsN2_0),.dout(w_dff_B_puRmXWhG3_0),.clk(gclk));
	jdff dff_B_5kNCBtc74_1(.din(n678),.dout(w_dff_B_5kNCBtc74_1),.clk(gclk));
	jdff dff_B_uoXHR67E5_1(.din(w_dff_B_5kNCBtc74_1),.dout(w_dff_B_uoXHR67E5_1),.clk(gclk));
	jdff dff_B_1ZwEeslb3_1(.din(w_dff_B_uoXHR67E5_1),.dout(w_dff_B_1ZwEeslb3_1),.clk(gclk));
	jdff dff_B_Vu1XErOu6_1(.din(w_dff_B_1ZwEeslb3_1),.dout(w_dff_B_Vu1XErOu6_1),.clk(gclk));
	jdff dff_B_S0oXXYtW8_1(.din(w_dff_B_Vu1XErOu6_1),.dout(w_dff_B_S0oXXYtW8_1),.clk(gclk));
	jdff dff_B_8hiwjcQm3_1(.din(w_dff_B_S0oXXYtW8_1),.dout(w_dff_B_8hiwjcQm3_1),.clk(gclk));
	jdff dff_B_VaCA9vCu2_1(.din(w_dff_B_8hiwjcQm3_1),.dout(w_dff_B_VaCA9vCu2_1),.clk(gclk));
	jdff dff_B_NEOb3VVp4_1(.din(w_dff_B_VaCA9vCu2_1),.dout(w_dff_B_NEOb3VVp4_1),.clk(gclk));
	jdff dff_B_uxmPXaA96_1(.din(w_dff_B_NEOb3VVp4_1),.dout(w_dff_B_uxmPXaA96_1),.clk(gclk));
	jdff dff_B_SeGm6zRR2_1(.din(w_dff_B_uxmPXaA96_1),.dout(w_dff_B_SeGm6zRR2_1),.clk(gclk));
	jdff dff_B_plgHfCGH5_1(.din(w_dff_B_SeGm6zRR2_1),.dout(w_dff_B_plgHfCGH5_1),.clk(gclk));
	jdff dff_B_C5jDYmwz1_1(.din(w_dff_B_plgHfCGH5_1),.dout(w_dff_B_C5jDYmwz1_1),.clk(gclk));
	jdff dff_B_VwM0htNJ5_1(.din(w_dff_B_C5jDYmwz1_1),.dout(w_dff_B_VwM0htNJ5_1),.clk(gclk));
	jdff dff_B_0JdZOWma5_1(.din(w_dff_B_VwM0htNJ5_1),.dout(w_dff_B_0JdZOWma5_1),.clk(gclk));
	jdff dff_B_wK7wchF66_1(.din(w_dff_B_0JdZOWma5_1),.dout(w_dff_B_wK7wchF66_1),.clk(gclk));
	jdff dff_B_tDKb11eW6_1(.din(w_dff_B_wK7wchF66_1),.dout(w_dff_B_tDKb11eW6_1),.clk(gclk));
	jdff dff_B_xLCAc80U8_1(.din(w_dff_B_tDKb11eW6_1),.dout(w_dff_B_xLCAc80U8_1),.clk(gclk));
	jdff dff_B_snmgibni4_1(.din(w_dff_B_xLCAc80U8_1),.dout(w_dff_B_snmgibni4_1),.clk(gclk));
	jdff dff_B_P3rbp7P50_1(.din(w_dff_B_snmgibni4_1),.dout(w_dff_B_P3rbp7P50_1),.clk(gclk));
	jdff dff_B_D5Y9nkM24_1(.din(w_dff_B_P3rbp7P50_1),.dout(w_dff_B_D5Y9nkM24_1),.clk(gclk));
	jdff dff_B_7esFzaJc1_1(.din(w_dff_B_D5Y9nkM24_1),.dout(w_dff_B_7esFzaJc1_1),.clk(gclk));
	jdff dff_B_Vj0rlalk2_1(.din(w_dff_B_7esFzaJc1_1),.dout(w_dff_B_Vj0rlalk2_1),.clk(gclk));
	jdff dff_B_6YqNFGIg7_1(.din(w_dff_B_Vj0rlalk2_1),.dout(w_dff_B_6YqNFGIg7_1),.clk(gclk));
	jdff dff_B_v0ep1tLh9_1(.din(w_dff_B_6YqNFGIg7_1),.dout(w_dff_B_v0ep1tLh9_1),.clk(gclk));
	jdff dff_B_dkWHpMiA5_1(.din(w_dff_B_v0ep1tLh9_1),.dout(w_dff_B_dkWHpMiA5_1),.clk(gclk));
	jdff dff_B_N6bZIXBS3_1(.din(w_dff_B_dkWHpMiA5_1),.dout(w_dff_B_N6bZIXBS3_1),.clk(gclk));
	jdff dff_B_Vw5v93c62_1(.din(w_dff_B_N6bZIXBS3_1),.dout(w_dff_B_Vw5v93c62_1),.clk(gclk));
	jdff dff_B_Y7f2ZDFI3_1(.din(w_dff_B_Vw5v93c62_1),.dout(w_dff_B_Y7f2ZDFI3_1),.clk(gclk));
	jdff dff_B_nw43XgZG2_1(.din(w_dff_B_Y7f2ZDFI3_1),.dout(w_dff_B_nw43XgZG2_1),.clk(gclk));
	jdff dff_B_2BrZbtDu9_1(.din(w_dff_B_nw43XgZG2_1),.dout(w_dff_B_2BrZbtDu9_1),.clk(gclk));
	jdff dff_B_tokFQjsw5_1(.din(w_dff_B_2BrZbtDu9_1),.dout(w_dff_B_tokFQjsw5_1),.clk(gclk));
	jdff dff_B_nulaadlk4_1(.din(w_dff_B_tokFQjsw5_1),.dout(w_dff_B_nulaadlk4_1),.clk(gclk));
	jdff dff_B_wUKrFFBA3_1(.din(w_dff_B_nulaadlk4_1),.dout(w_dff_B_wUKrFFBA3_1),.clk(gclk));
	jdff dff_B_V4imVhSE2_1(.din(w_dff_B_wUKrFFBA3_1),.dout(w_dff_B_V4imVhSE2_1),.clk(gclk));
	jdff dff_B_ifZ4tcSX1_1(.din(w_dff_B_V4imVhSE2_1),.dout(w_dff_B_ifZ4tcSX1_1),.clk(gclk));
	jdff dff_B_5B80bnKd4_1(.din(w_dff_B_ifZ4tcSX1_1),.dout(w_dff_B_5B80bnKd4_1),.clk(gclk));
	jdff dff_B_wtpp65Ik2_1(.din(w_dff_B_5B80bnKd4_1),.dout(w_dff_B_wtpp65Ik2_1),.clk(gclk));
	jdff dff_B_zkt4Jsye9_1(.din(w_dff_B_wtpp65Ik2_1),.dout(w_dff_B_zkt4Jsye9_1),.clk(gclk));
	jdff dff_B_QTuSFALZ7_1(.din(w_dff_B_zkt4Jsye9_1),.dout(w_dff_B_QTuSFALZ7_1),.clk(gclk));
	jdff dff_B_Fflv2MGN1_1(.din(w_dff_B_QTuSFALZ7_1),.dout(w_dff_B_Fflv2MGN1_1),.clk(gclk));
	jdff dff_B_gSOESurT3_1(.din(w_dff_B_Fflv2MGN1_1),.dout(w_dff_B_gSOESurT3_1),.clk(gclk));
	jdff dff_B_zLpnZT2N8_1(.din(w_dff_B_gSOESurT3_1),.dout(w_dff_B_zLpnZT2N8_1),.clk(gclk));
	jdff dff_B_MS6rJ1o08_1(.din(w_dff_B_zLpnZT2N8_1),.dout(w_dff_B_MS6rJ1o08_1),.clk(gclk));
	jdff dff_B_1bb3jT2z7_1(.din(w_dff_B_MS6rJ1o08_1),.dout(w_dff_B_1bb3jT2z7_1),.clk(gclk));
	jdff dff_B_UxfLqzNf8_1(.din(w_dff_B_1bb3jT2z7_1),.dout(w_dff_B_UxfLqzNf8_1),.clk(gclk));
	jdff dff_B_rvgwMEOG7_1(.din(w_dff_B_UxfLqzNf8_1),.dout(w_dff_B_rvgwMEOG7_1),.clk(gclk));
	jdff dff_B_ftd9imrv6_1(.din(w_dff_B_rvgwMEOG7_1),.dout(w_dff_B_ftd9imrv6_1),.clk(gclk));
	jdff dff_B_ITNKsc4Y9_1(.din(w_dff_B_ftd9imrv6_1),.dout(w_dff_B_ITNKsc4Y9_1),.clk(gclk));
	jdff dff_B_GecnHXzy9_1(.din(w_dff_B_ITNKsc4Y9_1),.dout(w_dff_B_GecnHXzy9_1),.clk(gclk));
	jdff dff_B_RYLpmxO94_0(.din(n679),.dout(w_dff_B_RYLpmxO94_0),.clk(gclk));
	jdff dff_B_G13H5dCi3_0(.din(w_dff_B_RYLpmxO94_0),.dout(w_dff_B_G13H5dCi3_0),.clk(gclk));
	jdff dff_B_ezjcyRii5_0(.din(w_dff_B_G13H5dCi3_0),.dout(w_dff_B_ezjcyRii5_0),.clk(gclk));
	jdff dff_B_XVFFCW5k8_0(.din(w_dff_B_ezjcyRii5_0),.dout(w_dff_B_XVFFCW5k8_0),.clk(gclk));
	jdff dff_B_1X2vffpK4_0(.din(w_dff_B_XVFFCW5k8_0),.dout(w_dff_B_1X2vffpK4_0),.clk(gclk));
	jdff dff_B_5quM9VZJ2_0(.din(w_dff_B_1X2vffpK4_0),.dout(w_dff_B_5quM9VZJ2_0),.clk(gclk));
	jdff dff_B_xqYvSQZX6_0(.din(w_dff_B_5quM9VZJ2_0),.dout(w_dff_B_xqYvSQZX6_0),.clk(gclk));
	jdff dff_B_OynyNYX33_0(.din(w_dff_B_xqYvSQZX6_0),.dout(w_dff_B_OynyNYX33_0),.clk(gclk));
	jdff dff_B_wmDOAMH98_0(.din(w_dff_B_OynyNYX33_0),.dout(w_dff_B_wmDOAMH98_0),.clk(gclk));
	jdff dff_B_ymvk5kmL8_0(.din(w_dff_B_wmDOAMH98_0),.dout(w_dff_B_ymvk5kmL8_0),.clk(gclk));
	jdff dff_B_jyUaxdDZ9_0(.din(w_dff_B_ymvk5kmL8_0),.dout(w_dff_B_jyUaxdDZ9_0),.clk(gclk));
	jdff dff_B_TwIaURru0_0(.din(w_dff_B_jyUaxdDZ9_0),.dout(w_dff_B_TwIaURru0_0),.clk(gclk));
	jdff dff_B_lVYmrqF10_0(.din(w_dff_B_TwIaURru0_0),.dout(w_dff_B_lVYmrqF10_0),.clk(gclk));
	jdff dff_B_jQ2558Mk1_0(.din(w_dff_B_lVYmrqF10_0),.dout(w_dff_B_jQ2558Mk1_0),.clk(gclk));
	jdff dff_B_96muY35c1_0(.din(w_dff_B_jQ2558Mk1_0),.dout(w_dff_B_96muY35c1_0),.clk(gclk));
	jdff dff_B_zC14Kwyq9_0(.din(w_dff_B_96muY35c1_0),.dout(w_dff_B_zC14Kwyq9_0),.clk(gclk));
	jdff dff_B_QnUjg5pl5_0(.din(w_dff_B_zC14Kwyq9_0),.dout(w_dff_B_QnUjg5pl5_0),.clk(gclk));
	jdff dff_B_Wn9SE4811_0(.din(w_dff_B_QnUjg5pl5_0),.dout(w_dff_B_Wn9SE4811_0),.clk(gclk));
	jdff dff_B_arigDJuU6_0(.din(w_dff_B_Wn9SE4811_0),.dout(w_dff_B_arigDJuU6_0),.clk(gclk));
	jdff dff_B_hHmelqxt8_0(.din(w_dff_B_arigDJuU6_0),.dout(w_dff_B_hHmelqxt8_0),.clk(gclk));
	jdff dff_B_wDalVPYk4_0(.din(w_dff_B_hHmelqxt8_0),.dout(w_dff_B_wDalVPYk4_0),.clk(gclk));
	jdff dff_B_XgFvN2AZ3_0(.din(w_dff_B_wDalVPYk4_0),.dout(w_dff_B_XgFvN2AZ3_0),.clk(gclk));
	jdff dff_B_Idhox2Iw6_0(.din(w_dff_B_XgFvN2AZ3_0),.dout(w_dff_B_Idhox2Iw6_0),.clk(gclk));
	jdff dff_B_5cvJRhJw0_0(.din(w_dff_B_Idhox2Iw6_0),.dout(w_dff_B_5cvJRhJw0_0),.clk(gclk));
	jdff dff_B_TYDBNPwG1_0(.din(w_dff_B_5cvJRhJw0_0),.dout(w_dff_B_TYDBNPwG1_0),.clk(gclk));
	jdff dff_B_46eipWmF1_0(.din(w_dff_B_TYDBNPwG1_0),.dout(w_dff_B_46eipWmF1_0),.clk(gclk));
	jdff dff_B_VQPO9YMH9_0(.din(w_dff_B_46eipWmF1_0),.dout(w_dff_B_VQPO9YMH9_0),.clk(gclk));
	jdff dff_B_nCrUplG55_0(.din(w_dff_B_VQPO9YMH9_0),.dout(w_dff_B_nCrUplG55_0),.clk(gclk));
	jdff dff_B_mise7VtT4_0(.din(w_dff_B_nCrUplG55_0),.dout(w_dff_B_mise7VtT4_0),.clk(gclk));
	jdff dff_B_9nz9xISJ3_0(.din(w_dff_B_mise7VtT4_0),.dout(w_dff_B_9nz9xISJ3_0),.clk(gclk));
	jdff dff_B_XEwqnxQC9_0(.din(w_dff_B_9nz9xISJ3_0),.dout(w_dff_B_XEwqnxQC9_0),.clk(gclk));
	jdff dff_B_9Y7rA5TP6_0(.din(w_dff_B_XEwqnxQC9_0),.dout(w_dff_B_9Y7rA5TP6_0),.clk(gclk));
	jdff dff_B_50PypCeG2_0(.din(w_dff_B_9Y7rA5TP6_0),.dout(w_dff_B_50PypCeG2_0),.clk(gclk));
	jdff dff_B_rqJwqihk6_0(.din(w_dff_B_50PypCeG2_0),.dout(w_dff_B_rqJwqihk6_0),.clk(gclk));
	jdff dff_B_fhUqZg6j4_0(.din(w_dff_B_rqJwqihk6_0),.dout(w_dff_B_fhUqZg6j4_0),.clk(gclk));
	jdff dff_B_3HJqArCw7_0(.din(w_dff_B_fhUqZg6j4_0),.dout(w_dff_B_3HJqArCw7_0),.clk(gclk));
	jdff dff_B_uEFjUHwe5_0(.din(w_dff_B_3HJqArCw7_0),.dout(w_dff_B_uEFjUHwe5_0),.clk(gclk));
	jdff dff_B_kYsVhlIg9_0(.din(w_dff_B_uEFjUHwe5_0),.dout(w_dff_B_kYsVhlIg9_0),.clk(gclk));
	jdff dff_B_gzPfgmdf1_0(.din(w_dff_B_kYsVhlIg9_0),.dout(w_dff_B_gzPfgmdf1_0),.clk(gclk));
	jdff dff_B_eQqM7EEQ8_0(.din(w_dff_B_gzPfgmdf1_0),.dout(w_dff_B_eQqM7EEQ8_0),.clk(gclk));
	jdff dff_B_zKUvKSTu6_0(.din(w_dff_B_eQqM7EEQ8_0),.dout(w_dff_B_zKUvKSTu6_0),.clk(gclk));
	jdff dff_B_H8PZzNAC0_0(.din(w_dff_B_zKUvKSTu6_0),.dout(w_dff_B_H8PZzNAC0_0),.clk(gclk));
	jdff dff_B_Rb4ms70y4_0(.din(w_dff_B_H8PZzNAC0_0),.dout(w_dff_B_Rb4ms70y4_0),.clk(gclk));
	jdff dff_B_uaqzDU7K0_0(.din(w_dff_B_Rb4ms70y4_0),.dout(w_dff_B_uaqzDU7K0_0),.clk(gclk));
	jdff dff_B_yvUUtoGq8_0(.din(w_dff_B_uaqzDU7K0_0),.dout(w_dff_B_yvUUtoGq8_0),.clk(gclk));
	jdff dff_B_6PmNXT3k8_0(.din(w_dff_B_yvUUtoGq8_0),.dout(w_dff_B_6PmNXT3k8_0),.clk(gclk));
	jdff dff_B_9D24XVkK7_0(.din(w_dff_B_6PmNXT3k8_0),.dout(w_dff_B_9D24XVkK7_0),.clk(gclk));
	jdff dff_B_5p3UXoCp3_0(.din(w_dff_B_9D24XVkK7_0),.dout(w_dff_B_5p3UXoCp3_0),.clk(gclk));
	jdff dff_B_CtINLd6Q5_0(.din(w_dff_B_5p3UXoCp3_0),.dout(w_dff_B_CtINLd6Q5_0),.clk(gclk));
	jdff dff_B_6sCSTLSj4_1(.din(n672),.dout(w_dff_B_6sCSTLSj4_1),.clk(gclk));
	jdff dff_B_GvGqxZ3V3_1(.din(w_dff_B_6sCSTLSj4_1),.dout(w_dff_B_GvGqxZ3V3_1),.clk(gclk));
	jdff dff_B_hWFjEYmV3_1(.din(w_dff_B_GvGqxZ3V3_1),.dout(w_dff_B_hWFjEYmV3_1),.clk(gclk));
	jdff dff_B_6crFkfLe6_1(.din(w_dff_B_hWFjEYmV3_1),.dout(w_dff_B_6crFkfLe6_1),.clk(gclk));
	jdff dff_B_DjMlEltp7_1(.din(w_dff_B_6crFkfLe6_1),.dout(w_dff_B_DjMlEltp7_1),.clk(gclk));
	jdff dff_B_Gry2k59O3_1(.din(w_dff_B_DjMlEltp7_1),.dout(w_dff_B_Gry2k59O3_1),.clk(gclk));
	jdff dff_B_VYsM1v2D8_1(.din(w_dff_B_Gry2k59O3_1),.dout(w_dff_B_VYsM1v2D8_1),.clk(gclk));
	jdff dff_B_VmyNWgjk3_1(.din(w_dff_B_VYsM1v2D8_1),.dout(w_dff_B_VmyNWgjk3_1),.clk(gclk));
	jdff dff_B_JDJFjqGW1_1(.din(w_dff_B_VmyNWgjk3_1),.dout(w_dff_B_JDJFjqGW1_1),.clk(gclk));
	jdff dff_B_DkBYT4ie2_1(.din(w_dff_B_JDJFjqGW1_1),.dout(w_dff_B_DkBYT4ie2_1),.clk(gclk));
	jdff dff_B_PwBl56if5_1(.din(w_dff_B_DkBYT4ie2_1),.dout(w_dff_B_PwBl56if5_1),.clk(gclk));
	jdff dff_B_yLKumY2s4_1(.din(w_dff_B_PwBl56if5_1),.dout(w_dff_B_yLKumY2s4_1),.clk(gclk));
	jdff dff_B_KLAVQKdh3_1(.din(w_dff_B_yLKumY2s4_1),.dout(w_dff_B_KLAVQKdh3_1),.clk(gclk));
	jdff dff_B_t4pfyRXO9_1(.din(w_dff_B_KLAVQKdh3_1),.dout(w_dff_B_t4pfyRXO9_1),.clk(gclk));
	jdff dff_B_Rqu0kexE4_1(.din(w_dff_B_t4pfyRXO9_1),.dout(w_dff_B_Rqu0kexE4_1),.clk(gclk));
	jdff dff_B_NIkRan838_1(.din(w_dff_B_Rqu0kexE4_1),.dout(w_dff_B_NIkRan838_1),.clk(gclk));
	jdff dff_B_31ln5hJh9_1(.din(w_dff_B_NIkRan838_1),.dout(w_dff_B_31ln5hJh9_1),.clk(gclk));
	jdff dff_B_99R7wNjY7_1(.din(w_dff_B_31ln5hJh9_1),.dout(w_dff_B_99R7wNjY7_1),.clk(gclk));
	jdff dff_B_Rj55s4yc2_1(.din(w_dff_B_99R7wNjY7_1),.dout(w_dff_B_Rj55s4yc2_1),.clk(gclk));
	jdff dff_B_FWEtqpvL3_1(.din(w_dff_B_Rj55s4yc2_1),.dout(w_dff_B_FWEtqpvL3_1),.clk(gclk));
	jdff dff_B_W78dtbey3_1(.din(w_dff_B_FWEtqpvL3_1),.dout(w_dff_B_W78dtbey3_1),.clk(gclk));
	jdff dff_B_pqhKhvzM5_1(.din(w_dff_B_W78dtbey3_1),.dout(w_dff_B_pqhKhvzM5_1),.clk(gclk));
	jdff dff_B_EEOq5RlS0_1(.din(w_dff_B_pqhKhvzM5_1),.dout(w_dff_B_EEOq5RlS0_1),.clk(gclk));
	jdff dff_B_WUkmjuyB8_1(.din(w_dff_B_EEOq5RlS0_1),.dout(w_dff_B_WUkmjuyB8_1),.clk(gclk));
	jdff dff_B_ExzLkwKL5_1(.din(w_dff_B_WUkmjuyB8_1),.dout(w_dff_B_ExzLkwKL5_1),.clk(gclk));
	jdff dff_B_wxpM6EWG3_1(.din(w_dff_B_ExzLkwKL5_1),.dout(w_dff_B_wxpM6EWG3_1),.clk(gclk));
	jdff dff_B_BePO5IXJ4_1(.din(w_dff_B_wxpM6EWG3_1),.dout(w_dff_B_BePO5IXJ4_1),.clk(gclk));
	jdff dff_B_5nJkuluL7_1(.din(w_dff_B_BePO5IXJ4_1),.dout(w_dff_B_5nJkuluL7_1),.clk(gclk));
	jdff dff_B_LOqAfdhc0_1(.din(w_dff_B_5nJkuluL7_1),.dout(w_dff_B_LOqAfdhc0_1),.clk(gclk));
	jdff dff_B_mc8q4U0a2_1(.din(w_dff_B_LOqAfdhc0_1),.dout(w_dff_B_mc8q4U0a2_1),.clk(gclk));
	jdff dff_B_oPu8Kb6S7_1(.din(w_dff_B_mc8q4U0a2_1),.dout(w_dff_B_oPu8Kb6S7_1),.clk(gclk));
	jdff dff_B_7C3ASDbp1_1(.din(w_dff_B_oPu8Kb6S7_1),.dout(w_dff_B_7C3ASDbp1_1),.clk(gclk));
	jdff dff_B_Yk31x2LH0_1(.din(w_dff_B_7C3ASDbp1_1),.dout(w_dff_B_Yk31x2LH0_1),.clk(gclk));
	jdff dff_B_k65tflB37_1(.din(w_dff_B_Yk31x2LH0_1),.dout(w_dff_B_k65tflB37_1),.clk(gclk));
	jdff dff_B_ufgvtTPv4_1(.din(w_dff_B_k65tflB37_1),.dout(w_dff_B_ufgvtTPv4_1),.clk(gclk));
	jdff dff_B_cifzNKpT5_1(.din(w_dff_B_ufgvtTPv4_1),.dout(w_dff_B_cifzNKpT5_1),.clk(gclk));
	jdff dff_B_xojATAs66_1(.din(w_dff_B_cifzNKpT5_1),.dout(w_dff_B_xojATAs66_1),.clk(gclk));
	jdff dff_B_2s4vnN7u1_1(.din(w_dff_B_xojATAs66_1),.dout(w_dff_B_2s4vnN7u1_1),.clk(gclk));
	jdff dff_B_3u3MEhQz3_1(.din(w_dff_B_2s4vnN7u1_1),.dout(w_dff_B_3u3MEhQz3_1),.clk(gclk));
	jdff dff_B_CrhhMABa3_1(.din(w_dff_B_3u3MEhQz3_1),.dout(w_dff_B_CrhhMABa3_1),.clk(gclk));
	jdff dff_B_6zXPqvjK6_1(.din(w_dff_B_CrhhMABa3_1),.dout(w_dff_B_6zXPqvjK6_1),.clk(gclk));
	jdff dff_B_ZvnD84cz9_1(.din(w_dff_B_6zXPqvjK6_1),.dout(w_dff_B_ZvnD84cz9_1),.clk(gclk));
	jdff dff_B_hFt9XGbI9_1(.din(w_dff_B_ZvnD84cz9_1),.dout(w_dff_B_hFt9XGbI9_1),.clk(gclk));
	jdff dff_B_I5dzgASW8_1(.din(w_dff_B_hFt9XGbI9_1),.dout(w_dff_B_I5dzgASW8_1),.clk(gclk));
	jdff dff_B_ap2KaO5W2_1(.din(w_dff_B_I5dzgASW8_1),.dout(w_dff_B_ap2KaO5W2_1),.clk(gclk));
	jdff dff_B_CWsNdAS21_1(.din(w_dff_B_ap2KaO5W2_1),.dout(w_dff_B_CWsNdAS21_1),.clk(gclk));
	jdff dff_B_w8Vn2nOt6_1(.din(w_dff_B_CWsNdAS21_1),.dout(w_dff_B_w8Vn2nOt6_1),.clk(gclk));
	jdff dff_B_jwcKYoSU1_1(.din(w_dff_B_w8Vn2nOt6_1),.dout(w_dff_B_jwcKYoSU1_1),.clk(gclk));
	jdff dff_B_40axs05m0_0(.din(n673),.dout(w_dff_B_40axs05m0_0),.clk(gclk));
	jdff dff_B_OffUMx7R8_0(.din(w_dff_B_40axs05m0_0),.dout(w_dff_B_OffUMx7R8_0),.clk(gclk));
	jdff dff_B_Q8B2xwor8_0(.din(w_dff_B_OffUMx7R8_0),.dout(w_dff_B_Q8B2xwor8_0),.clk(gclk));
	jdff dff_B_sGD3YZEY0_0(.din(w_dff_B_Q8B2xwor8_0),.dout(w_dff_B_sGD3YZEY0_0),.clk(gclk));
	jdff dff_B_kZ11lPUx2_0(.din(w_dff_B_sGD3YZEY0_0),.dout(w_dff_B_kZ11lPUx2_0),.clk(gclk));
	jdff dff_B_ISezBBuN8_0(.din(w_dff_B_kZ11lPUx2_0),.dout(w_dff_B_ISezBBuN8_0),.clk(gclk));
	jdff dff_B_taLFUeXC6_0(.din(w_dff_B_ISezBBuN8_0),.dout(w_dff_B_taLFUeXC6_0),.clk(gclk));
	jdff dff_B_IgyaCaAn1_0(.din(w_dff_B_taLFUeXC6_0),.dout(w_dff_B_IgyaCaAn1_0),.clk(gclk));
	jdff dff_B_XgiNsoNh7_0(.din(w_dff_B_IgyaCaAn1_0),.dout(w_dff_B_XgiNsoNh7_0),.clk(gclk));
	jdff dff_B_z3zWNLWx9_0(.din(w_dff_B_XgiNsoNh7_0),.dout(w_dff_B_z3zWNLWx9_0),.clk(gclk));
	jdff dff_B_CuBVRx4n9_0(.din(w_dff_B_z3zWNLWx9_0),.dout(w_dff_B_CuBVRx4n9_0),.clk(gclk));
	jdff dff_B_7Hc6tHMn0_0(.din(w_dff_B_CuBVRx4n9_0),.dout(w_dff_B_7Hc6tHMn0_0),.clk(gclk));
	jdff dff_B_IYDyJz1m5_0(.din(w_dff_B_7Hc6tHMn0_0),.dout(w_dff_B_IYDyJz1m5_0),.clk(gclk));
	jdff dff_B_fr9wnS0u6_0(.din(w_dff_B_IYDyJz1m5_0),.dout(w_dff_B_fr9wnS0u6_0),.clk(gclk));
	jdff dff_B_soMDuZBG4_0(.din(w_dff_B_fr9wnS0u6_0),.dout(w_dff_B_soMDuZBG4_0),.clk(gclk));
	jdff dff_B_h8BXpw9J3_0(.din(w_dff_B_soMDuZBG4_0),.dout(w_dff_B_h8BXpw9J3_0),.clk(gclk));
	jdff dff_B_RONKxCzt3_0(.din(w_dff_B_h8BXpw9J3_0),.dout(w_dff_B_RONKxCzt3_0),.clk(gclk));
	jdff dff_B_xpjWN0uD0_0(.din(w_dff_B_RONKxCzt3_0),.dout(w_dff_B_xpjWN0uD0_0),.clk(gclk));
	jdff dff_B_k0chVUju2_0(.din(w_dff_B_xpjWN0uD0_0),.dout(w_dff_B_k0chVUju2_0),.clk(gclk));
	jdff dff_B_aD44xSYH9_0(.din(w_dff_B_k0chVUju2_0),.dout(w_dff_B_aD44xSYH9_0),.clk(gclk));
	jdff dff_B_7hruGXbF7_0(.din(w_dff_B_aD44xSYH9_0),.dout(w_dff_B_7hruGXbF7_0),.clk(gclk));
	jdff dff_B_QZPvQEjj7_0(.din(w_dff_B_7hruGXbF7_0),.dout(w_dff_B_QZPvQEjj7_0),.clk(gclk));
	jdff dff_B_AGfo1Rsu2_0(.din(w_dff_B_QZPvQEjj7_0),.dout(w_dff_B_AGfo1Rsu2_0),.clk(gclk));
	jdff dff_B_d1aLTJp94_0(.din(w_dff_B_AGfo1Rsu2_0),.dout(w_dff_B_d1aLTJp94_0),.clk(gclk));
	jdff dff_B_fxd2ASEM6_0(.din(w_dff_B_d1aLTJp94_0),.dout(w_dff_B_fxd2ASEM6_0),.clk(gclk));
	jdff dff_B_8EJ4AQyt2_0(.din(w_dff_B_fxd2ASEM6_0),.dout(w_dff_B_8EJ4AQyt2_0),.clk(gclk));
	jdff dff_B_QVV9mnIC8_0(.din(w_dff_B_8EJ4AQyt2_0),.dout(w_dff_B_QVV9mnIC8_0),.clk(gclk));
	jdff dff_B_Buunm74Z4_0(.din(w_dff_B_QVV9mnIC8_0),.dout(w_dff_B_Buunm74Z4_0),.clk(gclk));
	jdff dff_B_CZLvVthy3_0(.din(w_dff_B_Buunm74Z4_0),.dout(w_dff_B_CZLvVthy3_0),.clk(gclk));
	jdff dff_B_uAu4QFrV7_0(.din(w_dff_B_CZLvVthy3_0),.dout(w_dff_B_uAu4QFrV7_0),.clk(gclk));
	jdff dff_B_36JBPEQP6_0(.din(w_dff_B_uAu4QFrV7_0),.dout(w_dff_B_36JBPEQP6_0),.clk(gclk));
	jdff dff_B_gpGrFkiB2_0(.din(w_dff_B_36JBPEQP6_0),.dout(w_dff_B_gpGrFkiB2_0),.clk(gclk));
	jdff dff_B_JE3xncqI2_0(.din(w_dff_B_gpGrFkiB2_0),.dout(w_dff_B_JE3xncqI2_0),.clk(gclk));
	jdff dff_B_lA9ksrmU5_0(.din(w_dff_B_JE3xncqI2_0),.dout(w_dff_B_lA9ksrmU5_0),.clk(gclk));
	jdff dff_B_rgWBQvSp3_0(.din(w_dff_B_lA9ksrmU5_0),.dout(w_dff_B_rgWBQvSp3_0),.clk(gclk));
	jdff dff_B_cH9MFqUT0_0(.din(w_dff_B_rgWBQvSp3_0),.dout(w_dff_B_cH9MFqUT0_0),.clk(gclk));
	jdff dff_B_ERfPkje79_0(.din(w_dff_B_cH9MFqUT0_0),.dout(w_dff_B_ERfPkje79_0),.clk(gclk));
	jdff dff_B_SzbEFIL33_0(.din(w_dff_B_ERfPkje79_0),.dout(w_dff_B_SzbEFIL33_0),.clk(gclk));
	jdff dff_B_z8ogwEuY9_0(.din(w_dff_B_SzbEFIL33_0),.dout(w_dff_B_z8ogwEuY9_0),.clk(gclk));
	jdff dff_B_xHe58wJT7_0(.din(w_dff_B_z8ogwEuY9_0),.dout(w_dff_B_xHe58wJT7_0),.clk(gclk));
	jdff dff_B_35IDh1Zl0_0(.din(w_dff_B_xHe58wJT7_0),.dout(w_dff_B_35IDh1Zl0_0),.clk(gclk));
	jdff dff_B_h8D3TgeQ2_0(.din(w_dff_B_35IDh1Zl0_0),.dout(w_dff_B_h8D3TgeQ2_0),.clk(gclk));
	jdff dff_B_i1O2QFby3_0(.din(w_dff_B_h8D3TgeQ2_0),.dout(w_dff_B_i1O2QFby3_0),.clk(gclk));
	jdff dff_B_dM1kPNpR2_0(.din(w_dff_B_i1O2QFby3_0),.dout(w_dff_B_dM1kPNpR2_0),.clk(gclk));
	jdff dff_B_uDBbSCPA7_0(.din(w_dff_B_dM1kPNpR2_0),.dout(w_dff_B_uDBbSCPA7_0),.clk(gclk));
	jdff dff_B_ms9K776m3_0(.din(w_dff_B_uDBbSCPA7_0),.dout(w_dff_B_ms9K776m3_0),.clk(gclk));
	jdff dff_B_VLbvT5nE1_0(.din(w_dff_B_ms9K776m3_0),.dout(w_dff_B_VLbvT5nE1_0),.clk(gclk));
	jdff dff_B_YAxWtq8t8_0(.din(w_dff_B_VLbvT5nE1_0),.dout(w_dff_B_YAxWtq8t8_0),.clk(gclk));
	jdff dff_B_vvWIz1QP5_1(.din(n666),.dout(w_dff_B_vvWIz1QP5_1),.clk(gclk));
	jdff dff_B_x6ed2YVm7_1(.din(w_dff_B_vvWIz1QP5_1),.dout(w_dff_B_x6ed2YVm7_1),.clk(gclk));
	jdff dff_B_vhBEouJ16_1(.din(w_dff_B_x6ed2YVm7_1),.dout(w_dff_B_vhBEouJ16_1),.clk(gclk));
	jdff dff_B_JOnOab7Y5_1(.din(w_dff_B_vhBEouJ16_1),.dout(w_dff_B_JOnOab7Y5_1),.clk(gclk));
	jdff dff_B_H8TNWflg5_1(.din(w_dff_B_JOnOab7Y5_1),.dout(w_dff_B_H8TNWflg5_1),.clk(gclk));
	jdff dff_B_rYuSiGpX3_1(.din(w_dff_B_H8TNWflg5_1),.dout(w_dff_B_rYuSiGpX3_1),.clk(gclk));
	jdff dff_B_PjNOFRsW3_1(.din(w_dff_B_rYuSiGpX3_1),.dout(w_dff_B_PjNOFRsW3_1),.clk(gclk));
	jdff dff_B_yzUMUqn91_1(.din(w_dff_B_PjNOFRsW3_1),.dout(w_dff_B_yzUMUqn91_1),.clk(gclk));
	jdff dff_B_MPCpsYqI3_1(.din(w_dff_B_yzUMUqn91_1),.dout(w_dff_B_MPCpsYqI3_1),.clk(gclk));
	jdff dff_B_NU2sOvR51_1(.din(w_dff_B_MPCpsYqI3_1),.dout(w_dff_B_NU2sOvR51_1),.clk(gclk));
	jdff dff_B_CKTlIbPr3_1(.din(w_dff_B_NU2sOvR51_1),.dout(w_dff_B_CKTlIbPr3_1),.clk(gclk));
	jdff dff_B_2Cj7x41M4_1(.din(w_dff_B_CKTlIbPr3_1),.dout(w_dff_B_2Cj7x41M4_1),.clk(gclk));
	jdff dff_B_FG7SWVwj6_1(.din(w_dff_B_2Cj7x41M4_1),.dout(w_dff_B_FG7SWVwj6_1),.clk(gclk));
	jdff dff_B_rR0cphWL9_1(.din(w_dff_B_FG7SWVwj6_1),.dout(w_dff_B_rR0cphWL9_1),.clk(gclk));
	jdff dff_B_1h989HLm3_1(.din(w_dff_B_rR0cphWL9_1),.dout(w_dff_B_1h989HLm3_1),.clk(gclk));
	jdff dff_B_QuJVjKsV6_1(.din(w_dff_B_1h989HLm3_1),.dout(w_dff_B_QuJVjKsV6_1),.clk(gclk));
	jdff dff_B_IKAiJwAl0_1(.din(w_dff_B_QuJVjKsV6_1),.dout(w_dff_B_IKAiJwAl0_1),.clk(gclk));
	jdff dff_B_WtPJZocd1_1(.din(w_dff_B_IKAiJwAl0_1),.dout(w_dff_B_WtPJZocd1_1),.clk(gclk));
	jdff dff_B_QAdpB0jX0_1(.din(w_dff_B_WtPJZocd1_1),.dout(w_dff_B_QAdpB0jX0_1),.clk(gclk));
	jdff dff_B_1Px8bGZx0_1(.din(w_dff_B_QAdpB0jX0_1),.dout(w_dff_B_1Px8bGZx0_1),.clk(gclk));
	jdff dff_B_vRPiREMc6_1(.din(w_dff_B_1Px8bGZx0_1),.dout(w_dff_B_vRPiREMc6_1),.clk(gclk));
	jdff dff_B_kBMyCMHf2_1(.din(w_dff_B_vRPiREMc6_1),.dout(w_dff_B_kBMyCMHf2_1),.clk(gclk));
	jdff dff_B_8Ezv7QT95_1(.din(w_dff_B_kBMyCMHf2_1),.dout(w_dff_B_8Ezv7QT95_1),.clk(gclk));
	jdff dff_B_sBBygfT39_1(.din(w_dff_B_8Ezv7QT95_1),.dout(w_dff_B_sBBygfT39_1),.clk(gclk));
	jdff dff_B_GW2KJw0R7_1(.din(w_dff_B_sBBygfT39_1),.dout(w_dff_B_GW2KJw0R7_1),.clk(gclk));
	jdff dff_B_jGursqEB5_1(.din(w_dff_B_GW2KJw0R7_1),.dout(w_dff_B_jGursqEB5_1),.clk(gclk));
	jdff dff_B_PQpomRoH7_1(.din(w_dff_B_jGursqEB5_1),.dout(w_dff_B_PQpomRoH7_1),.clk(gclk));
	jdff dff_B_Ge2ue2aj0_1(.din(w_dff_B_PQpomRoH7_1),.dout(w_dff_B_Ge2ue2aj0_1),.clk(gclk));
	jdff dff_B_p1WsVsb60_1(.din(w_dff_B_Ge2ue2aj0_1),.dout(w_dff_B_p1WsVsb60_1),.clk(gclk));
	jdff dff_B_ZNo9H01j1_1(.din(w_dff_B_p1WsVsb60_1),.dout(w_dff_B_ZNo9H01j1_1),.clk(gclk));
	jdff dff_B_Ty8hcaE66_1(.din(w_dff_B_ZNo9H01j1_1),.dout(w_dff_B_Ty8hcaE66_1),.clk(gclk));
	jdff dff_B_FZGIMHUy7_1(.din(w_dff_B_Ty8hcaE66_1),.dout(w_dff_B_FZGIMHUy7_1),.clk(gclk));
	jdff dff_B_qA0QAqjM5_1(.din(w_dff_B_FZGIMHUy7_1),.dout(w_dff_B_qA0QAqjM5_1),.clk(gclk));
	jdff dff_B_FHvAcDl31_1(.din(w_dff_B_qA0QAqjM5_1),.dout(w_dff_B_FHvAcDl31_1),.clk(gclk));
	jdff dff_B_0gOv2HX11_1(.din(w_dff_B_FHvAcDl31_1),.dout(w_dff_B_0gOv2HX11_1),.clk(gclk));
	jdff dff_B_l8qcYsiU9_1(.din(w_dff_B_0gOv2HX11_1),.dout(w_dff_B_l8qcYsiU9_1),.clk(gclk));
	jdff dff_B_WIxcTGWV3_1(.din(w_dff_B_l8qcYsiU9_1),.dout(w_dff_B_WIxcTGWV3_1),.clk(gclk));
	jdff dff_B_SKbqsVY74_1(.din(w_dff_B_WIxcTGWV3_1),.dout(w_dff_B_SKbqsVY74_1),.clk(gclk));
	jdff dff_B_GCQuWFux6_1(.din(w_dff_B_SKbqsVY74_1),.dout(w_dff_B_GCQuWFux6_1),.clk(gclk));
	jdff dff_B_x5IXtwpv7_1(.din(w_dff_B_GCQuWFux6_1),.dout(w_dff_B_x5IXtwpv7_1),.clk(gclk));
	jdff dff_B_2yyDiDP56_1(.din(w_dff_B_x5IXtwpv7_1),.dout(w_dff_B_2yyDiDP56_1),.clk(gclk));
	jdff dff_B_GsfZAp0v5_1(.din(w_dff_B_2yyDiDP56_1),.dout(w_dff_B_GsfZAp0v5_1),.clk(gclk));
	jdff dff_B_8Ynj0uPy0_1(.din(w_dff_B_GsfZAp0v5_1),.dout(w_dff_B_8Ynj0uPy0_1),.clk(gclk));
	jdff dff_B_2FLoPUoD0_1(.din(w_dff_B_8Ynj0uPy0_1),.dout(w_dff_B_2FLoPUoD0_1),.clk(gclk));
	jdff dff_B_RieSgn2L4_1(.din(w_dff_B_2FLoPUoD0_1),.dout(w_dff_B_RieSgn2L4_1),.clk(gclk));
	jdff dff_B_jyOn7VFb8_1(.din(w_dff_B_RieSgn2L4_1),.dout(w_dff_B_jyOn7VFb8_1),.clk(gclk));
	jdff dff_B_HGuNeMUK0_1(.din(w_dff_B_jyOn7VFb8_1),.dout(w_dff_B_HGuNeMUK0_1),.clk(gclk));
	jdff dff_B_X5L2oJc08_0(.din(n667),.dout(w_dff_B_X5L2oJc08_0),.clk(gclk));
	jdff dff_B_hsMdZii72_0(.din(w_dff_B_X5L2oJc08_0),.dout(w_dff_B_hsMdZii72_0),.clk(gclk));
	jdff dff_B_sFIILIqp7_0(.din(w_dff_B_hsMdZii72_0),.dout(w_dff_B_sFIILIqp7_0),.clk(gclk));
	jdff dff_B_KqsKhx3Y1_0(.din(w_dff_B_sFIILIqp7_0),.dout(w_dff_B_KqsKhx3Y1_0),.clk(gclk));
	jdff dff_B_uJogh1Xe0_0(.din(w_dff_B_KqsKhx3Y1_0),.dout(w_dff_B_uJogh1Xe0_0),.clk(gclk));
	jdff dff_B_wS9chUuM1_0(.din(w_dff_B_uJogh1Xe0_0),.dout(w_dff_B_wS9chUuM1_0),.clk(gclk));
	jdff dff_B_rPv7w3865_0(.din(w_dff_B_wS9chUuM1_0),.dout(w_dff_B_rPv7w3865_0),.clk(gclk));
	jdff dff_B_8KAfykP25_0(.din(w_dff_B_rPv7w3865_0),.dout(w_dff_B_8KAfykP25_0),.clk(gclk));
	jdff dff_B_NOPEF98n0_0(.din(w_dff_B_8KAfykP25_0),.dout(w_dff_B_NOPEF98n0_0),.clk(gclk));
	jdff dff_B_sH6WML8f9_0(.din(w_dff_B_NOPEF98n0_0),.dout(w_dff_B_sH6WML8f9_0),.clk(gclk));
	jdff dff_B_wWCohYwY7_0(.din(w_dff_B_sH6WML8f9_0),.dout(w_dff_B_wWCohYwY7_0),.clk(gclk));
	jdff dff_B_4KyL94eA2_0(.din(w_dff_B_wWCohYwY7_0),.dout(w_dff_B_4KyL94eA2_0),.clk(gclk));
	jdff dff_B_ayAxIPLi7_0(.din(w_dff_B_4KyL94eA2_0),.dout(w_dff_B_ayAxIPLi7_0),.clk(gclk));
	jdff dff_B_S1d0e5Lm2_0(.din(w_dff_B_ayAxIPLi7_0),.dout(w_dff_B_S1d0e5Lm2_0),.clk(gclk));
	jdff dff_B_SxZayiWL5_0(.din(w_dff_B_S1d0e5Lm2_0),.dout(w_dff_B_SxZayiWL5_0),.clk(gclk));
	jdff dff_B_cC3Lp0en3_0(.din(w_dff_B_SxZayiWL5_0),.dout(w_dff_B_cC3Lp0en3_0),.clk(gclk));
	jdff dff_B_YIIPcC1A9_0(.din(w_dff_B_cC3Lp0en3_0),.dout(w_dff_B_YIIPcC1A9_0),.clk(gclk));
	jdff dff_B_A4xCihqY4_0(.din(w_dff_B_YIIPcC1A9_0),.dout(w_dff_B_A4xCihqY4_0),.clk(gclk));
	jdff dff_B_3xONO7RM1_0(.din(w_dff_B_A4xCihqY4_0),.dout(w_dff_B_3xONO7RM1_0),.clk(gclk));
	jdff dff_B_Xepa6ujA6_0(.din(w_dff_B_3xONO7RM1_0),.dout(w_dff_B_Xepa6ujA6_0),.clk(gclk));
	jdff dff_B_LkWWh7pG9_0(.din(w_dff_B_Xepa6ujA6_0),.dout(w_dff_B_LkWWh7pG9_0),.clk(gclk));
	jdff dff_B_hr4JckW02_0(.din(w_dff_B_LkWWh7pG9_0),.dout(w_dff_B_hr4JckW02_0),.clk(gclk));
	jdff dff_B_yxJkppAV7_0(.din(w_dff_B_hr4JckW02_0),.dout(w_dff_B_yxJkppAV7_0),.clk(gclk));
	jdff dff_B_t4NlzVy80_0(.din(w_dff_B_yxJkppAV7_0),.dout(w_dff_B_t4NlzVy80_0),.clk(gclk));
	jdff dff_B_XRwplYNf4_0(.din(w_dff_B_t4NlzVy80_0),.dout(w_dff_B_XRwplYNf4_0),.clk(gclk));
	jdff dff_B_7mztHKZu6_0(.din(w_dff_B_XRwplYNf4_0),.dout(w_dff_B_7mztHKZu6_0),.clk(gclk));
	jdff dff_B_5AhiBGHR0_0(.din(w_dff_B_7mztHKZu6_0),.dout(w_dff_B_5AhiBGHR0_0),.clk(gclk));
	jdff dff_B_9G4rxd8p1_0(.din(w_dff_B_5AhiBGHR0_0),.dout(w_dff_B_9G4rxd8p1_0),.clk(gclk));
	jdff dff_B_sVtwLxFP0_0(.din(w_dff_B_9G4rxd8p1_0),.dout(w_dff_B_sVtwLxFP0_0),.clk(gclk));
	jdff dff_B_6uOiN1TZ0_0(.din(w_dff_B_sVtwLxFP0_0),.dout(w_dff_B_6uOiN1TZ0_0),.clk(gclk));
	jdff dff_B_23IPDeYb4_0(.din(w_dff_B_6uOiN1TZ0_0),.dout(w_dff_B_23IPDeYb4_0),.clk(gclk));
	jdff dff_B_8O8qpHJS1_0(.din(w_dff_B_23IPDeYb4_0),.dout(w_dff_B_8O8qpHJS1_0),.clk(gclk));
	jdff dff_B_GM8Q3bDK6_0(.din(w_dff_B_8O8qpHJS1_0),.dout(w_dff_B_GM8Q3bDK6_0),.clk(gclk));
	jdff dff_B_0RpHrqHE3_0(.din(w_dff_B_GM8Q3bDK6_0),.dout(w_dff_B_0RpHrqHE3_0),.clk(gclk));
	jdff dff_B_V7TIGBT59_0(.din(w_dff_B_0RpHrqHE3_0),.dout(w_dff_B_V7TIGBT59_0),.clk(gclk));
	jdff dff_B_2D6U3nw51_0(.din(w_dff_B_V7TIGBT59_0),.dout(w_dff_B_2D6U3nw51_0),.clk(gclk));
	jdff dff_B_Xp7snU9d4_0(.din(w_dff_B_2D6U3nw51_0),.dout(w_dff_B_Xp7snU9d4_0),.clk(gclk));
	jdff dff_B_so8Tqb4r7_0(.din(w_dff_B_Xp7snU9d4_0),.dout(w_dff_B_so8Tqb4r7_0),.clk(gclk));
	jdff dff_B_Maa3dE9Q0_0(.din(w_dff_B_so8Tqb4r7_0),.dout(w_dff_B_Maa3dE9Q0_0),.clk(gclk));
	jdff dff_B_u8uo5R6K2_0(.din(w_dff_B_Maa3dE9Q0_0),.dout(w_dff_B_u8uo5R6K2_0),.clk(gclk));
	jdff dff_B_RApRDQZK1_0(.din(w_dff_B_u8uo5R6K2_0),.dout(w_dff_B_RApRDQZK1_0),.clk(gclk));
	jdff dff_B_Kn0gZBDs8_0(.din(w_dff_B_RApRDQZK1_0),.dout(w_dff_B_Kn0gZBDs8_0),.clk(gclk));
	jdff dff_B_kizdjsid5_0(.din(w_dff_B_Kn0gZBDs8_0),.dout(w_dff_B_kizdjsid5_0),.clk(gclk));
	jdff dff_B_IgXKponO7_0(.din(w_dff_B_kizdjsid5_0),.dout(w_dff_B_IgXKponO7_0),.clk(gclk));
	jdff dff_B_YoVBKepe5_0(.din(w_dff_B_IgXKponO7_0),.dout(w_dff_B_YoVBKepe5_0),.clk(gclk));
	jdff dff_B_7FHPGv6J7_0(.din(w_dff_B_YoVBKepe5_0),.dout(w_dff_B_7FHPGv6J7_0),.clk(gclk));
	jdff dff_B_dL6uwy6j5_0(.din(w_dff_B_7FHPGv6J7_0),.dout(w_dff_B_dL6uwy6j5_0),.clk(gclk));
	jdff dff_B_RareMZ3a0_1(.din(n660),.dout(w_dff_B_RareMZ3a0_1),.clk(gclk));
	jdff dff_B_yF59gkoW3_1(.din(w_dff_B_RareMZ3a0_1),.dout(w_dff_B_yF59gkoW3_1),.clk(gclk));
	jdff dff_B_tBiJ8S9k1_1(.din(w_dff_B_yF59gkoW3_1),.dout(w_dff_B_tBiJ8S9k1_1),.clk(gclk));
	jdff dff_B_jLAeV3cH0_1(.din(w_dff_B_tBiJ8S9k1_1),.dout(w_dff_B_jLAeV3cH0_1),.clk(gclk));
	jdff dff_B_3wzp0HUu3_1(.din(w_dff_B_jLAeV3cH0_1),.dout(w_dff_B_3wzp0HUu3_1),.clk(gclk));
	jdff dff_B_CrgpEJ4p0_1(.din(w_dff_B_3wzp0HUu3_1),.dout(w_dff_B_CrgpEJ4p0_1),.clk(gclk));
	jdff dff_B_6Ja2co3F4_1(.din(w_dff_B_CrgpEJ4p0_1),.dout(w_dff_B_6Ja2co3F4_1),.clk(gclk));
	jdff dff_B_59DVj8Js9_1(.din(w_dff_B_6Ja2co3F4_1),.dout(w_dff_B_59DVj8Js9_1),.clk(gclk));
	jdff dff_B_bJyV7eUw5_1(.din(w_dff_B_59DVj8Js9_1),.dout(w_dff_B_bJyV7eUw5_1),.clk(gclk));
	jdff dff_B_3OZ1ouUr1_1(.din(w_dff_B_bJyV7eUw5_1),.dout(w_dff_B_3OZ1ouUr1_1),.clk(gclk));
	jdff dff_B_bYOqyUOC4_1(.din(w_dff_B_3OZ1ouUr1_1),.dout(w_dff_B_bYOqyUOC4_1),.clk(gclk));
	jdff dff_B_BNbpJa2r6_1(.din(w_dff_B_bYOqyUOC4_1),.dout(w_dff_B_BNbpJa2r6_1),.clk(gclk));
	jdff dff_B_gHbPwMYe9_1(.din(w_dff_B_BNbpJa2r6_1),.dout(w_dff_B_gHbPwMYe9_1),.clk(gclk));
	jdff dff_B_6gQnOMtJ9_1(.din(w_dff_B_gHbPwMYe9_1),.dout(w_dff_B_6gQnOMtJ9_1),.clk(gclk));
	jdff dff_B_HEfMyAge5_1(.din(w_dff_B_6gQnOMtJ9_1),.dout(w_dff_B_HEfMyAge5_1),.clk(gclk));
	jdff dff_B_gbJFsDfJ5_1(.din(w_dff_B_HEfMyAge5_1),.dout(w_dff_B_gbJFsDfJ5_1),.clk(gclk));
	jdff dff_B_40aohpb96_1(.din(w_dff_B_gbJFsDfJ5_1),.dout(w_dff_B_40aohpb96_1),.clk(gclk));
	jdff dff_B_IZQeTgDk9_1(.din(w_dff_B_40aohpb96_1),.dout(w_dff_B_IZQeTgDk9_1),.clk(gclk));
	jdff dff_B_FBiPRHqU8_1(.din(w_dff_B_IZQeTgDk9_1),.dout(w_dff_B_FBiPRHqU8_1),.clk(gclk));
	jdff dff_B_diTHVDpi4_1(.din(w_dff_B_FBiPRHqU8_1),.dout(w_dff_B_diTHVDpi4_1),.clk(gclk));
	jdff dff_B_vKbaXYpi3_1(.din(w_dff_B_diTHVDpi4_1),.dout(w_dff_B_vKbaXYpi3_1),.clk(gclk));
	jdff dff_B_cg8SRKwx1_1(.din(w_dff_B_vKbaXYpi3_1),.dout(w_dff_B_cg8SRKwx1_1),.clk(gclk));
	jdff dff_B_VRL8Nveg9_1(.din(w_dff_B_cg8SRKwx1_1),.dout(w_dff_B_VRL8Nveg9_1),.clk(gclk));
	jdff dff_B_SUNP9bmW7_1(.din(w_dff_B_VRL8Nveg9_1),.dout(w_dff_B_SUNP9bmW7_1),.clk(gclk));
	jdff dff_B_UCtUPBnI0_1(.din(w_dff_B_SUNP9bmW7_1),.dout(w_dff_B_UCtUPBnI0_1),.clk(gclk));
	jdff dff_B_UfQaruGv7_1(.din(w_dff_B_UCtUPBnI0_1),.dout(w_dff_B_UfQaruGv7_1),.clk(gclk));
	jdff dff_B_LkXJbTM55_1(.din(w_dff_B_UfQaruGv7_1),.dout(w_dff_B_LkXJbTM55_1),.clk(gclk));
	jdff dff_B_JFCnja7Y7_1(.din(w_dff_B_LkXJbTM55_1),.dout(w_dff_B_JFCnja7Y7_1),.clk(gclk));
	jdff dff_B_WeVK8C5h8_1(.din(w_dff_B_JFCnja7Y7_1),.dout(w_dff_B_WeVK8C5h8_1),.clk(gclk));
	jdff dff_B_lAsJRaTI5_1(.din(w_dff_B_WeVK8C5h8_1),.dout(w_dff_B_lAsJRaTI5_1),.clk(gclk));
	jdff dff_B_12mobeAb1_1(.din(w_dff_B_lAsJRaTI5_1),.dout(w_dff_B_12mobeAb1_1),.clk(gclk));
	jdff dff_B_zbkT3Di76_1(.din(w_dff_B_12mobeAb1_1),.dout(w_dff_B_zbkT3Di76_1),.clk(gclk));
	jdff dff_B_CRcalJ793_1(.din(w_dff_B_zbkT3Di76_1),.dout(w_dff_B_CRcalJ793_1),.clk(gclk));
	jdff dff_B_7eNX7ec42_1(.din(w_dff_B_CRcalJ793_1),.dout(w_dff_B_7eNX7ec42_1),.clk(gclk));
	jdff dff_B_lIez84FE3_1(.din(w_dff_B_7eNX7ec42_1),.dout(w_dff_B_lIez84FE3_1),.clk(gclk));
	jdff dff_B_P4nF0UWT6_1(.din(w_dff_B_lIez84FE3_1),.dout(w_dff_B_P4nF0UWT6_1),.clk(gclk));
	jdff dff_B_W62ryUpn4_1(.din(w_dff_B_P4nF0UWT6_1),.dout(w_dff_B_W62ryUpn4_1),.clk(gclk));
	jdff dff_B_mHjw1S9M1_1(.din(w_dff_B_W62ryUpn4_1),.dout(w_dff_B_mHjw1S9M1_1),.clk(gclk));
	jdff dff_B_oMqc1zsx4_1(.din(w_dff_B_mHjw1S9M1_1),.dout(w_dff_B_oMqc1zsx4_1),.clk(gclk));
	jdff dff_B_0Nh5DdFJ8_1(.din(w_dff_B_oMqc1zsx4_1),.dout(w_dff_B_0Nh5DdFJ8_1),.clk(gclk));
	jdff dff_B_aIL6VXuh6_1(.din(w_dff_B_0Nh5DdFJ8_1),.dout(w_dff_B_aIL6VXuh6_1),.clk(gclk));
	jdff dff_B_lmVL6hjy9_1(.din(w_dff_B_aIL6VXuh6_1),.dout(w_dff_B_lmVL6hjy9_1),.clk(gclk));
	jdff dff_B_gSQlFaGW5_1(.din(w_dff_B_lmVL6hjy9_1),.dout(w_dff_B_gSQlFaGW5_1),.clk(gclk));
	jdff dff_B_2fXr4ntQ1_1(.din(w_dff_B_gSQlFaGW5_1),.dout(w_dff_B_2fXr4ntQ1_1),.clk(gclk));
	jdff dff_B_dT5YuAQX7_1(.din(w_dff_B_2fXr4ntQ1_1),.dout(w_dff_B_dT5YuAQX7_1),.clk(gclk));
	jdff dff_B_ka8N4w5F3_1(.din(w_dff_B_dT5YuAQX7_1),.dout(w_dff_B_ka8N4w5F3_1),.clk(gclk));
	jdff dff_B_aBsTRinM6_0(.din(n661),.dout(w_dff_B_aBsTRinM6_0),.clk(gclk));
	jdff dff_B_4EqVSWda4_0(.din(w_dff_B_aBsTRinM6_0),.dout(w_dff_B_4EqVSWda4_0),.clk(gclk));
	jdff dff_B_yOsaRBXF0_0(.din(w_dff_B_4EqVSWda4_0),.dout(w_dff_B_yOsaRBXF0_0),.clk(gclk));
	jdff dff_B_Xj56PTnV0_0(.din(w_dff_B_yOsaRBXF0_0),.dout(w_dff_B_Xj56PTnV0_0),.clk(gclk));
	jdff dff_B_PXMx5Mmx9_0(.din(w_dff_B_Xj56PTnV0_0),.dout(w_dff_B_PXMx5Mmx9_0),.clk(gclk));
	jdff dff_B_xNgy5rF84_0(.din(w_dff_B_PXMx5Mmx9_0),.dout(w_dff_B_xNgy5rF84_0),.clk(gclk));
	jdff dff_B_8Ci4NS0g4_0(.din(w_dff_B_xNgy5rF84_0),.dout(w_dff_B_8Ci4NS0g4_0),.clk(gclk));
	jdff dff_B_9YgRv75p1_0(.din(w_dff_B_8Ci4NS0g4_0),.dout(w_dff_B_9YgRv75p1_0),.clk(gclk));
	jdff dff_B_OACoJPxt3_0(.din(w_dff_B_9YgRv75p1_0),.dout(w_dff_B_OACoJPxt3_0),.clk(gclk));
	jdff dff_B_TRn10SlH3_0(.din(w_dff_B_OACoJPxt3_0),.dout(w_dff_B_TRn10SlH3_0),.clk(gclk));
	jdff dff_B_icnd60Cb2_0(.din(w_dff_B_TRn10SlH3_0),.dout(w_dff_B_icnd60Cb2_0),.clk(gclk));
	jdff dff_B_0FwPjB7W8_0(.din(w_dff_B_icnd60Cb2_0),.dout(w_dff_B_0FwPjB7W8_0),.clk(gclk));
	jdff dff_B_vryRiryW3_0(.din(w_dff_B_0FwPjB7W8_0),.dout(w_dff_B_vryRiryW3_0),.clk(gclk));
	jdff dff_B_ZK0JBD3a4_0(.din(w_dff_B_vryRiryW3_0),.dout(w_dff_B_ZK0JBD3a4_0),.clk(gclk));
	jdff dff_B_e7eddv003_0(.din(w_dff_B_ZK0JBD3a4_0),.dout(w_dff_B_e7eddv003_0),.clk(gclk));
	jdff dff_B_FjTq0QQM7_0(.din(w_dff_B_e7eddv003_0),.dout(w_dff_B_FjTq0QQM7_0),.clk(gclk));
	jdff dff_B_IdUpPekU8_0(.din(w_dff_B_FjTq0QQM7_0),.dout(w_dff_B_IdUpPekU8_0),.clk(gclk));
	jdff dff_B_dOBM42Mt6_0(.din(w_dff_B_IdUpPekU8_0),.dout(w_dff_B_dOBM42Mt6_0),.clk(gclk));
	jdff dff_B_XjpTKGfm1_0(.din(w_dff_B_dOBM42Mt6_0),.dout(w_dff_B_XjpTKGfm1_0),.clk(gclk));
	jdff dff_B_yfMw7pnX1_0(.din(w_dff_B_XjpTKGfm1_0),.dout(w_dff_B_yfMw7pnX1_0),.clk(gclk));
	jdff dff_B_O6QePwCH2_0(.din(w_dff_B_yfMw7pnX1_0),.dout(w_dff_B_O6QePwCH2_0),.clk(gclk));
	jdff dff_B_zrIknAPE4_0(.din(w_dff_B_O6QePwCH2_0),.dout(w_dff_B_zrIknAPE4_0),.clk(gclk));
	jdff dff_B_kHdafHAP4_0(.din(w_dff_B_zrIknAPE4_0),.dout(w_dff_B_kHdafHAP4_0),.clk(gclk));
	jdff dff_B_8zBUV71a6_0(.din(w_dff_B_kHdafHAP4_0),.dout(w_dff_B_8zBUV71a6_0),.clk(gclk));
	jdff dff_B_wfWOYZJ37_0(.din(w_dff_B_8zBUV71a6_0),.dout(w_dff_B_wfWOYZJ37_0),.clk(gclk));
	jdff dff_B_KNhaQbf18_0(.din(w_dff_B_wfWOYZJ37_0),.dout(w_dff_B_KNhaQbf18_0),.clk(gclk));
	jdff dff_B_O3YF9qtD9_0(.din(w_dff_B_KNhaQbf18_0),.dout(w_dff_B_O3YF9qtD9_0),.clk(gclk));
	jdff dff_B_oP3PMArx1_0(.din(w_dff_B_O3YF9qtD9_0),.dout(w_dff_B_oP3PMArx1_0),.clk(gclk));
	jdff dff_B_ycfeH6QV9_0(.din(w_dff_B_oP3PMArx1_0),.dout(w_dff_B_ycfeH6QV9_0),.clk(gclk));
	jdff dff_B_zdHLg6hv5_0(.din(w_dff_B_ycfeH6QV9_0),.dout(w_dff_B_zdHLg6hv5_0),.clk(gclk));
	jdff dff_B_UmV4s7tZ3_0(.din(w_dff_B_zdHLg6hv5_0),.dout(w_dff_B_UmV4s7tZ3_0),.clk(gclk));
	jdff dff_B_1HiDBbvd4_0(.din(w_dff_B_UmV4s7tZ3_0),.dout(w_dff_B_1HiDBbvd4_0),.clk(gclk));
	jdff dff_B_JZZIy4KT8_0(.din(w_dff_B_1HiDBbvd4_0),.dout(w_dff_B_JZZIy4KT8_0),.clk(gclk));
	jdff dff_B_fjntXGqZ9_0(.din(w_dff_B_JZZIy4KT8_0),.dout(w_dff_B_fjntXGqZ9_0),.clk(gclk));
	jdff dff_B_vBqpgiy78_0(.din(w_dff_B_fjntXGqZ9_0),.dout(w_dff_B_vBqpgiy78_0),.clk(gclk));
	jdff dff_B_dW4CplXG6_0(.din(w_dff_B_vBqpgiy78_0),.dout(w_dff_B_dW4CplXG6_0),.clk(gclk));
	jdff dff_B_VASnbmaW8_0(.din(w_dff_B_dW4CplXG6_0),.dout(w_dff_B_VASnbmaW8_0),.clk(gclk));
	jdff dff_B_FGMHauze8_0(.din(w_dff_B_VASnbmaW8_0),.dout(w_dff_B_FGMHauze8_0),.clk(gclk));
	jdff dff_B_48aUyuVU1_0(.din(w_dff_B_FGMHauze8_0),.dout(w_dff_B_48aUyuVU1_0),.clk(gclk));
	jdff dff_B_JyRHmNJl6_0(.din(w_dff_B_48aUyuVU1_0),.dout(w_dff_B_JyRHmNJl6_0),.clk(gclk));
	jdff dff_B_60oyD4mx1_0(.din(w_dff_B_JyRHmNJl6_0),.dout(w_dff_B_60oyD4mx1_0),.clk(gclk));
	jdff dff_B_UcLgOXrH5_0(.din(w_dff_B_60oyD4mx1_0),.dout(w_dff_B_UcLgOXrH5_0),.clk(gclk));
	jdff dff_B_SxEj46qu5_0(.din(w_dff_B_UcLgOXrH5_0),.dout(w_dff_B_SxEj46qu5_0),.clk(gclk));
	jdff dff_B_6cpYQZsk3_0(.din(w_dff_B_SxEj46qu5_0),.dout(w_dff_B_6cpYQZsk3_0),.clk(gclk));
	jdff dff_B_8LNWvVGh4_0(.din(w_dff_B_6cpYQZsk3_0),.dout(w_dff_B_8LNWvVGh4_0),.clk(gclk));
	jdff dff_B_ZUFZvbyO9_0(.din(w_dff_B_8LNWvVGh4_0),.dout(w_dff_B_ZUFZvbyO9_0),.clk(gclk));
	jdff dff_B_BfJV4Ur19_1(.din(n654),.dout(w_dff_B_BfJV4Ur19_1),.clk(gclk));
	jdff dff_B_xjnpz65V7_1(.din(w_dff_B_BfJV4Ur19_1),.dout(w_dff_B_xjnpz65V7_1),.clk(gclk));
	jdff dff_B_4u32G6LM7_1(.din(w_dff_B_xjnpz65V7_1),.dout(w_dff_B_4u32G6LM7_1),.clk(gclk));
	jdff dff_B_PhsnOrBz1_1(.din(w_dff_B_4u32G6LM7_1),.dout(w_dff_B_PhsnOrBz1_1),.clk(gclk));
	jdff dff_B_n3k8eKwb9_1(.din(w_dff_B_PhsnOrBz1_1),.dout(w_dff_B_n3k8eKwb9_1),.clk(gclk));
	jdff dff_B_Bhppne3H4_1(.din(w_dff_B_n3k8eKwb9_1),.dout(w_dff_B_Bhppne3H4_1),.clk(gclk));
	jdff dff_B_BHZXVDlh5_1(.din(w_dff_B_Bhppne3H4_1),.dout(w_dff_B_BHZXVDlh5_1),.clk(gclk));
	jdff dff_B_3DZdZwSO7_1(.din(w_dff_B_BHZXVDlh5_1),.dout(w_dff_B_3DZdZwSO7_1),.clk(gclk));
	jdff dff_B_qgjwp6H59_1(.din(w_dff_B_3DZdZwSO7_1),.dout(w_dff_B_qgjwp6H59_1),.clk(gclk));
	jdff dff_B_FjISFoFn0_1(.din(w_dff_B_qgjwp6H59_1),.dout(w_dff_B_FjISFoFn0_1),.clk(gclk));
	jdff dff_B_eVP6afzg4_1(.din(w_dff_B_FjISFoFn0_1),.dout(w_dff_B_eVP6afzg4_1),.clk(gclk));
	jdff dff_B_dGAnLv7S1_1(.din(w_dff_B_eVP6afzg4_1),.dout(w_dff_B_dGAnLv7S1_1),.clk(gclk));
	jdff dff_B_wrltKf9t8_1(.din(w_dff_B_dGAnLv7S1_1),.dout(w_dff_B_wrltKf9t8_1),.clk(gclk));
	jdff dff_B_E6wfKDYf8_1(.din(w_dff_B_wrltKf9t8_1),.dout(w_dff_B_E6wfKDYf8_1),.clk(gclk));
	jdff dff_B_zstLw8Pf6_1(.din(w_dff_B_E6wfKDYf8_1),.dout(w_dff_B_zstLw8Pf6_1),.clk(gclk));
	jdff dff_B_iJZwrhS32_1(.din(w_dff_B_zstLw8Pf6_1),.dout(w_dff_B_iJZwrhS32_1),.clk(gclk));
	jdff dff_B_zW7vuYN68_1(.din(w_dff_B_iJZwrhS32_1),.dout(w_dff_B_zW7vuYN68_1),.clk(gclk));
	jdff dff_B_8qToVnRD6_1(.din(w_dff_B_zW7vuYN68_1),.dout(w_dff_B_8qToVnRD6_1),.clk(gclk));
	jdff dff_B_c3uE6Jvq8_1(.din(w_dff_B_8qToVnRD6_1),.dout(w_dff_B_c3uE6Jvq8_1),.clk(gclk));
	jdff dff_B_aFajiWuF4_1(.din(w_dff_B_c3uE6Jvq8_1),.dout(w_dff_B_aFajiWuF4_1),.clk(gclk));
	jdff dff_B_9SPTMo1L0_1(.din(w_dff_B_aFajiWuF4_1),.dout(w_dff_B_9SPTMo1L0_1),.clk(gclk));
	jdff dff_B_UkSdvZEm2_1(.din(w_dff_B_9SPTMo1L0_1),.dout(w_dff_B_UkSdvZEm2_1),.clk(gclk));
	jdff dff_B_KuA1hRWS2_1(.din(w_dff_B_UkSdvZEm2_1),.dout(w_dff_B_KuA1hRWS2_1),.clk(gclk));
	jdff dff_B_mQKcb8SE7_1(.din(w_dff_B_KuA1hRWS2_1),.dout(w_dff_B_mQKcb8SE7_1),.clk(gclk));
	jdff dff_B_tLUqMK891_1(.din(w_dff_B_mQKcb8SE7_1),.dout(w_dff_B_tLUqMK891_1),.clk(gclk));
	jdff dff_B_qsRDDkov8_1(.din(w_dff_B_tLUqMK891_1),.dout(w_dff_B_qsRDDkov8_1),.clk(gclk));
	jdff dff_B_g8KZL2Hr0_1(.din(w_dff_B_qsRDDkov8_1),.dout(w_dff_B_g8KZL2Hr0_1),.clk(gclk));
	jdff dff_B_qeGANq7a7_1(.din(w_dff_B_g8KZL2Hr0_1),.dout(w_dff_B_qeGANq7a7_1),.clk(gclk));
	jdff dff_B_MxjdNVv43_1(.din(w_dff_B_qeGANq7a7_1),.dout(w_dff_B_MxjdNVv43_1),.clk(gclk));
	jdff dff_B_dZSiIDYK9_1(.din(w_dff_B_MxjdNVv43_1),.dout(w_dff_B_dZSiIDYK9_1),.clk(gclk));
	jdff dff_B_5aDJs0GN8_1(.din(w_dff_B_dZSiIDYK9_1),.dout(w_dff_B_5aDJs0GN8_1),.clk(gclk));
	jdff dff_B_6T6hcWBO8_1(.din(w_dff_B_5aDJs0GN8_1),.dout(w_dff_B_6T6hcWBO8_1),.clk(gclk));
	jdff dff_B_bTpRRFzg5_1(.din(w_dff_B_6T6hcWBO8_1),.dout(w_dff_B_bTpRRFzg5_1),.clk(gclk));
	jdff dff_B_YGtQo8gn1_1(.din(w_dff_B_bTpRRFzg5_1),.dout(w_dff_B_YGtQo8gn1_1),.clk(gclk));
	jdff dff_B_zrDe780f4_1(.din(w_dff_B_YGtQo8gn1_1),.dout(w_dff_B_zrDe780f4_1),.clk(gclk));
	jdff dff_B_rxgdsmxm4_1(.din(w_dff_B_zrDe780f4_1),.dout(w_dff_B_rxgdsmxm4_1),.clk(gclk));
	jdff dff_B_oKnqqtqY3_1(.din(w_dff_B_rxgdsmxm4_1),.dout(w_dff_B_oKnqqtqY3_1),.clk(gclk));
	jdff dff_B_GvHDDkT62_1(.din(w_dff_B_oKnqqtqY3_1),.dout(w_dff_B_GvHDDkT62_1),.clk(gclk));
	jdff dff_B_UlL2W78Z6_1(.din(w_dff_B_GvHDDkT62_1),.dout(w_dff_B_UlL2W78Z6_1),.clk(gclk));
	jdff dff_B_V41fX9643_1(.din(w_dff_B_UlL2W78Z6_1),.dout(w_dff_B_V41fX9643_1),.clk(gclk));
	jdff dff_B_6bVTpYNH6_1(.din(w_dff_B_V41fX9643_1),.dout(w_dff_B_6bVTpYNH6_1),.clk(gclk));
	jdff dff_B_yOlqlKDM7_1(.din(w_dff_B_6bVTpYNH6_1),.dout(w_dff_B_yOlqlKDM7_1),.clk(gclk));
	jdff dff_B_QdvKYQ2L9_1(.din(w_dff_B_yOlqlKDM7_1),.dout(w_dff_B_QdvKYQ2L9_1),.clk(gclk));
	jdff dff_B_06brwXGZ0_1(.din(w_dff_B_QdvKYQ2L9_1),.dout(w_dff_B_06brwXGZ0_1),.clk(gclk));
	jdff dff_B_Fx8sXFkn9_1(.din(w_dff_B_06brwXGZ0_1),.dout(w_dff_B_Fx8sXFkn9_1),.clk(gclk));
	jdff dff_B_FbtI6Of34_0(.din(n655),.dout(w_dff_B_FbtI6Of34_0),.clk(gclk));
	jdff dff_B_XDIlVbMV0_0(.din(w_dff_B_FbtI6Of34_0),.dout(w_dff_B_XDIlVbMV0_0),.clk(gclk));
	jdff dff_B_eCaRibv90_0(.din(w_dff_B_XDIlVbMV0_0),.dout(w_dff_B_eCaRibv90_0),.clk(gclk));
	jdff dff_B_kW2IixvL6_0(.din(w_dff_B_eCaRibv90_0),.dout(w_dff_B_kW2IixvL6_0),.clk(gclk));
	jdff dff_B_LfgYQ0ge5_0(.din(w_dff_B_kW2IixvL6_0),.dout(w_dff_B_LfgYQ0ge5_0),.clk(gclk));
	jdff dff_B_E23eIArt9_0(.din(w_dff_B_LfgYQ0ge5_0),.dout(w_dff_B_E23eIArt9_0),.clk(gclk));
	jdff dff_B_uMppIBr96_0(.din(w_dff_B_E23eIArt9_0),.dout(w_dff_B_uMppIBr96_0),.clk(gclk));
	jdff dff_B_XoByUtor9_0(.din(w_dff_B_uMppIBr96_0),.dout(w_dff_B_XoByUtor9_0),.clk(gclk));
	jdff dff_B_N2Xmux2n4_0(.din(w_dff_B_XoByUtor9_0),.dout(w_dff_B_N2Xmux2n4_0),.clk(gclk));
	jdff dff_B_y7iCFvdQ0_0(.din(w_dff_B_N2Xmux2n4_0),.dout(w_dff_B_y7iCFvdQ0_0),.clk(gclk));
	jdff dff_B_ZZ2qEJM67_0(.din(w_dff_B_y7iCFvdQ0_0),.dout(w_dff_B_ZZ2qEJM67_0),.clk(gclk));
	jdff dff_B_WhCYHgX61_0(.din(w_dff_B_ZZ2qEJM67_0),.dout(w_dff_B_WhCYHgX61_0),.clk(gclk));
	jdff dff_B_fRebIAFe5_0(.din(w_dff_B_WhCYHgX61_0),.dout(w_dff_B_fRebIAFe5_0),.clk(gclk));
	jdff dff_B_GHVhWHSr4_0(.din(w_dff_B_fRebIAFe5_0),.dout(w_dff_B_GHVhWHSr4_0),.clk(gclk));
	jdff dff_B_Bxujhhbu5_0(.din(w_dff_B_GHVhWHSr4_0),.dout(w_dff_B_Bxujhhbu5_0),.clk(gclk));
	jdff dff_B_7Hpz5qb68_0(.din(w_dff_B_Bxujhhbu5_0),.dout(w_dff_B_7Hpz5qb68_0),.clk(gclk));
	jdff dff_B_Ccp5HXRm9_0(.din(w_dff_B_7Hpz5qb68_0),.dout(w_dff_B_Ccp5HXRm9_0),.clk(gclk));
	jdff dff_B_s72c2n8R6_0(.din(w_dff_B_Ccp5HXRm9_0),.dout(w_dff_B_s72c2n8R6_0),.clk(gclk));
	jdff dff_B_2DLnntdb6_0(.din(w_dff_B_s72c2n8R6_0),.dout(w_dff_B_2DLnntdb6_0),.clk(gclk));
	jdff dff_B_QDRaTnnQ7_0(.din(w_dff_B_2DLnntdb6_0),.dout(w_dff_B_QDRaTnnQ7_0),.clk(gclk));
	jdff dff_B_WFGXknLw9_0(.din(w_dff_B_QDRaTnnQ7_0),.dout(w_dff_B_WFGXknLw9_0),.clk(gclk));
	jdff dff_B_AUaRfcRm1_0(.din(w_dff_B_WFGXknLw9_0),.dout(w_dff_B_AUaRfcRm1_0),.clk(gclk));
	jdff dff_B_rXCzInwj3_0(.din(w_dff_B_AUaRfcRm1_0),.dout(w_dff_B_rXCzInwj3_0),.clk(gclk));
	jdff dff_B_yaLJiO3n9_0(.din(w_dff_B_rXCzInwj3_0),.dout(w_dff_B_yaLJiO3n9_0),.clk(gclk));
	jdff dff_B_5DQoXppv8_0(.din(w_dff_B_yaLJiO3n9_0),.dout(w_dff_B_5DQoXppv8_0),.clk(gclk));
	jdff dff_B_5s19uiwV6_0(.din(w_dff_B_5DQoXppv8_0),.dout(w_dff_B_5s19uiwV6_0),.clk(gclk));
	jdff dff_B_xuj8m10v6_0(.din(w_dff_B_5s19uiwV6_0),.dout(w_dff_B_xuj8m10v6_0),.clk(gclk));
	jdff dff_B_rlN7NpqB4_0(.din(w_dff_B_xuj8m10v6_0),.dout(w_dff_B_rlN7NpqB4_0),.clk(gclk));
	jdff dff_B_46Uwhuwb6_0(.din(w_dff_B_rlN7NpqB4_0),.dout(w_dff_B_46Uwhuwb6_0),.clk(gclk));
	jdff dff_B_z4UHXo5W6_0(.din(w_dff_B_46Uwhuwb6_0),.dout(w_dff_B_z4UHXo5W6_0),.clk(gclk));
	jdff dff_B_6dwXgyjx3_0(.din(w_dff_B_z4UHXo5W6_0),.dout(w_dff_B_6dwXgyjx3_0),.clk(gclk));
	jdff dff_B_YmFpfVVW8_0(.din(w_dff_B_6dwXgyjx3_0),.dout(w_dff_B_YmFpfVVW8_0),.clk(gclk));
	jdff dff_B_TU7GA8Qi2_0(.din(w_dff_B_YmFpfVVW8_0),.dout(w_dff_B_TU7GA8Qi2_0),.clk(gclk));
	jdff dff_B_W9Xb6OZx8_0(.din(w_dff_B_TU7GA8Qi2_0),.dout(w_dff_B_W9Xb6OZx8_0),.clk(gclk));
	jdff dff_B_2UNFf4Ty5_0(.din(w_dff_B_W9Xb6OZx8_0),.dout(w_dff_B_2UNFf4Ty5_0),.clk(gclk));
	jdff dff_B_IDcAj2xk5_0(.din(w_dff_B_2UNFf4Ty5_0),.dout(w_dff_B_IDcAj2xk5_0),.clk(gclk));
	jdff dff_B_IIK19u7o6_0(.din(w_dff_B_IDcAj2xk5_0),.dout(w_dff_B_IIK19u7o6_0),.clk(gclk));
	jdff dff_B_cgSfWJbn2_0(.din(w_dff_B_IIK19u7o6_0),.dout(w_dff_B_cgSfWJbn2_0),.clk(gclk));
	jdff dff_B_5uh1eMy41_0(.din(w_dff_B_cgSfWJbn2_0),.dout(w_dff_B_5uh1eMy41_0),.clk(gclk));
	jdff dff_B_ltZQHJzB0_0(.din(w_dff_B_5uh1eMy41_0),.dout(w_dff_B_ltZQHJzB0_0),.clk(gclk));
	jdff dff_B_picAWtcF3_0(.din(w_dff_B_ltZQHJzB0_0),.dout(w_dff_B_picAWtcF3_0),.clk(gclk));
	jdff dff_B_yOnKICW88_0(.din(w_dff_B_picAWtcF3_0),.dout(w_dff_B_yOnKICW88_0),.clk(gclk));
	jdff dff_B_AaGCz7o39_0(.din(w_dff_B_yOnKICW88_0),.dout(w_dff_B_AaGCz7o39_0),.clk(gclk));
	jdff dff_B_Tc3H8Sc58_0(.din(w_dff_B_AaGCz7o39_0),.dout(w_dff_B_Tc3H8Sc58_0),.clk(gclk));
	jdff dff_B_ru1ByfvL1_0(.din(w_dff_B_Tc3H8Sc58_0),.dout(w_dff_B_ru1ByfvL1_0),.clk(gclk));
	jdff dff_B_ZbhWhr9i0_1(.din(n648),.dout(w_dff_B_ZbhWhr9i0_1),.clk(gclk));
	jdff dff_B_pwsoJJEN3_1(.din(w_dff_B_ZbhWhr9i0_1),.dout(w_dff_B_pwsoJJEN3_1),.clk(gclk));
	jdff dff_B_wq6ka6iV3_1(.din(w_dff_B_pwsoJJEN3_1),.dout(w_dff_B_wq6ka6iV3_1),.clk(gclk));
	jdff dff_B_uAgzUDyg8_1(.din(w_dff_B_wq6ka6iV3_1),.dout(w_dff_B_uAgzUDyg8_1),.clk(gclk));
	jdff dff_B_AeRvJUhx5_1(.din(w_dff_B_uAgzUDyg8_1),.dout(w_dff_B_AeRvJUhx5_1),.clk(gclk));
	jdff dff_B_2CW2rMrE2_1(.din(w_dff_B_AeRvJUhx5_1),.dout(w_dff_B_2CW2rMrE2_1),.clk(gclk));
	jdff dff_B_5beuRPkf9_1(.din(w_dff_B_2CW2rMrE2_1),.dout(w_dff_B_5beuRPkf9_1),.clk(gclk));
	jdff dff_B_U3TaZbq12_1(.din(w_dff_B_5beuRPkf9_1),.dout(w_dff_B_U3TaZbq12_1),.clk(gclk));
	jdff dff_B_7XCG2brg3_1(.din(w_dff_B_U3TaZbq12_1),.dout(w_dff_B_7XCG2brg3_1),.clk(gclk));
	jdff dff_B_2IDYKDSB4_1(.din(w_dff_B_7XCG2brg3_1),.dout(w_dff_B_2IDYKDSB4_1),.clk(gclk));
	jdff dff_B_qv8EtgK93_1(.din(w_dff_B_2IDYKDSB4_1),.dout(w_dff_B_qv8EtgK93_1),.clk(gclk));
	jdff dff_B_OInE0V554_1(.din(w_dff_B_qv8EtgK93_1),.dout(w_dff_B_OInE0V554_1),.clk(gclk));
	jdff dff_B_I4qmYqrl8_1(.din(w_dff_B_OInE0V554_1),.dout(w_dff_B_I4qmYqrl8_1),.clk(gclk));
	jdff dff_B_FJ1p4NKB9_1(.din(w_dff_B_I4qmYqrl8_1),.dout(w_dff_B_FJ1p4NKB9_1),.clk(gclk));
	jdff dff_B_yTzjFn1Z3_1(.din(w_dff_B_FJ1p4NKB9_1),.dout(w_dff_B_yTzjFn1Z3_1),.clk(gclk));
	jdff dff_B_SRSGRlyT9_1(.din(w_dff_B_yTzjFn1Z3_1),.dout(w_dff_B_SRSGRlyT9_1),.clk(gclk));
	jdff dff_B_DSZxKQR17_1(.din(w_dff_B_SRSGRlyT9_1),.dout(w_dff_B_DSZxKQR17_1),.clk(gclk));
	jdff dff_B_cErlBgLi0_1(.din(w_dff_B_DSZxKQR17_1),.dout(w_dff_B_cErlBgLi0_1),.clk(gclk));
	jdff dff_B_iAiTcOsN1_1(.din(w_dff_B_cErlBgLi0_1),.dout(w_dff_B_iAiTcOsN1_1),.clk(gclk));
	jdff dff_B_UvuNRS5J0_1(.din(w_dff_B_iAiTcOsN1_1),.dout(w_dff_B_UvuNRS5J0_1),.clk(gclk));
	jdff dff_B_3Ojifvup9_1(.din(w_dff_B_UvuNRS5J0_1),.dout(w_dff_B_3Ojifvup9_1),.clk(gclk));
	jdff dff_B_IN6YxyS01_1(.din(w_dff_B_3Ojifvup9_1),.dout(w_dff_B_IN6YxyS01_1),.clk(gclk));
	jdff dff_B_riZB7D8v0_1(.din(w_dff_B_IN6YxyS01_1),.dout(w_dff_B_riZB7D8v0_1),.clk(gclk));
	jdff dff_B_zSBr4CkT5_1(.din(w_dff_B_riZB7D8v0_1),.dout(w_dff_B_zSBr4CkT5_1),.clk(gclk));
	jdff dff_B_w9foHQ6s1_1(.din(w_dff_B_zSBr4CkT5_1),.dout(w_dff_B_w9foHQ6s1_1),.clk(gclk));
	jdff dff_B_4LRWFXGT3_1(.din(w_dff_B_w9foHQ6s1_1),.dout(w_dff_B_4LRWFXGT3_1),.clk(gclk));
	jdff dff_B_O0b8v42C3_1(.din(w_dff_B_4LRWFXGT3_1),.dout(w_dff_B_O0b8v42C3_1),.clk(gclk));
	jdff dff_B_bYfmDYht4_1(.din(w_dff_B_O0b8v42C3_1),.dout(w_dff_B_bYfmDYht4_1),.clk(gclk));
	jdff dff_B_5qgNxNOJ5_1(.din(w_dff_B_bYfmDYht4_1),.dout(w_dff_B_5qgNxNOJ5_1),.clk(gclk));
	jdff dff_B_L9jk8hv28_1(.din(w_dff_B_5qgNxNOJ5_1),.dout(w_dff_B_L9jk8hv28_1),.clk(gclk));
	jdff dff_B_bf80tCGe1_1(.din(w_dff_B_L9jk8hv28_1),.dout(w_dff_B_bf80tCGe1_1),.clk(gclk));
	jdff dff_B_CICJpYsg8_1(.din(w_dff_B_bf80tCGe1_1),.dout(w_dff_B_CICJpYsg8_1),.clk(gclk));
	jdff dff_B_aSlR0yiB8_1(.din(w_dff_B_CICJpYsg8_1),.dout(w_dff_B_aSlR0yiB8_1),.clk(gclk));
	jdff dff_B_Ipg9G7pv1_1(.din(w_dff_B_aSlR0yiB8_1),.dout(w_dff_B_Ipg9G7pv1_1),.clk(gclk));
	jdff dff_B_OkRAWWVb1_1(.din(w_dff_B_Ipg9G7pv1_1),.dout(w_dff_B_OkRAWWVb1_1),.clk(gclk));
	jdff dff_B_WeMiE7JE1_1(.din(w_dff_B_OkRAWWVb1_1),.dout(w_dff_B_WeMiE7JE1_1),.clk(gclk));
	jdff dff_B_5BgT35oh5_1(.din(w_dff_B_WeMiE7JE1_1),.dout(w_dff_B_5BgT35oh5_1),.clk(gclk));
	jdff dff_B_Oyu48oAj2_1(.din(w_dff_B_5BgT35oh5_1),.dout(w_dff_B_Oyu48oAj2_1),.clk(gclk));
	jdff dff_B_uaEDwFjn2_1(.din(w_dff_B_Oyu48oAj2_1),.dout(w_dff_B_uaEDwFjn2_1),.clk(gclk));
	jdff dff_B_2RX2wqtp4_1(.din(w_dff_B_uaEDwFjn2_1),.dout(w_dff_B_2RX2wqtp4_1),.clk(gclk));
	jdff dff_B_DiaR3j2k7_1(.din(w_dff_B_2RX2wqtp4_1),.dout(w_dff_B_DiaR3j2k7_1),.clk(gclk));
	jdff dff_B_Yf4r0V2C1_1(.din(w_dff_B_DiaR3j2k7_1),.dout(w_dff_B_Yf4r0V2C1_1),.clk(gclk));
	jdff dff_B_OdLRh7Za6_1(.din(w_dff_B_Yf4r0V2C1_1),.dout(w_dff_B_OdLRh7Za6_1),.clk(gclk));
	jdff dff_B_y5N9hr4K5_1(.din(w_dff_B_OdLRh7Za6_1),.dout(w_dff_B_y5N9hr4K5_1),.clk(gclk));
	jdff dff_B_rkFLpgaS2_0(.din(n649),.dout(w_dff_B_rkFLpgaS2_0),.clk(gclk));
	jdff dff_B_S3LOZWvw8_0(.din(w_dff_B_rkFLpgaS2_0),.dout(w_dff_B_S3LOZWvw8_0),.clk(gclk));
	jdff dff_B_LoTvtAJc4_0(.din(w_dff_B_S3LOZWvw8_0),.dout(w_dff_B_LoTvtAJc4_0),.clk(gclk));
	jdff dff_B_d0CprS0L3_0(.din(w_dff_B_LoTvtAJc4_0),.dout(w_dff_B_d0CprS0L3_0),.clk(gclk));
	jdff dff_B_buPdR9c42_0(.din(w_dff_B_d0CprS0L3_0),.dout(w_dff_B_buPdR9c42_0),.clk(gclk));
	jdff dff_B_wDac1SNJ8_0(.din(w_dff_B_buPdR9c42_0),.dout(w_dff_B_wDac1SNJ8_0),.clk(gclk));
	jdff dff_B_JrZRhLJN3_0(.din(w_dff_B_wDac1SNJ8_0),.dout(w_dff_B_JrZRhLJN3_0),.clk(gclk));
	jdff dff_B_93tL2AYf2_0(.din(w_dff_B_JrZRhLJN3_0),.dout(w_dff_B_93tL2AYf2_0),.clk(gclk));
	jdff dff_B_YhpaIu4D4_0(.din(w_dff_B_93tL2AYf2_0),.dout(w_dff_B_YhpaIu4D4_0),.clk(gclk));
	jdff dff_B_q1a5rF7N6_0(.din(w_dff_B_YhpaIu4D4_0),.dout(w_dff_B_q1a5rF7N6_0),.clk(gclk));
	jdff dff_B_crQsYrUo4_0(.din(w_dff_B_q1a5rF7N6_0),.dout(w_dff_B_crQsYrUo4_0),.clk(gclk));
	jdff dff_B_4VnZWyum0_0(.din(w_dff_B_crQsYrUo4_0),.dout(w_dff_B_4VnZWyum0_0),.clk(gclk));
	jdff dff_B_vlxWcSOz7_0(.din(w_dff_B_4VnZWyum0_0),.dout(w_dff_B_vlxWcSOz7_0),.clk(gclk));
	jdff dff_B_sQ58d6Wc9_0(.din(w_dff_B_vlxWcSOz7_0),.dout(w_dff_B_sQ58d6Wc9_0),.clk(gclk));
	jdff dff_B_KCxSDtfF1_0(.din(w_dff_B_sQ58d6Wc9_0),.dout(w_dff_B_KCxSDtfF1_0),.clk(gclk));
	jdff dff_B_GkdOq5lE8_0(.din(w_dff_B_KCxSDtfF1_0),.dout(w_dff_B_GkdOq5lE8_0),.clk(gclk));
	jdff dff_B_N9cRcq5A6_0(.din(w_dff_B_GkdOq5lE8_0),.dout(w_dff_B_N9cRcq5A6_0),.clk(gclk));
	jdff dff_B_ivW5Zqpi7_0(.din(w_dff_B_N9cRcq5A6_0),.dout(w_dff_B_ivW5Zqpi7_0),.clk(gclk));
	jdff dff_B_Mmm72eLt8_0(.din(w_dff_B_ivW5Zqpi7_0),.dout(w_dff_B_Mmm72eLt8_0),.clk(gclk));
	jdff dff_B_cqGSFRGD7_0(.din(w_dff_B_Mmm72eLt8_0),.dout(w_dff_B_cqGSFRGD7_0),.clk(gclk));
	jdff dff_B_DT1w3ZyN0_0(.din(w_dff_B_cqGSFRGD7_0),.dout(w_dff_B_DT1w3ZyN0_0),.clk(gclk));
	jdff dff_B_1UFxYQH18_0(.din(w_dff_B_DT1w3ZyN0_0),.dout(w_dff_B_1UFxYQH18_0),.clk(gclk));
	jdff dff_B_CuM2w5TT6_0(.din(w_dff_B_1UFxYQH18_0),.dout(w_dff_B_CuM2w5TT6_0),.clk(gclk));
	jdff dff_B_nIyt3SmD3_0(.din(w_dff_B_CuM2w5TT6_0),.dout(w_dff_B_nIyt3SmD3_0),.clk(gclk));
	jdff dff_B_vq6JB6IU9_0(.din(w_dff_B_nIyt3SmD3_0),.dout(w_dff_B_vq6JB6IU9_0),.clk(gclk));
	jdff dff_B_Lbvj6yNV7_0(.din(w_dff_B_vq6JB6IU9_0),.dout(w_dff_B_Lbvj6yNV7_0),.clk(gclk));
	jdff dff_B_dLcS5xX39_0(.din(w_dff_B_Lbvj6yNV7_0),.dout(w_dff_B_dLcS5xX39_0),.clk(gclk));
	jdff dff_B_I3EZLtz33_0(.din(w_dff_B_dLcS5xX39_0),.dout(w_dff_B_I3EZLtz33_0),.clk(gclk));
	jdff dff_B_69D6oSmW9_0(.din(w_dff_B_I3EZLtz33_0),.dout(w_dff_B_69D6oSmW9_0),.clk(gclk));
	jdff dff_B_9mL590f38_0(.din(w_dff_B_69D6oSmW9_0),.dout(w_dff_B_9mL590f38_0),.clk(gclk));
	jdff dff_B_oRwYY0Nh0_0(.din(w_dff_B_9mL590f38_0),.dout(w_dff_B_oRwYY0Nh0_0),.clk(gclk));
	jdff dff_B_Bn0kH5WL1_0(.din(w_dff_B_oRwYY0Nh0_0),.dout(w_dff_B_Bn0kH5WL1_0),.clk(gclk));
	jdff dff_B_hgQsWDyx3_0(.din(w_dff_B_Bn0kH5WL1_0),.dout(w_dff_B_hgQsWDyx3_0),.clk(gclk));
	jdff dff_B_ReiD0qrT1_0(.din(w_dff_B_hgQsWDyx3_0),.dout(w_dff_B_ReiD0qrT1_0),.clk(gclk));
	jdff dff_B_al2HzM9O1_0(.din(w_dff_B_ReiD0qrT1_0),.dout(w_dff_B_al2HzM9O1_0),.clk(gclk));
	jdff dff_B_SlrMrmXS7_0(.din(w_dff_B_al2HzM9O1_0),.dout(w_dff_B_SlrMrmXS7_0),.clk(gclk));
	jdff dff_B_DCBYSJg66_0(.din(w_dff_B_SlrMrmXS7_0),.dout(w_dff_B_DCBYSJg66_0),.clk(gclk));
	jdff dff_B_lUAmwcSL1_0(.din(w_dff_B_DCBYSJg66_0),.dout(w_dff_B_lUAmwcSL1_0),.clk(gclk));
	jdff dff_B_Aug3b18x0_0(.din(w_dff_B_lUAmwcSL1_0),.dout(w_dff_B_Aug3b18x0_0),.clk(gclk));
	jdff dff_B_Tny9fVpg8_0(.din(w_dff_B_Aug3b18x0_0),.dout(w_dff_B_Tny9fVpg8_0),.clk(gclk));
	jdff dff_B_5AZs62he7_0(.din(w_dff_B_Tny9fVpg8_0),.dout(w_dff_B_5AZs62he7_0),.clk(gclk));
	jdff dff_B_ZzddWN548_0(.din(w_dff_B_5AZs62he7_0),.dout(w_dff_B_ZzddWN548_0),.clk(gclk));
	jdff dff_B_hy209J786_0(.din(w_dff_B_ZzddWN548_0),.dout(w_dff_B_hy209J786_0),.clk(gclk));
	jdff dff_B_XJ6b8ERc3_0(.din(w_dff_B_hy209J786_0),.dout(w_dff_B_XJ6b8ERc3_0),.clk(gclk));
	jdff dff_B_hmXEDbDG4_1(.din(n642),.dout(w_dff_B_hmXEDbDG4_1),.clk(gclk));
	jdff dff_B_tAKMLcDx5_1(.din(w_dff_B_hmXEDbDG4_1),.dout(w_dff_B_tAKMLcDx5_1),.clk(gclk));
	jdff dff_B_qcy2NM5A9_1(.din(w_dff_B_tAKMLcDx5_1),.dout(w_dff_B_qcy2NM5A9_1),.clk(gclk));
	jdff dff_B_nvNvYJlT6_1(.din(w_dff_B_qcy2NM5A9_1),.dout(w_dff_B_nvNvYJlT6_1),.clk(gclk));
	jdff dff_B_OldzLEIo1_1(.din(w_dff_B_nvNvYJlT6_1),.dout(w_dff_B_OldzLEIo1_1),.clk(gclk));
	jdff dff_B_rYqClixL7_1(.din(w_dff_B_OldzLEIo1_1),.dout(w_dff_B_rYqClixL7_1),.clk(gclk));
	jdff dff_B_VwjJ68u28_1(.din(w_dff_B_rYqClixL7_1),.dout(w_dff_B_VwjJ68u28_1),.clk(gclk));
	jdff dff_B_4kQ3BXYM6_1(.din(w_dff_B_VwjJ68u28_1),.dout(w_dff_B_4kQ3BXYM6_1),.clk(gclk));
	jdff dff_B_qZprjZLy9_1(.din(w_dff_B_4kQ3BXYM6_1),.dout(w_dff_B_qZprjZLy9_1),.clk(gclk));
	jdff dff_B_ZvKlv1NG2_1(.din(w_dff_B_qZprjZLy9_1),.dout(w_dff_B_ZvKlv1NG2_1),.clk(gclk));
	jdff dff_B_uPgYOZAa7_1(.din(w_dff_B_ZvKlv1NG2_1),.dout(w_dff_B_uPgYOZAa7_1),.clk(gclk));
	jdff dff_B_PWeIYkio6_1(.din(w_dff_B_uPgYOZAa7_1),.dout(w_dff_B_PWeIYkio6_1),.clk(gclk));
	jdff dff_B_evfM2W0p2_1(.din(w_dff_B_PWeIYkio6_1),.dout(w_dff_B_evfM2W0p2_1),.clk(gclk));
	jdff dff_B_XfqALNc12_1(.din(w_dff_B_evfM2W0p2_1),.dout(w_dff_B_XfqALNc12_1),.clk(gclk));
	jdff dff_B_zomaaGNg7_1(.din(w_dff_B_XfqALNc12_1),.dout(w_dff_B_zomaaGNg7_1),.clk(gclk));
	jdff dff_B_rwxtLz4s9_1(.din(w_dff_B_zomaaGNg7_1),.dout(w_dff_B_rwxtLz4s9_1),.clk(gclk));
	jdff dff_B_5TDEQuhY7_1(.din(w_dff_B_rwxtLz4s9_1),.dout(w_dff_B_5TDEQuhY7_1),.clk(gclk));
	jdff dff_B_kZhyqGCq0_1(.din(w_dff_B_5TDEQuhY7_1),.dout(w_dff_B_kZhyqGCq0_1),.clk(gclk));
	jdff dff_B_hvCzCf3a9_1(.din(w_dff_B_kZhyqGCq0_1),.dout(w_dff_B_hvCzCf3a9_1),.clk(gclk));
	jdff dff_B_TKJIU4lu4_1(.din(w_dff_B_hvCzCf3a9_1),.dout(w_dff_B_TKJIU4lu4_1),.clk(gclk));
	jdff dff_B_DW4uxPVp3_1(.din(w_dff_B_TKJIU4lu4_1),.dout(w_dff_B_DW4uxPVp3_1),.clk(gclk));
	jdff dff_B_sc1hreCE8_1(.din(w_dff_B_DW4uxPVp3_1),.dout(w_dff_B_sc1hreCE8_1),.clk(gclk));
	jdff dff_B_4Uyq7GMV3_1(.din(w_dff_B_sc1hreCE8_1),.dout(w_dff_B_4Uyq7GMV3_1),.clk(gclk));
	jdff dff_B_iAIZ3eEk3_1(.din(w_dff_B_4Uyq7GMV3_1),.dout(w_dff_B_iAIZ3eEk3_1),.clk(gclk));
	jdff dff_B_jpco5LcG1_1(.din(w_dff_B_iAIZ3eEk3_1),.dout(w_dff_B_jpco5LcG1_1),.clk(gclk));
	jdff dff_B_JLALGLXw4_1(.din(w_dff_B_jpco5LcG1_1),.dout(w_dff_B_JLALGLXw4_1),.clk(gclk));
	jdff dff_B_sNirE9If7_1(.din(w_dff_B_JLALGLXw4_1),.dout(w_dff_B_sNirE9If7_1),.clk(gclk));
	jdff dff_B_45hiEaMW8_1(.din(w_dff_B_sNirE9If7_1),.dout(w_dff_B_45hiEaMW8_1),.clk(gclk));
	jdff dff_B_OOFHBLuB8_1(.din(w_dff_B_45hiEaMW8_1),.dout(w_dff_B_OOFHBLuB8_1),.clk(gclk));
	jdff dff_B_BBfyzCDk5_1(.din(w_dff_B_OOFHBLuB8_1),.dout(w_dff_B_BBfyzCDk5_1),.clk(gclk));
	jdff dff_B_EfMLlRon4_1(.din(w_dff_B_BBfyzCDk5_1),.dout(w_dff_B_EfMLlRon4_1),.clk(gclk));
	jdff dff_B_GQ9mPjde4_1(.din(w_dff_B_EfMLlRon4_1),.dout(w_dff_B_GQ9mPjde4_1),.clk(gclk));
	jdff dff_B_ncShczgI2_1(.din(w_dff_B_GQ9mPjde4_1),.dout(w_dff_B_ncShczgI2_1),.clk(gclk));
	jdff dff_B_eqgTEXam7_1(.din(w_dff_B_ncShczgI2_1),.dout(w_dff_B_eqgTEXam7_1),.clk(gclk));
	jdff dff_B_ltCw1BIv3_1(.din(w_dff_B_eqgTEXam7_1),.dout(w_dff_B_ltCw1BIv3_1),.clk(gclk));
	jdff dff_B_zl72ZCTT2_1(.din(w_dff_B_ltCw1BIv3_1),.dout(w_dff_B_zl72ZCTT2_1),.clk(gclk));
	jdff dff_B_vI4GBiwP8_1(.din(w_dff_B_zl72ZCTT2_1),.dout(w_dff_B_vI4GBiwP8_1),.clk(gclk));
	jdff dff_B_lqeuXDbv6_1(.din(w_dff_B_vI4GBiwP8_1),.dout(w_dff_B_lqeuXDbv6_1),.clk(gclk));
	jdff dff_B_QDNHosOz1_1(.din(w_dff_B_lqeuXDbv6_1),.dout(w_dff_B_QDNHosOz1_1),.clk(gclk));
	jdff dff_B_94wIuLld1_1(.din(w_dff_B_QDNHosOz1_1),.dout(w_dff_B_94wIuLld1_1),.clk(gclk));
	jdff dff_B_RY0SM2dq1_1(.din(w_dff_B_94wIuLld1_1),.dout(w_dff_B_RY0SM2dq1_1),.clk(gclk));
	jdff dff_B_INBVpObJ2_1(.din(w_dff_B_RY0SM2dq1_1),.dout(w_dff_B_INBVpObJ2_1),.clk(gclk));
	jdff dff_B_OGZRqfWA9_1(.din(w_dff_B_INBVpObJ2_1),.dout(w_dff_B_OGZRqfWA9_1),.clk(gclk));
	jdff dff_B_VVBVUF222_0(.din(n643),.dout(w_dff_B_VVBVUF222_0),.clk(gclk));
	jdff dff_B_dJiUKVNg4_0(.din(w_dff_B_VVBVUF222_0),.dout(w_dff_B_dJiUKVNg4_0),.clk(gclk));
	jdff dff_B_sxj8NmoB9_0(.din(w_dff_B_dJiUKVNg4_0),.dout(w_dff_B_sxj8NmoB9_0),.clk(gclk));
	jdff dff_B_4CuSmZZ12_0(.din(w_dff_B_sxj8NmoB9_0),.dout(w_dff_B_4CuSmZZ12_0),.clk(gclk));
	jdff dff_B_4eXe4Rzb2_0(.din(w_dff_B_4CuSmZZ12_0),.dout(w_dff_B_4eXe4Rzb2_0),.clk(gclk));
	jdff dff_B_9qxlf1dl6_0(.din(w_dff_B_4eXe4Rzb2_0),.dout(w_dff_B_9qxlf1dl6_0),.clk(gclk));
	jdff dff_B_qZOEJsS60_0(.din(w_dff_B_9qxlf1dl6_0),.dout(w_dff_B_qZOEJsS60_0),.clk(gclk));
	jdff dff_B_7iZNVHLr6_0(.din(w_dff_B_qZOEJsS60_0),.dout(w_dff_B_7iZNVHLr6_0),.clk(gclk));
	jdff dff_B_8HD9x4128_0(.din(w_dff_B_7iZNVHLr6_0),.dout(w_dff_B_8HD9x4128_0),.clk(gclk));
	jdff dff_B_e47r6vrl8_0(.din(w_dff_B_8HD9x4128_0),.dout(w_dff_B_e47r6vrl8_0),.clk(gclk));
	jdff dff_B_uNUhQLKP7_0(.din(w_dff_B_e47r6vrl8_0),.dout(w_dff_B_uNUhQLKP7_0),.clk(gclk));
	jdff dff_B_GqCWByrM3_0(.din(w_dff_B_uNUhQLKP7_0),.dout(w_dff_B_GqCWByrM3_0),.clk(gclk));
	jdff dff_B_3mZkS0QV7_0(.din(w_dff_B_GqCWByrM3_0),.dout(w_dff_B_3mZkS0QV7_0),.clk(gclk));
	jdff dff_B_rH3stAxW8_0(.din(w_dff_B_3mZkS0QV7_0),.dout(w_dff_B_rH3stAxW8_0),.clk(gclk));
	jdff dff_B_eNzgpg0A5_0(.din(w_dff_B_rH3stAxW8_0),.dout(w_dff_B_eNzgpg0A5_0),.clk(gclk));
	jdff dff_B_j8Sjl2VU8_0(.din(w_dff_B_eNzgpg0A5_0),.dout(w_dff_B_j8Sjl2VU8_0),.clk(gclk));
	jdff dff_B_squWjeIf5_0(.din(w_dff_B_j8Sjl2VU8_0),.dout(w_dff_B_squWjeIf5_0),.clk(gclk));
	jdff dff_B_Un8OMywj5_0(.din(w_dff_B_squWjeIf5_0),.dout(w_dff_B_Un8OMywj5_0),.clk(gclk));
	jdff dff_B_nSBg6gC83_0(.din(w_dff_B_Un8OMywj5_0),.dout(w_dff_B_nSBg6gC83_0),.clk(gclk));
	jdff dff_B_HW9QDRPy6_0(.din(w_dff_B_nSBg6gC83_0),.dout(w_dff_B_HW9QDRPy6_0),.clk(gclk));
	jdff dff_B_KW0rY31m7_0(.din(w_dff_B_HW9QDRPy6_0),.dout(w_dff_B_KW0rY31m7_0),.clk(gclk));
	jdff dff_B_7xpzeyZY0_0(.din(w_dff_B_KW0rY31m7_0),.dout(w_dff_B_7xpzeyZY0_0),.clk(gclk));
	jdff dff_B_5fY9Roe13_0(.din(w_dff_B_7xpzeyZY0_0),.dout(w_dff_B_5fY9Roe13_0),.clk(gclk));
	jdff dff_B_EjbYz7756_0(.din(w_dff_B_5fY9Roe13_0),.dout(w_dff_B_EjbYz7756_0),.clk(gclk));
	jdff dff_B_fA27xfmz5_0(.din(w_dff_B_EjbYz7756_0),.dout(w_dff_B_fA27xfmz5_0),.clk(gclk));
	jdff dff_B_AFUcymdh8_0(.din(w_dff_B_fA27xfmz5_0),.dout(w_dff_B_AFUcymdh8_0),.clk(gclk));
	jdff dff_B_IyRtfTsA2_0(.din(w_dff_B_AFUcymdh8_0),.dout(w_dff_B_IyRtfTsA2_0),.clk(gclk));
	jdff dff_B_zciLAZl70_0(.din(w_dff_B_IyRtfTsA2_0),.dout(w_dff_B_zciLAZl70_0),.clk(gclk));
	jdff dff_B_UTBQFDlX6_0(.din(w_dff_B_zciLAZl70_0),.dout(w_dff_B_UTBQFDlX6_0),.clk(gclk));
	jdff dff_B_YXvOjyel5_0(.din(w_dff_B_UTBQFDlX6_0),.dout(w_dff_B_YXvOjyel5_0),.clk(gclk));
	jdff dff_B_Fcp0nyhg4_0(.din(w_dff_B_YXvOjyel5_0),.dout(w_dff_B_Fcp0nyhg4_0),.clk(gclk));
	jdff dff_B_i7pyVAgt8_0(.din(w_dff_B_Fcp0nyhg4_0),.dout(w_dff_B_i7pyVAgt8_0),.clk(gclk));
	jdff dff_B_K2PKQ5uq7_0(.din(w_dff_B_i7pyVAgt8_0),.dout(w_dff_B_K2PKQ5uq7_0),.clk(gclk));
	jdff dff_B_FoR2v05a5_0(.din(w_dff_B_K2PKQ5uq7_0),.dout(w_dff_B_FoR2v05a5_0),.clk(gclk));
	jdff dff_B_9SxyD6vQ9_0(.din(w_dff_B_FoR2v05a5_0),.dout(w_dff_B_9SxyD6vQ9_0),.clk(gclk));
	jdff dff_B_XafsW9UQ1_0(.din(w_dff_B_9SxyD6vQ9_0),.dout(w_dff_B_XafsW9UQ1_0),.clk(gclk));
	jdff dff_B_BTAE8Es11_0(.din(w_dff_B_XafsW9UQ1_0),.dout(w_dff_B_BTAE8Es11_0),.clk(gclk));
	jdff dff_B_yT7dIv8Q0_0(.din(w_dff_B_BTAE8Es11_0),.dout(w_dff_B_yT7dIv8Q0_0),.clk(gclk));
	jdff dff_B_OKsCZfTR4_0(.din(w_dff_B_yT7dIv8Q0_0),.dout(w_dff_B_OKsCZfTR4_0),.clk(gclk));
	jdff dff_B_y7gRlNEB5_0(.din(w_dff_B_OKsCZfTR4_0),.dout(w_dff_B_y7gRlNEB5_0),.clk(gclk));
	jdff dff_B_5T8yzaqJ1_0(.din(w_dff_B_y7gRlNEB5_0),.dout(w_dff_B_5T8yzaqJ1_0),.clk(gclk));
	jdff dff_B_ntLbGJVc0_0(.din(w_dff_B_5T8yzaqJ1_0),.dout(w_dff_B_ntLbGJVc0_0),.clk(gclk));
	jdff dff_B_O1mNMYi88_0(.din(w_dff_B_ntLbGJVc0_0),.dout(w_dff_B_O1mNMYi88_0),.clk(gclk));
	jdff dff_B_I7LqbT2f6_1(.din(n636),.dout(w_dff_B_I7LqbT2f6_1),.clk(gclk));
	jdff dff_B_wVR5WhD46_1(.din(w_dff_B_I7LqbT2f6_1),.dout(w_dff_B_wVR5WhD46_1),.clk(gclk));
	jdff dff_B_D7PpRXsQ3_1(.din(w_dff_B_wVR5WhD46_1),.dout(w_dff_B_D7PpRXsQ3_1),.clk(gclk));
	jdff dff_B_KagA3vx81_1(.din(w_dff_B_D7PpRXsQ3_1),.dout(w_dff_B_KagA3vx81_1),.clk(gclk));
	jdff dff_B_WS2gRnrE3_1(.din(w_dff_B_KagA3vx81_1),.dout(w_dff_B_WS2gRnrE3_1),.clk(gclk));
	jdff dff_B_diIbVVjn3_1(.din(w_dff_B_WS2gRnrE3_1),.dout(w_dff_B_diIbVVjn3_1),.clk(gclk));
	jdff dff_B_vBFGn19E8_1(.din(w_dff_B_diIbVVjn3_1),.dout(w_dff_B_vBFGn19E8_1),.clk(gclk));
	jdff dff_B_s9J8fvom2_1(.din(w_dff_B_vBFGn19E8_1),.dout(w_dff_B_s9J8fvom2_1),.clk(gclk));
	jdff dff_B_GdFp3fIg8_1(.din(w_dff_B_s9J8fvom2_1),.dout(w_dff_B_GdFp3fIg8_1),.clk(gclk));
	jdff dff_B_CLfn7nv39_1(.din(w_dff_B_GdFp3fIg8_1),.dout(w_dff_B_CLfn7nv39_1),.clk(gclk));
	jdff dff_B_9LbufJdN7_1(.din(w_dff_B_CLfn7nv39_1),.dout(w_dff_B_9LbufJdN7_1),.clk(gclk));
	jdff dff_B_HXBPWuK24_1(.din(w_dff_B_9LbufJdN7_1),.dout(w_dff_B_HXBPWuK24_1),.clk(gclk));
	jdff dff_B_Y0L3hPQ42_1(.din(w_dff_B_HXBPWuK24_1),.dout(w_dff_B_Y0L3hPQ42_1),.clk(gclk));
	jdff dff_B_QwcrBjxJ0_1(.din(w_dff_B_Y0L3hPQ42_1),.dout(w_dff_B_QwcrBjxJ0_1),.clk(gclk));
	jdff dff_B_AYkb6pPK8_1(.din(w_dff_B_QwcrBjxJ0_1),.dout(w_dff_B_AYkb6pPK8_1),.clk(gclk));
	jdff dff_B_UvpjWccQ2_1(.din(w_dff_B_AYkb6pPK8_1),.dout(w_dff_B_UvpjWccQ2_1),.clk(gclk));
	jdff dff_B_zfncn8f53_1(.din(w_dff_B_UvpjWccQ2_1),.dout(w_dff_B_zfncn8f53_1),.clk(gclk));
	jdff dff_B_EjYAWdsV3_1(.din(w_dff_B_zfncn8f53_1),.dout(w_dff_B_EjYAWdsV3_1),.clk(gclk));
	jdff dff_B_bNEs9cej4_1(.din(w_dff_B_EjYAWdsV3_1),.dout(w_dff_B_bNEs9cej4_1),.clk(gclk));
	jdff dff_B_woE3QMSV8_1(.din(w_dff_B_bNEs9cej4_1),.dout(w_dff_B_woE3QMSV8_1),.clk(gclk));
	jdff dff_B_vGS18eus3_1(.din(w_dff_B_woE3QMSV8_1),.dout(w_dff_B_vGS18eus3_1),.clk(gclk));
	jdff dff_B_BGuh95xX6_1(.din(w_dff_B_vGS18eus3_1),.dout(w_dff_B_BGuh95xX6_1),.clk(gclk));
	jdff dff_B_SKbrTr5H8_1(.din(w_dff_B_BGuh95xX6_1),.dout(w_dff_B_SKbrTr5H8_1),.clk(gclk));
	jdff dff_B_1dRHI08r1_1(.din(w_dff_B_SKbrTr5H8_1),.dout(w_dff_B_1dRHI08r1_1),.clk(gclk));
	jdff dff_B_W4yY2TYG2_1(.din(w_dff_B_1dRHI08r1_1),.dout(w_dff_B_W4yY2TYG2_1),.clk(gclk));
	jdff dff_B_2FBvsjGC4_1(.din(w_dff_B_W4yY2TYG2_1),.dout(w_dff_B_2FBvsjGC4_1),.clk(gclk));
	jdff dff_B_0eAzUOTC7_1(.din(w_dff_B_2FBvsjGC4_1),.dout(w_dff_B_0eAzUOTC7_1),.clk(gclk));
	jdff dff_B_mLwQ88MO4_1(.din(w_dff_B_0eAzUOTC7_1),.dout(w_dff_B_mLwQ88MO4_1),.clk(gclk));
	jdff dff_B_WeXoqRHL7_1(.din(w_dff_B_mLwQ88MO4_1),.dout(w_dff_B_WeXoqRHL7_1),.clk(gclk));
	jdff dff_B_5Ok4u67t8_1(.din(w_dff_B_WeXoqRHL7_1),.dout(w_dff_B_5Ok4u67t8_1),.clk(gclk));
	jdff dff_B_fd6fsVzN1_1(.din(w_dff_B_5Ok4u67t8_1),.dout(w_dff_B_fd6fsVzN1_1),.clk(gclk));
	jdff dff_B_ff2Mmcw55_1(.din(w_dff_B_fd6fsVzN1_1),.dout(w_dff_B_ff2Mmcw55_1),.clk(gclk));
	jdff dff_B_WHqckdFZ1_1(.din(w_dff_B_ff2Mmcw55_1),.dout(w_dff_B_WHqckdFZ1_1),.clk(gclk));
	jdff dff_B_A2aximwh1_1(.din(w_dff_B_WHqckdFZ1_1),.dout(w_dff_B_A2aximwh1_1),.clk(gclk));
	jdff dff_B_Y6BkQyQw2_1(.din(w_dff_B_A2aximwh1_1),.dout(w_dff_B_Y6BkQyQw2_1),.clk(gclk));
	jdff dff_B_hFmPcJDa1_1(.din(w_dff_B_Y6BkQyQw2_1),.dout(w_dff_B_hFmPcJDa1_1),.clk(gclk));
	jdff dff_B_Ii4Oanhf1_1(.din(w_dff_B_hFmPcJDa1_1),.dout(w_dff_B_Ii4Oanhf1_1),.clk(gclk));
	jdff dff_B_CpGhp91t1_1(.din(w_dff_B_Ii4Oanhf1_1),.dout(w_dff_B_CpGhp91t1_1),.clk(gclk));
	jdff dff_B_2twUHnhx1_1(.din(w_dff_B_CpGhp91t1_1),.dout(w_dff_B_2twUHnhx1_1),.clk(gclk));
	jdff dff_B_zIWJSRtM2_1(.din(w_dff_B_2twUHnhx1_1),.dout(w_dff_B_zIWJSRtM2_1),.clk(gclk));
	jdff dff_B_AkqcSZze2_1(.din(w_dff_B_zIWJSRtM2_1),.dout(w_dff_B_AkqcSZze2_1),.clk(gclk));
	jdff dff_B_JMCouiXX8_1(.din(w_dff_B_AkqcSZze2_1),.dout(w_dff_B_JMCouiXX8_1),.clk(gclk));
	jdff dff_B_AcSz1DMq5_0(.din(n637),.dout(w_dff_B_AcSz1DMq5_0),.clk(gclk));
	jdff dff_B_PJePDGCS2_0(.din(w_dff_B_AcSz1DMq5_0),.dout(w_dff_B_PJePDGCS2_0),.clk(gclk));
	jdff dff_B_NqHLJzGF9_0(.din(w_dff_B_PJePDGCS2_0),.dout(w_dff_B_NqHLJzGF9_0),.clk(gclk));
	jdff dff_B_il8JkgqN6_0(.din(w_dff_B_NqHLJzGF9_0),.dout(w_dff_B_il8JkgqN6_0),.clk(gclk));
	jdff dff_B_zQJPEKn48_0(.din(w_dff_B_il8JkgqN6_0),.dout(w_dff_B_zQJPEKn48_0),.clk(gclk));
	jdff dff_B_crfEaEZ47_0(.din(w_dff_B_zQJPEKn48_0),.dout(w_dff_B_crfEaEZ47_0),.clk(gclk));
	jdff dff_B_7zA5mFRp7_0(.din(w_dff_B_crfEaEZ47_0),.dout(w_dff_B_7zA5mFRp7_0),.clk(gclk));
	jdff dff_B_n6y0sVy43_0(.din(w_dff_B_7zA5mFRp7_0),.dout(w_dff_B_n6y0sVy43_0),.clk(gclk));
	jdff dff_B_KpbAV0gT4_0(.din(w_dff_B_n6y0sVy43_0),.dout(w_dff_B_KpbAV0gT4_0),.clk(gclk));
	jdff dff_B_pkI9WEZY4_0(.din(w_dff_B_KpbAV0gT4_0),.dout(w_dff_B_pkI9WEZY4_0),.clk(gclk));
	jdff dff_B_0fdd2xVV6_0(.din(w_dff_B_pkI9WEZY4_0),.dout(w_dff_B_0fdd2xVV6_0),.clk(gclk));
	jdff dff_B_5LduqPRo9_0(.din(w_dff_B_0fdd2xVV6_0),.dout(w_dff_B_5LduqPRo9_0),.clk(gclk));
	jdff dff_B_yPThiWtg6_0(.din(w_dff_B_5LduqPRo9_0),.dout(w_dff_B_yPThiWtg6_0),.clk(gclk));
	jdff dff_B_42s6Ek1s7_0(.din(w_dff_B_yPThiWtg6_0),.dout(w_dff_B_42s6Ek1s7_0),.clk(gclk));
	jdff dff_B_jINLYooY0_0(.din(w_dff_B_42s6Ek1s7_0),.dout(w_dff_B_jINLYooY0_0),.clk(gclk));
	jdff dff_B_H9n2s8wP1_0(.din(w_dff_B_jINLYooY0_0),.dout(w_dff_B_H9n2s8wP1_0),.clk(gclk));
	jdff dff_B_zlMEz8vm0_0(.din(w_dff_B_H9n2s8wP1_0),.dout(w_dff_B_zlMEz8vm0_0),.clk(gclk));
	jdff dff_B_OcQJchxO8_0(.din(w_dff_B_zlMEz8vm0_0),.dout(w_dff_B_OcQJchxO8_0),.clk(gclk));
	jdff dff_B_lXsVs8a26_0(.din(w_dff_B_OcQJchxO8_0),.dout(w_dff_B_lXsVs8a26_0),.clk(gclk));
	jdff dff_B_ufQptKRw5_0(.din(w_dff_B_lXsVs8a26_0),.dout(w_dff_B_ufQptKRw5_0),.clk(gclk));
	jdff dff_B_lfl0aAXB5_0(.din(w_dff_B_ufQptKRw5_0),.dout(w_dff_B_lfl0aAXB5_0),.clk(gclk));
	jdff dff_B_O1QkvmHl2_0(.din(w_dff_B_lfl0aAXB5_0),.dout(w_dff_B_O1QkvmHl2_0),.clk(gclk));
	jdff dff_B_mFnNs4YD8_0(.din(w_dff_B_O1QkvmHl2_0),.dout(w_dff_B_mFnNs4YD8_0),.clk(gclk));
	jdff dff_B_A8Lo3swX6_0(.din(w_dff_B_mFnNs4YD8_0),.dout(w_dff_B_A8Lo3swX6_0),.clk(gclk));
	jdff dff_B_LE03pELK4_0(.din(w_dff_B_A8Lo3swX6_0),.dout(w_dff_B_LE03pELK4_0),.clk(gclk));
	jdff dff_B_Lb21lxX88_0(.din(w_dff_B_LE03pELK4_0),.dout(w_dff_B_Lb21lxX88_0),.clk(gclk));
	jdff dff_B_1eUFobsA4_0(.din(w_dff_B_Lb21lxX88_0),.dout(w_dff_B_1eUFobsA4_0),.clk(gclk));
	jdff dff_B_5WtdonBp8_0(.din(w_dff_B_1eUFobsA4_0),.dout(w_dff_B_5WtdonBp8_0),.clk(gclk));
	jdff dff_B_vuYe2YEX1_0(.din(w_dff_B_5WtdonBp8_0),.dout(w_dff_B_vuYe2YEX1_0),.clk(gclk));
	jdff dff_B_Io1QzfOL0_0(.din(w_dff_B_vuYe2YEX1_0),.dout(w_dff_B_Io1QzfOL0_0),.clk(gclk));
	jdff dff_B_Q32EF3Z83_0(.din(w_dff_B_Io1QzfOL0_0),.dout(w_dff_B_Q32EF3Z83_0),.clk(gclk));
	jdff dff_B_sS1Du8u40_0(.din(w_dff_B_Q32EF3Z83_0),.dout(w_dff_B_sS1Du8u40_0),.clk(gclk));
	jdff dff_B_Ow6NRkMo4_0(.din(w_dff_B_sS1Du8u40_0),.dout(w_dff_B_Ow6NRkMo4_0),.clk(gclk));
	jdff dff_B_ew8IcJrQ3_0(.din(w_dff_B_Ow6NRkMo4_0),.dout(w_dff_B_ew8IcJrQ3_0),.clk(gclk));
	jdff dff_B_vgmPifxO3_0(.din(w_dff_B_ew8IcJrQ3_0),.dout(w_dff_B_vgmPifxO3_0),.clk(gclk));
	jdff dff_B_Cn1Ozxvh4_0(.din(w_dff_B_vgmPifxO3_0),.dout(w_dff_B_Cn1Ozxvh4_0),.clk(gclk));
	jdff dff_B_lzsM3vLa5_0(.din(w_dff_B_Cn1Ozxvh4_0),.dout(w_dff_B_lzsM3vLa5_0),.clk(gclk));
	jdff dff_B_mWy09Jvh2_0(.din(w_dff_B_lzsM3vLa5_0),.dout(w_dff_B_mWy09Jvh2_0),.clk(gclk));
	jdff dff_B_e3BiTXmW2_0(.din(w_dff_B_mWy09Jvh2_0),.dout(w_dff_B_e3BiTXmW2_0),.clk(gclk));
	jdff dff_B_v9og7iuP2_0(.din(w_dff_B_e3BiTXmW2_0),.dout(w_dff_B_v9og7iuP2_0),.clk(gclk));
	jdff dff_B_r5gEe0757_0(.din(w_dff_B_v9og7iuP2_0),.dout(w_dff_B_r5gEe0757_0),.clk(gclk));
	jdff dff_B_Fe0B8YFI0_0(.din(w_dff_B_r5gEe0757_0),.dout(w_dff_B_Fe0B8YFI0_0),.clk(gclk));
	jdff dff_B_LfvVBueY0_1(.din(n630),.dout(w_dff_B_LfvVBueY0_1),.clk(gclk));
	jdff dff_B_NcKvCmdt5_1(.din(w_dff_B_LfvVBueY0_1),.dout(w_dff_B_NcKvCmdt5_1),.clk(gclk));
	jdff dff_B_DJ6o65Lq3_1(.din(w_dff_B_NcKvCmdt5_1),.dout(w_dff_B_DJ6o65Lq3_1),.clk(gclk));
	jdff dff_B_q0Psu5Uy0_1(.din(w_dff_B_DJ6o65Lq3_1),.dout(w_dff_B_q0Psu5Uy0_1),.clk(gclk));
	jdff dff_B_Je1FYDtC3_1(.din(w_dff_B_q0Psu5Uy0_1),.dout(w_dff_B_Je1FYDtC3_1),.clk(gclk));
	jdff dff_B_iFxXbCNx8_1(.din(w_dff_B_Je1FYDtC3_1),.dout(w_dff_B_iFxXbCNx8_1),.clk(gclk));
	jdff dff_B_oC44ZmXv2_1(.din(w_dff_B_iFxXbCNx8_1),.dout(w_dff_B_oC44ZmXv2_1),.clk(gclk));
	jdff dff_B_uinjqs4z6_1(.din(w_dff_B_oC44ZmXv2_1),.dout(w_dff_B_uinjqs4z6_1),.clk(gclk));
	jdff dff_B_pDoJZss74_1(.din(w_dff_B_uinjqs4z6_1),.dout(w_dff_B_pDoJZss74_1),.clk(gclk));
	jdff dff_B_5SihKAo75_1(.din(w_dff_B_pDoJZss74_1),.dout(w_dff_B_5SihKAo75_1),.clk(gclk));
	jdff dff_B_JRksUubY9_1(.din(w_dff_B_5SihKAo75_1),.dout(w_dff_B_JRksUubY9_1),.clk(gclk));
	jdff dff_B_nJegQheD2_1(.din(w_dff_B_JRksUubY9_1),.dout(w_dff_B_nJegQheD2_1),.clk(gclk));
	jdff dff_B_h87hwmAm7_1(.din(w_dff_B_nJegQheD2_1),.dout(w_dff_B_h87hwmAm7_1),.clk(gclk));
	jdff dff_B_DB7syB5h6_1(.din(w_dff_B_h87hwmAm7_1),.dout(w_dff_B_DB7syB5h6_1),.clk(gclk));
	jdff dff_B_QQxYH7d35_1(.din(w_dff_B_DB7syB5h6_1),.dout(w_dff_B_QQxYH7d35_1),.clk(gclk));
	jdff dff_B_gWGgSwGM6_1(.din(w_dff_B_QQxYH7d35_1),.dout(w_dff_B_gWGgSwGM6_1),.clk(gclk));
	jdff dff_B_X5apSPjd9_1(.din(w_dff_B_gWGgSwGM6_1),.dout(w_dff_B_X5apSPjd9_1),.clk(gclk));
	jdff dff_B_8gCECxur4_1(.din(w_dff_B_X5apSPjd9_1),.dout(w_dff_B_8gCECxur4_1),.clk(gclk));
	jdff dff_B_6z21e0oO0_1(.din(w_dff_B_8gCECxur4_1),.dout(w_dff_B_6z21e0oO0_1),.clk(gclk));
	jdff dff_B_jdSjGdEz7_1(.din(w_dff_B_6z21e0oO0_1),.dout(w_dff_B_jdSjGdEz7_1),.clk(gclk));
	jdff dff_B_437FKpI84_1(.din(w_dff_B_jdSjGdEz7_1),.dout(w_dff_B_437FKpI84_1),.clk(gclk));
	jdff dff_B_wA7ZMEcc7_1(.din(w_dff_B_437FKpI84_1),.dout(w_dff_B_wA7ZMEcc7_1),.clk(gclk));
	jdff dff_B_H7zLB2vL5_1(.din(w_dff_B_wA7ZMEcc7_1),.dout(w_dff_B_H7zLB2vL5_1),.clk(gclk));
	jdff dff_B_ykok26La2_1(.din(w_dff_B_H7zLB2vL5_1),.dout(w_dff_B_ykok26La2_1),.clk(gclk));
	jdff dff_B_EsPOWioc0_1(.din(w_dff_B_ykok26La2_1),.dout(w_dff_B_EsPOWioc0_1),.clk(gclk));
	jdff dff_B_Kq9F65Lt1_1(.din(w_dff_B_EsPOWioc0_1),.dout(w_dff_B_Kq9F65Lt1_1),.clk(gclk));
	jdff dff_B_MkO2miZq2_1(.din(w_dff_B_Kq9F65Lt1_1),.dout(w_dff_B_MkO2miZq2_1),.clk(gclk));
	jdff dff_B_TElzeroM0_1(.din(w_dff_B_MkO2miZq2_1),.dout(w_dff_B_TElzeroM0_1),.clk(gclk));
	jdff dff_B_oQrqWhYX1_1(.din(w_dff_B_TElzeroM0_1),.dout(w_dff_B_oQrqWhYX1_1),.clk(gclk));
	jdff dff_B_iXFk4EJZ2_1(.din(w_dff_B_oQrqWhYX1_1),.dout(w_dff_B_iXFk4EJZ2_1),.clk(gclk));
	jdff dff_B_O8NN1KSx5_1(.din(w_dff_B_iXFk4EJZ2_1),.dout(w_dff_B_O8NN1KSx5_1),.clk(gclk));
	jdff dff_B_DM7PYOeZ4_1(.din(w_dff_B_O8NN1KSx5_1),.dout(w_dff_B_DM7PYOeZ4_1),.clk(gclk));
	jdff dff_B_9jHn0Qrs3_1(.din(w_dff_B_DM7PYOeZ4_1),.dout(w_dff_B_9jHn0Qrs3_1),.clk(gclk));
	jdff dff_B_xh44CqbF7_1(.din(w_dff_B_9jHn0Qrs3_1),.dout(w_dff_B_xh44CqbF7_1),.clk(gclk));
	jdff dff_B_4ChyFnB71_1(.din(w_dff_B_xh44CqbF7_1),.dout(w_dff_B_4ChyFnB71_1),.clk(gclk));
	jdff dff_B_lqlvHr5s5_1(.din(w_dff_B_4ChyFnB71_1),.dout(w_dff_B_lqlvHr5s5_1),.clk(gclk));
	jdff dff_B_aKvZTimR6_1(.din(w_dff_B_lqlvHr5s5_1),.dout(w_dff_B_aKvZTimR6_1),.clk(gclk));
	jdff dff_B_UfLN8bv23_1(.din(w_dff_B_aKvZTimR6_1),.dout(w_dff_B_UfLN8bv23_1),.clk(gclk));
	jdff dff_B_rNYfaluK9_1(.din(w_dff_B_UfLN8bv23_1),.dout(w_dff_B_rNYfaluK9_1),.clk(gclk));
	jdff dff_B_daPY71Er5_1(.din(w_dff_B_rNYfaluK9_1),.dout(w_dff_B_daPY71Er5_1),.clk(gclk));
	jdff dff_B_AyOrLbF03_1(.din(w_dff_B_daPY71Er5_1),.dout(w_dff_B_AyOrLbF03_1),.clk(gclk));
	jdff dff_B_8QmPIgxg7_0(.din(n631),.dout(w_dff_B_8QmPIgxg7_0),.clk(gclk));
	jdff dff_B_gdpXlBXN8_0(.din(w_dff_B_8QmPIgxg7_0),.dout(w_dff_B_gdpXlBXN8_0),.clk(gclk));
	jdff dff_B_AugFBj339_0(.din(w_dff_B_gdpXlBXN8_0),.dout(w_dff_B_AugFBj339_0),.clk(gclk));
	jdff dff_B_JC1E4JBT7_0(.din(w_dff_B_AugFBj339_0),.dout(w_dff_B_JC1E4JBT7_0),.clk(gclk));
	jdff dff_B_ymUm0FtD5_0(.din(w_dff_B_JC1E4JBT7_0),.dout(w_dff_B_ymUm0FtD5_0),.clk(gclk));
	jdff dff_B_57KJpRgz0_0(.din(w_dff_B_ymUm0FtD5_0),.dout(w_dff_B_57KJpRgz0_0),.clk(gclk));
	jdff dff_B_wtk4BUCI5_0(.din(w_dff_B_57KJpRgz0_0),.dout(w_dff_B_wtk4BUCI5_0),.clk(gclk));
	jdff dff_B_UpULRIn27_0(.din(w_dff_B_wtk4BUCI5_0),.dout(w_dff_B_UpULRIn27_0),.clk(gclk));
	jdff dff_B_AmpsyZsk8_0(.din(w_dff_B_UpULRIn27_0),.dout(w_dff_B_AmpsyZsk8_0),.clk(gclk));
	jdff dff_B_tmnkAl681_0(.din(w_dff_B_AmpsyZsk8_0),.dout(w_dff_B_tmnkAl681_0),.clk(gclk));
	jdff dff_B_JoB70bx69_0(.din(w_dff_B_tmnkAl681_0),.dout(w_dff_B_JoB70bx69_0),.clk(gclk));
	jdff dff_B_hMab1QwY0_0(.din(w_dff_B_JoB70bx69_0),.dout(w_dff_B_hMab1QwY0_0),.clk(gclk));
	jdff dff_B_4eDjRmk35_0(.din(w_dff_B_hMab1QwY0_0),.dout(w_dff_B_4eDjRmk35_0),.clk(gclk));
	jdff dff_B_iWtDPUc90_0(.din(w_dff_B_4eDjRmk35_0),.dout(w_dff_B_iWtDPUc90_0),.clk(gclk));
	jdff dff_B_qaMoqtoE5_0(.din(w_dff_B_iWtDPUc90_0),.dout(w_dff_B_qaMoqtoE5_0),.clk(gclk));
	jdff dff_B_RaTFKHR32_0(.din(w_dff_B_qaMoqtoE5_0),.dout(w_dff_B_RaTFKHR32_0),.clk(gclk));
	jdff dff_B_30aKGob80_0(.din(w_dff_B_RaTFKHR32_0),.dout(w_dff_B_30aKGob80_0),.clk(gclk));
	jdff dff_B_fErKBY4y9_0(.din(w_dff_B_30aKGob80_0),.dout(w_dff_B_fErKBY4y9_0),.clk(gclk));
	jdff dff_B_YzZSBsJV3_0(.din(w_dff_B_fErKBY4y9_0),.dout(w_dff_B_YzZSBsJV3_0),.clk(gclk));
	jdff dff_B_m6Ympzvr4_0(.din(w_dff_B_YzZSBsJV3_0),.dout(w_dff_B_m6Ympzvr4_0),.clk(gclk));
	jdff dff_B_2oURZFRQ9_0(.din(w_dff_B_m6Ympzvr4_0),.dout(w_dff_B_2oURZFRQ9_0),.clk(gclk));
	jdff dff_B_RtKZtlBg9_0(.din(w_dff_B_2oURZFRQ9_0),.dout(w_dff_B_RtKZtlBg9_0),.clk(gclk));
	jdff dff_B_mj71ook10_0(.din(w_dff_B_RtKZtlBg9_0),.dout(w_dff_B_mj71ook10_0),.clk(gclk));
	jdff dff_B_2mmi0acZ2_0(.din(w_dff_B_mj71ook10_0),.dout(w_dff_B_2mmi0acZ2_0),.clk(gclk));
	jdff dff_B_bbiEC2Of8_0(.din(w_dff_B_2mmi0acZ2_0),.dout(w_dff_B_bbiEC2Of8_0),.clk(gclk));
	jdff dff_B_COsaEQCG9_0(.din(w_dff_B_bbiEC2Of8_0),.dout(w_dff_B_COsaEQCG9_0),.clk(gclk));
	jdff dff_B_yFeoltQO1_0(.din(w_dff_B_COsaEQCG9_0),.dout(w_dff_B_yFeoltQO1_0),.clk(gclk));
	jdff dff_B_TCUhTIcm8_0(.din(w_dff_B_yFeoltQO1_0),.dout(w_dff_B_TCUhTIcm8_0),.clk(gclk));
	jdff dff_B_o364N6ic5_0(.din(w_dff_B_TCUhTIcm8_0),.dout(w_dff_B_o364N6ic5_0),.clk(gclk));
	jdff dff_B_KWOueVoT5_0(.din(w_dff_B_o364N6ic5_0),.dout(w_dff_B_KWOueVoT5_0),.clk(gclk));
	jdff dff_B_I8390tJR1_0(.din(w_dff_B_KWOueVoT5_0),.dout(w_dff_B_I8390tJR1_0),.clk(gclk));
	jdff dff_B_kJwWrDQw3_0(.din(w_dff_B_I8390tJR1_0),.dout(w_dff_B_kJwWrDQw3_0),.clk(gclk));
	jdff dff_B_RHzLpNHa0_0(.din(w_dff_B_kJwWrDQw3_0),.dout(w_dff_B_RHzLpNHa0_0),.clk(gclk));
	jdff dff_B_bDxRWC8G9_0(.din(w_dff_B_RHzLpNHa0_0),.dout(w_dff_B_bDxRWC8G9_0),.clk(gclk));
	jdff dff_B_DvLBN5eN1_0(.din(w_dff_B_bDxRWC8G9_0),.dout(w_dff_B_DvLBN5eN1_0),.clk(gclk));
	jdff dff_B_D78bRx178_0(.din(w_dff_B_DvLBN5eN1_0),.dout(w_dff_B_D78bRx178_0),.clk(gclk));
	jdff dff_B_6zdCY1st4_0(.din(w_dff_B_D78bRx178_0),.dout(w_dff_B_6zdCY1st4_0),.clk(gclk));
	jdff dff_B_jrGRcu648_0(.din(w_dff_B_6zdCY1st4_0),.dout(w_dff_B_jrGRcu648_0),.clk(gclk));
	jdff dff_B_OjIGXFHP6_0(.din(w_dff_B_jrGRcu648_0),.dout(w_dff_B_OjIGXFHP6_0),.clk(gclk));
	jdff dff_B_LpJVmWzl0_0(.din(w_dff_B_OjIGXFHP6_0),.dout(w_dff_B_LpJVmWzl0_0),.clk(gclk));
	jdff dff_B_Vysb7cc73_0(.din(w_dff_B_LpJVmWzl0_0),.dout(w_dff_B_Vysb7cc73_0),.clk(gclk));
	jdff dff_B_JtBXUdKo9_1(.din(n624),.dout(w_dff_B_JtBXUdKo9_1),.clk(gclk));
	jdff dff_B_tnuR8YWP5_1(.din(w_dff_B_JtBXUdKo9_1),.dout(w_dff_B_tnuR8YWP5_1),.clk(gclk));
	jdff dff_B_ylFQdDCL4_1(.din(w_dff_B_tnuR8YWP5_1),.dout(w_dff_B_ylFQdDCL4_1),.clk(gclk));
	jdff dff_B_FEWVQ50k5_1(.din(w_dff_B_ylFQdDCL4_1),.dout(w_dff_B_FEWVQ50k5_1),.clk(gclk));
	jdff dff_B_l6SyDGht7_1(.din(w_dff_B_FEWVQ50k5_1),.dout(w_dff_B_l6SyDGht7_1),.clk(gclk));
	jdff dff_B_NJVX5EQd2_1(.din(w_dff_B_l6SyDGht7_1),.dout(w_dff_B_NJVX5EQd2_1),.clk(gclk));
	jdff dff_B_Snv4rtsR1_1(.din(w_dff_B_NJVX5EQd2_1),.dout(w_dff_B_Snv4rtsR1_1),.clk(gclk));
	jdff dff_B_XGof5jkU7_1(.din(w_dff_B_Snv4rtsR1_1),.dout(w_dff_B_XGof5jkU7_1),.clk(gclk));
	jdff dff_B_lX3DDY6P2_1(.din(w_dff_B_XGof5jkU7_1),.dout(w_dff_B_lX3DDY6P2_1),.clk(gclk));
	jdff dff_B_xrqOj9PN6_1(.din(w_dff_B_lX3DDY6P2_1),.dout(w_dff_B_xrqOj9PN6_1),.clk(gclk));
	jdff dff_B_6ijP604D0_1(.din(w_dff_B_xrqOj9PN6_1),.dout(w_dff_B_6ijP604D0_1),.clk(gclk));
	jdff dff_B_DsvsmWQi6_1(.din(w_dff_B_6ijP604D0_1),.dout(w_dff_B_DsvsmWQi6_1),.clk(gclk));
	jdff dff_B_MNC9zpYz2_1(.din(w_dff_B_DsvsmWQi6_1),.dout(w_dff_B_MNC9zpYz2_1),.clk(gclk));
	jdff dff_B_Bny0fsYb5_1(.din(w_dff_B_MNC9zpYz2_1),.dout(w_dff_B_Bny0fsYb5_1),.clk(gclk));
	jdff dff_B_9e1uVB6s3_1(.din(w_dff_B_Bny0fsYb5_1),.dout(w_dff_B_9e1uVB6s3_1),.clk(gclk));
	jdff dff_B_loMNqfOv9_1(.din(w_dff_B_9e1uVB6s3_1),.dout(w_dff_B_loMNqfOv9_1),.clk(gclk));
	jdff dff_B_Y1r64aQ38_1(.din(w_dff_B_loMNqfOv9_1),.dout(w_dff_B_Y1r64aQ38_1),.clk(gclk));
	jdff dff_B_9qjEfqHL5_1(.din(w_dff_B_Y1r64aQ38_1),.dout(w_dff_B_9qjEfqHL5_1),.clk(gclk));
	jdff dff_B_1mpgSUft4_1(.din(w_dff_B_9qjEfqHL5_1),.dout(w_dff_B_1mpgSUft4_1),.clk(gclk));
	jdff dff_B_eZTibyd20_1(.din(w_dff_B_1mpgSUft4_1),.dout(w_dff_B_eZTibyd20_1),.clk(gclk));
	jdff dff_B_vnDv5Lrd5_1(.din(w_dff_B_eZTibyd20_1),.dout(w_dff_B_vnDv5Lrd5_1),.clk(gclk));
	jdff dff_B_XJpXZniX4_1(.din(w_dff_B_vnDv5Lrd5_1),.dout(w_dff_B_XJpXZniX4_1),.clk(gclk));
	jdff dff_B_j8My0uqp8_1(.din(w_dff_B_XJpXZniX4_1),.dout(w_dff_B_j8My0uqp8_1),.clk(gclk));
	jdff dff_B_CKDDbEDM3_1(.din(w_dff_B_j8My0uqp8_1),.dout(w_dff_B_CKDDbEDM3_1),.clk(gclk));
	jdff dff_B_YZortXJx0_1(.din(w_dff_B_CKDDbEDM3_1),.dout(w_dff_B_YZortXJx0_1),.clk(gclk));
	jdff dff_B_PZV5GHdW1_1(.din(w_dff_B_YZortXJx0_1),.dout(w_dff_B_PZV5GHdW1_1),.clk(gclk));
	jdff dff_B_J6hPIZzi6_1(.din(w_dff_B_PZV5GHdW1_1),.dout(w_dff_B_J6hPIZzi6_1),.clk(gclk));
	jdff dff_B_QuZ4fmUX1_1(.din(w_dff_B_J6hPIZzi6_1),.dout(w_dff_B_QuZ4fmUX1_1),.clk(gclk));
	jdff dff_B_nbjg4KOP4_1(.din(w_dff_B_QuZ4fmUX1_1),.dout(w_dff_B_nbjg4KOP4_1),.clk(gclk));
	jdff dff_B_LH6xMYq93_1(.din(w_dff_B_nbjg4KOP4_1),.dout(w_dff_B_LH6xMYq93_1),.clk(gclk));
	jdff dff_B_7kXgOwiy2_1(.din(w_dff_B_LH6xMYq93_1),.dout(w_dff_B_7kXgOwiy2_1),.clk(gclk));
	jdff dff_B_gocHhJhU6_1(.din(w_dff_B_7kXgOwiy2_1),.dout(w_dff_B_gocHhJhU6_1),.clk(gclk));
	jdff dff_B_4RytfaR86_1(.din(w_dff_B_gocHhJhU6_1),.dout(w_dff_B_4RytfaR86_1),.clk(gclk));
	jdff dff_B_wRNdkMcH9_1(.din(w_dff_B_4RytfaR86_1),.dout(w_dff_B_wRNdkMcH9_1),.clk(gclk));
	jdff dff_B_0GN34qzU1_1(.din(w_dff_B_wRNdkMcH9_1),.dout(w_dff_B_0GN34qzU1_1),.clk(gclk));
	jdff dff_B_LaLGX4Cn7_1(.din(w_dff_B_0GN34qzU1_1),.dout(w_dff_B_LaLGX4Cn7_1),.clk(gclk));
	jdff dff_B_Ihdgu3SC3_1(.din(w_dff_B_LaLGX4Cn7_1),.dout(w_dff_B_Ihdgu3SC3_1),.clk(gclk));
	jdff dff_B_NcT0vIXU4_1(.din(w_dff_B_Ihdgu3SC3_1),.dout(w_dff_B_NcT0vIXU4_1),.clk(gclk));
	jdff dff_B_2FaxzmXI9_1(.din(w_dff_B_NcT0vIXU4_1),.dout(w_dff_B_2FaxzmXI9_1),.clk(gclk));
	jdff dff_B_snRizMBV3_1(.din(w_dff_B_2FaxzmXI9_1),.dout(w_dff_B_snRizMBV3_1),.clk(gclk));
	jdff dff_B_o8mfxGyU6_0(.din(n625),.dout(w_dff_B_o8mfxGyU6_0),.clk(gclk));
	jdff dff_B_PUPElYb84_0(.din(w_dff_B_o8mfxGyU6_0),.dout(w_dff_B_PUPElYb84_0),.clk(gclk));
	jdff dff_B_dLpcJHua6_0(.din(w_dff_B_PUPElYb84_0),.dout(w_dff_B_dLpcJHua6_0),.clk(gclk));
	jdff dff_B_TkbtOCnL5_0(.din(w_dff_B_dLpcJHua6_0),.dout(w_dff_B_TkbtOCnL5_0),.clk(gclk));
	jdff dff_B_fDi3aK9J6_0(.din(w_dff_B_TkbtOCnL5_0),.dout(w_dff_B_fDi3aK9J6_0),.clk(gclk));
	jdff dff_B_Ul0Z20f02_0(.din(w_dff_B_fDi3aK9J6_0),.dout(w_dff_B_Ul0Z20f02_0),.clk(gclk));
	jdff dff_B_1sqn5kY48_0(.din(w_dff_B_Ul0Z20f02_0),.dout(w_dff_B_1sqn5kY48_0),.clk(gclk));
	jdff dff_B_zTtg9Q927_0(.din(w_dff_B_1sqn5kY48_0),.dout(w_dff_B_zTtg9Q927_0),.clk(gclk));
	jdff dff_B_AqwG4Rta1_0(.din(w_dff_B_zTtg9Q927_0),.dout(w_dff_B_AqwG4Rta1_0),.clk(gclk));
	jdff dff_B_poKcUpzJ3_0(.din(w_dff_B_AqwG4Rta1_0),.dout(w_dff_B_poKcUpzJ3_0),.clk(gclk));
	jdff dff_B_X6h0VplD7_0(.din(w_dff_B_poKcUpzJ3_0),.dout(w_dff_B_X6h0VplD7_0),.clk(gclk));
	jdff dff_B_RNKjgaXI1_0(.din(w_dff_B_X6h0VplD7_0),.dout(w_dff_B_RNKjgaXI1_0),.clk(gclk));
	jdff dff_B_oQRgSYB33_0(.din(w_dff_B_RNKjgaXI1_0),.dout(w_dff_B_oQRgSYB33_0),.clk(gclk));
	jdff dff_B_rm1TJM0X5_0(.din(w_dff_B_oQRgSYB33_0),.dout(w_dff_B_rm1TJM0X5_0),.clk(gclk));
	jdff dff_B_wKmXwpRf0_0(.din(w_dff_B_rm1TJM0X5_0),.dout(w_dff_B_wKmXwpRf0_0),.clk(gclk));
	jdff dff_B_iXGhHx0F6_0(.din(w_dff_B_wKmXwpRf0_0),.dout(w_dff_B_iXGhHx0F6_0),.clk(gclk));
	jdff dff_B_I4H8JLQ83_0(.din(w_dff_B_iXGhHx0F6_0),.dout(w_dff_B_I4H8JLQ83_0),.clk(gclk));
	jdff dff_B_xdM7t0hJ0_0(.din(w_dff_B_I4H8JLQ83_0),.dout(w_dff_B_xdM7t0hJ0_0),.clk(gclk));
	jdff dff_B_G7AG8Hem0_0(.din(w_dff_B_xdM7t0hJ0_0),.dout(w_dff_B_G7AG8Hem0_0),.clk(gclk));
	jdff dff_B_RWt0LnXB7_0(.din(w_dff_B_G7AG8Hem0_0),.dout(w_dff_B_RWt0LnXB7_0),.clk(gclk));
	jdff dff_B_U1BaAeiV1_0(.din(w_dff_B_RWt0LnXB7_0),.dout(w_dff_B_U1BaAeiV1_0),.clk(gclk));
	jdff dff_B_TAUiwysf0_0(.din(w_dff_B_U1BaAeiV1_0),.dout(w_dff_B_TAUiwysf0_0),.clk(gclk));
	jdff dff_B_m61JRhu45_0(.din(w_dff_B_TAUiwysf0_0),.dout(w_dff_B_m61JRhu45_0),.clk(gclk));
	jdff dff_B_D0X3Pn096_0(.din(w_dff_B_m61JRhu45_0),.dout(w_dff_B_D0X3Pn096_0),.clk(gclk));
	jdff dff_B_QdgAXuHb7_0(.din(w_dff_B_D0X3Pn096_0),.dout(w_dff_B_QdgAXuHb7_0),.clk(gclk));
	jdff dff_B_TMJA1A3w8_0(.din(w_dff_B_QdgAXuHb7_0),.dout(w_dff_B_TMJA1A3w8_0),.clk(gclk));
	jdff dff_B_XhNtbCfn9_0(.din(w_dff_B_TMJA1A3w8_0),.dout(w_dff_B_XhNtbCfn9_0),.clk(gclk));
	jdff dff_B_4zRtAuoH9_0(.din(w_dff_B_XhNtbCfn9_0),.dout(w_dff_B_4zRtAuoH9_0),.clk(gclk));
	jdff dff_B_dAH1Q7QK9_0(.din(w_dff_B_4zRtAuoH9_0),.dout(w_dff_B_dAH1Q7QK9_0),.clk(gclk));
	jdff dff_B_19RreQQs1_0(.din(w_dff_B_dAH1Q7QK9_0),.dout(w_dff_B_19RreQQs1_0),.clk(gclk));
	jdff dff_B_94366zT98_0(.din(w_dff_B_19RreQQs1_0),.dout(w_dff_B_94366zT98_0),.clk(gclk));
	jdff dff_B_juOMJ1AY3_0(.din(w_dff_B_94366zT98_0),.dout(w_dff_B_juOMJ1AY3_0),.clk(gclk));
	jdff dff_B_aA85Jycj4_0(.din(w_dff_B_juOMJ1AY3_0),.dout(w_dff_B_aA85Jycj4_0),.clk(gclk));
	jdff dff_B_5fCnl3QD9_0(.din(w_dff_B_aA85Jycj4_0),.dout(w_dff_B_5fCnl3QD9_0),.clk(gclk));
	jdff dff_B_qXgoHIwS3_0(.din(w_dff_B_5fCnl3QD9_0),.dout(w_dff_B_qXgoHIwS3_0),.clk(gclk));
	jdff dff_B_nBYX7AaE3_0(.din(w_dff_B_qXgoHIwS3_0),.dout(w_dff_B_nBYX7AaE3_0),.clk(gclk));
	jdff dff_B_7BmlLgs43_0(.din(w_dff_B_nBYX7AaE3_0),.dout(w_dff_B_7BmlLgs43_0),.clk(gclk));
	jdff dff_B_pBBtc8UM7_0(.din(w_dff_B_7BmlLgs43_0),.dout(w_dff_B_pBBtc8UM7_0),.clk(gclk));
	jdff dff_B_6O2Govit3_0(.din(w_dff_B_pBBtc8UM7_0),.dout(w_dff_B_6O2Govit3_0),.clk(gclk));
	jdff dff_B_v6JmAK7j4_0(.din(w_dff_B_6O2Govit3_0),.dout(w_dff_B_v6JmAK7j4_0),.clk(gclk));
	jdff dff_B_xzNs3A4M6_1(.din(n618),.dout(w_dff_B_xzNs3A4M6_1),.clk(gclk));
	jdff dff_B_s01y1Wtc1_1(.din(w_dff_B_xzNs3A4M6_1),.dout(w_dff_B_s01y1Wtc1_1),.clk(gclk));
	jdff dff_B_wCtWxCcz4_1(.din(w_dff_B_s01y1Wtc1_1),.dout(w_dff_B_wCtWxCcz4_1),.clk(gclk));
	jdff dff_B_8yP6upqU5_1(.din(w_dff_B_wCtWxCcz4_1),.dout(w_dff_B_8yP6upqU5_1),.clk(gclk));
	jdff dff_B_C5GJfc6h0_1(.din(w_dff_B_8yP6upqU5_1),.dout(w_dff_B_C5GJfc6h0_1),.clk(gclk));
	jdff dff_B_8tpjvD302_1(.din(w_dff_B_C5GJfc6h0_1),.dout(w_dff_B_8tpjvD302_1),.clk(gclk));
	jdff dff_B_qaTYaa3Z7_1(.din(w_dff_B_8tpjvD302_1),.dout(w_dff_B_qaTYaa3Z7_1),.clk(gclk));
	jdff dff_B_6DXjRWWV4_1(.din(w_dff_B_qaTYaa3Z7_1),.dout(w_dff_B_6DXjRWWV4_1),.clk(gclk));
	jdff dff_B_7yuGZxwu6_1(.din(w_dff_B_6DXjRWWV4_1),.dout(w_dff_B_7yuGZxwu6_1),.clk(gclk));
	jdff dff_B_irM2ab3R0_1(.din(w_dff_B_7yuGZxwu6_1),.dout(w_dff_B_irM2ab3R0_1),.clk(gclk));
	jdff dff_B_psde5juB8_1(.din(w_dff_B_irM2ab3R0_1),.dout(w_dff_B_psde5juB8_1),.clk(gclk));
	jdff dff_B_O2O1igCC1_1(.din(w_dff_B_psde5juB8_1),.dout(w_dff_B_O2O1igCC1_1),.clk(gclk));
	jdff dff_B_HJPnBiZm2_1(.din(w_dff_B_O2O1igCC1_1),.dout(w_dff_B_HJPnBiZm2_1),.clk(gclk));
	jdff dff_B_LQo44HpF2_1(.din(w_dff_B_HJPnBiZm2_1),.dout(w_dff_B_LQo44HpF2_1),.clk(gclk));
	jdff dff_B_n7IBoHt73_1(.din(w_dff_B_LQo44HpF2_1),.dout(w_dff_B_n7IBoHt73_1),.clk(gclk));
	jdff dff_B_Nb6mRhav0_1(.din(w_dff_B_n7IBoHt73_1),.dout(w_dff_B_Nb6mRhav0_1),.clk(gclk));
	jdff dff_B_iVfYt3Xp8_1(.din(w_dff_B_Nb6mRhav0_1),.dout(w_dff_B_iVfYt3Xp8_1),.clk(gclk));
	jdff dff_B_x1f5z0VI7_1(.din(w_dff_B_iVfYt3Xp8_1),.dout(w_dff_B_x1f5z0VI7_1),.clk(gclk));
	jdff dff_B_51nqEt9r5_1(.din(w_dff_B_x1f5z0VI7_1),.dout(w_dff_B_51nqEt9r5_1),.clk(gclk));
	jdff dff_B_HChZ5S6X1_1(.din(w_dff_B_51nqEt9r5_1),.dout(w_dff_B_HChZ5S6X1_1),.clk(gclk));
	jdff dff_B_KKocAJDS9_1(.din(w_dff_B_HChZ5S6X1_1),.dout(w_dff_B_KKocAJDS9_1),.clk(gclk));
	jdff dff_B_xANEwfpg5_1(.din(w_dff_B_KKocAJDS9_1),.dout(w_dff_B_xANEwfpg5_1),.clk(gclk));
	jdff dff_B_N9aBp7x86_1(.din(w_dff_B_xANEwfpg5_1),.dout(w_dff_B_N9aBp7x86_1),.clk(gclk));
	jdff dff_B_rjpQ0Vrr7_1(.din(w_dff_B_N9aBp7x86_1),.dout(w_dff_B_rjpQ0Vrr7_1),.clk(gclk));
	jdff dff_B_eVLvNr9U2_1(.din(w_dff_B_rjpQ0Vrr7_1),.dout(w_dff_B_eVLvNr9U2_1),.clk(gclk));
	jdff dff_B_wzZLjjXc3_1(.din(w_dff_B_eVLvNr9U2_1),.dout(w_dff_B_wzZLjjXc3_1),.clk(gclk));
	jdff dff_B_LCB8nkvn4_1(.din(w_dff_B_wzZLjjXc3_1),.dout(w_dff_B_LCB8nkvn4_1),.clk(gclk));
	jdff dff_B_IaVkYITB1_1(.din(w_dff_B_LCB8nkvn4_1),.dout(w_dff_B_IaVkYITB1_1),.clk(gclk));
	jdff dff_B_TJtf2OrS3_1(.din(w_dff_B_IaVkYITB1_1),.dout(w_dff_B_TJtf2OrS3_1),.clk(gclk));
	jdff dff_B_4shiWAZO0_1(.din(w_dff_B_TJtf2OrS3_1),.dout(w_dff_B_4shiWAZO0_1),.clk(gclk));
	jdff dff_B_TX61vdvN2_1(.din(w_dff_B_4shiWAZO0_1),.dout(w_dff_B_TX61vdvN2_1),.clk(gclk));
	jdff dff_B_NEYiPyj59_1(.din(w_dff_B_TX61vdvN2_1),.dout(w_dff_B_NEYiPyj59_1),.clk(gclk));
	jdff dff_B_wCBlSHfj3_1(.din(w_dff_B_NEYiPyj59_1),.dout(w_dff_B_wCBlSHfj3_1),.clk(gclk));
	jdff dff_B_gp754SI74_1(.din(w_dff_B_wCBlSHfj3_1),.dout(w_dff_B_gp754SI74_1),.clk(gclk));
	jdff dff_B_5KZNcjZo2_1(.din(w_dff_B_gp754SI74_1),.dout(w_dff_B_5KZNcjZo2_1),.clk(gclk));
	jdff dff_B_ojL8Y5TK5_1(.din(w_dff_B_5KZNcjZo2_1),.dout(w_dff_B_ojL8Y5TK5_1),.clk(gclk));
	jdff dff_B_URhAnzRc0_1(.din(w_dff_B_ojL8Y5TK5_1),.dout(w_dff_B_URhAnzRc0_1),.clk(gclk));
	jdff dff_B_84Hiap2m8_1(.din(w_dff_B_URhAnzRc0_1),.dout(w_dff_B_84Hiap2m8_1),.clk(gclk));
	jdff dff_B_1cZChDiV8_1(.din(w_dff_B_84Hiap2m8_1),.dout(w_dff_B_1cZChDiV8_1),.clk(gclk));
	jdff dff_B_i5VTpo2H0_0(.din(n619),.dout(w_dff_B_i5VTpo2H0_0),.clk(gclk));
	jdff dff_B_RQmDHBCp0_0(.din(w_dff_B_i5VTpo2H0_0),.dout(w_dff_B_RQmDHBCp0_0),.clk(gclk));
	jdff dff_B_rvxlBOtD2_0(.din(w_dff_B_RQmDHBCp0_0),.dout(w_dff_B_rvxlBOtD2_0),.clk(gclk));
	jdff dff_B_yqNj9LDA3_0(.din(w_dff_B_rvxlBOtD2_0),.dout(w_dff_B_yqNj9LDA3_0),.clk(gclk));
	jdff dff_B_RIATV5hH1_0(.din(w_dff_B_yqNj9LDA3_0),.dout(w_dff_B_RIATV5hH1_0),.clk(gclk));
	jdff dff_B_jMsOL3vp7_0(.din(w_dff_B_RIATV5hH1_0),.dout(w_dff_B_jMsOL3vp7_0),.clk(gclk));
	jdff dff_B_r9zowARR0_0(.din(w_dff_B_jMsOL3vp7_0),.dout(w_dff_B_r9zowARR0_0),.clk(gclk));
	jdff dff_B_Zg4iFbBX0_0(.din(w_dff_B_r9zowARR0_0),.dout(w_dff_B_Zg4iFbBX0_0),.clk(gclk));
	jdff dff_B_lCXmiMOp9_0(.din(w_dff_B_Zg4iFbBX0_0),.dout(w_dff_B_lCXmiMOp9_0),.clk(gclk));
	jdff dff_B_g4UFrxPP1_0(.din(w_dff_B_lCXmiMOp9_0),.dout(w_dff_B_g4UFrxPP1_0),.clk(gclk));
	jdff dff_B_jFPiEOD57_0(.din(w_dff_B_g4UFrxPP1_0),.dout(w_dff_B_jFPiEOD57_0),.clk(gclk));
	jdff dff_B_QMMJIS8c6_0(.din(w_dff_B_jFPiEOD57_0),.dout(w_dff_B_QMMJIS8c6_0),.clk(gclk));
	jdff dff_B_4lmsmhQq7_0(.din(w_dff_B_QMMJIS8c6_0),.dout(w_dff_B_4lmsmhQq7_0),.clk(gclk));
	jdff dff_B_bCrYGWew7_0(.din(w_dff_B_4lmsmhQq7_0),.dout(w_dff_B_bCrYGWew7_0),.clk(gclk));
	jdff dff_B_GK3lBu273_0(.din(w_dff_B_bCrYGWew7_0),.dout(w_dff_B_GK3lBu273_0),.clk(gclk));
	jdff dff_B_Bgr8ryv43_0(.din(w_dff_B_GK3lBu273_0),.dout(w_dff_B_Bgr8ryv43_0),.clk(gclk));
	jdff dff_B_0ltDi3rS8_0(.din(w_dff_B_Bgr8ryv43_0),.dout(w_dff_B_0ltDi3rS8_0),.clk(gclk));
	jdff dff_B_bedNWeIh6_0(.din(w_dff_B_0ltDi3rS8_0),.dout(w_dff_B_bedNWeIh6_0),.clk(gclk));
	jdff dff_B_CZhY63wi9_0(.din(w_dff_B_bedNWeIh6_0),.dout(w_dff_B_CZhY63wi9_0),.clk(gclk));
	jdff dff_B_6AxVyPtV2_0(.din(w_dff_B_CZhY63wi9_0),.dout(w_dff_B_6AxVyPtV2_0),.clk(gclk));
	jdff dff_B_o4vlHLg51_0(.din(w_dff_B_6AxVyPtV2_0),.dout(w_dff_B_o4vlHLg51_0),.clk(gclk));
	jdff dff_B_ejQ3axLP1_0(.din(w_dff_B_o4vlHLg51_0),.dout(w_dff_B_ejQ3axLP1_0),.clk(gclk));
	jdff dff_B_pj9IPYEV4_0(.din(w_dff_B_ejQ3axLP1_0),.dout(w_dff_B_pj9IPYEV4_0),.clk(gclk));
	jdff dff_B_YC3DZGqd5_0(.din(w_dff_B_pj9IPYEV4_0),.dout(w_dff_B_YC3DZGqd5_0),.clk(gclk));
	jdff dff_B_p7v87gs65_0(.din(w_dff_B_YC3DZGqd5_0),.dout(w_dff_B_p7v87gs65_0),.clk(gclk));
	jdff dff_B_Q1FbSoin3_0(.din(w_dff_B_p7v87gs65_0),.dout(w_dff_B_Q1FbSoin3_0),.clk(gclk));
	jdff dff_B_Isxlw9op1_0(.din(w_dff_B_Q1FbSoin3_0),.dout(w_dff_B_Isxlw9op1_0),.clk(gclk));
	jdff dff_B_GEdcbSpu6_0(.din(w_dff_B_Isxlw9op1_0),.dout(w_dff_B_GEdcbSpu6_0),.clk(gclk));
	jdff dff_B_9UGnkm8S6_0(.din(w_dff_B_GEdcbSpu6_0),.dout(w_dff_B_9UGnkm8S6_0),.clk(gclk));
	jdff dff_B_ul4Emnel7_0(.din(w_dff_B_9UGnkm8S6_0),.dout(w_dff_B_ul4Emnel7_0),.clk(gclk));
	jdff dff_B_mReWuBRi7_0(.din(w_dff_B_ul4Emnel7_0),.dout(w_dff_B_mReWuBRi7_0),.clk(gclk));
	jdff dff_B_80BJIkHo9_0(.din(w_dff_B_mReWuBRi7_0),.dout(w_dff_B_80BJIkHo9_0),.clk(gclk));
	jdff dff_B_qhgaY1TM3_0(.din(w_dff_B_80BJIkHo9_0),.dout(w_dff_B_qhgaY1TM3_0),.clk(gclk));
	jdff dff_B_h0ypPEU98_0(.din(w_dff_B_qhgaY1TM3_0),.dout(w_dff_B_h0ypPEU98_0),.clk(gclk));
	jdff dff_B_4waKMxF29_0(.din(w_dff_B_h0ypPEU98_0),.dout(w_dff_B_4waKMxF29_0),.clk(gclk));
	jdff dff_B_TAYMfE5T9_0(.din(w_dff_B_4waKMxF29_0),.dout(w_dff_B_TAYMfE5T9_0),.clk(gclk));
	jdff dff_B_CwvfHwiR1_0(.din(w_dff_B_TAYMfE5T9_0),.dout(w_dff_B_CwvfHwiR1_0),.clk(gclk));
	jdff dff_B_l4zQADy20_0(.din(w_dff_B_CwvfHwiR1_0),.dout(w_dff_B_l4zQADy20_0),.clk(gclk));
	jdff dff_B_GoygnPeZ7_0(.din(w_dff_B_l4zQADy20_0),.dout(w_dff_B_GoygnPeZ7_0),.clk(gclk));
	jdff dff_B_iOAW5AkF8_1(.din(n612),.dout(w_dff_B_iOAW5AkF8_1),.clk(gclk));
	jdff dff_B_9L0ukpX21_1(.din(w_dff_B_iOAW5AkF8_1),.dout(w_dff_B_9L0ukpX21_1),.clk(gclk));
	jdff dff_B_bwvSSOEo8_1(.din(w_dff_B_9L0ukpX21_1),.dout(w_dff_B_bwvSSOEo8_1),.clk(gclk));
	jdff dff_B_ROFAGxLi7_1(.din(w_dff_B_bwvSSOEo8_1),.dout(w_dff_B_ROFAGxLi7_1),.clk(gclk));
	jdff dff_B_jT6Ym0JL5_1(.din(w_dff_B_ROFAGxLi7_1),.dout(w_dff_B_jT6Ym0JL5_1),.clk(gclk));
	jdff dff_B_SqxwqfOG2_1(.din(w_dff_B_jT6Ym0JL5_1),.dout(w_dff_B_SqxwqfOG2_1),.clk(gclk));
	jdff dff_B_cLvbRdyC2_1(.din(w_dff_B_SqxwqfOG2_1),.dout(w_dff_B_cLvbRdyC2_1),.clk(gclk));
	jdff dff_B_7bK7jhrl1_1(.din(w_dff_B_cLvbRdyC2_1),.dout(w_dff_B_7bK7jhrl1_1),.clk(gclk));
	jdff dff_B_ckTpkfs12_1(.din(w_dff_B_7bK7jhrl1_1),.dout(w_dff_B_ckTpkfs12_1),.clk(gclk));
	jdff dff_B_Pb7DM3cE3_1(.din(w_dff_B_ckTpkfs12_1),.dout(w_dff_B_Pb7DM3cE3_1),.clk(gclk));
	jdff dff_B_3g2H9eTP3_1(.din(w_dff_B_Pb7DM3cE3_1),.dout(w_dff_B_3g2H9eTP3_1),.clk(gclk));
	jdff dff_B_coVYVmSq1_1(.din(w_dff_B_3g2H9eTP3_1),.dout(w_dff_B_coVYVmSq1_1),.clk(gclk));
	jdff dff_B_6odMHASB8_1(.din(w_dff_B_coVYVmSq1_1),.dout(w_dff_B_6odMHASB8_1),.clk(gclk));
	jdff dff_B_VFhPuvlR3_1(.din(w_dff_B_6odMHASB8_1),.dout(w_dff_B_VFhPuvlR3_1),.clk(gclk));
	jdff dff_B_u2oY7gAH2_1(.din(w_dff_B_VFhPuvlR3_1),.dout(w_dff_B_u2oY7gAH2_1),.clk(gclk));
	jdff dff_B_eNekqtlL6_1(.din(w_dff_B_u2oY7gAH2_1),.dout(w_dff_B_eNekqtlL6_1),.clk(gclk));
	jdff dff_B_0vTuaUAb2_1(.din(w_dff_B_eNekqtlL6_1),.dout(w_dff_B_0vTuaUAb2_1),.clk(gclk));
	jdff dff_B_bC4I7ru02_1(.din(w_dff_B_0vTuaUAb2_1),.dout(w_dff_B_bC4I7ru02_1),.clk(gclk));
	jdff dff_B_5uaozvxf7_1(.din(w_dff_B_bC4I7ru02_1),.dout(w_dff_B_5uaozvxf7_1),.clk(gclk));
	jdff dff_B_cZmWyixe1_1(.din(w_dff_B_5uaozvxf7_1),.dout(w_dff_B_cZmWyixe1_1),.clk(gclk));
	jdff dff_B_2Mq98epl1_1(.din(w_dff_B_cZmWyixe1_1),.dout(w_dff_B_2Mq98epl1_1),.clk(gclk));
	jdff dff_B_DVyKpPt54_1(.din(w_dff_B_2Mq98epl1_1),.dout(w_dff_B_DVyKpPt54_1),.clk(gclk));
	jdff dff_B_Ug8Xamma4_1(.din(w_dff_B_DVyKpPt54_1),.dout(w_dff_B_Ug8Xamma4_1),.clk(gclk));
	jdff dff_B_zWjkUzMy5_1(.din(w_dff_B_Ug8Xamma4_1),.dout(w_dff_B_zWjkUzMy5_1),.clk(gclk));
	jdff dff_B_LTJcstDk5_1(.din(w_dff_B_zWjkUzMy5_1),.dout(w_dff_B_LTJcstDk5_1),.clk(gclk));
	jdff dff_B_3tjs6x592_1(.din(w_dff_B_LTJcstDk5_1),.dout(w_dff_B_3tjs6x592_1),.clk(gclk));
	jdff dff_B_ONjHRyg59_1(.din(w_dff_B_3tjs6x592_1),.dout(w_dff_B_ONjHRyg59_1),.clk(gclk));
	jdff dff_B_9PreDRWH4_1(.din(w_dff_B_ONjHRyg59_1),.dout(w_dff_B_9PreDRWH4_1),.clk(gclk));
	jdff dff_B_xPSeyFCx0_1(.din(w_dff_B_9PreDRWH4_1),.dout(w_dff_B_xPSeyFCx0_1),.clk(gclk));
	jdff dff_B_xdN6Hr634_1(.din(w_dff_B_xPSeyFCx0_1),.dout(w_dff_B_xdN6Hr634_1),.clk(gclk));
	jdff dff_B_wNfL7A9v3_1(.din(w_dff_B_xdN6Hr634_1),.dout(w_dff_B_wNfL7A9v3_1),.clk(gclk));
	jdff dff_B_l18RPvVU6_1(.din(w_dff_B_wNfL7A9v3_1),.dout(w_dff_B_l18RPvVU6_1),.clk(gclk));
	jdff dff_B_TO7PzIaj3_1(.din(w_dff_B_l18RPvVU6_1),.dout(w_dff_B_TO7PzIaj3_1),.clk(gclk));
	jdff dff_B_bipiOQLK9_1(.din(w_dff_B_TO7PzIaj3_1),.dout(w_dff_B_bipiOQLK9_1),.clk(gclk));
	jdff dff_B_3s3EH4Fk3_1(.din(w_dff_B_bipiOQLK9_1),.dout(w_dff_B_3s3EH4Fk3_1),.clk(gclk));
	jdff dff_B_cycLBPrn5_1(.din(w_dff_B_3s3EH4Fk3_1),.dout(w_dff_B_cycLBPrn5_1),.clk(gclk));
	jdff dff_B_NHJKcyqZ4_1(.din(w_dff_B_cycLBPrn5_1),.dout(w_dff_B_NHJKcyqZ4_1),.clk(gclk));
	jdff dff_B_u1eB0U854_1(.din(w_dff_B_NHJKcyqZ4_1),.dout(w_dff_B_u1eB0U854_1),.clk(gclk));
	jdff dff_B_Z8jCkfZY6_0(.din(n613),.dout(w_dff_B_Z8jCkfZY6_0),.clk(gclk));
	jdff dff_B_Bt7Owyjw5_0(.din(w_dff_B_Z8jCkfZY6_0),.dout(w_dff_B_Bt7Owyjw5_0),.clk(gclk));
	jdff dff_B_TlvrmO933_0(.din(w_dff_B_Bt7Owyjw5_0),.dout(w_dff_B_TlvrmO933_0),.clk(gclk));
	jdff dff_B_LgIM5swc7_0(.din(w_dff_B_TlvrmO933_0),.dout(w_dff_B_LgIM5swc7_0),.clk(gclk));
	jdff dff_B_Cqf05TVk4_0(.din(w_dff_B_LgIM5swc7_0),.dout(w_dff_B_Cqf05TVk4_0),.clk(gclk));
	jdff dff_B_hD6wqKc17_0(.din(w_dff_B_Cqf05TVk4_0),.dout(w_dff_B_hD6wqKc17_0),.clk(gclk));
	jdff dff_B_aRhaC4cG6_0(.din(w_dff_B_hD6wqKc17_0),.dout(w_dff_B_aRhaC4cG6_0),.clk(gclk));
	jdff dff_B_3nAD1CKi8_0(.din(w_dff_B_aRhaC4cG6_0),.dout(w_dff_B_3nAD1CKi8_0),.clk(gclk));
	jdff dff_B_QOAJRXMM4_0(.din(w_dff_B_3nAD1CKi8_0),.dout(w_dff_B_QOAJRXMM4_0),.clk(gclk));
	jdff dff_B_76qjEiyE8_0(.din(w_dff_B_QOAJRXMM4_0),.dout(w_dff_B_76qjEiyE8_0),.clk(gclk));
	jdff dff_B_HRdRkrcI1_0(.din(w_dff_B_76qjEiyE8_0),.dout(w_dff_B_HRdRkrcI1_0),.clk(gclk));
	jdff dff_B_yhZHwnXK9_0(.din(w_dff_B_HRdRkrcI1_0),.dout(w_dff_B_yhZHwnXK9_0),.clk(gclk));
	jdff dff_B_B8um4RKu0_0(.din(w_dff_B_yhZHwnXK9_0),.dout(w_dff_B_B8um4RKu0_0),.clk(gclk));
	jdff dff_B_MBAOr4b09_0(.din(w_dff_B_B8um4RKu0_0),.dout(w_dff_B_MBAOr4b09_0),.clk(gclk));
	jdff dff_B_et7e8b3V1_0(.din(w_dff_B_MBAOr4b09_0),.dout(w_dff_B_et7e8b3V1_0),.clk(gclk));
	jdff dff_B_L0nYeOLq4_0(.din(w_dff_B_et7e8b3V1_0),.dout(w_dff_B_L0nYeOLq4_0),.clk(gclk));
	jdff dff_B_IqrIqAQr5_0(.din(w_dff_B_L0nYeOLq4_0),.dout(w_dff_B_IqrIqAQr5_0),.clk(gclk));
	jdff dff_B_UV6KRfwW4_0(.din(w_dff_B_IqrIqAQr5_0),.dout(w_dff_B_UV6KRfwW4_0),.clk(gclk));
	jdff dff_B_tFgU9Iza0_0(.din(w_dff_B_UV6KRfwW4_0),.dout(w_dff_B_tFgU9Iza0_0),.clk(gclk));
	jdff dff_B_L3DnhOEG3_0(.din(w_dff_B_tFgU9Iza0_0),.dout(w_dff_B_L3DnhOEG3_0),.clk(gclk));
	jdff dff_B_UsxwXYhk4_0(.din(w_dff_B_L3DnhOEG3_0),.dout(w_dff_B_UsxwXYhk4_0),.clk(gclk));
	jdff dff_B_zCxnUZ4G7_0(.din(w_dff_B_UsxwXYhk4_0),.dout(w_dff_B_zCxnUZ4G7_0),.clk(gclk));
	jdff dff_B_l5QxuTNN1_0(.din(w_dff_B_zCxnUZ4G7_0),.dout(w_dff_B_l5QxuTNN1_0),.clk(gclk));
	jdff dff_B_j8HtY50C2_0(.din(w_dff_B_l5QxuTNN1_0),.dout(w_dff_B_j8HtY50C2_0),.clk(gclk));
	jdff dff_B_A1hVmr8q2_0(.din(w_dff_B_j8HtY50C2_0),.dout(w_dff_B_A1hVmr8q2_0),.clk(gclk));
	jdff dff_B_b3bUlmRR2_0(.din(w_dff_B_A1hVmr8q2_0),.dout(w_dff_B_b3bUlmRR2_0),.clk(gclk));
	jdff dff_B_G1iaj4CP7_0(.din(w_dff_B_b3bUlmRR2_0),.dout(w_dff_B_G1iaj4CP7_0),.clk(gclk));
	jdff dff_B_8KVtQ9Jx0_0(.din(w_dff_B_G1iaj4CP7_0),.dout(w_dff_B_8KVtQ9Jx0_0),.clk(gclk));
	jdff dff_B_zVaeqir66_0(.din(w_dff_B_8KVtQ9Jx0_0),.dout(w_dff_B_zVaeqir66_0),.clk(gclk));
	jdff dff_B_X2EG9XJK3_0(.din(w_dff_B_zVaeqir66_0),.dout(w_dff_B_X2EG9XJK3_0),.clk(gclk));
	jdff dff_B_LD9DlGyG4_0(.din(w_dff_B_X2EG9XJK3_0),.dout(w_dff_B_LD9DlGyG4_0),.clk(gclk));
	jdff dff_B_wRbo9ZCb1_0(.din(w_dff_B_LD9DlGyG4_0),.dout(w_dff_B_wRbo9ZCb1_0),.clk(gclk));
	jdff dff_B_I2GqYFZV5_0(.din(w_dff_B_wRbo9ZCb1_0),.dout(w_dff_B_I2GqYFZV5_0),.clk(gclk));
	jdff dff_B_20nn7j327_0(.din(w_dff_B_I2GqYFZV5_0),.dout(w_dff_B_20nn7j327_0),.clk(gclk));
	jdff dff_B_m4ydpTvG5_0(.din(w_dff_B_20nn7j327_0),.dout(w_dff_B_m4ydpTvG5_0),.clk(gclk));
	jdff dff_B_4f0BJZaz9_0(.din(w_dff_B_m4ydpTvG5_0),.dout(w_dff_B_4f0BJZaz9_0),.clk(gclk));
	jdff dff_B_ccXyxJ5S1_0(.din(w_dff_B_4f0BJZaz9_0),.dout(w_dff_B_ccXyxJ5S1_0),.clk(gclk));
	jdff dff_B_wdau1vMx1_0(.din(w_dff_B_ccXyxJ5S1_0),.dout(w_dff_B_wdau1vMx1_0),.clk(gclk));
	jdff dff_B_f4hct7133_1(.din(n606),.dout(w_dff_B_f4hct7133_1),.clk(gclk));
	jdff dff_B_UXIyiguw6_1(.din(w_dff_B_f4hct7133_1),.dout(w_dff_B_UXIyiguw6_1),.clk(gclk));
	jdff dff_B_ozl04Lbd5_1(.din(w_dff_B_UXIyiguw6_1),.dout(w_dff_B_ozl04Lbd5_1),.clk(gclk));
	jdff dff_B_JJnQpDCe3_1(.din(w_dff_B_ozl04Lbd5_1),.dout(w_dff_B_JJnQpDCe3_1),.clk(gclk));
	jdff dff_B_20Iin53p2_1(.din(w_dff_B_JJnQpDCe3_1),.dout(w_dff_B_20Iin53p2_1),.clk(gclk));
	jdff dff_B_CPAQ9Htg8_1(.din(w_dff_B_20Iin53p2_1),.dout(w_dff_B_CPAQ9Htg8_1),.clk(gclk));
	jdff dff_B_bXOSEEV56_1(.din(w_dff_B_CPAQ9Htg8_1),.dout(w_dff_B_bXOSEEV56_1),.clk(gclk));
	jdff dff_B_mH2SAvxU1_1(.din(w_dff_B_bXOSEEV56_1),.dout(w_dff_B_mH2SAvxU1_1),.clk(gclk));
	jdff dff_B_MixDna5N6_1(.din(w_dff_B_mH2SAvxU1_1),.dout(w_dff_B_MixDna5N6_1),.clk(gclk));
	jdff dff_B_t8szfHZc6_1(.din(w_dff_B_MixDna5N6_1),.dout(w_dff_B_t8szfHZc6_1),.clk(gclk));
	jdff dff_B_lDBahBDa5_1(.din(w_dff_B_t8szfHZc6_1),.dout(w_dff_B_lDBahBDa5_1),.clk(gclk));
	jdff dff_B_Qc5i2W7l6_1(.din(w_dff_B_lDBahBDa5_1),.dout(w_dff_B_Qc5i2W7l6_1),.clk(gclk));
	jdff dff_B_jlMKZlRA4_1(.din(w_dff_B_Qc5i2W7l6_1),.dout(w_dff_B_jlMKZlRA4_1),.clk(gclk));
	jdff dff_B_HsOv0bM55_1(.din(w_dff_B_jlMKZlRA4_1),.dout(w_dff_B_HsOv0bM55_1),.clk(gclk));
	jdff dff_B_hcChzzT21_1(.din(w_dff_B_HsOv0bM55_1),.dout(w_dff_B_hcChzzT21_1),.clk(gclk));
	jdff dff_B_jOZWmHiB3_1(.din(w_dff_B_hcChzzT21_1),.dout(w_dff_B_jOZWmHiB3_1),.clk(gclk));
	jdff dff_B_6W51sSxp6_1(.din(w_dff_B_jOZWmHiB3_1),.dout(w_dff_B_6W51sSxp6_1),.clk(gclk));
	jdff dff_B_yVQvIEVZ7_1(.din(w_dff_B_6W51sSxp6_1),.dout(w_dff_B_yVQvIEVZ7_1),.clk(gclk));
	jdff dff_B_ctGeb99d9_1(.din(w_dff_B_yVQvIEVZ7_1),.dout(w_dff_B_ctGeb99d9_1),.clk(gclk));
	jdff dff_B_eUTnZ67z0_1(.din(w_dff_B_ctGeb99d9_1),.dout(w_dff_B_eUTnZ67z0_1),.clk(gclk));
	jdff dff_B_EEHIYTbk5_1(.din(w_dff_B_eUTnZ67z0_1),.dout(w_dff_B_EEHIYTbk5_1),.clk(gclk));
	jdff dff_B_jLjqArVF7_1(.din(w_dff_B_EEHIYTbk5_1),.dout(w_dff_B_jLjqArVF7_1),.clk(gclk));
	jdff dff_B_ycN4tM0G0_1(.din(w_dff_B_jLjqArVF7_1),.dout(w_dff_B_ycN4tM0G0_1),.clk(gclk));
	jdff dff_B_65HPNs7T0_1(.din(w_dff_B_ycN4tM0G0_1),.dout(w_dff_B_65HPNs7T0_1),.clk(gclk));
	jdff dff_B_2jEWg2ys7_1(.din(w_dff_B_65HPNs7T0_1),.dout(w_dff_B_2jEWg2ys7_1),.clk(gclk));
	jdff dff_B_ljjvTOLC3_1(.din(w_dff_B_2jEWg2ys7_1),.dout(w_dff_B_ljjvTOLC3_1),.clk(gclk));
	jdff dff_B_v3B2YGPr4_1(.din(w_dff_B_ljjvTOLC3_1),.dout(w_dff_B_v3B2YGPr4_1),.clk(gclk));
	jdff dff_B_IQ7KbHQ30_1(.din(w_dff_B_v3B2YGPr4_1),.dout(w_dff_B_IQ7KbHQ30_1),.clk(gclk));
	jdff dff_B_ihQOhxU36_1(.din(w_dff_B_IQ7KbHQ30_1),.dout(w_dff_B_ihQOhxU36_1),.clk(gclk));
	jdff dff_B_U1veCSAc6_1(.din(w_dff_B_ihQOhxU36_1),.dout(w_dff_B_U1veCSAc6_1),.clk(gclk));
	jdff dff_B_X53RkT039_1(.din(w_dff_B_U1veCSAc6_1),.dout(w_dff_B_X53RkT039_1),.clk(gclk));
	jdff dff_B_MRkHPJkR3_1(.din(w_dff_B_X53RkT039_1),.dout(w_dff_B_MRkHPJkR3_1),.clk(gclk));
	jdff dff_B_uxWcVFyM7_1(.din(w_dff_B_MRkHPJkR3_1),.dout(w_dff_B_uxWcVFyM7_1),.clk(gclk));
	jdff dff_B_pskpqPuo7_1(.din(w_dff_B_uxWcVFyM7_1),.dout(w_dff_B_pskpqPuo7_1),.clk(gclk));
	jdff dff_B_R3I60Yzp2_1(.din(w_dff_B_pskpqPuo7_1),.dout(w_dff_B_R3I60Yzp2_1),.clk(gclk));
	jdff dff_B_5fIXPGLI4_1(.din(w_dff_B_R3I60Yzp2_1),.dout(w_dff_B_5fIXPGLI4_1),.clk(gclk));
	jdff dff_B_S6RAvCjq6_1(.din(w_dff_B_5fIXPGLI4_1),.dout(w_dff_B_S6RAvCjq6_1),.clk(gclk));
	jdff dff_B_DmHFh1vJ1_0(.din(n607),.dout(w_dff_B_DmHFh1vJ1_0),.clk(gclk));
	jdff dff_B_VqROpL253_0(.din(w_dff_B_DmHFh1vJ1_0),.dout(w_dff_B_VqROpL253_0),.clk(gclk));
	jdff dff_B_jIHgcl5h1_0(.din(w_dff_B_VqROpL253_0),.dout(w_dff_B_jIHgcl5h1_0),.clk(gclk));
	jdff dff_B_Sgdhq7o45_0(.din(w_dff_B_jIHgcl5h1_0),.dout(w_dff_B_Sgdhq7o45_0),.clk(gclk));
	jdff dff_B_ilIt7LCa6_0(.din(w_dff_B_Sgdhq7o45_0),.dout(w_dff_B_ilIt7LCa6_0),.clk(gclk));
	jdff dff_B_R0DJgRiQ3_0(.din(w_dff_B_ilIt7LCa6_0),.dout(w_dff_B_R0DJgRiQ3_0),.clk(gclk));
	jdff dff_B_5R8mmLHp8_0(.din(w_dff_B_R0DJgRiQ3_0),.dout(w_dff_B_5R8mmLHp8_0),.clk(gclk));
	jdff dff_B_CguuiksR8_0(.din(w_dff_B_5R8mmLHp8_0),.dout(w_dff_B_CguuiksR8_0),.clk(gclk));
	jdff dff_B_FGXbcDCf4_0(.din(w_dff_B_CguuiksR8_0),.dout(w_dff_B_FGXbcDCf4_0),.clk(gclk));
	jdff dff_B_OqgE3CEy2_0(.din(w_dff_B_FGXbcDCf4_0),.dout(w_dff_B_OqgE3CEy2_0),.clk(gclk));
	jdff dff_B_ns4710rp3_0(.din(w_dff_B_OqgE3CEy2_0),.dout(w_dff_B_ns4710rp3_0),.clk(gclk));
	jdff dff_B_dyeMjlIy7_0(.din(w_dff_B_ns4710rp3_0),.dout(w_dff_B_dyeMjlIy7_0),.clk(gclk));
	jdff dff_B_CFUDoG6Z3_0(.din(w_dff_B_dyeMjlIy7_0),.dout(w_dff_B_CFUDoG6Z3_0),.clk(gclk));
	jdff dff_B_B0sOZkZM6_0(.din(w_dff_B_CFUDoG6Z3_0),.dout(w_dff_B_B0sOZkZM6_0),.clk(gclk));
	jdff dff_B_5gcYsIoH5_0(.din(w_dff_B_B0sOZkZM6_0),.dout(w_dff_B_5gcYsIoH5_0),.clk(gclk));
	jdff dff_B_xiOR2scU6_0(.din(w_dff_B_5gcYsIoH5_0),.dout(w_dff_B_xiOR2scU6_0),.clk(gclk));
	jdff dff_B_BzsR9TK23_0(.din(w_dff_B_xiOR2scU6_0),.dout(w_dff_B_BzsR9TK23_0),.clk(gclk));
	jdff dff_B_bhrvY4bm6_0(.din(w_dff_B_BzsR9TK23_0),.dout(w_dff_B_bhrvY4bm6_0),.clk(gclk));
	jdff dff_B_REKnead37_0(.din(w_dff_B_bhrvY4bm6_0),.dout(w_dff_B_REKnead37_0),.clk(gclk));
	jdff dff_B_1mNAH0Ly8_0(.din(w_dff_B_REKnead37_0),.dout(w_dff_B_1mNAH0Ly8_0),.clk(gclk));
	jdff dff_B_Auq973zI4_0(.din(w_dff_B_1mNAH0Ly8_0),.dout(w_dff_B_Auq973zI4_0),.clk(gclk));
	jdff dff_B_h3Z9Bh2Q6_0(.din(w_dff_B_Auq973zI4_0),.dout(w_dff_B_h3Z9Bh2Q6_0),.clk(gclk));
	jdff dff_B_ilqOOL8z3_0(.din(w_dff_B_h3Z9Bh2Q6_0),.dout(w_dff_B_ilqOOL8z3_0),.clk(gclk));
	jdff dff_B_J1VZ0xkc1_0(.din(w_dff_B_ilqOOL8z3_0),.dout(w_dff_B_J1VZ0xkc1_0),.clk(gclk));
	jdff dff_B_9DyUJqlf7_0(.din(w_dff_B_J1VZ0xkc1_0),.dout(w_dff_B_9DyUJqlf7_0),.clk(gclk));
	jdff dff_B_Otk4fYEB1_0(.din(w_dff_B_9DyUJqlf7_0),.dout(w_dff_B_Otk4fYEB1_0),.clk(gclk));
	jdff dff_B_dr9GPM9O7_0(.din(w_dff_B_Otk4fYEB1_0),.dout(w_dff_B_dr9GPM9O7_0),.clk(gclk));
	jdff dff_B_gskPMh415_0(.din(w_dff_B_dr9GPM9O7_0),.dout(w_dff_B_gskPMh415_0),.clk(gclk));
	jdff dff_B_BzhcQmsX5_0(.din(w_dff_B_gskPMh415_0),.dout(w_dff_B_BzhcQmsX5_0),.clk(gclk));
	jdff dff_B_tT4ya5nE6_0(.din(w_dff_B_BzhcQmsX5_0),.dout(w_dff_B_tT4ya5nE6_0),.clk(gclk));
	jdff dff_B_5Vz0mAoU0_0(.din(w_dff_B_tT4ya5nE6_0),.dout(w_dff_B_5Vz0mAoU0_0),.clk(gclk));
	jdff dff_B_BGDhAFpM9_0(.din(w_dff_B_5Vz0mAoU0_0),.dout(w_dff_B_BGDhAFpM9_0),.clk(gclk));
	jdff dff_B_YfzPuViz1_0(.din(w_dff_B_BGDhAFpM9_0),.dout(w_dff_B_YfzPuViz1_0),.clk(gclk));
	jdff dff_B_ZEuUTuhN9_0(.din(w_dff_B_YfzPuViz1_0),.dout(w_dff_B_ZEuUTuhN9_0),.clk(gclk));
	jdff dff_B_xR5NWHE36_0(.din(w_dff_B_ZEuUTuhN9_0),.dout(w_dff_B_xR5NWHE36_0),.clk(gclk));
	jdff dff_B_LviJle7c6_0(.din(w_dff_B_xR5NWHE36_0),.dout(w_dff_B_LviJle7c6_0),.clk(gclk));
	jdff dff_B_vt7Bt9w49_0(.din(w_dff_B_LviJle7c6_0),.dout(w_dff_B_vt7Bt9w49_0),.clk(gclk));
	jdff dff_B_h5xdW6Ka7_1(.din(n600),.dout(w_dff_B_h5xdW6Ka7_1),.clk(gclk));
	jdff dff_B_sMzxXgdl5_1(.din(w_dff_B_h5xdW6Ka7_1),.dout(w_dff_B_sMzxXgdl5_1),.clk(gclk));
	jdff dff_B_icuzylNk4_1(.din(w_dff_B_sMzxXgdl5_1),.dout(w_dff_B_icuzylNk4_1),.clk(gclk));
	jdff dff_B_52MpWRoQ2_1(.din(w_dff_B_icuzylNk4_1),.dout(w_dff_B_52MpWRoQ2_1),.clk(gclk));
	jdff dff_B_tt2ib7Qh9_1(.din(w_dff_B_52MpWRoQ2_1),.dout(w_dff_B_tt2ib7Qh9_1),.clk(gclk));
	jdff dff_B_UPDmu91F1_1(.din(w_dff_B_tt2ib7Qh9_1),.dout(w_dff_B_UPDmu91F1_1),.clk(gclk));
	jdff dff_B_HcO25vxE5_1(.din(w_dff_B_UPDmu91F1_1),.dout(w_dff_B_HcO25vxE5_1),.clk(gclk));
	jdff dff_B_jpD1P5a48_1(.din(w_dff_B_HcO25vxE5_1),.dout(w_dff_B_jpD1P5a48_1),.clk(gclk));
	jdff dff_B_qfrnzzyn2_1(.din(w_dff_B_jpD1P5a48_1),.dout(w_dff_B_qfrnzzyn2_1),.clk(gclk));
	jdff dff_B_MxZOwriT5_1(.din(w_dff_B_qfrnzzyn2_1),.dout(w_dff_B_MxZOwriT5_1),.clk(gclk));
	jdff dff_B_Hu6DelX76_1(.din(w_dff_B_MxZOwriT5_1),.dout(w_dff_B_Hu6DelX76_1),.clk(gclk));
	jdff dff_B_hQHzplWL8_1(.din(w_dff_B_Hu6DelX76_1),.dout(w_dff_B_hQHzplWL8_1),.clk(gclk));
	jdff dff_B_D4IoxlfC7_1(.din(w_dff_B_hQHzplWL8_1),.dout(w_dff_B_D4IoxlfC7_1),.clk(gclk));
	jdff dff_B_gFuvVzQ31_1(.din(w_dff_B_D4IoxlfC7_1),.dout(w_dff_B_gFuvVzQ31_1),.clk(gclk));
	jdff dff_B_7X2EEtLC2_1(.din(w_dff_B_gFuvVzQ31_1),.dout(w_dff_B_7X2EEtLC2_1),.clk(gclk));
	jdff dff_B_0cN8V0ev7_1(.din(w_dff_B_7X2EEtLC2_1),.dout(w_dff_B_0cN8V0ev7_1),.clk(gclk));
	jdff dff_B_kNX0wAeJ9_1(.din(w_dff_B_0cN8V0ev7_1),.dout(w_dff_B_kNX0wAeJ9_1),.clk(gclk));
	jdff dff_B_sWp3WGKN7_1(.din(w_dff_B_kNX0wAeJ9_1),.dout(w_dff_B_sWp3WGKN7_1),.clk(gclk));
	jdff dff_B_kKOGdNK46_1(.din(w_dff_B_sWp3WGKN7_1),.dout(w_dff_B_kKOGdNK46_1),.clk(gclk));
	jdff dff_B_KYBZSZZK0_1(.din(w_dff_B_kKOGdNK46_1),.dout(w_dff_B_KYBZSZZK0_1),.clk(gclk));
	jdff dff_B_VtTivnjq1_1(.din(w_dff_B_KYBZSZZK0_1),.dout(w_dff_B_VtTivnjq1_1),.clk(gclk));
	jdff dff_B_caDg5JJH9_1(.din(w_dff_B_VtTivnjq1_1),.dout(w_dff_B_caDg5JJH9_1),.clk(gclk));
	jdff dff_B_el37d9oH3_1(.din(w_dff_B_caDg5JJH9_1),.dout(w_dff_B_el37d9oH3_1),.clk(gclk));
	jdff dff_B_94qDdOOI4_1(.din(w_dff_B_el37d9oH3_1),.dout(w_dff_B_94qDdOOI4_1),.clk(gclk));
	jdff dff_B_bxI4QB295_1(.din(w_dff_B_94qDdOOI4_1),.dout(w_dff_B_bxI4QB295_1),.clk(gclk));
	jdff dff_B_lMWKw1qL3_1(.din(w_dff_B_bxI4QB295_1),.dout(w_dff_B_lMWKw1qL3_1),.clk(gclk));
	jdff dff_B_lpHH3xJE8_1(.din(w_dff_B_lMWKw1qL3_1),.dout(w_dff_B_lpHH3xJE8_1),.clk(gclk));
	jdff dff_B_xcIt5GSE5_1(.din(w_dff_B_lpHH3xJE8_1),.dout(w_dff_B_xcIt5GSE5_1),.clk(gclk));
	jdff dff_B_juPcgAlV9_1(.din(w_dff_B_xcIt5GSE5_1),.dout(w_dff_B_juPcgAlV9_1),.clk(gclk));
	jdff dff_B_p3GPETM53_1(.din(w_dff_B_juPcgAlV9_1),.dout(w_dff_B_p3GPETM53_1),.clk(gclk));
	jdff dff_B_z0YRF4gu7_1(.din(w_dff_B_p3GPETM53_1),.dout(w_dff_B_z0YRF4gu7_1),.clk(gclk));
	jdff dff_B_GX55SWVr3_1(.din(w_dff_B_z0YRF4gu7_1),.dout(w_dff_B_GX55SWVr3_1),.clk(gclk));
	jdff dff_B_pIXeCOyP1_1(.din(w_dff_B_GX55SWVr3_1),.dout(w_dff_B_pIXeCOyP1_1),.clk(gclk));
	jdff dff_B_ltcYCDCy1_1(.din(w_dff_B_pIXeCOyP1_1),.dout(w_dff_B_ltcYCDCy1_1),.clk(gclk));
	jdff dff_B_t23r44QK3_1(.din(w_dff_B_ltcYCDCy1_1),.dout(w_dff_B_t23r44QK3_1),.clk(gclk));
	jdff dff_B_ntOAyf159_1(.din(w_dff_B_t23r44QK3_1),.dout(w_dff_B_ntOAyf159_1),.clk(gclk));
	jdff dff_B_BA3uUTcD5_0(.din(n601),.dout(w_dff_B_BA3uUTcD5_0),.clk(gclk));
	jdff dff_B_IY37tbG36_0(.din(w_dff_B_BA3uUTcD5_0),.dout(w_dff_B_IY37tbG36_0),.clk(gclk));
	jdff dff_B_rX8QeA4w1_0(.din(w_dff_B_IY37tbG36_0),.dout(w_dff_B_rX8QeA4w1_0),.clk(gclk));
	jdff dff_B_UunReUbN6_0(.din(w_dff_B_rX8QeA4w1_0),.dout(w_dff_B_UunReUbN6_0),.clk(gclk));
	jdff dff_B_GO1xSD9R9_0(.din(w_dff_B_UunReUbN6_0),.dout(w_dff_B_GO1xSD9R9_0),.clk(gclk));
	jdff dff_B_QdCBvY8M0_0(.din(w_dff_B_GO1xSD9R9_0),.dout(w_dff_B_QdCBvY8M0_0),.clk(gclk));
	jdff dff_B_WYNtXSG78_0(.din(w_dff_B_QdCBvY8M0_0),.dout(w_dff_B_WYNtXSG78_0),.clk(gclk));
	jdff dff_B_vw1qRB0Y3_0(.din(w_dff_B_WYNtXSG78_0),.dout(w_dff_B_vw1qRB0Y3_0),.clk(gclk));
	jdff dff_B_21VJfEaJ9_0(.din(w_dff_B_vw1qRB0Y3_0),.dout(w_dff_B_21VJfEaJ9_0),.clk(gclk));
	jdff dff_B_cMFwrMor9_0(.din(w_dff_B_21VJfEaJ9_0),.dout(w_dff_B_cMFwrMor9_0),.clk(gclk));
	jdff dff_B_HypVbknO8_0(.din(w_dff_B_cMFwrMor9_0),.dout(w_dff_B_HypVbknO8_0),.clk(gclk));
	jdff dff_B_U6v6e7Ma9_0(.din(w_dff_B_HypVbknO8_0),.dout(w_dff_B_U6v6e7Ma9_0),.clk(gclk));
	jdff dff_B_7JABikK63_0(.din(w_dff_B_U6v6e7Ma9_0),.dout(w_dff_B_7JABikK63_0),.clk(gclk));
	jdff dff_B_Wcy97j6v0_0(.din(w_dff_B_7JABikK63_0),.dout(w_dff_B_Wcy97j6v0_0),.clk(gclk));
	jdff dff_B_wAZV1ICG5_0(.din(w_dff_B_Wcy97j6v0_0),.dout(w_dff_B_wAZV1ICG5_0),.clk(gclk));
	jdff dff_B_RnExXpTC8_0(.din(w_dff_B_wAZV1ICG5_0),.dout(w_dff_B_RnExXpTC8_0),.clk(gclk));
	jdff dff_B_M6EWYHAY4_0(.din(w_dff_B_RnExXpTC8_0),.dout(w_dff_B_M6EWYHAY4_0),.clk(gclk));
	jdff dff_B_ztlmdiCI5_0(.din(w_dff_B_M6EWYHAY4_0),.dout(w_dff_B_ztlmdiCI5_0),.clk(gclk));
	jdff dff_B_gOvI0Pqc2_0(.din(w_dff_B_ztlmdiCI5_0),.dout(w_dff_B_gOvI0Pqc2_0),.clk(gclk));
	jdff dff_B_BedvMGyv6_0(.din(w_dff_B_gOvI0Pqc2_0),.dout(w_dff_B_BedvMGyv6_0),.clk(gclk));
	jdff dff_B_12UjqWxY1_0(.din(w_dff_B_BedvMGyv6_0),.dout(w_dff_B_12UjqWxY1_0),.clk(gclk));
	jdff dff_B_Hr36akQr9_0(.din(w_dff_B_12UjqWxY1_0),.dout(w_dff_B_Hr36akQr9_0),.clk(gclk));
	jdff dff_B_9E4UyoDN3_0(.din(w_dff_B_Hr36akQr9_0),.dout(w_dff_B_9E4UyoDN3_0),.clk(gclk));
	jdff dff_B_KU25avqa7_0(.din(w_dff_B_9E4UyoDN3_0),.dout(w_dff_B_KU25avqa7_0),.clk(gclk));
	jdff dff_B_BvqJYc5o9_0(.din(w_dff_B_KU25avqa7_0),.dout(w_dff_B_BvqJYc5o9_0),.clk(gclk));
	jdff dff_B_g3pE7bqQ3_0(.din(w_dff_B_BvqJYc5o9_0),.dout(w_dff_B_g3pE7bqQ3_0),.clk(gclk));
	jdff dff_B_bjj7b4G76_0(.din(w_dff_B_g3pE7bqQ3_0),.dout(w_dff_B_bjj7b4G76_0),.clk(gclk));
	jdff dff_B_ts6zT4X01_0(.din(w_dff_B_bjj7b4G76_0),.dout(w_dff_B_ts6zT4X01_0),.clk(gclk));
	jdff dff_B_1WI8exoW7_0(.din(w_dff_B_ts6zT4X01_0),.dout(w_dff_B_1WI8exoW7_0),.clk(gclk));
	jdff dff_B_dQzew06Y4_0(.din(w_dff_B_1WI8exoW7_0),.dout(w_dff_B_dQzew06Y4_0),.clk(gclk));
	jdff dff_B_s5s1FNvm2_0(.din(w_dff_B_dQzew06Y4_0),.dout(w_dff_B_s5s1FNvm2_0),.clk(gclk));
	jdff dff_B_LTklb7IV9_0(.din(w_dff_B_s5s1FNvm2_0),.dout(w_dff_B_LTklb7IV9_0),.clk(gclk));
	jdff dff_B_3OBW9knB7_0(.din(w_dff_B_LTklb7IV9_0),.dout(w_dff_B_3OBW9knB7_0),.clk(gclk));
	jdff dff_B_ksPxZ7WT3_0(.din(w_dff_B_3OBW9knB7_0),.dout(w_dff_B_ksPxZ7WT3_0),.clk(gclk));
	jdff dff_B_T2Fc7qLA3_0(.din(w_dff_B_ksPxZ7WT3_0),.dout(w_dff_B_T2Fc7qLA3_0),.clk(gclk));
	jdff dff_B_Giv88Gjw1_0(.din(w_dff_B_T2Fc7qLA3_0),.dout(w_dff_B_Giv88Gjw1_0),.clk(gclk));
	jdff dff_B_RFleY3cT7_1(.din(n594),.dout(w_dff_B_RFleY3cT7_1),.clk(gclk));
	jdff dff_B_o0SdHfrv0_1(.din(w_dff_B_RFleY3cT7_1),.dout(w_dff_B_o0SdHfrv0_1),.clk(gclk));
	jdff dff_B_PKCgycnV4_1(.din(w_dff_B_o0SdHfrv0_1),.dout(w_dff_B_PKCgycnV4_1),.clk(gclk));
	jdff dff_B_n7CGMQ451_1(.din(w_dff_B_PKCgycnV4_1),.dout(w_dff_B_n7CGMQ451_1),.clk(gclk));
	jdff dff_B_aaMGmXGc4_1(.din(w_dff_B_n7CGMQ451_1),.dout(w_dff_B_aaMGmXGc4_1),.clk(gclk));
	jdff dff_B_n3t1iiLE1_1(.din(w_dff_B_aaMGmXGc4_1),.dout(w_dff_B_n3t1iiLE1_1),.clk(gclk));
	jdff dff_B_zoIudX5I5_1(.din(w_dff_B_n3t1iiLE1_1),.dout(w_dff_B_zoIudX5I5_1),.clk(gclk));
	jdff dff_B_0uGNVUpk4_1(.din(w_dff_B_zoIudX5I5_1),.dout(w_dff_B_0uGNVUpk4_1),.clk(gclk));
	jdff dff_B_N5OF68FT9_1(.din(w_dff_B_0uGNVUpk4_1),.dout(w_dff_B_N5OF68FT9_1),.clk(gclk));
	jdff dff_B_oxLipQWa5_1(.din(w_dff_B_N5OF68FT9_1),.dout(w_dff_B_oxLipQWa5_1),.clk(gclk));
	jdff dff_B_d3Tt3NNn6_1(.din(w_dff_B_oxLipQWa5_1),.dout(w_dff_B_d3Tt3NNn6_1),.clk(gclk));
	jdff dff_B_gLIVBpqf8_1(.din(w_dff_B_d3Tt3NNn6_1),.dout(w_dff_B_gLIVBpqf8_1),.clk(gclk));
	jdff dff_B_gLSRRrlu8_1(.din(w_dff_B_gLIVBpqf8_1),.dout(w_dff_B_gLSRRrlu8_1),.clk(gclk));
	jdff dff_B_DCCReXPn7_1(.din(w_dff_B_gLSRRrlu8_1),.dout(w_dff_B_DCCReXPn7_1),.clk(gclk));
	jdff dff_B_RhH8y4yo4_1(.din(w_dff_B_DCCReXPn7_1),.dout(w_dff_B_RhH8y4yo4_1),.clk(gclk));
	jdff dff_B_5kKUMZGE4_1(.din(w_dff_B_RhH8y4yo4_1),.dout(w_dff_B_5kKUMZGE4_1),.clk(gclk));
	jdff dff_B_Vy6giZbs8_1(.din(w_dff_B_5kKUMZGE4_1),.dout(w_dff_B_Vy6giZbs8_1),.clk(gclk));
	jdff dff_B_4HeTjNQa2_1(.din(w_dff_B_Vy6giZbs8_1),.dout(w_dff_B_4HeTjNQa2_1),.clk(gclk));
	jdff dff_B_jHqlPfIE7_1(.din(w_dff_B_4HeTjNQa2_1),.dout(w_dff_B_jHqlPfIE7_1),.clk(gclk));
	jdff dff_B_m88H5LkI7_1(.din(w_dff_B_jHqlPfIE7_1),.dout(w_dff_B_m88H5LkI7_1),.clk(gclk));
	jdff dff_B_NxU417Uu9_1(.din(w_dff_B_m88H5LkI7_1),.dout(w_dff_B_NxU417Uu9_1),.clk(gclk));
	jdff dff_B_K7fU8ITe9_1(.din(w_dff_B_NxU417Uu9_1),.dout(w_dff_B_K7fU8ITe9_1),.clk(gclk));
	jdff dff_B_QG2BfaTf6_1(.din(w_dff_B_K7fU8ITe9_1),.dout(w_dff_B_QG2BfaTf6_1),.clk(gclk));
	jdff dff_B_5V6RjaT84_1(.din(w_dff_B_QG2BfaTf6_1),.dout(w_dff_B_5V6RjaT84_1),.clk(gclk));
	jdff dff_B_wI1eJqcb0_1(.din(w_dff_B_5V6RjaT84_1),.dout(w_dff_B_wI1eJqcb0_1),.clk(gclk));
	jdff dff_B_ZPIO6g0O6_1(.din(w_dff_B_wI1eJqcb0_1),.dout(w_dff_B_ZPIO6g0O6_1),.clk(gclk));
	jdff dff_B_6hHLCboa5_1(.din(w_dff_B_ZPIO6g0O6_1),.dout(w_dff_B_6hHLCboa5_1),.clk(gclk));
	jdff dff_B_8UPRRRSB7_1(.din(w_dff_B_6hHLCboa5_1),.dout(w_dff_B_8UPRRRSB7_1),.clk(gclk));
	jdff dff_B_QkHjKDoB8_1(.din(w_dff_B_8UPRRRSB7_1),.dout(w_dff_B_QkHjKDoB8_1),.clk(gclk));
	jdff dff_B_4kZcQGWj4_1(.din(w_dff_B_QkHjKDoB8_1),.dout(w_dff_B_4kZcQGWj4_1),.clk(gclk));
	jdff dff_B_s8fbOKAE3_1(.din(w_dff_B_4kZcQGWj4_1),.dout(w_dff_B_s8fbOKAE3_1),.clk(gclk));
	jdff dff_B_TtdLCU858_1(.din(w_dff_B_s8fbOKAE3_1),.dout(w_dff_B_TtdLCU858_1),.clk(gclk));
	jdff dff_B_VY1D2qEV5_1(.din(w_dff_B_TtdLCU858_1),.dout(w_dff_B_VY1D2qEV5_1),.clk(gclk));
	jdff dff_B_9XkkEIKa9_1(.din(w_dff_B_VY1D2qEV5_1),.dout(w_dff_B_9XkkEIKa9_1),.clk(gclk));
	jdff dff_B_PbcuSyj41_1(.din(w_dff_B_9XkkEIKa9_1),.dout(w_dff_B_PbcuSyj41_1),.clk(gclk));
	jdff dff_B_Rqvx2lkt1_0(.din(n595),.dout(w_dff_B_Rqvx2lkt1_0),.clk(gclk));
	jdff dff_B_MUXDV8y82_0(.din(w_dff_B_Rqvx2lkt1_0),.dout(w_dff_B_MUXDV8y82_0),.clk(gclk));
	jdff dff_B_Hib5v7zF8_0(.din(w_dff_B_MUXDV8y82_0),.dout(w_dff_B_Hib5v7zF8_0),.clk(gclk));
	jdff dff_B_36deffBk1_0(.din(w_dff_B_Hib5v7zF8_0),.dout(w_dff_B_36deffBk1_0),.clk(gclk));
	jdff dff_B_Z4trfWgg6_0(.din(w_dff_B_36deffBk1_0),.dout(w_dff_B_Z4trfWgg6_0),.clk(gclk));
	jdff dff_B_w1i2sHnu1_0(.din(w_dff_B_Z4trfWgg6_0),.dout(w_dff_B_w1i2sHnu1_0),.clk(gclk));
	jdff dff_B_xJyfTY1R9_0(.din(w_dff_B_w1i2sHnu1_0),.dout(w_dff_B_xJyfTY1R9_0),.clk(gclk));
	jdff dff_B_nkW5Mc1L2_0(.din(w_dff_B_xJyfTY1R9_0),.dout(w_dff_B_nkW5Mc1L2_0),.clk(gclk));
	jdff dff_B_hr540QWz5_0(.din(w_dff_B_nkW5Mc1L2_0),.dout(w_dff_B_hr540QWz5_0),.clk(gclk));
	jdff dff_B_s5CVi2OT9_0(.din(w_dff_B_hr540QWz5_0),.dout(w_dff_B_s5CVi2OT9_0),.clk(gclk));
	jdff dff_B_Zrlwuc2h1_0(.din(w_dff_B_s5CVi2OT9_0),.dout(w_dff_B_Zrlwuc2h1_0),.clk(gclk));
	jdff dff_B_lk1kZ6Oj4_0(.din(w_dff_B_Zrlwuc2h1_0),.dout(w_dff_B_lk1kZ6Oj4_0),.clk(gclk));
	jdff dff_B_IoEansJ12_0(.din(w_dff_B_lk1kZ6Oj4_0),.dout(w_dff_B_IoEansJ12_0),.clk(gclk));
	jdff dff_B_vKcd36FX3_0(.din(w_dff_B_IoEansJ12_0),.dout(w_dff_B_vKcd36FX3_0),.clk(gclk));
	jdff dff_B_yPl8uL8o9_0(.din(w_dff_B_vKcd36FX3_0),.dout(w_dff_B_yPl8uL8o9_0),.clk(gclk));
	jdff dff_B_dxNMwbHM4_0(.din(w_dff_B_yPl8uL8o9_0),.dout(w_dff_B_dxNMwbHM4_0),.clk(gclk));
	jdff dff_B_1Bp3UrTf9_0(.din(w_dff_B_dxNMwbHM4_0),.dout(w_dff_B_1Bp3UrTf9_0),.clk(gclk));
	jdff dff_B_bdrTM9D63_0(.din(w_dff_B_1Bp3UrTf9_0),.dout(w_dff_B_bdrTM9D63_0),.clk(gclk));
	jdff dff_B_S2GLdNs63_0(.din(w_dff_B_bdrTM9D63_0),.dout(w_dff_B_S2GLdNs63_0),.clk(gclk));
	jdff dff_B_UogI0Y4z9_0(.din(w_dff_B_S2GLdNs63_0),.dout(w_dff_B_UogI0Y4z9_0),.clk(gclk));
	jdff dff_B_ZGwpUHiZ3_0(.din(w_dff_B_UogI0Y4z9_0),.dout(w_dff_B_ZGwpUHiZ3_0),.clk(gclk));
	jdff dff_B_AW74jYXA5_0(.din(w_dff_B_ZGwpUHiZ3_0),.dout(w_dff_B_AW74jYXA5_0),.clk(gclk));
	jdff dff_B_G1gWiONj5_0(.din(w_dff_B_AW74jYXA5_0),.dout(w_dff_B_G1gWiONj5_0),.clk(gclk));
	jdff dff_B_otHs145F4_0(.din(w_dff_B_G1gWiONj5_0),.dout(w_dff_B_otHs145F4_0),.clk(gclk));
	jdff dff_B_J6HEMNNZ1_0(.din(w_dff_B_otHs145F4_0),.dout(w_dff_B_J6HEMNNZ1_0),.clk(gclk));
	jdff dff_B_nzuQA4Fm8_0(.din(w_dff_B_J6HEMNNZ1_0),.dout(w_dff_B_nzuQA4Fm8_0),.clk(gclk));
	jdff dff_B_qK5Sdcws0_0(.din(w_dff_B_nzuQA4Fm8_0),.dout(w_dff_B_qK5Sdcws0_0),.clk(gclk));
	jdff dff_B_3OTtlZsH6_0(.din(w_dff_B_qK5Sdcws0_0),.dout(w_dff_B_3OTtlZsH6_0),.clk(gclk));
	jdff dff_B_U8xbl7qB7_0(.din(w_dff_B_3OTtlZsH6_0),.dout(w_dff_B_U8xbl7qB7_0),.clk(gclk));
	jdff dff_B_rwAlfQEC1_0(.din(w_dff_B_U8xbl7qB7_0),.dout(w_dff_B_rwAlfQEC1_0),.clk(gclk));
	jdff dff_B_WD8zd9KI8_0(.din(w_dff_B_rwAlfQEC1_0),.dout(w_dff_B_WD8zd9KI8_0),.clk(gclk));
	jdff dff_B_tgrF5Hzc9_0(.din(w_dff_B_WD8zd9KI8_0),.dout(w_dff_B_tgrF5Hzc9_0),.clk(gclk));
	jdff dff_B_NBNeCR8Y4_0(.din(w_dff_B_tgrF5Hzc9_0),.dout(w_dff_B_NBNeCR8Y4_0),.clk(gclk));
	jdff dff_B_UgeCLmEn2_0(.din(w_dff_B_NBNeCR8Y4_0),.dout(w_dff_B_UgeCLmEn2_0),.clk(gclk));
	jdff dff_B_N2n8UqAM7_0(.din(w_dff_B_UgeCLmEn2_0),.dout(w_dff_B_N2n8UqAM7_0),.clk(gclk));
	jdff dff_B_02b2xEfn2_1(.din(n588),.dout(w_dff_B_02b2xEfn2_1),.clk(gclk));
	jdff dff_B_gkzTkmCx1_1(.din(w_dff_B_02b2xEfn2_1),.dout(w_dff_B_gkzTkmCx1_1),.clk(gclk));
	jdff dff_B_jRWgKmn68_1(.din(w_dff_B_gkzTkmCx1_1),.dout(w_dff_B_jRWgKmn68_1),.clk(gclk));
	jdff dff_B_plYVua4g6_1(.din(w_dff_B_jRWgKmn68_1),.dout(w_dff_B_plYVua4g6_1),.clk(gclk));
	jdff dff_B_tjH0DXuC6_1(.din(w_dff_B_plYVua4g6_1),.dout(w_dff_B_tjH0DXuC6_1),.clk(gclk));
	jdff dff_B_Ipjlbscu2_1(.din(w_dff_B_tjH0DXuC6_1),.dout(w_dff_B_Ipjlbscu2_1),.clk(gclk));
	jdff dff_B_50Lqqz3j7_1(.din(w_dff_B_Ipjlbscu2_1),.dout(w_dff_B_50Lqqz3j7_1),.clk(gclk));
	jdff dff_B_oeLEYTe21_1(.din(w_dff_B_50Lqqz3j7_1),.dout(w_dff_B_oeLEYTe21_1),.clk(gclk));
	jdff dff_B_oomihasE2_1(.din(w_dff_B_oeLEYTe21_1),.dout(w_dff_B_oomihasE2_1),.clk(gclk));
	jdff dff_B_Una2FvI36_1(.din(w_dff_B_oomihasE2_1),.dout(w_dff_B_Una2FvI36_1),.clk(gclk));
	jdff dff_B_xASc30645_1(.din(w_dff_B_Una2FvI36_1),.dout(w_dff_B_xASc30645_1),.clk(gclk));
	jdff dff_B_ZSFXmSrz0_1(.din(w_dff_B_xASc30645_1),.dout(w_dff_B_ZSFXmSrz0_1),.clk(gclk));
	jdff dff_B_Klg170KV7_1(.din(w_dff_B_ZSFXmSrz0_1),.dout(w_dff_B_Klg170KV7_1),.clk(gclk));
	jdff dff_B_926dC0rJ0_1(.din(w_dff_B_Klg170KV7_1),.dout(w_dff_B_926dC0rJ0_1),.clk(gclk));
	jdff dff_B_FjgoKXaQ8_1(.din(w_dff_B_926dC0rJ0_1),.dout(w_dff_B_FjgoKXaQ8_1),.clk(gclk));
	jdff dff_B_FIntbdhJ6_1(.din(w_dff_B_FjgoKXaQ8_1),.dout(w_dff_B_FIntbdhJ6_1),.clk(gclk));
	jdff dff_B_RjS4d5lB5_1(.din(w_dff_B_FIntbdhJ6_1),.dout(w_dff_B_RjS4d5lB5_1),.clk(gclk));
	jdff dff_B_1Ct1ObmX7_1(.din(w_dff_B_RjS4d5lB5_1),.dout(w_dff_B_1Ct1ObmX7_1),.clk(gclk));
	jdff dff_B_RnbTfalx4_1(.din(w_dff_B_1Ct1ObmX7_1),.dout(w_dff_B_RnbTfalx4_1),.clk(gclk));
	jdff dff_B_BbDgaJkA2_1(.din(w_dff_B_RnbTfalx4_1),.dout(w_dff_B_BbDgaJkA2_1),.clk(gclk));
	jdff dff_B_A4O1rxU15_1(.din(w_dff_B_BbDgaJkA2_1),.dout(w_dff_B_A4O1rxU15_1),.clk(gclk));
	jdff dff_B_yYNvWGU08_1(.din(w_dff_B_A4O1rxU15_1),.dout(w_dff_B_yYNvWGU08_1),.clk(gclk));
	jdff dff_B_KuIDJd9f3_1(.din(w_dff_B_yYNvWGU08_1),.dout(w_dff_B_KuIDJd9f3_1),.clk(gclk));
	jdff dff_B_TdjAzBHD0_1(.din(w_dff_B_KuIDJd9f3_1),.dout(w_dff_B_TdjAzBHD0_1),.clk(gclk));
	jdff dff_B_CoN9U1CR8_1(.din(w_dff_B_TdjAzBHD0_1),.dout(w_dff_B_CoN9U1CR8_1),.clk(gclk));
	jdff dff_B_R2j7WGDG4_1(.din(w_dff_B_CoN9U1CR8_1),.dout(w_dff_B_R2j7WGDG4_1),.clk(gclk));
	jdff dff_B_A74IMyT57_1(.din(w_dff_B_R2j7WGDG4_1),.dout(w_dff_B_A74IMyT57_1),.clk(gclk));
	jdff dff_B_Ky1Ma0gz9_1(.din(w_dff_B_A74IMyT57_1),.dout(w_dff_B_Ky1Ma0gz9_1),.clk(gclk));
	jdff dff_B_IUzz9bHI1_1(.din(w_dff_B_Ky1Ma0gz9_1),.dout(w_dff_B_IUzz9bHI1_1),.clk(gclk));
	jdff dff_B_LLMWUEpr8_1(.din(w_dff_B_IUzz9bHI1_1),.dout(w_dff_B_LLMWUEpr8_1),.clk(gclk));
	jdff dff_B_bWlS1lQp9_1(.din(w_dff_B_LLMWUEpr8_1),.dout(w_dff_B_bWlS1lQp9_1),.clk(gclk));
	jdff dff_B_faX2aisv2_1(.din(w_dff_B_bWlS1lQp9_1),.dout(w_dff_B_faX2aisv2_1),.clk(gclk));
	jdff dff_B_RvlOhSxn9_1(.din(w_dff_B_faX2aisv2_1),.dout(w_dff_B_RvlOhSxn9_1),.clk(gclk));
	jdff dff_B_xBRXkssz2_1(.din(w_dff_B_RvlOhSxn9_1),.dout(w_dff_B_xBRXkssz2_1),.clk(gclk));
	jdff dff_B_jPjE4w566_0(.din(n589),.dout(w_dff_B_jPjE4w566_0),.clk(gclk));
	jdff dff_B_Ri33JLN58_0(.din(w_dff_B_jPjE4w566_0),.dout(w_dff_B_Ri33JLN58_0),.clk(gclk));
	jdff dff_B_qzVPKuyH0_0(.din(w_dff_B_Ri33JLN58_0),.dout(w_dff_B_qzVPKuyH0_0),.clk(gclk));
	jdff dff_B_Z9Wml6E79_0(.din(w_dff_B_qzVPKuyH0_0),.dout(w_dff_B_Z9Wml6E79_0),.clk(gclk));
	jdff dff_B_DpwaP6ej4_0(.din(w_dff_B_Z9Wml6E79_0),.dout(w_dff_B_DpwaP6ej4_0),.clk(gclk));
	jdff dff_B_FO1BGuR42_0(.din(w_dff_B_DpwaP6ej4_0),.dout(w_dff_B_FO1BGuR42_0),.clk(gclk));
	jdff dff_B_CGZ7jiuy1_0(.din(w_dff_B_FO1BGuR42_0),.dout(w_dff_B_CGZ7jiuy1_0),.clk(gclk));
	jdff dff_B_Zzm804cc2_0(.din(w_dff_B_CGZ7jiuy1_0),.dout(w_dff_B_Zzm804cc2_0),.clk(gclk));
	jdff dff_B_PQ69IjpM0_0(.din(w_dff_B_Zzm804cc2_0),.dout(w_dff_B_PQ69IjpM0_0),.clk(gclk));
	jdff dff_B_DNhqEuWv9_0(.din(w_dff_B_PQ69IjpM0_0),.dout(w_dff_B_DNhqEuWv9_0),.clk(gclk));
	jdff dff_B_ZLY8E1Ar3_0(.din(w_dff_B_DNhqEuWv9_0),.dout(w_dff_B_ZLY8E1Ar3_0),.clk(gclk));
	jdff dff_B_AbBPNhSW3_0(.din(w_dff_B_ZLY8E1Ar3_0),.dout(w_dff_B_AbBPNhSW3_0),.clk(gclk));
	jdff dff_B_g4mkXwWN6_0(.din(w_dff_B_AbBPNhSW3_0),.dout(w_dff_B_g4mkXwWN6_0),.clk(gclk));
	jdff dff_B_aAQAtjIZ1_0(.din(w_dff_B_g4mkXwWN6_0),.dout(w_dff_B_aAQAtjIZ1_0),.clk(gclk));
	jdff dff_B_lAOr0Neg3_0(.din(w_dff_B_aAQAtjIZ1_0),.dout(w_dff_B_lAOr0Neg3_0),.clk(gclk));
	jdff dff_B_PxYGi3lK2_0(.din(w_dff_B_lAOr0Neg3_0),.dout(w_dff_B_PxYGi3lK2_0),.clk(gclk));
	jdff dff_B_m9edO10P9_0(.din(w_dff_B_PxYGi3lK2_0),.dout(w_dff_B_m9edO10P9_0),.clk(gclk));
	jdff dff_B_8m53RdS99_0(.din(w_dff_B_m9edO10P9_0),.dout(w_dff_B_8m53RdS99_0),.clk(gclk));
	jdff dff_B_OqzuyDLw2_0(.din(w_dff_B_8m53RdS99_0),.dout(w_dff_B_OqzuyDLw2_0),.clk(gclk));
	jdff dff_B_87Cmlgxq5_0(.din(w_dff_B_OqzuyDLw2_0),.dout(w_dff_B_87Cmlgxq5_0),.clk(gclk));
	jdff dff_B_KwyDwHQw0_0(.din(w_dff_B_87Cmlgxq5_0),.dout(w_dff_B_KwyDwHQw0_0),.clk(gclk));
	jdff dff_B_Advn2Nhl0_0(.din(w_dff_B_KwyDwHQw0_0),.dout(w_dff_B_Advn2Nhl0_0),.clk(gclk));
	jdff dff_B_r1lyi1PS9_0(.din(w_dff_B_Advn2Nhl0_0),.dout(w_dff_B_r1lyi1PS9_0),.clk(gclk));
	jdff dff_B_sTmFQkDr7_0(.din(w_dff_B_r1lyi1PS9_0),.dout(w_dff_B_sTmFQkDr7_0),.clk(gclk));
	jdff dff_B_r2VTro4A7_0(.din(w_dff_B_sTmFQkDr7_0),.dout(w_dff_B_r2VTro4A7_0),.clk(gclk));
	jdff dff_B_YavBotb38_0(.din(w_dff_B_r2VTro4A7_0),.dout(w_dff_B_YavBotb38_0),.clk(gclk));
	jdff dff_B_J4vcTPkf5_0(.din(w_dff_B_YavBotb38_0),.dout(w_dff_B_J4vcTPkf5_0),.clk(gclk));
	jdff dff_B_CiejrLnL6_0(.din(w_dff_B_J4vcTPkf5_0),.dout(w_dff_B_CiejrLnL6_0),.clk(gclk));
	jdff dff_B_s0ABvs464_0(.din(w_dff_B_CiejrLnL6_0),.dout(w_dff_B_s0ABvs464_0),.clk(gclk));
	jdff dff_B_IXBbbxc29_0(.din(w_dff_B_s0ABvs464_0),.dout(w_dff_B_IXBbbxc29_0),.clk(gclk));
	jdff dff_B_aHx5w51h0_0(.din(w_dff_B_IXBbbxc29_0),.dout(w_dff_B_aHx5w51h0_0),.clk(gclk));
	jdff dff_B_mEZxTeOo9_0(.din(w_dff_B_aHx5w51h0_0),.dout(w_dff_B_mEZxTeOo9_0),.clk(gclk));
	jdff dff_B_iI1rlTwq7_0(.din(w_dff_B_mEZxTeOo9_0),.dout(w_dff_B_iI1rlTwq7_0),.clk(gclk));
	jdff dff_B_NuWicBqk2_0(.din(w_dff_B_iI1rlTwq7_0),.dout(w_dff_B_NuWicBqk2_0),.clk(gclk));
	jdff dff_B_02Ap5I3I2_1(.din(n582),.dout(w_dff_B_02Ap5I3I2_1),.clk(gclk));
	jdff dff_B_KMkF11mo1_1(.din(w_dff_B_02Ap5I3I2_1),.dout(w_dff_B_KMkF11mo1_1),.clk(gclk));
	jdff dff_B_wFI2wHrj4_1(.din(w_dff_B_KMkF11mo1_1),.dout(w_dff_B_wFI2wHrj4_1),.clk(gclk));
	jdff dff_B_l9DDrO862_1(.din(w_dff_B_wFI2wHrj4_1),.dout(w_dff_B_l9DDrO862_1),.clk(gclk));
	jdff dff_B_80uY3sSQ4_1(.din(w_dff_B_l9DDrO862_1),.dout(w_dff_B_80uY3sSQ4_1),.clk(gclk));
	jdff dff_B_zWWTpkUM0_1(.din(w_dff_B_80uY3sSQ4_1),.dout(w_dff_B_zWWTpkUM0_1),.clk(gclk));
	jdff dff_B_4hoZaLfJ4_1(.din(w_dff_B_zWWTpkUM0_1),.dout(w_dff_B_4hoZaLfJ4_1),.clk(gclk));
	jdff dff_B_64h7T9QD7_1(.din(w_dff_B_4hoZaLfJ4_1),.dout(w_dff_B_64h7T9QD7_1),.clk(gclk));
	jdff dff_B_6ZBuhXOA6_1(.din(w_dff_B_64h7T9QD7_1),.dout(w_dff_B_6ZBuhXOA6_1),.clk(gclk));
	jdff dff_B_M2iBSq8J2_1(.din(w_dff_B_6ZBuhXOA6_1),.dout(w_dff_B_M2iBSq8J2_1),.clk(gclk));
	jdff dff_B_Eujl7wjc8_1(.din(w_dff_B_M2iBSq8J2_1),.dout(w_dff_B_Eujl7wjc8_1),.clk(gclk));
	jdff dff_B_i60bOPkj2_1(.din(w_dff_B_Eujl7wjc8_1),.dout(w_dff_B_i60bOPkj2_1),.clk(gclk));
	jdff dff_B_F6HgQXgX6_1(.din(w_dff_B_i60bOPkj2_1),.dout(w_dff_B_F6HgQXgX6_1),.clk(gclk));
	jdff dff_B_wFnbaeXT9_1(.din(w_dff_B_F6HgQXgX6_1),.dout(w_dff_B_wFnbaeXT9_1),.clk(gclk));
	jdff dff_B_QfdSnFPW9_1(.din(w_dff_B_wFnbaeXT9_1),.dout(w_dff_B_QfdSnFPW9_1),.clk(gclk));
	jdff dff_B_UdEM3CIt5_1(.din(w_dff_B_QfdSnFPW9_1),.dout(w_dff_B_UdEM3CIt5_1),.clk(gclk));
	jdff dff_B_N8lCJAP71_1(.din(w_dff_B_UdEM3CIt5_1),.dout(w_dff_B_N8lCJAP71_1),.clk(gclk));
	jdff dff_B_9KpUejbz4_1(.din(w_dff_B_N8lCJAP71_1),.dout(w_dff_B_9KpUejbz4_1),.clk(gclk));
	jdff dff_B_u6uv26L64_1(.din(w_dff_B_9KpUejbz4_1),.dout(w_dff_B_u6uv26L64_1),.clk(gclk));
	jdff dff_B_gwihwOcj1_1(.din(w_dff_B_u6uv26L64_1),.dout(w_dff_B_gwihwOcj1_1),.clk(gclk));
	jdff dff_B_12ndL5kl2_1(.din(w_dff_B_gwihwOcj1_1),.dout(w_dff_B_12ndL5kl2_1),.clk(gclk));
	jdff dff_B_w7LtAWwv4_1(.din(w_dff_B_12ndL5kl2_1),.dout(w_dff_B_w7LtAWwv4_1),.clk(gclk));
	jdff dff_B_8DU8tLtq3_1(.din(w_dff_B_w7LtAWwv4_1),.dout(w_dff_B_8DU8tLtq3_1),.clk(gclk));
	jdff dff_B_ZQQIIxgW6_1(.din(w_dff_B_8DU8tLtq3_1),.dout(w_dff_B_ZQQIIxgW6_1),.clk(gclk));
	jdff dff_B_rHDfCPm65_1(.din(w_dff_B_ZQQIIxgW6_1),.dout(w_dff_B_rHDfCPm65_1),.clk(gclk));
	jdff dff_B_BLOZd5o33_1(.din(w_dff_B_rHDfCPm65_1),.dout(w_dff_B_BLOZd5o33_1),.clk(gclk));
	jdff dff_B_ybr6fgZm2_1(.din(w_dff_B_BLOZd5o33_1),.dout(w_dff_B_ybr6fgZm2_1),.clk(gclk));
	jdff dff_B_JfQCiZAS3_1(.din(w_dff_B_ybr6fgZm2_1),.dout(w_dff_B_JfQCiZAS3_1),.clk(gclk));
	jdff dff_B_vD1Xj51c1_1(.din(w_dff_B_JfQCiZAS3_1),.dout(w_dff_B_vD1Xj51c1_1),.clk(gclk));
	jdff dff_B_zqSHb1R55_1(.din(w_dff_B_vD1Xj51c1_1),.dout(w_dff_B_zqSHb1R55_1),.clk(gclk));
	jdff dff_B_zlZ0WpMP4_1(.din(w_dff_B_zqSHb1R55_1),.dout(w_dff_B_zlZ0WpMP4_1),.clk(gclk));
	jdff dff_B_anBghBRu9_1(.din(w_dff_B_zlZ0WpMP4_1),.dout(w_dff_B_anBghBRu9_1),.clk(gclk));
	jdff dff_B_D2kiPHXL3_1(.din(w_dff_B_anBghBRu9_1),.dout(w_dff_B_D2kiPHXL3_1),.clk(gclk));
	jdff dff_B_7RJiBTay1_0(.din(n583),.dout(w_dff_B_7RJiBTay1_0),.clk(gclk));
	jdff dff_B_VpafdGyq6_0(.din(w_dff_B_7RJiBTay1_0),.dout(w_dff_B_VpafdGyq6_0),.clk(gclk));
	jdff dff_B_LOxNFQMu9_0(.din(w_dff_B_VpafdGyq6_0),.dout(w_dff_B_LOxNFQMu9_0),.clk(gclk));
	jdff dff_B_xdQIF0Ce8_0(.din(w_dff_B_LOxNFQMu9_0),.dout(w_dff_B_xdQIF0Ce8_0),.clk(gclk));
	jdff dff_B_JhyBeqdV9_0(.din(w_dff_B_xdQIF0Ce8_0),.dout(w_dff_B_JhyBeqdV9_0),.clk(gclk));
	jdff dff_B_ypxhoOHo6_0(.din(w_dff_B_JhyBeqdV9_0),.dout(w_dff_B_ypxhoOHo6_0),.clk(gclk));
	jdff dff_B_RtYdGEuc6_0(.din(w_dff_B_ypxhoOHo6_0),.dout(w_dff_B_RtYdGEuc6_0),.clk(gclk));
	jdff dff_B_kCbcZnUt0_0(.din(w_dff_B_RtYdGEuc6_0),.dout(w_dff_B_kCbcZnUt0_0),.clk(gclk));
	jdff dff_B_JmmLgQQy9_0(.din(w_dff_B_kCbcZnUt0_0),.dout(w_dff_B_JmmLgQQy9_0),.clk(gclk));
	jdff dff_B_bud2Cav66_0(.din(w_dff_B_JmmLgQQy9_0),.dout(w_dff_B_bud2Cav66_0),.clk(gclk));
	jdff dff_B_Qacz87Np6_0(.din(w_dff_B_bud2Cav66_0),.dout(w_dff_B_Qacz87Np6_0),.clk(gclk));
	jdff dff_B_roIrZ3r95_0(.din(w_dff_B_Qacz87Np6_0),.dout(w_dff_B_roIrZ3r95_0),.clk(gclk));
	jdff dff_B_INQJCmsq4_0(.din(w_dff_B_roIrZ3r95_0),.dout(w_dff_B_INQJCmsq4_0),.clk(gclk));
	jdff dff_B_S2YUjpry2_0(.din(w_dff_B_INQJCmsq4_0),.dout(w_dff_B_S2YUjpry2_0),.clk(gclk));
	jdff dff_B_hQvhKyRF0_0(.din(w_dff_B_S2YUjpry2_0),.dout(w_dff_B_hQvhKyRF0_0),.clk(gclk));
	jdff dff_B_gBAv87676_0(.din(w_dff_B_hQvhKyRF0_0),.dout(w_dff_B_gBAv87676_0),.clk(gclk));
	jdff dff_B_eMJv1uhA0_0(.din(w_dff_B_gBAv87676_0),.dout(w_dff_B_eMJv1uhA0_0),.clk(gclk));
	jdff dff_B_pbKGzT0D2_0(.din(w_dff_B_eMJv1uhA0_0),.dout(w_dff_B_pbKGzT0D2_0),.clk(gclk));
	jdff dff_B_xy3halQ76_0(.din(w_dff_B_pbKGzT0D2_0),.dout(w_dff_B_xy3halQ76_0),.clk(gclk));
	jdff dff_B_R019oiuF3_0(.din(w_dff_B_xy3halQ76_0),.dout(w_dff_B_R019oiuF3_0),.clk(gclk));
	jdff dff_B_Esw8TCrc8_0(.din(w_dff_B_R019oiuF3_0),.dout(w_dff_B_Esw8TCrc8_0),.clk(gclk));
	jdff dff_B_wU4KaYnM5_0(.din(w_dff_B_Esw8TCrc8_0),.dout(w_dff_B_wU4KaYnM5_0),.clk(gclk));
	jdff dff_B_Gmqk0wQw5_0(.din(w_dff_B_wU4KaYnM5_0),.dout(w_dff_B_Gmqk0wQw5_0),.clk(gclk));
	jdff dff_B_38OZjszQ5_0(.din(w_dff_B_Gmqk0wQw5_0),.dout(w_dff_B_38OZjszQ5_0),.clk(gclk));
	jdff dff_B_QLzSVlP16_0(.din(w_dff_B_38OZjszQ5_0),.dout(w_dff_B_QLzSVlP16_0),.clk(gclk));
	jdff dff_B_YnqMNmTs9_0(.din(w_dff_B_QLzSVlP16_0),.dout(w_dff_B_YnqMNmTs9_0),.clk(gclk));
	jdff dff_B_rJLGgzlb4_0(.din(w_dff_B_YnqMNmTs9_0),.dout(w_dff_B_rJLGgzlb4_0),.clk(gclk));
	jdff dff_B_SmFLyRQE5_0(.din(w_dff_B_rJLGgzlb4_0),.dout(w_dff_B_SmFLyRQE5_0),.clk(gclk));
	jdff dff_B_Lqoqfaep2_0(.din(w_dff_B_SmFLyRQE5_0),.dout(w_dff_B_Lqoqfaep2_0),.clk(gclk));
	jdff dff_B_Nqo52NhK6_0(.din(w_dff_B_Lqoqfaep2_0),.dout(w_dff_B_Nqo52NhK6_0),.clk(gclk));
	jdff dff_B_4FBdH4nN3_0(.din(w_dff_B_Nqo52NhK6_0),.dout(w_dff_B_4FBdH4nN3_0),.clk(gclk));
	jdff dff_B_HZFIiVPS6_0(.din(w_dff_B_4FBdH4nN3_0),.dout(w_dff_B_HZFIiVPS6_0),.clk(gclk));
	jdff dff_B_76wrGEuj0_0(.din(w_dff_B_HZFIiVPS6_0),.dout(w_dff_B_76wrGEuj0_0),.clk(gclk));
	jdff dff_B_tcHJDcFR1_1(.din(n576),.dout(w_dff_B_tcHJDcFR1_1),.clk(gclk));
	jdff dff_B_9WZlktg52_1(.din(w_dff_B_tcHJDcFR1_1),.dout(w_dff_B_9WZlktg52_1),.clk(gclk));
	jdff dff_B_70J7M71a6_1(.din(w_dff_B_9WZlktg52_1),.dout(w_dff_B_70J7M71a6_1),.clk(gclk));
	jdff dff_B_0bNe4Y0s1_1(.din(w_dff_B_70J7M71a6_1),.dout(w_dff_B_0bNe4Y0s1_1),.clk(gclk));
	jdff dff_B_nL0y6gwC7_1(.din(w_dff_B_0bNe4Y0s1_1),.dout(w_dff_B_nL0y6gwC7_1),.clk(gclk));
	jdff dff_B_oLYZUBoU8_1(.din(w_dff_B_nL0y6gwC7_1),.dout(w_dff_B_oLYZUBoU8_1),.clk(gclk));
	jdff dff_B_8e33wE607_1(.din(w_dff_B_oLYZUBoU8_1),.dout(w_dff_B_8e33wE607_1),.clk(gclk));
	jdff dff_B_cwZcdbUu5_1(.din(w_dff_B_8e33wE607_1),.dout(w_dff_B_cwZcdbUu5_1),.clk(gclk));
	jdff dff_B_AZBe0AUB8_1(.din(w_dff_B_cwZcdbUu5_1),.dout(w_dff_B_AZBe0AUB8_1),.clk(gclk));
	jdff dff_B_Q8rdd7TP9_1(.din(w_dff_B_AZBe0AUB8_1),.dout(w_dff_B_Q8rdd7TP9_1),.clk(gclk));
	jdff dff_B_ihvEdK217_1(.din(w_dff_B_Q8rdd7TP9_1),.dout(w_dff_B_ihvEdK217_1),.clk(gclk));
	jdff dff_B_HKvyjCvR1_1(.din(w_dff_B_ihvEdK217_1),.dout(w_dff_B_HKvyjCvR1_1),.clk(gclk));
	jdff dff_B_AHs9aKfS6_1(.din(w_dff_B_HKvyjCvR1_1),.dout(w_dff_B_AHs9aKfS6_1),.clk(gclk));
	jdff dff_B_cL4iQgTA6_1(.din(w_dff_B_AHs9aKfS6_1),.dout(w_dff_B_cL4iQgTA6_1),.clk(gclk));
	jdff dff_B_bBfx54BQ6_1(.din(w_dff_B_cL4iQgTA6_1),.dout(w_dff_B_bBfx54BQ6_1),.clk(gclk));
	jdff dff_B_K7JRSSOa8_1(.din(w_dff_B_bBfx54BQ6_1),.dout(w_dff_B_K7JRSSOa8_1),.clk(gclk));
	jdff dff_B_Y4PA8f7k0_1(.din(w_dff_B_K7JRSSOa8_1),.dout(w_dff_B_Y4PA8f7k0_1),.clk(gclk));
	jdff dff_B_UrbgIzAO2_1(.din(w_dff_B_Y4PA8f7k0_1),.dout(w_dff_B_UrbgIzAO2_1),.clk(gclk));
	jdff dff_B_z7F38Wm55_1(.din(w_dff_B_UrbgIzAO2_1),.dout(w_dff_B_z7F38Wm55_1),.clk(gclk));
	jdff dff_B_M7kYfyXx9_1(.din(w_dff_B_z7F38Wm55_1),.dout(w_dff_B_M7kYfyXx9_1),.clk(gclk));
	jdff dff_B_3tsAD5WQ5_1(.din(w_dff_B_M7kYfyXx9_1),.dout(w_dff_B_3tsAD5WQ5_1),.clk(gclk));
	jdff dff_B_vt5r96si8_1(.din(w_dff_B_3tsAD5WQ5_1),.dout(w_dff_B_vt5r96si8_1),.clk(gclk));
	jdff dff_B_vo4VCx545_1(.din(w_dff_B_vt5r96si8_1),.dout(w_dff_B_vo4VCx545_1),.clk(gclk));
	jdff dff_B_6boj367I4_1(.din(w_dff_B_vo4VCx545_1),.dout(w_dff_B_6boj367I4_1),.clk(gclk));
	jdff dff_B_9lkMKfrF3_1(.din(w_dff_B_6boj367I4_1),.dout(w_dff_B_9lkMKfrF3_1),.clk(gclk));
	jdff dff_B_qCwmP2Bx2_1(.din(w_dff_B_9lkMKfrF3_1),.dout(w_dff_B_qCwmP2Bx2_1),.clk(gclk));
	jdff dff_B_SnPkuC3J6_1(.din(w_dff_B_qCwmP2Bx2_1),.dout(w_dff_B_SnPkuC3J6_1),.clk(gclk));
	jdff dff_B_nJDSxQzd6_1(.din(w_dff_B_SnPkuC3J6_1),.dout(w_dff_B_nJDSxQzd6_1),.clk(gclk));
	jdff dff_B_M8fpqb9M1_1(.din(w_dff_B_nJDSxQzd6_1),.dout(w_dff_B_M8fpqb9M1_1),.clk(gclk));
	jdff dff_B_r7PLsI4y8_1(.din(w_dff_B_M8fpqb9M1_1),.dout(w_dff_B_r7PLsI4y8_1),.clk(gclk));
	jdff dff_B_ObSE17NU7_1(.din(w_dff_B_r7PLsI4y8_1),.dout(w_dff_B_ObSE17NU7_1),.clk(gclk));
	jdff dff_B_vpzfAeXc3_1(.din(w_dff_B_ObSE17NU7_1),.dout(w_dff_B_vpzfAeXc3_1),.clk(gclk));
	jdff dff_B_LTNSCy3T5_0(.din(n577),.dout(w_dff_B_LTNSCy3T5_0),.clk(gclk));
	jdff dff_B_Kq8KMKH56_0(.din(w_dff_B_LTNSCy3T5_0),.dout(w_dff_B_Kq8KMKH56_0),.clk(gclk));
	jdff dff_B_j5jfyqWt5_0(.din(w_dff_B_Kq8KMKH56_0),.dout(w_dff_B_j5jfyqWt5_0),.clk(gclk));
	jdff dff_B_oZlHD0Yl6_0(.din(w_dff_B_j5jfyqWt5_0),.dout(w_dff_B_oZlHD0Yl6_0),.clk(gclk));
	jdff dff_B_HepHhI2P1_0(.din(w_dff_B_oZlHD0Yl6_0),.dout(w_dff_B_HepHhI2P1_0),.clk(gclk));
	jdff dff_B_8Efjhcm60_0(.din(w_dff_B_HepHhI2P1_0),.dout(w_dff_B_8Efjhcm60_0),.clk(gclk));
	jdff dff_B_ONwbUvE51_0(.din(w_dff_B_8Efjhcm60_0),.dout(w_dff_B_ONwbUvE51_0),.clk(gclk));
	jdff dff_B_VPLQHarR4_0(.din(w_dff_B_ONwbUvE51_0),.dout(w_dff_B_VPLQHarR4_0),.clk(gclk));
	jdff dff_B_lYpDM30S8_0(.din(w_dff_B_VPLQHarR4_0),.dout(w_dff_B_lYpDM30S8_0),.clk(gclk));
	jdff dff_B_gkWjX6SZ2_0(.din(w_dff_B_lYpDM30S8_0),.dout(w_dff_B_gkWjX6SZ2_0),.clk(gclk));
	jdff dff_B_xHe8vVaJ7_0(.din(w_dff_B_gkWjX6SZ2_0),.dout(w_dff_B_xHe8vVaJ7_0),.clk(gclk));
	jdff dff_B_yMdjtUHY0_0(.din(w_dff_B_xHe8vVaJ7_0),.dout(w_dff_B_yMdjtUHY0_0),.clk(gclk));
	jdff dff_B_NJJYcFd94_0(.din(w_dff_B_yMdjtUHY0_0),.dout(w_dff_B_NJJYcFd94_0),.clk(gclk));
	jdff dff_B_JYBt8lY52_0(.din(w_dff_B_NJJYcFd94_0),.dout(w_dff_B_JYBt8lY52_0),.clk(gclk));
	jdff dff_B_rjhanWVQ0_0(.din(w_dff_B_JYBt8lY52_0),.dout(w_dff_B_rjhanWVQ0_0),.clk(gclk));
	jdff dff_B_N8FOrpxZ3_0(.din(w_dff_B_rjhanWVQ0_0),.dout(w_dff_B_N8FOrpxZ3_0),.clk(gclk));
	jdff dff_B_1qRgo3sm0_0(.din(w_dff_B_N8FOrpxZ3_0),.dout(w_dff_B_1qRgo3sm0_0),.clk(gclk));
	jdff dff_B_ZehycAL99_0(.din(w_dff_B_1qRgo3sm0_0),.dout(w_dff_B_ZehycAL99_0),.clk(gclk));
	jdff dff_B_F8h5tk9C4_0(.din(w_dff_B_ZehycAL99_0),.dout(w_dff_B_F8h5tk9C4_0),.clk(gclk));
	jdff dff_B_xxiTipoX3_0(.din(w_dff_B_F8h5tk9C4_0),.dout(w_dff_B_xxiTipoX3_0),.clk(gclk));
	jdff dff_B_Z51J2Y152_0(.din(w_dff_B_xxiTipoX3_0),.dout(w_dff_B_Z51J2Y152_0),.clk(gclk));
	jdff dff_B_FSbsuUJ49_0(.din(w_dff_B_Z51J2Y152_0),.dout(w_dff_B_FSbsuUJ49_0),.clk(gclk));
	jdff dff_B_c2Ni1VaX3_0(.din(w_dff_B_FSbsuUJ49_0),.dout(w_dff_B_c2Ni1VaX3_0),.clk(gclk));
	jdff dff_B_hJYS97bM5_0(.din(w_dff_B_c2Ni1VaX3_0),.dout(w_dff_B_hJYS97bM5_0),.clk(gclk));
	jdff dff_B_uZPAnIg84_0(.din(w_dff_B_hJYS97bM5_0),.dout(w_dff_B_uZPAnIg84_0),.clk(gclk));
	jdff dff_B_rxbIYFOS9_0(.din(w_dff_B_uZPAnIg84_0),.dout(w_dff_B_rxbIYFOS9_0),.clk(gclk));
	jdff dff_B_pjsjn3Lx1_0(.din(w_dff_B_rxbIYFOS9_0),.dout(w_dff_B_pjsjn3Lx1_0),.clk(gclk));
	jdff dff_B_AXIT0TSo2_0(.din(w_dff_B_pjsjn3Lx1_0),.dout(w_dff_B_AXIT0TSo2_0),.clk(gclk));
	jdff dff_B_MJXNOGvL3_0(.din(w_dff_B_AXIT0TSo2_0),.dout(w_dff_B_MJXNOGvL3_0),.clk(gclk));
	jdff dff_B_LtvlIL626_0(.din(w_dff_B_MJXNOGvL3_0),.dout(w_dff_B_LtvlIL626_0),.clk(gclk));
	jdff dff_B_SOMmHbp60_0(.din(w_dff_B_LtvlIL626_0),.dout(w_dff_B_SOMmHbp60_0),.clk(gclk));
	jdff dff_B_cOSHsCTW4_0(.din(w_dff_B_SOMmHbp60_0),.dout(w_dff_B_cOSHsCTW4_0),.clk(gclk));
	jdff dff_B_samYFRy26_1(.din(n570),.dout(w_dff_B_samYFRy26_1),.clk(gclk));
	jdff dff_B_v8zPcZTW1_1(.din(w_dff_B_samYFRy26_1),.dout(w_dff_B_v8zPcZTW1_1),.clk(gclk));
	jdff dff_B_ckoCJW2f2_1(.din(w_dff_B_v8zPcZTW1_1),.dout(w_dff_B_ckoCJW2f2_1),.clk(gclk));
	jdff dff_B_UGRsZrVB2_1(.din(w_dff_B_ckoCJW2f2_1),.dout(w_dff_B_UGRsZrVB2_1),.clk(gclk));
	jdff dff_B_Z7KUzV076_1(.din(w_dff_B_UGRsZrVB2_1),.dout(w_dff_B_Z7KUzV076_1),.clk(gclk));
	jdff dff_B_7ie9hnnY2_1(.din(w_dff_B_Z7KUzV076_1),.dout(w_dff_B_7ie9hnnY2_1),.clk(gclk));
	jdff dff_B_aCNE0rnf2_1(.din(w_dff_B_7ie9hnnY2_1),.dout(w_dff_B_aCNE0rnf2_1),.clk(gclk));
	jdff dff_B_zi007nmq0_1(.din(w_dff_B_aCNE0rnf2_1),.dout(w_dff_B_zi007nmq0_1),.clk(gclk));
	jdff dff_B_zHr8XPjf7_1(.din(w_dff_B_zi007nmq0_1),.dout(w_dff_B_zHr8XPjf7_1),.clk(gclk));
	jdff dff_B_QVu79ELB2_1(.din(w_dff_B_zHr8XPjf7_1),.dout(w_dff_B_QVu79ELB2_1),.clk(gclk));
	jdff dff_B_rpOfhEHv6_1(.din(w_dff_B_QVu79ELB2_1),.dout(w_dff_B_rpOfhEHv6_1),.clk(gclk));
	jdff dff_B_kW7Ee0re6_1(.din(w_dff_B_rpOfhEHv6_1),.dout(w_dff_B_kW7Ee0re6_1),.clk(gclk));
	jdff dff_B_O1W0Lwt47_1(.din(w_dff_B_kW7Ee0re6_1),.dout(w_dff_B_O1W0Lwt47_1),.clk(gclk));
	jdff dff_B_5P8jtjQX2_1(.din(w_dff_B_O1W0Lwt47_1),.dout(w_dff_B_5P8jtjQX2_1),.clk(gclk));
	jdff dff_B_WIAfGV192_1(.din(w_dff_B_5P8jtjQX2_1),.dout(w_dff_B_WIAfGV192_1),.clk(gclk));
	jdff dff_B_PX7GPVOA0_1(.din(w_dff_B_WIAfGV192_1),.dout(w_dff_B_PX7GPVOA0_1),.clk(gclk));
	jdff dff_B_0idppEZJ3_1(.din(w_dff_B_PX7GPVOA0_1),.dout(w_dff_B_0idppEZJ3_1),.clk(gclk));
	jdff dff_B_XoIYF6co2_1(.din(w_dff_B_0idppEZJ3_1),.dout(w_dff_B_XoIYF6co2_1),.clk(gclk));
	jdff dff_B_c93rijkr7_1(.din(w_dff_B_XoIYF6co2_1),.dout(w_dff_B_c93rijkr7_1),.clk(gclk));
	jdff dff_B_2xgoZpIf0_1(.din(w_dff_B_c93rijkr7_1),.dout(w_dff_B_2xgoZpIf0_1),.clk(gclk));
	jdff dff_B_WyJIYZMM9_1(.din(w_dff_B_2xgoZpIf0_1),.dout(w_dff_B_WyJIYZMM9_1),.clk(gclk));
	jdff dff_B_9aIXKL2h6_1(.din(w_dff_B_WyJIYZMM9_1),.dout(w_dff_B_9aIXKL2h6_1),.clk(gclk));
	jdff dff_B_ArO8sxJ99_1(.din(w_dff_B_9aIXKL2h6_1),.dout(w_dff_B_ArO8sxJ99_1),.clk(gclk));
	jdff dff_B_B6nLJOJA8_1(.din(w_dff_B_ArO8sxJ99_1),.dout(w_dff_B_B6nLJOJA8_1),.clk(gclk));
	jdff dff_B_dlr1o53y1_1(.din(w_dff_B_B6nLJOJA8_1),.dout(w_dff_B_dlr1o53y1_1),.clk(gclk));
	jdff dff_B_s88bDLvV1_1(.din(w_dff_B_dlr1o53y1_1),.dout(w_dff_B_s88bDLvV1_1),.clk(gclk));
	jdff dff_B_jhR3FbZ11_1(.din(w_dff_B_s88bDLvV1_1),.dout(w_dff_B_jhR3FbZ11_1),.clk(gclk));
	jdff dff_B_Hu4pUPJp1_1(.din(w_dff_B_jhR3FbZ11_1),.dout(w_dff_B_Hu4pUPJp1_1),.clk(gclk));
	jdff dff_B_bEJ5Q8kn7_1(.din(w_dff_B_Hu4pUPJp1_1),.dout(w_dff_B_bEJ5Q8kn7_1),.clk(gclk));
	jdff dff_B_6b8ZfWk11_1(.din(w_dff_B_bEJ5Q8kn7_1),.dout(w_dff_B_6b8ZfWk11_1),.clk(gclk));
	jdff dff_B_MqGZ9eEe7_1(.din(w_dff_B_6b8ZfWk11_1),.dout(w_dff_B_MqGZ9eEe7_1),.clk(gclk));
	jdff dff_B_9Ggorrgr6_0(.din(n571),.dout(w_dff_B_9Ggorrgr6_0),.clk(gclk));
	jdff dff_B_ug1THLAA8_0(.din(w_dff_B_9Ggorrgr6_0),.dout(w_dff_B_ug1THLAA8_0),.clk(gclk));
	jdff dff_B_p2njF8Wy0_0(.din(w_dff_B_ug1THLAA8_0),.dout(w_dff_B_p2njF8Wy0_0),.clk(gclk));
	jdff dff_B_7BqpENEe4_0(.din(w_dff_B_p2njF8Wy0_0),.dout(w_dff_B_7BqpENEe4_0),.clk(gclk));
	jdff dff_B_VQ8RXdVW7_0(.din(w_dff_B_7BqpENEe4_0),.dout(w_dff_B_VQ8RXdVW7_0),.clk(gclk));
	jdff dff_B_m0Aee3JC2_0(.din(w_dff_B_VQ8RXdVW7_0),.dout(w_dff_B_m0Aee3JC2_0),.clk(gclk));
	jdff dff_B_5rh7trX38_0(.din(w_dff_B_m0Aee3JC2_0),.dout(w_dff_B_5rh7trX38_0),.clk(gclk));
	jdff dff_B_yGaqTppP6_0(.din(w_dff_B_5rh7trX38_0),.dout(w_dff_B_yGaqTppP6_0),.clk(gclk));
	jdff dff_B_eg2ny05c4_0(.din(w_dff_B_yGaqTppP6_0),.dout(w_dff_B_eg2ny05c4_0),.clk(gclk));
	jdff dff_B_0VrRwCMq1_0(.din(w_dff_B_eg2ny05c4_0),.dout(w_dff_B_0VrRwCMq1_0),.clk(gclk));
	jdff dff_B_s2sZnpMk3_0(.din(w_dff_B_0VrRwCMq1_0),.dout(w_dff_B_s2sZnpMk3_0),.clk(gclk));
	jdff dff_B_214eGyoe3_0(.din(w_dff_B_s2sZnpMk3_0),.dout(w_dff_B_214eGyoe3_0),.clk(gclk));
	jdff dff_B_YmbertBM1_0(.din(w_dff_B_214eGyoe3_0),.dout(w_dff_B_YmbertBM1_0),.clk(gclk));
	jdff dff_B_iNuIMc615_0(.din(w_dff_B_YmbertBM1_0),.dout(w_dff_B_iNuIMc615_0),.clk(gclk));
	jdff dff_B_UgRoswJS6_0(.din(w_dff_B_iNuIMc615_0),.dout(w_dff_B_UgRoswJS6_0),.clk(gclk));
	jdff dff_B_ol2PWX3g7_0(.din(w_dff_B_UgRoswJS6_0),.dout(w_dff_B_ol2PWX3g7_0),.clk(gclk));
	jdff dff_B_QqvKBaoG2_0(.din(w_dff_B_ol2PWX3g7_0),.dout(w_dff_B_QqvKBaoG2_0),.clk(gclk));
	jdff dff_B_1R9OOYbQ0_0(.din(w_dff_B_QqvKBaoG2_0),.dout(w_dff_B_1R9OOYbQ0_0),.clk(gclk));
	jdff dff_B_s3RzwFa12_0(.din(w_dff_B_1R9OOYbQ0_0),.dout(w_dff_B_s3RzwFa12_0),.clk(gclk));
	jdff dff_B_3BVcZBgW8_0(.din(w_dff_B_s3RzwFa12_0),.dout(w_dff_B_3BVcZBgW8_0),.clk(gclk));
	jdff dff_B_2G1Aa0kZ9_0(.din(w_dff_B_3BVcZBgW8_0),.dout(w_dff_B_2G1Aa0kZ9_0),.clk(gclk));
	jdff dff_B_45XYBINy1_0(.din(w_dff_B_2G1Aa0kZ9_0),.dout(w_dff_B_45XYBINy1_0),.clk(gclk));
	jdff dff_B_ynroTsRQ3_0(.din(w_dff_B_45XYBINy1_0),.dout(w_dff_B_ynroTsRQ3_0),.clk(gclk));
	jdff dff_B_EN9YDQum1_0(.din(w_dff_B_ynroTsRQ3_0),.dout(w_dff_B_EN9YDQum1_0),.clk(gclk));
	jdff dff_B_NkzF3NyE6_0(.din(w_dff_B_EN9YDQum1_0),.dout(w_dff_B_NkzF3NyE6_0),.clk(gclk));
	jdff dff_B_jhDoapJP3_0(.din(w_dff_B_NkzF3NyE6_0),.dout(w_dff_B_jhDoapJP3_0),.clk(gclk));
	jdff dff_B_ip3MrRlz8_0(.din(w_dff_B_jhDoapJP3_0),.dout(w_dff_B_ip3MrRlz8_0),.clk(gclk));
	jdff dff_B_1F86GwH13_0(.din(w_dff_B_ip3MrRlz8_0),.dout(w_dff_B_1F86GwH13_0),.clk(gclk));
	jdff dff_B_7JgE58Gx7_0(.din(w_dff_B_1F86GwH13_0),.dout(w_dff_B_7JgE58Gx7_0),.clk(gclk));
	jdff dff_B_ppIkGrU39_0(.din(w_dff_B_7JgE58Gx7_0),.dout(w_dff_B_ppIkGrU39_0),.clk(gclk));
	jdff dff_B_znPY8YBC7_0(.din(w_dff_B_ppIkGrU39_0),.dout(w_dff_B_znPY8YBC7_0),.clk(gclk));
	jdff dff_B_Cz4WtRxM5_1(.din(n564),.dout(w_dff_B_Cz4WtRxM5_1),.clk(gclk));
	jdff dff_B_hX4DDc072_1(.din(w_dff_B_Cz4WtRxM5_1),.dout(w_dff_B_hX4DDc072_1),.clk(gclk));
	jdff dff_B_vO4oC1wC1_1(.din(w_dff_B_hX4DDc072_1),.dout(w_dff_B_vO4oC1wC1_1),.clk(gclk));
	jdff dff_B_N4QkzRah0_1(.din(w_dff_B_vO4oC1wC1_1),.dout(w_dff_B_N4QkzRah0_1),.clk(gclk));
	jdff dff_B_noq5BmFc8_1(.din(w_dff_B_N4QkzRah0_1),.dout(w_dff_B_noq5BmFc8_1),.clk(gclk));
	jdff dff_B_wot6X4XY2_1(.din(w_dff_B_noq5BmFc8_1),.dout(w_dff_B_wot6X4XY2_1),.clk(gclk));
	jdff dff_B_SoZ8p6EM4_1(.din(w_dff_B_wot6X4XY2_1),.dout(w_dff_B_SoZ8p6EM4_1),.clk(gclk));
	jdff dff_B_AzSalxIW5_1(.din(w_dff_B_SoZ8p6EM4_1),.dout(w_dff_B_AzSalxIW5_1),.clk(gclk));
	jdff dff_B_8lhDmClm5_1(.din(w_dff_B_AzSalxIW5_1),.dout(w_dff_B_8lhDmClm5_1),.clk(gclk));
	jdff dff_B_upPOgiH16_1(.din(w_dff_B_8lhDmClm5_1),.dout(w_dff_B_upPOgiH16_1),.clk(gclk));
	jdff dff_B_vdn2loSW0_1(.din(w_dff_B_upPOgiH16_1),.dout(w_dff_B_vdn2loSW0_1),.clk(gclk));
	jdff dff_B_ovjpKjld3_1(.din(w_dff_B_vdn2loSW0_1),.dout(w_dff_B_ovjpKjld3_1),.clk(gclk));
	jdff dff_B_iF3FEifp1_1(.din(w_dff_B_ovjpKjld3_1),.dout(w_dff_B_iF3FEifp1_1),.clk(gclk));
	jdff dff_B_bCE7ygWT0_1(.din(w_dff_B_iF3FEifp1_1),.dout(w_dff_B_bCE7ygWT0_1),.clk(gclk));
	jdff dff_B_2WFUWllr6_1(.din(w_dff_B_bCE7ygWT0_1),.dout(w_dff_B_2WFUWllr6_1),.clk(gclk));
	jdff dff_B_Hn1ui6Rj0_1(.din(w_dff_B_2WFUWllr6_1),.dout(w_dff_B_Hn1ui6Rj0_1),.clk(gclk));
	jdff dff_B_6Ko2H74B0_1(.din(w_dff_B_Hn1ui6Rj0_1),.dout(w_dff_B_6Ko2H74B0_1),.clk(gclk));
	jdff dff_B_kOy0lbw30_1(.din(w_dff_B_6Ko2H74B0_1),.dout(w_dff_B_kOy0lbw30_1),.clk(gclk));
	jdff dff_B_v1EP3kgw5_1(.din(w_dff_B_kOy0lbw30_1),.dout(w_dff_B_v1EP3kgw5_1),.clk(gclk));
	jdff dff_B_9zav3DDa1_1(.din(w_dff_B_v1EP3kgw5_1),.dout(w_dff_B_9zav3DDa1_1),.clk(gclk));
	jdff dff_B_orFt2uhv8_1(.din(w_dff_B_9zav3DDa1_1),.dout(w_dff_B_orFt2uhv8_1),.clk(gclk));
	jdff dff_B_lOUweBA10_1(.din(w_dff_B_orFt2uhv8_1),.dout(w_dff_B_lOUweBA10_1),.clk(gclk));
	jdff dff_B_pAQzK9x95_1(.din(w_dff_B_lOUweBA10_1),.dout(w_dff_B_pAQzK9x95_1),.clk(gclk));
	jdff dff_B_4FvCS16N8_1(.din(w_dff_B_pAQzK9x95_1),.dout(w_dff_B_4FvCS16N8_1),.clk(gclk));
	jdff dff_B_KXpwsZS63_1(.din(w_dff_B_4FvCS16N8_1),.dout(w_dff_B_KXpwsZS63_1),.clk(gclk));
	jdff dff_B_kd2gB3L62_1(.din(w_dff_B_KXpwsZS63_1),.dout(w_dff_B_kd2gB3L62_1),.clk(gclk));
	jdff dff_B_QVdUCIrd3_1(.din(w_dff_B_kd2gB3L62_1),.dout(w_dff_B_QVdUCIrd3_1),.clk(gclk));
	jdff dff_B_Q3XMAHfH4_1(.din(w_dff_B_QVdUCIrd3_1),.dout(w_dff_B_Q3XMAHfH4_1),.clk(gclk));
	jdff dff_B_LTDwHoxl1_1(.din(w_dff_B_Q3XMAHfH4_1),.dout(w_dff_B_LTDwHoxl1_1),.clk(gclk));
	jdff dff_B_fYp7rwhu5_1(.din(w_dff_B_LTDwHoxl1_1),.dout(w_dff_B_fYp7rwhu5_1),.clk(gclk));
	jdff dff_B_KVAaujiM8_0(.din(n565),.dout(w_dff_B_KVAaujiM8_0),.clk(gclk));
	jdff dff_B_qau2pyoL4_0(.din(w_dff_B_KVAaujiM8_0),.dout(w_dff_B_qau2pyoL4_0),.clk(gclk));
	jdff dff_B_cERkMASt4_0(.din(w_dff_B_qau2pyoL4_0),.dout(w_dff_B_cERkMASt4_0),.clk(gclk));
	jdff dff_B_CL07I3La5_0(.din(w_dff_B_cERkMASt4_0),.dout(w_dff_B_CL07I3La5_0),.clk(gclk));
	jdff dff_B_VekVdwrf9_0(.din(w_dff_B_CL07I3La5_0),.dout(w_dff_B_VekVdwrf9_0),.clk(gclk));
	jdff dff_B_gw8GjGg32_0(.din(w_dff_B_VekVdwrf9_0),.dout(w_dff_B_gw8GjGg32_0),.clk(gclk));
	jdff dff_B_dIFaRqJ38_0(.din(w_dff_B_gw8GjGg32_0),.dout(w_dff_B_dIFaRqJ38_0),.clk(gclk));
	jdff dff_B_s0SY6L6P3_0(.din(w_dff_B_dIFaRqJ38_0),.dout(w_dff_B_s0SY6L6P3_0),.clk(gclk));
	jdff dff_B_xZqCvfWm9_0(.din(w_dff_B_s0SY6L6P3_0),.dout(w_dff_B_xZqCvfWm9_0),.clk(gclk));
	jdff dff_B_rR833kho1_0(.din(w_dff_B_xZqCvfWm9_0),.dout(w_dff_B_rR833kho1_0),.clk(gclk));
	jdff dff_B_f4Hjsnyc5_0(.din(w_dff_B_rR833kho1_0),.dout(w_dff_B_f4Hjsnyc5_0),.clk(gclk));
	jdff dff_B_HIFK3fD29_0(.din(w_dff_B_f4Hjsnyc5_0),.dout(w_dff_B_HIFK3fD29_0),.clk(gclk));
	jdff dff_B_7GAWPKnJ8_0(.din(w_dff_B_HIFK3fD29_0),.dout(w_dff_B_7GAWPKnJ8_0),.clk(gclk));
	jdff dff_B_pMq7HHim5_0(.din(w_dff_B_7GAWPKnJ8_0),.dout(w_dff_B_pMq7HHim5_0),.clk(gclk));
	jdff dff_B_Hpll6Zaz4_0(.din(w_dff_B_pMq7HHim5_0),.dout(w_dff_B_Hpll6Zaz4_0),.clk(gclk));
	jdff dff_B_3bOyimU30_0(.din(w_dff_B_Hpll6Zaz4_0),.dout(w_dff_B_3bOyimU30_0),.clk(gclk));
	jdff dff_B_0r66Rra19_0(.din(w_dff_B_3bOyimU30_0),.dout(w_dff_B_0r66Rra19_0),.clk(gclk));
	jdff dff_B_sc2CgKKH6_0(.din(w_dff_B_0r66Rra19_0),.dout(w_dff_B_sc2CgKKH6_0),.clk(gclk));
	jdff dff_B_bhTrfgfj9_0(.din(w_dff_B_sc2CgKKH6_0),.dout(w_dff_B_bhTrfgfj9_0),.clk(gclk));
	jdff dff_B_zBU8oC3W8_0(.din(w_dff_B_bhTrfgfj9_0),.dout(w_dff_B_zBU8oC3W8_0),.clk(gclk));
	jdff dff_B_Wp6clGhC6_0(.din(w_dff_B_zBU8oC3W8_0),.dout(w_dff_B_Wp6clGhC6_0),.clk(gclk));
	jdff dff_B_gyKCnTy02_0(.din(w_dff_B_Wp6clGhC6_0),.dout(w_dff_B_gyKCnTy02_0),.clk(gclk));
	jdff dff_B_mue6Cm2y2_0(.din(w_dff_B_gyKCnTy02_0),.dout(w_dff_B_mue6Cm2y2_0),.clk(gclk));
	jdff dff_B_sBWbgYsk6_0(.din(w_dff_B_mue6Cm2y2_0),.dout(w_dff_B_sBWbgYsk6_0),.clk(gclk));
	jdff dff_B_DobI48jM4_0(.din(w_dff_B_sBWbgYsk6_0),.dout(w_dff_B_DobI48jM4_0),.clk(gclk));
	jdff dff_B_Iae9FgpR7_0(.din(w_dff_B_DobI48jM4_0),.dout(w_dff_B_Iae9FgpR7_0),.clk(gclk));
	jdff dff_B_SW8NICzc1_0(.din(w_dff_B_Iae9FgpR7_0),.dout(w_dff_B_SW8NICzc1_0),.clk(gclk));
	jdff dff_B_jrdi6QfX3_0(.din(w_dff_B_SW8NICzc1_0),.dout(w_dff_B_jrdi6QfX3_0),.clk(gclk));
	jdff dff_B_FuBS1k7T9_0(.din(w_dff_B_jrdi6QfX3_0),.dout(w_dff_B_FuBS1k7T9_0),.clk(gclk));
	jdff dff_B_norHvl765_0(.din(w_dff_B_FuBS1k7T9_0),.dout(w_dff_B_norHvl765_0),.clk(gclk));
	jdff dff_B_M14cBlRa3_1(.din(n558),.dout(w_dff_B_M14cBlRa3_1),.clk(gclk));
	jdff dff_B_5uJWKH683_1(.din(w_dff_B_M14cBlRa3_1),.dout(w_dff_B_5uJWKH683_1),.clk(gclk));
	jdff dff_B_ORDz8jHr0_1(.din(w_dff_B_5uJWKH683_1),.dout(w_dff_B_ORDz8jHr0_1),.clk(gclk));
	jdff dff_B_Y9B4bwQp3_1(.din(w_dff_B_ORDz8jHr0_1),.dout(w_dff_B_Y9B4bwQp3_1),.clk(gclk));
	jdff dff_B_SXpLQFZD3_1(.din(w_dff_B_Y9B4bwQp3_1),.dout(w_dff_B_SXpLQFZD3_1),.clk(gclk));
	jdff dff_B_HVIgRfMF6_1(.din(w_dff_B_SXpLQFZD3_1),.dout(w_dff_B_HVIgRfMF6_1),.clk(gclk));
	jdff dff_B_9zRL7yZl3_1(.din(w_dff_B_HVIgRfMF6_1),.dout(w_dff_B_9zRL7yZl3_1),.clk(gclk));
	jdff dff_B_5P3N4tZX5_1(.din(w_dff_B_9zRL7yZl3_1),.dout(w_dff_B_5P3N4tZX5_1),.clk(gclk));
	jdff dff_B_1UtBCH3i9_1(.din(w_dff_B_5P3N4tZX5_1),.dout(w_dff_B_1UtBCH3i9_1),.clk(gclk));
	jdff dff_B_6qhYjcvS4_1(.din(w_dff_B_1UtBCH3i9_1),.dout(w_dff_B_6qhYjcvS4_1),.clk(gclk));
	jdff dff_B_yBwEhq9Y5_1(.din(w_dff_B_6qhYjcvS4_1),.dout(w_dff_B_yBwEhq9Y5_1),.clk(gclk));
	jdff dff_B_vKMEa47W2_1(.din(w_dff_B_yBwEhq9Y5_1),.dout(w_dff_B_vKMEa47W2_1),.clk(gclk));
	jdff dff_B_tSIC5Z2N9_1(.din(w_dff_B_vKMEa47W2_1),.dout(w_dff_B_tSIC5Z2N9_1),.clk(gclk));
	jdff dff_B_R4LvJLUz9_1(.din(w_dff_B_tSIC5Z2N9_1),.dout(w_dff_B_R4LvJLUz9_1),.clk(gclk));
	jdff dff_B_f4LXkT1g6_1(.din(w_dff_B_R4LvJLUz9_1),.dout(w_dff_B_f4LXkT1g6_1),.clk(gclk));
	jdff dff_B_k0qWQIyd3_1(.din(w_dff_B_f4LXkT1g6_1),.dout(w_dff_B_k0qWQIyd3_1),.clk(gclk));
	jdff dff_B_I3VXEj6g5_1(.din(w_dff_B_k0qWQIyd3_1),.dout(w_dff_B_I3VXEj6g5_1),.clk(gclk));
	jdff dff_B_nHVGy9fB0_1(.din(w_dff_B_I3VXEj6g5_1),.dout(w_dff_B_nHVGy9fB0_1),.clk(gclk));
	jdff dff_B_JLI54C3i4_1(.din(w_dff_B_nHVGy9fB0_1),.dout(w_dff_B_JLI54C3i4_1),.clk(gclk));
	jdff dff_B_6GlsA9Pl1_1(.din(w_dff_B_JLI54C3i4_1),.dout(w_dff_B_6GlsA9Pl1_1),.clk(gclk));
	jdff dff_B_baVt6ZSl9_1(.din(w_dff_B_6GlsA9Pl1_1),.dout(w_dff_B_baVt6ZSl9_1),.clk(gclk));
	jdff dff_B_3xuXNVe27_1(.din(w_dff_B_baVt6ZSl9_1),.dout(w_dff_B_3xuXNVe27_1),.clk(gclk));
	jdff dff_B_DytvXwob2_1(.din(w_dff_B_3xuXNVe27_1),.dout(w_dff_B_DytvXwob2_1),.clk(gclk));
	jdff dff_B_ddtiVxdK6_1(.din(w_dff_B_DytvXwob2_1),.dout(w_dff_B_ddtiVxdK6_1),.clk(gclk));
	jdff dff_B_bTFY9pP37_1(.din(w_dff_B_ddtiVxdK6_1),.dout(w_dff_B_bTFY9pP37_1),.clk(gclk));
	jdff dff_B_Z8zTQmtf6_1(.din(w_dff_B_bTFY9pP37_1),.dout(w_dff_B_Z8zTQmtf6_1),.clk(gclk));
	jdff dff_B_vlazR5UV4_1(.din(w_dff_B_Z8zTQmtf6_1),.dout(w_dff_B_vlazR5UV4_1),.clk(gclk));
	jdff dff_B_ycAvA3bo6_1(.din(w_dff_B_vlazR5UV4_1),.dout(w_dff_B_ycAvA3bo6_1),.clk(gclk));
	jdff dff_B_8BjQK9zd0_1(.din(w_dff_B_ycAvA3bo6_1),.dout(w_dff_B_8BjQK9zd0_1),.clk(gclk));
	jdff dff_B_K955MgLd2_0(.din(n559),.dout(w_dff_B_K955MgLd2_0),.clk(gclk));
	jdff dff_B_0bFrWliJ3_0(.din(w_dff_B_K955MgLd2_0),.dout(w_dff_B_0bFrWliJ3_0),.clk(gclk));
	jdff dff_B_u3xurdFd9_0(.din(w_dff_B_0bFrWliJ3_0),.dout(w_dff_B_u3xurdFd9_0),.clk(gclk));
	jdff dff_B_qEPqL1lz8_0(.din(w_dff_B_u3xurdFd9_0),.dout(w_dff_B_qEPqL1lz8_0),.clk(gclk));
	jdff dff_B_FRy9Sbe00_0(.din(w_dff_B_qEPqL1lz8_0),.dout(w_dff_B_FRy9Sbe00_0),.clk(gclk));
	jdff dff_B_usV5zQIJ5_0(.din(w_dff_B_FRy9Sbe00_0),.dout(w_dff_B_usV5zQIJ5_0),.clk(gclk));
	jdff dff_B_ZCAcNYzC6_0(.din(w_dff_B_usV5zQIJ5_0),.dout(w_dff_B_ZCAcNYzC6_0),.clk(gclk));
	jdff dff_B_mfWO26go4_0(.din(w_dff_B_ZCAcNYzC6_0),.dout(w_dff_B_mfWO26go4_0),.clk(gclk));
	jdff dff_B_7j8eGKHU3_0(.din(w_dff_B_mfWO26go4_0),.dout(w_dff_B_7j8eGKHU3_0),.clk(gclk));
	jdff dff_B_CReshun12_0(.din(w_dff_B_7j8eGKHU3_0),.dout(w_dff_B_CReshun12_0),.clk(gclk));
	jdff dff_B_6TAgUcO31_0(.din(w_dff_B_CReshun12_0),.dout(w_dff_B_6TAgUcO31_0),.clk(gclk));
	jdff dff_B_GjDh4VHQ9_0(.din(w_dff_B_6TAgUcO31_0),.dout(w_dff_B_GjDh4VHQ9_0),.clk(gclk));
	jdff dff_B_6hsWPD6h3_0(.din(w_dff_B_GjDh4VHQ9_0),.dout(w_dff_B_6hsWPD6h3_0),.clk(gclk));
	jdff dff_B_2SC8oVLH8_0(.din(w_dff_B_6hsWPD6h3_0),.dout(w_dff_B_2SC8oVLH8_0),.clk(gclk));
	jdff dff_B_ZpiByu876_0(.din(w_dff_B_2SC8oVLH8_0),.dout(w_dff_B_ZpiByu876_0),.clk(gclk));
	jdff dff_B_FzaFPmnd4_0(.din(w_dff_B_ZpiByu876_0),.dout(w_dff_B_FzaFPmnd4_0),.clk(gclk));
	jdff dff_B_EkXR9rup5_0(.din(w_dff_B_FzaFPmnd4_0),.dout(w_dff_B_EkXR9rup5_0),.clk(gclk));
	jdff dff_B_9EgvbX9c9_0(.din(w_dff_B_EkXR9rup5_0),.dout(w_dff_B_9EgvbX9c9_0),.clk(gclk));
	jdff dff_B_qGVosCTG1_0(.din(w_dff_B_9EgvbX9c9_0),.dout(w_dff_B_qGVosCTG1_0),.clk(gclk));
	jdff dff_B_1DYf3zti2_0(.din(w_dff_B_qGVosCTG1_0),.dout(w_dff_B_1DYf3zti2_0),.clk(gclk));
	jdff dff_B_k3atWQ127_0(.din(w_dff_B_1DYf3zti2_0),.dout(w_dff_B_k3atWQ127_0),.clk(gclk));
	jdff dff_B_KqOdcc988_0(.din(w_dff_B_k3atWQ127_0),.dout(w_dff_B_KqOdcc988_0),.clk(gclk));
	jdff dff_B_0ldvzPUH2_0(.din(w_dff_B_KqOdcc988_0),.dout(w_dff_B_0ldvzPUH2_0),.clk(gclk));
	jdff dff_B_VRpTGNTt2_0(.din(w_dff_B_0ldvzPUH2_0),.dout(w_dff_B_VRpTGNTt2_0),.clk(gclk));
	jdff dff_B_XRq1WP6W0_0(.din(w_dff_B_VRpTGNTt2_0),.dout(w_dff_B_XRq1WP6W0_0),.clk(gclk));
	jdff dff_B_STiWvv1c6_0(.din(w_dff_B_XRq1WP6W0_0),.dout(w_dff_B_STiWvv1c6_0),.clk(gclk));
	jdff dff_B_5GKmYqIk5_0(.din(w_dff_B_STiWvv1c6_0),.dout(w_dff_B_5GKmYqIk5_0),.clk(gclk));
	jdff dff_B_dxJBpCHf6_0(.din(w_dff_B_5GKmYqIk5_0),.dout(w_dff_B_dxJBpCHf6_0),.clk(gclk));
	jdff dff_B_qICniHxc5_0(.din(w_dff_B_dxJBpCHf6_0),.dout(w_dff_B_qICniHxc5_0),.clk(gclk));
	jdff dff_B_WwGsn7LM4_1(.din(n552),.dout(w_dff_B_WwGsn7LM4_1),.clk(gclk));
	jdff dff_B_f5ScmcyJ6_1(.din(w_dff_B_WwGsn7LM4_1),.dout(w_dff_B_f5ScmcyJ6_1),.clk(gclk));
	jdff dff_B_aCLgWyNj8_1(.din(w_dff_B_f5ScmcyJ6_1),.dout(w_dff_B_aCLgWyNj8_1),.clk(gclk));
	jdff dff_B_NSG7h4PV7_1(.din(w_dff_B_aCLgWyNj8_1),.dout(w_dff_B_NSG7h4PV7_1),.clk(gclk));
	jdff dff_B_Nm7SQCST1_1(.din(w_dff_B_NSG7h4PV7_1),.dout(w_dff_B_Nm7SQCST1_1),.clk(gclk));
	jdff dff_B_jHSFzABG5_1(.din(w_dff_B_Nm7SQCST1_1),.dout(w_dff_B_jHSFzABG5_1),.clk(gclk));
	jdff dff_B_pdZ06Urv9_1(.din(w_dff_B_jHSFzABG5_1),.dout(w_dff_B_pdZ06Urv9_1),.clk(gclk));
	jdff dff_B_nG97F2Ex8_1(.din(w_dff_B_pdZ06Urv9_1),.dout(w_dff_B_nG97F2Ex8_1),.clk(gclk));
	jdff dff_B_c7ZVKITz0_1(.din(w_dff_B_nG97F2Ex8_1),.dout(w_dff_B_c7ZVKITz0_1),.clk(gclk));
	jdff dff_B_Gt7NUnjt0_1(.din(w_dff_B_c7ZVKITz0_1),.dout(w_dff_B_Gt7NUnjt0_1),.clk(gclk));
	jdff dff_B_VbnvtDzw0_1(.din(w_dff_B_Gt7NUnjt0_1),.dout(w_dff_B_VbnvtDzw0_1),.clk(gclk));
	jdff dff_B_sCBkMioo1_1(.din(w_dff_B_VbnvtDzw0_1),.dout(w_dff_B_sCBkMioo1_1),.clk(gclk));
	jdff dff_B_mlholDQR6_1(.din(w_dff_B_sCBkMioo1_1),.dout(w_dff_B_mlholDQR6_1),.clk(gclk));
	jdff dff_B_ASDanwoZ2_1(.din(w_dff_B_mlholDQR6_1),.dout(w_dff_B_ASDanwoZ2_1),.clk(gclk));
	jdff dff_B_NmEhouA63_1(.din(w_dff_B_ASDanwoZ2_1),.dout(w_dff_B_NmEhouA63_1),.clk(gclk));
	jdff dff_B_puvOBG1g8_1(.din(w_dff_B_NmEhouA63_1),.dout(w_dff_B_puvOBG1g8_1),.clk(gclk));
	jdff dff_B_3ALvuP1T5_1(.din(w_dff_B_puvOBG1g8_1),.dout(w_dff_B_3ALvuP1T5_1),.clk(gclk));
	jdff dff_B_rA6yFVJI6_1(.din(w_dff_B_3ALvuP1T5_1),.dout(w_dff_B_rA6yFVJI6_1),.clk(gclk));
	jdff dff_B_4CQIpvhh0_1(.din(w_dff_B_rA6yFVJI6_1),.dout(w_dff_B_4CQIpvhh0_1),.clk(gclk));
	jdff dff_B_9rjun1La0_1(.din(w_dff_B_4CQIpvhh0_1),.dout(w_dff_B_9rjun1La0_1),.clk(gclk));
	jdff dff_B_OxW1yAXT0_1(.din(w_dff_B_9rjun1La0_1),.dout(w_dff_B_OxW1yAXT0_1),.clk(gclk));
	jdff dff_B_cKJveguF8_1(.din(w_dff_B_OxW1yAXT0_1),.dout(w_dff_B_cKJveguF8_1),.clk(gclk));
	jdff dff_B_tHXTKG4t0_1(.din(w_dff_B_cKJveguF8_1),.dout(w_dff_B_tHXTKG4t0_1),.clk(gclk));
	jdff dff_B_dQwJwBfQ7_1(.din(w_dff_B_tHXTKG4t0_1),.dout(w_dff_B_dQwJwBfQ7_1),.clk(gclk));
	jdff dff_B_OgDtmjCn6_1(.din(w_dff_B_dQwJwBfQ7_1),.dout(w_dff_B_OgDtmjCn6_1),.clk(gclk));
	jdff dff_B_ET19mGkv9_1(.din(w_dff_B_OgDtmjCn6_1),.dout(w_dff_B_ET19mGkv9_1),.clk(gclk));
	jdff dff_B_dbGglKDe6_1(.din(w_dff_B_ET19mGkv9_1),.dout(w_dff_B_dbGglKDe6_1),.clk(gclk));
	jdff dff_B_2YMJeXnr4_1(.din(w_dff_B_dbGglKDe6_1),.dout(w_dff_B_2YMJeXnr4_1),.clk(gclk));
	jdff dff_B_jB9dqKE43_0(.din(n553),.dout(w_dff_B_jB9dqKE43_0),.clk(gclk));
	jdff dff_B_Xa6ExE5U8_0(.din(w_dff_B_jB9dqKE43_0),.dout(w_dff_B_Xa6ExE5U8_0),.clk(gclk));
	jdff dff_B_Xe2eAvbj2_0(.din(w_dff_B_Xa6ExE5U8_0),.dout(w_dff_B_Xe2eAvbj2_0),.clk(gclk));
	jdff dff_B_utP8Au306_0(.din(w_dff_B_Xe2eAvbj2_0),.dout(w_dff_B_utP8Au306_0),.clk(gclk));
	jdff dff_B_pJQs1Bcx6_0(.din(w_dff_B_utP8Au306_0),.dout(w_dff_B_pJQs1Bcx6_0),.clk(gclk));
	jdff dff_B_7Z1s3hJ50_0(.din(w_dff_B_pJQs1Bcx6_0),.dout(w_dff_B_7Z1s3hJ50_0),.clk(gclk));
	jdff dff_B_2yVGrjXx0_0(.din(w_dff_B_7Z1s3hJ50_0),.dout(w_dff_B_2yVGrjXx0_0),.clk(gclk));
	jdff dff_B_PshY9lv55_0(.din(w_dff_B_2yVGrjXx0_0),.dout(w_dff_B_PshY9lv55_0),.clk(gclk));
	jdff dff_B_CkzlWNUu7_0(.din(w_dff_B_PshY9lv55_0),.dout(w_dff_B_CkzlWNUu7_0),.clk(gclk));
	jdff dff_B_XrQqis6x0_0(.din(w_dff_B_CkzlWNUu7_0),.dout(w_dff_B_XrQqis6x0_0),.clk(gclk));
	jdff dff_B_zd0ukQpz7_0(.din(w_dff_B_XrQqis6x0_0),.dout(w_dff_B_zd0ukQpz7_0),.clk(gclk));
	jdff dff_B_qB9AiSgF4_0(.din(w_dff_B_zd0ukQpz7_0),.dout(w_dff_B_qB9AiSgF4_0),.clk(gclk));
	jdff dff_B_6lqgn5wN8_0(.din(w_dff_B_qB9AiSgF4_0),.dout(w_dff_B_6lqgn5wN8_0),.clk(gclk));
	jdff dff_B_UurPIyiQ3_0(.din(w_dff_B_6lqgn5wN8_0),.dout(w_dff_B_UurPIyiQ3_0),.clk(gclk));
	jdff dff_B_AZTO00TC7_0(.din(w_dff_B_UurPIyiQ3_0),.dout(w_dff_B_AZTO00TC7_0),.clk(gclk));
	jdff dff_B_1zuWxfB68_0(.din(w_dff_B_AZTO00TC7_0),.dout(w_dff_B_1zuWxfB68_0),.clk(gclk));
	jdff dff_B_yVylfGHH5_0(.din(w_dff_B_1zuWxfB68_0),.dout(w_dff_B_yVylfGHH5_0),.clk(gclk));
	jdff dff_B_2pixfssf7_0(.din(w_dff_B_yVylfGHH5_0),.dout(w_dff_B_2pixfssf7_0),.clk(gclk));
	jdff dff_B_bqLpzn4O5_0(.din(w_dff_B_2pixfssf7_0),.dout(w_dff_B_bqLpzn4O5_0),.clk(gclk));
	jdff dff_B_cLRNaMk04_0(.din(w_dff_B_bqLpzn4O5_0),.dout(w_dff_B_cLRNaMk04_0),.clk(gclk));
	jdff dff_B_dWHjnBLA2_0(.din(w_dff_B_cLRNaMk04_0),.dout(w_dff_B_dWHjnBLA2_0),.clk(gclk));
	jdff dff_B_Sp28x1Ar4_0(.din(w_dff_B_dWHjnBLA2_0),.dout(w_dff_B_Sp28x1Ar4_0),.clk(gclk));
	jdff dff_B_STtDZsFd2_0(.din(w_dff_B_Sp28x1Ar4_0),.dout(w_dff_B_STtDZsFd2_0),.clk(gclk));
	jdff dff_B_k6gMftkm4_0(.din(w_dff_B_STtDZsFd2_0),.dout(w_dff_B_k6gMftkm4_0),.clk(gclk));
	jdff dff_B_v4YSt8vz1_0(.din(w_dff_B_k6gMftkm4_0),.dout(w_dff_B_v4YSt8vz1_0),.clk(gclk));
	jdff dff_B_mQg6QTo99_0(.din(w_dff_B_v4YSt8vz1_0),.dout(w_dff_B_mQg6QTo99_0),.clk(gclk));
	jdff dff_B_rAcpl1I21_0(.din(w_dff_B_mQg6QTo99_0),.dout(w_dff_B_rAcpl1I21_0),.clk(gclk));
	jdff dff_B_X8LY3C7p1_0(.din(w_dff_B_rAcpl1I21_0),.dout(w_dff_B_X8LY3C7p1_0),.clk(gclk));
	jdff dff_B_jEbGC2eA4_1(.din(n546),.dout(w_dff_B_jEbGC2eA4_1),.clk(gclk));
	jdff dff_B_N1xf8Rcn6_1(.din(w_dff_B_jEbGC2eA4_1),.dout(w_dff_B_N1xf8Rcn6_1),.clk(gclk));
	jdff dff_B_Muv2PFjB5_1(.din(w_dff_B_N1xf8Rcn6_1),.dout(w_dff_B_Muv2PFjB5_1),.clk(gclk));
	jdff dff_B_xw8Q4aK42_1(.din(w_dff_B_Muv2PFjB5_1),.dout(w_dff_B_xw8Q4aK42_1),.clk(gclk));
	jdff dff_B_p7z4SON57_1(.din(w_dff_B_xw8Q4aK42_1),.dout(w_dff_B_p7z4SON57_1),.clk(gclk));
	jdff dff_B_7jxHsP4f2_1(.din(w_dff_B_p7z4SON57_1),.dout(w_dff_B_7jxHsP4f2_1),.clk(gclk));
	jdff dff_B_ViqrtEds8_1(.din(w_dff_B_7jxHsP4f2_1),.dout(w_dff_B_ViqrtEds8_1),.clk(gclk));
	jdff dff_B_hPARAbyN5_1(.din(w_dff_B_ViqrtEds8_1),.dout(w_dff_B_hPARAbyN5_1),.clk(gclk));
	jdff dff_B_QjBjnzj84_1(.din(w_dff_B_hPARAbyN5_1),.dout(w_dff_B_QjBjnzj84_1),.clk(gclk));
	jdff dff_B_Yyp7tIBm2_1(.din(w_dff_B_QjBjnzj84_1),.dout(w_dff_B_Yyp7tIBm2_1),.clk(gclk));
	jdff dff_B_x3H8XNX06_1(.din(w_dff_B_Yyp7tIBm2_1),.dout(w_dff_B_x3H8XNX06_1),.clk(gclk));
	jdff dff_B_8EszFODT5_1(.din(w_dff_B_x3H8XNX06_1),.dout(w_dff_B_8EszFODT5_1),.clk(gclk));
	jdff dff_B_81DWx3yH1_1(.din(w_dff_B_8EszFODT5_1),.dout(w_dff_B_81DWx3yH1_1),.clk(gclk));
	jdff dff_B_DvNlnxOf2_1(.din(w_dff_B_81DWx3yH1_1),.dout(w_dff_B_DvNlnxOf2_1),.clk(gclk));
	jdff dff_B_pJ6Gmn2H1_1(.din(w_dff_B_DvNlnxOf2_1),.dout(w_dff_B_pJ6Gmn2H1_1),.clk(gclk));
	jdff dff_B_giWiqLOj7_1(.din(w_dff_B_pJ6Gmn2H1_1),.dout(w_dff_B_giWiqLOj7_1),.clk(gclk));
	jdff dff_B_UY4LD7Fn5_1(.din(w_dff_B_giWiqLOj7_1),.dout(w_dff_B_UY4LD7Fn5_1),.clk(gclk));
	jdff dff_B_Vp0VVceo5_1(.din(w_dff_B_UY4LD7Fn5_1),.dout(w_dff_B_Vp0VVceo5_1),.clk(gclk));
	jdff dff_B_0GsAUBrv1_1(.din(w_dff_B_Vp0VVceo5_1),.dout(w_dff_B_0GsAUBrv1_1),.clk(gclk));
	jdff dff_B_2QT99DA90_1(.din(w_dff_B_0GsAUBrv1_1),.dout(w_dff_B_2QT99DA90_1),.clk(gclk));
	jdff dff_B_6PQDSOM19_1(.din(w_dff_B_2QT99DA90_1),.dout(w_dff_B_6PQDSOM19_1),.clk(gclk));
	jdff dff_B_SKkqFQD85_1(.din(w_dff_B_6PQDSOM19_1),.dout(w_dff_B_SKkqFQD85_1),.clk(gclk));
	jdff dff_B_PZ5OFXo40_1(.din(w_dff_B_SKkqFQD85_1),.dout(w_dff_B_PZ5OFXo40_1),.clk(gclk));
	jdff dff_B_mcYUlvgW4_1(.din(w_dff_B_PZ5OFXo40_1),.dout(w_dff_B_mcYUlvgW4_1),.clk(gclk));
	jdff dff_B_W1aVsd749_1(.din(w_dff_B_mcYUlvgW4_1),.dout(w_dff_B_W1aVsd749_1),.clk(gclk));
	jdff dff_B_zPLs8g880_1(.din(w_dff_B_W1aVsd749_1),.dout(w_dff_B_zPLs8g880_1),.clk(gclk));
	jdff dff_B_UIEJM1lk8_1(.din(w_dff_B_zPLs8g880_1),.dout(w_dff_B_UIEJM1lk8_1),.clk(gclk));
	jdff dff_B_AWw7MNe60_0(.din(n547),.dout(w_dff_B_AWw7MNe60_0),.clk(gclk));
	jdff dff_B_kF1uaxWH8_0(.din(w_dff_B_AWw7MNe60_0),.dout(w_dff_B_kF1uaxWH8_0),.clk(gclk));
	jdff dff_B_a28HfzOT6_0(.din(w_dff_B_kF1uaxWH8_0),.dout(w_dff_B_a28HfzOT6_0),.clk(gclk));
	jdff dff_B_bUKqhQLd8_0(.din(w_dff_B_a28HfzOT6_0),.dout(w_dff_B_bUKqhQLd8_0),.clk(gclk));
	jdff dff_B_UAXnDc7f5_0(.din(w_dff_B_bUKqhQLd8_0),.dout(w_dff_B_UAXnDc7f5_0),.clk(gclk));
	jdff dff_B_EI4oPBKI2_0(.din(w_dff_B_UAXnDc7f5_0),.dout(w_dff_B_EI4oPBKI2_0),.clk(gclk));
	jdff dff_B_K9sMFS0A1_0(.din(w_dff_B_EI4oPBKI2_0),.dout(w_dff_B_K9sMFS0A1_0),.clk(gclk));
	jdff dff_B_Sg9hxv1q9_0(.din(w_dff_B_K9sMFS0A1_0),.dout(w_dff_B_Sg9hxv1q9_0),.clk(gclk));
	jdff dff_B_CMnCBKYk6_0(.din(w_dff_B_Sg9hxv1q9_0),.dout(w_dff_B_CMnCBKYk6_0),.clk(gclk));
	jdff dff_B_BbvIvvKF4_0(.din(w_dff_B_CMnCBKYk6_0),.dout(w_dff_B_BbvIvvKF4_0),.clk(gclk));
	jdff dff_B_4VpBNvBM1_0(.din(w_dff_B_BbvIvvKF4_0),.dout(w_dff_B_4VpBNvBM1_0),.clk(gclk));
	jdff dff_B_XYAcKEcw3_0(.din(w_dff_B_4VpBNvBM1_0),.dout(w_dff_B_XYAcKEcw3_0),.clk(gclk));
	jdff dff_B_K1Tmd6IG7_0(.din(w_dff_B_XYAcKEcw3_0),.dout(w_dff_B_K1Tmd6IG7_0),.clk(gclk));
	jdff dff_B_wAtzXDS95_0(.din(w_dff_B_K1Tmd6IG7_0),.dout(w_dff_B_wAtzXDS95_0),.clk(gclk));
	jdff dff_B_TNLldSDC0_0(.din(w_dff_B_wAtzXDS95_0),.dout(w_dff_B_TNLldSDC0_0),.clk(gclk));
	jdff dff_B_RWGFRdYC9_0(.din(w_dff_B_TNLldSDC0_0),.dout(w_dff_B_RWGFRdYC9_0),.clk(gclk));
	jdff dff_B_RAAQqzSZ3_0(.din(w_dff_B_RWGFRdYC9_0),.dout(w_dff_B_RAAQqzSZ3_0),.clk(gclk));
	jdff dff_B_DISV63gQ0_0(.din(w_dff_B_RAAQqzSZ3_0),.dout(w_dff_B_DISV63gQ0_0),.clk(gclk));
	jdff dff_B_DhzvxISg0_0(.din(w_dff_B_DISV63gQ0_0),.dout(w_dff_B_DhzvxISg0_0),.clk(gclk));
	jdff dff_B_sSsDZT0G4_0(.din(w_dff_B_DhzvxISg0_0),.dout(w_dff_B_sSsDZT0G4_0),.clk(gclk));
	jdff dff_B_QUxvVfjt7_0(.din(w_dff_B_sSsDZT0G4_0),.dout(w_dff_B_QUxvVfjt7_0),.clk(gclk));
	jdff dff_B_lDnu2xxq9_0(.din(w_dff_B_QUxvVfjt7_0),.dout(w_dff_B_lDnu2xxq9_0),.clk(gclk));
	jdff dff_B_CV1cKdzL0_0(.din(w_dff_B_lDnu2xxq9_0),.dout(w_dff_B_CV1cKdzL0_0),.clk(gclk));
	jdff dff_B_qhHkb7Ch0_0(.din(w_dff_B_CV1cKdzL0_0),.dout(w_dff_B_qhHkb7Ch0_0),.clk(gclk));
	jdff dff_B_euxuPu5B7_0(.din(w_dff_B_qhHkb7Ch0_0),.dout(w_dff_B_euxuPu5B7_0),.clk(gclk));
	jdff dff_B_9Xff2Fa12_0(.din(w_dff_B_euxuPu5B7_0),.dout(w_dff_B_9Xff2Fa12_0),.clk(gclk));
	jdff dff_B_d3Bc1Lmg9_0(.din(w_dff_B_9Xff2Fa12_0),.dout(w_dff_B_d3Bc1Lmg9_0),.clk(gclk));
	jdff dff_B_m47kjmmf6_1(.din(n540),.dout(w_dff_B_m47kjmmf6_1),.clk(gclk));
	jdff dff_B_zEKrbGf94_1(.din(w_dff_B_m47kjmmf6_1),.dout(w_dff_B_zEKrbGf94_1),.clk(gclk));
	jdff dff_B_H1UwU8lb9_1(.din(w_dff_B_zEKrbGf94_1),.dout(w_dff_B_H1UwU8lb9_1),.clk(gclk));
	jdff dff_B_cJefzE431_1(.din(w_dff_B_H1UwU8lb9_1),.dout(w_dff_B_cJefzE431_1),.clk(gclk));
	jdff dff_B_upxIZDjY4_1(.din(w_dff_B_cJefzE431_1),.dout(w_dff_B_upxIZDjY4_1),.clk(gclk));
	jdff dff_B_p0hMUHHl6_1(.din(w_dff_B_upxIZDjY4_1),.dout(w_dff_B_p0hMUHHl6_1),.clk(gclk));
	jdff dff_B_SD1wIlEX0_1(.din(w_dff_B_p0hMUHHl6_1),.dout(w_dff_B_SD1wIlEX0_1),.clk(gclk));
	jdff dff_B_UXLwP4lR4_1(.din(w_dff_B_SD1wIlEX0_1),.dout(w_dff_B_UXLwP4lR4_1),.clk(gclk));
	jdff dff_B_MsRu5ljh5_1(.din(w_dff_B_UXLwP4lR4_1),.dout(w_dff_B_MsRu5ljh5_1),.clk(gclk));
	jdff dff_B_aSlCRTCN1_1(.din(w_dff_B_MsRu5ljh5_1),.dout(w_dff_B_aSlCRTCN1_1),.clk(gclk));
	jdff dff_B_Yjl4ESYk8_1(.din(w_dff_B_aSlCRTCN1_1),.dout(w_dff_B_Yjl4ESYk8_1),.clk(gclk));
	jdff dff_B_jq0aeaTg8_1(.din(w_dff_B_Yjl4ESYk8_1),.dout(w_dff_B_jq0aeaTg8_1),.clk(gclk));
	jdff dff_B_mSQQUG2e5_1(.din(w_dff_B_jq0aeaTg8_1),.dout(w_dff_B_mSQQUG2e5_1),.clk(gclk));
	jdff dff_B_vmZPRSBL5_1(.din(w_dff_B_mSQQUG2e5_1),.dout(w_dff_B_vmZPRSBL5_1),.clk(gclk));
	jdff dff_B_W3oA2bFZ1_1(.din(w_dff_B_vmZPRSBL5_1),.dout(w_dff_B_W3oA2bFZ1_1),.clk(gclk));
	jdff dff_B_qhDGW6su6_1(.din(w_dff_B_W3oA2bFZ1_1),.dout(w_dff_B_qhDGW6su6_1),.clk(gclk));
	jdff dff_B_XrYy7vtE8_1(.din(w_dff_B_qhDGW6su6_1),.dout(w_dff_B_XrYy7vtE8_1),.clk(gclk));
	jdff dff_B_gTMcphaj8_1(.din(w_dff_B_XrYy7vtE8_1),.dout(w_dff_B_gTMcphaj8_1),.clk(gclk));
	jdff dff_B_LuUPDFaz9_1(.din(w_dff_B_gTMcphaj8_1),.dout(w_dff_B_LuUPDFaz9_1),.clk(gclk));
	jdff dff_B_eVAlL21p9_1(.din(w_dff_B_LuUPDFaz9_1),.dout(w_dff_B_eVAlL21p9_1),.clk(gclk));
	jdff dff_B_gGkGFiGi3_1(.din(w_dff_B_eVAlL21p9_1),.dout(w_dff_B_gGkGFiGi3_1),.clk(gclk));
	jdff dff_B_sYS25J7f9_1(.din(w_dff_B_gGkGFiGi3_1),.dout(w_dff_B_sYS25J7f9_1),.clk(gclk));
	jdff dff_B_YYnhOVjW6_1(.din(w_dff_B_sYS25J7f9_1),.dout(w_dff_B_YYnhOVjW6_1),.clk(gclk));
	jdff dff_B_qpi6SN8X2_1(.din(w_dff_B_YYnhOVjW6_1),.dout(w_dff_B_qpi6SN8X2_1),.clk(gclk));
	jdff dff_B_LQskBW503_1(.din(w_dff_B_qpi6SN8X2_1),.dout(w_dff_B_LQskBW503_1),.clk(gclk));
	jdff dff_B_YvVPAofT6_1(.din(w_dff_B_LQskBW503_1),.dout(w_dff_B_YvVPAofT6_1),.clk(gclk));
	jdff dff_B_6LkOjHvA7_0(.din(n541),.dout(w_dff_B_6LkOjHvA7_0),.clk(gclk));
	jdff dff_B_4XYmqwGw4_0(.din(w_dff_B_6LkOjHvA7_0),.dout(w_dff_B_4XYmqwGw4_0),.clk(gclk));
	jdff dff_B_iolOQF2d8_0(.din(w_dff_B_4XYmqwGw4_0),.dout(w_dff_B_iolOQF2d8_0),.clk(gclk));
	jdff dff_B_RnfMtriw1_0(.din(w_dff_B_iolOQF2d8_0),.dout(w_dff_B_RnfMtriw1_0),.clk(gclk));
	jdff dff_B_sUsicH7W0_0(.din(w_dff_B_RnfMtriw1_0),.dout(w_dff_B_sUsicH7W0_0),.clk(gclk));
	jdff dff_B_QJnco1Dq8_0(.din(w_dff_B_sUsicH7W0_0),.dout(w_dff_B_QJnco1Dq8_0),.clk(gclk));
	jdff dff_B_Hh5ikDDx5_0(.din(w_dff_B_QJnco1Dq8_0),.dout(w_dff_B_Hh5ikDDx5_0),.clk(gclk));
	jdff dff_B_IR9jkgZl4_0(.din(w_dff_B_Hh5ikDDx5_0),.dout(w_dff_B_IR9jkgZl4_0),.clk(gclk));
	jdff dff_B_scrGlXOA1_0(.din(w_dff_B_IR9jkgZl4_0),.dout(w_dff_B_scrGlXOA1_0),.clk(gclk));
	jdff dff_B_V1Yi3vbE7_0(.din(w_dff_B_scrGlXOA1_0),.dout(w_dff_B_V1Yi3vbE7_0),.clk(gclk));
	jdff dff_B_UobApmHn1_0(.din(w_dff_B_V1Yi3vbE7_0),.dout(w_dff_B_UobApmHn1_0),.clk(gclk));
	jdff dff_B_bePznbIU0_0(.din(w_dff_B_UobApmHn1_0),.dout(w_dff_B_bePznbIU0_0),.clk(gclk));
	jdff dff_B_wPzL3Mn84_0(.din(w_dff_B_bePznbIU0_0),.dout(w_dff_B_wPzL3Mn84_0),.clk(gclk));
	jdff dff_B_5s9X372m0_0(.din(w_dff_B_wPzL3Mn84_0),.dout(w_dff_B_5s9X372m0_0),.clk(gclk));
	jdff dff_B_g9XD0cEj8_0(.din(w_dff_B_5s9X372m0_0),.dout(w_dff_B_g9XD0cEj8_0),.clk(gclk));
	jdff dff_B_DRy4QOlE3_0(.din(w_dff_B_g9XD0cEj8_0),.dout(w_dff_B_DRy4QOlE3_0),.clk(gclk));
	jdff dff_B_p395qPK33_0(.din(w_dff_B_DRy4QOlE3_0),.dout(w_dff_B_p395qPK33_0),.clk(gclk));
	jdff dff_B_H9PsgRw26_0(.din(w_dff_B_p395qPK33_0),.dout(w_dff_B_H9PsgRw26_0),.clk(gclk));
	jdff dff_B_pXTfVs3i5_0(.din(w_dff_B_H9PsgRw26_0),.dout(w_dff_B_pXTfVs3i5_0),.clk(gclk));
	jdff dff_B_H3VVbSMP6_0(.din(w_dff_B_pXTfVs3i5_0),.dout(w_dff_B_H3VVbSMP6_0),.clk(gclk));
	jdff dff_B_FvACIz0R3_0(.din(w_dff_B_H3VVbSMP6_0),.dout(w_dff_B_FvACIz0R3_0),.clk(gclk));
	jdff dff_B_3u3wk3C94_0(.din(w_dff_B_FvACIz0R3_0),.dout(w_dff_B_3u3wk3C94_0),.clk(gclk));
	jdff dff_B_g8Cm3rJN0_0(.din(w_dff_B_3u3wk3C94_0),.dout(w_dff_B_g8Cm3rJN0_0),.clk(gclk));
	jdff dff_B_HIycXObK2_0(.din(w_dff_B_g8Cm3rJN0_0),.dout(w_dff_B_HIycXObK2_0),.clk(gclk));
	jdff dff_B_CT7QS0sv9_0(.din(w_dff_B_HIycXObK2_0),.dout(w_dff_B_CT7QS0sv9_0),.clk(gclk));
	jdff dff_B_bFwFmeEw7_0(.din(w_dff_B_CT7QS0sv9_0),.dout(w_dff_B_bFwFmeEw7_0),.clk(gclk));
	jdff dff_B_Wb0mxUq91_1(.din(n534),.dout(w_dff_B_Wb0mxUq91_1),.clk(gclk));
	jdff dff_B_WiO3QQhK2_1(.din(w_dff_B_Wb0mxUq91_1),.dout(w_dff_B_WiO3QQhK2_1),.clk(gclk));
	jdff dff_B_GYWvVFsF0_1(.din(w_dff_B_WiO3QQhK2_1),.dout(w_dff_B_GYWvVFsF0_1),.clk(gclk));
	jdff dff_B_qhkzfFXX1_1(.din(w_dff_B_GYWvVFsF0_1),.dout(w_dff_B_qhkzfFXX1_1),.clk(gclk));
	jdff dff_B_nylJwnYH2_1(.din(w_dff_B_qhkzfFXX1_1),.dout(w_dff_B_nylJwnYH2_1),.clk(gclk));
	jdff dff_B_pdQynfY53_1(.din(w_dff_B_nylJwnYH2_1),.dout(w_dff_B_pdQynfY53_1),.clk(gclk));
	jdff dff_B_FbVuU11Y5_1(.din(w_dff_B_pdQynfY53_1),.dout(w_dff_B_FbVuU11Y5_1),.clk(gclk));
	jdff dff_B_uEDEhPiX2_1(.din(w_dff_B_FbVuU11Y5_1),.dout(w_dff_B_uEDEhPiX2_1),.clk(gclk));
	jdff dff_B_VGYtJ86v7_1(.din(w_dff_B_uEDEhPiX2_1),.dout(w_dff_B_VGYtJ86v7_1),.clk(gclk));
	jdff dff_B_2QwbOco99_1(.din(w_dff_B_VGYtJ86v7_1),.dout(w_dff_B_2QwbOco99_1),.clk(gclk));
	jdff dff_B_B9VzruyW8_1(.din(w_dff_B_2QwbOco99_1),.dout(w_dff_B_B9VzruyW8_1),.clk(gclk));
	jdff dff_B_5l5KD6jS0_1(.din(w_dff_B_B9VzruyW8_1),.dout(w_dff_B_5l5KD6jS0_1),.clk(gclk));
	jdff dff_B_uhAMMFSz4_1(.din(w_dff_B_5l5KD6jS0_1),.dout(w_dff_B_uhAMMFSz4_1),.clk(gclk));
	jdff dff_B_WJ0QK7hy6_1(.din(w_dff_B_uhAMMFSz4_1),.dout(w_dff_B_WJ0QK7hy6_1),.clk(gclk));
	jdff dff_B_1URQWq077_1(.din(w_dff_B_WJ0QK7hy6_1),.dout(w_dff_B_1URQWq077_1),.clk(gclk));
	jdff dff_B_GTxav8wm7_1(.din(w_dff_B_1URQWq077_1),.dout(w_dff_B_GTxav8wm7_1),.clk(gclk));
	jdff dff_B_WDFwtscJ7_1(.din(w_dff_B_GTxav8wm7_1),.dout(w_dff_B_WDFwtscJ7_1),.clk(gclk));
	jdff dff_B_8qsrFrGL2_1(.din(w_dff_B_WDFwtscJ7_1),.dout(w_dff_B_8qsrFrGL2_1),.clk(gclk));
	jdff dff_B_Zm5x2N2B7_1(.din(w_dff_B_8qsrFrGL2_1),.dout(w_dff_B_Zm5x2N2B7_1),.clk(gclk));
	jdff dff_B_0pT00Q9e4_1(.din(w_dff_B_Zm5x2N2B7_1),.dout(w_dff_B_0pT00Q9e4_1),.clk(gclk));
	jdff dff_B_RzrTjCVQ8_1(.din(w_dff_B_0pT00Q9e4_1),.dout(w_dff_B_RzrTjCVQ8_1),.clk(gclk));
	jdff dff_B_QElwnxde8_1(.din(w_dff_B_RzrTjCVQ8_1),.dout(w_dff_B_QElwnxde8_1),.clk(gclk));
	jdff dff_B_fdLvrelX7_1(.din(w_dff_B_QElwnxde8_1),.dout(w_dff_B_fdLvrelX7_1),.clk(gclk));
	jdff dff_B_Gzqg4BA45_1(.din(w_dff_B_fdLvrelX7_1),.dout(w_dff_B_Gzqg4BA45_1),.clk(gclk));
	jdff dff_B_nk8Q4hzv5_1(.din(w_dff_B_Gzqg4BA45_1),.dout(w_dff_B_nk8Q4hzv5_1),.clk(gclk));
	jdff dff_B_db5T3eSR1_0(.din(n535),.dout(w_dff_B_db5T3eSR1_0),.clk(gclk));
	jdff dff_B_AYPQc4Vq2_0(.din(w_dff_B_db5T3eSR1_0),.dout(w_dff_B_AYPQc4Vq2_0),.clk(gclk));
	jdff dff_B_jHtMmMs17_0(.din(w_dff_B_AYPQc4Vq2_0),.dout(w_dff_B_jHtMmMs17_0),.clk(gclk));
	jdff dff_B_UHjYbtox8_0(.din(w_dff_B_jHtMmMs17_0),.dout(w_dff_B_UHjYbtox8_0),.clk(gclk));
	jdff dff_B_sYdTR8HW9_0(.din(w_dff_B_UHjYbtox8_0),.dout(w_dff_B_sYdTR8HW9_0),.clk(gclk));
	jdff dff_B_QPRMV83g6_0(.din(w_dff_B_sYdTR8HW9_0),.dout(w_dff_B_QPRMV83g6_0),.clk(gclk));
	jdff dff_B_TY2eUKX81_0(.din(w_dff_B_QPRMV83g6_0),.dout(w_dff_B_TY2eUKX81_0),.clk(gclk));
	jdff dff_B_duOTAfbj6_0(.din(w_dff_B_TY2eUKX81_0),.dout(w_dff_B_duOTAfbj6_0),.clk(gclk));
	jdff dff_B_0LrOqCnH6_0(.din(w_dff_B_duOTAfbj6_0),.dout(w_dff_B_0LrOqCnH6_0),.clk(gclk));
	jdff dff_B_G6daYLZo1_0(.din(w_dff_B_0LrOqCnH6_0),.dout(w_dff_B_G6daYLZo1_0),.clk(gclk));
	jdff dff_B_WT7QBB8j8_0(.din(w_dff_B_G6daYLZo1_0),.dout(w_dff_B_WT7QBB8j8_0),.clk(gclk));
	jdff dff_B_UXiN6msR9_0(.din(w_dff_B_WT7QBB8j8_0),.dout(w_dff_B_UXiN6msR9_0),.clk(gclk));
	jdff dff_B_z0k8JdLs2_0(.din(w_dff_B_UXiN6msR9_0),.dout(w_dff_B_z0k8JdLs2_0),.clk(gclk));
	jdff dff_B_tvfgLy9T5_0(.din(w_dff_B_z0k8JdLs2_0),.dout(w_dff_B_tvfgLy9T5_0),.clk(gclk));
	jdff dff_B_YBtL3Jbo1_0(.din(w_dff_B_tvfgLy9T5_0),.dout(w_dff_B_YBtL3Jbo1_0),.clk(gclk));
	jdff dff_B_xjmg3mpv1_0(.din(w_dff_B_YBtL3Jbo1_0),.dout(w_dff_B_xjmg3mpv1_0),.clk(gclk));
	jdff dff_B_vDtxa8cd9_0(.din(w_dff_B_xjmg3mpv1_0),.dout(w_dff_B_vDtxa8cd9_0),.clk(gclk));
	jdff dff_B_4e90aYLG8_0(.din(w_dff_B_vDtxa8cd9_0),.dout(w_dff_B_4e90aYLG8_0),.clk(gclk));
	jdff dff_B_i3Jja0yv6_0(.din(w_dff_B_4e90aYLG8_0),.dout(w_dff_B_i3Jja0yv6_0),.clk(gclk));
	jdff dff_B_HQalQ15v3_0(.din(w_dff_B_i3Jja0yv6_0),.dout(w_dff_B_HQalQ15v3_0),.clk(gclk));
	jdff dff_B_Q8dyLceV7_0(.din(w_dff_B_HQalQ15v3_0),.dout(w_dff_B_Q8dyLceV7_0),.clk(gclk));
	jdff dff_B_rBGac74U7_0(.din(w_dff_B_Q8dyLceV7_0),.dout(w_dff_B_rBGac74U7_0),.clk(gclk));
	jdff dff_B_f359shWt5_0(.din(w_dff_B_rBGac74U7_0),.dout(w_dff_B_f359shWt5_0),.clk(gclk));
	jdff dff_B_VuXxQXSH5_0(.din(w_dff_B_f359shWt5_0),.dout(w_dff_B_VuXxQXSH5_0),.clk(gclk));
	jdff dff_B_kc8HMq882_0(.din(w_dff_B_VuXxQXSH5_0),.dout(w_dff_B_kc8HMq882_0),.clk(gclk));
	jdff dff_B_AnRFY6P59_1(.din(n528),.dout(w_dff_B_AnRFY6P59_1),.clk(gclk));
	jdff dff_B_1ilWoncE7_1(.din(w_dff_B_AnRFY6P59_1),.dout(w_dff_B_1ilWoncE7_1),.clk(gclk));
	jdff dff_B_TtVvSwnO9_1(.din(w_dff_B_1ilWoncE7_1),.dout(w_dff_B_TtVvSwnO9_1),.clk(gclk));
	jdff dff_B_2e2GW7yY0_1(.din(w_dff_B_TtVvSwnO9_1),.dout(w_dff_B_2e2GW7yY0_1),.clk(gclk));
	jdff dff_B_XfbvT7Nc6_1(.din(w_dff_B_2e2GW7yY0_1),.dout(w_dff_B_XfbvT7Nc6_1),.clk(gclk));
	jdff dff_B_ahL5U5e97_1(.din(w_dff_B_XfbvT7Nc6_1),.dout(w_dff_B_ahL5U5e97_1),.clk(gclk));
	jdff dff_B_8pAs6gXb9_1(.din(w_dff_B_ahL5U5e97_1),.dout(w_dff_B_8pAs6gXb9_1),.clk(gclk));
	jdff dff_B_pzbWGiv33_1(.din(w_dff_B_8pAs6gXb9_1),.dout(w_dff_B_pzbWGiv33_1),.clk(gclk));
	jdff dff_B_zmTmNv9A8_1(.din(w_dff_B_pzbWGiv33_1),.dout(w_dff_B_zmTmNv9A8_1),.clk(gclk));
	jdff dff_B_SFd7vEGX0_1(.din(w_dff_B_zmTmNv9A8_1),.dout(w_dff_B_SFd7vEGX0_1),.clk(gclk));
	jdff dff_B_mPM0y6mF0_1(.din(w_dff_B_SFd7vEGX0_1),.dout(w_dff_B_mPM0y6mF0_1),.clk(gclk));
	jdff dff_B_Fg9q1f5W4_1(.din(w_dff_B_mPM0y6mF0_1),.dout(w_dff_B_Fg9q1f5W4_1),.clk(gclk));
	jdff dff_B_hby8E9yb4_1(.din(w_dff_B_Fg9q1f5W4_1),.dout(w_dff_B_hby8E9yb4_1),.clk(gclk));
	jdff dff_B_KO7H60of7_1(.din(w_dff_B_hby8E9yb4_1),.dout(w_dff_B_KO7H60of7_1),.clk(gclk));
	jdff dff_B_esIAVLEp6_1(.din(w_dff_B_KO7H60of7_1),.dout(w_dff_B_esIAVLEp6_1),.clk(gclk));
	jdff dff_B_NmX60Cay4_1(.din(w_dff_B_esIAVLEp6_1),.dout(w_dff_B_NmX60Cay4_1),.clk(gclk));
	jdff dff_B_VSgvxO1I9_1(.din(w_dff_B_NmX60Cay4_1),.dout(w_dff_B_VSgvxO1I9_1),.clk(gclk));
	jdff dff_B_XhQg9Mxx1_1(.din(w_dff_B_VSgvxO1I9_1),.dout(w_dff_B_XhQg9Mxx1_1),.clk(gclk));
	jdff dff_B_qHdW0Lby3_1(.din(w_dff_B_XhQg9Mxx1_1),.dout(w_dff_B_qHdW0Lby3_1),.clk(gclk));
	jdff dff_B_0rJbQZPN9_1(.din(w_dff_B_qHdW0Lby3_1),.dout(w_dff_B_0rJbQZPN9_1),.clk(gclk));
	jdff dff_B_UqtMZYYs4_1(.din(w_dff_B_0rJbQZPN9_1),.dout(w_dff_B_UqtMZYYs4_1),.clk(gclk));
	jdff dff_B_2STSG4oh5_1(.din(w_dff_B_UqtMZYYs4_1),.dout(w_dff_B_2STSG4oh5_1),.clk(gclk));
	jdff dff_B_FXFRtHln0_1(.din(w_dff_B_2STSG4oh5_1),.dout(w_dff_B_FXFRtHln0_1),.clk(gclk));
	jdff dff_B_mAYLtnxH0_1(.din(w_dff_B_FXFRtHln0_1),.dout(w_dff_B_mAYLtnxH0_1),.clk(gclk));
	jdff dff_B_ORB5OVYO5_0(.din(n529),.dout(w_dff_B_ORB5OVYO5_0),.clk(gclk));
	jdff dff_B_dsD3knkv5_0(.din(w_dff_B_ORB5OVYO5_0),.dout(w_dff_B_dsD3knkv5_0),.clk(gclk));
	jdff dff_B_rBiIlAy80_0(.din(w_dff_B_dsD3knkv5_0),.dout(w_dff_B_rBiIlAy80_0),.clk(gclk));
	jdff dff_B_0wGjaba27_0(.din(w_dff_B_rBiIlAy80_0),.dout(w_dff_B_0wGjaba27_0),.clk(gclk));
	jdff dff_B_RgCIjfmT8_0(.din(w_dff_B_0wGjaba27_0),.dout(w_dff_B_RgCIjfmT8_0),.clk(gclk));
	jdff dff_B_BQDcfmLy4_0(.din(w_dff_B_RgCIjfmT8_0),.dout(w_dff_B_BQDcfmLy4_0),.clk(gclk));
	jdff dff_B_xUWZgGL89_0(.din(w_dff_B_BQDcfmLy4_0),.dout(w_dff_B_xUWZgGL89_0),.clk(gclk));
	jdff dff_B_hsB7URDw7_0(.din(w_dff_B_xUWZgGL89_0),.dout(w_dff_B_hsB7URDw7_0),.clk(gclk));
	jdff dff_B_phT04UDP8_0(.din(w_dff_B_hsB7URDw7_0),.dout(w_dff_B_phT04UDP8_0),.clk(gclk));
	jdff dff_B_FQMjJqiN4_0(.din(w_dff_B_phT04UDP8_0),.dout(w_dff_B_FQMjJqiN4_0),.clk(gclk));
	jdff dff_B_C64ubjqN9_0(.din(w_dff_B_FQMjJqiN4_0),.dout(w_dff_B_C64ubjqN9_0),.clk(gclk));
	jdff dff_B_EUN409DQ7_0(.din(w_dff_B_C64ubjqN9_0),.dout(w_dff_B_EUN409DQ7_0),.clk(gclk));
	jdff dff_B_2dXi4wSe8_0(.din(w_dff_B_EUN409DQ7_0),.dout(w_dff_B_2dXi4wSe8_0),.clk(gclk));
	jdff dff_B_JCRcWhEw7_0(.din(w_dff_B_2dXi4wSe8_0),.dout(w_dff_B_JCRcWhEw7_0),.clk(gclk));
	jdff dff_B_3HENdVeT2_0(.din(w_dff_B_JCRcWhEw7_0),.dout(w_dff_B_3HENdVeT2_0),.clk(gclk));
	jdff dff_B_lutsWKzk8_0(.din(w_dff_B_3HENdVeT2_0),.dout(w_dff_B_lutsWKzk8_0),.clk(gclk));
	jdff dff_B_iXN2t8V27_0(.din(w_dff_B_lutsWKzk8_0),.dout(w_dff_B_iXN2t8V27_0),.clk(gclk));
	jdff dff_B_uft6ISGb8_0(.din(w_dff_B_iXN2t8V27_0),.dout(w_dff_B_uft6ISGb8_0),.clk(gclk));
	jdff dff_B_qNlsMg7G1_0(.din(w_dff_B_uft6ISGb8_0),.dout(w_dff_B_qNlsMg7G1_0),.clk(gclk));
	jdff dff_B_2PO0njAe1_0(.din(w_dff_B_qNlsMg7G1_0),.dout(w_dff_B_2PO0njAe1_0),.clk(gclk));
	jdff dff_B_PsqNBR7s9_0(.din(w_dff_B_2PO0njAe1_0),.dout(w_dff_B_PsqNBR7s9_0),.clk(gclk));
	jdff dff_B_7Ptke34g1_0(.din(w_dff_B_PsqNBR7s9_0),.dout(w_dff_B_7Ptke34g1_0),.clk(gclk));
	jdff dff_B_duuzWikO5_0(.din(w_dff_B_7Ptke34g1_0),.dout(w_dff_B_duuzWikO5_0),.clk(gclk));
	jdff dff_B_WEHr8swc1_0(.din(w_dff_B_duuzWikO5_0),.dout(w_dff_B_WEHr8swc1_0),.clk(gclk));
	jdff dff_B_7edgnBR81_1(.din(n522),.dout(w_dff_B_7edgnBR81_1),.clk(gclk));
	jdff dff_B_0MAQMHq53_1(.din(w_dff_B_7edgnBR81_1),.dout(w_dff_B_0MAQMHq53_1),.clk(gclk));
	jdff dff_B_QQdnpqgp6_1(.din(w_dff_B_0MAQMHq53_1),.dout(w_dff_B_QQdnpqgp6_1),.clk(gclk));
	jdff dff_B_piijkjuC6_1(.din(w_dff_B_QQdnpqgp6_1),.dout(w_dff_B_piijkjuC6_1),.clk(gclk));
	jdff dff_B_EqSLs5iI7_1(.din(w_dff_B_piijkjuC6_1),.dout(w_dff_B_EqSLs5iI7_1),.clk(gclk));
	jdff dff_B_3AwOmlqM8_1(.din(w_dff_B_EqSLs5iI7_1),.dout(w_dff_B_3AwOmlqM8_1),.clk(gclk));
	jdff dff_B_AGCKqSXE6_1(.din(w_dff_B_3AwOmlqM8_1),.dout(w_dff_B_AGCKqSXE6_1),.clk(gclk));
	jdff dff_B_flH8TDKj3_1(.din(w_dff_B_AGCKqSXE6_1),.dout(w_dff_B_flH8TDKj3_1),.clk(gclk));
	jdff dff_B_HR7UytV38_1(.din(w_dff_B_flH8TDKj3_1),.dout(w_dff_B_HR7UytV38_1),.clk(gclk));
	jdff dff_B_39c2frOG5_1(.din(w_dff_B_HR7UytV38_1),.dout(w_dff_B_39c2frOG5_1),.clk(gclk));
	jdff dff_B_CiMxmFWS0_1(.din(w_dff_B_39c2frOG5_1),.dout(w_dff_B_CiMxmFWS0_1),.clk(gclk));
	jdff dff_B_Duad9wHL9_1(.din(w_dff_B_CiMxmFWS0_1),.dout(w_dff_B_Duad9wHL9_1),.clk(gclk));
	jdff dff_B_mUQ0sMOW8_1(.din(w_dff_B_Duad9wHL9_1),.dout(w_dff_B_mUQ0sMOW8_1),.clk(gclk));
	jdff dff_B_xH0H4AfA9_1(.din(w_dff_B_mUQ0sMOW8_1),.dout(w_dff_B_xH0H4AfA9_1),.clk(gclk));
	jdff dff_B_MBpaSc8S3_1(.din(w_dff_B_xH0H4AfA9_1),.dout(w_dff_B_MBpaSc8S3_1),.clk(gclk));
	jdff dff_B_9VgXWMOX3_1(.din(w_dff_B_MBpaSc8S3_1),.dout(w_dff_B_9VgXWMOX3_1),.clk(gclk));
	jdff dff_B_rMCj5kZg9_1(.din(w_dff_B_9VgXWMOX3_1),.dout(w_dff_B_rMCj5kZg9_1),.clk(gclk));
	jdff dff_B_LEkqTHx12_1(.din(w_dff_B_rMCj5kZg9_1),.dout(w_dff_B_LEkqTHx12_1),.clk(gclk));
	jdff dff_B_8gaKvIj29_1(.din(w_dff_B_LEkqTHx12_1),.dout(w_dff_B_8gaKvIj29_1),.clk(gclk));
	jdff dff_B_IPopdG0o3_1(.din(w_dff_B_8gaKvIj29_1),.dout(w_dff_B_IPopdG0o3_1),.clk(gclk));
	jdff dff_B_CdY3vwIN9_1(.din(w_dff_B_IPopdG0o3_1),.dout(w_dff_B_CdY3vwIN9_1),.clk(gclk));
	jdff dff_B_QYAa0j5h3_1(.din(w_dff_B_CdY3vwIN9_1),.dout(w_dff_B_QYAa0j5h3_1),.clk(gclk));
	jdff dff_B_fxvTyWRy8_1(.din(w_dff_B_QYAa0j5h3_1),.dout(w_dff_B_fxvTyWRy8_1),.clk(gclk));
	jdff dff_B_VxcVUf7H5_0(.din(n523),.dout(w_dff_B_VxcVUf7H5_0),.clk(gclk));
	jdff dff_B_BJxiAccS9_0(.din(w_dff_B_VxcVUf7H5_0),.dout(w_dff_B_BJxiAccS9_0),.clk(gclk));
	jdff dff_B_vh1CGSU90_0(.din(w_dff_B_BJxiAccS9_0),.dout(w_dff_B_vh1CGSU90_0),.clk(gclk));
	jdff dff_B_qhTbMA485_0(.din(w_dff_B_vh1CGSU90_0),.dout(w_dff_B_qhTbMA485_0),.clk(gclk));
	jdff dff_B_gH3C0luF2_0(.din(w_dff_B_qhTbMA485_0),.dout(w_dff_B_gH3C0luF2_0),.clk(gclk));
	jdff dff_B_O6BkGu1Z7_0(.din(w_dff_B_gH3C0luF2_0),.dout(w_dff_B_O6BkGu1Z7_0),.clk(gclk));
	jdff dff_B_ubtcXv1d0_0(.din(w_dff_B_O6BkGu1Z7_0),.dout(w_dff_B_ubtcXv1d0_0),.clk(gclk));
	jdff dff_B_huwtojip9_0(.din(w_dff_B_ubtcXv1d0_0),.dout(w_dff_B_huwtojip9_0),.clk(gclk));
	jdff dff_B_wNLgOwHR6_0(.din(w_dff_B_huwtojip9_0),.dout(w_dff_B_wNLgOwHR6_0),.clk(gclk));
	jdff dff_B_yboVqc1q9_0(.din(w_dff_B_wNLgOwHR6_0),.dout(w_dff_B_yboVqc1q9_0),.clk(gclk));
	jdff dff_B_UTxHv5kQ9_0(.din(w_dff_B_yboVqc1q9_0),.dout(w_dff_B_UTxHv5kQ9_0),.clk(gclk));
	jdff dff_B_WGzj0TcJ3_0(.din(w_dff_B_UTxHv5kQ9_0),.dout(w_dff_B_WGzj0TcJ3_0),.clk(gclk));
	jdff dff_B_Io800KAz5_0(.din(w_dff_B_WGzj0TcJ3_0),.dout(w_dff_B_Io800KAz5_0),.clk(gclk));
	jdff dff_B_cjg6KSmO8_0(.din(w_dff_B_Io800KAz5_0),.dout(w_dff_B_cjg6KSmO8_0),.clk(gclk));
	jdff dff_B_nH0wW2JQ2_0(.din(w_dff_B_cjg6KSmO8_0),.dout(w_dff_B_nH0wW2JQ2_0),.clk(gclk));
	jdff dff_B_CGyoJYNY3_0(.din(w_dff_B_nH0wW2JQ2_0),.dout(w_dff_B_CGyoJYNY3_0),.clk(gclk));
	jdff dff_B_CjT98AnT2_0(.din(w_dff_B_CGyoJYNY3_0),.dout(w_dff_B_CjT98AnT2_0),.clk(gclk));
	jdff dff_B_NFjf6lvI5_0(.din(w_dff_B_CjT98AnT2_0),.dout(w_dff_B_NFjf6lvI5_0),.clk(gclk));
	jdff dff_B_mKaBape88_0(.din(w_dff_B_NFjf6lvI5_0),.dout(w_dff_B_mKaBape88_0),.clk(gclk));
	jdff dff_B_IG5BdfI66_0(.din(w_dff_B_mKaBape88_0),.dout(w_dff_B_IG5BdfI66_0),.clk(gclk));
	jdff dff_B_iCQC6N7R7_0(.din(w_dff_B_IG5BdfI66_0),.dout(w_dff_B_iCQC6N7R7_0),.clk(gclk));
	jdff dff_B_YCCdy70h4_0(.din(w_dff_B_iCQC6N7R7_0),.dout(w_dff_B_YCCdy70h4_0),.clk(gclk));
	jdff dff_B_vffmUHZP1_0(.din(w_dff_B_YCCdy70h4_0),.dout(w_dff_B_vffmUHZP1_0),.clk(gclk));
	jdff dff_B_DXhPNNpz1_1(.din(n516),.dout(w_dff_B_DXhPNNpz1_1),.clk(gclk));
	jdff dff_B_mTtX9v0t9_1(.din(w_dff_B_DXhPNNpz1_1),.dout(w_dff_B_mTtX9v0t9_1),.clk(gclk));
	jdff dff_B_Y2ANFewa3_1(.din(w_dff_B_mTtX9v0t9_1),.dout(w_dff_B_Y2ANFewa3_1),.clk(gclk));
	jdff dff_B_jgzopvEA0_1(.din(w_dff_B_Y2ANFewa3_1),.dout(w_dff_B_jgzopvEA0_1),.clk(gclk));
	jdff dff_B_Aq5Ikao38_1(.din(w_dff_B_jgzopvEA0_1),.dout(w_dff_B_Aq5Ikao38_1),.clk(gclk));
	jdff dff_B_UhfBFeYt6_1(.din(w_dff_B_Aq5Ikao38_1),.dout(w_dff_B_UhfBFeYt6_1),.clk(gclk));
	jdff dff_B_fHb0j4ew5_1(.din(w_dff_B_UhfBFeYt6_1),.dout(w_dff_B_fHb0j4ew5_1),.clk(gclk));
	jdff dff_B_hEoaFcUm6_1(.din(w_dff_B_fHb0j4ew5_1),.dout(w_dff_B_hEoaFcUm6_1),.clk(gclk));
	jdff dff_B_6JB7cQ9z3_1(.din(w_dff_B_hEoaFcUm6_1),.dout(w_dff_B_6JB7cQ9z3_1),.clk(gclk));
	jdff dff_B_jpBio3oi6_1(.din(w_dff_B_6JB7cQ9z3_1),.dout(w_dff_B_jpBio3oi6_1),.clk(gclk));
	jdff dff_B_cS71ko3Z0_1(.din(w_dff_B_jpBio3oi6_1),.dout(w_dff_B_cS71ko3Z0_1),.clk(gclk));
	jdff dff_B_tP12ks5X0_1(.din(w_dff_B_cS71ko3Z0_1),.dout(w_dff_B_tP12ks5X0_1),.clk(gclk));
	jdff dff_B_P0wl6mZ51_1(.din(w_dff_B_tP12ks5X0_1),.dout(w_dff_B_P0wl6mZ51_1),.clk(gclk));
	jdff dff_B_BeJoeIXj7_1(.din(w_dff_B_P0wl6mZ51_1),.dout(w_dff_B_BeJoeIXj7_1),.clk(gclk));
	jdff dff_B_79b0qMv45_1(.din(w_dff_B_BeJoeIXj7_1),.dout(w_dff_B_79b0qMv45_1),.clk(gclk));
	jdff dff_B_vnx7SaAd2_1(.din(w_dff_B_79b0qMv45_1),.dout(w_dff_B_vnx7SaAd2_1),.clk(gclk));
	jdff dff_B_Lk6oOYTe4_1(.din(w_dff_B_vnx7SaAd2_1),.dout(w_dff_B_Lk6oOYTe4_1),.clk(gclk));
	jdff dff_B_mL0PLyNd4_1(.din(w_dff_B_Lk6oOYTe4_1),.dout(w_dff_B_mL0PLyNd4_1),.clk(gclk));
	jdff dff_B_wFhZGdBy9_1(.din(w_dff_B_mL0PLyNd4_1),.dout(w_dff_B_wFhZGdBy9_1),.clk(gclk));
	jdff dff_B_O0Gb9j260_1(.din(w_dff_B_wFhZGdBy9_1),.dout(w_dff_B_O0Gb9j260_1),.clk(gclk));
	jdff dff_B_BMUS3aHp6_1(.din(w_dff_B_O0Gb9j260_1),.dout(w_dff_B_BMUS3aHp6_1),.clk(gclk));
	jdff dff_B_tOY8ECp76_1(.din(w_dff_B_BMUS3aHp6_1),.dout(w_dff_B_tOY8ECp76_1),.clk(gclk));
	jdff dff_B_GwfYFLQG5_0(.din(n517),.dout(w_dff_B_GwfYFLQG5_0),.clk(gclk));
	jdff dff_B_CS57lDA07_0(.din(w_dff_B_GwfYFLQG5_0),.dout(w_dff_B_CS57lDA07_0),.clk(gclk));
	jdff dff_B_By5F7GgY5_0(.din(w_dff_B_CS57lDA07_0),.dout(w_dff_B_By5F7GgY5_0),.clk(gclk));
	jdff dff_B_RtcdwQQd6_0(.din(w_dff_B_By5F7GgY5_0),.dout(w_dff_B_RtcdwQQd6_0),.clk(gclk));
	jdff dff_B_7Do5rFZp5_0(.din(w_dff_B_RtcdwQQd6_0),.dout(w_dff_B_7Do5rFZp5_0),.clk(gclk));
	jdff dff_B_WOqwXhkh7_0(.din(w_dff_B_7Do5rFZp5_0),.dout(w_dff_B_WOqwXhkh7_0),.clk(gclk));
	jdff dff_B_IxbFk8cI6_0(.din(w_dff_B_WOqwXhkh7_0),.dout(w_dff_B_IxbFk8cI6_0),.clk(gclk));
	jdff dff_B_0bOUT9uw7_0(.din(w_dff_B_IxbFk8cI6_0),.dout(w_dff_B_0bOUT9uw7_0),.clk(gclk));
	jdff dff_B_kwMH0CsE1_0(.din(w_dff_B_0bOUT9uw7_0),.dout(w_dff_B_kwMH0CsE1_0),.clk(gclk));
	jdff dff_B_jOj3r1vQ2_0(.din(w_dff_B_kwMH0CsE1_0),.dout(w_dff_B_jOj3r1vQ2_0),.clk(gclk));
	jdff dff_B_sfI0GuZh1_0(.din(w_dff_B_jOj3r1vQ2_0),.dout(w_dff_B_sfI0GuZh1_0),.clk(gclk));
	jdff dff_B_haoZ0fGm4_0(.din(w_dff_B_sfI0GuZh1_0),.dout(w_dff_B_haoZ0fGm4_0),.clk(gclk));
	jdff dff_B_QDtWVFUm6_0(.din(w_dff_B_haoZ0fGm4_0),.dout(w_dff_B_QDtWVFUm6_0),.clk(gclk));
	jdff dff_B_VSll0QuP2_0(.din(w_dff_B_QDtWVFUm6_0),.dout(w_dff_B_VSll0QuP2_0),.clk(gclk));
	jdff dff_B_s0KFDVXq0_0(.din(w_dff_B_VSll0QuP2_0),.dout(w_dff_B_s0KFDVXq0_0),.clk(gclk));
	jdff dff_B_lPBRUhZt3_0(.din(w_dff_B_s0KFDVXq0_0),.dout(w_dff_B_lPBRUhZt3_0),.clk(gclk));
	jdff dff_B_T52oUi9m8_0(.din(w_dff_B_lPBRUhZt3_0),.dout(w_dff_B_T52oUi9m8_0),.clk(gclk));
	jdff dff_B_QIfhqqZY6_0(.din(w_dff_B_T52oUi9m8_0),.dout(w_dff_B_QIfhqqZY6_0),.clk(gclk));
	jdff dff_B_h1TRqlBE7_0(.din(w_dff_B_QIfhqqZY6_0),.dout(w_dff_B_h1TRqlBE7_0),.clk(gclk));
	jdff dff_B_xxmYYP6a8_0(.din(w_dff_B_h1TRqlBE7_0),.dout(w_dff_B_xxmYYP6a8_0),.clk(gclk));
	jdff dff_B_y6CzhVen1_0(.din(w_dff_B_xxmYYP6a8_0),.dout(w_dff_B_y6CzhVen1_0),.clk(gclk));
	jdff dff_B_nKZIowO61_0(.din(w_dff_B_y6CzhVen1_0),.dout(w_dff_B_nKZIowO61_0),.clk(gclk));
	jdff dff_B_cnQQSUWE9_1(.din(n510),.dout(w_dff_B_cnQQSUWE9_1),.clk(gclk));
	jdff dff_B_oUTwsU4C2_1(.din(w_dff_B_cnQQSUWE9_1),.dout(w_dff_B_oUTwsU4C2_1),.clk(gclk));
	jdff dff_B_zlOAONAj5_1(.din(w_dff_B_oUTwsU4C2_1),.dout(w_dff_B_zlOAONAj5_1),.clk(gclk));
	jdff dff_B_IFtzdkkf5_1(.din(w_dff_B_zlOAONAj5_1),.dout(w_dff_B_IFtzdkkf5_1),.clk(gclk));
	jdff dff_B_Nu8LDJL90_1(.din(w_dff_B_IFtzdkkf5_1),.dout(w_dff_B_Nu8LDJL90_1),.clk(gclk));
	jdff dff_B_FvjXZquD1_1(.din(w_dff_B_Nu8LDJL90_1),.dout(w_dff_B_FvjXZquD1_1),.clk(gclk));
	jdff dff_B_FK3KUyQ09_1(.din(w_dff_B_FvjXZquD1_1),.dout(w_dff_B_FK3KUyQ09_1),.clk(gclk));
	jdff dff_B_ogbSYZp63_1(.din(w_dff_B_FK3KUyQ09_1),.dout(w_dff_B_ogbSYZp63_1),.clk(gclk));
	jdff dff_B_lR3wgXjs6_1(.din(w_dff_B_ogbSYZp63_1),.dout(w_dff_B_lR3wgXjs6_1),.clk(gclk));
	jdff dff_B_rnEWP2BY7_1(.din(w_dff_B_lR3wgXjs6_1),.dout(w_dff_B_rnEWP2BY7_1),.clk(gclk));
	jdff dff_B_nl7gEe5Z0_1(.din(w_dff_B_rnEWP2BY7_1),.dout(w_dff_B_nl7gEe5Z0_1),.clk(gclk));
	jdff dff_B_syBgmKT68_1(.din(w_dff_B_nl7gEe5Z0_1),.dout(w_dff_B_syBgmKT68_1),.clk(gclk));
	jdff dff_B_pvIK8Qgf1_1(.din(w_dff_B_syBgmKT68_1),.dout(w_dff_B_pvIK8Qgf1_1),.clk(gclk));
	jdff dff_B_ZPySYxyv9_1(.din(w_dff_B_pvIK8Qgf1_1),.dout(w_dff_B_ZPySYxyv9_1),.clk(gclk));
	jdff dff_B_1b9OPo4x8_1(.din(w_dff_B_ZPySYxyv9_1),.dout(w_dff_B_1b9OPo4x8_1),.clk(gclk));
	jdff dff_B_qAcmV4t20_1(.din(w_dff_B_1b9OPo4x8_1),.dout(w_dff_B_qAcmV4t20_1),.clk(gclk));
	jdff dff_B_8r8vNDIX4_1(.din(w_dff_B_qAcmV4t20_1),.dout(w_dff_B_8r8vNDIX4_1),.clk(gclk));
	jdff dff_B_zECH9nE16_1(.din(w_dff_B_8r8vNDIX4_1),.dout(w_dff_B_zECH9nE16_1),.clk(gclk));
	jdff dff_B_cXOIeajH7_1(.din(w_dff_B_zECH9nE16_1),.dout(w_dff_B_cXOIeajH7_1),.clk(gclk));
	jdff dff_B_GNMk3aiO0_1(.din(w_dff_B_cXOIeajH7_1),.dout(w_dff_B_GNMk3aiO0_1),.clk(gclk));
	jdff dff_B_k8b5cujs9_1(.din(w_dff_B_GNMk3aiO0_1),.dout(w_dff_B_k8b5cujs9_1),.clk(gclk));
	jdff dff_B_LhQmirqn3_0(.din(n511),.dout(w_dff_B_LhQmirqn3_0),.clk(gclk));
	jdff dff_B_3m5Josyl8_0(.din(w_dff_B_LhQmirqn3_0),.dout(w_dff_B_3m5Josyl8_0),.clk(gclk));
	jdff dff_B_MPMk29jj0_0(.din(w_dff_B_3m5Josyl8_0),.dout(w_dff_B_MPMk29jj0_0),.clk(gclk));
	jdff dff_B_Orp2IKKa9_0(.din(w_dff_B_MPMk29jj0_0),.dout(w_dff_B_Orp2IKKa9_0),.clk(gclk));
	jdff dff_B_hxwCphf05_0(.din(w_dff_B_Orp2IKKa9_0),.dout(w_dff_B_hxwCphf05_0),.clk(gclk));
	jdff dff_B_fXmjm7Bw7_0(.din(w_dff_B_hxwCphf05_0),.dout(w_dff_B_fXmjm7Bw7_0),.clk(gclk));
	jdff dff_B_Fg94zmG79_0(.din(w_dff_B_fXmjm7Bw7_0),.dout(w_dff_B_Fg94zmG79_0),.clk(gclk));
	jdff dff_B_Yarf2wHy0_0(.din(w_dff_B_Fg94zmG79_0),.dout(w_dff_B_Yarf2wHy0_0),.clk(gclk));
	jdff dff_B_xgEYqYuX6_0(.din(w_dff_B_Yarf2wHy0_0),.dout(w_dff_B_xgEYqYuX6_0),.clk(gclk));
	jdff dff_B_n4gDINIR7_0(.din(w_dff_B_xgEYqYuX6_0),.dout(w_dff_B_n4gDINIR7_0),.clk(gclk));
	jdff dff_B_IqiUbNfT0_0(.din(w_dff_B_n4gDINIR7_0),.dout(w_dff_B_IqiUbNfT0_0),.clk(gclk));
	jdff dff_B_n6VTFJq68_0(.din(w_dff_B_IqiUbNfT0_0),.dout(w_dff_B_n6VTFJq68_0),.clk(gclk));
	jdff dff_B_ieku2ZGi2_0(.din(w_dff_B_n6VTFJq68_0),.dout(w_dff_B_ieku2ZGi2_0),.clk(gclk));
	jdff dff_B_3GFJHEF15_0(.din(w_dff_B_ieku2ZGi2_0),.dout(w_dff_B_3GFJHEF15_0),.clk(gclk));
	jdff dff_B_FXOG0ofc5_0(.din(w_dff_B_3GFJHEF15_0),.dout(w_dff_B_FXOG0ofc5_0),.clk(gclk));
	jdff dff_B_kxgwOpN27_0(.din(w_dff_B_FXOG0ofc5_0),.dout(w_dff_B_kxgwOpN27_0),.clk(gclk));
	jdff dff_B_U8RnmLws4_0(.din(w_dff_B_kxgwOpN27_0),.dout(w_dff_B_U8RnmLws4_0),.clk(gclk));
	jdff dff_B_sCjKKZX31_0(.din(w_dff_B_U8RnmLws4_0),.dout(w_dff_B_sCjKKZX31_0),.clk(gclk));
	jdff dff_B_ZJUtsRPy0_0(.din(w_dff_B_sCjKKZX31_0),.dout(w_dff_B_ZJUtsRPy0_0),.clk(gclk));
	jdff dff_B_mO2p0KBo5_0(.din(w_dff_B_ZJUtsRPy0_0),.dout(w_dff_B_mO2p0KBo5_0),.clk(gclk));
	jdff dff_B_TpJykMPA5_0(.din(w_dff_B_mO2p0KBo5_0),.dout(w_dff_B_TpJykMPA5_0),.clk(gclk));
	jdff dff_B_xa5x4JPM2_1(.din(n504),.dout(w_dff_B_xa5x4JPM2_1),.clk(gclk));
	jdff dff_B_av4abSpH4_1(.din(w_dff_B_xa5x4JPM2_1),.dout(w_dff_B_av4abSpH4_1),.clk(gclk));
	jdff dff_B_7RVwqZRE9_1(.din(w_dff_B_av4abSpH4_1),.dout(w_dff_B_7RVwqZRE9_1),.clk(gclk));
	jdff dff_B_EpxKxves7_1(.din(w_dff_B_7RVwqZRE9_1),.dout(w_dff_B_EpxKxves7_1),.clk(gclk));
	jdff dff_B_dahhMMJK4_1(.din(w_dff_B_EpxKxves7_1),.dout(w_dff_B_dahhMMJK4_1),.clk(gclk));
	jdff dff_B_bTUnJ4mk9_1(.din(w_dff_B_dahhMMJK4_1),.dout(w_dff_B_bTUnJ4mk9_1),.clk(gclk));
	jdff dff_B_FtDA7Hzj1_1(.din(w_dff_B_bTUnJ4mk9_1),.dout(w_dff_B_FtDA7Hzj1_1),.clk(gclk));
	jdff dff_B_jVOJ518L1_1(.din(w_dff_B_FtDA7Hzj1_1),.dout(w_dff_B_jVOJ518L1_1),.clk(gclk));
	jdff dff_B_YrimiXEq6_1(.din(w_dff_B_jVOJ518L1_1),.dout(w_dff_B_YrimiXEq6_1),.clk(gclk));
	jdff dff_B_fwlunybC8_1(.din(w_dff_B_YrimiXEq6_1),.dout(w_dff_B_fwlunybC8_1),.clk(gclk));
	jdff dff_B_SRurwE5R8_1(.din(w_dff_B_fwlunybC8_1),.dout(w_dff_B_SRurwE5R8_1),.clk(gclk));
	jdff dff_B_pcsLQWjT7_1(.din(w_dff_B_SRurwE5R8_1),.dout(w_dff_B_pcsLQWjT7_1),.clk(gclk));
	jdff dff_B_I4OBEttl2_1(.din(w_dff_B_pcsLQWjT7_1),.dout(w_dff_B_I4OBEttl2_1),.clk(gclk));
	jdff dff_B_d9HUysRq7_1(.din(w_dff_B_I4OBEttl2_1),.dout(w_dff_B_d9HUysRq7_1),.clk(gclk));
	jdff dff_B_z3ugAY2a0_1(.din(w_dff_B_d9HUysRq7_1),.dout(w_dff_B_z3ugAY2a0_1),.clk(gclk));
	jdff dff_B_1lZkDcvQ6_1(.din(w_dff_B_z3ugAY2a0_1),.dout(w_dff_B_1lZkDcvQ6_1),.clk(gclk));
	jdff dff_B_3ZXPQKqH3_1(.din(w_dff_B_1lZkDcvQ6_1),.dout(w_dff_B_3ZXPQKqH3_1),.clk(gclk));
	jdff dff_B_k3RquIqD7_1(.din(w_dff_B_3ZXPQKqH3_1),.dout(w_dff_B_k3RquIqD7_1),.clk(gclk));
	jdff dff_B_LlQSbhOp9_1(.din(w_dff_B_k3RquIqD7_1),.dout(w_dff_B_LlQSbhOp9_1),.clk(gclk));
	jdff dff_B_wFlt2aWE8_1(.din(w_dff_B_LlQSbhOp9_1),.dout(w_dff_B_wFlt2aWE8_1),.clk(gclk));
	jdff dff_B_H3SsZrFy0_0(.din(n505),.dout(w_dff_B_H3SsZrFy0_0),.clk(gclk));
	jdff dff_B_H5otAfpI1_0(.din(w_dff_B_H3SsZrFy0_0),.dout(w_dff_B_H5otAfpI1_0),.clk(gclk));
	jdff dff_B_9b3gyfzp3_0(.din(w_dff_B_H5otAfpI1_0),.dout(w_dff_B_9b3gyfzp3_0),.clk(gclk));
	jdff dff_B_cVUdhSle8_0(.din(w_dff_B_9b3gyfzp3_0),.dout(w_dff_B_cVUdhSle8_0),.clk(gclk));
	jdff dff_B_E2LqWjd31_0(.din(w_dff_B_cVUdhSle8_0),.dout(w_dff_B_E2LqWjd31_0),.clk(gclk));
	jdff dff_B_iANMbePJ3_0(.din(w_dff_B_E2LqWjd31_0),.dout(w_dff_B_iANMbePJ3_0),.clk(gclk));
	jdff dff_B_204ll75a2_0(.din(w_dff_B_iANMbePJ3_0),.dout(w_dff_B_204ll75a2_0),.clk(gclk));
	jdff dff_B_Qpz3pLeL0_0(.din(w_dff_B_204ll75a2_0),.dout(w_dff_B_Qpz3pLeL0_0),.clk(gclk));
	jdff dff_B_RdFzMQdt7_0(.din(w_dff_B_Qpz3pLeL0_0),.dout(w_dff_B_RdFzMQdt7_0),.clk(gclk));
	jdff dff_B_nun3bSB21_0(.din(w_dff_B_RdFzMQdt7_0),.dout(w_dff_B_nun3bSB21_0),.clk(gclk));
	jdff dff_B_2oQtiWqH0_0(.din(w_dff_B_nun3bSB21_0),.dout(w_dff_B_2oQtiWqH0_0),.clk(gclk));
	jdff dff_B_D7yUlmOE0_0(.din(w_dff_B_2oQtiWqH0_0),.dout(w_dff_B_D7yUlmOE0_0),.clk(gclk));
	jdff dff_B_HjwDF7Qh8_0(.din(w_dff_B_D7yUlmOE0_0),.dout(w_dff_B_HjwDF7Qh8_0),.clk(gclk));
	jdff dff_B_lxJyeo6e9_0(.din(w_dff_B_HjwDF7Qh8_0),.dout(w_dff_B_lxJyeo6e9_0),.clk(gclk));
	jdff dff_B_Rptzv1ER2_0(.din(w_dff_B_lxJyeo6e9_0),.dout(w_dff_B_Rptzv1ER2_0),.clk(gclk));
	jdff dff_B_P6S8frr96_0(.din(w_dff_B_Rptzv1ER2_0),.dout(w_dff_B_P6S8frr96_0),.clk(gclk));
	jdff dff_B_sgXZrIhN5_0(.din(w_dff_B_P6S8frr96_0),.dout(w_dff_B_sgXZrIhN5_0),.clk(gclk));
	jdff dff_B_JPDt3g8i0_0(.din(w_dff_B_sgXZrIhN5_0),.dout(w_dff_B_JPDt3g8i0_0),.clk(gclk));
	jdff dff_B_RpyLTre07_0(.din(w_dff_B_JPDt3g8i0_0),.dout(w_dff_B_RpyLTre07_0),.clk(gclk));
	jdff dff_B_srqfiaFR0_0(.din(w_dff_B_RpyLTre07_0),.dout(w_dff_B_srqfiaFR0_0),.clk(gclk));
	jdff dff_B_7xK6EmhU6_1(.din(n498),.dout(w_dff_B_7xK6EmhU6_1),.clk(gclk));
	jdff dff_B_SPsZqQtm8_1(.din(w_dff_B_7xK6EmhU6_1),.dout(w_dff_B_SPsZqQtm8_1),.clk(gclk));
	jdff dff_B_imSWdBGf4_1(.din(w_dff_B_SPsZqQtm8_1),.dout(w_dff_B_imSWdBGf4_1),.clk(gclk));
	jdff dff_B_VGJaJ7kk0_1(.din(w_dff_B_imSWdBGf4_1),.dout(w_dff_B_VGJaJ7kk0_1),.clk(gclk));
	jdff dff_B_SGCN2dbh9_1(.din(w_dff_B_VGJaJ7kk0_1),.dout(w_dff_B_SGCN2dbh9_1),.clk(gclk));
	jdff dff_B_ZCKVZTnK8_1(.din(w_dff_B_SGCN2dbh9_1),.dout(w_dff_B_ZCKVZTnK8_1),.clk(gclk));
	jdff dff_B_jDUYEp0T5_1(.din(w_dff_B_ZCKVZTnK8_1),.dout(w_dff_B_jDUYEp0T5_1),.clk(gclk));
	jdff dff_B_Z3LhNeMH3_1(.din(w_dff_B_jDUYEp0T5_1),.dout(w_dff_B_Z3LhNeMH3_1),.clk(gclk));
	jdff dff_B_TqNQSCfI3_1(.din(w_dff_B_Z3LhNeMH3_1),.dout(w_dff_B_TqNQSCfI3_1),.clk(gclk));
	jdff dff_B_vBA2cLxo4_1(.din(w_dff_B_TqNQSCfI3_1),.dout(w_dff_B_vBA2cLxo4_1),.clk(gclk));
	jdff dff_B_fEmIoLXP6_1(.din(w_dff_B_vBA2cLxo4_1),.dout(w_dff_B_fEmIoLXP6_1),.clk(gclk));
	jdff dff_B_CysGEYLx3_1(.din(w_dff_B_fEmIoLXP6_1),.dout(w_dff_B_CysGEYLx3_1),.clk(gclk));
	jdff dff_B_ukjc9Gao2_1(.din(w_dff_B_CysGEYLx3_1),.dout(w_dff_B_ukjc9Gao2_1),.clk(gclk));
	jdff dff_B_sGVK40HI1_1(.din(w_dff_B_ukjc9Gao2_1),.dout(w_dff_B_sGVK40HI1_1),.clk(gclk));
	jdff dff_B_cdALOMMl5_1(.din(w_dff_B_sGVK40HI1_1),.dout(w_dff_B_cdALOMMl5_1),.clk(gclk));
	jdff dff_B_duGQQq2r0_1(.din(w_dff_B_cdALOMMl5_1),.dout(w_dff_B_duGQQq2r0_1),.clk(gclk));
	jdff dff_B_LwqrRRbV9_1(.din(w_dff_B_duGQQq2r0_1),.dout(w_dff_B_LwqrRRbV9_1),.clk(gclk));
	jdff dff_B_o61DiKme9_1(.din(w_dff_B_LwqrRRbV9_1),.dout(w_dff_B_o61DiKme9_1),.clk(gclk));
	jdff dff_B_eyYJitxH0_1(.din(w_dff_B_o61DiKme9_1),.dout(w_dff_B_eyYJitxH0_1),.clk(gclk));
	jdff dff_B_8w5aLc5T3_0(.din(n499),.dout(w_dff_B_8w5aLc5T3_0),.clk(gclk));
	jdff dff_B_gJywaFgx6_0(.din(w_dff_B_8w5aLc5T3_0),.dout(w_dff_B_gJywaFgx6_0),.clk(gclk));
	jdff dff_B_aBDAsdZZ9_0(.din(w_dff_B_gJywaFgx6_0),.dout(w_dff_B_aBDAsdZZ9_0),.clk(gclk));
	jdff dff_B_Q5n57uH98_0(.din(w_dff_B_aBDAsdZZ9_0),.dout(w_dff_B_Q5n57uH98_0),.clk(gclk));
	jdff dff_B_JCX5X2EQ6_0(.din(w_dff_B_Q5n57uH98_0),.dout(w_dff_B_JCX5X2EQ6_0),.clk(gclk));
	jdff dff_B_YMf9Wzeq2_0(.din(w_dff_B_JCX5X2EQ6_0),.dout(w_dff_B_YMf9Wzeq2_0),.clk(gclk));
	jdff dff_B_xxDpY2CJ6_0(.din(w_dff_B_YMf9Wzeq2_0),.dout(w_dff_B_xxDpY2CJ6_0),.clk(gclk));
	jdff dff_B_iWetE3sI0_0(.din(w_dff_B_xxDpY2CJ6_0),.dout(w_dff_B_iWetE3sI0_0),.clk(gclk));
	jdff dff_B_OFNgbhx92_0(.din(w_dff_B_iWetE3sI0_0),.dout(w_dff_B_OFNgbhx92_0),.clk(gclk));
	jdff dff_B_gMdIllk53_0(.din(w_dff_B_OFNgbhx92_0),.dout(w_dff_B_gMdIllk53_0),.clk(gclk));
	jdff dff_B_7jKOpOTx5_0(.din(w_dff_B_gMdIllk53_0),.dout(w_dff_B_7jKOpOTx5_0),.clk(gclk));
	jdff dff_B_SZvlTEXt2_0(.din(w_dff_B_7jKOpOTx5_0),.dout(w_dff_B_SZvlTEXt2_0),.clk(gclk));
	jdff dff_B_yW0M5Jdg2_0(.din(w_dff_B_SZvlTEXt2_0),.dout(w_dff_B_yW0M5Jdg2_0),.clk(gclk));
	jdff dff_B_glbPXlE80_0(.din(w_dff_B_yW0M5Jdg2_0),.dout(w_dff_B_glbPXlE80_0),.clk(gclk));
	jdff dff_B_iCpyig4C6_0(.din(w_dff_B_glbPXlE80_0),.dout(w_dff_B_iCpyig4C6_0),.clk(gclk));
	jdff dff_B_VkNIvHyH4_0(.din(w_dff_B_iCpyig4C6_0),.dout(w_dff_B_VkNIvHyH4_0),.clk(gclk));
	jdff dff_B_5aHwBBEa3_0(.din(w_dff_B_VkNIvHyH4_0),.dout(w_dff_B_5aHwBBEa3_0),.clk(gclk));
	jdff dff_B_TNHDgILC3_0(.din(w_dff_B_5aHwBBEa3_0),.dout(w_dff_B_TNHDgILC3_0),.clk(gclk));
	jdff dff_B_CcU9AiUi0_0(.din(w_dff_B_TNHDgILC3_0),.dout(w_dff_B_CcU9AiUi0_0),.clk(gclk));
	jdff dff_B_DsqcDONC2_1(.din(n492),.dout(w_dff_B_DsqcDONC2_1),.clk(gclk));
	jdff dff_B_qEY7xbD11_1(.din(w_dff_B_DsqcDONC2_1),.dout(w_dff_B_qEY7xbD11_1),.clk(gclk));
	jdff dff_B_AZSKonBw8_1(.din(w_dff_B_qEY7xbD11_1),.dout(w_dff_B_AZSKonBw8_1),.clk(gclk));
	jdff dff_B_T86nmV2p3_1(.din(w_dff_B_AZSKonBw8_1),.dout(w_dff_B_T86nmV2p3_1),.clk(gclk));
	jdff dff_B_1fBNeVli2_1(.din(w_dff_B_T86nmV2p3_1),.dout(w_dff_B_1fBNeVli2_1),.clk(gclk));
	jdff dff_B_82Rxo4n26_1(.din(w_dff_B_1fBNeVli2_1),.dout(w_dff_B_82Rxo4n26_1),.clk(gclk));
	jdff dff_B_99fEhW9B9_1(.din(w_dff_B_82Rxo4n26_1),.dout(w_dff_B_99fEhW9B9_1),.clk(gclk));
	jdff dff_B_M1gUdRdO6_1(.din(w_dff_B_99fEhW9B9_1),.dout(w_dff_B_M1gUdRdO6_1),.clk(gclk));
	jdff dff_B_idh8pFW65_1(.din(w_dff_B_M1gUdRdO6_1),.dout(w_dff_B_idh8pFW65_1),.clk(gclk));
	jdff dff_B_Ew5zMVam9_1(.din(w_dff_B_idh8pFW65_1),.dout(w_dff_B_Ew5zMVam9_1),.clk(gclk));
	jdff dff_B_hMLPG4LO5_1(.din(w_dff_B_Ew5zMVam9_1),.dout(w_dff_B_hMLPG4LO5_1),.clk(gclk));
	jdff dff_B_EEc5s4PX5_1(.din(w_dff_B_hMLPG4LO5_1),.dout(w_dff_B_EEc5s4PX5_1),.clk(gclk));
	jdff dff_B_qdyNlzfl1_1(.din(w_dff_B_EEc5s4PX5_1),.dout(w_dff_B_qdyNlzfl1_1),.clk(gclk));
	jdff dff_B_AW4wJHbW8_1(.din(w_dff_B_qdyNlzfl1_1),.dout(w_dff_B_AW4wJHbW8_1),.clk(gclk));
	jdff dff_B_lLRNHaXk1_1(.din(w_dff_B_AW4wJHbW8_1),.dout(w_dff_B_lLRNHaXk1_1),.clk(gclk));
	jdff dff_B_nUz2s5yt4_1(.din(w_dff_B_lLRNHaXk1_1),.dout(w_dff_B_nUz2s5yt4_1),.clk(gclk));
	jdff dff_B_pP5A4g558_1(.din(w_dff_B_nUz2s5yt4_1),.dout(w_dff_B_pP5A4g558_1),.clk(gclk));
	jdff dff_B_EWKSzcRm1_1(.din(w_dff_B_pP5A4g558_1),.dout(w_dff_B_EWKSzcRm1_1),.clk(gclk));
	jdff dff_B_qPGFOp2M9_0(.din(n493),.dout(w_dff_B_qPGFOp2M9_0),.clk(gclk));
	jdff dff_B_Q6xMljOf6_0(.din(w_dff_B_qPGFOp2M9_0),.dout(w_dff_B_Q6xMljOf6_0),.clk(gclk));
	jdff dff_B_TzODdsoK2_0(.din(w_dff_B_Q6xMljOf6_0),.dout(w_dff_B_TzODdsoK2_0),.clk(gclk));
	jdff dff_B_1HHyb4Xq0_0(.din(w_dff_B_TzODdsoK2_0),.dout(w_dff_B_1HHyb4Xq0_0),.clk(gclk));
	jdff dff_B_aGWFNs8B4_0(.din(w_dff_B_1HHyb4Xq0_0),.dout(w_dff_B_aGWFNs8B4_0),.clk(gclk));
	jdff dff_B_atTLjLDJ8_0(.din(w_dff_B_aGWFNs8B4_0),.dout(w_dff_B_atTLjLDJ8_0),.clk(gclk));
	jdff dff_B_akv8Vddd3_0(.din(w_dff_B_atTLjLDJ8_0),.dout(w_dff_B_akv8Vddd3_0),.clk(gclk));
	jdff dff_B_QOhnN9BP5_0(.din(w_dff_B_akv8Vddd3_0),.dout(w_dff_B_QOhnN9BP5_0),.clk(gclk));
	jdff dff_B_ak1MbCZO2_0(.din(w_dff_B_QOhnN9BP5_0),.dout(w_dff_B_ak1MbCZO2_0),.clk(gclk));
	jdff dff_B_eubY1vOU3_0(.din(w_dff_B_ak1MbCZO2_0),.dout(w_dff_B_eubY1vOU3_0),.clk(gclk));
	jdff dff_B_OeRke0uK6_0(.din(w_dff_B_eubY1vOU3_0),.dout(w_dff_B_OeRke0uK6_0),.clk(gclk));
	jdff dff_B_JX7VGQvK9_0(.din(w_dff_B_OeRke0uK6_0),.dout(w_dff_B_JX7VGQvK9_0),.clk(gclk));
	jdff dff_B_mOpQjRKP9_0(.din(w_dff_B_JX7VGQvK9_0),.dout(w_dff_B_mOpQjRKP9_0),.clk(gclk));
	jdff dff_B_upekkd5I8_0(.din(w_dff_B_mOpQjRKP9_0),.dout(w_dff_B_upekkd5I8_0),.clk(gclk));
	jdff dff_B_Vql2Za4h8_0(.din(w_dff_B_upekkd5I8_0),.dout(w_dff_B_Vql2Za4h8_0),.clk(gclk));
	jdff dff_B_QMvYmRMk4_0(.din(w_dff_B_Vql2Za4h8_0),.dout(w_dff_B_QMvYmRMk4_0),.clk(gclk));
	jdff dff_B_IGdmWZAf5_0(.din(w_dff_B_QMvYmRMk4_0),.dout(w_dff_B_IGdmWZAf5_0),.clk(gclk));
	jdff dff_B_bS2zNEr15_0(.din(w_dff_B_IGdmWZAf5_0),.dout(w_dff_B_bS2zNEr15_0),.clk(gclk));
	jdff dff_B_DtGIA1Qr8_1(.din(n486),.dout(w_dff_B_DtGIA1Qr8_1),.clk(gclk));
	jdff dff_B_TClm6Gwg8_1(.din(w_dff_B_DtGIA1Qr8_1),.dout(w_dff_B_TClm6Gwg8_1),.clk(gclk));
	jdff dff_B_cQPMdY607_1(.din(w_dff_B_TClm6Gwg8_1),.dout(w_dff_B_cQPMdY607_1),.clk(gclk));
	jdff dff_B_OWOQHXBv3_1(.din(w_dff_B_cQPMdY607_1),.dout(w_dff_B_OWOQHXBv3_1),.clk(gclk));
	jdff dff_B_zJjkWGXe6_1(.din(w_dff_B_OWOQHXBv3_1),.dout(w_dff_B_zJjkWGXe6_1),.clk(gclk));
	jdff dff_B_3jo62fHS0_1(.din(w_dff_B_zJjkWGXe6_1),.dout(w_dff_B_3jo62fHS0_1),.clk(gclk));
	jdff dff_B_hSUjpPmh8_1(.din(w_dff_B_3jo62fHS0_1),.dout(w_dff_B_hSUjpPmh8_1),.clk(gclk));
	jdff dff_B_Ub5VEuQF6_1(.din(w_dff_B_hSUjpPmh8_1),.dout(w_dff_B_Ub5VEuQF6_1),.clk(gclk));
	jdff dff_B_peaUIY4i2_1(.din(w_dff_B_Ub5VEuQF6_1),.dout(w_dff_B_peaUIY4i2_1),.clk(gclk));
	jdff dff_B_SW51JjHT7_1(.din(w_dff_B_peaUIY4i2_1),.dout(w_dff_B_SW51JjHT7_1),.clk(gclk));
	jdff dff_B_Lla3yk331_1(.din(w_dff_B_SW51JjHT7_1),.dout(w_dff_B_Lla3yk331_1),.clk(gclk));
	jdff dff_B_1PU1J8NF4_1(.din(w_dff_B_Lla3yk331_1),.dout(w_dff_B_1PU1J8NF4_1),.clk(gclk));
	jdff dff_B_RGGE4mWw1_1(.din(w_dff_B_1PU1J8NF4_1),.dout(w_dff_B_RGGE4mWw1_1),.clk(gclk));
	jdff dff_B_CQkr8GgQ9_1(.din(w_dff_B_RGGE4mWw1_1),.dout(w_dff_B_CQkr8GgQ9_1),.clk(gclk));
	jdff dff_B_ejvwjjJS3_1(.din(w_dff_B_CQkr8GgQ9_1),.dout(w_dff_B_ejvwjjJS3_1),.clk(gclk));
	jdff dff_B_aIm1Iwxd0_1(.din(w_dff_B_ejvwjjJS3_1),.dout(w_dff_B_aIm1Iwxd0_1),.clk(gclk));
	jdff dff_B_LxQ84mjb0_1(.din(w_dff_B_aIm1Iwxd0_1),.dout(w_dff_B_LxQ84mjb0_1),.clk(gclk));
	jdff dff_B_4cj0w4qp2_0(.din(n487),.dout(w_dff_B_4cj0w4qp2_0),.clk(gclk));
	jdff dff_B_ttfr3fBJ7_0(.din(w_dff_B_4cj0w4qp2_0),.dout(w_dff_B_ttfr3fBJ7_0),.clk(gclk));
	jdff dff_B_IjsRDjAf5_0(.din(w_dff_B_ttfr3fBJ7_0),.dout(w_dff_B_IjsRDjAf5_0),.clk(gclk));
	jdff dff_B_Q4n4QISs2_0(.din(w_dff_B_IjsRDjAf5_0),.dout(w_dff_B_Q4n4QISs2_0),.clk(gclk));
	jdff dff_B_UzWE0xuc0_0(.din(w_dff_B_Q4n4QISs2_0),.dout(w_dff_B_UzWE0xuc0_0),.clk(gclk));
	jdff dff_B_G8UOLQmu2_0(.din(w_dff_B_UzWE0xuc0_0),.dout(w_dff_B_G8UOLQmu2_0),.clk(gclk));
	jdff dff_B_SRkte2WQ7_0(.din(w_dff_B_G8UOLQmu2_0),.dout(w_dff_B_SRkte2WQ7_0),.clk(gclk));
	jdff dff_B_y7IBRBiF8_0(.din(w_dff_B_SRkte2WQ7_0),.dout(w_dff_B_y7IBRBiF8_0),.clk(gclk));
	jdff dff_B_XVFsoCZ73_0(.din(w_dff_B_y7IBRBiF8_0),.dout(w_dff_B_XVFsoCZ73_0),.clk(gclk));
	jdff dff_B_5geMDvRG6_0(.din(w_dff_B_XVFsoCZ73_0),.dout(w_dff_B_5geMDvRG6_0),.clk(gclk));
	jdff dff_B_StHB7Yd60_0(.din(w_dff_B_5geMDvRG6_0),.dout(w_dff_B_StHB7Yd60_0),.clk(gclk));
	jdff dff_B_AL3LKkyJ7_0(.din(w_dff_B_StHB7Yd60_0),.dout(w_dff_B_AL3LKkyJ7_0),.clk(gclk));
	jdff dff_B_lNiXWzoT9_0(.din(w_dff_B_AL3LKkyJ7_0),.dout(w_dff_B_lNiXWzoT9_0),.clk(gclk));
	jdff dff_B_I0pcZiVS8_0(.din(w_dff_B_lNiXWzoT9_0),.dout(w_dff_B_I0pcZiVS8_0),.clk(gclk));
	jdff dff_B_ylFPqo4h2_0(.din(w_dff_B_I0pcZiVS8_0),.dout(w_dff_B_ylFPqo4h2_0),.clk(gclk));
	jdff dff_B_UXzqSjqs2_0(.din(w_dff_B_ylFPqo4h2_0),.dout(w_dff_B_UXzqSjqs2_0),.clk(gclk));
	jdff dff_B_M2JhGCeu4_0(.din(w_dff_B_UXzqSjqs2_0),.dout(w_dff_B_M2JhGCeu4_0),.clk(gclk));
	jdff dff_B_5S7dBTMF2_1(.din(n480),.dout(w_dff_B_5S7dBTMF2_1),.clk(gclk));
	jdff dff_B_H66g06Jv7_1(.din(w_dff_B_5S7dBTMF2_1),.dout(w_dff_B_H66g06Jv7_1),.clk(gclk));
	jdff dff_B_eqgmM5eX7_1(.din(w_dff_B_H66g06Jv7_1),.dout(w_dff_B_eqgmM5eX7_1),.clk(gclk));
	jdff dff_B_nrlqClN77_1(.din(w_dff_B_eqgmM5eX7_1),.dout(w_dff_B_nrlqClN77_1),.clk(gclk));
	jdff dff_B_zDiHmWge8_1(.din(w_dff_B_nrlqClN77_1),.dout(w_dff_B_zDiHmWge8_1),.clk(gclk));
	jdff dff_B_3T24PzSq4_1(.din(w_dff_B_zDiHmWge8_1),.dout(w_dff_B_3T24PzSq4_1),.clk(gclk));
	jdff dff_B_6v6jhMIb4_1(.din(w_dff_B_3T24PzSq4_1),.dout(w_dff_B_6v6jhMIb4_1),.clk(gclk));
	jdff dff_B_9YuYCD3O9_1(.din(w_dff_B_6v6jhMIb4_1),.dout(w_dff_B_9YuYCD3O9_1),.clk(gclk));
	jdff dff_B_bUSViud42_1(.din(w_dff_B_9YuYCD3O9_1),.dout(w_dff_B_bUSViud42_1),.clk(gclk));
	jdff dff_B_egv2g8IU9_1(.din(w_dff_B_bUSViud42_1),.dout(w_dff_B_egv2g8IU9_1),.clk(gclk));
	jdff dff_B_Cvh92W7r2_1(.din(w_dff_B_egv2g8IU9_1),.dout(w_dff_B_Cvh92W7r2_1),.clk(gclk));
	jdff dff_B_mowFca6I7_1(.din(w_dff_B_Cvh92W7r2_1),.dout(w_dff_B_mowFca6I7_1),.clk(gclk));
	jdff dff_B_hZppC5Ry8_1(.din(w_dff_B_mowFca6I7_1),.dout(w_dff_B_hZppC5Ry8_1),.clk(gclk));
	jdff dff_B_buqsmvbG4_1(.din(w_dff_B_hZppC5Ry8_1),.dout(w_dff_B_buqsmvbG4_1),.clk(gclk));
	jdff dff_B_rZuwkguI5_1(.din(w_dff_B_buqsmvbG4_1),.dout(w_dff_B_rZuwkguI5_1),.clk(gclk));
	jdff dff_B_ghzowI0M3_1(.din(w_dff_B_rZuwkguI5_1),.dout(w_dff_B_ghzowI0M3_1),.clk(gclk));
	jdff dff_B_Gs3icwdR1_0(.din(n481),.dout(w_dff_B_Gs3icwdR1_0),.clk(gclk));
	jdff dff_B_2m4GT23m8_0(.din(w_dff_B_Gs3icwdR1_0),.dout(w_dff_B_2m4GT23m8_0),.clk(gclk));
	jdff dff_B_6fJxv6bY6_0(.din(w_dff_B_2m4GT23m8_0),.dout(w_dff_B_6fJxv6bY6_0),.clk(gclk));
	jdff dff_B_sBPeg4QF7_0(.din(w_dff_B_6fJxv6bY6_0),.dout(w_dff_B_sBPeg4QF7_0),.clk(gclk));
	jdff dff_B_DrHk8ME58_0(.din(w_dff_B_sBPeg4QF7_0),.dout(w_dff_B_DrHk8ME58_0),.clk(gclk));
	jdff dff_B_ge20eKXn4_0(.din(w_dff_B_DrHk8ME58_0),.dout(w_dff_B_ge20eKXn4_0),.clk(gclk));
	jdff dff_B_YzzD5oRv5_0(.din(w_dff_B_ge20eKXn4_0),.dout(w_dff_B_YzzD5oRv5_0),.clk(gclk));
	jdff dff_B_m4ChRGeD3_0(.din(w_dff_B_YzzD5oRv5_0),.dout(w_dff_B_m4ChRGeD3_0),.clk(gclk));
	jdff dff_B_tBNOCMDy4_0(.din(w_dff_B_m4ChRGeD3_0),.dout(w_dff_B_tBNOCMDy4_0),.clk(gclk));
	jdff dff_B_TKgZ6uI55_0(.din(w_dff_B_tBNOCMDy4_0),.dout(w_dff_B_TKgZ6uI55_0),.clk(gclk));
	jdff dff_B_Wq8VXjwJ4_0(.din(w_dff_B_TKgZ6uI55_0),.dout(w_dff_B_Wq8VXjwJ4_0),.clk(gclk));
	jdff dff_B_cyAFaND39_0(.din(w_dff_B_Wq8VXjwJ4_0),.dout(w_dff_B_cyAFaND39_0),.clk(gclk));
	jdff dff_B_cSwYfqwq8_0(.din(w_dff_B_cyAFaND39_0),.dout(w_dff_B_cSwYfqwq8_0),.clk(gclk));
	jdff dff_B_aBR3e6eT0_0(.din(w_dff_B_cSwYfqwq8_0),.dout(w_dff_B_aBR3e6eT0_0),.clk(gclk));
	jdff dff_B_w2W4jLg07_0(.din(w_dff_B_aBR3e6eT0_0),.dout(w_dff_B_w2W4jLg07_0),.clk(gclk));
	jdff dff_B_Ps1HkcOR8_0(.din(w_dff_B_w2W4jLg07_0),.dout(w_dff_B_Ps1HkcOR8_0),.clk(gclk));
	jdff dff_B_CUOXvnUc5_1(.din(n474),.dout(w_dff_B_CUOXvnUc5_1),.clk(gclk));
	jdff dff_B_HPfjBPEr9_1(.din(w_dff_B_CUOXvnUc5_1),.dout(w_dff_B_HPfjBPEr9_1),.clk(gclk));
	jdff dff_B_PGPELzGd7_1(.din(w_dff_B_HPfjBPEr9_1),.dout(w_dff_B_PGPELzGd7_1),.clk(gclk));
	jdff dff_B_Kb2hf6kc5_1(.din(w_dff_B_PGPELzGd7_1),.dout(w_dff_B_Kb2hf6kc5_1),.clk(gclk));
	jdff dff_B_sjwpyMU29_1(.din(w_dff_B_Kb2hf6kc5_1),.dout(w_dff_B_sjwpyMU29_1),.clk(gclk));
	jdff dff_B_tspZSzwa7_1(.din(w_dff_B_sjwpyMU29_1),.dout(w_dff_B_tspZSzwa7_1),.clk(gclk));
	jdff dff_B_NVQoXH6E9_1(.din(w_dff_B_tspZSzwa7_1),.dout(w_dff_B_NVQoXH6E9_1),.clk(gclk));
	jdff dff_B_YUo1Ygd56_1(.din(w_dff_B_NVQoXH6E9_1),.dout(w_dff_B_YUo1Ygd56_1),.clk(gclk));
	jdff dff_B_6Rm8qGhB8_1(.din(w_dff_B_YUo1Ygd56_1),.dout(w_dff_B_6Rm8qGhB8_1),.clk(gclk));
	jdff dff_B_lvZN4CVJ2_1(.din(w_dff_B_6Rm8qGhB8_1),.dout(w_dff_B_lvZN4CVJ2_1),.clk(gclk));
	jdff dff_B_gxtRfNv60_1(.din(w_dff_B_lvZN4CVJ2_1),.dout(w_dff_B_gxtRfNv60_1),.clk(gclk));
	jdff dff_B_ikB8jArh1_1(.din(w_dff_B_gxtRfNv60_1),.dout(w_dff_B_ikB8jArh1_1),.clk(gclk));
	jdff dff_B_odm2xBLw5_1(.din(w_dff_B_ikB8jArh1_1),.dout(w_dff_B_odm2xBLw5_1),.clk(gclk));
	jdff dff_B_m9q3uzCY6_1(.din(w_dff_B_odm2xBLw5_1),.dout(w_dff_B_m9q3uzCY6_1),.clk(gclk));
	jdff dff_B_ORoqjfaO4_1(.din(w_dff_B_m9q3uzCY6_1),.dout(w_dff_B_ORoqjfaO4_1),.clk(gclk));
	jdff dff_B_sXbzJ5Q78_0(.din(n475),.dout(w_dff_B_sXbzJ5Q78_0),.clk(gclk));
	jdff dff_B_rQsG1VQ11_0(.din(w_dff_B_sXbzJ5Q78_0),.dout(w_dff_B_rQsG1VQ11_0),.clk(gclk));
	jdff dff_B_gHa8KuJC1_0(.din(w_dff_B_rQsG1VQ11_0),.dout(w_dff_B_gHa8KuJC1_0),.clk(gclk));
	jdff dff_B_UTQABHOg7_0(.din(w_dff_B_gHa8KuJC1_0),.dout(w_dff_B_UTQABHOg7_0),.clk(gclk));
	jdff dff_B_AbJRHRrv1_0(.din(w_dff_B_UTQABHOg7_0),.dout(w_dff_B_AbJRHRrv1_0),.clk(gclk));
	jdff dff_B_46AXX8fY8_0(.din(w_dff_B_AbJRHRrv1_0),.dout(w_dff_B_46AXX8fY8_0),.clk(gclk));
	jdff dff_B_3z2JPzpZ4_0(.din(w_dff_B_46AXX8fY8_0),.dout(w_dff_B_3z2JPzpZ4_0),.clk(gclk));
	jdff dff_B_JTqh1Zvp5_0(.din(w_dff_B_3z2JPzpZ4_0),.dout(w_dff_B_JTqh1Zvp5_0),.clk(gclk));
	jdff dff_B_pi3yEozm0_0(.din(w_dff_B_JTqh1Zvp5_0),.dout(w_dff_B_pi3yEozm0_0),.clk(gclk));
	jdff dff_B_HQGS0GVA7_0(.din(w_dff_B_pi3yEozm0_0),.dout(w_dff_B_HQGS0GVA7_0),.clk(gclk));
	jdff dff_B_lO38nP6x1_0(.din(w_dff_B_HQGS0GVA7_0),.dout(w_dff_B_lO38nP6x1_0),.clk(gclk));
	jdff dff_B_sknHGjTq1_0(.din(w_dff_B_lO38nP6x1_0),.dout(w_dff_B_sknHGjTq1_0),.clk(gclk));
	jdff dff_B_phSHpzuI8_0(.din(w_dff_B_sknHGjTq1_0),.dout(w_dff_B_phSHpzuI8_0),.clk(gclk));
	jdff dff_B_YlwRzazy5_0(.din(w_dff_B_phSHpzuI8_0),.dout(w_dff_B_YlwRzazy5_0),.clk(gclk));
	jdff dff_B_Azuoeek25_0(.din(w_dff_B_YlwRzazy5_0),.dout(w_dff_B_Azuoeek25_0),.clk(gclk));
	jdff dff_B_hyJeNg6b4_1(.din(n468),.dout(w_dff_B_hyJeNg6b4_1),.clk(gclk));
	jdff dff_B_eiqVd13B5_1(.din(w_dff_B_hyJeNg6b4_1),.dout(w_dff_B_eiqVd13B5_1),.clk(gclk));
	jdff dff_B_zyDhBBD60_1(.din(w_dff_B_eiqVd13B5_1),.dout(w_dff_B_zyDhBBD60_1),.clk(gclk));
	jdff dff_B_Mi3poAXu6_1(.din(w_dff_B_zyDhBBD60_1),.dout(w_dff_B_Mi3poAXu6_1),.clk(gclk));
	jdff dff_B_gE4KwiDc3_1(.din(w_dff_B_Mi3poAXu6_1),.dout(w_dff_B_gE4KwiDc3_1),.clk(gclk));
	jdff dff_B_Ev1G5wgk2_1(.din(w_dff_B_gE4KwiDc3_1),.dout(w_dff_B_Ev1G5wgk2_1),.clk(gclk));
	jdff dff_B_fNerFjHe8_1(.din(w_dff_B_Ev1G5wgk2_1),.dout(w_dff_B_fNerFjHe8_1),.clk(gclk));
	jdff dff_B_Qe6Tvfbg1_1(.din(w_dff_B_fNerFjHe8_1),.dout(w_dff_B_Qe6Tvfbg1_1),.clk(gclk));
	jdff dff_B_vcXp2qKs8_1(.din(w_dff_B_Qe6Tvfbg1_1),.dout(w_dff_B_vcXp2qKs8_1),.clk(gclk));
	jdff dff_B_zpcHU6sG8_1(.din(w_dff_B_vcXp2qKs8_1),.dout(w_dff_B_zpcHU6sG8_1),.clk(gclk));
	jdff dff_B_XDopxJbJ5_1(.din(w_dff_B_zpcHU6sG8_1),.dout(w_dff_B_XDopxJbJ5_1),.clk(gclk));
	jdff dff_B_vbZvn9X06_1(.din(w_dff_B_XDopxJbJ5_1),.dout(w_dff_B_vbZvn9X06_1),.clk(gclk));
	jdff dff_B_WgGQvFyk8_1(.din(w_dff_B_vbZvn9X06_1),.dout(w_dff_B_WgGQvFyk8_1),.clk(gclk));
	jdff dff_B_LgXnSLIA1_1(.din(w_dff_B_WgGQvFyk8_1),.dout(w_dff_B_LgXnSLIA1_1),.clk(gclk));
	jdff dff_B_fEYIY6q44_0(.din(n469),.dout(w_dff_B_fEYIY6q44_0),.clk(gclk));
	jdff dff_B_kXVhlyVg4_0(.din(w_dff_B_fEYIY6q44_0),.dout(w_dff_B_kXVhlyVg4_0),.clk(gclk));
	jdff dff_B_kpZkyfY87_0(.din(w_dff_B_kXVhlyVg4_0),.dout(w_dff_B_kpZkyfY87_0),.clk(gclk));
	jdff dff_B_uy1hztZS6_0(.din(w_dff_B_kpZkyfY87_0),.dout(w_dff_B_uy1hztZS6_0),.clk(gclk));
	jdff dff_B_69c0OADM1_0(.din(w_dff_B_uy1hztZS6_0),.dout(w_dff_B_69c0OADM1_0),.clk(gclk));
	jdff dff_B_QJzL0RRy6_0(.din(w_dff_B_69c0OADM1_0),.dout(w_dff_B_QJzL0RRy6_0),.clk(gclk));
	jdff dff_B_ibk2HsTc8_0(.din(w_dff_B_QJzL0RRy6_0),.dout(w_dff_B_ibk2HsTc8_0),.clk(gclk));
	jdff dff_B_86zqUp2N9_0(.din(w_dff_B_ibk2HsTc8_0),.dout(w_dff_B_86zqUp2N9_0),.clk(gclk));
	jdff dff_B_OW9IdvrP2_0(.din(w_dff_B_86zqUp2N9_0),.dout(w_dff_B_OW9IdvrP2_0),.clk(gclk));
	jdff dff_B_2h6rtg9U0_0(.din(w_dff_B_OW9IdvrP2_0),.dout(w_dff_B_2h6rtg9U0_0),.clk(gclk));
	jdff dff_B_TDMm0ipE7_0(.din(w_dff_B_2h6rtg9U0_0),.dout(w_dff_B_TDMm0ipE7_0),.clk(gclk));
	jdff dff_B_FxCCraqz2_0(.din(w_dff_B_TDMm0ipE7_0),.dout(w_dff_B_FxCCraqz2_0),.clk(gclk));
	jdff dff_B_b858IeTD0_0(.din(w_dff_B_FxCCraqz2_0),.dout(w_dff_B_b858IeTD0_0),.clk(gclk));
	jdff dff_B_bY5KWRW79_0(.din(w_dff_B_b858IeTD0_0),.dout(w_dff_B_bY5KWRW79_0),.clk(gclk));
	jdff dff_B_EVgls9Hj2_1(.din(n462),.dout(w_dff_B_EVgls9Hj2_1),.clk(gclk));
	jdff dff_B_wKsM1TJx2_1(.din(w_dff_B_EVgls9Hj2_1),.dout(w_dff_B_wKsM1TJx2_1),.clk(gclk));
	jdff dff_B_llvWFGdo3_1(.din(w_dff_B_wKsM1TJx2_1),.dout(w_dff_B_llvWFGdo3_1),.clk(gclk));
	jdff dff_B_hNfCcbQL1_1(.din(w_dff_B_llvWFGdo3_1),.dout(w_dff_B_hNfCcbQL1_1),.clk(gclk));
	jdff dff_B_36yABsft3_1(.din(w_dff_B_hNfCcbQL1_1),.dout(w_dff_B_36yABsft3_1),.clk(gclk));
	jdff dff_B_FMp0B9V20_1(.din(w_dff_B_36yABsft3_1),.dout(w_dff_B_FMp0B9V20_1),.clk(gclk));
	jdff dff_B_p7VG3Aqa4_1(.din(w_dff_B_FMp0B9V20_1),.dout(w_dff_B_p7VG3Aqa4_1),.clk(gclk));
	jdff dff_B_YlZbSA8n2_1(.din(w_dff_B_p7VG3Aqa4_1),.dout(w_dff_B_YlZbSA8n2_1),.clk(gclk));
	jdff dff_B_GTIBmeFe0_1(.din(w_dff_B_YlZbSA8n2_1),.dout(w_dff_B_GTIBmeFe0_1),.clk(gclk));
	jdff dff_B_BjNPsRSJ7_1(.din(w_dff_B_GTIBmeFe0_1),.dout(w_dff_B_BjNPsRSJ7_1),.clk(gclk));
	jdff dff_B_4bEbYv7J7_1(.din(w_dff_B_BjNPsRSJ7_1),.dout(w_dff_B_4bEbYv7J7_1),.clk(gclk));
	jdff dff_B_lUDUU1OZ7_1(.din(w_dff_B_4bEbYv7J7_1),.dout(w_dff_B_lUDUU1OZ7_1),.clk(gclk));
	jdff dff_B_EbOdpOXS9_1(.din(w_dff_B_lUDUU1OZ7_1),.dout(w_dff_B_EbOdpOXS9_1),.clk(gclk));
	jdff dff_B_5CeuyEaX6_0(.din(n463),.dout(w_dff_B_5CeuyEaX6_0),.clk(gclk));
	jdff dff_B_a5tanuw44_0(.din(w_dff_B_5CeuyEaX6_0),.dout(w_dff_B_a5tanuw44_0),.clk(gclk));
	jdff dff_B_p1SXfKS10_0(.din(w_dff_B_a5tanuw44_0),.dout(w_dff_B_p1SXfKS10_0),.clk(gclk));
	jdff dff_B_yHilQjpp3_0(.din(w_dff_B_p1SXfKS10_0),.dout(w_dff_B_yHilQjpp3_0),.clk(gclk));
	jdff dff_B_RTwv84eT1_0(.din(w_dff_B_yHilQjpp3_0),.dout(w_dff_B_RTwv84eT1_0),.clk(gclk));
	jdff dff_B_sI2dhu6C0_0(.din(w_dff_B_RTwv84eT1_0),.dout(w_dff_B_sI2dhu6C0_0),.clk(gclk));
	jdff dff_B_s6pp4PGW1_0(.din(w_dff_B_sI2dhu6C0_0),.dout(w_dff_B_s6pp4PGW1_0),.clk(gclk));
	jdff dff_B_NlD4pJqc0_0(.din(w_dff_B_s6pp4PGW1_0),.dout(w_dff_B_NlD4pJqc0_0),.clk(gclk));
	jdff dff_B_1AX1uVCb8_0(.din(w_dff_B_NlD4pJqc0_0),.dout(w_dff_B_1AX1uVCb8_0),.clk(gclk));
	jdff dff_B_VugXbhlk9_0(.din(w_dff_B_1AX1uVCb8_0),.dout(w_dff_B_VugXbhlk9_0),.clk(gclk));
	jdff dff_B_q5dE9HBj3_0(.din(w_dff_B_VugXbhlk9_0),.dout(w_dff_B_q5dE9HBj3_0),.clk(gclk));
	jdff dff_B_RKWmxwpd3_0(.din(w_dff_B_q5dE9HBj3_0),.dout(w_dff_B_RKWmxwpd3_0),.clk(gclk));
	jdff dff_B_hz8fGERr9_0(.din(w_dff_B_RKWmxwpd3_0),.dout(w_dff_B_hz8fGERr9_0),.clk(gclk));
	jdff dff_B_xgqsNOXB1_1(.din(n456),.dout(w_dff_B_xgqsNOXB1_1),.clk(gclk));
	jdff dff_B_NWHntx2t2_1(.din(w_dff_B_xgqsNOXB1_1),.dout(w_dff_B_NWHntx2t2_1),.clk(gclk));
	jdff dff_B_AlPmFwRW4_1(.din(w_dff_B_NWHntx2t2_1),.dout(w_dff_B_AlPmFwRW4_1),.clk(gclk));
	jdff dff_B_2a8lfKA75_1(.din(w_dff_B_AlPmFwRW4_1),.dout(w_dff_B_2a8lfKA75_1),.clk(gclk));
	jdff dff_B_XxLjBnFw8_1(.din(w_dff_B_2a8lfKA75_1),.dout(w_dff_B_XxLjBnFw8_1),.clk(gclk));
	jdff dff_B_NBWtTwgR2_1(.din(w_dff_B_XxLjBnFw8_1),.dout(w_dff_B_NBWtTwgR2_1),.clk(gclk));
	jdff dff_B_Okr54iu12_1(.din(w_dff_B_NBWtTwgR2_1),.dout(w_dff_B_Okr54iu12_1),.clk(gclk));
	jdff dff_B_6Jsg1KBg1_1(.din(w_dff_B_Okr54iu12_1),.dout(w_dff_B_6Jsg1KBg1_1),.clk(gclk));
	jdff dff_B_g5zSm0bu7_1(.din(w_dff_B_6Jsg1KBg1_1),.dout(w_dff_B_g5zSm0bu7_1),.clk(gclk));
	jdff dff_B_FPt83beR7_1(.din(w_dff_B_g5zSm0bu7_1),.dout(w_dff_B_FPt83beR7_1),.clk(gclk));
	jdff dff_B_8JMvHWgE6_1(.din(w_dff_B_FPt83beR7_1),.dout(w_dff_B_8JMvHWgE6_1),.clk(gclk));
	jdff dff_B_Uziv0Vnv8_1(.din(w_dff_B_8JMvHWgE6_1),.dout(w_dff_B_Uziv0Vnv8_1),.clk(gclk));
	jdff dff_B_9AR7u68N2_0(.din(n457),.dout(w_dff_B_9AR7u68N2_0),.clk(gclk));
	jdff dff_B_TbnkcOLG4_0(.din(w_dff_B_9AR7u68N2_0),.dout(w_dff_B_TbnkcOLG4_0),.clk(gclk));
	jdff dff_B_RR9bi7VC1_0(.din(w_dff_B_TbnkcOLG4_0),.dout(w_dff_B_RR9bi7VC1_0),.clk(gclk));
	jdff dff_B_oT1a1THS1_0(.din(w_dff_B_RR9bi7VC1_0),.dout(w_dff_B_oT1a1THS1_0),.clk(gclk));
	jdff dff_B_uZLVjhAF8_0(.din(w_dff_B_oT1a1THS1_0),.dout(w_dff_B_uZLVjhAF8_0),.clk(gclk));
	jdff dff_B_DHQwpGTR8_0(.din(w_dff_B_uZLVjhAF8_0),.dout(w_dff_B_DHQwpGTR8_0),.clk(gclk));
	jdff dff_B_u02w9fFj6_0(.din(w_dff_B_DHQwpGTR8_0),.dout(w_dff_B_u02w9fFj6_0),.clk(gclk));
	jdff dff_B_sfoT66hB2_0(.din(w_dff_B_u02w9fFj6_0),.dout(w_dff_B_sfoT66hB2_0),.clk(gclk));
	jdff dff_B_dmAlHyGz0_0(.din(w_dff_B_sfoT66hB2_0),.dout(w_dff_B_dmAlHyGz0_0),.clk(gclk));
	jdff dff_B_8Ts70Iic0_0(.din(w_dff_B_dmAlHyGz0_0),.dout(w_dff_B_8Ts70Iic0_0),.clk(gclk));
	jdff dff_B_M0RIAs7T5_0(.din(w_dff_B_8Ts70Iic0_0),.dout(w_dff_B_M0RIAs7T5_0),.clk(gclk));
	jdff dff_B_PT2aeLqK8_0(.din(w_dff_B_M0RIAs7T5_0),.dout(w_dff_B_PT2aeLqK8_0),.clk(gclk));
	jdff dff_B_iK8IYRs33_1(.din(n450),.dout(w_dff_B_iK8IYRs33_1),.clk(gclk));
	jdff dff_B_RvBrkqoy3_1(.din(w_dff_B_iK8IYRs33_1),.dout(w_dff_B_RvBrkqoy3_1),.clk(gclk));
	jdff dff_B_b93Wd1dM7_1(.din(w_dff_B_RvBrkqoy3_1),.dout(w_dff_B_b93Wd1dM7_1),.clk(gclk));
	jdff dff_B_cL4TKsTY2_1(.din(w_dff_B_b93Wd1dM7_1),.dout(w_dff_B_cL4TKsTY2_1),.clk(gclk));
	jdff dff_B_8KTSPmul4_1(.din(w_dff_B_cL4TKsTY2_1),.dout(w_dff_B_8KTSPmul4_1),.clk(gclk));
	jdff dff_B_qcBfZHT42_1(.din(w_dff_B_8KTSPmul4_1),.dout(w_dff_B_qcBfZHT42_1),.clk(gclk));
	jdff dff_B_WgmbwlWN9_1(.din(w_dff_B_qcBfZHT42_1),.dout(w_dff_B_WgmbwlWN9_1),.clk(gclk));
	jdff dff_B_hl8ngWvW5_1(.din(w_dff_B_WgmbwlWN9_1),.dout(w_dff_B_hl8ngWvW5_1),.clk(gclk));
	jdff dff_B_gP2Ricw43_1(.din(w_dff_B_hl8ngWvW5_1),.dout(w_dff_B_gP2Ricw43_1),.clk(gclk));
	jdff dff_B_FeH8ThDA8_1(.din(w_dff_B_gP2Ricw43_1),.dout(w_dff_B_FeH8ThDA8_1),.clk(gclk));
	jdff dff_B_27LeE5x30_1(.din(w_dff_B_FeH8ThDA8_1),.dout(w_dff_B_27LeE5x30_1),.clk(gclk));
	jdff dff_B_WzittY0J2_0(.din(n451),.dout(w_dff_B_WzittY0J2_0),.clk(gclk));
	jdff dff_B_digy4ypN5_0(.din(w_dff_B_WzittY0J2_0),.dout(w_dff_B_digy4ypN5_0),.clk(gclk));
	jdff dff_B_IyXXLOIo4_0(.din(w_dff_B_digy4ypN5_0),.dout(w_dff_B_IyXXLOIo4_0),.clk(gclk));
	jdff dff_B_4SFULI4g1_0(.din(w_dff_B_IyXXLOIo4_0),.dout(w_dff_B_4SFULI4g1_0),.clk(gclk));
	jdff dff_B_NHHorC111_0(.din(w_dff_B_4SFULI4g1_0),.dout(w_dff_B_NHHorC111_0),.clk(gclk));
	jdff dff_B_Qu85MC6D7_0(.din(w_dff_B_NHHorC111_0),.dout(w_dff_B_Qu85MC6D7_0),.clk(gclk));
	jdff dff_B_CWlIy23N7_0(.din(w_dff_B_Qu85MC6D7_0),.dout(w_dff_B_CWlIy23N7_0),.clk(gclk));
	jdff dff_B_FXDHyn1B9_0(.din(w_dff_B_CWlIy23N7_0),.dout(w_dff_B_FXDHyn1B9_0),.clk(gclk));
	jdff dff_B_2pvDVzF08_0(.din(w_dff_B_FXDHyn1B9_0),.dout(w_dff_B_2pvDVzF08_0),.clk(gclk));
	jdff dff_B_kd5CM0fw2_0(.din(w_dff_B_2pvDVzF08_0),.dout(w_dff_B_kd5CM0fw2_0),.clk(gclk));
	jdff dff_B_nKJsQ9ti3_0(.din(w_dff_B_kd5CM0fw2_0),.dout(w_dff_B_nKJsQ9ti3_0),.clk(gclk));
	jdff dff_B_u8Aqn7YY6_1(.din(n444),.dout(w_dff_B_u8Aqn7YY6_1),.clk(gclk));
	jdff dff_B_2fzYDzLE3_1(.din(w_dff_B_u8Aqn7YY6_1),.dout(w_dff_B_2fzYDzLE3_1),.clk(gclk));
	jdff dff_B_61jnnUxf9_1(.din(w_dff_B_2fzYDzLE3_1),.dout(w_dff_B_61jnnUxf9_1),.clk(gclk));
	jdff dff_B_XVXDV8qX3_1(.din(w_dff_B_61jnnUxf9_1),.dout(w_dff_B_XVXDV8qX3_1),.clk(gclk));
	jdff dff_B_a7TVaVEo9_1(.din(w_dff_B_XVXDV8qX3_1),.dout(w_dff_B_a7TVaVEo9_1),.clk(gclk));
	jdff dff_B_Dp5bon0S1_1(.din(w_dff_B_a7TVaVEo9_1),.dout(w_dff_B_Dp5bon0S1_1),.clk(gclk));
	jdff dff_B_ME01Jysm8_1(.din(w_dff_B_Dp5bon0S1_1),.dout(w_dff_B_ME01Jysm8_1),.clk(gclk));
	jdff dff_B_hYK1Ehqo1_1(.din(w_dff_B_ME01Jysm8_1),.dout(w_dff_B_hYK1Ehqo1_1),.clk(gclk));
	jdff dff_B_C6X7E3jq9_1(.din(w_dff_B_hYK1Ehqo1_1),.dout(w_dff_B_C6X7E3jq9_1),.clk(gclk));
	jdff dff_B_o5sfoxtN0_1(.din(w_dff_B_C6X7E3jq9_1),.dout(w_dff_B_o5sfoxtN0_1),.clk(gclk));
	jdff dff_B_2CqZQwGP3_0(.din(n445),.dout(w_dff_B_2CqZQwGP3_0),.clk(gclk));
	jdff dff_B_Xidoqr8P2_0(.din(w_dff_B_2CqZQwGP3_0),.dout(w_dff_B_Xidoqr8P2_0),.clk(gclk));
	jdff dff_B_PbfwgGb02_0(.din(w_dff_B_Xidoqr8P2_0),.dout(w_dff_B_PbfwgGb02_0),.clk(gclk));
	jdff dff_B_HzSKeLUp3_0(.din(w_dff_B_PbfwgGb02_0),.dout(w_dff_B_HzSKeLUp3_0),.clk(gclk));
	jdff dff_B_t7oo0FTl8_0(.din(w_dff_B_HzSKeLUp3_0),.dout(w_dff_B_t7oo0FTl8_0),.clk(gclk));
	jdff dff_B_k5jTnxDk4_0(.din(w_dff_B_t7oo0FTl8_0),.dout(w_dff_B_k5jTnxDk4_0),.clk(gclk));
	jdff dff_B_0NEvZZis7_0(.din(w_dff_B_k5jTnxDk4_0),.dout(w_dff_B_0NEvZZis7_0),.clk(gclk));
	jdff dff_B_1UqxfKPV0_0(.din(w_dff_B_0NEvZZis7_0),.dout(w_dff_B_1UqxfKPV0_0),.clk(gclk));
	jdff dff_B_2VgunHW36_0(.din(w_dff_B_1UqxfKPV0_0),.dout(w_dff_B_2VgunHW36_0),.clk(gclk));
	jdff dff_B_njqcx4ts3_0(.din(w_dff_B_2VgunHW36_0),.dout(w_dff_B_njqcx4ts3_0),.clk(gclk));
	jdff dff_B_WZxvvIYD2_1(.din(n438),.dout(w_dff_B_WZxvvIYD2_1),.clk(gclk));
	jdff dff_B_TSlxqhxh6_1(.din(w_dff_B_WZxvvIYD2_1),.dout(w_dff_B_TSlxqhxh6_1),.clk(gclk));
	jdff dff_B_G7hfJw6t8_1(.din(w_dff_B_TSlxqhxh6_1),.dout(w_dff_B_G7hfJw6t8_1),.clk(gclk));
	jdff dff_B_KFMw82Hu5_1(.din(w_dff_B_G7hfJw6t8_1),.dout(w_dff_B_KFMw82Hu5_1),.clk(gclk));
	jdff dff_B_mfGu0USy7_1(.din(w_dff_B_KFMw82Hu5_1),.dout(w_dff_B_mfGu0USy7_1),.clk(gclk));
	jdff dff_B_Ds146Ekz3_1(.din(w_dff_B_mfGu0USy7_1),.dout(w_dff_B_Ds146Ekz3_1),.clk(gclk));
	jdff dff_B_42Jk9NQm2_1(.din(w_dff_B_Ds146Ekz3_1),.dout(w_dff_B_42Jk9NQm2_1),.clk(gclk));
	jdff dff_B_EbeYix8q6_1(.din(w_dff_B_42Jk9NQm2_1),.dout(w_dff_B_EbeYix8q6_1),.clk(gclk));
	jdff dff_B_uSgQnbDf2_1(.din(w_dff_B_EbeYix8q6_1),.dout(w_dff_B_uSgQnbDf2_1),.clk(gclk));
	jdff dff_B_vUH7yW4f1_0(.din(n439),.dout(w_dff_B_vUH7yW4f1_0),.clk(gclk));
	jdff dff_B_YJXgnpGf7_0(.din(w_dff_B_vUH7yW4f1_0),.dout(w_dff_B_YJXgnpGf7_0),.clk(gclk));
	jdff dff_B_iBuwANGT9_0(.din(w_dff_B_YJXgnpGf7_0),.dout(w_dff_B_iBuwANGT9_0),.clk(gclk));
	jdff dff_B_UhDLPyJA2_0(.din(w_dff_B_iBuwANGT9_0),.dout(w_dff_B_UhDLPyJA2_0),.clk(gclk));
	jdff dff_B_A5abHHqR5_0(.din(w_dff_B_UhDLPyJA2_0),.dout(w_dff_B_A5abHHqR5_0),.clk(gclk));
	jdff dff_B_7S0Ebel80_0(.din(w_dff_B_A5abHHqR5_0),.dout(w_dff_B_7S0Ebel80_0),.clk(gclk));
	jdff dff_B_cIvKwSkV4_0(.din(w_dff_B_7S0Ebel80_0),.dout(w_dff_B_cIvKwSkV4_0),.clk(gclk));
	jdff dff_B_hpnBngai8_0(.din(w_dff_B_cIvKwSkV4_0),.dout(w_dff_B_hpnBngai8_0),.clk(gclk));
	jdff dff_B_oTv1F9FH9_0(.din(w_dff_B_hpnBngai8_0),.dout(w_dff_B_oTv1F9FH9_0),.clk(gclk));
	jdff dff_B_2kSTW6Sd7_1(.din(n432),.dout(w_dff_B_2kSTW6Sd7_1),.clk(gclk));
	jdff dff_B_HihNYsOz6_1(.din(w_dff_B_2kSTW6Sd7_1),.dout(w_dff_B_HihNYsOz6_1),.clk(gclk));
	jdff dff_B_rwmtQSBt7_1(.din(w_dff_B_HihNYsOz6_1),.dout(w_dff_B_rwmtQSBt7_1),.clk(gclk));
	jdff dff_B_zGrYmkmI8_1(.din(w_dff_B_rwmtQSBt7_1),.dout(w_dff_B_zGrYmkmI8_1),.clk(gclk));
	jdff dff_B_C55HPewp1_1(.din(w_dff_B_zGrYmkmI8_1),.dout(w_dff_B_C55HPewp1_1),.clk(gclk));
	jdff dff_B_ydCb9c8S3_1(.din(w_dff_B_C55HPewp1_1),.dout(w_dff_B_ydCb9c8S3_1),.clk(gclk));
	jdff dff_B_fZ9qS8y43_1(.din(w_dff_B_ydCb9c8S3_1),.dout(w_dff_B_fZ9qS8y43_1),.clk(gclk));
	jdff dff_B_N7wdEcYt6_1(.din(w_dff_B_fZ9qS8y43_1),.dout(w_dff_B_N7wdEcYt6_1),.clk(gclk));
	jdff dff_B_vKddPc6J4_0(.din(n433),.dout(w_dff_B_vKddPc6J4_0),.clk(gclk));
	jdff dff_B_SFgyGw4V0_0(.din(w_dff_B_vKddPc6J4_0),.dout(w_dff_B_SFgyGw4V0_0),.clk(gclk));
	jdff dff_B_A2G2QvTk2_0(.din(w_dff_B_SFgyGw4V0_0),.dout(w_dff_B_A2G2QvTk2_0),.clk(gclk));
	jdff dff_B_9Td78AnT3_0(.din(w_dff_B_A2G2QvTk2_0),.dout(w_dff_B_9Td78AnT3_0),.clk(gclk));
	jdff dff_B_RaHIRqRo3_0(.din(w_dff_B_9Td78AnT3_0),.dout(w_dff_B_RaHIRqRo3_0),.clk(gclk));
	jdff dff_B_kXvKi1aH9_0(.din(w_dff_B_RaHIRqRo3_0),.dout(w_dff_B_kXvKi1aH9_0),.clk(gclk));
	jdff dff_B_Jh6s40yZ9_0(.din(w_dff_B_kXvKi1aH9_0),.dout(w_dff_B_Jh6s40yZ9_0),.clk(gclk));
	jdff dff_B_mJs1Nkki5_0(.din(w_dff_B_Jh6s40yZ9_0),.dout(w_dff_B_mJs1Nkki5_0),.clk(gclk));
	jdff dff_B_OB2obTJX4_1(.din(n426),.dout(w_dff_B_OB2obTJX4_1),.clk(gclk));
	jdff dff_B_zaoNu5t89_1(.din(w_dff_B_OB2obTJX4_1),.dout(w_dff_B_zaoNu5t89_1),.clk(gclk));
	jdff dff_B_vrBd0hBk1_1(.din(w_dff_B_zaoNu5t89_1),.dout(w_dff_B_vrBd0hBk1_1),.clk(gclk));
	jdff dff_B_yJ2vPBkx1_1(.din(w_dff_B_vrBd0hBk1_1),.dout(w_dff_B_yJ2vPBkx1_1),.clk(gclk));
	jdff dff_B_qcTM0oYr3_1(.din(w_dff_B_yJ2vPBkx1_1),.dout(w_dff_B_qcTM0oYr3_1),.clk(gclk));
	jdff dff_B_hRNmHLjc4_1(.din(w_dff_B_qcTM0oYr3_1),.dout(w_dff_B_hRNmHLjc4_1),.clk(gclk));
	jdff dff_B_hLXcHmzy9_1(.din(w_dff_B_hRNmHLjc4_1),.dout(w_dff_B_hLXcHmzy9_1),.clk(gclk));
	jdff dff_B_pxoEL8Ao6_0(.din(n427),.dout(w_dff_B_pxoEL8Ao6_0),.clk(gclk));
	jdff dff_B_u7GZB3fE3_0(.din(w_dff_B_pxoEL8Ao6_0),.dout(w_dff_B_u7GZB3fE3_0),.clk(gclk));
	jdff dff_B_VAKcFD7K6_0(.din(w_dff_B_u7GZB3fE3_0),.dout(w_dff_B_VAKcFD7K6_0),.clk(gclk));
	jdff dff_B_2mjUAZxI7_0(.din(w_dff_B_VAKcFD7K6_0),.dout(w_dff_B_2mjUAZxI7_0),.clk(gclk));
	jdff dff_B_1STAXDoW0_0(.din(w_dff_B_2mjUAZxI7_0),.dout(w_dff_B_1STAXDoW0_0),.clk(gclk));
	jdff dff_B_dTc5u5NJ3_0(.din(w_dff_B_1STAXDoW0_0),.dout(w_dff_B_dTc5u5NJ3_0),.clk(gclk));
	jdff dff_B_ct1c3ZgN9_0(.din(w_dff_B_dTc5u5NJ3_0),.dout(w_dff_B_ct1c3ZgN9_0),.clk(gclk));
	jdff dff_B_CHUBRtFA7_1(.din(n420),.dout(w_dff_B_CHUBRtFA7_1),.clk(gclk));
	jdff dff_B_n0X03tB08_1(.din(w_dff_B_CHUBRtFA7_1),.dout(w_dff_B_n0X03tB08_1),.clk(gclk));
	jdff dff_B_ASNfjgOR3_1(.din(w_dff_B_n0X03tB08_1),.dout(w_dff_B_ASNfjgOR3_1),.clk(gclk));
	jdff dff_B_GHlrtJBt5_1(.din(w_dff_B_ASNfjgOR3_1),.dout(w_dff_B_GHlrtJBt5_1),.clk(gclk));
	jdff dff_B_6Ozoswgv6_1(.din(w_dff_B_GHlrtJBt5_1),.dout(w_dff_B_6Ozoswgv6_1),.clk(gclk));
	jdff dff_B_7AXejlE29_1(.din(w_dff_B_6Ozoswgv6_1),.dout(w_dff_B_7AXejlE29_1),.clk(gclk));
	jdff dff_B_OW2MPfgS2_0(.din(n421),.dout(w_dff_B_OW2MPfgS2_0),.clk(gclk));
	jdff dff_B_8V7YNLIH4_0(.din(w_dff_B_OW2MPfgS2_0),.dout(w_dff_B_8V7YNLIH4_0),.clk(gclk));
	jdff dff_B_xLIWOsd62_0(.din(w_dff_B_8V7YNLIH4_0),.dout(w_dff_B_xLIWOsd62_0),.clk(gclk));
	jdff dff_B_pLV3pkIm4_0(.din(w_dff_B_xLIWOsd62_0),.dout(w_dff_B_pLV3pkIm4_0),.clk(gclk));
	jdff dff_B_BxtlValQ7_0(.din(w_dff_B_pLV3pkIm4_0),.dout(w_dff_B_BxtlValQ7_0),.clk(gclk));
	jdff dff_B_jwfquIHg2_0(.din(w_dff_B_BxtlValQ7_0),.dout(w_dff_B_jwfquIHg2_0),.clk(gclk));
	jdff dff_B_HuqhDjQS5_1(.din(n414),.dout(w_dff_B_HuqhDjQS5_1),.clk(gclk));
	jdff dff_B_IE6E3WZZ4_1(.din(w_dff_B_HuqhDjQS5_1),.dout(w_dff_B_IE6E3WZZ4_1),.clk(gclk));
	jdff dff_B_sMlnHecV2_1(.din(w_dff_B_IE6E3WZZ4_1),.dout(w_dff_B_sMlnHecV2_1),.clk(gclk));
	jdff dff_B_3RzBsZo46_1(.din(w_dff_B_sMlnHecV2_1),.dout(w_dff_B_3RzBsZo46_1),.clk(gclk));
	jdff dff_B_IAJMsY3O3_1(.din(w_dff_B_3RzBsZo46_1),.dout(w_dff_B_IAJMsY3O3_1),.clk(gclk));
	jdff dff_B_1XUtnL036_0(.din(n415),.dout(w_dff_B_1XUtnL036_0),.clk(gclk));
	jdff dff_B_dumKUOU95_0(.din(w_dff_B_1XUtnL036_0),.dout(w_dff_B_dumKUOU95_0),.clk(gclk));
	jdff dff_B_IhzeJ2iA2_0(.din(w_dff_B_dumKUOU95_0),.dout(w_dff_B_IhzeJ2iA2_0),.clk(gclk));
	jdff dff_B_6HLLPz0U0_0(.din(w_dff_B_IhzeJ2iA2_0),.dout(w_dff_B_6HLLPz0U0_0),.clk(gclk));
	jdff dff_B_D2KL4nNr1_0(.din(w_dff_B_6HLLPz0U0_0),.dout(w_dff_B_D2KL4nNr1_0),.clk(gclk));
	jdff dff_B_91yUkRCn4_1(.din(n408),.dout(w_dff_B_91yUkRCn4_1),.clk(gclk));
	jdff dff_B_fO5HpThl3_1(.din(w_dff_B_91yUkRCn4_1),.dout(w_dff_B_fO5HpThl3_1),.clk(gclk));
	jdff dff_B_nHghsEwQ6_1(.din(w_dff_B_fO5HpThl3_1),.dout(w_dff_B_nHghsEwQ6_1),.clk(gclk));
	jdff dff_B_9DVgFh9T1_1(.din(w_dff_B_nHghsEwQ6_1),.dout(w_dff_B_9DVgFh9T1_1),.clk(gclk));
	jdff dff_B_DBi1JzBL5_0(.din(n409),.dout(w_dff_B_DBi1JzBL5_0),.clk(gclk));
	jdff dff_B_OSgiaOyx3_0(.din(w_dff_B_DBi1JzBL5_0),.dout(w_dff_B_OSgiaOyx3_0),.clk(gclk));
	jdff dff_B_jpsm4AHP2_0(.din(w_dff_B_OSgiaOyx3_0),.dout(w_dff_B_jpsm4AHP2_0),.clk(gclk));
	jdff dff_B_NsJlHOhQ0_0(.din(w_dff_B_jpsm4AHP2_0),.dout(w_dff_B_NsJlHOhQ0_0),.clk(gclk));
	jdff dff_B_rrHAuH711_1(.din(n402),.dout(w_dff_B_rrHAuH711_1),.clk(gclk));
	jdff dff_B_AAX4DMaO0_1(.din(w_dff_B_rrHAuH711_1),.dout(w_dff_B_AAX4DMaO0_1),.clk(gclk));
	jdff dff_B_RYyduIeI2_1(.din(w_dff_B_AAX4DMaO0_1),.dout(w_dff_B_RYyduIeI2_1),.clk(gclk));
	jdff dff_B_U5MNQmS86_0(.din(n403),.dout(w_dff_B_U5MNQmS86_0),.clk(gclk));
	jdff dff_B_6rt9170L4_0(.din(w_dff_B_U5MNQmS86_0),.dout(w_dff_B_6rt9170L4_0),.clk(gclk));
	jdff dff_B_tOSk0HiB9_0(.din(w_dff_B_6rt9170L4_0),.dout(w_dff_B_tOSk0HiB9_0),.clk(gclk));
	jdff dff_B_q4293DRu4_1(.din(n396),.dout(w_dff_B_q4293DRu4_1),.clk(gclk));
	jdff dff_B_XC6XIR9e5_1(.din(w_dff_B_q4293DRu4_1),.dout(w_dff_B_XC6XIR9e5_1),.clk(gclk));
	jdff dff_B_yaQER63f8_0(.din(n397),.dout(w_dff_B_yaQER63f8_0),.clk(gclk));
	jdff dff_B_MevlBocM3_0(.din(w_dff_B_yaQER63f8_0),.dout(w_dff_B_MevlBocM3_0),.clk(gclk));
	jdff dff_B_bq66TJJL2_1(.din(n390),.dout(w_dff_B_bq66TJJL2_1),.clk(gclk));
	jdff dff_B_7v1bBDjM8_0(.din(n391),.dout(w_dff_B_7v1bBDjM8_0),.clk(gclk));
	jdff dff_A_i0Y4neCV3_2(.dout(w_dff_A_j9T031q05_0),.din(w_dff_A_i0Y4neCV3_2),.clk(gclk));
	jdff dff_A_j9T031q05_0(.dout(w_dff_A_vOiNMKYP3_0),.din(w_dff_A_j9T031q05_0),.clk(gclk));
	jdff dff_A_vOiNMKYP3_0(.dout(w_dff_A_g7jlr3ng4_0),.din(w_dff_A_vOiNMKYP3_0),.clk(gclk));
	jdff dff_A_g7jlr3ng4_0(.dout(w_dff_A_7xO2jXg01_0),.din(w_dff_A_g7jlr3ng4_0),.clk(gclk));
	jdff dff_A_7xO2jXg01_0(.dout(w_dff_A_iMKXw20r6_0),.din(w_dff_A_7xO2jXg01_0),.clk(gclk));
	jdff dff_A_iMKXw20r6_0(.dout(w_dff_A_MsCrJjMJ8_0),.din(w_dff_A_iMKXw20r6_0),.clk(gclk));
	jdff dff_A_MsCrJjMJ8_0(.dout(w_dff_A_4vHSuZu70_0),.din(w_dff_A_MsCrJjMJ8_0),.clk(gclk));
	jdff dff_A_4vHSuZu70_0(.dout(w_dff_A_WjGq4SrP5_0),.din(w_dff_A_4vHSuZu70_0),.clk(gclk));
	jdff dff_A_WjGq4SrP5_0(.dout(w_dff_A_UD7Fx71E9_0),.din(w_dff_A_WjGq4SrP5_0),.clk(gclk));
	jdff dff_A_UD7Fx71E9_0(.dout(w_dff_A_BlG5FfJJ3_0),.din(w_dff_A_UD7Fx71E9_0),.clk(gclk));
	jdff dff_A_BlG5FfJJ3_0(.dout(w_dff_A_u78ECBzG5_0),.din(w_dff_A_BlG5FfJJ3_0),.clk(gclk));
	jdff dff_A_u78ECBzG5_0(.dout(w_dff_A_IjlLUlhH9_0),.din(w_dff_A_u78ECBzG5_0),.clk(gclk));
	jdff dff_A_IjlLUlhH9_0(.dout(w_dff_A_DeVWj5dN4_0),.din(w_dff_A_IjlLUlhH9_0),.clk(gclk));
	jdff dff_A_DeVWj5dN4_0(.dout(w_dff_A_NGHM5wy50_0),.din(w_dff_A_DeVWj5dN4_0),.clk(gclk));
	jdff dff_A_NGHM5wy50_0(.dout(w_dff_A_fmaRaMD69_0),.din(w_dff_A_NGHM5wy50_0),.clk(gclk));
	jdff dff_A_fmaRaMD69_0(.dout(w_dff_A_1QE0PPCo6_0),.din(w_dff_A_fmaRaMD69_0),.clk(gclk));
	jdff dff_A_1QE0PPCo6_0(.dout(w_dff_A_MtM8rSW48_0),.din(w_dff_A_1QE0PPCo6_0),.clk(gclk));
	jdff dff_A_MtM8rSW48_0(.dout(w_dff_A_FVQJGeqJ3_0),.din(w_dff_A_MtM8rSW48_0),.clk(gclk));
	jdff dff_A_FVQJGeqJ3_0(.dout(w_dff_A_qyRq3uJQ5_0),.din(w_dff_A_FVQJGeqJ3_0),.clk(gclk));
	jdff dff_A_qyRq3uJQ5_0(.dout(w_dff_A_3jDPCLoI8_0),.din(w_dff_A_qyRq3uJQ5_0),.clk(gclk));
	jdff dff_A_3jDPCLoI8_0(.dout(w_dff_A_1hGM26PS8_0),.din(w_dff_A_3jDPCLoI8_0),.clk(gclk));
	jdff dff_A_1hGM26PS8_0(.dout(w_dff_A_BsNAX5yA1_0),.din(w_dff_A_1hGM26PS8_0),.clk(gclk));
	jdff dff_A_BsNAX5yA1_0(.dout(w_dff_A_BbLFrTpV2_0),.din(w_dff_A_BsNAX5yA1_0),.clk(gclk));
	jdff dff_A_BbLFrTpV2_0(.dout(w_dff_A_Br5jEmCl2_0),.din(w_dff_A_BbLFrTpV2_0),.clk(gclk));
	jdff dff_A_Br5jEmCl2_0(.dout(w_dff_A_5cjTzbmW6_0),.din(w_dff_A_Br5jEmCl2_0),.clk(gclk));
	jdff dff_A_5cjTzbmW6_0(.dout(w_dff_A_Q4HY9n4w0_0),.din(w_dff_A_5cjTzbmW6_0),.clk(gclk));
	jdff dff_A_Q4HY9n4w0_0(.dout(w_dff_A_KSDQi7Sr8_0),.din(w_dff_A_Q4HY9n4w0_0),.clk(gclk));
	jdff dff_A_KSDQi7Sr8_0(.dout(w_dff_A_9Esn0sSu7_0),.din(w_dff_A_KSDQi7Sr8_0),.clk(gclk));
	jdff dff_A_9Esn0sSu7_0(.dout(w_dff_A_NYjX1kI69_0),.din(w_dff_A_9Esn0sSu7_0),.clk(gclk));
	jdff dff_A_NYjX1kI69_0(.dout(w_dff_A_PAv4FYSN4_0),.din(w_dff_A_NYjX1kI69_0),.clk(gclk));
	jdff dff_A_PAv4FYSN4_0(.dout(w_dff_A_fZbm0Pb18_0),.din(w_dff_A_PAv4FYSN4_0),.clk(gclk));
	jdff dff_A_fZbm0Pb18_0(.dout(w_dff_A_CpTsBUrx7_0),.din(w_dff_A_fZbm0Pb18_0),.clk(gclk));
	jdff dff_A_CpTsBUrx7_0(.dout(w_dff_A_wpibraiv9_0),.din(w_dff_A_CpTsBUrx7_0),.clk(gclk));
	jdff dff_A_wpibraiv9_0(.dout(w_dff_A_YECaqBxJ3_0),.din(w_dff_A_wpibraiv9_0),.clk(gclk));
	jdff dff_A_YECaqBxJ3_0(.dout(w_dff_A_YvPcmbAA1_0),.din(w_dff_A_YECaqBxJ3_0),.clk(gclk));
	jdff dff_A_YvPcmbAA1_0(.dout(w_dff_A_h1bwGIX91_0),.din(w_dff_A_YvPcmbAA1_0),.clk(gclk));
	jdff dff_A_h1bwGIX91_0(.dout(w_dff_A_mytFLC8s0_0),.din(w_dff_A_h1bwGIX91_0),.clk(gclk));
	jdff dff_A_mytFLC8s0_0(.dout(w_dff_A_ChQHW2bi6_0),.din(w_dff_A_mytFLC8s0_0),.clk(gclk));
	jdff dff_A_ChQHW2bi6_0(.dout(w_dff_A_Bfpumz2I0_0),.din(w_dff_A_ChQHW2bi6_0),.clk(gclk));
	jdff dff_A_Bfpumz2I0_0(.dout(w_dff_A_AQlr7wG59_0),.din(w_dff_A_Bfpumz2I0_0),.clk(gclk));
	jdff dff_A_AQlr7wG59_0(.dout(w_dff_A_p3fLkJ6r9_0),.din(w_dff_A_AQlr7wG59_0),.clk(gclk));
	jdff dff_A_p3fLkJ6r9_0(.dout(w_dff_A_FfFHmd7v3_0),.din(w_dff_A_p3fLkJ6r9_0),.clk(gclk));
	jdff dff_A_FfFHmd7v3_0(.dout(w_dff_A_a5Oc9kr70_0),.din(w_dff_A_FfFHmd7v3_0),.clk(gclk));
	jdff dff_A_a5Oc9kr70_0(.dout(w_dff_A_Ra95uvKl2_0),.din(w_dff_A_a5Oc9kr70_0),.clk(gclk));
	jdff dff_A_Ra95uvKl2_0(.dout(w_dff_A_wQ78edMl3_0),.din(w_dff_A_Ra95uvKl2_0),.clk(gclk));
	jdff dff_A_wQ78edMl3_0(.dout(w_dff_A_lNWXIFlC6_0),.din(w_dff_A_wQ78edMl3_0),.clk(gclk));
	jdff dff_A_lNWXIFlC6_0(.dout(w_dff_A_EQajtwzB7_0),.din(w_dff_A_lNWXIFlC6_0),.clk(gclk));
	jdff dff_A_EQajtwzB7_0(.dout(w_dff_A_nS0N2j9E4_0),.din(w_dff_A_EQajtwzB7_0),.clk(gclk));
	jdff dff_A_nS0N2j9E4_0(.dout(w_dff_A_F7vrl6TH5_0),.din(w_dff_A_nS0N2j9E4_0),.clk(gclk));
	jdff dff_A_F7vrl6TH5_0(.dout(w_dff_A_F82sm3Qg5_0),.din(w_dff_A_F7vrl6TH5_0),.clk(gclk));
	jdff dff_A_F82sm3Qg5_0(.dout(w_dff_A_DWlzNtNs3_0),.din(w_dff_A_F82sm3Qg5_0),.clk(gclk));
	jdff dff_A_DWlzNtNs3_0(.dout(w_dff_A_lzKWaH0E2_0),.din(w_dff_A_DWlzNtNs3_0),.clk(gclk));
	jdff dff_A_lzKWaH0E2_0(.dout(w_dff_A_MdGhRnUY2_0),.din(w_dff_A_lzKWaH0E2_0),.clk(gclk));
	jdff dff_A_MdGhRnUY2_0(.dout(w_dff_A_QwkWUQC88_0),.din(w_dff_A_MdGhRnUY2_0),.clk(gclk));
	jdff dff_A_QwkWUQC88_0(.dout(w_dff_A_s16Kjcf04_0),.din(w_dff_A_QwkWUQC88_0),.clk(gclk));
	jdff dff_A_s16Kjcf04_0(.dout(w_dff_A_8C1R7pBF0_0),.din(w_dff_A_s16Kjcf04_0),.clk(gclk));
	jdff dff_A_8C1R7pBF0_0(.dout(w_dff_A_A698ntck9_0),.din(w_dff_A_8C1R7pBF0_0),.clk(gclk));
	jdff dff_A_A698ntck9_0(.dout(w_dff_A_XMpNqoHx8_0),.din(w_dff_A_A698ntck9_0),.clk(gclk));
	jdff dff_A_XMpNqoHx8_0(.dout(w_dff_A_mbphToWb7_0),.din(w_dff_A_XMpNqoHx8_0),.clk(gclk));
	jdff dff_A_mbphToWb7_0(.dout(w_dff_A_h8kgWcfH2_0),.din(w_dff_A_mbphToWb7_0),.clk(gclk));
	jdff dff_A_h8kgWcfH2_0(.dout(w_dff_A_wdiR9ZbH8_0),.din(w_dff_A_h8kgWcfH2_0),.clk(gclk));
	jdff dff_A_wdiR9ZbH8_0(.dout(w_dff_A_9aXA21gj8_0),.din(w_dff_A_wdiR9ZbH8_0),.clk(gclk));
	jdff dff_A_9aXA21gj8_0(.dout(w_dff_A_dllhdTsZ5_0),.din(w_dff_A_9aXA21gj8_0),.clk(gclk));
	jdff dff_A_dllhdTsZ5_0(.dout(w_dff_A_hkntw2iQ3_0),.din(w_dff_A_dllhdTsZ5_0),.clk(gclk));
	jdff dff_A_hkntw2iQ3_0(.dout(w_dff_A_F2R2oWU87_0),.din(w_dff_A_hkntw2iQ3_0),.clk(gclk));
	jdff dff_A_F2R2oWU87_0(.dout(w_dff_A_Yz94n4vv2_0),.din(w_dff_A_F2R2oWU87_0),.clk(gclk));
	jdff dff_A_Yz94n4vv2_0(.dout(w_dff_A_mW3QoIE34_0),.din(w_dff_A_Yz94n4vv2_0),.clk(gclk));
	jdff dff_A_mW3QoIE34_0(.dout(w_dff_A_p0NmxDOf5_0),.din(w_dff_A_mW3QoIE34_0),.clk(gclk));
	jdff dff_A_p0NmxDOf5_0(.dout(w_dff_A_hAjsqHFs7_0),.din(w_dff_A_p0NmxDOf5_0),.clk(gclk));
	jdff dff_A_hAjsqHFs7_0(.dout(w_dff_A_XSuWdF6A5_0),.din(w_dff_A_hAjsqHFs7_0),.clk(gclk));
	jdff dff_A_XSuWdF6A5_0(.dout(w_dff_A_oU0ETh9J1_0),.din(w_dff_A_XSuWdF6A5_0),.clk(gclk));
	jdff dff_A_oU0ETh9J1_0(.dout(w_dff_A_b8zCdsUw4_0),.din(w_dff_A_oU0ETh9J1_0),.clk(gclk));
	jdff dff_A_b8zCdsUw4_0(.dout(w_dff_A_tNUiQJeN7_0),.din(w_dff_A_b8zCdsUw4_0),.clk(gclk));
	jdff dff_A_tNUiQJeN7_0(.dout(w_dff_A_sBerItzw4_0),.din(w_dff_A_tNUiQJeN7_0),.clk(gclk));
	jdff dff_A_sBerItzw4_0(.dout(w_dff_A_Ck24AXEd6_0),.din(w_dff_A_sBerItzw4_0),.clk(gclk));
	jdff dff_A_Ck24AXEd6_0(.dout(w_dff_A_zLwlimAo0_0),.din(w_dff_A_Ck24AXEd6_0),.clk(gclk));
	jdff dff_A_zLwlimAo0_0(.dout(w_dff_A_q7N8tmnv2_0),.din(w_dff_A_zLwlimAo0_0),.clk(gclk));
	jdff dff_A_q7N8tmnv2_0(.dout(w_dff_A_s07mlbpA8_0),.din(w_dff_A_q7N8tmnv2_0),.clk(gclk));
	jdff dff_A_s07mlbpA8_0(.dout(w_dff_A_xN753xVm5_0),.din(w_dff_A_s07mlbpA8_0),.clk(gclk));
	jdff dff_A_xN753xVm5_0(.dout(w_dff_A_ltBC9pjb9_0),.din(w_dff_A_xN753xVm5_0),.clk(gclk));
	jdff dff_A_ltBC9pjb9_0(.dout(w_dff_A_rsthNRDN8_0),.din(w_dff_A_ltBC9pjb9_0),.clk(gclk));
	jdff dff_A_rsthNRDN8_0(.dout(w_dff_A_6VmHlJVB6_0),.din(w_dff_A_rsthNRDN8_0),.clk(gclk));
	jdff dff_A_6VmHlJVB6_0(.dout(w_dff_A_Rd7ZK2f16_0),.din(w_dff_A_6VmHlJVB6_0),.clk(gclk));
	jdff dff_A_Rd7ZK2f16_0(.dout(w_dff_A_MhIDTrRH2_0),.din(w_dff_A_Rd7ZK2f16_0),.clk(gclk));
	jdff dff_A_MhIDTrRH2_0(.dout(w_dff_A_2084AwKm7_0),.din(w_dff_A_MhIDTrRH2_0),.clk(gclk));
	jdff dff_A_2084AwKm7_0(.dout(w_dff_A_dyLYxj1m9_0),.din(w_dff_A_2084AwKm7_0),.clk(gclk));
	jdff dff_A_dyLYxj1m9_0(.dout(w_dff_A_r76cTSru5_0),.din(w_dff_A_dyLYxj1m9_0),.clk(gclk));
	jdff dff_A_r76cTSru5_0(.dout(w_dff_A_9upUtRfy7_0),.din(w_dff_A_r76cTSru5_0),.clk(gclk));
	jdff dff_A_9upUtRfy7_0(.dout(w_dff_A_R3GFswzi0_0),.din(w_dff_A_9upUtRfy7_0),.clk(gclk));
	jdff dff_A_R3GFswzi0_0(.dout(w_dff_A_qDpZEltD3_0),.din(w_dff_A_R3GFswzi0_0),.clk(gclk));
	jdff dff_A_qDpZEltD3_0(.dout(w_dff_A_tQ21VjHR8_0),.din(w_dff_A_qDpZEltD3_0),.clk(gclk));
	jdff dff_A_tQ21VjHR8_0(.dout(w_dff_A_APJkiJjk3_0),.din(w_dff_A_tQ21VjHR8_0),.clk(gclk));
	jdff dff_A_APJkiJjk3_0(.dout(w_dff_A_f0jsEngB0_0),.din(w_dff_A_APJkiJjk3_0),.clk(gclk));
	jdff dff_A_f0jsEngB0_0(.dout(w_dff_A_bj5kxm8C9_0),.din(w_dff_A_f0jsEngB0_0),.clk(gclk));
	jdff dff_A_bj5kxm8C9_0(.dout(w_dff_A_892gOQmY8_0),.din(w_dff_A_bj5kxm8C9_0),.clk(gclk));
	jdff dff_A_892gOQmY8_0(.dout(w_dff_A_CXFTnmf38_0),.din(w_dff_A_892gOQmY8_0),.clk(gclk));
	jdff dff_A_CXFTnmf38_0(.dout(w_dff_A_n5VIXJVX0_0),.din(w_dff_A_CXFTnmf38_0),.clk(gclk));
	jdff dff_A_n5VIXJVX0_0(.dout(w_dff_A_OvUzNb0a9_0),.din(w_dff_A_n5VIXJVX0_0),.clk(gclk));
	jdff dff_A_OvUzNb0a9_0(.dout(w_dff_A_3T7R4z2L7_0),.din(w_dff_A_OvUzNb0a9_0),.clk(gclk));
	jdff dff_A_3T7R4z2L7_0(.dout(w_dff_A_6hVGcGjn7_0),.din(w_dff_A_3T7R4z2L7_0),.clk(gclk));
	jdff dff_A_6hVGcGjn7_0(.dout(w_dff_A_1bs2MkNT3_0),.din(w_dff_A_6hVGcGjn7_0),.clk(gclk));
	jdff dff_A_1bs2MkNT3_0(.dout(w_dff_A_hq1hQlX82_0),.din(w_dff_A_1bs2MkNT3_0),.clk(gclk));
	jdff dff_A_hq1hQlX82_0(.dout(w_dff_A_K6RhxdqK9_0),.din(w_dff_A_hq1hQlX82_0),.clk(gclk));
	jdff dff_A_K6RhxdqK9_0(.dout(w_dff_A_lB4foRKx4_0),.din(w_dff_A_K6RhxdqK9_0),.clk(gclk));
	jdff dff_A_lB4foRKx4_0(.dout(w_dff_A_SyYyACrh3_0),.din(w_dff_A_lB4foRKx4_0),.clk(gclk));
	jdff dff_A_SyYyACrh3_0(.dout(w_dff_A_vrg7IbP29_0),.din(w_dff_A_SyYyACrh3_0),.clk(gclk));
	jdff dff_A_vrg7IbP29_0(.dout(w_dff_A_hw9WaR1E0_0),.din(w_dff_A_vrg7IbP29_0),.clk(gclk));
	jdff dff_A_hw9WaR1E0_0(.dout(w_dff_A_FnaEgvJL6_0),.din(w_dff_A_hw9WaR1E0_0),.clk(gclk));
	jdff dff_A_FnaEgvJL6_0(.dout(w_dff_A_L5GZFCwL1_0),.din(w_dff_A_FnaEgvJL6_0),.clk(gclk));
	jdff dff_A_L5GZFCwL1_0(.dout(w_dff_A_7Ge97Kqv7_0),.din(w_dff_A_L5GZFCwL1_0),.clk(gclk));
	jdff dff_A_7Ge97Kqv7_0(.dout(w_dff_A_5dlhIaId4_0),.din(w_dff_A_7Ge97Kqv7_0),.clk(gclk));
	jdff dff_A_5dlhIaId4_0(.dout(w_dff_A_kAsFlyjP4_0),.din(w_dff_A_5dlhIaId4_0),.clk(gclk));
	jdff dff_A_kAsFlyjP4_0(.dout(w_dff_A_TzGzpJ4C3_0),.din(w_dff_A_kAsFlyjP4_0),.clk(gclk));
	jdff dff_A_TzGzpJ4C3_0(.dout(w_dff_A_a3hY8lG88_0),.din(w_dff_A_TzGzpJ4C3_0),.clk(gclk));
	jdff dff_A_a3hY8lG88_0(.dout(w_dff_A_TtW8gwUa3_0),.din(w_dff_A_a3hY8lG88_0),.clk(gclk));
	jdff dff_A_TtW8gwUa3_0(.dout(w_dff_A_jJJCywzm0_0),.din(w_dff_A_TtW8gwUa3_0),.clk(gclk));
	jdff dff_A_jJJCywzm0_0(.dout(w_dff_A_3anXx5NG1_0),.din(w_dff_A_jJJCywzm0_0),.clk(gclk));
	jdff dff_A_3anXx5NG1_0(.dout(w_dff_A_LsjfsP1Y6_0),.din(w_dff_A_3anXx5NG1_0),.clk(gclk));
	jdff dff_A_LsjfsP1Y6_0(.dout(w_dff_A_crqbojAo4_0),.din(w_dff_A_LsjfsP1Y6_0),.clk(gclk));
	jdff dff_A_crqbojAo4_0(.dout(w_dff_A_jC9vxI7n8_0),.din(w_dff_A_crqbojAo4_0),.clk(gclk));
	jdff dff_A_jC9vxI7n8_0(.dout(w_dff_A_xxv6f08e9_0),.din(w_dff_A_jC9vxI7n8_0),.clk(gclk));
	jdff dff_A_xxv6f08e9_0(.dout(w_dff_A_IVoLt4XJ3_0),.din(w_dff_A_xxv6f08e9_0),.clk(gclk));
	jdff dff_A_IVoLt4XJ3_0(.dout(w_dff_A_vf1lBtKz5_0),.din(w_dff_A_IVoLt4XJ3_0),.clk(gclk));
	jdff dff_A_vf1lBtKz5_0(.dout(w_dff_A_jWt7kMj01_0),.din(w_dff_A_vf1lBtKz5_0),.clk(gclk));
	jdff dff_A_jWt7kMj01_0(.dout(w_dff_A_LsCziHwc8_0),.din(w_dff_A_jWt7kMj01_0),.clk(gclk));
	jdff dff_A_LsCziHwc8_0(.dout(w_dff_A_dYHDCUxr5_0),.din(w_dff_A_LsCziHwc8_0),.clk(gclk));
	jdff dff_A_dYHDCUxr5_0(.dout(f0),.din(w_dff_A_dYHDCUxr5_0),.clk(gclk));
	jdff dff_A_0HyOVMXh8_2(.dout(w_dff_A_3G23CtSw0_0),.din(w_dff_A_0HyOVMXh8_2),.clk(gclk));
	jdff dff_A_3G23CtSw0_0(.dout(w_dff_A_0nIw1xIb5_0),.din(w_dff_A_3G23CtSw0_0),.clk(gclk));
	jdff dff_A_0nIw1xIb5_0(.dout(w_dff_A_QYm95bez2_0),.din(w_dff_A_0nIw1xIb5_0),.clk(gclk));
	jdff dff_A_QYm95bez2_0(.dout(w_dff_A_own2PeE63_0),.din(w_dff_A_QYm95bez2_0),.clk(gclk));
	jdff dff_A_own2PeE63_0(.dout(w_dff_A_PnCakQKp7_0),.din(w_dff_A_own2PeE63_0),.clk(gclk));
	jdff dff_A_PnCakQKp7_0(.dout(w_dff_A_95eyG7NE0_0),.din(w_dff_A_PnCakQKp7_0),.clk(gclk));
	jdff dff_A_95eyG7NE0_0(.dout(w_dff_A_j6fh7tBp4_0),.din(w_dff_A_95eyG7NE0_0),.clk(gclk));
	jdff dff_A_j6fh7tBp4_0(.dout(w_dff_A_dCXANpXg1_0),.din(w_dff_A_j6fh7tBp4_0),.clk(gclk));
	jdff dff_A_dCXANpXg1_0(.dout(w_dff_A_6RytlC7I6_0),.din(w_dff_A_dCXANpXg1_0),.clk(gclk));
	jdff dff_A_6RytlC7I6_0(.dout(w_dff_A_Ai7zWDjI4_0),.din(w_dff_A_6RytlC7I6_0),.clk(gclk));
	jdff dff_A_Ai7zWDjI4_0(.dout(w_dff_A_dssNx9xZ2_0),.din(w_dff_A_Ai7zWDjI4_0),.clk(gclk));
	jdff dff_A_dssNx9xZ2_0(.dout(w_dff_A_X5qBjmyC9_0),.din(w_dff_A_dssNx9xZ2_0),.clk(gclk));
	jdff dff_A_X5qBjmyC9_0(.dout(w_dff_A_dXWKlv5p2_0),.din(w_dff_A_X5qBjmyC9_0),.clk(gclk));
	jdff dff_A_dXWKlv5p2_0(.dout(w_dff_A_caK9uQfT4_0),.din(w_dff_A_dXWKlv5p2_0),.clk(gclk));
	jdff dff_A_caK9uQfT4_0(.dout(w_dff_A_WgiQCrIh1_0),.din(w_dff_A_caK9uQfT4_0),.clk(gclk));
	jdff dff_A_WgiQCrIh1_0(.dout(w_dff_A_H2n7MluO8_0),.din(w_dff_A_WgiQCrIh1_0),.clk(gclk));
	jdff dff_A_H2n7MluO8_0(.dout(w_dff_A_lzT9a55J2_0),.din(w_dff_A_H2n7MluO8_0),.clk(gclk));
	jdff dff_A_lzT9a55J2_0(.dout(w_dff_A_ru8uTTJN4_0),.din(w_dff_A_lzT9a55J2_0),.clk(gclk));
	jdff dff_A_ru8uTTJN4_0(.dout(w_dff_A_8iTMwZxx2_0),.din(w_dff_A_ru8uTTJN4_0),.clk(gclk));
	jdff dff_A_8iTMwZxx2_0(.dout(w_dff_A_vclqBMNU4_0),.din(w_dff_A_8iTMwZxx2_0),.clk(gclk));
	jdff dff_A_vclqBMNU4_0(.dout(w_dff_A_u65A8I2k2_0),.din(w_dff_A_vclqBMNU4_0),.clk(gclk));
	jdff dff_A_u65A8I2k2_0(.dout(w_dff_A_40WVdttX2_0),.din(w_dff_A_u65A8I2k2_0),.clk(gclk));
	jdff dff_A_40WVdttX2_0(.dout(w_dff_A_vX7CEtcz9_0),.din(w_dff_A_40WVdttX2_0),.clk(gclk));
	jdff dff_A_vX7CEtcz9_0(.dout(w_dff_A_Sz6NsqZl6_0),.din(w_dff_A_vX7CEtcz9_0),.clk(gclk));
	jdff dff_A_Sz6NsqZl6_0(.dout(w_dff_A_JBr9KMOI3_0),.din(w_dff_A_Sz6NsqZl6_0),.clk(gclk));
	jdff dff_A_JBr9KMOI3_0(.dout(w_dff_A_O0W1wJmi4_0),.din(w_dff_A_JBr9KMOI3_0),.clk(gclk));
	jdff dff_A_O0W1wJmi4_0(.dout(w_dff_A_chSHBBma5_0),.din(w_dff_A_O0W1wJmi4_0),.clk(gclk));
	jdff dff_A_chSHBBma5_0(.dout(w_dff_A_tNvW27wX0_0),.din(w_dff_A_chSHBBma5_0),.clk(gclk));
	jdff dff_A_tNvW27wX0_0(.dout(w_dff_A_vL2PBhjs8_0),.din(w_dff_A_tNvW27wX0_0),.clk(gclk));
	jdff dff_A_vL2PBhjs8_0(.dout(w_dff_A_Li7ZzbTp0_0),.din(w_dff_A_vL2PBhjs8_0),.clk(gclk));
	jdff dff_A_Li7ZzbTp0_0(.dout(w_dff_A_CRD7aBrp1_0),.din(w_dff_A_Li7ZzbTp0_0),.clk(gclk));
	jdff dff_A_CRD7aBrp1_0(.dout(w_dff_A_85BVUYDg4_0),.din(w_dff_A_CRD7aBrp1_0),.clk(gclk));
	jdff dff_A_85BVUYDg4_0(.dout(w_dff_A_Ur617CXp1_0),.din(w_dff_A_85BVUYDg4_0),.clk(gclk));
	jdff dff_A_Ur617CXp1_0(.dout(w_dff_A_xR42W3dx1_0),.din(w_dff_A_Ur617CXp1_0),.clk(gclk));
	jdff dff_A_xR42W3dx1_0(.dout(w_dff_A_MUBBZAyu8_0),.din(w_dff_A_xR42W3dx1_0),.clk(gclk));
	jdff dff_A_MUBBZAyu8_0(.dout(w_dff_A_0IqHmckP5_0),.din(w_dff_A_MUBBZAyu8_0),.clk(gclk));
	jdff dff_A_0IqHmckP5_0(.dout(w_dff_A_mtVZU8B56_0),.din(w_dff_A_0IqHmckP5_0),.clk(gclk));
	jdff dff_A_mtVZU8B56_0(.dout(w_dff_A_yHrDEpg68_0),.din(w_dff_A_mtVZU8B56_0),.clk(gclk));
	jdff dff_A_yHrDEpg68_0(.dout(w_dff_A_1ED0imto9_0),.din(w_dff_A_yHrDEpg68_0),.clk(gclk));
	jdff dff_A_1ED0imto9_0(.dout(w_dff_A_nNi07eYW2_0),.din(w_dff_A_1ED0imto9_0),.clk(gclk));
	jdff dff_A_nNi07eYW2_0(.dout(w_dff_A_4Nomh9bM3_0),.din(w_dff_A_nNi07eYW2_0),.clk(gclk));
	jdff dff_A_4Nomh9bM3_0(.dout(w_dff_A_SQNXA9Wl9_0),.din(w_dff_A_4Nomh9bM3_0),.clk(gclk));
	jdff dff_A_SQNXA9Wl9_0(.dout(w_dff_A_irmpFzn86_0),.din(w_dff_A_SQNXA9Wl9_0),.clk(gclk));
	jdff dff_A_irmpFzn86_0(.dout(w_dff_A_WcITGojs6_0),.din(w_dff_A_irmpFzn86_0),.clk(gclk));
	jdff dff_A_WcITGojs6_0(.dout(w_dff_A_5CVuS75m4_0),.din(w_dff_A_WcITGojs6_0),.clk(gclk));
	jdff dff_A_5CVuS75m4_0(.dout(w_dff_A_xgR6y6b96_0),.din(w_dff_A_5CVuS75m4_0),.clk(gclk));
	jdff dff_A_xgR6y6b96_0(.dout(w_dff_A_UMmVYahG3_0),.din(w_dff_A_xgR6y6b96_0),.clk(gclk));
	jdff dff_A_UMmVYahG3_0(.dout(w_dff_A_t58Ms7ZG9_0),.din(w_dff_A_UMmVYahG3_0),.clk(gclk));
	jdff dff_A_t58Ms7ZG9_0(.dout(w_dff_A_9JTQdnKu9_0),.din(w_dff_A_t58Ms7ZG9_0),.clk(gclk));
	jdff dff_A_9JTQdnKu9_0(.dout(w_dff_A_noVY6HwB7_0),.din(w_dff_A_9JTQdnKu9_0),.clk(gclk));
	jdff dff_A_noVY6HwB7_0(.dout(w_dff_A_v1rMq7UA9_0),.din(w_dff_A_noVY6HwB7_0),.clk(gclk));
	jdff dff_A_v1rMq7UA9_0(.dout(w_dff_A_WExnmypd3_0),.din(w_dff_A_v1rMq7UA9_0),.clk(gclk));
	jdff dff_A_WExnmypd3_0(.dout(w_dff_A_RcP08nNg3_0),.din(w_dff_A_WExnmypd3_0),.clk(gclk));
	jdff dff_A_RcP08nNg3_0(.dout(w_dff_A_Z179FsCr8_0),.din(w_dff_A_RcP08nNg3_0),.clk(gclk));
	jdff dff_A_Z179FsCr8_0(.dout(w_dff_A_VOwnRV5i0_0),.din(w_dff_A_Z179FsCr8_0),.clk(gclk));
	jdff dff_A_VOwnRV5i0_0(.dout(w_dff_A_MGRIkIPv5_0),.din(w_dff_A_VOwnRV5i0_0),.clk(gclk));
	jdff dff_A_MGRIkIPv5_0(.dout(w_dff_A_B68fX2v50_0),.din(w_dff_A_MGRIkIPv5_0),.clk(gclk));
	jdff dff_A_B68fX2v50_0(.dout(w_dff_A_KqVPuXUG4_0),.din(w_dff_A_B68fX2v50_0),.clk(gclk));
	jdff dff_A_KqVPuXUG4_0(.dout(w_dff_A_9whzdQBg6_0),.din(w_dff_A_KqVPuXUG4_0),.clk(gclk));
	jdff dff_A_9whzdQBg6_0(.dout(w_dff_A_Cq0ZoSVK5_0),.din(w_dff_A_9whzdQBg6_0),.clk(gclk));
	jdff dff_A_Cq0ZoSVK5_0(.dout(w_dff_A_4ihd7n8u0_0),.din(w_dff_A_Cq0ZoSVK5_0),.clk(gclk));
	jdff dff_A_4ihd7n8u0_0(.dout(w_dff_A_uX8FinwS8_0),.din(w_dff_A_4ihd7n8u0_0),.clk(gclk));
	jdff dff_A_uX8FinwS8_0(.dout(w_dff_A_tbCkAZXf3_0),.din(w_dff_A_uX8FinwS8_0),.clk(gclk));
	jdff dff_A_tbCkAZXf3_0(.dout(w_dff_A_L9QagEZF0_0),.din(w_dff_A_tbCkAZXf3_0),.clk(gclk));
	jdff dff_A_L9QagEZF0_0(.dout(w_dff_A_Bd0HKDFY7_0),.din(w_dff_A_L9QagEZF0_0),.clk(gclk));
	jdff dff_A_Bd0HKDFY7_0(.dout(w_dff_A_LcE5VPro2_0),.din(w_dff_A_Bd0HKDFY7_0),.clk(gclk));
	jdff dff_A_LcE5VPro2_0(.dout(w_dff_A_BCS6BT2t9_0),.din(w_dff_A_LcE5VPro2_0),.clk(gclk));
	jdff dff_A_BCS6BT2t9_0(.dout(w_dff_A_O5mNMmaB9_0),.din(w_dff_A_BCS6BT2t9_0),.clk(gclk));
	jdff dff_A_O5mNMmaB9_0(.dout(w_dff_A_aqz37mCq3_0),.din(w_dff_A_O5mNMmaB9_0),.clk(gclk));
	jdff dff_A_aqz37mCq3_0(.dout(w_dff_A_g7eRWlGo3_0),.din(w_dff_A_aqz37mCq3_0),.clk(gclk));
	jdff dff_A_g7eRWlGo3_0(.dout(w_dff_A_Xqb01NrL2_0),.din(w_dff_A_g7eRWlGo3_0),.clk(gclk));
	jdff dff_A_Xqb01NrL2_0(.dout(w_dff_A_CLSGyjeC9_0),.din(w_dff_A_Xqb01NrL2_0),.clk(gclk));
	jdff dff_A_CLSGyjeC9_0(.dout(w_dff_A_S1Yusywy5_0),.din(w_dff_A_CLSGyjeC9_0),.clk(gclk));
	jdff dff_A_S1Yusywy5_0(.dout(w_dff_A_Sr2E2Dy67_0),.din(w_dff_A_S1Yusywy5_0),.clk(gclk));
	jdff dff_A_Sr2E2Dy67_0(.dout(w_dff_A_Juu2DPc14_0),.din(w_dff_A_Sr2E2Dy67_0),.clk(gclk));
	jdff dff_A_Juu2DPc14_0(.dout(w_dff_A_sFEwPaDj8_0),.din(w_dff_A_Juu2DPc14_0),.clk(gclk));
	jdff dff_A_sFEwPaDj8_0(.dout(w_dff_A_VzD49Oyz8_0),.din(w_dff_A_sFEwPaDj8_0),.clk(gclk));
	jdff dff_A_VzD49Oyz8_0(.dout(w_dff_A_ubPW59ec6_0),.din(w_dff_A_VzD49Oyz8_0),.clk(gclk));
	jdff dff_A_ubPW59ec6_0(.dout(w_dff_A_5rY6TR0a9_0),.din(w_dff_A_ubPW59ec6_0),.clk(gclk));
	jdff dff_A_5rY6TR0a9_0(.dout(w_dff_A_TRIlYsW30_0),.din(w_dff_A_5rY6TR0a9_0),.clk(gclk));
	jdff dff_A_TRIlYsW30_0(.dout(w_dff_A_6KJfzSC90_0),.din(w_dff_A_TRIlYsW30_0),.clk(gclk));
	jdff dff_A_6KJfzSC90_0(.dout(w_dff_A_dBw8ThP34_0),.din(w_dff_A_6KJfzSC90_0),.clk(gclk));
	jdff dff_A_dBw8ThP34_0(.dout(w_dff_A_r5IGKeUn0_0),.din(w_dff_A_dBw8ThP34_0),.clk(gclk));
	jdff dff_A_r5IGKeUn0_0(.dout(w_dff_A_Hy53EKJI8_0),.din(w_dff_A_r5IGKeUn0_0),.clk(gclk));
	jdff dff_A_Hy53EKJI8_0(.dout(w_dff_A_tpdXvOML4_0),.din(w_dff_A_Hy53EKJI8_0),.clk(gclk));
	jdff dff_A_tpdXvOML4_0(.dout(w_dff_A_va51BmCQ9_0),.din(w_dff_A_tpdXvOML4_0),.clk(gclk));
	jdff dff_A_va51BmCQ9_0(.dout(w_dff_A_YN7tNNay4_0),.din(w_dff_A_va51BmCQ9_0),.clk(gclk));
	jdff dff_A_YN7tNNay4_0(.dout(w_dff_A_imQL9fn46_0),.din(w_dff_A_YN7tNNay4_0),.clk(gclk));
	jdff dff_A_imQL9fn46_0(.dout(w_dff_A_396hJunk3_0),.din(w_dff_A_imQL9fn46_0),.clk(gclk));
	jdff dff_A_396hJunk3_0(.dout(w_dff_A_IVgNkzZM8_0),.din(w_dff_A_396hJunk3_0),.clk(gclk));
	jdff dff_A_IVgNkzZM8_0(.dout(w_dff_A_QCtLnjdX3_0),.din(w_dff_A_IVgNkzZM8_0),.clk(gclk));
	jdff dff_A_QCtLnjdX3_0(.dout(w_dff_A_1m1hyP6z8_0),.din(w_dff_A_QCtLnjdX3_0),.clk(gclk));
	jdff dff_A_1m1hyP6z8_0(.dout(w_dff_A_R7HV63Vw0_0),.din(w_dff_A_1m1hyP6z8_0),.clk(gclk));
	jdff dff_A_R7HV63Vw0_0(.dout(w_dff_A_TgzLISqZ2_0),.din(w_dff_A_R7HV63Vw0_0),.clk(gclk));
	jdff dff_A_TgzLISqZ2_0(.dout(w_dff_A_0NBdKgS54_0),.din(w_dff_A_TgzLISqZ2_0),.clk(gclk));
	jdff dff_A_0NBdKgS54_0(.dout(w_dff_A_19S5qRxr3_0),.din(w_dff_A_0NBdKgS54_0),.clk(gclk));
	jdff dff_A_19S5qRxr3_0(.dout(w_dff_A_PnlfMz8I5_0),.din(w_dff_A_19S5qRxr3_0),.clk(gclk));
	jdff dff_A_PnlfMz8I5_0(.dout(w_dff_A_EyVPaNEH4_0),.din(w_dff_A_PnlfMz8I5_0),.clk(gclk));
	jdff dff_A_EyVPaNEH4_0(.dout(w_dff_A_JLEnT9bs8_0),.din(w_dff_A_EyVPaNEH4_0),.clk(gclk));
	jdff dff_A_JLEnT9bs8_0(.dout(w_dff_A_EMfMitW65_0),.din(w_dff_A_JLEnT9bs8_0),.clk(gclk));
	jdff dff_A_EMfMitW65_0(.dout(w_dff_A_yZ71UeeG4_0),.din(w_dff_A_EMfMitW65_0),.clk(gclk));
	jdff dff_A_yZ71UeeG4_0(.dout(w_dff_A_bV8uCmZ90_0),.din(w_dff_A_yZ71UeeG4_0),.clk(gclk));
	jdff dff_A_bV8uCmZ90_0(.dout(w_dff_A_L75unZ0w2_0),.din(w_dff_A_bV8uCmZ90_0),.clk(gclk));
	jdff dff_A_L75unZ0w2_0(.dout(w_dff_A_V2N1sjSX9_0),.din(w_dff_A_L75unZ0w2_0),.clk(gclk));
	jdff dff_A_V2N1sjSX9_0(.dout(w_dff_A_QEKkZaOf6_0),.din(w_dff_A_V2N1sjSX9_0),.clk(gclk));
	jdff dff_A_QEKkZaOf6_0(.dout(w_dff_A_fbbg29LL4_0),.din(w_dff_A_QEKkZaOf6_0),.clk(gclk));
	jdff dff_A_fbbg29LL4_0(.dout(w_dff_A_tmdxY3We9_0),.din(w_dff_A_fbbg29LL4_0),.clk(gclk));
	jdff dff_A_tmdxY3We9_0(.dout(w_dff_A_Z5AYQiKM9_0),.din(w_dff_A_tmdxY3We9_0),.clk(gclk));
	jdff dff_A_Z5AYQiKM9_0(.dout(w_dff_A_RwuSfQ1A3_0),.din(w_dff_A_Z5AYQiKM9_0),.clk(gclk));
	jdff dff_A_RwuSfQ1A3_0(.dout(w_dff_A_xU7Yr7KA6_0),.din(w_dff_A_RwuSfQ1A3_0),.clk(gclk));
	jdff dff_A_xU7Yr7KA6_0(.dout(w_dff_A_GQwdU88m4_0),.din(w_dff_A_xU7Yr7KA6_0),.clk(gclk));
	jdff dff_A_GQwdU88m4_0(.dout(w_dff_A_SSoRjrpe6_0),.din(w_dff_A_GQwdU88m4_0),.clk(gclk));
	jdff dff_A_SSoRjrpe6_0(.dout(w_dff_A_Lqcg1Ngn9_0),.din(w_dff_A_SSoRjrpe6_0),.clk(gclk));
	jdff dff_A_Lqcg1Ngn9_0(.dout(w_dff_A_SGLJI8Q25_0),.din(w_dff_A_Lqcg1Ngn9_0),.clk(gclk));
	jdff dff_A_SGLJI8Q25_0(.dout(w_dff_A_WhjorSEl2_0),.din(w_dff_A_SGLJI8Q25_0),.clk(gclk));
	jdff dff_A_WhjorSEl2_0(.dout(w_dff_A_ajTaRkWl7_0),.din(w_dff_A_WhjorSEl2_0),.clk(gclk));
	jdff dff_A_ajTaRkWl7_0(.dout(w_dff_A_GPrw2l8F5_0),.din(w_dff_A_ajTaRkWl7_0),.clk(gclk));
	jdff dff_A_GPrw2l8F5_0(.dout(w_dff_A_6f4VSBjy6_0),.din(w_dff_A_GPrw2l8F5_0),.clk(gclk));
	jdff dff_A_6f4VSBjy6_0(.dout(w_dff_A_98OqeYdm1_0),.din(w_dff_A_6f4VSBjy6_0),.clk(gclk));
	jdff dff_A_98OqeYdm1_0(.dout(w_dff_A_pFjwNU4X6_0),.din(w_dff_A_98OqeYdm1_0),.clk(gclk));
	jdff dff_A_pFjwNU4X6_0(.dout(w_dff_A_KP3JqESX0_0),.din(w_dff_A_pFjwNU4X6_0),.clk(gclk));
	jdff dff_A_KP3JqESX0_0(.dout(w_dff_A_7m0DZKCr2_0),.din(w_dff_A_KP3JqESX0_0),.clk(gclk));
	jdff dff_A_7m0DZKCr2_0(.dout(w_dff_A_QFuhrs5q5_0),.din(w_dff_A_7m0DZKCr2_0),.clk(gclk));
	jdff dff_A_QFuhrs5q5_0(.dout(w_dff_A_V6W5MPpX4_0),.din(w_dff_A_QFuhrs5q5_0),.clk(gclk));
	jdff dff_A_V6W5MPpX4_0(.dout(w_dff_A_BhZgMGEA0_0),.din(w_dff_A_V6W5MPpX4_0),.clk(gclk));
	jdff dff_A_BhZgMGEA0_0(.dout(f1),.din(w_dff_A_BhZgMGEA0_0),.clk(gclk));
	jdff dff_A_BvD62S921_2(.dout(w_dff_A_gMz6Lb5D8_0),.din(w_dff_A_BvD62S921_2),.clk(gclk));
	jdff dff_A_gMz6Lb5D8_0(.dout(w_dff_A_yLtN7iw95_0),.din(w_dff_A_gMz6Lb5D8_0),.clk(gclk));
	jdff dff_A_yLtN7iw95_0(.dout(w_dff_A_IA3oxORP5_0),.din(w_dff_A_yLtN7iw95_0),.clk(gclk));
	jdff dff_A_IA3oxORP5_0(.dout(w_dff_A_AUiNijlD2_0),.din(w_dff_A_IA3oxORP5_0),.clk(gclk));
	jdff dff_A_AUiNijlD2_0(.dout(w_dff_A_zMekuf8x1_0),.din(w_dff_A_AUiNijlD2_0),.clk(gclk));
	jdff dff_A_zMekuf8x1_0(.dout(w_dff_A_C5IQIOJW6_0),.din(w_dff_A_zMekuf8x1_0),.clk(gclk));
	jdff dff_A_C5IQIOJW6_0(.dout(w_dff_A_j6WANsVL1_0),.din(w_dff_A_C5IQIOJW6_0),.clk(gclk));
	jdff dff_A_j6WANsVL1_0(.dout(w_dff_A_JUMS4rlL9_0),.din(w_dff_A_j6WANsVL1_0),.clk(gclk));
	jdff dff_A_JUMS4rlL9_0(.dout(w_dff_A_b7MWDKxD3_0),.din(w_dff_A_JUMS4rlL9_0),.clk(gclk));
	jdff dff_A_b7MWDKxD3_0(.dout(w_dff_A_L0p1xxS55_0),.din(w_dff_A_b7MWDKxD3_0),.clk(gclk));
	jdff dff_A_L0p1xxS55_0(.dout(w_dff_A_QPb7BxDj1_0),.din(w_dff_A_L0p1xxS55_0),.clk(gclk));
	jdff dff_A_QPb7BxDj1_0(.dout(w_dff_A_zQBw3Rtn4_0),.din(w_dff_A_QPb7BxDj1_0),.clk(gclk));
	jdff dff_A_zQBw3Rtn4_0(.dout(w_dff_A_La4d9nsL1_0),.din(w_dff_A_zQBw3Rtn4_0),.clk(gclk));
	jdff dff_A_La4d9nsL1_0(.dout(w_dff_A_FhHZAgEC8_0),.din(w_dff_A_La4d9nsL1_0),.clk(gclk));
	jdff dff_A_FhHZAgEC8_0(.dout(w_dff_A_m1qLRZr12_0),.din(w_dff_A_FhHZAgEC8_0),.clk(gclk));
	jdff dff_A_m1qLRZr12_0(.dout(w_dff_A_AOAbQvcI2_0),.din(w_dff_A_m1qLRZr12_0),.clk(gclk));
	jdff dff_A_AOAbQvcI2_0(.dout(w_dff_A_0frBFz460_0),.din(w_dff_A_AOAbQvcI2_0),.clk(gclk));
	jdff dff_A_0frBFz460_0(.dout(w_dff_A_FZdDIpnV1_0),.din(w_dff_A_0frBFz460_0),.clk(gclk));
	jdff dff_A_FZdDIpnV1_0(.dout(w_dff_A_pcJmtdQc1_0),.din(w_dff_A_FZdDIpnV1_0),.clk(gclk));
	jdff dff_A_pcJmtdQc1_0(.dout(w_dff_A_hi8IlDSj0_0),.din(w_dff_A_pcJmtdQc1_0),.clk(gclk));
	jdff dff_A_hi8IlDSj0_0(.dout(w_dff_A_6eUrlbcC0_0),.din(w_dff_A_hi8IlDSj0_0),.clk(gclk));
	jdff dff_A_6eUrlbcC0_0(.dout(w_dff_A_CiCKQe8J9_0),.din(w_dff_A_6eUrlbcC0_0),.clk(gclk));
	jdff dff_A_CiCKQe8J9_0(.dout(w_dff_A_uwkglmLH0_0),.din(w_dff_A_CiCKQe8J9_0),.clk(gclk));
	jdff dff_A_uwkglmLH0_0(.dout(w_dff_A_Fxxmc7iO8_0),.din(w_dff_A_uwkglmLH0_0),.clk(gclk));
	jdff dff_A_Fxxmc7iO8_0(.dout(w_dff_A_F57YYRhM2_0),.din(w_dff_A_Fxxmc7iO8_0),.clk(gclk));
	jdff dff_A_F57YYRhM2_0(.dout(w_dff_A_ChVRGd0L0_0),.din(w_dff_A_F57YYRhM2_0),.clk(gclk));
	jdff dff_A_ChVRGd0L0_0(.dout(w_dff_A_7IDO9qf89_0),.din(w_dff_A_ChVRGd0L0_0),.clk(gclk));
	jdff dff_A_7IDO9qf89_0(.dout(w_dff_A_34iojwkP1_0),.din(w_dff_A_7IDO9qf89_0),.clk(gclk));
	jdff dff_A_34iojwkP1_0(.dout(w_dff_A_DUHIAmDv9_0),.din(w_dff_A_34iojwkP1_0),.clk(gclk));
	jdff dff_A_DUHIAmDv9_0(.dout(w_dff_A_sDpan7jS9_0),.din(w_dff_A_DUHIAmDv9_0),.clk(gclk));
	jdff dff_A_sDpan7jS9_0(.dout(w_dff_A_WVVgc9Sf9_0),.din(w_dff_A_sDpan7jS9_0),.clk(gclk));
	jdff dff_A_WVVgc9Sf9_0(.dout(w_dff_A_53N0H0zX5_0),.din(w_dff_A_WVVgc9Sf9_0),.clk(gclk));
	jdff dff_A_53N0H0zX5_0(.dout(w_dff_A_6MXTdlQ91_0),.din(w_dff_A_53N0H0zX5_0),.clk(gclk));
	jdff dff_A_6MXTdlQ91_0(.dout(w_dff_A_C97PlHyO2_0),.din(w_dff_A_6MXTdlQ91_0),.clk(gclk));
	jdff dff_A_C97PlHyO2_0(.dout(w_dff_A_tLb5D9S65_0),.din(w_dff_A_C97PlHyO2_0),.clk(gclk));
	jdff dff_A_tLb5D9S65_0(.dout(w_dff_A_t7G32yOC5_0),.din(w_dff_A_tLb5D9S65_0),.clk(gclk));
	jdff dff_A_t7G32yOC5_0(.dout(w_dff_A_H54wYtCl3_0),.din(w_dff_A_t7G32yOC5_0),.clk(gclk));
	jdff dff_A_H54wYtCl3_0(.dout(w_dff_A_XfdL9HlW6_0),.din(w_dff_A_H54wYtCl3_0),.clk(gclk));
	jdff dff_A_XfdL9HlW6_0(.dout(w_dff_A_pIdsk8F65_0),.din(w_dff_A_XfdL9HlW6_0),.clk(gclk));
	jdff dff_A_pIdsk8F65_0(.dout(w_dff_A_ZMs4jKWp8_0),.din(w_dff_A_pIdsk8F65_0),.clk(gclk));
	jdff dff_A_ZMs4jKWp8_0(.dout(w_dff_A_nkNIQKSY4_0),.din(w_dff_A_ZMs4jKWp8_0),.clk(gclk));
	jdff dff_A_nkNIQKSY4_0(.dout(w_dff_A_0Fk5wTtC2_0),.din(w_dff_A_nkNIQKSY4_0),.clk(gclk));
	jdff dff_A_0Fk5wTtC2_0(.dout(w_dff_A_o4DQiZVa7_0),.din(w_dff_A_0Fk5wTtC2_0),.clk(gclk));
	jdff dff_A_o4DQiZVa7_0(.dout(w_dff_A_h1Jt0UWn1_0),.din(w_dff_A_o4DQiZVa7_0),.clk(gclk));
	jdff dff_A_h1Jt0UWn1_0(.dout(w_dff_A_GCnye3ZX9_0),.din(w_dff_A_h1Jt0UWn1_0),.clk(gclk));
	jdff dff_A_GCnye3ZX9_0(.dout(w_dff_A_7NPpwmKi3_0),.din(w_dff_A_GCnye3ZX9_0),.clk(gclk));
	jdff dff_A_7NPpwmKi3_0(.dout(w_dff_A_cfpTaVgI3_0),.din(w_dff_A_7NPpwmKi3_0),.clk(gclk));
	jdff dff_A_cfpTaVgI3_0(.dout(w_dff_A_ZAB4PPed8_0),.din(w_dff_A_cfpTaVgI3_0),.clk(gclk));
	jdff dff_A_ZAB4PPed8_0(.dout(w_dff_A_EJeNXIFi1_0),.din(w_dff_A_ZAB4PPed8_0),.clk(gclk));
	jdff dff_A_EJeNXIFi1_0(.dout(w_dff_A_X1nkO6wo0_0),.din(w_dff_A_EJeNXIFi1_0),.clk(gclk));
	jdff dff_A_X1nkO6wo0_0(.dout(w_dff_A_1RnWr8J29_0),.din(w_dff_A_X1nkO6wo0_0),.clk(gclk));
	jdff dff_A_1RnWr8J29_0(.dout(w_dff_A_nDsazNLQ9_0),.din(w_dff_A_1RnWr8J29_0),.clk(gclk));
	jdff dff_A_nDsazNLQ9_0(.dout(w_dff_A_3nqhLmj45_0),.din(w_dff_A_nDsazNLQ9_0),.clk(gclk));
	jdff dff_A_3nqhLmj45_0(.dout(w_dff_A_bN1SHJC38_0),.din(w_dff_A_3nqhLmj45_0),.clk(gclk));
	jdff dff_A_bN1SHJC38_0(.dout(w_dff_A_zME2Tpf04_0),.din(w_dff_A_bN1SHJC38_0),.clk(gclk));
	jdff dff_A_zME2Tpf04_0(.dout(w_dff_A_7k56kaHd7_0),.din(w_dff_A_zME2Tpf04_0),.clk(gclk));
	jdff dff_A_7k56kaHd7_0(.dout(w_dff_A_1hCIaHIB3_0),.din(w_dff_A_7k56kaHd7_0),.clk(gclk));
	jdff dff_A_1hCIaHIB3_0(.dout(w_dff_A_yngkKjXy7_0),.din(w_dff_A_1hCIaHIB3_0),.clk(gclk));
	jdff dff_A_yngkKjXy7_0(.dout(w_dff_A_xMFeIU907_0),.din(w_dff_A_yngkKjXy7_0),.clk(gclk));
	jdff dff_A_xMFeIU907_0(.dout(w_dff_A_HcXcIV3N6_0),.din(w_dff_A_xMFeIU907_0),.clk(gclk));
	jdff dff_A_HcXcIV3N6_0(.dout(w_dff_A_fR0Ob4G44_0),.din(w_dff_A_HcXcIV3N6_0),.clk(gclk));
	jdff dff_A_fR0Ob4G44_0(.dout(w_dff_A_2ykFKu2t5_0),.din(w_dff_A_fR0Ob4G44_0),.clk(gclk));
	jdff dff_A_2ykFKu2t5_0(.dout(w_dff_A_jm9LYl8C6_0),.din(w_dff_A_2ykFKu2t5_0),.clk(gclk));
	jdff dff_A_jm9LYl8C6_0(.dout(w_dff_A_tUp7NdTr2_0),.din(w_dff_A_jm9LYl8C6_0),.clk(gclk));
	jdff dff_A_tUp7NdTr2_0(.dout(w_dff_A_bwTsA3Q15_0),.din(w_dff_A_tUp7NdTr2_0),.clk(gclk));
	jdff dff_A_bwTsA3Q15_0(.dout(w_dff_A_eXAvG3xU4_0),.din(w_dff_A_bwTsA3Q15_0),.clk(gclk));
	jdff dff_A_eXAvG3xU4_0(.dout(w_dff_A_KDyacK611_0),.din(w_dff_A_eXAvG3xU4_0),.clk(gclk));
	jdff dff_A_KDyacK611_0(.dout(w_dff_A_jPiwoq8Q8_0),.din(w_dff_A_KDyacK611_0),.clk(gclk));
	jdff dff_A_jPiwoq8Q8_0(.dout(w_dff_A_fGDojP762_0),.din(w_dff_A_jPiwoq8Q8_0),.clk(gclk));
	jdff dff_A_fGDojP762_0(.dout(w_dff_A_VyoFmQkw5_0),.din(w_dff_A_fGDojP762_0),.clk(gclk));
	jdff dff_A_VyoFmQkw5_0(.dout(w_dff_A_T8khXwxt6_0),.din(w_dff_A_VyoFmQkw5_0),.clk(gclk));
	jdff dff_A_T8khXwxt6_0(.dout(w_dff_A_K73VURR94_0),.din(w_dff_A_T8khXwxt6_0),.clk(gclk));
	jdff dff_A_K73VURR94_0(.dout(w_dff_A_EUMWAIkn3_0),.din(w_dff_A_K73VURR94_0),.clk(gclk));
	jdff dff_A_EUMWAIkn3_0(.dout(w_dff_A_WEXHHw9z4_0),.din(w_dff_A_EUMWAIkn3_0),.clk(gclk));
	jdff dff_A_WEXHHw9z4_0(.dout(w_dff_A_eazaBLVO4_0),.din(w_dff_A_WEXHHw9z4_0),.clk(gclk));
	jdff dff_A_eazaBLVO4_0(.dout(w_dff_A_rjirzV5f0_0),.din(w_dff_A_eazaBLVO4_0),.clk(gclk));
	jdff dff_A_rjirzV5f0_0(.dout(w_dff_A_Czdqyu6Y0_0),.din(w_dff_A_rjirzV5f0_0),.clk(gclk));
	jdff dff_A_Czdqyu6Y0_0(.dout(w_dff_A_Z1Laxp9i4_0),.din(w_dff_A_Czdqyu6Y0_0),.clk(gclk));
	jdff dff_A_Z1Laxp9i4_0(.dout(w_dff_A_15Gtg2h36_0),.din(w_dff_A_Z1Laxp9i4_0),.clk(gclk));
	jdff dff_A_15Gtg2h36_0(.dout(w_dff_A_QpFTH8B80_0),.din(w_dff_A_15Gtg2h36_0),.clk(gclk));
	jdff dff_A_QpFTH8B80_0(.dout(w_dff_A_V9QrQztm9_0),.din(w_dff_A_QpFTH8B80_0),.clk(gclk));
	jdff dff_A_V9QrQztm9_0(.dout(w_dff_A_qRYXWz9X8_0),.din(w_dff_A_V9QrQztm9_0),.clk(gclk));
	jdff dff_A_qRYXWz9X8_0(.dout(w_dff_A_xFtAuA2J5_0),.din(w_dff_A_qRYXWz9X8_0),.clk(gclk));
	jdff dff_A_xFtAuA2J5_0(.dout(w_dff_A_fmsyS0um0_0),.din(w_dff_A_xFtAuA2J5_0),.clk(gclk));
	jdff dff_A_fmsyS0um0_0(.dout(w_dff_A_m9HoNS8u7_0),.din(w_dff_A_fmsyS0um0_0),.clk(gclk));
	jdff dff_A_m9HoNS8u7_0(.dout(w_dff_A_YY7pLLwB6_0),.din(w_dff_A_m9HoNS8u7_0),.clk(gclk));
	jdff dff_A_YY7pLLwB6_0(.dout(w_dff_A_pkQtA9eJ2_0),.din(w_dff_A_YY7pLLwB6_0),.clk(gclk));
	jdff dff_A_pkQtA9eJ2_0(.dout(w_dff_A_PCclndeQ9_0),.din(w_dff_A_pkQtA9eJ2_0),.clk(gclk));
	jdff dff_A_PCclndeQ9_0(.dout(w_dff_A_4kthRXsq7_0),.din(w_dff_A_PCclndeQ9_0),.clk(gclk));
	jdff dff_A_4kthRXsq7_0(.dout(w_dff_A_kNM1InUm8_0),.din(w_dff_A_4kthRXsq7_0),.clk(gclk));
	jdff dff_A_kNM1InUm8_0(.dout(w_dff_A_5LvdS70S0_0),.din(w_dff_A_kNM1InUm8_0),.clk(gclk));
	jdff dff_A_5LvdS70S0_0(.dout(w_dff_A_pK93onTu3_0),.din(w_dff_A_5LvdS70S0_0),.clk(gclk));
	jdff dff_A_pK93onTu3_0(.dout(w_dff_A_YX6yAdRf8_0),.din(w_dff_A_pK93onTu3_0),.clk(gclk));
	jdff dff_A_YX6yAdRf8_0(.dout(w_dff_A_rckmqZmE9_0),.din(w_dff_A_YX6yAdRf8_0),.clk(gclk));
	jdff dff_A_rckmqZmE9_0(.dout(w_dff_A_dZJDu4xZ9_0),.din(w_dff_A_rckmqZmE9_0),.clk(gclk));
	jdff dff_A_dZJDu4xZ9_0(.dout(w_dff_A_0jpG0GS89_0),.din(w_dff_A_dZJDu4xZ9_0),.clk(gclk));
	jdff dff_A_0jpG0GS89_0(.dout(w_dff_A_93fubIHx8_0),.din(w_dff_A_0jpG0GS89_0),.clk(gclk));
	jdff dff_A_93fubIHx8_0(.dout(w_dff_A_IuzcCOiA7_0),.din(w_dff_A_93fubIHx8_0),.clk(gclk));
	jdff dff_A_IuzcCOiA7_0(.dout(w_dff_A_ISeyzKuN8_0),.din(w_dff_A_IuzcCOiA7_0),.clk(gclk));
	jdff dff_A_ISeyzKuN8_0(.dout(w_dff_A_grOGOaF14_0),.din(w_dff_A_ISeyzKuN8_0),.clk(gclk));
	jdff dff_A_grOGOaF14_0(.dout(w_dff_A_ZzJuS0Wi2_0),.din(w_dff_A_grOGOaF14_0),.clk(gclk));
	jdff dff_A_ZzJuS0Wi2_0(.dout(w_dff_A_bPAKUw0p5_0),.din(w_dff_A_ZzJuS0Wi2_0),.clk(gclk));
	jdff dff_A_bPAKUw0p5_0(.dout(w_dff_A_VNSZvRpl0_0),.din(w_dff_A_bPAKUw0p5_0),.clk(gclk));
	jdff dff_A_VNSZvRpl0_0(.dout(w_dff_A_ab6HyjvL7_0),.din(w_dff_A_VNSZvRpl0_0),.clk(gclk));
	jdff dff_A_ab6HyjvL7_0(.dout(w_dff_A_95N8oCST4_0),.din(w_dff_A_ab6HyjvL7_0),.clk(gclk));
	jdff dff_A_95N8oCST4_0(.dout(w_dff_A_kDxktsP28_0),.din(w_dff_A_95N8oCST4_0),.clk(gclk));
	jdff dff_A_kDxktsP28_0(.dout(w_dff_A_k9lIUXm30_0),.din(w_dff_A_kDxktsP28_0),.clk(gclk));
	jdff dff_A_k9lIUXm30_0(.dout(w_dff_A_jpGpTGH53_0),.din(w_dff_A_k9lIUXm30_0),.clk(gclk));
	jdff dff_A_jpGpTGH53_0(.dout(w_dff_A_57lRtJJu5_0),.din(w_dff_A_jpGpTGH53_0),.clk(gclk));
	jdff dff_A_57lRtJJu5_0(.dout(w_dff_A_ozZC3i9t3_0),.din(w_dff_A_57lRtJJu5_0),.clk(gclk));
	jdff dff_A_ozZC3i9t3_0(.dout(w_dff_A_FL5FHqTE2_0),.din(w_dff_A_ozZC3i9t3_0),.clk(gclk));
	jdff dff_A_FL5FHqTE2_0(.dout(w_dff_A_ou4I5wYa1_0),.din(w_dff_A_FL5FHqTE2_0),.clk(gclk));
	jdff dff_A_ou4I5wYa1_0(.dout(w_dff_A_4lFlDF7p6_0),.din(w_dff_A_ou4I5wYa1_0),.clk(gclk));
	jdff dff_A_4lFlDF7p6_0(.dout(w_dff_A_bxIXJpTJ0_0),.din(w_dff_A_4lFlDF7p6_0),.clk(gclk));
	jdff dff_A_bxIXJpTJ0_0(.dout(w_dff_A_gTy9ccLO5_0),.din(w_dff_A_bxIXJpTJ0_0),.clk(gclk));
	jdff dff_A_gTy9ccLO5_0(.dout(w_dff_A_xDWTr75G7_0),.din(w_dff_A_gTy9ccLO5_0),.clk(gclk));
	jdff dff_A_xDWTr75G7_0(.dout(w_dff_A_MV3cRGsb8_0),.din(w_dff_A_xDWTr75G7_0),.clk(gclk));
	jdff dff_A_MV3cRGsb8_0(.dout(w_dff_A_plKD2YaN9_0),.din(w_dff_A_MV3cRGsb8_0),.clk(gclk));
	jdff dff_A_plKD2YaN9_0(.dout(w_dff_A_5a8Is8P98_0),.din(w_dff_A_plKD2YaN9_0),.clk(gclk));
	jdff dff_A_5a8Is8P98_0(.dout(w_dff_A_ZQfeTGbs4_0),.din(w_dff_A_5a8Is8P98_0),.clk(gclk));
	jdff dff_A_ZQfeTGbs4_0(.dout(w_dff_A_xLY0Q4XN2_0),.din(w_dff_A_ZQfeTGbs4_0),.clk(gclk));
	jdff dff_A_xLY0Q4XN2_0(.dout(w_dff_A_25MA11i46_0),.din(w_dff_A_xLY0Q4XN2_0),.clk(gclk));
	jdff dff_A_25MA11i46_0(.dout(w_dff_A_P1xX5SoN3_0),.din(w_dff_A_25MA11i46_0),.clk(gclk));
	jdff dff_A_P1xX5SoN3_0(.dout(w_dff_A_qRlywRaA1_0),.din(w_dff_A_P1xX5SoN3_0),.clk(gclk));
	jdff dff_A_qRlywRaA1_0(.dout(f2),.din(w_dff_A_qRlywRaA1_0),.clk(gclk));
	jdff dff_A_lRUw1Ruu2_2(.dout(w_dff_A_La1LKto64_0),.din(w_dff_A_lRUw1Ruu2_2),.clk(gclk));
	jdff dff_A_La1LKto64_0(.dout(w_dff_A_bdp3MxDE8_0),.din(w_dff_A_La1LKto64_0),.clk(gclk));
	jdff dff_A_bdp3MxDE8_0(.dout(w_dff_A_WqgofUlT6_0),.din(w_dff_A_bdp3MxDE8_0),.clk(gclk));
	jdff dff_A_WqgofUlT6_0(.dout(w_dff_A_HURVWnDK0_0),.din(w_dff_A_WqgofUlT6_0),.clk(gclk));
	jdff dff_A_HURVWnDK0_0(.dout(w_dff_A_tE3EP4Gv0_0),.din(w_dff_A_HURVWnDK0_0),.clk(gclk));
	jdff dff_A_tE3EP4Gv0_0(.dout(w_dff_A_aq0xns4Z7_0),.din(w_dff_A_tE3EP4Gv0_0),.clk(gclk));
	jdff dff_A_aq0xns4Z7_0(.dout(w_dff_A_3nR77eZh3_0),.din(w_dff_A_aq0xns4Z7_0),.clk(gclk));
	jdff dff_A_3nR77eZh3_0(.dout(w_dff_A_Ah14sbfU8_0),.din(w_dff_A_3nR77eZh3_0),.clk(gclk));
	jdff dff_A_Ah14sbfU8_0(.dout(w_dff_A_1WcRL1Tj4_0),.din(w_dff_A_Ah14sbfU8_0),.clk(gclk));
	jdff dff_A_1WcRL1Tj4_0(.dout(w_dff_A_ONCu3cv30_0),.din(w_dff_A_1WcRL1Tj4_0),.clk(gclk));
	jdff dff_A_ONCu3cv30_0(.dout(w_dff_A_KDg5tI2k3_0),.din(w_dff_A_ONCu3cv30_0),.clk(gclk));
	jdff dff_A_KDg5tI2k3_0(.dout(w_dff_A_235zJRRa7_0),.din(w_dff_A_KDg5tI2k3_0),.clk(gclk));
	jdff dff_A_235zJRRa7_0(.dout(w_dff_A_aOiZ6Bzx1_0),.din(w_dff_A_235zJRRa7_0),.clk(gclk));
	jdff dff_A_aOiZ6Bzx1_0(.dout(w_dff_A_FChoMAaX2_0),.din(w_dff_A_aOiZ6Bzx1_0),.clk(gclk));
	jdff dff_A_FChoMAaX2_0(.dout(w_dff_A_pCtOXO764_0),.din(w_dff_A_FChoMAaX2_0),.clk(gclk));
	jdff dff_A_pCtOXO764_0(.dout(w_dff_A_0h8zISNG9_0),.din(w_dff_A_pCtOXO764_0),.clk(gclk));
	jdff dff_A_0h8zISNG9_0(.dout(w_dff_A_fF46Ozse3_0),.din(w_dff_A_0h8zISNG9_0),.clk(gclk));
	jdff dff_A_fF46Ozse3_0(.dout(w_dff_A_gi1fmzJE6_0),.din(w_dff_A_fF46Ozse3_0),.clk(gclk));
	jdff dff_A_gi1fmzJE6_0(.dout(w_dff_A_gaqTL2bo9_0),.din(w_dff_A_gi1fmzJE6_0),.clk(gclk));
	jdff dff_A_gaqTL2bo9_0(.dout(w_dff_A_Ax5bWosD2_0),.din(w_dff_A_gaqTL2bo9_0),.clk(gclk));
	jdff dff_A_Ax5bWosD2_0(.dout(w_dff_A_ctSG34BC7_0),.din(w_dff_A_Ax5bWosD2_0),.clk(gclk));
	jdff dff_A_ctSG34BC7_0(.dout(w_dff_A_IaQmkzvh0_0),.din(w_dff_A_ctSG34BC7_0),.clk(gclk));
	jdff dff_A_IaQmkzvh0_0(.dout(w_dff_A_rgU0Bqgn6_0),.din(w_dff_A_IaQmkzvh0_0),.clk(gclk));
	jdff dff_A_rgU0Bqgn6_0(.dout(w_dff_A_hqA5agcV1_0),.din(w_dff_A_rgU0Bqgn6_0),.clk(gclk));
	jdff dff_A_hqA5agcV1_0(.dout(w_dff_A_h3XBLhf63_0),.din(w_dff_A_hqA5agcV1_0),.clk(gclk));
	jdff dff_A_h3XBLhf63_0(.dout(w_dff_A_G2k3SXBg8_0),.din(w_dff_A_h3XBLhf63_0),.clk(gclk));
	jdff dff_A_G2k3SXBg8_0(.dout(w_dff_A_3GpCjouF8_0),.din(w_dff_A_G2k3SXBg8_0),.clk(gclk));
	jdff dff_A_3GpCjouF8_0(.dout(w_dff_A_yHuxXgw80_0),.din(w_dff_A_3GpCjouF8_0),.clk(gclk));
	jdff dff_A_yHuxXgw80_0(.dout(w_dff_A_RRLV3ErP9_0),.din(w_dff_A_yHuxXgw80_0),.clk(gclk));
	jdff dff_A_RRLV3ErP9_0(.dout(w_dff_A_zj0CkmKh7_0),.din(w_dff_A_RRLV3ErP9_0),.clk(gclk));
	jdff dff_A_zj0CkmKh7_0(.dout(w_dff_A_lem8Aolv3_0),.din(w_dff_A_zj0CkmKh7_0),.clk(gclk));
	jdff dff_A_lem8Aolv3_0(.dout(w_dff_A_6Vmug3QF6_0),.din(w_dff_A_lem8Aolv3_0),.clk(gclk));
	jdff dff_A_6Vmug3QF6_0(.dout(w_dff_A_fDNILKEJ8_0),.din(w_dff_A_6Vmug3QF6_0),.clk(gclk));
	jdff dff_A_fDNILKEJ8_0(.dout(w_dff_A_9lTlUCnX7_0),.din(w_dff_A_fDNILKEJ8_0),.clk(gclk));
	jdff dff_A_9lTlUCnX7_0(.dout(w_dff_A_24lpbOJf9_0),.din(w_dff_A_9lTlUCnX7_0),.clk(gclk));
	jdff dff_A_24lpbOJf9_0(.dout(w_dff_A_kbYCQ5jM7_0),.din(w_dff_A_24lpbOJf9_0),.clk(gclk));
	jdff dff_A_kbYCQ5jM7_0(.dout(w_dff_A_Utn0vbNx7_0),.din(w_dff_A_kbYCQ5jM7_0),.clk(gclk));
	jdff dff_A_Utn0vbNx7_0(.dout(w_dff_A_ik0m86LA5_0),.din(w_dff_A_Utn0vbNx7_0),.clk(gclk));
	jdff dff_A_ik0m86LA5_0(.dout(w_dff_A_0bcUWQKt5_0),.din(w_dff_A_ik0m86LA5_0),.clk(gclk));
	jdff dff_A_0bcUWQKt5_0(.dout(w_dff_A_MiWzcOCo6_0),.din(w_dff_A_0bcUWQKt5_0),.clk(gclk));
	jdff dff_A_MiWzcOCo6_0(.dout(w_dff_A_o6g47jgN2_0),.din(w_dff_A_MiWzcOCo6_0),.clk(gclk));
	jdff dff_A_o6g47jgN2_0(.dout(w_dff_A_Ojr2sefc3_0),.din(w_dff_A_o6g47jgN2_0),.clk(gclk));
	jdff dff_A_Ojr2sefc3_0(.dout(w_dff_A_fpXtYxcH7_0),.din(w_dff_A_Ojr2sefc3_0),.clk(gclk));
	jdff dff_A_fpXtYxcH7_0(.dout(w_dff_A_tzuzDKzW6_0),.din(w_dff_A_fpXtYxcH7_0),.clk(gclk));
	jdff dff_A_tzuzDKzW6_0(.dout(w_dff_A_REThOIV03_0),.din(w_dff_A_tzuzDKzW6_0),.clk(gclk));
	jdff dff_A_REThOIV03_0(.dout(w_dff_A_nssv3Qjd3_0),.din(w_dff_A_REThOIV03_0),.clk(gclk));
	jdff dff_A_nssv3Qjd3_0(.dout(w_dff_A_9zVim3YN2_0),.din(w_dff_A_nssv3Qjd3_0),.clk(gclk));
	jdff dff_A_9zVim3YN2_0(.dout(w_dff_A_NzYZyxNE7_0),.din(w_dff_A_9zVim3YN2_0),.clk(gclk));
	jdff dff_A_NzYZyxNE7_0(.dout(w_dff_A_zwYNBsE24_0),.din(w_dff_A_NzYZyxNE7_0),.clk(gclk));
	jdff dff_A_zwYNBsE24_0(.dout(w_dff_A_hAQEzWNP0_0),.din(w_dff_A_zwYNBsE24_0),.clk(gclk));
	jdff dff_A_hAQEzWNP0_0(.dout(w_dff_A_8fjYSDN06_0),.din(w_dff_A_hAQEzWNP0_0),.clk(gclk));
	jdff dff_A_8fjYSDN06_0(.dout(w_dff_A_8nW0GRpX9_0),.din(w_dff_A_8fjYSDN06_0),.clk(gclk));
	jdff dff_A_8nW0GRpX9_0(.dout(w_dff_A_BMshOraN6_0),.din(w_dff_A_8nW0GRpX9_0),.clk(gclk));
	jdff dff_A_BMshOraN6_0(.dout(w_dff_A_0N8IAiOv9_0),.din(w_dff_A_BMshOraN6_0),.clk(gclk));
	jdff dff_A_0N8IAiOv9_0(.dout(w_dff_A_hahuCbq42_0),.din(w_dff_A_0N8IAiOv9_0),.clk(gclk));
	jdff dff_A_hahuCbq42_0(.dout(w_dff_A_6ykzNZKe3_0),.din(w_dff_A_hahuCbq42_0),.clk(gclk));
	jdff dff_A_6ykzNZKe3_0(.dout(w_dff_A_INdv5qFp5_0),.din(w_dff_A_6ykzNZKe3_0),.clk(gclk));
	jdff dff_A_INdv5qFp5_0(.dout(w_dff_A_duTSnfOO7_0),.din(w_dff_A_INdv5qFp5_0),.clk(gclk));
	jdff dff_A_duTSnfOO7_0(.dout(w_dff_A_nwTJnMl86_0),.din(w_dff_A_duTSnfOO7_0),.clk(gclk));
	jdff dff_A_nwTJnMl86_0(.dout(w_dff_A_V6AQytRS5_0),.din(w_dff_A_nwTJnMl86_0),.clk(gclk));
	jdff dff_A_V6AQytRS5_0(.dout(w_dff_A_Hl27t9hM6_0),.din(w_dff_A_V6AQytRS5_0),.clk(gclk));
	jdff dff_A_Hl27t9hM6_0(.dout(w_dff_A_dRyg1Mam4_0),.din(w_dff_A_Hl27t9hM6_0),.clk(gclk));
	jdff dff_A_dRyg1Mam4_0(.dout(w_dff_A_6FlbFwlC6_0),.din(w_dff_A_dRyg1Mam4_0),.clk(gclk));
	jdff dff_A_6FlbFwlC6_0(.dout(w_dff_A_v13qb5nq7_0),.din(w_dff_A_6FlbFwlC6_0),.clk(gclk));
	jdff dff_A_v13qb5nq7_0(.dout(w_dff_A_c6hh5IUo6_0),.din(w_dff_A_v13qb5nq7_0),.clk(gclk));
	jdff dff_A_c6hh5IUo6_0(.dout(w_dff_A_hbFtzmBo3_0),.din(w_dff_A_c6hh5IUo6_0),.clk(gclk));
	jdff dff_A_hbFtzmBo3_0(.dout(w_dff_A_kxGQXqtr9_0),.din(w_dff_A_hbFtzmBo3_0),.clk(gclk));
	jdff dff_A_kxGQXqtr9_0(.dout(w_dff_A_JDnZjqQp7_0),.din(w_dff_A_kxGQXqtr9_0),.clk(gclk));
	jdff dff_A_JDnZjqQp7_0(.dout(w_dff_A_fKgz4nob1_0),.din(w_dff_A_JDnZjqQp7_0),.clk(gclk));
	jdff dff_A_fKgz4nob1_0(.dout(w_dff_A_KkpAdIZ04_0),.din(w_dff_A_fKgz4nob1_0),.clk(gclk));
	jdff dff_A_KkpAdIZ04_0(.dout(w_dff_A_b6SKdcWb7_0),.din(w_dff_A_KkpAdIZ04_0),.clk(gclk));
	jdff dff_A_b6SKdcWb7_0(.dout(w_dff_A_i3payFii8_0),.din(w_dff_A_b6SKdcWb7_0),.clk(gclk));
	jdff dff_A_i3payFii8_0(.dout(w_dff_A_R6ME8LkR2_0),.din(w_dff_A_i3payFii8_0),.clk(gclk));
	jdff dff_A_R6ME8LkR2_0(.dout(w_dff_A_vHWmL4bY5_0),.din(w_dff_A_R6ME8LkR2_0),.clk(gclk));
	jdff dff_A_vHWmL4bY5_0(.dout(w_dff_A_fxuGvgar1_0),.din(w_dff_A_vHWmL4bY5_0),.clk(gclk));
	jdff dff_A_fxuGvgar1_0(.dout(w_dff_A_monQdnWv6_0),.din(w_dff_A_fxuGvgar1_0),.clk(gclk));
	jdff dff_A_monQdnWv6_0(.dout(w_dff_A_vYhJ3o3P3_0),.din(w_dff_A_monQdnWv6_0),.clk(gclk));
	jdff dff_A_vYhJ3o3P3_0(.dout(w_dff_A_qOYDpDCm0_0),.din(w_dff_A_vYhJ3o3P3_0),.clk(gclk));
	jdff dff_A_qOYDpDCm0_0(.dout(w_dff_A_PcI56gSH0_0),.din(w_dff_A_qOYDpDCm0_0),.clk(gclk));
	jdff dff_A_PcI56gSH0_0(.dout(w_dff_A_L7RLkWpq5_0),.din(w_dff_A_PcI56gSH0_0),.clk(gclk));
	jdff dff_A_L7RLkWpq5_0(.dout(w_dff_A_APOk7nlo8_0),.din(w_dff_A_L7RLkWpq5_0),.clk(gclk));
	jdff dff_A_APOk7nlo8_0(.dout(w_dff_A_V8oT1Aak0_0),.din(w_dff_A_APOk7nlo8_0),.clk(gclk));
	jdff dff_A_V8oT1Aak0_0(.dout(w_dff_A_6Wo7BBeT1_0),.din(w_dff_A_V8oT1Aak0_0),.clk(gclk));
	jdff dff_A_6Wo7BBeT1_0(.dout(w_dff_A_AVszMIfw3_0),.din(w_dff_A_6Wo7BBeT1_0),.clk(gclk));
	jdff dff_A_AVszMIfw3_0(.dout(w_dff_A_ndAAfpjO1_0),.din(w_dff_A_AVszMIfw3_0),.clk(gclk));
	jdff dff_A_ndAAfpjO1_0(.dout(w_dff_A_MycMRMU68_0),.din(w_dff_A_ndAAfpjO1_0),.clk(gclk));
	jdff dff_A_MycMRMU68_0(.dout(w_dff_A_o6KCc00R9_0),.din(w_dff_A_MycMRMU68_0),.clk(gclk));
	jdff dff_A_o6KCc00R9_0(.dout(w_dff_A_ElfwmsAm5_0),.din(w_dff_A_o6KCc00R9_0),.clk(gclk));
	jdff dff_A_ElfwmsAm5_0(.dout(w_dff_A_QncfXZiP9_0),.din(w_dff_A_ElfwmsAm5_0),.clk(gclk));
	jdff dff_A_QncfXZiP9_0(.dout(w_dff_A_cFHV3YQ45_0),.din(w_dff_A_QncfXZiP9_0),.clk(gclk));
	jdff dff_A_cFHV3YQ45_0(.dout(w_dff_A_OTrGdUVH8_0),.din(w_dff_A_cFHV3YQ45_0),.clk(gclk));
	jdff dff_A_OTrGdUVH8_0(.dout(w_dff_A_N2ERbr8I4_0),.din(w_dff_A_OTrGdUVH8_0),.clk(gclk));
	jdff dff_A_N2ERbr8I4_0(.dout(w_dff_A_ZIs4rbFq8_0),.din(w_dff_A_N2ERbr8I4_0),.clk(gclk));
	jdff dff_A_ZIs4rbFq8_0(.dout(w_dff_A_AZUEEfxO7_0),.din(w_dff_A_ZIs4rbFq8_0),.clk(gclk));
	jdff dff_A_AZUEEfxO7_0(.dout(w_dff_A_iLufhf6o8_0),.din(w_dff_A_AZUEEfxO7_0),.clk(gclk));
	jdff dff_A_iLufhf6o8_0(.dout(w_dff_A_MyMyPt571_0),.din(w_dff_A_iLufhf6o8_0),.clk(gclk));
	jdff dff_A_MyMyPt571_0(.dout(w_dff_A_tRzYee8n4_0),.din(w_dff_A_MyMyPt571_0),.clk(gclk));
	jdff dff_A_tRzYee8n4_0(.dout(w_dff_A_iYOAAS3t5_0),.din(w_dff_A_tRzYee8n4_0),.clk(gclk));
	jdff dff_A_iYOAAS3t5_0(.dout(w_dff_A_B8MDTUpb8_0),.din(w_dff_A_iYOAAS3t5_0),.clk(gclk));
	jdff dff_A_B8MDTUpb8_0(.dout(w_dff_A_IfozyU0f6_0),.din(w_dff_A_B8MDTUpb8_0),.clk(gclk));
	jdff dff_A_IfozyU0f6_0(.dout(w_dff_A_TeAQgpvl3_0),.din(w_dff_A_IfozyU0f6_0),.clk(gclk));
	jdff dff_A_TeAQgpvl3_0(.dout(w_dff_A_N8imk39S0_0),.din(w_dff_A_TeAQgpvl3_0),.clk(gclk));
	jdff dff_A_N8imk39S0_0(.dout(w_dff_A_SFT6a6JL3_0),.din(w_dff_A_N8imk39S0_0),.clk(gclk));
	jdff dff_A_SFT6a6JL3_0(.dout(w_dff_A_z2m4hU9P3_0),.din(w_dff_A_SFT6a6JL3_0),.clk(gclk));
	jdff dff_A_z2m4hU9P3_0(.dout(w_dff_A_zfpi0cDF6_0),.din(w_dff_A_z2m4hU9P3_0),.clk(gclk));
	jdff dff_A_zfpi0cDF6_0(.dout(w_dff_A_vG7Wtfqb2_0),.din(w_dff_A_zfpi0cDF6_0),.clk(gclk));
	jdff dff_A_vG7Wtfqb2_0(.dout(w_dff_A_Q6MQmU7a3_0),.din(w_dff_A_vG7Wtfqb2_0),.clk(gclk));
	jdff dff_A_Q6MQmU7a3_0(.dout(w_dff_A_kqxinkmM3_0),.din(w_dff_A_Q6MQmU7a3_0),.clk(gclk));
	jdff dff_A_kqxinkmM3_0(.dout(w_dff_A_27Y7HHIo6_0),.din(w_dff_A_kqxinkmM3_0),.clk(gclk));
	jdff dff_A_27Y7HHIo6_0(.dout(w_dff_A_GxAGMbpU9_0),.din(w_dff_A_27Y7HHIo6_0),.clk(gclk));
	jdff dff_A_GxAGMbpU9_0(.dout(w_dff_A_6mZaMQ2u8_0),.din(w_dff_A_GxAGMbpU9_0),.clk(gclk));
	jdff dff_A_6mZaMQ2u8_0(.dout(w_dff_A_OPV7AuyA9_0),.din(w_dff_A_6mZaMQ2u8_0),.clk(gclk));
	jdff dff_A_OPV7AuyA9_0(.dout(w_dff_A_Mvev92x47_0),.din(w_dff_A_OPV7AuyA9_0),.clk(gclk));
	jdff dff_A_Mvev92x47_0(.dout(w_dff_A_FSH3reNl4_0),.din(w_dff_A_Mvev92x47_0),.clk(gclk));
	jdff dff_A_FSH3reNl4_0(.dout(w_dff_A_LxDiXIh96_0),.din(w_dff_A_FSH3reNl4_0),.clk(gclk));
	jdff dff_A_LxDiXIh96_0(.dout(w_dff_A_mRkKIUyw0_0),.din(w_dff_A_LxDiXIh96_0),.clk(gclk));
	jdff dff_A_mRkKIUyw0_0(.dout(w_dff_A_4heoCdeK5_0),.din(w_dff_A_mRkKIUyw0_0),.clk(gclk));
	jdff dff_A_4heoCdeK5_0(.dout(w_dff_A_NrVXIPUz6_0),.din(w_dff_A_4heoCdeK5_0),.clk(gclk));
	jdff dff_A_NrVXIPUz6_0(.dout(w_dff_A_yDjtFI9Y3_0),.din(w_dff_A_NrVXIPUz6_0),.clk(gclk));
	jdff dff_A_yDjtFI9Y3_0(.dout(w_dff_A_1Bt2Y9695_0),.din(w_dff_A_yDjtFI9Y3_0),.clk(gclk));
	jdff dff_A_1Bt2Y9695_0(.dout(w_dff_A_U3ZrDMSm2_0),.din(w_dff_A_1Bt2Y9695_0),.clk(gclk));
	jdff dff_A_U3ZrDMSm2_0(.dout(w_dff_A_9yc2b15b4_0),.din(w_dff_A_U3ZrDMSm2_0),.clk(gclk));
	jdff dff_A_9yc2b15b4_0(.dout(w_dff_A_6mwv8tLa6_0),.din(w_dff_A_9yc2b15b4_0),.clk(gclk));
	jdff dff_A_6mwv8tLa6_0(.dout(f3),.din(w_dff_A_6mwv8tLa6_0),.clk(gclk));
	jdff dff_A_1VQG7qnR4_2(.dout(w_dff_A_5Fa9cNUP9_0),.din(w_dff_A_1VQG7qnR4_2),.clk(gclk));
	jdff dff_A_5Fa9cNUP9_0(.dout(w_dff_A_XszYuBZn6_0),.din(w_dff_A_5Fa9cNUP9_0),.clk(gclk));
	jdff dff_A_XszYuBZn6_0(.dout(w_dff_A_rYDI6ieU0_0),.din(w_dff_A_XszYuBZn6_0),.clk(gclk));
	jdff dff_A_rYDI6ieU0_0(.dout(w_dff_A_Mb7TeTvB7_0),.din(w_dff_A_rYDI6ieU0_0),.clk(gclk));
	jdff dff_A_Mb7TeTvB7_0(.dout(w_dff_A_7oPnku5t2_0),.din(w_dff_A_Mb7TeTvB7_0),.clk(gclk));
	jdff dff_A_7oPnku5t2_0(.dout(w_dff_A_zXBJKvOz5_0),.din(w_dff_A_7oPnku5t2_0),.clk(gclk));
	jdff dff_A_zXBJKvOz5_0(.dout(w_dff_A_L0Frk5Ii6_0),.din(w_dff_A_zXBJKvOz5_0),.clk(gclk));
	jdff dff_A_L0Frk5Ii6_0(.dout(w_dff_A_uumZ1lpo8_0),.din(w_dff_A_L0Frk5Ii6_0),.clk(gclk));
	jdff dff_A_uumZ1lpo8_0(.dout(w_dff_A_7xBWhwoN9_0),.din(w_dff_A_uumZ1lpo8_0),.clk(gclk));
	jdff dff_A_7xBWhwoN9_0(.dout(w_dff_A_ZkF2pzgP4_0),.din(w_dff_A_7xBWhwoN9_0),.clk(gclk));
	jdff dff_A_ZkF2pzgP4_0(.dout(w_dff_A_iNMcl5751_0),.din(w_dff_A_ZkF2pzgP4_0),.clk(gclk));
	jdff dff_A_iNMcl5751_0(.dout(w_dff_A_25m6uuBK2_0),.din(w_dff_A_iNMcl5751_0),.clk(gclk));
	jdff dff_A_25m6uuBK2_0(.dout(w_dff_A_jH9p5tME8_0),.din(w_dff_A_25m6uuBK2_0),.clk(gclk));
	jdff dff_A_jH9p5tME8_0(.dout(w_dff_A_FoMYKH7m5_0),.din(w_dff_A_jH9p5tME8_0),.clk(gclk));
	jdff dff_A_FoMYKH7m5_0(.dout(w_dff_A_QMiARZyX8_0),.din(w_dff_A_FoMYKH7m5_0),.clk(gclk));
	jdff dff_A_QMiARZyX8_0(.dout(w_dff_A_5a6wVnjT2_0),.din(w_dff_A_QMiARZyX8_0),.clk(gclk));
	jdff dff_A_5a6wVnjT2_0(.dout(w_dff_A_HjFceiDg1_0),.din(w_dff_A_5a6wVnjT2_0),.clk(gclk));
	jdff dff_A_HjFceiDg1_0(.dout(w_dff_A_77u0j4Uq4_0),.din(w_dff_A_HjFceiDg1_0),.clk(gclk));
	jdff dff_A_77u0j4Uq4_0(.dout(w_dff_A_sICGys189_0),.din(w_dff_A_77u0j4Uq4_0),.clk(gclk));
	jdff dff_A_sICGys189_0(.dout(w_dff_A_8WD7kccW5_0),.din(w_dff_A_sICGys189_0),.clk(gclk));
	jdff dff_A_8WD7kccW5_0(.dout(w_dff_A_XPVG3QX59_0),.din(w_dff_A_8WD7kccW5_0),.clk(gclk));
	jdff dff_A_XPVG3QX59_0(.dout(w_dff_A_5xDpoGie3_0),.din(w_dff_A_XPVG3QX59_0),.clk(gclk));
	jdff dff_A_5xDpoGie3_0(.dout(w_dff_A_fDdvouAS8_0),.din(w_dff_A_5xDpoGie3_0),.clk(gclk));
	jdff dff_A_fDdvouAS8_0(.dout(w_dff_A_CX8XH9k80_0),.din(w_dff_A_fDdvouAS8_0),.clk(gclk));
	jdff dff_A_CX8XH9k80_0(.dout(w_dff_A_wWsff6kH7_0),.din(w_dff_A_CX8XH9k80_0),.clk(gclk));
	jdff dff_A_wWsff6kH7_0(.dout(w_dff_A_tyOQC1gb4_0),.din(w_dff_A_wWsff6kH7_0),.clk(gclk));
	jdff dff_A_tyOQC1gb4_0(.dout(w_dff_A_JOM0hDP27_0),.din(w_dff_A_tyOQC1gb4_0),.clk(gclk));
	jdff dff_A_JOM0hDP27_0(.dout(w_dff_A_VxOcX4fM4_0),.din(w_dff_A_JOM0hDP27_0),.clk(gclk));
	jdff dff_A_VxOcX4fM4_0(.dout(w_dff_A_9XJ5I31a5_0),.din(w_dff_A_VxOcX4fM4_0),.clk(gclk));
	jdff dff_A_9XJ5I31a5_0(.dout(w_dff_A_vNiNP8Ud7_0),.din(w_dff_A_9XJ5I31a5_0),.clk(gclk));
	jdff dff_A_vNiNP8Ud7_0(.dout(w_dff_A_iFD7q3yd1_0),.din(w_dff_A_vNiNP8Ud7_0),.clk(gclk));
	jdff dff_A_iFD7q3yd1_0(.dout(w_dff_A_9lFpBAUQ4_0),.din(w_dff_A_iFD7q3yd1_0),.clk(gclk));
	jdff dff_A_9lFpBAUQ4_0(.dout(w_dff_A_j4kMoJ2N8_0),.din(w_dff_A_9lFpBAUQ4_0),.clk(gclk));
	jdff dff_A_j4kMoJ2N8_0(.dout(w_dff_A_koYqHtAr5_0),.din(w_dff_A_j4kMoJ2N8_0),.clk(gclk));
	jdff dff_A_koYqHtAr5_0(.dout(w_dff_A_j6EMyffI1_0),.din(w_dff_A_koYqHtAr5_0),.clk(gclk));
	jdff dff_A_j6EMyffI1_0(.dout(w_dff_A_deUhHxrn3_0),.din(w_dff_A_j6EMyffI1_0),.clk(gclk));
	jdff dff_A_deUhHxrn3_0(.dout(w_dff_A_iYXB5tPh6_0),.din(w_dff_A_deUhHxrn3_0),.clk(gclk));
	jdff dff_A_iYXB5tPh6_0(.dout(w_dff_A_jRDIlC7w5_0),.din(w_dff_A_iYXB5tPh6_0),.clk(gclk));
	jdff dff_A_jRDIlC7w5_0(.dout(w_dff_A_X1yj2HMP6_0),.din(w_dff_A_jRDIlC7w5_0),.clk(gclk));
	jdff dff_A_X1yj2HMP6_0(.dout(w_dff_A_J0VsU88V9_0),.din(w_dff_A_X1yj2HMP6_0),.clk(gclk));
	jdff dff_A_J0VsU88V9_0(.dout(w_dff_A_UJPKrkUT0_0),.din(w_dff_A_J0VsU88V9_0),.clk(gclk));
	jdff dff_A_UJPKrkUT0_0(.dout(w_dff_A_l0OsOiUk9_0),.din(w_dff_A_UJPKrkUT0_0),.clk(gclk));
	jdff dff_A_l0OsOiUk9_0(.dout(w_dff_A_Y7gaWkRM9_0),.din(w_dff_A_l0OsOiUk9_0),.clk(gclk));
	jdff dff_A_Y7gaWkRM9_0(.dout(w_dff_A_XgrdThwL7_0),.din(w_dff_A_Y7gaWkRM9_0),.clk(gclk));
	jdff dff_A_XgrdThwL7_0(.dout(w_dff_A_zukOVIFp0_0),.din(w_dff_A_XgrdThwL7_0),.clk(gclk));
	jdff dff_A_zukOVIFp0_0(.dout(w_dff_A_aMkd7sWD0_0),.din(w_dff_A_zukOVIFp0_0),.clk(gclk));
	jdff dff_A_aMkd7sWD0_0(.dout(w_dff_A_ynriJyoJ2_0),.din(w_dff_A_aMkd7sWD0_0),.clk(gclk));
	jdff dff_A_ynriJyoJ2_0(.dout(w_dff_A_JselGAOv0_0),.din(w_dff_A_ynriJyoJ2_0),.clk(gclk));
	jdff dff_A_JselGAOv0_0(.dout(w_dff_A_dhQ5W5hO5_0),.din(w_dff_A_JselGAOv0_0),.clk(gclk));
	jdff dff_A_dhQ5W5hO5_0(.dout(w_dff_A_3fFDjsAL8_0),.din(w_dff_A_dhQ5W5hO5_0),.clk(gclk));
	jdff dff_A_3fFDjsAL8_0(.dout(w_dff_A_2KmSNbko8_0),.din(w_dff_A_3fFDjsAL8_0),.clk(gclk));
	jdff dff_A_2KmSNbko8_0(.dout(w_dff_A_2ubffZrC5_0),.din(w_dff_A_2KmSNbko8_0),.clk(gclk));
	jdff dff_A_2ubffZrC5_0(.dout(w_dff_A_b2XEM6J21_0),.din(w_dff_A_2ubffZrC5_0),.clk(gclk));
	jdff dff_A_b2XEM6J21_0(.dout(w_dff_A_lqauPCNQ4_0),.din(w_dff_A_b2XEM6J21_0),.clk(gclk));
	jdff dff_A_lqauPCNQ4_0(.dout(w_dff_A_RLWv6Flx1_0),.din(w_dff_A_lqauPCNQ4_0),.clk(gclk));
	jdff dff_A_RLWv6Flx1_0(.dout(w_dff_A_ZUVhd7L38_0),.din(w_dff_A_RLWv6Flx1_0),.clk(gclk));
	jdff dff_A_ZUVhd7L38_0(.dout(w_dff_A_IejkbUIe2_0),.din(w_dff_A_ZUVhd7L38_0),.clk(gclk));
	jdff dff_A_IejkbUIe2_0(.dout(w_dff_A_wIRfZAe26_0),.din(w_dff_A_IejkbUIe2_0),.clk(gclk));
	jdff dff_A_wIRfZAe26_0(.dout(w_dff_A_IzkQeg2s2_0),.din(w_dff_A_wIRfZAe26_0),.clk(gclk));
	jdff dff_A_IzkQeg2s2_0(.dout(w_dff_A_N9cHApKK5_0),.din(w_dff_A_IzkQeg2s2_0),.clk(gclk));
	jdff dff_A_N9cHApKK5_0(.dout(w_dff_A_IhvCVoOx3_0),.din(w_dff_A_N9cHApKK5_0),.clk(gclk));
	jdff dff_A_IhvCVoOx3_0(.dout(w_dff_A_rWO4psWV7_0),.din(w_dff_A_IhvCVoOx3_0),.clk(gclk));
	jdff dff_A_rWO4psWV7_0(.dout(w_dff_A_mgZclAPZ3_0),.din(w_dff_A_rWO4psWV7_0),.clk(gclk));
	jdff dff_A_mgZclAPZ3_0(.dout(w_dff_A_y43MHAER3_0),.din(w_dff_A_mgZclAPZ3_0),.clk(gclk));
	jdff dff_A_y43MHAER3_0(.dout(w_dff_A_cnBx4Qn79_0),.din(w_dff_A_y43MHAER3_0),.clk(gclk));
	jdff dff_A_cnBx4Qn79_0(.dout(w_dff_A_6upFUy2T4_0),.din(w_dff_A_cnBx4Qn79_0),.clk(gclk));
	jdff dff_A_6upFUy2T4_0(.dout(w_dff_A_ab4oi3PL5_0),.din(w_dff_A_6upFUy2T4_0),.clk(gclk));
	jdff dff_A_ab4oi3PL5_0(.dout(w_dff_A_No1HjYZc6_0),.din(w_dff_A_ab4oi3PL5_0),.clk(gclk));
	jdff dff_A_No1HjYZc6_0(.dout(w_dff_A_BrZnQq3L7_0),.din(w_dff_A_No1HjYZc6_0),.clk(gclk));
	jdff dff_A_BrZnQq3L7_0(.dout(w_dff_A_NyZpidZa7_0),.din(w_dff_A_BrZnQq3L7_0),.clk(gclk));
	jdff dff_A_NyZpidZa7_0(.dout(w_dff_A_PZvrJR4n4_0),.din(w_dff_A_NyZpidZa7_0),.clk(gclk));
	jdff dff_A_PZvrJR4n4_0(.dout(w_dff_A_TzN4dReA4_0),.din(w_dff_A_PZvrJR4n4_0),.clk(gclk));
	jdff dff_A_TzN4dReA4_0(.dout(w_dff_A_HFSgiQ2O8_0),.din(w_dff_A_TzN4dReA4_0),.clk(gclk));
	jdff dff_A_HFSgiQ2O8_0(.dout(w_dff_A_Rk5annqX2_0),.din(w_dff_A_HFSgiQ2O8_0),.clk(gclk));
	jdff dff_A_Rk5annqX2_0(.dout(w_dff_A_MThSq39d1_0),.din(w_dff_A_Rk5annqX2_0),.clk(gclk));
	jdff dff_A_MThSq39d1_0(.dout(w_dff_A_loObXrDX8_0),.din(w_dff_A_MThSq39d1_0),.clk(gclk));
	jdff dff_A_loObXrDX8_0(.dout(w_dff_A_Re12mYPe0_0),.din(w_dff_A_loObXrDX8_0),.clk(gclk));
	jdff dff_A_Re12mYPe0_0(.dout(w_dff_A_sbmHq4qd3_0),.din(w_dff_A_Re12mYPe0_0),.clk(gclk));
	jdff dff_A_sbmHq4qd3_0(.dout(w_dff_A_GacHLWK03_0),.din(w_dff_A_sbmHq4qd3_0),.clk(gclk));
	jdff dff_A_GacHLWK03_0(.dout(w_dff_A_Rqd5EoRH3_0),.din(w_dff_A_GacHLWK03_0),.clk(gclk));
	jdff dff_A_Rqd5EoRH3_0(.dout(w_dff_A_VRTcxhZo9_0),.din(w_dff_A_Rqd5EoRH3_0),.clk(gclk));
	jdff dff_A_VRTcxhZo9_0(.dout(w_dff_A_mXfj60WY4_0),.din(w_dff_A_VRTcxhZo9_0),.clk(gclk));
	jdff dff_A_mXfj60WY4_0(.dout(w_dff_A_AGYcJ9yt6_0),.din(w_dff_A_mXfj60WY4_0),.clk(gclk));
	jdff dff_A_AGYcJ9yt6_0(.dout(w_dff_A_g5sCEzc00_0),.din(w_dff_A_AGYcJ9yt6_0),.clk(gclk));
	jdff dff_A_g5sCEzc00_0(.dout(w_dff_A_662Q5HJj8_0),.din(w_dff_A_g5sCEzc00_0),.clk(gclk));
	jdff dff_A_662Q5HJj8_0(.dout(w_dff_A_wMkIaqNk1_0),.din(w_dff_A_662Q5HJj8_0),.clk(gclk));
	jdff dff_A_wMkIaqNk1_0(.dout(w_dff_A_pYKCuL1D1_0),.din(w_dff_A_wMkIaqNk1_0),.clk(gclk));
	jdff dff_A_pYKCuL1D1_0(.dout(w_dff_A_OtkchGOg2_0),.din(w_dff_A_pYKCuL1D1_0),.clk(gclk));
	jdff dff_A_OtkchGOg2_0(.dout(w_dff_A_GteGHVar9_0),.din(w_dff_A_OtkchGOg2_0),.clk(gclk));
	jdff dff_A_GteGHVar9_0(.dout(w_dff_A_ewLSiq3B8_0),.din(w_dff_A_GteGHVar9_0),.clk(gclk));
	jdff dff_A_ewLSiq3B8_0(.dout(w_dff_A_DBsiDWtA6_0),.din(w_dff_A_ewLSiq3B8_0),.clk(gclk));
	jdff dff_A_DBsiDWtA6_0(.dout(w_dff_A_x2X0pvH39_0),.din(w_dff_A_DBsiDWtA6_0),.clk(gclk));
	jdff dff_A_x2X0pvH39_0(.dout(w_dff_A_y1iJf8Sb3_0),.din(w_dff_A_x2X0pvH39_0),.clk(gclk));
	jdff dff_A_y1iJf8Sb3_0(.dout(w_dff_A_J9sa2Ghz4_0),.din(w_dff_A_y1iJf8Sb3_0),.clk(gclk));
	jdff dff_A_J9sa2Ghz4_0(.dout(w_dff_A_SVoKgd9P2_0),.din(w_dff_A_J9sa2Ghz4_0),.clk(gclk));
	jdff dff_A_SVoKgd9P2_0(.dout(w_dff_A_h3Bnk4hO7_0),.din(w_dff_A_SVoKgd9P2_0),.clk(gclk));
	jdff dff_A_h3Bnk4hO7_0(.dout(w_dff_A_mBo9V4g62_0),.din(w_dff_A_h3Bnk4hO7_0),.clk(gclk));
	jdff dff_A_mBo9V4g62_0(.dout(w_dff_A_eEd3ROE53_0),.din(w_dff_A_mBo9V4g62_0),.clk(gclk));
	jdff dff_A_eEd3ROE53_0(.dout(w_dff_A_yZK3LxT81_0),.din(w_dff_A_eEd3ROE53_0),.clk(gclk));
	jdff dff_A_yZK3LxT81_0(.dout(w_dff_A_JXfeZ7db4_0),.din(w_dff_A_yZK3LxT81_0),.clk(gclk));
	jdff dff_A_JXfeZ7db4_0(.dout(w_dff_A_Xb6kUgQI5_0),.din(w_dff_A_JXfeZ7db4_0),.clk(gclk));
	jdff dff_A_Xb6kUgQI5_0(.dout(w_dff_A_WL7gqoW80_0),.din(w_dff_A_Xb6kUgQI5_0),.clk(gclk));
	jdff dff_A_WL7gqoW80_0(.dout(w_dff_A_e8WV26aU0_0),.din(w_dff_A_WL7gqoW80_0),.clk(gclk));
	jdff dff_A_e8WV26aU0_0(.dout(w_dff_A_00jNVlvt5_0),.din(w_dff_A_e8WV26aU0_0),.clk(gclk));
	jdff dff_A_00jNVlvt5_0(.dout(w_dff_A_GUGBYtzZ5_0),.din(w_dff_A_00jNVlvt5_0),.clk(gclk));
	jdff dff_A_GUGBYtzZ5_0(.dout(w_dff_A_i41Ga4qU9_0),.din(w_dff_A_GUGBYtzZ5_0),.clk(gclk));
	jdff dff_A_i41Ga4qU9_0(.dout(w_dff_A_XBBCXx695_0),.din(w_dff_A_i41Ga4qU9_0),.clk(gclk));
	jdff dff_A_XBBCXx695_0(.dout(w_dff_A_Qe5cWNkw4_0),.din(w_dff_A_XBBCXx695_0),.clk(gclk));
	jdff dff_A_Qe5cWNkw4_0(.dout(w_dff_A_6Flh009Z9_0),.din(w_dff_A_Qe5cWNkw4_0),.clk(gclk));
	jdff dff_A_6Flh009Z9_0(.dout(w_dff_A_E4APkXAG5_0),.din(w_dff_A_6Flh009Z9_0),.clk(gclk));
	jdff dff_A_E4APkXAG5_0(.dout(w_dff_A_asgeTDbE9_0),.din(w_dff_A_E4APkXAG5_0),.clk(gclk));
	jdff dff_A_asgeTDbE9_0(.dout(w_dff_A_UxgsX2GP6_0),.din(w_dff_A_asgeTDbE9_0),.clk(gclk));
	jdff dff_A_UxgsX2GP6_0(.dout(w_dff_A_ZT6miqI60_0),.din(w_dff_A_UxgsX2GP6_0),.clk(gclk));
	jdff dff_A_ZT6miqI60_0(.dout(w_dff_A_aSIs1bdk3_0),.din(w_dff_A_ZT6miqI60_0),.clk(gclk));
	jdff dff_A_aSIs1bdk3_0(.dout(w_dff_A_MV6fgJqE2_0),.din(w_dff_A_aSIs1bdk3_0),.clk(gclk));
	jdff dff_A_MV6fgJqE2_0(.dout(w_dff_A_0JsU6p5D3_0),.din(w_dff_A_MV6fgJqE2_0),.clk(gclk));
	jdff dff_A_0JsU6p5D3_0(.dout(w_dff_A_t2Ktl2Mx2_0),.din(w_dff_A_0JsU6p5D3_0),.clk(gclk));
	jdff dff_A_t2Ktl2Mx2_0(.dout(w_dff_A_MM7DwEUX2_0),.din(w_dff_A_t2Ktl2Mx2_0),.clk(gclk));
	jdff dff_A_MM7DwEUX2_0(.dout(w_dff_A_THFzVDnS6_0),.din(w_dff_A_MM7DwEUX2_0),.clk(gclk));
	jdff dff_A_THFzVDnS6_0(.dout(w_dff_A_3Qz4fLsn5_0),.din(w_dff_A_THFzVDnS6_0),.clk(gclk));
	jdff dff_A_3Qz4fLsn5_0(.dout(w_dff_A_Q0j0c46J3_0),.din(w_dff_A_3Qz4fLsn5_0),.clk(gclk));
	jdff dff_A_Q0j0c46J3_0(.dout(w_dff_A_IuqKgyK03_0),.din(w_dff_A_Q0j0c46J3_0),.clk(gclk));
	jdff dff_A_IuqKgyK03_0(.dout(f4),.din(w_dff_A_IuqKgyK03_0),.clk(gclk));
	jdff dff_A_IdkFl4Xp4_2(.dout(w_dff_A_7WOSKiuK6_0),.din(w_dff_A_IdkFl4Xp4_2),.clk(gclk));
	jdff dff_A_7WOSKiuK6_0(.dout(w_dff_A_whqaaO4I3_0),.din(w_dff_A_7WOSKiuK6_0),.clk(gclk));
	jdff dff_A_whqaaO4I3_0(.dout(w_dff_A_dWZmbI9c4_0),.din(w_dff_A_whqaaO4I3_0),.clk(gclk));
	jdff dff_A_dWZmbI9c4_0(.dout(w_dff_A_cLSxEBWv5_0),.din(w_dff_A_dWZmbI9c4_0),.clk(gclk));
	jdff dff_A_cLSxEBWv5_0(.dout(w_dff_A_js64y1LC4_0),.din(w_dff_A_cLSxEBWv5_0),.clk(gclk));
	jdff dff_A_js64y1LC4_0(.dout(w_dff_A_LmWZIKY74_0),.din(w_dff_A_js64y1LC4_0),.clk(gclk));
	jdff dff_A_LmWZIKY74_0(.dout(w_dff_A_0lvHdkUq6_0),.din(w_dff_A_LmWZIKY74_0),.clk(gclk));
	jdff dff_A_0lvHdkUq6_0(.dout(w_dff_A_k1VAt9Tt4_0),.din(w_dff_A_0lvHdkUq6_0),.clk(gclk));
	jdff dff_A_k1VAt9Tt4_0(.dout(w_dff_A_68DsUUIw2_0),.din(w_dff_A_k1VAt9Tt4_0),.clk(gclk));
	jdff dff_A_68DsUUIw2_0(.dout(w_dff_A_ZZVkgg8w2_0),.din(w_dff_A_68DsUUIw2_0),.clk(gclk));
	jdff dff_A_ZZVkgg8w2_0(.dout(w_dff_A_FYyBu26T7_0),.din(w_dff_A_ZZVkgg8w2_0),.clk(gclk));
	jdff dff_A_FYyBu26T7_0(.dout(w_dff_A_6ZGFAdw08_0),.din(w_dff_A_FYyBu26T7_0),.clk(gclk));
	jdff dff_A_6ZGFAdw08_0(.dout(w_dff_A_FYqQvUoA1_0),.din(w_dff_A_6ZGFAdw08_0),.clk(gclk));
	jdff dff_A_FYqQvUoA1_0(.dout(w_dff_A_NI6BFi2u9_0),.din(w_dff_A_FYqQvUoA1_0),.clk(gclk));
	jdff dff_A_NI6BFi2u9_0(.dout(w_dff_A_M1XSP2in8_0),.din(w_dff_A_NI6BFi2u9_0),.clk(gclk));
	jdff dff_A_M1XSP2in8_0(.dout(w_dff_A_CkbEmAKk1_0),.din(w_dff_A_M1XSP2in8_0),.clk(gclk));
	jdff dff_A_CkbEmAKk1_0(.dout(w_dff_A_Wtm3Bdwb3_0),.din(w_dff_A_CkbEmAKk1_0),.clk(gclk));
	jdff dff_A_Wtm3Bdwb3_0(.dout(w_dff_A_4RlHqDPm5_0),.din(w_dff_A_Wtm3Bdwb3_0),.clk(gclk));
	jdff dff_A_4RlHqDPm5_0(.dout(w_dff_A_WCIIhXIK5_0),.din(w_dff_A_4RlHqDPm5_0),.clk(gclk));
	jdff dff_A_WCIIhXIK5_0(.dout(w_dff_A_mzThEMH35_0),.din(w_dff_A_WCIIhXIK5_0),.clk(gclk));
	jdff dff_A_mzThEMH35_0(.dout(w_dff_A_RdHcBSkH5_0),.din(w_dff_A_mzThEMH35_0),.clk(gclk));
	jdff dff_A_RdHcBSkH5_0(.dout(w_dff_A_dCB1WaR64_0),.din(w_dff_A_RdHcBSkH5_0),.clk(gclk));
	jdff dff_A_dCB1WaR64_0(.dout(w_dff_A_KuwRXycy1_0),.din(w_dff_A_dCB1WaR64_0),.clk(gclk));
	jdff dff_A_KuwRXycy1_0(.dout(w_dff_A_ydza07DE2_0),.din(w_dff_A_KuwRXycy1_0),.clk(gclk));
	jdff dff_A_ydza07DE2_0(.dout(w_dff_A_imZOv0kF7_0),.din(w_dff_A_ydza07DE2_0),.clk(gclk));
	jdff dff_A_imZOv0kF7_0(.dout(w_dff_A_2j8Kcy691_0),.din(w_dff_A_imZOv0kF7_0),.clk(gclk));
	jdff dff_A_2j8Kcy691_0(.dout(w_dff_A_FaqfAlgy0_0),.din(w_dff_A_2j8Kcy691_0),.clk(gclk));
	jdff dff_A_FaqfAlgy0_0(.dout(w_dff_A_YggbqMBl2_0),.din(w_dff_A_FaqfAlgy0_0),.clk(gclk));
	jdff dff_A_YggbqMBl2_0(.dout(w_dff_A_8kmZQxlg9_0),.din(w_dff_A_YggbqMBl2_0),.clk(gclk));
	jdff dff_A_8kmZQxlg9_0(.dout(w_dff_A_AmeYctPz0_0),.din(w_dff_A_8kmZQxlg9_0),.clk(gclk));
	jdff dff_A_AmeYctPz0_0(.dout(w_dff_A_BCkLTDGX2_0),.din(w_dff_A_AmeYctPz0_0),.clk(gclk));
	jdff dff_A_BCkLTDGX2_0(.dout(w_dff_A_wn8ICb4d3_0),.din(w_dff_A_BCkLTDGX2_0),.clk(gclk));
	jdff dff_A_wn8ICb4d3_0(.dout(w_dff_A_0DNGrGX60_0),.din(w_dff_A_wn8ICb4d3_0),.clk(gclk));
	jdff dff_A_0DNGrGX60_0(.dout(w_dff_A_KkoH3SFT0_0),.din(w_dff_A_0DNGrGX60_0),.clk(gclk));
	jdff dff_A_KkoH3SFT0_0(.dout(w_dff_A_K0V2sZl95_0),.din(w_dff_A_KkoH3SFT0_0),.clk(gclk));
	jdff dff_A_K0V2sZl95_0(.dout(w_dff_A_b64RPAkx2_0),.din(w_dff_A_K0V2sZl95_0),.clk(gclk));
	jdff dff_A_b64RPAkx2_0(.dout(w_dff_A_i8Bw4ziX8_0),.din(w_dff_A_b64RPAkx2_0),.clk(gclk));
	jdff dff_A_i8Bw4ziX8_0(.dout(w_dff_A_LynwnBL54_0),.din(w_dff_A_i8Bw4ziX8_0),.clk(gclk));
	jdff dff_A_LynwnBL54_0(.dout(w_dff_A_pbUMnuaJ6_0),.din(w_dff_A_LynwnBL54_0),.clk(gclk));
	jdff dff_A_pbUMnuaJ6_0(.dout(w_dff_A_eenawJlp6_0),.din(w_dff_A_pbUMnuaJ6_0),.clk(gclk));
	jdff dff_A_eenawJlp6_0(.dout(w_dff_A_h68K7PFM5_0),.din(w_dff_A_eenawJlp6_0),.clk(gclk));
	jdff dff_A_h68K7PFM5_0(.dout(w_dff_A_MM1znDoQ2_0),.din(w_dff_A_h68K7PFM5_0),.clk(gclk));
	jdff dff_A_MM1znDoQ2_0(.dout(w_dff_A_wQnt1osF4_0),.din(w_dff_A_MM1znDoQ2_0),.clk(gclk));
	jdff dff_A_wQnt1osF4_0(.dout(w_dff_A_jBqP9Rno1_0),.din(w_dff_A_wQnt1osF4_0),.clk(gclk));
	jdff dff_A_jBqP9Rno1_0(.dout(w_dff_A_6SPblfPN8_0),.din(w_dff_A_jBqP9Rno1_0),.clk(gclk));
	jdff dff_A_6SPblfPN8_0(.dout(w_dff_A_Q4FfvqYs8_0),.din(w_dff_A_6SPblfPN8_0),.clk(gclk));
	jdff dff_A_Q4FfvqYs8_0(.dout(w_dff_A_MdaOHuhM2_0),.din(w_dff_A_Q4FfvqYs8_0),.clk(gclk));
	jdff dff_A_MdaOHuhM2_0(.dout(w_dff_A_yT3Zyqar2_0),.din(w_dff_A_MdaOHuhM2_0),.clk(gclk));
	jdff dff_A_yT3Zyqar2_0(.dout(w_dff_A_JBeftkVZ9_0),.din(w_dff_A_yT3Zyqar2_0),.clk(gclk));
	jdff dff_A_JBeftkVZ9_0(.dout(w_dff_A_80DNT7ja4_0),.din(w_dff_A_JBeftkVZ9_0),.clk(gclk));
	jdff dff_A_80DNT7ja4_0(.dout(w_dff_A_aYGx0Sx09_0),.din(w_dff_A_80DNT7ja4_0),.clk(gclk));
	jdff dff_A_aYGx0Sx09_0(.dout(w_dff_A_Za84DtOn4_0),.din(w_dff_A_aYGx0Sx09_0),.clk(gclk));
	jdff dff_A_Za84DtOn4_0(.dout(w_dff_A_CAfnn6Ln6_0),.din(w_dff_A_Za84DtOn4_0),.clk(gclk));
	jdff dff_A_CAfnn6Ln6_0(.dout(w_dff_A_iX3mfOFH4_0),.din(w_dff_A_CAfnn6Ln6_0),.clk(gclk));
	jdff dff_A_iX3mfOFH4_0(.dout(w_dff_A_GIAv927z8_0),.din(w_dff_A_iX3mfOFH4_0),.clk(gclk));
	jdff dff_A_GIAv927z8_0(.dout(w_dff_A_GJeHbi3J5_0),.din(w_dff_A_GIAv927z8_0),.clk(gclk));
	jdff dff_A_GJeHbi3J5_0(.dout(w_dff_A_AVEVBteC2_0),.din(w_dff_A_GJeHbi3J5_0),.clk(gclk));
	jdff dff_A_AVEVBteC2_0(.dout(w_dff_A_3owZC4ri1_0),.din(w_dff_A_AVEVBteC2_0),.clk(gclk));
	jdff dff_A_3owZC4ri1_0(.dout(w_dff_A_fsC9gKLw2_0),.din(w_dff_A_3owZC4ri1_0),.clk(gclk));
	jdff dff_A_fsC9gKLw2_0(.dout(w_dff_A_EWpfq3hw8_0),.din(w_dff_A_fsC9gKLw2_0),.clk(gclk));
	jdff dff_A_EWpfq3hw8_0(.dout(w_dff_A_qk84iQld3_0),.din(w_dff_A_EWpfq3hw8_0),.clk(gclk));
	jdff dff_A_qk84iQld3_0(.dout(w_dff_A_Wu21gRUj5_0),.din(w_dff_A_qk84iQld3_0),.clk(gclk));
	jdff dff_A_Wu21gRUj5_0(.dout(w_dff_A_0GjjQOdK3_0),.din(w_dff_A_Wu21gRUj5_0),.clk(gclk));
	jdff dff_A_0GjjQOdK3_0(.dout(w_dff_A_ug4j69FI0_0),.din(w_dff_A_0GjjQOdK3_0),.clk(gclk));
	jdff dff_A_ug4j69FI0_0(.dout(w_dff_A_fCZfGh1d4_0),.din(w_dff_A_ug4j69FI0_0),.clk(gclk));
	jdff dff_A_fCZfGh1d4_0(.dout(w_dff_A_NWCLG5AO6_0),.din(w_dff_A_fCZfGh1d4_0),.clk(gclk));
	jdff dff_A_NWCLG5AO6_0(.dout(w_dff_A_2ktIlevG8_0),.din(w_dff_A_NWCLG5AO6_0),.clk(gclk));
	jdff dff_A_2ktIlevG8_0(.dout(w_dff_A_ueVTdPtx1_0),.din(w_dff_A_2ktIlevG8_0),.clk(gclk));
	jdff dff_A_ueVTdPtx1_0(.dout(w_dff_A_LSNEDSnm8_0),.din(w_dff_A_ueVTdPtx1_0),.clk(gclk));
	jdff dff_A_LSNEDSnm8_0(.dout(w_dff_A_5xGXelTX6_0),.din(w_dff_A_LSNEDSnm8_0),.clk(gclk));
	jdff dff_A_5xGXelTX6_0(.dout(w_dff_A_bghyKuUI2_0),.din(w_dff_A_5xGXelTX6_0),.clk(gclk));
	jdff dff_A_bghyKuUI2_0(.dout(w_dff_A_E2i1ybhL0_0),.din(w_dff_A_bghyKuUI2_0),.clk(gclk));
	jdff dff_A_E2i1ybhL0_0(.dout(w_dff_A_EK1Gfz8W8_0),.din(w_dff_A_E2i1ybhL0_0),.clk(gclk));
	jdff dff_A_EK1Gfz8W8_0(.dout(w_dff_A_uLktFuWB3_0),.din(w_dff_A_EK1Gfz8W8_0),.clk(gclk));
	jdff dff_A_uLktFuWB3_0(.dout(w_dff_A_MAndBeXK5_0),.din(w_dff_A_uLktFuWB3_0),.clk(gclk));
	jdff dff_A_MAndBeXK5_0(.dout(w_dff_A_yYgzJu3u3_0),.din(w_dff_A_MAndBeXK5_0),.clk(gclk));
	jdff dff_A_yYgzJu3u3_0(.dout(w_dff_A_wqBpYfAS3_0),.din(w_dff_A_yYgzJu3u3_0),.clk(gclk));
	jdff dff_A_wqBpYfAS3_0(.dout(w_dff_A_Yj1onD7G7_0),.din(w_dff_A_wqBpYfAS3_0),.clk(gclk));
	jdff dff_A_Yj1onD7G7_0(.dout(w_dff_A_jkjdi0Vl0_0),.din(w_dff_A_Yj1onD7G7_0),.clk(gclk));
	jdff dff_A_jkjdi0Vl0_0(.dout(w_dff_A_KIVEmHgf9_0),.din(w_dff_A_jkjdi0Vl0_0),.clk(gclk));
	jdff dff_A_KIVEmHgf9_0(.dout(w_dff_A_386dJLEL3_0),.din(w_dff_A_KIVEmHgf9_0),.clk(gclk));
	jdff dff_A_386dJLEL3_0(.dout(w_dff_A_sHLcL5qa6_0),.din(w_dff_A_386dJLEL3_0),.clk(gclk));
	jdff dff_A_sHLcL5qa6_0(.dout(w_dff_A_24Glr9AA7_0),.din(w_dff_A_sHLcL5qa6_0),.clk(gclk));
	jdff dff_A_24Glr9AA7_0(.dout(w_dff_A_v1VNd8VQ7_0),.din(w_dff_A_24Glr9AA7_0),.clk(gclk));
	jdff dff_A_v1VNd8VQ7_0(.dout(w_dff_A_nvOXj3F57_0),.din(w_dff_A_v1VNd8VQ7_0),.clk(gclk));
	jdff dff_A_nvOXj3F57_0(.dout(w_dff_A_NTJ7VvsC7_0),.din(w_dff_A_nvOXj3F57_0),.clk(gclk));
	jdff dff_A_NTJ7VvsC7_0(.dout(w_dff_A_CQN2ArvX2_0),.din(w_dff_A_NTJ7VvsC7_0),.clk(gclk));
	jdff dff_A_CQN2ArvX2_0(.dout(w_dff_A_U0yJrItQ5_0),.din(w_dff_A_CQN2ArvX2_0),.clk(gclk));
	jdff dff_A_U0yJrItQ5_0(.dout(w_dff_A_rBEuEehq5_0),.din(w_dff_A_U0yJrItQ5_0),.clk(gclk));
	jdff dff_A_rBEuEehq5_0(.dout(w_dff_A_fn0Ukzzx7_0),.din(w_dff_A_rBEuEehq5_0),.clk(gclk));
	jdff dff_A_fn0Ukzzx7_0(.dout(w_dff_A_NUOEiGJw3_0),.din(w_dff_A_fn0Ukzzx7_0),.clk(gclk));
	jdff dff_A_NUOEiGJw3_0(.dout(w_dff_A_vNswGoVS3_0),.din(w_dff_A_NUOEiGJw3_0),.clk(gclk));
	jdff dff_A_vNswGoVS3_0(.dout(w_dff_A_Cg96wRru5_0),.din(w_dff_A_vNswGoVS3_0),.clk(gclk));
	jdff dff_A_Cg96wRru5_0(.dout(w_dff_A_36QFqgDz7_0),.din(w_dff_A_Cg96wRru5_0),.clk(gclk));
	jdff dff_A_36QFqgDz7_0(.dout(w_dff_A_RGa31G8G5_0),.din(w_dff_A_36QFqgDz7_0),.clk(gclk));
	jdff dff_A_RGa31G8G5_0(.dout(w_dff_A_YCPseZMm8_0),.din(w_dff_A_RGa31G8G5_0),.clk(gclk));
	jdff dff_A_YCPseZMm8_0(.dout(w_dff_A_UvlBsSF25_0),.din(w_dff_A_YCPseZMm8_0),.clk(gclk));
	jdff dff_A_UvlBsSF25_0(.dout(w_dff_A_kpiZTyzw1_0),.din(w_dff_A_UvlBsSF25_0),.clk(gclk));
	jdff dff_A_kpiZTyzw1_0(.dout(w_dff_A_ayqQ7A1i2_0),.din(w_dff_A_kpiZTyzw1_0),.clk(gclk));
	jdff dff_A_ayqQ7A1i2_0(.dout(w_dff_A_NjUHC57B1_0),.din(w_dff_A_ayqQ7A1i2_0),.clk(gclk));
	jdff dff_A_NjUHC57B1_0(.dout(w_dff_A_r2mKJ7wF9_0),.din(w_dff_A_NjUHC57B1_0),.clk(gclk));
	jdff dff_A_r2mKJ7wF9_0(.dout(w_dff_A_57AD0IWV2_0),.din(w_dff_A_r2mKJ7wF9_0),.clk(gclk));
	jdff dff_A_57AD0IWV2_0(.dout(w_dff_A_6P8UH6uW9_0),.din(w_dff_A_57AD0IWV2_0),.clk(gclk));
	jdff dff_A_6P8UH6uW9_0(.dout(w_dff_A_60bRszFd5_0),.din(w_dff_A_6P8UH6uW9_0),.clk(gclk));
	jdff dff_A_60bRszFd5_0(.dout(w_dff_A_8sKKRmnR2_0),.din(w_dff_A_60bRszFd5_0),.clk(gclk));
	jdff dff_A_8sKKRmnR2_0(.dout(w_dff_A_xV2v85oK2_0),.din(w_dff_A_8sKKRmnR2_0),.clk(gclk));
	jdff dff_A_xV2v85oK2_0(.dout(w_dff_A_DvCj09hQ3_0),.din(w_dff_A_xV2v85oK2_0),.clk(gclk));
	jdff dff_A_DvCj09hQ3_0(.dout(w_dff_A_I1weYQuB4_0),.din(w_dff_A_DvCj09hQ3_0),.clk(gclk));
	jdff dff_A_I1weYQuB4_0(.dout(w_dff_A_q27U2D9o8_0),.din(w_dff_A_I1weYQuB4_0),.clk(gclk));
	jdff dff_A_q27U2D9o8_0(.dout(w_dff_A_yPvM6QNu6_0),.din(w_dff_A_q27U2D9o8_0),.clk(gclk));
	jdff dff_A_yPvM6QNu6_0(.dout(w_dff_A_lvQAJwyq8_0),.din(w_dff_A_yPvM6QNu6_0),.clk(gclk));
	jdff dff_A_lvQAJwyq8_0(.dout(w_dff_A_uIAXNmT81_0),.din(w_dff_A_lvQAJwyq8_0),.clk(gclk));
	jdff dff_A_uIAXNmT81_0(.dout(w_dff_A_oHDaYBC27_0),.din(w_dff_A_uIAXNmT81_0),.clk(gclk));
	jdff dff_A_oHDaYBC27_0(.dout(w_dff_A_4WTwgyoU7_0),.din(w_dff_A_oHDaYBC27_0),.clk(gclk));
	jdff dff_A_4WTwgyoU7_0(.dout(w_dff_A_dz8QVQCV4_0),.din(w_dff_A_4WTwgyoU7_0),.clk(gclk));
	jdff dff_A_dz8QVQCV4_0(.dout(w_dff_A_Id0BBLu50_0),.din(w_dff_A_dz8QVQCV4_0),.clk(gclk));
	jdff dff_A_Id0BBLu50_0(.dout(w_dff_A_Yi8Wyf0m3_0),.din(w_dff_A_Id0BBLu50_0),.clk(gclk));
	jdff dff_A_Yi8Wyf0m3_0(.dout(w_dff_A_ZDKNtDlh6_0),.din(w_dff_A_Yi8Wyf0m3_0),.clk(gclk));
	jdff dff_A_ZDKNtDlh6_0(.dout(w_dff_A_F2IbXNIW0_0),.din(w_dff_A_ZDKNtDlh6_0),.clk(gclk));
	jdff dff_A_F2IbXNIW0_0(.dout(w_dff_A_u8FpD4uR5_0),.din(w_dff_A_F2IbXNIW0_0),.clk(gclk));
	jdff dff_A_u8FpD4uR5_0(.dout(w_dff_A_9oP0trCv0_0),.din(w_dff_A_u8FpD4uR5_0),.clk(gclk));
	jdff dff_A_9oP0trCv0_0(.dout(f5),.din(w_dff_A_9oP0trCv0_0),.clk(gclk));
	jdff dff_A_IFRtoXuS7_2(.dout(w_dff_A_dNM5ioeY8_0),.din(w_dff_A_IFRtoXuS7_2),.clk(gclk));
	jdff dff_A_dNM5ioeY8_0(.dout(w_dff_A_0ygzNt811_0),.din(w_dff_A_dNM5ioeY8_0),.clk(gclk));
	jdff dff_A_0ygzNt811_0(.dout(w_dff_A_EedsJ0zS4_0),.din(w_dff_A_0ygzNt811_0),.clk(gclk));
	jdff dff_A_EedsJ0zS4_0(.dout(w_dff_A_nR94jSnj8_0),.din(w_dff_A_EedsJ0zS4_0),.clk(gclk));
	jdff dff_A_nR94jSnj8_0(.dout(w_dff_A_eXjQiPQt7_0),.din(w_dff_A_nR94jSnj8_0),.clk(gclk));
	jdff dff_A_eXjQiPQt7_0(.dout(w_dff_A_OfoPCtRU5_0),.din(w_dff_A_eXjQiPQt7_0),.clk(gclk));
	jdff dff_A_OfoPCtRU5_0(.dout(w_dff_A_1HGnTNNH6_0),.din(w_dff_A_OfoPCtRU5_0),.clk(gclk));
	jdff dff_A_1HGnTNNH6_0(.dout(w_dff_A_H0D9fyRI8_0),.din(w_dff_A_1HGnTNNH6_0),.clk(gclk));
	jdff dff_A_H0D9fyRI8_0(.dout(w_dff_A_O8ywRI6V9_0),.din(w_dff_A_H0D9fyRI8_0),.clk(gclk));
	jdff dff_A_O8ywRI6V9_0(.dout(w_dff_A_2puUNEVy8_0),.din(w_dff_A_O8ywRI6V9_0),.clk(gclk));
	jdff dff_A_2puUNEVy8_0(.dout(w_dff_A_e63m2zQL1_0),.din(w_dff_A_2puUNEVy8_0),.clk(gclk));
	jdff dff_A_e63m2zQL1_0(.dout(w_dff_A_x7oyIXNW4_0),.din(w_dff_A_e63m2zQL1_0),.clk(gclk));
	jdff dff_A_x7oyIXNW4_0(.dout(w_dff_A_8k4OgaXM9_0),.din(w_dff_A_x7oyIXNW4_0),.clk(gclk));
	jdff dff_A_8k4OgaXM9_0(.dout(w_dff_A_GQZndfBN9_0),.din(w_dff_A_8k4OgaXM9_0),.clk(gclk));
	jdff dff_A_GQZndfBN9_0(.dout(w_dff_A_78akKty68_0),.din(w_dff_A_GQZndfBN9_0),.clk(gclk));
	jdff dff_A_78akKty68_0(.dout(w_dff_A_jDohhRzZ7_0),.din(w_dff_A_78akKty68_0),.clk(gclk));
	jdff dff_A_jDohhRzZ7_0(.dout(w_dff_A_sigLi1SZ7_0),.din(w_dff_A_jDohhRzZ7_0),.clk(gclk));
	jdff dff_A_sigLi1SZ7_0(.dout(w_dff_A_KyI08DTP9_0),.din(w_dff_A_sigLi1SZ7_0),.clk(gclk));
	jdff dff_A_KyI08DTP9_0(.dout(w_dff_A_ay1uCFuY0_0),.din(w_dff_A_KyI08DTP9_0),.clk(gclk));
	jdff dff_A_ay1uCFuY0_0(.dout(w_dff_A_PTBc4VHW4_0),.din(w_dff_A_ay1uCFuY0_0),.clk(gclk));
	jdff dff_A_PTBc4VHW4_0(.dout(w_dff_A_UhzCJEAI6_0),.din(w_dff_A_PTBc4VHW4_0),.clk(gclk));
	jdff dff_A_UhzCJEAI6_0(.dout(w_dff_A_wZntfqmn0_0),.din(w_dff_A_UhzCJEAI6_0),.clk(gclk));
	jdff dff_A_wZntfqmn0_0(.dout(w_dff_A_QiAw9Cso6_0),.din(w_dff_A_wZntfqmn0_0),.clk(gclk));
	jdff dff_A_QiAw9Cso6_0(.dout(w_dff_A_I2m3H2mn7_0),.din(w_dff_A_QiAw9Cso6_0),.clk(gclk));
	jdff dff_A_I2m3H2mn7_0(.dout(w_dff_A_qb9nrwjr8_0),.din(w_dff_A_I2m3H2mn7_0),.clk(gclk));
	jdff dff_A_qb9nrwjr8_0(.dout(w_dff_A_vxNMFwka9_0),.din(w_dff_A_qb9nrwjr8_0),.clk(gclk));
	jdff dff_A_vxNMFwka9_0(.dout(w_dff_A_lv50pEPm8_0),.din(w_dff_A_vxNMFwka9_0),.clk(gclk));
	jdff dff_A_lv50pEPm8_0(.dout(w_dff_A_QNnuq1g22_0),.din(w_dff_A_lv50pEPm8_0),.clk(gclk));
	jdff dff_A_QNnuq1g22_0(.dout(w_dff_A_Qdj1UiX54_0),.din(w_dff_A_QNnuq1g22_0),.clk(gclk));
	jdff dff_A_Qdj1UiX54_0(.dout(w_dff_A_iUDjuwIf4_0),.din(w_dff_A_Qdj1UiX54_0),.clk(gclk));
	jdff dff_A_iUDjuwIf4_0(.dout(w_dff_A_sRzHDofR2_0),.din(w_dff_A_iUDjuwIf4_0),.clk(gclk));
	jdff dff_A_sRzHDofR2_0(.dout(w_dff_A_lXIBZskz4_0),.din(w_dff_A_sRzHDofR2_0),.clk(gclk));
	jdff dff_A_lXIBZskz4_0(.dout(w_dff_A_ieKkynYu2_0),.din(w_dff_A_lXIBZskz4_0),.clk(gclk));
	jdff dff_A_ieKkynYu2_0(.dout(w_dff_A_GqLd6dGd4_0),.din(w_dff_A_ieKkynYu2_0),.clk(gclk));
	jdff dff_A_GqLd6dGd4_0(.dout(w_dff_A_yNASuVxS7_0),.din(w_dff_A_GqLd6dGd4_0),.clk(gclk));
	jdff dff_A_yNASuVxS7_0(.dout(w_dff_A_mpq0EkWt2_0),.din(w_dff_A_yNASuVxS7_0),.clk(gclk));
	jdff dff_A_mpq0EkWt2_0(.dout(w_dff_A_PzDfoN9w7_0),.din(w_dff_A_mpq0EkWt2_0),.clk(gclk));
	jdff dff_A_PzDfoN9w7_0(.dout(w_dff_A_79FKcPhC3_0),.din(w_dff_A_PzDfoN9w7_0),.clk(gclk));
	jdff dff_A_79FKcPhC3_0(.dout(w_dff_A_aAE1O8N46_0),.din(w_dff_A_79FKcPhC3_0),.clk(gclk));
	jdff dff_A_aAE1O8N46_0(.dout(w_dff_A_mL4QLLKf1_0),.din(w_dff_A_aAE1O8N46_0),.clk(gclk));
	jdff dff_A_mL4QLLKf1_0(.dout(w_dff_A_8nu04Mvj3_0),.din(w_dff_A_mL4QLLKf1_0),.clk(gclk));
	jdff dff_A_8nu04Mvj3_0(.dout(w_dff_A_dKUoN67J0_0),.din(w_dff_A_8nu04Mvj3_0),.clk(gclk));
	jdff dff_A_dKUoN67J0_0(.dout(w_dff_A_PWoB4sES5_0),.din(w_dff_A_dKUoN67J0_0),.clk(gclk));
	jdff dff_A_PWoB4sES5_0(.dout(w_dff_A_SSWeRzZ21_0),.din(w_dff_A_PWoB4sES5_0),.clk(gclk));
	jdff dff_A_SSWeRzZ21_0(.dout(w_dff_A_jUfcUwEM8_0),.din(w_dff_A_SSWeRzZ21_0),.clk(gclk));
	jdff dff_A_jUfcUwEM8_0(.dout(w_dff_A_dIno3LGr7_0),.din(w_dff_A_jUfcUwEM8_0),.clk(gclk));
	jdff dff_A_dIno3LGr7_0(.dout(w_dff_A_lLTkimK53_0),.din(w_dff_A_dIno3LGr7_0),.clk(gclk));
	jdff dff_A_lLTkimK53_0(.dout(w_dff_A_nDAF2WLG0_0),.din(w_dff_A_lLTkimK53_0),.clk(gclk));
	jdff dff_A_nDAF2WLG0_0(.dout(w_dff_A_H1RYwhUX7_0),.din(w_dff_A_nDAF2WLG0_0),.clk(gclk));
	jdff dff_A_H1RYwhUX7_0(.dout(w_dff_A_zREFLy8k6_0),.din(w_dff_A_H1RYwhUX7_0),.clk(gclk));
	jdff dff_A_zREFLy8k6_0(.dout(w_dff_A_KFr37E3a6_0),.din(w_dff_A_zREFLy8k6_0),.clk(gclk));
	jdff dff_A_KFr37E3a6_0(.dout(w_dff_A_UUGkqhtd8_0),.din(w_dff_A_KFr37E3a6_0),.clk(gclk));
	jdff dff_A_UUGkqhtd8_0(.dout(w_dff_A_bKg73B4J5_0),.din(w_dff_A_UUGkqhtd8_0),.clk(gclk));
	jdff dff_A_bKg73B4J5_0(.dout(w_dff_A_cT9CC3GP3_0),.din(w_dff_A_bKg73B4J5_0),.clk(gclk));
	jdff dff_A_cT9CC3GP3_0(.dout(w_dff_A_w2BcjzP62_0),.din(w_dff_A_cT9CC3GP3_0),.clk(gclk));
	jdff dff_A_w2BcjzP62_0(.dout(w_dff_A_uSPJcw9i8_0),.din(w_dff_A_w2BcjzP62_0),.clk(gclk));
	jdff dff_A_uSPJcw9i8_0(.dout(w_dff_A_UmoshPVG6_0),.din(w_dff_A_uSPJcw9i8_0),.clk(gclk));
	jdff dff_A_UmoshPVG6_0(.dout(w_dff_A_SjfTFShX6_0),.din(w_dff_A_UmoshPVG6_0),.clk(gclk));
	jdff dff_A_SjfTFShX6_0(.dout(w_dff_A_PtLRR8HG1_0),.din(w_dff_A_SjfTFShX6_0),.clk(gclk));
	jdff dff_A_PtLRR8HG1_0(.dout(w_dff_A_sJrkBDuJ7_0),.din(w_dff_A_PtLRR8HG1_0),.clk(gclk));
	jdff dff_A_sJrkBDuJ7_0(.dout(w_dff_A_6ggOcCn26_0),.din(w_dff_A_sJrkBDuJ7_0),.clk(gclk));
	jdff dff_A_6ggOcCn26_0(.dout(w_dff_A_AENC41aY6_0),.din(w_dff_A_6ggOcCn26_0),.clk(gclk));
	jdff dff_A_AENC41aY6_0(.dout(w_dff_A_4UL4ueNJ7_0),.din(w_dff_A_AENC41aY6_0),.clk(gclk));
	jdff dff_A_4UL4ueNJ7_0(.dout(w_dff_A_dk8ZWBl44_0),.din(w_dff_A_4UL4ueNJ7_0),.clk(gclk));
	jdff dff_A_dk8ZWBl44_0(.dout(w_dff_A_7wjnj2BV3_0),.din(w_dff_A_dk8ZWBl44_0),.clk(gclk));
	jdff dff_A_7wjnj2BV3_0(.dout(w_dff_A_phvBqXQN8_0),.din(w_dff_A_7wjnj2BV3_0),.clk(gclk));
	jdff dff_A_phvBqXQN8_0(.dout(w_dff_A_xgz9OHjq8_0),.din(w_dff_A_phvBqXQN8_0),.clk(gclk));
	jdff dff_A_xgz9OHjq8_0(.dout(w_dff_A_3npU9qCm6_0),.din(w_dff_A_xgz9OHjq8_0),.clk(gclk));
	jdff dff_A_3npU9qCm6_0(.dout(w_dff_A_8MquYxoq7_0),.din(w_dff_A_3npU9qCm6_0),.clk(gclk));
	jdff dff_A_8MquYxoq7_0(.dout(w_dff_A_pRYTgd5Y3_0),.din(w_dff_A_8MquYxoq7_0),.clk(gclk));
	jdff dff_A_pRYTgd5Y3_0(.dout(w_dff_A_QSxdLCdb2_0),.din(w_dff_A_pRYTgd5Y3_0),.clk(gclk));
	jdff dff_A_QSxdLCdb2_0(.dout(w_dff_A_0JuxbPDB7_0),.din(w_dff_A_QSxdLCdb2_0),.clk(gclk));
	jdff dff_A_0JuxbPDB7_0(.dout(w_dff_A_lZSBKMYh7_0),.din(w_dff_A_0JuxbPDB7_0),.clk(gclk));
	jdff dff_A_lZSBKMYh7_0(.dout(w_dff_A_UvC2xjUo2_0),.din(w_dff_A_lZSBKMYh7_0),.clk(gclk));
	jdff dff_A_UvC2xjUo2_0(.dout(w_dff_A_xceiiTia7_0),.din(w_dff_A_UvC2xjUo2_0),.clk(gclk));
	jdff dff_A_xceiiTia7_0(.dout(w_dff_A_cto6lBMf8_0),.din(w_dff_A_xceiiTia7_0),.clk(gclk));
	jdff dff_A_cto6lBMf8_0(.dout(w_dff_A_hzLgh0216_0),.din(w_dff_A_cto6lBMf8_0),.clk(gclk));
	jdff dff_A_hzLgh0216_0(.dout(w_dff_A_pQLE9Es92_0),.din(w_dff_A_hzLgh0216_0),.clk(gclk));
	jdff dff_A_pQLE9Es92_0(.dout(w_dff_A_8xlRWhvp6_0),.din(w_dff_A_pQLE9Es92_0),.clk(gclk));
	jdff dff_A_8xlRWhvp6_0(.dout(w_dff_A_3V3HZntB9_0),.din(w_dff_A_8xlRWhvp6_0),.clk(gclk));
	jdff dff_A_3V3HZntB9_0(.dout(w_dff_A_F5KFFyef7_0),.din(w_dff_A_3V3HZntB9_0),.clk(gclk));
	jdff dff_A_F5KFFyef7_0(.dout(w_dff_A_go6OBVaW8_0),.din(w_dff_A_F5KFFyef7_0),.clk(gclk));
	jdff dff_A_go6OBVaW8_0(.dout(w_dff_A_RX5tRT9m0_0),.din(w_dff_A_go6OBVaW8_0),.clk(gclk));
	jdff dff_A_RX5tRT9m0_0(.dout(w_dff_A_Be4yMm239_0),.din(w_dff_A_RX5tRT9m0_0),.clk(gclk));
	jdff dff_A_Be4yMm239_0(.dout(w_dff_A_uOdvJjvm4_0),.din(w_dff_A_Be4yMm239_0),.clk(gclk));
	jdff dff_A_uOdvJjvm4_0(.dout(w_dff_A_42nriZNs1_0),.din(w_dff_A_uOdvJjvm4_0),.clk(gclk));
	jdff dff_A_42nriZNs1_0(.dout(w_dff_A_ppgYe0Kr6_0),.din(w_dff_A_42nriZNs1_0),.clk(gclk));
	jdff dff_A_ppgYe0Kr6_0(.dout(w_dff_A_otdmyLKD7_0),.din(w_dff_A_ppgYe0Kr6_0),.clk(gclk));
	jdff dff_A_otdmyLKD7_0(.dout(w_dff_A_rWF4A0gh4_0),.din(w_dff_A_otdmyLKD7_0),.clk(gclk));
	jdff dff_A_rWF4A0gh4_0(.dout(w_dff_A_UwWgvn8a0_0),.din(w_dff_A_rWF4A0gh4_0),.clk(gclk));
	jdff dff_A_UwWgvn8a0_0(.dout(w_dff_A_w2czANKh2_0),.din(w_dff_A_UwWgvn8a0_0),.clk(gclk));
	jdff dff_A_w2czANKh2_0(.dout(w_dff_A_CJ26oO9q6_0),.din(w_dff_A_w2czANKh2_0),.clk(gclk));
	jdff dff_A_CJ26oO9q6_0(.dout(w_dff_A_jpbqLsyl6_0),.din(w_dff_A_CJ26oO9q6_0),.clk(gclk));
	jdff dff_A_jpbqLsyl6_0(.dout(w_dff_A_bHTNkRPH6_0),.din(w_dff_A_jpbqLsyl6_0),.clk(gclk));
	jdff dff_A_bHTNkRPH6_0(.dout(w_dff_A_tnzXvyKY8_0),.din(w_dff_A_bHTNkRPH6_0),.clk(gclk));
	jdff dff_A_tnzXvyKY8_0(.dout(w_dff_A_TSwnZtYR1_0),.din(w_dff_A_tnzXvyKY8_0),.clk(gclk));
	jdff dff_A_TSwnZtYR1_0(.dout(w_dff_A_q8ytKrrd2_0),.din(w_dff_A_TSwnZtYR1_0),.clk(gclk));
	jdff dff_A_q8ytKrrd2_0(.dout(w_dff_A_Ue1GZ5cq5_0),.din(w_dff_A_q8ytKrrd2_0),.clk(gclk));
	jdff dff_A_Ue1GZ5cq5_0(.dout(w_dff_A_Ywq21yhK5_0),.din(w_dff_A_Ue1GZ5cq5_0),.clk(gclk));
	jdff dff_A_Ywq21yhK5_0(.dout(w_dff_A_xG9KR7KU8_0),.din(w_dff_A_Ywq21yhK5_0),.clk(gclk));
	jdff dff_A_xG9KR7KU8_0(.dout(w_dff_A_lVxRtu1v4_0),.din(w_dff_A_xG9KR7KU8_0),.clk(gclk));
	jdff dff_A_lVxRtu1v4_0(.dout(w_dff_A_TZjE7A617_0),.din(w_dff_A_lVxRtu1v4_0),.clk(gclk));
	jdff dff_A_TZjE7A617_0(.dout(w_dff_A_hPOK1ZsB9_0),.din(w_dff_A_TZjE7A617_0),.clk(gclk));
	jdff dff_A_hPOK1ZsB9_0(.dout(w_dff_A_4j3yS4H37_0),.din(w_dff_A_hPOK1ZsB9_0),.clk(gclk));
	jdff dff_A_4j3yS4H37_0(.dout(w_dff_A_TluW0DJW4_0),.din(w_dff_A_4j3yS4H37_0),.clk(gclk));
	jdff dff_A_TluW0DJW4_0(.dout(w_dff_A_GnHab2jC0_0),.din(w_dff_A_TluW0DJW4_0),.clk(gclk));
	jdff dff_A_GnHab2jC0_0(.dout(w_dff_A_RfhKmTB59_0),.din(w_dff_A_GnHab2jC0_0),.clk(gclk));
	jdff dff_A_RfhKmTB59_0(.dout(w_dff_A_UJYzzDkr1_0),.din(w_dff_A_RfhKmTB59_0),.clk(gclk));
	jdff dff_A_UJYzzDkr1_0(.dout(w_dff_A_925rrjgO8_0),.din(w_dff_A_UJYzzDkr1_0),.clk(gclk));
	jdff dff_A_925rrjgO8_0(.dout(w_dff_A_a1tI1IAw9_0),.din(w_dff_A_925rrjgO8_0),.clk(gclk));
	jdff dff_A_a1tI1IAw9_0(.dout(w_dff_A_EWxKoSIP0_0),.din(w_dff_A_a1tI1IAw9_0),.clk(gclk));
	jdff dff_A_EWxKoSIP0_0(.dout(w_dff_A_t1uDvSzH4_0),.din(w_dff_A_EWxKoSIP0_0),.clk(gclk));
	jdff dff_A_t1uDvSzH4_0(.dout(w_dff_A_yyWyHS926_0),.din(w_dff_A_t1uDvSzH4_0),.clk(gclk));
	jdff dff_A_yyWyHS926_0(.dout(w_dff_A_Wdkx0ujD7_0),.din(w_dff_A_yyWyHS926_0),.clk(gclk));
	jdff dff_A_Wdkx0ujD7_0(.dout(w_dff_A_TYoTy2uZ8_0),.din(w_dff_A_Wdkx0ujD7_0),.clk(gclk));
	jdff dff_A_TYoTy2uZ8_0(.dout(w_dff_A_ZmqUekGv8_0),.din(w_dff_A_TYoTy2uZ8_0),.clk(gclk));
	jdff dff_A_ZmqUekGv8_0(.dout(w_dff_A_PCLwuSUy5_0),.din(w_dff_A_ZmqUekGv8_0),.clk(gclk));
	jdff dff_A_PCLwuSUy5_0(.dout(w_dff_A_iGyCGKtU5_0),.din(w_dff_A_PCLwuSUy5_0),.clk(gclk));
	jdff dff_A_iGyCGKtU5_0(.dout(w_dff_A_hnlozL1W4_0),.din(w_dff_A_iGyCGKtU5_0),.clk(gclk));
	jdff dff_A_hnlozL1W4_0(.dout(w_dff_A_yaVjxPvn7_0),.din(w_dff_A_hnlozL1W4_0),.clk(gclk));
	jdff dff_A_yaVjxPvn7_0(.dout(f6),.din(w_dff_A_yaVjxPvn7_0),.clk(gclk));
	jdff dff_A_sGoHlvcX8_2(.dout(w_dff_A_4W6QZxc78_0),.din(w_dff_A_sGoHlvcX8_2),.clk(gclk));
	jdff dff_A_4W6QZxc78_0(.dout(w_dff_A_egHFEAyw0_0),.din(w_dff_A_4W6QZxc78_0),.clk(gclk));
	jdff dff_A_egHFEAyw0_0(.dout(w_dff_A_xQncDKc42_0),.din(w_dff_A_egHFEAyw0_0),.clk(gclk));
	jdff dff_A_xQncDKc42_0(.dout(w_dff_A_g4eQNZOc3_0),.din(w_dff_A_xQncDKc42_0),.clk(gclk));
	jdff dff_A_g4eQNZOc3_0(.dout(w_dff_A_hOLSdc635_0),.din(w_dff_A_g4eQNZOc3_0),.clk(gclk));
	jdff dff_A_hOLSdc635_0(.dout(w_dff_A_fqYRsZHI8_0),.din(w_dff_A_hOLSdc635_0),.clk(gclk));
	jdff dff_A_fqYRsZHI8_0(.dout(w_dff_A_Jb19i3wQ9_0),.din(w_dff_A_fqYRsZHI8_0),.clk(gclk));
	jdff dff_A_Jb19i3wQ9_0(.dout(w_dff_A_kYfU3JQz5_0),.din(w_dff_A_Jb19i3wQ9_0),.clk(gclk));
	jdff dff_A_kYfU3JQz5_0(.dout(w_dff_A_8gRy1Co38_0),.din(w_dff_A_kYfU3JQz5_0),.clk(gclk));
	jdff dff_A_8gRy1Co38_0(.dout(w_dff_A_lVyFbCZS6_0),.din(w_dff_A_8gRy1Co38_0),.clk(gclk));
	jdff dff_A_lVyFbCZS6_0(.dout(w_dff_A_KQxBJq8i3_0),.din(w_dff_A_lVyFbCZS6_0),.clk(gclk));
	jdff dff_A_KQxBJq8i3_0(.dout(w_dff_A_dj9Kq0th5_0),.din(w_dff_A_KQxBJq8i3_0),.clk(gclk));
	jdff dff_A_dj9Kq0th5_0(.dout(w_dff_A_kCgK3GXG1_0),.din(w_dff_A_dj9Kq0th5_0),.clk(gclk));
	jdff dff_A_kCgK3GXG1_0(.dout(w_dff_A_U1RU7iWf1_0),.din(w_dff_A_kCgK3GXG1_0),.clk(gclk));
	jdff dff_A_U1RU7iWf1_0(.dout(w_dff_A_Q8udJ7bo7_0),.din(w_dff_A_U1RU7iWf1_0),.clk(gclk));
	jdff dff_A_Q8udJ7bo7_0(.dout(w_dff_A_nkJA41tR4_0),.din(w_dff_A_Q8udJ7bo7_0),.clk(gclk));
	jdff dff_A_nkJA41tR4_0(.dout(w_dff_A_8HcvDrca6_0),.din(w_dff_A_nkJA41tR4_0),.clk(gclk));
	jdff dff_A_8HcvDrca6_0(.dout(w_dff_A_ydAZef970_0),.din(w_dff_A_8HcvDrca6_0),.clk(gclk));
	jdff dff_A_ydAZef970_0(.dout(w_dff_A_P6LCG2DZ0_0),.din(w_dff_A_ydAZef970_0),.clk(gclk));
	jdff dff_A_P6LCG2DZ0_0(.dout(w_dff_A_nLTMRlbh1_0),.din(w_dff_A_P6LCG2DZ0_0),.clk(gclk));
	jdff dff_A_nLTMRlbh1_0(.dout(w_dff_A_n3ZpOXDP8_0),.din(w_dff_A_nLTMRlbh1_0),.clk(gclk));
	jdff dff_A_n3ZpOXDP8_0(.dout(w_dff_A_VdA4E3q73_0),.din(w_dff_A_n3ZpOXDP8_0),.clk(gclk));
	jdff dff_A_VdA4E3q73_0(.dout(w_dff_A_eBOsIbtN9_0),.din(w_dff_A_VdA4E3q73_0),.clk(gclk));
	jdff dff_A_eBOsIbtN9_0(.dout(w_dff_A_sRNozZAn6_0),.din(w_dff_A_eBOsIbtN9_0),.clk(gclk));
	jdff dff_A_sRNozZAn6_0(.dout(w_dff_A_SHwXN1RT1_0),.din(w_dff_A_sRNozZAn6_0),.clk(gclk));
	jdff dff_A_SHwXN1RT1_0(.dout(w_dff_A_cFyh7PrA6_0),.din(w_dff_A_SHwXN1RT1_0),.clk(gclk));
	jdff dff_A_cFyh7PrA6_0(.dout(w_dff_A_VskicEZp3_0),.din(w_dff_A_cFyh7PrA6_0),.clk(gclk));
	jdff dff_A_VskicEZp3_0(.dout(w_dff_A_IfunqZdA5_0),.din(w_dff_A_VskicEZp3_0),.clk(gclk));
	jdff dff_A_IfunqZdA5_0(.dout(w_dff_A_2RpfZK663_0),.din(w_dff_A_IfunqZdA5_0),.clk(gclk));
	jdff dff_A_2RpfZK663_0(.dout(w_dff_A_ZbZntsYK3_0),.din(w_dff_A_2RpfZK663_0),.clk(gclk));
	jdff dff_A_ZbZntsYK3_0(.dout(w_dff_A_v5ncrlI21_0),.din(w_dff_A_ZbZntsYK3_0),.clk(gclk));
	jdff dff_A_v5ncrlI21_0(.dout(w_dff_A_4eNYktAA3_0),.din(w_dff_A_v5ncrlI21_0),.clk(gclk));
	jdff dff_A_4eNYktAA3_0(.dout(w_dff_A_un74S38m7_0),.din(w_dff_A_4eNYktAA3_0),.clk(gclk));
	jdff dff_A_un74S38m7_0(.dout(w_dff_A_zM36sHxC7_0),.din(w_dff_A_un74S38m7_0),.clk(gclk));
	jdff dff_A_zM36sHxC7_0(.dout(w_dff_A_nCJAiT6V4_0),.din(w_dff_A_zM36sHxC7_0),.clk(gclk));
	jdff dff_A_nCJAiT6V4_0(.dout(w_dff_A_1mMAkSBq5_0),.din(w_dff_A_nCJAiT6V4_0),.clk(gclk));
	jdff dff_A_1mMAkSBq5_0(.dout(w_dff_A_qkvT121X8_0),.din(w_dff_A_1mMAkSBq5_0),.clk(gclk));
	jdff dff_A_qkvT121X8_0(.dout(w_dff_A_JMf8sMHM2_0),.din(w_dff_A_qkvT121X8_0),.clk(gclk));
	jdff dff_A_JMf8sMHM2_0(.dout(w_dff_A_93Ktuyfd4_0),.din(w_dff_A_JMf8sMHM2_0),.clk(gclk));
	jdff dff_A_93Ktuyfd4_0(.dout(w_dff_A_r1GFEXQe4_0),.din(w_dff_A_93Ktuyfd4_0),.clk(gclk));
	jdff dff_A_r1GFEXQe4_0(.dout(w_dff_A_6yJ42Ukp5_0),.din(w_dff_A_r1GFEXQe4_0),.clk(gclk));
	jdff dff_A_6yJ42Ukp5_0(.dout(w_dff_A_iNarG90M1_0),.din(w_dff_A_6yJ42Ukp5_0),.clk(gclk));
	jdff dff_A_iNarG90M1_0(.dout(w_dff_A_N3XvRgar4_0),.din(w_dff_A_iNarG90M1_0),.clk(gclk));
	jdff dff_A_N3XvRgar4_0(.dout(w_dff_A_XsHZS8VK4_0),.din(w_dff_A_N3XvRgar4_0),.clk(gclk));
	jdff dff_A_XsHZS8VK4_0(.dout(w_dff_A_0Cz0pDGs1_0),.din(w_dff_A_XsHZS8VK4_0),.clk(gclk));
	jdff dff_A_0Cz0pDGs1_0(.dout(w_dff_A_1Wr2h8cN8_0),.din(w_dff_A_0Cz0pDGs1_0),.clk(gclk));
	jdff dff_A_1Wr2h8cN8_0(.dout(w_dff_A_xRp3GTiY1_0),.din(w_dff_A_1Wr2h8cN8_0),.clk(gclk));
	jdff dff_A_xRp3GTiY1_0(.dout(w_dff_A_eHpDtK417_0),.din(w_dff_A_xRp3GTiY1_0),.clk(gclk));
	jdff dff_A_eHpDtK417_0(.dout(w_dff_A_ZVNAuxVq1_0),.din(w_dff_A_eHpDtK417_0),.clk(gclk));
	jdff dff_A_ZVNAuxVq1_0(.dout(w_dff_A_UO38ASv10_0),.din(w_dff_A_ZVNAuxVq1_0),.clk(gclk));
	jdff dff_A_UO38ASv10_0(.dout(w_dff_A_bB9O1liK7_0),.din(w_dff_A_UO38ASv10_0),.clk(gclk));
	jdff dff_A_bB9O1liK7_0(.dout(w_dff_A_lXbVM0Hc0_0),.din(w_dff_A_bB9O1liK7_0),.clk(gclk));
	jdff dff_A_lXbVM0Hc0_0(.dout(w_dff_A_AFab10RQ2_0),.din(w_dff_A_lXbVM0Hc0_0),.clk(gclk));
	jdff dff_A_AFab10RQ2_0(.dout(w_dff_A_ZwNktAb33_0),.din(w_dff_A_AFab10RQ2_0),.clk(gclk));
	jdff dff_A_ZwNktAb33_0(.dout(w_dff_A_sczRJfeQ8_0),.din(w_dff_A_ZwNktAb33_0),.clk(gclk));
	jdff dff_A_sczRJfeQ8_0(.dout(w_dff_A_ljBd9yWV3_0),.din(w_dff_A_sczRJfeQ8_0),.clk(gclk));
	jdff dff_A_ljBd9yWV3_0(.dout(w_dff_A_6EPYn6hh2_0),.din(w_dff_A_ljBd9yWV3_0),.clk(gclk));
	jdff dff_A_6EPYn6hh2_0(.dout(w_dff_A_sEQHXFxK6_0),.din(w_dff_A_6EPYn6hh2_0),.clk(gclk));
	jdff dff_A_sEQHXFxK6_0(.dout(w_dff_A_9BSO4exH9_0),.din(w_dff_A_sEQHXFxK6_0),.clk(gclk));
	jdff dff_A_9BSO4exH9_0(.dout(w_dff_A_g06sEK4S9_0),.din(w_dff_A_9BSO4exH9_0),.clk(gclk));
	jdff dff_A_g06sEK4S9_0(.dout(w_dff_A_YTQR9xzP1_0),.din(w_dff_A_g06sEK4S9_0),.clk(gclk));
	jdff dff_A_YTQR9xzP1_0(.dout(w_dff_A_zwNUoZ8I6_0),.din(w_dff_A_YTQR9xzP1_0),.clk(gclk));
	jdff dff_A_zwNUoZ8I6_0(.dout(w_dff_A_OwqRkI7r5_0),.din(w_dff_A_zwNUoZ8I6_0),.clk(gclk));
	jdff dff_A_OwqRkI7r5_0(.dout(w_dff_A_Xi4fSevg6_0),.din(w_dff_A_OwqRkI7r5_0),.clk(gclk));
	jdff dff_A_Xi4fSevg6_0(.dout(w_dff_A_SEvnLM3O7_0),.din(w_dff_A_Xi4fSevg6_0),.clk(gclk));
	jdff dff_A_SEvnLM3O7_0(.dout(w_dff_A_Af7rwO4Z3_0),.din(w_dff_A_SEvnLM3O7_0),.clk(gclk));
	jdff dff_A_Af7rwO4Z3_0(.dout(w_dff_A_cPeZ6SD53_0),.din(w_dff_A_Af7rwO4Z3_0),.clk(gclk));
	jdff dff_A_cPeZ6SD53_0(.dout(w_dff_A_5hx7B5lh3_0),.din(w_dff_A_cPeZ6SD53_0),.clk(gclk));
	jdff dff_A_5hx7B5lh3_0(.dout(w_dff_A_Q6Nl3oap9_0),.din(w_dff_A_5hx7B5lh3_0),.clk(gclk));
	jdff dff_A_Q6Nl3oap9_0(.dout(w_dff_A_zRuQDe172_0),.din(w_dff_A_Q6Nl3oap9_0),.clk(gclk));
	jdff dff_A_zRuQDe172_0(.dout(w_dff_A_grXBwiRm9_0),.din(w_dff_A_zRuQDe172_0),.clk(gclk));
	jdff dff_A_grXBwiRm9_0(.dout(w_dff_A_Sr2siA583_0),.din(w_dff_A_grXBwiRm9_0),.clk(gclk));
	jdff dff_A_Sr2siA583_0(.dout(w_dff_A_ESw6a8MQ7_0),.din(w_dff_A_Sr2siA583_0),.clk(gclk));
	jdff dff_A_ESw6a8MQ7_0(.dout(w_dff_A_4BjnqR7I0_0),.din(w_dff_A_ESw6a8MQ7_0),.clk(gclk));
	jdff dff_A_4BjnqR7I0_0(.dout(w_dff_A_cRTrEahq9_0),.din(w_dff_A_4BjnqR7I0_0),.clk(gclk));
	jdff dff_A_cRTrEahq9_0(.dout(w_dff_A_qmuqNwqD7_0),.din(w_dff_A_cRTrEahq9_0),.clk(gclk));
	jdff dff_A_qmuqNwqD7_0(.dout(w_dff_A_YLFiNG3B4_0),.din(w_dff_A_qmuqNwqD7_0),.clk(gclk));
	jdff dff_A_YLFiNG3B4_0(.dout(w_dff_A_J1xrbLhx1_0),.din(w_dff_A_YLFiNG3B4_0),.clk(gclk));
	jdff dff_A_J1xrbLhx1_0(.dout(w_dff_A_OGLOL5e16_0),.din(w_dff_A_J1xrbLhx1_0),.clk(gclk));
	jdff dff_A_OGLOL5e16_0(.dout(w_dff_A_NZ6qgRVI9_0),.din(w_dff_A_OGLOL5e16_0),.clk(gclk));
	jdff dff_A_NZ6qgRVI9_0(.dout(w_dff_A_yDktkIvR3_0),.din(w_dff_A_NZ6qgRVI9_0),.clk(gclk));
	jdff dff_A_yDktkIvR3_0(.dout(w_dff_A_6izQlhzq8_0),.din(w_dff_A_yDktkIvR3_0),.clk(gclk));
	jdff dff_A_6izQlhzq8_0(.dout(w_dff_A_7YKBEPnx5_0),.din(w_dff_A_6izQlhzq8_0),.clk(gclk));
	jdff dff_A_7YKBEPnx5_0(.dout(w_dff_A_IoSZqDpj8_0),.din(w_dff_A_7YKBEPnx5_0),.clk(gclk));
	jdff dff_A_IoSZqDpj8_0(.dout(w_dff_A_5EeVt9Zi0_0),.din(w_dff_A_IoSZqDpj8_0),.clk(gclk));
	jdff dff_A_5EeVt9Zi0_0(.dout(w_dff_A_XhSkDvQV1_0),.din(w_dff_A_5EeVt9Zi0_0),.clk(gclk));
	jdff dff_A_XhSkDvQV1_0(.dout(w_dff_A_TVkwsmJZ4_0),.din(w_dff_A_XhSkDvQV1_0),.clk(gclk));
	jdff dff_A_TVkwsmJZ4_0(.dout(w_dff_A_GNGWReUy8_0),.din(w_dff_A_TVkwsmJZ4_0),.clk(gclk));
	jdff dff_A_GNGWReUy8_0(.dout(w_dff_A_hsVe60Ms8_0),.din(w_dff_A_GNGWReUy8_0),.clk(gclk));
	jdff dff_A_hsVe60Ms8_0(.dout(w_dff_A_7KETfTpp2_0),.din(w_dff_A_hsVe60Ms8_0),.clk(gclk));
	jdff dff_A_7KETfTpp2_0(.dout(w_dff_A_QhwUvnqZ9_0),.din(w_dff_A_7KETfTpp2_0),.clk(gclk));
	jdff dff_A_QhwUvnqZ9_0(.dout(w_dff_A_FRo5TK4e1_0),.din(w_dff_A_QhwUvnqZ9_0),.clk(gclk));
	jdff dff_A_FRo5TK4e1_0(.dout(w_dff_A_t2taBbP39_0),.din(w_dff_A_FRo5TK4e1_0),.clk(gclk));
	jdff dff_A_t2taBbP39_0(.dout(w_dff_A_rheuBGEr4_0),.din(w_dff_A_t2taBbP39_0),.clk(gclk));
	jdff dff_A_rheuBGEr4_0(.dout(w_dff_A_rKnPW2378_0),.din(w_dff_A_rheuBGEr4_0),.clk(gclk));
	jdff dff_A_rKnPW2378_0(.dout(w_dff_A_DFP2rKdu3_0),.din(w_dff_A_rKnPW2378_0),.clk(gclk));
	jdff dff_A_DFP2rKdu3_0(.dout(w_dff_A_xuXzxhla2_0),.din(w_dff_A_DFP2rKdu3_0),.clk(gclk));
	jdff dff_A_xuXzxhla2_0(.dout(w_dff_A_sFJmA4jD6_0),.din(w_dff_A_xuXzxhla2_0),.clk(gclk));
	jdff dff_A_sFJmA4jD6_0(.dout(w_dff_A_oVxZavgL9_0),.din(w_dff_A_sFJmA4jD6_0),.clk(gclk));
	jdff dff_A_oVxZavgL9_0(.dout(w_dff_A_awQuYCXd9_0),.din(w_dff_A_oVxZavgL9_0),.clk(gclk));
	jdff dff_A_awQuYCXd9_0(.dout(w_dff_A_J4a8nY809_0),.din(w_dff_A_awQuYCXd9_0),.clk(gclk));
	jdff dff_A_J4a8nY809_0(.dout(w_dff_A_2FgvZGJk8_0),.din(w_dff_A_J4a8nY809_0),.clk(gclk));
	jdff dff_A_2FgvZGJk8_0(.dout(w_dff_A_KmD7Mh4p8_0),.din(w_dff_A_2FgvZGJk8_0),.clk(gclk));
	jdff dff_A_KmD7Mh4p8_0(.dout(w_dff_A_IjoCFhh39_0),.din(w_dff_A_KmD7Mh4p8_0),.clk(gclk));
	jdff dff_A_IjoCFhh39_0(.dout(w_dff_A_1RoD7IHH2_0),.din(w_dff_A_IjoCFhh39_0),.clk(gclk));
	jdff dff_A_1RoD7IHH2_0(.dout(w_dff_A_qfEw5MSI1_0),.din(w_dff_A_1RoD7IHH2_0),.clk(gclk));
	jdff dff_A_qfEw5MSI1_0(.dout(w_dff_A_bJGkmqbU5_0),.din(w_dff_A_qfEw5MSI1_0),.clk(gclk));
	jdff dff_A_bJGkmqbU5_0(.dout(w_dff_A_jXJoTtAM3_0),.din(w_dff_A_bJGkmqbU5_0),.clk(gclk));
	jdff dff_A_jXJoTtAM3_0(.dout(w_dff_A_Vg6NI2J61_0),.din(w_dff_A_jXJoTtAM3_0),.clk(gclk));
	jdff dff_A_Vg6NI2J61_0(.dout(w_dff_A_qDULmxVk6_0),.din(w_dff_A_Vg6NI2J61_0),.clk(gclk));
	jdff dff_A_qDULmxVk6_0(.dout(w_dff_A_LFMid0cB6_0),.din(w_dff_A_qDULmxVk6_0),.clk(gclk));
	jdff dff_A_LFMid0cB6_0(.dout(w_dff_A_2VakWFqR1_0),.din(w_dff_A_LFMid0cB6_0),.clk(gclk));
	jdff dff_A_2VakWFqR1_0(.dout(w_dff_A_7EZaGmYx2_0),.din(w_dff_A_2VakWFqR1_0),.clk(gclk));
	jdff dff_A_7EZaGmYx2_0(.dout(w_dff_A_R4ues0R64_0),.din(w_dff_A_7EZaGmYx2_0),.clk(gclk));
	jdff dff_A_R4ues0R64_0(.dout(w_dff_A_YG7bvOdM3_0),.din(w_dff_A_R4ues0R64_0),.clk(gclk));
	jdff dff_A_YG7bvOdM3_0(.dout(w_dff_A_MgyK0MRL9_0),.din(w_dff_A_YG7bvOdM3_0),.clk(gclk));
	jdff dff_A_MgyK0MRL9_0(.dout(w_dff_A_R7FH4fbX2_0),.din(w_dff_A_MgyK0MRL9_0),.clk(gclk));
	jdff dff_A_R7FH4fbX2_0(.dout(w_dff_A_58MSGd9a7_0),.din(w_dff_A_R7FH4fbX2_0),.clk(gclk));
	jdff dff_A_58MSGd9a7_0(.dout(w_dff_A_ZLwKLtJq3_0),.din(w_dff_A_58MSGd9a7_0),.clk(gclk));
	jdff dff_A_ZLwKLtJq3_0(.dout(f7),.din(w_dff_A_ZLwKLtJq3_0),.clk(gclk));
	jdff dff_A_hqBdsfmR3_2(.dout(w_dff_A_sWOG7FHo8_0),.din(w_dff_A_hqBdsfmR3_2),.clk(gclk));
	jdff dff_A_sWOG7FHo8_0(.dout(w_dff_A_k077Uut50_0),.din(w_dff_A_sWOG7FHo8_0),.clk(gclk));
	jdff dff_A_k077Uut50_0(.dout(w_dff_A_bADamjWn4_0),.din(w_dff_A_k077Uut50_0),.clk(gclk));
	jdff dff_A_bADamjWn4_0(.dout(w_dff_A_Q60y1mUk9_0),.din(w_dff_A_bADamjWn4_0),.clk(gclk));
	jdff dff_A_Q60y1mUk9_0(.dout(w_dff_A_1mVcQcAE2_0),.din(w_dff_A_Q60y1mUk9_0),.clk(gclk));
	jdff dff_A_1mVcQcAE2_0(.dout(w_dff_A_fe1zIwkf6_0),.din(w_dff_A_1mVcQcAE2_0),.clk(gclk));
	jdff dff_A_fe1zIwkf6_0(.dout(w_dff_A_0VUjgbwC6_0),.din(w_dff_A_fe1zIwkf6_0),.clk(gclk));
	jdff dff_A_0VUjgbwC6_0(.dout(w_dff_A_As6ONpT40_0),.din(w_dff_A_0VUjgbwC6_0),.clk(gclk));
	jdff dff_A_As6ONpT40_0(.dout(w_dff_A_xnxkpoyT4_0),.din(w_dff_A_As6ONpT40_0),.clk(gclk));
	jdff dff_A_xnxkpoyT4_0(.dout(w_dff_A_HMsgNolo4_0),.din(w_dff_A_xnxkpoyT4_0),.clk(gclk));
	jdff dff_A_HMsgNolo4_0(.dout(w_dff_A_gtfnUHQE7_0),.din(w_dff_A_HMsgNolo4_0),.clk(gclk));
	jdff dff_A_gtfnUHQE7_0(.dout(w_dff_A_A3i2bFjX6_0),.din(w_dff_A_gtfnUHQE7_0),.clk(gclk));
	jdff dff_A_A3i2bFjX6_0(.dout(w_dff_A_UbUe2Kf17_0),.din(w_dff_A_A3i2bFjX6_0),.clk(gclk));
	jdff dff_A_UbUe2Kf17_0(.dout(w_dff_A_U1S8mGzU5_0),.din(w_dff_A_UbUe2Kf17_0),.clk(gclk));
	jdff dff_A_U1S8mGzU5_0(.dout(w_dff_A_Z6zYKh7O3_0),.din(w_dff_A_U1S8mGzU5_0),.clk(gclk));
	jdff dff_A_Z6zYKh7O3_0(.dout(w_dff_A_ewdPHNFY3_0),.din(w_dff_A_Z6zYKh7O3_0),.clk(gclk));
	jdff dff_A_ewdPHNFY3_0(.dout(w_dff_A_yuhBwgqv6_0),.din(w_dff_A_ewdPHNFY3_0),.clk(gclk));
	jdff dff_A_yuhBwgqv6_0(.dout(w_dff_A_wl9MechG2_0),.din(w_dff_A_yuhBwgqv6_0),.clk(gclk));
	jdff dff_A_wl9MechG2_0(.dout(w_dff_A_yCspxLdO2_0),.din(w_dff_A_wl9MechG2_0),.clk(gclk));
	jdff dff_A_yCspxLdO2_0(.dout(w_dff_A_yaYyfitw1_0),.din(w_dff_A_yCspxLdO2_0),.clk(gclk));
	jdff dff_A_yaYyfitw1_0(.dout(w_dff_A_Xty69Cur9_0),.din(w_dff_A_yaYyfitw1_0),.clk(gclk));
	jdff dff_A_Xty69Cur9_0(.dout(w_dff_A_grMN48ne6_0),.din(w_dff_A_Xty69Cur9_0),.clk(gclk));
	jdff dff_A_grMN48ne6_0(.dout(w_dff_A_LROwg5h05_0),.din(w_dff_A_grMN48ne6_0),.clk(gclk));
	jdff dff_A_LROwg5h05_0(.dout(w_dff_A_Uhaay64q2_0),.din(w_dff_A_LROwg5h05_0),.clk(gclk));
	jdff dff_A_Uhaay64q2_0(.dout(w_dff_A_wmNJ4NLZ6_0),.din(w_dff_A_Uhaay64q2_0),.clk(gclk));
	jdff dff_A_wmNJ4NLZ6_0(.dout(w_dff_A_bpGILDte4_0),.din(w_dff_A_wmNJ4NLZ6_0),.clk(gclk));
	jdff dff_A_bpGILDte4_0(.dout(w_dff_A_yiPhruxa3_0),.din(w_dff_A_bpGILDte4_0),.clk(gclk));
	jdff dff_A_yiPhruxa3_0(.dout(w_dff_A_aC4K7Shp1_0),.din(w_dff_A_yiPhruxa3_0),.clk(gclk));
	jdff dff_A_aC4K7Shp1_0(.dout(w_dff_A_KB6IMC2P3_0),.din(w_dff_A_aC4K7Shp1_0),.clk(gclk));
	jdff dff_A_KB6IMC2P3_0(.dout(w_dff_A_HZmqnJB74_0),.din(w_dff_A_KB6IMC2P3_0),.clk(gclk));
	jdff dff_A_HZmqnJB74_0(.dout(w_dff_A_oyuTAxmT1_0),.din(w_dff_A_HZmqnJB74_0),.clk(gclk));
	jdff dff_A_oyuTAxmT1_0(.dout(w_dff_A_IflzbrZW3_0),.din(w_dff_A_oyuTAxmT1_0),.clk(gclk));
	jdff dff_A_IflzbrZW3_0(.dout(w_dff_A_xbGI44Ak3_0),.din(w_dff_A_IflzbrZW3_0),.clk(gclk));
	jdff dff_A_xbGI44Ak3_0(.dout(w_dff_A_fSU4pXCM5_0),.din(w_dff_A_xbGI44Ak3_0),.clk(gclk));
	jdff dff_A_fSU4pXCM5_0(.dout(w_dff_A_QQ0lJoft1_0),.din(w_dff_A_fSU4pXCM5_0),.clk(gclk));
	jdff dff_A_QQ0lJoft1_0(.dout(w_dff_A_JqtMtWun6_0),.din(w_dff_A_QQ0lJoft1_0),.clk(gclk));
	jdff dff_A_JqtMtWun6_0(.dout(w_dff_A_kv7h2Yzn8_0),.din(w_dff_A_JqtMtWun6_0),.clk(gclk));
	jdff dff_A_kv7h2Yzn8_0(.dout(w_dff_A_tKN3LHxy9_0),.din(w_dff_A_kv7h2Yzn8_0),.clk(gclk));
	jdff dff_A_tKN3LHxy9_0(.dout(w_dff_A_DsBILMrL1_0),.din(w_dff_A_tKN3LHxy9_0),.clk(gclk));
	jdff dff_A_DsBILMrL1_0(.dout(w_dff_A_33D6SsAU4_0),.din(w_dff_A_DsBILMrL1_0),.clk(gclk));
	jdff dff_A_33D6SsAU4_0(.dout(w_dff_A_hcMwm2DF9_0),.din(w_dff_A_33D6SsAU4_0),.clk(gclk));
	jdff dff_A_hcMwm2DF9_0(.dout(w_dff_A_bLdxEBzI7_0),.din(w_dff_A_hcMwm2DF9_0),.clk(gclk));
	jdff dff_A_bLdxEBzI7_0(.dout(w_dff_A_feBtEQQh4_0),.din(w_dff_A_bLdxEBzI7_0),.clk(gclk));
	jdff dff_A_feBtEQQh4_0(.dout(w_dff_A_6pYcdlUK1_0),.din(w_dff_A_feBtEQQh4_0),.clk(gclk));
	jdff dff_A_6pYcdlUK1_0(.dout(w_dff_A_YB4C5e1F9_0),.din(w_dff_A_6pYcdlUK1_0),.clk(gclk));
	jdff dff_A_YB4C5e1F9_0(.dout(w_dff_A_8OiCmwzk0_0),.din(w_dff_A_YB4C5e1F9_0),.clk(gclk));
	jdff dff_A_8OiCmwzk0_0(.dout(w_dff_A_rDGj7Q1i0_0),.din(w_dff_A_8OiCmwzk0_0),.clk(gclk));
	jdff dff_A_rDGj7Q1i0_0(.dout(w_dff_A_FxwGHjLl7_0),.din(w_dff_A_rDGj7Q1i0_0),.clk(gclk));
	jdff dff_A_FxwGHjLl7_0(.dout(w_dff_A_8mrxMDRD8_0),.din(w_dff_A_FxwGHjLl7_0),.clk(gclk));
	jdff dff_A_8mrxMDRD8_0(.dout(w_dff_A_w5XAm7Bf9_0),.din(w_dff_A_8mrxMDRD8_0),.clk(gclk));
	jdff dff_A_w5XAm7Bf9_0(.dout(w_dff_A_uhtTf1z16_0),.din(w_dff_A_w5XAm7Bf9_0),.clk(gclk));
	jdff dff_A_uhtTf1z16_0(.dout(w_dff_A_Hi1W0WRm2_0),.din(w_dff_A_uhtTf1z16_0),.clk(gclk));
	jdff dff_A_Hi1W0WRm2_0(.dout(w_dff_A_SZ4ePauA4_0),.din(w_dff_A_Hi1W0WRm2_0),.clk(gclk));
	jdff dff_A_SZ4ePauA4_0(.dout(w_dff_A_cYOgFdTT7_0),.din(w_dff_A_SZ4ePauA4_0),.clk(gclk));
	jdff dff_A_cYOgFdTT7_0(.dout(w_dff_A_zFO9lnkS7_0),.din(w_dff_A_cYOgFdTT7_0),.clk(gclk));
	jdff dff_A_zFO9lnkS7_0(.dout(w_dff_A_QnOwsA0K0_0),.din(w_dff_A_zFO9lnkS7_0),.clk(gclk));
	jdff dff_A_QnOwsA0K0_0(.dout(w_dff_A_yUI10Bf42_0),.din(w_dff_A_QnOwsA0K0_0),.clk(gclk));
	jdff dff_A_yUI10Bf42_0(.dout(w_dff_A_SbCVwLaa2_0),.din(w_dff_A_yUI10Bf42_0),.clk(gclk));
	jdff dff_A_SbCVwLaa2_0(.dout(w_dff_A_lK38vy6x5_0),.din(w_dff_A_SbCVwLaa2_0),.clk(gclk));
	jdff dff_A_lK38vy6x5_0(.dout(w_dff_A_435CGDln8_0),.din(w_dff_A_lK38vy6x5_0),.clk(gclk));
	jdff dff_A_435CGDln8_0(.dout(w_dff_A_mnr3JpNV6_0),.din(w_dff_A_435CGDln8_0),.clk(gclk));
	jdff dff_A_mnr3JpNV6_0(.dout(w_dff_A_IMd2R1Fa5_0),.din(w_dff_A_mnr3JpNV6_0),.clk(gclk));
	jdff dff_A_IMd2R1Fa5_0(.dout(w_dff_A_KrUrWVju1_0),.din(w_dff_A_IMd2R1Fa5_0),.clk(gclk));
	jdff dff_A_KrUrWVju1_0(.dout(w_dff_A_vWNn7eQH1_0),.din(w_dff_A_KrUrWVju1_0),.clk(gclk));
	jdff dff_A_vWNn7eQH1_0(.dout(w_dff_A_vP6t7DhO5_0),.din(w_dff_A_vWNn7eQH1_0),.clk(gclk));
	jdff dff_A_vP6t7DhO5_0(.dout(w_dff_A_muhXB0j46_0),.din(w_dff_A_vP6t7DhO5_0),.clk(gclk));
	jdff dff_A_muhXB0j46_0(.dout(w_dff_A_w15OVzbB4_0),.din(w_dff_A_muhXB0j46_0),.clk(gclk));
	jdff dff_A_w15OVzbB4_0(.dout(w_dff_A_bQyoU5vk1_0),.din(w_dff_A_w15OVzbB4_0),.clk(gclk));
	jdff dff_A_bQyoU5vk1_0(.dout(w_dff_A_tsgWoKuc9_0),.din(w_dff_A_bQyoU5vk1_0),.clk(gclk));
	jdff dff_A_tsgWoKuc9_0(.dout(w_dff_A_mMoeQG1x2_0),.din(w_dff_A_tsgWoKuc9_0),.clk(gclk));
	jdff dff_A_mMoeQG1x2_0(.dout(w_dff_A_GZeM7Lgj3_0),.din(w_dff_A_mMoeQG1x2_0),.clk(gclk));
	jdff dff_A_GZeM7Lgj3_0(.dout(w_dff_A_Tcs5UMHB1_0),.din(w_dff_A_GZeM7Lgj3_0),.clk(gclk));
	jdff dff_A_Tcs5UMHB1_0(.dout(w_dff_A_mVINKIeB2_0),.din(w_dff_A_Tcs5UMHB1_0),.clk(gclk));
	jdff dff_A_mVINKIeB2_0(.dout(w_dff_A_4yW2qVps5_0),.din(w_dff_A_mVINKIeB2_0),.clk(gclk));
	jdff dff_A_4yW2qVps5_0(.dout(w_dff_A_ioWvvnrU1_0),.din(w_dff_A_4yW2qVps5_0),.clk(gclk));
	jdff dff_A_ioWvvnrU1_0(.dout(w_dff_A_QVFiNPEC8_0),.din(w_dff_A_ioWvvnrU1_0),.clk(gclk));
	jdff dff_A_QVFiNPEC8_0(.dout(w_dff_A_Koe9jSw08_0),.din(w_dff_A_QVFiNPEC8_0),.clk(gclk));
	jdff dff_A_Koe9jSw08_0(.dout(w_dff_A_RCzhCTvV3_0),.din(w_dff_A_Koe9jSw08_0),.clk(gclk));
	jdff dff_A_RCzhCTvV3_0(.dout(w_dff_A_y0RdezRs4_0),.din(w_dff_A_RCzhCTvV3_0),.clk(gclk));
	jdff dff_A_y0RdezRs4_0(.dout(w_dff_A_IKfcsEwg4_0),.din(w_dff_A_y0RdezRs4_0),.clk(gclk));
	jdff dff_A_IKfcsEwg4_0(.dout(w_dff_A_MHankf090_0),.din(w_dff_A_IKfcsEwg4_0),.clk(gclk));
	jdff dff_A_MHankf090_0(.dout(w_dff_A_uvgGtS777_0),.din(w_dff_A_MHankf090_0),.clk(gclk));
	jdff dff_A_uvgGtS777_0(.dout(w_dff_A_jYvkSs9A3_0),.din(w_dff_A_uvgGtS777_0),.clk(gclk));
	jdff dff_A_jYvkSs9A3_0(.dout(w_dff_A_VSOwTyg44_0),.din(w_dff_A_jYvkSs9A3_0),.clk(gclk));
	jdff dff_A_VSOwTyg44_0(.dout(w_dff_A_ZpoxRcY69_0),.din(w_dff_A_VSOwTyg44_0),.clk(gclk));
	jdff dff_A_ZpoxRcY69_0(.dout(w_dff_A_k9ra6rwE2_0),.din(w_dff_A_ZpoxRcY69_0),.clk(gclk));
	jdff dff_A_k9ra6rwE2_0(.dout(w_dff_A_prvXHNpo0_0),.din(w_dff_A_k9ra6rwE2_0),.clk(gclk));
	jdff dff_A_prvXHNpo0_0(.dout(w_dff_A_dgwlu9WA5_0),.din(w_dff_A_prvXHNpo0_0),.clk(gclk));
	jdff dff_A_dgwlu9WA5_0(.dout(w_dff_A_uxnVYdDa8_0),.din(w_dff_A_dgwlu9WA5_0),.clk(gclk));
	jdff dff_A_uxnVYdDa8_0(.dout(w_dff_A_6LswrDbN6_0),.din(w_dff_A_uxnVYdDa8_0),.clk(gclk));
	jdff dff_A_6LswrDbN6_0(.dout(w_dff_A_GfsIvQtw0_0),.din(w_dff_A_6LswrDbN6_0),.clk(gclk));
	jdff dff_A_GfsIvQtw0_0(.dout(w_dff_A_KSLFMHLk7_0),.din(w_dff_A_GfsIvQtw0_0),.clk(gclk));
	jdff dff_A_KSLFMHLk7_0(.dout(w_dff_A_sQckYULF7_0),.din(w_dff_A_KSLFMHLk7_0),.clk(gclk));
	jdff dff_A_sQckYULF7_0(.dout(w_dff_A_OmyVFBLf8_0),.din(w_dff_A_sQckYULF7_0),.clk(gclk));
	jdff dff_A_OmyVFBLf8_0(.dout(w_dff_A_3Lb1IWRL3_0),.din(w_dff_A_OmyVFBLf8_0),.clk(gclk));
	jdff dff_A_3Lb1IWRL3_0(.dout(w_dff_A_NSTjunAr1_0),.din(w_dff_A_3Lb1IWRL3_0),.clk(gclk));
	jdff dff_A_NSTjunAr1_0(.dout(w_dff_A_BkhXo2AL4_0),.din(w_dff_A_NSTjunAr1_0),.clk(gclk));
	jdff dff_A_BkhXo2AL4_0(.dout(w_dff_A_xaEYEOJW9_0),.din(w_dff_A_BkhXo2AL4_0),.clk(gclk));
	jdff dff_A_xaEYEOJW9_0(.dout(w_dff_A_D4qYnBMC2_0),.din(w_dff_A_xaEYEOJW9_0),.clk(gclk));
	jdff dff_A_D4qYnBMC2_0(.dout(w_dff_A_w0dYMDYg0_0),.din(w_dff_A_D4qYnBMC2_0),.clk(gclk));
	jdff dff_A_w0dYMDYg0_0(.dout(w_dff_A_getjz7V28_0),.din(w_dff_A_w0dYMDYg0_0),.clk(gclk));
	jdff dff_A_getjz7V28_0(.dout(w_dff_A_7LpYKxFt5_0),.din(w_dff_A_getjz7V28_0),.clk(gclk));
	jdff dff_A_7LpYKxFt5_0(.dout(w_dff_A_28W5aH2K6_0),.din(w_dff_A_7LpYKxFt5_0),.clk(gclk));
	jdff dff_A_28W5aH2K6_0(.dout(w_dff_A_U5RnASk11_0),.din(w_dff_A_28W5aH2K6_0),.clk(gclk));
	jdff dff_A_U5RnASk11_0(.dout(w_dff_A_r0GVk2Pe7_0),.din(w_dff_A_U5RnASk11_0),.clk(gclk));
	jdff dff_A_r0GVk2Pe7_0(.dout(w_dff_A_TBVMeCGo8_0),.din(w_dff_A_r0GVk2Pe7_0),.clk(gclk));
	jdff dff_A_TBVMeCGo8_0(.dout(w_dff_A_ErTjsSXk7_0),.din(w_dff_A_TBVMeCGo8_0),.clk(gclk));
	jdff dff_A_ErTjsSXk7_0(.dout(w_dff_A_2OZLHZDr4_0),.din(w_dff_A_ErTjsSXk7_0),.clk(gclk));
	jdff dff_A_2OZLHZDr4_0(.dout(w_dff_A_2ZqmUP6w1_0),.din(w_dff_A_2OZLHZDr4_0),.clk(gclk));
	jdff dff_A_2ZqmUP6w1_0(.dout(w_dff_A_1riIuvg58_0),.din(w_dff_A_2ZqmUP6w1_0),.clk(gclk));
	jdff dff_A_1riIuvg58_0(.dout(w_dff_A_CBWZWl9S5_0),.din(w_dff_A_1riIuvg58_0),.clk(gclk));
	jdff dff_A_CBWZWl9S5_0(.dout(w_dff_A_sx9ATPQC2_0),.din(w_dff_A_CBWZWl9S5_0),.clk(gclk));
	jdff dff_A_sx9ATPQC2_0(.dout(w_dff_A_6OrMUFPu2_0),.din(w_dff_A_sx9ATPQC2_0),.clk(gclk));
	jdff dff_A_6OrMUFPu2_0(.dout(w_dff_A_kf5oJuF46_0),.din(w_dff_A_6OrMUFPu2_0),.clk(gclk));
	jdff dff_A_kf5oJuF46_0(.dout(w_dff_A_PFaQGYxK9_0),.din(w_dff_A_kf5oJuF46_0),.clk(gclk));
	jdff dff_A_PFaQGYxK9_0(.dout(w_dff_A_pPuynFWl5_0),.din(w_dff_A_PFaQGYxK9_0),.clk(gclk));
	jdff dff_A_pPuynFWl5_0(.dout(w_dff_A_XfMAWmc97_0),.din(w_dff_A_pPuynFWl5_0),.clk(gclk));
	jdff dff_A_XfMAWmc97_0(.dout(w_dff_A_gQEtfDcs9_0),.din(w_dff_A_XfMAWmc97_0),.clk(gclk));
	jdff dff_A_gQEtfDcs9_0(.dout(f8),.din(w_dff_A_gQEtfDcs9_0),.clk(gclk));
	jdff dff_A_TPd6RMHY6_2(.dout(w_dff_A_5qhc1AdK0_0),.din(w_dff_A_TPd6RMHY6_2),.clk(gclk));
	jdff dff_A_5qhc1AdK0_0(.dout(w_dff_A_oKwebBb92_0),.din(w_dff_A_5qhc1AdK0_0),.clk(gclk));
	jdff dff_A_oKwebBb92_0(.dout(w_dff_A_ELgAvyqV1_0),.din(w_dff_A_oKwebBb92_0),.clk(gclk));
	jdff dff_A_ELgAvyqV1_0(.dout(w_dff_A_Fo1cNxNA2_0),.din(w_dff_A_ELgAvyqV1_0),.clk(gclk));
	jdff dff_A_Fo1cNxNA2_0(.dout(w_dff_A_C4diHBCU1_0),.din(w_dff_A_Fo1cNxNA2_0),.clk(gclk));
	jdff dff_A_C4diHBCU1_0(.dout(w_dff_A_uG1H5xEk7_0),.din(w_dff_A_C4diHBCU1_0),.clk(gclk));
	jdff dff_A_uG1H5xEk7_0(.dout(w_dff_A_VjwGpPpD4_0),.din(w_dff_A_uG1H5xEk7_0),.clk(gclk));
	jdff dff_A_VjwGpPpD4_0(.dout(w_dff_A_oFbnVh4y7_0),.din(w_dff_A_VjwGpPpD4_0),.clk(gclk));
	jdff dff_A_oFbnVh4y7_0(.dout(w_dff_A_BGYlffrk1_0),.din(w_dff_A_oFbnVh4y7_0),.clk(gclk));
	jdff dff_A_BGYlffrk1_0(.dout(w_dff_A_Rvpn2TQb6_0),.din(w_dff_A_BGYlffrk1_0),.clk(gclk));
	jdff dff_A_Rvpn2TQb6_0(.dout(w_dff_A_TuUKr8CC7_0),.din(w_dff_A_Rvpn2TQb6_0),.clk(gclk));
	jdff dff_A_TuUKr8CC7_0(.dout(w_dff_A_Kr0BLb9U2_0),.din(w_dff_A_TuUKr8CC7_0),.clk(gclk));
	jdff dff_A_Kr0BLb9U2_0(.dout(w_dff_A_C8WuXlrQ4_0),.din(w_dff_A_Kr0BLb9U2_0),.clk(gclk));
	jdff dff_A_C8WuXlrQ4_0(.dout(w_dff_A_fJE7ZlUa4_0),.din(w_dff_A_C8WuXlrQ4_0),.clk(gclk));
	jdff dff_A_fJE7ZlUa4_0(.dout(w_dff_A_ng8tJ7AN0_0),.din(w_dff_A_fJE7ZlUa4_0),.clk(gclk));
	jdff dff_A_ng8tJ7AN0_0(.dout(w_dff_A_gTG3JZtX0_0),.din(w_dff_A_ng8tJ7AN0_0),.clk(gclk));
	jdff dff_A_gTG3JZtX0_0(.dout(w_dff_A_pdKGmA085_0),.din(w_dff_A_gTG3JZtX0_0),.clk(gclk));
	jdff dff_A_pdKGmA085_0(.dout(w_dff_A_9jyAnHEI8_0),.din(w_dff_A_pdKGmA085_0),.clk(gclk));
	jdff dff_A_9jyAnHEI8_0(.dout(w_dff_A_soDGOWyV4_0),.din(w_dff_A_9jyAnHEI8_0),.clk(gclk));
	jdff dff_A_soDGOWyV4_0(.dout(w_dff_A_J540FnmE3_0),.din(w_dff_A_soDGOWyV4_0),.clk(gclk));
	jdff dff_A_J540FnmE3_0(.dout(w_dff_A_oapD8LyZ5_0),.din(w_dff_A_J540FnmE3_0),.clk(gclk));
	jdff dff_A_oapD8LyZ5_0(.dout(w_dff_A_ekk7WLap6_0),.din(w_dff_A_oapD8LyZ5_0),.clk(gclk));
	jdff dff_A_ekk7WLap6_0(.dout(w_dff_A_odu7KFF12_0),.din(w_dff_A_ekk7WLap6_0),.clk(gclk));
	jdff dff_A_odu7KFF12_0(.dout(w_dff_A_5O5Xh0b56_0),.din(w_dff_A_odu7KFF12_0),.clk(gclk));
	jdff dff_A_5O5Xh0b56_0(.dout(w_dff_A_0dyfs50F7_0),.din(w_dff_A_5O5Xh0b56_0),.clk(gclk));
	jdff dff_A_0dyfs50F7_0(.dout(w_dff_A_8MJ5XxQ18_0),.din(w_dff_A_0dyfs50F7_0),.clk(gclk));
	jdff dff_A_8MJ5XxQ18_0(.dout(w_dff_A_YfwHMbUa5_0),.din(w_dff_A_8MJ5XxQ18_0),.clk(gclk));
	jdff dff_A_YfwHMbUa5_0(.dout(w_dff_A_4rG5yjCy7_0),.din(w_dff_A_YfwHMbUa5_0),.clk(gclk));
	jdff dff_A_4rG5yjCy7_0(.dout(w_dff_A_Xw86b9FC6_0),.din(w_dff_A_4rG5yjCy7_0),.clk(gclk));
	jdff dff_A_Xw86b9FC6_0(.dout(w_dff_A_Qs1lpwUU0_0),.din(w_dff_A_Xw86b9FC6_0),.clk(gclk));
	jdff dff_A_Qs1lpwUU0_0(.dout(w_dff_A_JiPUreyM7_0),.din(w_dff_A_Qs1lpwUU0_0),.clk(gclk));
	jdff dff_A_JiPUreyM7_0(.dout(w_dff_A_jvkWY0FK8_0),.din(w_dff_A_JiPUreyM7_0),.clk(gclk));
	jdff dff_A_jvkWY0FK8_0(.dout(w_dff_A_zUZYuJGC7_0),.din(w_dff_A_jvkWY0FK8_0),.clk(gclk));
	jdff dff_A_zUZYuJGC7_0(.dout(w_dff_A_wWAf9Xjw7_0),.din(w_dff_A_zUZYuJGC7_0),.clk(gclk));
	jdff dff_A_wWAf9Xjw7_0(.dout(w_dff_A_81tWg6aq9_0),.din(w_dff_A_wWAf9Xjw7_0),.clk(gclk));
	jdff dff_A_81tWg6aq9_0(.dout(w_dff_A_P0IYBxEW8_0),.din(w_dff_A_81tWg6aq9_0),.clk(gclk));
	jdff dff_A_P0IYBxEW8_0(.dout(w_dff_A_mrvY481p7_0),.din(w_dff_A_P0IYBxEW8_0),.clk(gclk));
	jdff dff_A_mrvY481p7_0(.dout(w_dff_A_vHQRbkbV7_0),.din(w_dff_A_mrvY481p7_0),.clk(gclk));
	jdff dff_A_vHQRbkbV7_0(.dout(w_dff_A_F0mOwgfQ5_0),.din(w_dff_A_vHQRbkbV7_0),.clk(gclk));
	jdff dff_A_F0mOwgfQ5_0(.dout(w_dff_A_yWa4bRM23_0),.din(w_dff_A_F0mOwgfQ5_0),.clk(gclk));
	jdff dff_A_yWa4bRM23_0(.dout(w_dff_A_yI9ITnt29_0),.din(w_dff_A_yWa4bRM23_0),.clk(gclk));
	jdff dff_A_yI9ITnt29_0(.dout(w_dff_A_nkufeQnA9_0),.din(w_dff_A_yI9ITnt29_0),.clk(gclk));
	jdff dff_A_nkufeQnA9_0(.dout(w_dff_A_nTY9AT0U0_0),.din(w_dff_A_nkufeQnA9_0),.clk(gclk));
	jdff dff_A_nTY9AT0U0_0(.dout(w_dff_A_S4GDwsci3_0),.din(w_dff_A_nTY9AT0U0_0),.clk(gclk));
	jdff dff_A_S4GDwsci3_0(.dout(w_dff_A_ZhhuA6U36_0),.din(w_dff_A_S4GDwsci3_0),.clk(gclk));
	jdff dff_A_ZhhuA6U36_0(.dout(w_dff_A_okZIWMFN2_0),.din(w_dff_A_ZhhuA6U36_0),.clk(gclk));
	jdff dff_A_okZIWMFN2_0(.dout(w_dff_A_MJUYoofZ8_0),.din(w_dff_A_okZIWMFN2_0),.clk(gclk));
	jdff dff_A_MJUYoofZ8_0(.dout(w_dff_A_bnwczqnS6_0),.din(w_dff_A_MJUYoofZ8_0),.clk(gclk));
	jdff dff_A_bnwczqnS6_0(.dout(w_dff_A_XhCA6d1Z8_0),.din(w_dff_A_bnwczqnS6_0),.clk(gclk));
	jdff dff_A_XhCA6d1Z8_0(.dout(w_dff_A_lYO78a6M6_0),.din(w_dff_A_XhCA6d1Z8_0),.clk(gclk));
	jdff dff_A_lYO78a6M6_0(.dout(w_dff_A_TEOSqEFu7_0),.din(w_dff_A_lYO78a6M6_0),.clk(gclk));
	jdff dff_A_TEOSqEFu7_0(.dout(w_dff_A_1vOBBOuH5_0),.din(w_dff_A_TEOSqEFu7_0),.clk(gclk));
	jdff dff_A_1vOBBOuH5_0(.dout(w_dff_A_RHaFhZBA5_0),.din(w_dff_A_1vOBBOuH5_0),.clk(gclk));
	jdff dff_A_RHaFhZBA5_0(.dout(w_dff_A_cAjkRbEU0_0),.din(w_dff_A_RHaFhZBA5_0),.clk(gclk));
	jdff dff_A_cAjkRbEU0_0(.dout(w_dff_A_a2hoNyqg4_0),.din(w_dff_A_cAjkRbEU0_0),.clk(gclk));
	jdff dff_A_a2hoNyqg4_0(.dout(w_dff_A_uIWdLd6w0_0),.din(w_dff_A_a2hoNyqg4_0),.clk(gclk));
	jdff dff_A_uIWdLd6w0_0(.dout(w_dff_A_bGLF6RKs0_0),.din(w_dff_A_uIWdLd6w0_0),.clk(gclk));
	jdff dff_A_bGLF6RKs0_0(.dout(w_dff_A_UOjJV8NZ0_0),.din(w_dff_A_bGLF6RKs0_0),.clk(gclk));
	jdff dff_A_UOjJV8NZ0_0(.dout(w_dff_A_gE4pJxjk0_0),.din(w_dff_A_UOjJV8NZ0_0),.clk(gclk));
	jdff dff_A_gE4pJxjk0_0(.dout(w_dff_A_ZvmtSwUG1_0),.din(w_dff_A_gE4pJxjk0_0),.clk(gclk));
	jdff dff_A_ZvmtSwUG1_0(.dout(w_dff_A_MXobBHJP2_0),.din(w_dff_A_ZvmtSwUG1_0),.clk(gclk));
	jdff dff_A_MXobBHJP2_0(.dout(w_dff_A_hebXh9ER7_0),.din(w_dff_A_MXobBHJP2_0),.clk(gclk));
	jdff dff_A_hebXh9ER7_0(.dout(w_dff_A_SRDDYPek9_0),.din(w_dff_A_hebXh9ER7_0),.clk(gclk));
	jdff dff_A_SRDDYPek9_0(.dout(w_dff_A_evICsUMv8_0),.din(w_dff_A_SRDDYPek9_0),.clk(gclk));
	jdff dff_A_evICsUMv8_0(.dout(w_dff_A_f3h2CkNv2_0),.din(w_dff_A_evICsUMv8_0),.clk(gclk));
	jdff dff_A_f3h2CkNv2_0(.dout(w_dff_A_iQBt9nmS5_0),.din(w_dff_A_f3h2CkNv2_0),.clk(gclk));
	jdff dff_A_iQBt9nmS5_0(.dout(w_dff_A_SziMIP2j1_0),.din(w_dff_A_iQBt9nmS5_0),.clk(gclk));
	jdff dff_A_SziMIP2j1_0(.dout(w_dff_A_UJJV25nb3_0),.din(w_dff_A_SziMIP2j1_0),.clk(gclk));
	jdff dff_A_UJJV25nb3_0(.dout(w_dff_A_uYoSwYDn7_0),.din(w_dff_A_UJJV25nb3_0),.clk(gclk));
	jdff dff_A_uYoSwYDn7_0(.dout(w_dff_A_ts7zJ5Tb7_0),.din(w_dff_A_uYoSwYDn7_0),.clk(gclk));
	jdff dff_A_ts7zJ5Tb7_0(.dout(w_dff_A_F6w6UlAx6_0),.din(w_dff_A_ts7zJ5Tb7_0),.clk(gclk));
	jdff dff_A_F6w6UlAx6_0(.dout(w_dff_A_sYp8UMwn9_0),.din(w_dff_A_F6w6UlAx6_0),.clk(gclk));
	jdff dff_A_sYp8UMwn9_0(.dout(w_dff_A_EJo59HU06_0),.din(w_dff_A_sYp8UMwn9_0),.clk(gclk));
	jdff dff_A_EJo59HU06_0(.dout(w_dff_A_pbbhVIpa0_0),.din(w_dff_A_EJo59HU06_0),.clk(gclk));
	jdff dff_A_pbbhVIpa0_0(.dout(w_dff_A_AFHu6rDq3_0),.din(w_dff_A_pbbhVIpa0_0),.clk(gclk));
	jdff dff_A_AFHu6rDq3_0(.dout(w_dff_A_sN6r5Psz8_0),.din(w_dff_A_AFHu6rDq3_0),.clk(gclk));
	jdff dff_A_sN6r5Psz8_0(.dout(w_dff_A_9zncHu7w2_0),.din(w_dff_A_sN6r5Psz8_0),.clk(gclk));
	jdff dff_A_9zncHu7w2_0(.dout(w_dff_A_Ixb7AvpI6_0),.din(w_dff_A_9zncHu7w2_0),.clk(gclk));
	jdff dff_A_Ixb7AvpI6_0(.dout(w_dff_A_d2qge45n1_0),.din(w_dff_A_Ixb7AvpI6_0),.clk(gclk));
	jdff dff_A_d2qge45n1_0(.dout(w_dff_A_gploWS1K6_0),.din(w_dff_A_d2qge45n1_0),.clk(gclk));
	jdff dff_A_gploWS1K6_0(.dout(w_dff_A_a1G9LEd90_0),.din(w_dff_A_gploWS1K6_0),.clk(gclk));
	jdff dff_A_a1G9LEd90_0(.dout(w_dff_A_VKvFcBOQ3_0),.din(w_dff_A_a1G9LEd90_0),.clk(gclk));
	jdff dff_A_VKvFcBOQ3_0(.dout(w_dff_A_kPzPb2ib5_0),.din(w_dff_A_VKvFcBOQ3_0),.clk(gclk));
	jdff dff_A_kPzPb2ib5_0(.dout(w_dff_A_KT5Pzb5p2_0),.din(w_dff_A_kPzPb2ib5_0),.clk(gclk));
	jdff dff_A_KT5Pzb5p2_0(.dout(w_dff_A_2UifLQiR5_0),.din(w_dff_A_KT5Pzb5p2_0),.clk(gclk));
	jdff dff_A_2UifLQiR5_0(.dout(w_dff_A_WOZEytYC2_0),.din(w_dff_A_2UifLQiR5_0),.clk(gclk));
	jdff dff_A_WOZEytYC2_0(.dout(w_dff_A_VKkH7hu57_0),.din(w_dff_A_WOZEytYC2_0),.clk(gclk));
	jdff dff_A_VKkH7hu57_0(.dout(w_dff_A_8ovRG4gm6_0),.din(w_dff_A_VKkH7hu57_0),.clk(gclk));
	jdff dff_A_8ovRG4gm6_0(.dout(w_dff_A_coIA58xT9_0),.din(w_dff_A_8ovRG4gm6_0),.clk(gclk));
	jdff dff_A_coIA58xT9_0(.dout(w_dff_A_5lQMfcsz7_0),.din(w_dff_A_coIA58xT9_0),.clk(gclk));
	jdff dff_A_5lQMfcsz7_0(.dout(w_dff_A_HydVFWFi0_0),.din(w_dff_A_5lQMfcsz7_0),.clk(gclk));
	jdff dff_A_HydVFWFi0_0(.dout(w_dff_A_cbBspt3o2_0),.din(w_dff_A_HydVFWFi0_0),.clk(gclk));
	jdff dff_A_cbBspt3o2_0(.dout(w_dff_A_Cug2ntA18_0),.din(w_dff_A_cbBspt3o2_0),.clk(gclk));
	jdff dff_A_Cug2ntA18_0(.dout(w_dff_A_JItWcIBc7_0),.din(w_dff_A_Cug2ntA18_0),.clk(gclk));
	jdff dff_A_JItWcIBc7_0(.dout(w_dff_A_YfheOsXd8_0),.din(w_dff_A_JItWcIBc7_0),.clk(gclk));
	jdff dff_A_YfheOsXd8_0(.dout(w_dff_A_bXFhU7yJ8_0),.din(w_dff_A_YfheOsXd8_0),.clk(gclk));
	jdff dff_A_bXFhU7yJ8_0(.dout(w_dff_A_fqp1ss0R2_0),.din(w_dff_A_bXFhU7yJ8_0),.clk(gclk));
	jdff dff_A_fqp1ss0R2_0(.dout(w_dff_A_aW1GduXA8_0),.din(w_dff_A_fqp1ss0R2_0),.clk(gclk));
	jdff dff_A_aW1GduXA8_0(.dout(w_dff_A_qgbVWWsa7_0),.din(w_dff_A_aW1GduXA8_0),.clk(gclk));
	jdff dff_A_qgbVWWsa7_0(.dout(w_dff_A_2dzkjre17_0),.din(w_dff_A_qgbVWWsa7_0),.clk(gclk));
	jdff dff_A_2dzkjre17_0(.dout(w_dff_A_ti3AE9Nx9_0),.din(w_dff_A_2dzkjre17_0),.clk(gclk));
	jdff dff_A_ti3AE9Nx9_0(.dout(w_dff_A_3PPjiAZw2_0),.din(w_dff_A_ti3AE9Nx9_0),.clk(gclk));
	jdff dff_A_3PPjiAZw2_0(.dout(w_dff_A_GblVuIFG4_0),.din(w_dff_A_3PPjiAZw2_0),.clk(gclk));
	jdff dff_A_GblVuIFG4_0(.dout(w_dff_A_orpG6eH67_0),.din(w_dff_A_GblVuIFG4_0),.clk(gclk));
	jdff dff_A_orpG6eH67_0(.dout(w_dff_A_AoYMz5245_0),.din(w_dff_A_orpG6eH67_0),.clk(gclk));
	jdff dff_A_AoYMz5245_0(.dout(w_dff_A_jP4YGIUT1_0),.din(w_dff_A_AoYMz5245_0),.clk(gclk));
	jdff dff_A_jP4YGIUT1_0(.dout(w_dff_A_B3R1hoNp8_0),.din(w_dff_A_jP4YGIUT1_0),.clk(gclk));
	jdff dff_A_B3R1hoNp8_0(.dout(w_dff_A_g0A8uaiE3_0),.din(w_dff_A_B3R1hoNp8_0),.clk(gclk));
	jdff dff_A_g0A8uaiE3_0(.dout(w_dff_A_Qqr0eMQf2_0),.din(w_dff_A_g0A8uaiE3_0),.clk(gclk));
	jdff dff_A_Qqr0eMQf2_0(.dout(w_dff_A_gk7QQ19M1_0),.din(w_dff_A_Qqr0eMQf2_0),.clk(gclk));
	jdff dff_A_gk7QQ19M1_0(.dout(w_dff_A_cICvejxt9_0),.din(w_dff_A_gk7QQ19M1_0),.clk(gclk));
	jdff dff_A_cICvejxt9_0(.dout(w_dff_A_g7qhwGua2_0),.din(w_dff_A_cICvejxt9_0),.clk(gclk));
	jdff dff_A_g7qhwGua2_0(.dout(w_dff_A_0YxtZ9R23_0),.din(w_dff_A_g7qhwGua2_0),.clk(gclk));
	jdff dff_A_0YxtZ9R23_0(.dout(w_dff_A_lmO3bB5r4_0),.din(w_dff_A_0YxtZ9R23_0),.clk(gclk));
	jdff dff_A_lmO3bB5r4_0(.dout(w_dff_A_Vn8QyEAP3_0),.din(w_dff_A_lmO3bB5r4_0),.clk(gclk));
	jdff dff_A_Vn8QyEAP3_0(.dout(w_dff_A_CCCqz7dS7_0),.din(w_dff_A_Vn8QyEAP3_0),.clk(gclk));
	jdff dff_A_CCCqz7dS7_0(.dout(w_dff_A_GSewm7ZW8_0),.din(w_dff_A_CCCqz7dS7_0),.clk(gclk));
	jdff dff_A_GSewm7ZW8_0(.dout(f9),.din(w_dff_A_GSewm7ZW8_0),.clk(gclk));
	jdff dff_A_K99ijCAz4_2(.dout(w_dff_A_jjVoD3AR3_0),.din(w_dff_A_K99ijCAz4_2),.clk(gclk));
	jdff dff_A_jjVoD3AR3_0(.dout(w_dff_A_760m2NFX7_0),.din(w_dff_A_jjVoD3AR3_0),.clk(gclk));
	jdff dff_A_760m2NFX7_0(.dout(w_dff_A_iu1oGKb55_0),.din(w_dff_A_760m2NFX7_0),.clk(gclk));
	jdff dff_A_iu1oGKb55_0(.dout(w_dff_A_Pb5Ssgcu6_0),.din(w_dff_A_iu1oGKb55_0),.clk(gclk));
	jdff dff_A_Pb5Ssgcu6_0(.dout(w_dff_A_Czh0R1hf9_0),.din(w_dff_A_Pb5Ssgcu6_0),.clk(gclk));
	jdff dff_A_Czh0R1hf9_0(.dout(w_dff_A_uMob2VTh3_0),.din(w_dff_A_Czh0R1hf9_0),.clk(gclk));
	jdff dff_A_uMob2VTh3_0(.dout(w_dff_A_4mW44HZk6_0),.din(w_dff_A_uMob2VTh3_0),.clk(gclk));
	jdff dff_A_4mW44HZk6_0(.dout(w_dff_A_awGgXWEf0_0),.din(w_dff_A_4mW44HZk6_0),.clk(gclk));
	jdff dff_A_awGgXWEf0_0(.dout(w_dff_A_Efs3Kc2K5_0),.din(w_dff_A_awGgXWEf0_0),.clk(gclk));
	jdff dff_A_Efs3Kc2K5_0(.dout(w_dff_A_KNXOpXvx0_0),.din(w_dff_A_Efs3Kc2K5_0),.clk(gclk));
	jdff dff_A_KNXOpXvx0_0(.dout(w_dff_A_XOKGgzQL0_0),.din(w_dff_A_KNXOpXvx0_0),.clk(gclk));
	jdff dff_A_XOKGgzQL0_0(.dout(w_dff_A_MvhTjEBJ9_0),.din(w_dff_A_XOKGgzQL0_0),.clk(gclk));
	jdff dff_A_MvhTjEBJ9_0(.dout(w_dff_A_aAZ6A1kX5_0),.din(w_dff_A_MvhTjEBJ9_0),.clk(gclk));
	jdff dff_A_aAZ6A1kX5_0(.dout(w_dff_A_IGLhGCm57_0),.din(w_dff_A_aAZ6A1kX5_0),.clk(gclk));
	jdff dff_A_IGLhGCm57_0(.dout(w_dff_A_B0VJY4VC9_0),.din(w_dff_A_IGLhGCm57_0),.clk(gclk));
	jdff dff_A_B0VJY4VC9_0(.dout(w_dff_A_UsEBKtdf5_0),.din(w_dff_A_B0VJY4VC9_0),.clk(gclk));
	jdff dff_A_UsEBKtdf5_0(.dout(w_dff_A_zHZPFIvM2_0),.din(w_dff_A_UsEBKtdf5_0),.clk(gclk));
	jdff dff_A_zHZPFIvM2_0(.dout(w_dff_A_vDSd9rkY7_0),.din(w_dff_A_zHZPFIvM2_0),.clk(gclk));
	jdff dff_A_vDSd9rkY7_0(.dout(w_dff_A_WYATVSAs8_0),.din(w_dff_A_vDSd9rkY7_0),.clk(gclk));
	jdff dff_A_WYATVSAs8_0(.dout(w_dff_A_jIQYJQWf5_0),.din(w_dff_A_WYATVSAs8_0),.clk(gclk));
	jdff dff_A_jIQYJQWf5_0(.dout(w_dff_A_SDmt4iOz2_0),.din(w_dff_A_jIQYJQWf5_0),.clk(gclk));
	jdff dff_A_SDmt4iOz2_0(.dout(w_dff_A_iKBXCCy35_0),.din(w_dff_A_SDmt4iOz2_0),.clk(gclk));
	jdff dff_A_iKBXCCy35_0(.dout(w_dff_A_8oz9Wyhx9_0),.din(w_dff_A_iKBXCCy35_0),.clk(gclk));
	jdff dff_A_8oz9Wyhx9_0(.dout(w_dff_A_5fPehC8h2_0),.din(w_dff_A_8oz9Wyhx9_0),.clk(gclk));
	jdff dff_A_5fPehC8h2_0(.dout(w_dff_A_q02Z14UO1_0),.din(w_dff_A_5fPehC8h2_0),.clk(gclk));
	jdff dff_A_q02Z14UO1_0(.dout(w_dff_A_k0u9xkPa3_0),.din(w_dff_A_q02Z14UO1_0),.clk(gclk));
	jdff dff_A_k0u9xkPa3_0(.dout(w_dff_A_A4EBHP5a6_0),.din(w_dff_A_k0u9xkPa3_0),.clk(gclk));
	jdff dff_A_A4EBHP5a6_0(.dout(w_dff_A_JXLuhsgi7_0),.din(w_dff_A_A4EBHP5a6_0),.clk(gclk));
	jdff dff_A_JXLuhsgi7_0(.dout(w_dff_A_fT2p0KIq1_0),.din(w_dff_A_JXLuhsgi7_0),.clk(gclk));
	jdff dff_A_fT2p0KIq1_0(.dout(w_dff_A_Y6hv9qId6_0),.din(w_dff_A_fT2p0KIq1_0),.clk(gclk));
	jdff dff_A_Y6hv9qId6_0(.dout(w_dff_A_mMrFIkb33_0),.din(w_dff_A_Y6hv9qId6_0),.clk(gclk));
	jdff dff_A_mMrFIkb33_0(.dout(w_dff_A_OkStu4Nd7_0),.din(w_dff_A_mMrFIkb33_0),.clk(gclk));
	jdff dff_A_OkStu4Nd7_0(.dout(w_dff_A_SRX7Yj785_0),.din(w_dff_A_OkStu4Nd7_0),.clk(gclk));
	jdff dff_A_SRX7Yj785_0(.dout(w_dff_A_diBiWOwM1_0),.din(w_dff_A_SRX7Yj785_0),.clk(gclk));
	jdff dff_A_diBiWOwM1_0(.dout(w_dff_A_joy2avoE4_0),.din(w_dff_A_diBiWOwM1_0),.clk(gclk));
	jdff dff_A_joy2avoE4_0(.dout(w_dff_A_6qUWlzKo3_0),.din(w_dff_A_joy2avoE4_0),.clk(gclk));
	jdff dff_A_6qUWlzKo3_0(.dout(w_dff_A_Nw2b6nGT1_0),.din(w_dff_A_6qUWlzKo3_0),.clk(gclk));
	jdff dff_A_Nw2b6nGT1_0(.dout(w_dff_A_pGLygNaG3_0),.din(w_dff_A_Nw2b6nGT1_0),.clk(gclk));
	jdff dff_A_pGLygNaG3_0(.dout(w_dff_A_h9KHelO10_0),.din(w_dff_A_pGLygNaG3_0),.clk(gclk));
	jdff dff_A_h9KHelO10_0(.dout(w_dff_A_1zDzRekS7_0),.din(w_dff_A_h9KHelO10_0),.clk(gclk));
	jdff dff_A_1zDzRekS7_0(.dout(w_dff_A_2y0DEzx67_0),.din(w_dff_A_1zDzRekS7_0),.clk(gclk));
	jdff dff_A_2y0DEzx67_0(.dout(w_dff_A_QShYQLxL0_0),.din(w_dff_A_2y0DEzx67_0),.clk(gclk));
	jdff dff_A_QShYQLxL0_0(.dout(w_dff_A_1pWeIyes3_0),.din(w_dff_A_QShYQLxL0_0),.clk(gclk));
	jdff dff_A_1pWeIyes3_0(.dout(w_dff_A_wBuutEON8_0),.din(w_dff_A_1pWeIyes3_0),.clk(gclk));
	jdff dff_A_wBuutEON8_0(.dout(w_dff_A_LHfcZzWz7_0),.din(w_dff_A_wBuutEON8_0),.clk(gclk));
	jdff dff_A_LHfcZzWz7_0(.dout(w_dff_A_GMAWCa3R2_0),.din(w_dff_A_LHfcZzWz7_0),.clk(gclk));
	jdff dff_A_GMAWCa3R2_0(.dout(w_dff_A_ktH5KyYO5_0),.din(w_dff_A_GMAWCa3R2_0),.clk(gclk));
	jdff dff_A_ktH5KyYO5_0(.dout(w_dff_A_yws4mdaT6_0),.din(w_dff_A_ktH5KyYO5_0),.clk(gclk));
	jdff dff_A_yws4mdaT6_0(.dout(w_dff_A_PulnezTO5_0),.din(w_dff_A_yws4mdaT6_0),.clk(gclk));
	jdff dff_A_PulnezTO5_0(.dout(w_dff_A_m9ajVUs85_0),.din(w_dff_A_PulnezTO5_0),.clk(gclk));
	jdff dff_A_m9ajVUs85_0(.dout(w_dff_A_ic4iOkUk1_0),.din(w_dff_A_m9ajVUs85_0),.clk(gclk));
	jdff dff_A_ic4iOkUk1_0(.dout(w_dff_A_L0Gnt5tY2_0),.din(w_dff_A_ic4iOkUk1_0),.clk(gclk));
	jdff dff_A_L0Gnt5tY2_0(.dout(w_dff_A_Vt3B8Vjt5_0),.din(w_dff_A_L0Gnt5tY2_0),.clk(gclk));
	jdff dff_A_Vt3B8Vjt5_0(.dout(w_dff_A_NE52HxQy2_0),.din(w_dff_A_Vt3B8Vjt5_0),.clk(gclk));
	jdff dff_A_NE52HxQy2_0(.dout(w_dff_A_0CpsxfaY4_0),.din(w_dff_A_NE52HxQy2_0),.clk(gclk));
	jdff dff_A_0CpsxfaY4_0(.dout(w_dff_A_7QVX24J51_0),.din(w_dff_A_0CpsxfaY4_0),.clk(gclk));
	jdff dff_A_7QVX24J51_0(.dout(w_dff_A_zgn1OfDh1_0),.din(w_dff_A_7QVX24J51_0),.clk(gclk));
	jdff dff_A_zgn1OfDh1_0(.dout(w_dff_A_KGSIwgul8_0),.din(w_dff_A_zgn1OfDh1_0),.clk(gclk));
	jdff dff_A_KGSIwgul8_0(.dout(w_dff_A_p7PSgJBZ2_0),.din(w_dff_A_KGSIwgul8_0),.clk(gclk));
	jdff dff_A_p7PSgJBZ2_0(.dout(w_dff_A_yv9LbyyV0_0),.din(w_dff_A_p7PSgJBZ2_0),.clk(gclk));
	jdff dff_A_yv9LbyyV0_0(.dout(w_dff_A_1VLkec4L8_0),.din(w_dff_A_yv9LbyyV0_0),.clk(gclk));
	jdff dff_A_1VLkec4L8_0(.dout(w_dff_A_ZhHCxTWs3_0),.din(w_dff_A_1VLkec4L8_0),.clk(gclk));
	jdff dff_A_ZhHCxTWs3_0(.dout(w_dff_A_hmLEYL4z4_0),.din(w_dff_A_ZhHCxTWs3_0),.clk(gclk));
	jdff dff_A_hmLEYL4z4_0(.dout(w_dff_A_ZfWKkrDK8_0),.din(w_dff_A_hmLEYL4z4_0),.clk(gclk));
	jdff dff_A_ZfWKkrDK8_0(.dout(w_dff_A_r3SQdPc77_0),.din(w_dff_A_ZfWKkrDK8_0),.clk(gclk));
	jdff dff_A_r3SQdPc77_0(.dout(w_dff_A_ORuSLANz5_0),.din(w_dff_A_r3SQdPc77_0),.clk(gclk));
	jdff dff_A_ORuSLANz5_0(.dout(w_dff_A_rFJeUEJU0_0),.din(w_dff_A_ORuSLANz5_0),.clk(gclk));
	jdff dff_A_rFJeUEJU0_0(.dout(w_dff_A_nGz2vt9n0_0),.din(w_dff_A_rFJeUEJU0_0),.clk(gclk));
	jdff dff_A_nGz2vt9n0_0(.dout(w_dff_A_zbZiWfSE7_0),.din(w_dff_A_nGz2vt9n0_0),.clk(gclk));
	jdff dff_A_zbZiWfSE7_0(.dout(w_dff_A_8ux4ot8R9_0),.din(w_dff_A_zbZiWfSE7_0),.clk(gclk));
	jdff dff_A_8ux4ot8R9_0(.dout(w_dff_A_xU0AWXYE5_0),.din(w_dff_A_8ux4ot8R9_0),.clk(gclk));
	jdff dff_A_xU0AWXYE5_0(.dout(w_dff_A_WCdDihVX1_0),.din(w_dff_A_xU0AWXYE5_0),.clk(gclk));
	jdff dff_A_WCdDihVX1_0(.dout(w_dff_A_XDqWUvbp7_0),.din(w_dff_A_WCdDihVX1_0),.clk(gclk));
	jdff dff_A_XDqWUvbp7_0(.dout(w_dff_A_4iZsL2TP3_0),.din(w_dff_A_XDqWUvbp7_0),.clk(gclk));
	jdff dff_A_4iZsL2TP3_0(.dout(w_dff_A_GGLarvz40_0),.din(w_dff_A_4iZsL2TP3_0),.clk(gclk));
	jdff dff_A_GGLarvz40_0(.dout(w_dff_A_ycCWEksQ1_0),.din(w_dff_A_GGLarvz40_0),.clk(gclk));
	jdff dff_A_ycCWEksQ1_0(.dout(w_dff_A_Pe75E43a6_0),.din(w_dff_A_ycCWEksQ1_0),.clk(gclk));
	jdff dff_A_Pe75E43a6_0(.dout(w_dff_A_SNd5FNiI3_0),.din(w_dff_A_Pe75E43a6_0),.clk(gclk));
	jdff dff_A_SNd5FNiI3_0(.dout(w_dff_A_fiMYGD467_0),.din(w_dff_A_SNd5FNiI3_0),.clk(gclk));
	jdff dff_A_fiMYGD467_0(.dout(w_dff_A_ZpZkZq6D0_0),.din(w_dff_A_fiMYGD467_0),.clk(gclk));
	jdff dff_A_ZpZkZq6D0_0(.dout(w_dff_A_Zdi3dTfX2_0),.din(w_dff_A_ZpZkZq6D0_0),.clk(gclk));
	jdff dff_A_Zdi3dTfX2_0(.dout(w_dff_A_mGmPoZMn2_0),.din(w_dff_A_Zdi3dTfX2_0),.clk(gclk));
	jdff dff_A_mGmPoZMn2_0(.dout(w_dff_A_hpHhMutO5_0),.din(w_dff_A_mGmPoZMn2_0),.clk(gclk));
	jdff dff_A_hpHhMutO5_0(.dout(w_dff_A_rZsGNHMR6_0),.din(w_dff_A_hpHhMutO5_0),.clk(gclk));
	jdff dff_A_rZsGNHMR6_0(.dout(w_dff_A_wHLYRihD5_0),.din(w_dff_A_rZsGNHMR6_0),.clk(gclk));
	jdff dff_A_wHLYRihD5_0(.dout(w_dff_A_fQ9m1BRv2_0),.din(w_dff_A_wHLYRihD5_0),.clk(gclk));
	jdff dff_A_fQ9m1BRv2_0(.dout(w_dff_A_582nucf89_0),.din(w_dff_A_fQ9m1BRv2_0),.clk(gclk));
	jdff dff_A_582nucf89_0(.dout(w_dff_A_8lCQdlDI3_0),.din(w_dff_A_582nucf89_0),.clk(gclk));
	jdff dff_A_8lCQdlDI3_0(.dout(w_dff_A_tAdABm3I0_0),.din(w_dff_A_8lCQdlDI3_0),.clk(gclk));
	jdff dff_A_tAdABm3I0_0(.dout(w_dff_A_L9hMv4S83_0),.din(w_dff_A_tAdABm3I0_0),.clk(gclk));
	jdff dff_A_L9hMv4S83_0(.dout(w_dff_A_XL0RG6jC6_0),.din(w_dff_A_L9hMv4S83_0),.clk(gclk));
	jdff dff_A_XL0RG6jC6_0(.dout(w_dff_A_YoNPNwg12_0),.din(w_dff_A_XL0RG6jC6_0),.clk(gclk));
	jdff dff_A_YoNPNwg12_0(.dout(w_dff_A_QswfTllp6_0),.din(w_dff_A_YoNPNwg12_0),.clk(gclk));
	jdff dff_A_QswfTllp6_0(.dout(w_dff_A_QBQbdsmn7_0),.din(w_dff_A_QswfTllp6_0),.clk(gclk));
	jdff dff_A_QBQbdsmn7_0(.dout(w_dff_A_XSgTPFmZ9_0),.din(w_dff_A_QBQbdsmn7_0),.clk(gclk));
	jdff dff_A_XSgTPFmZ9_0(.dout(w_dff_A_oTrKD4mT9_0),.din(w_dff_A_XSgTPFmZ9_0),.clk(gclk));
	jdff dff_A_oTrKD4mT9_0(.dout(w_dff_A_6ntrtNGS0_0),.din(w_dff_A_oTrKD4mT9_0),.clk(gclk));
	jdff dff_A_6ntrtNGS0_0(.dout(w_dff_A_Bt5YQ6nr5_0),.din(w_dff_A_6ntrtNGS0_0),.clk(gclk));
	jdff dff_A_Bt5YQ6nr5_0(.dout(w_dff_A_5UkpyXkc2_0),.din(w_dff_A_Bt5YQ6nr5_0),.clk(gclk));
	jdff dff_A_5UkpyXkc2_0(.dout(w_dff_A_kRMDWBnH1_0),.din(w_dff_A_5UkpyXkc2_0),.clk(gclk));
	jdff dff_A_kRMDWBnH1_0(.dout(w_dff_A_TWfXQ2Sl3_0),.din(w_dff_A_kRMDWBnH1_0),.clk(gclk));
	jdff dff_A_TWfXQ2Sl3_0(.dout(w_dff_A_TfOavHbc7_0),.din(w_dff_A_TWfXQ2Sl3_0),.clk(gclk));
	jdff dff_A_TfOavHbc7_0(.dout(w_dff_A_UPVyrwD12_0),.din(w_dff_A_TfOavHbc7_0),.clk(gclk));
	jdff dff_A_UPVyrwD12_0(.dout(w_dff_A_bSkYozi36_0),.din(w_dff_A_UPVyrwD12_0),.clk(gclk));
	jdff dff_A_bSkYozi36_0(.dout(w_dff_A_Jh2bbCCl4_0),.din(w_dff_A_bSkYozi36_0),.clk(gclk));
	jdff dff_A_Jh2bbCCl4_0(.dout(w_dff_A_LOhNhGVW7_0),.din(w_dff_A_Jh2bbCCl4_0),.clk(gclk));
	jdff dff_A_LOhNhGVW7_0(.dout(w_dff_A_ySUfGGmy5_0),.din(w_dff_A_LOhNhGVW7_0),.clk(gclk));
	jdff dff_A_ySUfGGmy5_0(.dout(w_dff_A_qqT8UNDI9_0),.din(w_dff_A_ySUfGGmy5_0),.clk(gclk));
	jdff dff_A_qqT8UNDI9_0(.dout(w_dff_A_6cVKGCjB0_0),.din(w_dff_A_qqT8UNDI9_0),.clk(gclk));
	jdff dff_A_6cVKGCjB0_0(.dout(w_dff_A_LvN6XhM73_0),.din(w_dff_A_6cVKGCjB0_0),.clk(gclk));
	jdff dff_A_LvN6XhM73_0(.dout(w_dff_A_jQgHP0PG2_0),.din(w_dff_A_LvN6XhM73_0),.clk(gclk));
	jdff dff_A_jQgHP0PG2_0(.dout(w_dff_A_qQcI16md6_0),.din(w_dff_A_jQgHP0PG2_0),.clk(gclk));
	jdff dff_A_qQcI16md6_0(.dout(w_dff_A_3ZXZ8AV16_0),.din(w_dff_A_qQcI16md6_0),.clk(gclk));
	jdff dff_A_3ZXZ8AV16_0(.dout(w_dff_A_ZOzEY6Re4_0),.din(w_dff_A_3ZXZ8AV16_0),.clk(gclk));
	jdff dff_A_ZOzEY6Re4_0(.dout(w_dff_A_LUoCgbM72_0),.din(w_dff_A_ZOzEY6Re4_0),.clk(gclk));
	jdff dff_A_LUoCgbM72_0(.dout(w_dff_A_HvvODXkS3_0),.din(w_dff_A_LUoCgbM72_0),.clk(gclk));
	jdff dff_A_HvvODXkS3_0(.dout(f10),.din(w_dff_A_HvvODXkS3_0),.clk(gclk));
	jdff dff_A_ZrWr9ERl4_2(.dout(w_dff_A_15HcQg9U7_0),.din(w_dff_A_ZrWr9ERl4_2),.clk(gclk));
	jdff dff_A_15HcQg9U7_0(.dout(w_dff_A_UgVoAuRx9_0),.din(w_dff_A_15HcQg9U7_0),.clk(gclk));
	jdff dff_A_UgVoAuRx9_0(.dout(w_dff_A_6bKLCRhg7_0),.din(w_dff_A_UgVoAuRx9_0),.clk(gclk));
	jdff dff_A_6bKLCRhg7_0(.dout(w_dff_A_HnbtIPTM7_0),.din(w_dff_A_6bKLCRhg7_0),.clk(gclk));
	jdff dff_A_HnbtIPTM7_0(.dout(w_dff_A_bNSqxWpw3_0),.din(w_dff_A_HnbtIPTM7_0),.clk(gclk));
	jdff dff_A_bNSqxWpw3_0(.dout(w_dff_A_yZdg2bYG1_0),.din(w_dff_A_bNSqxWpw3_0),.clk(gclk));
	jdff dff_A_yZdg2bYG1_0(.dout(w_dff_A_C7rHcHnE5_0),.din(w_dff_A_yZdg2bYG1_0),.clk(gclk));
	jdff dff_A_C7rHcHnE5_0(.dout(w_dff_A_aBedArzx6_0),.din(w_dff_A_C7rHcHnE5_0),.clk(gclk));
	jdff dff_A_aBedArzx6_0(.dout(w_dff_A_ihv0gZ9z8_0),.din(w_dff_A_aBedArzx6_0),.clk(gclk));
	jdff dff_A_ihv0gZ9z8_0(.dout(w_dff_A_7UajP3OS9_0),.din(w_dff_A_ihv0gZ9z8_0),.clk(gclk));
	jdff dff_A_7UajP3OS9_0(.dout(w_dff_A_ql6x8v0S3_0),.din(w_dff_A_7UajP3OS9_0),.clk(gclk));
	jdff dff_A_ql6x8v0S3_0(.dout(w_dff_A_4NZ6UZoi0_0),.din(w_dff_A_ql6x8v0S3_0),.clk(gclk));
	jdff dff_A_4NZ6UZoi0_0(.dout(w_dff_A_TFI8iHyh5_0),.din(w_dff_A_4NZ6UZoi0_0),.clk(gclk));
	jdff dff_A_TFI8iHyh5_0(.dout(w_dff_A_pXWqM8PU1_0),.din(w_dff_A_TFI8iHyh5_0),.clk(gclk));
	jdff dff_A_pXWqM8PU1_0(.dout(w_dff_A_MP4QBkco0_0),.din(w_dff_A_pXWqM8PU1_0),.clk(gclk));
	jdff dff_A_MP4QBkco0_0(.dout(w_dff_A_2hcH2NAN2_0),.din(w_dff_A_MP4QBkco0_0),.clk(gclk));
	jdff dff_A_2hcH2NAN2_0(.dout(w_dff_A_Zbo3kZsU8_0),.din(w_dff_A_2hcH2NAN2_0),.clk(gclk));
	jdff dff_A_Zbo3kZsU8_0(.dout(w_dff_A_8iylWzLJ3_0),.din(w_dff_A_Zbo3kZsU8_0),.clk(gclk));
	jdff dff_A_8iylWzLJ3_0(.dout(w_dff_A_qiiQj4bI9_0),.din(w_dff_A_8iylWzLJ3_0),.clk(gclk));
	jdff dff_A_qiiQj4bI9_0(.dout(w_dff_A_4F24Tn4b3_0),.din(w_dff_A_qiiQj4bI9_0),.clk(gclk));
	jdff dff_A_4F24Tn4b3_0(.dout(w_dff_A_02mVP7GQ0_0),.din(w_dff_A_4F24Tn4b3_0),.clk(gclk));
	jdff dff_A_02mVP7GQ0_0(.dout(w_dff_A_rTUjMI7x2_0),.din(w_dff_A_02mVP7GQ0_0),.clk(gclk));
	jdff dff_A_rTUjMI7x2_0(.dout(w_dff_A_EyhoHLkS2_0),.din(w_dff_A_rTUjMI7x2_0),.clk(gclk));
	jdff dff_A_EyhoHLkS2_0(.dout(w_dff_A_bpx99x1V6_0),.din(w_dff_A_EyhoHLkS2_0),.clk(gclk));
	jdff dff_A_bpx99x1V6_0(.dout(w_dff_A_7leawFfC3_0),.din(w_dff_A_bpx99x1V6_0),.clk(gclk));
	jdff dff_A_7leawFfC3_0(.dout(w_dff_A_VJA0fGUk6_0),.din(w_dff_A_7leawFfC3_0),.clk(gclk));
	jdff dff_A_VJA0fGUk6_0(.dout(w_dff_A_qJeP7gsc4_0),.din(w_dff_A_VJA0fGUk6_0),.clk(gclk));
	jdff dff_A_qJeP7gsc4_0(.dout(w_dff_A_9JithcuB7_0),.din(w_dff_A_qJeP7gsc4_0),.clk(gclk));
	jdff dff_A_9JithcuB7_0(.dout(w_dff_A_Xprvgxjm3_0),.din(w_dff_A_9JithcuB7_0),.clk(gclk));
	jdff dff_A_Xprvgxjm3_0(.dout(w_dff_A_YiEK16rm4_0),.din(w_dff_A_Xprvgxjm3_0),.clk(gclk));
	jdff dff_A_YiEK16rm4_0(.dout(w_dff_A_fYv0izgo3_0),.din(w_dff_A_YiEK16rm4_0),.clk(gclk));
	jdff dff_A_fYv0izgo3_0(.dout(w_dff_A_3dcNZQKF6_0),.din(w_dff_A_fYv0izgo3_0),.clk(gclk));
	jdff dff_A_3dcNZQKF6_0(.dout(w_dff_A_yEf3t1Fx3_0),.din(w_dff_A_3dcNZQKF6_0),.clk(gclk));
	jdff dff_A_yEf3t1Fx3_0(.dout(w_dff_A_hOFFA0jj0_0),.din(w_dff_A_yEf3t1Fx3_0),.clk(gclk));
	jdff dff_A_hOFFA0jj0_0(.dout(w_dff_A_fBuzkhkP4_0),.din(w_dff_A_hOFFA0jj0_0),.clk(gclk));
	jdff dff_A_fBuzkhkP4_0(.dout(w_dff_A_5iiAkiTO5_0),.din(w_dff_A_fBuzkhkP4_0),.clk(gclk));
	jdff dff_A_5iiAkiTO5_0(.dout(w_dff_A_W9OkXWNG4_0),.din(w_dff_A_5iiAkiTO5_0),.clk(gclk));
	jdff dff_A_W9OkXWNG4_0(.dout(w_dff_A_kHYDAXqZ8_0),.din(w_dff_A_W9OkXWNG4_0),.clk(gclk));
	jdff dff_A_kHYDAXqZ8_0(.dout(w_dff_A_gbD6eOfb5_0),.din(w_dff_A_kHYDAXqZ8_0),.clk(gclk));
	jdff dff_A_gbD6eOfb5_0(.dout(w_dff_A_YOzaICmi4_0),.din(w_dff_A_gbD6eOfb5_0),.clk(gclk));
	jdff dff_A_YOzaICmi4_0(.dout(w_dff_A_vpE0DHAH5_0),.din(w_dff_A_YOzaICmi4_0),.clk(gclk));
	jdff dff_A_vpE0DHAH5_0(.dout(w_dff_A_wS7BklKo3_0),.din(w_dff_A_vpE0DHAH5_0),.clk(gclk));
	jdff dff_A_wS7BklKo3_0(.dout(w_dff_A_jzKdHl3s1_0),.din(w_dff_A_wS7BklKo3_0),.clk(gclk));
	jdff dff_A_jzKdHl3s1_0(.dout(w_dff_A_epCTTsWm8_0),.din(w_dff_A_jzKdHl3s1_0),.clk(gclk));
	jdff dff_A_epCTTsWm8_0(.dout(w_dff_A_9HpT1eWw8_0),.din(w_dff_A_epCTTsWm8_0),.clk(gclk));
	jdff dff_A_9HpT1eWw8_0(.dout(w_dff_A_nCzWPstu1_0),.din(w_dff_A_9HpT1eWw8_0),.clk(gclk));
	jdff dff_A_nCzWPstu1_0(.dout(w_dff_A_SUSXpkHA8_0),.din(w_dff_A_nCzWPstu1_0),.clk(gclk));
	jdff dff_A_SUSXpkHA8_0(.dout(w_dff_A_0VmBQBJr8_0),.din(w_dff_A_SUSXpkHA8_0),.clk(gclk));
	jdff dff_A_0VmBQBJr8_0(.dout(w_dff_A_bFYvkhAP3_0),.din(w_dff_A_0VmBQBJr8_0),.clk(gclk));
	jdff dff_A_bFYvkhAP3_0(.dout(w_dff_A_IxllTX1D4_0),.din(w_dff_A_bFYvkhAP3_0),.clk(gclk));
	jdff dff_A_IxllTX1D4_0(.dout(w_dff_A_ePPRqBus1_0),.din(w_dff_A_IxllTX1D4_0),.clk(gclk));
	jdff dff_A_ePPRqBus1_0(.dout(w_dff_A_fb60NbWI2_0),.din(w_dff_A_ePPRqBus1_0),.clk(gclk));
	jdff dff_A_fb60NbWI2_0(.dout(w_dff_A_pSZQOTxJ4_0),.din(w_dff_A_fb60NbWI2_0),.clk(gclk));
	jdff dff_A_pSZQOTxJ4_0(.dout(w_dff_A_dC2NcBKJ1_0),.din(w_dff_A_pSZQOTxJ4_0),.clk(gclk));
	jdff dff_A_dC2NcBKJ1_0(.dout(w_dff_A_JrCTLoXY6_0),.din(w_dff_A_dC2NcBKJ1_0),.clk(gclk));
	jdff dff_A_JrCTLoXY6_0(.dout(w_dff_A_SkJD0Apt5_0),.din(w_dff_A_JrCTLoXY6_0),.clk(gclk));
	jdff dff_A_SkJD0Apt5_0(.dout(w_dff_A_yIkeT2ln9_0),.din(w_dff_A_SkJD0Apt5_0),.clk(gclk));
	jdff dff_A_yIkeT2ln9_0(.dout(w_dff_A_S6bOPlNl4_0),.din(w_dff_A_yIkeT2ln9_0),.clk(gclk));
	jdff dff_A_S6bOPlNl4_0(.dout(w_dff_A_axCSck3S7_0),.din(w_dff_A_S6bOPlNl4_0),.clk(gclk));
	jdff dff_A_axCSck3S7_0(.dout(w_dff_A_cK4FlwEo1_0),.din(w_dff_A_axCSck3S7_0),.clk(gclk));
	jdff dff_A_cK4FlwEo1_0(.dout(w_dff_A_wUOK7QKQ4_0),.din(w_dff_A_cK4FlwEo1_0),.clk(gclk));
	jdff dff_A_wUOK7QKQ4_0(.dout(w_dff_A_10TaH3VO1_0),.din(w_dff_A_wUOK7QKQ4_0),.clk(gclk));
	jdff dff_A_10TaH3VO1_0(.dout(w_dff_A_J2CPWDlv9_0),.din(w_dff_A_10TaH3VO1_0),.clk(gclk));
	jdff dff_A_J2CPWDlv9_0(.dout(w_dff_A_hpt6nDx61_0),.din(w_dff_A_J2CPWDlv9_0),.clk(gclk));
	jdff dff_A_hpt6nDx61_0(.dout(w_dff_A_unztLCtB1_0),.din(w_dff_A_hpt6nDx61_0),.clk(gclk));
	jdff dff_A_unztLCtB1_0(.dout(w_dff_A_1zCq4sQO2_0),.din(w_dff_A_unztLCtB1_0),.clk(gclk));
	jdff dff_A_1zCq4sQO2_0(.dout(w_dff_A_dFoNTzyt0_0),.din(w_dff_A_1zCq4sQO2_0),.clk(gclk));
	jdff dff_A_dFoNTzyt0_0(.dout(w_dff_A_1bn6RTcI0_0),.din(w_dff_A_dFoNTzyt0_0),.clk(gclk));
	jdff dff_A_1bn6RTcI0_0(.dout(w_dff_A_fE1ekTHR0_0),.din(w_dff_A_1bn6RTcI0_0),.clk(gclk));
	jdff dff_A_fE1ekTHR0_0(.dout(w_dff_A_6wjvUxBG5_0),.din(w_dff_A_fE1ekTHR0_0),.clk(gclk));
	jdff dff_A_6wjvUxBG5_0(.dout(w_dff_A_tsagRu9B4_0),.din(w_dff_A_6wjvUxBG5_0),.clk(gclk));
	jdff dff_A_tsagRu9B4_0(.dout(w_dff_A_nbLw0WLj6_0),.din(w_dff_A_tsagRu9B4_0),.clk(gclk));
	jdff dff_A_nbLw0WLj6_0(.dout(w_dff_A_qVOIaLGz1_0),.din(w_dff_A_nbLw0WLj6_0),.clk(gclk));
	jdff dff_A_qVOIaLGz1_0(.dout(w_dff_A_pQj4XA6F6_0),.din(w_dff_A_qVOIaLGz1_0),.clk(gclk));
	jdff dff_A_pQj4XA6F6_0(.dout(w_dff_A_lenHzLJi4_0),.din(w_dff_A_pQj4XA6F6_0),.clk(gclk));
	jdff dff_A_lenHzLJi4_0(.dout(w_dff_A_eEBgcmwB1_0),.din(w_dff_A_lenHzLJi4_0),.clk(gclk));
	jdff dff_A_eEBgcmwB1_0(.dout(w_dff_A_dNFtxpV62_0),.din(w_dff_A_eEBgcmwB1_0),.clk(gclk));
	jdff dff_A_dNFtxpV62_0(.dout(w_dff_A_EZCKI5Vp6_0),.din(w_dff_A_dNFtxpV62_0),.clk(gclk));
	jdff dff_A_EZCKI5Vp6_0(.dout(w_dff_A_TlBzjPzF9_0),.din(w_dff_A_EZCKI5Vp6_0),.clk(gclk));
	jdff dff_A_TlBzjPzF9_0(.dout(w_dff_A_DZcnUb4g1_0),.din(w_dff_A_TlBzjPzF9_0),.clk(gclk));
	jdff dff_A_DZcnUb4g1_0(.dout(w_dff_A_5T5pFwlh1_0),.din(w_dff_A_DZcnUb4g1_0),.clk(gclk));
	jdff dff_A_5T5pFwlh1_0(.dout(w_dff_A_pNhYQ22y8_0),.din(w_dff_A_5T5pFwlh1_0),.clk(gclk));
	jdff dff_A_pNhYQ22y8_0(.dout(w_dff_A_rr4vJImw4_0),.din(w_dff_A_pNhYQ22y8_0),.clk(gclk));
	jdff dff_A_rr4vJImw4_0(.dout(w_dff_A_rfMzGpFH8_0),.din(w_dff_A_rr4vJImw4_0),.clk(gclk));
	jdff dff_A_rfMzGpFH8_0(.dout(w_dff_A_RblJ08sR7_0),.din(w_dff_A_rfMzGpFH8_0),.clk(gclk));
	jdff dff_A_RblJ08sR7_0(.dout(w_dff_A_eRWA5Weh2_0),.din(w_dff_A_RblJ08sR7_0),.clk(gclk));
	jdff dff_A_eRWA5Weh2_0(.dout(w_dff_A_bUCnsmSF5_0),.din(w_dff_A_eRWA5Weh2_0),.clk(gclk));
	jdff dff_A_bUCnsmSF5_0(.dout(w_dff_A_3G2OhcFT1_0),.din(w_dff_A_bUCnsmSF5_0),.clk(gclk));
	jdff dff_A_3G2OhcFT1_0(.dout(w_dff_A_ZbdzZVdS4_0),.din(w_dff_A_3G2OhcFT1_0),.clk(gclk));
	jdff dff_A_ZbdzZVdS4_0(.dout(w_dff_A_k3DCA6SB9_0),.din(w_dff_A_ZbdzZVdS4_0),.clk(gclk));
	jdff dff_A_k3DCA6SB9_0(.dout(w_dff_A_ET9lZcgD0_0),.din(w_dff_A_k3DCA6SB9_0),.clk(gclk));
	jdff dff_A_ET9lZcgD0_0(.dout(w_dff_A_OQNcGgK65_0),.din(w_dff_A_ET9lZcgD0_0),.clk(gclk));
	jdff dff_A_OQNcGgK65_0(.dout(w_dff_A_QG532PEa1_0),.din(w_dff_A_OQNcGgK65_0),.clk(gclk));
	jdff dff_A_QG532PEa1_0(.dout(w_dff_A_XNzX6bgo5_0),.din(w_dff_A_QG532PEa1_0),.clk(gclk));
	jdff dff_A_XNzX6bgo5_0(.dout(w_dff_A_7ZavvGFy8_0),.din(w_dff_A_XNzX6bgo5_0),.clk(gclk));
	jdff dff_A_7ZavvGFy8_0(.dout(w_dff_A_jltbk1ix3_0),.din(w_dff_A_7ZavvGFy8_0),.clk(gclk));
	jdff dff_A_jltbk1ix3_0(.dout(w_dff_A_o3bY3S3Y3_0),.din(w_dff_A_jltbk1ix3_0),.clk(gclk));
	jdff dff_A_o3bY3S3Y3_0(.dout(w_dff_A_H0hyyIro3_0),.din(w_dff_A_o3bY3S3Y3_0),.clk(gclk));
	jdff dff_A_H0hyyIro3_0(.dout(w_dff_A_uoAR7BSt3_0),.din(w_dff_A_H0hyyIro3_0),.clk(gclk));
	jdff dff_A_uoAR7BSt3_0(.dout(w_dff_A_ZIn0HoNO2_0),.din(w_dff_A_uoAR7BSt3_0),.clk(gclk));
	jdff dff_A_ZIn0HoNO2_0(.dout(w_dff_A_B9WWfpk30_0),.din(w_dff_A_ZIn0HoNO2_0),.clk(gclk));
	jdff dff_A_B9WWfpk30_0(.dout(w_dff_A_FO6D9ciQ6_0),.din(w_dff_A_B9WWfpk30_0),.clk(gclk));
	jdff dff_A_FO6D9ciQ6_0(.dout(w_dff_A_b3l3KliC4_0),.din(w_dff_A_FO6D9ciQ6_0),.clk(gclk));
	jdff dff_A_b3l3KliC4_0(.dout(w_dff_A_UYf7O8Tk2_0),.din(w_dff_A_b3l3KliC4_0),.clk(gclk));
	jdff dff_A_UYf7O8Tk2_0(.dout(w_dff_A_7aOcJt900_0),.din(w_dff_A_UYf7O8Tk2_0),.clk(gclk));
	jdff dff_A_7aOcJt900_0(.dout(w_dff_A_6bqglOVK8_0),.din(w_dff_A_7aOcJt900_0),.clk(gclk));
	jdff dff_A_6bqglOVK8_0(.dout(w_dff_A_AHXZk2rw1_0),.din(w_dff_A_6bqglOVK8_0),.clk(gclk));
	jdff dff_A_AHXZk2rw1_0(.dout(w_dff_A_dKkO9qPk8_0),.din(w_dff_A_AHXZk2rw1_0),.clk(gclk));
	jdff dff_A_dKkO9qPk8_0(.dout(w_dff_A_ZQNDci8i0_0),.din(w_dff_A_dKkO9qPk8_0),.clk(gclk));
	jdff dff_A_ZQNDci8i0_0(.dout(w_dff_A_oN8lrO2u9_0),.din(w_dff_A_ZQNDci8i0_0),.clk(gclk));
	jdff dff_A_oN8lrO2u9_0(.dout(w_dff_A_B0zb1x6Q7_0),.din(w_dff_A_oN8lrO2u9_0),.clk(gclk));
	jdff dff_A_B0zb1x6Q7_0(.dout(w_dff_A_PivgCzWd9_0),.din(w_dff_A_B0zb1x6Q7_0),.clk(gclk));
	jdff dff_A_PivgCzWd9_0(.dout(w_dff_A_QE7SKFjN1_0),.din(w_dff_A_PivgCzWd9_0),.clk(gclk));
	jdff dff_A_QE7SKFjN1_0(.dout(w_dff_A_ZFs8B1zb2_0),.din(w_dff_A_QE7SKFjN1_0),.clk(gclk));
	jdff dff_A_ZFs8B1zb2_0(.dout(w_dff_A_5DUOrROx7_0),.din(w_dff_A_ZFs8B1zb2_0),.clk(gclk));
	jdff dff_A_5DUOrROx7_0(.dout(f11),.din(w_dff_A_5DUOrROx7_0),.clk(gclk));
	jdff dff_A_fR6FTcm21_2(.dout(w_dff_A_y7WhSNYQ7_0),.din(w_dff_A_fR6FTcm21_2),.clk(gclk));
	jdff dff_A_y7WhSNYQ7_0(.dout(w_dff_A_6z1nnNHl4_0),.din(w_dff_A_y7WhSNYQ7_0),.clk(gclk));
	jdff dff_A_6z1nnNHl4_0(.dout(w_dff_A_XaOXOBOL0_0),.din(w_dff_A_6z1nnNHl4_0),.clk(gclk));
	jdff dff_A_XaOXOBOL0_0(.dout(w_dff_A_fodcdQKs6_0),.din(w_dff_A_XaOXOBOL0_0),.clk(gclk));
	jdff dff_A_fodcdQKs6_0(.dout(w_dff_A_7BXV6UXY4_0),.din(w_dff_A_fodcdQKs6_0),.clk(gclk));
	jdff dff_A_7BXV6UXY4_0(.dout(w_dff_A_tm0QLkmT1_0),.din(w_dff_A_7BXV6UXY4_0),.clk(gclk));
	jdff dff_A_tm0QLkmT1_0(.dout(w_dff_A_fZ3G0fIF0_0),.din(w_dff_A_tm0QLkmT1_0),.clk(gclk));
	jdff dff_A_fZ3G0fIF0_0(.dout(w_dff_A_sihbW0vt7_0),.din(w_dff_A_fZ3G0fIF0_0),.clk(gclk));
	jdff dff_A_sihbW0vt7_0(.dout(w_dff_A_SVDLCNvx2_0),.din(w_dff_A_sihbW0vt7_0),.clk(gclk));
	jdff dff_A_SVDLCNvx2_0(.dout(w_dff_A_6wDwT20S0_0),.din(w_dff_A_SVDLCNvx2_0),.clk(gclk));
	jdff dff_A_6wDwT20S0_0(.dout(w_dff_A_bmPmeZCt2_0),.din(w_dff_A_6wDwT20S0_0),.clk(gclk));
	jdff dff_A_bmPmeZCt2_0(.dout(w_dff_A_7RF50jCU8_0),.din(w_dff_A_bmPmeZCt2_0),.clk(gclk));
	jdff dff_A_7RF50jCU8_0(.dout(w_dff_A_zAJRgU9d4_0),.din(w_dff_A_7RF50jCU8_0),.clk(gclk));
	jdff dff_A_zAJRgU9d4_0(.dout(w_dff_A_3ToLIOZR1_0),.din(w_dff_A_zAJRgU9d4_0),.clk(gclk));
	jdff dff_A_3ToLIOZR1_0(.dout(w_dff_A_ikKcsmME0_0),.din(w_dff_A_3ToLIOZR1_0),.clk(gclk));
	jdff dff_A_ikKcsmME0_0(.dout(w_dff_A_I3KAtPI58_0),.din(w_dff_A_ikKcsmME0_0),.clk(gclk));
	jdff dff_A_I3KAtPI58_0(.dout(w_dff_A_LCDkvxGM6_0),.din(w_dff_A_I3KAtPI58_0),.clk(gclk));
	jdff dff_A_LCDkvxGM6_0(.dout(w_dff_A_WzzIVol07_0),.din(w_dff_A_LCDkvxGM6_0),.clk(gclk));
	jdff dff_A_WzzIVol07_0(.dout(w_dff_A_IaCWVXSM4_0),.din(w_dff_A_WzzIVol07_0),.clk(gclk));
	jdff dff_A_IaCWVXSM4_0(.dout(w_dff_A_nP8h33mC4_0),.din(w_dff_A_IaCWVXSM4_0),.clk(gclk));
	jdff dff_A_nP8h33mC4_0(.dout(w_dff_A_trIiBRfK7_0),.din(w_dff_A_nP8h33mC4_0),.clk(gclk));
	jdff dff_A_trIiBRfK7_0(.dout(w_dff_A_FbYro3jv7_0),.din(w_dff_A_trIiBRfK7_0),.clk(gclk));
	jdff dff_A_FbYro3jv7_0(.dout(w_dff_A_TS5kjr0u8_0),.din(w_dff_A_FbYro3jv7_0),.clk(gclk));
	jdff dff_A_TS5kjr0u8_0(.dout(w_dff_A_2jmUOqW10_0),.din(w_dff_A_TS5kjr0u8_0),.clk(gclk));
	jdff dff_A_2jmUOqW10_0(.dout(w_dff_A_IYyeKXR31_0),.din(w_dff_A_2jmUOqW10_0),.clk(gclk));
	jdff dff_A_IYyeKXR31_0(.dout(w_dff_A_lqPIHeOr2_0),.din(w_dff_A_IYyeKXR31_0),.clk(gclk));
	jdff dff_A_lqPIHeOr2_0(.dout(w_dff_A_AwcBvLbG3_0),.din(w_dff_A_lqPIHeOr2_0),.clk(gclk));
	jdff dff_A_AwcBvLbG3_0(.dout(w_dff_A_5w7Gfoom7_0),.din(w_dff_A_AwcBvLbG3_0),.clk(gclk));
	jdff dff_A_5w7Gfoom7_0(.dout(w_dff_A_GZnb6yT07_0),.din(w_dff_A_5w7Gfoom7_0),.clk(gclk));
	jdff dff_A_GZnb6yT07_0(.dout(w_dff_A_U3YbTNFS4_0),.din(w_dff_A_GZnb6yT07_0),.clk(gclk));
	jdff dff_A_U3YbTNFS4_0(.dout(w_dff_A_8j1E2ceg7_0),.din(w_dff_A_U3YbTNFS4_0),.clk(gclk));
	jdff dff_A_8j1E2ceg7_0(.dout(w_dff_A_SbMbh9sX0_0),.din(w_dff_A_8j1E2ceg7_0),.clk(gclk));
	jdff dff_A_SbMbh9sX0_0(.dout(w_dff_A_dnfJeEbh7_0),.din(w_dff_A_SbMbh9sX0_0),.clk(gclk));
	jdff dff_A_dnfJeEbh7_0(.dout(w_dff_A_dvvq5irm7_0),.din(w_dff_A_dnfJeEbh7_0),.clk(gclk));
	jdff dff_A_dvvq5irm7_0(.dout(w_dff_A_iGp2IYsb1_0),.din(w_dff_A_dvvq5irm7_0),.clk(gclk));
	jdff dff_A_iGp2IYsb1_0(.dout(w_dff_A_584jK6gU6_0),.din(w_dff_A_iGp2IYsb1_0),.clk(gclk));
	jdff dff_A_584jK6gU6_0(.dout(w_dff_A_iaokvyBS5_0),.din(w_dff_A_584jK6gU6_0),.clk(gclk));
	jdff dff_A_iaokvyBS5_0(.dout(w_dff_A_B2cji4F71_0),.din(w_dff_A_iaokvyBS5_0),.clk(gclk));
	jdff dff_A_B2cji4F71_0(.dout(w_dff_A_IHyt1oMD4_0),.din(w_dff_A_B2cji4F71_0),.clk(gclk));
	jdff dff_A_IHyt1oMD4_0(.dout(w_dff_A_kllMZS7q3_0),.din(w_dff_A_IHyt1oMD4_0),.clk(gclk));
	jdff dff_A_kllMZS7q3_0(.dout(w_dff_A_NJSNWmYt1_0),.din(w_dff_A_kllMZS7q3_0),.clk(gclk));
	jdff dff_A_NJSNWmYt1_0(.dout(w_dff_A_9n9jj4344_0),.din(w_dff_A_NJSNWmYt1_0),.clk(gclk));
	jdff dff_A_9n9jj4344_0(.dout(w_dff_A_FoO0ayB03_0),.din(w_dff_A_9n9jj4344_0),.clk(gclk));
	jdff dff_A_FoO0ayB03_0(.dout(w_dff_A_j6Ts3P5a0_0),.din(w_dff_A_FoO0ayB03_0),.clk(gclk));
	jdff dff_A_j6Ts3P5a0_0(.dout(w_dff_A_P99ZzB4Y7_0),.din(w_dff_A_j6Ts3P5a0_0),.clk(gclk));
	jdff dff_A_P99ZzB4Y7_0(.dout(w_dff_A_75W9U8704_0),.din(w_dff_A_P99ZzB4Y7_0),.clk(gclk));
	jdff dff_A_75W9U8704_0(.dout(w_dff_A_c1z5pt989_0),.din(w_dff_A_75W9U8704_0),.clk(gclk));
	jdff dff_A_c1z5pt989_0(.dout(w_dff_A_PPjWTK8L3_0),.din(w_dff_A_c1z5pt989_0),.clk(gclk));
	jdff dff_A_PPjWTK8L3_0(.dout(w_dff_A_6SzfAzzR1_0),.din(w_dff_A_PPjWTK8L3_0),.clk(gclk));
	jdff dff_A_6SzfAzzR1_0(.dout(w_dff_A_sWS2HhKH6_0),.din(w_dff_A_6SzfAzzR1_0),.clk(gclk));
	jdff dff_A_sWS2HhKH6_0(.dout(w_dff_A_tRTxfeMJ1_0),.din(w_dff_A_sWS2HhKH6_0),.clk(gclk));
	jdff dff_A_tRTxfeMJ1_0(.dout(w_dff_A_BxW6PY2o8_0),.din(w_dff_A_tRTxfeMJ1_0),.clk(gclk));
	jdff dff_A_BxW6PY2o8_0(.dout(w_dff_A_EHoXfIBY4_0),.din(w_dff_A_BxW6PY2o8_0),.clk(gclk));
	jdff dff_A_EHoXfIBY4_0(.dout(w_dff_A_1J4FoOdO4_0),.din(w_dff_A_EHoXfIBY4_0),.clk(gclk));
	jdff dff_A_1J4FoOdO4_0(.dout(w_dff_A_gAqIS2lD5_0),.din(w_dff_A_1J4FoOdO4_0),.clk(gclk));
	jdff dff_A_gAqIS2lD5_0(.dout(w_dff_A_xCvvQE6d4_0),.din(w_dff_A_gAqIS2lD5_0),.clk(gclk));
	jdff dff_A_xCvvQE6d4_0(.dout(w_dff_A_R8kdQ0IK5_0),.din(w_dff_A_xCvvQE6d4_0),.clk(gclk));
	jdff dff_A_R8kdQ0IK5_0(.dout(w_dff_A_lTAphZi96_0),.din(w_dff_A_R8kdQ0IK5_0),.clk(gclk));
	jdff dff_A_lTAphZi96_0(.dout(w_dff_A_5Swu2wGt3_0),.din(w_dff_A_lTAphZi96_0),.clk(gclk));
	jdff dff_A_5Swu2wGt3_0(.dout(w_dff_A_OlcjcwmA3_0),.din(w_dff_A_5Swu2wGt3_0),.clk(gclk));
	jdff dff_A_OlcjcwmA3_0(.dout(w_dff_A_LNM75Euf6_0),.din(w_dff_A_OlcjcwmA3_0),.clk(gclk));
	jdff dff_A_LNM75Euf6_0(.dout(w_dff_A_cPrvOmTY3_0),.din(w_dff_A_LNM75Euf6_0),.clk(gclk));
	jdff dff_A_cPrvOmTY3_0(.dout(w_dff_A_058Cf25e8_0),.din(w_dff_A_cPrvOmTY3_0),.clk(gclk));
	jdff dff_A_058Cf25e8_0(.dout(w_dff_A_KDS1bbSl9_0),.din(w_dff_A_058Cf25e8_0),.clk(gclk));
	jdff dff_A_KDS1bbSl9_0(.dout(w_dff_A_YNJYXBCF9_0),.din(w_dff_A_KDS1bbSl9_0),.clk(gclk));
	jdff dff_A_YNJYXBCF9_0(.dout(w_dff_A_xleCjhWi7_0),.din(w_dff_A_YNJYXBCF9_0),.clk(gclk));
	jdff dff_A_xleCjhWi7_0(.dout(w_dff_A_rq4jptBu8_0),.din(w_dff_A_xleCjhWi7_0),.clk(gclk));
	jdff dff_A_rq4jptBu8_0(.dout(w_dff_A_UaFuHvic3_0),.din(w_dff_A_rq4jptBu8_0),.clk(gclk));
	jdff dff_A_UaFuHvic3_0(.dout(w_dff_A_9QAQU2qe9_0),.din(w_dff_A_UaFuHvic3_0),.clk(gclk));
	jdff dff_A_9QAQU2qe9_0(.dout(w_dff_A_Y4dGORsR3_0),.din(w_dff_A_9QAQU2qe9_0),.clk(gclk));
	jdff dff_A_Y4dGORsR3_0(.dout(w_dff_A_aY0ry2Gg2_0),.din(w_dff_A_Y4dGORsR3_0),.clk(gclk));
	jdff dff_A_aY0ry2Gg2_0(.dout(w_dff_A_ldrmDmAz6_0),.din(w_dff_A_aY0ry2Gg2_0),.clk(gclk));
	jdff dff_A_ldrmDmAz6_0(.dout(w_dff_A_4ql2nkjp8_0),.din(w_dff_A_ldrmDmAz6_0),.clk(gclk));
	jdff dff_A_4ql2nkjp8_0(.dout(w_dff_A_Iht7PWfw9_0),.din(w_dff_A_4ql2nkjp8_0),.clk(gclk));
	jdff dff_A_Iht7PWfw9_0(.dout(w_dff_A_5LtbLBHI5_0),.din(w_dff_A_Iht7PWfw9_0),.clk(gclk));
	jdff dff_A_5LtbLBHI5_0(.dout(w_dff_A_UUERqg471_0),.din(w_dff_A_5LtbLBHI5_0),.clk(gclk));
	jdff dff_A_UUERqg471_0(.dout(w_dff_A_iKFmuGJR0_0),.din(w_dff_A_UUERqg471_0),.clk(gclk));
	jdff dff_A_iKFmuGJR0_0(.dout(w_dff_A_GdrE35gt8_0),.din(w_dff_A_iKFmuGJR0_0),.clk(gclk));
	jdff dff_A_GdrE35gt8_0(.dout(w_dff_A_pJSrhPX42_0),.din(w_dff_A_GdrE35gt8_0),.clk(gclk));
	jdff dff_A_pJSrhPX42_0(.dout(w_dff_A_3h1DO1Y98_0),.din(w_dff_A_pJSrhPX42_0),.clk(gclk));
	jdff dff_A_3h1DO1Y98_0(.dout(w_dff_A_kB1qCdO48_0),.din(w_dff_A_3h1DO1Y98_0),.clk(gclk));
	jdff dff_A_kB1qCdO48_0(.dout(w_dff_A_tciRGW9O9_0),.din(w_dff_A_kB1qCdO48_0),.clk(gclk));
	jdff dff_A_tciRGW9O9_0(.dout(w_dff_A_1IZjxcza9_0),.din(w_dff_A_tciRGW9O9_0),.clk(gclk));
	jdff dff_A_1IZjxcza9_0(.dout(w_dff_A_EelNvNHN2_0),.din(w_dff_A_1IZjxcza9_0),.clk(gclk));
	jdff dff_A_EelNvNHN2_0(.dout(w_dff_A_tRxX3MST2_0),.din(w_dff_A_EelNvNHN2_0),.clk(gclk));
	jdff dff_A_tRxX3MST2_0(.dout(w_dff_A_NjMjIRqf6_0),.din(w_dff_A_tRxX3MST2_0),.clk(gclk));
	jdff dff_A_NjMjIRqf6_0(.dout(w_dff_A_MSuLK1OP9_0),.din(w_dff_A_NjMjIRqf6_0),.clk(gclk));
	jdff dff_A_MSuLK1OP9_0(.dout(w_dff_A_7MM59aGF9_0),.din(w_dff_A_MSuLK1OP9_0),.clk(gclk));
	jdff dff_A_7MM59aGF9_0(.dout(w_dff_A_X3Qqwu5C6_0),.din(w_dff_A_7MM59aGF9_0),.clk(gclk));
	jdff dff_A_X3Qqwu5C6_0(.dout(w_dff_A_epdSzUUA3_0),.din(w_dff_A_X3Qqwu5C6_0),.clk(gclk));
	jdff dff_A_epdSzUUA3_0(.dout(w_dff_A_UKxYtE504_0),.din(w_dff_A_epdSzUUA3_0),.clk(gclk));
	jdff dff_A_UKxYtE504_0(.dout(w_dff_A_G6vb3wgD2_0),.din(w_dff_A_UKxYtE504_0),.clk(gclk));
	jdff dff_A_G6vb3wgD2_0(.dout(w_dff_A_jvt5CBJk3_0),.din(w_dff_A_G6vb3wgD2_0),.clk(gclk));
	jdff dff_A_jvt5CBJk3_0(.dout(w_dff_A_cqwQ3lgT8_0),.din(w_dff_A_jvt5CBJk3_0),.clk(gclk));
	jdff dff_A_cqwQ3lgT8_0(.dout(w_dff_A_PWeN0vfI1_0),.din(w_dff_A_cqwQ3lgT8_0),.clk(gclk));
	jdff dff_A_PWeN0vfI1_0(.dout(w_dff_A_30WlPK1O7_0),.din(w_dff_A_PWeN0vfI1_0),.clk(gclk));
	jdff dff_A_30WlPK1O7_0(.dout(w_dff_A_KjMxXW2Z7_0),.din(w_dff_A_30WlPK1O7_0),.clk(gclk));
	jdff dff_A_KjMxXW2Z7_0(.dout(w_dff_A_rWHmgSme1_0),.din(w_dff_A_KjMxXW2Z7_0),.clk(gclk));
	jdff dff_A_rWHmgSme1_0(.dout(w_dff_A_GKLPcDGC0_0),.din(w_dff_A_rWHmgSme1_0),.clk(gclk));
	jdff dff_A_GKLPcDGC0_0(.dout(w_dff_A_I863mCVa7_0),.din(w_dff_A_GKLPcDGC0_0),.clk(gclk));
	jdff dff_A_I863mCVa7_0(.dout(w_dff_A_na5gntbZ1_0),.din(w_dff_A_I863mCVa7_0),.clk(gclk));
	jdff dff_A_na5gntbZ1_0(.dout(w_dff_A_yD6dehP53_0),.din(w_dff_A_na5gntbZ1_0),.clk(gclk));
	jdff dff_A_yD6dehP53_0(.dout(w_dff_A_HNdbQz9a0_0),.din(w_dff_A_yD6dehP53_0),.clk(gclk));
	jdff dff_A_HNdbQz9a0_0(.dout(w_dff_A_JgLAJzPS0_0),.din(w_dff_A_HNdbQz9a0_0),.clk(gclk));
	jdff dff_A_JgLAJzPS0_0(.dout(w_dff_A_HT3oSSMJ1_0),.din(w_dff_A_JgLAJzPS0_0),.clk(gclk));
	jdff dff_A_HT3oSSMJ1_0(.dout(w_dff_A_HT34WWlX5_0),.din(w_dff_A_HT3oSSMJ1_0),.clk(gclk));
	jdff dff_A_HT34WWlX5_0(.dout(w_dff_A_cBHBIEwD0_0),.din(w_dff_A_HT34WWlX5_0),.clk(gclk));
	jdff dff_A_cBHBIEwD0_0(.dout(w_dff_A_hZAJBVeo9_0),.din(w_dff_A_cBHBIEwD0_0),.clk(gclk));
	jdff dff_A_hZAJBVeo9_0(.dout(w_dff_A_9HjBetnd0_0),.din(w_dff_A_hZAJBVeo9_0),.clk(gclk));
	jdff dff_A_9HjBetnd0_0(.dout(w_dff_A_oATdPfMO9_0),.din(w_dff_A_9HjBetnd0_0),.clk(gclk));
	jdff dff_A_oATdPfMO9_0(.dout(w_dff_A_VuFtPo5K3_0),.din(w_dff_A_oATdPfMO9_0),.clk(gclk));
	jdff dff_A_VuFtPo5K3_0(.dout(w_dff_A_dGceOg5Q2_0),.din(w_dff_A_VuFtPo5K3_0),.clk(gclk));
	jdff dff_A_dGceOg5Q2_0(.dout(w_dff_A_rI8AILxN3_0),.din(w_dff_A_dGceOg5Q2_0),.clk(gclk));
	jdff dff_A_rI8AILxN3_0(.dout(w_dff_A_LMG2NbA00_0),.din(w_dff_A_rI8AILxN3_0),.clk(gclk));
	jdff dff_A_LMG2NbA00_0(.dout(f12),.din(w_dff_A_LMG2NbA00_0),.clk(gclk));
	jdff dff_A_4btOcuhR0_2(.dout(w_dff_A_hXttFBOs2_0),.din(w_dff_A_4btOcuhR0_2),.clk(gclk));
	jdff dff_A_hXttFBOs2_0(.dout(w_dff_A_NvtMBi6u3_0),.din(w_dff_A_hXttFBOs2_0),.clk(gclk));
	jdff dff_A_NvtMBi6u3_0(.dout(w_dff_A_03ZgzymL3_0),.din(w_dff_A_NvtMBi6u3_0),.clk(gclk));
	jdff dff_A_03ZgzymL3_0(.dout(w_dff_A_y94CJZe51_0),.din(w_dff_A_03ZgzymL3_0),.clk(gclk));
	jdff dff_A_y94CJZe51_0(.dout(w_dff_A_oYuZa7Dx0_0),.din(w_dff_A_y94CJZe51_0),.clk(gclk));
	jdff dff_A_oYuZa7Dx0_0(.dout(w_dff_A_hoG73kf65_0),.din(w_dff_A_oYuZa7Dx0_0),.clk(gclk));
	jdff dff_A_hoG73kf65_0(.dout(w_dff_A_cuhbW1WL3_0),.din(w_dff_A_hoG73kf65_0),.clk(gclk));
	jdff dff_A_cuhbW1WL3_0(.dout(w_dff_A_m8zZi9If8_0),.din(w_dff_A_cuhbW1WL3_0),.clk(gclk));
	jdff dff_A_m8zZi9If8_0(.dout(w_dff_A_PD4rlpDZ4_0),.din(w_dff_A_m8zZi9If8_0),.clk(gclk));
	jdff dff_A_PD4rlpDZ4_0(.dout(w_dff_A_UZk2ijKF5_0),.din(w_dff_A_PD4rlpDZ4_0),.clk(gclk));
	jdff dff_A_UZk2ijKF5_0(.dout(w_dff_A_m7OtoNr67_0),.din(w_dff_A_UZk2ijKF5_0),.clk(gclk));
	jdff dff_A_m7OtoNr67_0(.dout(w_dff_A_mcqoY2Nm9_0),.din(w_dff_A_m7OtoNr67_0),.clk(gclk));
	jdff dff_A_mcqoY2Nm9_0(.dout(w_dff_A_Yx0d6Ig68_0),.din(w_dff_A_mcqoY2Nm9_0),.clk(gclk));
	jdff dff_A_Yx0d6Ig68_0(.dout(w_dff_A_4GUKwdtm9_0),.din(w_dff_A_Yx0d6Ig68_0),.clk(gclk));
	jdff dff_A_4GUKwdtm9_0(.dout(w_dff_A_Js0auYev8_0),.din(w_dff_A_4GUKwdtm9_0),.clk(gclk));
	jdff dff_A_Js0auYev8_0(.dout(w_dff_A_jH6ElGOA3_0),.din(w_dff_A_Js0auYev8_0),.clk(gclk));
	jdff dff_A_jH6ElGOA3_0(.dout(w_dff_A_iINnE84N6_0),.din(w_dff_A_jH6ElGOA3_0),.clk(gclk));
	jdff dff_A_iINnE84N6_0(.dout(w_dff_A_oXY8KzHG9_0),.din(w_dff_A_iINnE84N6_0),.clk(gclk));
	jdff dff_A_oXY8KzHG9_0(.dout(w_dff_A_wSsS3qDZ9_0),.din(w_dff_A_oXY8KzHG9_0),.clk(gclk));
	jdff dff_A_wSsS3qDZ9_0(.dout(w_dff_A_Tk2tLxqK3_0),.din(w_dff_A_wSsS3qDZ9_0),.clk(gclk));
	jdff dff_A_Tk2tLxqK3_0(.dout(w_dff_A_YHSGDYhC2_0),.din(w_dff_A_Tk2tLxqK3_0),.clk(gclk));
	jdff dff_A_YHSGDYhC2_0(.dout(w_dff_A_nxc5s4eE8_0),.din(w_dff_A_YHSGDYhC2_0),.clk(gclk));
	jdff dff_A_nxc5s4eE8_0(.dout(w_dff_A_C9PjyOXE4_0),.din(w_dff_A_nxc5s4eE8_0),.clk(gclk));
	jdff dff_A_C9PjyOXE4_0(.dout(w_dff_A_shMjUDjF5_0),.din(w_dff_A_C9PjyOXE4_0),.clk(gclk));
	jdff dff_A_shMjUDjF5_0(.dout(w_dff_A_WLnTsOxJ1_0),.din(w_dff_A_shMjUDjF5_0),.clk(gclk));
	jdff dff_A_WLnTsOxJ1_0(.dout(w_dff_A_Ke7AJq487_0),.din(w_dff_A_WLnTsOxJ1_0),.clk(gclk));
	jdff dff_A_Ke7AJq487_0(.dout(w_dff_A_IK6Sb2gW9_0),.din(w_dff_A_Ke7AJq487_0),.clk(gclk));
	jdff dff_A_IK6Sb2gW9_0(.dout(w_dff_A_CROxuNKx5_0),.din(w_dff_A_IK6Sb2gW9_0),.clk(gclk));
	jdff dff_A_CROxuNKx5_0(.dout(w_dff_A_6pD50PzY3_0),.din(w_dff_A_CROxuNKx5_0),.clk(gclk));
	jdff dff_A_6pD50PzY3_0(.dout(w_dff_A_DZ94IGi22_0),.din(w_dff_A_6pD50PzY3_0),.clk(gclk));
	jdff dff_A_DZ94IGi22_0(.dout(w_dff_A_Q5TRQSnK2_0),.din(w_dff_A_DZ94IGi22_0),.clk(gclk));
	jdff dff_A_Q5TRQSnK2_0(.dout(w_dff_A_qySVJRl90_0),.din(w_dff_A_Q5TRQSnK2_0),.clk(gclk));
	jdff dff_A_qySVJRl90_0(.dout(w_dff_A_oTrtil7C2_0),.din(w_dff_A_qySVJRl90_0),.clk(gclk));
	jdff dff_A_oTrtil7C2_0(.dout(w_dff_A_awa57HLB7_0),.din(w_dff_A_oTrtil7C2_0),.clk(gclk));
	jdff dff_A_awa57HLB7_0(.dout(w_dff_A_ZWbfvXf69_0),.din(w_dff_A_awa57HLB7_0),.clk(gclk));
	jdff dff_A_ZWbfvXf69_0(.dout(w_dff_A_hX1HJ0Sl6_0),.din(w_dff_A_ZWbfvXf69_0),.clk(gclk));
	jdff dff_A_hX1HJ0Sl6_0(.dout(w_dff_A_paQmIG9L8_0),.din(w_dff_A_hX1HJ0Sl6_0),.clk(gclk));
	jdff dff_A_paQmIG9L8_0(.dout(w_dff_A_wkUkTNpX6_0),.din(w_dff_A_paQmIG9L8_0),.clk(gclk));
	jdff dff_A_wkUkTNpX6_0(.dout(w_dff_A_959lsYZv3_0),.din(w_dff_A_wkUkTNpX6_0),.clk(gclk));
	jdff dff_A_959lsYZv3_0(.dout(w_dff_A_dkQiuSUf5_0),.din(w_dff_A_959lsYZv3_0),.clk(gclk));
	jdff dff_A_dkQiuSUf5_0(.dout(w_dff_A_KtPPWwrf5_0),.din(w_dff_A_dkQiuSUf5_0),.clk(gclk));
	jdff dff_A_KtPPWwrf5_0(.dout(w_dff_A_MN2bDWSH3_0),.din(w_dff_A_KtPPWwrf5_0),.clk(gclk));
	jdff dff_A_MN2bDWSH3_0(.dout(w_dff_A_CTxRTJUc4_0),.din(w_dff_A_MN2bDWSH3_0),.clk(gclk));
	jdff dff_A_CTxRTJUc4_0(.dout(w_dff_A_ppYLMWDX7_0),.din(w_dff_A_CTxRTJUc4_0),.clk(gclk));
	jdff dff_A_ppYLMWDX7_0(.dout(w_dff_A_gOKEH9Mi3_0),.din(w_dff_A_ppYLMWDX7_0),.clk(gclk));
	jdff dff_A_gOKEH9Mi3_0(.dout(w_dff_A_lwFhZSV63_0),.din(w_dff_A_gOKEH9Mi3_0),.clk(gclk));
	jdff dff_A_lwFhZSV63_0(.dout(w_dff_A_lFXtpmMq2_0),.din(w_dff_A_lwFhZSV63_0),.clk(gclk));
	jdff dff_A_lFXtpmMq2_0(.dout(w_dff_A_5IykvP8q6_0),.din(w_dff_A_lFXtpmMq2_0),.clk(gclk));
	jdff dff_A_5IykvP8q6_0(.dout(w_dff_A_D9s2Wfyp0_0),.din(w_dff_A_5IykvP8q6_0),.clk(gclk));
	jdff dff_A_D9s2Wfyp0_0(.dout(w_dff_A_903UcYyy5_0),.din(w_dff_A_D9s2Wfyp0_0),.clk(gclk));
	jdff dff_A_903UcYyy5_0(.dout(w_dff_A_MADuVCyn5_0),.din(w_dff_A_903UcYyy5_0),.clk(gclk));
	jdff dff_A_MADuVCyn5_0(.dout(w_dff_A_WJgNyte32_0),.din(w_dff_A_MADuVCyn5_0),.clk(gclk));
	jdff dff_A_WJgNyte32_0(.dout(w_dff_A_9PASpTxr3_0),.din(w_dff_A_WJgNyte32_0),.clk(gclk));
	jdff dff_A_9PASpTxr3_0(.dout(w_dff_A_ZgXvYBUH0_0),.din(w_dff_A_9PASpTxr3_0),.clk(gclk));
	jdff dff_A_ZgXvYBUH0_0(.dout(w_dff_A_dnv5g5VS8_0),.din(w_dff_A_ZgXvYBUH0_0),.clk(gclk));
	jdff dff_A_dnv5g5VS8_0(.dout(w_dff_A_vr9q5a4S4_0),.din(w_dff_A_dnv5g5VS8_0),.clk(gclk));
	jdff dff_A_vr9q5a4S4_0(.dout(w_dff_A_7q12eyA13_0),.din(w_dff_A_vr9q5a4S4_0),.clk(gclk));
	jdff dff_A_7q12eyA13_0(.dout(w_dff_A_OjjTLHzT5_0),.din(w_dff_A_7q12eyA13_0),.clk(gclk));
	jdff dff_A_OjjTLHzT5_0(.dout(w_dff_A_BaVuN3mm1_0),.din(w_dff_A_OjjTLHzT5_0),.clk(gclk));
	jdff dff_A_BaVuN3mm1_0(.dout(w_dff_A_9VScVT5G7_0),.din(w_dff_A_BaVuN3mm1_0),.clk(gclk));
	jdff dff_A_9VScVT5G7_0(.dout(w_dff_A_yCVnoLKQ1_0),.din(w_dff_A_9VScVT5G7_0),.clk(gclk));
	jdff dff_A_yCVnoLKQ1_0(.dout(w_dff_A_iSAmVDXf0_0),.din(w_dff_A_yCVnoLKQ1_0),.clk(gclk));
	jdff dff_A_iSAmVDXf0_0(.dout(w_dff_A_09faWQrZ7_0),.din(w_dff_A_iSAmVDXf0_0),.clk(gclk));
	jdff dff_A_09faWQrZ7_0(.dout(w_dff_A_Z3QjOCNN7_0),.din(w_dff_A_09faWQrZ7_0),.clk(gclk));
	jdff dff_A_Z3QjOCNN7_0(.dout(w_dff_A_iQgFg42F6_0),.din(w_dff_A_Z3QjOCNN7_0),.clk(gclk));
	jdff dff_A_iQgFg42F6_0(.dout(w_dff_A_WMZk7W2y7_0),.din(w_dff_A_iQgFg42F6_0),.clk(gclk));
	jdff dff_A_WMZk7W2y7_0(.dout(w_dff_A_oVGfMUpW3_0),.din(w_dff_A_WMZk7W2y7_0),.clk(gclk));
	jdff dff_A_oVGfMUpW3_0(.dout(w_dff_A_gmPSRknr4_0),.din(w_dff_A_oVGfMUpW3_0),.clk(gclk));
	jdff dff_A_gmPSRknr4_0(.dout(w_dff_A_FbCGl2cr6_0),.din(w_dff_A_gmPSRknr4_0),.clk(gclk));
	jdff dff_A_FbCGl2cr6_0(.dout(w_dff_A_O8zju9cV9_0),.din(w_dff_A_FbCGl2cr6_0),.clk(gclk));
	jdff dff_A_O8zju9cV9_0(.dout(w_dff_A_3wkPSCpg4_0),.din(w_dff_A_O8zju9cV9_0),.clk(gclk));
	jdff dff_A_3wkPSCpg4_0(.dout(w_dff_A_u5nLHFer9_0),.din(w_dff_A_3wkPSCpg4_0),.clk(gclk));
	jdff dff_A_u5nLHFer9_0(.dout(w_dff_A_mGWophlX7_0),.din(w_dff_A_u5nLHFer9_0),.clk(gclk));
	jdff dff_A_mGWophlX7_0(.dout(w_dff_A_D8zotPIB7_0),.din(w_dff_A_mGWophlX7_0),.clk(gclk));
	jdff dff_A_D8zotPIB7_0(.dout(w_dff_A_ZOKX4UXf0_0),.din(w_dff_A_D8zotPIB7_0),.clk(gclk));
	jdff dff_A_ZOKX4UXf0_0(.dout(w_dff_A_EMskCxFE2_0),.din(w_dff_A_ZOKX4UXf0_0),.clk(gclk));
	jdff dff_A_EMskCxFE2_0(.dout(w_dff_A_SSE4Bm1T4_0),.din(w_dff_A_EMskCxFE2_0),.clk(gclk));
	jdff dff_A_SSE4Bm1T4_0(.dout(w_dff_A_Whknq80S8_0),.din(w_dff_A_SSE4Bm1T4_0),.clk(gclk));
	jdff dff_A_Whknq80S8_0(.dout(w_dff_A_kf3sdHL45_0),.din(w_dff_A_Whknq80S8_0),.clk(gclk));
	jdff dff_A_kf3sdHL45_0(.dout(w_dff_A_sqeAyzXR3_0),.din(w_dff_A_kf3sdHL45_0),.clk(gclk));
	jdff dff_A_sqeAyzXR3_0(.dout(w_dff_A_hNqkMtzr7_0),.din(w_dff_A_sqeAyzXR3_0),.clk(gclk));
	jdff dff_A_hNqkMtzr7_0(.dout(w_dff_A_ZDeP8kxK7_0),.din(w_dff_A_hNqkMtzr7_0),.clk(gclk));
	jdff dff_A_ZDeP8kxK7_0(.dout(w_dff_A_ZE0cJZ223_0),.din(w_dff_A_ZDeP8kxK7_0),.clk(gclk));
	jdff dff_A_ZE0cJZ223_0(.dout(w_dff_A_iXdsnQH82_0),.din(w_dff_A_ZE0cJZ223_0),.clk(gclk));
	jdff dff_A_iXdsnQH82_0(.dout(w_dff_A_Rgooxdmk6_0),.din(w_dff_A_iXdsnQH82_0),.clk(gclk));
	jdff dff_A_Rgooxdmk6_0(.dout(w_dff_A_FRqZLU7g3_0),.din(w_dff_A_Rgooxdmk6_0),.clk(gclk));
	jdff dff_A_FRqZLU7g3_0(.dout(w_dff_A_WkppzNmy0_0),.din(w_dff_A_FRqZLU7g3_0),.clk(gclk));
	jdff dff_A_WkppzNmy0_0(.dout(w_dff_A_OLWEjz9g8_0),.din(w_dff_A_WkppzNmy0_0),.clk(gclk));
	jdff dff_A_OLWEjz9g8_0(.dout(w_dff_A_q8xt3tDc8_0),.din(w_dff_A_OLWEjz9g8_0),.clk(gclk));
	jdff dff_A_q8xt3tDc8_0(.dout(w_dff_A_WLIDP5Zz4_0),.din(w_dff_A_q8xt3tDc8_0),.clk(gclk));
	jdff dff_A_WLIDP5Zz4_0(.dout(w_dff_A_GNTGMBKc9_0),.din(w_dff_A_WLIDP5Zz4_0),.clk(gclk));
	jdff dff_A_GNTGMBKc9_0(.dout(w_dff_A_sHjPr8Sp6_0),.din(w_dff_A_GNTGMBKc9_0),.clk(gclk));
	jdff dff_A_sHjPr8Sp6_0(.dout(w_dff_A_wMIC8CQo7_0),.din(w_dff_A_sHjPr8Sp6_0),.clk(gclk));
	jdff dff_A_wMIC8CQo7_0(.dout(w_dff_A_HYOM6pDn3_0),.din(w_dff_A_wMIC8CQo7_0),.clk(gclk));
	jdff dff_A_HYOM6pDn3_0(.dout(w_dff_A_DcSnrUzy5_0),.din(w_dff_A_HYOM6pDn3_0),.clk(gclk));
	jdff dff_A_DcSnrUzy5_0(.dout(w_dff_A_d8TqntnM0_0),.din(w_dff_A_DcSnrUzy5_0),.clk(gclk));
	jdff dff_A_d8TqntnM0_0(.dout(w_dff_A_9KmiWiT92_0),.din(w_dff_A_d8TqntnM0_0),.clk(gclk));
	jdff dff_A_9KmiWiT92_0(.dout(w_dff_A_CT2Q01WD5_0),.din(w_dff_A_9KmiWiT92_0),.clk(gclk));
	jdff dff_A_CT2Q01WD5_0(.dout(w_dff_A_AN1R04cO2_0),.din(w_dff_A_CT2Q01WD5_0),.clk(gclk));
	jdff dff_A_AN1R04cO2_0(.dout(w_dff_A_V85UJkYn6_0),.din(w_dff_A_AN1R04cO2_0),.clk(gclk));
	jdff dff_A_V85UJkYn6_0(.dout(w_dff_A_bP85bTp89_0),.din(w_dff_A_V85UJkYn6_0),.clk(gclk));
	jdff dff_A_bP85bTp89_0(.dout(w_dff_A_JyAypsUK6_0),.din(w_dff_A_bP85bTp89_0),.clk(gclk));
	jdff dff_A_JyAypsUK6_0(.dout(w_dff_A_T9KwLQ7H4_0),.din(w_dff_A_JyAypsUK6_0),.clk(gclk));
	jdff dff_A_T9KwLQ7H4_0(.dout(w_dff_A_1GdOwlCq2_0),.din(w_dff_A_T9KwLQ7H4_0),.clk(gclk));
	jdff dff_A_1GdOwlCq2_0(.dout(w_dff_A_7Vw4aZnR7_0),.din(w_dff_A_1GdOwlCq2_0),.clk(gclk));
	jdff dff_A_7Vw4aZnR7_0(.dout(w_dff_A_WU4B3Z2E4_0),.din(w_dff_A_7Vw4aZnR7_0),.clk(gclk));
	jdff dff_A_WU4B3Z2E4_0(.dout(w_dff_A_Nde80F1o6_0),.din(w_dff_A_WU4B3Z2E4_0),.clk(gclk));
	jdff dff_A_Nde80F1o6_0(.dout(w_dff_A_E2eAmiMl8_0),.din(w_dff_A_Nde80F1o6_0),.clk(gclk));
	jdff dff_A_E2eAmiMl8_0(.dout(w_dff_A_911xVSQE4_0),.din(w_dff_A_E2eAmiMl8_0),.clk(gclk));
	jdff dff_A_911xVSQE4_0(.dout(w_dff_A_SYbQqYQ70_0),.din(w_dff_A_911xVSQE4_0),.clk(gclk));
	jdff dff_A_SYbQqYQ70_0(.dout(w_dff_A_AUQl2ueY1_0),.din(w_dff_A_SYbQqYQ70_0),.clk(gclk));
	jdff dff_A_AUQl2ueY1_0(.dout(w_dff_A_PkaHEOyh8_0),.din(w_dff_A_AUQl2ueY1_0),.clk(gclk));
	jdff dff_A_PkaHEOyh8_0(.dout(w_dff_A_I02I6plj8_0),.din(w_dff_A_PkaHEOyh8_0),.clk(gclk));
	jdff dff_A_I02I6plj8_0(.dout(f13),.din(w_dff_A_I02I6plj8_0),.clk(gclk));
	jdff dff_A_KPqmqRhW5_2(.dout(w_dff_A_SgEdjVGx2_0),.din(w_dff_A_KPqmqRhW5_2),.clk(gclk));
	jdff dff_A_SgEdjVGx2_0(.dout(w_dff_A_HetkYEha4_0),.din(w_dff_A_SgEdjVGx2_0),.clk(gclk));
	jdff dff_A_HetkYEha4_0(.dout(w_dff_A_FH4ChRH80_0),.din(w_dff_A_HetkYEha4_0),.clk(gclk));
	jdff dff_A_FH4ChRH80_0(.dout(w_dff_A_3cukWHsP5_0),.din(w_dff_A_FH4ChRH80_0),.clk(gclk));
	jdff dff_A_3cukWHsP5_0(.dout(w_dff_A_hm9tdfo84_0),.din(w_dff_A_3cukWHsP5_0),.clk(gclk));
	jdff dff_A_hm9tdfo84_0(.dout(w_dff_A_abnwBoSd5_0),.din(w_dff_A_hm9tdfo84_0),.clk(gclk));
	jdff dff_A_abnwBoSd5_0(.dout(w_dff_A_KyhkWLMK4_0),.din(w_dff_A_abnwBoSd5_0),.clk(gclk));
	jdff dff_A_KyhkWLMK4_0(.dout(w_dff_A_mB5zRLED2_0),.din(w_dff_A_KyhkWLMK4_0),.clk(gclk));
	jdff dff_A_mB5zRLED2_0(.dout(w_dff_A_MtOVPXtJ6_0),.din(w_dff_A_mB5zRLED2_0),.clk(gclk));
	jdff dff_A_MtOVPXtJ6_0(.dout(w_dff_A_vx89dJhg2_0),.din(w_dff_A_MtOVPXtJ6_0),.clk(gclk));
	jdff dff_A_vx89dJhg2_0(.dout(w_dff_A_mApcxBhK0_0),.din(w_dff_A_vx89dJhg2_0),.clk(gclk));
	jdff dff_A_mApcxBhK0_0(.dout(w_dff_A_1Bw9t0Vv9_0),.din(w_dff_A_mApcxBhK0_0),.clk(gclk));
	jdff dff_A_1Bw9t0Vv9_0(.dout(w_dff_A_WUYuQ3Ax1_0),.din(w_dff_A_1Bw9t0Vv9_0),.clk(gclk));
	jdff dff_A_WUYuQ3Ax1_0(.dout(w_dff_A_tE06Q4IP3_0),.din(w_dff_A_WUYuQ3Ax1_0),.clk(gclk));
	jdff dff_A_tE06Q4IP3_0(.dout(w_dff_A_t6Yvze558_0),.din(w_dff_A_tE06Q4IP3_0),.clk(gclk));
	jdff dff_A_t6Yvze558_0(.dout(w_dff_A_vnJpdQZV7_0),.din(w_dff_A_t6Yvze558_0),.clk(gclk));
	jdff dff_A_vnJpdQZV7_0(.dout(w_dff_A_kw3bRMWl0_0),.din(w_dff_A_vnJpdQZV7_0),.clk(gclk));
	jdff dff_A_kw3bRMWl0_0(.dout(w_dff_A_3SqsgBYE9_0),.din(w_dff_A_kw3bRMWl0_0),.clk(gclk));
	jdff dff_A_3SqsgBYE9_0(.dout(w_dff_A_OtfD1YTa1_0),.din(w_dff_A_3SqsgBYE9_0),.clk(gclk));
	jdff dff_A_OtfD1YTa1_0(.dout(w_dff_A_vrtYWndX5_0),.din(w_dff_A_OtfD1YTa1_0),.clk(gclk));
	jdff dff_A_vrtYWndX5_0(.dout(w_dff_A_czRBBvUL5_0),.din(w_dff_A_vrtYWndX5_0),.clk(gclk));
	jdff dff_A_czRBBvUL5_0(.dout(w_dff_A_vRp4RSR39_0),.din(w_dff_A_czRBBvUL5_0),.clk(gclk));
	jdff dff_A_vRp4RSR39_0(.dout(w_dff_A_IGtA3qJy1_0),.din(w_dff_A_vRp4RSR39_0),.clk(gclk));
	jdff dff_A_IGtA3qJy1_0(.dout(w_dff_A_jKrfyg6H5_0),.din(w_dff_A_IGtA3qJy1_0),.clk(gclk));
	jdff dff_A_jKrfyg6H5_0(.dout(w_dff_A_0muZVTpA4_0),.din(w_dff_A_jKrfyg6H5_0),.clk(gclk));
	jdff dff_A_0muZVTpA4_0(.dout(w_dff_A_lPGHCTwF3_0),.din(w_dff_A_0muZVTpA4_0),.clk(gclk));
	jdff dff_A_lPGHCTwF3_0(.dout(w_dff_A_PK428G8O8_0),.din(w_dff_A_lPGHCTwF3_0),.clk(gclk));
	jdff dff_A_PK428G8O8_0(.dout(w_dff_A_CTONW30k7_0),.din(w_dff_A_PK428G8O8_0),.clk(gclk));
	jdff dff_A_CTONW30k7_0(.dout(w_dff_A_qEYXtEOp1_0),.din(w_dff_A_CTONW30k7_0),.clk(gclk));
	jdff dff_A_qEYXtEOp1_0(.dout(w_dff_A_EdgR7YUl9_0),.din(w_dff_A_qEYXtEOp1_0),.clk(gclk));
	jdff dff_A_EdgR7YUl9_0(.dout(w_dff_A_aqlmcIsW4_0),.din(w_dff_A_EdgR7YUl9_0),.clk(gclk));
	jdff dff_A_aqlmcIsW4_0(.dout(w_dff_A_5TzlW5AR2_0),.din(w_dff_A_aqlmcIsW4_0),.clk(gclk));
	jdff dff_A_5TzlW5AR2_0(.dout(w_dff_A_D39lk0xg3_0),.din(w_dff_A_5TzlW5AR2_0),.clk(gclk));
	jdff dff_A_D39lk0xg3_0(.dout(w_dff_A_UM0DZMHy4_0),.din(w_dff_A_D39lk0xg3_0),.clk(gclk));
	jdff dff_A_UM0DZMHy4_0(.dout(w_dff_A_2JFILxsC6_0),.din(w_dff_A_UM0DZMHy4_0),.clk(gclk));
	jdff dff_A_2JFILxsC6_0(.dout(w_dff_A_NEVK5IJE1_0),.din(w_dff_A_2JFILxsC6_0),.clk(gclk));
	jdff dff_A_NEVK5IJE1_0(.dout(w_dff_A_zyzHFxkr2_0),.din(w_dff_A_NEVK5IJE1_0),.clk(gclk));
	jdff dff_A_zyzHFxkr2_0(.dout(w_dff_A_xlZHsfPf5_0),.din(w_dff_A_zyzHFxkr2_0),.clk(gclk));
	jdff dff_A_xlZHsfPf5_0(.dout(w_dff_A_vEICNVV24_0),.din(w_dff_A_xlZHsfPf5_0),.clk(gclk));
	jdff dff_A_vEICNVV24_0(.dout(w_dff_A_iuatYexV2_0),.din(w_dff_A_vEICNVV24_0),.clk(gclk));
	jdff dff_A_iuatYexV2_0(.dout(w_dff_A_rKCpqKrG3_0),.din(w_dff_A_iuatYexV2_0),.clk(gclk));
	jdff dff_A_rKCpqKrG3_0(.dout(w_dff_A_CqEKkPbK0_0),.din(w_dff_A_rKCpqKrG3_0),.clk(gclk));
	jdff dff_A_CqEKkPbK0_0(.dout(w_dff_A_TQXV4JQl7_0),.din(w_dff_A_CqEKkPbK0_0),.clk(gclk));
	jdff dff_A_TQXV4JQl7_0(.dout(w_dff_A_UabOpz156_0),.din(w_dff_A_TQXV4JQl7_0),.clk(gclk));
	jdff dff_A_UabOpz156_0(.dout(w_dff_A_5HSLAxjs0_0),.din(w_dff_A_UabOpz156_0),.clk(gclk));
	jdff dff_A_5HSLAxjs0_0(.dout(w_dff_A_74n0dB3u6_0),.din(w_dff_A_5HSLAxjs0_0),.clk(gclk));
	jdff dff_A_74n0dB3u6_0(.dout(w_dff_A_yFPpCaQx4_0),.din(w_dff_A_74n0dB3u6_0),.clk(gclk));
	jdff dff_A_yFPpCaQx4_0(.dout(w_dff_A_c4edFJCv7_0),.din(w_dff_A_yFPpCaQx4_0),.clk(gclk));
	jdff dff_A_c4edFJCv7_0(.dout(w_dff_A_lDQQ5RYS4_0),.din(w_dff_A_c4edFJCv7_0),.clk(gclk));
	jdff dff_A_lDQQ5RYS4_0(.dout(w_dff_A_XnkbO31U1_0),.din(w_dff_A_lDQQ5RYS4_0),.clk(gclk));
	jdff dff_A_XnkbO31U1_0(.dout(w_dff_A_DzICmh9B7_0),.din(w_dff_A_XnkbO31U1_0),.clk(gclk));
	jdff dff_A_DzICmh9B7_0(.dout(w_dff_A_dcAgGSrA6_0),.din(w_dff_A_DzICmh9B7_0),.clk(gclk));
	jdff dff_A_dcAgGSrA6_0(.dout(w_dff_A_K2pbJSQb0_0),.din(w_dff_A_dcAgGSrA6_0),.clk(gclk));
	jdff dff_A_K2pbJSQb0_0(.dout(w_dff_A_GQwykDTQ5_0),.din(w_dff_A_K2pbJSQb0_0),.clk(gclk));
	jdff dff_A_GQwykDTQ5_0(.dout(w_dff_A_EXnHnrBS4_0),.din(w_dff_A_GQwykDTQ5_0),.clk(gclk));
	jdff dff_A_EXnHnrBS4_0(.dout(w_dff_A_v9AW4DIs7_0),.din(w_dff_A_EXnHnrBS4_0),.clk(gclk));
	jdff dff_A_v9AW4DIs7_0(.dout(w_dff_A_HNUIv0sg7_0),.din(w_dff_A_v9AW4DIs7_0),.clk(gclk));
	jdff dff_A_HNUIv0sg7_0(.dout(w_dff_A_dfeB26CL8_0),.din(w_dff_A_HNUIv0sg7_0),.clk(gclk));
	jdff dff_A_dfeB26CL8_0(.dout(w_dff_A_SqOiAhrx1_0),.din(w_dff_A_dfeB26CL8_0),.clk(gclk));
	jdff dff_A_SqOiAhrx1_0(.dout(w_dff_A_s8GkfFRS9_0),.din(w_dff_A_SqOiAhrx1_0),.clk(gclk));
	jdff dff_A_s8GkfFRS9_0(.dout(w_dff_A_UNxOZJac6_0),.din(w_dff_A_s8GkfFRS9_0),.clk(gclk));
	jdff dff_A_UNxOZJac6_0(.dout(w_dff_A_NjGcVTVh4_0),.din(w_dff_A_UNxOZJac6_0),.clk(gclk));
	jdff dff_A_NjGcVTVh4_0(.dout(w_dff_A_Xi0GEigo5_0),.din(w_dff_A_NjGcVTVh4_0),.clk(gclk));
	jdff dff_A_Xi0GEigo5_0(.dout(w_dff_A_hCSux4bt4_0),.din(w_dff_A_Xi0GEigo5_0),.clk(gclk));
	jdff dff_A_hCSux4bt4_0(.dout(w_dff_A_Q0QoWgoU9_0),.din(w_dff_A_hCSux4bt4_0),.clk(gclk));
	jdff dff_A_Q0QoWgoU9_0(.dout(w_dff_A_6Ey0CQTk8_0),.din(w_dff_A_Q0QoWgoU9_0),.clk(gclk));
	jdff dff_A_6Ey0CQTk8_0(.dout(w_dff_A_DezHMF1g1_0),.din(w_dff_A_6Ey0CQTk8_0),.clk(gclk));
	jdff dff_A_DezHMF1g1_0(.dout(w_dff_A_tzD4vyM12_0),.din(w_dff_A_DezHMF1g1_0),.clk(gclk));
	jdff dff_A_tzD4vyM12_0(.dout(w_dff_A_H186WLXv5_0),.din(w_dff_A_tzD4vyM12_0),.clk(gclk));
	jdff dff_A_H186WLXv5_0(.dout(w_dff_A_nmNhH4aX5_0),.din(w_dff_A_H186WLXv5_0),.clk(gclk));
	jdff dff_A_nmNhH4aX5_0(.dout(w_dff_A_CGWHNEyM2_0),.din(w_dff_A_nmNhH4aX5_0),.clk(gclk));
	jdff dff_A_CGWHNEyM2_0(.dout(w_dff_A_pSnjdBT06_0),.din(w_dff_A_CGWHNEyM2_0),.clk(gclk));
	jdff dff_A_pSnjdBT06_0(.dout(w_dff_A_YukesCli4_0),.din(w_dff_A_pSnjdBT06_0),.clk(gclk));
	jdff dff_A_YukesCli4_0(.dout(w_dff_A_f9DTe8DA1_0),.din(w_dff_A_YukesCli4_0),.clk(gclk));
	jdff dff_A_f9DTe8DA1_0(.dout(w_dff_A_F5QjwUTG0_0),.din(w_dff_A_f9DTe8DA1_0),.clk(gclk));
	jdff dff_A_F5QjwUTG0_0(.dout(w_dff_A_SxUiaafq4_0),.din(w_dff_A_F5QjwUTG0_0),.clk(gclk));
	jdff dff_A_SxUiaafq4_0(.dout(w_dff_A_D5JkIpho2_0),.din(w_dff_A_SxUiaafq4_0),.clk(gclk));
	jdff dff_A_D5JkIpho2_0(.dout(w_dff_A_f53AXXp54_0),.din(w_dff_A_D5JkIpho2_0),.clk(gclk));
	jdff dff_A_f53AXXp54_0(.dout(w_dff_A_8hkLduPJ5_0),.din(w_dff_A_f53AXXp54_0),.clk(gclk));
	jdff dff_A_8hkLduPJ5_0(.dout(w_dff_A_TbkNVXXF9_0),.din(w_dff_A_8hkLduPJ5_0),.clk(gclk));
	jdff dff_A_TbkNVXXF9_0(.dout(w_dff_A_9B3bhSv31_0),.din(w_dff_A_TbkNVXXF9_0),.clk(gclk));
	jdff dff_A_9B3bhSv31_0(.dout(w_dff_A_0NWDLrLV9_0),.din(w_dff_A_9B3bhSv31_0),.clk(gclk));
	jdff dff_A_0NWDLrLV9_0(.dout(w_dff_A_CdA1pW6V7_0),.din(w_dff_A_0NWDLrLV9_0),.clk(gclk));
	jdff dff_A_CdA1pW6V7_0(.dout(w_dff_A_dP6BUQ6o9_0),.din(w_dff_A_CdA1pW6V7_0),.clk(gclk));
	jdff dff_A_dP6BUQ6o9_0(.dout(w_dff_A_zwJ9pYKE7_0),.din(w_dff_A_dP6BUQ6o9_0),.clk(gclk));
	jdff dff_A_zwJ9pYKE7_0(.dout(w_dff_A_pHlrahvY2_0),.din(w_dff_A_zwJ9pYKE7_0),.clk(gclk));
	jdff dff_A_pHlrahvY2_0(.dout(w_dff_A_4BsRjjQK7_0),.din(w_dff_A_pHlrahvY2_0),.clk(gclk));
	jdff dff_A_4BsRjjQK7_0(.dout(w_dff_A_5RTGDfZC7_0),.din(w_dff_A_4BsRjjQK7_0),.clk(gclk));
	jdff dff_A_5RTGDfZC7_0(.dout(w_dff_A_BkQHaBjS7_0),.din(w_dff_A_5RTGDfZC7_0),.clk(gclk));
	jdff dff_A_BkQHaBjS7_0(.dout(w_dff_A_c8tUtC9C0_0),.din(w_dff_A_BkQHaBjS7_0),.clk(gclk));
	jdff dff_A_c8tUtC9C0_0(.dout(w_dff_A_b9qcIKjf4_0),.din(w_dff_A_c8tUtC9C0_0),.clk(gclk));
	jdff dff_A_b9qcIKjf4_0(.dout(w_dff_A_ijFYYkgr2_0),.din(w_dff_A_b9qcIKjf4_0),.clk(gclk));
	jdff dff_A_ijFYYkgr2_0(.dout(w_dff_A_VW6FtWRb6_0),.din(w_dff_A_ijFYYkgr2_0),.clk(gclk));
	jdff dff_A_VW6FtWRb6_0(.dout(w_dff_A_jpkbdgbo6_0),.din(w_dff_A_VW6FtWRb6_0),.clk(gclk));
	jdff dff_A_jpkbdgbo6_0(.dout(w_dff_A_fHGKWQYF2_0),.din(w_dff_A_jpkbdgbo6_0),.clk(gclk));
	jdff dff_A_fHGKWQYF2_0(.dout(w_dff_A_WmNQ3cQ84_0),.din(w_dff_A_fHGKWQYF2_0),.clk(gclk));
	jdff dff_A_WmNQ3cQ84_0(.dout(w_dff_A_efv7ck776_0),.din(w_dff_A_WmNQ3cQ84_0),.clk(gclk));
	jdff dff_A_efv7ck776_0(.dout(w_dff_A_Trn2HCBl7_0),.din(w_dff_A_efv7ck776_0),.clk(gclk));
	jdff dff_A_Trn2HCBl7_0(.dout(w_dff_A_iPbWYITl4_0),.din(w_dff_A_Trn2HCBl7_0),.clk(gclk));
	jdff dff_A_iPbWYITl4_0(.dout(w_dff_A_p483Fs4E8_0),.din(w_dff_A_iPbWYITl4_0),.clk(gclk));
	jdff dff_A_p483Fs4E8_0(.dout(w_dff_A_3xps0bi00_0),.din(w_dff_A_p483Fs4E8_0),.clk(gclk));
	jdff dff_A_3xps0bi00_0(.dout(w_dff_A_96dI2mB01_0),.din(w_dff_A_3xps0bi00_0),.clk(gclk));
	jdff dff_A_96dI2mB01_0(.dout(w_dff_A_9BsK8oIj7_0),.din(w_dff_A_96dI2mB01_0),.clk(gclk));
	jdff dff_A_9BsK8oIj7_0(.dout(w_dff_A_mcXaiTRj5_0),.din(w_dff_A_9BsK8oIj7_0),.clk(gclk));
	jdff dff_A_mcXaiTRj5_0(.dout(w_dff_A_oRANdWsb5_0),.din(w_dff_A_mcXaiTRj5_0),.clk(gclk));
	jdff dff_A_oRANdWsb5_0(.dout(w_dff_A_UFtg8Tvl1_0),.din(w_dff_A_oRANdWsb5_0),.clk(gclk));
	jdff dff_A_UFtg8Tvl1_0(.dout(w_dff_A_Ge4dLXhI6_0),.din(w_dff_A_UFtg8Tvl1_0),.clk(gclk));
	jdff dff_A_Ge4dLXhI6_0(.dout(w_dff_A_yucONrb61_0),.din(w_dff_A_Ge4dLXhI6_0),.clk(gclk));
	jdff dff_A_yucONrb61_0(.dout(w_dff_A_16ubPdRp1_0),.din(w_dff_A_yucONrb61_0),.clk(gclk));
	jdff dff_A_16ubPdRp1_0(.dout(w_dff_A_6Y58dUmr3_0),.din(w_dff_A_16ubPdRp1_0),.clk(gclk));
	jdff dff_A_6Y58dUmr3_0(.dout(w_dff_A_IB8T7nYI1_0),.din(w_dff_A_6Y58dUmr3_0),.clk(gclk));
	jdff dff_A_IB8T7nYI1_0(.dout(w_dff_A_QpC3Hlss6_0),.din(w_dff_A_IB8T7nYI1_0),.clk(gclk));
	jdff dff_A_QpC3Hlss6_0(.dout(f14),.din(w_dff_A_QpC3Hlss6_0),.clk(gclk));
	jdff dff_A_3a83FO075_2(.dout(w_dff_A_R5ZzPwYw2_0),.din(w_dff_A_3a83FO075_2),.clk(gclk));
	jdff dff_A_R5ZzPwYw2_0(.dout(w_dff_A_unp3g2o18_0),.din(w_dff_A_R5ZzPwYw2_0),.clk(gclk));
	jdff dff_A_unp3g2o18_0(.dout(w_dff_A_eYMK1qX39_0),.din(w_dff_A_unp3g2o18_0),.clk(gclk));
	jdff dff_A_eYMK1qX39_0(.dout(w_dff_A_EaUr1SQN4_0),.din(w_dff_A_eYMK1qX39_0),.clk(gclk));
	jdff dff_A_EaUr1SQN4_0(.dout(w_dff_A_NuzNO3OM4_0),.din(w_dff_A_EaUr1SQN4_0),.clk(gclk));
	jdff dff_A_NuzNO3OM4_0(.dout(w_dff_A_sfNFdMeh4_0),.din(w_dff_A_NuzNO3OM4_0),.clk(gclk));
	jdff dff_A_sfNFdMeh4_0(.dout(w_dff_A_3j91GzBb3_0),.din(w_dff_A_sfNFdMeh4_0),.clk(gclk));
	jdff dff_A_3j91GzBb3_0(.dout(w_dff_A_N2MMRaGm8_0),.din(w_dff_A_3j91GzBb3_0),.clk(gclk));
	jdff dff_A_N2MMRaGm8_0(.dout(w_dff_A_DZP6L6OB8_0),.din(w_dff_A_N2MMRaGm8_0),.clk(gclk));
	jdff dff_A_DZP6L6OB8_0(.dout(w_dff_A_pk7boYRo2_0),.din(w_dff_A_DZP6L6OB8_0),.clk(gclk));
	jdff dff_A_pk7boYRo2_0(.dout(w_dff_A_3qZArAa61_0),.din(w_dff_A_pk7boYRo2_0),.clk(gclk));
	jdff dff_A_3qZArAa61_0(.dout(w_dff_A_tDox3vvh5_0),.din(w_dff_A_3qZArAa61_0),.clk(gclk));
	jdff dff_A_tDox3vvh5_0(.dout(w_dff_A_cNGGygDf1_0),.din(w_dff_A_tDox3vvh5_0),.clk(gclk));
	jdff dff_A_cNGGygDf1_0(.dout(w_dff_A_IGh0fp031_0),.din(w_dff_A_cNGGygDf1_0),.clk(gclk));
	jdff dff_A_IGh0fp031_0(.dout(w_dff_A_WdwOJxi03_0),.din(w_dff_A_IGh0fp031_0),.clk(gclk));
	jdff dff_A_WdwOJxi03_0(.dout(w_dff_A_NL3YWKon8_0),.din(w_dff_A_WdwOJxi03_0),.clk(gclk));
	jdff dff_A_NL3YWKon8_0(.dout(w_dff_A_gjwROSFG1_0),.din(w_dff_A_NL3YWKon8_0),.clk(gclk));
	jdff dff_A_gjwROSFG1_0(.dout(w_dff_A_4JmmDfE36_0),.din(w_dff_A_gjwROSFG1_0),.clk(gclk));
	jdff dff_A_4JmmDfE36_0(.dout(w_dff_A_WeoA5Rhf4_0),.din(w_dff_A_4JmmDfE36_0),.clk(gclk));
	jdff dff_A_WeoA5Rhf4_0(.dout(w_dff_A_loOnmAaY9_0),.din(w_dff_A_WeoA5Rhf4_0),.clk(gclk));
	jdff dff_A_loOnmAaY9_0(.dout(w_dff_A_YSxOoQvQ5_0),.din(w_dff_A_loOnmAaY9_0),.clk(gclk));
	jdff dff_A_YSxOoQvQ5_0(.dout(w_dff_A_lHSMrh6f6_0),.din(w_dff_A_YSxOoQvQ5_0),.clk(gclk));
	jdff dff_A_lHSMrh6f6_0(.dout(w_dff_A_M8U3bskl4_0),.din(w_dff_A_lHSMrh6f6_0),.clk(gclk));
	jdff dff_A_M8U3bskl4_0(.dout(w_dff_A_87QjXuSx7_0),.din(w_dff_A_M8U3bskl4_0),.clk(gclk));
	jdff dff_A_87QjXuSx7_0(.dout(w_dff_A_59sXhw6V9_0),.din(w_dff_A_87QjXuSx7_0),.clk(gclk));
	jdff dff_A_59sXhw6V9_0(.dout(w_dff_A_jpEupxkm3_0),.din(w_dff_A_59sXhw6V9_0),.clk(gclk));
	jdff dff_A_jpEupxkm3_0(.dout(w_dff_A_4PHBpZHu2_0),.din(w_dff_A_jpEupxkm3_0),.clk(gclk));
	jdff dff_A_4PHBpZHu2_0(.dout(w_dff_A_VTL1HRAQ7_0),.din(w_dff_A_4PHBpZHu2_0),.clk(gclk));
	jdff dff_A_VTL1HRAQ7_0(.dout(w_dff_A_t9adHGTj8_0),.din(w_dff_A_VTL1HRAQ7_0),.clk(gclk));
	jdff dff_A_t9adHGTj8_0(.dout(w_dff_A_i9JuflxC9_0),.din(w_dff_A_t9adHGTj8_0),.clk(gclk));
	jdff dff_A_i9JuflxC9_0(.dout(w_dff_A_PE6HJHdD0_0),.din(w_dff_A_i9JuflxC9_0),.clk(gclk));
	jdff dff_A_PE6HJHdD0_0(.dout(w_dff_A_K49rF0yR2_0),.din(w_dff_A_PE6HJHdD0_0),.clk(gclk));
	jdff dff_A_K49rF0yR2_0(.dout(w_dff_A_d0fHLS2q5_0),.din(w_dff_A_K49rF0yR2_0),.clk(gclk));
	jdff dff_A_d0fHLS2q5_0(.dout(w_dff_A_MDIZ812e6_0),.din(w_dff_A_d0fHLS2q5_0),.clk(gclk));
	jdff dff_A_MDIZ812e6_0(.dout(w_dff_A_sG4CTWPm4_0),.din(w_dff_A_MDIZ812e6_0),.clk(gclk));
	jdff dff_A_sG4CTWPm4_0(.dout(w_dff_A_7xy2MAdt6_0),.din(w_dff_A_sG4CTWPm4_0),.clk(gclk));
	jdff dff_A_7xy2MAdt6_0(.dout(w_dff_A_e3Ng8x4E9_0),.din(w_dff_A_7xy2MAdt6_0),.clk(gclk));
	jdff dff_A_e3Ng8x4E9_0(.dout(w_dff_A_edfSKao57_0),.din(w_dff_A_e3Ng8x4E9_0),.clk(gclk));
	jdff dff_A_edfSKao57_0(.dout(w_dff_A_83GvkYMm0_0),.din(w_dff_A_edfSKao57_0),.clk(gclk));
	jdff dff_A_83GvkYMm0_0(.dout(w_dff_A_f7suxt9F0_0),.din(w_dff_A_83GvkYMm0_0),.clk(gclk));
	jdff dff_A_f7suxt9F0_0(.dout(w_dff_A_owo9Ua9h9_0),.din(w_dff_A_f7suxt9F0_0),.clk(gclk));
	jdff dff_A_owo9Ua9h9_0(.dout(w_dff_A_RwQSpl3F0_0),.din(w_dff_A_owo9Ua9h9_0),.clk(gclk));
	jdff dff_A_RwQSpl3F0_0(.dout(w_dff_A_sveZIsL14_0),.din(w_dff_A_RwQSpl3F0_0),.clk(gclk));
	jdff dff_A_sveZIsL14_0(.dout(w_dff_A_vwk37Yfm0_0),.din(w_dff_A_sveZIsL14_0),.clk(gclk));
	jdff dff_A_vwk37Yfm0_0(.dout(w_dff_A_7bz1RmbR8_0),.din(w_dff_A_vwk37Yfm0_0),.clk(gclk));
	jdff dff_A_7bz1RmbR8_0(.dout(w_dff_A_GIx2hT7U5_0),.din(w_dff_A_7bz1RmbR8_0),.clk(gclk));
	jdff dff_A_GIx2hT7U5_0(.dout(w_dff_A_1bKXmKbl0_0),.din(w_dff_A_GIx2hT7U5_0),.clk(gclk));
	jdff dff_A_1bKXmKbl0_0(.dout(w_dff_A_a9df2deA1_0),.din(w_dff_A_1bKXmKbl0_0),.clk(gclk));
	jdff dff_A_a9df2deA1_0(.dout(w_dff_A_4DD8ByeP8_0),.din(w_dff_A_a9df2deA1_0),.clk(gclk));
	jdff dff_A_4DD8ByeP8_0(.dout(w_dff_A_HvTO4E3w0_0),.din(w_dff_A_4DD8ByeP8_0),.clk(gclk));
	jdff dff_A_HvTO4E3w0_0(.dout(w_dff_A_i6CM3pXk4_0),.din(w_dff_A_HvTO4E3w0_0),.clk(gclk));
	jdff dff_A_i6CM3pXk4_0(.dout(w_dff_A_Zwph8O7S6_0),.din(w_dff_A_i6CM3pXk4_0),.clk(gclk));
	jdff dff_A_Zwph8O7S6_0(.dout(w_dff_A_4KREGJ5L7_0),.din(w_dff_A_Zwph8O7S6_0),.clk(gclk));
	jdff dff_A_4KREGJ5L7_0(.dout(w_dff_A_nFH0Xs6i1_0),.din(w_dff_A_4KREGJ5L7_0),.clk(gclk));
	jdff dff_A_nFH0Xs6i1_0(.dout(w_dff_A_CrnPe1sW4_0),.din(w_dff_A_nFH0Xs6i1_0),.clk(gclk));
	jdff dff_A_CrnPe1sW4_0(.dout(w_dff_A_ABcuLraL3_0),.din(w_dff_A_CrnPe1sW4_0),.clk(gclk));
	jdff dff_A_ABcuLraL3_0(.dout(w_dff_A_msE5VSQQ4_0),.din(w_dff_A_ABcuLraL3_0),.clk(gclk));
	jdff dff_A_msE5VSQQ4_0(.dout(w_dff_A_tjiL7swM1_0),.din(w_dff_A_msE5VSQQ4_0),.clk(gclk));
	jdff dff_A_tjiL7swM1_0(.dout(w_dff_A_Urgu16Ef1_0),.din(w_dff_A_tjiL7swM1_0),.clk(gclk));
	jdff dff_A_Urgu16Ef1_0(.dout(w_dff_A_RceBeY541_0),.din(w_dff_A_Urgu16Ef1_0),.clk(gclk));
	jdff dff_A_RceBeY541_0(.dout(w_dff_A_IvFCHQvF9_0),.din(w_dff_A_RceBeY541_0),.clk(gclk));
	jdff dff_A_IvFCHQvF9_0(.dout(w_dff_A_k891ORud8_0),.din(w_dff_A_IvFCHQvF9_0),.clk(gclk));
	jdff dff_A_k891ORud8_0(.dout(w_dff_A_kz74VQLS6_0),.din(w_dff_A_k891ORud8_0),.clk(gclk));
	jdff dff_A_kz74VQLS6_0(.dout(w_dff_A_fqgSZzc77_0),.din(w_dff_A_kz74VQLS6_0),.clk(gclk));
	jdff dff_A_fqgSZzc77_0(.dout(w_dff_A_fafwZQnB2_0),.din(w_dff_A_fqgSZzc77_0),.clk(gclk));
	jdff dff_A_fafwZQnB2_0(.dout(w_dff_A_tiMs8Q3l6_0),.din(w_dff_A_fafwZQnB2_0),.clk(gclk));
	jdff dff_A_tiMs8Q3l6_0(.dout(w_dff_A_ogkJcjLT2_0),.din(w_dff_A_tiMs8Q3l6_0),.clk(gclk));
	jdff dff_A_ogkJcjLT2_0(.dout(w_dff_A_C4X5lUbO2_0),.din(w_dff_A_ogkJcjLT2_0),.clk(gclk));
	jdff dff_A_C4X5lUbO2_0(.dout(w_dff_A_rNeKw7dI1_0),.din(w_dff_A_C4X5lUbO2_0),.clk(gclk));
	jdff dff_A_rNeKw7dI1_0(.dout(w_dff_A_8UcDCQ3i0_0),.din(w_dff_A_rNeKw7dI1_0),.clk(gclk));
	jdff dff_A_8UcDCQ3i0_0(.dout(w_dff_A_E8tb1b9J8_0),.din(w_dff_A_8UcDCQ3i0_0),.clk(gclk));
	jdff dff_A_E8tb1b9J8_0(.dout(w_dff_A_xndHYYXf6_0),.din(w_dff_A_E8tb1b9J8_0),.clk(gclk));
	jdff dff_A_xndHYYXf6_0(.dout(w_dff_A_gUB4rCDK7_0),.din(w_dff_A_xndHYYXf6_0),.clk(gclk));
	jdff dff_A_gUB4rCDK7_0(.dout(w_dff_A_tptklpjh5_0),.din(w_dff_A_gUB4rCDK7_0),.clk(gclk));
	jdff dff_A_tptklpjh5_0(.dout(w_dff_A_Jn8tbMwm5_0),.din(w_dff_A_tptklpjh5_0),.clk(gclk));
	jdff dff_A_Jn8tbMwm5_0(.dout(w_dff_A_w2Ir4HAT0_0),.din(w_dff_A_Jn8tbMwm5_0),.clk(gclk));
	jdff dff_A_w2Ir4HAT0_0(.dout(w_dff_A_wGQeSFoD1_0),.din(w_dff_A_w2Ir4HAT0_0),.clk(gclk));
	jdff dff_A_wGQeSFoD1_0(.dout(w_dff_A_wxSmVvdS0_0),.din(w_dff_A_wGQeSFoD1_0),.clk(gclk));
	jdff dff_A_wxSmVvdS0_0(.dout(w_dff_A_b6tAiDf00_0),.din(w_dff_A_wxSmVvdS0_0),.clk(gclk));
	jdff dff_A_b6tAiDf00_0(.dout(w_dff_A_CHbzrRqv8_0),.din(w_dff_A_b6tAiDf00_0),.clk(gclk));
	jdff dff_A_CHbzrRqv8_0(.dout(w_dff_A_fvvU2Bu84_0),.din(w_dff_A_CHbzrRqv8_0),.clk(gclk));
	jdff dff_A_fvvU2Bu84_0(.dout(w_dff_A_toWNEzfK3_0),.din(w_dff_A_fvvU2Bu84_0),.clk(gclk));
	jdff dff_A_toWNEzfK3_0(.dout(w_dff_A_fPSmFcHY0_0),.din(w_dff_A_toWNEzfK3_0),.clk(gclk));
	jdff dff_A_fPSmFcHY0_0(.dout(w_dff_A_7BnloomA7_0),.din(w_dff_A_fPSmFcHY0_0),.clk(gclk));
	jdff dff_A_7BnloomA7_0(.dout(w_dff_A_eUc7EgCD2_0),.din(w_dff_A_7BnloomA7_0),.clk(gclk));
	jdff dff_A_eUc7EgCD2_0(.dout(w_dff_A_pNNbcazj4_0),.din(w_dff_A_eUc7EgCD2_0),.clk(gclk));
	jdff dff_A_pNNbcazj4_0(.dout(w_dff_A_YkKEgnKf8_0),.din(w_dff_A_pNNbcazj4_0),.clk(gclk));
	jdff dff_A_YkKEgnKf8_0(.dout(w_dff_A_dKuJHMS67_0),.din(w_dff_A_YkKEgnKf8_0),.clk(gclk));
	jdff dff_A_dKuJHMS67_0(.dout(w_dff_A_zCf0S6xz3_0),.din(w_dff_A_dKuJHMS67_0),.clk(gclk));
	jdff dff_A_zCf0S6xz3_0(.dout(w_dff_A_5IgKgJGL1_0),.din(w_dff_A_zCf0S6xz3_0),.clk(gclk));
	jdff dff_A_5IgKgJGL1_0(.dout(w_dff_A_AOmInIwT4_0),.din(w_dff_A_5IgKgJGL1_0),.clk(gclk));
	jdff dff_A_AOmInIwT4_0(.dout(w_dff_A_BX8cZWal2_0),.din(w_dff_A_AOmInIwT4_0),.clk(gclk));
	jdff dff_A_BX8cZWal2_0(.dout(w_dff_A_8zXJQ6Xx0_0),.din(w_dff_A_BX8cZWal2_0),.clk(gclk));
	jdff dff_A_8zXJQ6Xx0_0(.dout(w_dff_A_iKuApldO0_0),.din(w_dff_A_8zXJQ6Xx0_0),.clk(gclk));
	jdff dff_A_iKuApldO0_0(.dout(w_dff_A_VBo9wto11_0),.din(w_dff_A_iKuApldO0_0),.clk(gclk));
	jdff dff_A_VBo9wto11_0(.dout(w_dff_A_rLAOYLtl7_0),.din(w_dff_A_VBo9wto11_0),.clk(gclk));
	jdff dff_A_rLAOYLtl7_0(.dout(w_dff_A_vnaebWSB6_0),.din(w_dff_A_rLAOYLtl7_0),.clk(gclk));
	jdff dff_A_vnaebWSB6_0(.dout(w_dff_A_PQ6lY9By3_0),.din(w_dff_A_vnaebWSB6_0),.clk(gclk));
	jdff dff_A_PQ6lY9By3_0(.dout(w_dff_A_IbySE8iU2_0),.din(w_dff_A_PQ6lY9By3_0),.clk(gclk));
	jdff dff_A_IbySE8iU2_0(.dout(w_dff_A_DjASBRg76_0),.din(w_dff_A_IbySE8iU2_0),.clk(gclk));
	jdff dff_A_DjASBRg76_0(.dout(w_dff_A_a6Yv4szI3_0),.din(w_dff_A_DjASBRg76_0),.clk(gclk));
	jdff dff_A_a6Yv4szI3_0(.dout(w_dff_A_Z7QZXcGI3_0),.din(w_dff_A_a6Yv4szI3_0),.clk(gclk));
	jdff dff_A_Z7QZXcGI3_0(.dout(w_dff_A_ijbCtb7n5_0),.din(w_dff_A_Z7QZXcGI3_0),.clk(gclk));
	jdff dff_A_ijbCtb7n5_0(.dout(w_dff_A_vGTkiiCQ3_0),.din(w_dff_A_ijbCtb7n5_0),.clk(gclk));
	jdff dff_A_vGTkiiCQ3_0(.dout(w_dff_A_Fh9HDm058_0),.din(w_dff_A_vGTkiiCQ3_0),.clk(gclk));
	jdff dff_A_Fh9HDm058_0(.dout(w_dff_A_b9HBXwYE4_0),.din(w_dff_A_Fh9HDm058_0),.clk(gclk));
	jdff dff_A_b9HBXwYE4_0(.dout(w_dff_A_pR7WgH8F8_0),.din(w_dff_A_b9HBXwYE4_0),.clk(gclk));
	jdff dff_A_pR7WgH8F8_0(.dout(w_dff_A_HWlffA8n1_0),.din(w_dff_A_pR7WgH8F8_0),.clk(gclk));
	jdff dff_A_HWlffA8n1_0(.dout(w_dff_A_V2ySCPy10_0),.din(w_dff_A_HWlffA8n1_0),.clk(gclk));
	jdff dff_A_V2ySCPy10_0(.dout(w_dff_A_d1KRSa3g7_0),.din(w_dff_A_V2ySCPy10_0),.clk(gclk));
	jdff dff_A_d1KRSa3g7_0(.dout(w_dff_A_V3pZY9iN1_0),.din(w_dff_A_d1KRSa3g7_0),.clk(gclk));
	jdff dff_A_V3pZY9iN1_0(.dout(f15),.din(w_dff_A_V3pZY9iN1_0),.clk(gclk));
	jdff dff_A_LnRVlKwa4_2(.dout(w_dff_A_GK17Zi180_0),.din(w_dff_A_LnRVlKwa4_2),.clk(gclk));
	jdff dff_A_GK17Zi180_0(.dout(w_dff_A_lW9ue4Dn2_0),.din(w_dff_A_GK17Zi180_0),.clk(gclk));
	jdff dff_A_lW9ue4Dn2_0(.dout(w_dff_A_BE9RXxIO3_0),.din(w_dff_A_lW9ue4Dn2_0),.clk(gclk));
	jdff dff_A_BE9RXxIO3_0(.dout(w_dff_A_ixFFjpir3_0),.din(w_dff_A_BE9RXxIO3_0),.clk(gclk));
	jdff dff_A_ixFFjpir3_0(.dout(w_dff_A_AJc7r0aX4_0),.din(w_dff_A_ixFFjpir3_0),.clk(gclk));
	jdff dff_A_AJc7r0aX4_0(.dout(w_dff_A_uEnheoL41_0),.din(w_dff_A_AJc7r0aX4_0),.clk(gclk));
	jdff dff_A_uEnheoL41_0(.dout(w_dff_A_daE6IegH4_0),.din(w_dff_A_uEnheoL41_0),.clk(gclk));
	jdff dff_A_daE6IegH4_0(.dout(w_dff_A_vpGSQ5t40_0),.din(w_dff_A_daE6IegH4_0),.clk(gclk));
	jdff dff_A_vpGSQ5t40_0(.dout(w_dff_A_06lDjxKk2_0),.din(w_dff_A_vpGSQ5t40_0),.clk(gclk));
	jdff dff_A_06lDjxKk2_0(.dout(w_dff_A_QeflJm1n3_0),.din(w_dff_A_06lDjxKk2_0),.clk(gclk));
	jdff dff_A_QeflJm1n3_0(.dout(w_dff_A_Jz3tUiPJ3_0),.din(w_dff_A_QeflJm1n3_0),.clk(gclk));
	jdff dff_A_Jz3tUiPJ3_0(.dout(w_dff_A_vVpFV9RF8_0),.din(w_dff_A_Jz3tUiPJ3_0),.clk(gclk));
	jdff dff_A_vVpFV9RF8_0(.dout(w_dff_A_iUb9M4Mt3_0),.din(w_dff_A_vVpFV9RF8_0),.clk(gclk));
	jdff dff_A_iUb9M4Mt3_0(.dout(w_dff_A_UpoWBSax6_0),.din(w_dff_A_iUb9M4Mt3_0),.clk(gclk));
	jdff dff_A_UpoWBSax6_0(.dout(w_dff_A_NAlYSviQ2_0),.din(w_dff_A_UpoWBSax6_0),.clk(gclk));
	jdff dff_A_NAlYSviQ2_0(.dout(w_dff_A_DxhC7mnd2_0),.din(w_dff_A_NAlYSviQ2_0),.clk(gclk));
	jdff dff_A_DxhC7mnd2_0(.dout(w_dff_A_cUSAUAH70_0),.din(w_dff_A_DxhC7mnd2_0),.clk(gclk));
	jdff dff_A_cUSAUAH70_0(.dout(w_dff_A_Q9WX1Wb54_0),.din(w_dff_A_cUSAUAH70_0),.clk(gclk));
	jdff dff_A_Q9WX1Wb54_0(.dout(w_dff_A_GfLPjbmh9_0),.din(w_dff_A_Q9WX1Wb54_0),.clk(gclk));
	jdff dff_A_GfLPjbmh9_0(.dout(w_dff_A_gSi30ZFL0_0),.din(w_dff_A_GfLPjbmh9_0),.clk(gclk));
	jdff dff_A_gSi30ZFL0_0(.dout(w_dff_A_BqiiYC0T5_0),.din(w_dff_A_gSi30ZFL0_0),.clk(gclk));
	jdff dff_A_BqiiYC0T5_0(.dout(w_dff_A_YzG78xio8_0),.din(w_dff_A_BqiiYC0T5_0),.clk(gclk));
	jdff dff_A_YzG78xio8_0(.dout(w_dff_A_VLOdgHGE5_0),.din(w_dff_A_YzG78xio8_0),.clk(gclk));
	jdff dff_A_VLOdgHGE5_0(.dout(w_dff_A_dCxFqYyP6_0),.din(w_dff_A_VLOdgHGE5_0),.clk(gclk));
	jdff dff_A_dCxFqYyP6_0(.dout(w_dff_A_BMzsJ6o49_0),.din(w_dff_A_dCxFqYyP6_0),.clk(gclk));
	jdff dff_A_BMzsJ6o49_0(.dout(w_dff_A_gIkgkHOE3_0),.din(w_dff_A_BMzsJ6o49_0),.clk(gclk));
	jdff dff_A_gIkgkHOE3_0(.dout(w_dff_A_38zmTKvG5_0),.din(w_dff_A_gIkgkHOE3_0),.clk(gclk));
	jdff dff_A_38zmTKvG5_0(.dout(w_dff_A_AQbHBeld3_0),.din(w_dff_A_38zmTKvG5_0),.clk(gclk));
	jdff dff_A_AQbHBeld3_0(.dout(w_dff_A_utVQxiDS8_0),.din(w_dff_A_AQbHBeld3_0),.clk(gclk));
	jdff dff_A_utVQxiDS8_0(.dout(w_dff_A_8GKWIRTR2_0),.din(w_dff_A_utVQxiDS8_0),.clk(gclk));
	jdff dff_A_8GKWIRTR2_0(.dout(w_dff_A_JccYcWe10_0),.din(w_dff_A_8GKWIRTR2_0),.clk(gclk));
	jdff dff_A_JccYcWe10_0(.dout(w_dff_A_JFnIfDDo6_0),.din(w_dff_A_JccYcWe10_0),.clk(gclk));
	jdff dff_A_JFnIfDDo6_0(.dout(w_dff_A_0npYbGSR7_0),.din(w_dff_A_JFnIfDDo6_0),.clk(gclk));
	jdff dff_A_0npYbGSR7_0(.dout(w_dff_A_E3ewEzc74_0),.din(w_dff_A_0npYbGSR7_0),.clk(gclk));
	jdff dff_A_E3ewEzc74_0(.dout(w_dff_A_z2wogqZx3_0),.din(w_dff_A_E3ewEzc74_0),.clk(gclk));
	jdff dff_A_z2wogqZx3_0(.dout(w_dff_A_zefGtloA3_0),.din(w_dff_A_z2wogqZx3_0),.clk(gclk));
	jdff dff_A_zefGtloA3_0(.dout(w_dff_A_jxbUBYPm1_0),.din(w_dff_A_zefGtloA3_0),.clk(gclk));
	jdff dff_A_jxbUBYPm1_0(.dout(w_dff_A_qSkxmWZR6_0),.din(w_dff_A_jxbUBYPm1_0),.clk(gclk));
	jdff dff_A_qSkxmWZR6_0(.dout(w_dff_A_RijoFnLp3_0),.din(w_dff_A_qSkxmWZR6_0),.clk(gclk));
	jdff dff_A_RijoFnLp3_0(.dout(w_dff_A_XFr3uI0x3_0),.din(w_dff_A_RijoFnLp3_0),.clk(gclk));
	jdff dff_A_XFr3uI0x3_0(.dout(w_dff_A_crkcGPVa3_0),.din(w_dff_A_XFr3uI0x3_0),.clk(gclk));
	jdff dff_A_crkcGPVa3_0(.dout(w_dff_A_wmX7xsHM9_0),.din(w_dff_A_crkcGPVa3_0),.clk(gclk));
	jdff dff_A_wmX7xsHM9_0(.dout(w_dff_A_6NvJomrV2_0),.din(w_dff_A_wmX7xsHM9_0),.clk(gclk));
	jdff dff_A_6NvJomrV2_0(.dout(w_dff_A_VGtyecpn9_0),.din(w_dff_A_6NvJomrV2_0),.clk(gclk));
	jdff dff_A_VGtyecpn9_0(.dout(w_dff_A_MC0aPK002_0),.din(w_dff_A_VGtyecpn9_0),.clk(gclk));
	jdff dff_A_MC0aPK002_0(.dout(w_dff_A_QsANbYHm3_0),.din(w_dff_A_MC0aPK002_0),.clk(gclk));
	jdff dff_A_QsANbYHm3_0(.dout(w_dff_A_FvPki2c32_0),.din(w_dff_A_QsANbYHm3_0),.clk(gclk));
	jdff dff_A_FvPki2c32_0(.dout(w_dff_A_i3SnkOgy5_0),.din(w_dff_A_FvPki2c32_0),.clk(gclk));
	jdff dff_A_i3SnkOgy5_0(.dout(w_dff_A_MUwsc3Zd2_0),.din(w_dff_A_i3SnkOgy5_0),.clk(gclk));
	jdff dff_A_MUwsc3Zd2_0(.dout(w_dff_A_aQ2v3rbt2_0),.din(w_dff_A_MUwsc3Zd2_0),.clk(gclk));
	jdff dff_A_aQ2v3rbt2_0(.dout(w_dff_A_azkOg4LF7_0),.din(w_dff_A_aQ2v3rbt2_0),.clk(gclk));
	jdff dff_A_azkOg4LF7_0(.dout(w_dff_A_dS4JQigv7_0),.din(w_dff_A_azkOg4LF7_0),.clk(gclk));
	jdff dff_A_dS4JQigv7_0(.dout(w_dff_A_bRfeQZ0Q2_0),.din(w_dff_A_dS4JQigv7_0),.clk(gclk));
	jdff dff_A_bRfeQZ0Q2_0(.dout(w_dff_A_3AuhCwAT9_0),.din(w_dff_A_bRfeQZ0Q2_0),.clk(gclk));
	jdff dff_A_3AuhCwAT9_0(.dout(w_dff_A_2KtKK2LF4_0),.din(w_dff_A_3AuhCwAT9_0),.clk(gclk));
	jdff dff_A_2KtKK2LF4_0(.dout(w_dff_A_mFvcxgRC2_0),.din(w_dff_A_2KtKK2LF4_0),.clk(gclk));
	jdff dff_A_mFvcxgRC2_0(.dout(w_dff_A_Xub2dLhQ8_0),.din(w_dff_A_mFvcxgRC2_0),.clk(gclk));
	jdff dff_A_Xub2dLhQ8_0(.dout(w_dff_A_S9fstQr57_0),.din(w_dff_A_Xub2dLhQ8_0),.clk(gclk));
	jdff dff_A_S9fstQr57_0(.dout(w_dff_A_EbOiH5BD5_0),.din(w_dff_A_S9fstQr57_0),.clk(gclk));
	jdff dff_A_EbOiH5BD5_0(.dout(w_dff_A_DViXWFGQ6_0),.din(w_dff_A_EbOiH5BD5_0),.clk(gclk));
	jdff dff_A_DViXWFGQ6_0(.dout(w_dff_A_N9AWNA2D5_0),.din(w_dff_A_DViXWFGQ6_0),.clk(gclk));
	jdff dff_A_N9AWNA2D5_0(.dout(w_dff_A_xi5hklZm5_0),.din(w_dff_A_N9AWNA2D5_0),.clk(gclk));
	jdff dff_A_xi5hklZm5_0(.dout(w_dff_A_jZbA6zbg0_0),.din(w_dff_A_xi5hklZm5_0),.clk(gclk));
	jdff dff_A_jZbA6zbg0_0(.dout(w_dff_A_sPo61Znb1_0),.din(w_dff_A_jZbA6zbg0_0),.clk(gclk));
	jdff dff_A_sPo61Znb1_0(.dout(w_dff_A_IZ3BHVys4_0),.din(w_dff_A_sPo61Znb1_0),.clk(gclk));
	jdff dff_A_IZ3BHVys4_0(.dout(w_dff_A_fshhcu145_0),.din(w_dff_A_IZ3BHVys4_0),.clk(gclk));
	jdff dff_A_fshhcu145_0(.dout(w_dff_A_o8F1Q50S3_0),.din(w_dff_A_fshhcu145_0),.clk(gclk));
	jdff dff_A_o8F1Q50S3_0(.dout(w_dff_A_azSwqbDW3_0),.din(w_dff_A_o8F1Q50S3_0),.clk(gclk));
	jdff dff_A_azSwqbDW3_0(.dout(w_dff_A_jXDBjFuD2_0),.din(w_dff_A_azSwqbDW3_0),.clk(gclk));
	jdff dff_A_jXDBjFuD2_0(.dout(w_dff_A_9EwgyWNC7_0),.din(w_dff_A_jXDBjFuD2_0),.clk(gclk));
	jdff dff_A_9EwgyWNC7_0(.dout(w_dff_A_gNkFYLLe6_0),.din(w_dff_A_9EwgyWNC7_0),.clk(gclk));
	jdff dff_A_gNkFYLLe6_0(.dout(w_dff_A_Dkc77BML4_0),.din(w_dff_A_gNkFYLLe6_0),.clk(gclk));
	jdff dff_A_Dkc77BML4_0(.dout(w_dff_A_zVH8nU5U0_0),.din(w_dff_A_Dkc77BML4_0),.clk(gclk));
	jdff dff_A_zVH8nU5U0_0(.dout(w_dff_A_MeA5eeRx0_0),.din(w_dff_A_zVH8nU5U0_0),.clk(gclk));
	jdff dff_A_MeA5eeRx0_0(.dout(w_dff_A_TcuLzh6s8_0),.din(w_dff_A_MeA5eeRx0_0),.clk(gclk));
	jdff dff_A_TcuLzh6s8_0(.dout(w_dff_A_nkMtUgND0_0),.din(w_dff_A_TcuLzh6s8_0),.clk(gclk));
	jdff dff_A_nkMtUgND0_0(.dout(w_dff_A_oMBxkO476_0),.din(w_dff_A_nkMtUgND0_0),.clk(gclk));
	jdff dff_A_oMBxkO476_0(.dout(w_dff_A_TYV4Z4B59_0),.din(w_dff_A_oMBxkO476_0),.clk(gclk));
	jdff dff_A_TYV4Z4B59_0(.dout(w_dff_A_M8y88Keo2_0),.din(w_dff_A_TYV4Z4B59_0),.clk(gclk));
	jdff dff_A_M8y88Keo2_0(.dout(w_dff_A_wfUlKs3q1_0),.din(w_dff_A_M8y88Keo2_0),.clk(gclk));
	jdff dff_A_wfUlKs3q1_0(.dout(w_dff_A_Z1NBHCMx2_0),.din(w_dff_A_wfUlKs3q1_0),.clk(gclk));
	jdff dff_A_Z1NBHCMx2_0(.dout(w_dff_A_CBSOZ4se8_0),.din(w_dff_A_Z1NBHCMx2_0),.clk(gclk));
	jdff dff_A_CBSOZ4se8_0(.dout(w_dff_A_CJCdGsZp1_0),.din(w_dff_A_CBSOZ4se8_0),.clk(gclk));
	jdff dff_A_CJCdGsZp1_0(.dout(w_dff_A_yfK9XDiI3_0),.din(w_dff_A_CJCdGsZp1_0),.clk(gclk));
	jdff dff_A_yfK9XDiI3_0(.dout(w_dff_A_xsbLQR2Z2_0),.din(w_dff_A_yfK9XDiI3_0),.clk(gclk));
	jdff dff_A_xsbLQR2Z2_0(.dout(w_dff_A_afvFzpEu6_0),.din(w_dff_A_xsbLQR2Z2_0),.clk(gclk));
	jdff dff_A_afvFzpEu6_0(.dout(w_dff_A_8gKV97629_0),.din(w_dff_A_afvFzpEu6_0),.clk(gclk));
	jdff dff_A_8gKV97629_0(.dout(w_dff_A_4B0Q3ecX3_0),.din(w_dff_A_8gKV97629_0),.clk(gclk));
	jdff dff_A_4B0Q3ecX3_0(.dout(w_dff_A_McgJoamV3_0),.din(w_dff_A_4B0Q3ecX3_0),.clk(gclk));
	jdff dff_A_McgJoamV3_0(.dout(w_dff_A_nWNxZivz4_0),.din(w_dff_A_McgJoamV3_0),.clk(gclk));
	jdff dff_A_nWNxZivz4_0(.dout(w_dff_A_pjIBkap30_0),.din(w_dff_A_nWNxZivz4_0),.clk(gclk));
	jdff dff_A_pjIBkap30_0(.dout(w_dff_A_Tv38rjXd5_0),.din(w_dff_A_pjIBkap30_0),.clk(gclk));
	jdff dff_A_Tv38rjXd5_0(.dout(w_dff_A_BbUfIVL53_0),.din(w_dff_A_Tv38rjXd5_0),.clk(gclk));
	jdff dff_A_BbUfIVL53_0(.dout(w_dff_A_Dpw7lItZ4_0),.din(w_dff_A_BbUfIVL53_0),.clk(gclk));
	jdff dff_A_Dpw7lItZ4_0(.dout(w_dff_A_LvQWLnqK0_0),.din(w_dff_A_Dpw7lItZ4_0),.clk(gclk));
	jdff dff_A_LvQWLnqK0_0(.dout(w_dff_A_pe22L4Xn7_0),.din(w_dff_A_LvQWLnqK0_0),.clk(gclk));
	jdff dff_A_pe22L4Xn7_0(.dout(w_dff_A_cfbyEwWr9_0),.din(w_dff_A_pe22L4Xn7_0),.clk(gclk));
	jdff dff_A_cfbyEwWr9_0(.dout(w_dff_A_VDMuFJSj8_0),.din(w_dff_A_cfbyEwWr9_0),.clk(gclk));
	jdff dff_A_VDMuFJSj8_0(.dout(w_dff_A_pOvi5AFl4_0),.din(w_dff_A_VDMuFJSj8_0),.clk(gclk));
	jdff dff_A_pOvi5AFl4_0(.dout(w_dff_A_aenLQ3jJ3_0),.din(w_dff_A_pOvi5AFl4_0),.clk(gclk));
	jdff dff_A_aenLQ3jJ3_0(.dout(w_dff_A_E53xgmrV7_0),.din(w_dff_A_aenLQ3jJ3_0),.clk(gclk));
	jdff dff_A_E53xgmrV7_0(.dout(w_dff_A_H3iOXkfp6_0),.din(w_dff_A_E53xgmrV7_0),.clk(gclk));
	jdff dff_A_H3iOXkfp6_0(.dout(w_dff_A_gN7IGKPd0_0),.din(w_dff_A_H3iOXkfp6_0),.clk(gclk));
	jdff dff_A_gN7IGKPd0_0(.dout(w_dff_A_Jt9BIdY34_0),.din(w_dff_A_gN7IGKPd0_0),.clk(gclk));
	jdff dff_A_Jt9BIdY34_0(.dout(w_dff_A_eVtOGUf78_0),.din(w_dff_A_Jt9BIdY34_0),.clk(gclk));
	jdff dff_A_eVtOGUf78_0(.dout(w_dff_A_8bU3y6LR7_0),.din(w_dff_A_eVtOGUf78_0),.clk(gclk));
	jdff dff_A_8bU3y6LR7_0(.dout(w_dff_A_WdVxd6TF5_0),.din(w_dff_A_8bU3y6LR7_0),.clk(gclk));
	jdff dff_A_WdVxd6TF5_0(.dout(w_dff_A_TlbkNLvE8_0),.din(w_dff_A_WdVxd6TF5_0),.clk(gclk));
	jdff dff_A_TlbkNLvE8_0(.dout(w_dff_A_XhSVAIJU8_0),.din(w_dff_A_TlbkNLvE8_0),.clk(gclk));
	jdff dff_A_XhSVAIJU8_0(.dout(w_dff_A_bMqwp1pC8_0),.din(w_dff_A_XhSVAIJU8_0),.clk(gclk));
	jdff dff_A_bMqwp1pC8_0(.dout(f16),.din(w_dff_A_bMqwp1pC8_0),.clk(gclk));
	jdff dff_A_xWMjmKJE2_2(.dout(w_dff_A_DkJMFBsl0_0),.din(w_dff_A_xWMjmKJE2_2),.clk(gclk));
	jdff dff_A_DkJMFBsl0_0(.dout(w_dff_A_eRpe2XwF9_0),.din(w_dff_A_DkJMFBsl0_0),.clk(gclk));
	jdff dff_A_eRpe2XwF9_0(.dout(w_dff_A_xYvshyNj1_0),.din(w_dff_A_eRpe2XwF9_0),.clk(gclk));
	jdff dff_A_xYvshyNj1_0(.dout(w_dff_A_7L2wVWA19_0),.din(w_dff_A_xYvshyNj1_0),.clk(gclk));
	jdff dff_A_7L2wVWA19_0(.dout(w_dff_A_ntlnEkbs6_0),.din(w_dff_A_7L2wVWA19_0),.clk(gclk));
	jdff dff_A_ntlnEkbs6_0(.dout(w_dff_A_YhBG0bmk5_0),.din(w_dff_A_ntlnEkbs6_0),.clk(gclk));
	jdff dff_A_YhBG0bmk5_0(.dout(w_dff_A_L9buB5Kh1_0),.din(w_dff_A_YhBG0bmk5_0),.clk(gclk));
	jdff dff_A_L9buB5Kh1_0(.dout(w_dff_A_m7YZYDBO0_0),.din(w_dff_A_L9buB5Kh1_0),.clk(gclk));
	jdff dff_A_m7YZYDBO0_0(.dout(w_dff_A_mdTfVhnM0_0),.din(w_dff_A_m7YZYDBO0_0),.clk(gclk));
	jdff dff_A_mdTfVhnM0_0(.dout(w_dff_A_dGB1DOfZ8_0),.din(w_dff_A_mdTfVhnM0_0),.clk(gclk));
	jdff dff_A_dGB1DOfZ8_0(.dout(w_dff_A_j7Jxdgcg1_0),.din(w_dff_A_dGB1DOfZ8_0),.clk(gclk));
	jdff dff_A_j7Jxdgcg1_0(.dout(w_dff_A_VsohchKp2_0),.din(w_dff_A_j7Jxdgcg1_0),.clk(gclk));
	jdff dff_A_VsohchKp2_0(.dout(w_dff_A_nm58TXz85_0),.din(w_dff_A_VsohchKp2_0),.clk(gclk));
	jdff dff_A_nm58TXz85_0(.dout(w_dff_A_6V0Sn0jg2_0),.din(w_dff_A_nm58TXz85_0),.clk(gclk));
	jdff dff_A_6V0Sn0jg2_0(.dout(w_dff_A_yTKuAOOy3_0),.din(w_dff_A_6V0Sn0jg2_0),.clk(gclk));
	jdff dff_A_yTKuAOOy3_0(.dout(w_dff_A_YuarT5dq3_0),.din(w_dff_A_yTKuAOOy3_0),.clk(gclk));
	jdff dff_A_YuarT5dq3_0(.dout(w_dff_A_ypgxAohj8_0),.din(w_dff_A_YuarT5dq3_0),.clk(gclk));
	jdff dff_A_ypgxAohj8_0(.dout(w_dff_A_Cj4NbuNv3_0),.din(w_dff_A_ypgxAohj8_0),.clk(gclk));
	jdff dff_A_Cj4NbuNv3_0(.dout(w_dff_A_obf4KN2F3_0),.din(w_dff_A_Cj4NbuNv3_0),.clk(gclk));
	jdff dff_A_obf4KN2F3_0(.dout(w_dff_A_DepMQ3AP1_0),.din(w_dff_A_obf4KN2F3_0),.clk(gclk));
	jdff dff_A_DepMQ3AP1_0(.dout(w_dff_A_54Ip8c1M8_0),.din(w_dff_A_DepMQ3AP1_0),.clk(gclk));
	jdff dff_A_54Ip8c1M8_0(.dout(w_dff_A_VafUtmqL6_0),.din(w_dff_A_54Ip8c1M8_0),.clk(gclk));
	jdff dff_A_VafUtmqL6_0(.dout(w_dff_A_EwmlLQ6J8_0),.din(w_dff_A_VafUtmqL6_0),.clk(gclk));
	jdff dff_A_EwmlLQ6J8_0(.dout(w_dff_A_OMJ54ela6_0),.din(w_dff_A_EwmlLQ6J8_0),.clk(gclk));
	jdff dff_A_OMJ54ela6_0(.dout(w_dff_A_dmZJhJio1_0),.din(w_dff_A_OMJ54ela6_0),.clk(gclk));
	jdff dff_A_dmZJhJio1_0(.dout(w_dff_A_MTfHFV5n7_0),.din(w_dff_A_dmZJhJio1_0),.clk(gclk));
	jdff dff_A_MTfHFV5n7_0(.dout(w_dff_A_HYYEK37L1_0),.din(w_dff_A_MTfHFV5n7_0),.clk(gclk));
	jdff dff_A_HYYEK37L1_0(.dout(w_dff_A_vQ5WQZWB1_0),.din(w_dff_A_HYYEK37L1_0),.clk(gclk));
	jdff dff_A_vQ5WQZWB1_0(.dout(w_dff_A_rerBWFOs2_0),.din(w_dff_A_vQ5WQZWB1_0),.clk(gclk));
	jdff dff_A_rerBWFOs2_0(.dout(w_dff_A_JTqmsg9W8_0),.din(w_dff_A_rerBWFOs2_0),.clk(gclk));
	jdff dff_A_JTqmsg9W8_0(.dout(w_dff_A_olKsJiUt0_0),.din(w_dff_A_JTqmsg9W8_0),.clk(gclk));
	jdff dff_A_olKsJiUt0_0(.dout(w_dff_A_zhWekP025_0),.din(w_dff_A_olKsJiUt0_0),.clk(gclk));
	jdff dff_A_zhWekP025_0(.dout(w_dff_A_Xo1T2vJN0_0),.din(w_dff_A_zhWekP025_0),.clk(gclk));
	jdff dff_A_Xo1T2vJN0_0(.dout(w_dff_A_IUeXKzG53_0),.din(w_dff_A_Xo1T2vJN0_0),.clk(gclk));
	jdff dff_A_IUeXKzG53_0(.dout(w_dff_A_bWo59w982_0),.din(w_dff_A_IUeXKzG53_0),.clk(gclk));
	jdff dff_A_bWo59w982_0(.dout(w_dff_A_V6IQTE7s5_0),.din(w_dff_A_bWo59w982_0),.clk(gclk));
	jdff dff_A_V6IQTE7s5_0(.dout(w_dff_A_d29VOzQS2_0),.din(w_dff_A_V6IQTE7s5_0),.clk(gclk));
	jdff dff_A_d29VOzQS2_0(.dout(w_dff_A_g0NGThwQ6_0),.din(w_dff_A_d29VOzQS2_0),.clk(gclk));
	jdff dff_A_g0NGThwQ6_0(.dout(w_dff_A_5IJPJmME5_0),.din(w_dff_A_g0NGThwQ6_0),.clk(gclk));
	jdff dff_A_5IJPJmME5_0(.dout(w_dff_A_n3zITi9s8_0),.din(w_dff_A_5IJPJmME5_0),.clk(gclk));
	jdff dff_A_n3zITi9s8_0(.dout(w_dff_A_NG8jV5401_0),.din(w_dff_A_n3zITi9s8_0),.clk(gclk));
	jdff dff_A_NG8jV5401_0(.dout(w_dff_A_bm2zZj0w4_0),.din(w_dff_A_NG8jV5401_0),.clk(gclk));
	jdff dff_A_bm2zZj0w4_0(.dout(w_dff_A_sbe9cv5T4_0),.din(w_dff_A_bm2zZj0w4_0),.clk(gclk));
	jdff dff_A_sbe9cv5T4_0(.dout(w_dff_A_WuyrlZ9q5_0),.din(w_dff_A_sbe9cv5T4_0),.clk(gclk));
	jdff dff_A_WuyrlZ9q5_0(.dout(w_dff_A_NnwocXyi6_0),.din(w_dff_A_WuyrlZ9q5_0),.clk(gclk));
	jdff dff_A_NnwocXyi6_0(.dout(w_dff_A_U5PCJfn73_0),.din(w_dff_A_NnwocXyi6_0),.clk(gclk));
	jdff dff_A_U5PCJfn73_0(.dout(w_dff_A_YM0Hm7P92_0),.din(w_dff_A_U5PCJfn73_0),.clk(gclk));
	jdff dff_A_YM0Hm7P92_0(.dout(w_dff_A_pzdTgPyN8_0),.din(w_dff_A_YM0Hm7P92_0),.clk(gclk));
	jdff dff_A_pzdTgPyN8_0(.dout(w_dff_A_5p6oRS8A0_0),.din(w_dff_A_pzdTgPyN8_0),.clk(gclk));
	jdff dff_A_5p6oRS8A0_0(.dout(w_dff_A_ozu1WvW45_0),.din(w_dff_A_5p6oRS8A0_0),.clk(gclk));
	jdff dff_A_ozu1WvW45_0(.dout(w_dff_A_DvLvGVYE7_0),.din(w_dff_A_ozu1WvW45_0),.clk(gclk));
	jdff dff_A_DvLvGVYE7_0(.dout(w_dff_A_kw1oR4ST3_0),.din(w_dff_A_DvLvGVYE7_0),.clk(gclk));
	jdff dff_A_kw1oR4ST3_0(.dout(w_dff_A_0NnmIXzU9_0),.din(w_dff_A_kw1oR4ST3_0),.clk(gclk));
	jdff dff_A_0NnmIXzU9_0(.dout(w_dff_A_oVjXKx4p9_0),.din(w_dff_A_0NnmIXzU9_0),.clk(gclk));
	jdff dff_A_oVjXKx4p9_0(.dout(w_dff_A_X3R2WtyE0_0),.din(w_dff_A_oVjXKx4p9_0),.clk(gclk));
	jdff dff_A_X3R2WtyE0_0(.dout(w_dff_A_Ir5YRAR96_0),.din(w_dff_A_X3R2WtyE0_0),.clk(gclk));
	jdff dff_A_Ir5YRAR96_0(.dout(w_dff_A_02kA5U2F1_0),.din(w_dff_A_Ir5YRAR96_0),.clk(gclk));
	jdff dff_A_02kA5U2F1_0(.dout(w_dff_A_Z5HPi5Ou3_0),.din(w_dff_A_02kA5U2F1_0),.clk(gclk));
	jdff dff_A_Z5HPi5Ou3_0(.dout(w_dff_A_FDiGOMEP9_0),.din(w_dff_A_Z5HPi5Ou3_0),.clk(gclk));
	jdff dff_A_FDiGOMEP9_0(.dout(w_dff_A_ElnAZ9DI8_0),.din(w_dff_A_FDiGOMEP9_0),.clk(gclk));
	jdff dff_A_ElnAZ9DI8_0(.dout(w_dff_A_By2I0aJz1_0),.din(w_dff_A_ElnAZ9DI8_0),.clk(gclk));
	jdff dff_A_By2I0aJz1_0(.dout(w_dff_A_PASuZudb7_0),.din(w_dff_A_By2I0aJz1_0),.clk(gclk));
	jdff dff_A_PASuZudb7_0(.dout(w_dff_A_E3JSNpSC3_0),.din(w_dff_A_PASuZudb7_0),.clk(gclk));
	jdff dff_A_E3JSNpSC3_0(.dout(w_dff_A_5bCIY7b58_0),.din(w_dff_A_E3JSNpSC3_0),.clk(gclk));
	jdff dff_A_5bCIY7b58_0(.dout(w_dff_A_ZoejADoS4_0),.din(w_dff_A_5bCIY7b58_0),.clk(gclk));
	jdff dff_A_ZoejADoS4_0(.dout(w_dff_A_8DNFPTKt0_0),.din(w_dff_A_ZoejADoS4_0),.clk(gclk));
	jdff dff_A_8DNFPTKt0_0(.dout(w_dff_A_jnB6bsRC0_0),.din(w_dff_A_8DNFPTKt0_0),.clk(gclk));
	jdff dff_A_jnB6bsRC0_0(.dout(w_dff_A_sbXDQhRO6_0),.din(w_dff_A_jnB6bsRC0_0),.clk(gclk));
	jdff dff_A_sbXDQhRO6_0(.dout(w_dff_A_oFQ072T27_0),.din(w_dff_A_sbXDQhRO6_0),.clk(gclk));
	jdff dff_A_oFQ072T27_0(.dout(w_dff_A_bLN9Z6Uf8_0),.din(w_dff_A_oFQ072T27_0),.clk(gclk));
	jdff dff_A_bLN9Z6Uf8_0(.dout(w_dff_A_zjLxCi0u5_0),.din(w_dff_A_bLN9Z6Uf8_0),.clk(gclk));
	jdff dff_A_zjLxCi0u5_0(.dout(w_dff_A_r9vIrRWV2_0),.din(w_dff_A_zjLxCi0u5_0),.clk(gclk));
	jdff dff_A_r9vIrRWV2_0(.dout(w_dff_A_zPvoC2co9_0),.din(w_dff_A_r9vIrRWV2_0),.clk(gclk));
	jdff dff_A_zPvoC2co9_0(.dout(w_dff_A_lVeMbgJN4_0),.din(w_dff_A_zPvoC2co9_0),.clk(gclk));
	jdff dff_A_lVeMbgJN4_0(.dout(w_dff_A_XvciFmFD8_0),.din(w_dff_A_lVeMbgJN4_0),.clk(gclk));
	jdff dff_A_XvciFmFD8_0(.dout(w_dff_A_lPrlWIuJ9_0),.din(w_dff_A_XvciFmFD8_0),.clk(gclk));
	jdff dff_A_lPrlWIuJ9_0(.dout(w_dff_A_IasE0Rks4_0),.din(w_dff_A_lPrlWIuJ9_0),.clk(gclk));
	jdff dff_A_IasE0Rks4_0(.dout(w_dff_A_VWjgA6Ef2_0),.din(w_dff_A_IasE0Rks4_0),.clk(gclk));
	jdff dff_A_VWjgA6Ef2_0(.dout(w_dff_A_DbaijFgF9_0),.din(w_dff_A_VWjgA6Ef2_0),.clk(gclk));
	jdff dff_A_DbaijFgF9_0(.dout(w_dff_A_H6dru41O1_0),.din(w_dff_A_DbaijFgF9_0),.clk(gclk));
	jdff dff_A_H6dru41O1_0(.dout(w_dff_A_3GNLmASH0_0),.din(w_dff_A_H6dru41O1_0),.clk(gclk));
	jdff dff_A_3GNLmASH0_0(.dout(w_dff_A_Q2SslOAA9_0),.din(w_dff_A_3GNLmASH0_0),.clk(gclk));
	jdff dff_A_Q2SslOAA9_0(.dout(w_dff_A_vKmCJMEw4_0),.din(w_dff_A_Q2SslOAA9_0),.clk(gclk));
	jdff dff_A_vKmCJMEw4_0(.dout(w_dff_A_q8dPJcMt0_0),.din(w_dff_A_vKmCJMEw4_0),.clk(gclk));
	jdff dff_A_q8dPJcMt0_0(.dout(w_dff_A_OvWTKkgz4_0),.din(w_dff_A_q8dPJcMt0_0),.clk(gclk));
	jdff dff_A_OvWTKkgz4_0(.dout(w_dff_A_WTyIX9jb5_0),.din(w_dff_A_OvWTKkgz4_0),.clk(gclk));
	jdff dff_A_WTyIX9jb5_0(.dout(w_dff_A_OADpagla0_0),.din(w_dff_A_WTyIX9jb5_0),.clk(gclk));
	jdff dff_A_OADpagla0_0(.dout(w_dff_A_FUwEQ77B5_0),.din(w_dff_A_OADpagla0_0),.clk(gclk));
	jdff dff_A_FUwEQ77B5_0(.dout(w_dff_A_pX6Q9gKC1_0),.din(w_dff_A_FUwEQ77B5_0),.clk(gclk));
	jdff dff_A_pX6Q9gKC1_0(.dout(w_dff_A_Gjdp805S9_0),.din(w_dff_A_pX6Q9gKC1_0),.clk(gclk));
	jdff dff_A_Gjdp805S9_0(.dout(w_dff_A_LniBg7fT7_0),.din(w_dff_A_Gjdp805S9_0),.clk(gclk));
	jdff dff_A_LniBg7fT7_0(.dout(w_dff_A_JaJrjXgB0_0),.din(w_dff_A_LniBg7fT7_0),.clk(gclk));
	jdff dff_A_JaJrjXgB0_0(.dout(w_dff_A_qF9wrIKC8_0),.din(w_dff_A_JaJrjXgB0_0),.clk(gclk));
	jdff dff_A_qF9wrIKC8_0(.dout(w_dff_A_kEawaRxa6_0),.din(w_dff_A_qF9wrIKC8_0),.clk(gclk));
	jdff dff_A_kEawaRxa6_0(.dout(w_dff_A_XZr9GQfw1_0),.din(w_dff_A_kEawaRxa6_0),.clk(gclk));
	jdff dff_A_XZr9GQfw1_0(.dout(w_dff_A_jpdcxZII7_0),.din(w_dff_A_XZr9GQfw1_0),.clk(gclk));
	jdff dff_A_jpdcxZII7_0(.dout(w_dff_A_rqyXRseC1_0),.din(w_dff_A_jpdcxZII7_0),.clk(gclk));
	jdff dff_A_rqyXRseC1_0(.dout(w_dff_A_EVc1WssU0_0),.din(w_dff_A_rqyXRseC1_0),.clk(gclk));
	jdff dff_A_EVc1WssU0_0(.dout(w_dff_A_PmvkQFem2_0),.din(w_dff_A_EVc1WssU0_0),.clk(gclk));
	jdff dff_A_PmvkQFem2_0(.dout(w_dff_A_9qVp0lul8_0),.din(w_dff_A_PmvkQFem2_0),.clk(gclk));
	jdff dff_A_9qVp0lul8_0(.dout(w_dff_A_WgOfwrNZ0_0),.din(w_dff_A_9qVp0lul8_0),.clk(gclk));
	jdff dff_A_WgOfwrNZ0_0(.dout(w_dff_A_EhHxeAZK8_0),.din(w_dff_A_WgOfwrNZ0_0),.clk(gclk));
	jdff dff_A_EhHxeAZK8_0(.dout(w_dff_A_25Va3Ja75_0),.din(w_dff_A_EhHxeAZK8_0),.clk(gclk));
	jdff dff_A_25Va3Ja75_0(.dout(w_dff_A_Awe5Cts26_0),.din(w_dff_A_25Va3Ja75_0),.clk(gclk));
	jdff dff_A_Awe5Cts26_0(.dout(w_dff_A_uNrlZAZy5_0),.din(w_dff_A_Awe5Cts26_0),.clk(gclk));
	jdff dff_A_uNrlZAZy5_0(.dout(w_dff_A_qWAggIwb1_0),.din(w_dff_A_uNrlZAZy5_0),.clk(gclk));
	jdff dff_A_qWAggIwb1_0(.dout(w_dff_A_UxmRffia0_0),.din(w_dff_A_qWAggIwb1_0),.clk(gclk));
	jdff dff_A_UxmRffia0_0(.dout(w_dff_A_v0QMzmHJ8_0),.din(w_dff_A_UxmRffia0_0),.clk(gclk));
	jdff dff_A_v0QMzmHJ8_0(.dout(w_dff_A_1VMuFBuy4_0),.din(w_dff_A_v0QMzmHJ8_0),.clk(gclk));
	jdff dff_A_1VMuFBuy4_0(.dout(f17),.din(w_dff_A_1VMuFBuy4_0),.clk(gclk));
	jdff dff_A_0NVR8Dal9_2(.dout(w_dff_A_TOmvvoze0_0),.din(w_dff_A_0NVR8Dal9_2),.clk(gclk));
	jdff dff_A_TOmvvoze0_0(.dout(w_dff_A_TJfhYb0O1_0),.din(w_dff_A_TOmvvoze0_0),.clk(gclk));
	jdff dff_A_TJfhYb0O1_0(.dout(w_dff_A_40TqYhct7_0),.din(w_dff_A_TJfhYb0O1_0),.clk(gclk));
	jdff dff_A_40TqYhct7_0(.dout(w_dff_A_Skvnf2ON2_0),.din(w_dff_A_40TqYhct7_0),.clk(gclk));
	jdff dff_A_Skvnf2ON2_0(.dout(w_dff_A_nO7DapF13_0),.din(w_dff_A_Skvnf2ON2_0),.clk(gclk));
	jdff dff_A_nO7DapF13_0(.dout(w_dff_A_8SgC1x9o9_0),.din(w_dff_A_nO7DapF13_0),.clk(gclk));
	jdff dff_A_8SgC1x9o9_0(.dout(w_dff_A_XFjIpT4g5_0),.din(w_dff_A_8SgC1x9o9_0),.clk(gclk));
	jdff dff_A_XFjIpT4g5_0(.dout(w_dff_A_CHOiVaJH3_0),.din(w_dff_A_XFjIpT4g5_0),.clk(gclk));
	jdff dff_A_CHOiVaJH3_0(.dout(w_dff_A_EQ8jbN8w5_0),.din(w_dff_A_CHOiVaJH3_0),.clk(gclk));
	jdff dff_A_EQ8jbN8w5_0(.dout(w_dff_A_P37psMpY6_0),.din(w_dff_A_EQ8jbN8w5_0),.clk(gclk));
	jdff dff_A_P37psMpY6_0(.dout(w_dff_A_753iWZkq8_0),.din(w_dff_A_P37psMpY6_0),.clk(gclk));
	jdff dff_A_753iWZkq8_0(.dout(w_dff_A_Ary1l48t2_0),.din(w_dff_A_753iWZkq8_0),.clk(gclk));
	jdff dff_A_Ary1l48t2_0(.dout(w_dff_A_feVFlSEw9_0),.din(w_dff_A_Ary1l48t2_0),.clk(gclk));
	jdff dff_A_feVFlSEw9_0(.dout(w_dff_A_ISOWXJsA6_0),.din(w_dff_A_feVFlSEw9_0),.clk(gclk));
	jdff dff_A_ISOWXJsA6_0(.dout(w_dff_A_GHdujyMQ9_0),.din(w_dff_A_ISOWXJsA6_0),.clk(gclk));
	jdff dff_A_GHdujyMQ9_0(.dout(w_dff_A_96SLxyII2_0),.din(w_dff_A_GHdujyMQ9_0),.clk(gclk));
	jdff dff_A_96SLxyII2_0(.dout(w_dff_A_GjciuaJ36_0),.din(w_dff_A_96SLxyII2_0),.clk(gclk));
	jdff dff_A_GjciuaJ36_0(.dout(w_dff_A_3l9Pyy6i2_0),.din(w_dff_A_GjciuaJ36_0),.clk(gclk));
	jdff dff_A_3l9Pyy6i2_0(.dout(w_dff_A_hyth8iQW3_0),.din(w_dff_A_3l9Pyy6i2_0),.clk(gclk));
	jdff dff_A_hyth8iQW3_0(.dout(w_dff_A_5oR0vOOk1_0),.din(w_dff_A_hyth8iQW3_0),.clk(gclk));
	jdff dff_A_5oR0vOOk1_0(.dout(w_dff_A_nV2GqiOP5_0),.din(w_dff_A_5oR0vOOk1_0),.clk(gclk));
	jdff dff_A_nV2GqiOP5_0(.dout(w_dff_A_hzttibKQ1_0),.din(w_dff_A_nV2GqiOP5_0),.clk(gclk));
	jdff dff_A_hzttibKQ1_0(.dout(w_dff_A_imLKk0GV8_0),.din(w_dff_A_hzttibKQ1_0),.clk(gclk));
	jdff dff_A_imLKk0GV8_0(.dout(w_dff_A_VVAacT5S3_0),.din(w_dff_A_imLKk0GV8_0),.clk(gclk));
	jdff dff_A_VVAacT5S3_0(.dout(w_dff_A_vhxvB4Ou2_0),.din(w_dff_A_VVAacT5S3_0),.clk(gclk));
	jdff dff_A_vhxvB4Ou2_0(.dout(w_dff_A_sDNlSzfV3_0),.din(w_dff_A_vhxvB4Ou2_0),.clk(gclk));
	jdff dff_A_sDNlSzfV3_0(.dout(w_dff_A_elwENFas5_0),.din(w_dff_A_sDNlSzfV3_0),.clk(gclk));
	jdff dff_A_elwENFas5_0(.dout(w_dff_A_NPrINVDs1_0),.din(w_dff_A_elwENFas5_0),.clk(gclk));
	jdff dff_A_NPrINVDs1_0(.dout(w_dff_A_pmABDIji3_0),.din(w_dff_A_NPrINVDs1_0),.clk(gclk));
	jdff dff_A_pmABDIji3_0(.dout(w_dff_A_liuXLDjP6_0),.din(w_dff_A_pmABDIji3_0),.clk(gclk));
	jdff dff_A_liuXLDjP6_0(.dout(w_dff_A_BdY8vhzM2_0),.din(w_dff_A_liuXLDjP6_0),.clk(gclk));
	jdff dff_A_BdY8vhzM2_0(.dout(w_dff_A_PyFFHFsP3_0),.din(w_dff_A_BdY8vhzM2_0),.clk(gclk));
	jdff dff_A_PyFFHFsP3_0(.dout(w_dff_A_7fXEossO1_0),.din(w_dff_A_PyFFHFsP3_0),.clk(gclk));
	jdff dff_A_7fXEossO1_0(.dout(w_dff_A_pIAhj8wx5_0),.din(w_dff_A_7fXEossO1_0),.clk(gclk));
	jdff dff_A_pIAhj8wx5_0(.dout(w_dff_A_RlDydzZl0_0),.din(w_dff_A_pIAhj8wx5_0),.clk(gclk));
	jdff dff_A_RlDydzZl0_0(.dout(w_dff_A_KS40lmps3_0),.din(w_dff_A_RlDydzZl0_0),.clk(gclk));
	jdff dff_A_KS40lmps3_0(.dout(w_dff_A_lCu3HYrF7_0),.din(w_dff_A_KS40lmps3_0),.clk(gclk));
	jdff dff_A_lCu3HYrF7_0(.dout(w_dff_A_RboOhAq06_0),.din(w_dff_A_lCu3HYrF7_0),.clk(gclk));
	jdff dff_A_RboOhAq06_0(.dout(w_dff_A_lJOf4rp12_0),.din(w_dff_A_RboOhAq06_0),.clk(gclk));
	jdff dff_A_lJOf4rp12_0(.dout(w_dff_A_ay8oj7dI7_0),.din(w_dff_A_lJOf4rp12_0),.clk(gclk));
	jdff dff_A_ay8oj7dI7_0(.dout(w_dff_A_1lKNpT6U8_0),.din(w_dff_A_ay8oj7dI7_0),.clk(gclk));
	jdff dff_A_1lKNpT6U8_0(.dout(w_dff_A_Zgo8m8nF6_0),.din(w_dff_A_1lKNpT6U8_0),.clk(gclk));
	jdff dff_A_Zgo8m8nF6_0(.dout(w_dff_A_WlivYmsQ1_0),.din(w_dff_A_Zgo8m8nF6_0),.clk(gclk));
	jdff dff_A_WlivYmsQ1_0(.dout(w_dff_A_rWIXssFJ6_0),.din(w_dff_A_WlivYmsQ1_0),.clk(gclk));
	jdff dff_A_rWIXssFJ6_0(.dout(w_dff_A_O5Joij324_0),.din(w_dff_A_rWIXssFJ6_0),.clk(gclk));
	jdff dff_A_O5Joij324_0(.dout(w_dff_A_joFGlk3w6_0),.din(w_dff_A_O5Joij324_0),.clk(gclk));
	jdff dff_A_joFGlk3w6_0(.dout(w_dff_A_D4Z40p0y1_0),.din(w_dff_A_joFGlk3w6_0),.clk(gclk));
	jdff dff_A_D4Z40p0y1_0(.dout(w_dff_A_bVLZghZy9_0),.din(w_dff_A_D4Z40p0y1_0),.clk(gclk));
	jdff dff_A_bVLZghZy9_0(.dout(w_dff_A_NNAFmcZQ7_0),.din(w_dff_A_bVLZghZy9_0),.clk(gclk));
	jdff dff_A_NNAFmcZQ7_0(.dout(w_dff_A_orrABZaF8_0),.din(w_dff_A_NNAFmcZQ7_0),.clk(gclk));
	jdff dff_A_orrABZaF8_0(.dout(w_dff_A_Z6bh4OCV3_0),.din(w_dff_A_orrABZaF8_0),.clk(gclk));
	jdff dff_A_Z6bh4OCV3_0(.dout(w_dff_A_rMCwQX3i9_0),.din(w_dff_A_Z6bh4OCV3_0),.clk(gclk));
	jdff dff_A_rMCwQX3i9_0(.dout(w_dff_A_W8z0B9583_0),.din(w_dff_A_rMCwQX3i9_0),.clk(gclk));
	jdff dff_A_W8z0B9583_0(.dout(w_dff_A_6jgMqxPI5_0),.din(w_dff_A_W8z0B9583_0),.clk(gclk));
	jdff dff_A_6jgMqxPI5_0(.dout(w_dff_A_if9xx1hj8_0),.din(w_dff_A_6jgMqxPI5_0),.clk(gclk));
	jdff dff_A_if9xx1hj8_0(.dout(w_dff_A_u5eysuuu2_0),.din(w_dff_A_if9xx1hj8_0),.clk(gclk));
	jdff dff_A_u5eysuuu2_0(.dout(w_dff_A_o4m5kJR06_0),.din(w_dff_A_u5eysuuu2_0),.clk(gclk));
	jdff dff_A_o4m5kJR06_0(.dout(w_dff_A_2UwW5H9A9_0),.din(w_dff_A_o4m5kJR06_0),.clk(gclk));
	jdff dff_A_2UwW5H9A9_0(.dout(w_dff_A_V5watVz60_0),.din(w_dff_A_2UwW5H9A9_0),.clk(gclk));
	jdff dff_A_V5watVz60_0(.dout(w_dff_A_VZO3lMIw3_0),.din(w_dff_A_V5watVz60_0),.clk(gclk));
	jdff dff_A_VZO3lMIw3_0(.dout(w_dff_A_ItVFv0Rj3_0),.din(w_dff_A_VZO3lMIw3_0),.clk(gclk));
	jdff dff_A_ItVFv0Rj3_0(.dout(w_dff_A_3yisev2b6_0),.din(w_dff_A_ItVFv0Rj3_0),.clk(gclk));
	jdff dff_A_3yisev2b6_0(.dout(w_dff_A_KBTOBMpK8_0),.din(w_dff_A_3yisev2b6_0),.clk(gclk));
	jdff dff_A_KBTOBMpK8_0(.dout(w_dff_A_c9kv7l3X8_0),.din(w_dff_A_KBTOBMpK8_0),.clk(gclk));
	jdff dff_A_c9kv7l3X8_0(.dout(w_dff_A_ubitWyl53_0),.din(w_dff_A_c9kv7l3X8_0),.clk(gclk));
	jdff dff_A_ubitWyl53_0(.dout(w_dff_A_O8refhWl5_0),.din(w_dff_A_ubitWyl53_0),.clk(gclk));
	jdff dff_A_O8refhWl5_0(.dout(w_dff_A_EIX1avql9_0),.din(w_dff_A_O8refhWl5_0),.clk(gclk));
	jdff dff_A_EIX1avql9_0(.dout(w_dff_A_xfh00RZ62_0),.din(w_dff_A_EIX1avql9_0),.clk(gclk));
	jdff dff_A_xfh00RZ62_0(.dout(w_dff_A_oK5ygvzo9_0),.din(w_dff_A_xfh00RZ62_0),.clk(gclk));
	jdff dff_A_oK5ygvzo9_0(.dout(w_dff_A_7v9Wf43s3_0),.din(w_dff_A_oK5ygvzo9_0),.clk(gclk));
	jdff dff_A_7v9Wf43s3_0(.dout(w_dff_A_zAzllwME4_0),.din(w_dff_A_7v9Wf43s3_0),.clk(gclk));
	jdff dff_A_zAzllwME4_0(.dout(w_dff_A_Z4izq7vp3_0),.din(w_dff_A_zAzllwME4_0),.clk(gclk));
	jdff dff_A_Z4izq7vp3_0(.dout(w_dff_A_zQu47Bh95_0),.din(w_dff_A_Z4izq7vp3_0),.clk(gclk));
	jdff dff_A_zQu47Bh95_0(.dout(w_dff_A_SdGxpUpS2_0),.din(w_dff_A_zQu47Bh95_0),.clk(gclk));
	jdff dff_A_SdGxpUpS2_0(.dout(w_dff_A_QumTBtFd0_0),.din(w_dff_A_SdGxpUpS2_0),.clk(gclk));
	jdff dff_A_QumTBtFd0_0(.dout(w_dff_A_Y61zjZ820_0),.din(w_dff_A_QumTBtFd0_0),.clk(gclk));
	jdff dff_A_Y61zjZ820_0(.dout(w_dff_A_TWfwnIWv2_0),.din(w_dff_A_Y61zjZ820_0),.clk(gclk));
	jdff dff_A_TWfwnIWv2_0(.dout(w_dff_A_HMKdSwET0_0),.din(w_dff_A_TWfwnIWv2_0),.clk(gclk));
	jdff dff_A_HMKdSwET0_0(.dout(w_dff_A_vx4Y2RsJ8_0),.din(w_dff_A_HMKdSwET0_0),.clk(gclk));
	jdff dff_A_vx4Y2RsJ8_0(.dout(w_dff_A_AQ955nqT1_0),.din(w_dff_A_vx4Y2RsJ8_0),.clk(gclk));
	jdff dff_A_AQ955nqT1_0(.dout(w_dff_A_srhVHj253_0),.din(w_dff_A_AQ955nqT1_0),.clk(gclk));
	jdff dff_A_srhVHj253_0(.dout(w_dff_A_hbHulm8i7_0),.din(w_dff_A_srhVHj253_0),.clk(gclk));
	jdff dff_A_hbHulm8i7_0(.dout(w_dff_A_c55O5gyO6_0),.din(w_dff_A_hbHulm8i7_0),.clk(gclk));
	jdff dff_A_c55O5gyO6_0(.dout(w_dff_A_Cg7tF7AY1_0),.din(w_dff_A_c55O5gyO6_0),.clk(gclk));
	jdff dff_A_Cg7tF7AY1_0(.dout(w_dff_A_KgTGfBXg1_0),.din(w_dff_A_Cg7tF7AY1_0),.clk(gclk));
	jdff dff_A_KgTGfBXg1_0(.dout(w_dff_A_5orPkeyk6_0),.din(w_dff_A_KgTGfBXg1_0),.clk(gclk));
	jdff dff_A_5orPkeyk6_0(.dout(w_dff_A_AReFv5yH3_0),.din(w_dff_A_5orPkeyk6_0),.clk(gclk));
	jdff dff_A_AReFv5yH3_0(.dout(w_dff_A_UD8aM2XE4_0),.din(w_dff_A_AReFv5yH3_0),.clk(gclk));
	jdff dff_A_UD8aM2XE4_0(.dout(w_dff_A_4jtmBBXC2_0),.din(w_dff_A_UD8aM2XE4_0),.clk(gclk));
	jdff dff_A_4jtmBBXC2_0(.dout(w_dff_A_oXPoMipA6_0),.din(w_dff_A_4jtmBBXC2_0),.clk(gclk));
	jdff dff_A_oXPoMipA6_0(.dout(w_dff_A_Axfa65bU2_0),.din(w_dff_A_oXPoMipA6_0),.clk(gclk));
	jdff dff_A_Axfa65bU2_0(.dout(w_dff_A_WsrByzpk8_0),.din(w_dff_A_Axfa65bU2_0),.clk(gclk));
	jdff dff_A_WsrByzpk8_0(.dout(w_dff_A_uDueegk10_0),.din(w_dff_A_WsrByzpk8_0),.clk(gclk));
	jdff dff_A_uDueegk10_0(.dout(w_dff_A_lpwNtV4M6_0),.din(w_dff_A_uDueegk10_0),.clk(gclk));
	jdff dff_A_lpwNtV4M6_0(.dout(w_dff_A_aK4I4rg72_0),.din(w_dff_A_lpwNtV4M6_0),.clk(gclk));
	jdff dff_A_aK4I4rg72_0(.dout(w_dff_A_ujGyJ2Zj2_0),.din(w_dff_A_aK4I4rg72_0),.clk(gclk));
	jdff dff_A_ujGyJ2Zj2_0(.dout(w_dff_A_r8ob65RH6_0),.din(w_dff_A_ujGyJ2Zj2_0),.clk(gclk));
	jdff dff_A_r8ob65RH6_0(.dout(w_dff_A_TlFtjFoC9_0),.din(w_dff_A_r8ob65RH6_0),.clk(gclk));
	jdff dff_A_TlFtjFoC9_0(.dout(w_dff_A_LxbOVs2i8_0),.din(w_dff_A_TlFtjFoC9_0),.clk(gclk));
	jdff dff_A_LxbOVs2i8_0(.dout(w_dff_A_2JmFVYJO4_0),.din(w_dff_A_LxbOVs2i8_0),.clk(gclk));
	jdff dff_A_2JmFVYJO4_0(.dout(w_dff_A_WcGcB9Zg8_0),.din(w_dff_A_2JmFVYJO4_0),.clk(gclk));
	jdff dff_A_WcGcB9Zg8_0(.dout(w_dff_A_yMd3x3Gg2_0),.din(w_dff_A_WcGcB9Zg8_0),.clk(gclk));
	jdff dff_A_yMd3x3Gg2_0(.dout(w_dff_A_N5rLyz2h2_0),.din(w_dff_A_yMd3x3Gg2_0),.clk(gclk));
	jdff dff_A_N5rLyz2h2_0(.dout(w_dff_A_b718xl0k7_0),.din(w_dff_A_N5rLyz2h2_0),.clk(gclk));
	jdff dff_A_b718xl0k7_0(.dout(w_dff_A_yBtdBJDA7_0),.din(w_dff_A_b718xl0k7_0),.clk(gclk));
	jdff dff_A_yBtdBJDA7_0(.dout(w_dff_A_BUXDYlMr2_0),.din(w_dff_A_yBtdBJDA7_0),.clk(gclk));
	jdff dff_A_BUXDYlMr2_0(.dout(w_dff_A_EKQCWszx3_0),.din(w_dff_A_BUXDYlMr2_0),.clk(gclk));
	jdff dff_A_EKQCWszx3_0(.dout(w_dff_A_1sh2seEG3_0),.din(w_dff_A_EKQCWszx3_0),.clk(gclk));
	jdff dff_A_1sh2seEG3_0(.dout(f18),.din(w_dff_A_1sh2seEG3_0),.clk(gclk));
	jdff dff_A_Bp4ITOiF1_2(.dout(w_dff_A_jvMhEy0w4_0),.din(w_dff_A_Bp4ITOiF1_2),.clk(gclk));
	jdff dff_A_jvMhEy0w4_0(.dout(w_dff_A_puiqbAQJ0_0),.din(w_dff_A_jvMhEy0w4_0),.clk(gclk));
	jdff dff_A_puiqbAQJ0_0(.dout(w_dff_A_7OyJ08e32_0),.din(w_dff_A_puiqbAQJ0_0),.clk(gclk));
	jdff dff_A_7OyJ08e32_0(.dout(w_dff_A_K9STGv5v8_0),.din(w_dff_A_7OyJ08e32_0),.clk(gclk));
	jdff dff_A_K9STGv5v8_0(.dout(w_dff_A_hc21YYuw8_0),.din(w_dff_A_K9STGv5v8_0),.clk(gclk));
	jdff dff_A_hc21YYuw8_0(.dout(w_dff_A_cK8QsWnQ6_0),.din(w_dff_A_hc21YYuw8_0),.clk(gclk));
	jdff dff_A_cK8QsWnQ6_0(.dout(w_dff_A_pqJQEVZj6_0),.din(w_dff_A_cK8QsWnQ6_0),.clk(gclk));
	jdff dff_A_pqJQEVZj6_0(.dout(w_dff_A_Ve5qVmpp5_0),.din(w_dff_A_pqJQEVZj6_0),.clk(gclk));
	jdff dff_A_Ve5qVmpp5_0(.dout(w_dff_A_m1YTylw03_0),.din(w_dff_A_Ve5qVmpp5_0),.clk(gclk));
	jdff dff_A_m1YTylw03_0(.dout(w_dff_A_G9UEDFcj5_0),.din(w_dff_A_m1YTylw03_0),.clk(gclk));
	jdff dff_A_G9UEDFcj5_0(.dout(w_dff_A_hNduPF7j8_0),.din(w_dff_A_G9UEDFcj5_0),.clk(gclk));
	jdff dff_A_hNduPF7j8_0(.dout(w_dff_A_Pcauvq6G2_0),.din(w_dff_A_hNduPF7j8_0),.clk(gclk));
	jdff dff_A_Pcauvq6G2_0(.dout(w_dff_A_SeaAQBJf7_0),.din(w_dff_A_Pcauvq6G2_0),.clk(gclk));
	jdff dff_A_SeaAQBJf7_0(.dout(w_dff_A_rC2d8dQ85_0),.din(w_dff_A_SeaAQBJf7_0),.clk(gclk));
	jdff dff_A_rC2d8dQ85_0(.dout(w_dff_A_m8Ls7nyl0_0),.din(w_dff_A_rC2d8dQ85_0),.clk(gclk));
	jdff dff_A_m8Ls7nyl0_0(.dout(w_dff_A_nqunztJd7_0),.din(w_dff_A_m8Ls7nyl0_0),.clk(gclk));
	jdff dff_A_nqunztJd7_0(.dout(w_dff_A_m6k4tKll4_0),.din(w_dff_A_nqunztJd7_0),.clk(gclk));
	jdff dff_A_m6k4tKll4_0(.dout(w_dff_A_yZxNEeS50_0),.din(w_dff_A_m6k4tKll4_0),.clk(gclk));
	jdff dff_A_yZxNEeS50_0(.dout(w_dff_A_DiBA0nA22_0),.din(w_dff_A_yZxNEeS50_0),.clk(gclk));
	jdff dff_A_DiBA0nA22_0(.dout(w_dff_A_XRJDC3bM5_0),.din(w_dff_A_DiBA0nA22_0),.clk(gclk));
	jdff dff_A_XRJDC3bM5_0(.dout(w_dff_A_6CoknTaN6_0),.din(w_dff_A_XRJDC3bM5_0),.clk(gclk));
	jdff dff_A_6CoknTaN6_0(.dout(w_dff_A_qTtQNH2l9_0),.din(w_dff_A_6CoknTaN6_0),.clk(gclk));
	jdff dff_A_qTtQNH2l9_0(.dout(w_dff_A_30UqPXbZ2_0),.din(w_dff_A_qTtQNH2l9_0),.clk(gclk));
	jdff dff_A_30UqPXbZ2_0(.dout(w_dff_A_yzdiOauz1_0),.din(w_dff_A_30UqPXbZ2_0),.clk(gclk));
	jdff dff_A_yzdiOauz1_0(.dout(w_dff_A_EGFE87tl0_0),.din(w_dff_A_yzdiOauz1_0),.clk(gclk));
	jdff dff_A_EGFE87tl0_0(.dout(w_dff_A_9GPV57NR4_0),.din(w_dff_A_EGFE87tl0_0),.clk(gclk));
	jdff dff_A_9GPV57NR4_0(.dout(w_dff_A_DCyGSsyH7_0),.din(w_dff_A_9GPV57NR4_0),.clk(gclk));
	jdff dff_A_DCyGSsyH7_0(.dout(w_dff_A_J7K5a11g6_0),.din(w_dff_A_DCyGSsyH7_0),.clk(gclk));
	jdff dff_A_J7K5a11g6_0(.dout(w_dff_A_JMdkWgCK1_0),.din(w_dff_A_J7K5a11g6_0),.clk(gclk));
	jdff dff_A_JMdkWgCK1_0(.dout(w_dff_A_uQewDmo25_0),.din(w_dff_A_JMdkWgCK1_0),.clk(gclk));
	jdff dff_A_uQewDmo25_0(.dout(w_dff_A_ryzdhsBi2_0),.din(w_dff_A_uQewDmo25_0),.clk(gclk));
	jdff dff_A_ryzdhsBi2_0(.dout(w_dff_A_8sXp3TtB0_0),.din(w_dff_A_ryzdhsBi2_0),.clk(gclk));
	jdff dff_A_8sXp3TtB0_0(.dout(w_dff_A_iR67T7ca6_0),.din(w_dff_A_8sXp3TtB0_0),.clk(gclk));
	jdff dff_A_iR67T7ca6_0(.dout(w_dff_A_5xm66XVX3_0),.din(w_dff_A_iR67T7ca6_0),.clk(gclk));
	jdff dff_A_5xm66XVX3_0(.dout(w_dff_A_L2ZpyEHo1_0),.din(w_dff_A_5xm66XVX3_0),.clk(gclk));
	jdff dff_A_L2ZpyEHo1_0(.dout(w_dff_A_J5C6ccrW5_0),.din(w_dff_A_L2ZpyEHo1_0),.clk(gclk));
	jdff dff_A_J5C6ccrW5_0(.dout(w_dff_A_5OHCCJXW4_0),.din(w_dff_A_J5C6ccrW5_0),.clk(gclk));
	jdff dff_A_5OHCCJXW4_0(.dout(w_dff_A_7jfb9PZq1_0),.din(w_dff_A_5OHCCJXW4_0),.clk(gclk));
	jdff dff_A_7jfb9PZq1_0(.dout(w_dff_A_6IHFroO32_0),.din(w_dff_A_7jfb9PZq1_0),.clk(gclk));
	jdff dff_A_6IHFroO32_0(.dout(w_dff_A_4KQsbQom0_0),.din(w_dff_A_6IHFroO32_0),.clk(gclk));
	jdff dff_A_4KQsbQom0_0(.dout(w_dff_A_6u5Tfjln1_0),.din(w_dff_A_4KQsbQom0_0),.clk(gclk));
	jdff dff_A_6u5Tfjln1_0(.dout(w_dff_A_el4kXqXE6_0),.din(w_dff_A_6u5Tfjln1_0),.clk(gclk));
	jdff dff_A_el4kXqXE6_0(.dout(w_dff_A_cTMl91cR1_0),.din(w_dff_A_el4kXqXE6_0),.clk(gclk));
	jdff dff_A_cTMl91cR1_0(.dout(w_dff_A_cdypmyVO9_0),.din(w_dff_A_cTMl91cR1_0),.clk(gclk));
	jdff dff_A_cdypmyVO9_0(.dout(w_dff_A_pg18zwdY9_0),.din(w_dff_A_cdypmyVO9_0),.clk(gclk));
	jdff dff_A_pg18zwdY9_0(.dout(w_dff_A_1RWiZGir1_0),.din(w_dff_A_pg18zwdY9_0),.clk(gclk));
	jdff dff_A_1RWiZGir1_0(.dout(w_dff_A_Yqaqp5Sk0_0),.din(w_dff_A_1RWiZGir1_0),.clk(gclk));
	jdff dff_A_Yqaqp5Sk0_0(.dout(w_dff_A_1NlbArOp3_0),.din(w_dff_A_Yqaqp5Sk0_0),.clk(gclk));
	jdff dff_A_1NlbArOp3_0(.dout(w_dff_A_VrEsTOyr9_0),.din(w_dff_A_1NlbArOp3_0),.clk(gclk));
	jdff dff_A_VrEsTOyr9_0(.dout(w_dff_A_ij3597uh2_0),.din(w_dff_A_VrEsTOyr9_0),.clk(gclk));
	jdff dff_A_ij3597uh2_0(.dout(w_dff_A_LJrcCYPh6_0),.din(w_dff_A_ij3597uh2_0),.clk(gclk));
	jdff dff_A_LJrcCYPh6_0(.dout(w_dff_A_DUX6RMZG2_0),.din(w_dff_A_LJrcCYPh6_0),.clk(gclk));
	jdff dff_A_DUX6RMZG2_0(.dout(w_dff_A_ojpIOoXX6_0),.din(w_dff_A_DUX6RMZG2_0),.clk(gclk));
	jdff dff_A_ojpIOoXX6_0(.dout(w_dff_A_vCU6N5y40_0),.din(w_dff_A_ojpIOoXX6_0),.clk(gclk));
	jdff dff_A_vCU6N5y40_0(.dout(w_dff_A_RgvLKoKM6_0),.din(w_dff_A_vCU6N5y40_0),.clk(gclk));
	jdff dff_A_RgvLKoKM6_0(.dout(w_dff_A_g8Oi2kgh1_0),.din(w_dff_A_RgvLKoKM6_0),.clk(gclk));
	jdff dff_A_g8Oi2kgh1_0(.dout(w_dff_A_nq8tb7K39_0),.din(w_dff_A_g8Oi2kgh1_0),.clk(gclk));
	jdff dff_A_nq8tb7K39_0(.dout(w_dff_A_ymovtUPC6_0),.din(w_dff_A_nq8tb7K39_0),.clk(gclk));
	jdff dff_A_ymovtUPC6_0(.dout(w_dff_A_gs5PXvFi5_0),.din(w_dff_A_ymovtUPC6_0),.clk(gclk));
	jdff dff_A_gs5PXvFi5_0(.dout(w_dff_A_jouTIX5H4_0),.din(w_dff_A_gs5PXvFi5_0),.clk(gclk));
	jdff dff_A_jouTIX5H4_0(.dout(w_dff_A_x00fOAnh5_0),.din(w_dff_A_jouTIX5H4_0),.clk(gclk));
	jdff dff_A_x00fOAnh5_0(.dout(w_dff_A_qwQib3Cc3_0),.din(w_dff_A_x00fOAnh5_0),.clk(gclk));
	jdff dff_A_qwQib3Cc3_0(.dout(w_dff_A_3qVRkpfc8_0),.din(w_dff_A_qwQib3Cc3_0),.clk(gclk));
	jdff dff_A_3qVRkpfc8_0(.dout(w_dff_A_Djd8YOcl7_0),.din(w_dff_A_3qVRkpfc8_0),.clk(gclk));
	jdff dff_A_Djd8YOcl7_0(.dout(w_dff_A_7VSZ3mKu9_0),.din(w_dff_A_Djd8YOcl7_0),.clk(gclk));
	jdff dff_A_7VSZ3mKu9_0(.dout(w_dff_A_0dP8F4lu6_0),.din(w_dff_A_7VSZ3mKu9_0),.clk(gclk));
	jdff dff_A_0dP8F4lu6_0(.dout(w_dff_A_91S9c9Zg9_0),.din(w_dff_A_0dP8F4lu6_0),.clk(gclk));
	jdff dff_A_91S9c9Zg9_0(.dout(w_dff_A_scFQk9JK8_0),.din(w_dff_A_91S9c9Zg9_0),.clk(gclk));
	jdff dff_A_scFQk9JK8_0(.dout(w_dff_A_38WyhstZ1_0),.din(w_dff_A_scFQk9JK8_0),.clk(gclk));
	jdff dff_A_38WyhstZ1_0(.dout(w_dff_A_EBnWxIgM4_0),.din(w_dff_A_38WyhstZ1_0),.clk(gclk));
	jdff dff_A_EBnWxIgM4_0(.dout(w_dff_A_ZWMmg8BO0_0),.din(w_dff_A_EBnWxIgM4_0),.clk(gclk));
	jdff dff_A_ZWMmg8BO0_0(.dout(w_dff_A_htbS2hd94_0),.din(w_dff_A_ZWMmg8BO0_0),.clk(gclk));
	jdff dff_A_htbS2hd94_0(.dout(w_dff_A_B99DhVL18_0),.din(w_dff_A_htbS2hd94_0),.clk(gclk));
	jdff dff_A_B99DhVL18_0(.dout(w_dff_A_tq71fueL5_0),.din(w_dff_A_B99DhVL18_0),.clk(gclk));
	jdff dff_A_tq71fueL5_0(.dout(w_dff_A_BvJn82Ka8_0),.din(w_dff_A_tq71fueL5_0),.clk(gclk));
	jdff dff_A_BvJn82Ka8_0(.dout(w_dff_A_dEFFalXI5_0),.din(w_dff_A_BvJn82Ka8_0),.clk(gclk));
	jdff dff_A_dEFFalXI5_0(.dout(w_dff_A_HC7qwXAW2_0),.din(w_dff_A_dEFFalXI5_0),.clk(gclk));
	jdff dff_A_HC7qwXAW2_0(.dout(w_dff_A_GoYp4wky2_0),.din(w_dff_A_HC7qwXAW2_0),.clk(gclk));
	jdff dff_A_GoYp4wky2_0(.dout(w_dff_A_LkpETppz5_0),.din(w_dff_A_GoYp4wky2_0),.clk(gclk));
	jdff dff_A_LkpETppz5_0(.dout(w_dff_A_im0SIaHK6_0),.din(w_dff_A_LkpETppz5_0),.clk(gclk));
	jdff dff_A_im0SIaHK6_0(.dout(w_dff_A_JnZ8YA4g9_0),.din(w_dff_A_im0SIaHK6_0),.clk(gclk));
	jdff dff_A_JnZ8YA4g9_0(.dout(w_dff_A_x7cJdx304_0),.din(w_dff_A_JnZ8YA4g9_0),.clk(gclk));
	jdff dff_A_x7cJdx304_0(.dout(w_dff_A_weVeiff28_0),.din(w_dff_A_x7cJdx304_0),.clk(gclk));
	jdff dff_A_weVeiff28_0(.dout(w_dff_A_v3kfMOSZ9_0),.din(w_dff_A_weVeiff28_0),.clk(gclk));
	jdff dff_A_v3kfMOSZ9_0(.dout(w_dff_A_VnI56l6h0_0),.din(w_dff_A_v3kfMOSZ9_0),.clk(gclk));
	jdff dff_A_VnI56l6h0_0(.dout(w_dff_A_TeswHEfx1_0),.din(w_dff_A_VnI56l6h0_0),.clk(gclk));
	jdff dff_A_TeswHEfx1_0(.dout(w_dff_A_3AM0Dykc1_0),.din(w_dff_A_TeswHEfx1_0),.clk(gclk));
	jdff dff_A_3AM0Dykc1_0(.dout(w_dff_A_s8HIqjjZ9_0),.din(w_dff_A_3AM0Dykc1_0),.clk(gclk));
	jdff dff_A_s8HIqjjZ9_0(.dout(w_dff_A_POiu1HVf9_0),.din(w_dff_A_s8HIqjjZ9_0),.clk(gclk));
	jdff dff_A_POiu1HVf9_0(.dout(w_dff_A_iD2LdKTY9_0),.din(w_dff_A_POiu1HVf9_0),.clk(gclk));
	jdff dff_A_iD2LdKTY9_0(.dout(w_dff_A_7twhiEC58_0),.din(w_dff_A_iD2LdKTY9_0),.clk(gclk));
	jdff dff_A_7twhiEC58_0(.dout(w_dff_A_LfWqBv3s9_0),.din(w_dff_A_7twhiEC58_0),.clk(gclk));
	jdff dff_A_LfWqBv3s9_0(.dout(w_dff_A_NXIQYlJs4_0),.din(w_dff_A_LfWqBv3s9_0),.clk(gclk));
	jdff dff_A_NXIQYlJs4_0(.dout(w_dff_A_a7MwbyCF7_0),.din(w_dff_A_NXIQYlJs4_0),.clk(gclk));
	jdff dff_A_a7MwbyCF7_0(.dout(w_dff_A_qDSEG6sJ3_0),.din(w_dff_A_a7MwbyCF7_0),.clk(gclk));
	jdff dff_A_qDSEG6sJ3_0(.dout(w_dff_A_R2IheBoY1_0),.din(w_dff_A_qDSEG6sJ3_0),.clk(gclk));
	jdff dff_A_R2IheBoY1_0(.dout(w_dff_A_qQ7bp2U02_0),.din(w_dff_A_R2IheBoY1_0),.clk(gclk));
	jdff dff_A_qQ7bp2U02_0(.dout(w_dff_A_O8aSecI10_0),.din(w_dff_A_qQ7bp2U02_0),.clk(gclk));
	jdff dff_A_O8aSecI10_0(.dout(w_dff_A_2IWgLiww5_0),.din(w_dff_A_O8aSecI10_0),.clk(gclk));
	jdff dff_A_2IWgLiww5_0(.dout(w_dff_A_1J7GUhos8_0),.din(w_dff_A_2IWgLiww5_0),.clk(gclk));
	jdff dff_A_1J7GUhos8_0(.dout(w_dff_A_Vbg1HtEm6_0),.din(w_dff_A_1J7GUhos8_0),.clk(gclk));
	jdff dff_A_Vbg1HtEm6_0(.dout(w_dff_A_8nBXHZve6_0),.din(w_dff_A_Vbg1HtEm6_0),.clk(gclk));
	jdff dff_A_8nBXHZve6_0(.dout(w_dff_A_IU0ZPoAs6_0),.din(w_dff_A_8nBXHZve6_0),.clk(gclk));
	jdff dff_A_IU0ZPoAs6_0(.dout(w_dff_A_45yVBPQW0_0),.din(w_dff_A_IU0ZPoAs6_0),.clk(gclk));
	jdff dff_A_45yVBPQW0_0(.dout(w_dff_A_VpiuJnI57_0),.din(w_dff_A_45yVBPQW0_0),.clk(gclk));
	jdff dff_A_VpiuJnI57_0(.dout(w_dff_A_pUbe4B8Y8_0),.din(w_dff_A_VpiuJnI57_0),.clk(gclk));
	jdff dff_A_pUbe4B8Y8_0(.dout(w_dff_A_vNKOVZgK2_0),.din(w_dff_A_pUbe4B8Y8_0),.clk(gclk));
	jdff dff_A_vNKOVZgK2_0(.dout(f19),.din(w_dff_A_vNKOVZgK2_0),.clk(gclk));
	jdff dff_A_UvvGn9rX2_2(.dout(w_dff_A_8qGKI0RE0_0),.din(w_dff_A_UvvGn9rX2_2),.clk(gclk));
	jdff dff_A_8qGKI0RE0_0(.dout(w_dff_A_wZEg82Zz8_0),.din(w_dff_A_8qGKI0RE0_0),.clk(gclk));
	jdff dff_A_wZEg82Zz8_0(.dout(w_dff_A_mncMAK0q7_0),.din(w_dff_A_wZEg82Zz8_0),.clk(gclk));
	jdff dff_A_mncMAK0q7_0(.dout(w_dff_A_lGkx8MuB8_0),.din(w_dff_A_mncMAK0q7_0),.clk(gclk));
	jdff dff_A_lGkx8MuB8_0(.dout(w_dff_A_UIzdue6V0_0),.din(w_dff_A_lGkx8MuB8_0),.clk(gclk));
	jdff dff_A_UIzdue6V0_0(.dout(w_dff_A_gLD5VCrV3_0),.din(w_dff_A_UIzdue6V0_0),.clk(gclk));
	jdff dff_A_gLD5VCrV3_0(.dout(w_dff_A_gi3QU3QK9_0),.din(w_dff_A_gLD5VCrV3_0),.clk(gclk));
	jdff dff_A_gi3QU3QK9_0(.dout(w_dff_A_uLKcvOBz3_0),.din(w_dff_A_gi3QU3QK9_0),.clk(gclk));
	jdff dff_A_uLKcvOBz3_0(.dout(w_dff_A_4FTt6KVL3_0),.din(w_dff_A_uLKcvOBz3_0),.clk(gclk));
	jdff dff_A_4FTt6KVL3_0(.dout(w_dff_A_cVuFZiSb1_0),.din(w_dff_A_4FTt6KVL3_0),.clk(gclk));
	jdff dff_A_cVuFZiSb1_0(.dout(w_dff_A_IUTnGK8V2_0),.din(w_dff_A_cVuFZiSb1_0),.clk(gclk));
	jdff dff_A_IUTnGK8V2_0(.dout(w_dff_A_C3rhQdvh8_0),.din(w_dff_A_IUTnGK8V2_0),.clk(gclk));
	jdff dff_A_C3rhQdvh8_0(.dout(w_dff_A_8Zpd6bTi0_0),.din(w_dff_A_C3rhQdvh8_0),.clk(gclk));
	jdff dff_A_8Zpd6bTi0_0(.dout(w_dff_A_h4tYWMGz7_0),.din(w_dff_A_8Zpd6bTi0_0),.clk(gclk));
	jdff dff_A_h4tYWMGz7_0(.dout(w_dff_A_zubNrUp77_0),.din(w_dff_A_h4tYWMGz7_0),.clk(gclk));
	jdff dff_A_zubNrUp77_0(.dout(w_dff_A_FTlVkIkD3_0),.din(w_dff_A_zubNrUp77_0),.clk(gclk));
	jdff dff_A_FTlVkIkD3_0(.dout(w_dff_A_G5w5MOZf8_0),.din(w_dff_A_FTlVkIkD3_0),.clk(gclk));
	jdff dff_A_G5w5MOZf8_0(.dout(w_dff_A_iTK3nIE62_0),.din(w_dff_A_G5w5MOZf8_0),.clk(gclk));
	jdff dff_A_iTK3nIE62_0(.dout(w_dff_A_w0SUd0hn6_0),.din(w_dff_A_iTK3nIE62_0),.clk(gclk));
	jdff dff_A_w0SUd0hn6_0(.dout(w_dff_A_rr4a6nIK1_0),.din(w_dff_A_w0SUd0hn6_0),.clk(gclk));
	jdff dff_A_rr4a6nIK1_0(.dout(w_dff_A_JKnHVHzs3_0),.din(w_dff_A_rr4a6nIK1_0),.clk(gclk));
	jdff dff_A_JKnHVHzs3_0(.dout(w_dff_A_wT7ix1Px7_0),.din(w_dff_A_JKnHVHzs3_0),.clk(gclk));
	jdff dff_A_wT7ix1Px7_0(.dout(w_dff_A_QWACnWA75_0),.din(w_dff_A_wT7ix1Px7_0),.clk(gclk));
	jdff dff_A_QWACnWA75_0(.dout(w_dff_A_4elQGf0A5_0),.din(w_dff_A_QWACnWA75_0),.clk(gclk));
	jdff dff_A_4elQGf0A5_0(.dout(w_dff_A_3EDvDyQh8_0),.din(w_dff_A_4elQGf0A5_0),.clk(gclk));
	jdff dff_A_3EDvDyQh8_0(.dout(w_dff_A_4H2rBl3T7_0),.din(w_dff_A_3EDvDyQh8_0),.clk(gclk));
	jdff dff_A_4H2rBl3T7_0(.dout(w_dff_A_xaEvi8XX3_0),.din(w_dff_A_4H2rBl3T7_0),.clk(gclk));
	jdff dff_A_xaEvi8XX3_0(.dout(w_dff_A_AFE4a6kQ6_0),.din(w_dff_A_xaEvi8XX3_0),.clk(gclk));
	jdff dff_A_AFE4a6kQ6_0(.dout(w_dff_A_4LrasE4A6_0),.din(w_dff_A_AFE4a6kQ6_0),.clk(gclk));
	jdff dff_A_4LrasE4A6_0(.dout(w_dff_A_AbuQaFpq7_0),.din(w_dff_A_4LrasE4A6_0),.clk(gclk));
	jdff dff_A_AbuQaFpq7_0(.dout(w_dff_A_n6VYAloR6_0),.din(w_dff_A_AbuQaFpq7_0),.clk(gclk));
	jdff dff_A_n6VYAloR6_0(.dout(w_dff_A_8C69epkn0_0),.din(w_dff_A_n6VYAloR6_0),.clk(gclk));
	jdff dff_A_8C69epkn0_0(.dout(w_dff_A_6sCTv7YC9_0),.din(w_dff_A_8C69epkn0_0),.clk(gclk));
	jdff dff_A_6sCTv7YC9_0(.dout(w_dff_A_fvWKkfVd2_0),.din(w_dff_A_6sCTv7YC9_0),.clk(gclk));
	jdff dff_A_fvWKkfVd2_0(.dout(w_dff_A_Ps6BVgVk1_0),.din(w_dff_A_fvWKkfVd2_0),.clk(gclk));
	jdff dff_A_Ps6BVgVk1_0(.dout(w_dff_A_EgPX5KQE0_0),.din(w_dff_A_Ps6BVgVk1_0),.clk(gclk));
	jdff dff_A_EgPX5KQE0_0(.dout(w_dff_A_E7idzcbD4_0),.din(w_dff_A_EgPX5KQE0_0),.clk(gclk));
	jdff dff_A_E7idzcbD4_0(.dout(w_dff_A_YZ4GsjPS8_0),.din(w_dff_A_E7idzcbD4_0),.clk(gclk));
	jdff dff_A_YZ4GsjPS8_0(.dout(w_dff_A_oH7Srzv53_0),.din(w_dff_A_YZ4GsjPS8_0),.clk(gclk));
	jdff dff_A_oH7Srzv53_0(.dout(w_dff_A_oxZpepLt2_0),.din(w_dff_A_oH7Srzv53_0),.clk(gclk));
	jdff dff_A_oxZpepLt2_0(.dout(w_dff_A_AmMRAFFv3_0),.din(w_dff_A_oxZpepLt2_0),.clk(gclk));
	jdff dff_A_AmMRAFFv3_0(.dout(w_dff_A_mrpUq6Z82_0),.din(w_dff_A_AmMRAFFv3_0),.clk(gclk));
	jdff dff_A_mrpUq6Z82_0(.dout(w_dff_A_nRjCnJhy4_0),.din(w_dff_A_mrpUq6Z82_0),.clk(gclk));
	jdff dff_A_nRjCnJhy4_0(.dout(w_dff_A_n3nWSkU31_0),.din(w_dff_A_nRjCnJhy4_0),.clk(gclk));
	jdff dff_A_n3nWSkU31_0(.dout(w_dff_A_rUNMMlhJ6_0),.din(w_dff_A_n3nWSkU31_0),.clk(gclk));
	jdff dff_A_rUNMMlhJ6_0(.dout(w_dff_A_SKnDkxxv6_0),.din(w_dff_A_rUNMMlhJ6_0),.clk(gclk));
	jdff dff_A_SKnDkxxv6_0(.dout(w_dff_A_kAlCYB6y2_0),.din(w_dff_A_SKnDkxxv6_0),.clk(gclk));
	jdff dff_A_kAlCYB6y2_0(.dout(w_dff_A_Iqo0yklh8_0),.din(w_dff_A_kAlCYB6y2_0),.clk(gclk));
	jdff dff_A_Iqo0yklh8_0(.dout(w_dff_A_zMWDgjx27_0),.din(w_dff_A_Iqo0yklh8_0),.clk(gclk));
	jdff dff_A_zMWDgjx27_0(.dout(w_dff_A_A0xLaTrl7_0),.din(w_dff_A_zMWDgjx27_0),.clk(gclk));
	jdff dff_A_A0xLaTrl7_0(.dout(w_dff_A_HfKHwlDi5_0),.din(w_dff_A_A0xLaTrl7_0),.clk(gclk));
	jdff dff_A_HfKHwlDi5_0(.dout(w_dff_A_iDy24gsk4_0),.din(w_dff_A_HfKHwlDi5_0),.clk(gclk));
	jdff dff_A_iDy24gsk4_0(.dout(w_dff_A_KfmWXslX6_0),.din(w_dff_A_iDy24gsk4_0),.clk(gclk));
	jdff dff_A_KfmWXslX6_0(.dout(w_dff_A_psXl9lrP8_0),.din(w_dff_A_KfmWXslX6_0),.clk(gclk));
	jdff dff_A_psXl9lrP8_0(.dout(w_dff_A_zvymgTgE2_0),.din(w_dff_A_psXl9lrP8_0),.clk(gclk));
	jdff dff_A_zvymgTgE2_0(.dout(w_dff_A_vm4ecouK0_0),.din(w_dff_A_zvymgTgE2_0),.clk(gclk));
	jdff dff_A_vm4ecouK0_0(.dout(w_dff_A_iFKsiyEU8_0),.din(w_dff_A_vm4ecouK0_0),.clk(gclk));
	jdff dff_A_iFKsiyEU8_0(.dout(w_dff_A_tYvWPRNK3_0),.din(w_dff_A_iFKsiyEU8_0),.clk(gclk));
	jdff dff_A_tYvWPRNK3_0(.dout(w_dff_A_JahjJTGg0_0),.din(w_dff_A_tYvWPRNK3_0),.clk(gclk));
	jdff dff_A_JahjJTGg0_0(.dout(w_dff_A_KwwizCYN5_0),.din(w_dff_A_JahjJTGg0_0),.clk(gclk));
	jdff dff_A_KwwizCYN5_0(.dout(w_dff_A_VOgAkZLq2_0),.din(w_dff_A_KwwizCYN5_0),.clk(gclk));
	jdff dff_A_VOgAkZLq2_0(.dout(w_dff_A_ReRfwaqf9_0),.din(w_dff_A_VOgAkZLq2_0),.clk(gclk));
	jdff dff_A_ReRfwaqf9_0(.dout(w_dff_A_8lXzZFzS5_0),.din(w_dff_A_ReRfwaqf9_0),.clk(gclk));
	jdff dff_A_8lXzZFzS5_0(.dout(w_dff_A_kV1xeooL7_0),.din(w_dff_A_8lXzZFzS5_0),.clk(gclk));
	jdff dff_A_kV1xeooL7_0(.dout(w_dff_A_Ug59nff18_0),.din(w_dff_A_kV1xeooL7_0),.clk(gclk));
	jdff dff_A_Ug59nff18_0(.dout(w_dff_A_dljAIf8o1_0),.din(w_dff_A_Ug59nff18_0),.clk(gclk));
	jdff dff_A_dljAIf8o1_0(.dout(w_dff_A_90qzFw8Z0_0),.din(w_dff_A_dljAIf8o1_0),.clk(gclk));
	jdff dff_A_90qzFw8Z0_0(.dout(w_dff_A_cwBFOqul1_0),.din(w_dff_A_90qzFw8Z0_0),.clk(gclk));
	jdff dff_A_cwBFOqul1_0(.dout(w_dff_A_qzhBt72e5_0),.din(w_dff_A_cwBFOqul1_0),.clk(gclk));
	jdff dff_A_qzhBt72e5_0(.dout(w_dff_A_jZLHhsEk4_0),.din(w_dff_A_qzhBt72e5_0),.clk(gclk));
	jdff dff_A_jZLHhsEk4_0(.dout(w_dff_A_blQi8cHc4_0),.din(w_dff_A_jZLHhsEk4_0),.clk(gclk));
	jdff dff_A_blQi8cHc4_0(.dout(w_dff_A_jR5xStDa0_0),.din(w_dff_A_blQi8cHc4_0),.clk(gclk));
	jdff dff_A_jR5xStDa0_0(.dout(w_dff_A_7dgUCgTw7_0),.din(w_dff_A_jR5xStDa0_0),.clk(gclk));
	jdff dff_A_7dgUCgTw7_0(.dout(w_dff_A_CUVlYVML3_0),.din(w_dff_A_7dgUCgTw7_0),.clk(gclk));
	jdff dff_A_CUVlYVML3_0(.dout(w_dff_A_g6xHjmhg3_0),.din(w_dff_A_CUVlYVML3_0),.clk(gclk));
	jdff dff_A_g6xHjmhg3_0(.dout(w_dff_A_9wBVthNS5_0),.din(w_dff_A_g6xHjmhg3_0),.clk(gclk));
	jdff dff_A_9wBVthNS5_0(.dout(w_dff_A_HWuUvGrz7_0),.din(w_dff_A_9wBVthNS5_0),.clk(gclk));
	jdff dff_A_HWuUvGrz7_0(.dout(w_dff_A_KgwQzC4l7_0),.din(w_dff_A_HWuUvGrz7_0),.clk(gclk));
	jdff dff_A_KgwQzC4l7_0(.dout(w_dff_A_MHZkWSvw5_0),.din(w_dff_A_KgwQzC4l7_0),.clk(gclk));
	jdff dff_A_MHZkWSvw5_0(.dout(w_dff_A_UGOO3Pty4_0),.din(w_dff_A_MHZkWSvw5_0),.clk(gclk));
	jdff dff_A_UGOO3Pty4_0(.dout(w_dff_A_d8Av83NJ8_0),.din(w_dff_A_UGOO3Pty4_0),.clk(gclk));
	jdff dff_A_d8Av83NJ8_0(.dout(w_dff_A_rFsdYm2n6_0),.din(w_dff_A_d8Av83NJ8_0),.clk(gclk));
	jdff dff_A_rFsdYm2n6_0(.dout(w_dff_A_q1h92xXi7_0),.din(w_dff_A_rFsdYm2n6_0),.clk(gclk));
	jdff dff_A_q1h92xXi7_0(.dout(w_dff_A_PqUmnpAS6_0),.din(w_dff_A_q1h92xXi7_0),.clk(gclk));
	jdff dff_A_PqUmnpAS6_0(.dout(w_dff_A_gfZByBoH1_0),.din(w_dff_A_PqUmnpAS6_0),.clk(gclk));
	jdff dff_A_gfZByBoH1_0(.dout(w_dff_A_Ze3Tq36k7_0),.din(w_dff_A_gfZByBoH1_0),.clk(gclk));
	jdff dff_A_Ze3Tq36k7_0(.dout(w_dff_A_Y9kY4jDj7_0),.din(w_dff_A_Ze3Tq36k7_0),.clk(gclk));
	jdff dff_A_Y9kY4jDj7_0(.dout(w_dff_A_Ta9DDjfu9_0),.din(w_dff_A_Y9kY4jDj7_0),.clk(gclk));
	jdff dff_A_Ta9DDjfu9_0(.dout(w_dff_A_FVsT9Xjy5_0),.din(w_dff_A_Ta9DDjfu9_0),.clk(gclk));
	jdff dff_A_FVsT9Xjy5_0(.dout(w_dff_A_B3dhimzS7_0),.din(w_dff_A_FVsT9Xjy5_0),.clk(gclk));
	jdff dff_A_B3dhimzS7_0(.dout(w_dff_A_k6yMc0VY5_0),.din(w_dff_A_B3dhimzS7_0),.clk(gclk));
	jdff dff_A_k6yMc0VY5_0(.dout(w_dff_A_MRHDy74K5_0),.din(w_dff_A_k6yMc0VY5_0),.clk(gclk));
	jdff dff_A_MRHDy74K5_0(.dout(w_dff_A_Jb5HEV1x5_0),.din(w_dff_A_MRHDy74K5_0),.clk(gclk));
	jdff dff_A_Jb5HEV1x5_0(.dout(w_dff_A_s3YVPPW46_0),.din(w_dff_A_Jb5HEV1x5_0),.clk(gclk));
	jdff dff_A_s3YVPPW46_0(.dout(w_dff_A_c6QvyV1A1_0),.din(w_dff_A_s3YVPPW46_0),.clk(gclk));
	jdff dff_A_c6QvyV1A1_0(.dout(w_dff_A_atiBqafO7_0),.din(w_dff_A_c6QvyV1A1_0),.clk(gclk));
	jdff dff_A_atiBqafO7_0(.dout(w_dff_A_HFVpFWCU2_0),.din(w_dff_A_atiBqafO7_0),.clk(gclk));
	jdff dff_A_HFVpFWCU2_0(.dout(w_dff_A_viN9fqdh0_0),.din(w_dff_A_HFVpFWCU2_0),.clk(gclk));
	jdff dff_A_viN9fqdh0_0(.dout(w_dff_A_4vPXxwVj5_0),.din(w_dff_A_viN9fqdh0_0),.clk(gclk));
	jdff dff_A_4vPXxwVj5_0(.dout(w_dff_A_89L2DePF6_0),.din(w_dff_A_4vPXxwVj5_0),.clk(gclk));
	jdff dff_A_89L2DePF6_0(.dout(w_dff_A_WBX00K669_0),.din(w_dff_A_89L2DePF6_0),.clk(gclk));
	jdff dff_A_WBX00K669_0(.dout(w_dff_A_FesiCaIL4_0),.din(w_dff_A_WBX00K669_0),.clk(gclk));
	jdff dff_A_FesiCaIL4_0(.dout(w_dff_A_nAGDZfi66_0),.din(w_dff_A_FesiCaIL4_0),.clk(gclk));
	jdff dff_A_nAGDZfi66_0(.dout(w_dff_A_KE3h50LS1_0),.din(w_dff_A_nAGDZfi66_0),.clk(gclk));
	jdff dff_A_KE3h50LS1_0(.dout(w_dff_A_bgW4cfhb5_0),.din(w_dff_A_KE3h50LS1_0),.clk(gclk));
	jdff dff_A_bgW4cfhb5_0(.dout(w_dff_A_gT40v9Uv7_0),.din(w_dff_A_bgW4cfhb5_0),.clk(gclk));
	jdff dff_A_gT40v9Uv7_0(.dout(f20),.din(w_dff_A_gT40v9Uv7_0),.clk(gclk));
	jdff dff_A_lCHLbsXY9_2(.dout(w_dff_A_5pd3pxCd0_0),.din(w_dff_A_lCHLbsXY9_2),.clk(gclk));
	jdff dff_A_5pd3pxCd0_0(.dout(w_dff_A_izdYvg859_0),.din(w_dff_A_5pd3pxCd0_0),.clk(gclk));
	jdff dff_A_izdYvg859_0(.dout(w_dff_A_Rnq3BGaR9_0),.din(w_dff_A_izdYvg859_0),.clk(gclk));
	jdff dff_A_Rnq3BGaR9_0(.dout(w_dff_A_xLXJHLSE6_0),.din(w_dff_A_Rnq3BGaR9_0),.clk(gclk));
	jdff dff_A_xLXJHLSE6_0(.dout(w_dff_A_hmZBM0wt7_0),.din(w_dff_A_xLXJHLSE6_0),.clk(gclk));
	jdff dff_A_hmZBM0wt7_0(.dout(w_dff_A_csFKwb7y5_0),.din(w_dff_A_hmZBM0wt7_0),.clk(gclk));
	jdff dff_A_csFKwb7y5_0(.dout(w_dff_A_b3HbDjZj1_0),.din(w_dff_A_csFKwb7y5_0),.clk(gclk));
	jdff dff_A_b3HbDjZj1_0(.dout(w_dff_A_mtH9pT4D9_0),.din(w_dff_A_b3HbDjZj1_0),.clk(gclk));
	jdff dff_A_mtH9pT4D9_0(.dout(w_dff_A_DAeIv3Tt1_0),.din(w_dff_A_mtH9pT4D9_0),.clk(gclk));
	jdff dff_A_DAeIv3Tt1_0(.dout(w_dff_A_1X6Bji5v1_0),.din(w_dff_A_DAeIv3Tt1_0),.clk(gclk));
	jdff dff_A_1X6Bji5v1_0(.dout(w_dff_A_da7VZ5i46_0),.din(w_dff_A_1X6Bji5v1_0),.clk(gclk));
	jdff dff_A_da7VZ5i46_0(.dout(w_dff_A_Efcg6eXY2_0),.din(w_dff_A_da7VZ5i46_0),.clk(gclk));
	jdff dff_A_Efcg6eXY2_0(.dout(w_dff_A_igECOkQg8_0),.din(w_dff_A_Efcg6eXY2_0),.clk(gclk));
	jdff dff_A_igECOkQg8_0(.dout(w_dff_A_xT9E5Qgl6_0),.din(w_dff_A_igECOkQg8_0),.clk(gclk));
	jdff dff_A_xT9E5Qgl6_0(.dout(w_dff_A_sWHgN6M18_0),.din(w_dff_A_xT9E5Qgl6_0),.clk(gclk));
	jdff dff_A_sWHgN6M18_0(.dout(w_dff_A_6x1RHjpr7_0),.din(w_dff_A_sWHgN6M18_0),.clk(gclk));
	jdff dff_A_6x1RHjpr7_0(.dout(w_dff_A_u4KgYuln5_0),.din(w_dff_A_6x1RHjpr7_0),.clk(gclk));
	jdff dff_A_u4KgYuln5_0(.dout(w_dff_A_txc1f1B08_0),.din(w_dff_A_u4KgYuln5_0),.clk(gclk));
	jdff dff_A_txc1f1B08_0(.dout(w_dff_A_J1rU6GpA4_0),.din(w_dff_A_txc1f1B08_0),.clk(gclk));
	jdff dff_A_J1rU6GpA4_0(.dout(w_dff_A_PGt4U0254_0),.din(w_dff_A_J1rU6GpA4_0),.clk(gclk));
	jdff dff_A_PGt4U0254_0(.dout(w_dff_A_eRyfysyt0_0),.din(w_dff_A_PGt4U0254_0),.clk(gclk));
	jdff dff_A_eRyfysyt0_0(.dout(w_dff_A_PMs9oPPU5_0),.din(w_dff_A_eRyfysyt0_0),.clk(gclk));
	jdff dff_A_PMs9oPPU5_0(.dout(w_dff_A_S2133bGj5_0),.din(w_dff_A_PMs9oPPU5_0),.clk(gclk));
	jdff dff_A_S2133bGj5_0(.dout(w_dff_A_UXqeLZWi2_0),.din(w_dff_A_S2133bGj5_0),.clk(gclk));
	jdff dff_A_UXqeLZWi2_0(.dout(w_dff_A_OevOKfvM9_0),.din(w_dff_A_UXqeLZWi2_0),.clk(gclk));
	jdff dff_A_OevOKfvM9_0(.dout(w_dff_A_WM6lGyIs4_0),.din(w_dff_A_OevOKfvM9_0),.clk(gclk));
	jdff dff_A_WM6lGyIs4_0(.dout(w_dff_A_2ldw2KTm9_0),.din(w_dff_A_WM6lGyIs4_0),.clk(gclk));
	jdff dff_A_2ldw2KTm9_0(.dout(w_dff_A_3R25R7Af4_0),.din(w_dff_A_2ldw2KTm9_0),.clk(gclk));
	jdff dff_A_3R25R7Af4_0(.dout(w_dff_A_J0OSiSBk0_0),.din(w_dff_A_3R25R7Af4_0),.clk(gclk));
	jdff dff_A_J0OSiSBk0_0(.dout(w_dff_A_RyVAaV5H7_0),.din(w_dff_A_J0OSiSBk0_0),.clk(gclk));
	jdff dff_A_RyVAaV5H7_0(.dout(w_dff_A_KdelyN9K4_0),.din(w_dff_A_RyVAaV5H7_0),.clk(gclk));
	jdff dff_A_KdelyN9K4_0(.dout(w_dff_A_KmxVKamR8_0),.din(w_dff_A_KdelyN9K4_0),.clk(gclk));
	jdff dff_A_KmxVKamR8_0(.dout(w_dff_A_u6FvbWQy9_0),.din(w_dff_A_KmxVKamR8_0),.clk(gclk));
	jdff dff_A_u6FvbWQy9_0(.dout(w_dff_A_ejHZVtyW7_0),.din(w_dff_A_u6FvbWQy9_0),.clk(gclk));
	jdff dff_A_ejHZVtyW7_0(.dout(w_dff_A_Q2r438ol0_0),.din(w_dff_A_ejHZVtyW7_0),.clk(gclk));
	jdff dff_A_Q2r438ol0_0(.dout(w_dff_A_RFrBKZ1D2_0),.din(w_dff_A_Q2r438ol0_0),.clk(gclk));
	jdff dff_A_RFrBKZ1D2_0(.dout(w_dff_A_3kqEJFzN1_0),.din(w_dff_A_RFrBKZ1D2_0),.clk(gclk));
	jdff dff_A_3kqEJFzN1_0(.dout(w_dff_A_U2hHdySL3_0),.din(w_dff_A_3kqEJFzN1_0),.clk(gclk));
	jdff dff_A_U2hHdySL3_0(.dout(w_dff_A_B185ummz5_0),.din(w_dff_A_U2hHdySL3_0),.clk(gclk));
	jdff dff_A_B185ummz5_0(.dout(w_dff_A_Vt4CpBhV9_0),.din(w_dff_A_B185ummz5_0),.clk(gclk));
	jdff dff_A_Vt4CpBhV9_0(.dout(w_dff_A_IWSCJtX40_0),.din(w_dff_A_Vt4CpBhV9_0),.clk(gclk));
	jdff dff_A_IWSCJtX40_0(.dout(w_dff_A_gk2j205J0_0),.din(w_dff_A_IWSCJtX40_0),.clk(gclk));
	jdff dff_A_gk2j205J0_0(.dout(w_dff_A_a0GYr0En4_0),.din(w_dff_A_gk2j205J0_0),.clk(gclk));
	jdff dff_A_a0GYr0En4_0(.dout(w_dff_A_v1KTRN0H7_0),.din(w_dff_A_a0GYr0En4_0),.clk(gclk));
	jdff dff_A_v1KTRN0H7_0(.dout(w_dff_A_C0WmJupj1_0),.din(w_dff_A_v1KTRN0H7_0),.clk(gclk));
	jdff dff_A_C0WmJupj1_0(.dout(w_dff_A_m1omsexu0_0),.din(w_dff_A_C0WmJupj1_0),.clk(gclk));
	jdff dff_A_m1omsexu0_0(.dout(w_dff_A_UhxrpWp47_0),.din(w_dff_A_m1omsexu0_0),.clk(gclk));
	jdff dff_A_UhxrpWp47_0(.dout(w_dff_A_42kPPQaw7_0),.din(w_dff_A_UhxrpWp47_0),.clk(gclk));
	jdff dff_A_42kPPQaw7_0(.dout(w_dff_A_IfHcsQ6I8_0),.din(w_dff_A_42kPPQaw7_0),.clk(gclk));
	jdff dff_A_IfHcsQ6I8_0(.dout(w_dff_A_hIWv5xfW4_0),.din(w_dff_A_IfHcsQ6I8_0),.clk(gclk));
	jdff dff_A_hIWv5xfW4_0(.dout(w_dff_A_SDFz8boM9_0),.din(w_dff_A_hIWv5xfW4_0),.clk(gclk));
	jdff dff_A_SDFz8boM9_0(.dout(w_dff_A_gjvaAsRC3_0),.din(w_dff_A_SDFz8boM9_0),.clk(gclk));
	jdff dff_A_gjvaAsRC3_0(.dout(w_dff_A_RSnX1Ozu6_0),.din(w_dff_A_gjvaAsRC3_0),.clk(gclk));
	jdff dff_A_RSnX1Ozu6_0(.dout(w_dff_A_FJ2goiww9_0),.din(w_dff_A_RSnX1Ozu6_0),.clk(gclk));
	jdff dff_A_FJ2goiww9_0(.dout(w_dff_A_kAO5oVl70_0),.din(w_dff_A_FJ2goiww9_0),.clk(gclk));
	jdff dff_A_kAO5oVl70_0(.dout(w_dff_A_VyA3rdJQ5_0),.din(w_dff_A_kAO5oVl70_0),.clk(gclk));
	jdff dff_A_VyA3rdJQ5_0(.dout(w_dff_A_RWsENUmU9_0),.din(w_dff_A_VyA3rdJQ5_0),.clk(gclk));
	jdff dff_A_RWsENUmU9_0(.dout(w_dff_A_1iGcRfvK9_0),.din(w_dff_A_RWsENUmU9_0),.clk(gclk));
	jdff dff_A_1iGcRfvK9_0(.dout(w_dff_A_ewafylVO7_0),.din(w_dff_A_1iGcRfvK9_0),.clk(gclk));
	jdff dff_A_ewafylVO7_0(.dout(w_dff_A_bu0qEqds3_0),.din(w_dff_A_ewafylVO7_0),.clk(gclk));
	jdff dff_A_bu0qEqds3_0(.dout(w_dff_A_83a87D6G6_0),.din(w_dff_A_bu0qEqds3_0),.clk(gclk));
	jdff dff_A_83a87D6G6_0(.dout(w_dff_A_9jMDtlyG7_0),.din(w_dff_A_83a87D6G6_0),.clk(gclk));
	jdff dff_A_9jMDtlyG7_0(.dout(w_dff_A_j0h2hltR9_0),.din(w_dff_A_9jMDtlyG7_0),.clk(gclk));
	jdff dff_A_j0h2hltR9_0(.dout(w_dff_A_dPTtqRAw3_0),.din(w_dff_A_j0h2hltR9_0),.clk(gclk));
	jdff dff_A_dPTtqRAw3_0(.dout(w_dff_A_vTbSlqOB8_0),.din(w_dff_A_dPTtqRAw3_0),.clk(gclk));
	jdff dff_A_vTbSlqOB8_0(.dout(w_dff_A_tsBUC5qc9_0),.din(w_dff_A_vTbSlqOB8_0),.clk(gclk));
	jdff dff_A_tsBUC5qc9_0(.dout(w_dff_A_WbpGKj4t4_0),.din(w_dff_A_tsBUC5qc9_0),.clk(gclk));
	jdff dff_A_WbpGKj4t4_0(.dout(w_dff_A_ArDe8fKK7_0),.din(w_dff_A_WbpGKj4t4_0),.clk(gclk));
	jdff dff_A_ArDe8fKK7_0(.dout(w_dff_A_UNmXbe9h8_0),.din(w_dff_A_ArDe8fKK7_0),.clk(gclk));
	jdff dff_A_UNmXbe9h8_0(.dout(w_dff_A_9uWF6XgJ1_0),.din(w_dff_A_UNmXbe9h8_0),.clk(gclk));
	jdff dff_A_9uWF6XgJ1_0(.dout(w_dff_A_ABs5pq959_0),.din(w_dff_A_9uWF6XgJ1_0),.clk(gclk));
	jdff dff_A_ABs5pq959_0(.dout(w_dff_A_WGMF3nzx0_0),.din(w_dff_A_ABs5pq959_0),.clk(gclk));
	jdff dff_A_WGMF3nzx0_0(.dout(w_dff_A_IHkl6Zr74_0),.din(w_dff_A_WGMF3nzx0_0),.clk(gclk));
	jdff dff_A_IHkl6Zr74_0(.dout(w_dff_A_DN5ZxBeK5_0),.din(w_dff_A_IHkl6Zr74_0),.clk(gclk));
	jdff dff_A_DN5ZxBeK5_0(.dout(w_dff_A_KhAGHMYt3_0),.din(w_dff_A_DN5ZxBeK5_0),.clk(gclk));
	jdff dff_A_KhAGHMYt3_0(.dout(w_dff_A_FhHNseIR4_0),.din(w_dff_A_KhAGHMYt3_0),.clk(gclk));
	jdff dff_A_FhHNseIR4_0(.dout(w_dff_A_vjBGIUKh4_0),.din(w_dff_A_FhHNseIR4_0),.clk(gclk));
	jdff dff_A_vjBGIUKh4_0(.dout(w_dff_A_QHQv3pTk9_0),.din(w_dff_A_vjBGIUKh4_0),.clk(gclk));
	jdff dff_A_QHQv3pTk9_0(.dout(w_dff_A_ix0FDSO22_0),.din(w_dff_A_QHQv3pTk9_0),.clk(gclk));
	jdff dff_A_ix0FDSO22_0(.dout(w_dff_A_QPBq49vp8_0),.din(w_dff_A_ix0FDSO22_0),.clk(gclk));
	jdff dff_A_QPBq49vp8_0(.dout(w_dff_A_Ok8pvOZ99_0),.din(w_dff_A_QPBq49vp8_0),.clk(gclk));
	jdff dff_A_Ok8pvOZ99_0(.dout(w_dff_A_RRr3kmrq1_0),.din(w_dff_A_Ok8pvOZ99_0),.clk(gclk));
	jdff dff_A_RRr3kmrq1_0(.dout(w_dff_A_RCd0t5l57_0),.din(w_dff_A_RRr3kmrq1_0),.clk(gclk));
	jdff dff_A_RCd0t5l57_0(.dout(w_dff_A_UfZNiuRo8_0),.din(w_dff_A_RCd0t5l57_0),.clk(gclk));
	jdff dff_A_UfZNiuRo8_0(.dout(w_dff_A_ULDYjV6J5_0),.din(w_dff_A_UfZNiuRo8_0),.clk(gclk));
	jdff dff_A_ULDYjV6J5_0(.dout(w_dff_A_qO7GpZOl8_0),.din(w_dff_A_ULDYjV6J5_0),.clk(gclk));
	jdff dff_A_qO7GpZOl8_0(.dout(w_dff_A_fUmXCxD37_0),.din(w_dff_A_qO7GpZOl8_0),.clk(gclk));
	jdff dff_A_fUmXCxD37_0(.dout(w_dff_A_8b28aMpw2_0),.din(w_dff_A_fUmXCxD37_0),.clk(gclk));
	jdff dff_A_8b28aMpw2_0(.dout(w_dff_A_hfGCvspW4_0),.din(w_dff_A_8b28aMpw2_0),.clk(gclk));
	jdff dff_A_hfGCvspW4_0(.dout(w_dff_A_8gZjpzUU4_0),.din(w_dff_A_hfGCvspW4_0),.clk(gclk));
	jdff dff_A_8gZjpzUU4_0(.dout(w_dff_A_gKELwUX22_0),.din(w_dff_A_8gZjpzUU4_0),.clk(gclk));
	jdff dff_A_gKELwUX22_0(.dout(w_dff_A_PyKsbI6B2_0),.din(w_dff_A_gKELwUX22_0),.clk(gclk));
	jdff dff_A_PyKsbI6B2_0(.dout(w_dff_A_woH1tcJQ1_0),.din(w_dff_A_PyKsbI6B2_0),.clk(gclk));
	jdff dff_A_woH1tcJQ1_0(.dout(w_dff_A_7mvaKFp77_0),.din(w_dff_A_woH1tcJQ1_0),.clk(gclk));
	jdff dff_A_7mvaKFp77_0(.dout(w_dff_A_eECTUFPl2_0),.din(w_dff_A_7mvaKFp77_0),.clk(gclk));
	jdff dff_A_eECTUFPl2_0(.dout(w_dff_A_HZ4hGMrp8_0),.din(w_dff_A_eECTUFPl2_0),.clk(gclk));
	jdff dff_A_HZ4hGMrp8_0(.dout(w_dff_A_XqSGPLTf6_0),.din(w_dff_A_HZ4hGMrp8_0),.clk(gclk));
	jdff dff_A_XqSGPLTf6_0(.dout(w_dff_A_g7joznxS5_0),.din(w_dff_A_XqSGPLTf6_0),.clk(gclk));
	jdff dff_A_g7joznxS5_0(.dout(w_dff_A_kCotj0PF2_0),.din(w_dff_A_g7joznxS5_0),.clk(gclk));
	jdff dff_A_kCotj0PF2_0(.dout(w_dff_A_oGC5CTXB7_0),.din(w_dff_A_kCotj0PF2_0),.clk(gclk));
	jdff dff_A_oGC5CTXB7_0(.dout(w_dff_A_vuLBUkkB2_0),.din(w_dff_A_oGC5CTXB7_0),.clk(gclk));
	jdff dff_A_vuLBUkkB2_0(.dout(w_dff_A_galTre5O3_0),.din(w_dff_A_vuLBUkkB2_0),.clk(gclk));
	jdff dff_A_galTre5O3_0(.dout(w_dff_A_tOPjkisW3_0),.din(w_dff_A_galTre5O3_0),.clk(gclk));
	jdff dff_A_tOPjkisW3_0(.dout(w_dff_A_d1ZSvvVt7_0),.din(w_dff_A_tOPjkisW3_0),.clk(gclk));
	jdff dff_A_d1ZSvvVt7_0(.dout(w_dff_A_ArwO2Kdi0_0),.din(w_dff_A_d1ZSvvVt7_0),.clk(gclk));
	jdff dff_A_ArwO2Kdi0_0(.dout(f21),.din(w_dff_A_ArwO2Kdi0_0),.clk(gclk));
	jdff dff_A_bwlIPVrT6_2(.dout(w_dff_A_8FzXY3168_0),.din(w_dff_A_bwlIPVrT6_2),.clk(gclk));
	jdff dff_A_8FzXY3168_0(.dout(w_dff_A_A6vbtUuC7_0),.din(w_dff_A_8FzXY3168_0),.clk(gclk));
	jdff dff_A_A6vbtUuC7_0(.dout(w_dff_A_HM2WTPae1_0),.din(w_dff_A_A6vbtUuC7_0),.clk(gclk));
	jdff dff_A_HM2WTPae1_0(.dout(w_dff_A_tyIBQehs4_0),.din(w_dff_A_HM2WTPae1_0),.clk(gclk));
	jdff dff_A_tyIBQehs4_0(.dout(w_dff_A_WlOGOG2d7_0),.din(w_dff_A_tyIBQehs4_0),.clk(gclk));
	jdff dff_A_WlOGOG2d7_0(.dout(w_dff_A_hWB6KHfc7_0),.din(w_dff_A_WlOGOG2d7_0),.clk(gclk));
	jdff dff_A_hWB6KHfc7_0(.dout(w_dff_A_FAqR5UKH3_0),.din(w_dff_A_hWB6KHfc7_0),.clk(gclk));
	jdff dff_A_FAqR5UKH3_0(.dout(w_dff_A_vmz8Sacf3_0),.din(w_dff_A_FAqR5UKH3_0),.clk(gclk));
	jdff dff_A_vmz8Sacf3_0(.dout(w_dff_A_5DryWorU4_0),.din(w_dff_A_vmz8Sacf3_0),.clk(gclk));
	jdff dff_A_5DryWorU4_0(.dout(w_dff_A_kdmAfC7Z2_0),.din(w_dff_A_5DryWorU4_0),.clk(gclk));
	jdff dff_A_kdmAfC7Z2_0(.dout(w_dff_A_PDTG4Lyu3_0),.din(w_dff_A_kdmAfC7Z2_0),.clk(gclk));
	jdff dff_A_PDTG4Lyu3_0(.dout(w_dff_A_GVbLDY1S5_0),.din(w_dff_A_PDTG4Lyu3_0),.clk(gclk));
	jdff dff_A_GVbLDY1S5_0(.dout(w_dff_A_8KN4RRSD1_0),.din(w_dff_A_GVbLDY1S5_0),.clk(gclk));
	jdff dff_A_8KN4RRSD1_0(.dout(w_dff_A_f4brMCd86_0),.din(w_dff_A_8KN4RRSD1_0),.clk(gclk));
	jdff dff_A_f4brMCd86_0(.dout(w_dff_A_DEthHJvO7_0),.din(w_dff_A_f4brMCd86_0),.clk(gclk));
	jdff dff_A_DEthHJvO7_0(.dout(w_dff_A_OhHAtnqY5_0),.din(w_dff_A_DEthHJvO7_0),.clk(gclk));
	jdff dff_A_OhHAtnqY5_0(.dout(w_dff_A_cS62FSNa3_0),.din(w_dff_A_OhHAtnqY5_0),.clk(gclk));
	jdff dff_A_cS62FSNa3_0(.dout(w_dff_A_479AbONi3_0),.din(w_dff_A_cS62FSNa3_0),.clk(gclk));
	jdff dff_A_479AbONi3_0(.dout(w_dff_A_pJXoKSvf1_0),.din(w_dff_A_479AbONi3_0),.clk(gclk));
	jdff dff_A_pJXoKSvf1_0(.dout(w_dff_A_PTaAt3HY8_0),.din(w_dff_A_pJXoKSvf1_0),.clk(gclk));
	jdff dff_A_PTaAt3HY8_0(.dout(w_dff_A_C9sVdWhH5_0),.din(w_dff_A_PTaAt3HY8_0),.clk(gclk));
	jdff dff_A_C9sVdWhH5_0(.dout(w_dff_A_n8rPqkCb9_0),.din(w_dff_A_C9sVdWhH5_0),.clk(gclk));
	jdff dff_A_n8rPqkCb9_0(.dout(w_dff_A_qiCgNgwo3_0),.din(w_dff_A_n8rPqkCb9_0),.clk(gclk));
	jdff dff_A_qiCgNgwo3_0(.dout(w_dff_A_5TEwIZ6n8_0),.din(w_dff_A_qiCgNgwo3_0),.clk(gclk));
	jdff dff_A_5TEwIZ6n8_0(.dout(w_dff_A_0LSKHq6e7_0),.din(w_dff_A_5TEwIZ6n8_0),.clk(gclk));
	jdff dff_A_0LSKHq6e7_0(.dout(w_dff_A_fWBXEgeT7_0),.din(w_dff_A_0LSKHq6e7_0),.clk(gclk));
	jdff dff_A_fWBXEgeT7_0(.dout(w_dff_A_OAO0GRfY1_0),.din(w_dff_A_fWBXEgeT7_0),.clk(gclk));
	jdff dff_A_OAO0GRfY1_0(.dout(w_dff_A_uHDcmhm02_0),.din(w_dff_A_OAO0GRfY1_0),.clk(gclk));
	jdff dff_A_uHDcmhm02_0(.dout(w_dff_A_2E8jZQuZ7_0),.din(w_dff_A_uHDcmhm02_0),.clk(gclk));
	jdff dff_A_2E8jZQuZ7_0(.dout(w_dff_A_2rVGI5XN3_0),.din(w_dff_A_2E8jZQuZ7_0),.clk(gclk));
	jdff dff_A_2rVGI5XN3_0(.dout(w_dff_A_iu0JGMa19_0),.din(w_dff_A_2rVGI5XN3_0),.clk(gclk));
	jdff dff_A_iu0JGMa19_0(.dout(w_dff_A_Fjw2Ypi53_0),.din(w_dff_A_iu0JGMa19_0),.clk(gclk));
	jdff dff_A_Fjw2Ypi53_0(.dout(w_dff_A_SLd5HLax5_0),.din(w_dff_A_Fjw2Ypi53_0),.clk(gclk));
	jdff dff_A_SLd5HLax5_0(.dout(w_dff_A_kQ2WuSwu9_0),.din(w_dff_A_SLd5HLax5_0),.clk(gclk));
	jdff dff_A_kQ2WuSwu9_0(.dout(w_dff_A_RgpQF4Kq8_0),.din(w_dff_A_kQ2WuSwu9_0),.clk(gclk));
	jdff dff_A_RgpQF4Kq8_0(.dout(w_dff_A_zETwFmI94_0),.din(w_dff_A_RgpQF4Kq8_0),.clk(gclk));
	jdff dff_A_zETwFmI94_0(.dout(w_dff_A_0D30lWH01_0),.din(w_dff_A_zETwFmI94_0),.clk(gclk));
	jdff dff_A_0D30lWH01_0(.dout(w_dff_A_IfvT1kZq6_0),.din(w_dff_A_0D30lWH01_0),.clk(gclk));
	jdff dff_A_IfvT1kZq6_0(.dout(w_dff_A_pqMGsv5r8_0),.din(w_dff_A_IfvT1kZq6_0),.clk(gclk));
	jdff dff_A_pqMGsv5r8_0(.dout(w_dff_A_lkIyvNq03_0),.din(w_dff_A_pqMGsv5r8_0),.clk(gclk));
	jdff dff_A_lkIyvNq03_0(.dout(w_dff_A_4Fxy4zKq1_0),.din(w_dff_A_lkIyvNq03_0),.clk(gclk));
	jdff dff_A_4Fxy4zKq1_0(.dout(w_dff_A_TE1MwDsW3_0),.din(w_dff_A_4Fxy4zKq1_0),.clk(gclk));
	jdff dff_A_TE1MwDsW3_0(.dout(w_dff_A_okusVvoe8_0),.din(w_dff_A_TE1MwDsW3_0),.clk(gclk));
	jdff dff_A_okusVvoe8_0(.dout(w_dff_A_O0H93BUF7_0),.din(w_dff_A_okusVvoe8_0),.clk(gclk));
	jdff dff_A_O0H93BUF7_0(.dout(w_dff_A_9FL475L33_0),.din(w_dff_A_O0H93BUF7_0),.clk(gclk));
	jdff dff_A_9FL475L33_0(.dout(w_dff_A_giBoKNlS9_0),.din(w_dff_A_9FL475L33_0),.clk(gclk));
	jdff dff_A_giBoKNlS9_0(.dout(w_dff_A_M5zGQe7H2_0),.din(w_dff_A_giBoKNlS9_0),.clk(gclk));
	jdff dff_A_M5zGQe7H2_0(.dout(w_dff_A_C8dMslQp0_0),.din(w_dff_A_M5zGQe7H2_0),.clk(gclk));
	jdff dff_A_C8dMslQp0_0(.dout(w_dff_A_SSgz4MOR5_0),.din(w_dff_A_C8dMslQp0_0),.clk(gclk));
	jdff dff_A_SSgz4MOR5_0(.dout(w_dff_A_BXKlKgrx6_0),.din(w_dff_A_SSgz4MOR5_0),.clk(gclk));
	jdff dff_A_BXKlKgrx6_0(.dout(w_dff_A_P9FQj71Z8_0),.din(w_dff_A_BXKlKgrx6_0),.clk(gclk));
	jdff dff_A_P9FQj71Z8_0(.dout(w_dff_A_Yw7D2DO90_0),.din(w_dff_A_P9FQj71Z8_0),.clk(gclk));
	jdff dff_A_Yw7D2DO90_0(.dout(w_dff_A_Ooc3W83r8_0),.din(w_dff_A_Yw7D2DO90_0),.clk(gclk));
	jdff dff_A_Ooc3W83r8_0(.dout(w_dff_A_YKupuHdO1_0),.din(w_dff_A_Ooc3W83r8_0),.clk(gclk));
	jdff dff_A_YKupuHdO1_0(.dout(w_dff_A_O4BJ1L9Y0_0),.din(w_dff_A_YKupuHdO1_0),.clk(gclk));
	jdff dff_A_O4BJ1L9Y0_0(.dout(w_dff_A_IAQ9ylwU0_0),.din(w_dff_A_O4BJ1L9Y0_0),.clk(gclk));
	jdff dff_A_IAQ9ylwU0_0(.dout(w_dff_A_g58qylQv7_0),.din(w_dff_A_IAQ9ylwU0_0),.clk(gclk));
	jdff dff_A_g58qylQv7_0(.dout(w_dff_A_cmqRq9ll9_0),.din(w_dff_A_g58qylQv7_0),.clk(gclk));
	jdff dff_A_cmqRq9ll9_0(.dout(w_dff_A_fJqLOD2P9_0),.din(w_dff_A_cmqRq9ll9_0),.clk(gclk));
	jdff dff_A_fJqLOD2P9_0(.dout(w_dff_A_biog2G9A6_0),.din(w_dff_A_fJqLOD2P9_0),.clk(gclk));
	jdff dff_A_biog2G9A6_0(.dout(w_dff_A_6sZx2PC66_0),.din(w_dff_A_biog2G9A6_0),.clk(gclk));
	jdff dff_A_6sZx2PC66_0(.dout(w_dff_A_x1WcYlPQ0_0),.din(w_dff_A_6sZx2PC66_0),.clk(gclk));
	jdff dff_A_x1WcYlPQ0_0(.dout(w_dff_A_O4guebVd9_0),.din(w_dff_A_x1WcYlPQ0_0),.clk(gclk));
	jdff dff_A_O4guebVd9_0(.dout(w_dff_A_9DOVMoJo9_0),.din(w_dff_A_O4guebVd9_0),.clk(gclk));
	jdff dff_A_9DOVMoJo9_0(.dout(w_dff_A_NFWUJqb86_0),.din(w_dff_A_9DOVMoJo9_0),.clk(gclk));
	jdff dff_A_NFWUJqb86_0(.dout(w_dff_A_wHv1RlhK1_0),.din(w_dff_A_NFWUJqb86_0),.clk(gclk));
	jdff dff_A_wHv1RlhK1_0(.dout(w_dff_A_ZIxYcDhK3_0),.din(w_dff_A_wHv1RlhK1_0),.clk(gclk));
	jdff dff_A_ZIxYcDhK3_0(.dout(w_dff_A_LCoKL0Ld5_0),.din(w_dff_A_ZIxYcDhK3_0),.clk(gclk));
	jdff dff_A_LCoKL0Ld5_0(.dout(w_dff_A_kXkge0Qz3_0),.din(w_dff_A_LCoKL0Ld5_0),.clk(gclk));
	jdff dff_A_kXkge0Qz3_0(.dout(w_dff_A_ZFNKyjxw1_0),.din(w_dff_A_kXkge0Qz3_0),.clk(gclk));
	jdff dff_A_ZFNKyjxw1_0(.dout(w_dff_A_r4XED1Wz4_0),.din(w_dff_A_ZFNKyjxw1_0),.clk(gclk));
	jdff dff_A_r4XED1Wz4_0(.dout(w_dff_A_QdUAVXYu7_0),.din(w_dff_A_r4XED1Wz4_0),.clk(gclk));
	jdff dff_A_QdUAVXYu7_0(.dout(w_dff_A_KtnQqaVm6_0),.din(w_dff_A_QdUAVXYu7_0),.clk(gclk));
	jdff dff_A_KtnQqaVm6_0(.dout(w_dff_A_m6aHDcbn9_0),.din(w_dff_A_KtnQqaVm6_0),.clk(gclk));
	jdff dff_A_m6aHDcbn9_0(.dout(w_dff_A_De8Moz1T5_0),.din(w_dff_A_m6aHDcbn9_0),.clk(gclk));
	jdff dff_A_De8Moz1T5_0(.dout(w_dff_A_PanXAJOA6_0),.din(w_dff_A_De8Moz1T5_0),.clk(gclk));
	jdff dff_A_PanXAJOA6_0(.dout(w_dff_A_y90BUh0h2_0),.din(w_dff_A_PanXAJOA6_0),.clk(gclk));
	jdff dff_A_y90BUh0h2_0(.dout(w_dff_A_hF4kyPRr1_0),.din(w_dff_A_y90BUh0h2_0),.clk(gclk));
	jdff dff_A_hF4kyPRr1_0(.dout(w_dff_A_4MD2y8Ik0_0),.din(w_dff_A_hF4kyPRr1_0),.clk(gclk));
	jdff dff_A_4MD2y8Ik0_0(.dout(w_dff_A_EjK1JFvn1_0),.din(w_dff_A_4MD2y8Ik0_0),.clk(gclk));
	jdff dff_A_EjK1JFvn1_0(.dout(w_dff_A_GDqZ6AHT0_0),.din(w_dff_A_EjK1JFvn1_0),.clk(gclk));
	jdff dff_A_GDqZ6AHT0_0(.dout(w_dff_A_rA8UT6oB1_0),.din(w_dff_A_GDqZ6AHT0_0),.clk(gclk));
	jdff dff_A_rA8UT6oB1_0(.dout(w_dff_A_GHux770v4_0),.din(w_dff_A_rA8UT6oB1_0),.clk(gclk));
	jdff dff_A_GHux770v4_0(.dout(w_dff_A_fUOA2d2I4_0),.din(w_dff_A_GHux770v4_0),.clk(gclk));
	jdff dff_A_fUOA2d2I4_0(.dout(w_dff_A_3rFeyepe7_0),.din(w_dff_A_fUOA2d2I4_0),.clk(gclk));
	jdff dff_A_3rFeyepe7_0(.dout(w_dff_A_QxMgPICO1_0),.din(w_dff_A_3rFeyepe7_0),.clk(gclk));
	jdff dff_A_QxMgPICO1_0(.dout(w_dff_A_1L4XGj2E6_0),.din(w_dff_A_QxMgPICO1_0),.clk(gclk));
	jdff dff_A_1L4XGj2E6_0(.dout(w_dff_A_lzFKR7sV0_0),.din(w_dff_A_1L4XGj2E6_0),.clk(gclk));
	jdff dff_A_lzFKR7sV0_0(.dout(w_dff_A_I3oSY4fj2_0),.din(w_dff_A_lzFKR7sV0_0),.clk(gclk));
	jdff dff_A_I3oSY4fj2_0(.dout(w_dff_A_JQcrzHkQ3_0),.din(w_dff_A_I3oSY4fj2_0),.clk(gclk));
	jdff dff_A_JQcrzHkQ3_0(.dout(w_dff_A_pUp2hiZi9_0),.din(w_dff_A_JQcrzHkQ3_0),.clk(gclk));
	jdff dff_A_pUp2hiZi9_0(.dout(w_dff_A_hEbO0vre1_0),.din(w_dff_A_pUp2hiZi9_0),.clk(gclk));
	jdff dff_A_hEbO0vre1_0(.dout(w_dff_A_xUjPFYO97_0),.din(w_dff_A_hEbO0vre1_0),.clk(gclk));
	jdff dff_A_xUjPFYO97_0(.dout(w_dff_A_9N7vfbIU5_0),.din(w_dff_A_xUjPFYO97_0),.clk(gclk));
	jdff dff_A_9N7vfbIU5_0(.dout(w_dff_A_1BnerdXf2_0),.din(w_dff_A_9N7vfbIU5_0),.clk(gclk));
	jdff dff_A_1BnerdXf2_0(.dout(w_dff_A_pgrUrioX3_0),.din(w_dff_A_1BnerdXf2_0),.clk(gclk));
	jdff dff_A_pgrUrioX3_0(.dout(w_dff_A_Xjqc7oiz3_0),.din(w_dff_A_pgrUrioX3_0),.clk(gclk));
	jdff dff_A_Xjqc7oiz3_0(.dout(w_dff_A_RzMdwBna3_0),.din(w_dff_A_Xjqc7oiz3_0),.clk(gclk));
	jdff dff_A_RzMdwBna3_0(.dout(w_dff_A_d0zoPeGb8_0),.din(w_dff_A_RzMdwBna3_0),.clk(gclk));
	jdff dff_A_d0zoPeGb8_0(.dout(w_dff_A_kPT4fht42_0),.din(w_dff_A_d0zoPeGb8_0),.clk(gclk));
	jdff dff_A_kPT4fht42_0(.dout(w_dff_A_a2phIt3T8_0),.din(w_dff_A_kPT4fht42_0),.clk(gclk));
	jdff dff_A_a2phIt3T8_0(.dout(w_dff_A_g3gFHxxZ7_0),.din(w_dff_A_a2phIt3T8_0),.clk(gclk));
	jdff dff_A_g3gFHxxZ7_0(.dout(w_dff_A_gR2LLfUO8_0),.din(w_dff_A_g3gFHxxZ7_0),.clk(gclk));
	jdff dff_A_gR2LLfUO8_0(.dout(w_dff_A_akm2I8wf7_0),.din(w_dff_A_gR2LLfUO8_0),.clk(gclk));
	jdff dff_A_akm2I8wf7_0(.dout(f22),.din(w_dff_A_akm2I8wf7_0),.clk(gclk));
	jdff dff_A_SzoSoT3h7_2(.dout(w_dff_A_LXu8MeCK4_0),.din(w_dff_A_SzoSoT3h7_2),.clk(gclk));
	jdff dff_A_LXu8MeCK4_0(.dout(w_dff_A_PVWHarOq6_0),.din(w_dff_A_LXu8MeCK4_0),.clk(gclk));
	jdff dff_A_PVWHarOq6_0(.dout(w_dff_A_vifkcGun8_0),.din(w_dff_A_PVWHarOq6_0),.clk(gclk));
	jdff dff_A_vifkcGun8_0(.dout(w_dff_A_MdeSnA3n3_0),.din(w_dff_A_vifkcGun8_0),.clk(gclk));
	jdff dff_A_MdeSnA3n3_0(.dout(w_dff_A_vqkNSrdK9_0),.din(w_dff_A_MdeSnA3n3_0),.clk(gclk));
	jdff dff_A_vqkNSrdK9_0(.dout(w_dff_A_mF9lCjQ08_0),.din(w_dff_A_vqkNSrdK9_0),.clk(gclk));
	jdff dff_A_mF9lCjQ08_0(.dout(w_dff_A_Iyd8w0tZ1_0),.din(w_dff_A_mF9lCjQ08_0),.clk(gclk));
	jdff dff_A_Iyd8w0tZ1_0(.dout(w_dff_A_TeFjgyX76_0),.din(w_dff_A_Iyd8w0tZ1_0),.clk(gclk));
	jdff dff_A_TeFjgyX76_0(.dout(w_dff_A_YHZd3Amb7_0),.din(w_dff_A_TeFjgyX76_0),.clk(gclk));
	jdff dff_A_YHZd3Amb7_0(.dout(w_dff_A_GIadcR8T8_0),.din(w_dff_A_YHZd3Amb7_0),.clk(gclk));
	jdff dff_A_GIadcR8T8_0(.dout(w_dff_A_dtlDCxQZ1_0),.din(w_dff_A_GIadcR8T8_0),.clk(gclk));
	jdff dff_A_dtlDCxQZ1_0(.dout(w_dff_A_xpG3ulbz0_0),.din(w_dff_A_dtlDCxQZ1_0),.clk(gclk));
	jdff dff_A_xpG3ulbz0_0(.dout(w_dff_A_imuh9k5R6_0),.din(w_dff_A_xpG3ulbz0_0),.clk(gclk));
	jdff dff_A_imuh9k5R6_0(.dout(w_dff_A_IfgThEwV6_0),.din(w_dff_A_imuh9k5R6_0),.clk(gclk));
	jdff dff_A_IfgThEwV6_0(.dout(w_dff_A_IRrpS1iv1_0),.din(w_dff_A_IfgThEwV6_0),.clk(gclk));
	jdff dff_A_IRrpS1iv1_0(.dout(w_dff_A_jD2jZJ493_0),.din(w_dff_A_IRrpS1iv1_0),.clk(gclk));
	jdff dff_A_jD2jZJ493_0(.dout(w_dff_A_p1HjCQLw3_0),.din(w_dff_A_jD2jZJ493_0),.clk(gclk));
	jdff dff_A_p1HjCQLw3_0(.dout(w_dff_A_jCV2xufZ5_0),.din(w_dff_A_p1HjCQLw3_0),.clk(gclk));
	jdff dff_A_jCV2xufZ5_0(.dout(w_dff_A_qykpVwGV0_0),.din(w_dff_A_jCV2xufZ5_0),.clk(gclk));
	jdff dff_A_qykpVwGV0_0(.dout(w_dff_A_qB5FPRrW5_0),.din(w_dff_A_qykpVwGV0_0),.clk(gclk));
	jdff dff_A_qB5FPRrW5_0(.dout(w_dff_A_owfNYa9D9_0),.din(w_dff_A_qB5FPRrW5_0),.clk(gclk));
	jdff dff_A_owfNYa9D9_0(.dout(w_dff_A_mIU6Bse73_0),.din(w_dff_A_owfNYa9D9_0),.clk(gclk));
	jdff dff_A_mIU6Bse73_0(.dout(w_dff_A_2DbPMeuB7_0),.din(w_dff_A_mIU6Bse73_0),.clk(gclk));
	jdff dff_A_2DbPMeuB7_0(.dout(w_dff_A_bW4x1qXE8_0),.din(w_dff_A_2DbPMeuB7_0),.clk(gclk));
	jdff dff_A_bW4x1qXE8_0(.dout(w_dff_A_bY11Q5mg8_0),.din(w_dff_A_bW4x1qXE8_0),.clk(gclk));
	jdff dff_A_bY11Q5mg8_0(.dout(w_dff_A_BAEbRGrc1_0),.din(w_dff_A_bY11Q5mg8_0),.clk(gclk));
	jdff dff_A_BAEbRGrc1_0(.dout(w_dff_A_ASg1x7au3_0),.din(w_dff_A_BAEbRGrc1_0),.clk(gclk));
	jdff dff_A_ASg1x7au3_0(.dout(w_dff_A_gDgu3THB4_0),.din(w_dff_A_ASg1x7au3_0),.clk(gclk));
	jdff dff_A_gDgu3THB4_0(.dout(w_dff_A_BDvUB8TI5_0),.din(w_dff_A_gDgu3THB4_0),.clk(gclk));
	jdff dff_A_BDvUB8TI5_0(.dout(w_dff_A_jYfVz6oW2_0),.din(w_dff_A_BDvUB8TI5_0),.clk(gclk));
	jdff dff_A_jYfVz6oW2_0(.dout(w_dff_A_a8l5C6Ap1_0),.din(w_dff_A_jYfVz6oW2_0),.clk(gclk));
	jdff dff_A_a8l5C6Ap1_0(.dout(w_dff_A_8R47zttB4_0),.din(w_dff_A_a8l5C6Ap1_0),.clk(gclk));
	jdff dff_A_8R47zttB4_0(.dout(w_dff_A_G4aae9Zw2_0),.din(w_dff_A_8R47zttB4_0),.clk(gclk));
	jdff dff_A_G4aae9Zw2_0(.dout(w_dff_A_sW7Q7Knw0_0),.din(w_dff_A_G4aae9Zw2_0),.clk(gclk));
	jdff dff_A_sW7Q7Knw0_0(.dout(w_dff_A_2JXXtMpv3_0),.din(w_dff_A_sW7Q7Knw0_0),.clk(gclk));
	jdff dff_A_2JXXtMpv3_0(.dout(w_dff_A_kJ7juJXl2_0),.din(w_dff_A_2JXXtMpv3_0),.clk(gclk));
	jdff dff_A_kJ7juJXl2_0(.dout(w_dff_A_wxOnMeeI0_0),.din(w_dff_A_kJ7juJXl2_0),.clk(gclk));
	jdff dff_A_wxOnMeeI0_0(.dout(w_dff_A_ODt5AzzS7_0),.din(w_dff_A_wxOnMeeI0_0),.clk(gclk));
	jdff dff_A_ODt5AzzS7_0(.dout(w_dff_A_KcJqTdHP8_0),.din(w_dff_A_ODt5AzzS7_0),.clk(gclk));
	jdff dff_A_KcJqTdHP8_0(.dout(w_dff_A_kWPWQpGd3_0),.din(w_dff_A_KcJqTdHP8_0),.clk(gclk));
	jdff dff_A_kWPWQpGd3_0(.dout(w_dff_A_3TjJOnOC7_0),.din(w_dff_A_kWPWQpGd3_0),.clk(gclk));
	jdff dff_A_3TjJOnOC7_0(.dout(w_dff_A_sgXkth8x3_0),.din(w_dff_A_3TjJOnOC7_0),.clk(gclk));
	jdff dff_A_sgXkth8x3_0(.dout(w_dff_A_7eD9rVRi0_0),.din(w_dff_A_sgXkth8x3_0),.clk(gclk));
	jdff dff_A_7eD9rVRi0_0(.dout(w_dff_A_4cms8jLp0_0),.din(w_dff_A_7eD9rVRi0_0),.clk(gclk));
	jdff dff_A_4cms8jLp0_0(.dout(w_dff_A_KWhctdji3_0),.din(w_dff_A_4cms8jLp0_0),.clk(gclk));
	jdff dff_A_KWhctdji3_0(.dout(w_dff_A_QBDjBpOu8_0),.din(w_dff_A_KWhctdji3_0),.clk(gclk));
	jdff dff_A_QBDjBpOu8_0(.dout(w_dff_A_TgFxIp3s3_0),.din(w_dff_A_QBDjBpOu8_0),.clk(gclk));
	jdff dff_A_TgFxIp3s3_0(.dout(w_dff_A_6iBUmoJf0_0),.din(w_dff_A_TgFxIp3s3_0),.clk(gclk));
	jdff dff_A_6iBUmoJf0_0(.dout(w_dff_A_aejISBg08_0),.din(w_dff_A_6iBUmoJf0_0),.clk(gclk));
	jdff dff_A_aejISBg08_0(.dout(w_dff_A_uOcqpVc64_0),.din(w_dff_A_aejISBg08_0),.clk(gclk));
	jdff dff_A_uOcqpVc64_0(.dout(w_dff_A_ArBlX3jn0_0),.din(w_dff_A_uOcqpVc64_0),.clk(gclk));
	jdff dff_A_ArBlX3jn0_0(.dout(w_dff_A_klpiuytj8_0),.din(w_dff_A_ArBlX3jn0_0),.clk(gclk));
	jdff dff_A_klpiuytj8_0(.dout(w_dff_A_o56JiOSW0_0),.din(w_dff_A_klpiuytj8_0),.clk(gclk));
	jdff dff_A_o56JiOSW0_0(.dout(w_dff_A_gyPJsgey1_0),.din(w_dff_A_o56JiOSW0_0),.clk(gclk));
	jdff dff_A_gyPJsgey1_0(.dout(w_dff_A_kWZIIHBJ2_0),.din(w_dff_A_gyPJsgey1_0),.clk(gclk));
	jdff dff_A_kWZIIHBJ2_0(.dout(w_dff_A_IpEj3raU0_0),.din(w_dff_A_kWZIIHBJ2_0),.clk(gclk));
	jdff dff_A_IpEj3raU0_0(.dout(w_dff_A_YmNhCS0B9_0),.din(w_dff_A_IpEj3raU0_0),.clk(gclk));
	jdff dff_A_YmNhCS0B9_0(.dout(w_dff_A_CCATSn5H4_0),.din(w_dff_A_YmNhCS0B9_0),.clk(gclk));
	jdff dff_A_CCATSn5H4_0(.dout(w_dff_A_CGOYnW5O9_0),.din(w_dff_A_CCATSn5H4_0),.clk(gclk));
	jdff dff_A_CGOYnW5O9_0(.dout(w_dff_A_7LiUCqHo5_0),.din(w_dff_A_CGOYnW5O9_0),.clk(gclk));
	jdff dff_A_7LiUCqHo5_0(.dout(w_dff_A_9sODmkT92_0),.din(w_dff_A_7LiUCqHo5_0),.clk(gclk));
	jdff dff_A_9sODmkT92_0(.dout(w_dff_A_7KUhGUFr0_0),.din(w_dff_A_9sODmkT92_0),.clk(gclk));
	jdff dff_A_7KUhGUFr0_0(.dout(w_dff_A_oi1zJ8CS5_0),.din(w_dff_A_7KUhGUFr0_0),.clk(gclk));
	jdff dff_A_oi1zJ8CS5_0(.dout(w_dff_A_eKZGL1246_0),.din(w_dff_A_oi1zJ8CS5_0),.clk(gclk));
	jdff dff_A_eKZGL1246_0(.dout(w_dff_A_FsmKzGuw4_0),.din(w_dff_A_eKZGL1246_0),.clk(gclk));
	jdff dff_A_FsmKzGuw4_0(.dout(w_dff_A_AFrjmDBM4_0),.din(w_dff_A_FsmKzGuw4_0),.clk(gclk));
	jdff dff_A_AFrjmDBM4_0(.dout(w_dff_A_Gw0mfJZS8_0),.din(w_dff_A_AFrjmDBM4_0),.clk(gclk));
	jdff dff_A_Gw0mfJZS8_0(.dout(w_dff_A_6tpPbB2I3_0),.din(w_dff_A_Gw0mfJZS8_0),.clk(gclk));
	jdff dff_A_6tpPbB2I3_0(.dout(w_dff_A_0lWJ2Xti3_0),.din(w_dff_A_6tpPbB2I3_0),.clk(gclk));
	jdff dff_A_0lWJ2Xti3_0(.dout(w_dff_A_t4W4Gd1K1_0),.din(w_dff_A_0lWJ2Xti3_0),.clk(gclk));
	jdff dff_A_t4W4Gd1K1_0(.dout(w_dff_A_iyPVEQDl4_0),.din(w_dff_A_t4W4Gd1K1_0),.clk(gclk));
	jdff dff_A_iyPVEQDl4_0(.dout(w_dff_A_QZ18hAHR0_0),.din(w_dff_A_iyPVEQDl4_0),.clk(gclk));
	jdff dff_A_QZ18hAHR0_0(.dout(w_dff_A_2DG7GwYF4_0),.din(w_dff_A_QZ18hAHR0_0),.clk(gclk));
	jdff dff_A_2DG7GwYF4_0(.dout(w_dff_A_VoWJFzLW5_0),.din(w_dff_A_2DG7GwYF4_0),.clk(gclk));
	jdff dff_A_VoWJFzLW5_0(.dout(w_dff_A_zkdlMpUx4_0),.din(w_dff_A_VoWJFzLW5_0),.clk(gclk));
	jdff dff_A_zkdlMpUx4_0(.dout(w_dff_A_3OQZIldj0_0),.din(w_dff_A_zkdlMpUx4_0),.clk(gclk));
	jdff dff_A_3OQZIldj0_0(.dout(w_dff_A_4z0tI5rq0_0),.din(w_dff_A_3OQZIldj0_0),.clk(gclk));
	jdff dff_A_4z0tI5rq0_0(.dout(w_dff_A_vPiJCUxB6_0),.din(w_dff_A_4z0tI5rq0_0),.clk(gclk));
	jdff dff_A_vPiJCUxB6_0(.dout(w_dff_A_funNv0lY2_0),.din(w_dff_A_vPiJCUxB6_0),.clk(gclk));
	jdff dff_A_funNv0lY2_0(.dout(w_dff_A_6M6BaDUw3_0),.din(w_dff_A_funNv0lY2_0),.clk(gclk));
	jdff dff_A_6M6BaDUw3_0(.dout(w_dff_A_CoDM5QjP2_0),.din(w_dff_A_6M6BaDUw3_0),.clk(gclk));
	jdff dff_A_CoDM5QjP2_0(.dout(w_dff_A_EYDQ1SN71_0),.din(w_dff_A_CoDM5QjP2_0),.clk(gclk));
	jdff dff_A_EYDQ1SN71_0(.dout(w_dff_A_ekhQo3kf1_0),.din(w_dff_A_EYDQ1SN71_0),.clk(gclk));
	jdff dff_A_ekhQo3kf1_0(.dout(w_dff_A_RynvRZny4_0),.din(w_dff_A_ekhQo3kf1_0),.clk(gclk));
	jdff dff_A_RynvRZny4_0(.dout(w_dff_A_TKbnUnwF1_0),.din(w_dff_A_RynvRZny4_0),.clk(gclk));
	jdff dff_A_TKbnUnwF1_0(.dout(w_dff_A_WTAQeAF97_0),.din(w_dff_A_TKbnUnwF1_0),.clk(gclk));
	jdff dff_A_WTAQeAF97_0(.dout(w_dff_A_mnZVhNVH6_0),.din(w_dff_A_WTAQeAF97_0),.clk(gclk));
	jdff dff_A_mnZVhNVH6_0(.dout(w_dff_A_QQcMw8Fl8_0),.din(w_dff_A_mnZVhNVH6_0),.clk(gclk));
	jdff dff_A_QQcMw8Fl8_0(.dout(w_dff_A_HTZAA6WZ7_0),.din(w_dff_A_QQcMw8Fl8_0),.clk(gclk));
	jdff dff_A_HTZAA6WZ7_0(.dout(w_dff_A_1OmNtLNt8_0),.din(w_dff_A_HTZAA6WZ7_0),.clk(gclk));
	jdff dff_A_1OmNtLNt8_0(.dout(w_dff_A_8xAFlvmf0_0),.din(w_dff_A_1OmNtLNt8_0),.clk(gclk));
	jdff dff_A_8xAFlvmf0_0(.dout(w_dff_A_xWTpfVgj4_0),.din(w_dff_A_8xAFlvmf0_0),.clk(gclk));
	jdff dff_A_xWTpfVgj4_0(.dout(w_dff_A_GLwGk8Zm5_0),.din(w_dff_A_xWTpfVgj4_0),.clk(gclk));
	jdff dff_A_GLwGk8Zm5_0(.dout(w_dff_A_UjABIs6o9_0),.din(w_dff_A_GLwGk8Zm5_0),.clk(gclk));
	jdff dff_A_UjABIs6o9_0(.dout(w_dff_A_jhWgGv0K1_0),.din(w_dff_A_UjABIs6o9_0),.clk(gclk));
	jdff dff_A_jhWgGv0K1_0(.dout(w_dff_A_DWIOOwgf4_0),.din(w_dff_A_jhWgGv0K1_0),.clk(gclk));
	jdff dff_A_DWIOOwgf4_0(.dout(w_dff_A_wAvlJOGm1_0),.din(w_dff_A_DWIOOwgf4_0),.clk(gclk));
	jdff dff_A_wAvlJOGm1_0(.dout(w_dff_A_3DiWJpNI4_0),.din(w_dff_A_wAvlJOGm1_0),.clk(gclk));
	jdff dff_A_3DiWJpNI4_0(.dout(w_dff_A_Si5NIZHx2_0),.din(w_dff_A_3DiWJpNI4_0),.clk(gclk));
	jdff dff_A_Si5NIZHx2_0(.dout(w_dff_A_HHgAH7bn6_0),.din(w_dff_A_Si5NIZHx2_0),.clk(gclk));
	jdff dff_A_HHgAH7bn6_0(.dout(w_dff_A_fKfOJnKl3_0),.din(w_dff_A_HHgAH7bn6_0),.clk(gclk));
	jdff dff_A_fKfOJnKl3_0(.dout(w_dff_A_Aun1bA194_0),.din(w_dff_A_fKfOJnKl3_0),.clk(gclk));
	jdff dff_A_Aun1bA194_0(.dout(w_dff_A_VMJTXdB51_0),.din(w_dff_A_Aun1bA194_0),.clk(gclk));
	jdff dff_A_VMJTXdB51_0(.dout(f23),.din(w_dff_A_VMJTXdB51_0),.clk(gclk));
	jdff dff_A_ejqy7DXE0_2(.dout(w_dff_A_W9qGWd5L5_0),.din(w_dff_A_ejqy7DXE0_2),.clk(gclk));
	jdff dff_A_W9qGWd5L5_0(.dout(w_dff_A_ggFuGkP97_0),.din(w_dff_A_W9qGWd5L5_0),.clk(gclk));
	jdff dff_A_ggFuGkP97_0(.dout(w_dff_A_BVcr5RcT9_0),.din(w_dff_A_ggFuGkP97_0),.clk(gclk));
	jdff dff_A_BVcr5RcT9_0(.dout(w_dff_A_PNMtgzvZ3_0),.din(w_dff_A_BVcr5RcT9_0),.clk(gclk));
	jdff dff_A_PNMtgzvZ3_0(.dout(w_dff_A_9EZohE6J0_0),.din(w_dff_A_PNMtgzvZ3_0),.clk(gclk));
	jdff dff_A_9EZohE6J0_0(.dout(w_dff_A_Y7RBP92s3_0),.din(w_dff_A_9EZohE6J0_0),.clk(gclk));
	jdff dff_A_Y7RBP92s3_0(.dout(w_dff_A_lWHrxWO81_0),.din(w_dff_A_Y7RBP92s3_0),.clk(gclk));
	jdff dff_A_lWHrxWO81_0(.dout(w_dff_A_1sFEfer31_0),.din(w_dff_A_lWHrxWO81_0),.clk(gclk));
	jdff dff_A_1sFEfer31_0(.dout(w_dff_A_ViTw3MGF1_0),.din(w_dff_A_1sFEfer31_0),.clk(gclk));
	jdff dff_A_ViTw3MGF1_0(.dout(w_dff_A_kymaJul48_0),.din(w_dff_A_ViTw3MGF1_0),.clk(gclk));
	jdff dff_A_kymaJul48_0(.dout(w_dff_A_fUzRDZZ14_0),.din(w_dff_A_kymaJul48_0),.clk(gclk));
	jdff dff_A_fUzRDZZ14_0(.dout(w_dff_A_QK7TvgVu8_0),.din(w_dff_A_fUzRDZZ14_0),.clk(gclk));
	jdff dff_A_QK7TvgVu8_0(.dout(w_dff_A_KOdloJ791_0),.din(w_dff_A_QK7TvgVu8_0),.clk(gclk));
	jdff dff_A_KOdloJ791_0(.dout(w_dff_A_L7sNwnTe5_0),.din(w_dff_A_KOdloJ791_0),.clk(gclk));
	jdff dff_A_L7sNwnTe5_0(.dout(w_dff_A_MuG62oUz0_0),.din(w_dff_A_L7sNwnTe5_0),.clk(gclk));
	jdff dff_A_MuG62oUz0_0(.dout(w_dff_A_dRlNogGM5_0),.din(w_dff_A_MuG62oUz0_0),.clk(gclk));
	jdff dff_A_dRlNogGM5_0(.dout(w_dff_A_X46SUInS2_0),.din(w_dff_A_dRlNogGM5_0),.clk(gclk));
	jdff dff_A_X46SUInS2_0(.dout(w_dff_A_xZYRmbfw9_0),.din(w_dff_A_X46SUInS2_0),.clk(gclk));
	jdff dff_A_xZYRmbfw9_0(.dout(w_dff_A_LYTxWNRW4_0),.din(w_dff_A_xZYRmbfw9_0),.clk(gclk));
	jdff dff_A_LYTxWNRW4_0(.dout(w_dff_A_bf0aTqXI7_0),.din(w_dff_A_LYTxWNRW4_0),.clk(gclk));
	jdff dff_A_bf0aTqXI7_0(.dout(w_dff_A_aCxSvOX66_0),.din(w_dff_A_bf0aTqXI7_0),.clk(gclk));
	jdff dff_A_aCxSvOX66_0(.dout(w_dff_A_cIsj3QxJ3_0),.din(w_dff_A_aCxSvOX66_0),.clk(gclk));
	jdff dff_A_cIsj3QxJ3_0(.dout(w_dff_A_J9hs0yzB5_0),.din(w_dff_A_cIsj3QxJ3_0),.clk(gclk));
	jdff dff_A_J9hs0yzB5_0(.dout(w_dff_A_vQAFlWTx8_0),.din(w_dff_A_J9hs0yzB5_0),.clk(gclk));
	jdff dff_A_vQAFlWTx8_0(.dout(w_dff_A_m3L4hsq31_0),.din(w_dff_A_vQAFlWTx8_0),.clk(gclk));
	jdff dff_A_m3L4hsq31_0(.dout(w_dff_A_KtCpX6E49_0),.din(w_dff_A_m3L4hsq31_0),.clk(gclk));
	jdff dff_A_KtCpX6E49_0(.dout(w_dff_A_Fx8sSX2J7_0),.din(w_dff_A_KtCpX6E49_0),.clk(gclk));
	jdff dff_A_Fx8sSX2J7_0(.dout(w_dff_A_0aKUwqfo4_0),.din(w_dff_A_Fx8sSX2J7_0),.clk(gclk));
	jdff dff_A_0aKUwqfo4_0(.dout(w_dff_A_rUdDsgZT2_0),.din(w_dff_A_0aKUwqfo4_0),.clk(gclk));
	jdff dff_A_rUdDsgZT2_0(.dout(w_dff_A_ZzRGaad17_0),.din(w_dff_A_rUdDsgZT2_0),.clk(gclk));
	jdff dff_A_ZzRGaad17_0(.dout(w_dff_A_hyzJehtM7_0),.din(w_dff_A_ZzRGaad17_0),.clk(gclk));
	jdff dff_A_hyzJehtM7_0(.dout(w_dff_A_FVIX3Ia43_0),.din(w_dff_A_hyzJehtM7_0),.clk(gclk));
	jdff dff_A_FVIX3Ia43_0(.dout(w_dff_A_bI80vFUL4_0),.din(w_dff_A_FVIX3Ia43_0),.clk(gclk));
	jdff dff_A_bI80vFUL4_0(.dout(w_dff_A_WwcYynn03_0),.din(w_dff_A_bI80vFUL4_0),.clk(gclk));
	jdff dff_A_WwcYynn03_0(.dout(w_dff_A_3SeYvBSO4_0),.din(w_dff_A_WwcYynn03_0),.clk(gclk));
	jdff dff_A_3SeYvBSO4_0(.dout(w_dff_A_dvq20nJy5_0),.din(w_dff_A_3SeYvBSO4_0),.clk(gclk));
	jdff dff_A_dvq20nJy5_0(.dout(w_dff_A_V0TiymFn5_0),.din(w_dff_A_dvq20nJy5_0),.clk(gclk));
	jdff dff_A_V0TiymFn5_0(.dout(w_dff_A_InSpKmGW0_0),.din(w_dff_A_V0TiymFn5_0),.clk(gclk));
	jdff dff_A_InSpKmGW0_0(.dout(w_dff_A_vKNoR8dw6_0),.din(w_dff_A_InSpKmGW0_0),.clk(gclk));
	jdff dff_A_vKNoR8dw6_0(.dout(w_dff_A_bgz3aLVs5_0),.din(w_dff_A_vKNoR8dw6_0),.clk(gclk));
	jdff dff_A_bgz3aLVs5_0(.dout(w_dff_A_33If5CeM2_0),.din(w_dff_A_bgz3aLVs5_0),.clk(gclk));
	jdff dff_A_33If5CeM2_0(.dout(w_dff_A_Yl1H3zSP4_0),.din(w_dff_A_33If5CeM2_0),.clk(gclk));
	jdff dff_A_Yl1H3zSP4_0(.dout(w_dff_A_YSGDg2aq6_0),.din(w_dff_A_Yl1H3zSP4_0),.clk(gclk));
	jdff dff_A_YSGDg2aq6_0(.dout(w_dff_A_yRgScSfz9_0),.din(w_dff_A_YSGDg2aq6_0),.clk(gclk));
	jdff dff_A_yRgScSfz9_0(.dout(w_dff_A_emNbOSB58_0),.din(w_dff_A_yRgScSfz9_0),.clk(gclk));
	jdff dff_A_emNbOSB58_0(.dout(w_dff_A_0joguT0n8_0),.din(w_dff_A_emNbOSB58_0),.clk(gclk));
	jdff dff_A_0joguT0n8_0(.dout(w_dff_A_e95w1D3H2_0),.din(w_dff_A_0joguT0n8_0),.clk(gclk));
	jdff dff_A_e95w1D3H2_0(.dout(w_dff_A_7oxaZ6G89_0),.din(w_dff_A_e95w1D3H2_0),.clk(gclk));
	jdff dff_A_7oxaZ6G89_0(.dout(w_dff_A_PsMZRVYY6_0),.din(w_dff_A_7oxaZ6G89_0),.clk(gclk));
	jdff dff_A_PsMZRVYY6_0(.dout(w_dff_A_3jfRZvRo2_0),.din(w_dff_A_PsMZRVYY6_0),.clk(gclk));
	jdff dff_A_3jfRZvRo2_0(.dout(w_dff_A_L1gTztii4_0),.din(w_dff_A_3jfRZvRo2_0),.clk(gclk));
	jdff dff_A_L1gTztii4_0(.dout(w_dff_A_mZvLRIe05_0),.din(w_dff_A_L1gTztii4_0),.clk(gclk));
	jdff dff_A_mZvLRIe05_0(.dout(w_dff_A_2zqT3RIj3_0),.din(w_dff_A_mZvLRIe05_0),.clk(gclk));
	jdff dff_A_2zqT3RIj3_0(.dout(w_dff_A_bwyy7mFv5_0),.din(w_dff_A_2zqT3RIj3_0),.clk(gclk));
	jdff dff_A_bwyy7mFv5_0(.dout(w_dff_A_QiJKv5Qp0_0),.din(w_dff_A_bwyy7mFv5_0),.clk(gclk));
	jdff dff_A_QiJKv5Qp0_0(.dout(w_dff_A_bc5x8CLy1_0),.din(w_dff_A_QiJKv5Qp0_0),.clk(gclk));
	jdff dff_A_bc5x8CLy1_0(.dout(w_dff_A_CYhoSLiY4_0),.din(w_dff_A_bc5x8CLy1_0),.clk(gclk));
	jdff dff_A_CYhoSLiY4_0(.dout(w_dff_A_H1dQJ4ez0_0),.din(w_dff_A_CYhoSLiY4_0),.clk(gclk));
	jdff dff_A_H1dQJ4ez0_0(.dout(w_dff_A_IFsKeohE3_0),.din(w_dff_A_H1dQJ4ez0_0),.clk(gclk));
	jdff dff_A_IFsKeohE3_0(.dout(w_dff_A_ouXkB9Sb2_0),.din(w_dff_A_IFsKeohE3_0),.clk(gclk));
	jdff dff_A_ouXkB9Sb2_0(.dout(w_dff_A_V0XTjOvB4_0),.din(w_dff_A_ouXkB9Sb2_0),.clk(gclk));
	jdff dff_A_V0XTjOvB4_0(.dout(w_dff_A_k1r1iZuP7_0),.din(w_dff_A_V0XTjOvB4_0),.clk(gclk));
	jdff dff_A_k1r1iZuP7_0(.dout(w_dff_A_7RQ14DhJ7_0),.din(w_dff_A_k1r1iZuP7_0),.clk(gclk));
	jdff dff_A_7RQ14DhJ7_0(.dout(w_dff_A_8iuAEy5I8_0),.din(w_dff_A_7RQ14DhJ7_0),.clk(gclk));
	jdff dff_A_8iuAEy5I8_0(.dout(w_dff_A_RHyheddQ1_0),.din(w_dff_A_8iuAEy5I8_0),.clk(gclk));
	jdff dff_A_RHyheddQ1_0(.dout(w_dff_A_e8wzgcAC0_0),.din(w_dff_A_RHyheddQ1_0),.clk(gclk));
	jdff dff_A_e8wzgcAC0_0(.dout(w_dff_A_vkPOIoEu2_0),.din(w_dff_A_e8wzgcAC0_0),.clk(gclk));
	jdff dff_A_vkPOIoEu2_0(.dout(w_dff_A_LnAJKT816_0),.din(w_dff_A_vkPOIoEu2_0),.clk(gclk));
	jdff dff_A_LnAJKT816_0(.dout(w_dff_A_ZaC6eVBr4_0),.din(w_dff_A_LnAJKT816_0),.clk(gclk));
	jdff dff_A_ZaC6eVBr4_0(.dout(w_dff_A_EWZwgFVi5_0),.din(w_dff_A_ZaC6eVBr4_0),.clk(gclk));
	jdff dff_A_EWZwgFVi5_0(.dout(w_dff_A_DhLQcXRh7_0),.din(w_dff_A_EWZwgFVi5_0),.clk(gclk));
	jdff dff_A_DhLQcXRh7_0(.dout(w_dff_A_2V8rt1eX1_0),.din(w_dff_A_DhLQcXRh7_0),.clk(gclk));
	jdff dff_A_2V8rt1eX1_0(.dout(w_dff_A_98aflCDi5_0),.din(w_dff_A_2V8rt1eX1_0),.clk(gclk));
	jdff dff_A_98aflCDi5_0(.dout(w_dff_A_qf0SAwA50_0),.din(w_dff_A_98aflCDi5_0),.clk(gclk));
	jdff dff_A_qf0SAwA50_0(.dout(w_dff_A_vtUIdmVH0_0),.din(w_dff_A_qf0SAwA50_0),.clk(gclk));
	jdff dff_A_vtUIdmVH0_0(.dout(w_dff_A_4KwMGY9a7_0),.din(w_dff_A_vtUIdmVH0_0),.clk(gclk));
	jdff dff_A_4KwMGY9a7_0(.dout(w_dff_A_aBb5MOyb7_0),.din(w_dff_A_4KwMGY9a7_0),.clk(gclk));
	jdff dff_A_aBb5MOyb7_0(.dout(w_dff_A_DD5cBLyN5_0),.din(w_dff_A_aBb5MOyb7_0),.clk(gclk));
	jdff dff_A_DD5cBLyN5_0(.dout(w_dff_A_Lg4EKZAv1_0),.din(w_dff_A_DD5cBLyN5_0),.clk(gclk));
	jdff dff_A_Lg4EKZAv1_0(.dout(w_dff_A_NkcCgnAP7_0),.din(w_dff_A_Lg4EKZAv1_0),.clk(gclk));
	jdff dff_A_NkcCgnAP7_0(.dout(w_dff_A_uQb8QUWy7_0),.din(w_dff_A_NkcCgnAP7_0),.clk(gclk));
	jdff dff_A_uQb8QUWy7_0(.dout(w_dff_A_S4Zgh2Bs1_0),.din(w_dff_A_uQb8QUWy7_0),.clk(gclk));
	jdff dff_A_S4Zgh2Bs1_0(.dout(w_dff_A_K7UdTQ9A0_0),.din(w_dff_A_S4Zgh2Bs1_0),.clk(gclk));
	jdff dff_A_K7UdTQ9A0_0(.dout(w_dff_A_HirujnNS7_0),.din(w_dff_A_K7UdTQ9A0_0),.clk(gclk));
	jdff dff_A_HirujnNS7_0(.dout(w_dff_A_ZVRApH6F5_0),.din(w_dff_A_HirujnNS7_0),.clk(gclk));
	jdff dff_A_ZVRApH6F5_0(.dout(w_dff_A_UqiPodn99_0),.din(w_dff_A_ZVRApH6F5_0),.clk(gclk));
	jdff dff_A_UqiPodn99_0(.dout(w_dff_A_Isp1yFap2_0),.din(w_dff_A_UqiPodn99_0),.clk(gclk));
	jdff dff_A_Isp1yFap2_0(.dout(w_dff_A_n6pbBf6Z1_0),.din(w_dff_A_Isp1yFap2_0),.clk(gclk));
	jdff dff_A_n6pbBf6Z1_0(.dout(w_dff_A_EH6GaQiO8_0),.din(w_dff_A_n6pbBf6Z1_0),.clk(gclk));
	jdff dff_A_EH6GaQiO8_0(.dout(w_dff_A_B6MKY3l67_0),.din(w_dff_A_EH6GaQiO8_0),.clk(gclk));
	jdff dff_A_B6MKY3l67_0(.dout(w_dff_A_Rxo852FK5_0),.din(w_dff_A_B6MKY3l67_0),.clk(gclk));
	jdff dff_A_Rxo852FK5_0(.dout(w_dff_A_2k5F1CB89_0),.din(w_dff_A_Rxo852FK5_0),.clk(gclk));
	jdff dff_A_2k5F1CB89_0(.dout(w_dff_A_tJBO9hAc8_0),.din(w_dff_A_2k5F1CB89_0),.clk(gclk));
	jdff dff_A_tJBO9hAc8_0(.dout(w_dff_A_oNekGLhW2_0),.din(w_dff_A_tJBO9hAc8_0),.clk(gclk));
	jdff dff_A_oNekGLhW2_0(.dout(w_dff_A_Ao97cxID1_0),.din(w_dff_A_oNekGLhW2_0),.clk(gclk));
	jdff dff_A_Ao97cxID1_0(.dout(w_dff_A_I8fmg2eM1_0),.din(w_dff_A_Ao97cxID1_0),.clk(gclk));
	jdff dff_A_I8fmg2eM1_0(.dout(w_dff_A_Byqdnubd4_0),.din(w_dff_A_I8fmg2eM1_0),.clk(gclk));
	jdff dff_A_Byqdnubd4_0(.dout(w_dff_A_jRUa5FoK4_0),.din(w_dff_A_Byqdnubd4_0),.clk(gclk));
	jdff dff_A_jRUa5FoK4_0(.dout(w_dff_A_ymB7fdEt0_0),.din(w_dff_A_jRUa5FoK4_0),.clk(gclk));
	jdff dff_A_ymB7fdEt0_0(.dout(w_dff_A_uKaxxzL60_0),.din(w_dff_A_ymB7fdEt0_0),.clk(gclk));
	jdff dff_A_uKaxxzL60_0(.dout(w_dff_A_yQiRHdtT6_0),.din(w_dff_A_uKaxxzL60_0),.clk(gclk));
	jdff dff_A_yQiRHdtT6_0(.dout(w_dff_A_lRdahrlG0_0),.din(w_dff_A_yQiRHdtT6_0),.clk(gclk));
	jdff dff_A_lRdahrlG0_0(.dout(f24),.din(w_dff_A_lRdahrlG0_0),.clk(gclk));
	jdff dff_A_0nEZ1YGf2_2(.dout(w_dff_A_XpUQpVdN7_0),.din(w_dff_A_0nEZ1YGf2_2),.clk(gclk));
	jdff dff_A_XpUQpVdN7_0(.dout(w_dff_A_5thKmnai7_0),.din(w_dff_A_XpUQpVdN7_0),.clk(gclk));
	jdff dff_A_5thKmnai7_0(.dout(w_dff_A_n8SdQJkF4_0),.din(w_dff_A_5thKmnai7_0),.clk(gclk));
	jdff dff_A_n8SdQJkF4_0(.dout(w_dff_A_z2uBN0HD1_0),.din(w_dff_A_n8SdQJkF4_0),.clk(gclk));
	jdff dff_A_z2uBN0HD1_0(.dout(w_dff_A_uZ0XBi0R4_0),.din(w_dff_A_z2uBN0HD1_0),.clk(gclk));
	jdff dff_A_uZ0XBi0R4_0(.dout(w_dff_A_Piisp0vd7_0),.din(w_dff_A_uZ0XBi0R4_0),.clk(gclk));
	jdff dff_A_Piisp0vd7_0(.dout(w_dff_A_t59uKDX81_0),.din(w_dff_A_Piisp0vd7_0),.clk(gclk));
	jdff dff_A_t59uKDX81_0(.dout(w_dff_A_cvH13HmV0_0),.din(w_dff_A_t59uKDX81_0),.clk(gclk));
	jdff dff_A_cvH13HmV0_0(.dout(w_dff_A_G2JPCfLJ4_0),.din(w_dff_A_cvH13HmV0_0),.clk(gclk));
	jdff dff_A_G2JPCfLJ4_0(.dout(w_dff_A_LDlLZ7Ya8_0),.din(w_dff_A_G2JPCfLJ4_0),.clk(gclk));
	jdff dff_A_LDlLZ7Ya8_0(.dout(w_dff_A_CZNR46Kc9_0),.din(w_dff_A_LDlLZ7Ya8_0),.clk(gclk));
	jdff dff_A_CZNR46Kc9_0(.dout(w_dff_A_JycQkhvU5_0),.din(w_dff_A_CZNR46Kc9_0),.clk(gclk));
	jdff dff_A_JycQkhvU5_0(.dout(w_dff_A_ESgeG3L03_0),.din(w_dff_A_JycQkhvU5_0),.clk(gclk));
	jdff dff_A_ESgeG3L03_0(.dout(w_dff_A_lgBszO8L4_0),.din(w_dff_A_ESgeG3L03_0),.clk(gclk));
	jdff dff_A_lgBszO8L4_0(.dout(w_dff_A_qyI2Er4q2_0),.din(w_dff_A_lgBszO8L4_0),.clk(gclk));
	jdff dff_A_qyI2Er4q2_0(.dout(w_dff_A_HTx9f88E5_0),.din(w_dff_A_qyI2Er4q2_0),.clk(gclk));
	jdff dff_A_HTx9f88E5_0(.dout(w_dff_A_siduIdft4_0),.din(w_dff_A_HTx9f88E5_0),.clk(gclk));
	jdff dff_A_siduIdft4_0(.dout(w_dff_A_LcJTspSp3_0),.din(w_dff_A_siduIdft4_0),.clk(gclk));
	jdff dff_A_LcJTspSp3_0(.dout(w_dff_A_C3kAR2FE0_0),.din(w_dff_A_LcJTspSp3_0),.clk(gclk));
	jdff dff_A_C3kAR2FE0_0(.dout(w_dff_A_Zz4CQQak3_0),.din(w_dff_A_C3kAR2FE0_0),.clk(gclk));
	jdff dff_A_Zz4CQQak3_0(.dout(w_dff_A_iuF9XDjk1_0),.din(w_dff_A_Zz4CQQak3_0),.clk(gclk));
	jdff dff_A_iuF9XDjk1_0(.dout(w_dff_A_AruhJiPA3_0),.din(w_dff_A_iuF9XDjk1_0),.clk(gclk));
	jdff dff_A_AruhJiPA3_0(.dout(w_dff_A_9sxbnDaN2_0),.din(w_dff_A_AruhJiPA3_0),.clk(gclk));
	jdff dff_A_9sxbnDaN2_0(.dout(w_dff_A_OyjrpZtk1_0),.din(w_dff_A_9sxbnDaN2_0),.clk(gclk));
	jdff dff_A_OyjrpZtk1_0(.dout(w_dff_A_QbxKWqba6_0),.din(w_dff_A_OyjrpZtk1_0),.clk(gclk));
	jdff dff_A_QbxKWqba6_0(.dout(w_dff_A_Q9vYBh663_0),.din(w_dff_A_QbxKWqba6_0),.clk(gclk));
	jdff dff_A_Q9vYBh663_0(.dout(w_dff_A_2Hs9V9YX4_0),.din(w_dff_A_Q9vYBh663_0),.clk(gclk));
	jdff dff_A_2Hs9V9YX4_0(.dout(w_dff_A_K1c8lOqV3_0),.din(w_dff_A_2Hs9V9YX4_0),.clk(gclk));
	jdff dff_A_K1c8lOqV3_0(.dout(w_dff_A_XQrGES744_0),.din(w_dff_A_K1c8lOqV3_0),.clk(gclk));
	jdff dff_A_XQrGES744_0(.dout(w_dff_A_mOFz25wK9_0),.din(w_dff_A_XQrGES744_0),.clk(gclk));
	jdff dff_A_mOFz25wK9_0(.dout(w_dff_A_LiVm21O92_0),.din(w_dff_A_mOFz25wK9_0),.clk(gclk));
	jdff dff_A_LiVm21O92_0(.dout(w_dff_A_E6f6xOtF7_0),.din(w_dff_A_LiVm21O92_0),.clk(gclk));
	jdff dff_A_E6f6xOtF7_0(.dout(w_dff_A_tS6CCnjV3_0),.din(w_dff_A_E6f6xOtF7_0),.clk(gclk));
	jdff dff_A_tS6CCnjV3_0(.dout(w_dff_A_XNF6ZSNS0_0),.din(w_dff_A_tS6CCnjV3_0),.clk(gclk));
	jdff dff_A_XNF6ZSNS0_0(.dout(w_dff_A_fiiYCJKr0_0),.din(w_dff_A_XNF6ZSNS0_0),.clk(gclk));
	jdff dff_A_fiiYCJKr0_0(.dout(w_dff_A_9eUdAo6S2_0),.din(w_dff_A_fiiYCJKr0_0),.clk(gclk));
	jdff dff_A_9eUdAo6S2_0(.dout(w_dff_A_0JQKAZh02_0),.din(w_dff_A_9eUdAo6S2_0),.clk(gclk));
	jdff dff_A_0JQKAZh02_0(.dout(w_dff_A_8ToBNj5J8_0),.din(w_dff_A_0JQKAZh02_0),.clk(gclk));
	jdff dff_A_8ToBNj5J8_0(.dout(w_dff_A_BVLiAXXL2_0),.din(w_dff_A_8ToBNj5J8_0),.clk(gclk));
	jdff dff_A_BVLiAXXL2_0(.dout(w_dff_A_CYUuieAQ3_0),.din(w_dff_A_BVLiAXXL2_0),.clk(gclk));
	jdff dff_A_CYUuieAQ3_0(.dout(w_dff_A_TqA6t0059_0),.din(w_dff_A_CYUuieAQ3_0),.clk(gclk));
	jdff dff_A_TqA6t0059_0(.dout(w_dff_A_sQrLNdjJ9_0),.din(w_dff_A_TqA6t0059_0),.clk(gclk));
	jdff dff_A_sQrLNdjJ9_0(.dout(w_dff_A_ZaJ6jopY8_0),.din(w_dff_A_sQrLNdjJ9_0),.clk(gclk));
	jdff dff_A_ZaJ6jopY8_0(.dout(w_dff_A_VuPzxNaY5_0),.din(w_dff_A_ZaJ6jopY8_0),.clk(gclk));
	jdff dff_A_VuPzxNaY5_0(.dout(w_dff_A_ciMS16dp8_0),.din(w_dff_A_VuPzxNaY5_0),.clk(gclk));
	jdff dff_A_ciMS16dp8_0(.dout(w_dff_A_Az1NZDsQ0_0),.din(w_dff_A_ciMS16dp8_0),.clk(gclk));
	jdff dff_A_Az1NZDsQ0_0(.dout(w_dff_A_SNYxVHDd6_0),.din(w_dff_A_Az1NZDsQ0_0),.clk(gclk));
	jdff dff_A_SNYxVHDd6_0(.dout(w_dff_A_fOppy9ci6_0),.din(w_dff_A_SNYxVHDd6_0),.clk(gclk));
	jdff dff_A_fOppy9ci6_0(.dout(w_dff_A_PM4uTAe31_0),.din(w_dff_A_fOppy9ci6_0),.clk(gclk));
	jdff dff_A_PM4uTAe31_0(.dout(w_dff_A_KAdNvwF04_0),.din(w_dff_A_PM4uTAe31_0),.clk(gclk));
	jdff dff_A_KAdNvwF04_0(.dout(w_dff_A_pYFBSyyQ3_0),.din(w_dff_A_KAdNvwF04_0),.clk(gclk));
	jdff dff_A_pYFBSyyQ3_0(.dout(w_dff_A_gE1KLIn52_0),.din(w_dff_A_pYFBSyyQ3_0),.clk(gclk));
	jdff dff_A_gE1KLIn52_0(.dout(w_dff_A_j15LUhPb0_0),.din(w_dff_A_gE1KLIn52_0),.clk(gclk));
	jdff dff_A_j15LUhPb0_0(.dout(w_dff_A_IzFGJGlB4_0),.din(w_dff_A_j15LUhPb0_0),.clk(gclk));
	jdff dff_A_IzFGJGlB4_0(.dout(w_dff_A_9ih4B6lu8_0),.din(w_dff_A_IzFGJGlB4_0),.clk(gclk));
	jdff dff_A_9ih4B6lu8_0(.dout(w_dff_A_4pfPp2v81_0),.din(w_dff_A_9ih4B6lu8_0),.clk(gclk));
	jdff dff_A_4pfPp2v81_0(.dout(w_dff_A_4UTkAK6z4_0),.din(w_dff_A_4pfPp2v81_0),.clk(gclk));
	jdff dff_A_4UTkAK6z4_0(.dout(w_dff_A_ac8uZy296_0),.din(w_dff_A_4UTkAK6z4_0),.clk(gclk));
	jdff dff_A_ac8uZy296_0(.dout(w_dff_A_lxtRVMAD0_0),.din(w_dff_A_ac8uZy296_0),.clk(gclk));
	jdff dff_A_lxtRVMAD0_0(.dout(w_dff_A_Sf8lL5I23_0),.din(w_dff_A_lxtRVMAD0_0),.clk(gclk));
	jdff dff_A_Sf8lL5I23_0(.dout(w_dff_A_kwuv0SpU5_0),.din(w_dff_A_Sf8lL5I23_0),.clk(gclk));
	jdff dff_A_kwuv0SpU5_0(.dout(w_dff_A_joiyyHKD8_0),.din(w_dff_A_kwuv0SpU5_0),.clk(gclk));
	jdff dff_A_joiyyHKD8_0(.dout(w_dff_A_2KleqGgU8_0),.din(w_dff_A_joiyyHKD8_0),.clk(gclk));
	jdff dff_A_2KleqGgU8_0(.dout(w_dff_A_poGmEZQK4_0),.din(w_dff_A_2KleqGgU8_0),.clk(gclk));
	jdff dff_A_poGmEZQK4_0(.dout(w_dff_A_6QcNXvES6_0),.din(w_dff_A_poGmEZQK4_0),.clk(gclk));
	jdff dff_A_6QcNXvES6_0(.dout(w_dff_A_IxqDbUPP0_0),.din(w_dff_A_6QcNXvES6_0),.clk(gclk));
	jdff dff_A_IxqDbUPP0_0(.dout(w_dff_A_ElvEYsr06_0),.din(w_dff_A_IxqDbUPP0_0),.clk(gclk));
	jdff dff_A_ElvEYsr06_0(.dout(w_dff_A_b953PdWO9_0),.din(w_dff_A_ElvEYsr06_0),.clk(gclk));
	jdff dff_A_b953PdWO9_0(.dout(w_dff_A_AfY7WRZe5_0),.din(w_dff_A_b953PdWO9_0),.clk(gclk));
	jdff dff_A_AfY7WRZe5_0(.dout(w_dff_A_4dCduNFl5_0),.din(w_dff_A_AfY7WRZe5_0),.clk(gclk));
	jdff dff_A_4dCduNFl5_0(.dout(w_dff_A_r11WoBd07_0),.din(w_dff_A_4dCduNFl5_0),.clk(gclk));
	jdff dff_A_r11WoBd07_0(.dout(w_dff_A_IcebyBVR6_0),.din(w_dff_A_r11WoBd07_0),.clk(gclk));
	jdff dff_A_IcebyBVR6_0(.dout(w_dff_A_cw0ijJ1f5_0),.din(w_dff_A_IcebyBVR6_0),.clk(gclk));
	jdff dff_A_cw0ijJ1f5_0(.dout(w_dff_A_Wkt1B6bc8_0),.din(w_dff_A_cw0ijJ1f5_0),.clk(gclk));
	jdff dff_A_Wkt1B6bc8_0(.dout(w_dff_A_l7zRAedK6_0),.din(w_dff_A_Wkt1B6bc8_0),.clk(gclk));
	jdff dff_A_l7zRAedK6_0(.dout(w_dff_A_cRCBYTGX2_0),.din(w_dff_A_l7zRAedK6_0),.clk(gclk));
	jdff dff_A_cRCBYTGX2_0(.dout(w_dff_A_6fQmR3Kw0_0),.din(w_dff_A_cRCBYTGX2_0),.clk(gclk));
	jdff dff_A_6fQmR3Kw0_0(.dout(w_dff_A_pTfgEiJ99_0),.din(w_dff_A_6fQmR3Kw0_0),.clk(gclk));
	jdff dff_A_pTfgEiJ99_0(.dout(w_dff_A_JkVtL0DQ6_0),.din(w_dff_A_pTfgEiJ99_0),.clk(gclk));
	jdff dff_A_JkVtL0DQ6_0(.dout(w_dff_A_uJ4KZjgh4_0),.din(w_dff_A_JkVtL0DQ6_0),.clk(gclk));
	jdff dff_A_uJ4KZjgh4_0(.dout(w_dff_A_QrqrotYQ9_0),.din(w_dff_A_uJ4KZjgh4_0),.clk(gclk));
	jdff dff_A_QrqrotYQ9_0(.dout(w_dff_A_i14hUG3K5_0),.din(w_dff_A_QrqrotYQ9_0),.clk(gclk));
	jdff dff_A_i14hUG3K5_0(.dout(w_dff_A_TEveETai2_0),.din(w_dff_A_i14hUG3K5_0),.clk(gclk));
	jdff dff_A_TEveETai2_0(.dout(w_dff_A_k1wJ2nx67_0),.din(w_dff_A_TEveETai2_0),.clk(gclk));
	jdff dff_A_k1wJ2nx67_0(.dout(w_dff_A_0HSHNax31_0),.din(w_dff_A_k1wJ2nx67_0),.clk(gclk));
	jdff dff_A_0HSHNax31_0(.dout(w_dff_A_dJYTji9n6_0),.din(w_dff_A_0HSHNax31_0),.clk(gclk));
	jdff dff_A_dJYTji9n6_0(.dout(w_dff_A_ZCqFWlPC1_0),.din(w_dff_A_dJYTji9n6_0),.clk(gclk));
	jdff dff_A_ZCqFWlPC1_0(.dout(w_dff_A_g7sfD5oQ3_0),.din(w_dff_A_ZCqFWlPC1_0),.clk(gclk));
	jdff dff_A_g7sfD5oQ3_0(.dout(w_dff_A_N2RzlP2m1_0),.din(w_dff_A_g7sfD5oQ3_0),.clk(gclk));
	jdff dff_A_N2RzlP2m1_0(.dout(w_dff_A_aEDIY8A09_0),.din(w_dff_A_N2RzlP2m1_0),.clk(gclk));
	jdff dff_A_aEDIY8A09_0(.dout(w_dff_A_symwYzaY6_0),.din(w_dff_A_aEDIY8A09_0),.clk(gclk));
	jdff dff_A_symwYzaY6_0(.dout(w_dff_A_Nlm5jXQU7_0),.din(w_dff_A_symwYzaY6_0),.clk(gclk));
	jdff dff_A_Nlm5jXQU7_0(.dout(w_dff_A_bRV5paq16_0),.din(w_dff_A_Nlm5jXQU7_0),.clk(gclk));
	jdff dff_A_bRV5paq16_0(.dout(w_dff_A_GvoORiBG0_0),.din(w_dff_A_bRV5paq16_0),.clk(gclk));
	jdff dff_A_GvoORiBG0_0(.dout(w_dff_A_LZe8Cn5W9_0),.din(w_dff_A_GvoORiBG0_0),.clk(gclk));
	jdff dff_A_LZe8Cn5W9_0(.dout(w_dff_A_s4pctpVC2_0),.din(w_dff_A_LZe8Cn5W9_0),.clk(gclk));
	jdff dff_A_s4pctpVC2_0(.dout(w_dff_A_yyPkTCU93_0),.din(w_dff_A_s4pctpVC2_0),.clk(gclk));
	jdff dff_A_yyPkTCU93_0(.dout(w_dff_A_SesGA1bx1_0),.din(w_dff_A_yyPkTCU93_0),.clk(gclk));
	jdff dff_A_SesGA1bx1_0(.dout(w_dff_A_uEVqlit24_0),.din(w_dff_A_SesGA1bx1_0),.clk(gclk));
	jdff dff_A_uEVqlit24_0(.dout(w_dff_A_W90yQBs47_0),.din(w_dff_A_uEVqlit24_0),.clk(gclk));
	jdff dff_A_W90yQBs47_0(.dout(w_dff_A_x3X9er1E3_0),.din(w_dff_A_W90yQBs47_0),.clk(gclk));
	jdff dff_A_x3X9er1E3_0(.dout(f25),.din(w_dff_A_x3X9er1E3_0),.clk(gclk));
	jdff dff_A_M4eemYt31_2(.dout(w_dff_A_AwhbLbvS6_0),.din(w_dff_A_M4eemYt31_2),.clk(gclk));
	jdff dff_A_AwhbLbvS6_0(.dout(w_dff_A_rSr6SRMx2_0),.din(w_dff_A_AwhbLbvS6_0),.clk(gclk));
	jdff dff_A_rSr6SRMx2_0(.dout(w_dff_A_SmA2fzwJ5_0),.din(w_dff_A_rSr6SRMx2_0),.clk(gclk));
	jdff dff_A_SmA2fzwJ5_0(.dout(w_dff_A_5rHiVLHD0_0),.din(w_dff_A_SmA2fzwJ5_0),.clk(gclk));
	jdff dff_A_5rHiVLHD0_0(.dout(w_dff_A_bmCnJbg39_0),.din(w_dff_A_5rHiVLHD0_0),.clk(gclk));
	jdff dff_A_bmCnJbg39_0(.dout(w_dff_A_mPkeNnAl7_0),.din(w_dff_A_bmCnJbg39_0),.clk(gclk));
	jdff dff_A_mPkeNnAl7_0(.dout(w_dff_A_ow920u5m8_0),.din(w_dff_A_mPkeNnAl7_0),.clk(gclk));
	jdff dff_A_ow920u5m8_0(.dout(w_dff_A_EIR3NQ3l0_0),.din(w_dff_A_ow920u5m8_0),.clk(gclk));
	jdff dff_A_EIR3NQ3l0_0(.dout(w_dff_A_47tVZ46P3_0),.din(w_dff_A_EIR3NQ3l0_0),.clk(gclk));
	jdff dff_A_47tVZ46P3_0(.dout(w_dff_A_8DzQKIKq7_0),.din(w_dff_A_47tVZ46P3_0),.clk(gclk));
	jdff dff_A_8DzQKIKq7_0(.dout(w_dff_A_IJqun7Xu4_0),.din(w_dff_A_8DzQKIKq7_0),.clk(gclk));
	jdff dff_A_IJqun7Xu4_0(.dout(w_dff_A_0bdPYpd87_0),.din(w_dff_A_IJqun7Xu4_0),.clk(gclk));
	jdff dff_A_0bdPYpd87_0(.dout(w_dff_A_4iyrtd2z5_0),.din(w_dff_A_0bdPYpd87_0),.clk(gclk));
	jdff dff_A_4iyrtd2z5_0(.dout(w_dff_A_aX7UIuPX4_0),.din(w_dff_A_4iyrtd2z5_0),.clk(gclk));
	jdff dff_A_aX7UIuPX4_0(.dout(w_dff_A_1gQezk1d7_0),.din(w_dff_A_aX7UIuPX4_0),.clk(gclk));
	jdff dff_A_1gQezk1d7_0(.dout(w_dff_A_CbxhIpxn5_0),.din(w_dff_A_1gQezk1d7_0),.clk(gclk));
	jdff dff_A_CbxhIpxn5_0(.dout(w_dff_A_wfJAe4av2_0),.din(w_dff_A_CbxhIpxn5_0),.clk(gclk));
	jdff dff_A_wfJAe4av2_0(.dout(w_dff_A_UMDqXr348_0),.din(w_dff_A_wfJAe4av2_0),.clk(gclk));
	jdff dff_A_UMDqXr348_0(.dout(w_dff_A_pr0ZCi2E3_0),.din(w_dff_A_UMDqXr348_0),.clk(gclk));
	jdff dff_A_pr0ZCi2E3_0(.dout(w_dff_A_W0E2eudA5_0),.din(w_dff_A_pr0ZCi2E3_0),.clk(gclk));
	jdff dff_A_W0E2eudA5_0(.dout(w_dff_A_jvXVb8bu4_0),.din(w_dff_A_W0E2eudA5_0),.clk(gclk));
	jdff dff_A_jvXVb8bu4_0(.dout(w_dff_A_A4t18bvA2_0),.din(w_dff_A_jvXVb8bu4_0),.clk(gclk));
	jdff dff_A_A4t18bvA2_0(.dout(w_dff_A_NPMz15Gh0_0),.din(w_dff_A_A4t18bvA2_0),.clk(gclk));
	jdff dff_A_NPMz15Gh0_0(.dout(w_dff_A_j3DzRLm82_0),.din(w_dff_A_NPMz15Gh0_0),.clk(gclk));
	jdff dff_A_j3DzRLm82_0(.dout(w_dff_A_CRZMfwm49_0),.din(w_dff_A_j3DzRLm82_0),.clk(gclk));
	jdff dff_A_CRZMfwm49_0(.dout(w_dff_A_Jtu5BTpk1_0),.din(w_dff_A_CRZMfwm49_0),.clk(gclk));
	jdff dff_A_Jtu5BTpk1_0(.dout(w_dff_A_gBldQUzH8_0),.din(w_dff_A_Jtu5BTpk1_0),.clk(gclk));
	jdff dff_A_gBldQUzH8_0(.dout(w_dff_A_v7uE4mJ59_0),.din(w_dff_A_gBldQUzH8_0),.clk(gclk));
	jdff dff_A_v7uE4mJ59_0(.dout(w_dff_A_Ep5WBgiY6_0),.din(w_dff_A_v7uE4mJ59_0),.clk(gclk));
	jdff dff_A_Ep5WBgiY6_0(.dout(w_dff_A_IXnFGN1c5_0),.din(w_dff_A_Ep5WBgiY6_0),.clk(gclk));
	jdff dff_A_IXnFGN1c5_0(.dout(w_dff_A_gkPPHvL01_0),.din(w_dff_A_IXnFGN1c5_0),.clk(gclk));
	jdff dff_A_gkPPHvL01_0(.dout(w_dff_A_5IEqqgjo9_0),.din(w_dff_A_gkPPHvL01_0),.clk(gclk));
	jdff dff_A_5IEqqgjo9_0(.dout(w_dff_A_qpDgwJBG4_0),.din(w_dff_A_5IEqqgjo9_0),.clk(gclk));
	jdff dff_A_qpDgwJBG4_0(.dout(w_dff_A_3Gxms4ll2_0),.din(w_dff_A_qpDgwJBG4_0),.clk(gclk));
	jdff dff_A_3Gxms4ll2_0(.dout(w_dff_A_jEq3sh0o6_0),.din(w_dff_A_3Gxms4ll2_0),.clk(gclk));
	jdff dff_A_jEq3sh0o6_0(.dout(w_dff_A_6DiZT4nb9_0),.din(w_dff_A_jEq3sh0o6_0),.clk(gclk));
	jdff dff_A_6DiZT4nb9_0(.dout(w_dff_A_lnjxgXyp8_0),.din(w_dff_A_6DiZT4nb9_0),.clk(gclk));
	jdff dff_A_lnjxgXyp8_0(.dout(w_dff_A_uIFJt6je6_0),.din(w_dff_A_lnjxgXyp8_0),.clk(gclk));
	jdff dff_A_uIFJt6je6_0(.dout(w_dff_A_72ADBfXj2_0),.din(w_dff_A_uIFJt6je6_0),.clk(gclk));
	jdff dff_A_72ADBfXj2_0(.dout(w_dff_A_FsRRNwpR8_0),.din(w_dff_A_72ADBfXj2_0),.clk(gclk));
	jdff dff_A_FsRRNwpR8_0(.dout(w_dff_A_lvE2aJxj2_0),.din(w_dff_A_FsRRNwpR8_0),.clk(gclk));
	jdff dff_A_lvE2aJxj2_0(.dout(w_dff_A_xxvSkDpq0_0),.din(w_dff_A_lvE2aJxj2_0),.clk(gclk));
	jdff dff_A_xxvSkDpq0_0(.dout(w_dff_A_BQ0CF9jx4_0),.din(w_dff_A_xxvSkDpq0_0),.clk(gclk));
	jdff dff_A_BQ0CF9jx4_0(.dout(w_dff_A_VO8oeS5O6_0),.din(w_dff_A_BQ0CF9jx4_0),.clk(gclk));
	jdff dff_A_VO8oeS5O6_0(.dout(w_dff_A_qYblETKR2_0),.din(w_dff_A_VO8oeS5O6_0),.clk(gclk));
	jdff dff_A_qYblETKR2_0(.dout(w_dff_A_h5e7WUCW0_0),.din(w_dff_A_qYblETKR2_0),.clk(gclk));
	jdff dff_A_h5e7WUCW0_0(.dout(w_dff_A_0YyHPbH77_0),.din(w_dff_A_h5e7WUCW0_0),.clk(gclk));
	jdff dff_A_0YyHPbH77_0(.dout(w_dff_A_do74JSrz6_0),.din(w_dff_A_0YyHPbH77_0),.clk(gclk));
	jdff dff_A_do74JSrz6_0(.dout(w_dff_A_H4O3llyJ9_0),.din(w_dff_A_do74JSrz6_0),.clk(gclk));
	jdff dff_A_H4O3llyJ9_0(.dout(w_dff_A_hjpWyEbc5_0),.din(w_dff_A_H4O3llyJ9_0),.clk(gclk));
	jdff dff_A_hjpWyEbc5_0(.dout(w_dff_A_qoroFDrB1_0),.din(w_dff_A_hjpWyEbc5_0),.clk(gclk));
	jdff dff_A_qoroFDrB1_0(.dout(w_dff_A_teEdXXph2_0),.din(w_dff_A_qoroFDrB1_0),.clk(gclk));
	jdff dff_A_teEdXXph2_0(.dout(w_dff_A_adhHJpla8_0),.din(w_dff_A_teEdXXph2_0),.clk(gclk));
	jdff dff_A_adhHJpla8_0(.dout(w_dff_A_68o9WCJt7_0),.din(w_dff_A_adhHJpla8_0),.clk(gclk));
	jdff dff_A_68o9WCJt7_0(.dout(w_dff_A_5TlTkyEc5_0),.din(w_dff_A_68o9WCJt7_0),.clk(gclk));
	jdff dff_A_5TlTkyEc5_0(.dout(w_dff_A_VMd8OwCf6_0),.din(w_dff_A_5TlTkyEc5_0),.clk(gclk));
	jdff dff_A_VMd8OwCf6_0(.dout(w_dff_A_cDe528kn5_0),.din(w_dff_A_VMd8OwCf6_0),.clk(gclk));
	jdff dff_A_cDe528kn5_0(.dout(w_dff_A_OA3KMFzw5_0),.din(w_dff_A_cDe528kn5_0),.clk(gclk));
	jdff dff_A_OA3KMFzw5_0(.dout(w_dff_A_ORsblvhe9_0),.din(w_dff_A_OA3KMFzw5_0),.clk(gclk));
	jdff dff_A_ORsblvhe9_0(.dout(w_dff_A_QlqjVhUC7_0),.din(w_dff_A_ORsblvhe9_0),.clk(gclk));
	jdff dff_A_QlqjVhUC7_0(.dout(w_dff_A_OcZ2RIcp8_0),.din(w_dff_A_QlqjVhUC7_0),.clk(gclk));
	jdff dff_A_OcZ2RIcp8_0(.dout(w_dff_A_YWlqxvnI8_0),.din(w_dff_A_OcZ2RIcp8_0),.clk(gclk));
	jdff dff_A_YWlqxvnI8_0(.dout(w_dff_A_tSju8ERv6_0),.din(w_dff_A_YWlqxvnI8_0),.clk(gclk));
	jdff dff_A_tSju8ERv6_0(.dout(w_dff_A_l3p1HFJs9_0),.din(w_dff_A_tSju8ERv6_0),.clk(gclk));
	jdff dff_A_l3p1HFJs9_0(.dout(w_dff_A_LCy2irS62_0),.din(w_dff_A_l3p1HFJs9_0),.clk(gclk));
	jdff dff_A_LCy2irS62_0(.dout(w_dff_A_S2HXu8WE8_0),.din(w_dff_A_LCy2irS62_0),.clk(gclk));
	jdff dff_A_S2HXu8WE8_0(.dout(w_dff_A_lGd6oMyr3_0),.din(w_dff_A_S2HXu8WE8_0),.clk(gclk));
	jdff dff_A_lGd6oMyr3_0(.dout(w_dff_A_nZMV21yo1_0),.din(w_dff_A_lGd6oMyr3_0),.clk(gclk));
	jdff dff_A_nZMV21yo1_0(.dout(w_dff_A_2dDEbAuI8_0),.din(w_dff_A_nZMV21yo1_0),.clk(gclk));
	jdff dff_A_2dDEbAuI8_0(.dout(w_dff_A_mvSkrnOo8_0),.din(w_dff_A_2dDEbAuI8_0),.clk(gclk));
	jdff dff_A_mvSkrnOo8_0(.dout(w_dff_A_JDqeIWOB3_0),.din(w_dff_A_mvSkrnOo8_0),.clk(gclk));
	jdff dff_A_JDqeIWOB3_0(.dout(w_dff_A_zLa4xw4d8_0),.din(w_dff_A_JDqeIWOB3_0),.clk(gclk));
	jdff dff_A_zLa4xw4d8_0(.dout(w_dff_A_NHTmnWzZ6_0),.din(w_dff_A_zLa4xw4d8_0),.clk(gclk));
	jdff dff_A_NHTmnWzZ6_0(.dout(w_dff_A_kBywAWeH1_0),.din(w_dff_A_NHTmnWzZ6_0),.clk(gclk));
	jdff dff_A_kBywAWeH1_0(.dout(w_dff_A_s41c1RUy2_0),.din(w_dff_A_kBywAWeH1_0),.clk(gclk));
	jdff dff_A_s41c1RUy2_0(.dout(w_dff_A_Pow3qPc02_0),.din(w_dff_A_s41c1RUy2_0),.clk(gclk));
	jdff dff_A_Pow3qPc02_0(.dout(w_dff_A_YZtryBzI5_0),.din(w_dff_A_Pow3qPc02_0),.clk(gclk));
	jdff dff_A_YZtryBzI5_0(.dout(w_dff_A_ThqVqPIM1_0),.din(w_dff_A_YZtryBzI5_0),.clk(gclk));
	jdff dff_A_ThqVqPIM1_0(.dout(w_dff_A_N18mvCOA7_0),.din(w_dff_A_ThqVqPIM1_0),.clk(gclk));
	jdff dff_A_N18mvCOA7_0(.dout(w_dff_A_dCrDcmGc0_0),.din(w_dff_A_N18mvCOA7_0),.clk(gclk));
	jdff dff_A_dCrDcmGc0_0(.dout(w_dff_A_NFr1gWhT7_0),.din(w_dff_A_dCrDcmGc0_0),.clk(gclk));
	jdff dff_A_NFr1gWhT7_0(.dout(w_dff_A_jSzvHIwD2_0),.din(w_dff_A_NFr1gWhT7_0),.clk(gclk));
	jdff dff_A_jSzvHIwD2_0(.dout(w_dff_A_bZEafMQb4_0),.din(w_dff_A_jSzvHIwD2_0),.clk(gclk));
	jdff dff_A_bZEafMQb4_0(.dout(w_dff_A_CrFqYhE37_0),.din(w_dff_A_bZEafMQb4_0),.clk(gclk));
	jdff dff_A_CrFqYhE37_0(.dout(w_dff_A_uz0G5zVt6_0),.din(w_dff_A_CrFqYhE37_0),.clk(gclk));
	jdff dff_A_uz0G5zVt6_0(.dout(w_dff_A_5YEyLRgp1_0),.din(w_dff_A_uz0G5zVt6_0),.clk(gclk));
	jdff dff_A_5YEyLRgp1_0(.dout(w_dff_A_une5EDtn3_0),.din(w_dff_A_5YEyLRgp1_0),.clk(gclk));
	jdff dff_A_une5EDtn3_0(.dout(w_dff_A_HHmjhqcT3_0),.din(w_dff_A_une5EDtn3_0),.clk(gclk));
	jdff dff_A_HHmjhqcT3_0(.dout(w_dff_A_ABjHjKIJ1_0),.din(w_dff_A_HHmjhqcT3_0),.clk(gclk));
	jdff dff_A_ABjHjKIJ1_0(.dout(w_dff_A_L3Vo3gBg8_0),.din(w_dff_A_ABjHjKIJ1_0),.clk(gclk));
	jdff dff_A_L3Vo3gBg8_0(.dout(w_dff_A_AWlYYlg03_0),.din(w_dff_A_L3Vo3gBg8_0),.clk(gclk));
	jdff dff_A_AWlYYlg03_0(.dout(w_dff_A_JPX9N0WJ6_0),.din(w_dff_A_AWlYYlg03_0),.clk(gclk));
	jdff dff_A_JPX9N0WJ6_0(.dout(w_dff_A_19a4yM0v1_0),.din(w_dff_A_JPX9N0WJ6_0),.clk(gclk));
	jdff dff_A_19a4yM0v1_0(.dout(w_dff_A_eVPz5MYC9_0),.din(w_dff_A_19a4yM0v1_0),.clk(gclk));
	jdff dff_A_eVPz5MYC9_0(.dout(w_dff_A_GGaeYQ9t8_0),.din(w_dff_A_eVPz5MYC9_0),.clk(gclk));
	jdff dff_A_GGaeYQ9t8_0(.dout(w_dff_A_JgsCMeoa0_0),.din(w_dff_A_GGaeYQ9t8_0),.clk(gclk));
	jdff dff_A_JgsCMeoa0_0(.dout(w_dff_A_kAXY9dL53_0),.din(w_dff_A_JgsCMeoa0_0),.clk(gclk));
	jdff dff_A_kAXY9dL53_0(.dout(w_dff_A_2Ly2Dkto3_0),.din(w_dff_A_kAXY9dL53_0),.clk(gclk));
	jdff dff_A_2Ly2Dkto3_0(.dout(w_dff_A_flgrYN4N1_0),.din(w_dff_A_2Ly2Dkto3_0),.clk(gclk));
	jdff dff_A_flgrYN4N1_0(.dout(w_dff_A_DGVT5jvk5_0),.din(w_dff_A_flgrYN4N1_0),.clk(gclk));
	jdff dff_A_DGVT5jvk5_0(.dout(f26),.din(w_dff_A_DGVT5jvk5_0),.clk(gclk));
	jdff dff_A_JIss0YJB5_2(.dout(w_dff_A_dFCI4bb25_0),.din(w_dff_A_JIss0YJB5_2),.clk(gclk));
	jdff dff_A_dFCI4bb25_0(.dout(w_dff_A_GFVnMEX32_0),.din(w_dff_A_dFCI4bb25_0),.clk(gclk));
	jdff dff_A_GFVnMEX32_0(.dout(w_dff_A_PdhYMYTa6_0),.din(w_dff_A_GFVnMEX32_0),.clk(gclk));
	jdff dff_A_PdhYMYTa6_0(.dout(w_dff_A_uwY7OENu0_0),.din(w_dff_A_PdhYMYTa6_0),.clk(gclk));
	jdff dff_A_uwY7OENu0_0(.dout(w_dff_A_DwBmud3r9_0),.din(w_dff_A_uwY7OENu0_0),.clk(gclk));
	jdff dff_A_DwBmud3r9_0(.dout(w_dff_A_QcemS1tT2_0),.din(w_dff_A_DwBmud3r9_0),.clk(gclk));
	jdff dff_A_QcemS1tT2_0(.dout(w_dff_A_dF2stYhj8_0),.din(w_dff_A_QcemS1tT2_0),.clk(gclk));
	jdff dff_A_dF2stYhj8_0(.dout(w_dff_A_QEWyKXxR0_0),.din(w_dff_A_dF2stYhj8_0),.clk(gclk));
	jdff dff_A_QEWyKXxR0_0(.dout(w_dff_A_BP5s2Fs15_0),.din(w_dff_A_QEWyKXxR0_0),.clk(gclk));
	jdff dff_A_BP5s2Fs15_0(.dout(w_dff_A_sCdy9pmJ7_0),.din(w_dff_A_BP5s2Fs15_0),.clk(gclk));
	jdff dff_A_sCdy9pmJ7_0(.dout(w_dff_A_BAY9jtZM7_0),.din(w_dff_A_sCdy9pmJ7_0),.clk(gclk));
	jdff dff_A_BAY9jtZM7_0(.dout(w_dff_A_3DrsgkwA4_0),.din(w_dff_A_BAY9jtZM7_0),.clk(gclk));
	jdff dff_A_3DrsgkwA4_0(.dout(w_dff_A_O7FILHmv1_0),.din(w_dff_A_3DrsgkwA4_0),.clk(gclk));
	jdff dff_A_O7FILHmv1_0(.dout(w_dff_A_dCCpwe6g4_0),.din(w_dff_A_O7FILHmv1_0),.clk(gclk));
	jdff dff_A_dCCpwe6g4_0(.dout(w_dff_A_ccFSYTPt6_0),.din(w_dff_A_dCCpwe6g4_0),.clk(gclk));
	jdff dff_A_ccFSYTPt6_0(.dout(w_dff_A_z7sxxBzn0_0),.din(w_dff_A_ccFSYTPt6_0),.clk(gclk));
	jdff dff_A_z7sxxBzn0_0(.dout(w_dff_A_WiuD2U8K2_0),.din(w_dff_A_z7sxxBzn0_0),.clk(gclk));
	jdff dff_A_WiuD2U8K2_0(.dout(w_dff_A_NDPKldIP0_0),.din(w_dff_A_WiuD2U8K2_0),.clk(gclk));
	jdff dff_A_NDPKldIP0_0(.dout(w_dff_A_uv4kS5KF2_0),.din(w_dff_A_NDPKldIP0_0),.clk(gclk));
	jdff dff_A_uv4kS5KF2_0(.dout(w_dff_A_EInzX4nG2_0),.din(w_dff_A_uv4kS5KF2_0),.clk(gclk));
	jdff dff_A_EInzX4nG2_0(.dout(w_dff_A_SXRDNqca6_0),.din(w_dff_A_EInzX4nG2_0),.clk(gclk));
	jdff dff_A_SXRDNqca6_0(.dout(w_dff_A_UeQg360x7_0),.din(w_dff_A_SXRDNqca6_0),.clk(gclk));
	jdff dff_A_UeQg360x7_0(.dout(w_dff_A_nmm01ZeL2_0),.din(w_dff_A_UeQg360x7_0),.clk(gclk));
	jdff dff_A_nmm01ZeL2_0(.dout(w_dff_A_T7UI2LqQ6_0),.din(w_dff_A_nmm01ZeL2_0),.clk(gclk));
	jdff dff_A_T7UI2LqQ6_0(.dout(w_dff_A_lFapPDyx4_0),.din(w_dff_A_T7UI2LqQ6_0),.clk(gclk));
	jdff dff_A_lFapPDyx4_0(.dout(w_dff_A_UKtNuHeG7_0),.din(w_dff_A_lFapPDyx4_0),.clk(gclk));
	jdff dff_A_UKtNuHeG7_0(.dout(w_dff_A_mz5OpgzS5_0),.din(w_dff_A_UKtNuHeG7_0),.clk(gclk));
	jdff dff_A_mz5OpgzS5_0(.dout(w_dff_A_djjwCMzg8_0),.din(w_dff_A_mz5OpgzS5_0),.clk(gclk));
	jdff dff_A_djjwCMzg8_0(.dout(w_dff_A_0jpo4vPB3_0),.din(w_dff_A_djjwCMzg8_0),.clk(gclk));
	jdff dff_A_0jpo4vPB3_0(.dout(w_dff_A_V90F3OSd8_0),.din(w_dff_A_0jpo4vPB3_0),.clk(gclk));
	jdff dff_A_V90F3OSd8_0(.dout(w_dff_A_renxw8Dy1_0),.din(w_dff_A_V90F3OSd8_0),.clk(gclk));
	jdff dff_A_renxw8Dy1_0(.dout(w_dff_A_yJ4zkDVc7_0),.din(w_dff_A_renxw8Dy1_0),.clk(gclk));
	jdff dff_A_yJ4zkDVc7_0(.dout(w_dff_A_vaM0UJ282_0),.din(w_dff_A_yJ4zkDVc7_0),.clk(gclk));
	jdff dff_A_vaM0UJ282_0(.dout(w_dff_A_O8PSyLRJ1_0),.din(w_dff_A_vaM0UJ282_0),.clk(gclk));
	jdff dff_A_O8PSyLRJ1_0(.dout(w_dff_A_Y7eQ8eLF1_0),.din(w_dff_A_O8PSyLRJ1_0),.clk(gclk));
	jdff dff_A_Y7eQ8eLF1_0(.dout(w_dff_A_58NvqY4K1_0),.din(w_dff_A_Y7eQ8eLF1_0),.clk(gclk));
	jdff dff_A_58NvqY4K1_0(.dout(w_dff_A_fa3M0Vwx4_0),.din(w_dff_A_58NvqY4K1_0),.clk(gclk));
	jdff dff_A_fa3M0Vwx4_0(.dout(w_dff_A_L4fIWzaq4_0),.din(w_dff_A_fa3M0Vwx4_0),.clk(gclk));
	jdff dff_A_L4fIWzaq4_0(.dout(w_dff_A_4hDSqpYX9_0),.din(w_dff_A_L4fIWzaq4_0),.clk(gclk));
	jdff dff_A_4hDSqpYX9_0(.dout(w_dff_A_69heILq08_0),.din(w_dff_A_4hDSqpYX9_0),.clk(gclk));
	jdff dff_A_69heILq08_0(.dout(w_dff_A_lDrRWOtQ4_0),.din(w_dff_A_69heILq08_0),.clk(gclk));
	jdff dff_A_lDrRWOtQ4_0(.dout(w_dff_A_iUBY8FeP4_0),.din(w_dff_A_lDrRWOtQ4_0),.clk(gclk));
	jdff dff_A_iUBY8FeP4_0(.dout(w_dff_A_TIR4IRzl3_0),.din(w_dff_A_iUBY8FeP4_0),.clk(gclk));
	jdff dff_A_TIR4IRzl3_0(.dout(w_dff_A_JDijeVCl4_0),.din(w_dff_A_TIR4IRzl3_0),.clk(gclk));
	jdff dff_A_JDijeVCl4_0(.dout(w_dff_A_vKPhDFbO0_0),.din(w_dff_A_JDijeVCl4_0),.clk(gclk));
	jdff dff_A_vKPhDFbO0_0(.dout(w_dff_A_6ns2hWIN5_0),.din(w_dff_A_vKPhDFbO0_0),.clk(gclk));
	jdff dff_A_6ns2hWIN5_0(.dout(w_dff_A_Na6CQS4z7_0),.din(w_dff_A_6ns2hWIN5_0),.clk(gclk));
	jdff dff_A_Na6CQS4z7_0(.dout(w_dff_A_tXYMzNL66_0),.din(w_dff_A_Na6CQS4z7_0),.clk(gclk));
	jdff dff_A_tXYMzNL66_0(.dout(w_dff_A_E54WVSOc3_0),.din(w_dff_A_tXYMzNL66_0),.clk(gclk));
	jdff dff_A_E54WVSOc3_0(.dout(w_dff_A_BSKt0ocr1_0),.din(w_dff_A_E54WVSOc3_0),.clk(gclk));
	jdff dff_A_BSKt0ocr1_0(.dout(w_dff_A_dHs4lF3q7_0),.din(w_dff_A_BSKt0ocr1_0),.clk(gclk));
	jdff dff_A_dHs4lF3q7_0(.dout(w_dff_A_0fw8tlyi2_0),.din(w_dff_A_dHs4lF3q7_0),.clk(gclk));
	jdff dff_A_0fw8tlyi2_0(.dout(w_dff_A_Ilb9BIp96_0),.din(w_dff_A_0fw8tlyi2_0),.clk(gclk));
	jdff dff_A_Ilb9BIp96_0(.dout(w_dff_A_IAU5FW1b1_0),.din(w_dff_A_Ilb9BIp96_0),.clk(gclk));
	jdff dff_A_IAU5FW1b1_0(.dout(w_dff_A_idXBsFgP0_0),.din(w_dff_A_IAU5FW1b1_0),.clk(gclk));
	jdff dff_A_idXBsFgP0_0(.dout(w_dff_A_EcQN55hq3_0),.din(w_dff_A_idXBsFgP0_0),.clk(gclk));
	jdff dff_A_EcQN55hq3_0(.dout(w_dff_A_LHHL1ujd8_0),.din(w_dff_A_EcQN55hq3_0),.clk(gclk));
	jdff dff_A_LHHL1ujd8_0(.dout(w_dff_A_piItm0YG7_0),.din(w_dff_A_LHHL1ujd8_0),.clk(gclk));
	jdff dff_A_piItm0YG7_0(.dout(w_dff_A_uzv6tZZ44_0),.din(w_dff_A_piItm0YG7_0),.clk(gclk));
	jdff dff_A_uzv6tZZ44_0(.dout(w_dff_A_07i9yxNv3_0),.din(w_dff_A_uzv6tZZ44_0),.clk(gclk));
	jdff dff_A_07i9yxNv3_0(.dout(w_dff_A_mX6H77rn3_0),.din(w_dff_A_07i9yxNv3_0),.clk(gclk));
	jdff dff_A_mX6H77rn3_0(.dout(w_dff_A_p7gXbnKb1_0),.din(w_dff_A_mX6H77rn3_0),.clk(gclk));
	jdff dff_A_p7gXbnKb1_0(.dout(w_dff_A_b46PmH9S7_0),.din(w_dff_A_p7gXbnKb1_0),.clk(gclk));
	jdff dff_A_b46PmH9S7_0(.dout(w_dff_A_DwpVE6mL5_0),.din(w_dff_A_b46PmH9S7_0),.clk(gclk));
	jdff dff_A_DwpVE6mL5_0(.dout(w_dff_A_915szK9h8_0),.din(w_dff_A_DwpVE6mL5_0),.clk(gclk));
	jdff dff_A_915szK9h8_0(.dout(w_dff_A_lQtbeT7y7_0),.din(w_dff_A_915szK9h8_0),.clk(gclk));
	jdff dff_A_lQtbeT7y7_0(.dout(w_dff_A_MJ0uYOoe6_0),.din(w_dff_A_lQtbeT7y7_0),.clk(gclk));
	jdff dff_A_MJ0uYOoe6_0(.dout(w_dff_A_FNQX1sKs5_0),.din(w_dff_A_MJ0uYOoe6_0),.clk(gclk));
	jdff dff_A_FNQX1sKs5_0(.dout(w_dff_A_jnRz40jd9_0),.din(w_dff_A_FNQX1sKs5_0),.clk(gclk));
	jdff dff_A_jnRz40jd9_0(.dout(w_dff_A_OnAJmf9o9_0),.din(w_dff_A_jnRz40jd9_0),.clk(gclk));
	jdff dff_A_OnAJmf9o9_0(.dout(w_dff_A_knavpqI26_0),.din(w_dff_A_OnAJmf9o9_0),.clk(gclk));
	jdff dff_A_knavpqI26_0(.dout(w_dff_A_kQK27dXJ2_0),.din(w_dff_A_knavpqI26_0),.clk(gclk));
	jdff dff_A_kQK27dXJ2_0(.dout(w_dff_A_l7Fvddct6_0),.din(w_dff_A_kQK27dXJ2_0),.clk(gclk));
	jdff dff_A_l7Fvddct6_0(.dout(w_dff_A_le0X9G589_0),.din(w_dff_A_l7Fvddct6_0),.clk(gclk));
	jdff dff_A_le0X9G589_0(.dout(w_dff_A_jphLi6kC3_0),.din(w_dff_A_le0X9G589_0),.clk(gclk));
	jdff dff_A_jphLi6kC3_0(.dout(w_dff_A_ZygH8nJ06_0),.din(w_dff_A_jphLi6kC3_0),.clk(gclk));
	jdff dff_A_ZygH8nJ06_0(.dout(w_dff_A_SYgmEh182_0),.din(w_dff_A_ZygH8nJ06_0),.clk(gclk));
	jdff dff_A_SYgmEh182_0(.dout(w_dff_A_1jPWKSFF8_0),.din(w_dff_A_SYgmEh182_0),.clk(gclk));
	jdff dff_A_1jPWKSFF8_0(.dout(w_dff_A_O9VFiXuI4_0),.din(w_dff_A_1jPWKSFF8_0),.clk(gclk));
	jdff dff_A_O9VFiXuI4_0(.dout(w_dff_A_KvTgUuRd4_0),.din(w_dff_A_O9VFiXuI4_0),.clk(gclk));
	jdff dff_A_KvTgUuRd4_0(.dout(w_dff_A_TbFnflIP9_0),.din(w_dff_A_KvTgUuRd4_0),.clk(gclk));
	jdff dff_A_TbFnflIP9_0(.dout(w_dff_A_shMaAjZz3_0),.din(w_dff_A_TbFnflIP9_0),.clk(gclk));
	jdff dff_A_shMaAjZz3_0(.dout(w_dff_A_yDHJuRpm3_0),.din(w_dff_A_shMaAjZz3_0),.clk(gclk));
	jdff dff_A_yDHJuRpm3_0(.dout(w_dff_A_4V0cJoRk8_0),.din(w_dff_A_yDHJuRpm3_0),.clk(gclk));
	jdff dff_A_4V0cJoRk8_0(.dout(w_dff_A_UNa3qPhz6_0),.din(w_dff_A_4V0cJoRk8_0),.clk(gclk));
	jdff dff_A_UNa3qPhz6_0(.dout(w_dff_A_fv0KZ2QH1_0),.din(w_dff_A_UNa3qPhz6_0),.clk(gclk));
	jdff dff_A_fv0KZ2QH1_0(.dout(w_dff_A_DBhMB6uc9_0),.din(w_dff_A_fv0KZ2QH1_0),.clk(gclk));
	jdff dff_A_DBhMB6uc9_0(.dout(w_dff_A_tZewAjMR5_0),.din(w_dff_A_DBhMB6uc9_0),.clk(gclk));
	jdff dff_A_tZewAjMR5_0(.dout(w_dff_A_DYovrw3X8_0),.din(w_dff_A_tZewAjMR5_0),.clk(gclk));
	jdff dff_A_DYovrw3X8_0(.dout(w_dff_A_Mek4U3ad6_0),.din(w_dff_A_DYovrw3X8_0),.clk(gclk));
	jdff dff_A_Mek4U3ad6_0(.dout(w_dff_A_VQLu4bnW8_0),.din(w_dff_A_Mek4U3ad6_0),.clk(gclk));
	jdff dff_A_VQLu4bnW8_0(.dout(w_dff_A_b5cjhAkL5_0),.din(w_dff_A_VQLu4bnW8_0),.clk(gclk));
	jdff dff_A_b5cjhAkL5_0(.dout(w_dff_A_JArkOiN17_0),.din(w_dff_A_b5cjhAkL5_0),.clk(gclk));
	jdff dff_A_JArkOiN17_0(.dout(w_dff_A_7MLLdLaI6_0),.din(w_dff_A_JArkOiN17_0),.clk(gclk));
	jdff dff_A_7MLLdLaI6_0(.dout(w_dff_A_MNkbdDQn4_0),.din(w_dff_A_7MLLdLaI6_0),.clk(gclk));
	jdff dff_A_MNkbdDQn4_0(.dout(w_dff_A_wzovpAgm6_0),.din(w_dff_A_MNkbdDQn4_0),.clk(gclk));
	jdff dff_A_wzovpAgm6_0(.dout(w_dff_A_U7lON1Fz3_0),.din(w_dff_A_wzovpAgm6_0),.clk(gclk));
	jdff dff_A_U7lON1Fz3_0(.dout(w_dff_A_biKLaRG36_0),.din(w_dff_A_U7lON1Fz3_0),.clk(gclk));
	jdff dff_A_biKLaRG36_0(.dout(w_dff_A_8lnx8x7n9_0),.din(w_dff_A_biKLaRG36_0),.clk(gclk));
	jdff dff_A_8lnx8x7n9_0(.dout(f27),.din(w_dff_A_8lnx8x7n9_0),.clk(gclk));
	jdff dff_A_7BbhU6Rh4_2(.dout(w_dff_A_LfqjixaV1_0),.din(w_dff_A_7BbhU6Rh4_2),.clk(gclk));
	jdff dff_A_LfqjixaV1_0(.dout(w_dff_A_CzG9471b4_0),.din(w_dff_A_LfqjixaV1_0),.clk(gclk));
	jdff dff_A_CzG9471b4_0(.dout(w_dff_A_r9azPEcN4_0),.din(w_dff_A_CzG9471b4_0),.clk(gclk));
	jdff dff_A_r9azPEcN4_0(.dout(w_dff_A_Pdgj5oec8_0),.din(w_dff_A_r9azPEcN4_0),.clk(gclk));
	jdff dff_A_Pdgj5oec8_0(.dout(w_dff_A_Q2gWDUY78_0),.din(w_dff_A_Pdgj5oec8_0),.clk(gclk));
	jdff dff_A_Q2gWDUY78_0(.dout(w_dff_A_ptNq7EdW8_0),.din(w_dff_A_Q2gWDUY78_0),.clk(gclk));
	jdff dff_A_ptNq7EdW8_0(.dout(w_dff_A_UdO4ShWI5_0),.din(w_dff_A_ptNq7EdW8_0),.clk(gclk));
	jdff dff_A_UdO4ShWI5_0(.dout(w_dff_A_ubKkkyBH8_0),.din(w_dff_A_UdO4ShWI5_0),.clk(gclk));
	jdff dff_A_ubKkkyBH8_0(.dout(w_dff_A_tP9rBEk95_0),.din(w_dff_A_ubKkkyBH8_0),.clk(gclk));
	jdff dff_A_tP9rBEk95_0(.dout(w_dff_A_JUBlxMuu0_0),.din(w_dff_A_tP9rBEk95_0),.clk(gclk));
	jdff dff_A_JUBlxMuu0_0(.dout(w_dff_A_rTagaEW07_0),.din(w_dff_A_JUBlxMuu0_0),.clk(gclk));
	jdff dff_A_rTagaEW07_0(.dout(w_dff_A_Gwi2Ek4F6_0),.din(w_dff_A_rTagaEW07_0),.clk(gclk));
	jdff dff_A_Gwi2Ek4F6_0(.dout(w_dff_A_mWuA76ee5_0),.din(w_dff_A_Gwi2Ek4F6_0),.clk(gclk));
	jdff dff_A_mWuA76ee5_0(.dout(w_dff_A_hRvtBTWC3_0),.din(w_dff_A_mWuA76ee5_0),.clk(gclk));
	jdff dff_A_hRvtBTWC3_0(.dout(w_dff_A_9NKhObai5_0),.din(w_dff_A_hRvtBTWC3_0),.clk(gclk));
	jdff dff_A_9NKhObai5_0(.dout(w_dff_A_ms7K6n391_0),.din(w_dff_A_9NKhObai5_0),.clk(gclk));
	jdff dff_A_ms7K6n391_0(.dout(w_dff_A_2pCs6kaU2_0),.din(w_dff_A_ms7K6n391_0),.clk(gclk));
	jdff dff_A_2pCs6kaU2_0(.dout(w_dff_A_VcXGayQJ3_0),.din(w_dff_A_2pCs6kaU2_0),.clk(gclk));
	jdff dff_A_VcXGayQJ3_0(.dout(w_dff_A_Xomayz0X0_0),.din(w_dff_A_VcXGayQJ3_0),.clk(gclk));
	jdff dff_A_Xomayz0X0_0(.dout(w_dff_A_4zi2NolQ5_0),.din(w_dff_A_Xomayz0X0_0),.clk(gclk));
	jdff dff_A_4zi2NolQ5_0(.dout(w_dff_A_EDA33RRY5_0),.din(w_dff_A_4zi2NolQ5_0),.clk(gclk));
	jdff dff_A_EDA33RRY5_0(.dout(w_dff_A_EOLFbbpO6_0),.din(w_dff_A_EDA33RRY5_0),.clk(gclk));
	jdff dff_A_EOLFbbpO6_0(.dout(w_dff_A_wRLglZug3_0),.din(w_dff_A_EOLFbbpO6_0),.clk(gclk));
	jdff dff_A_wRLglZug3_0(.dout(w_dff_A_mAvKB8PR2_0),.din(w_dff_A_wRLglZug3_0),.clk(gclk));
	jdff dff_A_mAvKB8PR2_0(.dout(w_dff_A_6siqoi348_0),.din(w_dff_A_mAvKB8PR2_0),.clk(gclk));
	jdff dff_A_6siqoi348_0(.dout(w_dff_A_aXlJ4mY71_0),.din(w_dff_A_6siqoi348_0),.clk(gclk));
	jdff dff_A_aXlJ4mY71_0(.dout(w_dff_A_pjUxnIH16_0),.din(w_dff_A_aXlJ4mY71_0),.clk(gclk));
	jdff dff_A_pjUxnIH16_0(.dout(w_dff_A_GLfpGtGX4_0),.din(w_dff_A_pjUxnIH16_0),.clk(gclk));
	jdff dff_A_GLfpGtGX4_0(.dout(w_dff_A_c4LuTLzM0_0),.din(w_dff_A_GLfpGtGX4_0),.clk(gclk));
	jdff dff_A_c4LuTLzM0_0(.dout(w_dff_A_BAqqw0lj6_0),.din(w_dff_A_c4LuTLzM0_0),.clk(gclk));
	jdff dff_A_BAqqw0lj6_0(.dout(w_dff_A_g8teRVBZ3_0),.din(w_dff_A_BAqqw0lj6_0),.clk(gclk));
	jdff dff_A_g8teRVBZ3_0(.dout(w_dff_A_vxhYtxqg9_0),.din(w_dff_A_g8teRVBZ3_0),.clk(gclk));
	jdff dff_A_vxhYtxqg9_0(.dout(w_dff_A_b8AYPQMS8_0),.din(w_dff_A_vxhYtxqg9_0),.clk(gclk));
	jdff dff_A_b8AYPQMS8_0(.dout(w_dff_A_SSDggxQG5_0),.din(w_dff_A_b8AYPQMS8_0),.clk(gclk));
	jdff dff_A_SSDggxQG5_0(.dout(w_dff_A_WPudK0A88_0),.din(w_dff_A_SSDggxQG5_0),.clk(gclk));
	jdff dff_A_WPudK0A88_0(.dout(w_dff_A_KCBKK5vs7_0),.din(w_dff_A_WPudK0A88_0),.clk(gclk));
	jdff dff_A_KCBKK5vs7_0(.dout(w_dff_A_7oTS1dvG8_0),.din(w_dff_A_KCBKK5vs7_0),.clk(gclk));
	jdff dff_A_7oTS1dvG8_0(.dout(w_dff_A_LJMblzin1_0),.din(w_dff_A_7oTS1dvG8_0),.clk(gclk));
	jdff dff_A_LJMblzin1_0(.dout(w_dff_A_YqGI9qVV9_0),.din(w_dff_A_LJMblzin1_0),.clk(gclk));
	jdff dff_A_YqGI9qVV9_0(.dout(w_dff_A_96B7wQuc6_0),.din(w_dff_A_YqGI9qVV9_0),.clk(gclk));
	jdff dff_A_96B7wQuc6_0(.dout(w_dff_A_lxNJOSC74_0),.din(w_dff_A_96B7wQuc6_0),.clk(gclk));
	jdff dff_A_lxNJOSC74_0(.dout(w_dff_A_QVdlgMqI3_0),.din(w_dff_A_lxNJOSC74_0),.clk(gclk));
	jdff dff_A_QVdlgMqI3_0(.dout(w_dff_A_X3plMJtd9_0),.din(w_dff_A_QVdlgMqI3_0),.clk(gclk));
	jdff dff_A_X3plMJtd9_0(.dout(w_dff_A_Jk0J2XwE4_0),.din(w_dff_A_X3plMJtd9_0),.clk(gclk));
	jdff dff_A_Jk0J2XwE4_0(.dout(w_dff_A_OdOqU9Bt2_0),.din(w_dff_A_Jk0J2XwE4_0),.clk(gclk));
	jdff dff_A_OdOqU9Bt2_0(.dout(w_dff_A_rIEtuhjR9_0),.din(w_dff_A_OdOqU9Bt2_0),.clk(gclk));
	jdff dff_A_rIEtuhjR9_0(.dout(w_dff_A_p3Obv0Sw7_0),.din(w_dff_A_rIEtuhjR9_0),.clk(gclk));
	jdff dff_A_p3Obv0Sw7_0(.dout(w_dff_A_T2tSucid8_0),.din(w_dff_A_p3Obv0Sw7_0),.clk(gclk));
	jdff dff_A_T2tSucid8_0(.dout(w_dff_A_RU3Ti26G0_0),.din(w_dff_A_T2tSucid8_0),.clk(gclk));
	jdff dff_A_RU3Ti26G0_0(.dout(w_dff_A_kHFJTMML4_0),.din(w_dff_A_RU3Ti26G0_0),.clk(gclk));
	jdff dff_A_kHFJTMML4_0(.dout(w_dff_A_SHxhsyGG1_0),.din(w_dff_A_kHFJTMML4_0),.clk(gclk));
	jdff dff_A_SHxhsyGG1_0(.dout(w_dff_A_g72auxyq1_0),.din(w_dff_A_SHxhsyGG1_0),.clk(gclk));
	jdff dff_A_g72auxyq1_0(.dout(w_dff_A_j3Hgo9yH8_0),.din(w_dff_A_g72auxyq1_0),.clk(gclk));
	jdff dff_A_j3Hgo9yH8_0(.dout(w_dff_A_3iuzaVec6_0),.din(w_dff_A_j3Hgo9yH8_0),.clk(gclk));
	jdff dff_A_3iuzaVec6_0(.dout(w_dff_A_an3tkXxa8_0),.din(w_dff_A_3iuzaVec6_0),.clk(gclk));
	jdff dff_A_an3tkXxa8_0(.dout(w_dff_A_6PciCPRA1_0),.din(w_dff_A_an3tkXxa8_0),.clk(gclk));
	jdff dff_A_6PciCPRA1_0(.dout(w_dff_A_T998yKGk5_0),.din(w_dff_A_6PciCPRA1_0),.clk(gclk));
	jdff dff_A_T998yKGk5_0(.dout(w_dff_A_iBNgGZqc7_0),.din(w_dff_A_T998yKGk5_0),.clk(gclk));
	jdff dff_A_iBNgGZqc7_0(.dout(w_dff_A_Wx6HAjrJ9_0),.din(w_dff_A_iBNgGZqc7_0),.clk(gclk));
	jdff dff_A_Wx6HAjrJ9_0(.dout(w_dff_A_AmtJ0Lvy4_0),.din(w_dff_A_Wx6HAjrJ9_0),.clk(gclk));
	jdff dff_A_AmtJ0Lvy4_0(.dout(w_dff_A_iLT03WhG6_0),.din(w_dff_A_AmtJ0Lvy4_0),.clk(gclk));
	jdff dff_A_iLT03WhG6_0(.dout(w_dff_A_cCFA310V2_0),.din(w_dff_A_iLT03WhG6_0),.clk(gclk));
	jdff dff_A_cCFA310V2_0(.dout(w_dff_A_3BkecCwr9_0),.din(w_dff_A_cCFA310V2_0),.clk(gclk));
	jdff dff_A_3BkecCwr9_0(.dout(w_dff_A_TD3hJ0WH6_0),.din(w_dff_A_3BkecCwr9_0),.clk(gclk));
	jdff dff_A_TD3hJ0WH6_0(.dout(w_dff_A_La7zAyyV0_0),.din(w_dff_A_TD3hJ0WH6_0),.clk(gclk));
	jdff dff_A_La7zAyyV0_0(.dout(w_dff_A_WkkvUzwc0_0),.din(w_dff_A_La7zAyyV0_0),.clk(gclk));
	jdff dff_A_WkkvUzwc0_0(.dout(w_dff_A_MgnvXWx85_0),.din(w_dff_A_WkkvUzwc0_0),.clk(gclk));
	jdff dff_A_MgnvXWx85_0(.dout(w_dff_A_gahUMigD7_0),.din(w_dff_A_MgnvXWx85_0),.clk(gclk));
	jdff dff_A_gahUMigD7_0(.dout(w_dff_A_xLjB74ZW7_0),.din(w_dff_A_gahUMigD7_0),.clk(gclk));
	jdff dff_A_xLjB74ZW7_0(.dout(w_dff_A_FOiBFNYk7_0),.din(w_dff_A_xLjB74ZW7_0),.clk(gclk));
	jdff dff_A_FOiBFNYk7_0(.dout(w_dff_A_fIS3s7qB9_0),.din(w_dff_A_FOiBFNYk7_0),.clk(gclk));
	jdff dff_A_fIS3s7qB9_0(.dout(w_dff_A_1BufGXZm1_0),.din(w_dff_A_fIS3s7qB9_0),.clk(gclk));
	jdff dff_A_1BufGXZm1_0(.dout(w_dff_A_B1CbZCMp7_0),.din(w_dff_A_1BufGXZm1_0),.clk(gclk));
	jdff dff_A_B1CbZCMp7_0(.dout(w_dff_A_scuF2Pnb9_0),.din(w_dff_A_B1CbZCMp7_0),.clk(gclk));
	jdff dff_A_scuF2Pnb9_0(.dout(w_dff_A_W4kKV87n5_0),.din(w_dff_A_scuF2Pnb9_0),.clk(gclk));
	jdff dff_A_W4kKV87n5_0(.dout(w_dff_A_0qtbZQjT4_0),.din(w_dff_A_W4kKV87n5_0),.clk(gclk));
	jdff dff_A_0qtbZQjT4_0(.dout(w_dff_A_0wX0dJp43_0),.din(w_dff_A_0qtbZQjT4_0),.clk(gclk));
	jdff dff_A_0wX0dJp43_0(.dout(w_dff_A_N6EuIn5d5_0),.din(w_dff_A_0wX0dJp43_0),.clk(gclk));
	jdff dff_A_N6EuIn5d5_0(.dout(w_dff_A_mBWVEsDc6_0),.din(w_dff_A_N6EuIn5d5_0),.clk(gclk));
	jdff dff_A_mBWVEsDc6_0(.dout(w_dff_A_wyw8CGco8_0),.din(w_dff_A_mBWVEsDc6_0),.clk(gclk));
	jdff dff_A_wyw8CGco8_0(.dout(w_dff_A_XIoD1hcd4_0),.din(w_dff_A_wyw8CGco8_0),.clk(gclk));
	jdff dff_A_XIoD1hcd4_0(.dout(w_dff_A_0L0o0DIo3_0),.din(w_dff_A_XIoD1hcd4_0),.clk(gclk));
	jdff dff_A_0L0o0DIo3_0(.dout(w_dff_A_7zhPa08u0_0),.din(w_dff_A_0L0o0DIo3_0),.clk(gclk));
	jdff dff_A_7zhPa08u0_0(.dout(w_dff_A_GDXXn1gl2_0),.din(w_dff_A_7zhPa08u0_0),.clk(gclk));
	jdff dff_A_GDXXn1gl2_0(.dout(w_dff_A_bYiZELNT2_0),.din(w_dff_A_GDXXn1gl2_0),.clk(gclk));
	jdff dff_A_bYiZELNT2_0(.dout(w_dff_A_tJV84ufY1_0),.din(w_dff_A_bYiZELNT2_0),.clk(gclk));
	jdff dff_A_tJV84ufY1_0(.dout(w_dff_A_Nd6E7wDl2_0),.din(w_dff_A_tJV84ufY1_0),.clk(gclk));
	jdff dff_A_Nd6E7wDl2_0(.dout(w_dff_A_gUiLEGFE7_0),.din(w_dff_A_Nd6E7wDl2_0),.clk(gclk));
	jdff dff_A_gUiLEGFE7_0(.dout(w_dff_A_W0ruTNHa6_0),.din(w_dff_A_gUiLEGFE7_0),.clk(gclk));
	jdff dff_A_W0ruTNHa6_0(.dout(w_dff_A_GbwNOgds9_0),.din(w_dff_A_W0ruTNHa6_0),.clk(gclk));
	jdff dff_A_GbwNOgds9_0(.dout(w_dff_A_Yx9e2PyO5_0),.din(w_dff_A_GbwNOgds9_0),.clk(gclk));
	jdff dff_A_Yx9e2PyO5_0(.dout(w_dff_A_SW6Hhg3R3_0),.din(w_dff_A_Yx9e2PyO5_0),.clk(gclk));
	jdff dff_A_SW6Hhg3R3_0(.dout(w_dff_A_OMKRgBxR8_0),.din(w_dff_A_SW6Hhg3R3_0),.clk(gclk));
	jdff dff_A_OMKRgBxR8_0(.dout(w_dff_A_QOgItMQH7_0),.din(w_dff_A_OMKRgBxR8_0),.clk(gclk));
	jdff dff_A_QOgItMQH7_0(.dout(w_dff_A_cqMWJ4D96_0),.din(w_dff_A_QOgItMQH7_0),.clk(gclk));
	jdff dff_A_cqMWJ4D96_0(.dout(w_dff_A_kNwMTneU3_0),.din(w_dff_A_cqMWJ4D96_0),.clk(gclk));
	jdff dff_A_kNwMTneU3_0(.dout(w_dff_A_pQd90E2v8_0),.din(w_dff_A_kNwMTneU3_0),.clk(gclk));
	jdff dff_A_pQd90E2v8_0(.dout(w_dff_A_RaNHooAH3_0),.din(w_dff_A_pQd90E2v8_0),.clk(gclk));
	jdff dff_A_RaNHooAH3_0(.dout(f28),.din(w_dff_A_RaNHooAH3_0),.clk(gclk));
	jdff dff_A_MfypuXxv4_2(.dout(w_dff_A_zdOlqrlj4_0),.din(w_dff_A_MfypuXxv4_2),.clk(gclk));
	jdff dff_A_zdOlqrlj4_0(.dout(w_dff_A_42fAdlNi0_0),.din(w_dff_A_zdOlqrlj4_0),.clk(gclk));
	jdff dff_A_42fAdlNi0_0(.dout(w_dff_A_p9M1fOqB7_0),.din(w_dff_A_42fAdlNi0_0),.clk(gclk));
	jdff dff_A_p9M1fOqB7_0(.dout(w_dff_A_aundsJR19_0),.din(w_dff_A_p9M1fOqB7_0),.clk(gclk));
	jdff dff_A_aundsJR19_0(.dout(w_dff_A_jlRrOq8l8_0),.din(w_dff_A_aundsJR19_0),.clk(gclk));
	jdff dff_A_jlRrOq8l8_0(.dout(w_dff_A_57Jc3TMY4_0),.din(w_dff_A_jlRrOq8l8_0),.clk(gclk));
	jdff dff_A_57Jc3TMY4_0(.dout(w_dff_A_fBVi7L3t4_0),.din(w_dff_A_57Jc3TMY4_0),.clk(gclk));
	jdff dff_A_fBVi7L3t4_0(.dout(w_dff_A_TQQ8eY0j7_0),.din(w_dff_A_fBVi7L3t4_0),.clk(gclk));
	jdff dff_A_TQQ8eY0j7_0(.dout(w_dff_A_cQ2JmozW7_0),.din(w_dff_A_TQQ8eY0j7_0),.clk(gclk));
	jdff dff_A_cQ2JmozW7_0(.dout(w_dff_A_3jynR71t7_0),.din(w_dff_A_cQ2JmozW7_0),.clk(gclk));
	jdff dff_A_3jynR71t7_0(.dout(w_dff_A_QEwdM94c7_0),.din(w_dff_A_3jynR71t7_0),.clk(gclk));
	jdff dff_A_QEwdM94c7_0(.dout(w_dff_A_a2MCaISr1_0),.din(w_dff_A_QEwdM94c7_0),.clk(gclk));
	jdff dff_A_a2MCaISr1_0(.dout(w_dff_A_malu6XMK8_0),.din(w_dff_A_a2MCaISr1_0),.clk(gclk));
	jdff dff_A_malu6XMK8_0(.dout(w_dff_A_IEqFLfRv0_0),.din(w_dff_A_malu6XMK8_0),.clk(gclk));
	jdff dff_A_IEqFLfRv0_0(.dout(w_dff_A_RBHYtUxk6_0),.din(w_dff_A_IEqFLfRv0_0),.clk(gclk));
	jdff dff_A_RBHYtUxk6_0(.dout(w_dff_A_iRyGJHqH5_0),.din(w_dff_A_RBHYtUxk6_0),.clk(gclk));
	jdff dff_A_iRyGJHqH5_0(.dout(w_dff_A_ZZbYLUlh6_0),.din(w_dff_A_iRyGJHqH5_0),.clk(gclk));
	jdff dff_A_ZZbYLUlh6_0(.dout(w_dff_A_QDjTkkt51_0),.din(w_dff_A_ZZbYLUlh6_0),.clk(gclk));
	jdff dff_A_QDjTkkt51_0(.dout(w_dff_A_I3djsEor7_0),.din(w_dff_A_QDjTkkt51_0),.clk(gclk));
	jdff dff_A_I3djsEor7_0(.dout(w_dff_A_wFNrXV636_0),.din(w_dff_A_I3djsEor7_0),.clk(gclk));
	jdff dff_A_wFNrXV636_0(.dout(w_dff_A_QzkpQ2G45_0),.din(w_dff_A_wFNrXV636_0),.clk(gclk));
	jdff dff_A_QzkpQ2G45_0(.dout(w_dff_A_lXLczKgJ3_0),.din(w_dff_A_QzkpQ2G45_0),.clk(gclk));
	jdff dff_A_lXLczKgJ3_0(.dout(w_dff_A_j4EINsUi7_0),.din(w_dff_A_lXLczKgJ3_0),.clk(gclk));
	jdff dff_A_j4EINsUi7_0(.dout(w_dff_A_h5xR87ZD9_0),.din(w_dff_A_j4EINsUi7_0),.clk(gclk));
	jdff dff_A_h5xR87ZD9_0(.dout(w_dff_A_E7yf5PqQ5_0),.din(w_dff_A_h5xR87ZD9_0),.clk(gclk));
	jdff dff_A_E7yf5PqQ5_0(.dout(w_dff_A_bpHb6z6x1_0),.din(w_dff_A_E7yf5PqQ5_0),.clk(gclk));
	jdff dff_A_bpHb6z6x1_0(.dout(w_dff_A_9ijk4KA32_0),.din(w_dff_A_bpHb6z6x1_0),.clk(gclk));
	jdff dff_A_9ijk4KA32_0(.dout(w_dff_A_i49vIbw44_0),.din(w_dff_A_9ijk4KA32_0),.clk(gclk));
	jdff dff_A_i49vIbw44_0(.dout(w_dff_A_N45sGNyX9_0),.din(w_dff_A_i49vIbw44_0),.clk(gclk));
	jdff dff_A_N45sGNyX9_0(.dout(w_dff_A_qX3iKmqT5_0),.din(w_dff_A_N45sGNyX9_0),.clk(gclk));
	jdff dff_A_qX3iKmqT5_0(.dout(w_dff_A_0mLib3Ic1_0),.din(w_dff_A_qX3iKmqT5_0),.clk(gclk));
	jdff dff_A_0mLib3Ic1_0(.dout(w_dff_A_3zze6v4u0_0),.din(w_dff_A_0mLib3Ic1_0),.clk(gclk));
	jdff dff_A_3zze6v4u0_0(.dout(w_dff_A_0noVYfVc3_0),.din(w_dff_A_3zze6v4u0_0),.clk(gclk));
	jdff dff_A_0noVYfVc3_0(.dout(w_dff_A_JsOfsVKn6_0),.din(w_dff_A_0noVYfVc3_0),.clk(gclk));
	jdff dff_A_JsOfsVKn6_0(.dout(w_dff_A_keJyqdro0_0),.din(w_dff_A_JsOfsVKn6_0),.clk(gclk));
	jdff dff_A_keJyqdro0_0(.dout(w_dff_A_Rl8vP1is3_0),.din(w_dff_A_keJyqdro0_0),.clk(gclk));
	jdff dff_A_Rl8vP1is3_0(.dout(w_dff_A_KR1HlduH4_0),.din(w_dff_A_Rl8vP1is3_0),.clk(gclk));
	jdff dff_A_KR1HlduH4_0(.dout(w_dff_A_yt6d0OFb4_0),.din(w_dff_A_KR1HlduH4_0),.clk(gclk));
	jdff dff_A_yt6d0OFb4_0(.dout(w_dff_A_JCZDrZux9_0),.din(w_dff_A_yt6d0OFb4_0),.clk(gclk));
	jdff dff_A_JCZDrZux9_0(.dout(w_dff_A_qk3nEWK17_0),.din(w_dff_A_JCZDrZux9_0),.clk(gclk));
	jdff dff_A_qk3nEWK17_0(.dout(w_dff_A_Z9KNJgDX7_0),.din(w_dff_A_qk3nEWK17_0),.clk(gclk));
	jdff dff_A_Z9KNJgDX7_0(.dout(w_dff_A_drbAPcoA8_0),.din(w_dff_A_Z9KNJgDX7_0),.clk(gclk));
	jdff dff_A_drbAPcoA8_0(.dout(w_dff_A_Qh0Fs5Pk3_0),.din(w_dff_A_drbAPcoA8_0),.clk(gclk));
	jdff dff_A_Qh0Fs5Pk3_0(.dout(w_dff_A_XeMNdYYl4_0),.din(w_dff_A_Qh0Fs5Pk3_0),.clk(gclk));
	jdff dff_A_XeMNdYYl4_0(.dout(w_dff_A_7kClTru31_0),.din(w_dff_A_XeMNdYYl4_0),.clk(gclk));
	jdff dff_A_7kClTru31_0(.dout(w_dff_A_3DXMF5qy5_0),.din(w_dff_A_7kClTru31_0),.clk(gclk));
	jdff dff_A_3DXMF5qy5_0(.dout(w_dff_A_aV71sszD9_0),.din(w_dff_A_3DXMF5qy5_0),.clk(gclk));
	jdff dff_A_aV71sszD9_0(.dout(w_dff_A_LzAA1TkY3_0),.din(w_dff_A_aV71sszD9_0),.clk(gclk));
	jdff dff_A_LzAA1TkY3_0(.dout(w_dff_A_Fdw45Z5A7_0),.din(w_dff_A_LzAA1TkY3_0),.clk(gclk));
	jdff dff_A_Fdw45Z5A7_0(.dout(w_dff_A_cn5LbfD82_0),.din(w_dff_A_Fdw45Z5A7_0),.clk(gclk));
	jdff dff_A_cn5LbfD82_0(.dout(w_dff_A_s8eDJzvw0_0),.din(w_dff_A_cn5LbfD82_0),.clk(gclk));
	jdff dff_A_s8eDJzvw0_0(.dout(w_dff_A_fF8YfCvq9_0),.din(w_dff_A_s8eDJzvw0_0),.clk(gclk));
	jdff dff_A_fF8YfCvq9_0(.dout(w_dff_A_mVi9qIpC7_0),.din(w_dff_A_fF8YfCvq9_0),.clk(gclk));
	jdff dff_A_mVi9qIpC7_0(.dout(w_dff_A_UOAuhCY19_0),.din(w_dff_A_mVi9qIpC7_0),.clk(gclk));
	jdff dff_A_UOAuhCY19_0(.dout(w_dff_A_ixGzX1ZG5_0),.din(w_dff_A_UOAuhCY19_0),.clk(gclk));
	jdff dff_A_ixGzX1ZG5_0(.dout(w_dff_A_xjvzFRTM7_0),.din(w_dff_A_ixGzX1ZG5_0),.clk(gclk));
	jdff dff_A_xjvzFRTM7_0(.dout(w_dff_A_3TgUbAwo5_0),.din(w_dff_A_xjvzFRTM7_0),.clk(gclk));
	jdff dff_A_3TgUbAwo5_0(.dout(w_dff_A_IOBOnBpN0_0),.din(w_dff_A_3TgUbAwo5_0),.clk(gclk));
	jdff dff_A_IOBOnBpN0_0(.dout(w_dff_A_aZHK1LBo3_0),.din(w_dff_A_IOBOnBpN0_0),.clk(gclk));
	jdff dff_A_aZHK1LBo3_0(.dout(w_dff_A_UlPb7xGx1_0),.din(w_dff_A_aZHK1LBo3_0),.clk(gclk));
	jdff dff_A_UlPb7xGx1_0(.dout(w_dff_A_3iSZb6iK8_0),.din(w_dff_A_UlPb7xGx1_0),.clk(gclk));
	jdff dff_A_3iSZb6iK8_0(.dout(w_dff_A_wIa54FeD1_0),.din(w_dff_A_3iSZb6iK8_0),.clk(gclk));
	jdff dff_A_wIa54FeD1_0(.dout(w_dff_A_NcGd930p7_0),.din(w_dff_A_wIa54FeD1_0),.clk(gclk));
	jdff dff_A_NcGd930p7_0(.dout(w_dff_A_Kf3VFY2b2_0),.din(w_dff_A_NcGd930p7_0),.clk(gclk));
	jdff dff_A_Kf3VFY2b2_0(.dout(w_dff_A_N3bVx1ge8_0),.din(w_dff_A_Kf3VFY2b2_0),.clk(gclk));
	jdff dff_A_N3bVx1ge8_0(.dout(w_dff_A_B8Vtbp0b0_0),.din(w_dff_A_N3bVx1ge8_0),.clk(gclk));
	jdff dff_A_B8Vtbp0b0_0(.dout(w_dff_A_duyq20ZB4_0),.din(w_dff_A_B8Vtbp0b0_0),.clk(gclk));
	jdff dff_A_duyq20ZB4_0(.dout(w_dff_A_Kl1xbcvj7_0),.din(w_dff_A_duyq20ZB4_0),.clk(gclk));
	jdff dff_A_Kl1xbcvj7_0(.dout(w_dff_A_ZpfVUx930_0),.din(w_dff_A_Kl1xbcvj7_0),.clk(gclk));
	jdff dff_A_ZpfVUx930_0(.dout(w_dff_A_p8UVQvug3_0),.din(w_dff_A_ZpfVUx930_0),.clk(gclk));
	jdff dff_A_p8UVQvug3_0(.dout(w_dff_A_C4bcxwWo5_0),.din(w_dff_A_p8UVQvug3_0),.clk(gclk));
	jdff dff_A_C4bcxwWo5_0(.dout(w_dff_A_XulejHAB3_0),.din(w_dff_A_C4bcxwWo5_0),.clk(gclk));
	jdff dff_A_XulejHAB3_0(.dout(w_dff_A_VsEKWqlu7_0),.din(w_dff_A_XulejHAB3_0),.clk(gclk));
	jdff dff_A_VsEKWqlu7_0(.dout(w_dff_A_eVRwYDbN9_0),.din(w_dff_A_VsEKWqlu7_0),.clk(gclk));
	jdff dff_A_eVRwYDbN9_0(.dout(w_dff_A_mWXkjwms5_0),.din(w_dff_A_eVRwYDbN9_0),.clk(gclk));
	jdff dff_A_mWXkjwms5_0(.dout(w_dff_A_v5ozceBS8_0),.din(w_dff_A_mWXkjwms5_0),.clk(gclk));
	jdff dff_A_v5ozceBS8_0(.dout(w_dff_A_0f6rSJEj0_0),.din(w_dff_A_v5ozceBS8_0),.clk(gclk));
	jdff dff_A_0f6rSJEj0_0(.dout(w_dff_A_g9mNr2lb5_0),.din(w_dff_A_0f6rSJEj0_0),.clk(gclk));
	jdff dff_A_g9mNr2lb5_0(.dout(w_dff_A_amNppAe01_0),.din(w_dff_A_g9mNr2lb5_0),.clk(gclk));
	jdff dff_A_amNppAe01_0(.dout(w_dff_A_fHmNsu873_0),.din(w_dff_A_amNppAe01_0),.clk(gclk));
	jdff dff_A_fHmNsu873_0(.dout(w_dff_A_u8klzVdW5_0),.din(w_dff_A_fHmNsu873_0),.clk(gclk));
	jdff dff_A_u8klzVdW5_0(.dout(w_dff_A_MXTUzSFv4_0),.din(w_dff_A_u8klzVdW5_0),.clk(gclk));
	jdff dff_A_MXTUzSFv4_0(.dout(w_dff_A_RWccJ74E2_0),.din(w_dff_A_MXTUzSFv4_0),.clk(gclk));
	jdff dff_A_RWccJ74E2_0(.dout(w_dff_A_lEp38xPX1_0),.din(w_dff_A_RWccJ74E2_0),.clk(gclk));
	jdff dff_A_lEp38xPX1_0(.dout(w_dff_A_UgxBCfoA6_0),.din(w_dff_A_lEp38xPX1_0),.clk(gclk));
	jdff dff_A_UgxBCfoA6_0(.dout(w_dff_A_EGnWsPIg8_0),.din(w_dff_A_UgxBCfoA6_0),.clk(gclk));
	jdff dff_A_EGnWsPIg8_0(.dout(w_dff_A_iQZxSYWs6_0),.din(w_dff_A_EGnWsPIg8_0),.clk(gclk));
	jdff dff_A_iQZxSYWs6_0(.dout(w_dff_A_y9gAim2U1_0),.din(w_dff_A_iQZxSYWs6_0),.clk(gclk));
	jdff dff_A_y9gAim2U1_0(.dout(w_dff_A_St7HXQh97_0),.din(w_dff_A_y9gAim2U1_0),.clk(gclk));
	jdff dff_A_St7HXQh97_0(.dout(w_dff_A_RXPWyulM1_0),.din(w_dff_A_St7HXQh97_0),.clk(gclk));
	jdff dff_A_RXPWyulM1_0(.dout(w_dff_A_9vfmBxph2_0),.din(w_dff_A_RXPWyulM1_0),.clk(gclk));
	jdff dff_A_9vfmBxph2_0(.dout(w_dff_A_lX9CmjXJ9_0),.din(w_dff_A_9vfmBxph2_0),.clk(gclk));
	jdff dff_A_lX9CmjXJ9_0(.dout(w_dff_A_rWTbbxb21_0),.din(w_dff_A_lX9CmjXJ9_0),.clk(gclk));
	jdff dff_A_rWTbbxb21_0(.dout(w_dff_A_a3s3Pj7Q9_0),.din(w_dff_A_rWTbbxb21_0),.clk(gclk));
	jdff dff_A_a3s3Pj7Q9_0(.dout(w_dff_A_Q5uI4hct1_0),.din(w_dff_A_a3s3Pj7Q9_0),.clk(gclk));
	jdff dff_A_Q5uI4hct1_0(.dout(w_dff_A_Qwv4GP0i3_0),.din(w_dff_A_Q5uI4hct1_0),.clk(gclk));
	jdff dff_A_Qwv4GP0i3_0(.dout(w_dff_A_P9WI9vn16_0),.din(w_dff_A_Qwv4GP0i3_0),.clk(gclk));
	jdff dff_A_P9WI9vn16_0(.dout(f29),.din(w_dff_A_P9WI9vn16_0),.clk(gclk));
	jdff dff_A_m45eyEAd4_2(.dout(w_dff_A_Wx2kalZ99_0),.din(w_dff_A_m45eyEAd4_2),.clk(gclk));
	jdff dff_A_Wx2kalZ99_0(.dout(w_dff_A_EvLJEHTp5_0),.din(w_dff_A_Wx2kalZ99_0),.clk(gclk));
	jdff dff_A_EvLJEHTp5_0(.dout(w_dff_A_XlS8aBvx3_0),.din(w_dff_A_EvLJEHTp5_0),.clk(gclk));
	jdff dff_A_XlS8aBvx3_0(.dout(w_dff_A_v0r4CZtO2_0),.din(w_dff_A_XlS8aBvx3_0),.clk(gclk));
	jdff dff_A_v0r4CZtO2_0(.dout(w_dff_A_Penvwuy62_0),.din(w_dff_A_v0r4CZtO2_0),.clk(gclk));
	jdff dff_A_Penvwuy62_0(.dout(w_dff_A_RT75uAev7_0),.din(w_dff_A_Penvwuy62_0),.clk(gclk));
	jdff dff_A_RT75uAev7_0(.dout(w_dff_A_1P7i1joJ7_0),.din(w_dff_A_RT75uAev7_0),.clk(gclk));
	jdff dff_A_1P7i1joJ7_0(.dout(w_dff_A_PoWmjduH7_0),.din(w_dff_A_1P7i1joJ7_0),.clk(gclk));
	jdff dff_A_PoWmjduH7_0(.dout(w_dff_A_QoIRXqco0_0),.din(w_dff_A_PoWmjduH7_0),.clk(gclk));
	jdff dff_A_QoIRXqco0_0(.dout(w_dff_A_ziKmwNuf6_0),.din(w_dff_A_QoIRXqco0_0),.clk(gclk));
	jdff dff_A_ziKmwNuf6_0(.dout(w_dff_A_Iito4yRU6_0),.din(w_dff_A_ziKmwNuf6_0),.clk(gclk));
	jdff dff_A_Iito4yRU6_0(.dout(w_dff_A_vJsyDuPA2_0),.din(w_dff_A_Iito4yRU6_0),.clk(gclk));
	jdff dff_A_vJsyDuPA2_0(.dout(w_dff_A_CpnoYG6B6_0),.din(w_dff_A_vJsyDuPA2_0),.clk(gclk));
	jdff dff_A_CpnoYG6B6_0(.dout(w_dff_A_1jpseo286_0),.din(w_dff_A_CpnoYG6B6_0),.clk(gclk));
	jdff dff_A_1jpseo286_0(.dout(w_dff_A_nLWBu4Cq4_0),.din(w_dff_A_1jpseo286_0),.clk(gclk));
	jdff dff_A_nLWBu4Cq4_0(.dout(w_dff_A_bAqmkQ7I7_0),.din(w_dff_A_nLWBu4Cq4_0),.clk(gclk));
	jdff dff_A_bAqmkQ7I7_0(.dout(w_dff_A_uluriX6K5_0),.din(w_dff_A_bAqmkQ7I7_0),.clk(gclk));
	jdff dff_A_uluriX6K5_0(.dout(w_dff_A_RstTxIl16_0),.din(w_dff_A_uluriX6K5_0),.clk(gclk));
	jdff dff_A_RstTxIl16_0(.dout(w_dff_A_9f3Ev0xc5_0),.din(w_dff_A_RstTxIl16_0),.clk(gclk));
	jdff dff_A_9f3Ev0xc5_0(.dout(w_dff_A_MNhZlhs06_0),.din(w_dff_A_9f3Ev0xc5_0),.clk(gclk));
	jdff dff_A_MNhZlhs06_0(.dout(w_dff_A_5FB3KJOx8_0),.din(w_dff_A_MNhZlhs06_0),.clk(gclk));
	jdff dff_A_5FB3KJOx8_0(.dout(w_dff_A_JVTUOxxr4_0),.din(w_dff_A_5FB3KJOx8_0),.clk(gclk));
	jdff dff_A_JVTUOxxr4_0(.dout(w_dff_A_V1OTSyzX4_0),.din(w_dff_A_JVTUOxxr4_0),.clk(gclk));
	jdff dff_A_V1OTSyzX4_0(.dout(w_dff_A_4OoHZF5N3_0),.din(w_dff_A_V1OTSyzX4_0),.clk(gclk));
	jdff dff_A_4OoHZF5N3_0(.dout(w_dff_A_vXNH0Y9J2_0),.din(w_dff_A_4OoHZF5N3_0),.clk(gclk));
	jdff dff_A_vXNH0Y9J2_0(.dout(w_dff_A_hvv1rbL06_0),.din(w_dff_A_vXNH0Y9J2_0),.clk(gclk));
	jdff dff_A_hvv1rbL06_0(.dout(w_dff_A_dvYP2lsa1_0),.din(w_dff_A_hvv1rbL06_0),.clk(gclk));
	jdff dff_A_dvYP2lsa1_0(.dout(w_dff_A_ARgXA8Kr9_0),.din(w_dff_A_dvYP2lsa1_0),.clk(gclk));
	jdff dff_A_ARgXA8Kr9_0(.dout(w_dff_A_Us18klBO3_0),.din(w_dff_A_ARgXA8Kr9_0),.clk(gclk));
	jdff dff_A_Us18klBO3_0(.dout(w_dff_A_Bz56m29g8_0),.din(w_dff_A_Us18klBO3_0),.clk(gclk));
	jdff dff_A_Bz56m29g8_0(.dout(w_dff_A_buRIKoaZ1_0),.din(w_dff_A_Bz56m29g8_0),.clk(gclk));
	jdff dff_A_buRIKoaZ1_0(.dout(w_dff_A_VAWnMiBM9_0),.din(w_dff_A_buRIKoaZ1_0),.clk(gclk));
	jdff dff_A_VAWnMiBM9_0(.dout(w_dff_A_cv5Zs6vR2_0),.din(w_dff_A_VAWnMiBM9_0),.clk(gclk));
	jdff dff_A_cv5Zs6vR2_0(.dout(w_dff_A_757iSOvs6_0),.din(w_dff_A_cv5Zs6vR2_0),.clk(gclk));
	jdff dff_A_757iSOvs6_0(.dout(w_dff_A_vs1lzyKN0_0),.din(w_dff_A_757iSOvs6_0),.clk(gclk));
	jdff dff_A_vs1lzyKN0_0(.dout(w_dff_A_snFj8Xpl5_0),.din(w_dff_A_vs1lzyKN0_0),.clk(gclk));
	jdff dff_A_snFj8Xpl5_0(.dout(w_dff_A_rtq30XW18_0),.din(w_dff_A_snFj8Xpl5_0),.clk(gclk));
	jdff dff_A_rtq30XW18_0(.dout(w_dff_A_x0DbNDtM6_0),.din(w_dff_A_rtq30XW18_0),.clk(gclk));
	jdff dff_A_x0DbNDtM6_0(.dout(w_dff_A_346KtL4V2_0),.din(w_dff_A_x0DbNDtM6_0),.clk(gclk));
	jdff dff_A_346KtL4V2_0(.dout(w_dff_A_xWrAODEW4_0),.din(w_dff_A_346KtL4V2_0),.clk(gclk));
	jdff dff_A_xWrAODEW4_0(.dout(w_dff_A_NsReiRRY4_0),.din(w_dff_A_xWrAODEW4_0),.clk(gclk));
	jdff dff_A_NsReiRRY4_0(.dout(w_dff_A_HnZohz3y1_0),.din(w_dff_A_NsReiRRY4_0),.clk(gclk));
	jdff dff_A_HnZohz3y1_0(.dout(w_dff_A_BT3erJOD0_0),.din(w_dff_A_HnZohz3y1_0),.clk(gclk));
	jdff dff_A_BT3erJOD0_0(.dout(w_dff_A_TboxvwgO8_0),.din(w_dff_A_BT3erJOD0_0),.clk(gclk));
	jdff dff_A_TboxvwgO8_0(.dout(w_dff_A_NO6JhiHs4_0),.din(w_dff_A_TboxvwgO8_0),.clk(gclk));
	jdff dff_A_NO6JhiHs4_0(.dout(w_dff_A_sdL7SRKG8_0),.din(w_dff_A_NO6JhiHs4_0),.clk(gclk));
	jdff dff_A_sdL7SRKG8_0(.dout(w_dff_A_AHAq9gor6_0),.din(w_dff_A_sdL7SRKG8_0),.clk(gclk));
	jdff dff_A_AHAq9gor6_0(.dout(w_dff_A_iBGnvnJm3_0),.din(w_dff_A_AHAq9gor6_0),.clk(gclk));
	jdff dff_A_iBGnvnJm3_0(.dout(w_dff_A_SPMYRRwN1_0),.din(w_dff_A_iBGnvnJm3_0),.clk(gclk));
	jdff dff_A_SPMYRRwN1_0(.dout(w_dff_A_UET1ivrO7_0),.din(w_dff_A_SPMYRRwN1_0),.clk(gclk));
	jdff dff_A_UET1ivrO7_0(.dout(w_dff_A_oBLNfSXw3_0),.din(w_dff_A_UET1ivrO7_0),.clk(gclk));
	jdff dff_A_oBLNfSXw3_0(.dout(w_dff_A_wHq79Frn5_0),.din(w_dff_A_oBLNfSXw3_0),.clk(gclk));
	jdff dff_A_wHq79Frn5_0(.dout(w_dff_A_ADugQLl23_0),.din(w_dff_A_wHq79Frn5_0),.clk(gclk));
	jdff dff_A_ADugQLl23_0(.dout(w_dff_A_SmTcV4mc6_0),.din(w_dff_A_ADugQLl23_0),.clk(gclk));
	jdff dff_A_SmTcV4mc6_0(.dout(w_dff_A_IXIcvFv44_0),.din(w_dff_A_SmTcV4mc6_0),.clk(gclk));
	jdff dff_A_IXIcvFv44_0(.dout(w_dff_A_o8PPN4bL5_0),.din(w_dff_A_IXIcvFv44_0),.clk(gclk));
	jdff dff_A_o8PPN4bL5_0(.dout(w_dff_A_heM0Ijud4_0),.din(w_dff_A_o8PPN4bL5_0),.clk(gclk));
	jdff dff_A_heM0Ijud4_0(.dout(w_dff_A_wO4uCGDJ5_0),.din(w_dff_A_heM0Ijud4_0),.clk(gclk));
	jdff dff_A_wO4uCGDJ5_0(.dout(w_dff_A_1MrudNvZ3_0),.din(w_dff_A_wO4uCGDJ5_0),.clk(gclk));
	jdff dff_A_1MrudNvZ3_0(.dout(w_dff_A_t7LQzEWn2_0),.din(w_dff_A_1MrudNvZ3_0),.clk(gclk));
	jdff dff_A_t7LQzEWn2_0(.dout(w_dff_A_ILTVRGTn0_0),.din(w_dff_A_t7LQzEWn2_0),.clk(gclk));
	jdff dff_A_ILTVRGTn0_0(.dout(w_dff_A_JNX0A4MM6_0),.din(w_dff_A_ILTVRGTn0_0),.clk(gclk));
	jdff dff_A_JNX0A4MM6_0(.dout(w_dff_A_PAEzTRqn5_0),.din(w_dff_A_JNX0A4MM6_0),.clk(gclk));
	jdff dff_A_PAEzTRqn5_0(.dout(w_dff_A_ybZFxMBl2_0),.din(w_dff_A_PAEzTRqn5_0),.clk(gclk));
	jdff dff_A_ybZFxMBl2_0(.dout(w_dff_A_jrz5Vp8X8_0),.din(w_dff_A_ybZFxMBl2_0),.clk(gclk));
	jdff dff_A_jrz5Vp8X8_0(.dout(w_dff_A_9BSXmlwp0_0),.din(w_dff_A_jrz5Vp8X8_0),.clk(gclk));
	jdff dff_A_9BSXmlwp0_0(.dout(w_dff_A_b3eRhrYR7_0),.din(w_dff_A_9BSXmlwp0_0),.clk(gclk));
	jdff dff_A_b3eRhrYR7_0(.dout(w_dff_A_A2gXLhvE6_0),.din(w_dff_A_b3eRhrYR7_0),.clk(gclk));
	jdff dff_A_A2gXLhvE6_0(.dout(w_dff_A_9ko22dCP5_0),.din(w_dff_A_A2gXLhvE6_0),.clk(gclk));
	jdff dff_A_9ko22dCP5_0(.dout(w_dff_A_Mc04vk5y2_0),.din(w_dff_A_9ko22dCP5_0),.clk(gclk));
	jdff dff_A_Mc04vk5y2_0(.dout(w_dff_A_D4EhNa4Z4_0),.din(w_dff_A_Mc04vk5y2_0),.clk(gclk));
	jdff dff_A_D4EhNa4Z4_0(.dout(w_dff_A_I8X08HfC5_0),.din(w_dff_A_D4EhNa4Z4_0),.clk(gclk));
	jdff dff_A_I8X08HfC5_0(.dout(w_dff_A_CUzDiWlv2_0),.din(w_dff_A_I8X08HfC5_0),.clk(gclk));
	jdff dff_A_CUzDiWlv2_0(.dout(w_dff_A_mP6rND1o0_0),.din(w_dff_A_CUzDiWlv2_0),.clk(gclk));
	jdff dff_A_mP6rND1o0_0(.dout(w_dff_A_0EGG93Ll7_0),.din(w_dff_A_mP6rND1o0_0),.clk(gclk));
	jdff dff_A_0EGG93Ll7_0(.dout(w_dff_A_tg31B4vn7_0),.din(w_dff_A_0EGG93Ll7_0),.clk(gclk));
	jdff dff_A_tg31B4vn7_0(.dout(w_dff_A_ADCqHYX24_0),.din(w_dff_A_tg31B4vn7_0),.clk(gclk));
	jdff dff_A_ADCqHYX24_0(.dout(w_dff_A_hUd96aIE0_0),.din(w_dff_A_ADCqHYX24_0),.clk(gclk));
	jdff dff_A_hUd96aIE0_0(.dout(w_dff_A_d6y7TEOy1_0),.din(w_dff_A_hUd96aIE0_0),.clk(gclk));
	jdff dff_A_d6y7TEOy1_0(.dout(w_dff_A_PIVki6Pr5_0),.din(w_dff_A_d6y7TEOy1_0),.clk(gclk));
	jdff dff_A_PIVki6Pr5_0(.dout(w_dff_A_sSpUrxNE5_0),.din(w_dff_A_PIVki6Pr5_0),.clk(gclk));
	jdff dff_A_sSpUrxNE5_0(.dout(w_dff_A_sqMkZJiv2_0),.din(w_dff_A_sSpUrxNE5_0),.clk(gclk));
	jdff dff_A_sqMkZJiv2_0(.dout(w_dff_A_BJ6vWbrU0_0),.din(w_dff_A_sqMkZJiv2_0),.clk(gclk));
	jdff dff_A_BJ6vWbrU0_0(.dout(w_dff_A_LogdoRNP9_0),.din(w_dff_A_BJ6vWbrU0_0),.clk(gclk));
	jdff dff_A_LogdoRNP9_0(.dout(w_dff_A_LFxHf0T66_0),.din(w_dff_A_LogdoRNP9_0),.clk(gclk));
	jdff dff_A_LFxHf0T66_0(.dout(w_dff_A_8im5i1fx1_0),.din(w_dff_A_LFxHf0T66_0),.clk(gclk));
	jdff dff_A_8im5i1fx1_0(.dout(w_dff_A_wb0OGDCr6_0),.din(w_dff_A_8im5i1fx1_0),.clk(gclk));
	jdff dff_A_wb0OGDCr6_0(.dout(w_dff_A_a9tlW0gb4_0),.din(w_dff_A_wb0OGDCr6_0),.clk(gclk));
	jdff dff_A_a9tlW0gb4_0(.dout(w_dff_A_gXPX3UOS7_0),.din(w_dff_A_a9tlW0gb4_0),.clk(gclk));
	jdff dff_A_gXPX3UOS7_0(.dout(w_dff_A_qjwJ2l7P5_0),.din(w_dff_A_gXPX3UOS7_0),.clk(gclk));
	jdff dff_A_qjwJ2l7P5_0(.dout(w_dff_A_KQr5rPeX5_0),.din(w_dff_A_qjwJ2l7P5_0),.clk(gclk));
	jdff dff_A_KQr5rPeX5_0(.dout(w_dff_A_q30YGg2D0_0),.din(w_dff_A_KQr5rPeX5_0),.clk(gclk));
	jdff dff_A_q30YGg2D0_0(.dout(w_dff_A_ypL7O0d37_0),.din(w_dff_A_q30YGg2D0_0),.clk(gclk));
	jdff dff_A_ypL7O0d37_0(.dout(w_dff_A_PvH6dXMl1_0),.din(w_dff_A_ypL7O0d37_0),.clk(gclk));
	jdff dff_A_PvH6dXMl1_0(.dout(w_dff_A_L37lSGjN8_0),.din(w_dff_A_PvH6dXMl1_0),.clk(gclk));
	jdff dff_A_L37lSGjN8_0(.dout(w_dff_A_2iosBtlP0_0),.din(w_dff_A_L37lSGjN8_0),.clk(gclk));
	jdff dff_A_2iosBtlP0_0(.dout(f30),.din(w_dff_A_2iosBtlP0_0),.clk(gclk));
	jdff dff_A_HDJk7IDG5_2(.dout(w_dff_A_1KMSk5ni1_0),.din(w_dff_A_HDJk7IDG5_2),.clk(gclk));
	jdff dff_A_1KMSk5ni1_0(.dout(w_dff_A_LBQ3UZQS9_0),.din(w_dff_A_1KMSk5ni1_0),.clk(gclk));
	jdff dff_A_LBQ3UZQS9_0(.dout(w_dff_A_iIf5jTlO5_0),.din(w_dff_A_LBQ3UZQS9_0),.clk(gclk));
	jdff dff_A_iIf5jTlO5_0(.dout(w_dff_A_tkt2TCsn4_0),.din(w_dff_A_iIf5jTlO5_0),.clk(gclk));
	jdff dff_A_tkt2TCsn4_0(.dout(w_dff_A_QQpFWzS42_0),.din(w_dff_A_tkt2TCsn4_0),.clk(gclk));
	jdff dff_A_QQpFWzS42_0(.dout(w_dff_A_PSWnTCZk3_0),.din(w_dff_A_QQpFWzS42_0),.clk(gclk));
	jdff dff_A_PSWnTCZk3_0(.dout(w_dff_A_F4svAYcv1_0),.din(w_dff_A_PSWnTCZk3_0),.clk(gclk));
	jdff dff_A_F4svAYcv1_0(.dout(w_dff_A_Xv5YH3f47_0),.din(w_dff_A_F4svAYcv1_0),.clk(gclk));
	jdff dff_A_Xv5YH3f47_0(.dout(w_dff_A_v5s7pVLT7_0),.din(w_dff_A_Xv5YH3f47_0),.clk(gclk));
	jdff dff_A_v5s7pVLT7_0(.dout(w_dff_A_ZL25zWmZ5_0),.din(w_dff_A_v5s7pVLT7_0),.clk(gclk));
	jdff dff_A_ZL25zWmZ5_0(.dout(w_dff_A_52hs2BNB6_0),.din(w_dff_A_ZL25zWmZ5_0),.clk(gclk));
	jdff dff_A_52hs2BNB6_0(.dout(w_dff_A_Va2DCOu51_0),.din(w_dff_A_52hs2BNB6_0),.clk(gclk));
	jdff dff_A_Va2DCOu51_0(.dout(w_dff_A_6LX25aEP9_0),.din(w_dff_A_Va2DCOu51_0),.clk(gclk));
	jdff dff_A_6LX25aEP9_0(.dout(w_dff_A_hRtGsuXF9_0),.din(w_dff_A_6LX25aEP9_0),.clk(gclk));
	jdff dff_A_hRtGsuXF9_0(.dout(w_dff_A_RWPh9Knb3_0),.din(w_dff_A_hRtGsuXF9_0),.clk(gclk));
	jdff dff_A_RWPh9Knb3_0(.dout(w_dff_A_zyqUGTLi3_0),.din(w_dff_A_RWPh9Knb3_0),.clk(gclk));
	jdff dff_A_zyqUGTLi3_0(.dout(w_dff_A_Jgwcf05p3_0),.din(w_dff_A_zyqUGTLi3_0),.clk(gclk));
	jdff dff_A_Jgwcf05p3_0(.dout(w_dff_A_hwqlJh622_0),.din(w_dff_A_Jgwcf05p3_0),.clk(gclk));
	jdff dff_A_hwqlJh622_0(.dout(w_dff_A_jdzatfsk0_0),.din(w_dff_A_hwqlJh622_0),.clk(gclk));
	jdff dff_A_jdzatfsk0_0(.dout(w_dff_A_A9VfYmQc4_0),.din(w_dff_A_jdzatfsk0_0),.clk(gclk));
	jdff dff_A_A9VfYmQc4_0(.dout(w_dff_A_8LbLg9rS0_0),.din(w_dff_A_A9VfYmQc4_0),.clk(gclk));
	jdff dff_A_8LbLg9rS0_0(.dout(w_dff_A_Oz9q12bm0_0),.din(w_dff_A_8LbLg9rS0_0),.clk(gclk));
	jdff dff_A_Oz9q12bm0_0(.dout(w_dff_A_C8PnyTQS7_0),.din(w_dff_A_Oz9q12bm0_0),.clk(gclk));
	jdff dff_A_C8PnyTQS7_0(.dout(w_dff_A_Ku3Iad2r5_0),.din(w_dff_A_C8PnyTQS7_0),.clk(gclk));
	jdff dff_A_Ku3Iad2r5_0(.dout(w_dff_A_DqvvcaWd6_0),.din(w_dff_A_Ku3Iad2r5_0),.clk(gclk));
	jdff dff_A_DqvvcaWd6_0(.dout(w_dff_A_LN1mXno33_0),.din(w_dff_A_DqvvcaWd6_0),.clk(gclk));
	jdff dff_A_LN1mXno33_0(.dout(w_dff_A_xdNAfvfx0_0),.din(w_dff_A_LN1mXno33_0),.clk(gclk));
	jdff dff_A_xdNAfvfx0_0(.dout(w_dff_A_VLLhdAlN0_0),.din(w_dff_A_xdNAfvfx0_0),.clk(gclk));
	jdff dff_A_VLLhdAlN0_0(.dout(w_dff_A_8tA0gMe51_0),.din(w_dff_A_VLLhdAlN0_0),.clk(gclk));
	jdff dff_A_8tA0gMe51_0(.dout(w_dff_A_XKr94d6V6_0),.din(w_dff_A_8tA0gMe51_0),.clk(gclk));
	jdff dff_A_XKr94d6V6_0(.dout(w_dff_A_yQpU0N8V2_0),.din(w_dff_A_XKr94d6V6_0),.clk(gclk));
	jdff dff_A_yQpU0N8V2_0(.dout(w_dff_A_I2tGDJvr7_0),.din(w_dff_A_yQpU0N8V2_0),.clk(gclk));
	jdff dff_A_I2tGDJvr7_0(.dout(w_dff_A_4CUjPcWF2_0),.din(w_dff_A_I2tGDJvr7_0),.clk(gclk));
	jdff dff_A_4CUjPcWF2_0(.dout(w_dff_A_7vczdNd62_0),.din(w_dff_A_4CUjPcWF2_0),.clk(gclk));
	jdff dff_A_7vczdNd62_0(.dout(w_dff_A_Tfn1NlVW9_0),.din(w_dff_A_7vczdNd62_0),.clk(gclk));
	jdff dff_A_Tfn1NlVW9_0(.dout(w_dff_A_IcjXBsl08_0),.din(w_dff_A_Tfn1NlVW9_0),.clk(gclk));
	jdff dff_A_IcjXBsl08_0(.dout(w_dff_A_sf6HM8qM6_0),.din(w_dff_A_IcjXBsl08_0),.clk(gclk));
	jdff dff_A_sf6HM8qM6_0(.dout(w_dff_A_ANAj00bb7_0),.din(w_dff_A_sf6HM8qM6_0),.clk(gclk));
	jdff dff_A_ANAj00bb7_0(.dout(w_dff_A_Vu4xvi6C5_0),.din(w_dff_A_ANAj00bb7_0),.clk(gclk));
	jdff dff_A_Vu4xvi6C5_0(.dout(w_dff_A_P3IcNp4f3_0),.din(w_dff_A_Vu4xvi6C5_0),.clk(gclk));
	jdff dff_A_P3IcNp4f3_0(.dout(w_dff_A_RooPtbgS0_0),.din(w_dff_A_P3IcNp4f3_0),.clk(gclk));
	jdff dff_A_RooPtbgS0_0(.dout(w_dff_A_H6FfmfWI9_0),.din(w_dff_A_RooPtbgS0_0),.clk(gclk));
	jdff dff_A_H6FfmfWI9_0(.dout(w_dff_A_1yy10Jbe9_0),.din(w_dff_A_H6FfmfWI9_0),.clk(gclk));
	jdff dff_A_1yy10Jbe9_0(.dout(w_dff_A_lsjMGliR7_0),.din(w_dff_A_1yy10Jbe9_0),.clk(gclk));
	jdff dff_A_lsjMGliR7_0(.dout(w_dff_A_rgfsf5Yy5_0),.din(w_dff_A_lsjMGliR7_0),.clk(gclk));
	jdff dff_A_rgfsf5Yy5_0(.dout(w_dff_A_jr8yS74M4_0),.din(w_dff_A_rgfsf5Yy5_0),.clk(gclk));
	jdff dff_A_jr8yS74M4_0(.dout(w_dff_A_HVcr2GXv0_0),.din(w_dff_A_jr8yS74M4_0),.clk(gclk));
	jdff dff_A_HVcr2GXv0_0(.dout(w_dff_A_tdYKs75q0_0),.din(w_dff_A_HVcr2GXv0_0),.clk(gclk));
	jdff dff_A_tdYKs75q0_0(.dout(w_dff_A_QVztt8No4_0),.din(w_dff_A_tdYKs75q0_0),.clk(gclk));
	jdff dff_A_QVztt8No4_0(.dout(w_dff_A_9fYhtoq06_0),.din(w_dff_A_QVztt8No4_0),.clk(gclk));
	jdff dff_A_9fYhtoq06_0(.dout(w_dff_A_x0KInFsh7_0),.din(w_dff_A_9fYhtoq06_0),.clk(gclk));
	jdff dff_A_x0KInFsh7_0(.dout(w_dff_A_BCufJ05V9_0),.din(w_dff_A_x0KInFsh7_0),.clk(gclk));
	jdff dff_A_BCufJ05V9_0(.dout(w_dff_A_bdueen1P7_0),.din(w_dff_A_BCufJ05V9_0),.clk(gclk));
	jdff dff_A_bdueen1P7_0(.dout(w_dff_A_tUX7ATe30_0),.din(w_dff_A_bdueen1P7_0),.clk(gclk));
	jdff dff_A_tUX7ATe30_0(.dout(w_dff_A_C9jqr3F16_0),.din(w_dff_A_tUX7ATe30_0),.clk(gclk));
	jdff dff_A_C9jqr3F16_0(.dout(w_dff_A_Lft4Y8zd6_0),.din(w_dff_A_C9jqr3F16_0),.clk(gclk));
	jdff dff_A_Lft4Y8zd6_0(.dout(w_dff_A_h6lxUglG7_0),.din(w_dff_A_Lft4Y8zd6_0),.clk(gclk));
	jdff dff_A_h6lxUglG7_0(.dout(w_dff_A_DOeJSmlX8_0),.din(w_dff_A_h6lxUglG7_0),.clk(gclk));
	jdff dff_A_DOeJSmlX8_0(.dout(w_dff_A_DaUJHaia9_0),.din(w_dff_A_DOeJSmlX8_0),.clk(gclk));
	jdff dff_A_DaUJHaia9_0(.dout(w_dff_A_1pd9r7Lz1_0),.din(w_dff_A_DaUJHaia9_0),.clk(gclk));
	jdff dff_A_1pd9r7Lz1_0(.dout(w_dff_A_Zt2DUzCI9_0),.din(w_dff_A_1pd9r7Lz1_0),.clk(gclk));
	jdff dff_A_Zt2DUzCI9_0(.dout(w_dff_A_yAguPVvr3_0),.din(w_dff_A_Zt2DUzCI9_0),.clk(gclk));
	jdff dff_A_yAguPVvr3_0(.dout(w_dff_A_HD5dY2QX6_0),.din(w_dff_A_yAguPVvr3_0),.clk(gclk));
	jdff dff_A_HD5dY2QX6_0(.dout(w_dff_A_C8Vla8lD6_0),.din(w_dff_A_HD5dY2QX6_0),.clk(gclk));
	jdff dff_A_C8Vla8lD6_0(.dout(w_dff_A_aTsiJJrv4_0),.din(w_dff_A_C8Vla8lD6_0),.clk(gclk));
	jdff dff_A_aTsiJJrv4_0(.dout(w_dff_A_9mqD6HUG9_0),.din(w_dff_A_aTsiJJrv4_0),.clk(gclk));
	jdff dff_A_9mqD6HUG9_0(.dout(w_dff_A_Iw5anqG08_0),.din(w_dff_A_9mqD6HUG9_0),.clk(gclk));
	jdff dff_A_Iw5anqG08_0(.dout(w_dff_A_X4pmaQtB5_0),.din(w_dff_A_Iw5anqG08_0),.clk(gclk));
	jdff dff_A_X4pmaQtB5_0(.dout(w_dff_A_IPFAysBJ2_0),.din(w_dff_A_X4pmaQtB5_0),.clk(gclk));
	jdff dff_A_IPFAysBJ2_0(.dout(w_dff_A_KmQYMo2f8_0),.din(w_dff_A_IPFAysBJ2_0),.clk(gclk));
	jdff dff_A_KmQYMo2f8_0(.dout(w_dff_A_kSpLcaRg0_0),.din(w_dff_A_KmQYMo2f8_0),.clk(gclk));
	jdff dff_A_kSpLcaRg0_0(.dout(w_dff_A_gwo3cl2g1_0),.din(w_dff_A_kSpLcaRg0_0),.clk(gclk));
	jdff dff_A_gwo3cl2g1_0(.dout(w_dff_A_RNmscOtN0_0),.din(w_dff_A_gwo3cl2g1_0),.clk(gclk));
	jdff dff_A_RNmscOtN0_0(.dout(w_dff_A_e21daD3A5_0),.din(w_dff_A_RNmscOtN0_0),.clk(gclk));
	jdff dff_A_e21daD3A5_0(.dout(w_dff_A_FL5nlnuk2_0),.din(w_dff_A_e21daD3A5_0),.clk(gclk));
	jdff dff_A_FL5nlnuk2_0(.dout(w_dff_A_mF38GD9n2_0),.din(w_dff_A_FL5nlnuk2_0),.clk(gclk));
	jdff dff_A_mF38GD9n2_0(.dout(w_dff_A_MCCRLRZ42_0),.din(w_dff_A_mF38GD9n2_0),.clk(gclk));
	jdff dff_A_MCCRLRZ42_0(.dout(w_dff_A_Q6wfGJAf8_0),.din(w_dff_A_MCCRLRZ42_0),.clk(gclk));
	jdff dff_A_Q6wfGJAf8_0(.dout(w_dff_A_SDIwXHON3_0),.din(w_dff_A_Q6wfGJAf8_0),.clk(gclk));
	jdff dff_A_SDIwXHON3_0(.dout(w_dff_A_xzUct8pV1_0),.din(w_dff_A_SDIwXHON3_0),.clk(gclk));
	jdff dff_A_xzUct8pV1_0(.dout(w_dff_A_ZVXFcrWg6_0),.din(w_dff_A_xzUct8pV1_0),.clk(gclk));
	jdff dff_A_ZVXFcrWg6_0(.dout(w_dff_A_NjyRr0XE5_0),.din(w_dff_A_ZVXFcrWg6_0),.clk(gclk));
	jdff dff_A_NjyRr0XE5_0(.dout(w_dff_A_qi0spAow0_0),.din(w_dff_A_NjyRr0XE5_0),.clk(gclk));
	jdff dff_A_qi0spAow0_0(.dout(w_dff_A_IKJdRuNe5_0),.din(w_dff_A_qi0spAow0_0),.clk(gclk));
	jdff dff_A_IKJdRuNe5_0(.dout(w_dff_A_tyFnN7DZ0_0),.din(w_dff_A_IKJdRuNe5_0),.clk(gclk));
	jdff dff_A_tyFnN7DZ0_0(.dout(w_dff_A_qmyFeJwd2_0),.din(w_dff_A_tyFnN7DZ0_0),.clk(gclk));
	jdff dff_A_qmyFeJwd2_0(.dout(w_dff_A_pqhGVZIS8_0),.din(w_dff_A_qmyFeJwd2_0),.clk(gclk));
	jdff dff_A_pqhGVZIS8_0(.dout(w_dff_A_040MvXAb1_0),.din(w_dff_A_pqhGVZIS8_0),.clk(gclk));
	jdff dff_A_040MvXAb1_0(.dout(w_dff_A_DIwhYRBt6_0),.din(w_dff_A_040MvXAb1_0),.clk(gclk));
	jdff dff_A_DIwhYRBt6_0(.dout(w_dff_A_LtSWvQew5_0),.din(w_dff_A_DIwhYRBt6_0),.clk(gclk));
	jdff dff_A_LtSWvQew5_0(.dout(w_dff_A_4zHkLZ1s7_0),.din(w_dff_A_LtSWvQew5_0),.clk(gclk));
	jdff dff_A_4zHkLZ1s7_0(.dout(w_dff_A_urxoGnKd6_0),.din(w_dff_A_4zHkLZ1s7_0),.clk(gclk));
	jdff dff_A_urxoGnKd6_0(.dout(w_dff_A_f51uoYlA1_0),.din(w_dff_A_urxoGnKd6_0),.clk(gclk));
	jdff dff_A_f51uoYlA1_0(.dout(w_dff_A_gf7ecoOt2_0),.din(w_dff_A_f51uoYlA1_0),.clk(gclk));
	jdff dff_A_gf7ecoOt2_0(.dout(w_dff_A_hY9hUxCJ7_0),.din(w_dff_A_gf7ecoOt2_0),.clk(gclk));
	jdff dff_A_hY9hUxCJ7_0(.dout(f31),.din(w_dff_A_hY9hUxCJ7_0),.clk(gclk));
	jdff dff_A_Vbwd5rP60_2(.dout(w_dff_A_acguHRy91_0),.din(w_dff_A_Vbwd5rP60_2),.clk(gclk));
	jdff dff_A_acguHRy91_0(.dout(w_dff_A_eWBgmLM32_0),.din(w_dff_A_acguHRy91_0),.clk(gclk));
	jdff dff_A_eWBgmLM32_0(.dout(w_dff_A_JSH2BpPH9_0),.din(w_dff_A_eWBgmLM32_0),.clk(gclk));
	jdff dff_A_JSH2BpPH9_0(.dout(w_dff_A_HMEXUphm2_0),.din(w_dff_A_JSH2BpPH9_0),.clk(gclk));
	jdff dff_A_HMEXUphm2_0(.dout(w_dff_A_bcVfDLXc9_0),.din(w_dff_A_HMEXUphm2_0),.clk(gclk));
	jdff dff_A_bcVfDLXc9_0(.dout(w_dff_A_5WXv0ir40_0),.din(w_dff_A_bcVfDLXc9_0),.clk(gclk));
	jdff dff_A_5WXv0ir40_0(.dout(w_dff_A_qFOHSeqv5_0),.din(w_dff_A_5WXv0ir40_0),.clk(gclk));
	jdff dff_A_qFOHSeqv5_0(.dout(w_dff_A_ghqATLCH7_0),.din(w_dff_A_qFOHSeqv5_0),.clk(gclk));
	jdff dff_A_ghqATLCH7_0(.dout(w_dff_A_jtc57SmF2_0),.din(w_dff_A_ghqATLCH7_0),.clk(gclk));
	jdff dff_A_jtc57SmF2_0(.dout(w_dff_A_TxwVwgWQ2_0),.din(w_dff_A_jtc57SmF2_0),.clk(gclk));
	jdff dff_A_TxwVwgWQ2_0(.dout(w_dff_A_YJb9zqtS3_0),.din(w_dff_A_TxwVwgWQ2_0),.clk(gclk));
	jdff dff_A_YJb9zqtS3_0(.dout(w_dff_A_clURgq829_0),.din(w_dff_A_YJb9zqtS3_0),.clk(gclk));
	jdff dff_A_clURgq829_0(.dout(w_dff_A_B9nmkbPJ4_0),.din(w_dff_A_clURgq829_0),.clk(gclk));
	jdff dff_A_B9nmkbPJ4_0(.dout(w_dff_A_2k5Gk8BW7_0),.din(w_dff_A_B9nmkbPJ4_0),.clk(gclk));
	jdff dff_A_2k5Gk8BW7_0(.dout(w_dff_A_xhVLUZNi0_0),.din(w_dff_A_2k5Gk8BW7_0),.clk(gclk));
	jdff dff_A_xhVLUZNi0_0(.dout(w_dff_A_Eq0bb39p0_0),.din(w_dff_A_xhVLUZNi0_0),.clk(gclk));
	jdff dff_A_Eq0bb39p0_0(.dout(w_dff_A_lZWxKl9K6_0),.din(w_dff_A_Eq0bb39p0_0),.clk(gclk));
	jdff dff_A_lZWxKl9K6_0(.dout(w_dff_A_Bkm471TL8_0),.din(w_dff_A_lZWxKl9K6_0),.clk(gclk));
	jdff dff_A_Bkm471TL8_0(.dout(w_dff_A_mbXB2Dlq7_0),.din(w_dff_A_Bkm471TL8_0),.clk(gclk));
	jdff dff_A_mbXB2Dlq7_0(.dout(w_dff_A_8cDSucz92_0),.din(w_dff_A_mbXB2Dlq7_0),.clk(gclk));
	jdff dff_A_8cDSucz92_0(.dout(w_dff_A_zH2D31n48_0),.din(w_dff_A_8cDSucz92_0),.clk(gclk));
	jdff dff_A_zH2D31n48_0(.dout(w_dff_A_IllvKo8r0_0),.din(w_dff_A_zH2D31n48_0),.clk(gclk));
	jdff dff_A_IllvKo8r0_0(.dout(w_dff_A_F20VDSIx8_0),.din(w_dff_A_IllvKo8r0_0),.clk(gclk));
	jdff dff_A_F20VDSIx8_0(.dout(w_dff_A_Gy8blDOL3_0),.din(w_dff_A_F20VDSIx8_0),.clk(gclk));
	jdff dff_A_Gy8blDOL3_0(.dout(w_dff_A_R4YmRgQh0_0),.din(w_dff_A_Gy8blDOL3_0),.clk(gclk));
	jdff dff_A_R4YmRgQh0_0(.dout(w_dff_A_ZdZ8LIVF8_0),.din(w_dff_A_R4YmRgQh0_0),.clk(gclk));
	jdff dff_A_ZdZ8LIVF8_0(.dout(w_dff_A_lYwOT3XD6_0),.din(w_dff_A_ZdZ8LIVF8_0),.clk(gclk));
	jdff dff_A_lYwOT3XD6_0(.dout(w_dff_A_8NbSjTYQ0_0),.din(w_dff_A_lYwOT3XD6_0),.clk(gclk));
	jdff dff_A_8NbSjTYQ0_0(.dout(w_dff_A_8zrlZBVF5_0),.din(w_dff_A_8NbSjTYQ0_0),.clk(gclk));
	jdff dff_A_8zrlZBVF5_0(.dout(w_dff_A_f4lrLZTC3_0),.din(w_dff_A_8zrlZBVF5_0),.clk(gclk));
	jdff dff_A_f4lrLZTC3_0(.dout(w_dff_A_gDeO2G2C8_0),.din(w_dff_A_f4lrLZTC3_0),.clk(gclk));
	jdff dff_A_gDeO2G2C8_0(.dout(w_dff_A_FYGNwlxr1_0),.din(w_dff_A_gDeO2G2C8_0),.clk(gclk));
	jdff dff_A_FYGNwlxr1_0(.dout(w_dff_A_pfDFAsdz6_0),.din(w_dff_A_FYGNwlxr1_0),.clk(gclk));
	jdff dff_A_pfDFAsdz6_0(.dout(w_dff_A_zhWHKqVw6_0),.din(w_dff_A_pfDFAsdz6_0),.clk(gclk));
	jdff dff_A_zhWHKqVw6_0(.dout(w_dff_A_nxdqapsb6_0),.din(w_dff_A_zhWHKqVw6_0),.clk(gclk));
	jdff dff_A_nxdqapsb6_0(.dout(w_dff_A_9Ifi4L7F7_0),.din(w_dff_A_nxdqapsb6_0),.clk(gclk));
	jdff dff_A_9Ifi4L7F7_0(.dout(w_dff_A_e6CBJ4h21_0),.din(w_dff_A_9Ifi4L7F7_0),.clk(gclk));
	jdff dff_A_e6CBJ4h21_0(.dout(w_dff_A_PyiqqjOK3_0),.din(w_dff_A_e6CBJ4h21_0),.clk(gclk));
	jdff dff_A_PyiqqjOK3_0(.dout(w_dff_A_0aj8yugc3_0),.din(w_dff_A_PyiqqjOK3_0),.clk(gclk));
	jdff dff_A_0aj8yugc3_0(.dout(w_dff_A_Kbk3X0P69_0),.din(w_dff_A_0aj8yugc3_0),.clk(gclk));
	jdff dff_A_Kbk3X0P69_0(.dout(w_dff_A_ZFyWwRUf5_0),.din(w_dff_A_Kbk3X0P69_0),.clk(gclk));
	jdff dff_A_ZFyWwRUf5_0(.dout(w_dff_A_LjKvTvfa8_0),.din(w_dff_A_ZFyWwRUf5_0),.clk(gclk));
	jdff dff_A_LjKvTvfa8_0(.dout(w_dff_A_pKhsl2lB8_0),.din(w_dff_A_LjKvTvfa8_0),.clk(gclk));
	jdff dff_A_pKhsl2lB8_0(.dout(w_dff_A_mg62jM3S4_0),.din(w_dff_A_pKhsl2lB8_0),.clk(gclk));
	jdff dff_A_mg62jM3S4_0(.dout(w_dff_A_AAqXqg4v1_0),.din(w_dff_A_mg62jM3S4_0),.clk(gclk));
	jdff dff_A_AAqXqg4v1_0(.dout(w_dff_A_7y4CXdXA3_0),.din(w_dff_A_AAqXqg4v1_0),.clk(gclk));
	jdff dff_A_7y4CXdXA3_0(.dout(w_dff_A_VeG9PlFa4_0),.din(w_dff_A_7y4CXdXA3_0),.clk(gclk));
	jdff dff_A_VeG9PlFa4_0(.dout(w_dff_A_VHCXykxR6_0),.din(w_dff_A_VeG9PlFa4_0),.clk(gclk));
	jdff dff_A_VHCXykxR6_0(.dout(w_dff_A_r2eJsA1e5_0),.din(w_dff_A_VHCXykxR6_0),.clk(gclk));
	jdff dff_A_r2eJsA1e5_0(.dout(w_dff_A_lyLOCxks8_0),.din(w_dff_A_r2eJsA1e5_0),.clk(gclk));
	jdff dff_A_lyLOCxks8_0(.dout(w_dff_A_NKwRdkeW2_0),.din(w_dff_A_lyLOCxks8_0),.clk(gclk));
	jdff dff_A_NKwRdkeW2_0(.dout(w_dff_A_pb51qD7V7_0),.din(w_dff_A_NKwRdkeW2_0),.clk(gclk));
	jdff dff_A_pb51qD7V7_0(.dout(w_dff_A_Dh9H56nq3_0),.din(w_dff_A_pb51qD7V7_0),.clk(gclk));
	jdff dff_A_Dh9H56nq3_0(.dout(w_dff_A_e3fK55SL2_0),.din(w_dff_A_Dh9H56nq3_0),.clk(gclk));
	jdff dff_A_e3fK55SL2_0(.dout(w_dff_A_aSqW5MCq7_0),.din(w_dff_A_e3fK55SL2_0),.clk(gclk));
	jdff dff_A_aSqW5MCq7_0(.dout(w_dff_A_FIlD0ynx6_0),.din(w_dff_A_aSqW5MCq7_0),.clk(gclk));
	jdff dff_A_FIlD0ynx6_0(.dout(w_dff_A_1jOcEIC86_0),.din(w_dff_A_FIlD0ynx6_0),.clk(gclk));
	jdff dff_A_1jOcEIC86_0(.dout(w_dff_A_ErHwsI9U1_0),.din(w_dff_A_1jOcEIC86_0),.clk(gclk));
	jdff dff_A_ErHwsI9U1_0(.dout(w_dff_A_E0UGvoOz7_0),.din(w_dff_A_ErHwsI9U1_0),.clk(gclk));
	jdff dff_A_E0UGvoOz7_0(.dout(w_dff_A_b4I4O6NT4_0),.din(w_dff_A_E0UGvoOz7_0),.clk(gclk));
	jdff dff_A_b4I4O6NT4_0(.dout(w_dff_A_Qvjglidr8_0),.din(w_dff_A_b4I4O6NT4_0),.clk(gclk));
	jdff dff_A_Qvjglidr8_0(.dout(w_dff_A_7hICxZOP3_0),.din(w_dff_A_Qvjglidr8_0),.clk(gclk));
	jdff dff_A_7hICxZOP3_0(.dout(w_dff_A_b3ZCy4If2_0),.din(w_dff_A_7hICxZOP3_0),.clk(gclk));
	jdff dff_A_b3ZCy4If2_0(.dout(w_dff_A_iNXygzty4_0),.din(w_dff_A_b3ZCy4If2_0),.clk(gclk));
	jdff dff_A_iNXygzty4_0(.dout(w_dff_A_I6CWKPnt2_0),.din(w_dff_A_iNXygzty4_0),.clk(gclk));
	jdff dff_A_I6CWKPnt2_0(.dout(w_dff_A_Ij6AZunJ7_0),.din(w_dff_A_I6CWKPnt2_0),.clk(gclk));
	jdff dff_A_Ij6AZunJ7_0(.dout(w_dff_A_J8aEbPPM5_0),.din(w_dff_A_Ij6AZunJ7_0),.clk(gclk));
	jdff dff_A_J8aEbPPM5_0(.dout(w_dff_A_8LEMS8j92_0),.din(w_dff_A_J8aEbPPM5_0),.clk(gclk));
	jdff dff_A_8LEMS8j92_0(.dout(w_dff_A_zuTy6rDg4_0),.din(w_dff_A_8LEMS8j92_0),.clk(gclk));
	jdff dff_A_zuTy6rDg4_0(.dout(w_dff_A_lMoM9Gie5_0),.din(w_dff_A_zuTy6rDg4_0),.clk(gclk));
	jdff dff_A_lMoM9Gie5_0(.dout(w_dff_A_63TjIIhN6_0),.din(w_dff_A_lMoM9Gie5_0),.clk(gclk));
	jdff dff_A_63TjIIhN6_0(.dout(w_dff_A_9U3JIBlW5_0),.din(w_dff_A_63TjIIhN6_0),.clk(gclk));
	jdff dff_A_9U3JIBlW5_0(.dout(w_dff_A_dOXYVYLk3_0),.din(w_dff_A_9U3JIBlW5_0),.clk(gclk));
	jdff dff_A_dOXYVYLk3_0(.dout(w_dff_A_iQkxLnZO6_0),.din(w_dff_A_dOXYVYLk3_0),.clk(gclk));
	jdff dff_A_iQkxLnZO6_0(.dout(w_dff_A_e9uXjCFR8_0),.din(w_dff_A_iQkxLnZO6_0),.clk(gclk));
	jdff dff_A_e9uXjCFR8_0(.dout(w_dff_A_D1x8SWGG8_0),.din(w_dff_A_e9uXjCFR8_0),.clk(gclk));
	jdff dff_A_D1x8SWGG8_0(.dout(w_dff_A_EN0b0VM04_0),.din(w_dff_A_D1x8SWGG8_0),.clk(gclk));
	jdff dff_A_EN0b0VM04_0(.dout(w_dff_A_hOUe51KZ0_0),.din(w_dff_A_EN0b0VM04_0),.clk(gclk));
	jdff dff_A_hOUe51KZ0_0(.dout(w_dff_A_RASIn91O7_0),.din(w_dff_A_hOUe51KZ0_0),.clk(gclk));
	jdff dff_A_RASIn91O7_0(.dout(w_dff_A_C5xiiUX07_0),.din(w_dff_A_RASIn91O7_0),.clk(gclk));
	jdff dff_A_C5xiiUX07_0(.dout(w_dff_A_5ocXhG7j9_0),.din(w_dff_A_C5xiiUX07_0),.clk(gclk));
	jdff dff_A_5ocXhG7j9_0(.dout(w_dff_A_lrIdjV6O5_0),.din(w_dff_A_5ocXhG7j9_0),.clk(gclk));
	jdff dff_A_lrIdjV6O5_0(.dout(w_dff_A_v27JInPy5_0),.din(w_dff_A_lrIdjV6O5_0),.clk(gclk));
	jdff dff_A_v27JInPy5_0(.dout(w_dff_A_JwrjPW391_0),.din(w_dff_A_v27JInPy5_0),.clk(gclk));
	jdff dff_A_JwrjPW391_0(.dout(w_dff_A_b3eubL1g9_0),.din(w_dff_A_JwrjPW391_0),.clk(gclk));
	jdff dff_A_b3eubL1g9_0(.dout(w_dff_A_SVuujN5B0_0),.din(w_dff_A_b3eubL1g9_0),.clk(gclk));
	jdff dff_A_SVuujN5B0_0(.dout(w_dff_A_clOeg2UJ0_0),.din(w_dff_A_SVuujN5B0_0),.clk(gclk));
	jdff dff_A_clOeg2UJ0_0(.dout(w_dff_A_IQkFWOGN0_0),.din(w_dff_A_clOeg2UJ0_0),.clk(gclk));
	jdff dff_A_IQkFWOGN0_0(.dout(w_dff_A_VZcJ0Hsj1_0),.din(w_dff_A_IQkFWOGN0_0),.clk(gclk));
	jdff dff_A_VZcJ0Hsj1_0(.dout(w_dff_A_371ihWaD5_0),.din(w_dff_A_VZcJ0Hsj1_0),.clk(gclk));
	jdff dff_A_371ihWaD5_0(.dout(w_dff_A_l6xAvpDk0_0),.din(w_dff_A_371ihWaD5_0),.clk(gclk));
	jdff dff_A_l6xAvpDk0_0(.dout(w_dff_A_YGN7U03v6_0),.din(w_dff_A_l6xAvpDk0_0),.clk(gclk));
	jdff dff_A_YGN7U03v6_0(.dout(w_dff_A_PR52G4kM5_0),.din(w_dff_A_YGN7U03v6_0),.clk(gclk));
	jdff dff_A_PR52G4kM5_0(.dout(w_dff_A_xGcvzYlW6_0),.din(w_dff_A_PR52G4kM5_0),.clk(gclk));
	jdff dff_A_xGcvzYlW6_0(.dout(f32),.din(w_dff_A_xGcvzYlW6_0),.clk(gclk));
	jdff dff_A_AA7idxgZ2_2(.dout(w_dff_A_IXmzJoD52_0),.din(w_dff_A_AA7idxgZ2_2),.clk(gclk));
	jdff dff_A_IXmzJoD52_0(.dout(w_dff_A_SUiDWMsI0_0),.din(w_dff_A_IXmzJoD52_0),.clk(gclk));
	jdff dff_A_SUiDWMsI0_0(.dout(w_dff_A_8ttcsU1w2_0),.din(w_dff_A_SUiDWMsI0_0),.clk(gclk));
	jdff dff_A_8ttcsU1w2_0(.dout(w_dff_A_BtjTE1X13_0),.din(w_dff_A_8ttcsU1w2_0),.clk(gclk));
	jdff dff_A_BtjTE1X13_0(.dout(w_dff_A_iIJyQgKl8_0),.din(w_dff_A_BtjTE1X13_0),.clk(gclk));
	jdff dff_A_iIJyQgKl8_0(.dout(w_dff_A_4BgOiuQ80_0),.din(w_dff_A_iIJyQgKl8_0),.clk(gclk));
	jdff dff_A_4BgOiuQ80_0(.dout(w_dff_A_ar2v2KAu2_0),.din(w_dff_A_4BgOiuQ80_0),.clk(gclk));
	jdff dff_A_ar2v2KAu2_0(.dout(w_dff_A_OI9oBg3b5_0),.din(w_dff_A_ar2v2KAu2_0),.clk(gclk));
	jdff dff_A_OI9oBg3b5_0(.dout(w_dff_A_Fvd5Iqva9_0),.din(w_dff_A_OI9oBg3b5_0),.clk(gclk));
	jdff dff_A_Fvd5Iqva9_0(.dout(w_dff_A_e4DhpLi45_0),.din(w_dff_A_Fvd5Iqva9_0),.clk(gclk));
	jdff dff_A_e4DhpLi45_0(.dout(w_dff_A_AdpjdJE36_0),.din(w_dff_A_e4DhpLi45_0),.clk(gclk));
	jdff dff_A_AdpjdJE36_0(.dout(w_dff_A_uAxjzFmT5_0),.din(w_dff_A_AdpjdJE36_0),.clk(gclk));
	jdff dff_A_uAxjzFmT5_0(.dout(w_dff_A_oiCFDegG8_0),.din(w_dff_A_uAxjzFmT5_0),.clk(gclk));
	jdff dff_A_oiCFDegG8_0(.dout(w_dff_A_LZFLbM197_0),.din(w_dff_A_oiCFDegG8_0),.clk(gclk));
	jdff dff_A_LZFLbM197_0(.dout(w_dff_A_DDdq2hdP1_0),.din(w_dff_A_LZFLbM197_0),.clk(gclk));
	jdff dff_A_DDdq2hdP1_0(.dout(w_dff_A_4swA2f0R9_0),.din(w_dff_A_DDdq2hdP1_0),.clk(gclk));
	jdff dff_A_4swA2f0R9_0(.dout(w_dff_A_pD2JoyfP9_0),.din(w_dff_A_4swA2f0R9_0),.clk(gclk));
	jdff dff_A_pD2JoyfP9_0(.dout(w_dff_A_JkLgDBAh7_0),.din(w_dff_A_pD2JoyfP9_0),.clk(gclk));
	jdff dff_A_JkLgDBAh7_0(.dout(w_dff_A_6atLCMun9_0),.din(w_dff_A_JkLgDBAh7_0),.clk(gclk));
	jdff dff_A_6atLCMun9_0(.dout(w_dff_A_FzUfkCb47_0),.din(w_dff_A_6atLCMun9_0),.clk(gclk));
	jdff dff_A_FzUfkCb47_0(.dout(w_dff_A_s28azhb96_0),.din(w_dff_A_FzUfkCb47_0),.clk(gclk));
	jdff dff_A_s28azhb96_0(.dout(w_dff_A_BKabnSNy7_0),.din(w_dff_A_s28azhb96_0),.clk(gclk));
	jdff dff_A_BKabnSNy7_0(.dout(w_dff_A_abzSJv9j8_0),.din(w_dff_A_BKabnSNy7_0),.clk(gclk));
	jdff dff_A_abzSJv9j8_0(.dout(w_dff_A_moYeier78_0),.din(w_dff_A_abzSJv9j8_0),.clk(gclk));
	jdff dff_A_moYeier78_0(.dout(w_dff_A_3rJjjKxc2_0),.din(w_dff_A_moYeier78_0),.clk(gclk));
	jdff dff_A_3rJjjKxc2_0(.dout(w_dff_A_nXxWogiK6_0),.din(w_dff_A_3rJjjKxc2_0),.clk(gclk));
	jdff dff_A_nXxWogiK6_0(.dout(w_dff_A_pYxWmkhq9_0),.din(w_dff_A_nXxWogiK6_0),.clk(gclk));
	jdff dff_A_pYxWmkhq9_0(.dout(w_dff_A_9I0NvBXT3_0),.din(w_dff_A_pYxWmkhq9_0),.clk(gclk));
	jdff dff_A_9I0NvBXT3_0(.dout(w_dff_A_BSRWfDZO2_0),.din(w_dff_A_9I0NvBXT3_0),.clk(gclk));
	jdff dff_A_BSRWfDZO2_0(.dout(w_dff_A_Rqpj8eeM9_0),.din(w_dff_A_BSRWfDZO2_0),.clk(gclk));
	jdff dff_A_Rqpj8eeM9_0(.dout(w_dff_A_D1MWBfai8_0),.din(w_dff_A_Rqpj8eeM9_0),.clk(gclk));
	jdff dff_A_D1MWBfai8_0(.dout(w_dff_A_ylUcUOKr0_0),.din(w_dff_A_D1MWBfai8_0),.clk(gclk));
	jdff dff_A_ylUcUOKr0_0(.dout(w_dff_A_7HtJzcqB7_0),.din(w_dff_A_ylUcUOKr0_0),.clk(gclk));
	jdff dff_A_7HtJzcqB7_0(.dout(w_dff_A_RGHXKlFs4_0),.din(w_dff_A_7HtJzcqB7_0),.clk(gclk));
	jdff dff_A_RGHXKlFs4_0(.dout(w_dff_A_h7P5aI7x7_0),.din(w_dff_A_RGHXKlFs4_0),.clk(gclk));
	jdff dff_A_h7P5aI7x7_0(.dout(w_dff_A_smmsHfTa6_0),.din(w_dff_A_h7P5aI7x7_0),.clk(gclk));
	jdff dff_A_smmsHfTa6_0(.dout(w_dff_A_EyUiVyjx5_0),.din(w_dff_A_smmsHfTa6_0),.clk(gclk));
	jdff dff_A_EyUiVyjx5_0(.dout(w_dff_A_e4bPu2DX3_0),.din(w_dff_A_EyUiVyjx5_0),.clk(gclk));
	jdff dff_A_e4bPu2DX3_0(.dout(w_dff_A_3sr77xXo2_0),.din(w_dff_A_e4bPu2DX3_0),.clk(gclk));
	jdff dff_A_3sr77xXo2_0(.dout(w_dff_A_DDofauw05_0),.din(w_dff_A_3sr77xXo2_0),.clk(gclk));
	jdff dff_A_DDofauw05_0(.dout(w_dff_A_uB5FBS4F3_0),.din(w_dff_A_DDofauw05_0),.clk(gclk));
	jdff dff_A_uB5FBS4F3_0(.dout(w_dff_A_IiNkcaVJ4_0),.din(w_dff_A_uB5FBS4F3_0),.clk(gclk));
	jdff dff_A_IiNkcaVJ4_0(.dout(w_dff_A_BjqJnB1N6_0),.din(w_dff_A_IiNkcaVJ4_0),.clk(gclk));
	jdff dff_A_BjqJnB1N6_0(.dout(w_dff_A_RHqTVs6M4_0),.din(w_dff_A_BjqJnB1N6_0),.clk(gclk));
	jdff dff_A_RHqTVs6M4_0(.dout(w_dff_A_ziibFKak8_0),.din(w_dff_A_RHqTVs6M4_0),.clk(gclk));
	jdff dff_A_ziibFKak8_0(.dout(w_dff_A_obMBmyXc1_0),.din(w_dff_A_ziibFKak8_0),.clk(gclk));
	jdff dff_A_obMBmyXc1_0(.dout(w_dff_A_WxsrymzD2_0),.din(w_dff_A_obMBmyXc1_0),.clk(gclk));
	jdff dff_A_WxsrymzD2_0(.dout(w_dff_A_H1viYh4t5_0),.din(w_dff_A_WxsrymzD2_0),.clk(gclk));
	jdff dff_A_H1viYh4t5_0(.dout(w_dff_A_OfYT7qSR0_0),.din(w_dff_A_H1viYh4t5_0),.clk(gclk));
	jdff dff_A_OfYT7qSR0_0(.dout(w_dff_A_0DiFCaFh0_0),.din(w_dff_A_OfYT7qSR0_0),.clk(gclk));
	jdff dff_A_0DiFCaFh0_0(.dout(w_dff_A_f98SiEhU9_0),.din(w_dff_A_0DiFCaFh0_0),.clk(gclk));
	jdff dff_A_f98SiEhU9_0(.dout(w_dff_A_iomll8mg2_0),.din(w_dff_A_f98SiEhU9_0),.clk(gclk));
	jdff dff_A_iomll8mg2_0(.dout(w_dff_A_pd95cPaR6_0),.din(w_dff_A_iomll8mg2_0),.clk(gclk));
	jdff dff_A_pd95cPaR6_0(.dout(w_dff_A_NAWgwRXy1_0),.din(w_dff_A_pd95cPaR6_0),.clk(gclk));
	jdff dff_A_NAWgwRXy1_0(.dout(w_dff_A_zS2cQVBn4_0),.din(w_dff_A_NAWgwRXy1_0),.clk(gclk));
	jdff dff_A_zS2cQVBn4_0(.dout(w_dff_A_8LnUQHd07_0),.din(w_dff_A_zS2cQVBn4_0),.clk(gclk));
	jdff dff_A_8LnUQHd07_0(.dout(w_dff_A_J6dmwfBt1_0),.din(w_dff_A_8LnUQHd07_0),.clk(gclk));
	jdff dff_A_J6dmwfBt1_0(.dout(w_dff_A_f5mH1I341_0),.din(w_dff_A_J6dmwfBt1_0),.clk(gclk));
	jdff dff_A_f5mH1I341_0(.dout(w_dff_A_SnITCqxm0_0),.din(w_dff_A_f5mH1I341_0),.clk(gclk));
	jdff dff_A_SnITCqxm0_0(.dout(w_dff_A_1wiy9psF6_0),.din(w_dff_A_SnITCqxm0_0),.clk(gclk));
	jdff dff_A_1wiy9psF6_0(.dout(w_dff_A_b7nmvzCl5_0),.din(w_dff_A_1wiy9psF6_0),.clk(gclk));
	jdff dff_A_b7nmvzCl5_0(.dout(w_dff_A_B24VU6qr8_0),.din(w_dff_A_b7nmvzCl5_0),.clk(gclk));
	jdff dff_A_B24VU6qr8_0(.dout(w_dff_A_BKMY13M98_0),.din(w_dff_A_B24VU6qr8_0),.clk(gclk));
	jdff dff_A_BKMY13M98_0(.dout(w_dff_A_bGXrTSQm1_0),.din(w_dff_A_BKMY13M98_0),.clk(gclk));
	jdff dff_A_bGXrTSQm1_0(.dout(w_dff_A_0gfJ2qsd5_0),.din(w_dff_A_bGXrTSQm1_0),.clk(gclk));
	jdff dff_A_0gfJ2qsd5_0(.dout(w_dff_A_qwMrHx5C7_0),.din(w_dff_A_0gfJ2qsd5_0),.clk(gclk));
	jdff dff_A_qwMrHx5C7_0(.dout(w_dff_A_X7FPCX4q5_0),.din(w_dff_A_qwMrHx5C7_0),.clk(gclk));
	jdff dff_A_X7FPCX4q5_0(.dout(w_dff_A_o07PCTzF8_0),.din(w_dff_A_X7FPCX4q5_0),.clk(gclk));
	jdff dff_A_o07PCTzF8_0(.dout(w_dff_A_Yk0FZKU76_0),.din(w_dff_A_o07PCTzF8_0),.clk(gclk));
	jdff dff_A_Yk0FZKU76_0(.dout(w_dff_A_FlwsofEx2_0),.din(w_dff_A_Yk0FZKU76_0),.clk(gclk));
	jdff dff_A_FlwsofEx2_0(.dout(w_dff_A_OnR1Doqj1_0),.din(w_dff_A_FlwsofEx2_0),.clk(gclk));
	jdff dff_A_OnR1Doqj1_0(.dout(w_dff_A_2he1DkqY1_0),.din(w_dff_A_OnR1Doqj1_0),.clk(gclk));
	jdff dff_A_2he1DkqY1_0(.dout(w_dff_A_F0QLvxFp8_0),.din(w_dff_A_2he1DkqY1_0),.clk(gclk));
	jdff dff_A_F0QLvxFp8_0(.dout(w_dff_A_doVAtjvv4_0),.din(w_dff_A_F0QLvxFp8_0),.clk(gclk));
	jdff dff_A_doVAtjvv4_0(.dout(w_dff_A_YNwZFz0b5_0),.din(w_dff_A_doVAtjvv4_0),.clk(gclk));
	jdff dff_A_YNwZFz0b5_0(.dout(w_dff_A_iiS1uhtG2_0),.din(w_dff_A_YNwZFz0b5_0),.clk(gclk));
	jdff dff_A_iiS1uhtG2_0(.dout(w_dff_A_mSnl7QXm0_0),.din(w_dff_A_iiS1uhtG2_0),.clk(gclk));
	jdff dff_A_mSnl7QXm0_0(.dout(w_dff_A_qtMP3eTI2_0),.din(w_dff_A_mSnl7QXm0_0),.clk(gclk));
	jdff dff_A_qtMP3eTI2_0(.dout(w_dff_A_8gSwC1OM6_0),.din(w_dff_A_qtMP3eTI2_0),.clk(gclk));
	jdff dff_A_8gSwC1OM6_0(.dout(w_dff_A_4vJTNDWE6_0),.din(w_dff_A_8gSwC1OM6_0),.clk(gclk));
	jdff dff_A_4vJTNDWE6_0(.dout(w_dff_A_BXTRr1C68_0),.din(w_dff_A_4vJTNDWE6_0),.clk(gclk));
	jdff dff_A_BXTRr1C68_0(.dout(w_dff_A_byH2M9Em8_0),.din(w_dff_A_BXTRr1C68_0),.clk(gclk));
	jdff dff_A_byH2M9Em8_0(.dout(w_dff_A_DCC8dUoA2_0),.din(w_dff_A_byH2M9Em8_0),.clk(gclk));
	jdff dff_A_DCC8dUoA2_0(.dout(w_dff_A_mW4mUuKi0_0),.din(w_dff_A_DCC8dUoA2_0),.clk(gclk));
	jdff dff_A_mW4mUuKi0_0(.dout(w_dff_A_RG18yxmP6_0),.din(w_dff_A_mW4mUuKi0_0),.clk(gclk));
	jdff dff_A_RG18yxmP6_0(.dout(w_dff_A_YrIiJjdx1_0),.din(w_dff_A_RG18yxmP6_0),.clk(gclk));
	jdff dff_A_YrIiJjdx1_0(.dout(w_dff_A_7RQJdfYD5_0),.din(w_dff_A_YrIiJjdx1_0),.clk(gclk));
	jdff dff_A_7RQJdfYD5_0(.dout(w_dff_A_rELg6bc66_0),.din(w_dff_A_7RQJdfYD5_0),.clk(gclk));
	jdff dff_A_rELg6bc66_0(.dout(w_dff_A_GRm0XSQP3_0),.din(w_dff_A_rELg6bc66_0),.clk(gclk));
	jdff dff_A_GRm0XSQP3_0(.dout(w_dff_A_ecCi7hRr4_0),.din(w_dff_A_GRm0XSQP3_0),.clk(gclk));
	jdff dff_A_ecCi7hRr4_0(.dout(w_dff_A_LXFfsDD52_0),.din(w_dff_A_ecCi7hRr4_0),.clk(gclk));
	jdff dff_A_LXFfsDD52_0(.dout(w_dff_A_VcVhUY0c1_0),.din(w_dff_A_LXFfsDD52_0),.clk(gclk));
	jdff dff_A_VcVhUY0c1_0(.dout(w_dff_A_rOMkywIm4_0),.din(w_dff_A_VcVhUY0c1_0),.clk(gclk));
	jdff dff_A_rOMkywIm4_0(.dout(f33),.din(w_dff_A_rOMkywIm4_0),.clk(gclk));
	jdff dff_A_RzzGmYzn3_2(.dout(w_dff_A_dBfSA6ub2_0),.din(w_dff_A_RzzGmYzn3_2),.clk(gclk));
	jdff dff_A_dBfSA6ub2_0(.dout(w_dff_A_XVUpZ1zt4_0),.din(w_dff_A_dBfSA6ub2_0),.clk(gclk));
	jdff dff_A_XVUpZ1zt4_0(.dout(w_dff_A_ujn4DM6Y2_0),.din(w_dff_A_XVUpZ1zt4_0),.clk(gclk));
	jdff dff_A_ujn4DM6Y2_0(.dout(w_dff_A_l1mlQqA58_0),.din(w_dff_A_ujn4DM6Y2_0),.clk(gclk));
	jdff dff_A_l1mlQqA58_0(.dout(w_dff_A_muVwVuO97_0),.din(w_dff_A_l1mlQqA58_0),.clk(gclk));
	jdff dff_A_muVwVuO97_0(.dout(w_dff_A_3CqjXeza9_0),.din(w_dff_A_muVwVuO97_0),.clk(gclk));
	jdff dff_A_3CqjXeza9_0(.dout(w_dff_A_qSonBavG7_0),.din(w_dff_A_3CqjXeza9_0),.clk(gclk));
	jdff dff_A_qSonBavG7_0(.dout(w_dff_A_jMbSoduW0_0),.din(w_dff_A_qSonBavG7_0),.clk(gclk));
	jdff dff_A_jMbSoduW0_0(.dout(w_dff_A_TqndA2fP0_0),.din(w_dff_A_jMbSoduW0_0),.clk(gclk));
	jdff dff_A_TqndA2fP0_0(.dout(w_dff_A_5wxTBUxl4_0),.din(w_dff_A_TqndA2fP0_0),.clk(gclk));
	jdff dff_A_5wxTBUxl4_0(.dout(w_dff_A_S6H1fwlD7_0),.din(w_dff_A_5wxTBUxl4_0),.clk(gclk));
	jdff dff_A_S6H1fwlD7_0(.dout(w_dff_A_K6qO0xqR0_0),.din(w_dff_A_S6H1fwlD7_0),.clk(gclk));
	jdff dff_A_K6qO0xqR0_0(.dout(w_dff_A_im83zL383_0),.din(w_dff_A_K6qO0xqR0_0),.clk(gclk));
	jdff dff_A_im83zL383_0(.dout(w_dff_A_9DOqdkgc0_0),.din(w_dff_A_im83zL383_0),.clk(gclk));
	jdff dff_A_9DOqdkgc0_0(.dout(w_dff_A_WJCw94Aj0_0),.din(w_dff_A_9DOqdkgc0_0),.clk(gclk));
	jdff dff_A_WJCw94Aj0_0(.dout(w_dff_A_KWN1dpvq2_0),.din(w_dff_A_WJCw94Aj0_0),.clk(gclk));
	jdff dff_A_KWN1dpvq2_0(.dout(w_dff_A_kxCmcfCc4_0),.din(w_dff_A_KWN1dpvq2_0),.clk(gclk));
	jdff dff_A_kxCmcfCc4_0(.dout(w_dff_A_lHHp85zP6_0),.din(w_dff_A_kxCmcfCc4_0),.clk(gclk));
	jdff dff_A_lHHp85zP6_0(.dout(w_dff_A_BYrGi2QE3_0),.din(w_dff_A_lHHp85zP6_0),.clk(gclk));
	jdff dff_A_BYrGi2QE3_0(.dout(w_dff_A_zk1BHnw74_0),.din(w_dff_A_BYrGi2QE3_0),.clk(gclk));
	jdff dff_A_zk1BHnw74_0(.dout(w_dff_A_64r3MPyM1_0),.din(w_dff_A_zk1BHnw74_0),.clk(gclk));
	jdff dff_A_64r3MPyM1_0(.dout(w_dff_A_m3JAd3kv5_0),.din(w_dff_A_64r3MPyM1_0),.clk(gclk));
	jdff dff_A_m3JAd3kv5_0(.dout(w_dff_A_0coZ5S9K5_0),.din(w_dff_A_m3JAd3kv5_0),.clk(gclk));
	jdff dff_A_0coZ5S9K5_0(.dout(w_dff_A_QB0Ew6V78_0),.din(w_dff_A_0coZ5S9K5_0),.clk(gclk));
	jdff dff_A_QB0Ew6V78_0(.dout(w_dff_A_5iNSLTx45_0),.din(w_dff_A_QB0Ew6V78_0),.clk(gclk));
	jdff dff_A_5iNSLTx45_0(.dout(w_dff_A_bYHfNVbu0_0),.din(w_dff_A_5iNSLTx45_0),.clk(gclk));
	jdff dff_A_bYHfNVbu0_0(.dout(w_dff_A_iJkKEHDC9_0),.din(w_dff_A_bYHfNVbu0_0),.clk(gclk));
	jdff dff_A_iJkKEHDC9_0(.dout(w_dff_A_pCb7MVQY4_0),.din(w_dff_A_iJkKEHDC9_0),.clk(gclk));
	jdff dff_A_pCb7MVQY4_0(.dout(w_dff_A_0A1tRegP0_0),.din(w_dff_A_pCb7MVQY4_0),.clk(gclk));
	jdff dff_A_0A1tRegP0_0(.dout(w_dff_A_7IqpVO0B0_0),.din(w_dff_A_0A1tRegP0_0),.clk(gclk));
	jdff dff_A_7IqpVO0B0_0(.dout(w_dff_A_AW8ITODf7_0),.din(w_dff_A_7IqpVO0B0_0),.clk(gclk));
	jdff dff_A_AW8ITODf7_0(.dout(w_dff_A_fqASo0au1_0),.din(w_dff_A_AW8ITODf7_0),.clk(gclk));
	jdff dff_A_fqASo0au1_0(.dout(w_dff_A_me17I2Uh7_0),.din(w_dff_A_fqASo0au1_0),.clk(gclk));
	jdff dff_A_me17I2Uh7_0(.dout(w_dff_A_SHmfCT5H6_0),.din(w_dff_A_me17I2Uh7_0),.clk(gclk));
	jdff dff_A_SHmfCT5H6_0(.dout(w_dff_A_XnnE3lZb4_0),.din(w_dff_A_SHmfCT5H6_0),.clk(gclk));
	jdff dff_A_XnnE3lZb4_0(.dout(w_dff_A_CAYP4COO3_0),.din(w_dff_A_XnnE3lZb4_0),.clk(gclk));
	jdff dff_A_CAYP4COO3_0(.dout(w_dff_A_vT7dtpOs6_0),.din(w_dff_A_CAYP4COO3_0),.clk(gclk));
	jdff dff_A_vT7dtpOs6_0(.dout(w_dff_A_0CCWzmD37_0),.din(w_dff_A_vT7dtpOs6_0),.clk(gclk));
	jdff dff_A_0CCWzmD37_0(.dout(w_dff_A_rtpnFsbC4_0),.din(w_dff_A_0CCWzmD37_0),.clk(gclk));
	jdff dff_A_rtpnFsbC4_0(.dout(w_dff_A_CNta6gfV7_0),.din(w_dff_A_rtpnFsbC4_0),.clk(gclk));
	jdff dff_A_CNta6gfV7_0(.dout(w_dff_A_h1jEWET94_0),.din(w_dff_A_CNta6gfV7_0),.clk(gclk));
	jdff dff_A_h1jEWET94_0(.dout(w_dff_A_PRPja86B6_0),.din(w_dff_A_h1jEWET94_0),.clk(gclk));
	jdff dff_A_PRPja86B6_0(.dout(w_dff_A_XmzsLt3A5_0),.din(w_dff_A_PRPja86B6_0),.clk(gclk));
	jdff dff_A_XmzsLt3A5_0(.dout(w_dff_A_4s28Zs3r3_0),.din(w_dff_A_XmzsLt3A5_0),.clk(gclk));
	jdff dff_A_4s28Zs3r3_0(.dout(w_dff_A_6DZhO1yC4_0),.din(w_dff_A_4s28Zs3r3_0),.clk(gclk));
	jdff dff_A_6DZhO1yC4_0(.dout(w_dff_A_J8SHmDK24_0),.din(w_dff_A_6DZhO1yC4_0),.clk(gclk));
	jdff dff_A_J8SHmDK24_0(.dout(w_dff_A_Kfi0iQGv1_0),.din(w_dff_A_J8SHmDK24_0),.clk(gclk));
	jdff dff_A_Kfi0iQGv1_0(.dout(w_dff_A_lRlRaB3M2_0),.din(w_dff_A_Kfi0iQGv1_0),.clk(gclk));
	jdff dff_A_lRlRaB3M2_0(.dout(w_dff_A_Duc2nt1T2_0),.din(w_dff_A_lRlRaB3M2_0),.clk(gclk));
	jdff dff_A_Duc2nt1T2_0(.dout(w_dff_A_tQeUDxrn0_0),.din(w_dff_A_Duc2nt1T2_0),.clk(gclk));
	jdff dff_A_tQeUDxrn0_0(.dout(w_dff_A_uXAl6YYf0_0),.din(w_dff_A_tQeUDxrn0_0),.clk(gclk));
	jdff dff_A_uXAl6YYf0_0(.dout(w_dff_A_F9UTqTjf7_0),.din(w_dff_A_uXAl6YYf0_0),.clk(gclk));
	jdff dff_A_F9UTqTjf7_0(.dout(w_dff_A_ktsnwwmm6_0),.din(w_dff_A_F9UTqTjf7_0),.clk(gclk));
	jdff dff_A_ktsnwwmm6_0(.dout(w_dff_A_yTS93qct5_0),.din(w_dff_A_ktsnwwmm6_0),.clk(gclk));
	jdff dff_A_yTS93qct5_0(.dout(w_dff_A_EkQB7zjQ9_0),.din(w_dff_A_yTS93qct5_0),.clk(gclk));
	jdff dff_A_EkQB7zjQ9_0(.dout(w_dff_A_tQ0JowUq0_0),.din(w_dff_A_EkQB7zjQ9_0),.clk(gclk));
	jdff dff_A_tQ0JowUq0_0(.dout(w_dff_A_PVT7U1Ql3_0),.din(w_dff_A_tQ0JowUq0_0),.clk(gclk));
	jdff dff_A_PVT7U1Ql3_0(.dout(w_dff_A_sSql4X0H4_0),.din(w_dff_A_PVT7U1Ql3_0),.clk(gclk));
	jdff dff_A_sSql4X0H4_0(.dout(w_dff_A_Umyqc3P18_0),.din(w_dff_A_sSql4X0H4_0),.clk(gclk));
	jdff dff_A_Umyqc3P18_0(.dout(w_dff_A_cbI1DzSd1_0),.din(w_dff_A_Umyqc3P18_0),.clk(gclk));
	jdff dff_A_cbI1DzSd1_0(.dout(w_dff_A_caKcpMok2_0),.din(w_dff_A_cbI1DzSd1_0),.clk(gclk));
	jdff dff_A_caKcpMok2_0(.dout(w_dff_A_LUG9mbHN3_0),.din(w_dff_A_caKcpMok2_0),.clk(gclk));
	jdff dff_A_LUG9mbHN3_0(.dout(w_dff_A_TxDL49bF2_0),.din(w_dff_A_LUG9mbHN3_0),.clk(gclk));
	jdff dff_A_TxDL49bF2_0(.dout(w_dff_A_ArgMUspD6_0),.din(w_dff_A_TxDL49bF2_0),.clk(gclk));
	jdff dff_A_ArgMUspD6_0(.dout(w_dff_A_d8aAiL6X2_0),.din(w_dff_A_ArgMUspD6_0),.clk(gclk));
	jdff dff_A_d8aAiL6X2_0(.dout(w_dff_A_PSF79s9m0_0),.din(w_dff_A_d8aAiL6X2_0),.clk(gclk));
	jdff dff_A_PSF79s9m0_0(.dout(w_dff_A_jPrwRqPh1_0),.din(w_dff_A_PSF79s9m0_0),.clk(gclk));
	jdff dff_A_jPrwRqPh1_0(.dout(w_dff_A_yJ53mRLy5_0),.din(w_dff_A_jPrwRqPh1_0),.clk(gclk));
	jdff dff_A_yJ53mRLy5_0(.dout(w_dff_A_14G7cpxf1_0),.din(w_dff_A_yJ53mRLy5_0),.clk(gclk));
	jdff dff_A_14G7cpxf1_0(.dout(w_dff_A_SD4vpAb10_0),.din(w_dff_A_14G7cpxf1_0),.clk(gclk));
	jdff dff_A_SD4vpAb10_0(.dout(w_dff_A_PfqZXFCM0_0),.din(w_dff_A_SD4vpAb10_0),.clk(gclk));
	jdff dff_A_PfqZXFCM0_0(.dout(w_dff_A_aIEP0Nlq5_0),.din(w_dff_A_PfqZXFCM0_0),.clk(gclk));
	jdff dff_A_aIEP0Nlq5_0(.dout(w_dff_A_Jyw4jyqW7_0),.din(w_dff_A_aIEP0Nlq5_0),.clk(gclk));
	jdff dff_A_Jyw4jyqW7_0(.dout(w_dff_A_SCuselYG2_0),.din(w_dff_A_Jyw4jyqW7_0),.clk(gclk));
	jdff dff_A_SCuselYG2_0(.dout(w_dff_A_7Z92uT2d2_0),.din(w_dff_A_SCuselYG2_0),.clk(gclk));
	jdff dff_A_7Z92uT2d2_0(.dout(w_dff_A_2j4uVMqg2_0),.din(w_dff_A_7Z92uT2d2_0),.clk(gclk));
	jdff dff_A_2j4uVMqg2_0(.dout(w_dff_A_0fuoSUpE0_0),.din(w_dff_A_2j4uVMqg2_0),.clk(gclk));
	jdff dff_A_0fuoSUpE0_0(.dout(w_dff_A_PLux0Fem7_0),.din(w_dff_A_0fuoSUpE0_0),.clk(gclk));
	jdff dff_A_PLux0Fem7_0(.dout(w_dff_A_sZAgWQbQ5_0),.din(w_dff_A_PLux0Fem7_0),.clk(gclk));
	jdff dff_A_sZAgWQbQ5_0(.dout(w_dff_A_ST7RWL082_0),.din(w_dff_A_sZAgWQbQ5_0),.clk(gclk));
	jdff dff_A_ST7RWL082_0(.dout(w_dff_A_miTjf7vK9_0),.din(w_dff_A_ST7RWL082_0),.clk(gclk));
	jdff dff_A_miTjf7vK9_0(.dout(w_dff_A_QJTWqxwc1_0),.din(w_dff_A_miTjf7vK9_0),.clk(gclk));
	jdff dff_A_QJTWqxwc1_0(.dout(w_dff_A_yI6rIQoi0_0),.din(w_dff_A_QJTWqxwc1_0),.clk(gclk));
	jdff dff_A_yI6rIQoi0_0(.dout(w_dff_A_naKFjRhr9_0),.din(w_dff_A_yI6rIQoi0_0),.clk(gclk));
	jdff dff_A_naKFjRhr9_0(.dout(w_dff_A_g43cBc1v4_0),.din(w_dff_A_naKFjRhr9_0),.clk(gclk));
	jdff dff_A_g43cBc1v4_0(.dout(w_dff_A_hpfzuxVx6_0),.din(w_dff_A_g43cBc1v4_0),.clk(gclk));
	jdff dff_A_hpfzuxVx6_0(.dout(w_dff_A_JDOqkfEf8_0),.din(w_dff_A_hpfzuxVx6_0),.clk(gclk));
	jdff dff_A_JDOqkfEf8_0(.dout(w_dff_A_gU9MVpxj7_0),.din(w_dff_A_JDOqkfEf8_0),.clk(gclk));
	jdff dff_A_gU9MVpxj7_0(.dout(w_dff_A_egeb3Qdl9_0),.din(w_dff_A_gU9MVpxj7_0),.clk(gclk));
	jdff dff_A_egeb3Qdl9_0(.dout(w_dff_A_BiyTWZcm5_0),.din(w_dff_A_egeb3Qdl9_0),.clk(gclk));
	jdff dff_A_BiyTWZcm5_0(.dout(w_dff_A_X1eUhFJm8_0),.din(w_dff_A_BiyTWZcm5_0),.clk(gclk));
	jdff dff_A_X1eUhFJm8_0(.dout(w_dff_A_Ilp4LSRo3_0),.din(w_dff_A_X1eUhFJm8_0),.clk(gclk));
	jdff dff_A_Ilp4LSRo3_0(.dout(f34),.din(w_dff_A_Ilp4LSRo3_0),.clk(gclk));
	jdff dff_A_tKTU1hRn7_2(.dout(w_dff_A_Ch2Oc2vb5_0),.din(w_dff_A_tKTU1hRn7_2),.clk(gclk));
	jdff dff_A_Ch2Oc2vb5_0(.dout(w_dff_A_nEGB37bK5_0),.din(w_dff_A_Ch2Oc2vb5_0),.clk(gclk));
	jdff dff_A_nEGB37bK5_0(.dout(w_dff_A_ZiGXwpii3_0),.din(w_dff_A_nEGB37bK5_0),.clk(gclk));
	jdff dff_A_ZiGXwpii3_0(.dout(w_dff_A_Q8VRtOFn1_0),.din(w_dff_A_ZiGXwpii3_0),.clk(gclk));
	jdff dff_A_Q8VRtOFn1_0(.dout(w_dff_A_VHdbFjJo8_0),.din(w_dff_A_Q8VRtOFn1_0),.clk(gclk));
	jdff dff_A_VHdbFjJo8_0(.dout(w_dff_A_hObWfp1Q2_0),.din(w_dff_A_VHdbFjJo8_0),.clk(gclk));
	jdff dff_A_hObWfp1Q2_0(.dout(w_dff_A_tpi6swYx9_0),.din(w_dff_A_hObWfp1Q2_0),.clk(gclk));
	jdff dff_A_tpi6swYx9_0(.dout(w_dff_A_wlGiXxif3_0),.din(w_dff_A_tpi6swYx9_0),.clk(gclk));
	jdff dff_A_wlGiXxif3_0(.dout(w_dff_A_ujbI0SNB8_0),.din(w_dff_A_wlGiXxif3_0),.clk(gclk));
	jdff dff_A_ujbI0SNB8_0(.dout(w_dff_A_DliQZfyC6_0),.din(w_dff_A_ujbI0SNB8_0),.clk(gclk));
	jdff dff_A_DliQZfyC6_0(.dout(w_dff_A_fOcyHfS14_0),.din(w_dff_A_DliQZfyC6_0),.clk(gclk));
	jdff dff_A_fOcyHfS14_0(.dout(w_dff_A_NFEmeulP6_0),.din(w_dff_A_fOcyHfS14_0),.clk(gclk));
	jdff dff_A_NFEmeulP6_0(.dout(w_dff_A_RO69BTiY7_0),.din(w_dff_A_NFEmeulP6_0),.clk(gclk));
	jdff dff_A_RO69BTiY7_0(.dout(w_dff_A_URj2PuUt2_0),.din(w_dff_A_RO69BTiY7_0),.clk(gclk));
	jdff dff_A_URj2PuUt2_0(.dout(w_dff_A_7Jdxw4nk7_0),.din(w_dff_A_URj2PuUt2_0),.clk(gclk));
	jdff dff_A_7Jdxw4nk7_0(.dout(w_dff_A_TzpHA0bX3_0),.din(w_dff_A_7Jdxw4nk7_0),.clk(gclk));
	jdff dff_A_TzpHA0bX3_0(.dout(w_dff_A_bzazDJTk5_0),.din(w_dff_A_TzpHA0bX3_0),.clk(gclk));
	jdff dff_A_bzazDJTk5_0(.dout(w_dff_A_eE9Ur35R2_0),.din(w_dff_A_bzazDJTk5_0),.clk(gclk));
	jdff dff_A_eE9Ur35R2_0(.dout(w_dff_A_LJpxmHmg6_0),.din(w_dff_A_eE9Ur35R2_0),.clk(gclk));
	jdff dff_A_LJpxmHmg6_0(.dout(w_dff_A_aS182kDO4_0),.din(w_dff_A_LJpxmHmg6_0),.clk(gclk));
	jdff dff_A_aS182kDO4_0(.dout(w_dff_A_0iGgeNPM6_0),.din(w_dff_A_aS182kDO4_0),.clk(gclk));
	jdff dff_A_0iGgeNPM6_0(.dout(w_dff_A_btKxdY4I0_0),.din(w_dff_A_0iGgeNPM6_0),.clk(gclk));
	jdff dff_A_btKxdY4I0_0(.dout(w_dff_A_0z5DsSvY5_0),.din(w_dff_A_btKxdY4I0_0),.clk(gclk));
	jdff dff_A_0z5DsSvY5_0(.dout(w_dff_A_TIZn6i9V6_0),.din(w_dff_A_0z5DsSvY5_0),.clk(gclk));
	jdff dff_A_TIZn6i9V6_0(.dout(w_dff_A_bIGOQxb50_0),.din(w_dff_A_TIZn6i9V6_0),.clk(gclk));
	jdff dff_A_bIGOQxb50_0(.dout(w_dff_A_rsTvC55X9_0),.din(w_dff_A_bIGOQxb50_0),.clk(gclk));
	jdff dff_A_rsTvC55X9_0(.dout(w_dff_A_fAX1yO723_0),.din(w_dff_A_rsTvC55X9_0),.clk(gclk));
	jdff dff_A_fAX1yO723_0(.dout(w_dff_A_AWg4IurG0_0),.din(w_dff_A_fAX1yO723_0),.clk(gclk));
	jdff dff_A_AWg4IurG0_0(.dout(w_dff_A_vZOxgZKa5_0),.din(w_dff_A_AWg4IurG0_0),.clk(gclk));
	jdff dff_A_vZOxgZKa5_0(.dout(w_dff_A_SHEgAk5h7_0),.din(w_dff_A_vZOxgZKa5_0),.clk(gclk));
	jdff dff_A_SHEgAk5h7_0(.dout(w_dff_A_sf0PebLT0_0),.din(w_dff_A_SHEgAk5h7_0),.clk(gclk));
	jdff dff_A_sf0PebLT0_0(.dout(w_dff_A_kQl7OQ3c1_0),.din(w_dff_A_sf0PebLT0_0),.clk(gclk));
	jdff dff_A_kQl7OQ3c1_0(.dout(w_dff_A_ADZ85spc2_0),.din(w_dff_A_kQl7OQ3c1_0),.clk(gclk));
	jdff dff_A_ADZ85spc2_0(.dout(w_dff_A_LorQSN5d3_0),.din(w_dff_A_ADZ85spc2_0),.clk(gclk));
	jdff dff_A_LorQSN5d3_0(.dout(w_dff_A_rEbafI8f1_0),.din(w_dff_A_LorQSN5d3_0),.clk(gclk));
	jdff dff_A_rEbafI8f1_0(.dout(w_dff_A_JpdLi8XN8_0),.din(w_dff_A_rEbafI8f1_0),.clk(gclk));
	jdff dff_A_JpdLi8XN8_0(.dout(w_dff_A_EH7Uq0tc1_0),.din(w_dff_A_JpdLi8XN8_0),.clk(gclk));
	jdff dff_A_EH7Uq0tc1_0(.dout(w_dff_A_hYcRuqmh7_0),.din(w_dff_A_EH7Uq0tc1_0),.clk(gclk));
	jdff dff_A_hYcRuqmh7_0(.dout(w_dff_A_GrHDx2OA1_0),.din(w_dff_A_hYcRuqmh7_0),.clk(gclk));
	jdff dff_A_GrHDx2OA1_0(.dout(w_dff_A_Ua3RxwqY9_0),.din(w_dff_A_GrHDx2OA1_0),.clk(gclk));
	jdff dff_A_Ua3RxwqY9_0(.dout(w_dff_A_5nrNoENL2_0),.din(w_dff_A_Ua3RxwqY9_0),.clk(gclk));
	jdff dff_A_5nrNoENL2_0(.dout(w_dff_A_u4BwEYyt4_0),.din(w_dff_A_5nrNoENL2_0),.clk(gclk));
	jdff dff_A_u4BwEYyt4_0(.dout(w_dff_A_rr7t9NPn8_0),.din(w_dff_A_u4BwEYyt4_0),.clk(gclk));
	jdff dff_A_rr7t9NPn8_0(.dout(w_dff_A_M0ZSeS8F3_0),.din(w_dff_A_rr7t9NPn8_0),.clk(gclk));
	jdff dff_A_M0ZSeS8F3_0(.dout(w_dff_A_hNN00mLk6_0),.din(w_dff_A_M0ZSeS8F3_0),.clk(gclk));
	jdff dff_A_hNN00mLk6_0(.dout(w_dff_A_LFaK89Zb7_0),.din(w_dff_A_hNN00mLk6_0),.clk(gclk));
	jdff dff_A_LFaK89Zb7_0(.dout(w_dff_A_TPKgoR8J2_0),.din(w_dff_A_LFaK89Zb7_0),.clk(gclk));
	jdff dff_A_TPKgoR8J2_0(.dout(w_dff_A_g8p3WKfb4_0),.din(w_dff_A_TPKgoR8J2_0),.clk(gclk));
	jdff dff_A_g8p3WKfb4_0(.dout(w_dff_A_cuh9UZAW3_0),.din(w_dff_A_g8p3WKfb4_0),.clk(gclk));
	jdff dff_A_cuh9UZAW3_0(.dout(w_dff_A_EJB30njP4_0),.din(w_dff_A_cuh9UZAW3_0),.clk(gclk));
	jdff dff_A_EJB30njP4_0(.dout(w_dff_A_Bf6PewtZ0_0),.din(w_dff_A_EJB30njP4_0),.clk(gclk));
	jdff dff_A_Bf6PewtZ0_0(.dout(w_dff_A_kF9UhB5E9_0),.din(w_dff_A_Bf6PewtZ0_0),.clk(gclk));
	jdff dff_A_kF9UhB5E9_0(.dout(w_dff_A_tAcKHAuS4_0),.din(w_dff_A_kF9UhB5E9_0),.clk(gclk));
	jdff dff_A_tAcKHAuS4_0(.dout(w_dff_A_vioj2Pha6_0),.din(w_dff_A_tAcKHAuS4_0),.clk(gclk));
	jdff dff_A_vioj2Pha6_0(.dout(w_dff_A_CStbZH4x4_0),.din(w_dff_A_vioj2Pha6_0),.clk(gclk));
	jdff dff_A_CStbZH4x4_0(.dout(w_dff_A_3rH5S1gQ1_0),.din(w_dff_A_CStbZH4x4_0),.clk(gclk));
	jdff dff_A_3rH5S1gQ1_0(.dout(w_dff_A_a63eicb86_0),.din(w_dff_A_3rH5S1gQ1_0),.clk(gclk));
	jdff dff_A_a63eicb86_0(.dout(w_dff_A_6fDPp9Ko2_0),.din(w_dff_A_a63eicb86_0),.clk(gclk));
	jdff dff_A_6fDPp9Ko2_0(.dout(w_dff_A_xXjgOvOx6_0),.din(w_dff_A_6fDPp9Ko2_0),.clk(gclk));
	jdff dff_A_xXjgOvOx6_0(.dout(w_dff_A_qsEblaWp6_0),.din(w_dff_A_xXjgOvOx6_0),.clk(gclk));
	jdff dff_A_qsEblaWp6_0(.dout(w_dff_A_VE8F3smc3_0),.din(w_dff_A_qsEblaWp6_0),.clk(gclk));
	jdff dff_A_VE8F3smc3_0(.dout(w_dff_A_7dyisAIS6_0),.din(w_dff_A_VE8F3smc3_0),.clk(gclk));
	jdff dff_A_7dyisAIS6_0(.dout(w_dff_A_BlMmpKU17_0),.din(w_dff_A_7dyisAIS6_0),.clk(gclk));
	jdff dff_A_BlMmpKU17_0(.dout(w_dff_A_UmSf4Fxd1_0),.din(w_dff_A_BlMmpKU17_0),.clk(gclk));
	jdff dff_A_UmSf4Fxd1_0(.dout(w_dff_A_m9VmeOCU6_0),.din(w_dff_A_UmSf4Fxd1_0),.clk(gclk));
	jdff dff_A_m9VmeOCU6_0(.dout(w_dff_A_JDSlJP507_0),.din(w_dff_A_m9VmeOCU6_0),.clk(gclk));
	jdff dff_A_JDSlJP507_0(.dout(w_dff_A_kwUMshQW9_0),.din(w_dff_A_JDSlJP507_0),.clk(gclk));
	jdff dff_A_kwUMshQW9_0(.dout(w_dff_A_H1DIgAo81_0),.din(w_dff_A_kwUMshQW9_0),.clk(gclk));
	jdff dff_A_H1DIgAo81_0(.dout(w_dff_A_cDG6dHMF3_0),.din(w_dff_A_H1DIgAo81_0),.clk(gclk));
	jdff dff_A_cDG6dHMF3_0(.dout(w_dff_A_wTl97SuH3_0),.din(w_dff_A_cDG6dHMF3_0),.clk(gclk));
	jdff dff_A_wTl97SuH3_0(.dout(w_dff_A_fOBCRBWX0_0),.din(w_dff_A_wTl97SuH3_0),.clk(gclk));
	jdff dff_A_fOBCRBWX0_0(.dout(w_dff_A_UW2g8f6K7_0),.din(w_dff_A_fOBCRBWX0_0),.clk(gclk));
	jdff dff_A_UW2g8f6K7_0(.dout(w_dff_A_Jzq2nXK18_0),.din(w_dff_A_UW2g8f6K7_0),.clk(gclk));
	jdff dff_A_Jzq2nXK18_0(.dout(w_dff_A_qML8P6q92_0),.din(w_dff_A_Jzq2nXK18_0),.clk(gclk));
	jdff dff_A_qML8P6q92_0(.dout(w_dff_A_rNbqGuBL8_0),.din(w_dff_A_qML8P6q92_0),.clk(gclk));
	jdff dff_A_rNbqGuBL8_0(.dout(w_dff_A_IJbS29KA6_0),.din(w_dff_A_rNbqGuBL8_0),.clk(gclk));
	jdff dff_A_IJbS29KA6_0(.dout(w_dff_A_VpMBkWWc6_0),.din(w_dff_A_IJbS29KA6_0),.clk(gclk));
	jdff dff_A_VpMBkWWc6_0(.dout(w_dff_A_VXEiqVYQ0_0),.din(w_dff_A_VpMBkWWc6_0),.clk(gclk));
	jdff dff_A_VXEiqVYQ0_0(.dout(w_dff_A_J3s55izY0_0),.din(w_dff_A_VXEiqVYQ0_0),.clk(gclk));
	jdff dff_A_J3s55izY0_0(.dout(w_dff_A_lBsBNlMg3_0),.din(w_dff_A_J3s55izY0_0),.clk(gclk));
	jdff dff_A_lBsBNlMg3_0(.dout(w_dff_A_KGShAaPC6_0),.din(w_dff_A_lBsBNlMg3_0),.clk(gclk));
	jdff dff_A_KGShAaPC6_0(.dout(w_dff_A_iYupWikI9_0),.din(w_dff_A_KGShAaPC6_0),.clk(gclk));
	jdff dff_A_iYupWikI9_0(.dout(w_dff_A_Ky1TfkKH7_0),.din(w_dff_A_iYupWikI9_0),.clk(gclk));
	jdff dff_A_Ky1TfkKH7_0(.dout(w_dff_A_yg6YV2HR6_0),.din(w_dff_A_Ky1TfkKH7_0),.clk(gclk));
	jdff dff_A_yg6YV2HR6_0(.dout(w_dff_A_daVDB4VH8_0),.din(w_dff_A_yg6YV2HR6_0),.clk(gclk));
	jdff dff_A_daVDB4VH8_0(.dout(w_dff_A_tW5EWCgl4_0),.din(w_dff_A_daVDB4VH8_0),.clk(gclk));
	jdff dff_A_tW5EWCgl4_0(.dout(w_dff_A_0Yg2Inx50_0),.din(w_dff_A_tW5EWCgl4_0),.clk(gclk));
	jdff dff_A_0Yg2Inx50_0(.dout(w_dff_A_araptS9w7_0),.din(w_dff_A_0Yg2Inx50_0),.clk(gclk));
	jdff dff_A_araptS9w7_0(.dout(w_dff_A_qtWGmOkL9_0),.din(w_dff_A_araptS9w7_0),.clk(gclk));
	jdff dff_A_qtWGmOkL9_0(.dout(w_dff_A_MsxhfmAU1_0),.din(w_dff_A_qtWGmOkL9_0),.clk(gclk));
	jdff dff_A_MsxhfmAU1_0(.dout(w_dff_A_WB1oNc4C1_0),.din(w_dff_A_MsxhfmAU1_0),.clk(gclk));
	jdff dff_A_WB1oNc4C1_0(.dout(f35),.din(w_dff_A_WB1oNc4C1_0),.clk(gclk));
	jdff dff_A_F7Oq80ij2_2(.dout(w_dff_A_bvG6h68p8_0),.din(w_dff_A_F7Oq80ij2_2),.clk(gclk));
	jdff dff_A_bvG6h68p8_0(.dout(w_dff_A_kKbT802A6_0),.din(w_dff_A_bvG6h68p8_0),.clk(gclk));
	jdff dff_A_kKbT802A6_0(.dout(w_dff_A_TicpFAni1_0),.din(w_dff_A_kKbT802A6_0),.clk(gclk));
	jdff dff_A_TicpFAni1_0(.dout(w_dff_A_e1ZMROkg9_0),.din(w_dff_A_TicpFAni1_0),.clk(gclk));
	jdff dff_A_e1ZMROkg9_0(.dout(w_dff_A_xtQuLvzQ0_0),.din(w_dff_A_e1ZMROkg9_0),.clk(gclk));
	jdff dff_A_xtQuLvzQ0_0(.dout(w_dff_A_FyNeBQTy3_0),.din(w_dff_A_xtQuLvzQ0_0),.clk(gclk));
	jdff dff_A_FyNeBQTy3_0(.dout(w_dff_A_ajSyLEgZ9_0),.din(w_dff_A_FyNeBQTy3_0),.clk(gclk));
	jdff dff_A_ajSyLEgZ9_0(.dout(w_dff_A_UuGRcLn26_0),.din(w_dff_A_ajSyLEgZ9_0),.clk(gclk));
	jdff dff_A_UuGRcLn26_0(.dout(w_dff_A_0GLxM1s98_0),.din(w_dff_A_UuGRcLn26_0),.clk(gclk));
	jdff dff_A_0GLxM1s98_0(.dout(w_dff_A_uyO9Rpkf1_0),.din(w_dff_A_0GLxM1s98_0),.clk(gclk));
	jdff dff_A_uyO9Rpkf1_0(.dout(w_dff_A_EeGEq80i9_0),.din(w_dff_A_uyO9Rpkf1_0),.clk(gclk));
	jdff dff_A_EeGEq80i9_0(.dout(w_dff_A_5Pbfy8tK5_0),.din(w_dff_A_EeGEq80i9_0),.clk(gclk));
	jdff dff_A_5Pbfy8tK5_0(.dout(w_dff_A_GlZW5Kgo0_0),.din(w_dff_A_5Pbfy8tK5_0),.clk(gclk));
	jdff dff_A_GlZW5Kgo0_0(.dout(w_dff_A_wrqmMmbC5_0),.din(w_dff_A_GlZW5Kgo0_0),.clk(gclk));
	jdff dff_A_wrqmMmbC5_0(.dout(w_dff_A_L6InOzRZ7_0),.din(w_dff_A_wrqmMmbC5_0),.clk(gclk));
	jdff dff_A_L6InOzRZ7_0(.dout(w_dff_A_h48qxO9F9_0),.din(w_dff_A_L6InOzRZ7_0),.clk(gclk));
	jdff dff_A_h48qxO9F9_0(.dout(w_dff_A_SEgcmIzs9_0),.din(w_dff_A_h48qxO9F9_0),.clk(gclk));
	jdff dff_A_SEgcmIzs9_0(.dout(w_dff_A_PVqVZHZZ2_0),.din(w_dff_A_SEgcmIzs9_0),.clk(gclk));
	jdff dff_A_PVqVZHZZ2_0(.dout(w_dff_A_Dt7Yzrww5_0),.din(w_dff_A_PVqVZHZZ2_0),.clk(gclk));
	jdff dff_A_Dt7Yzrww5_0(.dout(w_dff_A_0fVxvMb70_0),.din(w_dff_A_Dt7Yzrww5_0),.clk(gclk));
	jdff dff_A_0fVxvMb70_0(.dout(w_dff_A_pMf4uDEF6_0),.din(w_dff_A_0fVxvMb70_0),.clk(gclk));
	jdff dff_A_pMf4uDEF6_0(.dout(w_dff_A_knFVBxyb9_0),.din(w_dff_A_pMf4uDEF6_0),.clk(gclk));
	jdff dff_A_knFVBxyb9_0(.dout(w_dff_A_BypINXjO1_0),.din(w_dff_A_knFVBxyb9_0),.clk(gclk));
	jdff dff_A_BypINXjO1_0(.dout(w_dff_A_w2M4RpAV5_0),.din(w_dff_A_BypINXjO1_0),.clk(gclk));
	jdff dff_A_w2M4RpAV5_0(.dout(w_dff_A_w4BLgTFP6_0),.din(w_dff_A_w2M4RpAV5_0),.clk(gclk));
	jdff dff_A_w4BLgTFP6_0(.dout(w_dff_A_hkIpvIyN3_0),.din(w_dff_A_w4BLgTFP6_0),.clk(gclk));
	jdff dff_A_hkIpvIyN3_0(.dout(w_dff_A_by0cmANi0_0),.din(w_dff_A_hkIpvIyN3_0),.clk(gclk));
	jdff dff_A_by0cmANi0_0(.dout(w_dff_A_gKUxMeCj6_0),.din(w_dff_A_by0cmANi0_0),.clk(gclk));
	jdff dff_A_gKUxMeCj6_0(.dout(w_dff_A_yIdPt0dq0_0),.din(w_dff_A_gKUxMeCj6_0),.clk(gclk));
	jdff dff_A_yIdPt0dq0_0(.dout(w_dff_A_k6mVzKPC9_0),.din(w_dff_A_yIdPt0dq0_0),.clk(gclk));
	jdff dff_A_k6mVzKPC9_0(.dout(w_dff_A_OGdVz8h07_0),.din(w_dff_A_k6mVzKPC9_0),.clk(gclk));
	jdff dff_A_OGdVz8h07_0(.dout(w_dff_A_JR1LEqV33_0),.din(w_dff_A_OGdVz8h07_0),.clk(gclk));
	jdff dff_A_JR1LEqV33_0(.dout(w_dff_A_oA4uXYQI7_0),.din(w_dff_A_JR1LEqV33_0),.clk(gclk));
	jdff dff_A_oA4uXYQI7_0(.dout(w_dff_A_YeIbYm5q5_0),.din(w_dff_A_oA4uXYQI7_0),.clk(gclk));
	jdff dff_A_YeIbYm5q5_0(.dout(w_dff_A_Fad9lO6K7_0),.din(w_dff_A_YeIbYm5q5_0),.clk(gclk));
	jdff dff_A_Fad9lO6K7_0(.dout(w_dff_A_fP4VwOhA7_0),.din(w_dff_A_Fad9lO6K7_0),.clk(gclk));
	jdff dff_A_fP4VwOhA7_0(.dout(w_dff_A_wPGXAP1T8_0),.din(w_dff_A_fP4VwOhA7_0),.clk(gclk));
	jdff dff_A_wPGXAP1T8_0(.dout(w_dff_A_X5uy6Ul89_0),.din(w_dff_A_wPGXAP1T8_0),.clk(gclk));
	jdff dff_A_X5uy6Ul89_0(.dout(w_dff_A_5MU8qTkR3_0),.din(w_dff_A_X5uy6Ul89_0),.clk(gclk));
	jdff dff_A_5MU8qTkR3_0(.dout(w_dff_A_mta8aeIC9_0),.din(w_dff_A_5MU8qTkR3_0),.clk(gclk));
	jdff dff_A_mta8aeIC9_0(.dout(w_dff_A_lCezDUmS6_0),.din(w_dff_A_mta8aeIC9_0),.clk(gclk));
	jdff dff_A_lCezDUmS6_0(.dout(w_dff_A_GE9EpR9Y7_0),.din(w_dff_A_lCezDUmS6_0),.clk(gclk));
	jdff dff_A_GE9EpR9Y7_0(.dout(w_dff_A_gbC5Q28i4_0),.din(w_dff_A_GE9EpR9Y7_0),.clk(gclk));
	jdff dff_A_gbC5Q28i4_0(.dout(w_dff_A_oOrZQhdc6_0),.din(w_dff_A_gbC5Q28i4_0),.clk(gclk));
	jdff dff_A_oOrZQhdc6_0(.dout(w_dff_A_MshdEHUA3_0),.din(w_dff_A_oOrZQhdc6_0),.clk(gclk));
	jdff dff_A_MshdEHUA3_0(.dout(w_dff_A_GTVZegty5_0),.din(w_dff_A_MshdEHUA3_0),.clk(gclk));
	jdff dff_A_GTVZegty5_0(.dout(w_dff_A_upm7cW246_0),.din(w_dff_A_GTVZegty5_0),.clk(gclk));
	jdff dff_A_upm7cW246_0(.dout(w_dff_A_sFSjVZGK3_0),.din(w_dff_A_upm7cW246_0),.clk(gclk));
	jdff dff_A_sFSjVZGK3_0(.dout(w_dff_A_Hs4VEL4d4_0),.din(w_dff_A_sFSjVZGK3_0),.clk(gclk));
	jdff dff_A_Hs4VEL4d4_0(.dout(w_dff_A_sOsttbQ18_0),.din(w_dff_A_Hs4VEL4d4_0),.clk(gclk));
	jdff dff_A_sOsttbQ18_0(.dout(w_dff_A_YYe81kyk5_0),.din(w_dff_A_sOsttbQ18_0),.clk(gclk));
	jdff dff_A_YYe81kyk5_0(.dout(w_dff_A_9BGgxj7j8_0),.din(w_dff_A_YYe81kyk5_0),.clk(gclk));
	jdff dff_A_9BGgxj7j8_0(.dout(w_dff_A_vhGKTBuB6_0),.din(w_dff_A_9BGgxj7j8_0),.clk(gclk));
	jdff dff_A_vhGKTBuB6_0(.dout(w_dff_A_GNCaruMB7_0),.din(w_dff_A_vhGKTBuB6_0),.clk(gclk));
	jdff dff_A_GNCaruMB7_0(.dout(w_dff_A_xye2GpFu8_0),.din(w_dff_A_GNCaruMB7_0),.clk(gclk));
	jdff dff_A_xye2GpFu8_0(.dout(w_dff_A_q4ossp9T8_0),.din(w_dff_A_xye2GpFu8_0),.clk(gclk));
	jdff dff_A_q4ossp9T8_0(.dout(w_dff_A_gQtgonkD1_0),.din(w_dff_A_q4ossp9T8_0),.clk(gclk));
	jdff dff_A_gQtgonkD1_0(.dout(w_dff_A_AbmdYSKy3_0),.din(w_dff_A_gQtgonkD1_0),.clk(gclk));
	jdff dff_A_AbmdYSKy3_0(.dout(w_dff_A_NB4PiZFN3_0),.din(w_dff_A_AbmdYSKy3_0),.clk(gclk));
	jdff dff_A_NB4PiZFN3_0(.dout(w_dff_A_qTodR5Bt9_0),.din(w_dff_A_NB4PiZFN3_0),.clk(gclk));
	jdff dff_A_qTodR5Bt9_0(.dout(w_dff_A_Wt4m43OV1_0),.din(w_dff_A_qTodR5Bt9_0),.clk(gclk));
	jdff dff_A_Wt4m43OV1_0(.dout(w_dff_A_tRnFLsr66_0),.din(w_dff_A_Wt4m43OV1_0),.clk(gclk));
	jdff dff_A_tRnFLsr66_0(.dout(w_dff_A_QTLzNcJ88_0),.din(w_dff_A_tRnFLsr66_0),.clk(gclk));
	jdff dff_A_QTLzNcJ88_0(.dout(w_dff_A_wMLmqWG17_0),.din(w_dff_A_QTLzNcJ88_0),.clk(gclk));
	jdff dff_A_wMLmqWG17_0(.dout(w_dff_A_eZVlgkM91_0),.din(w_dff_A_wMLmqWG17_0),.clk(gclk));
	jdff dff_A_eZVlgkM91_0(.dout(w_dff_A_CQOseGOU6_0),.din(w_dff_A_eZVlgkM91_0),.clk(gclk));
	jdff dff_A_CQOseGOU6_0(.dout(w_dff_A_7TdwLPkn1_0),.din(w_dff_A_CQOseGOU6_0),.clk(gclk));
	jdff dff_A_7TdwLPkn1_0(.dout(w_dff_A_NCc31cjr8_0),.din(w_dff_A_7TdwLPkn1_0),.clk(gclk));
	jdff dff_A_NCc31cjr8_0(.dout(w_dff_A_KRXCyJt87_0),.din(w_dff_A_NCc31cjr8_0),.clk(gclk));
	jdff dff_A_KRXCyJt87_0(.dout(w_dff_A_GkQWWBe95_0),.din(w_dff_A_KRXCyJt87_0),.clk(gclk));
	jdff dff_A_GkQWWBe95_0(.dout(w_dff_A_mkdNoieO8_0),.din(w_dff_A_GkQWWBe95_0),.clk(gclk));
	jdff dff_A_mkdNoieO8_0(.dout(w_dff_A_qGr3qz6b0_0),.din(w_dff_A_mkdNoieO8_0),.clk(gclk));
	jdff dff_A_qGr3qz6b0_0(.dout(w_dff_A_9hMEaNkN1_0),.din(w_dff_A_qGr3qz6b0_0),.clk(gclk));
	jdff dff_A_9hMEaNkN1_0(.dout(w_dff_A_L6ecBm7o4_0),.din(w_dff_A_9hMEaNkN1_0),.clk(gclk));
	jdff dff_A_L6ecBm7o4_0(.dout(w_dff_A_TivH4GlN0_0),.din(w_dff_A_L6ecBm7o4_0),.clk(gclk));
	jdff dff_A_TivH4GlN0_0(.dout(w_dff_A_vdxWXSlF0_0),.din(w_dff_A_TivH4GlN0_0),.clk(gclk));
	jdff dff_A_vdxWXSlF0_0(.dout(w_dff_A_MelRwXzO6_0),.din(w_dff_A_vdxWXSlF0_0),.clk(gclk));
	jdff dff_A_MelRwXzO6_0(.dout(w_dff_A_BR0LuR3Q9_0),.din(w_dff_A_MelRwXzO6_0),.clk(gclk));
	jdff dff_A_BR0LuR3Q9_0(.dout(w_dff_A_N1YXJyvb9_0),.din(w_dff_A_BR0LuR3Q9_0),.clk(gclk));
	jdff dff_A_N1YXJyvb9_0(.dout(w_dff_A_gnlIbS416_0),.din(w_dff_A_N1YXJyvb9_0),.clk(gclk));
	jdff dff_A_gnlIbS416_0(.dout(w_dff_A_lkE8GRpU2_0),.din(w_dff_A_gnlIbS416_0),.clk(gclk));
	jdff dff_A_lkE8GRpU2_0(.dout(w_dff_A_XOL0iivq7_0),.din(w_dff_A_lkE8GRpU2_0),.clk(gclk));
	jdff dff_A_XOL0iivq7_0(.dout(w_dff_A_5Gv1WFMd0_0),.din(w_dff_A_XOL0iivq7_0),.clk(gclk));
	jdff dff_A_5Gv1WFMd0_0(.dout(w_dff_A_nv1F8qll0_0),.din(w_dff_A_5Gv1WFMd0_0),.clk(gclk));
	jdff dff_A_nv1F8qll0_0(.dout(w_dff_A_t7giiDop1_0),.din(w_dff_A_nv1F8qll0_0),.clk(gclk));
	jdff dff_A_t7giiDop1_0(.dout(w_dff_A_Io4Iw7zF1_0),.din(w_dff_A_t7giiDop1_0),.clk(gclk));
	jdff dff_A_Io4Iw7zF1_0(.dout(w_dff_A_I3u4EcEE3_0),.din(w_dff_A_Io4Iw7zF1_0),.clk(gclk));
	jdff dff_A_I3u4EcEE3_0(.dout(w_dff_A_DdJUbF8B1_0),.din(w_dff_A_I3u4EcEE3_0),.clk(gclk));
	jdff dff_A_DdJUbF8B1_0(.dout(w_dff_A_IJBDKL7L4_0),.din(w_dff_A_DdJUbF8B1_0),.clk(gclk));
	jdff dff_A_IJBDKL7L4_0(.dout(w_dff_A_FK59F2FA3_0),.din(w_dff_A_IJBDKL7L4_0),.clk(gclk));
	jdff dff_A_FK59F2FA3_0(.dout(f36),.din(w_dff_A_FK59F2FA3_0),.clk(gclk));
	jdff dff_A_nym5NQ194_2(.dout(w_dff_A_z8rrjKwU6_0),.din(w_dff_A_nym5NQ194_2),.clk(gclk));
	jdff dff_A_z8rrjKwU6_0(.dout(w_dff_A_I4QKR9tw3_0),.din(w_dff_A_z8rrjKwU6_0),.clk(gclk));
	jdff dff_A_I4QKR9tw3_0(.dout(w_dff_A_Qkr7HnZx3_0),.din(w_dff_A_I4QKR9tw3_0),.clk(gclk));
	jdff dff_A_Qkr7HnZx3_0(.dout(w_dff_A_3eRx8es30_0),.din(w_dff_A_Qkr7HnZx3_0),.clk(gclk));
	jdff dff_A_3eRx8es30_0(.dout(w_dff_A_qreLIVrI2_0),.din(w_dff_A_3eRx8es30_0),.clk(gclk));
	jdff dff_A_qreLIVrI2_0(.dout(w_dff_A_DMbCWc4Y4_0),.din(w_dff_A_qreLIVrI2_0),.clk(gclk));
	jdff dff_A_DMbCWc4Y4_0(.dout(w_dff_A_wG63FlUr6_0),.din(w_dff_A_DMbCWc4Y4_0),.clk(gclk));
	jdff dff_A_wG63FlUr6_0(.dout(w_dff_A_qL5P0RMW8_0),.din(w_dff_A_wG63FlUr6_0),.clk(gclk));
	jdff dff_A_qL5P0RMW8_0(.dout(w_dff_A_2bR3qjOS5_0),.din(w_dff_A_qL5P0RMW8_0),.clk(gclk));
	jdff dff_A_2bR3qjOS5_0(.dout(w_dff_A_LFSaiEVS3_0),.din(w_dff_A_2bR3qjOS5_0),.clk(gclk));
	jdff dff_A_LFSaiEVS3_0(.dout(w_dff_A_HlvMhO3J8_0),.din(w_dff_A_LFSaiEVS3_0),.clk(gclk));
	jdff dff_A_HlvMhO3J8_0(.dout(w_dff_A_RMJfd49g2_0),.din(w_dff_A_HlvMhO3J8_0),.clk(gclk));
	jdff dff_A_RMJfd49g2_0(.dout(w_dff_A_CYTDBucW7_0),.din(w_dff_A_RMJfd49g2_0),.clk(gclk));
	jdff dff_A_CYTDBucW7_0(.dout(w_dff_A_SodQK0h88_0),.din(w_dff_A_CYTDBucW7_0),.clk(gclk));
	jdff dff_A_SodQK0h88_0(.dout(w_dff_A_S8cMXxxy9_0),.din(w_dff_A_SodQK0h88_0),.clk(gclk));
	jdff dff_A_S8cMXxxy9_0(.dout(w_dff_A_K5EtG5RS6_0),.din(w_dff_A_S8cMXxxy9_0),.clk(gclk));
	jdff dff_A_K5EtG5RS6_0(.dout(w_dff_A_artkEDXD3_0),.din(w_dff_A_K5EtG5RS6_0),.clk(gclk));
	jdff dff_A_artkEDXD3_0(.dout(w_dff_A_Vly9DdtO7_0),.din(w_dff_A_artkEDXD3_0),.clk(gclk));
	jdff dff_A_Vly9DdtO7_0(.dout(w_dff_A_1kFvQbYh5_0),.din(w_dff_A_Vly9DdtO7_0),.clk(gclk));
	jdff dff_A_1kFvQbYh5_0(.dout(w_dff_A_XEVR1Y7w9_0),.din(w_dff_A_1kFvQbYh5_0),.clk(gclk));
	jdff dff_A_XEVR1Y7w9_0(.dout(w_dff_A_ZPbTvxwl7_0),.din(w_dff_A_XEVR1Y7w9_0),.clk(gclk));
	jdff dff_A_ZPbTvxwl7_0(.dout(w_dff_A_BOSLCrtr8_0),.din(w_dff_A_ZPbTvxwl7_0),.clk(gclk));
	jdff dff_A_BOSLCrtr8_0(.dout(w_dff_A_DHHMuR2n9_0),.din(w_dff_A_BOSLCrtr8_0),.clk(gclk));
	jdff dff_A_DHHMuR2n9_0(.dout(w_dff_A_qj7VCTNE5_0),.din(w_dff_A_DHHMuR2n9_0),.clk(gclk));
	jdff dff_A_qj7VCTNE5_0(.dout(w_dff_A_n0SqvMtf9_0),.din(w_dff_A_qj7VCTNE5_0),.clk(gclk));
	jdff dff_A_n0SqvMtf9_0(.dout(w_dff_A_gA2cuz2X1_0),.din(w_dff_A_n0SqvMtf9_0),.clk(gclk));
	jdff dff_A_gA2cuz2X1_0(.dout(w_dff_A_bYe5LaRl5_0),.din(w_dff_A_gA2cuz2X1_0),.clk(gclk));
	jdff dff_A_bYe5LaRl5_0(.dout(w_dff_A_LTMo0VBu4_0),.din(w_dff_A_bYe5LaRl5_0),.clk(gclk));
	jdff dff_A_LTMo0VBu4_0(.dout(w_dff_A_3KheANi86_0),.din(w_dff_A_LTMo0VBu4_0),.clk(gclk));
	jdff dff_A_3KheANi86_0(.dout(w_dff_A_JdqDOIb96_0),.din(w_dff_A_3KheANi86_0),.clk(gclk));
	jdff dff_A_JdqDOIb96_0(.dout(w_dff_A_V9D0exUG8_0),.din(w_dff_A_JdqDOIb96_0),.clk(gclk));
	jdff dff_A_V9D0exUG8_0(.dout(w_dff_A_43DpmDBQ5_0),.din(w_dff_A_V9D0exUG8_0),.clk(gclk));
	jdff dff_A_43DpmDBQ5_0(.dout(w_dff_A_8g3R5jU41_0),.din(w_dff_A_43DpmDBQ5_0),.clk(gclk));
	jdff dff_A_8g3R5jU41_0(.dout(w_dff_A_medKfdVW2_0),.din(w_dff_A_8g3R5jU41_0),.clk(gclk));
	jdff dff_A_medKfdVW2_0(.dout(w_dff_A_tMBVcawi7_0),.din(w_dff_A_medKfdVW2_0),.clk(gclk));
	jdff dff_A_tMBVcawi7_0(.dout(w_dff_A_Qb1M4P9u9_0),.din(w_dff_A_tMBVcawi7_0),.clk(gclk));
	jdff dff_A_Qb1M4P9u9_0(.dout(w_dff_A_d2p1vxxE4_0),.din(w_dff_A_Qb1M4P9u9_0),.clk(gclk));
	jdff dff_A_d2p1vxxE4_0(.dout(w_dff_A_yOyycVXV7_0),.din(w_dff_A_d2p1vxxE4_0),.clk(gclk));
	jdff dff_A_yOyycVXV7_0(.dout(w_dff_A_nyf4qYJ29_0),.din(w_dff_A_yOyycVXV7_0),.clk(gclk));
	jdff dff_A_nyf4qYJ29_0(.dout(w_dff_A_ODP5KXIC3_0),.din(w_dff_A_nyf4qYJ29_0),.clk(gclk));
	jdff dff_A_ODP5KXIC3_0(.dout(w_dff_A_8nOVQr7W5_0),.din(w_dff_A_ODP5KXIC3_0),.clk(gclk));
	jdff dff_A_8nOVQr7W5_0(.dout(w_dff_A_pfXDxnML3_0),.din(w_dff_A_8nOVQr7W5_0),.clk(gclk));
	jdff dff_A_pfXDxnML3_0(.dout(w_dff_A_qP8o6VDr9_0),.din(w_dff_A_pfXDxnML3_0),.clk(gclk));
	jdff dff_A_qP8o6VDr9_0(.dout(w_dff_A_LkUz6N6u9_0),.din(w_dff_A_qP8o6VDr9_0),.clk(gclk));
	jdff dff_A_LkUz6N6u9_0(.dout(w_dff_A_nlAmtiG30_0),.din(w_dff_A_LkUz6N6u9_0),.clk(gclk));
	jdff dff_A_nlAmtiG30_0(.dout(w_dff_A_MaaPbLPz7_0),.din(w_dff_A_nlAmtiG30_0),.clk(gclk));
	jdff dff_A_MaaPbLPz7_0(.dout(w_dff_A_7mtMJiAr6_0),.din(w_dff_A_MaaPbLPz7_0),.clk(gclk));
	jdff dff_A_7mtMJiAr6_0(.dout(w_dff_A_M5zgZ8059_0),.din(w_dff_A_7mtMJiAr6_0),.clk(gclk));
	jdff dff_A_M5zgZ8059_0(.dout(w_dff_A_H2KMaoOE6_0),.din(w_dff_A_M5zgZ8059_0),.clk(gclk));
	jdff dff_A_H2KMaoOE6_0(.dout(w_dff_A_GMgvfOpi1_0),.din(w_dff_A_H2KMaoOE6_0),.clk(gclk));
	jdff dff_A_GMgvfOpi1_0(.dout(w_dff_A_ggWpBlY67_0),.din(w_dff_A_GMgvfOpi1_0),.clk(gclk));
	jdff dff_A_ggWpBlY67_0(.dout(w_dff_A_nKF4HeOX3_0),.din(w_dff_A_ggWpBlY67_0),.clk(gclk));
	jdff dff_A_nKF4HeOX3_0(.dout(w_dff_A_hr0nIN654_0),.din(w_dff_A_nKF4HeOX3_0),.clk(gclk));
	jdff dff_A_hr0nIN654_0(.dout(w_dff_A_E8388oFY9_0),.din(w_dff_A_hr0nIN654_0),.clk(gclk));
	jdff dff_A_E8388oFY9_0(.dout(w_dff_A_IMqEEpQW4_0),.din(w_dff_A_E8388oFY9_0),.clk(gclk));
	jdff dff_A_IMqEEpQW4_0(.dout(w_dff_A_54XMmjVF9_0),.din(w_dff_A_IMqEEpQW4_0),.clk(gclk));
	jdff dff_A_54XMmjVF9_0(.dout(w_dff_A_3MGLJkYM7_0),.din(w_dff_A_54XMmjVF9_0),.clk(gclk));
	jdff dff_A_3MGLJkYM7_0(.dout(w_dff_A_l27ASzcF2_0),.din(w_dff_A_3MGLJkYM7_0),.clk(gclk));
	jdff dff_A_l27ASzcF2_0(.dout(w_dff_A_IXlO26rX6_0),.din(w_dff_A_l27ASzcF2_0),.clk(gclk));
	jdff dff_A_IXlO26rX6_0(.dout(w_dff_A_jiV4oIti1_0),.din(w_dff_A_IXlO26rX6_0),.clk(gclk));
	jdff dff_A_jiV4oIti1_0(.dout(w_dff_A_IthNF00f4_0),.din(w_dff_A_jiV4oIti1_0),.clk(gclk));
	jdff dff_A_IthNF00f4_0(.dout(w_dff_A_A0HzUWp40_0),.din(w_dff_A_IthNF00f4_0),.clk(gclk));
	jdff dff_A_A0HzUWp40_0(.dout(w_dff_A_I4rSGf2Q4_0),.din(w_dff_A_A0HzUWp40_0),.clk(gclk));
	jdff dff_A_I4rSGf2Q4_0(.dout(w_dff_A_EMnpFW7I4_0),.din(w_dff_A_I4rSGf2Q4_0),.clk(gclk));
	jdff dff_A_EMnpFW7I4_0(.dout(w_dff_A_SPFTZNXB6_0),.din(w_dff_A_EMnpFW7I4_0),.clk(gclk));
	jdff dff_A_SPFTZNXB6_0(.dout(w_dff_A_YHKBeXrG2_0),.din(w_dff_A_SPFTZNXB6_0),.clk(gclk));
	jdff dff_A_YHKBeXrG2_0(.dout(w_dff_A_xoIaY69s6_0),.din(w_dff_A_YHKBeXrG2_0),.clk(gclk));
	jdff dff_A_xoIaY69s6_0(.dout(w_dff_A_GTIU1wQ27_0),.din(w_dff_A_xoIaY69s6_0),.clk(gclk));
	jdff dff_A_GTIU1wQ27_0(.dout(w_dff_A_2cuCh8Y87_0),.din(w_dff_A_GTIU1wQ27_0),.clk(gclk));
	jdff dff_A_2cuCh8Y87_0(.dout(w_dff_A_vo8qKwrs9_0),.din(w_dff_A_2cuCh8Y87_0),.clk(gclk));
	jdff dff_A_vo8qKwrs9_0(.dout(w_dff_A_PfDLiwR91_0),.din(w_dff_A_vo8qKwrs9_0),.clk(gclk));
	jdff dff_A_PfDLiwR91_0(.dout(w_dff_A_aQ8ttUdW6_0),.din(w_dff_A_PfDLiwR91_0),.clk(gclk));
	jdff dff_A_aQ8ttUdW6_0(.dout(w_dff_A_Y00BZPE67_0),.din(w_dff_A_aQ8ttUdW6_0),.clk(gclk));
	jdff dff_A_Y00BZPE67_0(.dout(w_dff_A_FVU385FV6_0),.din(w_dff_A_Y00BZPE67_0),.clk(gclk));
	jdff dff_A_FVU385FV6_0(.dout(w_dff_A_28daTBMc4_0),.din(w_dff_A_FVU385FV6_0),.clk(gclk));
	jdff dff_A_28daTBMc4_0(.dout(w_dff_A_azsgFpCz9_0),.din(w_dff_A_28daTBMc4_0),.clk(gclk));
	jdff dff_A_azsgFpCz9_0(.dout(w_dff_A_MQptl2Hn9_0),.din(w_dff_A_azsgFpCz9_0),.clk(gclk));
	jdff dff_A_MQptl2Hn9_0(.dout(w_dff_A_BHMXI4SY3_0),.din(w_dff_A_MQptl2Hn9_0),.clk(gclk));
	jdff dff_A_BHMXI4SY3_0(.dout(w_dff_A_Cj3jlpbe7_0),.din(w_dff_A_BHMXI4SY3_0),.clk(gclk));
	jdff dff_A_Cj3jlpbe7_0(.dout(w_dff_A_wvFR0Uve3_0),.din(w_dff_A_Cj3jlpbe7_0),.clk(gclk));
	jdff dff_A_wvFR0Uve3_0(.dout(w_dff_A_JgJPasJh5_0),.din(w_dff_A_wvFR0Uve3_0),.clk(gclk));
	jdff dff_A_JgJPasJh5_0(.dout(w_dff_A_N6lR6jMC6_0),.din(w_dff_A_JgJPasJh5_0),.clk(gclk));
	jdff dff_A_N6lR6jMC6_0(.dout(w_dff_A_hhYbkQx20_0),.din(w_dff_A_N6lR6jMC6_0),.clk(gclk));
	jdff dff_A_hhYbkQx20_0(.dout(w_dff_A_wKjpYrWy5_0),.din(w_dff_A_hhYbkQx20_0),.clk(gclk));
	jdff dff_A_wKjpYrWy5_0(.dout(w_dff_A_ZeZ8qDSk1_0),.din(w_dff_A_wKjpYrWy5_0),.clk(gclk));
	jdff dff_A_ZeZ8qDSk1_0(.dout(w_dff_A_J2mufkAo7_0),.din(w_dff_A_ZeZ8qDSk1_0),.clk(gclk));
	jdff dff_A_J2mufkAo7_0(.dout(w_dff_A_dB4bUQiS8_0),.din(w_dff_A_J2mufkAo7_0),.clk(gclk));
	jdff dff_A_dB4bUQiS8_0(.dout(w_dff_A_JnsKETaU9_0),.din(w_dff_A_dB4bUQiS8_0),.clk(gclk));
	jdff dff_A_JnsKETaU9_0(.dout(w_dff_A_PXMtGslz3_0),.din(w_dff_A_JnsKETaU9_0),.clk(gclk));
	jdff dff_A_PXMtGslz3_0(.dout(f37),.din(w_dff_A_PXMtGslz3_0),.clk(gclk));
	jdff dff_A_4Rn8acWn9_2(.dout(w_dff_A_9ym0hURn8_0),.din(w_dff_A_4Rn8acWn9_2),.clk(gclk));
	jdff dff_A_9ym0hURn8_0(.dout(w_dff_A_yvKFYDyW6_0),.din(w_dff_A_9ym0hURn8_0),.clk(gclk));
	jdff dff_A_yvKFYDyW6_0(.dout(w_dff_A_rB3bBYAo8_0),.din(w_dff_A_yvKFYDyW6_0),.clk(gclk));
	jdff dff_A_rB3bBYAo8_0(.dout(w_dff_A_oPNcd0GF2_0),.din(w_dff_A_rB3bBYAo8_0),.clk(gclk));
	jdff dff_A_oPNcd0GF2_0(.dout(w_dff_A_NGB2M9Hx0_0),.din(w_dff_A_oPNcd0GF2_0),.clk(gclk));
	jdff dff_A_NGB2M9Hx0_0(.dout(w_dff_A_WbLPtOR91_0),.din(w_dff_A_NGB2M9Hx0_0),.clk(gclk));
	jdff dff_A_WbLPtOR91_0(.dout(w_dff_A_Tan51rf57_0),.din(w_dff_A_WbLPtOR91_0),.clk(gclk));
	jdff dff_A_Tan51rf57_0(.dout(w_dff_A_9LDDF9eD7_0),.din(w_dff_A_Tan51rf57_0),.clk(gclk));
	jdff dff_A_9LDDF9eD7_0(.dout(w_dff_A_oZC6NZOM0_0),.din(w_dff_A_9LDDF9eD7_0),.clk(gclk));
	jdff dff_A_oZC6NZOM0_0(.dout(w_dff_A_K9CinZsf7_0),.din(w_dff_A_oZC6NZOM0_0),.clk(gclk));
	jdff dff_A_K9CinZsf7_0(.dout(w_dff_A_DSjOBXel1_0),.din(w_dff_A_K9CinZsf7_0),.clk(gclk));
	jdff dff_A_DSjOBXel1_0(.dout(w_dff_A_ycxBJLah5_0),.din(w_dff_A_DSjOBXel1_0),.clk(gclk));
	jdff dff_A_ycxBJLah5_0(.dout(w_dff_A_wxiRA0pH7_0),.din(w_dff_A_ycxBJLah5_0),.clk(gclk));
	jdff dff_A_wxiRA0pH7_0(.dout(w_dff_A_mrlzsnng6_0),.din(w_dff_A_wxiRA0pH7_0),.clk(gclk));
	jdff dff_A_mrlzsnng6_0(.dout(w_dff_A_eTtNNSoP9_0),.din(w_dff_A_mrlzsnng6_0),.clk(gclk));
	jdff dff_A_eTtNNSoP9_0(.dout(w_dff_A_XsOaRDLz0_0),.din(w_dff_A_eTtNNSoP9_0),.clk(gclk));
	jdff dff_A_XsOaRDLz0_0(.dout(w_dff_A_vJWiNudq2_0),.din(w_dff_A_XsOaRDLz0_0),.clk(gclk));
	jdff dff_A_vJWiNudq2_0(.dout(w_dff_A_LS9J4qHz0_0),.din(w_dff_A_vJWiNudq2_0),.clk(gclk));
	jdff dff_A_LS9J4qHz0_0(.dout(w_dff_A_kakepyhG6_0),.din(w_dff_A_LS9J4qHz0_0),.clk(gclk));
	jdff dff_A_kakepyhG6_0(.dout(w_dff_A_gO8O1W7W3_0),.din(w_dff_A_kakepyhG6_0),.clk(gclk));
	jdff dff_A_gO8O1W7W3_0(.dout(w_dff_A_gVSjW9hB3_0),.din(w_dff_A_gO8O1W7W3_0),.clk(gclk));
	jdff dff_A_gVSjW9hB3_0(.dout(w_dff_A_tLv7LdDn5_0),.din(w_dff_A_gVSjW9hB3_0),.clk(gclk));
	jdff dff_A_tLv7LdDn5_0(.dout(w_dff_A_kDbAWkJD9_0),.din(w_dff_A_tLv7LdDn5_0),.clk(gclk));
	jdff dff_A_kDbAWkJD9_0(.dout(w_dff_A_VVQFFhE27_0),.din(w_dff_A_kDbAWkJD9_0),.clk(gclk));
	jdff dff_A_VVQFFhE27_0(.dout(w_dff_A_Q6keX4yH6_0),.din(w_dff_A_VVQFFhE27_0),.clk(gclk));
	jdff dff_A_Q6keX4yH6_0(.dout(w_dff_A_QxCZyVeY1_0),.din(w_dff_A_Q6keX4yH6_0),.clk(gclk));
	jdff dff_A_QxCZyVeY1_0(.dout(w_dff_A_pYp2jd4T7_0),.din(w_dff_A_QxCZyVeY1_0),.clk(gclk));
	jdff dff_A_pYp2jd4T7_0(.dout(w_dff_A_gefk1dwu5_0),.din(w_dff_A_pYp2jd4T7_0),.clk(gclk));
	jdff dff_A_gefk1dwu5_0(.dout(w_dff_A_mDn3iTYk4_0),.din(w_dff_A_gefk1dwu5_0),.clk(gclk));
	jdff dff_A_mDn3iTYk4_0(.dout(w_dff_A_vqwfpaBb5_0),.din(w_dff_A_mDn3iTYk4_0),.clk(gclk));
	jdff dff_A_vqwfpaBb5_0(.dout(w_dff_A_Y56fIn5Q0_0),.din(w_dff_A_vqwfpaBb5_0),.clk(gclk));
	jdff dff_A_Y56fIn5Q0_0(.dout(w_dff_A_2T2wMx4o9_0),.din(w_dff_A_Y56fIn5Q0_0),.clk(gclk));
	jdff dff_A_2T2wMx4o9_0(.dout(w_dff_A_X156pY411_0),.din(w_dff_A_2T2wMx4o9_0),.clk(gclk));
	jdff dff_A_X156pY411_0(.dout(w_dff_A_dgAWoQu22_0),.din(w_dff_A_X156pY411_0),.clk(gclk));
	jdff dff_A_dgAWoQu22_0(.dout(w_dff_A_n9Uuorpr4_0),.din(w_dff_A_dgAWoQu22_0),.clk(gclk));
	jdff dff_A_n9Uuorpr4_0(.dout(w_dff_A_JKTKpB1N1_0),.din(w_dff_A_n9Uuorpr4_0),.clk(gclk));
	jdff dff_A_JKTKpB1N1_0(.dout(w_dff_A_K3aRhSSR0_0),.din(w_dff_A_JKTKpB1N1_0),.clk(gclk));
	jdff dff_A_K3aRhSSR0_0(.dout(w_dff_A_NoKsbhUR5_0),.din(w_dff_A_K3aRhSSR0_0),.clk(gclk));
	jdff dff_A_NoKsbhUR5_0(.dout(w_dff_A_xenreQ6W3_0),.din(w_dff_A_NoKsbhUR5_0),.clk(gclk));
	jdff dff_A_xenreQ6W3_0(.dout(w_dff_A_vQwwAsJD1_0),.din(w_dff_A_xenreQ6W3_0),.clk(gclk));
	jdff dff_A_vQwwAsJD1_0(.dout(w_dff_A_SU4m2x337_0),.din(w_dff_A_vQwwAsJD1_0),.clk(gclk));
	jdff dff_A_SU4m2x337_0(.dout(w_dff_A_1PygVFLS0_0),.din(w_dff_A_SU4m2x337_0),.clk(gclk));
	jdff dff_A_1PygVFLS0_0(.dout(w_dff_A_pF3xXOZR0_0),.din(w_dff_A_1PygVFLS0_0),.clk(gclk));
	jdff dff_A_pF3xXOZR0_0(.dout(w_dff_A_EiAoH38c6_0),.din(w_dff_A_pF3xXOZR0_0),.clk(gclk));
	jdff dff_A_EiAoH38c6_0(.dout(w_dff_A_IiF9nW1Z6_0),.din(w_dff_A_EiAoH38c6_0),.clk(gclk));
	jdff dff_A_IiF9nW1Z6_0(.dout(w_dff_A_jWIFUvVH0_0),.din(w_dff_A_IiF9nW1Z6_0),.clk(gclk));
	jdff dff_A_jWIFUvVH0_0(.dout(w_dff_A_JrEEMHtX9_0),.din(w_dff_A_jWIFUvVH0_0),.clk(gclk));
	jdff dff_A_JrEEMHtX9_0(.dout(w_dff_A_0H0kz2tT0_0),.din(w_dff_A_JrEEMHtX9_0),.clk(gclk));
	jdff dff_A_0H0kz2tT0_0(.dout(w_dff_A_6FBUCSAl3_0),.din(w_dff_A_0H0kz2tT0_0),.clk(gclk));
	jdff dff_A_6FBUCSAl3_0(.dout(w_dff_A_r3JLqB512_0),.din(w_dff_A_6FBUCSAl3_0),.clk(gclk));
	jdff dff_A_r3JLqB512_0(.dout(w_dff_A_l4bRaizl6_0),.din(w_dff_A_r3JLqB512_0),.clk(gclk));
	jdff dff_A_l4bRaizl6_0(.dout(w_dff_A_zJMehraY4_0),.din(w_dff_A_l4bRaizl6_0),.clk(gclk));
	jdff dff_A_zJMehraY4_0(.dout(w_dff_A_SRFL3jk26_0),.din(w_dff_A_zJMehraY4_0),.clk(gclk));
	jdff dff_A_SRFL3jk26_0(.dout(w_dff_A_quz5vkU68_0),.din(w_dff_A_SRFL3jk26_0),.clk(gclk));
	jdff dff_A_quz5vkU68_0(.dout(w_dff_A_j5hplv7a5_0),.din(w_dff_A_quz5vkU68_0),.clk(gclk));
	jdff dff_A_j5hplv7a5_0(.dout(w_dff_A_dLDI33Zv4_0),.din(w_dff_A_j5hplv7a5_0),.clk(gclk));
	jdff dff_A_dLDI33Zv4_0(.dout(w_dff_A_YOUNvOLs8_0),.din(w_dff_A_dLDI33Zv4_0),.clk(gclk));
	jdff dff_A_YOUNvOLs8_0(.dout(w_dff_A_sjtAweMc6_0),.din(w_dff_A_YOUNvOLs8_0),.clk(gclk));
	jdff dff_A_sjtAweMc6_0(.dout(w_dff_A_M2WtbFEk0_0),.din(w_dff_A_sjtAweMc6_0),.clk(gclk));
	jdff dff_A_M2WtbFEk0_0(.dout(w_dff_A_uMYP7TBh0_0),.din(w_dff_A_M2WtbFEk0_0),.clk(gclk));
	jdff dff_A_uMYP7TBh0_0(.dout(w_dff_A_75g1qZ7J7_0),.din(w_dff_A_uMYP7TBh0_0),.clk(gclk));
	jdff dff_A_75g1qZ7J7_0(.dout(w_dff_A_weRWmR114_0),.din(w_dff_A_75g1qZ7J7_0),.clk(gclk));
	jdff dff_A_weRWmR114_0(.dout(w_dff_A_tLhWpRaf3_0),.din(w_dff_A_weRWmR114_0),.clk(gclk));
	jdff dff_A_tLhWpRaf3_0(.dout(w_dff_A_CpyKdXUj2_0),.din(w_dff_A_tLhWpRaf3_0),.clk(gclk));
	jdff dff_A_CpyKdXUj2_0(.dout(w_dff_A_3n6zaMjq7_0),.din(w_dff_A_CpyKdXUj2_0),.clk(gclk));
	jdff dff_A_3n6zaMjq7_0(.dout(w_dff_A_OeMeC6hR8_0),.din(w_dff_A_3n6zaMjq7_0),.clk(gclk));
	jdff dff_A_OeMeC6hR8_0(.dout(w_dff_A_VVtjRuJU5_0),.din(w_dff_A_OeMeC6hR8_0),.clk(gclk));
	jdff dff_A_VVtjRuJU5_0(.dout(w_dff_A_jt50o2VL2_0),.din(w_dff_A_VVtjRuJU5_0),.clk(gclk));
	jdff dff_A_jt50o2VL2_0(.dout(w_dff_A_arD3n7N57_0),.din(w_dff_A_jt50o2VL2_0),.clk(gclk));
	jdff dff_A_arD3n7N57_0(.dout(w_dff_A_KkJXCeBg6_0),.din(w_dff_A_arD3n7N57_0),.clk(gclk));
	jdff dff_A_KkJXCeBg6_0(.dout(w_dff_A_CwQrxJiv6_0),.din(w_dff_A_KkJXCeBg6_0),.clk(gclk));
	jdff dff_A_CwQrxJiv6_0(.dout(w_dff_A_m6Z1D3HT6_0),.din(w_dff_A_CwQrxJiv6_0),.clk(gclk));
	jdff dff_A_m6Z1D3HT6_0(.dout(w_dff_A_KPaFgBGL2_0),.din(w_dff_A_m6Z1D3HT6_0),.clk(gclk));
	jdff dff_A_KPaFgBGL2_0(.dout(w_dff_A_jpVJqQs63_0),.din(w_dff_A_KPaFgBGL2_0),.clk(gclk));
	jdff dff_A_jpVJqQs63_0(.dout(w_dff_A_gLpbDhbH4_0),.din(w_dff_A_jpVJqQs63_0),.clk(gclk));
	jdff dff_A_gLpbDhbH4_0(.dout(w_dff_A_x7EIawcx8_0),.din(w_dff_A_gLpbDhbH4_0),.clk(gclk));
	jdff dff_A_x7EIawcx8_0(.dout(w_dff_A_RHxXTx2I8_0),.din(w_dff_A_x7EIawcx8_0),.clk(gclk));
	jdff dff_A_RHxXTx2I8_0(.dout(w_dff_A_0nPt8unl8_0),.din(w_dff_A_RHxXTx2I8_0),.clk(gclk));
	jdff dff_A_0nPt8unl8_0(.dout(w_dff_A_pH3EjJnN6_0),.din(w_dff_A_0nPt8unl8_0),.clk(gclk));
	jdff dff_A_pH3EjJnN6_0(.dout(w_dff_A_459ve60a5_0),.din(w_dff_A_pH3EjJnN6_0),.clk(gclk));
	jdff dff_A_459ve60a5_0(.dout(w_dff_A_UGa98vKo1_0),.din(w_dff_A_459ve60a5_0),.clk(gclk));
	jdff dff_A_UGa98vKo1_0(.dout(w_dff_A_mbKVm1rI9_0),.din(w_dff_A_UGa98vKo1_0),.clk(gclk));
	jdff dff_A_mbKVm1rI9_0(.dout(w_dff_A_I10fOUxm7_0),.din(w_dff_A_mbKVm1rI9_0),.clk(gclk));
	jdff dff_A_I10fOUxm7_0(.dout(w_dff_A_zmyJ6ohw2_0),.din(w_dff_A_I10fOUxm7_0),.clk(gclk));
	jdff dff_A_zmyJ6ohw2_0(.dout(w_dff_A_ulqR7j5G3_0),.din(w_dff_A_zmyJ6ohw2_0),.clk(gclk));
	jdff dff_A_ulqR7j5G3_0(.dout(w_dff_A_5NYrJ0xk2_0),.din(w_dff_A_ulqR7j5G3_0),.clk(gclk));
	jdff dff_A_5NYrJ0xk2_0(.dout(w_dff_A_7qSoFryb6_0),.din(w_dff_A_5NYrJ0xk2_0),.clk(gclk));
	jdff dff_A_7qSoFryb6_0(.dout(w_dff_A_fi0uRMCN2_0),.din(w_dff_A_7qSoFryb6_0),.clk(gclk));
	jdff dff_A_fi0uRMCN2_0(.dout(f38),.din(w_dff_A_fi0uRMCN2_0),.clk(gclk));
	jdff dff_A_f746W3Pr1_2(.dout(w_dff_A_E1Mfhl4N4_0),.din(w_dff_A_f746W3Pr1_2),.clk(gclk));
	jdff dff_A_E1Mfhl4N4_0(.dout(w_dff_A_nAJmMpoC7_0),.din(w_dff_A_E1Mfhl4N4_0),.clk(gclk));
	jdff dff_A_nAJmMpoC7_0(.dout(w_dff_A_2IQuxUlC9_0),.din(w_dff_A_nAJmMpoC7_0),.clk(gclk));
	jdff dff_A_2IQuxUlC9_0(.dout(w_dff_A_GFnFqxHF0_0),.din(w_dff_A_2IQuxUlC9_0),.clk(gclk));
	jdff dff_A_GFnFqxHF0_0(.dout(w_dff_A_HZzxVe5R7_0),.din(w_dff_A_GFnFqxHF0_0),.clk(gclk));
	jdff dff_A_HZzxVe5R7_0(.dout(w_dff_A_xIPXtjfh6_0),.din(w_dff_A_HZzxVe5R7_0),.clk(gclk));
	jdff dff_A_xIPXtjfh6_0(.dout(w_dff_A_RXBPeT6X3_0),.din(w_dff_A_xIPXtjfh6_0),.clk(gclk));
	jdff dff_A_RXBPeT6X3_0(.dout(w_dff_A_FspnMCwp2_0),.din(w_dff_A_RXBPeT6X3_0),.clk(gclk));
	jdff dff_A_FspnMCwp2_0(.dout(w_dff_A_Gxfb6Dm70_0),.din(w_dff_A_FspnMCwp2_0),.clk(gclk));
	jdff dff_A_Gxfb6Dm70_0(.dout(w_dff_A_PyzkpODJ4_0),.din(w_dff_A_Gxfb6Dm70_0),.clk(gclk));
	jdff dff_A_PyzkpODJ4_0(.dout(w_dff_A_zMxAzMzW4_0),.din(w_dff_A_PyzkpODJ4_0),.clk(gclk));
	jdff dff_A_zMxAzMzW4_0(.dout(w_dff_A_N89C6uF51_0),.din(w_dff_A_zMxAzMzW4_0),.clk(gclk));
	jdff dff_A_N89C6uF51_0(.dout(w_dff_A_U2YbtVln0_0),.din(w_dff_A_N89C6uF51_0),.clk(gclk));
	jdff dff_A_U2YbtVln0_0(.dout(w_dff_A_LTjzwddC6_0),.din(w_dff_A_U2YbtVln0_0),.clk(gclk));
	jdff dff_A_LTjzwddC6_0(.dout(w_dff_A_s7wbO6Lb9_0),.din(w_dff_A_LTjzwddC6_0),.clk(gclk));
	jdff dff_A_s7wbO6Lb9_0(.dout(w_dff_A_RsstR8tj8_0),.din(w_dff_A_s7wbO6Lb9_0),.clk(gclk));
	jdff dff_A_RsstR8tj8_0(.dout(w_dff_A_H2ew9FRo0_0),.din(w_dff_A_RsstR8tj8_0),.clk(gclk));
	jdff dff_A_H2ew9FRo0_0(.dout(w_dff_A_5lX0hUKw1_0),.din(w_dff_A_H2ew9FRo0_0),.clk(gclk));
	jdff dff_A_5lX0hUKw1_0(.dout(w_dff_A_cyLsIclr2_0),.din(w_dff_A_5lX0hUKw1_0),.clk(gclk));
	jdff dff_A_cyLsIclr2_0(.dout(w_dff_A_JhO5zw7r0_0),.din(w_dff_A_cyLsIclr2_0),.clk(gclk));
	jdff dff_A_JhO5zw7r0_0(.dout(w_dff_A_Uy8oZC2A1_0),.din(w_dff_A_JhO5zw7r0_0),.clk(gclk));
	jdff dff_A_Uy8oZC2A1_0(.dout(w_dff_A_kgBQQ83n1_0),.din(w_dff_A_Uy8oZC2A1_0),.clk(gclk));
	jdff dff_A_kgBQQ83n1_0(.dout(w_dff_A_r8NL11tE5_0),.din(w_dff_A_kgBQQ83n1_0),.clk(gclk));
	jdff dff_A_r8NL11tE5_0(.dout(w_dff_A_8dAtUHwX9_0),.din(w_dff_A_r8NL11tE5_0),.clk(gclk));
	jdff dff_A_8dAtUHwX9_0(.dout(w_dff_A_p51L4Dw08_0),.din(w_dff_A_8dAtUHwX9_0),.clk(gclk));
	jdff dff_A_p51L4Dw08_0(.dout(w_dff_A_cH12S2Tx8_0),.din(w_dff_A_p51L4Dw08_0),.clk(gclk));
	jdff dff_A_cH12S2Tx8_0(.dout(w_dff_A_Y3Kn1imC6_0),.din(w_dff_A_cH12S2Tx8_0),.clk(gclk));
	jdff dff_A_Y3Kn1imC6_0(.dout(w_dff_A_3RkeztCx5_0),.din(w_dff_A_Y3Kn1imC6_0),.clk(gclk));
	jdff dff_A_3RkeztCx5_0(.dout(w_dff_A_wdQkdX3V4_0),.din(w_dff_A_3RkeztCx5_0),.clk(gclk));
	jdff dff_A_wdQkdX3V4_0(.dout(w_dff_A_Jnch4fUi1_0),.din(w_dff_A_wdQkdX3V4_0),.clk(gclk));
	jdff dff_A_Jnch4fUi1_0(.dout(w_dff_A_z6PWRfF86_0),.din(w_dff_A_Jnch4fUi1_0),.clk(gclk));
	jdff dff_A_z6PWRfF86_0(.dout(w_dff_A_EwKBplcw3_0),.din(w_dff_A_z6PWRfF86_0),.clk(gclk));
	jdff dff_A_EwKBplcw3_0(.dout(w_dff_A_l9ADmwb05_0),.din(w_dff_A_EwKBplcw3_0),.clk(gclk));
	jdff dff_A_l9ADmwb05_0(.dout(w_dff_A_AFILsLV16_0),.din(w_dff_A_l9ADmwb05_0),.clk(gclk));
	jdff dff_A_AFILsLV16_0(.dout(w_dff_A_fqef3RN83_0),.din(w_dff_A_AFILsLV16_0),.clk(gclk));
	jdff dff_A_fqef3RN83_0(.dout(w_dff_A_0NBBSGke1_0),.din(w_dff_A_fqef3RN83_0),.clk(gclk));
	jdff dff_A_0NBBSGke1_0(.dout(w_dff_A_epF3FsQ92_0),.din(w_dff_A_0NBBSGke1_0),.clk(gclk));
	jdff dff_A_epF3FsQ92_0(.dout(w_dff_A_RoRATiEh5_0),.din(w_dff_A_epF3FsQ92_0),.clk(gclk));
	jdff dff_A_RoRATiEh5_0(.dout(w_dff_A_1VL2fA4n8_0),.din(w_dff_A_RoRATiEh5_0),.clk(gclk));
	jdff dff_A_1VL2fA4n8_0(.dout(w_dff_A_pkrC71cH4_0),.din(w_dff_A_1VL2fA4n8_0),.clk(gclk));
	jdff dff_A_pkrC71cH4_0(.dout(w_dff_A_rl4ed3tV0_0),.din(w_dff_A_pkrC71cH4_0),.clk(gclk));
	jdff dff_A_rl4ed3tV0_0(.dout(w_dff_A_nzrpFkXX7_0),.din(w_dff_A_rl4ed3tV0_0),.clk(gclk));
	jdff dff_A_nzrpFkXX7_0(.dout(w_dff_A_1h4k5g802_0),.din(w_dff_A_nzrpFkXX7_0),.clk(gclk));
	jdff dff_A_1h4k5g802_0(.dout(w_dff_A_hPVc5LxE5_0),.din(w_dff_A_1h4k5g802_0),.clk(gclk));
	jdff dff_A_hPVc5LxE5_0(.dout(w_dff_A_CxjkIRIS8_0),.din(w_dff_A_hPVc5LxE5_0),.clk(gclk));
	jdff dff_A_CxjkIRIS8_0(.dout(w_dff_A_yC9zI7aD6_0),.din(w_dff_A_CxjkIRIS8_0),.clk(gclk));
	jdff dff_A_yC9zI7aD6_0(.dout(w_dff_A_Z8kFUtuq4_0),.din(w_dff_A_yC9zI7aD6_0),.clk(gclk));
	jdff dff_A_Z8kFUtuq4_0(.dout(w_dff_A_c8DXcmZi7_0),.din(w_dff_A_Z8kFUtuq4_0),.clk(gclk));
	jdff dff_A_c8DXcmZi7_0(.dout(w_dff_A_wdUWkAd01_0),.din(w_dff_A_c8DXcmZi7_0),.clk(gclk));
	jdff dff_A_wdUWkAd01_0(.dout(w_dff_A_0sYeAFDC2_0),.din(w_dff_A_wdUWkAd01_0),.clk(gclk));
	jdff dff_A_0sYeAFDC2_0(.dout(w_dff_A_ckcRrgRj0_0),.din(w_dff_A_0sYeAFDC2_0),.clk(gclk));
	jdff dff_A_ckcRrgRj0_0(.dout(w_dff_A_t9wIPvBX3_0),.din(w_dff_A_ckcRrgRj0_0),.clk(gclk));
	jdff dff_A_t9wIPvBX3_0(.dout(w_dff_A_Kabk8kkV2_0),.din(w_dff_A_t9wIPvBX3_0),.clk(gclk));
	jdff dff_A_Kabk8kkV2_0(.dout(w_dff_A_gpdwEzTC9_0),.din(w_dff_A_Kabk8kkV2_0),.clk(gclk));
	jdff dff_A_gpdwEzTC9_0(.dout(w_dff_A_D4QrJoqY0_0),.din(w_dff_A_gpdwEzTC9_0),.clk(gclk));
	jdff dff_A_D4QrJoqY0_0(.dout(w_dff_A_w2rtCkcZ5_0),.din(w_dff_A_D4QrJoqY0_0),.clk(gclk));
	jdff dff_A_w2rtCkcZ5_0(.dout(w_dff_A_NnX9lT930_0),.din(w_dff_A_w2rtCkcZ5_0),.clk(gclk));
	jdff dff_A_NnX9lT930_0(.dout(w_dff_A_S1DvLhHm1_0),.din(w_dff_A_NnX9lT930_0),.clk(gclk));
	jdff dff_A_S1DvLhHm1_0(.dout(w_dff_A_iEoEVDmH4_0),.din(w_dff_A_S1DvLhHm1_0),.clk(gclk));
	jdff dff_A_iEoEVDmH4_0(.dout(w_dff_A_7gGC4gM24_0),.din(w_dff_A_iEoEVDmH4_0),.clk(gclk));
	jdff dff_A_7gGC4gM24_0(.dout(w_dff_A_kqH80jDy3_0),.din(w_dff_A_7gGC4gM24_0),.clk(gclk));
	jdff dff_A_kqH80jDy3_0(.dout(w_dff_A_UPhesf4B9_0),.din(w_dff_A_kqH80jDy3_0),.clk(gclk));
	jdff dff_A_UPhesf4B9_0(.dout(w_dff_A_oppNHXX38_0),.din(w_dff_A_UPhesf4B9_0),.clk(gclk));
	jdff dff_A_oppNHXX38_0(.dout(w_dff_A_aWjCQfwP4_0),.din(w_dff_A_oppNHXX38_0),.clk(gclk));
	jdff dff_A_aWjCQfwP4_0(.dout(w_dff_A_bsVY1f6c5_0),.din(w_dff_A_aWjCQfwP4_0),.clk(gclk));
	jdff dff_A_bsVY1f6c5_0(.dout(w_dff_A_qOnrAXDp1_0),.din(w_dff_A_bsVY1f6c5_0),.clk(gclk));
	jdff dff_A_qOnrAXDp1_0(.dout(w_dff_A_591tFOw36_0),.din(w_dff_A_qOnrAXDp1_0),.clk(gclk));
	jdff dff_A_591tFOw36_0(.dout(w_dff_A_9sf7j4QP6_0),.din(w_dff_A_591tFOw36_0),.clk(gclk));
	jdff dff_A_9sf7j4QP6_0(.dout(w_dff_A_sjwMV4JZ0_0),.din(w_dff_A_9sf7j4QP6_0),.clk(gclk));
	jdff dff_A_sjwMV4JZ0_0(.dout(w_dff_A_NK0Uaf4n7_0),.din(w_dff_A_sjwMV4JZ0_0),.clk(gclk));
	jdff dff_A_NK0Uaf4n7_0(.dout(w_dff_A_OGGO79F78_0),.din(w_dff_A_NK0Uaf4n7_0),.clk(gclk));
	jdff dff_A_OGGO79F78_0(.dout(w_dff_A_8pWyg9LJ3_0),.din(w_dff_A_OGGO79F78_0),.clk(gclk));
	jdff dff_A_8pWyg9LJ3_0(.dout(w_dff_A_1BWoCeRx2_0),.din(w_dff_A_8pWyg9LJ3_0),.clk(gclk));
	jdff dff_A_1BWoCeRx2_0(.dout(w_dff_A_ZSsTMc9r7_0),.din(w_dff_A_1BWoCeRx2_0),.clk(gclk));
	jdff dff_A_ZSsTMc9r7_0(.dout(w_dff_A_1acBxVBM3_0),.din(w_dff_A_ZSsTMc9r7_0),.clk(gclk));
	jdff dff_A_1acBxVBM3_0(.dout(w_dff_A_aFoE6i4s8_0),.din(w_dff_A_1acBxVBM3_0),.clk(gclk));
	jdff dff_A_aFoE6i4s8_0(.dout(w_dff_A_k9hEVnLb9_0),.din(w_dff_A_aFoE6i4s8_0),.clk(gclk));
	jdff dff_A_k9hEVnLb9_0(.dout(w_dff_A_p1Bx8YHV3_0),.din(w_dff_A_k9hEVnLb9_0),.clk(gclk));
	jdff dff_A_p1Bx8YHV3_0(.dout(w_dff_A_mWnRbqn53_0),.din(w_dff_A_p1Bx8YHV3_0),.clk(gclk));
	jdff dff_A_mWnRbqn53_0(.dout(w_dff_A_HeGKQYiV1_0),.din(w_dff_A_mWnRbqn53_0),.clk(gclk));
	jdff dff_A_HeGKQYiV1_0(.dout(w_dff_A_jJQY80bG2_0),.din(w_dff_A_HeGKQYiV1_0),.clk(gclk));
	jdff dff_A_jJQY80bG2_0(.dout(w_dff_A_2VATXkln2_0),.din(w_dff_A_jJQY80bG2_0),.clk(gclk));
	jdff dff_A_2VATXkln2_0(.dout(w_dff_A_V24kuI7C0_0),.din(w_dff_A_2VATXkln2_0),.clk(gclk));
	jdff dff_A_V24kuI7C0_0(.dout(w_dff_A_ZAAuTILi3_0),.din(w_dff_A_V24kuI7C0_0),.clk(gclk));
	jdff dff_A_ZAAuTILi3_0(.dout(w_dff_A_mpexeJvC7_0),.din(w_dff_A_ZAAuTILi3_0),.clk(gclk));
	jdff dff_A_mpexeJvC7_0(.dout(w_dff_A_XgAcfQmd8_0),.din(w_dff_A_mpexeJvC7_0),.clk(gclk));
	jdff dff_A_XgAcfQmd8_0(.dout(w_dff_A_if8icmPh1_0),.din(w_dff_A_XgAcfQmd8_0),.clk(gclk));
	jdff dff_A_if8icmPh1_0(.dout(f39),.din(w_dff_A_if8icmPh1_0),.clk(gclk));
	jdff dff_A_m6wDD8ja6_2(.dout(w_dff_A_BHl71OzP6_0),.din(w_dff_A_m6wDD8ja6_2),.clk(gclk));
	jdff dff_A_BHl71OzP6_0(.dout(w_dff_A_S4GDVtfe7_0),.din(w_dff_A_BHl71OzP6_0),.clk(gclk));
	jdff dff_A_S4GDVtfe7_0(.dout(w_dff_A_cRmTUQN44_0),.din(w_dff_A_S4GDVtfe7_0),.clk(gclk));
	jdff dff_A_cRmTUQN44_0(.dout(w_dff_A_uWQhdzul9_0),.din(w_dff_A_cRmTUQN44_0),.clk(gclk));
	jdff dff_A_uWQhdzul9_0(.dout(w_dff_A_a5vYoFVz5_0),.din(w_dff_A_uWQhdzul9_0),.clk(gclk));
	jdff dff_A_a5vYoFVz5_0(.dout(w_dff_A_rnPYtGdE9_0),.din(w_dff_A_a5vYoFVz5_0),.clk(gclk));
	jdff dff_A_rnPYtGdE9_0(.dout(w_dff_A_NLeXx2aM6_0),.din(w_dff_A_rnPYtGdE9_0),.clk(gclk));
	jdff dff_A_NLeXx2aM6_0(.dout(w_dff_A_MB8CsnD64_0),.din(w_dff_A_NLeXx2aM6_0),.clk(gclk));
	jdff dff_A_MB8CsnD64_0(.dout(w_dff_A_o9waanZ98_0),.din(w_dff_A_MB8CsnD64_0),.clk(gclk));
	jdff dff_A_o9waanZ98_0(.dout(w_dff_A_83Q7eVzm6_0),.din(w_dff_A_o9waanZ98_0),.clk(gclk));
	jdff dff_A_83Q7eVzm6_0(.dout(w_dff_A_MhHoKnEJ1_0),.din(w_dff_A_83Q7eVzm6_0),.clk(gclk));
	jdff dff_A_MhHoKnEJ1_0(.dout(w_dff_A_qZx5AP5s3_0),.din(w_dff_A_MhHoKnEJ1_0),.clk(gclk));
	jdff dff_A_qZx5AP5s3_0(.dout(w_dff_A_6gVuoz968_0),.din(w_dff_A_qZx5AP5s3_0),.clk(gclk));
	jdff dff_A_6gVuoz968_0(.dout(w_dff_A_clfWsd9i5_0),.din(w_dff_A_6gVuoz968_0),.clk(gclk));
	jdff dff_A_clfWsd9i5_0(.dout(w_dff_A_4IrE0puv3_0),.din(w_dff_A_clfWsd9i5_0),.clk(gclk));
	jdff dff_A_4IrE0puv3_0(.dout(w_dff_A_7yK4No5Y2_0),.din(w_dff_A_4IrE0puv3_0),.clk(gclk));
	jdff dff_A_7yK4No5Y2_0(.dout(w_dff_A_NNZst9LK6_0),.din(w_dff_A_7yK4No5Y2_0),.clk(gclk));
	jdff dff_A_NNZst9LK6_0(.dout(w_dff_A_fS440rFR4_0),.din(w_dff_A_NNZst9LK6_0),.clk(gclk));
	jdff dff_A_fS440rFR4_0(.dout(w_dff_A_2n9xBBUw3_0),.din(w_dff_A_fS440rFR4_0),.clk(gclk));
	jdff dff_A_2n9xBBUw3_0(.dout(w_dff_A_DgkeoheS6_0),.din(w_dff_A_2n9xBBUw3_0),.clk(gclk));
	jdff dff_A_DgkeoheS6_0(.dout(w_dff_A_ZONus89Q2_0),.din(w_dff_A_DgkeoheS6_0),.clk(gclk));
	jdff dff_A_ZONus89Q2_0(.dout(w_dff_A_RXs2uRQk6_0),.din(w_dff_A_ZONus89Q2_0),.clk(gclk));
	jdff dff_A_RXs2uRQk6_0(.dout(w_dff_A_iMfpHmTI1_0),.din(w_dff_A_RXs2uRQk6_0),.clk(gclk));
	jdff dff_A_iMfpHmTI1_0(.dout(w_dff_A_NGEBiC2z9_0),.din(w_dff_A_iMfpHmTI1_0),.clk(gclk));
	jdff dff_A_NGEBiC2z9_0(.dout(w_dff_A_XofUm5kU4_0),.din(w_dff_A_NGEBiC2z9_0),.clk(gclk));
	jdff dff_A_XofUm5kU4_0(.dout(w_dff_A_EQsX8gc47_0),.din(w_dff_A_XofUm5kU4_0),.clk(gclk));
	jdff dff_A_EQsX8gc47_0(.dout(w_dff_A_bX8uZ8OQ0_0),.din(w_dff_A_EQsX8gc47_0),.clk(gclk));
	jdff dff_A_bX8uZ8OQ0_0(.dout(w_dff_A_XthixKrH0_0),.din(w_dff_A_bX8uZ8OQ0_0),.clk(gclk));
	jdff dff_A_XthixKrH0_0(.dout(w_dff_A_mg4tjIf27_0),.din(w_dff_A_XthixKrH0_0),.clk(gclk));
	jdff dff_A_mg4tjIf27_0(.dout(w_dff_A_7CHxDIrY9_0),.din(w_dff_A_mg4tjIf27_0),.clk(gclk));
	jdff dff_A_7CHxDIrY9_0(.dout(w_dff_A_YJUfiYMX4_0),.din(w_dff_A_7CHxDIrY9_0),.clk(gclk));
	jdff dff_A_YJUfiYMX4_0(.dout(w_dff_A_MDdt7uyp0_0),.din(w_dff_A_YJUfiYMX4_0),.clk(gclk));
	jdff dff_A_MDdt7uyp0_0(.dout(w_dff_A_NoRviJwv3_0),.din(w_dff_A_MDdt7uyp0_0),.clk(gclk));
	jdff dff_A_NoRviJwv3_0(.dout(w_dff_A_bcLj5S4W0_0),.din(w_dff_A_NoRviJwv3_0),.clk(gclk));
	jdff dff_A_bcLj5S4W0_0(.dout(w_dff_A_iE0weS3a2_0),.din(w_dff_A_bcLj5S4W0_0),.clk(gclk));
	jdff dff_A_iE0weS3a2_0(.dout(w_dff_A_OPQnamKv6_0),.din(w_dff_A_iE0weS3a2_0),.clk(gclk));
	jdff dff_A_OPQnamKv6_0(.dout(w_dff_A_AAQLtQEV3_0),.din(w_dff_A_OPQnamKv6_0),.clk(gclk));
	jdff dff_A_AAQLtQEV3_0(.dout(w_dff_A_zoQbiNIp2_0),.din(w_dff_A_AAQLtQEV3_0),.clk(gclk));
	jdff dff_A_zoQbiNIp2_0(.dout(w_dff_A_QY7m5XD97_0),.din(w_dff_A_zoQbiNIp2_0),.clk(gclk));
	jdff dff_A_QY7m5XD97_0(.dout(w_dff_A_IltStdH92_0),.din(w_dff_A_QY7m5XD97_0),.clk(gclk));
	jdff dff_A_IltStdH92_0(.dout(w_dff_A_ZmXyIiqy5_0),.din(w_dff_A_IltStdH92_0),.clk(gclk));
	jdff dff_A_ZmXyIiqy5_0(.dout(w_dff_A_qZMfuUDk2_0),.din(w_dff_A_ZmXyIiqy5_0),.clk(gclk));
	jdff dff_A_qZMfuUDk2_0(.dout(w_dff_A_GsGgvVHS6_0),.din(w_dff_A_qZMfuUDk2_0),.clk(gclk));
	jdff dff_A_GsGgvVHS6_0(.dout(w_dff_A_wLewi5y66_0),.din(w_dff_A_GsGgvVHS6_0),.clk(gclk));
	jdff dff_A_wLewi5y66_0(.dout(w_dff_A_4PdaJDLe5_0),.din(w_dff_A_wLewi5y66_0),.clk(gclk));
	jdff dff_A_4PdaJDLe5_0(.dout(w_dff_A_CxMkWETV2_0),.din(w_dff_A_4PdaJDLe5_0),.clk(gclk));
	jdff dff_A_CxMkWETV2_0(.dout(w_dff_A_MNSEKAZY8_0),.din(w_dff_A_CxMkWETV2_0),.clk(gclk));
	jdff dff_A_MNSEKAZY8_0(.dout(w_dff_A_CIxn2oFn2_0),.din(w_dff_A_MNSEKAZY8_0),.clk(gclk));
	jdff dff_A_CIxn2oFn2_0(.dout(w_dff_A_sXMgN7PZ6_0),.din(w_dff_A_CIxn2oFn2_0),.clk(gclk));
	jdff dff_A_sXMgN7PZ6_0(.dout(w_dff_A_KwnQ1ZhS6_0),.din(w_dff_A_sXMgN7PZ6_0),.clk(gclk));
	jdff dff_A_KwnQ1ZhS6_0(.dout(w_dff_A_1MX8UB0b3_0),.din(w_dff_A_KwnQ1ZhS6_0),.clk(gclk));
	jdff dff_A_1MX8UB0b3_0(.dout(w_dff_A_PFFVTUPD0_0),.din(w_dff_A_1MX8UB0b3_0),.clk(gclk));
	jdff dff_A_PFFVTUPD0_0(.dout(w_dff_A_Rl1XKOgL6_0),.din(w_dff_A_PFFVTUPD0_0),.clk(gclk));
	jdff dff_A_Rl1XKOgL6_0(.dout(w_dff_A_G2ptjs5y9_0),.din(w_dff_A_Rl1XKOgL6_0),.clk(gclk));
	jdff dff_A_G2ptjs5y9_0(.dout(w_dff_A_m7hKvn1g7_0),.din(w_dff_A_G2ptjs5y9_0),.clk(gclk));
	jdff dff_A_m7hKvn1g7_0(.dout(w_dff_A_mKaa2Wjo9_0),.din(w_dff_A_m7hKvn1g7_0),.clk(gclk));
	jdff dff_A_mKaa2Wjo9_0(.dout(w_dff_A_iAXsZpMl6_0),.din(w_dff_A_mKaa2Wjo9_0),.clk(gclk));
	jdff dff_A_iAXsZpMl6_0(.dout(w_dff_A_oNiRWPRy6_0),.din(w_dff_A_iAXsZpMl6_0),.clk(gclk));
	jdff dff_A_oNiRWPRy6_0(.dout(w_dff_A_XiOtLwJA8_0),.din(w_dff_A_oNiRWPRy6_0),.clk(gclk));
	jdff dff_A_XiOtLwJA8_0(.dout(w_dff_A_w8IQmPQa7_0),.din(w_dff_A_XiOtLwJA8_0),.clk(gclk));
	jdff dff_A_w8IQmPQa7_0(.dout(w_dff_A_DoDLtp033_0),.din(w_dff_A_w8IQmPQa7_0),.clk(gclk));
	jdff dff_A_DoDLtp033_0(.dout(w_dff_A_ErMBmMqg0_0),.din(w_dff_A_DoDLtp033_0),.clk(gclk));
	jdff dff_A_ErMBmMqg0_0(.dout(w_dff_A_VtrilmPI6_0),.din(w_dff_A_ErMBmMqg0_0),.clk(gclk));
	jdff dff_A_VtrilmPI6_0(.dout(w_dff_A_nes9wCju9_0),.din(w_dff_A_VtrilmPI6_0),.clk(gclk));
	jdff dff_A_nes9wCju9_0(.dout(w_dff_A_aSF9Ppk55_0),.din(w_dff_A_nes9wCju9_0),.clk(gclk));
	jdff dff_A_aSF9Ppk55_0(.dout(w_dff_A_RfruNhaw6_0),.din(w_dff_A_aSF9Ppk55_0),.clk(gclk));
	jdff dff_A_RfruNhaw6_0(.dout(w_dff_A_9wL3LaY63_0),.din(w_dff_A_RfruNhaw6_0),.clk(gclk));
	jdff dff_A_9wL3LaY63_0(.dout(w_dff_A_ZIXCrHd76_0),.din(w_dff_A_9wL3LaY63_0),.clk(gclk));
	jdff dff_A_ZIXCrHd76_0(.dout(w_dff_A_5CPZt2DX2_0),.din(w_dff_A_ZIXCrHd76_0),.clk(gclk));
	jdff dff_A_5CPZt2DX2_0(.dout(w_dff_A_JjvqSUFo5_0),.din(w_dff_A_5CPZt2DX2_0),.clk(gclk));
	jdff dff_A_JjvqSUFo5_0(.dout(w_dff_A_ki65u2I14_0),.din(w_dff_A_JjvqSUFo5_0),.clk(gclk));
	jdff dff_A_ki65u2I14_0(.dout(w_dff_A_fMg8iQoO7_0),.din(w_dff_A_ki65u2I14_0),.clk(gclk));
	jdff dff_A_fMg8iQoO7_0(.dout(w_dff_A_Z7rjPR5j1_0),.din(w_dff_A_fMg8iQoO7_0),.clk(gclk));
	jdff dff_A_Z7rjPR5j1_0(.dout(w_dff_A_fUzznTMX5_0),.din(w_dff_A_Z7rjPR5j1_0),.clk(gclk));
	jdff dff_A_fUzznTMX5_0(.dout(w_dff_A_DKGdcBaW3_0),.din(w_dff_A_fUzznTMX5_0),.clk(gclk));
	jdff dff_A_DKGdcBaW3_0(.dout(w_dff_A_jEmefuQ65_0),.din(w_dff_A_DKGdcBaW3_0),.clk(gclk));
	jdff dff_A_jEmefuQ65_0(.dout(w_dff_A_DfENg6Lk5_0),.din(w_dff_A_jEmefuQ65_0),.clk(gclk));
	jdff dff_A_DfENg6Lk5_0(.dout(w_dff_A_GrHit8J09_0),.din(w_dff_A_DfENg6Lk5_0),.clk(gclk));
	jdff dff_A_GrHit8J09_0(.dout(w_dff_A_C22bGiM54_0),.din(w_dff_A_GrHit8J09_0),.clk(gclk));
	jdff dff_A_C22bGiM54_0(.dout(w_dff_A_wn6vPOZK6_0),.din(w_dff_A_C22bGiM54_0),.clk(gclk));
	jdff dff_A_wn6vPOZK6_0(.dout(w_dff_A_hioXIX2W7_0),.din(w_dff_A_wn6vPOZK6_0),.clk(gclk));
	jdff dff_A_hioXIX2W7_0(.dout(w_dff_A_TtlENguc7_0),.din(w_dff_A_hioXIX2W7_0),.clk(gclk));
	jdff dff_A_TtlENguc7_0(.dout(w_dff_A_S0rUy7ha6_0),.din(w_dff_A_TtlENguc7_0),.clk(gclk));
	jdff dff_A_S0rUy7ha6_0(.dout(w_dff_A_MARckjvl6_0),.din(w_dff_A_S0rUy7ha6_0),.clk(gclk));
	jdff dff_A_MARckjvl6_0(.dout(w_dff_A_Uie4O28Q1_0),.din(w_dff_A_MARckjvl6_0),.clk(gclk));
	jdff dff_A_Uie4O28Q1_0(.dout(w_dff_A_0pMDkLN33_0),.din(w_dff_A_Uie4O28Q1_0),.clk(gclk));
	jdff dff_A_0pMDkLN33_0(.dout(f40),.din(w_dff_A_0pMDkLN33_0),.clk(gclk));
	jdff dff_A_6JBK2nPW1_2(.dout(w_dff_A_Ig44NJbk9_0),.din(w_dff_A_6JBK2nPW1_2),.clk(gclk));
	jdff dff_A_Ig44NJbk9_0(.dout(w_dff_A_LRmVccAH5_0),.din(w_dff_A_Ig44NJbk9_0),.clk(gclk));
	jdff dff_A_LRmVccAH5_0(.dout(w_dff_A_Am39zBpf9_0),.din(w_dff_A_LRmVccAH5_0),.clk(gclk));
	jdff dff_A_Am39zBpf9_0(.dout(w_dff_A_q6bkMG3r5_0),.din(w_dff_A_Am39zBpf9_0),.clk(gclk));
	jdff dff_A_q6bkMG3r5_0(.dout(w_dff_A_ofzib6Ux9_0),.din(w_dff_A_q6bkMG3r5_0),.clk(gclk));
	jdff dff_A_ofzib6Ux9_0(.dout(w_dff_A_7zVHYnFG1_0),.din(w_dff_A_ofzib6Ux9_0),.clk(gclk));
	jdff dff_A_7zVHYnFG1_0(.dout(w_dff_A_9GPFFWsn2_0),.din(w_dff_A_7zVHYnFG1_0),.clk(gclk));
	jdff dff_A_9GPFFWsn2_0(.dout(w_dff_A_RwRYpOlV1_0),.din(w_dff_A_9GPFFWsn2_0),.clk(gclk));
	jdff dff_A_RwRYpOlV1_0(.dout(w_dff_A_eUeSG9P08_0),.din(w_dff_A_RwRYpOlV1_0),.clk(gclk));
	jdff dff_A_eUeSG9P08_0(.dout(w_dff_A_XahTCvEH2_0),.din(w_dff_A_eUeSG9P08_0),.clk(gclk));
	jdff dff_A_XahTCvEH2_0(.dout(w_dff_A_eElY7Vk07_0),.din(w_dff_A_XahTCvEH2_0),.clk(gclk));
	jdff dff_A_eElY7Vk07_0(.dout(w_dff_A_CFuzPRoq3_0),.din(w_dff_A_eElY7Vk07_0),.clk(gclk));
	jdff dff_A_CFuzPRoq3_0(.dout(w_dff_A_HCXVOM8T0_0),.din(w_dff_A_CFuzPRoq3_0),.clk(gclk));
	jdff dff_A_HCXVOM8T0_0(.dout(w_dff_A_dmlUJlRM8_0),.din(w_dff_A_HCXVOM8T0_0),.clk(gclk));
	jdff dff_A_dmlUJlRM8_0(.dout(w_dff_A_0BVAuxGp3_0),.din(w_dff_A_dmlUJlRM8_0),.clk(gclk));
	jdff dff_A_0BVAuxGp3_0(.dout(w_dff_A_9SlYBCUY1_0),.din(w_dff_A_0BVAuxGp3_0),.clk(gclk));
	jdff dff_A_9SlYBCUY1_0(.dout(w_dff_A_6E7u8WM83_0),.din(w_dff_A_9SlYBCUY1_0),.clk(gclk));
	jdff dff_A_6E7u8WM83_0(.dout(w_dff_A_GGuJuZlR5_0),.din(w_dff_A_6E7u8WM83_0),.clk(gclk));
	jdff dff_A_GGuJuZlR5_0(.dout(w_dff_A_MTP2Fc0D0_0),.din(w_dff_A_GGuJuZlR5_0),.clk(gclk));
	jdff dff_A_MTP2Fc0D0_0(.dout(w_dff_A_TzeoYon48_0),.din(w_dff_A_MTP2Fc0D0_0),.clk(gclk));
	jdff dff_A_TzeoYon48_0(.dout(w_dff_A_wVUOj4Hb5_0),.din(w_dff_A_TzeoYon48_0),.clk(gclk));
	jdff dff_A_wVUOj4Hb5_0(.dout(w_dff_A_bxlmQx078_0),.din(w_dff_A_wVUOj4Hb5_0),.clk(gclk));
	jdff dff_A_bxlmQx078_0(.dout(w_dff_A_0yjJIeKB8_0),.din(w_dff_A_bxlmQx078_0),.clk(gclk));
	jdff dff_A_0yjJIeKB8_0(.dout(w_dff_A_pIANq9rP9_0),.din(w_dff_A_0yjJIeKB8_0),.clk(gclk));
	jdff dff_A_pIANq9rP9_0(.dout(w_dff_A_vniFLQhn9_0),.din(w_dff_A_pIANq9rP9_0),.clk(gclk));
	jdff dff_A_vniFLQhn9_0(.dout(w_dff_A_HLNnf8aX0_0),.din(w_dff_A_vniFLQhn9_0),.clk(gclk));
	jdff dff_A_HLNnf8aX0_0(.dout(w_dff_A_SUcwoulU3_0),.din(w_dff_A_HLNnf8aX0_0),.clk(gclk));
	jdff dff_A_SUcwoulU3_0(.dout(w_dff_A_bzGrdG5L8_0),.din(w_dff_A_SUcwoulU3_0),.clk(gclk));
	jdff dff_A_bzGrdG5L8_0(.dout(w_dff_A_3trIzNcl2_0),.din(w_dff_A_bzGrdG5L8_0),.clk(gclk));
	jdff dff_A_3trIzNcl2_0(.dout(w_dff_A_6wlYvITz1_0),.din(w_dff_A_3trIzNcl2_0),.clk(gclk));
	jdff dff_A_6wlYvITz1_0(.dout(w_dff_A_RFj2KSND7_0),.din(w_dff_A_6wlYvITz1_0),.clk(gclk));
	jdff dff_A_RFj2KSND7_0(.dout(w_dff_A_aYNYGUpa4_0),.din(w_dff_A_RFj2KSND7_0),.clk(gclk));
	jdff dff_A_aYNYGUpa4_0(.dout(w_dff_A_9VJhQXUh0_0),.din(w_dff_A_aYNYGUpa4_0),.clk(gclk));
	jdff dff_A_9VJhQXUh0_0(.dout(w_dff_A_xvgY8m9d7_0),.din(w_dff_A_9VJhQXUh0_0),.clk(gclk));
	jdff dff_A_xvgY8m9d7_0(.dout(w_dff_A_ernyu3e28_0),.din(w_dff_A_xvgY8m9d7_0),.clk(gclk));
	jdff dff_A_ernyu3e28_0(.dout(w_dff_A_4uFfwBbG9_0),.din(w_dff_A_ernyu3e28_0),.clk(gclk));
	jdff dff_A_4uFfwBbG9_0(.dout(w_dff_A_mckkwymu8_0),.din(w_dff_A_4uFfwBbG9_0),.clk(gclk));
	jdff dff_A_mckkwymu8_0(.dout(w_dff_A_weLrtYMy0_0),.din(w_dff_A_mckkwymu8_0),.clk(gclk));
	jdff dff_A_weLrtYMy0_0(.dout(w_dff_A_vRFb8hrF5_0),.din(w_dff_A_weLrtYMy0_0),.clk(gclk));
	jdff dff_A_vRFb8hrF5_0(.dout(w_dff_A_GP5KH0aN7_0),.din(w_dff_A_vRFb8hrF5_0),.clk(gclk));
	jdff dff_A_GP5KH0aN7_0(.dout(w_dff_A_0YryPYix4_0),.din(w_dff_A_GP5KH0aN7_0),.clk(gclk));
	jdff dff_A_0YryPYix4_0(.dout(w_dff_A_Idl9YaUA0_0),.din(w_dff_A_0YryPYix4_0),.clk(gclk));
	jdff dff_A_Idl9YaUA0_0(.dout(w_dff_A_YuSX56it9_0),.din(w_dff_A_Idl9YaUA0_0),.clk(gclk));
	jdff dff_A_YuSX56it9_0(.dout(w_dff_A_RNJFjpIk6_0),.din(w_dff_A_YuSX56it9_0),.clk(gclk));
	jdff dff_A_RNJFjpIk6_0(.dout(w_dff_A_p0UhPUEZ0_0),.din(w_dff_A_RNJFjpIk6_0),.clk(gclk));
	jdff dff_A_p0UhPUEZ0_0(.dout(w_dff_A_HNCAy7Cb2_0),.din(w_dff_A_p0UhPUEZ0_0),.clk(gclk));
	jdff dff_A_HNCAy7Cb2_0(.dout(w_dff_A_SqR5GScA3_0),.din(w_dff_A_HNCAy7Cb2_0),.clk(gclk));
	jdff dff_A_SqR5GScA3_0(.dout(w_dff_A_zCCKVcRW1_0),.din(w_dff_A_SqR5GScA3_0),.clk(gclk));
	jdff dff_A_zCCKVcRW1_0(.dout(w_dff_A_Qevygbzi0_0),.din(w_dff_A_zCCKVcRW1_0),.clk(gclk));
	jdff dff_A_Qevygbzi0_0(.dout(w_dff_A_pGSbur8B1_0),.din(w_dff_A_Qevygbzi0_0),.clk(gclk));
	jdff dff_A_pGSbur8B1_0(.dout(w_dff_A_JXc14ZzH6_0),.din(w_dff_A_pGSbur8B1_0),.clk(gclk));
	jdff dff_A_JXc14ZzH6_0(.dout(w_dff_A_Xa9PaJDy1_0),.din(w_dff_A_JXc14ZzH6_0),.clk(gclk));
	jdff dff_A_Xa9PaJDy1_0(.dout(w_dff_A_JodmWguB4_0),.din(w_dff_A_Xa9PaJDy1_0),.clk(gclk));
	jdff dff_A_JodmWguB4_0(.dout(w_dff_A_1VCMknYK8_0),.din(w_dff_A_JodmWguB4_0),.clk(gclk));
	jdff dff_A_1VCMknYK8_0(.dout(w_dff_A_xPOqCAD35_0),.din(w_dff_A_1VCMknYK8_0),.clk(gclk));
	jdff dff_A_xPOqCAD35_0(.dout(w_dff_A_JGEFaSEz3_0),.din(w_dff_A_xPOqCAD35_0),.clk(gclk));
	jdff dff_A_JGEFaSEz3_0(.dout(w_dff_A_bTiUZa0d0_0),.din(w_dff_A_JGEFaSEz3_0),.clk(gclk));
	jdff dff_A_bTiUZa0d0_0(.dout(w_dff_A_bFtFCiV93_0),.din(w_dff_A_bTiUZa0d0_0),.clk(gclk));
	jdff dff_A_bFtFCiV93_0(.dout(w_dff_A_JDnTg7Wy2_0),.din(w_dff_A_bFtFCiV93_0),.clk(gclk));
	jdff dff_A_JDnTg7Wy2_0(.dout(w_dff_A_0xGYnvYT9_0),.din(w_dff_A_JDnTg7Wy2_0),.clk(gclk));
	jdff dff_A_0xGYnvYT9_0(.dout(w_dff_A_Rx2AkfOZ7_0),.din(w_dff_A_0xGYnvYT9_0),.clk(gclk));
	jdff dff_A_Rx2AkfOZ7_0(.dout(w_dff_A_Id7s039g1_0),.din(w_dff_A_Rx2AkfOZ7_0),.clk(gclk));
	jdff dff_A_Id7s039g1_0(.dout(w_dff_A_FeHNKsXG8_0),.din(w_dff_A_Id7s039g1_0),.clk(gclk));
	jdff dff_A_FeHNKsXG8_0(.dout(w_dff_A_373RZLtH2_0),.din(w_dff_A_FeHNKsXG8_0),.clk(gclk));
	jdff dff_A_373RZLtH2_0(.dout(w_dff_A_cy6TiKAY7_0),.din(w_dff_A_373RZLtH2_0),.clk(gclk));
	jdff dff_A_cy6TiKAY7_0(.dout(w_dff_A_zqHffu1C6_0),.din(w_dff_A_cy6TiKAY7_0),.clk(gclk));
	jdff dff_A_zqHffu1C6_0(.dout(w_dff_A_yBIXVU8B0_0),.din(w_dff_A_zqHffu1C6_0),.clk(gclk));
	jdff dff_A_yBIXVU8B0_0(.dout(w_dff_A_hohG6Ava7_0),.din(w_dff_A_yBIXVU8B0_0),.clk(gclk));
	jdff dff_A_hohG6Ava7_0(.dout(w_dff_A_YrozW7jp0_0),.din(w_dff_A_hohG6Ava7_0),.clk(gclk));
	jdff dff_A_YrozW7jp0_0(.dout(w_dff_A_ozpiGovK3_0),.din(w_dff_A_YrozW7jp0_0),.clk(gclk));
	jdff dff_A_ozpiGovK3_0(.dout(w_dff_A_dqAuvGf84_0),.din(w_dff_A_ozpiGovK3_0),.clk(gclk));
	jdff dff_A_dqAuvGf84_0(.dout(w_dff_A_MjaYf2H42_0),.din(w_dff_A_dqAuvGf84_0),.clk(gclk));
	jdff dff_A_MjaYf2H42_0(.dout(w_dff_A_fh10UvDM3_0),.din(w_dff_A_MjaYf2H42_0),.clk(gclk));
	jdff dff_A_fh10UvDM3_0(.dout(w_dff_A_GftTKNNO5_0),.din(w_dff_A_fh10UvDM3_0),.clk(gclk));
	jdff dff_A_GftTKNNO5_0(.dout(w_dff_A_LOkLnOjh0_0),.din(w_dff_A_GftTKNNO5_0),.clk(gclk));
	jdff dff_A_LOkLnOjh0_0(.dout(w_dff_A_vKPllyVC5_0),.din(w_dff_A_LOkLnOjh0_0),.clk(gclk));
	jdff dff_A_vKPllyVC5_0(.dout(w_dff_A_d0RxXPR64_0),.din(w_dff_A_vKPllyVC5_0),.clk(gclk));
	jdff dff_A_d0RxXPR64_0(.dout(w_dff_A_QvVkHKpg3_0),.din(w_dff_A_d0RxXPR64_0),.clk(gclk));
	jdff dff_A_QvVkHKpg3_0(.dout(w_dff_A_GaRmSQ3Z4_0),.din(w_dff_A_QvVkHKpg3_0),.clk(gclk));
	jdff dff_A_GaRmSQ3Z4_0(.dout(w_dff_A_MLa1aEM94_0),.din(w_dff_A_GaRmSQ3Z4_0),.clk(gclk));
	jdff dff_A_MLa1aEM94_0(.dout(w_dff_A_npUhE63i2_0),.din(w_dff_A_MLa1aEM94_0),.clk(gclk));
	jdff dff_A_npUhE63i2_0(.dout(w_dff_A_h3uBRfXY5_0),.din(w_dff_A_npUhE63i2_0),.clk(gclk));
	jdff dff_A_h3uBRfXY5_0(.dout(w_dff_A_UrcCR59f5_0),.din(w_dff_A_h3uBRfXY5_0),.clk(gclk));
	jdff dff_A_UrcCR59f5_0(.dout(w_dff_A_wWJe65Pb1_0),.din(w_dff_A_UrcCR59f5_0),.clk(gclk));
	jdff dff_A_wWJe65Pb1_0(.dout(w_dff_A_j2CmVjSk5_0),.din(w_dff_A_wWJe65Pb1_0),.clk(gclk));
	jdff dff_A_j2CmVjSk5_0(.dout(f41),.din(w_dff_A_j2CmVjSk5_0),.clk(gclk));
	jdff dff_A_09ujqjlu8_2(.dout(w_dff_A_be74fz819_0),.din(w_dff_A_09ujqjlu8_2),.clk(gclk));
	jdff dff_A_be74fz819_0(.dout(w_dff_A_I8xteb4F9_0),.din(w_dff_A_be74fz819_0),.clk(gclk));
	jdff dff_A_I8xteb4F9_0(.dout(w_dff_A_VGF7z3iy1_0),.din(w_dff_A_I8xteb4F9_0),.clk(gclk));
	jdff dff_A_VGF7z3iy1_0(.dout(w_dff_A_sDZi5Mfg2_0),.din(w_dff_A_VGF7z3iy1_0),.clk(gclk));
	jdff dff_A_sDZi5Mfg2_0(.dout(w_dff_A_tbda1U0P4_0),.din(w_dff_A_sDZi5Mfg2_0),.clk(gclk));
	jdff dff_A_tbda1U0P4_0(.dout(w_dff_A_MufNjFSd8_0),.din(w_dff_A_tbda1U0P4_0),.clk(gclk));
	jdff dff_A_MufNjFSd8_0(.dout(w_dff_A_DlmJ5lzi0_0),.din(w_dff_A_MufNjFSd8_0),.clk(gclk));
	jdff dff_A_DlmJ5lzi0_0(.dout(w_dff_A_WVLj8wRy6_0),.din(w_dff_A_DlmJ5lzi0_0),.clk(gclk));
	jdff dff_A_WVLj8wRy6_0(.dout(w_dff_A_xtE0Ueya9_0),.din(w_dff_A_WVLj8wRy6_0),.clk(gclk));
	jdff dff_A_xtE0Ueya9_0(.dout(w_dff_A_bjSse2pa1_0),.din(w_dff_A_xtE0Ueya9_0),.clk(gclk));
	jdff dff_A_bjSse2pa1_0(.dout(w_dff_A_hoWIJ4us4_0),.din(w_dff_A_bjSse2pa1_0),.clk(gclk));
	jdff dff_A_hoWIJ4us4_0(.dout(w_dff_A_upKxRkym8_0),.din(w_dff_A_hoWIJ4us4_0),.clk(gclk));
	jdff dff_A_upKxRkym8_0(.dout(w_dff_A_RJCqsJvr3_0),.din(w_dff_A_upKxRkym8_0),.clk(gclk));
	jdff dff_A_RJCqsJvr3_0(.dout(w_dff_A_nzmIOttB8_0),.din(w_dff_A_RJCqsJvr3_0),.clk(gclk));
	jdff dff_A_nzmIOttB8_0(.dout(w_dff_A_UeRAWBye8_0),.din(w_dff_A_nzmIOttB8_0),.clk(gclk));
	jdff dff_A_UeRAWBye8_0(.dout(w_dff_A_kiyyZw0H3_0),.din(w_dff_A_UeRAWBye8_0),.clk(gclk));
	jdff dff_A_kiyyZw0H3_0(.dout(w_dff_A_JCNxAO7s4_0),.din(w_dff_A_kiyyZw0H3_0),.clk(gclk));
	jdff dff_A_JCNxAO7s4_0(.dout(w_dff_A_SEjjlhd79_0),.din(w_dff_A_JCNxAO7s4_0),.clk(gclk));
	jdff dff_A_SEjjlhd79_0(.dout(w_dff_A_dPGrPTZq1_0),.din(w_dff_A_SEjjlhd79_0),.clk(gclk));
	jdff dff_A_dPGrPTZq1_0(.dout(w_dff_A_pXA8IV9V3_0),.din(w_dff_A_dPGrPTZq1_0),.clk(gclk));
	jdff dff_A_pXA8IV9V3_0(.dout(w_dff_A_CKqMEaNF6_0),.din(w_dff_A_pXA8IV9V3_0),.clk(gclk));
	jdff dff_A_CKqMEaNF6_0(.dout(w_dff_A_aQhVcq0b3_0),.din(w_dff_A_CKqMEaNF6_0),.clk(gclk));
	jdff dff_A_aQhVcq0b3_0(.dout(w_dff_A_hRhEXDo67_0),.din(w_dff_A_aQhVcq0b3_0),.clk(gclk));
	jdff dff_A_hRhEXDo67_0(.dout(w_dff_A_LrdEYM1a5_0),.din(w_dff_A_hRhEXDo67_0),.clk(gclk));
	jdff dff_A_LrdEYM1a5_0(.dout(w_dff_A_AjIxpUJS5_0),.din(w_dff_A_LrdEYM1a5_0),.clk(gclk));
	jdff dff_A_AjIxpUJS5_0(.dout(w_dff_A_BnDQLnGE7_0),.din(w_dff_A_AjIxpUJS5_0),.clk(gclk));
	jdff dff_A_BnDQLnGE7_0(.dout(w_dff_A_Jnzh4Z970_0),.din(w_dff_A_BnDQLnGE7_0),.clk(gclk));
	jdff dff_A_Jnzh4Z970_0(.dout(w_dff_A_LIVMCQeI7_0),.din(w_dff_A_Jnzh4Z970_0),.clk(gclk));
	jdff dff_A_LIVMCQeI7_0(.dout(w_dff_A_9bO3gilc0_0),.din(w_dff_A_LIVMCQeI7_0),.clk(gclk));
	jdff dff_A_9bO3gilc0_0(.dout(w_dff_A_91CtK90a0_0),.din(w_dff_A_9bO3gilc0_0),.clk(gclk));
	jdff dff_A_91CtK90a0_0(.dout(w_dff_A_0V7efWrM5_0),.din(w_dff_A_91CtK90a0_0),.clk(gclk));
	jdff dff_A_0V7efWrM5_0(.dout(w_dff_A_KO6zhEyl8_0),.din(w_dff_A_0V7efWrM5_0),.clk(gclk));
	jdff dff_A_KO6zhEyl8_0(.dout(w_dff_A_zgXRiywV5_0),.din(w_dff_A_KO6zhEyl8_0),.clk(gclk));
	jdff dff_A_zgXRiywV5_0(.dout(w_dff_A_zGfviu9u3_0),.din(w_dff_A_zgXRiywV5_0),.clk(gclk));
	jdff dff_A_zGfviu9u3_0(.dout(w_dff_A_66rZtyR85_0),.din(w_dff_A_zGfviu9u3_0),.clk(gclk));
	jdff dff_A_66rZtyR85_0(.dout(w_dff_A_CLw6JZE77_0),.din(w_dff_A_66rZtyR85_0),.clk(gclk));
	jdff dff_A_CLw6JZE77_0(.dout(w_dff_A_tO3ncZsQ3_0),.din(w_dff_A_CLw6JZE77_0),.clk(gclk));
	jdff dff_A_tO3ncZsQ3_0(.dout(w_dff_A_zhxgy1SI9_0),.din(w_dff_A_tO3ncZsQ3_0),.clk(gclk));
	jdff dff_A_zhxgy1SI9_0(.dout(w_dff_A_F02IGJHi6_0),.din(w_dff_A_zhxgy1SI9_0),.clk(gclk));
	jdff dff_A_F02IGJHi6_0(.dout(w_dff_A_vlgSZwsw9_0),.din(w_dff_A_F02IGJHi6_0),.clk(gclk));
	jdff dff_A_vlgSZwsw9_0(.dout(w_dff_A_QvmUDdwW1_0),.din(w_dff_A_vlgSZwsw9_0),.clk(gclk));
	jdff dff_A_QvmUDdwW1_0(.dout(w_dff_A_qs5sUFd54_0),.din(w_dff_A_QvmUDdwW1_0),.clk(gclk));
	jdff dff_A_qs5sUFd54_0(.dout(w_dff_A_tvvEPsvj5_0),.din(w_dff_A_qs5sUFd54_0),.clk(gclk));
	jdff dff_A_tvvEPsvj5_0(.dout(w_dff_A_m2rz8ZOa0_0),.din(w_dff_A_tvvEPsvj5_0),.clk(gclk));
	jdff dff_A_m2rz8ZOa0_0(.dout(w_dff_A_7b5xt8Jb6_0),.din(w_dff_A_m2rz8ZOa0_0),.clk(gclk));
	jdff dff_A_7b5xt8Jb6_0(.dout(w_dff_A_RMLMDYql2_0),.din(w_dff_A_7b5xt8Jb6_0),.clk(gclk));
	jdff dff_A_RMLMDYql2_0(.dout(w_dff_A_RxVrpxhD1_0),.din(w_dff_A_RMLMDYql2_0),.clk(gclk));
	jdff dff_A_RxVrpxhD1_0(.dout(w_dff_A_KsCP3sLU8_0),.din(w_dff_A_RxVrpxhD1_0),.clk(gclk));
	jdff dff_A_KsCP3sLU8_0(.dout(w_dff_A_CgPlzuhz8_0),.din(w_dff_A_KsCP3sLU8_0),.clk(gclk));
	jdff dff_A_CgPlzuhz8_0(.dout(w_dff_A_cNLxJw9X6_0),.din(w_dff_A_CgPlzuhz8_0),.clk(gclk));
	jdff dff_A_cNLxJw9X6_0(.dout(w_dff_A_fniQDc2H5_0),.din(w_dff_A_cNLxJw9X6_0),.clk(gclk));
	jdff dff_A_fniQDc2H5_0(.dout(w_dff_A_9xlETZAD4_0),.din(w_dff_A_fniQDc2H5_0),.clk(gclk));
	jdff dff_A_9xlETZAD4_0(.dout(w_dff_A_JL50S49p1_0),.din(w_dff_A_9xlETZAD4_0),.clk(gclk));
	jdff dff_A_JL50S49p1_0(.dout(w_dff_A_MlwASfw96_0),.din(w_dff_A_JL50S49p1_0),.clk(gclk));
	jdff dff_A_MlwASfw96_0(.dout(w_dff_A_dygkZ9gN4_0),.din(w_dff_A_MlwASfw96_0),.clk(gclk));
	jdff dff_A_dygkZ9gN4_0(.dout(w_dff_A_7NS9T6Ij1_0),.din(w_dff_A_dygkZ9gN4_0),.clk(gclk));
	jdff dff_A_7NS9T6Ij1_0(.dout(w_dff_A_ArA2uCLg4_0),.din(w_dff_A_7NS9T6Ij1_0),.clk(gclk));
	jdff dff_A_ArA2uCLg4_0(.dout(w_dff_A_jCK4P6Gw0_0),.din(w_dff_A_ArA2uCLg4_0),.clk(gclk));
	jdff dff_A_jCK4P6Gw0_0(.dout(w_dff_A_V7HGuMDS9_0),.din(w_dff_A_jCK4P6Gw0_0),.clk(gclk));
	jdff dff_A_V7HGuMDS9_0(.dout(w_dff_A_LCFq9c2U4_0),.din(w_dff_A_V7HGuMDS9_0),.clk(gclk));
	jdff dff_A_LCFq9c2U4_0(.dout(w_dff_A_RhWuPDMP0_0),.din(w_dff_A_LCFq9c2U4_0),.clk(gclk));
	jdff dff_A_RhWuPDMP0_0(.dout(w_dff_A_UrqmSOGO9_0),.din(w_dff_A_RhWuPDMP0_0),.clk(gclk));
	jdff dff_A_UrqmSOGO9_0(.dout(w_dff_A_B6kVDOoH6_0),.din(w_dff_A_UrqmSOGO9_0),.clk(gclk));
	jdff dff_A_B6kVDOoH6_0(.dout(w_dff_A_u49tUYXQ0_0),.din(w_dff_A_B6kVDOoH6_0),.clk(gclk));
	jdff dff_A_u49tUYXQ0_0(.dout(w_dff_A_VSIPmh6y8_0),.din(w_dff_A_u49tUYXQ0_0),.clk(gclk));
	jdff dff_A_VSIPmh6y8_0(.dout(w_dff_A_OAqUtPXc4_0),.din(w_dff_A_VSIPmh6y8_0),.clk(gclk));
	jdff dff_A_OAqUtPXc4_0(.dout(w_dff_A_OFsA9OWJ8_0),.din(w_dff_A_OAqUtPXc4_0),.clk(gclk));
	jdff dff_A_OFsA9OWJ8_0(.dout(w_dff_A_ic1PIJyN5_0),.din(w_dff_A_OFsA9OWJ8_0),.clk(gclk));
	jdff dff_A_ic1PIJyN5_0(.dout(w_dff_A_zckYKGVP9_0),.din(w_dff_A_ic1PIJyN5_0),.clk(gclk));
	jdff dff_A_zckYKGVP9_0(.dout(w_dff_A_vdsyRhqH3_0),.din(w_dff_A_zckYKGVP9_0),.clk(gclk));
	jdff dff_A_vdsyRhqH3_0(.dout(w_dff_A_zp7XrHna3_0),.din(w_dff_A_vdsyRhqH3_0),.clk(gclk));
	jdff dff_A_zp7XrHna3_0(.dout(w_dff_A_CvWdVhc81_0),.din(w_dff_A_zp7XrHna3_0),.clk(gclk));
	jdff dff_A_CvWdVhc81_0(.dout(w_dff_A_30dp7QUw0_0),.din(w_dff_A_CvWdVhc81_0),.clk(gclk));
	jdff dff_A_30dp7QUw0_0(.dout(w_dff_A_JYfTop5S5_0),.din(w_dff_A_30dp7QUw0_0),.clk(gclk));
	jdff dff_A_JYfTop5S5_0(.dout(w_dff_A_CTAMHKIb9_0),.din(w_dff_A_JYfTop5S5_0),.clk(gclk));
	jdff dff_A_CTAMHKIb9_0(.dout(w_dff_A_3NHchMO86_0),.din(w_dff_A_CTAMHKIb9_0),.clk(gclk));
	jdff dff_A_3NHchMO86_0(.dout(w_dff_A_YhkumKvG9_0),.din(w_dff_A_3NHchMO86_0),.clk(gclk));
	jdff dff_A_YhkumKvG9_0(.dout(w_dff_A_8gLtMPJH2_0),.din(w_dff_A_YhkumKvG9_0),.clk(gclk));
	jdff dff_A_8gLtMPJH2_0(.dout(w_dff_A_1KkeRVA44_0),.din(w_dff_A_8gLtMPJH2_0),.clk(gclk));
	jdff dff_A_1KkeRVA44_0(.dout(w_dff_A_E6sukExO1_0),.din(w_dff_A_1KkeRVA44_0),.clk(gclk));
	jdff dff_A_E6sukExO1_0(.dout(w_dff_A_muRFRCui3_0),.din(w_dff_A_E6sukExO1_0),.clk(gclk));
	jdff dff_A_muRFRCui3_0(.dout(w_dff_A_ouyj3V846_0),.din(w_dff_A_muRFRCui3_0),.clk(gclk));
	jdff dff_A_ouyj3V846_0(.dout(w_dff_A_pwOQZeRs9_0),.din(w_dff_A_ouyj3V846_0),.clk(gclk));
	jdff dff_A_pwOQZeRs9_0(.dout(w_dff_A_mr6hoPYX7_0),.din(w_dff_A_pwOQZeRs9_0),.clk(gclk));
	jdff dff_A_mr6hoPYX7_0(.dout(f42),.din(w_dff_A_mr6hoPYX7_0),.clk(gclk));
	jdff dff_A_I2YmvXsD7_2(.dout(w_dff_A_iwwCAYjP4_0),.din(w_dff_A_I2YmvXsD7_2),.clk(gclk));
	jdff dff_A_iwwCAYjP4_0(.dout(w_dff_A_9p7EbxrT3_0),.din(w_dff_A_iwwCAYjP4_0),.clk(gclk));
	jdff dff_A_9p7EbxrT3_0(.dout(w_dff_A_mBoupQAV6_0),.din(w_dff_A_9p7EbxrT3_0),.clk(gclk));
	jdff dff_A_mBoupQAV6_0(.dout(w_dff_A_dazKTbJF6_0),.din(w_dff_A_mBoupQAV6_0),.clk(gclk));
	jdff dff_A_dazKTbJF6_0(.dout(w_dff_A_YV3D9fTu4_0),.din(w_dff_A_dazKTbJF6_0),.clk(gclk));
	jdff dff_A_YV3D9fTu4_0(.dout(w_dff_A_5ICCUItY9_0),.din(w_dff_A_YV3D9fTu4_0),.clk(gclk));
	jdff dff_A_5ICCUItY9_0(.dout(w_dff_A_KAtL8Svj9_0),.din(w_dff_A_5ICCUItY9_0),.clk(gclk));
	jdff dff_A_KAtL8Svj9_0(.dout(w_dff_A_o0tbN3Rf5_0),.din(w_dff_A_KAtL8Svj9_0),.clk(gclk));
	jdff dff_A_o0tbN3Rf5_0(.dout(w_dff_A_3aglvj2B9_0),.din(w_dff_A_o0tbN3Rf5_0),.clk(gclk));
	jdff dff_A_3aglvj2B9_0(.dout(w_dff_A_0QZOk1Tt1_0),.din(w_dff_A_3aglvj2B9_0),.clk(gclk));
	jdff dff_A_0QZOk1Tt1_0(.dout(w_dff_A_RlsEu0s89_0),.din(w_dff_A_0QZOk1Tt1_0),.clk(gclk));
	jdff dff_A_RlsEu0s89_0(.dout(w_dff_A_mrf5lEzd8_0),.din(w_dff_A_RlsEu0s89_0),.clk(gclk));
	jdff dff_A_mrf5lEzd8_0(.dout(w_dff_A_K7n24jrx6_0),.din(w_dff_A_mrf5lEzd8_0),.clk(gclk));
	jdff dff_A_K7n24jrx6_0(.dout(w_dff_A_KhX8Zs792_0),.din(w_dff_A_K7n24jrx6_0),.clk(gclk));
	jdff dff_A_KhX8Zs792_0(.dout(w_dff_A_8XcG8xDf8_0),.din(w_dff_A_KhX8Zs792_0),.clk(gclk));
	jdff dff_A_8XcG8xDf8_0(.dout(w_dff_A_fRkOhPgT2_0),.din(w_dff_A_8XcG8xDf8_0),.clk(gclk));
	jdff dff_A_fRkOhPgT2_0(.dout(w_dff_A_1Aflo9lq5_0),.din(w_dff_A_fRkOhPgT2_0),.clk(gclk));
	jdff dff_A_1Aflo9lq5_0(.dout(w_dff_A_Z1ZPN1hd9_0),.din(w_dff_A_1Aflo9lq5_0),.clk(gclk));
	jdff dff_A_Z1ZPN1hd9_0(.dout(w_dff_A_Aj3mC7Yq8_0),.din(w_dff_A_Z1ZPN1hd9_0),.clk(gclk));
	jdff dff_A_Aj3mC7Yq8_0(.dout(w_dff_A_ctIBh6Wp8_0),.din(w_dff_A_Aj3mC7Yq8_0),.clk(gclk));
	jdff dff_A_ctIBh6Wp8_0(.dout(w_dff_A_zuvrfReM5_0),.din(w_dff_A_ctIBh6Wp8_0),.clk(gclk));
	jdff dff_A_zuvrfReM5_0(.dout(w_dff_A_xOdwzxux1_0),.din(w_dff_A_zuvrfReM5_0),.clk(gclk));
	jdff dff_A_xOdwzxux1_0(.dout(w_dff_A_IVGsGoaU6_0),.din(w_dff_A_xOdwzxux1_0),.clk(gclk));
	jdff dff_A_IVGsGoaU6_0(.dout(w_dff_A_0WhriuVL4_0),.din(w_dff_A_IVGsGoaU6_0),.clk(gclk));
	jdff dff_A_0WhriuVL4_0(.dout(w_dff_A_CQDIP57e0_0),.din(w_dff_A_0WhriuVL4_0),.clk(gclk));
	jdff dff_A_CQDIP57e0_0(.dout(w_dff_A_jTXsJJre9_0),.din(w_dff_A_CQDIP57e0_0),.clk(gclk));
	jdff dff_A_jTXsJJre9_0(.dout(w_dff_A_ivmbgxt15_0),.din(w_dff_A_jTXsJJre9_0),.clk(gclk));
	jdff dff_A_ivmbgxt15_0(.dout(w_dff_A_oF0LvA588_0),.din(w_dff_A_ivmbgxt15_0),.clk(gclk));
	jdff dff_A_oF0LvA588_0(.dout(w_dff_A_YaiEmU210_0),.din(w_dff_A_oF0LvA588_0),.clk(gclk));
	jdff dff_A_YaiEmU210_0(.dout(w_dff_A_ePXmgAeT0_0),.din(w_dff_A_YaiEmU210_0),.clk(gclk));
	jdff dff_A_ePXmgAeT0_0(.dout(w_dff_A_CrFaqAzs6_0),.din(w_dff_A_ePXmgAeT0_0),.clk(gclk));
	jdff dff_A_CrFaqAzs6_0(.dout(w_dff_A_sd9WIwLu6_0),.din(w_dff_A_CrFaqAzs6_0),.clk(gclk));
	jdff dff_A_sd9WIwLu6_0(.dout(w_dff_A_cyhdTi2s7_0),.din(w_dff_A_sd9WIwLu6_0),.clk(gclk));
	jdff dff_A_cyhdTi2s7_0(.dout(w_dff_A_Ebrbe4Ro5_0),.din(w_dff_A_cyhdTi2s7_0),.clk(gclk));
	jdff dff_A_Ebrbe4Ro5_0(.dout(w_dff_A_oUJM2Xul3_0),.din(w_dff_A_Ebrbe4Ro5_0),.clk(gclk));
	jdff dff_A_oUJM2Xul3_0(.dout(w_dff_A_BbnissWg5_0),.din(w_dff_A_oUJM2Xul3_0),.clk(gclk));
	jdff dff_A_BbnissWg5_0(.dout(w_dff_A_EG7x2Eyy4_0),.din(w_dff_A_BbnissWg5_0),.clk(gclk));
	jdff dff_A_EG7x2Eyy4_0(.dout(w_dff_A_wV8ZhxCo5_0),.din(w_dff_A_EG7x2Eyy4_0),.clk(gclk));
	jdff dff_A_wV8ZhxCo5_0(.dout(w_dff_A_47GtF05j5_0),.din(w_dff_A_wV8ZhxCo5_0),.clk(gclk));
	jdff dff_A_47GtF05j5_0(.dout(w_dff_A_loQ3y2CI1_0),.din(w_dff_A_47GtF05j5_0),.clk(gclk));
	jdff dff_A_loQ3y2CI1_0(.dout(w_dff_A_8PssS20B1_0),.din(w_dff_A_loQ3y2CI1_0),.clk(gclk));
	jdff dff_A_8PssS20B1_0(.dout(w_dff_A_dxvju1Yp4_0),.din(w_dff_A_8PssS20B1_0),.clk(gclk));
	jdff dff_A_dxvju1Yp4_0(.dout(w_dff_A_5GFDt7Em0_0),.din(w_dff_A_dxvju1Yp4_0),.clk(gclk));
	jdff dff_A_5GFDt7Em0_0(.dout(w_dff_A_vf1L7Tlg0_0),.din(w_dff_A_5GFDt7Em0_0),.clk(gclk));
	jdff dff_A_vf1L7Tlg0_0(.dout(w_dff_A_jMxMaCax5_0),.din(w_dff_A_vf1L7Tlg0_0),.clk(gclk));
	jdff dff_A_jMxMaCax5_0(.dout(w_dff_A_y0aBSAA14_0),.din(w_dff_A_jMxMaCax5_0),.clk(gclk));
	jdff dff_A_y0aBSAA14_0(.dout(w_dff_A_UcENqhBs2_0),.din(w_dff_A_y0aBSAA14_0),.clk(gclk));
	jdff dff_A_UcENqhBs2_0(.dout(w_dff_A_8i7DLpwY8_0),.din(w_dff_A_UcENqhBs2_0),.clk(gclk));
	jdff dff_A_8i7DLpwY8_0(.dout(w_dff_A_lLY9jVsG9_0),.din(w_dff_A_8i7DLpwY8_0),.clk(gclk));
	jdff dff_A_lLY9jVsG9_0(.dout(w_dff_A_KVDN2Mls1_0),.din(w_dff_A_lLY9jVsG9_0),.clk(gclk));
	jdff dff_A_KVDN2Mls1_0(.dout(w_dff_A_68UTzHBK5_0),.din(w_dff_A_KVDN2Mls1_0),.clk(gclk));
	jdff dff_A_68UTzHBK5_0(.dout(w_dff_A_4qDqqGwG1_0),.din(w_dff_A_68UTzHBK5_0),.clk(gclk));
	jdff dff_A_4qDqqGwG1_0(.dout(w_dff_A_kHXU97Lc7_0),.din(w_dff_A_4qDqqGwG1_0),.clk(gclk));
	jdff dff_A_kHXU97Lc7_0(.dout(w_dff_A_XpPYjHLw5_0),.din(w_dff_A_kHXU97Lc7_0),.clk(gclk));
	jdff dff_A_XpPYjHLw5_0(.dout(w_dff_A_flJKFsXs7_0),.din(w_dff_A_XpPYjHLw5_0),.clk(gclk));
	jdff dff_A_flJKFsXs7_0(.dout(w_dff_A_D7MGyajg3_0),.din(w_dff_A_flJKFsXs7_0),.clk(gclk));
	jdff dff_A_D7MGyajg3_0(.dout(w_dff_A_phhfLAtf2_0),.din(w_dff_A_D7MGyajg3_0),.clk(gclk));
	jdff dff_A_phhfLAtf2_0(.dout(w_dff_A_lEEZB3fQ8_0),.din(w_dff_A_phhfLAtf2_0),.clk(gclk));
	jdff dff_A_lEEZB3fQ8_0(.dout(w_dff_A_KDeHjTUE0_0),.din(w_dff_A_lEEZB3fQ8_0),.clk(gclk));
	jdff dff_A_KDeHjTUE0_0(.dout(w_dff_A_Bbf8bry06_0),.din(w_dff_A_KDeHjTUE0_0),.clk(gclk));
	jdff dff_A_Bbf8bry06_0(.dout(w_dff_A_bohYFnGH5_0),.din(w_dff_A_Bbf8bry06_0),.clk(gclk));
	jdff dff_A_bohYFnGH5_0(.dout(w_dff_A_EicDp3dW2_0),.din(w_dff_A_bohYFnGH5_0),.clk(gclk));
	jdff dff_A_EicDp3dW2_0(.dout(w_dff_A_gRCiM6iH3_0),.din(w_dff_A_EicDp3dW2_0),.clk(gclk));
	jdff dff_A_gRCiM6iH3_0(.dout(w_dff_A_P87bsD3U0_0),.din(w_dff_A_gRCiM6iH3_0),.clk(gclk));
	jdff dff_A_P87bsD3U0_0(.dout(w_dff_A_58f8sd3p0_0),.din(w_dff_A_P87bsD3U0_0),.clk(gclk));
	jdff dff_A_58f8sd3p0_0(.dout(w_dff_A_YhN4a1Q65_0),.din(w_dff_A_58f8sd3p0_0),.clk(gclk));
	jdff dff_A_YhN4a1Q65_0(.dout(w_dff_A_egnquzXW2_0),.din(w_dff_A_YhN4a1Q65_0),.clk(gclk));
	jdff dff_A_egnquzXW2_0(.dout(w_dff_A_dXhZkiuG8_0),.din(w_dff_A_egnquzXW2_0),.clk(gclk));
	jdff dff_A_dXhZkiuG8_0(.dout(w_dff_A_JHVMi7LS0_0),.din(w_dff_A_dXhZkiuG8_0),.clk(gclk));
	jdff dff_A_JHVMi7LS0_0(.dout(w_dff_A_QzZnwF7e5_0),.din(w_dff_A_JHVMi7LS0_0),.clk(gclk));
	jdff dff_A_QzZnwF7e5_0(.dout(w_dff_A_6HgVXsN02_0),.din(w_dff_A_QzZnwF7e5_0),.clk(gclk));
	jdff dff_A_6HgVXsN02_0(.dout(w_dff_A_hbakRN0M2_0),.din(w_dff_A_6HgVXsN02_0),.clk(gclk));
	jdff dff_A_hbakRN0M2_0(.dout(w_dff_A_QAEXknsg6_0),.din(w_dff_A_hbakRN0M2_0),.clk(gclk));
	jdff dff_A_QAEXknsg6_0(.dout(w_dff_A_QnYlALgD3_0),.din(w_dff_A_QAEXknsg6_0),.clk(gclk));
	jdff dff_A_QnYlALgD3_0(.dout(w_dff_A_J769Eo012_0),.din(w_dff_A_QnYlALgD3_0),.clk(gclk));
	jdff dff_A_J769Eo012_0(.dout(w_dff_A_dIiHWuHW0_0),.din(w_dff_A_J769Eo012_0),.clk(gclk));
	jdff dff_A_dIiHWuHW0_0(.dout(w_dff_A_awPYj27s3_0),.din(w_dff_A_dIiHWuHW0_0),.clk(gclk));
	jdff dff_A_awPYj27s3_0(.dout(w_dff_A_6RgqpFib8_0),.din(w_dff_A_awPYj27s3_0),.clk(gclk));
	jdff dff_A_6RgqpFib8_0(.dout(w_dff_A_FgVjMgpT8_0),.din(w_dff_A_6RgqpFib8_0),.clk(gclk));
	jdff dff_A_FgVjMgpT8_0(.dout(w_dff_A_Fhux8ibn9_0),.din(w_dff_A_FgVjMgpT8_0),.clk(gclk));
	jdff dff_A_Fhux8ibn9_0(.dout(w_dff_A_ExWud07P6_0),.din(w_dff_A_Fhux8ibn9_0),.clk(gclk));
	jdff dff_A_ExWud07P6_0(.dout(w_dff_A_yDKO6jnY6_0),.din(w_dff_A_ExWud07P6_0),.clk(gclk));
	jdff dff_A_yDKO6jnY6_0(.dout(w_dff_A_i9TXfYjA3_0),.din(w_dff_A_yDKO6jnY6_0),.clk(gclk));
	jdff dff_A_i9TXfYjA3_0(.dout(f43),.din(w_dff_A_i9TXfYjA3_0),.clk(gclk));
	jdff dff_A_QwZFXhVA9_2(.dout(w_dff_A_nvkloFpO9_0),.din(w_dff_A_QwZFXhVA9_2),.clk(gclk));
	jdff dff_A_nvkloFpO9_0(.dout(w_dff_A_LbIgM0Sr3_0),.din(w_dff_A_nvkloFpO9_0),.clk(gclk));
	jdff dff_A_LbIgM0Sr3_0(.dout(w_dff_A_H0iNvINO7_0),.din(w_dff_A_LbIgM0Sr3_0),.clk(gclk));
	jdff dff_A_H0iNvINO7_0(.dout(w_dff_A_RundX8An2_0),.din(w_dff_A_H0iNvINO7_0),.clk(gclk));
	jdff dff_A_RundX8An2_0(.dout(w_dff_A_9rxmYfdH1_0),.din(w_dff_A_RundX8An2_0),.clk(gclk));
	jdff dff_A_9rxmYfdH1_0(.dout(w_dff_A_xFel332I6_0),.din(w_dff_A_9rxmYfdH1_0),.clk(gclk));
	jdff dff_A_xFel332I6_0(.dout(w_dff_A_af9wKAWX3_0),.din(w_dff_A_xFel332I6_0),.clk(gclk));
	jdff dff_A_af9wKAWX3_0(.dout(w_dff_A_YsM1BgCH8_0),.din(w_dff_A_af9wKAWX3_0),.clk(gclk));
	jdff dff_A_YsM1BgCH8_0(.dout(w_dff_A_GadyavqL7_0),.din(w_dff_A_YsM1BgCH8_0),.clk(gclk));
	jdff dff_A_GadyavqL7_0(.dout(w_dff_A_xEiZUlON1_0),.din(w_dff_A_GadyavqL7_0),.clk(gclk));
	jdff dff_A_xEiZUlON1_0(.dout(w_dff_A_mUMsLDWr3_0),.din(w_dff_A_xEiZUlON1_0),.clk(gclk));
	jdff dff_A_mUMsLDWr3_0(.dout(w_dff_A_ZVXD2CPn3_0),.din(w_dff_A_mUMsLDWr3_0),.clk(gclk));
	jdff dff_A_ZVXD2CPn3_0(.dout(w_dff_A_JSxkZfCp4_0),.din(w_dff_A_ZVXD2CPn3_0),.clk(gclk));
	jdff dff_A_JSxkZfCp4_0(.dout(w_dff_A_AmTlAO325_0),.din(w_dff_A_JSxkZfCp4_0),.clk(gclk));
	jdff dff_A_AmTlAO325_0(.dout(w_dff_A_Pvxw8xvc6_0),.din(w_dff_A_AmTlAO325_0),.clk(gclk));
	jdff dff_A_Pvxw8xvc6_0(.dout(w_dff_A_81QK1hPd9_0),.din(w_dff_A_Pvxw8xvc6_0),.clk(gclk));
	jdff dff_A_81QK1hPd9_0(.dout(w_dff_A_GOB7TVp82_0),.din(w_dff_A_81QK1hPd9_0),.clk(gclk));
	jdff dff_A_GOB7TVp82_0(.dout(w_dff_A_Yli3KqZy3_0),.din(w_dff_A_GOB7TVp82_0),.clk(gclk));
	jdff dff_A_Yli3KqZy3_0(.dout(w_dff_A_yfOL9Q0B2_0),.din(w_dff_A_Yli3KqZy3_0),.clk(gclk));
	jdff dff_A_yfOL9Q0B2_0(.dout(w_dff_A_vLarxcGg2_0),.din(w_dff_A_yfOL9Q0B2_0),.clk(gclk));
	jdff dff_A_vLarxcGg2_0(.dout(w_dff_A_xe0yl61c4_0),.din(w_dff_A_vLarxcGg2_0),.clk(gclk));
	jdff dff_A_xe0yl61c4_0(.dout(w_dff_A_uTizlrAL6_0),.din(w_dff_A_xe0yl61c4_0),.clk(gclk));
	jdff dff_A_uTizlrAL6_0(.dout(w_dff_A_ku1iD0Y45_0),.din(w_dff_A_uTizlrAL6_0),.clk(gclk));
	jdff dff_A_ku1iD0Y45_0(.dout(w_dff_A_EGR2RRYy4_0),.din(w_dff_A_ku1iD0Y45_0),.clk(gclk));
	jdff dff_A_EGR2RRYy4_0(.dout(w_dff_A_Zcrx2RQa9_0),.din(w_dff_A_EGR2RRYy4_0),.clk(gclk));
	jdff dff_A_Zcrx2RQa9_0(.dout(w_dff_A_s9LAINHP7_0),.din(w_dff_A_Zcrx2RQa9_0),.clk(gclk));
	jdff dff_A_s9LAINHP7_0(.dout(w_dff_A_2z9xenZG0_0),.din(w_dff_A_s9LAINHP7_0),.clk(gclk));
	jdff dff_A_2z9xenZG0_0(.dout(w_dff_A_NoDevIiG5_0),.din(w_dff_A_2z9xenZG0_0),.clk(gclk));
	jdff dff_A_NoDevIiG5_0(.dout(w_dff_A_KuJ735h86_0),.din(w_dff_A_NoDevIiG5_0),.clk(gclk));
	jdff dff_A_KuJ735h86_0(.dout(w_dff_A_aQ3KPV1F1_0),.din(w_dff_A_KuJ735h86_0),.clk(gclk));
	jdff dff_A_aQ3KPV1F1_0(.dout(w_dff_A_B6ElxsZl8_0),.din(w_dff_A_aQ3KPV1F1_0),.clk(gclk));
	jdff dff_A_B6ElxsZl8_0(.dout(w_dff_A_b7mtH4VV7_0),.din(w_dff_A_B6ElxsZl8_0),.clk(gclk));
	jdff dff_A_b7mtH4VV7_0(.dout(w_dff_A_q3qkhjU29_0),.din(w_dff_A_b7mtH4VV7_0),.clk(gclk));
	jdff dff_A_q3qkhjU29_0(.dout(w_dff_A_4u9iplea2_0),.din(w_dff_A_q3qkhjU29_0),.clk(gclk));
	jdff dff_A_4u9iplea2_0(.dout(w_dff_A_9EGFBIGa0_0),.din(w_dff_A_4u9iplea2_0),.clk(gclk));
	jdff dff_A_9EGFBIGa0_0(.dout(w_dff_A_K4YooPV45_0),.din(w_dff_A_9EGFBIGa0_0),.clk(gclk));
	jdff dff_A_K4YooPV45_0(.dout(w_dff_A_l7cCkc5d2_0),.din(w_dff_A_K4YooPV45_0),.clk(gclk));
	jdff dff_A_l7cCkc5d2_0(.dout(w_dff_A_sOC4NZV84_0),.din(w_dff_A_l7cCkc5d2_0),.clk(gclk));
	jdff dff_A_sOC4NZV84_0(.dout(w_dff_A_PuxORUE67_0),.din(w_dff_A_sOC4NZV84_0),.clk(gclk));
	jdff dff_A_PuxORUE67_0(.dout(w_dff_A_CDTko9DL1_0),.din(w_dff_A_PuxORUE67_0),.clk(gclk));
	jdff dff_A_CDTko9DL1_0(.dout(w_dff_A_WFz45bpl7_0),.din(w_dff_A_CDTko9DL1_0),.clk(gclk));
	jdff dff_A_WFz45bpl7_0(.dout(w_dff_A_boFmAM0m4_0),.din(w_dff_A_WFz45bpl7_0),.clk(gclk));
	jdff dff_A_boFmAM0m4_0(.dout(w_dff_A_acxQhCmO9_0),.din(w_dff_A_boFmAM0m4_0),.clk(gclk));
	jdff dff_A_acxQhCmO9_0(.dout(w_dff_A_blJxPUGY0_0),.din(w_dff_A_acxQhCmO9_0),.clk(gclk));
	jdff dff_A_blJxPUGY0_0(.dout(w_dff_A_Aig1CN4X5_0),.din(w_dff_A_blJxPUGY0_0),.clk(gclk));
	jdff dff_A_Aig1CN4X5_0(.dout(w_dff_A_VbChy4NS9_0),.din(w_dff_A_Aig1CN4X5_0),.clk(gclk));
	jdff dff_A_VbChy4NS9_0(.dout(w_dff_A_hDHVBNZY4_0),.din(w_dff_A_VbChy4NS9_0),.clk(gclk));
	jdff dff_A_hDHVBNZY4_0(.dout(w_dff_A_iOHFtmFf5_0),.din(w_dff_A_hDHVBNZY4_0),.clk(gclk));
	jdff dff_A_iOHFtmFf5_0(.dout(w_dff_A_2MTiY6nB1_0),.din(w_dff_A_iOHFtmFf5_0),.clk(gclk));
	jdff dff_A_2MTiY6nB1_0(.dout(w_dff_A_1n4N6PNy0_0),.din(w_dff_A_2MTiY6nB1_0),.clk(gclk));
	jdff dff_A_1n4N6PNy0_0(.dout(w_dff_A_BctyuwEo3_0),.din(w_dff_A_1n4N6PNy0_0),.clk(gclk));
	jdff dff_A_BctyuwEo3_0(.dout(w_dff_A_TNhBJMbf5_0),.din(w_dff_A_BctyuwEo3_0),.clk(gclk));
	jdff dff_A_TNhBJMbf5_0(.dout(w_dff_A_xUUKkhNU0_0),.din(w_dff_A_TNhBJMbf5_0),.clk(gclk));
	jdff dff_A_xUUKkhNU0_0(.dout(w_dff_A_6orM6LHi7_0),.din(w_dff_A_xUUKkhNU0_0),.clk(gclk));
	jdff dff_A_6orM6LHi7_0(.dout(w_dff_A_MwbP0iqd2_0),.din(w_dff_A_6orM6LHi7_0),.clk(gclk));
	jdff dff_A_MwbP0iqd2_0(.dout(w_dff_A_CljpVI755_0),.din(w_dff_A_MwbP0iqd2_0),.clk(gclk));
	jdff dff_A_CljpVI755_0(.dout(w_dff_A_XZcBWpOe8_0),.din(w_dff_A_CljpVI755_0),.clk(gclk));
	jdff dff_A_XZcBWpOe8_0(.dout(w_dff_A_N6QmLFWO4_0),.din(w_dff_A_XZcBWpOe8_0),.clk(gclk));
	jdff dff_A_N6QmLFWO4_0(.dout(w_dff_A_9XtA2kaC0_0),.din(w_dff_A_N6QmLFWO4_0),.clk(gclk));
	jdff dff_A_9XtA2kaC0_0(.dout(w_dff_A_jhlepn2y3_0),.din(w_dff_A_9XtA2kaC0_0),.clk(gclk));
	jdff dff_A_jhlepn2y3_0(.dout(w_dff_A_hjDgVkUM7_0),.din(w_dff_A_jhlepn2y3_0),.clk(gclk));
	jdff dff_A_hjDgVkUM7_0(.dout(w_dff_A_m1JHBSk70_0),.din(w_dff_A_hjDgVkUM7_0),.clk(gclk));
	jdff dff_A_m1JHBSk70_0(.dout(w_dff_A_IunuhWCv9_0),.din(w_dff_A_m1JHBSk70_0),.clk(gclk));
	jdff dff_A_IunuhWCv9_0(.dout(w_dff_A_y8jHW5686_0),.din(w_dff_A_IunuhWCv9_0),.clk(gclk));
	jdff dff_A_y8jHW5686_0(.dout(w_dff_A_aWhpgFXZ8_0),.din(w_dff_A_y8jHW5686_0),.clk(gclk));
	jdff dff_A_aWhpgFXZ8_0(.dout(w_dff_A_Ze0Tjzul6_0),.din(w_dff_A_aWhpgFXZ8_0),.clk(gclk));
	jdff dff_A_Ze0Tjzul6_0(.dout(w_dff_A_Tvg1wBCr4_0),.din(w_dff_A_Ze0Tjzul6_0),.clk(gclk));
	jdff dff_A_Tvg1wBCr4_0(.dout(w_dff_A_GvUqMuMM9_0),.din(w_dff_A_Tvg1wBCr4_0),.clk(gclk));
	jdff dff_A_GvUqMuMM9_0(.dout(w_dff_A_PgcqJA811_0),.din(w_dff_A_GvUqMuMM9_0),.clk(gclk));
	jdff dff_A_PgcqJA811_0(.dout(w_dff_A_51nk0jiv9_0),.din(w_dff_A_PgcqJA811_0),.clk(gclk));
	jdff dff_A_51nk0jiv9_0(.dout(w_dff_A_QLhtEXxF2_0),.din(w_dff_A_51nk0jiv9_0),.clk(gclk));
	jdff dff_A_QLhtEXxF2_0(.dout(w_dff_A_EQqmmGRC4_0),.din(w_dff_A_QLhtEXxF2_0),.clk(gclk));
	jdff dff_A_EQqmmGRC4_0(.dout(w_dff_A_PNHhgyPK1_0),.din(w_dff_A_EQqmmGRC4_0),.clk(gclk));
	jdff dff_A_PNHhgyPK1_0(.dout(w_dff_A_NAGUwB5e0_0),.din(w_dff_A_PNHhgyPK1_0),.clk(gclk));
	jdff dff_A_NAGUwB5e0_0(.dout(w_dff_A_AkjmE9m44_0),.din(w_dff_A_NAGUwB5e0_0),.clk(gclk));
	jdff dff_A_AkjmE9m44_0(.dout(w_dff_A_PJpTeiGq5_0),.din(w_dff_A_AkjmE9m44_0),.clk(gclk));
	jdff dff_A_PJpTeiGq5_0(.dout(w_dff_A_pss17xV59_0),.din(w_dff_A_PJpTeiGq5_0),.clk(gclk));
	jdff dff_A_pss17xV59_0(.dout(w_dff_A_Q9GGttvB4_0),.din(w_dff_A_pss17xV59_0),.clk(gclk));
	jdff dff_A_Q9GGttvB4_0(.dout(w_dff_A_wP2gzpTS6_0),.din(w_dff_A_Q9GGttvB4_0),.clk(gclk));
	jdff dff_A_wP2gzpTS6_0(.dout(w_dff_A_sDTcExYP1_0),.din(w_dff_A_wP2gzpTS6_0),.clk(gclk));
	jdff dff_A_sDTcExYP1_0(.dout(w_dff_A_spfe5KAf1_0),.din(w_dff_A_sDTcExYP1_0),.clk(gclk));
	jdff dff_A_spfe5KAf1_0(.dout(w_dff_A_liL365568_0),.din(w_dff_A_spfe5KAf1_0),.clk(gclk));
	jdff dff_A_liL365568_0(.dout(f44),.din(w_dff_A_liL365568_0),.clk(gclk));
	jdff dff_A_VA8FezrL8_2(.dout(w_dff_A_b226qRnN3_0),.din(w_dff_A_VA8FezrL8_2),.clk(gclk));
	jdff dff_A_b226qRnN3_0(.dout(w_dff_A_pZPQjE2g3_0),.din(w_dff_A_b226qRnN3_0),.clk(gclk));
	jdff dff_A_pZPQjE2g3_0(.dout(w_dff_A_8iIdkfKF8_0),.din(w_dff_A_pZPQjE2g3_0),.clk(gclk));
	jdff dff_A_8iIdkfKF8_0(.dout(w_dff_A_o1GZ0zij0_0),.din(w_dff_A_8iIdkfKF8_0),.clk(gclk));
	jdff dff_A_o1GZ0zij0_0(.dout(w_dff_A_if8Baa843_0),.din(w_dff_A_o1GZ0zij0_0),.clk(gclk));
	jdff dff_A_if8Baa843_0(.dout(w_dff_A_UAz8SeHi6_0),.din(w_dff_A_if8Baa843_0),.clk(gclk));
	jdff dff_A_UAz8SeHi6_0(.dout(w_dff_A_sg4Csuqz8_0),.din(w_dff_A_UAz8SeHi6_0),.clk(gclk));
	jdff dff_A_sg4Csuqz8_0(.dout(w_dff_A_4o1VsA5K8_0),.din(w_dff_A_sg4Csuqz8_0),.clk(gclk));
	jdff dff_A_4o1VsA5K8_0(.dout(w_dff_A_iCI7vs3b9_0),.din(w_dff_A_4o1VsA5K8_0),.clk(gclk));
	jdff dff_A_iCI7vs3b9_0(.dout(w_dff_A_UMYRLIK44_0),.din(w_dff_A_iCI7vs3b9_0),.clk(gclk));
	jdff dff_A_UMYRLIK44_0(.dout(w_dff_A_oYqbKALq1_0),.din(w_dff_A_UMYRLIK44_0),.clk(gclk));
	jdff dff_A_oYqbKALq1_0(.dout(w_dff_A_y2unAVqf9_0),.din(w_dff_A_oYqbKALq1_0),.clk(gclk));
	jdff dff_A_y2unAVqf9_0(.dout(w_dff_A_gI3iWxhH5_0),.din(w_dff_A_y2unAVqf9_0),.clk(gclk));
	jdff dff_A_gI3iWxhH5_0(.dout(w_dff_A_wMP0kDfA4_0),.din(w_dff_A_gI3iWxhH5_0),.clk(gclk));
	jdff dff_A_wMP0kDfA4_0(.dout(w_dff_A_aYdScR2t7_0),.din(w_dff_A_wMP0kDfA4_0),.clk(gclk));
	jdff dff_A_aYdScR2t7_0(.dout(w_dff_A_XCCaEhXv4_0),.din(w_dff_A_aYdScR2t7_0),.clk(gclk));
	jdff dff_A_XCCaEhXv4_0(.dout(w_dff_A_1uG86Qwl6_0),.din(w_dff_A_XCCaEhXv4_0),.clk(gclk));
	jdff dff_A_1uG86Qwl6_0(.dout(w_dff_A_xRbjSe2j1_0),.din(w_dff_A_1uG86Qwl6_0),.clk(gclk));
	jdff dff_A_xRbjSe2j1_0(.dout(w_dff_A_SmxzjB9o1_0),.din(w_dff_A_xRbjSe2j1_0),.clk(gclk));
	jdff dff_A_SmxzjB9o1_0(.dout(w_dff_A_OPR2Dgfc7_0),.din(w_dff_A_SmxzjB9o1_0),.clk(gclk));
	jdff dff_A_OPR2Dgfc7_0(.dout(w_dff_A_2g2TVycB8_0),.din(w_dff_A_OPR2Dgfc7_0),.clk(gclk));
	jdff dff_A_2g2TVycB8_0(.dout(w_dff_A_vIvx6jIH3_0),.din(w_dff_A_2g2TVycB8_0),.clk(gclk));
	jdff dff_A_vIvx6jIH3_0(.dout(w_dff_A_eRmnPQA45_0),.din(w_dff_A_vIvx6jIH3_0),.clk(gclk));
	jdff dff_A_eRmnPQA45_0(.dout(w_dff_A_zz7xbobE6_0),.din(w_dff_A_eRmnPQA45_0),.clk(gclk));
	jdff dff_A_zz7xbobE6_0(.dout(w_dff_A_GNkl9cSO1_0),.din(w_dff_A_zz7xbobE6_0),.clk(gclk));
	jdff dff_A_GNkl9cSO1_0(.dout(w_dff_A_dLlbPJj91_0),.din(w_dff_A_GNkl9cSO1_0),.clk(gclk));
	jdff dff_A_dLlbPJj91_0(.dout(w_dff_A_HsZ4XLDi9_0),.din(w_dff_A_dLlbPJj91_0),.clk(gclk));
	jdff dff_A_HsZ4XLDi9_0(.dout(w_dff_A_lnF6INVy1_0),.din(w_dff_A_HsZ4XLDi9_0),.clk(gclk));
	jdff dff_A_lnF6INVy1_0(.dout(w_dff_A_PtH2FU308_0),.din(w_dff_A_lnF6INVy1_0),.clk(gclk));
	jdff dff_A_PtH2FU308_0(.dout(w_dff_A_bLRHLw6I0_0),.din(w_dff_A_PtH2FU308_0),.clk(gclk));
	jdff dff_A_bLRHLw6I0_0(.dout(w_dff_A_qTs8cf0U2_0),.din(w_dff_A_bLRHLw6I0_0),.clk(gclk));
	jdff dff_A_qTs8cf0U2_0(.dout(w_dff_A_4AX9puio9_0),.din(w_dff_A_qTs8cf0U2_0),.clk(gclk));
	jdff dff_A_4AX9puio9_0(.dout(w_dff_A_gJHyPL2e9_0),.din(w_dff_A_4AX9puio9_0),.clk(gclk));
	jdff dff_A_gJHyPL2e9_0(.dout(w_dff_A_WisRR6O13_0),.din(w_dff_A_gJHyPL2e9_0),.clk(gclk));
	jdff dff_A_WisRR6O13_0(.dout(w_dff_A_19Do98xE4_0),.din(w_dff_A_WisRR6O13_0),.clk(gclk));
	jdff dff_A_19Do98xE4_0(.dout(w_dff_A_kczk54597_0),.din(w_dff_A_19Do98xE4_0),.clk(gclk));
	jdff dff_A_kczk54597_0(.dout(w_dff_A_myTyPijs6_0),.din(w_dff_A_kczk54597_0),.clk(gclk));
	jdff dff_A_myTyPijs6_0(.dout(w_dff_A_4kvYeWPA1_0),.din(w_dff_A_myTyPijs6_0),.clk(gclk));
	jdff dff_A_4kvYeWPA1_0(.dout(w_dff_A_S9e7LfMG8_0),.din(w_dff_A_4kvYeWPA1_0),.clk(gclk));
	jdff dff_A_S9e7LfMG8_0(.dout(w_dff_A_XgxjNJ0K7_0),.din(w_dff_A_S9e7LfMG8_0),.clk(gclk));
	jdff dff_A_XgxjNJ0K7_0(.dout(w_dff_A_FKlQSajr2_0),.din(w_dff_A_XgxjNJ0K7_0),.clk(gclk));
	jdff dff_A_FKlQSajr2_0(.dout(w_dff_A_xedhvIKq8_0),.din(w_dff_A_FKlQSajr2_0),.clk(gclk));
	jdff dff_A_xedhvIKq8_0(.dout(w_dff_A_LvhQ5N1D1_0),.din(w_dff_A_xedhvIKq8_0),.clk(gclk));
	jdff dff_A_LvhQ5N1D1_0(.dout(w_dff_A_LtTvRMsL8_0),.din(w_dff_A_LvhQ5N1D1_0),.clk(gclk));
	jdff dff_A_LtTvRMsL8_0(.dout(w_dff_A_w4u5U6lP8_0),.din(w_dff_A_LtTvRMsL8_0),.clk(gclk));
	jdff dff_A_w4u5U6lP8_0(.dout(w_dff_A_4SoVkHw83_0),.din(w_dff_A_w4u5U6lP8_0),.clk(gclk));
	jdff dff_A_4SoVkHw83_0(.dout(w_dff_A_uI1Xt1Ht0_0),.din(w_dff_A_4SoVkHw83_0),.clk(gclk));
	jdff dff_A_uI1Xt1Ht0_0(.dout(w_dff_A_2xt2lJfA0_0),.din(w_dff_A_uI1Xt1Ht0_0),.clk(gclk));
	jdff dff_A_2xt2lJfA0_0(.dout(w_dff_A_VJFz8Uom7_0),.din(w_dff_A_2xt2lJfA0_0),.clk(gclk));
	jdff dff_A_VJFz8Uom7_0(.dout(w_dff_A_4mVtzz5I9_0),.din(w_dff_A_VJFz8Uom7_0),.clk(gclk));
	jdff dff_A_4mVtzz5I9_0(.dout(w_dff_A_Jh0Pbxth0_0),.din(w_dff_A_4mVtzz5I9_0),.clk(gclk));
	jdff dff_A_Jh0Pbxth0_0(.dout(w_dff_A_ep2o8L4k1_0),.din(w_dff_A_Jh0Pbxth0_0),.clk(gclk));
	jdff dff_A_ep2o8L4k1_0(.dout(w_dff_A_ZfGnjXiW7_0),.din(w_dff_A_ep2o8L4k1_0),.clk(gclk));
	jdff dff_A_ZfGnjXiW7_0(.dout(w_dff_A_pWPCIsz71_0),.din(w_dff_A_ZfGnjXiW7_0),.clk(gclk));
	jdff dff_A_pWPCIsz71_0(.dout(w_dff_A_catsBTZK1_0),.din(w_dff_A_pWPCIsz71_0),.clk(gclk));
	jdff dff_A_catsBTZK1_0(.dout(w_dff_A_mlRZ4bO28_0),.din(w_dff_A_catsBTZK1_0),.clk(gclk));
	jdff dff_A_mlRZ4bO28_0(.dout(w_dff_A_CTOicfeF0_0),.din(w_dff_A_mlRZ4bO28_0),.clk(gclk));
	jdff dff_A_CTOicfeF0_0(.dout(w_dff_A_TJ5n8bcQ7_0),.din(w_dff_A_CTOicfeF0_0),.clk(gclk));
	jdff dff_A_TJ5n8bcQ7_0(.dout(w_dff_A_laPYLZzS2_0),.din(w_dff_A_TJ5n8bcQ7_0),.clk(gclk));
	jdff dff_A_laPYLZzS2_0(.dout(w_dff_A_4FOur9j23_0),.din(w_dff_A_laPYLZzS2_0),.clk(gclk));
	jdff dff_A_4FOur9j23_0(.dout(w_dff_A_Sf8DfBWg5_0),.din(w_dff_A_4FOur9j23_0),.clk(gclk));
	jdff dff_A_Sf8DfBWg5_0(.dout(w_dff_A_zbu4IAnq0_0),.din(w_dff_A_Sf8DfBWg5_0),.clk(gclk));
	jdff dff_A_zbu4IAnq0_0(.dout(w_dff_A_58knblez0_0),.din(w_dff_A_zbu4IAnq0_0),.clk(gclk));
	jdff dff_A_58knblez0_0(.dout(w_dff_A_1rYtvV0Z8_0),.din(w_dff_A_58knblez0_0),.clk(gclk));
	jdff dff_A_1rYtvV0Z8_0(.dout(w_dff_A_F8kjRSmg6_0),.din(w_dff_A_1rYtvV0Z8_0),.clk(gclk));
	jdff dff_A_F8kjRSmg6_0(.dout(w_dff_A_lPw9gapI9_0),.din(w_dff_A_F8kjRSmg6_0),.clk(gclk));
	jdff dff_A_lPw9gapI9_0(.dout(w_dff_A_dfkK1r7m6_0),.din(w_dff_A_lPw9gapI9_0),.clk(gclk));
	jdff dff_A_dfkK1r7m6_0(.dout(w_dff_A_SeZGPuyv4_0),.din(w_dff_A_dfkK1r7m6_0),.clk(gclk));
	jdff dff_A_SeZGPuyv4_0(.dout(w_dff_A_HZStFoNn9_0),.din(w_dff_A_SeZGPuyv4_0),.clk(gclk));
	jdff dff_A_HZStFoNn9_0(.dout(w_dff_A_KIP5wquy5_0),.din(w_dff_A_HZStFoNn9_0),.clk(gclk));
	jdff dff_A_KIP5wquy5_0(.dout(w_dff_A_HXrZOhLr9_0),.din(w_dff_A_KIP5wquy5_0),.clk(gclk));
	jdff dff_A_HXrZOhLr9_0(.dout(w_dff_A_Znn79pgt7_0),.din(w_dff_A_HXrZOhLr9_0),.clk(gclk));
	jdff dff_A_Znn79pgt7_0(.dout(w_dff_A_3sEmRykW0_0),.din(w_dff_A_Znn79pgt7_0),.clk(gclk));
	jdff dff_A_3sEmRykW0_0(.dout(w_dff_A_Qlwi5kWE7_0),.din(w_dff_A_3sEmRykW0_0),.clk(gclk));
	jdff dff_A_Qlwi5kWE7_0(.dout(w_dff_A_6t05PBfO9_0),.din(w_dff_A_Qlwi5kWE7_0),.clk(gclk));
	jdff dff_A_6t05PBfO9_0(.dout(w_dff_A_hNUpVLeR7_0),.din(w_dff_A_6t05PBfO9_0),.clk(gclk));
	jdff dff_A_hNUpVLeR7_0(.dout(w_dff_A_9yqlOFht4_0),.din(w_dff_A_hNUpVLeR7_0),.clk(gclk));
	jdff dff_A_9yqlOFht4_0(.dout(w_dff_A_pskIfvvL5_0),.din(w_dff_A_9yqlOFht4_0),.clk(gclk));
	jdff dff_A_pskIfvvL5_0(.dout(w_dff_A_6FTNQ2Kh1_0),.din(w_dff_A_pskIfvvL5_0),.clk(gclk));
	jdff dff_A_6FTNQ2Kh1_0(.dout(w_dff_A_uhHD4lyL4_0),.din(w_dff_A_6FTNQ2Kh1_0),.clk(gclk));
	jdff dff_A_uhHD4lyL4_0(.dout(w_dff_A_aDYoSPHZ4_0),.din(w_dff_A_uhHD4lyL4_0),.clk(gclk));
	jdff dff_A_aDYoSPHZ4_0(.dout(f45),.din(w_dff_A_aDYoSPHZ4_0),.clk(gclk));
	jdff dff_A_HG05Fu3s6_2(.dout(w_dff_A_1Y3ZXEOD9_0),.din(w_dff_A_HG05Fu3s6_2),.clk(gclk));
	jdff dff_A_1Y3ZXEOD9_0(.dout(w_dff_A_rsaC8EOD4_0),.din(w_dff_A_1Y3ZXEOD9_0),.clk(gclk));
	jdff dff_A_rsaC8EOD4_0(.dout(w_dff_A_yJa8GiY56_0),.din(w_dff_A_rsaC8EOD4_0),.clk(gclk));
	jdff dff_A_yJa8GiY56_0(.dout(w_dff_A_d2U2JZ351_0),.din(w_dff_A_yJa8GiY56_0),.clk(gclk));
	jdff dff_A_d2U2JZ351_0(.dout(w_dff_A_eiabcs987_0),.din(w_dff_A_d2U2JZ351_0),.clk(gclk));
	jdff dff_A_eiabcs987_0(.dout(w_dff_A_oT8JnhJB9_0),.din(w_dff_A_eiabcs987_0),.clk(gclk));
	jdff dff_A_oT8JnhJB9_0(.dout(w_dff_A_4O6DHlfK5_0),.din(w_dff_A_oT8JnhJB9_0),.clk(gclk));
	jdff dff_A_4O6DHlfK5_0(.dout(w_dff_A_Axp9Kb249_0),.din(w_dff_A_4O6DHlfK5_0),.clk(gclk));
	jdff dff_A_Axp9Kb249_0(.dout(w_dff_A_JtWxbxBH8_0),.din(w_dff_A_Axp9Kb249_0),.clk(gclk));
	jdff dff_A_JtWxbxBH8_0(.dout(w_dff_A_BNiSuHog3_0),.din(w_dff_A_JtWxbxBH8_0),.clk(gclk));
	jdff dff_A_BNiSuHog3_0(.dout(w_dff_A_Itc1YIAW7_0),.din(w_dff_A_BNiSuHog3_0),.clk(gclk));
	jdff dff_A_Itc1YIAW7_0(.dout(w_dff_A_YKCK1I1K7_0),.din(w_dff_A_Itc1YIAW7_0),.clk(gclk));
	jdff dff_A_YKCK1I1K7_0(.dout(w_dff_A_JjPsMhjR4_0),.din(w_dff_A_YKCK1I1K7_0),.clk(gclk));
	jdff dff_A_JjPsMhjR4_0(.dout(w_dff_A_vSPqQAyF0_0),.din(w_dff_A_JjPsMhjR4_0),.clk(gclk));
	jdff dff_A_vSPqQAyF0_0(.dout(w_dff_A_m9NmUZsP0_0),.din(w_dff_A_vSPqQAyF0_0),.clk(gclk));
	jdff dff_A_m9NmUZsP0_0(.dout(w_dff_A_WCnoFlRp1_0),.din(w_dff_A_m9NmUZsP0_0),.clk(gclk));
	jdff dff_A_WCnoFlRp1_0(.dout(w_dff_A_q1nV2qLW9_0),.din(w_dff_A_WCnoFlRp1_0),.clk(gclk));
	jdff dff_A_q1nV2qLW9_0(.dout(w_dff_A_QYTzw6fn8_0),.din(w_dff_A_q1nV2qLW9_0),.clk(gclk));
	jdff dff_A_QYTzw6fn8_0(.dout(w_dff_A_3b2N48St1_0),.din(w_dff_A_QYTzw6fn8_0),.clk(gclk));
	jdff dff_A_3b2N48St1_0(.dout(w_dff_A_QvS2scxK0_0),.din(w_dff_A_3b2N48St1_0),.clk(gclk));
	jdff dff_A_QvS2scxK0_0(.dout(w_dff_A_cj63GRbJ6_0),.din(w_dff_A_QvS2scxK0_0),.clk(gclk));
	jdff dff_A_cj63GRbJ6_0(.dout(w_dff_A_qGrn4L5R4_0),.din(w_dff_A_cj63GRbJ6_0),.clk(gclk));
	jdff dff_A_qGrn4L5R4_0(.dout(w_dff_A_nTSRAmSa6_0),.din(w_dff_A_qGrn4L5R4_0),.clk(gclk));
	jdff dff_A_nTSRAmSa6_0(.dout(w_dff_A_BOoo0Xz64_0),.din(w_dff_A_nTSRAmSa6_0),.clk(gclk));
	jdff dff_A_BOoo0Xz64_0(.dout(w_dff_A_7q1MmhDE7_0),.din(w_dff_A_BOoo0Xz64_0),.clk(gclk));
	jdff dff_A_7q1MmhDE7_0(.dout(w_dff_A_pbsXAUVu7_0),.din(w_dff_A_7q1MmhDE7_0),.clk(gclk));
	jdff dff_A_pbsXAUVu7_0(.dout(w_dff_A_NNkfLj2L5_0),.din(w_dff_A_pbsXAUVu7_0),.clk(gclk));
	jdff dff_A_NNkfLj2L5_0(.dout(w_dff_A_JSNZxt6X2_0),.din(w_dff_A_NNkfLj2L5_0),.clk(gclk));
	jdff dff_A_JSNZxt6X2_0(.dout(w_dff_A_UjzPN8SU4_0),.din(w_dff_A_JSNZxt6X2_0),.clk(gclk));
	jdff dff_A_UjzPN8SU4_0(.dout(w_dff_A_qEJrqRI55_0),.din(w_dff_A_UjzPN8SU4_0),.clk(gclk));
	jdff dff_A_qEJrqRI55_0(.dout(w_dff_A_38cUQZwu9_0),.din(w_dff_A_qEJrqRI55_0),.clk(gclk));
	jdff dff_A_38cUQZwu9_0(.dout(w_dff_A_cfAXH0Q49_0),.din(w_dff_A_38cUQZwu9_0),.clk(gclk));
	jdff dff_A_cfAXH0Q49_0(.dout(w_dff_A_ezuQ3fGf2_0),.din(w_dff_A_cfAXH0Q49_0),.clk(gclk));
	jdff dff_A_ezuQ3fGf2_0(.dout(w_dff_A_7hofpAoX7_0),.din(w_dff_A_ezuQ3fGf2_0),.clk(gclk));
	jdff dff_A_7hofpAoX7_0(.dout(w_dff_A_44GbYigZ9_0),.din(w_dff_A_7hofpAoX7_0),.clk(gclk));
	jdff dff_A_44GbYigZ9_0(.dout(w_dff_A_17OAx2DH4_0),.din(w_dff_A_44GbYigZ9_0),.clk(gclk));
	jdff dff_A_17OAx2DH4_0(.dout(w_dff_A_8TO0W6bo3_0),.din(w_dff_A_17OAx2DH4_0),.clk(gclk));
	jdff dff_A_8TO0W6bo3_0(.dout(w_dff_A_fczQbtFl7_0),.din(w_dff_A_8TO0W6bo3_0),.clk(gclk));
	jdff dff_A_fczQbtFl7_0(.dout(w_dff_A_NdHswp9u8_0),.din(w_dff_A_fczQbtFl7_0),.clk(gclk));
	jdff dff_A_NdHswp9u8_0(.dout(w_dff_A_yEneimwF9_0),.din(w_dff_A_NdHswp9u8_0),.clk(gclk));
	jdff dff_A_yEneimwF9_0(.dout(w_dff_A_4owuKtWK4_0),.din(w_dff_A_yEneimwF9_0),.clk(gclk));
	jdff dff_A_4owuKtWK4_0(.dout(w_dff_A_RwptPYlL4_0),.din(w_dff_A_4owuKtWK4_0),.clk(gclk));
	jdff dff_A_RwptPYlL4_0(.dout(w_dff_A_LDHXtFyS9_0),.din(w_dff_A_RwptPYlL4_0),.clk(gclk));
	jdff dff_A_LDHXtFyS9_0(.dout(w_dff_A_7dAVMnmv3_0),.din(w_dff_A_LDHXtFyS9_0),.clk(gclk));
	jdff dff_A_7dAVMnmv3_0(.dout(w_dff_A_orhT70XV3_0),.din(w_dff_A_7dAVMnmv3_0),.clk(gclk));
	jdff dff_A_orhT70XV3_0(.dout(w_dff_A_GHWlDHQF7_0),.din(w_dff_A_orhT70XV3_0),.clk(gclk));
	jdff dff_A_GHWlDHQF7_0(.dout(w_dff_A_F0gPMduf0_0),.din(w_dff_A_GHWlDHQF7_0),.clk(gclk));
	jdff dff_A_F0gPMduf0_0(.dout(w_dff_A_Kh7bOlBZ0_0),.din(w_dff_A_F0gPMduf0_0),.clk(gclk));
	jdff dff_A_Kh7bOlBZ0_0(.dout(w_dff_A_4SMjnric5_0),.din(w_dff_A_Kh7bOlBZ0_0),.clk(gclk));
	jdff dff_A_4SMjnric5_0(.dout(w_dff_A_HEtPXXun2_0),.din(w_dff_A_4SMjnric5_0),.clk(gclk));
	jdff dff_A_HEtPXXun2_0(.dout(w_dff_A_hU4xo7TJ9_0),.din(w_dff_A_HEtPXXun2_0),.clk(gclk));
	jdff dff_A_hU4xo7TJ9_0(.dout(w_dff_A_cNq82MEO3_0),.din(w_dff_A_hU4xo7TJ9_0),.clk(gclk));
	jdff dff_A_cNq82MEO3_0(.dout(w_dff_A_v9ERO0Hi2_0),.din(w_dff_A_cNq82MEO3_0),.clk(gclk));
	jdff dff_A_v9ERO0Hi2_0(.dout(w_dff_A_p6fawIhc5_0),.din(w_dff_A_v9ERO0Hi2_0),.clk(gclk));
	jdff dff_A_p6fawIhc5_0(.dout(w_dff_A_xjzdKE530_0),.din(w_dff_A_p6fawIhc5_0),.clk(gclk));
	jdff dff_A_xjzdKE530_0(.dout(w_dff_A_72mGvg8Z2_0),.din(w_dff_A_xjzdKE530_0),.clk(gclk));
	jdff dff_A_72mGvg8Z2_0(.dout(w_dff_A_aZYbpUCt3_0),.din(w_dff_A_72mGvg8Z2_0),.clk(gclk));
	jdff dff_A_aZYbpUCt3_0(.dout(w_dff_A_ISOq6j5g6_0),.din(w_dff_A_aZYbpUCt3_0),.clk(gclk));
	jdff dff_A_ISOq6j5g6_0(.dout(w_dff_A_wHy9NTg48_0),.din(w_dff_A_ISOq6j5g6_0),.clk(gclk));
	jdff dff_A_wHy9NTg48_0(.dout(w_dff_A_ko4ok0sf2_0),.din(w_dff_A_wHy9NTg48_0),.clk(gclk));
	jdff dff_A_ko4ok0sf2_0(.dout(w_dff_A_U4Jpn1HQ1_0),.din(w_dff_A_ko4ok0sf2_0),.clk(gclk));
	jdff dff_A_U4Jpn1HQ1_0(.dout(w_dff_A_ymMe0Kz95_0),.din(w_dff_A_U4Jpn1HQ1_0),.clk(gclk));
	jdff dff_A_ymMe0Kz95_0(.dout(w_dff_A_4g7pn8cp7_0),.din(w_dff_A_ymMe0Kz95_0),.clk(gclk));
	jdff dff_A_4g7pn8cp7_0(.dout(w_dff_A_h9ctqVME7_0),.din(w_dff_A_4g7pn8cp7_0),.clk(gclk));
	jdff dff_A_h9ctqVME7_0(.dout(w_dff_A_AIfM2gNc4_0),.din(w_dff_A_h9ctqVME7_0),.clk(gclk));
	jdff dff_A_AIfM2gNc4_0(.dout(w_dff_A_Q59DK8NO1_0),.din(w_dff_A_AIfM2gNc4_0),.clk(gclk));
	jdff dff_A_Q59DK8NO1_0(.dout(w_dff_A_KdUAUdq19_0),.din(w_dff_A_Q59DK8NO1_0),.clk(gclk));
	jdff dff_A_KdUAUdq19_0(.dout(w_dff_A_FX5IWUoc2_0),.din(w_dff_A_KdUAUdq19_0),.clk(gclk));
	jdff dff_A_FX5IWUoc2_0(.dout(w_dff_A_q7cZZz3O8_0),.din(w_dff_A_FX5IWUoc2_0),.clk(gclk));
	jdff dff_A_q7cZZz3O8_0(.dout(w_dff_A_3On6WqYB1_0),.din(w_dff_A_q7cZZz3O8_0),.clk(gclk));
	jdff dff_A_3On6WqYB1_0(.dout(w_dff_A_63tcd6cp9_0),.din(w_dff_A_3On6WqYB1_0),.clk(gclk));
	jdff dff_A_63tcd6cp9_0(.dout(w_dff_A_7iAXgQrL4_0),.din(w_dff_A_63tcd6cp9_0),.clk(gclk));
	jdff dff_A_7iAXgQrL4_0(.dout(w_dff_A_2JdxGfgq4_0),.din(w_dff_A_7iAXgQrL4_0),.clk(gclk));
	jdff dff_A_2JdxGfgq4_0(.dout(w_dff_A_LycyT0BB9_0),.din(w_dff_A_2JdxGfgq4_0),.clk(gclk));
	jdff dff_A_LycyT0BB9_0(.dout(w_dff_A_B1YASNI46_0),.din(w_dff_A_LycyT0BB9_0),.clk(gclk));
	jdff dff_A_B1YASNI46_0(.dout(w_dff_A_lQ5xWwDV2_0),.din(w_dff_A_B1YASNI46_0),.clk(gclk));
	jdff dff_A_lQ5xWwDV2_0(.dout(w_dff_A_UQL8PhEg0_0),.din(w_dff_A_lQ5xWwDV2_0),.clk(gclk));
	jdff dff_A_UQL8PhEg0_0(.dout(w_dff_A_dqLrMj3M3_0),.din(w_dff_A_UQL8PhEg0_0),.clk(gclk));
	jdff dff_A_dqLrMj3M3_0(.dout(w_dff_A_cSsadq7C0_0),.din(w_dff_A_dqLrMj3M3_0),.clk(gclk));
	jdff dff_A_cSsadq7C0_0(.dout(w_dff_A_WLW2og5L4_0),.din(w_dff_A_cSsadq7C0_0),.clk(gclk));
	jdff dff_A_WLW2og5L4_0(.dout(f46),.din(w_dff_A_WLW2og5L4_0),.clk(gclk));
	jdff dff_A_AIhCfEsq4_2(.dout(w_dff_A_Mcd8r44t0_0),.din(w_dff_A_AIhCfEsq4_2),.clk(gclk));
	jdff dff_A_Mcd8r44t0_0(.dout(w_dff_A_Qz76Zm9s4_0),.din(w_dff_A_Mcd8r44t0_0),.clk(gclk));
	jdff dff_A_Qz76Zm9s4_0(.dout(w_dff_A_2G23Zo3b2_0),.din(w_dff_A_Qz76Zm9s4_0),.clk(gclk));
	jdff dff_A_2G23Zo3b2_0(.dout(w_dff_A_pwAFPXiY0_0),.din(w_dff_A_2G23Zo3b2_0),.clk(gclk));
	jdff dff_A_pwAFPXiY0_0(.dout(w_dff_A_VJQ4SxBm8_0),.din(w_dff_A_pwAFPXiY0_0),.clk(gclk));
	jdff dff_A_VJQ4SxBm8_0(.dout(w_dff_A_LBYLBaZf6_0),.din(w_dff_A_VJQ4SxBm8_0),.clk(gclk));
	jdff dff_A_LBYLBaZf6_0(.dout(w_dff_A_npyf1nAS8_0),.din(w_dff_A_LBYLBaZf6_0),.clk(gclk));
	jdff dff_A_npyf1nAS8_0(.dout(w_dff_A_x4ZsDeE40_0),.din(w_dff_A_npyf1nAS8_0),.clk(gclk));
	jdff dff_A_x4ZsDeE40_0(.dout(w_dff_A_pb2gld0l1_0),.din(w_dff_A_x4ZsDeE40_0),.clk(gclk));
	jdff dff_A_pb2gld0l1_0(.dout(w_dff_A_m0P8Dk0L5_0),.din(w_dff_A_pb2gld0l1_0),.clk(gclk));
	jdff dff_A_m0P8Dk0L5_0(.dout(w_dff_A_LKxYA0WB2_0),.din(w_dff_A_m0P8Dk0L5_0),.clk(gclk));
	jdff dff_A_LKxYA0WB2_0(.dout(w_dff_A_MJpTqKJE0_0),.din(w_dff_A_LKxYA0WB2_0),.clk(gclk));
	jdff dff_A_MJpTqKJE0_0(.dout(w_dff_A_k1udsWbK9_0),.din(w_dff_A_MJpTqKJE0_0),.clk(gclk));
	jdff dff_A_k1udsWbK9_0(.dout(w_dff_A_oWtbHikt8_0),.din(w_dff_A_k1udsWbK9_0),.clk(gclk));
	jdff dff_A_oWtbHikt8_0(.dout(w_dff_A_QUJegnHs2_0),.din(w_dff_A_oWtbHikt8_0),.clk(gclk));
	jdff dff_A_QUJegnHs2_0(.dout(w_dff_A_BPIXwtwp8_0),.din(w_dff_A_QUJegnHs2_0),.clk(gclk));
	jdff dff_A_BPIXwtwp8_0(.dout(w_dff_A_11srEgQN9_0),.din(w_dff_A_BPIXwtwp8_0),.clk(gclk));
	jdff dff_A_11srEgQN9_0(.dout(w_dff_A_DbDtTKK26_0),.din(w_dff_A_11srEgQN9_0),.clk(gclk));
	jdff dff_A_DbDtTKK26_0(.dout(w_dff_A_uztct3wy2_0),.din(w_dff_A_DbDtTKK26_0),.clk(gclk));
	jdff dff_A_uztct3wy2_0(.dout(w_dff_A_IsPJJbj62_0),.din(w_dff_A_uztct3wy2_0),.clk(gclk));
	jdff dff_A_IsPJJbj62_0(.dout(w_dff_A_ulaPoL4U6_0),.din(w_dff_A_IsPJJbj62_0),.clk(gclk));
	jdff dff_A_ulaPoL4U6_0(.dout(w_dff_A_JEDaHwzL6_0),.din(w_dff_A_ulaPoL4U6_0),.clk(gclk));
	jdff dff_A_JEDaHwzL6_0(.dout(w_dff_A_XgUakTwu2_0),.din(w_dff_A_JEDaHwzL6_0),.clk(gclk));
	jdff dff_A_XgUakTwu2_0(.dout(w_dff_A_yVBiuFpG4_0),.din(w_dff_A_XgUakTwu2_0),.clk(gclk));
	jdff dff_A_yVBiuFpG4_0(.dout(w_dff_A_Zkot34Qt5_0),.din(w_dff_A_yVBiuFpG4_0),.clk(gclk));
	jdff dff_A_Zkot34Qt5_0(.dout(w_dff_A_GuYhh4d83_0),.din(w_dff_A_Zkot34Qt5_0),.clk(gclk));
	jdff dff_A_GuYhh4d83_0(.dout(w_dff_A_pzCSfwi07_0),.din(w_dff_A_GuYhh4d83_0),.clk(gclk));
	jdff dff_A_pzCSfwi07_0(.dout(w_dff_A_AqDyW98h9_0),.din(w_dff_A_pzCSfwi07_0),.clk(gclk));
	jdff dff_A_AqDyW98h9_0(.dout(w_dff_A_aXjtoTK27_0),.din(w_dff_A_AqDyW98h9_0),.clk(gclk));
	jdff dff_A_aXjtoTK27_0(.dout(w_dff_A_CyR4yuNj0_0),.din(w_dff_A_aXjtoTK27_0),.clk(gclk));
	jdff dff_A_CyR4yuNj0_0(.dout(w_dff_A_JnkblOjK9_0),.din(w_dff_A_CyR4yuNj0_0),.clk(gclk));
	jdff dff_A_JnkblOjK9_0(.dout(w_dff_A_CY9bIOQj4_0),.din(w_dff_A_JnkblOjK9_0),.clk(gclk));
	jdff dff_A_CY9bIOQj4_0(.dout(w_dff_A_eKWNEgVB3_0),.din(w_dff_A_CY9bIOQj4_0),.clk(gclk));
	jdff dff_A_eKWNEgVB3_0(.dout(w_dff_A_axhDMKbh6_0),.din(w_dff_A_eKWNEgVB3_0),.clk(gclk));
	jdff dff_A_axhDMKbh6_0(.dout(w_dff_A_Fz6TVdNW7_0),.din(w_dff_A_axhDMKbh6_0),.clk(gclk));
	jdff dff_A_Fz6TVdNW7_0(.dout(w_dff_A_Dr6sawMl5_0),.din(w_dff_A_Fz6TVdNW7_0),.clk(gclk));
	jdff dff_A_Dr6sawMl5_0(.dout(w_dff_A_I2VRxduo4_0),.din(w_dff_A_Dr6sawMl5_0),.clk(gclk));
	jdff dff_A_I2VRxduo4_0(.dout(w_dff_A_Go1GYNxA0_0),.din(w_dff_A_I2VRxduo4_0),.clk(gclk));
	jdff dff_A_Go1GYNxA0_0(.dout(w_dff_A_y8QegFjn5_0),.din(w_dff_A_Go1GYNxA0_0),.clk(gclk));
	jdff dff_A_y8QegFjn5_0(.dout(w_dff_A_TLN9vnk87_0),.din(w_dff_A_y8QegFjn5_0),.clk(gclk));
	jdff dff_A_TLN9vnk87_0(.dout(w_dff_A_Uq4FoVBv9_0),.din(w_dff_A_TLN9vnk87_0),.clk(gclk));
	jdff dff_A_Uq4FoVBv9_0(.dout(w_dff_A_W2W9dNqC7_0),.din(w_dff_A_Uq4FoVBv9_0),.clk(gclk));
	jdff dff_A_W2W9dNqC7_0(.dout(w_dff_A_x2objUkJ2_0),.din(w_dff_A_W2W9dNqC7_0),.clk(gclk));
	jdff dff_A_x2objUkJ2_0(.dout(w_dff_A_H9VUiw3e3_0),.din(w_dff_A_x2objUkJ2_0),.clk(gclk));
	jdff dff_A_H9VUiw3e3_0(.dout(w_dff_A_ZoFSIXa75_0),.din(w_dff_A_H9VUiw3e3_0),.clk(gclk));
	jdff dff_A_ZoFSIXa75_0(.dout(w_dff_A_396Ek8fd9_0),.din(w_dff_A_ZoFSIXa75_0),.clk(gclk));
	jdff dff_A_396Ek8fd9_0(.dout(w_dff_A_uqgLOtsS9_0),.din(w_dff_A_396Ek8fd9_0),.clk(gclk));
	jdff dff_A_uqgLOtsS9_0(.dout(w_dff_A_QeEHURnA2_0),.din(w_dff_A_uqgLOtsS9_0),.clk(gclk));
	jdff dff_A_QeEHURnA2_0(.dout(w_dff_A_BYUnO9Sh1_0),.din(w_dff_A_QeEHURnA2_0),.clk(gclk));
	jdff dff_A_BYUnO9Sh1_0(.dout(w_dff_A_3HYrIsu11_0),.din(w_dff_A_BYUnO9Sh1_0),.clk(gclk));
	jdff dff_A_3HYrIsu11_0(.dout(w_dff_A_1Cox9EfY1_0),.din(w_dff_A_3HYrIsu11_0),.clk(gclk));
	jdff dff_A_1Cox9EfY1_0(.dout(w_dff_A_vHYudDBo5_0),.din(w_dff_A_1Cox9EfY1_0),.clk(gclk));
	jdff dff_A_vHYudDBo5_0(.dout(w_dff_A_YqHoSDXs5_0),.din(w_dff_A_vHYudDBo5_0),.clk(gclk));
	jdff dff_A_YqHoSDXs5_0(.dout(w_dff_A_9790vaaC0_0),.din(w_dff_A_YqHoSDXs5_0),.clk(gclk));
	jdff dff_A_9790vaaC0_0(.dout(w_dff_A_gvXChzq40_0),.din(w_dff_A_9790vaaC0_0),.clk(gclk));
	jdff dff_A_gvXChzq40_0(.dout(w_dff_A_T56Os9rB3_0),.din(w_dff_A_gvXChzq40_0),.clk(gclk));
	jdff dff_A_T56Os9rB3_0(.dout(w_dff_A_7x7hpyfc0_0),.din(w_dff_A_T56Os9rB3_0),.clk(gclk));
	jdff dff_A_7x7hpyfc0_0(.dout(w_dff_A_4VmKR2rn3_0),.din(w_dff_A_7x7hpyfc0_0),.clk(gclk));
	jdff dff_A_4VmKR2rn3_0(.dout(w_dff_A_6pZ9RTP72_0),.din(w_dff_A_4VmKR2rn3_0),.clk(gclk));
	jdff dff_A_6pZ9RTP72_0(.dout(w_dff_A_qXLvXRzj6_0),.din(w_dff_A_6pZ9RTP72_0),.clk(gclk));
	jdff dff_A_qXLvXRzj6_0(.dout(w_dff_A_o8iW57Rc1_0),.din(w_dff_A_qXLvXRzj6_0),.clk(gclk));
	jdff dff_A_o8iW57Rc1_0(.dout(w_dff_A_4cUt3PnS1_0),.din(w_dff_A_o8iW57Rc1_0),.clk(gclk));
	jdff dff_A_4cUt3PnS1_0(.dout(w_dff_A_oa0VrNQq6_0),.din(w_dff_A_4cUt3PnS1_0),.clk(gclk));
	jdff dff_A_oa0VrNQq6_0(.dout(w_dff_A_be0FEAY46_0),.din(w_dff_A_oa0VrNQq6_0),.clk(gclk));
	jdff dff_A_be0FEAY46_0(.dout(w_dff_A_uTgQXcrR3_0),.din(w_dff_A_be0FEAY46_0),.clk(gclk));
	jdff dff_A_uTgQXcrR3_0(.dout(w_dff_A_0xZV8J2l9_0),.din(w_dff_A_uTgQXcrR3_0),.clk(gclk));
	jdff dff_A_0xZV8J2l9_0(.dout(w_dff_A_o13xOGmh6_0),.din(w_dff_A_0xZV8J2l9_0),.clk(gclk));
	jdff dff_A_o13xOGmh6_0(.dout(w_dff_A_GgOvRwNH3_0),.din(w_dff_A_o13xOGmh6_0),.clk(gclk));
	jdff dff_A_GgOvRwNH3_0(.dout(w_dff_A_n1h1dw9K3_0),.din(w_dff_A_GgOvRwNH3_0),.clk(gclk));
	jdff dff_A_n1h1dw9K3_0(.dout(w_dff_A_lVS80qA86_0),.din(w_dff_A_n1h1dw9K3_0),.clk(gclk));
	jdff dff_A_lVS80qA86_0(.dout(w_dff_A_fk6lzoKa2_0),.din(w_dff_A_lVS80qA86_0),.clk(gclk));
	jdff dff_A_fk6lzoKa2_0(.dout(w_dff_A_BEdpB4C30_0),.din(w_dff_A_fk6lzoKa2_0),.clk(gclk));
	jdff dff_A_BEdpB4C30_0(.dout(w_dff_A_b1dLA96G0_0),.din(w_dff_A_BEdpB4C30_0),.clk(gclk));
	jdff dff_A_b1dLA96G0_0(.dout(w_dff_A_QR4EX62S0_0),.din(w_dff_A_b1dLA96G0_0),.clk(gclk));
	jdff dff_A_QR4EX62S0_0(.dout(w_dff_A_MFAyzbx46_0),.din(w_dff_A_QR4EX62S0_0),.clk(gclk));
	jdff dff_A_MFAyzbx46_0(.dout(w_dff_A_GVp1UVPk7_0),.din(w_dff_A_MFAyzbx46_0),.clk(gclk));
	jdff dff_A_GVp1UVPk7_0(.dout(w_dff_A_PM5ZtlQD7_0),.din(w_dff_A_GVp1UVPk7_0),.clk(gclk));
	jdff dff_A_PM5ZtlQD7_0(.dout(w_dff_A_2ycVZnh81_0),.din(w_dff_A_PM5ZtlQD7_0),.clk(gclk));
	jdff dff_A_2ycVZnh81_0(.dout(w_dff_A_tQit25iN5_0),.din(w_dff_A_2ycVZnh81_0),.clk(gclk));
	jdff dff_A_tQit25iN5_0(.dout(f47),.din(w_dff_A_tQit25iN5_0),.clk(gclk));
	jdff dff_A_aJxExRy15_2(.dout(w_dff_A_NJQV6SZi2_0),.din(w_dff_A_aJxExRy15_2),.clk(gclk));
	jdff dff_A_NJQV6SZi2_0(.dout(w_dff_A_MhBca7KV1_0),.din(w_dff_A_NJQV6SZi2_0),.clk(gclk));
	jdff dff_A_MhBca7KV1_0(.dout(w_dff_A_9OlWWsqQ2_0),.din(w_dff_A_MhBca7KV1_0),.clk(gclk));
	jdff dff_A_9OlWWsqQ2_0(.dout(w_dff_A_Zqv09oBS6_0),.din(w_dff_A_9OlWWsqQ2_0),.clk(gclk));
	jdff dff_A_Zqv09oBS6_0(.dout(w_dff_A_VVASM3SG2_0),.din(w_dff_A_Zqv09oBS6_0),.clk(gclk));
	jdff dff_A_VVASM3SG2_0(.dout(w_dff_A_YVPc6j3h6_0),.din(w_dff_A_VVASM3SG2_0),.clk(gclk));
	jdff dff_A_YVPc6j3h6_0(.dout(w_dff_A_0z8fme2q7_0),.din(w_dff_A_YVPc6j3h6_0),.clk(gclk));
	jdff dff_A_0z8fme2q7_0(.dout(w_dff_A_nGHTJf3E0_0),.din(w_dff_A_0z8fme2q7_0),.clk(gclk));
	jdff dff_A_nGHTJf3E0_0(.dout(w_dff_A_JdMdHrXo9_0),.din(w_dff_A_nGHTJf3E0_0),.clk(gclk));
	jdff dff_A_JdMdHrXo9_0(.dout(w_dff_A_CjQsWB2y3_0),.din(w_dff_A_JdMdHrXo9_0),.clk(gclk));
	jdff dff_A_CjQsWB2y3_0(.dout(w_dff_A_61ToQZPn3_0),.din(w_dff_A_CjQsWB2y3_0),.clk(gclk));
	jdff dff_A_61ToQZPn3_0(.dout(w_dff_A_7HDDk0Ny2_0),.din(w_dff_A_61ToQZPn3_0),.clk(gclk));
	jdff dff_A_7HDDk0Ny2_0(.dout(w_dff_A_CA81cROY1_0),.din(w_dff_A_7HDDk0Ny2_0),.clk(gclk));
	jdff dff_A_CA81cROY1_0(.dout(w_dff_A_jDJVLSTG9_0),.din(w_dff_A_CA81cROY1_0),.clk(gclk));
	jdff dff_A_jDJVLSTG9_0(.dout(w_dff_A_Dukm22Qj1_0),.din(w_dff_A_jDJVLSTG9_0),.clk(gclk));
	jdff dff_A_Dukm22Qj1_0(.dout(w_dff_A_5wF390iD5_0),.din(w_dff_A_Dukm22Qj1_0),.clk(gclk));
	jdff dff_A_5wF390iD5_0(.dout(w_dff_A_XGe4BT3r3_0),.din(w_dff_A_5wF390iD5_0),.clk(gclk));
	jdff dff_A_XGe4BT3r3_0(.dout(w_dff_A_RedMbgfE6_0),.din(w_dff_A_XGe4BT3r3_0),.clk(gclk));
	jdff dff_A_RedMbgfE6_0(.dout(w_dff_A_yORgae439_0),.din(w_dff_A_RedMbgfE6_0),.clk(gclk));
	jdff dff_A_yORgae439_0(.dout(w_dff_A_2c5OQJUM8_0),.din(w_dff_A_yORgae439_0),.clk(gclk));
	jdff dff_A_2c5OQJUM8_0(.dout(w_dff_A_uumfmRZn3_0),.din(w_dff_A_2c5OQJUM8_0),.clk(gclk));
	jdff dff_A_uumfmRZn3_0(.dout(w_dff_A_aAakDUJN0_0),.din(w_dff_A_uumfmRZn3_0),.clk(gclk));
	jdff dff_A_aAakDUJN0_0(.dout(w_dff_A_fl4wvd8T3_0),.din(w_dff_A_aAakDUJN0_0),.clk(gclk));
	jdff dff_A_fl4wvd8T3_0(.dout(w_dff_A_kQ5Oqr6u0_0),.din(w_dff_A_fl4wvd8T3_0),.clk(gclk));
	jdff dff_A_kQ5Oqr6u0_0(.dout(w_dff_A_lrb8EH9h7_0),.din(w_dff_A_kQ5Oqr6u0_0),.clk(gclk));
	jdff dff_A_lrb8EH9h7_0(.dout(w_dff_A_SBhgyTjs2_0),.din(w_dff_A_lrb8EH9h7_0),.clk(gclk));
	jdff dff_A_SBhgyTjs2_0(.dout(w_dff_A_zq4e2W0W9_0),.din(w_dff_A_SBhgyTjs2_0),.clk(gclk));
	jdff dff_A_zq4e2W0W9_0(.dout(w_dff_A_6gFVf2vb0_0),.din(w_dff_A_zq4e2W0W9_0),.clk(gclk));
	jdff dff_A_6gFVf2vb0_0(.dout(w_dff_A_VAGS6w1e8_0),.din(w_dff_A_6gFVf2vb0_0),.clk(gclk));
	jdff dff_A_VAGS6w1e8_0(.dout(w_dff_A_p8DQ8MmW0_0),.din(w_dff_A_VAGS6w1e8_0),.clk(gclk));
	jdff dff_A_p8DQ8MmW0_0(.dout(w_dff_A_SaFZpYw31_0),.din(w_dff_A_p8DQ8MmW0_0),.clk(gclk));
	jdff dff_A_SaFZpYw31_0(.dout(w_dff_A_2schEaM23_0),.din(w_dff_A_SaFZpYw31_0),.clk(gclk));
	jdff dff_A_2schEaM23_0(.dout(w_dff_A_WVuOI4ok0_0),.din(w_dff_A_2schEaM23_0),.clk(gclk));
	jdff dff_A_WVuOI4ok0_0(.dout(w_dff_A_ZAWf4ALq5_0),.din(w_dff_A_WVuOI4ok0_0),.clk(gclk));
	jdff dff_A_ZAWf4ALq5_0(.dout(w_dff_A_toFNROMF5_0),.din(w_dff_A_ZAWf4ALq5_0),.clk(gclk));
	jdff dff_A_toFNROMF5_0(.dout(w_dff_A_OL7lrtJo9_0),.din(w_dff_A_toFNROMF5_0),.clk(gclk));
	jdff dff_A_OL7lrtJo9_0(.dout(w_dff_A_FJXgFxuv3_0),.din(w_dff_A_OL7lrtJo9_0),.clk(gclk));
	jdff dff_A_FJXgFxuv3_0(.dout(w_dff_A_hnOh2mkZ4_0),.din(w_dff_A_FJXgFxuv3_0),.clk(gclk));
	jdff dff_A_hnOh2mkZ4_0(.dout(w_dff_A_fsZYiXue4_0),.din(w_dff_A_hnOh2mkZ4_0),.clk(gclk));
	jdff dff_A_fsZYiXue4_0(.dout(w_dff_A_i19eDR6q7_0),.din(w_dff_A_fsZYiXue4_0),.clk(gclk));
	jdff dff_A_i19eDR6q7_0(.dout(w_dff_A_f8MnNG2o7_0),.din(w_dff_A_i19eDR6q7_0),.clk(gclk));
	jdff dff_A_f8MnNG2o7_0(.dout(w_dff_A_Rc2w68Zs3_0),.din(w_dff_A_f8MnNG2o7_0),.clk(gclk));
	jdff dff_A_Rc2w68Zs3_0(.dout(w_dff_A_Ng4GBPnK8_0),.din(w_dff_A_Rc2w68Zs3_0),.clk(gclk));
	jdff dff_A_Ng4GBPnK8_0(.dout(w_dff_A_SZzkyurj3_0),.din(w_dff_A_Ng4GBPnK8_0),.clk(gclk));
	jdff dff_A_SZzkyurj3_0(.dout(w_dff_A_sTSzT9z68_0),.din(w_dff_A_SZzkyurj3_0),.clk(gclk));
	jdff dff_A_sTSzT9z68_0(.dout(w_dff_A_i1cHP5Pz3_0),.din(w_dff_A_sTSzT9z68_0),.clk(gclk));
	jdff dff_A_i1cHP5Pz3_0(.dout(w_dff_A_ZOeMV3mx5_0),.din(w_dff_A_i1cHP5Pz3_0),.clk(gclk));
	jdff dff_A_ZOeMV3mx5_0(.dout(w_dff_A_BVmgYYX16_0),.din(w_dff_A_ZOeMV3mx5_0),.clk(gclk));
	jdff dff_A_BVmgYYX16_0(.dout(w_dff_A_Dcy9FYHD4_0),.din(w_dff_A_BVmgYYX16_0),.clk(gclk));
	jdff dff_A_Dcy9FYHD4_0(.dout(w_dff_A_53TW0JYo5_0),.din(w_dff_A_Dcy9FYHD4_0),.clk(gclk));
	jdff dff_A_53TW0JYo5_0(.dout(w_dff_A_kD4t3t1u3_0),.din(w_dff_A_53TW0JYo5_0),.clk(gclk));
	jdff dff_A_kD4t3t1u3_0(.dout(w_dff_A_MjW4Y4X77_0),.din(w_dff_A_kD4t3t1u3_0),.clk(gclk));
	jdff dff_A_MjW4Y4X77_0(.dout(w_dff_A_jset7Hrp4_0),.din(w_dff_A_MjW4Y4X77_0),.clk(gclk));
	jdff dff_A_jset7Hrp4_0(.dout(w_dff_A_bo5hM1YX6_0),.din(w_dff_A_jset7Hrp4_0),.clk(gclk));
	jdff dff_A_bo5hM1YX6_0(.dout(w_dff_A_OeEAXBqx7_0),.din(w_dff_A_bo5hM1YX6_0),.clk(gclk));
	jdff dff_A_OeEAXBqx7_0(.dout(w_dff_A_gvOndYL90_0),.din(w_dff_A_OeEAXBqx7_0),.clk(gclk));
	jdff dff_A_gvOndYL90_0(.dout(w_dff_A_Sv6v8ZMG7_0),.din(w_dff_A_gvOndYL90_0),.clk(gclk));
	jdff dff_A_Sv6v8ZMG7_0(.dout(w_dff_A_SgPoUcIc4_0),.din(w_dff_A_Sv6v8ZMG7_0),.clk(gclk));
	jdff dff_A_SgPoUcIc4_0(.dout(w_dff_A_t5CxSU6p2_0),.din(w_dff_A_SgPoUcIc4_0),.clk(gclk));
	jdff dff_A_t5CxSU6p2_0(.dout(w_dff_A_2sxTJBzf2_0),.din(w_dff_A_t5CxSU6p2_0),.clk(gclk));
	jdff dff_A_2sxTJBzf2_0(.dout(w_dff_A_SCp9anKm5_0),.din(w_dff_A_2sxTJBzf2_0),.clk(gclk));
	jdff dff_A_SCp9anKm5_0(.dout(w_dff_A_SilJIt3L9_0),.din(w_dff_A_SCp9anKm5_0),.clk(gclk));
	jdff dff_A_SilJIt3L9_0(.dout(w_dff_A_jdVbzgzD8_0),.din(w_dff_A_SilJIt3L9_0),.clk(gclk));
	jdff dff_A_jdVbzgzD8_0(.dout(w_dff_A_Z2UORUHY9_0),.din(w_dff_A_jdVbzgzD8_0),.clk(gclk));
	jdff dff_A_Z2UORUHY9_0(.dout(w_dff_A_HV3OpqiV2_0),.din(w_dff_A_Z2UORUHY9_0),.clk(gclk));
	jdff dff_A_HV3OpqiV2_0(.dout(w_dff_A_sTbfWvpH0_0),.din(w_dff_A_HV3OpqiV2_0),.clk(gclk));
	jdff dff_A_sTbfWvpH0_0(.dout(w_dff_A_WIHKVHEv6_0),.din(w_dff_A_sTbfWvpH0_0),.clk(gclk));
	jdff dff_A_WIHKVHEv6_0(.dout(w_dff_A_vYxh0iqH1_0),.din(w_dff_A_WIHKVHEv6_0),.clk(gclk));
	jdff dff_A_vYxh0iqH1_0(.dout(w_dff_A_CKoeG2LA3_0),.din(w_dff_A_vYxh0iqH1_0),.clk(gclk));
	jdff dff_A_CKoeG2LA3_0(.dout(w_dff_A_Ajoa1CTr4_0),.din(w_dff_A_CKoeG2LA3_0),.clk(gclk));
	jdff dff_A_Ajoa1CTr4_0(.dout(w_dff_A_0E6OY1vP3_0),.din(w_dff_A_Ajoa1CTr4_0),.clk(gclk));
	jdff dff_A_0E6OY1vP3_0(.dout(w_dff_A_BSzPQ1cr8_0),.din(w_dff_A_0E6OY1vP3_0),.clk(gclk));
	jdff dff_A_BSzPQ1cr8_0(.dout(w_dff_A_GODjdHIs6_0),.din(w_dff_A_BSzPQ1cr8_0),.clk(gclk));
	jdff dff_A_GODjdHIs6_0(.dout(w_dff_A_vsh7Yx6j7_0),.din(w_dff_A_GODjdHIs6_0),.clk(gclk));
	jdff dff_A_vsh7Yx6j7_0(.dout(w_dff_A_iLtnmXgW9_0),.din(w_dff_A_vsh7Yx6j7_0),.clk(gclk));
	jdff dff_A_iLtnmXgW9_0(.dout(w_dff_A_tQSgV8Ht4_0),.din(w_dff_A_iLtnmXgW9_0),.clk(gclk));
	jdff dff_A_tQSgV8Ht4_0(.dout(w_dff_A_aDglIXsz2_0),.din(w_dff_A_tQSgV8Ht4_0),.clk(gclk));
	jdff dff_A_aDglIXsz2_0(.dout(w_dff_A_tpByKxB19_0),.din(w_dff_A_aDglIXsz2_0),.clk(gclk));
	jdff dff_A_tpByKxB19_0(.dout(f48),.din(w_dff_A_tpByKxB19_0),.clk(gclk));
	jdff dff_A_3mKSz1HS2_2(.dout(w_dff_A_Ayv7Ppx06_0),.din(w_dff_A_3mKSz1HS2_2),.clk(gclk));
	jdff dff_A_Ayv7Ppx06_0(.dout(w_dff_A_VRZQs1TI6_0),.din(w_dff_A_Ayv7Ppx06_0),.clk(gclk));
	jdff dff_A_VRZQs1TI6_0(.dout(w_dff_A_qsKJ5qbk2_0),.din(w_dff_A_VRZQs1TI6_0),.clk(gclk));
	jdff dff_A_qsKJ5qbk2_0(.dout(w_dff_A_1HZKPwpJ8_0),.din(w_dff_A_qsKJ5qbk2_0),.clk(gclk));
	jdff dff_A_1HZKPwpJ8_0(.dout(w_dff_A_dYhEOeAy8_0),.din(w_dff_A_1HZKPwpJ8_0),.clk(gclk));
	jdff dff_A_dYhEOeAy8_0(.dout(w_dff_A_RSd7YNyE2_0),.din(w_dff_A_dYhEOeAy8_0),.clk(gclk));
	jdff dff_A_RSd7YNyE2_0(.dout(w_dff_A_A9abrbx92_0),.din(w_dff_A_RSd7YNyE2_0),.clk(gclk));
	jdff dff_A_A9abrbx92_0(.dout(w_dff_A_Rf4Lq1LW1_0),.din(w_dff_A_A9abrbx92_0),.clk(gclk));
	jdff dff_A_Rf4Lq1LW1_0(.dout(w_dff_A_hjLywgXr8_0),.din(w_dff_A_Rf4Lq1LW1_0),.clk(gclk));
	jdff dff_A_hjLywgXr8_0(.dout(w_dff_A_ww7T9sFt0_0),.din(w_dff_A_hjLywgXr8_0),.clk(gclk));
	jdff dff_A_ww7T9sFt0_0(.dout(w_dff_A_rSdSHtaX5_0),.din(w_dff_A_ww7T9sFt0_0),.clk(gclk));
	jdff dff_A_rSdSHtaX5_0(.dout(w_dff_A_I55otHc79_0),.din(w_dff_A_rSdSHtaX5_0),.clk(gclk));
	jdff dff_A_I55otHc79_0(.dout(w_dff_A_m6HZRIDq8_0),.din(w_dff_A_I55otHc79_0),.clk(gclk));
	jdff dff_A_m6HZRIDq8_0(.dout(w_dff_A_0GsZJ3Mb8_0),.din(w_dff_A_m6HZRIDq8_0),.clk(gclk));
	jdff dff_A_0GsZJ3Mb8_0(.dout(w_dff_A_0pK4sGkm1_0),.din(w_dff_A_0GsZJ3Mb8_0),.clk(gclk));
	jdff dff_A_0pK4sGkm1_0(.dout(w_dff_A_hyf7lwvX0_0),.din(w_dff_A_0pK4sGkm1_0),.clk(gclk));
	jdff dff_A_hyf7lwvX0_0(.dout(w_dff_A_HvcpWl597_0),.din(w_dff_A_hyf7lwvX0_0),.clk(gclk));
	jdff dff_A_HvcpWl597_0(.dout(w_dff_A_rJki5nAi1_0),.din(w_dff_A_HvcpWl597_0),.clk(gclk));
	jdff dff_A_rJki5nAi1_0(.dout(w_dff_A_9VJqhq2B5_0),.din(w_dff_A_rJki5nAi1_0),.clk(gclk));
	jdff dff_A_9VJqhq2B5_0(.dout(w_dff_A_BdMtPa6c2_0),.din(w_dff_A_9VJqhq2B5_0),.clk(gclk));
	jdff dff_A_BdMtPa6c2_0(.dout(w_dff_A_NZQ6XDaE5_0),.din(w_dff_A_BdMtPa6c2_0),.clk(gclk));
	jdff dff_A_NZQ6XDaE5_0(.dout(w_dff_A_JptcqQKJ8_0),.din(w_dff_A_NZQ6XDaE5_0),.clk(gclk));
	jdff dff_A_JptcqQKJ8_0(.dout(w_dff_A_LqMDoJNm5_0),.din(w_dff_A_JptcqQKJ8_0),.clk(gclk));
	jdff dff_A_LqMDoJNm5_0(.dout(w_dff_A_q90xRDts9_0),.din(w_dff_A_LqMDoJNm5_0),.clk(gclk));
	jdff dff_A_q90xRDts9_0(.dout(w_dff_A_TpJpQaKf0_0),.din(w_dff_A_q90xRDts9_0),.clk(gclk));
	jdff dff_A_TpJpQaKf0_0(.dout(w_dff_A_orumTqvT2_0),.din(w_dff_A_TpJpQaKf0_0),.clk(gclk));
	jdff dff_A_orumTqvT2_0(.dout(w_dff_A_7xJ4e79C4_0),.din(w_dff_A_orumTqvT2_0),.clk(gclk));
	jdff dff_A_7xJ4e79C4_0(.dout(w_dff_A_5B6tToZH1_0),.din(w_dff_A_7xJ4e79C4_0),.clk(gclk));
	jdff dff_A_5B6tToZH1_0(.dout(w_dff_A_qYJIAWMz3_0),.din(w_dff_A_5B6tToZH1_0),.clk(gclk));
	jdff dff_A_qYJIAWMz3_0(.dout(w_dff_A_xHpIpZJQ9_0),.din(w_dff_A_qYJIAWMz3_0),.clk(gclk));
	jdff dff_A_xHpIpZJQ9_0(.dout(w_dff_A_4qI47ELd3_0),.din(w_dff_A_xHpIpZJQ9_0),.clk(gclk));
	jdff dff_A_4qI47ELd3_0(.dout(w_dff_A_aEUSdggI8_0),.din(w_dff_A_4qI47ELd3_0),.clk(gclk));
	jdff dff_A_aEUSdggI8_0(.dout(w_dff_A_9MjpSZ2L5_0),.din(w_dff_A_aEUSdggI8_0),.clk(gclk));
	jdff dff_A_9MjpSZ2L5_0(.dout(w_dff_A_mJdFMrsI5_0),.din(w_dff_A_9MjpSZ2L5_0),.clk(gclk));
	jdff dff_A_mJdFMrsI5_0(.dout(w_dff_A_GVM2uqUo8_0),.din(w_dff_A_mJdFMrsI5_0),.clk(gclk));
	jdff dff_A_GVM2uqUo8_0(.dout(w_dff_A_FCk9xpC88_0),.din(w_dff_A_GVM2uqUo8_0),.clk(gclk));
	jdff dff_A_FCk9xpC88_0(.dout(w_dff_A_yVTWZZlE3_0),.din(w_dff_A_FCk9xpC88_0),.clk(gclk));
	jdff dff_A_yVTWZZlE3_0(.dout(w_dff_A_BwnN4wyZ6_0),.din(w_dff_A_yVTWZZlE3_0),.clk(gclk));
	jdff dff_A_BwnN4wyZ6_0(.dout(w_dff_A_zsLCgcyH6_0),.din(w_dff_A_BwnN4wyZ6_0),.clk(gclk));
	jdff dff_A_zsLCgcyH6_0(.dout(w_dff_A_QJ9RmIWD8_0),.din(w_dff_A_zsLCgcyH6_0),.clk(gclk));
	jdff dff_A_QJ9RmIWD8_0(.dout(w_dff_A_CnvvP1RT2_0),.din(w_dff_A_QJ9RmIWD8_0),.clk(gclk));
	jdff dff_A_CnvvP1RT2_0(.dout(w_dff_A_lloiz32N1_0),.din(w_dff_A_CnvvP1RT2_0),.clk(gclk));
	jdff dff_A_lloiz32N1_0(.dout(w_dff_A_pmP8KUow4_0),.din(w_dff_A_lloiz32N1_0),.clk(gclk));
	jdff dff_A_pmP8KUow4_0(.dout(w_dff_A_FPm68tqi3_0),.din(w_dff_A_pmP8KUow4_0),.clk(gclk));
	jdff dff_A_FPm68tqi3_0(.dout(w_dff_A_PuULeQOX4_0),.din(w_dff_A_FPm68tqi3_0),.clk(gclk));
	jdff dff_A_PuULeQOX4_0(.dout(w_dff_A_oVV6jfYC5_0),.din(w_dff_A_PuULeQOX4_0),.clk(gclk));
	jdff dff_A_oVV6jfYC5_0(.dout(w_dff_A_F38qtnoU0_0),.din(w_dff_A_oVV6jfYC5_0),.clk(gclk));
	jdff dff_A_F38qtnoU0_0(.dout(w_dff_A_QboQC8Am2_0),.din(w_dff_A_F38qtnoU0_0),.clk(gclk));
	jdff dff_A_QboQC8Am2_0(.dout(w_dff_A_nG0DJOaO2_0),.din(w_dff_A_QboQC8Am2_0),.clk(gclk));
	jdff dff_A_nG0DJOaO2_0(.dout(w_dff_A_J4pwPtEZ7_0),.din(w_dff_A_nG0DJOaO2_0),.clk(gclk));
	jdff dff_A_J4pwPtEZ7_0(.dout(w_dff_A_L3RBCFh35_0),.din(w_dff_A_J4pwPtEZ7_0),.clk(gclk));
	jdff dff_A_L3RBCFh35_0(.dout(w_dff_A_hIz7n9vM4_0),.din(w_dff_A_L3RBCFh35_0),.clk(gclk));
	jdff dff_A_hIz7n9vM4_0(.dout(w_dff_A_AbiGTZzy0_0),.din(w_dff_A_hIz7n9vM4_0),.clk(gclk));
	jdff dff_A_AbiGTZzy0_0(.dout(w_dff_A_Qbl7wfZu4_0),.din(w_dff_A_AbiGTZzy0_0),.clk(gclk));
	jdff dff_A_Qbl7wfZu4_0(.dout(w_dff_A_r6IAGJNV0_0),.din(w_dff_A_Qbl7wfZu4_0),.clk(gclk));
	jdff dff_A_r6IAGJNV0_0(.dout(w_dff_A_5tez9fPY8_0),.din(w_dff_A_r6IAGJNV0_0),.clk(gclk));
	jdff dff_A_5tez9fPY8_0(.dout(w_dff_A_4Rk2jIV46_0),.din(w_dff_A_5tez9fPY8_0),.clk(gclk));
	jdff dff_A_4Rk2jIV46_0(.dout(w_dff_A_WKEXg25Z4_0),.din(w_dff_A_4Rk2jIV46_0),.clk(gclk));
	jdff dff_A_WKEXg25Z4_0(.dout(w_dff_A_VU38RyNS6_0),.din(w_dff_A_WKEXg25Z4_0),.clk(gclk));
	jdff dff_A_VU38RyNS6_0(.dout(w_dff_A_EiwL64n56_0),.din(w_dff_A_VU38RyNS6_0),.clk(gclk));
	jdff dff_A_EiwL64n56_0(.dout(w_dff_A_uhc33KPv8_0),.din(w_dff_A_EiwL64n56_0),.clk(gclk));
	jdff dff_A_uhc33KPv8_0(.dout(w_dff_A_JwDn17xS7_0),.din(w_dff_A_uhc33KPv8_0),.clk(gclk));
	jdff dff_A_JwDn17xS7_0(.dout(w_dff_A_2U74uBbJ9_0),.din(w_dff_A_JwDn17xS7_0),.clk(gclk));
	jdff dff_A_2U74uBbJ9_0(.dout(w_dff_A_rpX69VDC6_0),.din(w_dff_A_2U74uBbJ9_0),.clk(gclk));
	jdff dff_A_rpX69VDC6_0(.dout(w_dff_A_E4GIdYLV5_0),.din(w_dff_A_rpX69VDC6_0),.clk(gclk));
	jdff dff_A_E4GIdYLV5_0(.dout(w_dff_A_6WTvRgv09_0),.din(w_dff_A_E4GIdYLV5_0),.clk(gclk));
	jdff dff_A_6WTvRgv09_0(.dout(w_dff_A_4Yw9ASMd9_0),.din(w_dff_A_6WTvRgv09_0),.clk(gclk));
	jdff dff_A_4Yw9ASMd9_0(.dout(w_dff_A_gzOCrBSk3_0),.din(w_dff_A_4Yw9ASMd9_0),.clk(gclk));
	jdff dff_A_gzOCrBSk3_0(.dout(w_dff_A_6EzLwRpF3_0),.din(w_dff_A_gzOCrBSk3_0),.clk(gclk));
	jdff dff_A_6EzLwRpF3_0(.dout(w_dff_A_Jaj8X0jw9_0),.din(w_dff_A_6EzLwRpF3_0),.clk(gclk));
	jdff dff_A_Jaj8X0jw9_0(.dout(w_dff_A_rwzbeZNn0_0),.din(w_dff_A_Jaj8X0jw9_0),.clk(gclk));
	jdff dff_A_rwzbeZNn0_0(.dout(w_dff_A_b67luegq1_0),.din(w_dff_A_rwzbeZNn0_0),.clk(gclk));
	jdff dff_A_b67luegq1_0(.dout(w_dff_A_MC6t3PqP5_0),.din(w_dff_A_b67luegq1_0),.clk(gclk));
	jdff dff_A_MC6t3PqP5_0(.dout(w_dff_A_NqoWYY8r9_0),.din(w_dff_A_MC6t3PqP5_0),.clk(gclk));
	jdff dff_A_NqoWYY8r9_0(.dout(w_dff_A_MIjE16wO4_0),.din(w_dff_A_NqoWYY8r9_0),.clk(gclk));
	jdff dff_A_MIjE16wO4_0(.dout(w_dff_A_P2YgcVvb8_0),.din(w_dff_A_MIjE16wO4_0),.clk(gclk));
	jdff dff_A_P2YgcVvb8_0(.dout(w_dff_A_Tr8mwIHU2_0),.din(w_dff_A_P2YgcVvb8_0),.clk(gclk));
	jdff dff_A_Tr8mwIHU2_0(.dout(f49),.din(w_dff_A_Tr8mwIHU2_0),.clk(gclk));
	jdff dff_A_s2adAl7P4_2(.dout(w_dff_A_p9e74CQN8_0),.din(w_dff_A_s2adAl7P4_2),.clk(gclk));
	jdff dff_A_p9e74CQN8_0(.dout(w_dff_A_nPiZY0MH4_0),.din(w_dff_A_p9e74CQN8_0),.clk(gclk));
	jdff dff_A_nPiZY0MH4_0(.dout(w_dff_A_dzEbedML5_0),.din(w_dff_A_nPiZY0MH4_0),.clk(gclk));
	jdff dff_A_dzEbedML5_0(.dout(w_dff_A_NOpDgdU14_0),.din(w_dff_A_dzEbedML5_0),.clk(gclk));
	jdff dff_A_NOpDgdU14_0(.dout(w_dff_A_lXzMcDau3_0),.din(w_dff_A_NOpDgdU14_0),.clk(gclk));
	jdff dff_A_lXzMcDau3_0(.dout(w_dff_A_VYRVjvVu5_0),.din(w_dff_A_lXzMcDau3_0),.clk(gclk));
	jdff dff_A_VYRVjvVu5_0(.dout(w_dff_A_xGtHPyAS5_0),.din(w_dff_A_VYRVjvVu5_0),.clk(gclk));
	jdff dff_A_xGtHPyAS5_0(.dout(w_dff_A_w1U5qlyc9_0),.din(w_dff_A_xGtHPyAS5_0),.clk(gclk));
	jdff dff_A_w1U5qlyc9_0(.dout(w_dff_A_E43w3Iwf1_0),.din(w_dff_A_w1U5qlyc9_0),.clk(gclk));
	jdff dff_A_E43w3Iwf1_0(.dout(w_dff_A_OqgKUni50_0),.din(w_dff_A_E43w3Iwf1_0),.clk(gclk));
	jdff dff_A_OqgKUni50_0(.dout(w_dff_A_aIvvBTVq1_0),.din(w_dff_A_OqgKUni50_0),.clk(gclk));
	jdff dff_A_aIvvBTVq1_0(.dout(w_dff_A_lodkKEjr8_0),.din(w_dff_A_aIvvBTVq1_0),.clk(gclk));
	jdff dff_A_lodkKEjr8_0(.dout(w_dff_A_1oWgng8M0_0),.din(w_dff_A_lodkKEjr8_0),.clk(gclk));
	jdff dff_A_1oWgng8M0_0(.dout(w_dff_A_Mt25iuGA4_0),.din(w_dff_A_1oWgng8M0_0),.clk(gclk));
	jdff dff_A_Mt25iuGA4_0(.dout(w_dff_A_uamHzhzN6_0),.din(w_dff_A_Mt25iuGA4_0),.clk(gclk));
	jdff dff_A_uamHzhzN6_0(.dout(w_dff_A_3t3oRcwu8_0),.din(w_dff_A_uamHzhzN6_0),.clk(gclk));
	jdff dff_A_3t3oRcwu8_0(.dout(w_dff_A_P9yYoLt63_0),.din(w_dff_A_3t3oRcwu8_0),.clk(gclk));
	jdff dff_A_P9yYoLt63_0(.dout(w_dff_A_iuz09znQ0_0),.din(w_dff_A_P9yYoLt63_0),.clk(gclk));
	jdff dff_A_iuz09znQ0_0(.dout(w_dff_A_eMwdA4SH8_0),.din(w_dff_A_iuz09znQ0_0),.clk(gclk));
	jdff dff_A_eMwdA4SH8_0(.dout(w_dff_A_axXOLZgR8_0),.din(w_dff_A_eMwdA4SH8_0),.clk(gclk));
	jdff dff_A_axXOLZgR8_0(.dout(w_dff_A_9X9chWfX8_0),.din(w_dff_A_axXOLZgR8_0),.clk(gclk));
	jdff dff_A_9X9chWfX8_0(.dout(w_dff_A_DYOmGE027_0),.din(w_dff_A_9X9chWfX8_0),.clk(gclk));
	jdff dff_A_DYOmGE027_0(.dout(w_dff_A_J8qY0DHt8_0),.din(w_dff_A_DYOmGE027_0),.clk(gclk));
	jdff dff_A_J8qY0DHt8_0(.dout(w_dff_A_3Lz4mhlJ9_0),.din(w_dff_A_J8qY0DHt8_0),.clk(gclk));
	jdff dff_A_3Lz4mhlJ9_0(.dout(w_dff_A_UMUx6kGP8_0),.din(w_dff_A_3Lz4mhlJ9_0),.clk(gclk));
	jdff dff_A_UMUx6kGP8_0(.dout(w_dff_A_mNB4LWA62_0),.din(w_dff_A_UMUx6kGP8_0),.clk(gclk));
	jdff dff_A_mNB4LWA62_0(.dout(w_dff_A_0cpTtEaZ6_0),.din(w_dff_A_mNB4LWA62_0),.clk(gclk));
	jdff dff_A_0cpTtEaZ6_0(.dout(w_dff_A_VLKZEIgi1_0),.din(w_dff_A_0cpTtEaZ6_0),.clk(gclk));
	jdff dff_A_VLKZEIgi1_0(.dout(w_dff_A_ftD70KiW2_0),.din(w_dff_A_VLKZEIgi1_0),.clk(gclk));
	jdff dff_A_ftD70KiW2_0(.dout(w_dff_A_76xFgNlE8_0),.din(w_dff_A_ftD70KiW2_0),.clk(gclk));
	jdff dff_A_76xFgNlE8_0(.dout(w_dff_A_7okjH4Kb2_0),.din(w_dff_A_76xFgNlE8_0),.clk(gclk));
	jdff dff_A_7okjH4Kb2_0(.dout(w_dff_A_fxSkxYUh1_0),.din(w_dff_A_7okjH4Kb2_0),.clk(gclk));
	jdff dff_A_fxSkxYUh1_0(.dout(w_dff_A_wST5657d5_0),.din(w_dff_A_fxSkxYUh1_0),.clk(gclk));
	jdff dff_A_wST5657d5_0(.dout(w_dff_A_nBRekPHZ8_0),.din(w_dff_A_wST5657d5_0),.clk(gclk));
	jdff dff_A_nBRekPHZ8_0(.dout(w_dff_A_mb2ngAR64_0),.din(w_dff_A_nBRekPHZ8_0),.clk(gclk));
	jdff dff_A_mb2ngAR64_0(.dout(w_dff_A_5KIViX3l8_0),.din(w_dff_A_mb2ngAR64_0),.clk(gclk));
	jdff dff_A_5KIViX3l8_0(.dout(w_dff_A_AGWHZpDO6_0),.din(w_dff_A_5KIViX3l8_0),.clk(gclk));
	jdff dff_A_AGWHZpDO6_0(.dout(w_dff_A_zMLwvWqH8_0),.din(w_dff_A_AGWHZpDO6_0),.clk(gclk));
	jdff dff_A_zMLwvWqH8_0(.dout(w_dff_A_qd6bs8PP5_0),.din(w_dff_A_zMLwvWqH8_0),.clk(gclk));
	jdff dff_A_qd6bs8PP5_0(.dout(w_dff_A_P2Ro2ra41_0),.din(w_dff_A_qd6bs8PP5_0),.clk(gclk));
	jdff dff_A_P2Ro2ra41_0(.dout(w_dff_A_2xv3eXLA9_0),.din(w_dff_A_P2Ro2ra41_0),.clk(gclk));
	jdff dff_A_2xv3eXLA9_0(.dout(w_dff_A_Mnry7XKU8_0),.din(w_dff_A_2xv3eXLA9_0),.clk(gclk));
	jdff dff_A_Mnry7XKU8_0(.dout(w_dff_A_Nxp6sLEB9_0),.din(w_dff_A_Mnry7XKU8_0),.clk(gclk));
	jdff dff_A_Nxp6sLEB9_0(.dout(w_dff_A_2Ad0xBuh4_0),.din(w_dff_A_Nxp6sLEB9_0),.clk(gclk));
	jdff dff_A_2Ad0xBuh4_0(.dout(w_dff_A_PlYmFzEy7_0),.din(w_dff_A_2Ad0xBuh4_0),.clk(gclk));
	jdff dff_A_PlYmFzEy7_0(.dout(w_dff_A_xgwGsZFZ7_0),.din(w_dff_A_PlYmFzEy7_0),.clk(gclk));
	jdff dff_A_xgwGsZFZ7_0(.dout(w_dff_A_3yhwGmLo8_0),.din(w_dff_A_xgwGsZFZ7_0),.clk(gclk));
	jdff dff_A_3yhwGmLo8_0(.dout(w_dff_A_Vz30GvIZ3_0),.din(w_dff_A_3yhwGmLo8_0),.clk(gclk));
	jdff dff_A_Vz30GvIZ3_0(.dout(w_dff_A_7DQC3X7E3_0),.din(w_dff_A_Vz30GvIZ3_0),.clk(gclk));
	jdff dff_A_7DQC3X7E3_0(.dout(w_dff_A_zb6EAGno7_0),.din(w_dff_A_7DQC3X7E3_0),.clk(gclk));
	jdff dff_A_zb6EAGno7_0(.dout(w_dff_A_RPUJQJwf1_0),.din(w_dff_A_zb6EAGno7_0),.clk(gclk));
	jdff dff_A_RPUJQJwf1_0(.dout(w_dff_A_Wfq44m7z6_0),.din(w_dff_A_RPUJQJwf1_0),.clk(gclk));
	jdff dff_A_Wfq44m7z6_0(.dout(w_dff_A_2P7uytly9_0),.din(w_dff_A_Wfq44m7z6_0),.clk(gclk));
	jdff dff_A_2P7uytly9_0(.dout(w_dff_A_XfE6Rlyr3_0),.din(w_dff_A_2P7uytly9_0),.clk(gclk));
	jdff dff_A_XfE6Rlyr3_0(.dout(w_dff_A_xDalQPYM0_0),.din(w_dff_A_XfE6Rlyr3_0),.clk(gclk));
	jdff dff_A_xDalQPYM0_0(.dout(w_dff_A_OtFyS5E27_0),.din(w_dff_A_xDalQPYM0_0),.clk(gclk));
	jdff dff_A_OtFyS5E27_0(.dout(w_dff_A_pIqfvuvg1_0),.din(w_dff_A_OtFyS5E27_0),.clk(gclk));
	jdff dff_A_pIqfvuvg1_0(.dout(w_dff_A_aTfSc5CN2_0),.din(w_dff_A_pIqfvuvg1_0),.clk(gclk));
	jdff dff_A_aTfSc5CN2_0(.dout(w_dff_A_unE3wgMZ3_0),.din(w_dff_A_aTfSc5CN2_0),.clk(gclk));
	jdff dff_A_unE3wgMZ3_0(.dout(w_dff_A_vs8e6brq8_0),.din(w_dff_A_unE3wgMZ3_0),.clk(gclk));
	jdff dff_A_vs8e6brq8_0(.dout(w_dff_A_IoCGsAx39_0),.din(w_dff_A_vs8e6brq8_0),.clk(gclk));
	jdff dff_A_IoCGsAx39_0(.dout(w_dff_A_TPugt1ud5_0),.din(w_dff_A_IoCGsAx39_0),.clk(gclk));
	jdff dff_A_TPugt1ud5_0(.dout(w_dff_A_RoiPUm8A4_0),.din(w_dff_A_TPugt1ud5_0),.clk(gclk));
	jdff dff_A_RoiPUm8A4_0(.dout(w_dff_A_wBzyuGAx4_0),.din(w_dff_A_RoiPUm8A4_0),.clk(gclk));
	jdff dff_A_wBzyuGAx4_0(.dout(w_dff_A_ZzMkZ7tJ5_0),.din(w_dff_A_wBzyuGAx4_0),.clk(gclk));
	jdff dff_A_ZzMkZ7tJ5_0(.dout(w_dff_A_gi9R00dn4_0),.din(w_dff_A_ZzMkZ7tJ5_0),.clk(gclk));
	jdff dff_A_gi9R00dn4_0(.dout(w_dff_A_jT6H4wEd8_0),.din(w_dff_A_gi9R00dn4_0),.clk(gclk));
	jdff dff_A_jT6H4wEd8_0(.dout(w_dff_A_c5sFRDUV9_0),.din(w_dff_A_jT6H4wEd8_0),.clk(gclk));
	jdff dff_A_c5sFRDUV9_0(.dout(w_dff_A_4QgCc8kE3_0),.din(w_dff_A_c5sFRDUV9_0),.clk(gclk));
	jdff dff_A_4QgCc8kE3_0(.dout(w_dff_A_maY7meEX3_0),.din(w_dff_A_4QgCc8kE3_0),.clk(gclk));
	jdff dff_A_maY7meEX3_0(.dout(w_dff_A_SmiJYLCg8_0),.din(w_dff_A_maY7meEX3_0),.clk(gclk));
	jdff dff_A_SmiJYLCg8_0(.dout(w_dff_A_WAI2As8U6_0),.din(w_dff_A_SmiJYLCg8_0),.clk(gclk));
	jdff dff_A_WAI2As8U6_0(.dout(w_dff_A_cg1LW6JN5_0),.din(w_dff_A_WAI2As8U6_0),.clk(gclk));
	jdff dff_A_cg1LW6JN5_0(.dout(w_dff_A_fLyeR8lw5_0),.din(w_dff_A_cg1LW6JN5_0),.clk(gclk));
	jdff dff_A_fLyeR8lw5_0(.dout(w_dff_A_msZXrXJB8_0),.din(w_dff_A_fLyeR8lw5_0),.clk(gclk));
	jdff dff_A_msZXrXJB8_0(.dout(w_dff_A_1EaWz1YO0_0),.din(w_dff_A_msZXrXJB8_0),.clk(gclk));
	jdff dff_A_1EaWz1YO0_0(.dout(f50),.din(w_dff_A_1EaWz1YO0_0),.clk(gclk));
	jdff dff_A_FVUuRbF61_2(.dout(w_dff_A_za6uKTJo8_0),.din(w_dff_A_FVUuRbF61_2),.clk(gclk));
	jdff dff_A_za6uKTJo8_0(.dout(w_dff_A_C1vBaGHQ0_0),.din(w_dff_A_za6uKTJo8_0),.clk(gclk));
	jdff dff_A_C1vBaGHQ0_0(.dout(w_dff_A_yy1oYe0Q9_0),.din(w_dff_A_C1vBaGHQ0_0),.clk(gclk));
	jdff dff_A_yy1oYe0Q9_0(.dout(w_dff_A_Ka45KprM5_0),.din(w_dff_A_yy1oYe0Q9_0),.clk(gclk));
	jdff dff_A_Ka45KprM5_0(.dout(w_dff_A_1v5LnPC65_0),.din(w_dff_A_Ka45KprM5_0),.clk(gclk));
	jdff dff_A_1v5LnPC65_0(.dout(w_dff_A_99xxFQsX7_0),.din(w_dff_A_1v5LnPC65_0),.clk(gclk));
	jdff dff_A_99xxFQsX7_0(.dout(w_dff_A_0V0sCq0t5_0),.din(w_dff_A_99xxFQsX7_0),.clk(gclk));
	jdff dff_A_0V0sCq0t5_0(.dout(w_dff_A_xRnN0fqv0_0),.din(w_dff_A_0V0sCq0t5_0),.clk(gclk));
	jdff dff_A_xRnN0fqv0_0(.dout(w_dff_A_3w4Bxij31_0),.din(w_dff_A_xRnN0fqv0_0),.clk(gclk));
	jdff dff_A_3w4Bxij31_0(.dout(w_dff_A_y8L2Rgy94_0),.din(w_dff_A_3w4Bxij31_0),.clk(gclk));
	jdff dff_A_y8L2Rgy94_0(.dout(w_dff_A_bHjadYxX0_0),.din(w_dff_A_y8L2Rgy94_0),.clk(gclk));
	jdff dff_A_bHjadYxX0_0(.dout(w_dff_A_vwBaucBK1_0),.din(w_dff_A_bHjadYxX0_0),.clk(gclk));
	jdff dff_A_vwBaucBK1_0(.dout(w_dff_A_hRggI1r32_0),.din(w_dff_A_vwBaucBK1_0),.clk(gclk));
	jdff dff_A_hRggI1r32_0(.dout(w_dff_A_SpUHXYxh5_0),.din(w_dff_A_hRggI1r32_0),.clk(gclk));
	jdff dff_A_SpUHXYxh5_0(.dout(w_dff_A_OZDyMNbJ0_0),.din(w_dff_A_SpUHXYxh5_0),.clk(gclk));
	jdff dff_A_OZDyMNbJ0_0(.dout(w_dff_A_hscaPDxD1_0),.din(w_dff_A_OZDyMNbJ0_0),.clk(gclk));
	jdff dff_A_hscaPDxD1_0(.dout(w_dff_A_oIPBw6n24_0),.din(w_dff_A_hscaPDxD1_0),.clk(gclk));
	jdff dff_A_oIPBw6n24_0(.dout(w_dff_A_ZrTDPSko0_0),.din(w_dff_A_oIPBw6n24_0),.clk(gclk));
	jdff dff_A_ZrTDPSko0_0(.dout(w_dff_A_jISupvsL9_0),.din(w_dff_A_ZrTDPSko0_0),.clk(gclk));
	jdff dff_A_jISupvsL9_0(.dout(w_dff_A_Z6Wte2wt5_0),.din(w_dff_A_jISupvsL9_0),.clk(gclk));
	jdff dff_A_Z6Wte2wt5_0(.dout(w_dff_A_DMbG3TAN0_0),.din(w_dff_A_Z6Wte2wt5_0),.clk(gclk));
	jdff dff_A_DMbG3TAN0_0(.dout(w_dff_A_ty99He0M5_0),.din(w_dff_A_DMbG3TAN0_0),.clk(gclk));
	jdff dff_A_ty99He0M5_0(.dout(w_dff_A_FpQrcYFN9_0),.din(w_dff_A_ty99He0M5_0),.clk(gclk));
	jdff dff_A_FpQrcYFN9_0(.dout(w_dff_A_eTyRV7Uv1_0),.din(w_dff_A_FpQrcYFN9_0),.clk(gclk));
	jdff dff_A_eTyRV7Uv1_0(.dout(w_dff_A_9tQgvxoD1_0),.din(w_dff_A_eTyRV7Uv1_0),.clk(gclk));
	jdff dff_A_9tQgvxoD1_0(.dout(w_dff_A_uKFy8WHt6_0),.din(w_dff_A_9tQgvxoD1_0),.clk(gclk));
	jdff dff_A_uKFy8WHt6_0(.dout(w_dff_A_FaUFIllK8_0),.din(w_dff_A_uKFy8WHt6_0),.clk(gclk));
	jdff dff_A_FaUFIllK8_0(.dout(w_dff_A_r3Jz7kyX5_0),.din(w_dff_A_FaUFIllK8_0),.clk(gclk));
	jdff dff_A_r3Jz7kyX5_0(.dout(w_dff_A_DPpqnHGu3_0),.din(w_dff_A_r3Jz7kyX5_0),.clk(gclk));
	jdff dff_A_DPpqnHGu3_0(.dout(w_dff_A_sJ8FYyXE7_0),.din(w_dff_A_DPpqnHGu3_0),.clk(gclk));
	jdff dff_A_sJ8FYyXE7_0(.dout(w_dff_A_fkBJLsLl2_0),.din(w_dff_A_sJ8FYyXE7_0),.clk(gclk));
	jdff dff_A_fkBJLsLl2_0(.dout(w_dff_A_uInRUfya7_0),.din(w_dff_A_fkBJLsLl2_0),.clk(gclk));
	jdff dff_A_uInRUfya7_0(.dout(w_dff_A_AZHjDvnt3_0),.din(w_dff_A_uInRUfya7_0),.clk(gclk));
	jdff dff_A_AZHjDvnt3_0(.dout(w_dff_A_LFFSWndL4_0),.din(w_dff_A_AZHjDvnt3_0),.clk(gclk));
	jdff dff_A_LFFSWndL4_0(.dout(w_dff_A_uwP9rW7q0_0),.din(w_dff_A_LFFSWndL4_0),.clk(gclk));
	jdff dff_A_uwP9rW7q0_0(.dout(w_dff_A_iTMrYELx1_0),.din(w_dff_A_uwP9rW7q0_0),.clk(gclk));
	jdff dff_A_iTMrYELx1_0(.dout(w_dff_A_dKru4FVS3_0),.din(w_dff_A_iTMrYELx1_0),.clk(gclk));
	jdff dff_A_dKru4FVS3_0(.dout(w_dff_A_gc6PomZM1_0),.din(w_dff_A_dKru4FVS3_0),.clk(gclk));
	jdff dff_A_gc6PomZM1_0(.dout(w_dff_A_wgS1mZES9_0),.din(w_dff_A_gc6PomZM1_0),.clk(gclk));
	jdff dff_A_wgS1mZES9_0(.dout(w_dff_A_A7ogKbe88_0),.din(w_dff_A_wgS1mZES9_0),.clk(gclk));
	jdff dff_A_A7ogKbe88_0(.dout(w_dff_A_GGEAhZFD1_0),.din(w_dff_A_A7ogKbe88_0),.clk(gclk));
	jdff dff_A_GGEAhZFD1_0(.dout(w_dff_A_EMU3bqyG5_0),.din(w_dff_A_GGEAhZFD1_0),.clk(gclk));
	jdff dff_A_EMU3bqyG5_0(.dout(w_dff_A_sZdgB3DU9_0),.din(w_dff_A_EMU3bqyG5_0),.clk(gclk));
	jdff dff_A_sZdgB3DU9_0(.dout(w_dff_A_qh8CFvTP9_0),.din(w_dff_A_sZdgB3DU9_0),.clk(gclk));
	jdff dff_A_qh8CFvTP9_0(.dout(w_dff_A_Oa0Eoz0O7_0),.din(w_dff_A_qh8CFvTP9_0),.clk(gclk));
	jdff dff_A_Oa0Eoz0O7_0(.dout(w_dff_A_F4vtuYJg5_0),.din(w_dff_A_Oa0Eoz0O7_0),.clk(gclk));
	jdff dff_A_F4vtuYJg5_0(.dout(w_dff_A_C1QnvXea3_0),.din(w_dff_A_F4vtuYJg5_0),.clk(gclk));
	jdff dff_A_C1QnvXea3_0(.dout(w_dff_A_Z0XmoKy22_0),.din(w_dff_A_C1QnvXea3_0),.clk(gclk));
	jdff dff_A_Z0XmoKy22_0(.dout(w_dff_A_mLieapSf5_0),.din(w_dff_A_Z0XmoKy22_0),.clk(gclk));
	jdff dff_A_mLieapSf5_0(.dout(w_dff_A_wki21UKd6_0),.din(w_dff_A_mLieapSf5_0),.clk(gclk));
	jdff dff_A_wki21UKd6_0(.dout(w_dff_A_V2QxSvUa3_0),.din(w_dff_A_wki21UKd6_0),.clk(gclk));
	jdff dff_A_V2QxSvUa3_0(.dout(w_dff_A_3SMUQ99Y2_0),.din(w_dff_A_V2QxSvUa3_0),.clk(gclk));
	jdff dff_A_3SMUQ99Y2_0(.dout(w_dff_A_NTZvkYIE1_0),.din(w_dff_A_3SMUQ99Y2_0),.clk(gclk));
	jdff dff_A_NTZvkYIE1_0(.dout(w_dff_A_v6gqwMek3_0),.din(w_dff_A_NTZvkYIE1_0),.clk(gclk));
	jdff dff_A_v6gqwMek3_0(.dout(w_dff_A_P5UemhMJ4_0),.din(w_dff_A_v6gqwMek3_0),.clk(gclk));
	jdff dff_A_P5UemhMJ4_0(.dout(w_dff_A_rAzB2KhL6_0),.din(w_dff_A_P5UemhMJ4_0),.clk(gclk));
	jdff dff_A_rAzB2KhL6_0(.dout(w_dff_A_BXZ6q2DB4_0),.din(w_dff_A_rAzB2KhL6_0),.clk(gclk));
	jdff dff_A_BXZ6q2DB4_0(.dout(w_dff_A_iMMJWG2L5_0),.din(w_dff_A_BXZ6q2DB4_0),.clk(gclk));
	jdff dff_A_iMMJWG2L5_0(.dout(w_dff_A_zhj8ihkX4_0),.din(w_dff_A_iMMJWG2L5_0),.clk(gclk));
	jdff dff_A_zhj8ihkX4_0(.dout(w_dff_A_kZ7tR5Vs6_0),.din(w_dff_A_zhj8ihkX4_0),.clk(gclk));
	jdff dff_A_kZ7tR5Vs6_0(.dout(w_dff_A_J25sRFb05_0),.din(w_dff_A_kZ7tR5Vs6_0),.clk(gclk));
	jdff dff_A_J25sRFb05_0(.dout(w_dff_A_qTXuH1Rl1_0),.din(w_dff_A_J25sRFb05_0),.clk(gclk));
	jdff dff_A_qTXuH1Rl1_0(.dout(w_dff_A_wJzBZD5p8_0),.din(w_dff_A_qTXuH1Rl1_0),.clk(gclk));
	jdff dff_A_wJzBZD5p8_0(.dout(w_dff_A_o6BtxZ6k7_0),.din(w_dff_A_wJzBZD5p8_0),.clk(gclk));
	jdff dff_A_o6BtxZ6k7_0(.dout(w_dff_A_DGm31C3J9_0),.din(w_dff_A_o6BtxZ6k7_0),.clk(gclk));
	jdff dff_A_DGm31C3J9_0(.dout(w_dff_A_XvQxqeEL5_0),.din(w_dff_A_DGm31C3J9_0),.clk(gclk));
	jdff dff_A_XvQxqeEL5_0(.dout(w_dff_A_tyEDMw7H2_0),.din(w_dff_A_XvQxqeEL5_0),.clk(gclk));
	jdff dff_A_tyEDMw7H2_0(.dout(w_dff_A_lS2OuWMh8_0),.din(w_dff_A_tyEDMw7H2_0),.clk(gclk));
	jdff dff_A_lS2OuWMh8_0(.dout(w_dff_A_AiLT5bqw0_0),.din(w_dff_A_lS2OuWMh8_0),.clk(gclk));
	jdff dff_A_AiLT5bqw0_0(.dout(w_dff_A_oZeBMBU93_0),.din(w_dff_A_AiLT5bqw0_0),.clk(gclk));
	jdff dff_A_oZeBMBU93_0(.dout(w_dff_A_RCoLPb1E4_0),.din(w_dff_A_oZeBMBU93_0),.clk(gclk));
	jdff dff_A_RCoLPb1E4_0(.dout(w_dff_A_8aHZwmOH9_0),.din(w_dff_A_RCoLPb1E4_0),.clk(gclk));
	jdff dff_A_8aHZwmOH9_0(.dout(w_dff_A_6p1zyRIY9_0),.din(w_dff_A_8aHZwmOH9_0),.clk(gclk));
	jdff dff_A_6p1zyRIY9_0(.dout(w_dff_A_gEO0PD3S4_0),.din(w_dff_A_6p1zyRIY9_0),.clk(gclk));
	jdff dff_A_gEO0PD3S4_0(.dout(w_dff_A_t0EGDvpx4_0),.din(w_dff_A_gEO0PD3S4_0),.clk(gclk));
	jdff dff_A_t0EGDvpx4_0(.dout(f51),.din(w_dff_A_t0EGDvpx4_0),.clk(gclk));
	jdff dff_A_G7GNSuM17_2(.dout(w_dff_A_l1Vh7YgW6_0),.din(w_dff_A_G7GNSuM17_2),.clk(gclk));
	jdff dff_A_l1Vh7YgW6_0(.dout(w_dff_A_YRgofBZ27_0),.din(w_dff_A_l1Vh7YgW6_0),.clk(gclk));
	jdff dff_A_YRgofBZ27_0(.dout(w_dff_A_t781VRLc6_0),.din(w_dff_A_YRgofBZ27_0),.clk(gclk));
	jdff dff_A_t781VRLc6_0(.dout(w_dff_A_OpGV8T1d9_0),.din(w_dff_A_t781VRLc6_0),.clk(gclk));
	jdff dff_A_OpGV8T1d9_0(.dout(w_dff_A_ZZI8jzxH0_0),.din(w_dff_A_OpGV8T1d9_0),.clk(gclk));
	jdff dff_A_ZZI8jzxH0_0(.dout(w_dff_A_BTmzGfix2_0),.din(w_dff_A_ZZI8jzxH0_0),.clk(gclk));
	jdff dff_A_BTmzGfix2_0(.dout(w_dff_A_iMOunIXD4_0),.din(w_dff_A_BTmzGfix2_0),.clk(gclk));
	jdff dff_A_iMOunIXD4_0(.dout(w_dff_A_uZkFKS1K2_0),.din(w_dff_A_iMOunIXD4_0),.clk(gclk));
	jdff dff_A_uZkFKS1K2_0(.dout(w_dff_A_7qGuwbAV7_0),.din(w_dff_A_uZkFKS1K2_0),.clk(gclk));
	jdff dff_A_7qGuwbAV7_0(.dout(w_dff_A_dVrQ63pj9_0),.din(w_dff_A_7qGuwbAV7_0),.clk(gclk));
	jdff dff_A_dVrQ63pj9_0(.dout(w_dff_A_EiR4OOmW4_0),.din(w_dff_A_dVrQ63pj9_0),.clk(gclk));
	jdff dff_A_EiR4OOmW4_0(.dout(w_dff_A_2wySulYn7_0),.din(w_dff_A_EiR4OOmW4_0),.clk(gclk));
	jdff dff_A_2wySulYn7_0(.dout(w_dff_A_FyJTiNBa6_0),.din(w_dff_A_2wySulYn7_0),.clk(gclk));
	jdff dff_A_FyJTiNBa6_0(.dout(w_dff_A_POP8tHOu1_0),.din(w_dff_A_FyJTiNBa6_0),.clk(gclk));
	jdff dff_A_POP8tHOu1_0(.dout(w_dff_A_09a3uzDm5_0),.din(w_dff_A_POP8tHOu1_0),.clk(gclk));
	jdff dff_A_09a3uzDm5_0(.dout(w_dff_A_86xese044_0),.din(w_dff_A_09a3uzDm5_0),.clk(gclk));
	jdff dff_A_86xese044_0(.dout(w_dff_A_wvbbBwei4_0),.din(w_dff_A_86xese044_0),.clk(gclk));
	jdff dff_A_wvbbBwei4_0(.dout(w_dff_A_QaWOJcub3_0),.din(w_dff_A_wvbbBwei4_0),.clk(gclk));
	jdff dff_A_QaWOJcub3_0(.dout(w_dff_A_G7bYDsnd0_0),.din(w_dff_A_QaWOJcub3_0),.clk(gclk));
	jdff dff_A_G7bYDsnd0_0(.dout(w_dff_A_ge6JoBjL4_0),.din(w_dff_A_G7bYDsnd0_0),.clk(gclk));
	jdff dff_A_ge6JoBjL4_0(.dout(w_dff_A_iXzRamAH7_0),.din(w_dff_A_ge6JoBjL4_0),.clk(gclk));
	jdff dff_A_iXzRamAH7_0(.dout(w_dff_A_YWdabcHF9_0),.din(w_dff_A_iXzRamAH7_0),.clk(gclk));
	jdff dff_A_YWdabcHF9_0(.dout(w_dff_A_kZ4PPs6C3_0),.din(w_dff_A_YWdabcHF9_0),.clk(gclk));
	jdff dff_A_kZ4PPs6C3_0(.dout(w_dff_A_hjCbWuiG0_0),.din(w_dff_A_kZ4PPs6C3_0),.clk(gclk));
	jdff dff_A_hjCbWuiG0_0(.dout(w_dff_A_zIAZchVZ0_0),.din(w_dff_A_hjCbWuiG0_0),.clk(gclk));
	jdff dff_A_zIAZchVZ0_0(.dout(w_dff_A_6k73NZF09_0),.din(w_dff_A_zIAZchVZ0_0),.clk(gclk));
	jdff dff_A_6k73NZF09_0(.dout(w_dff_A_u39syC7A8_0),.din(w_dff_A_6k73NZF09_0),.clk(gclk));
	jdff dff_A_u39syC7A8_0(.dout(w_dff_A_DLjQm3Yl1_0),.din(w_dff_A_u39syC7A8_0),.clk(gclk));
	jdff dff_A_DLjQm3Yl1_0(.dout(w_dff_A_cghGQbgO7_0),.din(w_dff_A_DLjQm3Yl1_0),.clk(gclk));
	jdff dff_A_cghGQbgO7_0(.dout(w_dff_A_BSLORxXU8_0),.din(w_dff_A_cghGQbgO7_0),.clk(gclk));
	jdff dff_A_BSLORxXU8_0(.dout(w_dff_A_t89g5p5Z7_0),.din(w_dff_A_BSLORxXU8_0),.clk(gclk));
	jdff dff_A_t89g5p5Z7_0(.dout(w_dff_A_jwDQdgv20_0),.din(w_dff_A_t89g5p5Z7_0),.clk(gclk));
	jdff dff_A_jwDQdgv20_0(.dout(w_dff_A_SSNR797D2_0),.din(w_dff_A_jwDQdgv20_0),.clk(gclk));
	jdff dff_A_SSNR797D2_0(.dout(w_dff_A_OdDu2nXl1_0),.din(w_dff_A_SSNR797D2_0),.clk(gclk));
	jdff dff_A_OdDu2nXl1_0(.dout(w_dff_A_xp0xzVgW6_0),.din(w_dff_A_OdDu2nXl1_0),.clk(gclk));
	jdff dff_A_xp0xzVgW6_0(.dout(w_dff_A_3UVpfIHH2_0),.din(w_dff_A_xp0xzVgW6_0),.clk(gclk));
	jdff dff_A_3UVpfIHH2_0(.dout(w_dff_A_eWAChmSl3_0),.din(w_dff_A_3UVpfIHH2_0),.clk(gclk));
	jdff dff_A_eWAChmSl3_0(.dout(w_dff_A_B2x0OPTf8_0),.din(w_dff_A_eWAChmSl3_0),.clk(gclk));
	jdff dff_A_B2x0OPTf8_0(.dout(w_dff_A_svCp7Kuf3_0),.din(w_dff_A_B2x0OPTf8_0),.clk(gclk));
	jdff dff_A_svCp7Kuf3_0(.dout(w_dff_A_3Y9U3X1j0_0),.din(w_dff_A_svCp7Kuf3_0),.clk(gclk));
	jdff dff_A_3Y9U3X1j0_0(.dout(w_dff_A_BlOuYw4O7_0),.din(w_dff_A_3Y9U3X1j0_0),.clk(gclk));
	jdff dff_A_BlOuYw4O7_0(.dout(w_dff_A_UiZeewtW8_0),.din(w_dff_A_BlOuYw4O7_0),.clk(gclk));
	jdff dff_A_UiZeewtW8_0(.dout(w_dff_A_G9vZRCnT1_0),.din(w_dff_A_UiZeewtW8_0),.clk(gclk));
	jdff dff_A_G9vZRCnT1_0(.dout(w_dff_A_pdE64WSt8_0),.din(w_dff_A_G9vZRCnT1_0),.clk(gclk));
	jdff dff_A_pdE64WSt8_0(.dout(w_dff_A_a8wci0QL2_0),.din(w_dff_A_pdE64WSt8_0),.clk(gclk));
	jdff dff_A_a8wci0QL2_0(.dout(w_dff_A_HVtc20pM6_0),.din(w_dff_A_a8wci0QL2_0),.clk(gclk));
	jdff dff_A_HVtc20pM6_0(.dout(w_dff_A_HoqDBzTy0_0),.din(w_dff_A_HVtc20pM6_0),.clk(gclk));
	jdff dff_A_HoqDBzTy0_0(.dout(w_dff_A_rvGeCKCp4_0),.din(w_dff_A_HoqDBzTy0_0),.clk(gclk));
	jdff dff_A_rvGeCKCp4_0(.dout(w_dff_A_5lX71WQ05_0),.din(w_dff_A_rvGeCKCp4_0),.clk(gclk));
	jdff dff_A_5lX71WQ05_0(.dout(w_dff_A_lRr46IbB3_0),.din(w_dff_A_5lX71WQ05_0),.clk(gclk));
	jdff dff_A_lRr46IbB3_0(.dout(w_dff_A_D2B9kVQh6_0),.din(w_dff_A_lRr46IbB3_0),.clk(gclk));
	jdff dff_A_D2B9kVQh6_0(.dout(w_dff_A_Ng1EtVUH7_0),.din(w_dff_A_D2B9kVQh6_0),.clk(gclk));
	jdff dff_A_Ng1EtVUH7_0(.dout(w_dff_A_6TU938Al0_0),.din(w_dff_A_Ng1EtVUH7_0),.clk(gclk));
	jdff dff_A_6TU938Al0_0(.dout(w_dff_A_cjivnYUC6_0),.din(w_dff_A_6TU938Al0_0),.clk(gclk));
	jdff dff_A_cjivnYUC6_0(.dout(w_dff_A_ph7VmcbG0_0),.din(w_dff_A_cjivnYUC6_0),.clk(gclk));
	jdff dff_A_ph7VmcbG0_0(.dout(w_dff_A_psBOdpLB2_0),.din(w_dff_A_ph7VmcbG0_0),.clk(gclk));
	jdff dff_A_psBOdpLB2_0(.dout(w_dff_A_5wUvn2Aa6_0),.din(w_dff_A_psBOdpLB2_0),.clk(gclk));
	jdff dff_A_5wUvn2Aa6_0(.dout(w_dff_A_o5aCjrWi9_0),.din(w_dff_A_5wUvn2Aa6_0),.clk(gclk));
	jdff dff_A_o5aCjrWi9_0(.dout(w_dff_A_yX64Na0j3_0),.din(w_dff_A_o5aCjrWi9_0),.clk(gclk));
	jdff dff_A_yX64Na0j3_0(.dout(w_dff_A_ybwSwN4q5_0),.din(w_dff_A_yX64Na0j3_0),.clk(gclk));
	jdff dff_A_ybwSwN4q5_0(.dout(w_dff_A_eqIXxdOv3_0),.din(w_dff_A_ybwSwN4q5_0),.clk(gclk));
	jdff dff_A_eqIXxdOv3_0(.dout(w_dff_A_EMdEozSn7_0),.din(w_dff_A_eqIXxdOv3_0),.clk(gclk));
	jdff dff_A_EMdEozSn7_0(.dout(w_dff_A_EqCpjty86_0),.din(w_dff_A_EMdEozSn7_0),.clk(gclk));
	jdff dff_A_EqCpjty86_0(.dout(w_dff_A_qJzw7aX38_0),.din(w_dff_A_EqCpjty86_0),.clk(gclk));
	jdff dff_A_qJzw7aX38_0(.dout(w_dff_A_Ih6dXHZ23_0),.din(w_dff_A_qJzw7aX38_0),.clk(gclk));
	jdff dff_A_Ih6dXHZ23_0(.dout(w_dff_A_dWAEoDRf8_0),.din(w_dff_A_Ih6dXHZ23_0),.clk(gclk));
	jdff dff_A_dWAEoDRf8_0(.dout(w_dff_A_ExzG3lhp8_0),.din(w_dff_A_dWAEoDRf8_0),.clk(gclk));
	jdff dff_A_ExzG3lhp8_0(.dout(w_dff_A_gmVidBMn2_0),.din(w_dff_A_ExzG3lhp8_0),.clk(gclk));
	jdff dff_A_gmVidBMn2_0(.dout(w_dff_A_ge5HwoRn0_0),.din(w_dff_A_gmVidBMn2_0),.clk(gclk));
	jdff dff_A_ge5HwoRn0_0(.dout(w_dff_A_2zNkM9dH8_0),.din(w_dff_A_ge5HwoRn0_0),.clk(gclk));
	jdff dff_A_2zNkM9dH8_0(.dout(w_dff_A_YJ1UD6012_0),.din(w_dff_A_2zNkM9dH8_0),.clk(gclk));
	jdff dff_A_YJ1UD6012_0(.dout(w_dff_A_xg3ILKV69_0),.din(w_dff_A_YJ1UD6012_0),.clk(gclk));
	jdff dff_A_xg3ILKV69_0(.dout(w_dff_A_hekdlsy96_0),.din(w_dff_A_xg3ILKV69_0),.clk(gclk));
	jdff dff_A_hekdlsy96_0(.dout(w_dff_A_ZkGIJPPY3_0),.din(w_dff_A_hekdlsy96_0),.clk(gclk));
	jdff dff_A_ZkGIJPPY3_0(.dout(f52),.din(w_dff_A_ZkGIJPPY3_0),.clk(gclk));
	jdff dff_A_J9A7hwTx6_2(.dout(w_dff_A_OT3GK1AG8_0),.din(w_dff_A_J9A7hwTx6_2),.clk(gclk));
	jdff dff_A_OT3GK1AG8_0(.dout(w_dff_A_z88WRpUP4_0),.din(w_dff_A_OT3GK1AG8_0),.clk(gclk));
	jdff dff_A_z88WRpUP4_0(.dout(w_dff_A_6aCdpau06_0),.din(w_dff_A_z88WRpUP4_0),.clk(gclk));
	jdff dff_A_6aCdpau06_0(.dout(w_dff_A_Z2SxVOMq0_0),.din(w_dff_A_6aCdpau06_0),.clk(gclk));
	jdff dff_A_Z2SxVOMq0_0(.dout(w_dff_A_t9pJlqlj0_0),.din(w_dff_A_Z2SxVOMq0_0),.clk(gclk));
	jdff dff_A_t9pJlqlj0_0(.dout(w_dff_A_mBrLKQAS5_0),.din(w_dff_A_t9pJlqlj0_0),.clk(gclk));
	jdff dff_A_mBrLKQAS5_0(.dout(w_dff_A_pPYqN8QY9_0),.din(w_dff_A_mBrLKQAS5_0),.clk(gclk));
	jdff dff_A_pPYqN8QY9_0(.dout(w_dff_A_nDxfWVzy4_0),.din(w_dff_A_pPYqN8QY9_0),.clk(gclk));
	jdff dff_A_nDxfWVzy4_0(.dout(w_dff_A_aKs1sSID5_0),.din(w_dff_A_nDxfWVzy4_0),.clk(gclk));
	jdff dff_A_aKs1sSID5_0(.dout(w_dff_A_SaDtsbVW5_0),.din(w_dff_A_aKs1sSID5_0),.clk(gclk));
	jdff dff_A_SaDtsbVW5_0(.dout(w_dff_A_rskkAhRw5_0),.din(w_dff_A_SaDtsbVW5_0),.clk(gclk));
	jdff dff_A_rskkAhRw5_0(.dout(w_dff_A_d16tCrGm7_0),.din(w_dff_A_rskkAhRw5_0),.clk(gclk));
	jdff dff_A_d16tCrGm7_0(.dout(w_dff_A_RrPLuR4w6_0),.din(w_dff_A_d16tCrGm7_0),.clk(gclk));
	jdff dff_A_RrPLuR4w6_0(.dout(w_dff_A_JPkdiDbF3_0),.din(w_dff_A_RrPLuR4w6_0),.clk(gclk));
	jdff dff_A_JPkdiDbF3_0(.dout(w_dff_A_CIZG3EZr5_0),.din(w_dff_A_JPkdiDbF3_0),.clk(gclk));
	jdff dff_A_CIZG3EZr5_0(.dout(w_dff_A_HrWvwZoa3_0),.din(w_dff_A_CIZG3EZr5_0),.clk(gclk));
	jdff dff_A_HrWvwZoa3_0(.dout(w_dff_A_T6keuIcK0_0),.din(w_dff_A_HrWvwZoa3_0),.clk(gclk));
	jdff dff_A_T6keuIcK0_0(.dout(w_dff_A_byhhlgXr4_0),.din(w_dff_A_T6keuIcK0_0),.clk(gclk));
	jdff dff_A_byhhlgXr4_0(.dout(w_dff_A_HQtRgNkz1_0),.din(w_dff_A_byhhlgXr4_0),.clk(gclk));
	jdff dff_A_HQtRgNkz1_0(.dout(w_dff_A_REKRK8Lc4_0),.din(w_dff_A_HQtRgNkz1_0),.clk(gclk));
	jdff dff_A_REKRK8Lc4_0(.dout(w_dff_A_mHslQZmo1_0),.din(w_dff_A_REKRK8Lc4_0),.clk(gclk));
	jdff dff_A_mHslQZmo1_0(.dout(w_dff_A_LPYnCjel0_0),.din(w_dff_A_mHslQZmo1_0),.clk(gclk));
	jdff dff_A_LPYnCjel0_0(.dout(w_dff_A_aiC8ujeM9_0),.din(w_dff_A_LPYnCjel0_0),.clk(gclk));
	jdff dff_A_aiC8ujeM9_0(.dout(w_dff_A_npbiUpmV7_0),.din(w_dff_A_aiC8ujeM9_0),.clk(gclk));
	jdff dff_A_npbiUpmV7_0(.dout(w_dff_A_WLuGQe8X5_0),.din(w_dff_A_npbiUpmV7_0),.clk(gclk));
	jdff dff_A_WLuGQe8X5_0(.dout(w_dff_A_ARD4GBYd6_0),.din(w_dff_A_WLuGQe8X5_0),.clk(gclk));
	jdff dff_A_ARD4GBYd6_0(.dout(w_dff_A_6vOwHz3W0_0),.din(w_dff_A_ARD4GBYd6_0),.clk(gclk));
	jdff dff_A_6vOwHz3W0_0(.dout(w_dff_A_1mVz9cx33_0),.din(w_dff_A_6vOwHz3W0_0),.clk(gclk));
	jdff dff_A_1mVz9cx33_0(.dout(w_dff_A_CezH1A4P9_0),.din(w_dff_A_1mVz9cx33_0),.clk(gclk));
	jdff dff_A_CezH1A4P9_0(.dout(w_dff_A_WkD4XFm68_0),.din(w_dff_A_CezH1A4P9_0),.clk(gclk));
	jdff dff_A_WkD4XFm68_0(.dout(w_dff_A_egb0vbE24_0),.din(w_dff_A_WkD4XFm68_0),.clk(gclk));
	jdff dff_A_egb0vbE24_0(.dout(w_dff_A_mUUSMgpW1_0),.din(w_dff_A_egb0vbE24_0),.clk(gclk));
	jdff dff_A_mUUSMgpW1_0(.dout(w_dff_A_tplcAAZk3_0),.din(w_dff_A_mUUSMgpW1_0),.clk(gclk));
	jdff dff_A_tplcAAZk3_0(.dout(w_dff_A_cugwLUWM2_0),.din(w_dff_A_tplcAAZk3_0),.clk(gclk));
	jdff dff_A_cugwLUWM2_0(.dout(w_dff_A_gCBjj5To0_0),.din(w_dff_A_cugwLUWM2_0),.clk(gclk));
	jdff dff_A_gCBjj5To0_0(.dout(w_dff_A_jS5ZeMDw7_0),.din(w_dff_A_gCBjj5To0_0),.clk(gclk));
	jdff dff_A_jS5ZeMDw7_0(.dout(w_dff_A_Kc14vn7P7_0),.din(w_dff_A_jS5ZeMDw7_0),.clk(gclk));
	jdff dff_A_Kc14vn7P7_0(.dout(w_dff_A_ieTvplCn3_0),.din(w_dff_A_Kc14vn7P7_0),.clk(gclk));
	jdff dff_A_ieTvplCn3_0(.dout(w_dff_A_prZETgUx6_0),.din(w_dff_A_ieTvplCn3_0),.clk(gclk));
	jdff dff_A_prZETgUx6_0(.dout(w_dff_A_CfTi23LL4_0),.din(w_dff_A_prZETgUx6_0),.clk(gclk));
	jdff dff_A_CfTi23LL4_0(.dout(w_dff_A_W5YcOg6s9_0),.din(w_dff_A_CfTi23LL4_0),.clk(gclk));
	jdff dff_A_W5YcOg6s9_0(.dout(w_dff_A_Y1xhP8IX0_0),.din(w_dff_A_W5YcOg6s9_0),.clk(gclk));
	jdff dff_A_Y1xhP8IX0_0(.dout(w_dff_A_i1ZkUOO01_0),.din(w_dff_A_Y1xhP8IX0_0),.clk(gclk));
	jdff dff_A_i1ZkUOO01_0(.dout(w_dff_A_ZpMOjCMn8_0),.din(w_dff_A_i1ZkUOO01_0),.clk(gclk));
	jdff dff_A_ZpMOjCMn8_0(.dout(w_dff_A_pdcznA3U1_0),.din(w_dff_A_ZpMOjCMn8_0),.clk(gclk));
	jdff dff_A_pdcznA3U1_0(.dout(w_dff_A_90PSYUac0_0),.din(w_dff_A_pdcznA3U1_0),.clk(gclk));
	jdff dff_A_90PSYUac0_0(.dout(w_dff_A_vYZoLNUU9_0),.din(w_dff_A_90PSYUac0_0),.clk(gclk));
	jdff dff_A_vYZoLNUU9_0(.dout(w_dff_A_clk9LFOM3_0),.din(w_dff_A_vYZoLNUU9_0),.clk(gclk));
	jdff dff_A_clk9LFOM3_0(.dout(w_dff_A_SiZXybuQ0_0),.din(w_dff_A_clk9LFOM3_0),.clk(gclk));
	jdff dff_A_SiZXybuQ0_0(.dout(w_dff_A_zX62wHPB0_0),.din(w_dff_A_SiZXybuQ0_0),.clk(gclk));
	jdff dff_A_zX62wHPB0_0(.dout(w_dff_A_LDuhTvzO4_0),.din(w_dff_A_zX62wHPB0_0),.clk(gclk));
	jdff dff_A_LDuhTvzO4_0(.dout(w_dff_A_utt3HlAP6_0),.din(w_dff_A_LDuhTvzO4_0),.clk(gclk));
	jdff dff_A_utt3HlAP6_0(.dout(w_dff_A_0kol8nHv1_0),.din(w_dff_A_utt3HlAP6_0),.clk(gclk));
	jdff dff_A_0kol8nHv1_0(.dout(w_dff_A_1dTZoTcV6_0),.din(w_dff_A_0kol8nHv1_0),.clk(gclk));
	jdff dff_A_1dTZoTcV6_0(.dout(w_dff_A_prsExu7H8_0),.din(w_dff_A_1dTZoTcV6_0),.clk(gclk));
	jdff dff_A_prsExu7H8_0(.dout(w_dff_A_qpW5m0wq7_0),.din(w_dff_A_prsExu7H8_0),.clk(gclk));
	jdff dff_A_qpW5m0wq7_0(.dout(w_dff_A_oLgD2FYp6_0),.din(w_dff_A_qpW5m0wq7_0),.clk(gclk));
	jdff dff_A_oLgD2FYp6_0(.dout(w_dff_A_tFvLmla28_0),.din(w_dff_A_oLgD2FYp6_0),.clk(gclk));
	jdff dff_A_tFvLmla28_0(.dout(w_dff_A_astKMbRC9_0),.din(w_dff_A_tFvLmla28_0),.clk(gclk));
	jdff dff_A_astKMbRC9_0(.dout(w_dff_A_DR0N3oYZ3_0),.din(w_dff_A_astKMbRC9_0),.clk(gclk));
	jdff dff_A_DR0N3oYZ3_0(.dout(w_dff_A_6ervdhKj7_0),.din(w_dff_A_DR0N3oYZ3_0),.clk(gclk));
	jdff dff_A_6ervdhKj7_0(.dout(w_dff_A_YDBDD9XM0_0),.din(w_dff_A_6ervdhKj7_0),.clk(gclk));
	jdff dff_A_YDBDD9XM0_0(.dout(w_dff_A_szJk4oae9_0),.din(w_dff_A_YDBDD9XM0_0),.clk(gclk));
	jdff dff_A_szJk4oae9_0(.dout(w_dff_A_dzOdhbct6_0),.din(w_dff_A_szJk4oae9_0),.clk(gclk));
	jdff dff_A_dzOdhbct6_0(.dout(w_dff_A_Z9iGPVmW6_0),.din(w_dff_A_dzOdhbct6_0),.clk(gclk));
	jdff dff_A_Z9iGPVmW6_0(.dout(w_dff_A_WReiHmMH0_0),.din(w_dff_A_Z9iGPVmW6_0),.clk(gclk));
	jdff dff_A_WReiHmMH0_0(.dout(w_dff_A_1PpJj5r82_0),.din(w_dff_A_WReiHmMH0_0),.clk(gclk));
	jdff dff_A_1PpJj5r82_0(.dout(w_dff_A_H7MVETaQ9_0),.din(w_dff_A_1PpJj5r82_0),.clk(gclk));
	jdff dff_A_H7MVETaQ9_0(.dout(w_dff_A_bfht0aHI1_0),.din(w_dff_A_H7MVETaQ9_0),.clk(gclk));
	jdff dff_A_bfht0aHI1_0(.dout(w_dff_A_yDaHJsnz9_0),.din(w_dff_A_bfht0aHI1_0),.clk(gclk));
	jdff dff_A_yDaHJsnz9_0(.dout(w_dff_A_pn6SeXyP7_0),.din(w_dff_A_yDaHJsnz9_0),.clk(gclk));
	jdff dff_A_pn6SeXyP7_0(.dout(w_dff_A_9SIcFGXG8_0),.din(w_dff_A_pn6SeXyP7_0),.clk(gclk));
	jdff dff_A_9SIcFGXG8_0(.dout(w_dff_A_PdGDE0w11_0),.din(w_dff_A_9SIcFGXG8_0),.clk(gclk));
	jdff dff_A_PdGDE0w11_0(.dout(f53),.din(w_dff_A_PdGDE0w11_0),.clk(gclk));
	jdff dff_A_VAnnSBRN8_2(.dout(w_dff_A_9dclbZFg8_0),.din(w_dff_A_VAnnSBRN8_2),.clk(gclk));
	jdff dff_A_9dclbZFg8_0(.dout(w_dff_A_H1Vz3KZD4_0),.din(w_dff_A_9dclbZFg8_0),.clk(gclk));
	jdff dff_A_H1Vz3KZD4_0(.dout(w_dff_A_714oKhDN7_0),.din(w_dff_A_H1Vz3KZD4_0),.clk(gclk));
	jdff dff_A_714oKhDN7_0(.dout(w_dff_A_Dbo2qgqC8_0),.din(w_dff_A_714oKhDN7_0),.clk(gclk));
	jdff dff_A_Dbo2qgqC8_0(.dout(w_dff_A_knKqIHwR8_0),.din(w_dff_A_Dbo2qgqC8_0),.clk(gclk));
	jdff dff_A_knKqIHwR8_0(.dout(w_dff_A_HLs8llKn5_0),.din(w_dff_A_knKqIHwR8_0),.clk(gclk));
	jdff dff_A_HLs8llKn5_0(.dout(w_dff_A_wjyhKIaP9_0),.din(w_dff_A_HLs8llKn5_0),.clk(gclk));
	jdff dff_A_wjyhKIaP9_0(.dout(w_dff_A_dlGzekG65_0),.din(w_dff_A_wjyhKIaP9_0),.clk(gclk));
	jdff dff_A_dlGzekG65_0(.dout(w_dff_A_44mmG9RV8_0),.din(w_dff_A_dlGzekG65_0),.clk(gclk));
	jdff dff_A_44mmG9RV8_0(.dout(w_dff_A_4KtgLMUH1_0),.din(w_dff_A_44mmG9RV8_0),.clk(gclk));
	jdff dff_A_4KtgLMUH1_0(.dout(w_dff_A_5Y1m7mUl0_0),.din(w_dff_A_4KtgLMUH1_0),.clk(gclk));
	jdff dff_A_5Y1m7mUl0_0(.dout(w_dff_A_TrnfOlBA5_0),.din(w_dff_A_5Y1m7mUl0_0),.clk(gclk));
	jdff dff_A_TrnfOlBA5_0(.dout(w_dff_A_9Q3mkgmn8_0),.din(w_dff_A_TrnfOlBA5_0),.clk(gclk));
	jdff dff_A_9Q3mkgmn8_0(.dout(w_dff_A_TWfIS3Y48_0),.din(w_dff_A_9Q3mkgmn8_0),.clk(gclk));
	jdff dff_A_TWfIS3Y48_0(.dout(w_dff_A_3OYjzytK3_0),.din(w_dff_A_TWfIS3Y48_0),.clk(gclk));
	jdff dff_A_3OYjzytK3_0(.dout(w_dff_A_b28BH3sI6_0),.din(w_dff_A_3OYjzytK3_0),.clk(gclk));
	jdff dff_A_b28BH3sI6_0(.dout(w_dff_A_dfu5OI8d7_0),.din(w_dff_A_b28BH3sI6_0),.clk(gclk));
	jdff dff_A_dfu5OI8d7_0(.dout(w_dff_A_FLLW9SZi4_0),.din(w_dff_A_dfu5OI8d7_0),.clk(gclk));
	jdff dff_A_FLLW9SZi4_0(.dout(w_dff_A_eurZLrOl5_0),.din(w_dff_A_FLLW9SZi4_0),.clk(gclk));
	jdff dff_A_eurZLrOl5_0(.dout(w_dff_A_J4lRUlM41_0),.din(w_dff_A_eurZLrOl5_0),.clk(gclk));
	jdff dff_A_J4lRUlM41_0(.dout(w_dff_A_FH8Jbixz1_0),.din(w_dff_A_J4lRUlM41_0),.clk(gclk));
	jdff dff_A_FH8Jbixz1_0(.dout(w_dff_A_AU04OJJb4_0),.din(w_dff_A_FH8Jbixz1_0),.clk(gclk));
	jdff dff_A_AU04OJJb4_0(.dout(w_dff_A_z1Ip7aOA5_0),.din(w_dff_A_AU04OJJb4_0),.clk(gclk));
	jdff dff_A_z1Ip7aOA5_0(.dout(w_dff_A_3rq6zMSZ4_0),.din(w_dff_A_z1Ip7aOA5_0),.clk(gclk));
	jdff dff_A_3rq6zMSZ4_0(.dout(w_dff_A_1FgSU8u30_0),.din(w_dff_A_3rq6zMSZ4_0),.clk(gclk));
	jdff dff_A_1FgSU8u30_0(.dout(w_dff_A_nU5DdzsQ8_0),.din(w_dff_A_1FgSU8u30_0),.clk(gclk));
	jdff dff_A_nU5DdzsQ8_0(.dout(w_dff_A_jHgPgV3P6_0),.din(w_dff_A_nU5DdzsQ8_0),.clk(gclk));
	jdff dff_A_jHgPgV3P6_0(.dout(w_dff_A_f78FGPY04_0),.din(w_dff_A_jHgPgV3P6_0),.clk(gclk));
	jdff dff_A_f78FGPY04_0(.dout(w_dff_A_xxjc11Jw2_0),.din(w_dff_A_f78FGPY04_0),.clk(gclk));
	jdff dff_A_xxjc11Jw2_0(.dout(w_dff_A_pHY3wEVz0_0),.din(w_dff_A_xxjc11Jw2_0),.clk(gclk));
	jdff dff_A_pHY3wEVz0_0(.dout(w_dff_A_woeJLyyP5_0),.din(w_dff_A_pHY3wEVz0_0),.clk(gclk));
	jdff dff_A_woeJLyyP5_0(.dout(w_dff_A_shKRasrK3_0),.din(w_dff_A_woeJLyyP5_0),.clk(gclk));
	jdff dff_A_shKRasrK3_0(.dout(w_dff_A_e4VjbQK76_0),.din(w_dff_A_shKRasrK3_0),.clk(gclk));
	jdff dff_A_e4VjbQK76_0(.dout(w_dff_A_laEcLmxb5_0),.din(w_dff_A_e4VjbQK76_0),.clk(gclk));
	jdff dff_A_laEcLmxb5_0(.dout(w_dff_A_VnS7i1n47_0),.din(w_dff_A_laEcLmxb5_0),.clk(gclk));
	jdff dff_A_VnS7i1n47_0(.dout(w_dff_A_gYlyyBcP4_0),.din(w_dff_A_VnS7i1n47_0),.clk(gclk));
	jdff dff_A_gYlyyBcP4_0(.dout(w_dff_A_gnzT7elK8_0),.din(w_dff_A_gYlyyBcP4_0),.clk(gclk));
	jdff dff_A_gnzT7elK8_0(.dout(w_dff_A_KT063OkY9_0),.din(w_dff_A_gnzT7elK8_0),.clk(gclk));
	jdff dff_A_KT063OkY9_0(.dout(w_dff_A_REvm0Ti38_0),.din(w_dff_A_KT063OkY9_0),.clk(gclk));
	jdff dff_A_REvm0Ti38_0(.dout(w_dff_A_hEIdsQBR7_0),.din(w_dff_A_REvm0Ti38_0),.clk(gclk));
	jdff dff_A_hEIdsQBR7_0(.dout(w_dff_A_lrxGnw5p6_0),.din(w_dff_A_hEIdsQBR7_0),.clk(gclk));
	jdff dff_A_lrxGnw5p6_0(.dout(w_dff_A_NksPVsVY1_0),.din(w_dff_A_lrxGnw5p6_0),.clk(gclk));
	jdff dff_A_NksPVsVY1_0(.dout(w_dff_A_B0e1tjFT2_0),.din(w_dff_A_NksPVsVY1_0),.clk(gclk));
	jdff dff_A_B0e1tjFT2_0(.dout(w_dff_A_wGAb6cgj5_0),.din(w_dff_A_B0e1tjFT2_0),.clk(gclk));
	jdff dff_A_wGAb6cgj5_0(.dout(w_dff_A_kOvwD4EN1_0),.din(w_dff_A_wGAb6cgj5_0),.clk(gclk));
	jdff dff_A_kOvwD4EN1_0(.dout(w_dff_A_xXh45aOw1_0),.din(w_dff_A_kOvwD4EN1_0),.clk(gclk));
	jdff dff_A_xXh45aOw1_0(.dout(w_dff_A_F7myeWuA9_0),.din(w_dff_A_xXh45aOw1_0),.clk(gclk));
	jdff dff_A_F7myeWuA9_0(.dout(w_dff_A_NzAkOC3J2_0),.din(w_dff_A_F7myeWuA9_0),.clk(gclk));
	jdff dff_A_NzAkOC3J2_0(.dout(w_dff_A_lHMY5O9U2_0),.din(w_dff_A_NzAkOC3J2_0),.clk(gclk));
	jdff dff_A_lHMY5O9U2_0(.dout(w_dff_A_WaprlTOm8_0),.din(w_dff_A_lHMY5O9U2_0),.clk(gclk));
	jdff dff_A_WaprlTOm8_0(.dout(w_dff_A_Z9V70P7D1_0),.din(w_dff_A_WaprlTOm8_0),.clk(gclk));
	jdff dff_A_Z9V70P7D1_0(.dout(w_dff_A_FoIMywaP6_0),.din(w_dff_A_Z9V70P7D1_0),.clk(gclk));
	jdff dff_A_FoIMywaP6_0(.dout(w_dff_A_aUiQH5065_0),.din(w_dff_A_FoIMywaP6_0),.clk(gclk));
	jdff dff_A_aUiQH5065_0(.dout(w_dff_A_UaEBNyVD6_0),.din(w_dff_A_aUiQH5065_0),.clk(gclk));
	jdff dff_A_UaEBNyVD6_0(.dout(w_dff_A_v8xBNfep9_0),.din(w_dff_A_UaEBNyVD6_0),.clk(gclk));
	jdff dff_A_v8xBNfep9_0(.dout(w_dff_A_6TCBvEZt0_0),.din(w_dff_A_v8xBNfep9_0),.clk(gclk));
	jdff dff_A_6TCBvEZt0_0(.dout(w_dff_A_UGYMim0V1_0),.din(w_dff_A_6TCBvEZt0_0),.clk(gclk));
	jdff dff_A_UGYMim0V1_0(.dout(w_dff_A_2PjSqNPD0_0),.din(w_dff_A_UGYMim0V1_0),.clk(gclk));
	jdff dff_A_2PjSqNPD0_0(.dout(w_dff_A_ELfXi9OM0_0),.din(w_dff_A_2PjSqNPD0_0),.clk(gclk));
	jdff dff_A_ELfXi9OM0_0(.dout(w_dff_A_ScjEGo8T7_0),.din(w_dff_A_ELfXi9OM0_0),.clk(gclk));
	jdff dff_A_ScjEGo8T7_0(.dout(w_dff_A_yLQPyHP65_0),.din(w_dff_A_ScjEGo8T7_0),.clk(gclk));
	jdff dff_A_yLQPyHP65_0(.dout(w_dff_A_h5Z40Nx32_0),.din(w_dff_A_yLQPyHP65_0),.clk(gclk));
	jdff dff_A_h5Z40Nx32_0(.dout(w_dff_A_e6FpgkT84_0),.din(w_dff_A_h5Z40Nx32_0),.clk(gclk));
	jdff dff_A_e6FpgkT84_0(.dout(w_dff_A_271WHuu79_0),.din(w_dff_A_e6FpgkT84_0),.clk(gclk));
	jdff dff_A_271WHuu79_0(.dout(w_dff_A_hZJlLi9b2_0),.din(w_dff_A_271WHuu79_0),.clk(gclk));
	jdff dff_A_hZJlLi9b2_0(.dout(w_dff_A_gr1AarT87_0),.din(w_dff_A_hZJlLi9b2_0),.clk(gclk));
	jdff dff_A_gr1AarT87_0(.dout(w_dff_A_ZsrDp5Hb4_0),.din(w_dff_A_gr1AarT87_0),.clk(gclk));
	jdff dff_A_ZsrDp5Hb4_0(.dout(w_dff_A_r7TiYwRb5_0),.din(w_dff_A_ZsrDp5Hb4_0),.clk(gclk));
	jdff dff_A_r7TiYwRb5_0(.dout(w_dff_A_wQc4N6F10_0),.din(w_dff_A_r7TiYwRb5_0),.clk(gclk));
	jdff dff_A_wQc4N6F10_0(.dout(w_dff_A_w0TpfyKX6_0),.din(w_dff_A_wQc4N6F10_0),.clk(gclk));
	jdff dff_A_w0TpfyKX6_0(.dout(w_dff_A_i00tNIAk7_0),.din(w_dff_A_w0TpfyKX6_0),.clk(gclk));
	jdff dff_A_i00tNIAk7_0(.dout(w_dff_A_ayUQ4M2B4_0),.din(w_dff_A_i00tNIAk7_0),.clk(gclk));
	jdff dff_A_ayUQ4M2B4_0(.dout(f54),.din(w_dff_A_ayUQ4M2B4_0),.clk(gclk));
	jdff dff_A_w2HyVyOp2_2(.dout(w_dff_A_dEgH3gZa5_0),.din(w_dff_A_w2HyVyOp2_2),.clk(gclk));
	jdff dff_A_dEgH3gZa5_0(.dout(w_dff_A_e3EN56Ug9_0),.din(w_dff_A_dEgH3gZa5_0),.clk(gclk));
	jdff dff_A_e3EN56Ug9_0(.dout(w_dff_A_MGsqM0QD9_0),.din(w_dff_A_e3EN56Ug9_0),.clk(gclk));
	jdff dff_A_MGsqM0QD9_0(.dout(w_dff_A_424vlOw97_0),.din(w_dff_A_MGsqM0QD9_0),.clk(gclk));
	jdff dff_A_424vlOw97_0(.dout(w_dff_A_vqFXGeDc9_0),.din(w_dff_A_424vlOw97_0),.clk(gclk));
	jdff dff_A_vqFXGeDc9_0(.dout(w_dff_A_fxeMHGBj1_0),.din(w_dff_A_vqFXGeDc9_0),.clk(gclk));
	jdff dff_A_fxeMHGBj1_0(.dout(w_dff_A_5eCmOOrO8_0),.din(w_dff_A_fxeMHGBj1_0),.clk(gclk));
	jdff dff_A_5eCmOOrO8_0(.dout(w_dff_A_fCnjqpdM9_0),.din(w_dff_A_5eCmOOrO8_0),.clk(gclk));
	jdff dff_A_fCnjqpdM9_0(.dout(w_dff_A_SP5xCAOO3_0),.din(w_dff_A_fCnjqpdM9_0),.clk(gclk));
	jdff dff_A_SP5xCAOO3_0(.dout(w_dff_A_nOCCSmuC9_0),.din(w_dff_A_SP5xCAOO3_0),.clk(gclk));
	jdff dff_A_nOCCSmuC9_0(.dout(w_dff_A_4y19yrRB2_0),.din(w_dff_A_nOCCSmuC9_0),.clk(gclk));
	jdff dff_A_4y19yrRB2_0(.dout(w_dff_A_cn1xMRgu8_0),.din(w_dff_A_4y19yrRB2_0),.clk(gclk));
	jdff dff_A_cn1xMRgu8_0(.dout(w_dff_A_lHLZynKs6_0),.din(w_dff_A_cn1xMRgu8_0),.clk(gclk));
	jdff dff_A_lHLZynKs6_0(.dout(w_dff_A_FBWUylAB6_0),.din(w_dff_A_lHLZynKs6_0),.clk(gclk));
	jdff dff_A_FBWUylAB6_0(.dout(w_dff_A_hlnueaBz6_0),.din(w_dff_A_FBWUylAB6_0),.clk(gclk));
	jdff dff_A_hlnueaBz6_0(.dout(w_dff_A_fC7LxQrg5_0),.din(w_dff_A_hlnueaBz6_0),.clk(gclk));
	jdff dff_A_fC7LxQrg5_0(.dout(w_dff_A_pbo0JmI97_0),.din(w_dff_A_fC7LxQrg5_0),.clk(gclk));
	jdff dff_A_pbo0JmI97_0(.dout(w_dff_A_WtUhihMP7_0),.din(w_dff_A_pbo0JmI97_0),.clk(gclk));
	jdff dff_A_WtUhihMP7_0(.dout(w_dff_A_5IlrSkiZ1_0),.din(w_dff_A_WtUhihMP7_0),.clk(gclk));
	jdff dff_A_5IlrSkiZ1_0(.dout(w_dff_A_eOyP6tTM9_0),.din(w_dff_A_5IlrSkiZ1_0),.clk(gclk));
	jdff dff_A_eOyP6tTM9_0(.dout(w_dff_A_wIKtdQ1K0_0),.din(w_dff_A_eOyP6tTM9_0),.clk(gclk));
	jdff dff_A_wIKtdQ1K0_0(.dout(w_dff_A_cnW6YU3B0_0),.din(w_dff_A_wIKtdQ1K0_0),.clk(gclk));
	jdff dff_A_cnW6YU3B0_0(.dout(w_dff_A_DNneq2c38_0),.din(w_dff_A_cnW6YU3B0_0),.clk(gclk));
	jdff dff_A_DNneq2c38_0(.dout(w_dff_A_vTKNXfgK2_0),.din(w_dff_A_DNneq2c38_0),.clk(gclk));
	jdff dff_A_vTKNXfgK2_0(.dout(w_dff_A_ETAzq8d28_0),.din(w_dff_A_vTKNXfgK2_0),.clk(gclk));
	jdff dff_A_ETAzq8d28_0(.dout(w_dff_A_wRj2UmGg4_0),.din(w_dff_A_ETAzq8d28_0),.clk(gclk));
	jdff dff_A_wRj2UmGg4_0(.dout(w_dff_A_TezxDVX47_0),.din(w_dff_A_wRj2UmGg4_0),.clk(gclk));
	jdff dff_A_TezxDVX47_0(.dout(w_dff_A_CiubDuNg1_0),.din(w_dff_A_TezxDVX47_0),.clk(gclk));
	jdff dff_A_CiubDuNg1_0(.dout(w_dff_A_6839GalW5_0),.din(w_dff_A_CiubDuNg1_0),.clk(gclk));
	jdff dff_A_6839GalW5_0(.dout(w_dff_A_JZiKi63P2_0),.din(w_dff_A_6839GalW5_0),.clk(gclk));
	jdff dff_A_JZiKi63P2_0(.dout(w_dff_A_UmeOw9qz5_0),.din(w_dff_A_JZiKi63P2_0),.clk(gclk));
	jdff dff_A_UmeOw9qz5_0(.dout(w_dff_A_om6LMqsY6_0),.din(w_dff_A_UmeOw9qz5_0),.clk(gclk));
	jdff dff_A_om6LMqsY6_0(.dout(w_dff_A_pnKXDrFZ2_0),.din(w_dff_A_om6LMqsY6_0),.clk(gclk));
	jdff dff_A_pnKXDrFZ2_0(.dout(w_dff_A_EkvWhy9c1_0),.din(w_dff_A_pnKXDrFZ2_0),.clk(gclk));
	jdff dff_A_EkvWhy9c1_0(.dout(w_dff_A_McuKVLE19_0),.din(w_dff_A_EkvWhy9c1_0),.clk(gclk));
	jdff dff_A_McuKVLE19_0(.dout(w_dff_A_O2c9yV886_0),.din(w_dff_A_McuKVLE19_0),.clk(gclk));
	jdff dff_A_O2c9yV886_0(.dout(w_dff_A_vmS1Tf6j7_0),.din(w_dff_A_O2c9yV886_0),.clk(gclk));
	jdff dff_A_vmS1Tf6j7_0(.dout(w_dff_A_BcQnvUUK0_0),.din(w_dff_A_vmS1Tf6j7_0),.clk(gclk));
	jdff dff_A_BcQnvUUK0_0(.dout(w_dff_A_XxhYinKL9_0),.din(w_dff_A_BcQnvUUK0_0),.clk(gclk));
	jdff dff_A_XxhYinKL9_0(.dout(w_dff_A_jmScHiG65_0),.din(w_dff_A_XxhYinKL9_0),.clk(gclk));
	jdff dff_A_jmScHiG65_0(.dout(w_dff_A_6HrDtJvH1_0),.din(w_dff_A_jmScHiG65_0),.clk(gclk));
	jdff dff_A_6HrDtJvH1_0(.dout(w_dff_A_EeofwH1E4_0),.din(w_dff_A_6HrDtJvH1_0),.clk(gclk));
	jdff dff_A_EeofwH1E4_0(.dout(w_dff_A_qMNdxDAx8_0),.din(w_dff_A_EeofwH1E4_0),.clk(gclk));
	jdff dff_A_qMNdxDAx8_0(.dout(w_dff_A_sRnl4iWS2_0),.din(w_dff_A_qMNdxDAx8_0),.clk(gclk));
	jdff dff_A_sRnl4iWS2_0(.dout(w_dff_A_Gov2DavA1_0),.din(w_dff_A_sRnl4iWS2_0),.clk(gclk));
	jdff dff_A_Gov2DavA1_0(.dout(w_dff_A_1x2YLxUC5_0),.din(w_dff_A_Gov2DavA1_0),.clk(gclk));
	jdff dff_A_1x2YLxUC5_0(.dout(w_dff_A_qHqQcl8L5_0),.din(w_dff_A_1x2YLxUC5_0),.clk(gclk));
	jdff dff_A_qHqQcl8L5_0(.dout(w_dff_A_AaPLH0O98_0),.din(w_dff_A_qHqQcl8L5_0),.clk(gclk));
	jdff dff_A_AaPLH0O98_0(.dout(w_dff_A_zDreKGMw3_0),.din(w_dff_A_AaPLH0O98_0),.clk(gclk));
	jdff dff_A_zDreKGMw3_0(.dout(w_dff_A_1B5uHCIJ5_0),.din(w_dff_A_zDreKGMw3_0),.clk(gclk));
	jdff dff_A_1B5uHCIJ5_0(.dout(w_dff_A_obB3jffj7_0),.din(w_dff_A_1B5uHCIJ5_0),.clk(gclk));
	jdff dff_A_obB3jffj7_0(.dout(w_dff_A_2inXgvHr5_0),.din(w_dff_A_obB3jffj7_0),.clk(gclk));
	jdff dff_A_2inXgvHr5_0(.dout(w_dff_A_zMQsW4rp5_0),.din(w_dff_A_2inXgvHr5_0),.clk(gclk));
	jdff dff_A_zMQsW4rp5_0(.dout(w_dff_A_kDzuObk15_0),.din(w_dff_A_zMQsW4rp5_0),.clk(gclk));
	jdff dff_A_kDzuObk15_0(.dout(w_dff_A_gM8rTyx33_0),.din(w_dff_A_kDzuObk15_0),.clk(gclk));
	jdff dff_A_gM8rTyx33_0(.dout(w_dff_A_3KhK7FKk4_0),.din(w_dff_A_gM8rTyx33_0),.clk(gclk));
	jdff dff_A_3KhK7FKk4_0(.dout(w_dff_A_YHo9eLPz9_0),.din(w_dff_A_3KhK7FKk4_0),.clk(gclk));
	jdff dff_A_YHo9eLPz9_0(.dout(w_dff_A_B3mL47Ol0_0),.din(w_dff_A_YHo9eLPz9_0),.clk(gclk));
	jdff dff_A_B3mL47Ol0_0(.dout(w_dff_A_UIose7X75_0),.din(w_dff_A_B3mL47Ol0_0),.clk(gclk));
	jdff dff_A_UIose7X75_0(.dout(w_dff_A_6knHOhdi5_0),.din(w_dff_A_UIose7X75_0),.clk(gclk));
	jdff dff_A_6knHOhdi5_0(.dout(w_dff_A_ujgxaduW8_0),.din(w_dff_A_6knHOhdi5_0),.clk(gclk));
	jdff dff_A_ujgxaduW8_0(.dout(w_dff_A_zdrczSWU2_0),.din(w_dff_A_ujgxaduW8_0),.clk(gclk));
	jdff dff_A_zdrczSWU2_0(.dout(w_dff_A_nEf6vn7y6_0),.din(w_dff_A_zdrczSWU2_0),.clk(gclk));
	jdff dff_A_nEf6vn7y6_0(.dout(w_dff_A_XuxYCQog7_0),.din(w_dff_A_nEf6vn7y6_0),.clk(gclk));
	jdff dff_A_XuxYCQog7_0(.dout(w_dff_A_lT651o3w4_0),.din(w_dff_A_XuxYCQog7_0),.clk(gclk));
	jdff dff_A_lT651o3w4_0(.dout(w_dff_A_mTAZ184J2_0),.din(w_dff_A_lT651o3w4_0),.clk(gclk));
	jdff dff_A_mTAZ184J2_0(.dout(w_dff_A_NzAA6erK0_0),.din(w_dff_A_mTAZ184J2_0),.clk(gclk));
	jdff dff_A_NzAA6erK0_0(.dout(w_dff_A_CI7tv4nR2_0),.din(w_dff_A_NzAA6erK0_0),.clk(gclk));
	jdff dff_A_CI7tv4nR2_0(.dout(w_dff_A_Q2dUOvdm8_0),.din(w_dff_A_CI7tv4nR2_0),.clk(gclk));
	jdff dff_A_Q2dUOvdm8_0(.dout(w_dff_A_QUCKT1qY1_0),.din(w_dff_A_Q2dUOvdm8_0),.clk(gclk));
	jdff dff_A_QUCKT1qY1_0(.dout(w_dff_A_XfBcr8Xc9_0),.din(w_dff_A_QUCKT1qY1_0),.clk(gclk));
	jdff dff_A_XfBcr8Xc9_0(.dout(f55),.din(w_dff_A_XfBcr8Xc9_0),.clk(gclk));
	jdff dff_A_0ifBWpOE0_2(.dout(w_dff_A_Rmu6IeBp3_0),.din(w_dff_A_0ifBWpOE0_2),.clk(gclk));
	jdff dff_A_Rmu6IeBp3_0(.dout(w_dff_A_c13PA3Mc0_0),.din(w_dff_A_Rmu6IeBp3_0),.clk(gclk));
	jdff dff_A_c13PA3Mc0_0(.dout(w_dff_A_ayPpK3iw9_0),.din(w_dff_A_c13PA3Mc0_0),.clk(gclk));
	jdff dff_A_ayPpK3iw9_0(.dout(w_dff_A_zVD5pPD83_0),.din(w_dff_A_ayPpK3iw9_0),.clk(gclk));
	jdff dff_A_zVD5pPD83_0(.dout(w_dff_A_qhCPedcf8_0),.din(w_dff_A_zVD5pPD83_0),.clk(gclk));
	jdff dff_A_qhCPedcf8_0(.dout(w_dff_A_5mdW9eA25_0),.din(w_dff_A_qhCPedcf8_0),.clk(gclk));
	jdff dff_A_5mdW9eA25_0(.dout(w_dff_A_dL6WfK9L7_0),.din(w_dff_A_5mdW9eA25_0),.clk(gclk));
	jdff dff_A_dL6WfK9L7_0(.dout(w_dff_A_SpbtbmWe6_0),.din(w_dff_A_dL6WfK9L7_0),.clk(gclk));
	jdff dff_A_SpbtbmWe6_0(.dout(w_dff_A_hbuPn93z3_0),.din(w_dff_A_SpbtbmWe6_0),.clk(gclk));
	jdff dff_A_hbuPn93z3_0(.dout(w_dff_A_PMldSt8j0_0),.din(w_dff_A_hbuPn93z3_0),.clk(gclk));
	jdff dff_A_PMldSt8j0_0(.dout(w_dff_A_0xgDCn5z7_0),.din(w_dff_A_PMldSt8j0_0),.clk(gclk));
	jdff dff_A_0xgDCn5z7_0(.dout(w_dff_A_c9ANKgon7_0),.din(w_dff_A_0xgDCn5z7_0),.clk(gclk));
	jdff dff_A_c9ANKgon7_0(.dout(w_dff_A_DzYvff6t7_0),.din(w_dff_A_c9ANKgon7_0),.clk(gclk));
	jdff dff_A_DzYvff6t7_0(.dout(w_dff_A_dLsKJYNz0_0),.din(w_dff_A_DzYvff6t7_0),.clk(gclk));
	jdff dff_A_dLsKJYNz0_0(.dout(w_dff_A_546VhKMd2_0),.din(w_dff_A_dLsKJYNz0_0),.clk(gclk));
	jdff dff_A_546VhKMd2_0(.dout(w_dff_A_2fvITQwY3_0),.din(w_dff_A_546VhKMd2_0),.clk(gclk));
	jdff dff_A_2fvITQwY3_0(.dout(w_dff_A_VM0zCInD4_0),.din(w_dff_A_2fvITQwY3_0),.clk(gclk));
	jdff dff_A_VM0zCInD4_0(.dout(w_dff_A_qRs64vNu7_0),.din(w_dff_A_VM0zCInD4_0),.clk(gclk));
	jdff dff_A_qRs64vNu7_0(.dout(w_dff_A_tLRrioN56_0),.din(w_dff_A_qRs64vNu7_0),.clk(gclk));
	jdff dff_A_tLRrioN56_0(.dout(w_dff_A_oLi9KfmR3_0),.din(w_dff_A_tLRrioN56_0),.clk(gclk));
	jdff dff_A_oLi9KfmR3_0(.dout(w_dff_A_qOumC5p46_0),.din(w_dff_A_oLi9KfmR3_0),.clk(gclk));
	jdff dff_A_qOumC5p46_0(.dout(w_dff_A_zc5VxotV5_0),.din(w_dff_A_qOumC5p46_0),.clk(gclk));
	jdff dff_A_zc5VxotV5_0(.dout(w_dff_A_t6hlBMUT9_0),.din(w_dff_A_zc5VxotV5_0),.clk(gclk));
	jdff dff_A_t6hlBMUT9_0(.dout(w_dff_A_4lpClHmY8_0),.din(w_dff_A_t6hlBMUT9_0),.clk(gclk));
	jdff dff_A_4lpClHmY8_0(.dout(w_dff_A_GDcdsuGN7_0),.din(w_dff_A_4lpClHmY8_0),.clk(gclk));
	jdff dff_A_GDcdsuGN7_0(.dout(w_dff_A_CnGQY7IH6_0),.din(w_dff_A_GDcdsuGN7_0),.clk(gclk));
	jdff dff_A_CnGQY7IH6_0(.dout(w_dff_A_IEP2ywln1_0),.din(w_dff_A_CnGQY7IH6_0),.clk(gclk));
	jdff dff_A_IEP2ywln1_0(.dout(w_dff_A_HVl97lFC3_0),.din(w_dff_A_IEP2ywln1_0),.clk(gclk));
	jdff dff_A_HVl97lFC3_0(.dout(w_dff_A_9pPqOvsr4_0),.din(w_dff_A_HVl97lFC3_0),.clk(gclk));
	jdff dff_A_9pPqOvsr4_0(.dout(w_dff_A_Ds1Iroqm5_0),.din(w_dff_A_9pPqOvsr4_0),.clk(gclk));
	jdff dff_A_Ds1Iroqm5_0(.dout(w_dff_A_a4mejR9R5_0),.din(w_dff_A_Ds1Iroqm5_0),.clk(gclk));
	jdff dff_A_a4mejR9R5_0(.dout(w_dff_A_Lw9Wm6ZG2_0),.din(w_dff_A_a4mejR9R5_0),.clk(gclk));
	jdff dff_A_Lw9Wm6ZG2_0(.dout(w_dff_A_Qji9yAsW6_0),.din(w_dff_A_Lw9Wm6ZG2_0),.clk(gclk));
	jdff dff_A_Qji9yAsW6_0(.dout(w_dff_A_kE8lqlHy4_0),.din(w_dff_A_Qji9yAsW6_0),.clk(gclk));
	jdff dff_A_kE8lqlHy4_0(.dout(w_dff_A_xTIwdaok7_0),.din(w_dff_A_kE8lqlHy4_0),.clk(gclk));
	jdff dff_A_xTIwdaok7_0(.dout(w_dff_A_xLxeiD2W4_0),.din(w_dff_A_xTIwdaok7_0),.clk(gclk));
	jdff dff_A_xLxeiD2W4_0(.dout(w_dff_A_NpK5X4pA4_0),.din(w_dff_A_xLxeiD2W4_0),.clk(gclk));
	jdff dff_A_NpK5X4pA4_0(.dout(w_dff_A_wrZW0Lw43_0),.din(w_dff_A_NpK5X4pA4_0),.clk(gclk));
	jdff dff_A_wrZW0Lw43_0(.dout(w_dff_A_iOxkUXdF8_0),.din(w_dff_A_wrZW0Lw43_0),.clk(gclk));
	jdff dff_A_iOxkUXdF8_0(.dout(w_dff_A_NSdiEKXq9_0),.din(w_dff_A_iOxkUXdF8_0),.clk(gclk));
	jdff dff_A_NSdiEKXq9_0(.dout(w_dff_A_F632qRFm3_0),.din(w_dff_A_NSdiEKXq9_0),.clk(gclk));
	jdff dff_A_F632qRFm3_0(.dout(w_dff_A_5oZFBbjY8_0),.din(w_dff_A_F632qRFm3_0),.clk(gclk));
	jdff dff_A_5oZFBbjY8_0(.dout(w_dff_A_a2vEkte32_0),.din(w_dff_A_5oZFBbjY8_0),.clk(gclk));
	jdff dff_A_a2vEkte32_0(.dout(w_dff_A_N7jT3wYM6_0),.din(w_dff_A_a2vEkte32_0),.clk(gclk));
	jdff dff_A_N7jT3wYM6_0(.dout(w_dff_A_aleX8rro6_0),.din(w_dff_A_N7jT3wYM6_0),.clk(gclk));
	jdff dff_A_aleX8rro6_0(.dout(w_dff_A_MsPL2tlL5_0),.din(w_dff_A_aleX8rro6_0),.clk(gclk));
	jdff dff_A_MsPL2tlL5_0(.dout(w_dff_A_YJjFLiKR5_0),.din(w_dff_A_MsPL2tlL5_0),.clk(gclk));
	jdff dff_A_YJjFLiKR5_0(.dout(w_dff_A_wKeEnhlP8_0),.din(w_dff_A_YJjFLiKR5_0),.clk(gclk));
	jdff dff_A_wKeEnhlP8_0(.dout(w_dff_A_5hmPO68u9_0),.din(w_dff_A_wKeEnhlP8_0),.clk(gclk));
	jdff dff_A_5hmPO68u9_0(.dout(w_dff_A_URqIKR3N9_0),.din(w_dff_A_5hmPO68u9_0),.clk(gclk));
	jdff dff_A_URqIKR3N9_0(.dout(w_dff_A_b9MSUZHG0_0),.din(w_dff_A_URqIKR3N9_0),.clk(gclk));
	jdff dff_A_b9MSUZHG0_0(.dout(w_dff_A_llSMmZCC9_0),.din(w_dff_A_b9MSUZHG0_0),.clk(gclk));
	jdff dff_A_llSMmZCC9_0(.dout(w_dff_A_ViMwEsyT2_0),.din(w_dff_A_llSMmZCC9_0),.clk(gclk));
	jdff dff_A_ViMwEsyT2_0(.dout(w_dff_A_6DwsPHkN2_0),.din(w_dff_A_ViMwEsyT2_0),.clk(gclk));
	jdff dff_A_6DwsPHkN2_0(.dout(w_dff_A_qjpDKxOh4_0),.din(w_dff_A_6DwsPHkN2_0),.clk(gclk));
	jdff dff_A_qjpDKxOh4_0(.dout(w_dff_A_h17dLYDX7_0),.din(w_dff_A_qjpDKxOh4_0),.clk(gclk));
	jdff dff_A_h17dLYDX7_0(.dout(w_dff_A_qOY04Bby5_0),.din(w_dff_A_h17dLYDX7_0),.clk(gclk));
	jdff dff_A_qOY04Bby5_0(.dout(w_dff_A_KPm0xNmJ3_0),.din(w_dff_A_qOY04Bby5_0),.clk(gclk));
	jdff dff_A_KPm0xNmJ3_0(.dout(w_dff_A_ImRMMbb36_0),.din(w_dff_A_KPm0xNmJ3_0),.clk(gclk));
	jdff dff_A_ImRMMbb36_0(.dout(w_dff_A_l1gWUlAh7_0),.din(w_dff_A_ImRMMbb36_0),.clk(gclk));
	jdff dff_A_l1gWUlAh7_0(.dout(w_dff_A_fJAhGCsV8_0),.din(w_dff_A_l1gWUlAh7_0),.clk(gclk));
	jdff dff_A_fJAhGCsV8_0(.dout(w_dff_A_GOtZUZXK5_0),.din(w_dff_A_fJAhGCsV8_0),.clk(gclk));
	jdff dff_A_GOtZUZXK5_0(.dout(w_dff_A_hZuXznYA9_0),.din(w_dff_A_GOtZUZXK5_0),.clk(gclk));
	jdff dff_A_hZuXznYA9_0(.dout(w_dff_A_sL6QDJKH0_0),.din(w_dff_A_hZuXznYA9_0),.clk(gclk));
	jdff dff_A_sL6QDJKH0_0(.dout(w_dff_A_DtTSog067_0),.din(w_dff_A_sL6QDJKH0_0),.clk(gclk));
	jdff dff_A_DtTSog067_0(.dout(w_dff_A_tbGC8tld8_0),.din(w_dff_A_DtTSog067_0),.clk(gclk));
	jdff dff_A_tbGC8tld8_0(.dout(w_dff_A_64JxdCda3_0),.din(w_dff_A_tbGC8tld8_0),.clk(gclk));
	jdff dff_A_64JxdCda3_0(.dout(w_dff_A_WeCI0N5o2_0),.din(w_dff_A_64JxdCda3_0),.clk(gclk));
	jdff dff_A_WeCI0N5o2_0(.dout(w_dff_A_mJuGf5gD4_0),.din(w_dff_A_WeCI0N5o2_0),.clk(gclk));
	jdff dff_A_mJuGf5gD4_0(.dout(w_dff_A_IvTJn8Y02_0),.din(w_dff_A_mJuGf5gD4_0),.clk(gclk));
	jdff dff_A_IvTJn8Y02_0(.dout(f56),.din(w_dff_A_IvTJn8Y02_0),.clk(gclk));
	jdff dff_A_INrlTL4v6_2(.dout(w_dff_A_dzJBt3XK3_0),.din(w_dff_A_INrlTL4v6_2),.clk(gclk));
	jdff dff_A_dzJBt3XK3_0(.dout(w_dff_A_Vr2TkBZ93_0),.din(w_dff_A_dzJBt3XK3_0),.clk(gclk));
	jdff dff_A_Vr2TkBZ93_0(.dout(w_dff_A_Flr0wM298_0),.din(w_dff_A_Vr2TkBZ93_0),.clk(gclk));
	jdff dff_A_Flr0wM298_0(.dout(w_dff_A_Kc2qisMs5_0),.din(w_dff_A_Flr0wM298_0),.clk(gclk));
	jdff dff_A_Kc2qisMs5_0(.dout(w_dff_A_E2dKC4Xb7_0),.din(w_dff_A_Kc2qisMs5_0),.clk(gclk));
	jdff dff_A_E2dKC4Xb7_0(.dout(w_dff_A_n5ZDpFvC7_0),.din(w_dff_A_E2dKC4Xb7_0),.clk(gclk));
	jdff dff_A_n5ZDpFvC7_0(.dout(w_dff_A_2R71b5u67_0),.din(w_dff_A_n5ZDpFvC7_0),.clk(gclk));
	jdff dff_A_2R71b5u67_0(.dout(w_dff_A_Oqrq1htL2_0),.din(w_dff_A_2R71b5u67_0),.clk(gclk));
	jdff dff_A_Oqrq1htL2_0(.dout(w_dff_A_sHi9szqV5_0),.din(w_dff_A_Oqrq1htL2_0),.clk(gclk));
	jdff dff_A_sHi9szqV5_0(.dout(w_dff_A_YAPjvI9S1_0),.din(w_dff_A_sHi9szqV5_0),.clk(gclk));
	jdff dff_A_YAPjvI9S1_0(.dout(w_dff_A_nQ6HQWd80_0),.din(w_dff_A_YAPjvI9S1_0),.clk(gclk));
	jdff dff_A_nQ6HQWd80_0(.dout(w_dff_A_iXgVBlFM2_0),.din(w_dff_A_nQ6HQWd80_0),.clk(gclk));
	jdff dff_A_iXgVBlFM2_0(.dout(w_dff_A_444c1OEZ5_0),.din(w_dff_A_iXgVBlFM2_0),.clk(gclk));
	jdff dff_A_444c1OEZ5_0(.dout(w_dff_A_JLHjEdjq5_0),.din(w_dff_A_444c1OEZ5_0),.clk(gclk));
	jdff dff_A_JLHjEdjq5_0(.dout(w_dff_A_MUAHkjCu1_0),.din(w_dff_A_JLHjEdjq5_0),.clk(gclk));
	jdff dff_A_MUAHkjCu1_0(.dout(w_dff_A_7XJAZRSW1_0),.din(w_dff_A_MUAHkjCu1_0),.clk(gclk));
	jdff dff_A_7XJAZRSW1_0(.dout(w_dff_A_5Je0kVlb2_0),.din(w_dff_A_7XJAZRSW1_0),.clk(gclk));
	jdff dff_A_5Je0kVlb2_0(.dout(w_dff_A_UY1BCc0f6_0),.din(w_dff_A_5Je0kVlb2_0),.clk(gclk));
	jdff dff_A_UY1BCc0f6_0(.dout(w_dff_A_eQQGW6GA3_0),.din(w_dff_A_UY1BCc0f6_0),.clk(gclk));
	jdff dff_A_eQQGW6GA3_0(.dout(w_dff_A_ZxoQJk0A0_0),.din(w_dff_A_eQQGW6GA3_0),.clk(gclk));
	jdff dff_A_ZxoQJk0A0_0(.dout(w_dff_A_p3P2CgPH2_0),.din(w_dff_A_ZxoQJk0A0_0),.clk(gclk));
	jdff dff_A_p3P2CgPH2_0(.dout(w_dff_A_IUk9R3nt1_0),.din(w_dff_A_p3P2CgPH2_0),.clk(gclk));
	jdff dff_A_IUk9R3nt1_0(.dout(w_dff_A_Zna0LaSe0_0),.din(w_dff_A_IUk9R3nt1_0),.clk(gclk));
	jdff dff_A_Zna0LaSe0_0(.dout(w_dff_A_Y59SHbD43_0),.din(w_dff_A_Zna0LaSe0_0),.clk(gclk));
	jdff dff_A_Y59SHbD43_0(.dout(w_dff_A_lpdVdwYS8_0),.din(w_dff_A_Y59SHbD43_0),.clk(gclk));
	jdff dff_A_lpdVdwYS8_0(.dout(w_dff_A_wDZmmeic0_0),.din(w_dff_A_lpdVdwYS8_0),.clk(gclk));
	jdff dff_A_wDZmmeic0_0(.dout(w_dff_A_C0U5MoLj7_0),.din(w_dff_A_wDZmmeic0_0),.clk(gclk));
	jdff dff_A_C0U5MoLj7_0(.dout(w_dff_A_gNRhiPIO4_0),.din(w_dff_A_C0U5MoLj7_0),.clk(gclk));
	jdff dff_A_gNRhiPIO4_0(.dout(w_dff_A_lRndsGCf1_0),.din(w_dff_A_gNRhiPIO4_0),.clk(gclk));
	jdff dff_A_lRndsGCf1_0(.dout(w_dff_A_FchBVqcv4_0),.din(w_dff_A_lRndsGCf1_0),.clk(gclk));
	jdff dff_A_FchBVqcv4_0(.dout(w_dff_A_xRP8DBtF8_0),.din(w_dff_A_FchBVqcv4_0),.clk(gclk));
	jdff dff_A_xRP8DBtF8_0(.dout(w_dff_A_ySjBwn3y9_0),.din(w_dff_A_xRP8DBtF8_0),.clk(gclk));
	jdff dff_A_ySjBwn3y9_0(.dout(w_dff_A_hlCxXxgl1_0),.din(w_dff_A_ySjBwn3y9_0),.clk(gclk));
	jdff dff_A_hlCxXxgl1_0(.dout(w_dff_A_TYLYzYKD6_0),.din(w_dff_A_hlCxXxgl1_0),.clk(gclk));
	jdff dff_A_TYLYzYKD6_0(.dout(w_dff_A_YZ6lbGs56_0),.din(w_dff_A_TYLYzYKD6_0),.clk(gclk));
	jdff dff_A_YZ6lbGs56_0(.dout(w_dff_A_N3zUviHw5_0),.din(w_dff_A_YZ6lbGs56_0),.clk(gclk));
	jdff dff_A_N3zUviHw5_0(.dout(w_dff_A_pTv2ymDG2_0),.din(w_dff_A_N3zUviHw5_0),.clk(gclk));
	jdff dff_A_pTv2ymDG2_0(.dout(w_dff_A_265Slivm5_0),.din(w_dff_A_pTv2ymDG2_0),.clk(gclk));
	jdff dff_A_265Slivm5_0(.dout(w_dff_A_YhOHnR7d2_0),.din(w_dff_A_265Slivm5_0),.clk(gclk));
	jdff dff_A_YhOHnR7d2_0(.dout(w_dff_A_kPPJ7LfZ7_0),.din(w_dff_A_YhOHnR7d2_0),.clk(gclk));
	jdff dff_A_kPPJ7LfZ7_0(.dout(w_dff_A_bJQdLUD66_0),.din(w_dff_A_kPPJ7LfZ7_0),.clk(gclk));
	jdff dff_A_bJQdLUD66_0(.dout(w_dff_A_fUKoKbHh6_0),.din(w_dff_A_bJQdLUD66_0),.clk(gclk));
	jdff dff_A_fUKoKbHh6_0(.dout(w_dff_A_jVbtG9B81_0),.din(w_dff_A_fUKoKbHh6_0),.clk(gclk));
	jdff dff_A_jVbtG9B81_0(.dout(w_dff_A_a3rkbpN66_0),.din(w_dff_A_jVbtG9B81_0),.clk(gclk));
	jdff dff_A_a3rkbpN66_0(.dout(w_dff_A_HV3QeVWQ7_0),.din(w_dff_A_a3rkbpN66_0),.clk(gclk));
	jdff dff_A_HV3QeVWQ7_0(.dout(w_dff_A_msFJJVRT6_0),.din(w_dff_A_HV3QeVWQ7_0),.clk(gclk));
	jdff dff_A_msFJJVRT6_0(.dout(w_dff_A_duC2MSQt9_0),.din(w_dff_A_msFJJVRT6_0),.clk(gclk));
	jdff dff_A_duC2MSQt9_0(.dout(w_dff_A_9fyzrEba9_0),.din(w_dff_A_duC2MSQt9_0),.clk(gclk));
	jdff dff_A_9fyzrEba9_0(.dout(w_dff_A_WfR8fa7O6_0),.din(w_dff_A_9fyzrEba9_0),.clk(gclk));
	jdff dff_A_WfR8fa7O6_0(.dout(w_dff_A_SO0ETjHd5_0),.din(w_dff_A_WfR8fa7O6_0),.clk(gclk));
	jdff dff_A_SO0ETjHd5_0(.dout(w_dff_A_GpAnB8xc4_0),.din(w_dff_A_SO0ETjHd5_0),.clk(gclk));
	jdff dff_A_GpAnB8xc4_0(.dout(w_dff_A_oGlMQOfk5_0),.din(w_dff_A_GpAnB8xc4_0),.clk(gclk));
	jdff dff_A_oGlMQOfk5_0(.dout(w_dff_A_apJ3dJcE4_0),.din(w_dff_A_oGlMQOfk5_0),.clk(gclk));
	jdff dff_A_apJ3dJcE4_0(.dout(w_dff_A_170vd5ct5_0),.din(w_dff_A_apJ3dJcE4_0),.clk(gclk));
	jdff dff_A_170vd5ct5_0(.dout(w_dff_A_Tvp8A8RG7_0),.din(w_dff_A_170vd5ct5_0),.clk(gclk));
	jdff dff_A_Tvp8A8RG7_0(.dout(w_dff_A_8Mxb0QGd8_0),.din(w_dff_A_Tvp8A8RG7_0),.clk(gclk));
	jdff dff_A_8Mxb0QGd8_0(.dout(w_dff_A_OFto8a2a2_0),.din(w_dff_A_8Mxb0QGd8_0),.clk(gclk));
	jdff dff_A_OFto8a2a2_0(.dout(w_dff_A_925AHoRn1_0),.din(w_dff_A_OFto8a2a2_0),.clk(gclk));
	jdff dff_A_925AHoRn1_0(.dout(w_dff_A_rS0iKfSZ9_0),.din(w_dff_A_925AHoRn1_0),.clk(gclk));
	jdff dff_A_rS0iKfSZ9_0(.dout(w_dff_A_OUfcnEjW0_0),.din(w_dff_A_rS0iKfSZ9_0),.clk(gclk));
	jdff dff_A_OUfcnEjW0_0(.dout(w_dff_A_ldx1rHEh9_0),.din(w_dff_A_OUfcnEjW0_0),.clk(gclk));
	jdff dff_A_ldx1rHEh9_0(.dout(w_dff_A_PZgLZaZI0_0),.din(w_dff_A_ldx1rHEh9_0),.clk(gclk));
	jdff dff_A_PZgLZaZI0_0(.dout(w_dff_A_CInfOAQj1_0),.din(w_dff_A_PZgLZaZI0_0),.clk(gclk));
	jdff dff_A_CInfOAQj1_0(.dout(w_dff_A_yTNymAn70_0),.din(w_dff_A_CInfOAQj1_0),.clk(gclk));
	jdff dff_A_yTNymAn70_0(.dout(w_dff_A_RzedOrNj5_0),.din(w_dff_A_yTNymAn70_0),.clk(gclk));
	jdff dff_A_RzedOrNj5_0(.dout(w_dff_A_GEHMCHoa3_0),.din(w_dff_A_RzedOrNj5_0),.clk(gclk));
	jdff dff_A_GEHMCHoa3_0(.dout(w_dff_A_ddrCs4lg1_0),.din(w_dff_A_GEHMCHoa3_0),.clk(gclk));
	jdff dff_A_ddrCs4lg1_0(.dout(w_dff_A_vNi7B1Gi5_0),.din(w_dff_A_ddrCs4lg1_0),.clk(gclk));
	jdff dff_A_vNi7B1Gi5_0(.dout(w_dff_A_t1ePrhYd1_0),.din(w_dff_A_vNi7B1Gi5_0),.clk(gclk));
	jdff dff_A_t1ePrhYd1_0(.dout(f57),.din(w_dff_A_t1ePrhYd1_0),.clk(gclk));
	jdff dff_A_IAZs4o3E0_2(.dout(w_dff_A_ItinrNbG6_0),.din(w_dff_A_IAZs4o3E0_2),.clk(gclk));
	jdff dff_A_ItinrNbG6_0(.dout(w_dff_A_4Abqw0o03_0),.din(w_dff_A_ItinrNbG6_0),.clk(gclk));
	jdff dff_A_4Abqw0o03_0(.dout(w_dff_A_RO8TXVEV8_0),.din(w_dff_A_4Abqw0o03_0),.clk(gclk));
	jdff dff_A_RO8TXVEV8_0(.dout(w_dff_A_b4iNdPyV0_0),.din(w_dff_A_RO8TXVEV8_0),.clk(gclk));
	jdff dff_A_b4iNdPyV0_0(.dout(w_dff_A_RQdxJYaD5_0),.din(w_dff_A_b4iNdPyV0_0),.clk(gclk));
	jdff dff_A_RQdxJYaD5_0(.dout(w_dff_A_gbjOaIdn4_0),.din(w_dff_A_RQdxJYaD5_0),.clk(gclk));
	jdff dff_A_gbjOaIdn4_0(.dout(w_dff_A_64MVXsYw9_0),.din(w_dff_A_gbjOaIdn4_0),.clk(gclk));
	jdff dff_A_64MVXsYw9_0(.dout(w_dff_A_pgHrHjs61_0),.din(w_dff_A_64MVXsYw9_0),.clk(gclk));
	jdff dff_A_pgHrHjs61_0(.dout(w_dff_A_bOH4RhaY2_0),.din(w_dff_A_pgHrHjs61_0),.clk(gclk));
	jdff dff_A_bOH4RhaY2_0(.dout(w_dff_A_LBoqBJPW2_0),.din(w_dff_A_bOH4RhaY2_0),.clk(gclk));
	jdff dff_A_LBoqBJPW2_0(.dout(w_dff_A_2BYgK6QY3_0),.din(w_dff_A_LBoqBJPW2_0),.clk(gclk));
	jdff dff_A_2BYgK6QY3_0(.dout(w_dff_A_QFF96nlz6_0),.din(w_dff_A_2BYgK6QY3_0),.clk(gclk));
	jdff dff_A_QFF96nlz6_0(.dout(w_dff_A_4H0prr0p5_0),.din(w_dff_A_QFF96nlz6_0),.clk(gclk));
	jdff dff_A_4H0prr0p5_0(.dout(w_dff_A_q6uyiPbh9_0),.din(w_dff_A_4H0prr0p5_0),.clk(gclk));
	jdff dff_A_q6uyiPbh9_0(.dout(w_dff_A_g0egDFDs4_0),.din(w_dff_A_q6uyiPbh9_0),.clk(gclk));
	jdff dff_A_g0egDFDs4_0(.dout(w_dff_A_j0XC9rSh5_0),.din(w_dff_A_g0egDFDs4_0),.clk(gclk));
	jdff dff_A_j0XC9rSh5_0(.dout(w_dff_A_2l2u3Yf81_0),.din(w_dff_A_j0XC9rSh5_0),.clk(gclk));
	jdff dff_A_2l2u3Yf81_0(.dout(w_dff_A_oOWWJo2F3_0),.din(w_dff_A_2l2u3Yf81_0),.clk(gclk));
	jdff dff_A_oOWWJo2F3_0(.dout(w_dff_A_plnOhLod1_0),.din(w_dff_A_oOWWJo2F3_0),.clk(gclk));
	jdff dff_A_plnOhLod1_0(.dout(w_dff_A_oOP4xdlA8_0),.din(w_dff_A_plnOhLod1_0),.clk(gclk));
	jdff dff_A_oOP4xdlA8_0(.dout(w_dff_A_kjq3835h5_0),.din(w_dff_A_oOP4xdlA8_0),.clk(gclk));
	jdff dff_A_kjq3835h5_0(.dout(w_dff_A_Ggb9Bo7a0_0),.din(w_dff_A_kjq3835h5_0),.clk(gclk));
	jdff dff_A_Ggb9Bo7a0_0(.dout(w_dff_A_SfBCPdp25_0),.din(w_dff_A_Ggb9Bo7a0_0),.clk(gclk));
	jdff dff_A_SfBCPdp25_0(.dout(w_dff_A_de5F7q3x7_0),.din(w_dff_A_SfBCPdp25_0),.clk(gclk));
	jdff dff_A_de5F7q3x7_0(.dout(w_dff_A_YquGHsyh8_0),.din(w_dff_A_de5F7q3x7_0),.clk(gclk));
	jdff dff_A_YquGHsyh8_0(.dout(w_dff_A_woFHH4tr9_0),.din(w_dff_A_YquGHsyh8_0),.clk(gclk));
	jdff dff_A_woFHH4tr9_0(.dout(w_dff_A_oyGr7D3X5_0),.din(w_dff_A_woFHH4tr9_0),.clk(gclk));
	jdff dff_A_oyGr7D3X5_0(.dout(w_dff_A_Ckd77GBL9_0),.din(w_dff_A_oyGr7D3X5_0),.clk(gclk));
	jdff dff_A_Ckd77GBL9_0(.dout(w_dff_A_otg2TxFE9_0),.din(w_dff_A_Ckd77GBL9_0),.clk(gclk));
	jdff dff_A_otg2TxFE9_0(.dout(w_dff_A_1YtZ9VoF9_0),.din(w_dff_A_otg2TxFE9_0),.clk(gclk));
	jdff dff_A_1YtZ9VoF9_0(.dout(w_dff_A_UFa0VRPK7_0),.din(w_dff_A_1YtZ9VoF9_0),.clk(gclk));
	jdff dff_A_UFa0VRPK7_0(.dout(w_dff_A_y2Cpwbtj9_0),.din(w_dff_A_UFa0VRPK7_0),.clk(gclk));
	jdff dff_A_y2Cpwbtj9_0(.dout(w_dff_A_z2CMdxhl6_0),.din(w_dff_A_y2Cpwbtj9_0),.clk(gclk));
	jdff dff_A_z2CMdxhl6_0(.dout(w_dff_A_dsoI6mN01_0),.din(w_dff_A_z2CMdxhl6_0),.clk(gclk));
	jdff dff_A_dsoI6mN01_0(.dout(w_dff_A_SXfYOpZi7_0),.din(w_dff_A_dsoI6mN01_0),.clk(gclk));
	jdff dff_A_SXfYOpZi7_0(.dout(w_dff_A_VbfBQ0OQ0_0),.din(w_dff_A_SXfYOpZi7_0),.clk(gclk));
	jdff dff_A_VbfBQ0OQ0_0(.dout(w_dff_A_Hpj35L0u4_0),.din(w_dff_A_VbfBQ0OQ0_0),.clk(gclk));
	jdff dff_A_Hpj35L0u4_0(.dout(w_dff_A_pZrId7J13_0),.din(w_dff_A_Hpj35L0u4_0),.clk(gclk));
	jdff dff_A_pZrId7J13_0(.dout(w_dff_A_swZSLd5s3_0),.din(w_dff_A_pZrId7J13_0),.clk(gclk));
	jdff dff_A_swZSLd5s3_0(.dout(w_dff_A_APbaCdFl8_0),.din(w_dff_A_swZSLd5s3_0),.clk(gclk));
	jdff dff_A_APbaCdFl8_0(.dout(w_dff_A_jq9MgPEF3_0),.din(w_dff_A_APbaCdFl8_0),.clk(gclk));
	jdff dff_A_jq9MgPEF3_0(.dout(w_dff_A_bjLtbmY60_0),.din(w_dff_A_jq9MgPEF3_0),.clk(gclk));
	jdff dff_A_bjLtbmY60_0(.dout(w_dff_A_JBBcEA4Z7_0),.din(w_dff_A_bjLtbmY60_0),.clk(gclk));
	jdff dff_A_JBBcEA4Z7_0(.dout(w_dff_A_a7ZLB98X2_0),.din(w_dff_A_JBBcEA4Z7_0),.clk(gclk));
	jdff dff_A_a7ZLB98X2_0(.dout(w_dff_A_iJJYMslN2_0),.din(w_dff_A_a7ZLB98X2_0),.clk(gclk));
	jdff dff_A_iJJYMslN2_0(.dout(w_dff_A_o1BmuXI45_0),.din(w_dff_A_iJJYMslN2_0),.clk(gclk));
	jdff dff_A_o1BmuXI45_0(.dout(w_dff_A_qtGxJDtF0_0),.din(w_dff_A_o1BmuXI45_0),.clk(gclk));
	jdff dff_A_qtGxJDtF0_0(.dout(w_dff_A_7dFCxesR8_0),.din(w_dff_A_qtGxJDtF0_0),.clk(gclk));
	jdff dff_A_7dFCxesR8_0(.dout(w_dff_A_ZY7bDPDY5_0),.din(w_dff_A_7dFCxesR8_0),.clk(gclk));
	jdff dff_A_ZY7bDPDY5_0(.dout(w_dff_A_CglyVY7S2_0),.din(w_dff_A_ZY7bDPDY5_0),.clk(gclk));
	jdff dff_A_CglyVY7S2_0(.dout(w_dff_A_OUuJVZMo4_0),.din(w_dff_A_CglyVY7S2_0),.clk(gclk));
	jdff dff_A_OUuJVZMo4_0(.dout(w_dff_A_KeMazQGi9_0),.din(w_dff_A_OUuJVZMo4_0),.clk(gclk));
	jdff dff_A_KeMazQGi9_0(.dout(w_dff_A_SCOSbgDQ3_0),.din(w_dff_A_KeMazQGi9_0),.clk(gclk));
	jdff dff_A_SCOSbgDQ3_0(.dout(w_dff_A_0whYsXA34_0),.din(w_dff_A_SCOSbgDQ3_0),.clk(gclk));
	jdff dff_A_0whYsXA34_0(.dout(w_dff_A_Wj0ClU7E4_0),.din(w_dff_A_0whYsXA34_0),.clk(gclk));
	jdff dff_A_Wj0ClU7E4_0(.dout(w_dff_A_2GVeQnEa6_0),.din(w_dff_A_Wj0ClU7E4_0),.clk(gclk));
	jdff dff_A_2GVeQnEa6_0(.dout(w_dff_A_Usl54Erk1_0),.din(w_dff_A_2GVeQnEa6_0),.clk(gclk));
	jdff dff_A_Usl54Erk1_0(.dout(w_dff_A_1wMbp6Lr0_0),.din(w_dff_A_Usl54Erk1_0),.clk(gclk));
	jdff dff_A_1wMbp6Lr0_0(.dout(w_dff_A_2UqSuI3a2_0),.din(w_dff_A_1wMbp6Lr0_0),.clk(gclk));
	jdff dff_A_2UqSuI3a2_0(.dout(w_dff_A_8AN3YywG6_0),.din(w_dff_A_2UqSuI3a2_0),.clk(gclk));
	jdff dff_A_8AN3YywG6_0(.dout(w_dff_A_Qj5uX7bo9_0),.din(w_dff_A_8AN3YywG6_0),.clk(gclk));
	jdff dff_A_Qj5uX7bo9_0(.dout(w_dff_A_zhklAO6a8_0),.din(w_dff_A_Qj5uX7bo9_0),.clk(gclk));
	jdff dff_A_zhklAO6a8_0(.dout(w_dff_A_Ld80DM2H1_0),.din(w_dff_A_zhklAO6a8_0),.clk(gclk));
	jdff dff_A_Ld80DM2H1_0(.dout(w_dff_A_68qUDKBA9_0),.din(w_dff_A_Ld80DM2H1_0),.clk(gclk));
	jdff dff_A_68qUDKBA9_0(.dout(w_dff_A_J5JLUTcn0_0),.din(w_dff_A_68qUDKBA9_0),.clk(gclk));
	jdff dff_A_J5JLUTcn0_0(.dout(w_dff_A_D3oyc61M9_0),.din(w_dff_A_J5JLUTcn0_0),.clk(gclk));
	jdff dff_A_D3oyc61M9_0(.dout(w_dff_A_MeCNDPEa6_0),.din(w_dff_A_D3oyc61M9_0),.clk(gclk));
	jdff dff_A_MeCNDPEa6_0(.dout(w_dff_A_dFfcmXB78_0),.din(w_dff_A_MeCNDPEa6_0),.clk(gclk));
	jdff dff_A_dFfcmXB78_0(.dout(f58),.din(w_dff_A_dFfcmXB78_0),.clk(gclk));
	jdff dff_A_bZXjmX1T8_2(.dout(w_dff_A_J0OfzNGE4_0),.din(w_dff_A_bZXjmX1T8_2),.clk(gclk));
	jdff dff_A_J0OfzNGE4_0(.dout(w_dff_A_YxbWi1fC4_0),.din(w_dff_A_J0OfzNGE4_0),.clk(gclk));
	jdff dff_A_YxbWi1fC4_0(.dout(w_dff_A_ijb0lVcg0_0),.din(w_dff_A_YxbWi1fC4_0),.clk(gclk));
	jdff dff_A_ijb0lVcg0_0(.dout(w_dff_A_pAz3CRnI9_0),.din(w_dff_A_ijb0lVcg0_0),.clk(gclk));
	jdff dff_A_pAz3CRnI9_0(.dout(w_dff_A_RJoTSTKc7_0),.din(w_dff_A_pAz3CRnI9_0),.clk(gclk));
	jdff dff_A_RJoTSTKc7_0(.dout(w_dff_A_ojppQPfy7_0),.din(w_dff_A_RJoTSTKc7_0),.clk(gclk));
	jdff dff_A_ojppQPfy7_0(.dout(w_dff_A_whTb4Wka5_0),.din(w_dff_A_ojppQPfy7_0),.clk(gclk));
	jdff dff_A_whTb4Wka5_0(.dout(w_dff_A_auNV7sAo0_0),.din(w_dff_A_whTb4Wka5_0),.clk(gclk));
	jdff dff_A_auNV7sAo0_0(.dout(w_dff_A_kEL4YbMu6_0),.din(w_dff_A_auNV7sAo0_0),.clk(gclk));
	jdff dff_A_kEL4YbMu6_0(.dout(w_dff_A_rblVoy0h1_0),.din(w_dff_A_kEL4YbMu6_0),.clk(gclk));
	jdff dff_A_rblVoy0h1_0(.dout(w_dff_A_9LhXojvx8_0),.din(w_dff_A_rblVoy0h1_0),.clk(gclk));
	jdff dff_A_9LhXojvx8_0(.dout(w_dff_A_iCOWJdkT5_0),.din(w_dff_A_9LhXojvx8_0),.clk(gclk));
	jdff dff_A_iCOWJdkT5_0(.dout(w_dff_A_jJ5Qlu4Y8_0),.din(w_dff_A_iCOWJdkT5_0),.clk(gclk));
	jdff dff_A_jJ5Qlu4Y8_0(.dout(w_dff_A_wuSrx01o9_0),.din(w_dff_A_jJ5Qlu4Y8_0),.clk(gclk));
	jdff dff_A_wuSrx01o9_0(.dout(w_dff_A_PmWPTiZU2_0),.din(w_dff_A_wuSrx01o9_0),.clk(gclk));
	jdff dff_A_PmWPTiZU2_0(.dout(w_dff_A_BxlJGkPT7_0),.din(w_dff_A_PmWPTiZU2_0),.clk(gclk));
	jdff dff_A_BxlJGkPT7_0(.dout(w_dff_A_yZvDAxEX4_0),.din(w_dff_A_BxlJGkPT7_0),.clk(gclk));
	jdff dff_A_yZvDAxEX4_0(.dout(w_dff_A_bPdAc6T62_0),.din(w_dff_A_yZvDAxEX4_0),.clk(gclk));
	jdff dff_A_bPdAc6T62_0(.dout(w_dff_A_eHi8f8rP6_0),.din(w_dff_A_bPdAc6T62_0),.clk(gclk));
	jdff dff_A_eHi8f8rP6_0(.dout(w_dff_A_KaaP93St6_0),.din(w_dff_A_eHi8f8rP6_0),.clk(gclk));
	jdff dff_A_KaaP93St6_0(.dout(w_dff_A_rEQf91VJ5_0),.din(w_dff_A_KaaP93St6_0),.clk(gclk));
	jdff dff_A_rEQf91VJ5_0(.dout(w_dff_A_YAN38V8C2_0),.din(w_dff_A_rEQf91VJ5_0),.clk(gclk));
	jdff dff_A_YAN38V8C2_0(.dout(w_dff_A_cZOdT8la7_0),.din(w_dff_A_YAN38V8C2_0),.clk(gclk));
	jdff dff_A_cZOdT8la7_0(.dout(w_dff_A_ekVHlDMz7_0),.din(w_dff_A_cZOdT8la7_0),.clk(gclk));
	jdff dff_A_ekVHlDMz7_0(.dout(w_dff_A_gOBp3VlD1_0),.din(w_dff_A_ekVHlDMz7_0),.clk(gclk));
	jdff dff_A_gOBp3VlD1_0(.dout(w_dff_A_EIOPK32F7_0),.din(w_dff_A_gOBp3VlD1_0),.clk(gclk));
	jdff dff_A_EIOPK32F7_0(.dout(w_dff_A_wsehX8vH1_0),.din(w_dff_A_EIOPK32F7_0),.clk(gclk));
	jdff dff_A_wsehX8vH1_0(.dout(w_dff_A_EXdmOgX76_0),.din(w_dff_A_wsehX8vH1_0),.clk(gclk));
	jdff dff_A_EXdmOgX76_0(.dout(w_dff_A_pD8UYqFN8_0),.din(w_dff_A_EXdmOgX76_0),.clk(gclk));
	jdff dff_A_pD8UYqFN8_0(.dout(w_dff_A_5HkGXnDh4_0),.din(w_dff_A_pD8UYqFN8_0),.clk(gclk));
	jdff dff_A_5HkGXnDh4_0(.dout(w_dff_A_6mbR5O7N0_0),.din(w_dff_A_5HkGXnDh4_0),.clk(gclk));
	jdff dff_A_6mbR5O7N0_0(.dout(w_dff_A_k0MGrKmU1_0),.din(w_dff_A_6mbR5O7N0_0),.clk(gclk));
	jdff dff_A_k0MGrKmU1_0(.dout(w_dff_A_jEGbxiky3_0),.din(w_dff_A_k0MGrKmU1_0),.clk(gclk));
	jdff dff_A_jEGbxiky3_0(.dout(w_dff_A_tYzpPAIH3_0),.din(w_dff_A_jEGbxiky3_0),.clk(gclk));
	jdff dff_A_tYzpPAIH3_0(.dout(w_dff_A_wnoqg8Av2_0),.din(w_dff_A_tYzpPAIH3_0),.clk(gclk));
	jdff dff_A_wnoqg8Av2_0(.dout(w_dff_A_Q8slLJEZ5_0),.din(w_dff_A_wnoqg8Av2_0),.clk(gclk));
	jdff dff_A_Q8slLJEZ5_0(.dout(w_dff_A_alHIAczq5_0),.din(w_dff_A_Q8slLJEZ5_0),.clk(gclk));
	jdff dff_A_alHIAczq5_0(.dout(w_dff_A_GF0mvWa02_0),.din(w_dff_A_alHIAczq5_0),.clk(gclk));
	jdff dff_A_GF0mvWa02_0(.dout(w_dff_A_f9u2wKKo3_0),.din(w_dff_A_GF0mvWa02_0),.clk(gclk));
	jdff dff_A_f9u2wKKo3_0(.dout(w_dff_A_a6ZncgSM3_0),.din(w_dff_A_f9u2wKKo3_0),.clk(gclk));
	jdff dff_A_a6ZncgSM3_0(.dout(w_dff_A_vMU3Xfbq8_0),.din(w_dff_A_a6ZncgSM3_0),.clk(gclk));
	jdff dff_A_vMU3Xfbq8_0(.dout(w_dff_A_0qqEFaxx2_0),.din(w_dff_A_vMU3Xfbq8_0),.clk(gclk));
	jdff dff_A_0qqEFaxx2_0(.dout(w_dff_A_jsaQSO5d6_0),.din(w_dff_A_0qqEFaxx2_0),.clk(gclk));
	jdff dff_A_jsaQSO5d6_0(.dout(w_dff_A_DLeea00d6_0),.din(w_dff_A_jsaQSO5d6_0),.clk(gclk));
	jdff dff_A_DLeea00d6_0(.dout(w_dff_A_fsUUoAD81_0),.din(w_dff_A_DLeea00d6_0),.clk(gclk));
	jdff dff_A_fsUUoAD81_0(.dout(w_dff_A_AFyNESGA8_0),.din(w_dff_A_fsUUoAD81_0),.clk(gclk));
	jdff dff_A_AFyNESGA8_0(.dout(w_dff_A_Hrp0jJln5_0),.din(w_dff_A_AFyNESGA8_0),.clk(gclk));
	jdff dff_A_Hrp0jJln5_0(.dout(w_dff_A_M8Sx6SPF5_0),.din(w_dff_A_Hrp0jJln5_0),.clk(gclk));
	jdff dff_A_M8Sx6SPF5_0(.dout(w_dff_A_P0sRalXm7_0),.din(w_dff_A_M8Sx6SPF5_0),.clk(gclk));
	jdff dff_A_P0sRalXm7_0(.dout(w_dff_A_5CAqbjeG2_0),.din(w_dff_A_P0sRalXm7_0),.clk(gclk));
	jdff dff_A_5CAqbjeG2_0(.dout(w_dff_A_se3ZFNKb6_0),.din(w_dff_A_5CAqbjeG2_0),.clk(gclk));
	jdff dff_A_se3ZFNKb6_0(.dout(w_dff_A_93317jFh2_0),.din(w_dff_A_se3ZFNKb6_0),.clk(gclk));
	jdff dff_A_93317jFh2_0(.dout(w_dff_A_D3bY47Lm8_0),.din(w_dff_A_93317jFh2_0),.clk(gclk));
	jdff dff_A_D3bY47Lm8_0(.dout(w_dff_A_ezXm4KjA9_0),.din(w_dff_A_D3bY47Lm8_0),.clk(gclk));
	jdff dff_A_ezXm4KjA9_0(.dout(w_dff_A_mgudidAW3_0),.din(w_dff_A_ezXm4KjA9_0),.clk(gclk));
	jdff dff_A_mgudidAW3_0(.dout(w_dff_A_RXtlG59c6_0),.din(w_dff_A_mgudidAW3_0),.clk(gclk));
	jdff dff_A_RXtlG59c6_0(.dout(w_dff_A_RsBttq8o1_0),.din(w_dff_A_RXtlG59c6_0),.clk(gclk));
	jdff dff_A_RsBttq8o1_0(.dout(w_dff_A_IFH0cgii4_0),.din(w_dff_A_RsBttq8o1_0),.clk(gclk));
	jdff dff_A_IFH0cgii4_0(.dout(w_dff_A_WqwQnJIn4_0),.din(w_dff_A_IFH0cgii4_0),.clk(gclk));
	jdff dff_A_WqwQnJIn4_0(.dout(w_dff_A_EMUHb9yI1_0),.din(w_dff_A_WqwQnJIn4_0),.clk(gclk));
	jdff dff_A_EMUHb9yI1_0(.dout(w_dff_A_OaT702BY1_0),.din(w_dff_A_EMUHb9yI1_0),.clk(gclk));
	jdff dff_A_OaT702BY1_0(.dout(w_dff_A_MPEtOBkU2_0),.din(w_dff_A_OaT702BY1_0),.clk(gclk));
	jdff dff_A_MPEtOBkU2_0(.dout(w_dff_A_obS70QOw1_0),.din(w_dff_A_MPEtOBkU2_0),.clk(gclk));
	jdff dff_A_obS70QOw1_0(.dout(w_dff_A_mJo0oCdy0_0),.din(w_dff_A_obS70QOw1_0),.clk(gclk));
	jdff dff_A_mJo0oCdy0_0(.dout(w_dff_A_LXYObhyu6_0),.din(w_dff_A_mJo0oCdy0_0),.clk(gclk));
	jdff dff_A_LXYObhyu6_0(.dout(w_dff_A_IA2TyC683_0),.din(w_dff_A_LXYObhyu6_0),.clk(gclk));
	jdff dff_A_IA2TyC683_0(.dout(w_dff_A_eCTgGWm33_0),.din(w_dff_A_IA2TyC683_0),.clk(gclk));
	jdff dff_A_eCTgGWm33_0(.dout(f59),.din(w_dff_A_eCTgGWm33_0),.clk(gclk));
	jdff dff_A_73F8XiAD0_2(.dout(w_dff_A_iPKVGkco1_0),.din(w_dff_A_73F8XiAD0_2),.clk(gclk));
	jdff dff_A_iPKVGkco1_0(.dout(w_dff_A_6nfmMa9U8_0),.din(w_dff_A_iPKVGkco1_0),.clk(gclk));
	jdff dff_A_6nfmMa9U8_0(.dout(w_dff_A_rLBPzbBR9_0),.din(w_dff_A_6nfmMa9U8_0),.clk(gclk));
	jdff dff_A_rLBPzbBR9_0(.dout(w_dff_A_rtDu19XC0_0),.din(w_dff_A_rLBPzbBR9_0),.clk(gclk));
	jdff dff_A_rtDu19XC0_0(.dout(w_dff_A_XfQEC6OM4_0),.din(w_dff_A_rtDu19XC0_0),.clk(gclk));
	jdff dff_A_XfQEC6OM4_0(.dout(w_dff_A_CB6r4lDG5_0),.din(w_dff_A_XfQEC6OM4_0),.clk(gclk));
	jdff dff_A_CB6r4lDG5_0(.dout(w_dff_A_f9s9udqi9_0),.din(w_dff_A_CB6r4lDG5_0),.clk(gclk));
	jdff dff_A_f9s9udqi9_0(.dout(w_dff_A_0vRYqZP50_0),.din(w_dff_A_f9s9udqi9_0),.clk(gclk));
	jdff dff_A_0vRYqZP50_0(.dout(w_dff_A_vVkDP0P28_0),.din(w_dff_A_0vRYqZP50_0),.clk(gclk));
	jdff dff_A_vVkDP0P28_0(.dout(w_dff_A_61KF65Qe4_0),.din(w_dff_A_vVkDP0P28_0),.clk(gclk));
	jdff dff_A_61KF65Qe4_0(.dout(w_dff_A_6F1CRKmN5_0),.din(w_dff_A_61KF65Qe4_0),.clk(gclk));
	jdff dff_A_6F1CRKmN5_0(.dout(w_dff_A_LhGzkaqS7_0),.din(w_dff_A_6F1CRKmN5_0),.clk(gclk));
	jdff dff_A_LhGzkaqS7_0(.dout(w_dff_A_P9jAgzKT0_0),.din(w_dff_A_LhGzkaqS7_0),.clk(gclk));
	jdff dff_A_P9jAgzKT0_0(.dout(w_dff_A_SWzMbmyQ7_0),.din(w_dff_A_P9jAgzKT0_0),.clk(gclk));
	jdff dff_A_SWzMbmyQ7_0(.dout(w_dff_A_d1FGqUiP2_0),.din(w_dff_A_SWzMbmyQ7_0),.clk(gclk));
	jdff dff_A_d1FGqUiP2_0(.dout(w_dff_A_gPVPJXCs1_0),.din(w_dff_A_d1FGqUiP2_0),.clk(gclk));
	jdff dff_A_gPVPJXCs1_0(.dout(w_dff_A_w1hs2DSQ8_0),.din(w_dff_A_gPVPJXCs1_0),.clk(gclk));
	jdff dff_A_w1hs2DSQ8_0(.dout(w_dff_A_TjBlvOuY0_0),.din(w_dff_A_w1hs2DSQ8_0),.clk(gclk));
	jdff dff_A_TjBlvOuY0_0(.dout(w_dff_A_HXYImnU18_0),.din(w_dff_A_TjBlvOuY0_0),.clk(gclk));
	jdff dff_A_HXYImnU18_0(.dout(w_dff_A_XpaLSiGt5_0),.din(w_dff_A_HXYImnU18_0),.clk(gclk));
	jdff dff_A_XpaLSiGt5_0(.dout(w_dff_A_PUf5IYiC5_0),.din(w_dff_A_XpaLSiGt5_0),.clk(gclk));
	jdff dff_A_PUf5IYiC5_0(.dout(w_dff_A_Mer49gxn2_0),.din(w_dff_A_PUf5IYiC5_0),.clk(gclk));
	jdff dff_A_Mer49gxn2_0(.dout(w_dff_A_qi5lk1194_0),.din(w_dff_A_Mer49gxn2_0),.clk(gclk));
	jdff dff_A_qi5lk1194_0(.dout(w_dff_A_zSOTXPk00_0),.din(w_dff_A_qi5lk1194_0),.clk(gclk));
	jdff dff_A_zSOTXPk00_0(.dout(w_dff_A_w7WMnjLN2_0),.din(w_dff_A_zSOTXPk00_0),.clk(gclk));
	jdff dff_A_w7WMnjLN2_0(.dout(w_dff_A_adGmR87B9_0),.din(w_dff_A_w7WMnjLN2_0),.clk(gclk));
	jdff dff_A_adGmR87B9_0(.dout(w_dff_A_KZBXlJhR1_0),.din(w_dff_A_adGmR87B9_0),.clk(gclk));
	jdff dff_A_KZBXlJhR1_0(.dout(w_dff_A_jjFgBrHF1_0),.din(w_dff_A_KZBXlJhR1_0),.clk(gclk));
	jdff dff_A_jjFgBrHF1_0(.dout(w_dff_A_2V4vMHZg3_0),.din(w_dff_A_jjFgBrHF1_0),.clk(gclk));
	jdff dff_A_2V4vMHZg3_0(.dout(w_dff_A_4NmUx1zy8_0),.din(w_dff_A_2V4vMHZg3_0),.clk(gclk));
	jdff dff_A_4NmUx1zy8_0(.dout(w_dff_A_f3UNqLF68_0),.din(w_dff_A_4NmUx1zy8_0),.clk(gclk));
	jdff dff_A_f3UNqLF68_0(.dout(w_dff_A_1TkdnhK27_0),.din(w_dff_A_f3UNqLF68_0),.clk(gclk));
	jdff dff_A_1TkdnhK27_0(.dout(w_dff_A_7mtasAMM5_0),.din(w_dff_A_1TkdnhK27_0),.clk(gclk));
	jdff dff_A_7mtasAMM5_0(.dout(w_dff_A_vuUWrtzl7_0),.din(w_dff_A_7mtasAMM5_0),.clk(gclk));
	jdff dff_A_vuUWrtzl7_0(.dout(w_dff_A_hvqVntsB3_0),.din(w_dff_A_vuUWrtzl7_0),.clk(gclk));
	jdff dff_A_hvqVntsB3_0(.dout(w_dff_A_xn4A3gjX9_0),.din(w_dff_A_hvqVntsB3_0),.clk(gclk));
	jdff dff_A_xn4A3gjX9_0(.dout(w_dff_A_LGA0xfO45_0),.din(w_dff_A_xn4A3gjX9_0),.clk(gclk));
	jdff dff_A_LGA0xfO45_0(.dout(w_dff_A_xl2lWlZv4_0),.din(w_dff_A_LGA0xfO45_0),.clk(gclk));
	jdff dff_A_xl2lWlZv4_0(.dout(w_dff_A_RyB0ER9j9_0),.din(w_dff_A_xl2lWlZv4_0),.clk(gclk));
	jdff dff_A_RyB0ER9j9_0(.dout(w_dff_A_GmkmoVbC6_0),.din(w_dff_A_RyB0ER9j9_0),.clk(gclk));
	jdff dff_A_GmkmoVbC6_0(.dout(w_dff_A_Lo3cqPBt5_0),.din(w_dff_A_GmkmoVbC6_0),.clk(gclk));
	jdff dff_A_Lo3cqPBt5_0(.dout(w_dff_A_lUViqljC5_0),.din(w_dff_A_Lo3cqPBt5_0),.clk(gclk));
	jdff dff_A_lUViqljC5_0(.dout(w_dff_A_ToIZSpra2_0),.din(w_dff_A_lUViqljC5_0),.clk(gclk));
	jdff dff_A_ToIZSpra2_0(.dout(w_dff_A_xgU7Kr8u0_0),.din(w_dff_A_ToIZSpra2_0),.clk(gclk));
	jdff dff_A_xgU7Kr8u0_0(.dout(w_dff_A_ma8E5OHg5_0),.din(w_dff_A_xgU7Kr8u0_0),.clk(gclk));
	jdff dff_A_ma8E5OHg5_0(.dout(w_dff_A_ga3vZeMV5_0),.din(w_dff_A_ma8E5OHg5_0),.clk(gclk));
	jdff dff_A_ga3vZeMV5_0(.dout(w_dff_A_or1Aq6e42_0),.din(w_dff_A_ga3vZeMV5_0),.clk(gclk));
	jdff dff_A_or1Aq6e42_0(.dout(w_dff_A_96S3lsn00_0),.din(w_dff_A_or1Aq6e42_0),.clk(gclk));
	jdff dff_A_96S3lsn00_0(.dout(w_dff_A_FVslTOr77_0),.din(w_dff_A_96S3lsn00_0),.clk(gclk));
	jdff dff_A_FVslTOr77_0(.dout(w_dff_A_xtPfsbII4_0),.din(w_dff_A_FVslTOr77_0),.clk(gclk));
	jdff dff_A_xtPfsbII4_0(.dout(w_dff_A_b5iJ6r5u9_0),.din(w_dff_A_xtPfsbII4_0),.clk(gclk));
	jdff dff_A_b5iJ6r5u9_0(.dout(w_dff_A_BaUTZo9B0_0),.din(w_dff_A_b5iJ6r5u9_0),.clk(gclk));
	jdff dff_A_BaUTZo9B0_0(.dout(w_dff_A_hy3GACAm2_0),.din(w_dff_A_BaUTZo9B0_0),.clk(gclk));
	jdff dff_A_hy3GACAm2_0(.dout(w_dff_A_qsYpd8yx8_0),.din(w_dff_A_hy3GACAm2_0),.clk(gclk));
	jdff dff_A_qsYpd8yx8_0(.dout(w_dff_A_lfpFRE3U9_0),.din(w_dff_A_qsYpd8yx8_0),.clk(gclk));
	jdff dff_A_lfpFRE3U9_0(.dout(w_dff_A_y67T9QrJ9_0),.din(w_dff_A_lfpFRE3U9_0),.clk(gclk));
	jdff dff_A_y67T9QrJ9_0(.dout(w_dff_A_iTEsgKpP0_0),.din(w_dff_A_y67T9QrJ9_0),.clk(gclk));
	jdff dff_A_iTEsgKpP0_0(.dout(w_dff_A_aNKI4mui0_0),.din(w_dff_A_iTEsgKpP0_0),.clk(gclk));
	jdff dff_A_aNKI4mui0_0(.dout(w_dff_A_3z6DXO5Y2_0),.din(w_dff_A_aNKI4mui0_0),.clk(gclk));
	jdff dff_A_3z6DXO5Y2_0(.dout(w_dff_A_8S6W1afs5_0),.din(w_dff_A_3z6DXO5Y2_0),.clk(gclk));
	jdff dff_A_8S6W1afs5_0(.dout(w_dff_A_InSWDsT87_0),.din(w_dff_A_8S6W1afs5_0),.clk(gclk));
	jdff dff_A_InSWDsT87_0(.dout(w_dff_A_Gw5uphno0_0),.din(w_dff_A_InSWDsT87_0),.clk(gclk));
	jdff dff_A_Gw5uphno0_0(.dout(w_dff_A_3eXJ7f2T9_0),.din(w_dff_A_Gw5uphno0_0),.clk(gclk));
	jdff dff_A_3eXJ7f2T9_0(.dout(w_dff_A_CcjBL7KS9_0),.din(w_dff_A_3eXJ7f2T9_0),.clk(gclk));
	jdff dff_A_CcjBL7KS9_0(.dout(w_dff_A_PQ2jiEph5_0),.din(w_dff_A_CcjBL7KS9_0),.clk(gclk));
	jdff dff_A_PQ2jiEph5_0(.dout(w_dff_A_4laSHGJN4_0),.din(w_dff_A_PQ2jiEph5_0),.clk(gclk));
	jdff dff_A_4laSHGJN4_0(.dout(f60),.din(w_dff_A_4laSHGJN4_0),.clk(gclk));
	jdff dff_A_cbJx3cUU7_2(.dout(w_dff_A_kN1bSLPi0_0),.din(w_dff_A_cbJx3cUU7_2),.clk(gclk));
	jdff dff_A_kN1bSLPi0_0(.dout(w_dff_A_pU53Tzbz8_0),.din(w_dff_A_kN1bSLPi0_0),.clk(gclk));
	jdff dff_A_pU53Tzbz8_0(.dout(w_dff_A_fHXVlomx4_0),.din(w_dff_A_pU53Tzbz8_0),.clk(gclk));
	jdff dff_A_fHXVlomx4_0(.dout(w_dff_A_9lMNg9097_0),.din(w_dff_A_fHXVlomx4_0),.clk(gclk));
	jdff dff_A_9lMNg9097_0(.dout(w_dff_A_r5qrXXzZ8_0),.din(w_dff_A_9lMNg9097_0),.clk(gclk));
	jdff dff_A_r5qrXXzZ8_0(.dout(w_dff_A_NNhvWYBd5_0),.din(w_dff_A_r5qrXXzZ8_0),.clk(gclk));
	jdff dff_A_NNhvWYBd5_0(.dout(w_dff_A_BW8ScAn92_0),.din(w_dff_A_NNhvWYBd5_0),.clk(gclk));
	jdff dff_A_BW8ScAn92_0(.dout(w_dff_A_H7YuW3Io4_0),.din(w_dff_A_BW8ScAn92_0),.clk(gclk));
	jdff dff_A_H7YuW3Io4_0(.dout(w_dff_A_jyqamt6N6_0),.din(w_dff_A_H7YuW3Io4_0),.clk(gclk));
	jdff dff_A_jyqamt6N6_0(.dout(w_dff_A_CklLsOyq2_0),.din(w_dff_A_jyqamt6N6_0),.clk(gclk));
	jdff dff_A_CklLsOyq2_0(.dout(w_dff_A_6CPpkvLh9_0),.din(w_dff_A_CklLsOyq2_0),.clk(gclk));
	jdff dff_A_6CPpkvLh9_0(.dout(w_dff_A_Wm95GZbe9_0),.din(w_dff_A_6CPpkvLh9_0),.clk(gclk));
	jdff dff_A_Wm95GZbe9_0(.dout(w_dff_A_OrJ1VE671_0),.din(w_dff_A_Wm95GZbe9_0),.clk(gclk));
	jdff dff_A_OrJ1VE671_0(.dout(w_dff_A_O0jiO9VO5_0),.din(w_dff_A_OrJ1VE671_0),.clk(gclk));
	jdff dff_A_O0jiO9VO5_0(.dout(w_dff_A_vDd1nOyy4_0),.din(w_dff_A_O0jiO9VO5_0),.clk(gclk));
	jdff dff_A_vDd1nOyy4_0(.dout(w_dff_A_mhtgDgWK5_0),.din(w_dff_A_vDd1nOyy4_0),.clk(gclk));
	jdff dff_A_mhtgDgWK5_0(.dout(w_dff_A_rPLaUmXr4_0),.din(w_dff_A_mhtgDgWK5_0),.clk(gclk));
	jdff dff_A_rPLaUmXr4_0(.dout(w_dff_A_Agwmk0Xn6_0),.din(w_dff_A_rPLaUmXr4_0),.clk(gclk));
	jdff dff_A_Agwmk0Xn6_0(.dout(w_dff_A_YFC8JQ6b7_0),.din(w_dff_A_Agwmk0Xn6_0),.clk(gclk));
	jdff dff_A_YFC8JQ6b7_0(.dout(w_dff_A_ihtAkP0y8_0),.din(w_dff_A_YFC8JQ6b7_0),.clk(gclk));
	jdff dff_A_ihtAkP0y8_0(.dout(w_dff_A_5BBIUexo6_0),.din(w_dff_A_ihtAkP0y8_0),.clk(gclk));
	jdff dff_A_5BBIUexo6_0(.dout(w_dff_A_zKqflDUK0_0),.din(w_dff_A_5BBIUexo6_0),.clk(gclk));
	jdff dff_A_zKqflDUK0_0(.dout(w_dff_A_D3kO9vDW6_0),.din(w_dff_A_zKqflDUK0_0),.clk(gclk));
	jdff dff_A_D3kO9vDW6_0(.dout(w_dff_A_MDB4X0DZ7_0),.din(w_dff_A_D3kO9vDW6_0),.clk(gclk));
	jdff dff_A_MDB4X0DZ7_0(.dout(w_dff_A_VKvh9Ose0_0),.din(w_dff_A_MDB4X0DZ7_0),.clk(gclk));
	jdff dff_A_VKvh9Ose0_0(.dout(w_dff_A_s4cSdd4I1_0),.din(w_dff_A_VKvh9Ose0_0),.clk(gclk));
	jdff dff_A_s4cSdd4I1_0(.dout(w_dff_A_nm3nGpql9_0),.din(w_dff_A_s4cSdd4I1_0),.clk(gclk));
	jdff dff_A_nm3nGpql9_0(.dout(w_dff_A_i93jo2NR1_0),.din(w_dff_A_nm3nGpql9_0),.clk(gclk));
	jdff dff_A_i93jo2NR1_0(.dout(w_dff_A_fM9oUSDX1_0),.din(w_dff_A_i93jo2NR1_0),.clk(gclk));
	jdff dff_A_fM9oUSDX1_0(.dout(w_dff_A_YzMm3uIC9_0),.din(w_dff_A_fM9oUSDX1_0),.clk(gclk));
	jdff dff_A_YzMm3uIC9_0(.dout(w_dff_A_JXKbEr9G1_0),.din(w_dff_A_YzMm3uIC9_0),.clk(gclk));
	jdff dff_A_JXKbEr9G1_0(.dout(w_dff_A_pSJFC5g39_0),.din(w_dff_A_JXKbEr9G1_0),.clk(gclk));
	jdff dff_A_pSJFC5g39_0(.dout(w_dff_A_D1zuIqrG5_0),.din(w_dff_A_pSJFC5g39_0),.clk(gclk));
	jdff dff_A_D1zuIqrG5_0(.dout(w_dff_A_xL28KK234_0),.din(w_dff_A_D1zuIqrG5_0),.clk(gclk));
	jdff dff_A_xL28KK234_0(.dout(w_dff_A_lvTNrHnY2_0),.din(w_dff_A_xL28KK234_0),.clk(gclk));
	jdff dff_A_lvTNrHnY2_0(.dout(w_dff_A_e1D8fWgY0_0),.din(w_dff_A_lvTNrHnY2_0),.clk(gclk));
	jdff dff_A_e1D8fWgY0_0(.dout(w_dff_A_3ac4XeuC1_0),.din(w_dff_A_e1D8fWgY0_0),.clk(gclk));
	jdff dff_A_3ac4XeuC1_0(.dout(w_dff_A_bKSR799b3_0),.din(w_dff_A_3ac4XeuC1_0),.clk(gclk));
	jdff dff_A_bKSR799b3_0(.dout(w_dff_A_PkaK4fsu9_0),.din(w_dff_A_bKSR799b3_0),.clk(gclk));
	jdff dff_A_PkaK4fsu9_0(.dout(w_dff_A_CD6IEukq8_0),.din(w_dff_A_PkaK4fsu9_0),.clk(gclk));
	jdff dff_A_CD6IEukq8_0(.dout(w_dff_A_IHOJ7yki6_0),.din(w_dff_A_CD6IEukq8_0),.clk(gclk));
	jdff dff_A_IHOJ7yki6_0(.dout(w_dff_A_vMFXKzEU7_0),.din(w_dff_A_IHOJ7yki6_0),.clk(gclk));
	jdff dff_A_vMFXKzEU7_0(.dout(w_dff_A_HPDvgGPZ5_0),.din(w_dff_A_vMFXKzEU7_0),.clk(gclk));
	jdff dff_A_HPDvgGPZ5_0(.dout(w_dff_A_NE76jVWk7_0),.din(w_dff_A_HPDvgGPZ5_0),.clk(gclk));
	jdff dff_A_NE76jVWk7_0(.dout(w_dff_A_huvqzPo59_0),.din(w_dff_A_NE76jVWk7_0),.clk(gclk));
	jdff dff_A_huvqzPo59_0(.dout(w_dff_A_WYyDuJiZ8_0),.din(w_dff_A_huvqzPo59_0),.clk(gclk));
	jdff dff_A_WYyDuJiZ8_0(.dout(w_dff_A_9SEdrZrT9_0),.din(w_dff_A_WYyDuJiZ8_0),.clk(gclk));
	jdff dff_A_9SEdrZrT9_0(.dout(w_dff_A_zUuFTNIx7_0),.din(w_dff_A_9SEdrZrT9_0),.clk(gclk));
	jdff dff_A_zUuFTNIx7_0(.dout(w_dff_A_IvIvHytR2_0),.din(w_dff_A_zUuFTNIx7_0),.clk(gclk));
	jdff dff_A_IvIvHytR2_0(.dout(w_dff_A_dqathm1m8_0),.din(w_dff_A_IvIvHytR2_0),.clk(gclk));
	jdff dff_A_dqathm1m8_0(.dout(w_dff_A_hKuATZ0h5_0),.din(w_dff_A_dqathm1m8_0),.clk(gclk));
	jdff dff_A_hKuATZ0h5_0(.dout(w_dff_A_TbdAxbTg1_0),.din(w_dff_A_hKuATZ0h5_0),.clk(gclk));
	jdff dff_A_TbdAxbTg1_0(.dout(w_dff_A_UafSs2yk8_0),.din(w_dff_A_TbdAxbTg1_0),.clk(gclk));
	jdff dff_A_UafSs2yk8_0(.dout(w_dff_A_xejBHwc88_0),.din(w_dff_A_UafSs2yk8_0),.clk(gclk));
	jdff dff_A_xejBHwc88_0(.dout(w_dff_A_npyi6nsg2_0),.din(w_dff_A_xejBHwc88_0),.clk(gclk));
	jdff dff_A_npyi6nsg2_0(.dout(w_dff_A_6HR8vrRl8_0),.din(w_dff_A_npyi6nsg2_0),.clk(gclk));
	jdff dff_A_6HR8vrRl8_0(.dout(w_dff_A_ObTwPOA53_0),.din(w_dff_A_6HR8vrRl8_0),.clk(gclk));
	jdff dff_A_ObTwPOA53_0(.dout(w_dff_A_Gd7G0SPF3_0),.din(w_dff_A_ObTwPOA53_0),.clk(gclk));
	jdff dff_A_Gd7G0SPF3_0(.dout(w_dff_A_p921a5Ff0_0),.din(w_dff_A_Gd7G0SPF3_0),.clk(gclk));
	jdff dff_A_p921a5Ff0_0(.dout(w_dff_A_FWzLRRfM1_0),.din(w_dff_A_p921a5Ff0_0),.clk(gclk));
	jdff dff_A_FWzLRRfM1_0(.dout(w_dff_A_7iw3XPmD2_0),.din(w_dff_A_FWzLRRfM1_0),.clk(gclk));
	jdff dff_A_7iw3XPmD2_0(.dout(w_dff_A_nMFdD3i91_0),.din(w_dff_A_7iw3XPmD2_0),.clk(gclk));
	jdff dff_A_nMFdD3i91_0(.dout(w_dff_A_KoRukcaO3_0),.din(w_dff_A_nMFdD3i91_0),.clk(gclk));
	jdff dff_A_KoRukcaO3_0(.dout(w_dff_A_78UlX4T87_0),.din(w_dff_A_KoRukcaO3_0),.clk(gclk));
	jdff dff_A_78UlX4T87_0(.dout(w_dff_A_XAZwDoNk6_0),.din(w_dff_A_78UlX4T87_0),.clk(gclk));
	jdff dff_A_XAZwDoNk6_0(.dout(f61),.din(w_dff_A_XAZwDoNk6_0),.clk(gclk));
	jdff dff_A_9pd4SMnz2_2(.dout(w_dff_A_9PfmIkxi1_0),.din(w_dff_A_9pd4SMnz2_2),.clk(gclk));
	jdff dff_A_9PfmIkxi1_0(.dout(w_dff_A_gnBGN4Av4_0),.din(w_dff_A_9PfmIkxi1_0),.clk(gclk));
	jdff dff_A_gnBGN4Av4_0(.dout(w_dff_A_tnAvPrj45_0),.din(w_dff_A_gnBGN4Av4_0),.clk(gclk));
	jdff dff_A_tnAvPrj45_0(.dout(w_dff_A_6frgHy4c3_0),.din(w_dff_A_tnAvPrj45_0),.clk(gclk));
	jdff dff_A_6frgHy4c3_0(.dout(w_dff_A_UC3MrkNQ4_0),.din(w_dff_A_6frgHy4c3_0),.clk(gclk));
	jdff dff_A_UC3MrkNQ4_0(.dout(w_dff_A_jwBoS0RU2_0),.din(w_dff_A_UC3MrkNQ4_0),.clk(gclk));
	jdff dff_A_jwBoS0RU2_0(.dout(w_dff_A_DAUUFlDO5_0),.din(w_dff_A_jwBoS0RU2_0),.clk(gclk));
	jdff dff_A_DAUUFlDO5_0(.dout(w_dff_A_D7LneTQU1_0),.din(w_dff_A_DAUUFlDO5_0),.clk(gclk));
	jdff dff_A_D7LneTQU1_0(.dout(w_dff_A_GZv5SRhw9_0),.din(w_dff_A_D7LneTQU1_0),.clk(gclk));
	jdff dff_A_GZv5SRhw9_0(.dout(w_dff_A_5ONaDWk54_0),.din(w_dff_A_GZv5SRhw9_0),.clk(gclk));
	jdff dff_A_5ONaDWk54_0(.dout(w_dff_A_y8c5hkjk6_0),.din(w_dff_A_5ONaDWk54_0),.clk(gclk));
	jdff dff_A_y8c5hkjk6_0(.dout(w_dff_A_DRixAHwj6_0),.din(w_dff_A_y8c5hkjk6_0),.clk(gclk));
	jdff dff_A_DRixAHwj6_0(.dout(w_dff_A_WmqDGt3E9_0),.din(w_dff_A_DRixAHwj6_0),.clk(gclk));
	jdff dff_A_WmqDGt3E9_0(.dout(w_dff_A_kjyaosTa3_0),.din(w_dff_A_WmqDGt3E9_0),.clk(gclk));
	jdff dff_A_kjyaosTa3_0(.dout(w_dff_A_FLcztQVR8_0),.din(w_dff_A_kjyaosTa3_0),.clk(gclk));
	jdff dff_A_FLcztQVR8_0(.dout(w_dff_A_o7EYSRrV1_0),.din(w_dff_A_FLcztQVR8_0),.clk(gclk));
	jdff dff_A_o7EYSRrV1_0(.dout(w_dff_A_k0BcLd351_0),.din(w_dff_A_o7EYSRrV1_0),.clk(gclk));
	jdff dff_A_k0BcLd351_0(.dout(w_dff_A_vAsdVf9t2_0),.din(w_dff_A_k0BcLd351_0),.clk(gclk));
	jdff dff_A_vAsdVf9t2_0(.dout(w_dff_A_Wpxldu1u5_0),.din(w_dff_A_vAsdVf9t2_0),.clk(gclk));
	jdff dff_A_Wpxldu1u5_0(.dout(w_dff_A_DsxfHCAe8_0),.din(w_dff_A_Wpxldu1u5_0),.clk(gclk));
	jdff dff_A_DsxfHCAe8_0(.dout(w_dff_A_A0VIBD6f3_0),.din(w_dff_A_DsxfHCAe8_0),.clk(gclk));
	jdff dff_A_A0VIBD6f3_0(.dout(w_dff_A_D9LoGEHc7_0),.din(w_dff_A_A0VIBD6f3_0),.clk(gclk));
	jdff dff_A_D9LoGEHc7_0(.dout(w_dff_A_3QJY9zSq4_0),.din(w_dff_A_D9LoGEHc7_0),.clk(gclk));
	jdff dff_A_3QJY9zSq4_0(.dout(w_dff_A_SHrOD7al1_0),.din(w_dff_A_3QJY9zSq4_0),.clk(gclk));
	jdff dff_A_SHrOD7al1_0(.dout(w_dff_A_KSJ6qf754_0),.din(w_dff_A_SHrOD7al1_0),.clk(gclk));
	jdff dff_A_KSJ6qf754_0(.dout(w_dff_A_9R7PCgSB1_0),.din(w_dff_A_KSJ6qf754_0),.clk(gclk));
	jdff dff_A_9R7PCgSB1_0(.dout(w_dff_A_cNqTuilG0_0),.din(w_dff_A_9R7PCgSB1_0),.clk(gclk));
	jdff dff_A_cNqTuilG0_0(.dout(w_dff_A_ueFnkmeT1_0),.din(w_dff_A_cNqTuilG0_0),.clk(gclk));
	jdff dff_A_ueFnkmeT1_0(.dout(w_dff_A_ItioFyrS9_0),.din(w_dff_A_ueFnkmeT1_0),.clk(gclk));
	jdff dff_A_ItioFyrS9_0(.dout(w_dff_A_ef6IySI54_0),.din(w_dff_A_ItioFyrS9_0),.clk(gclk));
	jdff dff_A_ef6IySI54_0(.dout(w_dff_A_S5c0VLsR1_0),.din(w_dff_A_ef6IySI54_0),.clk(gclk));
	jdff dff_A_S5c0VLsR1_0(.dout(w_dff_A_rkSGiJT10_0),.din(w_dff_A_S5c0VLsR1_0),.clk(gclk));
	jdff dff_A_rkSGiJT10_0(.dout(w_dff_A_Rk3Hp52T3_0),.din(w_dff_A_rkSGiJT10_0),.clk(gclk));
	jdff dff_A_Rk3Hp52T3_0(.dout(w_dff_A_GU2CYuYu2_0),.din(w_dff_A_Rk3Hp52T3_0),.clk(gclk));
	jdff dff_A_GU2CYuYu2_0(.dout(w_dff_A_pxNQ3lJG6_0),.din(w_dff_A_GU2CYuYu2_0),.clk(gclk));
	jdff dff_A_pxNQ3lJG6_0(.dout(w_dff_A_ACfNOD8U5_0),.din(w_dff_A_pxNQ3lJG6_0),.clk(gclk));
	jdff dff_A_ACfNOD8U5_0(.dout(w_dff_A_BP3jpmuq8_0),.din(w_dff_A_ACfNOD8U5_0),.clk(gclk));
	jdff dff_A_BP3jpmuq8_0(.dout(w_dff_A_o197X08U4_0),.din(w_dff_A_BP3jpmuq8_0),.clk(gclk));
	jdff dff_A_o197X08U4_0(.dout(w_dff_A_IRKI83st1_0),.din(w_dff_A_o197X08U4_0),.clk(gclk));
	jdff dff_A_IRKI83st1_0(.dout(w_dff_A_6FcKrCVq1_0),.din(w_dff_A_IRKI83st1_0),.clk(gclk));
	jdff dff_A_6FcKrCVq1_0(.dout(w_dff_A_hyPT4sqK1_0),.din(w_dff_A_6FcKrCVq1_0),.clk(gclk));
	jdff dff_A_hyPT4sqK1_0(.dout(w_dff_A_J4PWYUh44_0),.din(w_dff_A_hyPT4sqK1_0),.clk(gclk));
	jdff dff_A_J4PWYUh44_0(.dout(w_dff_A_QMvEQTq83_0),.din(w_dff_A_J4PWYUh44_0),.clk(gclk));
	jdff dff_A_QMvEQTq83_0(.dout(w_dff_A_3B312j3m4_0),.din(w_dff_A_QMvEQTq83_0),.clk(gclk));
	jdff dff_A_3B312j3m4_0(.dout(w_dff_A_ML8REE182_0),.din(w_dff_A_3B312j3m4_0),.clk(gclk));
	jdff dff_A_ML8REE182_0(.dout(w_dff_A_JNRb510u1_0),.din(w_dff_A_ML8REE182_0),.clk(gclk));
	jdff dff_A_JNRb510u1_0(.dout(w_dff_A_ffVbLAbd2_0),.din(w_dff_A_JNRb510u1_0),.clk(gclk));
	jdff dff_A_ffVbLAbd2_0(.dout(w_dff_A_1c3odY0u9_0),.din(w_dff_A_ffVbLAbd2_0),.clk(gclk));
	jdff dff_A_1c3odY0u9_0(.dout(w_dff_A_OS0Gssdy5_0),.din(w_dff_A_1c3odY0u9_0),.clk(gclk));
	jdff dff_A_OS0Gssdy5_0(.dout(w_dff_A_zAO9MmO81_0),.din(w_dff_A_OS0Gssdy5_0),.clk(gclk));
	jdff dff_A_zAO9MmO81_0(.dout(w_dff_A_pRkvoXdJ9_0),.din(w_dff_A_zAO9MmO81_0),.clk(gclk));
	jdff dff_A_pRkvoXdJ9_0(.dout(w_dff_A_Ft8LhTns2_0),.din(w_dff_A_pRkvoXdJ9_0),.clk(gclk));
	jdff dff_A_Ft8LhTns2_0(.dout(w_dff_A_oytcSXHT7_0),.din(w_dff_A_Ft8LhTns2_0),.clk(gclk));
	jdff dff_A_oytcSXHT7_0(.dout(w_dff_A_mTsLmeyk1_0),.din(w_dff_A_oytcSXHT7_0),.clk(gclk));
	jdff dff_A_mTsLmeyk1_0(.dout(w_dff_A_IeRSX9aG3_0),.din(w_dff_A_mTsLmeyk1_0),.clk(gclk));
	jdff dff_A_IeRSX9aG3_0(.dout(w_dff_A_flvMSnwk1_0),.din(w_dff_A_IeRSX9aG3_0),.clk(gclk));
	jdff dff_A_flvMSnwk1_0(.dout(w_dff_A_4o8JhBtq6_0),.din(w_dff_A_flvMSnwk1_0),.clk(gclk));
	jdff dff_A_4o8JhBtq6_0(.dout(w_dff_A_RLhGQEcn3_0),.din(w_dff_A_4o8JhBtq6_0),.clk(gclk));
	jdff dff_A_RLhGQEcn3_0(.dout(w_dff_A_00lUY1g44_0),.din(w_dff_A_RLhGQEcn3_0),.clk(gclk));
	jdff dff_A_00lUY1g44_0(.dout(w_dff_A_RAQDISZA9_0),.din(w_dff_A_00lUY1g44_0),.clk(gclk));
	jdff dff_A_RAQDISZA9_0(.dout(w_dff_A_dyfR1rfK6_0),.din(w_dff_A_RAQDISZA9_0),.clk(gclk));
	jdff dff_A_dyfR1rfK6_0(.dout(w_dff_A_mLvQVxo51_0),.din(w_dff_A_dyfR1rfK6_0),.clk(gclk));
	jdff dff_A_mLvQVxo51_0(.dout(w_dff_A_DvKJ7lzu8_0),.din(w_dff_A_mLvQVxo51_0),.clk(gclk));
	jdff dff_A_DvKJ7lzu8_0(.dout(w_dff_A_F60rCu3e1_0),.din(w_dff_A_DvKJ7lzu8_0),.clk(gclk));
	jdff dff_A_F60rCu3e1_0(.dout(f62),.din(w_dff_A_F60rCu3e1_0),.clk(gclk));
	jdff dff_A_was1nG0s4_2(.dout(w_dff_A_4FCaNSnF5_0),.din(w_dff_A_was1nG0s4_2),.clk(gclk));
	jdff dff_A_4FCaNSnF5_0(.dout(w_dff_A_sYQ3v8rF5_0),.din(w_dff_A_4FCaNSnF5_0),.clk(gclk));
	jdff dff_A_sYQ3v8rF5_0(.dout(w_dff_A_qcCGrghB4_0),.din(w_dff_A_sYQ3v8rF5_0),.clk(gclk));
	jdff dff_A_qcCGrghB4_0(.dout(w_dff_A_vqWtrOhV2_0),.din(w_dff_A_qcCGrghB4_0),.clk(gclk));
	jdff dff_A_vqWtrOhV2_0(.dout(w_dff_A_GaEtTw5l1_0),.din(w_dff_A_vqWtrOhV2_0),.clk(gclk));
	jdff dff_A_GaEtTw5l1_0(.dout(w_dff_A_nmfPLLqq2_0),.din(w_dff_A_GaEtTw5l1_0),.clk(gclk));
	jdff dff_A_nmfPLLqq2_0(.dout(w_dff_A_x4vz5G3h7_0),.din(w_dff_A_nmfPLLqq2_0),.clk(gclk));
	jdff dff_A_x4vz5G3h7_0(.dout(w_dff_A_XBV70oQG5_0),.din(w_dff_A_x4vz5G3h7_0),.clk(gclk));
	jdff dff_A_XBV70oQG5_0(.dout(w_dff_A_swgCIWAw8_0),.din(w_dff_A_XBV70oQG5_0),.clk(gclk));
	jdff dff_A_swgCIWAw8_0(.dout(w_dff_A_mqJpZsjQ7_0),.din(w_dff_A_swgCIWAw8_0),.clk(gclk));
	jdff dff_A_mqJpZsjQ7_0(.dout(w_dff_A_aqiF1x5N2_0),.din(w_dff_A_mqJpZsjQ7_0),.clk(gclk));
	jdff dff_A_aqiF1x5N2_0(.dout(w_dff_A_WyWQDoRG2_0),.din(w_dff_A_aqiF1x5N2_0),.clk(gclk));
	jdff dff_A_WyWQDoRG2_0(.dout(w_dff_A_lclP3gQt2_0),.din(w_dff_A_WyWQDoRG2_0),.clk(gclk));
	jdff dff_A_lclP3gQt2_0(.dout(w_dff_A_K44fYD4X4_0),.din(w_dff_A_lclP3gQt2_0),.clk(gclk));
	jdff dff_A_K44fYD4X4_0(.dout(w_dff_A_9NVRQDrT2_0),.din(w_dff_A_K44fYD4X4_0),.clk(gclk));
	jdff dff_A_9NVRQDrT2_0(.dout(w_dff_A_6eKjYWIg9_0),.din(w_dff_A_9NVRQDrT2_0),.clk(gclk));
	jdff dff_A_6eKjYWIg9_0(.dout(w_dff_A_fRvKaxiS3_0),.din(w_dff_A_6eKjYWIg9_0),.clk(gclk));
	jdff dff_A_fRvKaxiS3_0(.dout(w_dff_A_z7fDSSEg3_0),.din(w_dff_A_fRvKaxiS3_0),.clk(gclk));
	jdff dff_A_z7fDSSEg3_0(.dout(w_dff_A_02JCHMu74_0),.din(w_dff_A_z7fDSSEg3_0),.clk(gclk));
	jdff dff_A_02JCHMu74_0(.dout(w_dff_A_BZFTdOfS3_0),.din(w_dff_A_02JCHMu74_0),.clk(gclk));
	jdff dff_A_BZFTdOfS3_0(.dout(w_dff_A_cAvlbuaf4_0),.din(w_dff_A_BZFTdOfS3_0),.clk(gclk));
	jdff dff_A_cAvlbuaf4_0(.dout(w_dff_A_IzU5Us0H6_0),.din(w_dff_A_cAvlbuaf4_0),.clk(gclk));
	jdff dff_A_IzU5Us0H6_0(.dout(w_dff_A_ImNjsGOR8_0),.din(w_dff_A_IzU5Us0H6_0),.clk(gclk));
	jdff dff_A_ImNjsGOR8_0(.dout(w_dff_A_N7K6viDq1_0),.din(w_dff_A_ImNjsGOR8_0),.clk(gclk));
	jdff dff_A_N7K6viDq1_0(.dout(w_dff_A_zNqy6v5z2_0),.din(w_dff_A_N7K6viDq1_0),.clk(gclk));
	jdff dff_A_zNqy6v5z2_0(.dout(w_dff_A_cpJQcQWt8_0),.din(w_dff_A_zNqy6v5z2_0),.clk(gclk));
	jdff dff_A_cpJQcQWt8_0(.dout(w_dff_A_qtfGvc608_0),.din(w_dff_A_cpJQcQWt8_0),.clk(gclk));
	jdff dff_A_qtfGvc608_0(.dout(w_dff_A_Tsx8jgau7_0),.din(w_dff_A_qtfGvc608_0),.clk(gclk));
	jdff dff_A_Tsx8jgau7_0(.dout(w_dff_A_edBHmIUS6_0),.din(w_dff_A_Tsx8jgau7_0),.clk(gclk));
	jdff dff_A_edBHmIUS6_0(.dout(w_dff_A_BmyhuMAs1_0),.din(w_dff_A_edBHmIUS6_0),.clk(gclk));
	jdff dff_A_BmyhuMAs1_0(.dout(w_dff_A_Vq2RT1fi4_0),.din(w_dff_A_BmyhuMAs1_0),.clk(gclk));
	jdff dff_A_Vq2RT1fi4_0(.dout(w_dff_A_7yvtcHVA1_0),.din(w_dff_A_Vq2RT1fi4_0),.clk(gclk));
	jdff dff_A_7yvtcHVA1_0(.dout(w_dff_A_VIOSofcj5_0),.din(w_dff_A_7yvtcHVA1_0),.clk(gclk));
	jdff dff_A_VIOSofcj5_0(.dout(w_dff_A_SWBjya4A5_0),.din(w_dff_A_VIOSofcj5_0),.clk(gclk));
	jdff dff_A_SWBjya4A5_0(.dout(w_dff_A_dwoItiIv1_0),.din(w_dff_A_SWBjya4A5_0),.clk(gclk));
	jdff dff_A_dwoItiIv1_0(.dout(w_dff_A_VnNfcXQ54_0),.din(w_dff_A_dwoItiIv1_0),.clk(gclk));
	jdff dff_A_VnNfcXQ54_0(.dout(w_dff_A_mgEdXRmX7_0),.din(w_dff_A_VnNfcXQ54_0),.clk(gclk));
	jdff dff_A_mgEdXRmX7_0(.dout(w_dff_A_XMGpYcXb6_0),.din(w_dff_A_mgEdXRmX7_0),.clk(gclk));
	jdff dff_A_XMGpYcXb6_0(.dout(w_dff_A_eVRl7QfR7_0),.din(w_dff_A_XMGpYcXb6_0),.clk(gclk));
	jdff dff_A_eVRl7QfR7_0(.dout(w_dff_A_lz2spGC57_0),.din(w_dff_A_eVRl7QfR7_0),.clk(gclk));
	jdff dff_A_lz2spGC57_0(.dout(w_dff_A_Y7GSdF3e7_0),.din(w_dff_A_lz2spGC57_0),.clk(gclk));
	jdff dff_A_Y7GSdF3e7_0(.dout(w_dff_A_7A8A5mft1_0),.din(w_dff_A_Y7GSdF3e7_0),.clk(gclk));
	jdff dff_A_7A8A5mft1_0(.dout(w_dff_A_P69w1Sok6_0),.din(w_dff_A_7A8A5mft1_0),.clk(gclk));
	jdff dff_A_P69w1Sok6_0(.dout(w_dff_A_Yio3Fn8R3_0),.din(w_dff_A_P69w1Sok6_0),.clk(gclk));
	jdff dff_A_Yio3Fn8R3_0(.dout(w_dff_A_cy6FQlo22_0),.din(w_dff_A_Yio3Fn8R3_0),.clk(gclk));
	jdff dff_A_cy6FQlo22_0(.dout(w_dff_A_ZMOegiTE0_0),.din(w_dff_A_cy6FQlo22_0),.clk(gclk));
	jdff dff_A_ZMOegiTE0_0(.dout(w_dff_A_r8X4Wh9u7_0),.din(w_dff_A_ZMOegiTE0_0),.clk(gclk));
	jdff dff_A_r8X4Wh9u7_0(.dout(w_dff_A_AZVzxgdu0_0),.din(w_dff_A_r8X4Wh9u7_0),.clk(gclk));
	jdff dff_A_AZVzxgdu0_0(.dout(w_dff_A_2ummRGDO3_0),.din(w_dff_A_AZVzxgdu0_0),.clk(gclk));
	jdff dff_A_2ummRGDO3_0(.dout(w_dff_A_umWVonQZ5_0),.din(w_dff_A_2ummRGDO3_0),.clk(gclk));
	jdff dff_A_umWVonQZ5_0(.dout(w_dff_A_bXrxUx4F1_0),.din(w_dff_A_umWVonQZ5_0),.clk(gclk));
	jdff dff_A_bXrxUx4F1_0(.dout(w_dff_A_qP4DiCFE7_0),.din(w_dff_A_bXrxUx4F1_0),.clk(gclk));
	jdff dff_A_qP4DiCFE7_0(.dout(w_dff_A_rXVWxa8g6_0),.din(w_dff_A_qP4DiCFE7_0),.clk(gclk));
	jdff dff_A_rXVWxa8g6_0(.dout(w_dff_A_jSx6AQGo9_0),.din(w_dff_A_rXVWxa8g6_0),.clk(gclk));
	jdff dff_A_jSx6AQGo9_0(.dout(w_dff_A_4riuOLE45_0),.din(w_dff_A_jSx6AQGo9_0),.clk(gclk));
	jdff dff_A_4riuOLE45_0(.dout(w_dff_A_p9D2YWv37_0),.din(w_dff_A_4riuOLE45_0),.clk(gclk));
	jdff dff_A_p9D2YWv37_0(.dout(w_dff_A_wzPmPtWd8_0),.din(w_dff_A_p9D2YWv37_0),.clk(gclk));
	jdff dff_A_wzPmPtWd8_0(.dout(w_dff_A_MNTDk6jt7_0),.din(w_dff_A_wzPmPtWd8_0),.clk(gclk));
	jdff dff_A_MNTDk6jt7_0(.dout(w_dff_A_gCGFNWpA0_0),.din(w_dff_A_MNTDk6jt7_0),.clk(gclk));
	jdff dff_A_gCGFNWpA0_0(.dout(w_dff_A_VvXUNJJr1_0),.din(w_dff_A_gCGFNWpA0_0),.clk(gclk));
	jdff dff_A_VvXUNJJr1_0(.dout(w_dff_A_lwpUp4NK5_0),.din(w_dff_A_VvXUNJJr1_0),.clk(gclk));
	jdff dff_A_lwpUp4NK5_0(.dout(w_dff_A_2zudnWq70_0),.din(w_dff_A_lwpUp4NK5_0),.clk(gclk));
	jdff dff_A_2zudnWq70_0(.dout(w_dff_A_YGHgvoIb8_0),.din(w_dff_A_2zudnWq70_0),.clk(gclk));
	jdff dff_A_YGHgvoIb8_0(.dout(f63),.din(w_dff_A_YGHgvoIb8_0),.clk(gclk));
	jdff dff_A_fVeXfF3y3_2(.dout(w_dff_A_o1WbTIJ53_0),.din(w_dff_A_fVeXfF3y3_2),.clk(gclk));
	jdff dff_A_o1WbTIJ53_0(.dout(w_dff_A_4eEuNoo61_0),.din(w_dff_A_o1WbTIJ53_0),.clk(gclk));
	jdff dff_A_4eEuNoo61_0(.dout(w_dff_A_72v3frcJ4_0),.din(w_dff_A_4eEuNoo61_0),.clk(gclk));
	jdff dff_A_72v3frcJ4_0(.dout(w_dff_A_kZg1QiDS8_0),.din(w_dff_A_72v3frcJ4_0),.clk(gclk));
	jdff dff_A_kZg1QiDS8_0(.dout(w_dff_A_mednfuaS8_0),.din(w_dff_A_kZg1QiDS8_0),.clk(gclk));
	jdff dff_A_mednfuaS8_0(.dout(w_dff_A_sY1vGI651_0),.din(w_dff_A_mednfuaS8_0),.clk(gclk));
	jdff dff_A_sY1vGI651_0(.dout(w_dff_A_rJL7EMod6_0),.din(w_dff_A_sY1vGI651_0),.clk(gclk));
	jdff dff_A_rJL7EMod6_0(.dout(w_dff_A_5MfCJlFm8_0),.din(w_dff_A_rJL7EMod6_0),.clk(gclk));
	jdff dff_A_5MfCJlFm8_0(.dout(w_dff_A_8GWrTFld8_0),.din(w_dff_A_5MfCJlFm8_0),.clk(gclk));
	jdff dff_A_8GWrTFld8_0(.dout(w_dff_A_gpSTQkSQ4_0),.din(w_dff_A_8GWrTFld8_0),.clk(gclk));
	jdff dff_A_gpSTQkSQ4_0(.dout(w_dff_A_lSEFbcnH4_0),.din(w_dff_A_gpSTQkSQ4_0),.clk(gclk));
	jdff dff_A_lSEFbcnH4_0(.dout(w_dff_A_4SzqUtKF6_0),.din(w_dff_A_lSEFbcnH4_0),.clk(gclk));
	jdff dff_A_4SzqUtKF6_0(.dout(w_dff_A_ZI9dAyYC3_0),.din(w_dff_A_4SzqUtKF6_0),.clk(gclk));
	jdff dff_A_ZI9dAyYC3_0(.dout(w_dff_A_dAmQL6R87_0),.din(w_dff_A_ZI9dAyYC3_0),.clk(gclk));
	jdff dff_A_dAmQL6R87_0(.dout(w_dff_A_D2u1fAc26_0),.din(w_dff_A_dAmQL6R87_0),.clk(gclk));
	jdff dff_A_D2u1fAc26_0(.dout(w_dff_A_wYVFaF601_0),.din(w_dff_A_D2u1fAc26_0),.clk(gclk));
	jdff dff_A_wYVFaF601_0(.dout(w_dff_A_2fVY5uF90_0),.din(w_dff_A_wYVFaF601_0),.clk(gclk));
	jdff dff_A_2fVY5uF90_0(.dout(w_dff_A_d7CVs3OQ2_0),.din(w_dff_A_2fVY5uF90_0),.clk(gclk));
	jdff dff_A_d7CVs3OQ2_0(.dout(w_dff_A_Juhqcp5p3_0),.din(w_dff_A_d7CVs3OQ2_0),.clk(gclk));
	jdff dff_A_Juhqcp5p3_0(.dout(w_dff_A_jdno4zPP3_0),.din(w_dff_A_Juhqcp5p3_0),.clk(gclk));
	jdff dff_A_jdno4zPP3_0(.dout(w_dff_A_yeIoEjSc1_0),.din(w_dff_A_jdno4zPP3_0),.clk(gclk));
	jdff dff_A_yeIoEjSc1_0(.dout(w_dff_A_qf7H07IF0_0),.din(w_dff_A_yeIoEjSc1_0),.clk(gclk));
	jdff dff_A_qf7H07IF0_0(.dout(w_dff_A_eIEnfp250_0),.din(w_dff_A_qf7H07IF0_0),.clk(gclk));
	jdff dff_A_eIEnfp250_0(.dout(w_dff_A_pACpSUQN8_0),.din(w_dff_A_eIEnfp250_0),.clk(gclk));
	jdff dff_A_pACpSUQN8_0(.dout(w_dff_A_0k2YviDZ5_0),.din(w_dff_A_pACpSUQN8_0),.clk(gclk));
	jdff dff_A_0k2YviDZ5_0(.dout(w_dff_A_pZYcFIXx1_0),.din(w_dff_A_0k2YviDZ5_0),.clk(gclk));
	jdff dff_A_pZYcFIXx1_0(.dout(w_dff_A_yC5XCXIo3_0),.din(w_dff_A_pZYcFIXx1_0),.clk(gclk));
	jdff dff_A_yC5XCXIo3_0(.dout(w_dff_A_Oupxy7zq7_0),.din(w_dff_A_yC5XCXIo3_0),.clk(gclk));
	jdff dff_A_Oupxy7zq7_0(.dout(w_dff_A_zfJQipgK6_0),.din(w_dff_A_Oupxy7zq7_0),.clk(gclk));
	jdff dff_A_zfJQipgK6_0(.dout(w_dff_A_PjOAOSvb3_0),.din(w_dff_A_zfJQipgK6_0),.clk(gclk));
	jdff dff_A_PjOAOSvb3_0(.dout(w_dff_A_ZM5WpisM4_0),.din(w_dff_A_PjOAOSvb3_0),.clk(gclk));
	jdff dff_A_ZM5WpisM4_0(.dout(w_dff_A_38XLV76J4_0),.din(w_dff_A_ZM5WpisM4_0),.clk(gclk));
	jdff dff_A_38XLV76J4_0(.dout(w_dff_A_C0jI8AXB2_0),.din(w_dff_A_38XLV76J4_0),.clk(gclk));
	jdff dff_A_C0jI8AXB2_0(.dout(w_dff_A_85cmRc3R2_0),.din(w_dff_A_C0jI8AXB2_0),.clk(gclk));
	jdff dff_A_85cmRc3R2_0(.dout(w_dff_A_50UOJVWl2_0),.din(w_dff_A_85cmRc3R2_0),.clk(gclk));
	jdff dff_A_50UOJVWl2_0(.dout(w_dff_A_DLG9CSI75_0),.din(w_dff_A_50UOJVWl2_0),.clk(gclk));
	jdff dff_A_DLG9CSI75_0(.dout(w_dff_A_sV7XXod07_0),.din(w_dff_A_DLG9CSI75_0),.clk(gclk));
	jdff dff_A_sV7XXod07_0(.dout(w_dff_A_Ib9ubb7Y3_0),.din(w_dff_A_sV7XXod07_0),.clk(gclk));
	jdff dff_A_Ib9ubb7Y3_0(.dout(w_dff_A_z6Bo6U7Z8_0),.din(w_dff_A_Ib9ubb7Y3_0),.clk(gclk));
	jdff dff_A_z6Bo6U7Z8_0(.dout(w_dff_A_b2Zd016Q4_0),.din(w_dff_A_z6Bo6U7Z8_0),.clk(gclk));
	jdff dff_A_b2Zd016Q4_0(.dout(w_dff_A_fcRqM66B9_0),.din(w_dff_A_b2Zd016Q4_0),.clk(gclk));
	jdff dff_A_fcRqM66B9_0(.dout(w_dff_A_ermp00R91_0),.din(w_dff_A_fcRqM66B9_0),.clk(gclk));
	jdff dff_A_ermp00R91_0(.dout(w_dff_A_WUqcmPqk2_0),.din(w_dff_A_ermp00R91_0),.clk(gclk));
	jdff dff_A_WUqcmPqk2_0(.dout(w_dff_A_CwN7wier7_0),.din(w_dff_A_WUqcmPqk2_0),.clk(gclk));
	jdff dff_A_CwN7wier7_0(.dout(w_dff_A_c5Mig13r5_0),.din(w_dff_A_CwN7wier7_0),.clk(gclk));
	jdff dff_A_c5Mig13r5_0(.dout(w_dff_A_G76WnMkG0_0),.din(w_dff_A_c5Mig13r5_0),.clk(gclk));
	jdff dff_A_G76WnMkG0_0(.dout(w_dff_A_NJSYByyM6_0),.din(w_dff_A_G76WnMkG0_0),.clk(gclk));
	jdff dff_A_NJSYByyM6_0(.dout(w_dff_A_iFj29ikR8_0),.din(w_dff_A_NJSYByyM6_0),.clk(gclk));
	jdff dff_A_iFj29ikR8_0(.dout(w_dff_A_SYIDHwaH8_0),.din(w_dff_A_iFj29ikR8_0),.clk(gclk));
	jdff dff_A_SYIDHwaH8_0(.dout(w_dff_A_1CylodWj4_0),.din(w_dff_A_SYIDHwaH8_0),.clk(gclk));
	jdff dff_A_1CylodWj4_0(.dout(w_dff_A_zcawgL1s4_0),.din(w_dff_A_1CylodWj4_0),.clk(gclk));
	jdff dff_A_zcawgL1s4_0(.dout(w_dff_A_9NCRn5P10_0),.din(w_dff_A_zcawgL1s4_0),.clk(gclk));
	jdff dff_A_9NCRn5P10_0(.dout(w_dff_A_a0EdeibP0_0),.din(w_dff_A_9NCRn5P10_0),.clk(gclk));
	jdff dff_A_a0EdeibP0_0(.dout(w_dff_A_Nw1pbC711_0),.din(w_dff_A_a0EdeibP0_0),.clk(gclk));
	jdff dff_A_Nw1pbC711_0(.dout(w_dff_A_3Exa6QLI5_0),.din(w_dff_A_Nw1pbC711_0),.clk(gclk));
	jdff dff_A_3Exa6QLI5_0(.dout(w_dff_A_1Uup38GA0_0),.din(w_dff_A_3Exa6QLI5_0),.clk(gclk));
	jdff dff_A_1Uup38GA0_0(.dout(w_dff_A_e3Y5oSoZ5_0),.din(w_dff_A_1Uup38GA0_0),.clk(gclk));
	jdff dff_A_e3Y5oSoZ5_0(.dout(w_dff_A_C3SSud2Z7_0),.din(w_dff_A_e3Y5oSoZ5_0),.clk(gclk));
	jdff dff_A_C3SSud2Z7_0(.dout(w_dff_A_KgomdcfT8_0),.din(w_dff_A_C3SSud2Z7_0),.clk(gclk));
	jdff dff_A_KgomdcfT8_0(.dout(w_dff_A_67JOcsvH6_0),.din(w_dff_A_KgomdcfT8_0),.clk(gclk));
	jdff dff_A_67JOcsvH6_0(.dout(w_dff_A_cpxzsT6Z9_0),.din(w_dff_A_67JOcsvH6_0),.clk(gclk));
	jdff dff_A_cpxzsT6Z9_0(.dout(w_dff_A_wS98UYih4_0),.din(w_dff_A_cpxzsT6Z9_0),.clk(gclk));
	jdff dff_A_wS98UYih4_0(.dout(f64),.din(w_dff_A_wS98UYih4_0),.clk(gclk));
	jdff dff_A_apv54JrL0_2(.dout(w_dff_A_dBAk415Y4_0),.din(w_dff_A_apv54JrL0_2),.clk(gclk));
	jdff dff_A_dBAk415Y4_0(.dout(w_dff_A_laIz5X6W5_0),.din(w_dff_A_dBAk415Y4_0),.clk(gclk));
	jdff dff_A_laIz5X6W5_0(.dout(w_dff_A_IRpYVF7F6_0),.din(w_dff_A_laIz5X6W5_0),.clk(gclk));
	jdff dff_A_IRpYVF7F6_0(.dout(w_dff_A_RxKwzf739_0),.din(w_dff_A_IRpYVF7F6_0),.clk(gclk));
	jdff dff_A_RxKwzf739_0(.dout(w_dff_A_2S5r6X6P3_0),.din(w_dff_A_RxKwzf739_0),.clk(gclk));
	jdff dff_A_2S5r6X6P3_0(.dout(w_dff_A_3Us7mh066_0),.din(w_dff_A_2S5r6X6P3_0),.clk(gclk));
	jdff dff_A_3Us7mh066_0(.dout(w_dff_A_CvCHQFPK6_0),.din(w_dff_A_3Us7mh066_0),.clk(gclk));
	jdff dff_A_CvCHQFPK6_0(.dout(w_dff_A_zw0oIhC57_0),.din(w_dff_A_CvCHQFPK6_0),.clk(gclk));
	jdff dff_A_zw0oIhC57_0(.dout(w_dff_A_h2ZRzyZK2_0),.din(w_dff_A_zw0oIhC57_0),.clk(gclk));
	jdff dff_A_h2ZRzyZK2_0(.dout(w_dff_A_AJkqN9Z77_0),.din(w_dff_A_h2ZRzyZK2_0),.clk(gclk));
	jdff dff_A_AJkqN9Z77_0(.dout(w_dff_A_UW7QAg7Q5_0),.din(w_dff_A_AJkqN9Z77_0),.clk(gclk));
	jdff dff_A_UW7QAg7Q5_0(.dout(w_dff_A_jXKBgfSv4_0),.din(w_dff_A_UW7QAg7Q5_0),.clk(gclk));
	jdff dff_A_jXKBgfSv4_0(.dout(w_dff_A_7uW6PcDh4_0),.din(w_dff_A_jXKBgfSv4_0),.clk(gclk));
	jdff dff_A_7uW6PcDh4_0(.dout(w_dff_A_uNczXrg00_0),.din(w_dff_A_7uW6PcDh4_0),.clk(gclk));
	jdff dff_A_uNczXrg00_0(.dout(w_dff_A_WmkES23T9_0),.din(w_dff_A_uNczXrg00_0),.clk(gclk));
	jdff dff_A_WmkES23T9_0(.dout(w_dff_A_TCzmEIA36_0),.din(w_dff_A_WmkES23T9_0),.clk(gclk));
	jdff dff_A_TCzmEIA36_0(.dout(w_dff_A_wyR3Q9Rc4_0),.din(w_dff_A_TCzmEIA36_0),.clk(gclk));
	jdff dff_A_wyR3Q9Rc4_0(.dout(w_dff_A_b6xjJOkB0_0),.din(w_dff_A_wyR3Q9Rc4_0),.clk(gclk));
	jdff dff_A_b6xjJOkB0_0(.dout(w_dff_A_Ayg9xbJf4_0),.din(w_dff_A_b6xjJOkB0_0),.clk(gclk));
	jdff dff_A_Ayg9xbJf4_0(.dout(w_dff_A_0dCwa6hS4_0),.din(w_dff_A_Ayg9xbJf4_0),.clk(gclk));
	jdff dff_A_0dCwa6hS4_0(.dout(w_dff_A_9C0bhD3t7_0),.din(w_dff_A_0dCwa6hS4_0),.clk(gclk));
	jdff dff_A_9C0bhD3t7_0(.dout(w_dff_A_xUTFGiiT1_0),.din(w_dff_A_9C0bhD3t7_0),.clk(gclk));
	jdff dff_A_xUTFGiiT1_0(.dout(w_dff_A_ytRNEqYc2_0),.din(w_dff_A_xUTFGiiT1_0),.clk(gclk));
	jdff dff_A_ytRNEqYc2_0(.dout(w_dff_A_04owxQqU3_0),.din(w_dff_A_ytRNEqYc2_0),.clk(gclk));
	jdff dff_A_04owxQqU3_0(.dout(w_dff_A_nN3yAUis8_0),.din(w_dff_A_04owxQqU3_0),.clk(gclk));
	jdff dff_A_nN3yAUis8_0(.dout(w_dff_A_0mEhRKRq8_0),.din(w_dff_A_nN3yAUis8_0),.clk(gclk));
	jdff dff_A_0mEhRKRq8_0(.dout(w_dff_A_MTpXKLcC3_0),.din(w_dff_A_0mEhRKRq8_0),.clk(gclk));
	jdff dff_A_MTpXKLcC3_0(.dout(w_dff_A_Ydmwoqxb1_0),.din(w_dff_A_MTpXKLcC3_0),.clk(gclk));
	jdff dff_A_Ydmwoqxb1_0(.dout(w_dff_A_v40fqtLM3_0),.din(w_dff_A_Ydmwoqxb1_0),.clk(gclk));
	jdff dff_A_v40fqtLM3_0(.dout(w_dff_A_CVsD3srr9_0),.din(w_dff_A_v40fqtLM3_0),.clk(gclk));
	jdff dff_A_CVsD3srr9_0(.dout(w_dff_A_i8WMIx4R4_0),.din(w_dff_A_CVsD3srr9_0),.clk(gclk));
	jdff dff_A_i8WMIx4R4_0(.dout(w_dff_A_7AXU1di97_0),.din(w_dff_A_i8WMIx4R4_0),.clk(gclk));
	jdff dff_A_7AXU1di97_0(.dout(w_dff_A_3MNZvNFh3_0),.din(w_dff_A_7AXU1di97_0),.clk(gclk));
	jdff dff_A_3MNZvNFh3_0(.dout(w_dff_A_CObArfJD6_0),.din(w_dff_A_3MNZvNFh3_0),.clk(gclk));
	jdff dff_A_CObArfJD6_0(.dout(w_dff_A_Hi4dpTD43_0),.din(w_dff_A_CObArfJD6_0),.clk(gclk));
	jdff dff_A_Hi4dpTD43_0(.dout(w_dff_A_Tr95Q3F94_0),.din(w_dff_A_Hi4dpTD43_0),.clk(gclk));
	jdff dff_A_Tr95Q3F94_0(.dout(w_dff_A_o17VLYLF1_0),.din(w_dff_A_Tr95Q3F94_0),.clk(gclk));
	jdff dff_A_o17VLYLF1_0(.dout(w_dff_A_CjEBfkaa9_0),.din(w_dff_A_o17VLYLF1_0),.clk(gclk));
	jdff dff_A_CjEBfkaa9_0(.dout(w_dff_A_JUnIpInf4_0),.din(w_dff_A_CjEBfkaa9_0),.clk(gclk));
	jdff dff_A_JUnIpInf4_0(.dout(w_dff_A_YF1KtEL77_0),.din(w_dff_A_JUnIpInf4_0),.clk(gclk));
	jdff dff_A_YF1KtEL77_0(.dout(w_dff_A_URGOLNDV3_0),.din(w_dff_A_YF1KtEL77_0),.clk(gclk));
	jdff dff_A_URGOLNDV3_0(.dout(w_dff_A_MMghgGcf7_0),.din(w_dff_A_URGOLNDV3_0),.clk(gclk));
	jdff dff_A_MMghgGcf7_0(.dout(w_dff_A_di2VmveN6_0),.din(w_dff_A_MMghgGcf7_0),.clk(gclk));
	jdff dff_A_di2VmveN6_0(.dout(w_dff_A_AFgb8HMT2_0),.din(w_dff_A_di2VmveN6_0),.clk(gclk));
	jdff dff_A_AFgb8HMT2_0(.dout(w_dff_A_yIC4WPEG8_0),.din(w_dff_A_AFgb8HMT2_0),.clk(gclk));
	jdff dff_A_yIC4WPEG8_0(.dout(w_dff_A_yNyn99U82_0),.din(w_dff_A_yIC4WPEG8_0),.clk(gclk));
	jdff dff_A_yNyn99U82_0(.dout(w_dff_A_0dWn8Spw9_0),.din(w_dff_A_yNyn99U82_0),.clk(gclk));
	jdff dff_A_0dWn8Spw9_0(.dout(w_dff_A_FPxhwbtW1_0),.din(w_dff_A_0dWn8Spw9_0),.clk(gclk));
	jdff dff_A_FPxhwbtW1_0(.dout(w_dff_A_qatcRyM88_0),.din(w_dff_A_FPxhwbtW1_0),.clk(gclk));
	jdff dff_A_qatcRyM88_0(.dout(w_dff_A_F043k6ju5_0),.din(w_dff_A_qatcRyM88_0),.clk(gclk));
	jdff dff_A_F043k6ju5_0(.dout(w_dff_A_rJWNtSpD6_0),.din(w_dff_A_F043k6ju5_0),.clk(gclk));
	jdff dff_A_rJWNtSpD6_0(.dout(w_dff_A_uZNWG3zu3_0),.din(w_dff_A_rJWNtSpD6_0),.clk(gclk));
	jdff dff_A_uZNWG3zu3_0(.dout(w_dff_A_1DIb0yIg8_0),.din(w_dff_A_uZNWG3zu3_0),.clk(gclk));
	jdff dff_A_1DIb0yIg8_0(.dout(w_dff_A_ZPEldzRF0_0),.din(w_dff_A_1DIb0yIg8_0),.clk(gclk));
	jdff dff_A_ZPEldzRF0_0(.dout(w_dff_A_bEHjzTA55_0),.din(w_dff_A_ZPEldzRF0_0),.clk(gclk));
	jdff dff_A_bEHjzTA55_0(.dout(w_dff_A_BrBKtJlW8_0),.din(w_dff_A_bEHjzTA55_0),.clk(gclk));
	jdff dff_A_BrBKtJlW8_0(.dout(w_dff_A_fDLHVQoQ9_0),.din(w_dff_A_BrBKtJlW8_0),.clk(gclk));
	jdff dff_A_fDLHVQoQ9_0(.dout(w_dff_A_S3Nt75zP6_0),.din(w_dff_A_fDLHVQoQ9_0),.clk(gclk));
	jdff dff_A_S3Nt75zP6_0(.dout(w_dff_A_xsOYTMRG8_0),.din(w_dff_A_S3Nt75zP6_0),.clk(gclk));
	jdff dff_A_xsOYTMRG8_0(.dout(w_dff_A_YUpDGpAj9_0),.din(w_dff_A_xsOYTMRG8_0),.clk(gclk));
	jdff dff_A_YUpDGpAj9_0(.dout(w_dff_A_W18ZItLa2_0),.din(w_dff_A_YUpDGpAj9_0),.clk(gclk));
	jdff dff_A_W18ZItLa2_0(.dout(f65),.din(w_dff_A_W18ZItLa2_0),.clk(gclk));
	jdff dff_A_u9JR45Q39_2(.dout(w_dff_A_a7kPmvzC1_0),.din(w_dff_A_u9JR45Q39_2),.clk(gclk));
	jdff dff_A_a7kPmvzC1_0(.dout(w_dff_A_7FNMHEa77_0),.din(w_dff_A_a7kPmvzC1_0),.clk(gclk));
	jdff dff_A_7FNMHEa77_0(.dout(w_dff_A_Qwgnt3vg5_0),.din(w_dff_A_7FNMHEa77_0),.clk(gclk));
	jdff dff_A_Qwgnt3vg5_0(.dout(w_dff_A_p3SR5rm08_0),.din(w_dff_A_Qwgnt3vg5_0),.clk(gclk));
	jdff dff_A_p3SR5rm08_0(.dout(w_dff_A_bAfZdBgC4_0),.din(w_dff_A_p3SR5rm08_0),.clk(gclk));
	jdff dff_A_bAfZdBgC4_0(.dout(w_dff_A_ZcmVLl2Z3_0),.din(w_dff_A_bAfZdBgC4_0),.clk(gclk));
	jdff dff_A_ZcmVLl2Z3_0(.dout(w_dff_A_GXhe9woH1_0),.din(w_dff_A_ZcmVLl2Z3_0),.clk(gclk));
	jdff dff_A_GXhe9woH1_0(.dout(w_dff_A_iZykjJyM7_0),.din(w_dff_A_GXhe9woH1_0),.clk(gclk));
	jdff dff_A_iZykjJyM7_0(.dout(w_dff_A_16kHkLPy9_0),.din(w_dff_A_iZykjJyM7_0),.clk(gclk));
	jdff dff_A_16kHkLPy9_0(.dout(w_dff_A_saj9RMhn5_0),.din(w_dff_A_16kHkLPy9_0),.clk(gclk));
	jdff dff_A_saj9RMhn5_0(.dout(w_dff_A_Y3xeWqjd5_0),.din(w_dff_A_saj9RMhn5_0),.clk(gclk));
	jdff dff_A_Y3xeWqjd5_0(.dout(w_dff_A_oXRebKbp3_0),.din(w_dff_A_Y3xeWqjd5_0),.clk(gclk));
	jdff dff_A_oXRebKbp3_0(.dout(w_dff_A_4aQmSl5r0_0),.din(w_dff_A_oXRebKbp3_0),.clk(gclk));
	jdff dff_A_4aQmSl5r0_0(.dout(w_dff_A_IGXyLNWA5_0),.din(w_dff_A_4aQmSl5r0_0),.clk(gclk));
	jdff dff_A_IGXyLNWA5_0(.dout(w_dff_A_i3ZYYbKD0_0),.din(w_dff_A_IGXyLNWA5_0),.clk(gclk));
	jdff dff_A_i3ZYYbKD0_0(.dout(w_dff_A_PT6v9qWd7_0),.din(w_dff_A_i3ZYYbKD0_0),.clk(gclk));
	jdff dff_A_PT6v9qWd7_0(.dout(w_dff_A_1JHiii4c8_0),.din(w_dff_A_PT6v9qWd7_0),.clk(gclk));
	jdff dff_A_1JHiii4c8_0(.dout(w_dff_A_DVPtnxHP0_0),.din(w_dff_A_1JHiii4c8_0),.clk(gclk));
	jdff dff_A_DVPtnxHP0_0(.dout(w_dff_A_gUQf8DSC8_0),.din(w_dff_A_DVPtnxHP0_0),.clk(gclk));
	jdff dff_A_gUQf8DSC8_0(.dout(w_dff_A_0Mnqp26m1_0),.din(w_dff_A_gUQf8DSC8_0),.clk(gclk));
	jdff dff_A_0Mnqp26m1_0(.dout(w_dff_A_rlTXzyAW9_0),.din(w_dff_A_0Mnqp26m1_0),.clk(gclk));
	jdff dff_A_rlTXzyAW9_0(.dout(w_dff_A_QfBEi23Q6_0),.din(w_dff_A_rlTXzyAW9_0),.clk(gclk));
	jdff dff_A_QfBEi23Q6_0(.dout(w_dff_A_mDtT5sAP9_0),.din(w_dff_A_QfBEi23Q6_0),.clk(gclk));
	jdff dff_A_mDtT5sAP9_0(.dout(w_dff_A_9w8IdPq26_0),.din(w_dff_A_mDtT5sAP9_0),.clk(gclk));
	jdff dff_A_9w8IdPq26_0(.dout(w_dff_A_fhqoxttH0_0),.din(w_dff_A_9w8IdPq26_0),.clk(gclk));
	jdff dff_A_fhqoxttH0_0(.dout(w_dff_A_d0Uepe1X4_0),.din(w_dff_A_fhqoxttH0_0),.clk(gclk));
	jdff dff_A_d0Uepe1X4_0(.dout(w_dff_A_WCzqahEH2_0),.din(w_dff_A_d0Uepe1X4_0),.clk(gclk));
	jdff dff_A_WCzqahEH2_0(.dout(w_dff_A_uV48ueqp1_0),.din(w_dff_A_WCzqahEH2_0),.clk(gclk));
	jdff dff_A_uV48ueqp1_0(.dout(w_dff_A_OESZUosL8_0),.din(w_dff_A_uV48ueqp1_0),.clk(gclk));
	jdff dff_A_OESZUosL8_0(.dout(w_dff_A_FKwp4Rvw4_0),.din(w_dff_A_OESZUosL8_0),.clk(gclk));
	jdff dff_A_FKwp4Rvw4_0(.dout(w_dff_A_4S07OXcP6_0),.din(w_dff_A_FKwp4Rvw4_0),.clk(gclk));
	jdff dff_A_4S07OXcP6_0(.dout(w_dff_A_GinmoGLY6_0),.din(w_dff_A_4S07OXcP6_0),.clk(gclk));
	jdff dff_A_GinmoGLY6_0(.dout(w_dff_A_9JNqIL4L4_0),.din(w_dff_A_GinmoGLY6_0),.clk(gclk));
	jdff dff_A_9JNqIL4L4_0(.dout(w_dff_A_wtsJNKpU2_0),.din(w_dff_A_9JNqIL4L4_0),.clk(gclk));
	jdff dff_A_wtsJNKpU2_0(.dout(w_dff_A_F1ZE7YzQ0_0),.din(w_dff_A_wtsJNKpU2_0),.clk(gclk));
	jdff dff_A_F1ZE7YzQ0_0(.dout(w_dff_A_mDd66k3u4_0),.din(w_dff_A_F1ZE7YzQ0_0),.clk(gclk));
	jdff dff_A_mDd66k3u4_0(.dout(w_dff_A_Qt2fUqli2_0),.din(w_dff_A_mDd66k3u4_0),.clk(gclk));
	jdff dff_A_Qt2fUqli2_0(.dout(w_dff_A_MnWZZulQ5_0),.din(w_dff_A_Qt2fUqli2_0),.clk(gclk));
	jdff dff_A_MnWZZulQ5_0(.dout(w_dff_A_ZUUa9zWM5_0),.din(w_dff_A_MnWZZulQ5_0),.clk(gclk));
	jdff dff_A_ZUUa9zWM5_0(.dout(w_dff_A_5TU1mqak4_0),.din(w_dff_A_ZUUa9zWM5_0),.clk(gclk));
	jdff dff_A_5TU1mqak4_0(.dout(w_dff_A_gDAlXsIW5_0),.din(w_dff_A_5TU1mqak4_0),.clk(gclk));
	jdff dff_A_gDAlXsIW5_0(.dout(w_dff_A_Ht03QWsm3_0),.din(w_dff_A_gDAlXsIW5_0),.clk(gclk));
	jdff dff_A_Ht03QWsm3_0(.dout(w_dff_A_DEwoiM0B5_0),.din(w_dff_A_Ht03QWsm3_0),.clk(gclk));
	jdff dff_A_DEwoiM0B5_0(.dout(w_dff_A_HnCVEyRa4_0),.din(w_dff_A_DEwoiM0B5_0),.clk(gclk));
	jdff dff_A_HnCVEyRa4_0(.dout(w_dff_A_6ACEfJDP4_0),.din(w_dff_A_HnCVEyRa4_0),.clk(gclk));
	jdff dff_A_6ACEfJDP4_0(.dout(w_dff_A_6DQffS4r7_0),.din(w_dff_A_6ACEfJDP4_0),.clk(gclk));
	jdff dff_A_6DQffS4r7_0(.dout(w_dff_A_rX2JkSeX4_0),.din(w_dff_A_6DQffS4r7_0),.clk(gclk));
	jdff dff_A_rX2JkSeX4_0(.dout(w_dff_A_TMJkF1bT0_0),.din(w_dff_A_rX2JkSeX4_0),.clk(gclk));
	jdff dff_A_TMJkF1bT0_0(.dout(w_dff_A_epTUJaUk7_0),.din(w_dff_A_TMJkF1bT0_0),.clk(gclk));
	jdff dff_A_epTUJaUk7_0(.dout(w_dff_A_vLvb4JyL5_0),.din(w_dff_A_epTUJaUk7_0),.clk(gclk));
	jdff dff_A_vLvb4JyL5_0(.dout(w_dff_A_1QrB1juE3_0),.din(w_dff_A_vLvb4JyL5_0),.clk(gclk));
	jdff dff_A_1QrB1juE3_0(.dout(w_dff_A_NSQRscGH1_0),.din(w_dff_A_1QrB1juE3_0),.clk(gclk));
	jdff dff_A_NSQRscGH1_0(.dout(w_dff_A_zutMZV7w2_0),.din(w_dff_A_NSQRscGH1_0),.clk(gclk));
	jdff dff_A_zutMZV7w2_0(.dout(w_dff_A_xqok4ro61_0),.din(w_dff_A_zutMZV7w2_0),.clk(gclk));
	jdff dff_A_xqok4ro61_0(.dout(w_dff_A_wQidtS463_0),.din(w_dff_A_xqok4ro61_0),.clk(gclk));
	jdff dff_A_wQidtS463_0(.dout(w_dff_A_2ldpwheP1_0),.din(w_dff_A_wQidtS463_0),.clk(gclk));
	jdff dff_A_2ldpwheP1_0(.dout(w_dff_A_DzL73d7t1_0),.din(w_dff_A_2ldpwheP1_0),.clk(gclk));
	jdff dff_A_DzL73d7t1_0(.dout(w_dff_A_aayfAdcH5_0),.din(w_dff_A_DzL73d7t1_0),.clk(gclk));
	jdff dff_A_aayfAdcH5_0(.dout(w_dff_A_d3nXRxgJ1_0),.din(w_dff_A_aayfAdcH5_0),.clk(gclk));
	jdff dff_A_d3nXRxgJ1_0(.dout(w_dff_A_9ozywqgS9_0),.din(w_dff_A_d3nXRxgJ1_0),.clk(gclk));
	jdff dff_A_9ozywqgS9_0(.dout(f66),.din(w_dff_A_9ozywqgS9_0),.clk(gclk));
	jdff dff_A_Z4pRlS9P8_2(.dout(w_dff_A_T6Ac4q6P4_0),.din(w_dff_A_Z4pRlS9P8_2),.clk(gclk));
	jdff dff_A_T6Ac4q6P4_0(.dout(w_dff_A_e7T8cfxq1_0),.din(w_dff_A_T6Ac4q6P4_0),.clk(gclk));
	jdff dff_A_e7T8cfxq1_0(.dout(w_dff_A_IrLFQIPX6_0),.din(w_dff_A_e7T8cfxq1_0),.clk(gclk));
	jdff dff_A_IrLFQIPX6_0(.dout(w_dff_A_A4JRQDsT1_0),.din(w_dff_A_IrLFQIPX6_0),.clk(gclk));
	jdff dff_A_A4JRQDsT1_0(.dout(w_dff_A_VZFsfBxM0_0),.din(w_dff_A_A4JRQDsT1_0),.clk(gclk));
	jdff dff_A_VZFsfBxM0_0(.dout(w_dff_A_6lua5B5g5_0),.din(w_dff_A_VZFsfBxM0_0),.clk(gclk));
	jdff dff_A_6lua5B5g5_0(.dout(w_dff_A_ql2yu8Hy8_0),.din(w_dff_A_6lua5B5g5_0),.clk(gclk));
	jdff dff_A_ql2yu8Hy8_0(.dout(w_dff_A_bhHMrDYy8_0),.din(w_dff_A_ql2yu8Hy8_0),.clk(gclk));
	jdff dff_A_bhHMrDYy8_0(.dout(w_dff_A_T3eqOZBl7_0),.din(w_dff_A_bhHMrDYy8_0),.clk(gclk));
	jdff dff_A_T3eqOZBl7_0(.dout(w_dff_A_hH2QfJjq6_0),.din(w_dff_A_T3eqOZBl7_0),.clk(gclk));
	jdff dff_A_hH2QfJjq6_0(.dout(w_dff_A_9NDLG0688_0),.din(w_dff_A_hH2QfJjq6_0),.clk(gclk));
	jdff dff_A_9NDLG0688_0(.dout(w_dff_A_nl88IL6c8_0),.din(w_dff_A_9NDLG0688_0),.clk(gclk));
	jdff dff_A_nl88IL6c8_0(.dout(w_dff_A_HxzuLJOW6_0),.din(w_dff_A_nl88IL6c8_0),.clk(gclk));
	jdff dff_A_HxzuLJOW6_0(.dout(w_dff_A_yeY0su3y6_0),.din(w_dff_A_HxzuLJOW6_0),.clk(gclk));
	jdff dff_A_yeY0su3y6_0(.dout(w_dff_A_8oeH0eZr5_0),.din(w_dff_A_yeY0su3y6_0),.clk(gclk));
	jdff dff_A_8oeH0eZr5_0(.dout(w_dff_A_8qJNKg2A8_0),.din(w_dff_A_8oeH0eZr5_0),.clk(gclk));
	jdff dff_A_8qJNKg2A8_0(.dout(w_dff_A_JihLZUbE8_0),.din(w_dff_A_8qJNKg2A8_0),.clk(gclk));
	jdff dff_A_JihLZUbE8_0(.dout(w_dff_A_SBqhS0Rm0_0),.din(w_dff_A_JihLZUbE8_0),.clk(gclk));
	jdff dff_A_SBqhS0Rm0_0(.dout(w_dff_A_CmpFw6cr6_0),.din(w_dff_A_SBqhS0Rm0_0),.clk(gclk));
	jdff dff_A_CmpFw6cr6_0(.dout(w_dff_A_OKZJTjQH0_0),.din(w_dff_A_CmpFw6cr6_0),.clk(gclk));
	jdff dff_A_OKZJTjQH0_0(.dout(w_dff_A_OsKbSxXn3_0),.din(w_dff_A_OKZJTjQH0_0),.clk(gclk));
	jdff dff_A_OsKbSxXn3_0(.dout(w_dff_A_fdp4NZXr5_0),.din(w_dff_A_OsKbSxXn3_0),.clk(gclk));
	jdff dff_A_fdp4NZXr5_0(.dout(w_dff_A_3EEOslsn8_0),.din(w_dff_A_fdp4NZXr5_0),.clk(gclk));
	jdff dff_A_3EEOslsn8_0(.dout(w_dff_A_fAtbWiGN6_0),.din(w_dff_A_3EEOslsn8_0),.clk(gclk));
	jdff dff_A_fAtbWiGN6_0(.dout(w_dff_A_gCvvaal76_0),.din(w_dff_A_fAtbWiGN6_0),.clk(gclk));
	jdff dff_A_gCvvaal76_0(.dout(w_dff_A_gnFjCrWj2_0),.din(w_dff_A_gCvvaal76_0),.clk(gclk));
	jdff dff_A_gnFjCrWj2_0(.dout(w_dff_A_pnErWyHg1_0),.din(w_dff_A_gnFjCrWj2_0),.clk(gclk));
	jdff dff_A_pnErWyHg1_0(.dout(w_dff_A_8B1TxZJ64_0),.din(w_dff_A_pnErWyHg1_0),.clk(gclk));
	jdff dff_A_8B1TxZJ64_0(.dout(w_dff_A_hOBxosRT4_0),.din(w_dff_A_8B1TxZJ64_0),.clk(gclk));
	jdff dff_A_hOBxosRT4_0(.dout(w_dff_A_wZB0b1xB6_0),.din(w_dff_A_hOBxosRT4_0),.clk(gclk));
	jdff dff_A_wZB0b1xB6_0(.dout(w_dff_A_nXNxlDSO0_0),.din(w_dff_A_wZB0b1xB6_0),.clk(gclk));
	jdff dff_A_nXNxlDSO0_0(.dout(w_dff_A_5U1Qd4AU7_0),.din(w_dff_A_nXNxlDSO0_0),.clk(gclk));
	jdff dff_A_5U1Qd4AU7_0(.dout(w_dff_A_pRm0Pu0r9_0),.din(w_dff_A_5U1Qd4AU7_0),.clk(gclk));
	jdff dff_A_pRm0Pu0r9_0(.dout(w_dff_A_Rq4vNT679_0),.din(w_dff_A_pRm0Pu0r9_0),.clk(gclk));
	jdff dff_A_Rq4vNT679_0(.dout(w_dff_A_odVIc5ZV1_0),.din(w_dff_A_Rq4vNT679_0),.clk(gclk));
	jdff dff_A_odVIc5ZV1_0(.dout(w_dff_A_7BoI3UZc9_0),.din(w_dff_A_odVIc5ZV1_0),.clk(gclk));
	jdff dff_A_7BoI3UZc9_0(.dout(w_dff_A_PkAvAav43_0),.din(w_dff_A_7BoI3UZc9_0),.clk(gclk));
	jdff dff_A_PkAvAav43_0(.dout(w_dff_A_SWqQ5eqI6_0),.din(w_dff_A_PkAvAav43_0),.clk(gclk));
	jdff dff_A_SWqQ5eqI6_0(.dout(w_dff_A_e3fmwp449_0),.din(w_dff_A_SWqQ5eqI6_0),.clk(gclk));
	jdff dff_A_e3fmwp449_0(.dout(w_dff_A_MVXNSLyo2_0),.din(w_dff_A_e3fmwp449_0),.clk(gclk));
	jdff dff_A_MVXNSLyo2_0(.dout(w_dff_A_VnSc2x1S6_0),.din(w_dff_A_MVXNSLyo2_0),.clk(gclk));
	jdff dff_A_VnSc2x1S6_0(.dout(w_dff_A_wie0GAka4_0),.din(w_dff_A_VnSc2x1S6_0),.clk(gclk));
	jdff dff_A_wie0GAka4_0(.dout(w_dff_A_u7h5RBDN1_0),.din(w_dff_A_wie0GAka4_0),.clk(gclk));
	jdff dff_A_u7h5RBDN1_0(.dout(w_dff_A_OhoNtRXj1_0),.din(w_dff_A_u7h5RBDN1_0),.clk(gclk));
	jdff dff_A_OhoNtRXj1_0(.dout(w_dff_A_F8UnrKcz5_0),.din(w_dff_A_OhoNtRXj1_0),.clk(gclk));
	jdff dff_A_F8UnrKcz5_0(.dout(w_dff_A_0eBV2Zsm0_0),.din(w_dff_A_F8UnrKcz5_0),.clk(gclk));
	jdff dff_A_0eBV2Zsm0_0(.dout(w_dff_A_klwVrK1f0_0),.din(w_dff_A_0eBV2Zsm0_0),.clk(gclk));
	jdff dff_A_klwVrK1f0_0(.dout(w_dff_A_mCCNTPrw8_0),.din(w_dff_A_klwVrK1f0_0),.clk(gclk));
	jdff dff_A_mCCNTPrw8_0(.dout(w_dff_A_bB1MRMHH5_0),.din(w_dff_A_mCCNTPrw8_0),.clk(gclk));
	jdff dff_A_bB1MRMHH5_0(.dout(w_dff_A_ptbj28cO4_0),.din(w_dff_A_bB1MRMHH5_0),.clk(gclk));
	jdff dff_A_ptbj28cO4_0(.dout(w_dff_A_E3KHyVyE3_0),.din(w_dff_A_ptbj28cO4_0),.clk(gclk));
	jdff dff_A_E3KHyVyE3_0(.dout(w_dff_A_1zBUEotC4_0),.din(w_dff_A_E3KHyVyE3_0),.clk(gclk));
	jdff dff_A_1zBUEotC4_0(.dout(w_dff_A_pm7rt7Lx9_0),.din(w_dff_A_1zBUEotC4_0),.clk(gclk));
	jdff dff_A_pm7rt7Lx9_0(.dout(w_dff_A_XRa3pBrd2_0),.din(w_dff_A_pm7rt7Lx9_0),.clk(gclk));
	jdff dff_A_XRa3pBrd2_0(.dout(w_dff_A_dpu9OwYR6_0),.din(w_dff_A_XRa3pBrd2_0),.clk(gclk));
	jdff dff_A_dpu9OwYR6_0(.dout(w_dff_A_NUyaeWkZ0_0),.din(w_dff_A_dpu9OwYR6_0),.clk(gclk));
	jdff dff_A_NUyaeWkZ0_0(.dout(w_dff_A_oL8BaBJh7_0),.din(w_dff_A_NUyaeWkZ0_0),.clk(gclk));
	jdff dff_A_oL8BaBJh7_0(.dout(w_dff_A_Pf3ReiLo4_0),.din(w_dff_A_oL8BaBJh7_0),.clk(gclk));
	jdff dff_A_Pf3ReiLo4_0(.dout(w_dff_A_4mB0fYKv9_0),.din(w_dff_A_Pf3ReiLo4_0),.clk(gclk));
	jdff dff_A_4mB0fYKv9_0(.dout(f67),.din(w_dff_A_4mB0fYKv9_0),.clk(gclk));
	jdff dff_A_RBUkAX7b8_2(.dout(w_dff_A_RqmSUKBW9_0),.din(w_dff_A_RBUkAX7b8_2),.clk(gclk));
	jdff dff_A_RqmSUKBW9_0(.dout(w_dff_A_k3slauRu1_0),.din(w_dff_A_RqmSUKBW9_0),.clk(gclk));
	jdff dff_A_k3slauRu1_0(.dout(w_dff_A_GOpyHYSR9_0),.din(w_dff_A_k3slauRu1_0),.clk(gclk));
	jdff dff_A_GOpyHYSR9_0(.dout(w_dff_A_8hxzPRz46_0),.din(w_dff_A_GOpyHYSR9_0),.clk(gclk));
	jdff dff_A_8hxzPRz46_0(.dout(w_dff_A_QQYRPL7l8_0),.din(w_dff_A_8hxzPRz46_0),.clk(gclk));
	jdff dff_A_QQYRPL7l8_0(.dout(w_dff_A_z0ZztFCX1_0),.din(w_dff_A_QQYRPL7l8_0),.clk(gclk));
	jdff dff_A_z0ZztFCX1_0(.dout(w_dff_A_IYRw5uzD3_0),.din(w_dff_A_z0ZztFCX1_0),.clk(gclk));
	jdff dff_A_IYRw5uzD3_0(.dout(w_dff_A_hTuqk3668_0),.din(w_dff_A_IYRw5uzD3_0),.clk(gclk));
	jdff dff_A_hTuqk3668_0(.dout(w_dff_A_HxuQcyJS4_0),.din(w_dff_A_hTuqk3668_0),.clk(gclk));
	jdff dff_A_HxuQcyJS4_0(.dout(w_dff_A_DtjwSTAQ8_0),.din(w_dff_A_HxuQcyJS4_0),.clk(gclk));
	jdff dff_A_DtjwSTAQ8_0(.dout(w_dff_A_91SPmLkQ8_0),.din(w_dff_A_DtjwSTAQ8_0),.clk(gclk));
	jdff dff_A_91SPmLkQ8_0(.dout(w_dff_A_BgtOKDIh5_0),.din(w_dff_A_91SPmLkQ8_0),.clk(gclk));
	jdff dff_A_BgtOKDIh5_0(.dout(w_dff_A_BrDzreaM9_0),.din(w_dff_A_BgtOKDIh5_0),.clk(gclk));
	jdff dff_A_BrDzreaM9_0(.dout(w_dff_A_6HFMtDfJ2_0),.din(w_dff_A_BrDzreaM9_0),.clk(gclk));
	jdff dff_A_6HFMtDfJ2_0(.dout(w_dff_A_RAbNNNLW2_0),.din(w_dff_A_6HFMtDfJ2_0),.clk(gclk));
	jdff dff_A_RAbNNNLW2_0(.dout(w_dff_A_bukx1VUX6_0),.din(w_dff_A_RAbNNNLW2_0),.clk(gclk));
	jdff dff_A_bukx1VUX6_0(.dout(w_dff_A_5rsQSmNv9_0),.din(w_dff_A_bukx1VUX6_0),.clk(gclk));
	jdff dff_A_5rsQSmNv9_0(.dout(w_dff_A_fRTuTzJI9_0),.din(w_dff_A_5rsQSmNv9_0),.clk(gclk));
	jdff dff_A_fRTuTzJI9_0(.dout(w_dff_A_Yz5CW6DV2_0),.din(w_dff_A_fRTuTzJI9_0),.clk(gclk));
	jdff dff_A_Yz5CW6DV2_0(.dout(w_dff_A_dhICiPAr9_0),.din(w_dff_A_Yz5CW6DV2_0),.clk(gclk));
	jdff dff_A_dhICiPAr9_0(.dout(w_dff_A_2o5QjwcZ0_0),.din(w_dff_A_dhICiPAr9_0),.clk(gclk));
	jdff dff_A_2o5QjwcZ0_0(.dout(w_dff_A_EWVIJrGP1_0),.din(w_dff_A_2o5QjwcZ0_0),.clk(gclk));
	jdff dff_A_EWVIJrGP1_0(.dout(w_dff_A_b3HXEpiv9_0),.din(w_dff_A_EWVIJrGP1_0),.clk(gclk));
	jdff dff_A_b3HXEpiv9_0(.dout(w_dff_A_W0wvWbet7_0),.din(w_dff_A_b3HXEpiv9_0),.clk(gclk));
	jdff dff_A_W0wvWbet7_0(.dout(w_dff_A_B31JlHjo7_0),.din(w_dff_A_W0wvWbet7_0),.clk(gclk));
	jdff dff_A_B31JlHjo7_0(.dout(w_dff_A_zLAhlYtw6_0),.din(w_dff_A_B31JlHjo7_0),.clk(gclk));
	jdff dff_A_zLAhlYtw6_0(.dout(w_dff_A_izwGJfV66_0),.din(w_dff_A_zLAhlYtw6_0),.clk(gclk));
	jdff dff_A_izwGJfV66_0(.dout(w_dff_A_b9yXsjgx3_0),.din(w_dff_A_izwGJfV66_0),.clk(gclk));
	jdff dff_A_b9yXsjgx3_0(.dout(w_dff_A_kj1KkzTv0_0),.din(w_dff_A_b9yXsjgx3_0),.clk(gclk));
	jdff dff_A_kj1KkzTv0_0(.dout(w_dff_A_HgO7x0Lc8_0),.din(w_dff_A_kj1KkzTv0_0),.clk(gclk));
	jdff dff_A_HgO7x0Lc8_0(.dout(w_dff_A_u7WqldW85_0),.din(w_dff_A_HgO7x0Lc8_0),.clk(gclk));
	jdff dff_A_u7WqldW85_0(.dout(w_dff_A_50gaQkM69_0),.din(w_dff_A_u7WqldW85_0),.clk(gclk));
	jdff dff_A_50gaQkM69_0(.dout(w_dff_A_ZKlQ6WzA5_0),.din(w_dff_A_50gaQkM69_0),.clk(gclk));
	jdff dff_A_ZKlQ6WzA5_0(.dout(w_dff_A_KUMl4IoR8_0),.din(w_dff_A_ZKlQ6WzA5_0),.clk(gclk));
	jdff dff_A_KUMl4IoR8_0(.dout(w_dff_A_XgqRKVkx9_0),.din(w_dff_A_KUMl4IoR8_0),.clk(gclk));
	jdff dff_A_XgqRKVkx9_0(.dout(w_dff_A_iCEoBT3I6_0),.din(w_dff_A_XgqRKVkx9_0),.clk(gclk));
	jdff dff_A_iCEoBT3I6_0(.dout(w_dff_A_hjkRxXNl3_0),.din(w_dff_A_iCEoBT3I6_0),.clk(gclk));
	jdff dff_A_hjkRxXNl3_0(.dout(w_dff_A_GSPv2VuK4_0),.din(w_dff_A_hjkRxXNl3_0),.clk(gclk));
	jdff dff_A_GSPv2VuK4_0(.dout(w_dff_A_06bO7B0w1_0),.din(w_dff_A_GSPv2VuK4_0),.clk(gclk));
	jdff dff_A_06bO7B0w1_0(.dout(w_dff_A_zpECHwwR8_0),.din(w_dff_A_06bO7B0w1_0),.clk(gclk));
	jdff dff_A_zpECHwwR8_0(.dout(w_dff_A_Shfwh0Ce9_0),.din(w_dff_A_zpECHwwR8_0),.clk(gclk));
	jdff dff_A_Shfwh0Ce9_0(.dout(w_dff_A_wu1vCQuc4_0),.din(w_dff_A_Shfwh0Ce9_0),.clk(gclk));
	jdff dff_A_wu1vCQuc4_0(.dout(w_dff_A_0TV2RpM41_0),.din(w_dff_A_wu1vCQuc4_0),.clk(gclk));
	jdff dff_A_0TV2RpM41_0(.dout(w_dff_A_pB849hJ15_0),.din(w_dff_A_0TV2RpM41_0),.clk(gclk));
	jdff dff_A_pB849hJ15_0(.dout(w_dff_A_fjVHhmRR4_0),.din(w_dff_A_pB849hJ15_0),.clk(gclk));
	jdff dff_A_fjVHhmRR4_0(.dout(w_dff_A_5HcNXxXi3_0),.din(w_dff_A_fjVHhmRR4_0),.clk(gclk));
	jdff dff_A_5HcNXxXi3_0(.dout(w_dff_A_bTgzmGKw0_0),.din(w_dff_A_5HcNXxXi3_0),.clk(gclk));
	jdff dff_A_bTgzmGKw0_0(.dout(w_dff_A_ANew8Hpr0_0),.din(w_dff_A_bTgzmGKw0_0),.clk(gclk));
	jdff dff_A_ANew8Hpr0_0(.dout(w_dff_A_gfOrLxGB4_0),.din(w_dff_A_ANew8Hpr0_0),.clk(gclk));
	jdff dff_A_gfOrLxGB4_0(.dout(w_dff_A_gkg8OXmv0_0),.din(w_dff_A_gfOrLxGB4_0),.clk(gclk));
	jdff dff_A_gkg8OXmv0_0(.dout(w_dff_A_qDRJvr5m6_0),.din(w_dff_A_gkg8OXmv0_0),.clk(gclk));
	jdff dff_A_qDRJvr5m6_0(.dout(w_dff_A_8gqkAWhr3_0),.din(w_dff_A_qDRJvr5m6_0),.clk(gclk));
	jdff dff_A_8gqkAWhr3_0(.dout(w_dff_A_ciX2eJ1s5_0),.din(w_dff_A_8gqkAWhr3_0),.clk(gclk));
	jdff dff_A_ciX2eJ1s5_0(.dout(w_dff_A_sGm9nNKc4_0),.din(w_dff_A_ciX2eJ1s5_0),.clk(gclk));
	jdff dff_A_sGm9nNKc4_0(.dout(w_dff_A_Op5Zb9bh7_0),.din(w_dff_A_sGm9nNKc4_0),.clk(gclk));
	jdff dff_A_Op5Zb9bh7_0(.dout(w_dff_A_rouTpG8B3_0),.din(w_dff_A_Op5Zb9bh7_0),.clk(gclk));
	jdff dff_A_rouTpG8B3_0(.dout(w_dff_A_JrVaruuE8_0),.din(w_dff_A_rouTpG8B3_0),.clk(gclk));
	jdff dff_A_JrVaruuE8_0(.dout(w_dff_A_PnCdcSrA3_0),.din(w_dff_A_JrVaruuE8_0),.clk(gclk));
	jdff dff_A_PnCdcSrA3_0(.dout(f68),.din(w_dff_A_PnCdcSrA3_0),.clk(gclk));
	jdff dff_A_VF0Og0Ap9_2(.dout(w_dff_A_nXroSYXR2_0),.din(w_dff_A_VF0Og0Ap9_2),.clk(gclk));
	jdff dff_A_nXroSYXR2_0(.dout(w_dff_A_aK1T7m2b4_0),.din(w_dff_A_nXroSYXR2_0),.clk(gclk));
	jdff dff_A_aK1T7m2b4_0(.dout(w_dff_A_qDJPqAJt3_0),.din(w_dff_A_aK1T7m2b4_0),.clk(gclk));
	jdff dff_A_qDJPqAJt3_0(.dout(w_dff_A_FWJnlYk33_0),.din(w_dff_A_qDJPqAJt3_0),.clk(gclk));
	jdff dff_A_FWJnlYk33_0(.dout(w_dff_A_OmtCMLWa8_0),.din(w_dff_A_FWJnlYk33_0),.clk(gclk));
	jdff dff_A_OmtCMLWa8_0(.dout(w_dff_A_H2wdNp3t5_0),.din(w_dff_A_OmtCMLWa8_0),.clk(gclk));
	jdff dff_A_H2wdNp3t5_0(.dout(w_dff_A_TGmNPq249_0),.din(w_dff_A_H2wdNp3t5_0),.clk(gclk));
	jdff dff_A_TGmNPq249_0(.dout(w_dff_A_wX6PvLmZ4_0),.din(w_dff_A_TGmNPq249_0),.clk(gclk));
	jdff dff_A_wX6PvLmZ4_0(.dout(w_dff_A_Q9EfKqwD2_0),.din(w_dff_A_wX6PvLmZ4_0),.clk(gclk));
	jdff dff_A_Q9EfKqwD2_0(.dout(w_dff_A_EOea4nGB1_0),.din(w_dff_A_Q9EfKqwD2_0),.clk(gclk));
	jdff dff_A_EOea4nGB1_0(.dout(w_dff_A_JXFJdGuC6_0),.din(w_dff_A_EOea4nGB1_0),.clk(gclk));
	jdff dff_A_JXFJdGuC6_0(.dout(w_dff_A_95LZ5gRE2_0),.din(w_dff_A_JXFJdGuC6_0),.clk(gclk));
	jdff dff_A_95LZ5gRE2_0(.dout(w_dff_A_VEyQvFaV5_0),.din(w_dff_A_95LZ5gRE2_0),.clk(gclk));
	jdff dff_A_VEyQvFaV5_0(.dout(w_dff_A_v4u7p8A44_0),.din(w_dff_A_VEyQvFaV5_0),.clk(gclk));
	jdff dff_A_v4u7p8A44_0(.dout(w_dff_A_71B6alZp2_0),.din(w_dff_A_v4u7p8A44_0),.clk(gclk));
	jdff dff_A_71B6alZp2_0(.dout(w_dff_A_RVmWBXHU7_0),.din(w_dff_A_71B6alZp2_0),.clk(gclk));
	jdff dff_A_RVmWBXHU7_0(.dout(w_dff_A_HjRXXXPB7_0),.din(w_dff_A_RVmWBXHU7_0),.clk(gclk));
	jdff dff_A_HjRXXXPB7_0(.dout(w_dff_A_0xwNUpSI0_0),.din(w_dff_A_HjRXXXPB7_0),.clk(gclk));
	jdff dff_A_0xwNUpSI0_0(.dout(w_dff_A_tbiT7czn9_0),.din(w_dff_A_0xwNUpSI0_0),.clk(gclk));
	jdff dff_A_tbiT7czn9_0(.dout(w_dff_A_2g3snXTF8_0),.din(w_dff_A_tbiT7czn9_0),.clk(gclk));
	jdff dff_A_2g3snXTF8_0(.dout(w_dff_A_7LsueYe93_0),.din(w_dff_A_2g3snXTF8_0),.clk(gclk));
	jdff dff_A_7LsueYe93_0(.dout(w_dff_A_cXZ7DTNB5_0),.din(w_dff_A_7LsueYe93_0),.clk(gclk));
	jdff dff_A_cXZ7DTNB5_0(.dout(w_dff_A_rpyI8TVa0_0),.din(w_dff_A_cXZ7DTNB5_0),.clk(gclk));
	jdff dff_A_rpyI8TVa0_0(.dout(w_dff_A_BUDM2W8v1_0),.din(w_dff_A_rpyI8TVa0_0),.clk(gclk));
	jdff dff_A_BUDM2W8v1_0(.dout(w_dff_A_QilB8ZQ87_0),.din(w_dff_A_BUDM2W8v1_0),.clk(gclk));
	jdff dff_A_QilB8ZQ87_0(.dout(w_dff_A_rMMBb6jS4_0),.din(w_dff_A_QilB8ZQ87_0),.clk(gclk));
	jdff dff_A_rMMBb6jS4_0(.dout(w_dff_A_axOLZP2J1_0),.din(w_dff_A_rMMBb6jS4_0),.clk(gclk));
	jdff dff_A_axOLZP2J1_0(.dout(w_dff_A_85XXMsKB6_0),.din(w_dff_A_axOLZP2J1_0),.clk(gclk));
	jdff dff_A_85XXMsKB6_0(.dout(w_dff_A_cqnHyzI32_0),.din(w_dff_A_85XXMsKB6_0),.clk(gclk));
	jdff dff_A_cqnHyzI32_0(.dout(w_dff_A_gyDLYRcc6_0),.din(w_dff_A_cqnHyzI32_0),.clk(gclk));
	jdff dff_A_gyDLYRcc6_0(.dout(w_dff_A_t3uaLxwH3_0),.din(w_dff_A_gyDLYRcc6_0),.clk(gclk));
	jdff dff_A_t3uaLxwH3_0(.dout(w_dff_A_3LQGQ5d49_0),.din(w_dff_A_t3uaLxwH3_0),.clk(gclk));
	jdff dff_A_3LQGQ5d49_0(.dout(w_dff_A_TmS3uBVf2_0),.din(w_dff_A_3LQGQ5d49_0),.clk(gclk));
	jdff dff_A_TmS3uBVf2_0(.dout(w_dff_A_xqstLM2H5_0),.din(w_dff_A_TmS3uBVf2_0),.clk(gclk));
	jdff dff_A_xqstLM2H5_0(.dout(w_dff_A_CZQzgRln7_0),.din(w_dff_A_xqstLM2H5_0),.clk(gclk));
	jdff dff_A_CZQzgRln7_0(.dout(w_dff_A_k3Jti8gx8_0),.din(w_dff_A_CZQzgRln7_0),.clk(gclk));
	jdff dff_A_k3Jti8gx8_0(.dout(w_dff_A_qhgXhkMW8_0),.din(w_dff_A_k3Jti8gx8_0),.clk(gclk));
	jdff dff_A_qhgXhkMW8_0(.dout(w_dff_A_2J8ko5oa0_0),.din(w_dff_A_qhgXhkMW8_0),.clk(gclk));
	jdff dff_A_2J8ko5oa0_0(.dout(w_dff_A_q4P4oeuS3_0),.din(w_dff_A_2J8ko5oa0_0),.clk(gclk));
	jdff dff_A_q4P4oeuS3_0(.dout(w_dff_A_Zg312tyK9_0),.din(w_dff_A_q4P4oeuS3_0),.clk(gclk));
	jdff dff_A_Zg312tyK9_0(.dout(w_dff_A_NmfKAelC5_0),.din(w_dff_A_Zg312tyK9_0),.clk(gclk));
	jdff dff_A_NmfKAelC5_0(.dout(w_dff_A_5UUxAp4w6_0),.din(w_dff_A_NmfKAelC5_0),.clk(gclk));
	jdff dff_A_5UUxAp4w6_0(.dout(w_dff_A_nit1TOWV1_0),.din(w_dff_A_5UUxAp4w6_0),.clk(gclk));
	jdff dff_A_nit1TOWV1_0(.dout(w_dff_A_10If2VMj9_0),.din(w_dff_A_nit1TOWV1_0),.clk(gclk));
	jdff dff_A_10If2VMj9_0(.dout(w_dff_A_KSeGRj1L7_0),.din(w_dff_A_10If2VMj9_0),.clk(gclk));
	jdff dff_A_KSeGRj1L7_0(.dout(w_dff_A_8I7X3FGR3_0),.din(w_dff_A_KSeGRj1L7_0),.clk(gclk));
	jdff dff_A_8I7X3FGR3_0(.dout(w_dff_A_jbfB4KMr5_0),.din(w_dff_A_8I7X3FGR3_0),.clk(gclk));
	jdff dff_A_jbfB4KMr5_0(.dout(w_dff_A_WC0wZdX67_0),.din(w_dff_A_jbfB4KMr5_0),.clk(gclk));
	jdff dff_A_WC0wZdX67_0(.dout(w_dff_A_xLg8XN027_0),.din(w_dff_A_WC0wZdX67_0),.clk(gclk));
	jdff dff_A_xLg8XN027_0(.dout(w_dff_A_TNLK19AJ3_0),.din(w_dff_A_xLg8XN027_0),.clk(gclk));
	jdff dff_A_TNLK19AJ3_0(.dout(w_dff_A_H8Waqkww6_0),.din(w_dff_A_TNLK19AJ3_0),.clk(gclk));
	jdff dff_A_H8Waqkww6_0(.dout(w_dff_A_1aZCad728_0),.din(w_dff_A_H8Waqkww6_0),.clk(gclk));
	jdff dff_A_1aZCad728_0(.dout(w_dff_A_hv5F2UiU6_0),.din(w_dff_A_1aZCad728_0),.clk(gclk));
	jdff dff_A_hv5F2UiU6_0(.dout(w_dff_A_MGBGWR1K2_0),.din(w_dff_A_hv5F2UiU6_0),.clk(gclk));
	jdff dff_A_MGBGWR1K2_0(.dout(w_dff_A_dowjjR7S7_0),.din(w_dff_A_MGBGWR1K2_0),.clk(gclk));
	jdff dff_A_dowjjR7S7_0(.dout(w_dff_A_Qcl0AmRC5_0),.din(w_dff_A_dowjjR7S7_0),.clk(gclk));
	jdff dff_A_Qcl0AmRC5_0(.dout(w_dff_A_BrfBedkC6_0),.din(w_dff_A_Qcl0AmRC5_0),.clk(gclk));
	jdff dff_A_BrfBedkC6_0(.dout(f69),.din(w_dff_A_BrfBedkC6_0),.clk(gclk));
	jdff dff_A_uaH4n4Vl7_2(.dout(w_dff_A_Hq5zPYQD9_0),.din(w_dff_A_uaH4n4Vl7_2),.clk(gclk));
	jdff dff_A_Hq5zPYQD9_0(.dout(w_dff_A_Pecahs0b8_0),.din(w_dff_A_Hq5zPYQD9_0),.clk(gclk));
	jdff dff_A_Pecahs0b8_0(.dout(w_dff_A_gnoytxa32_0),.din(w_dff_A_Pecahs0b8_0),.clk(gclk));
	jdff dff_A_gnoytxa32_0(.dout(w_dff_A_KzdkcyGv7_0),.din(w_dff_A_gnoytxa32_0),.clk(gclk));
	jdff dff_A_KzdkcyGv7_0(.dout(w_dff_A_hhdyFl8l3_0),.din(w_dff_A_KzdkcyGv7_0),.clk(gclk));
	jdff dff_A_hhdyFl8l3_0(.dout(w_dff_A_a814e7N81_0),.din(w_dff_A_hhdyFl8l3_0),.clk(gclk));
	jdff dff_A_a814e7N81_0(.dout(w_dff_A_dsfP5vaW0_0),.din(w_dff_A_a814e7N81_0),.clk(gclk));
	jdff dff_A_dsfP5vaW0_0(.dout(w_dff_A_Ja7mqpbw9_0),.din(w_dff_A_dsfP5vaW0_0),.clk(gclk));
	jdff dff_A_Ja7mqpbw9_0(.dout(w_dff_A_NV2Dn7d30_0),.din(w_dff_A_Ja7mqpbw9_0),.clk(gclk));
	jdff dff_A_NV2Dn7d30_0(.dout(w_dff_A_rYk6j1yo4_0),.din(w_dff_A_NV2Dn7d30_0),.clk(gclk));
	jdff dff_A_rYk6j1yo4_0(.dout(w_dff_A_ZyjSC7Iw3_0),.din(w_dff_A_rYk6j1yo4_0),.clk(gclk));
	jdff dff_A_ZyjSC7Iw3_0(.dout(w_dff_A_4InucV121_0),.din(w_dff_A_ZyjSC7Iw3_0),.clk(gclk));
	jdff dff_A_4InucV121_0(.dout(w_dff_A_QpiFVyba8_0),.din(w_dff_A_4InucV121_0),.clk(gclk));
	jdff dff_A_QpiFVyba8_0(.dout(w_dff_A_QTfQJtRn0_0),.din(w_dff_A_QpiFVyba8_0),.clk(gclk));
	jdff dff_A_QTfQJtRn0_0(.dout(w_dff_A_NsEimduf1_0),.din(w_dff_A_QTfQJtRn0_0),.clk(gclk));
	jdff dff_A_NsEimduf1_0(.dout(w_dff_A_hwrVZa7V8_0),.din(w_dff_A_NsEimduf1_0),.clk(gclk));
	jdff dff_A_hwrVZa7V8_0(.dout(w_dff_A_AbMD8cxu8_0),.din(w_dff_A_hwrVZa7V8_0),.clk(gclk));
	jdff dff_A_AbMD8cxu8_0(.dout(w_dff_A_hqNDzVSf2_0),.din(w_dff_A_AbMD8cxu8_0),.clk(gclk));
	jdff dff_A_hqNDzVSf2_0(.dout(w_dff_A_uXz3jG643_0),.din(w_dff_A_hqNDzVSf2_0),.clk(gclk));
	jdff dff_A_uXz3jG643_0(.dout(w_dff_A_onf41rlz9_0),.din(w_dff_A_uXz3jG643_0),.clk(gclk));
	jdff dff_A_onf41rlz9_0(.dout(w_dff_A_dL6cUK7B6_0),.din(w_dff_A_onf41rlz9_0),.clk(gclk));
	jdff dff_A_dL6cUK7B6_0(.dout(w_dff_A_weIgDyLp5_0),.din(w_dff_A_dL6cUK7B6_0),.clk(gclk));
	jdff dff_A_weIgDyLp5_0(.dout(w_dff_A_XRZlYPQ88_0),.din(w_dff_A_weIgDyLp5_0),.clk(gclk));
	jdff dff_A_XRZlYPQ88_0(.dout(w_dff_A_HkakeBHP5_0),.din(w_dff_A_XRZlYPQ88_0),.clk(gclk));
	jdff dff_A_HkakeBHP5_0(.dout(w_dff_A_KT1eTXe82_0),.din(w_dff_A_HkakeBHP5_0),.clk(gclk));
	jdff dff_A_KT1eTXe82_0(.dout(w_dff_A_14p1WUOo1_0),.din(w_dff_A_KT1eTXe82_0),.clk(gclk));
	jdff dff_A_14p1WUOo1_0(.dout(w_dff_A_MtXNWzBZ7_0),.din(w_dff_A_14p1WUOo1_0),.clk(gclk));
	jdff dff_A_MtXNWzBZ7_0(.dout(w_dff_A_E4ejwqDF9_0),.din(w_dff_A_MtXNWzBZ7_0),.clk(gclk));
	jdff dff_A_E4ejwqDF9_0(.dout(w_dff_A_yYu0LAmn5_0),.din(w_dff_A_E4ejwqDF9_0),.clk(gclk));
	jdff dff_A_yYu0LAmn5_0(.dout(w_dff_A_zwhA3urF5_0),.din(w_dff_A_yYu0LAmn5_0),.clk(gclk));
	jdff dff_A_zwhA3urF5_0(.dout(w_dff_A_y3iSHKgA9_0),.din(w_dff_A_zwhA3urF5_0),.clk(gclk));
	jdff dff_A_y3iSHKgA9_0(.dout(w_dff_A_ElFiynBr4_0),.din(w_dff_A_y3iSHKgA9_0),.clk(gclk));
	jdff dff_A_ElFiynBr4_0(.dout(w_dff_A_bW1f51vt8_0),.din(w_dff_A_ElFiynBr4_0),.clk(gclk));
	jdff dff_A_bW1f51vt8_0(.dout(w_dff_A_kszowhPr5_0),.din(w_dff_A_bW1f51vt8_0),.clk(gclk));
	jdff dff_A_kszowhPr5_0(.dout(w_dff_A_mTHsZxYA7_0),.din(w_dff_A_kszowhPr5_0),.clk(gclk));
	jdff dff_A_mTHsZxYA7_0(.dout(w_dff_A_hu4Fzncz4_0),.din(w_dff_A_mTHsZxYA7_0),.clk(gclk));
	jdff dff_A_hu4Fzncz4_0(.dout(w_dff_A_Q1edSFGu6_0),.din(w_dff_A_hu4Fzncz4_0),.clk(gclk));
	jdff dff_A_Q1edSFGu6_0(.dout(w_dff_A_LD2x6Hs68_0),.din(w_dff_A_Q1edSFGu6_0),.clk(gclk));
	jdff dff_A_LD2x6Hs68_0(.dout(w_dff_A_27Foccp19_0),.din(w_dff_A_LD2x6Hs68_0),.clk(gclk));
	jdff dff_A_27Foccp19_0(.dout(w_dff_A_SnhIeawK0_0),.din(w_dff_A_27Foccp19_0),.clk(gclk));
	jdff dff_A_SnhIeawK0_0(.dout(w_dff_A_5933i80A5_0),.din(w_dff_A_SnhIeawK0_0),.clk(gclk));
	jdff dff_A_5933i80A5_0(.dout(w_dff_A_4yDJceyl1_0),.din(w_dff_A_5933i80A5_0),.clk(gclk));
	jdff dff_A_4yDJceyl1_0(.dout(w_dff_A_banPibvB0_0),.din(w_dff_A_4yDJceyl1_0),.clk(gclk));
	jdff dff_A_banPibvB0_0(.dout(w_dff_A_VcmAb1kX0_0),.din(w_dff_A_banPibvB0_0),.clk(gclk));
	jdff dff_A_VcmAb1kX0_0(.dout(w_dff_A_T4DsH9M93_0),.din(w_dff_A_VcmAb1kX0_0),.clk(gclk));
	jdff dff_A_T4DsH9M93_0(.dout(w_dff_A_JseL2veh6_0),.din(w_dff_A_T4DsH9M93_0),.clk(gclk));
	jdff dff_A_JseL2veh6_0(.dout(w_dff_A_ObIID1MB1_0),.din(w_dff_A_JseL2veh6_0),.clk(gclk));
	jdff dff_A_ObIID1MB1_0(.dout(w_dff_A_jRrr0lXe2_0),.din(w_dff_A_ObIID1MB1_0),.clk(gclk));
	jdff dff_A_jRrr0lXe2_0(.dout(w_dff_A_2QTABo543_0),.din(w_dff_A_jRrr0lXe2_0),.clk(gclk));
	jdff dff_A_2QTABo543_0(.dout(w_dff_A_JkhXQLb51_0),.din(w_dff_A_2QTABo543_0),.clk(gclk));
	jdff dff_A_JkhXQLb51_0(.dout(w_dff_A_u9L4L54q2_0),.din(w_dff_A_JkhXQLb51_0),.clk(gclk));
	jdff dff_A_u9L4L54q2_0(.dout(w_dff_A_KK3uU43V2_0),.din(w_dff_A_u9L4L54q2_0),.clk(gclk));
	jdff dff_A_KK3uU43V2_0(.dout(w_dff_A_ZSPUFDMw5_0),.din(w_dff_A_KK3uU43V2_0),.clk(gclk));
	jdff dff_A_ZSPUFDMw5_0(.dout(w_dff_A_OfVv51LF4_0),.din(w_dff_A_ZSPUFDMw5_0),.clk(gclk));
	jdff dff_A_OfVv51LF4_0(.dout(w_dff_A_AMHXt1sX3_0),.din(w_dff_A_OfVv51LF4_0),.clk(gclk));
	jdff dff_A_AMHXt1sX3_0(.dout(w_dff_A_wtn1PM5s4_0),.din(w_dff_A_AMHXt1sX3_0),.clk(gclk));
	jdff dff_A_wtn1PM5s4_0(.dout(f70),.din(w_dff_A_wtn1PM5s4_0),.clk(gclk));
	jdff dff_A_25rg4D9y4_2(.dout(w_dff_A_gMaUZ1Jh2_0),.din(w_dff_A_25rg4D9y4_2),.clk(gclk));
	jdff dff_A_gMaUZ1Jh2_0(.dout(w_dff_A_QDtMMZLA4_0),.din(w_dff_A_gMaUZ1Jh2_0),.clk(gclk));
	jdff dff_A_QDtMMZLA4_0(.dout(w_dff_A_z3ckPqi00_0),.din(w_dff_A_QDtMMZLA4_0),.clk(gclk));
	jdff dff_A_z3ckPqi00_0(.dout(w_dff_A_bENZVi647_0),.din(w_dff_A_z3ckPqi00_0),.clk(gclk));
	jdff dff_A_bENZVi647_0(.dout(w_dff_A_vUWQXntf0_0),.din(w_dff_A_bENZVi647_0),.clk(gclk));
	jdff dff_A_vUWQXntf0_0(.dout(w_dff_A_pmwqGBGK4_0),.din(w_dff_A_vUWQXntf0_0),.clk(gclk));
	jdff dff_A_pmwqGBGK4_0(.dout(w_dff_A_vefyXECb7_0),.din(w_dff_A_pmwqGBGK4_0),.clk(gclk));
	jdff dff_A_vefyXECb7_0(.dout(w_dff_A_sPN1vKtc6_0),.din(w_dff_A_vefyXECb7_0),.clk(gclk));
	jdff dff_A_sPN1vKtc6_0(.dout(w_dff_A_HEiSK3Hi9_0),.din(w_dff_A_sPN1vKtc6_0),.clk(gclk));
	jdff dff_A_HEiSK3Hi9_0(.dout(w_dff_A_IwfVey4W3_0),.din(w_dff_A_HEiSK3Hi9_0),.clk(gclk));
	jdff dff_A_IwfVey4W3_0(.dout(w_dff_A_bY9n5lJI0_0),.din(w_dff_A_IwfVey4W3_0),.clk(gclk));
	jdff dff_A_bY9n5lJI0_0(.dout(w_dff_A_NnrB3y8e7_0),.din(w_dff_A_bY9n5lJI0_0),.clk(gclk));
	jdff dff_A_NnrB3y8e7_0(.dout(w_dff_A_P3m1j59o6_0),.din(w_dff_A_NnrB3y8e7_0),.clk(gclk));
	jdff dff_A_P3m1j59o6_0(.dout(w_dff_A_FCy7iKye6_0),.din(w_dff_A_P3m1j59o6_0),.clk(gclk));
	jdff dff_A_FCy7iKye6_0(.dout(w_dff_A_2kk1vipH4_0),.din(w_dff_A_FCy7iKye6_0),.clk(gclk));
	jdff dff_A_2kk1vipH4_0(.dout(w_dff_A_RQC1bsqx4_0),.din(w_dff_A_2kk1vipH4_0),.clk(gclk));
	jdff dff_A_RQC1bsqx4_0(.dout(w_dff_A_MbW3SaUX7_0),.din(w_dff_A_RQC1bsqx4_0),.clk(gclk));
	jdff dff_A_MbW3SaUX7_0(.dout(w_dff_A_fkQ1ghpz0_0),.din(w_dff_A_MbW3SaUX7_0),.clk(gclk));
	jdff dff_A_fkQ1ghpz0_0(.dout(w_dff_A_fFssae2R6_0),.din(w_dff_A_fkQ1ghpz0_0),.clk(gclk));
	jdff dff_A_fFssae2R6_0(.dout(w_dff_A_ZnOTxnJF5_0),.din(w_dff_A_fFssae2R6_0),.clk(gclk));
	jdff dff_A_ZnOTxnJF5_0(.dout(w_dff_A_vC8adhUD8_0),.din(w_dff_A_ZnOTxnJF5_0),.clk(gclk));
	jdff dff_A_vC8adhUD8_0(.dout(w_dff_A_Qf1RcdE39_0),.din(w_dff_A_vC8adhUD8_0),.clk(gclk));
	jdff dff_A_Qf1RcdE39_0(.dout(w_dff_A_aDTZ1pvD4_0),.din(w_dff_A_Qf1RcdE39_0),.clk(gclk));
	jdff dff_A_aDTZ1pvD4_0(.dout(w_dff_A_eJiRy7R26_0),.din(w_dff_A_aDTZ1pvD4_0),.clk(gclk));
	jdff dff_A_eJiRy7R26_0(.dout(w_dff_A_yIJEqPa52_0),.din(w_dff_A_eJiRy7R26_0),.clk(gclk));
	jdff dff_A_yIJEqPa52_0(.dout(w_dff_A_fYxJTW1N1_0),.din(w_dff_A_yIJEqPa52_0),.clk(gclk));
	jdff dff_A_fYxJTW1N1_0(.dout(w_dff_A_mAVxwpLn9_0),.din(w_dff_A_fYxJTW1N1_0),.clk(gclk));
	jdff dff_A_mAVxwpLn9_0(.dout(w_dff_A_vc5pq8HC2_0),.din(w_dff_A_mAVxwpLn9_0),.clk(gclk));
	jdff dff_A_vc5pq8HC2_0(.dout(w_dff_A_M2WDqZ791_0),.din(w_dff_A_vc5pq8HC2_0),.clk(gclk));
	jdff dff_A_M2WDqZ791_0(.dout(w_dff_A_jLVdDsl13_0),.din(w_dff_A_M2WDqZ791_0),.clk(gclk));
	jdff dff_A_jLVdDsl13_0(.dout(w_dff_A_cSQmsN7w0_0),.din(w_dff_A_jLVdDsl13_0),.clk(gclk));
	jdff dff_A_cSQmsN7w0_0(.dout(w_dff_A_f7kUYoyW4_0),.din(w_dff_A_cSQmsN7w0_0),.clk(gclk));
	jdff dff_A_f7kUYoyW4_0(.dout(w_dff_A_dWnrxnrF5_0),.din(w_dff_A_f7kUYoyW4_0),.clk(gclk));
	jdff dff_A_dWnrxnrF5_0(.dout(w_dff_A_fNU093Xm9_0),.din(w_dff_A_dWnrxnrF5_0),.clk(gclk));
	jdff dff_A_fNU093Xm9_0(.dout(w_dff_A_L03vf5bo3_0),.din(w_dff_A_fNU093Xm9_0),.clk(gclk));
	jdff dff_A_L03vf5bo3_0(.dout(w_dff_A_2vfH541f0_0),.din(w_dff_A_L03vf5bo3_0),.clk(gclk));
	jdff dff_A_2vfH541f0_0(.dout(w_dff_A_VilYtPz80_0),.din(w_dff_A_2vfH541f0_0),.clk(gclk));
	jdff dff_A_VilYtPz80_0(.dout(w_dff_A_ktQotUcz1_0),.din(w_dff_A_VilYtPz80_0),.clk(gclk));
	jdff dff_A_ktQotUcz1_0(.dout(w_dff_A_mHBWCIWG5_0),.din(w_dff_A_ktQotUcz1_0),.clk(gclk));
	jdff dff_A_mHBWCIWG5_0(.dout(w_dff_A_qNZugnpd2_0),.din(w_dff_A_mHBWCIWG5_0),.clk(gclk));
	jdff dff_A_qNZugnpd2_0(.dout(w_dff_A_flTF9aTV4_0),.din(w_dff_A_qNZugnpd2_0),.clk(gclk));
	jdff dff_A_flTF9aTV4_0(.dout(w_dff_A_OKoF0kGo8_0),.din(w_dff_A_flTF9aTV4_0),.clk(gclk));
	jdff dff_A_OKoF0kGo8_0(.dout(w_dff_A_Ez745p549_0),.din(w_dff_A_OKoF0kGo8_0),.clk(gclk));
	jdff dff_A_Ez745p549_0(.dout(w_dff_A_dJ4jmv8Z2_0),.din(w_dff_A_Ez745p549_0),.clk(gclk));
	jdff dff_A_dJ4jmv8Z2_0(.dout(w_dff_A_zfrwsumQ8_0),.din(w_dff_A_dJ4jmv8Z2_0),.clk(gclk));
	jdff dff_A_zfrwsumQ8_0(.dout(w_dff_A_H9fWrUxV1_0),.din(w_dff_A_zfrwsumQ8_0),.clk(gclk));
	jdff dff_A_H9fWrUxV1_0(.dout(w_dff_A_ODj0rsdq4_0),.din(w_dff_A_H9fWrUxV1_0),.clk(gclk));
	jdff dff_A_ODj0rsdq4_0(.dout(w_dff_A_IyOT4q7o7_0),.din(w_dff_A_ODj0rsdq4_0),.clk(gclk));
	jdff dff_A_IyOT4q7o7_0(.dout(w_dff_A_jMp5qYgI5_0),.din(w_dff_A_IyOT4q7o7_0),.clk(gclk));
	jdff dff_A_jMp5qYgI5_0(.dout(w_dff_A_glD8vUMN1_0),.din(w_dff_A_jMp5qYgI5_0),.clk(gclk));
	jdff dff_A_glD8vUMN1_0(.dout(w_dff_A_0GrgOJQn6_0),.din(w_dff_A_glD8vUMN1_0),.clk(gclk));
	jdff dff_A_0GrgOJQn6_0(.dout(w_dff_A_8EHSVeXd8_0),.din(w_dff_A_0GrgOJQn6_0),.clk(gclk));
	jdff dff_A_8EHSVeXd8_0(.dout(w_dff_A_EwOzXb3T5_0),.din(w_dff_A_8EHSVeXd8_0),.clk(gclk));
	jdff dff_A_EwOzXb3T5_0(.dout(w_dff_A_CbmndSSj4_0),.din(w_dff_A_EwOzXb3T5_0),.clk(gclk));
	jdff dff_A_CbmndSSj4_0(.dout(w_dff_A_iMzLpSO62_0),.din(w_dff_A_CbmndSSj4_0),.clk(gclk));
	jdff dff_A_iMzLpSO62_0(.dout(f71),.din(w_dff_A_iMzLpSO62_0),.clk(gclk));
	jdff dff_A_DAfWDgLl4_2(.dout(w_dff_A_ormSNGoe1_0),.din(w_dff_A_DAfWDgLl4_2),.clk(gclk));
	jdff dff_A_ormSNGoe1_0(.dout(w_dff_A_A4LRAPuQ9_0),.din(w_dff_A_ormSNGoe1_0),.clk(gclk));
	jdff dff_A_A4LRAPuQ9_0(.dout(w_dff_A_82FIWrjE3_0),.din(w_dff_A_A4LRAPuQ9_0),.clk(gclk));
	jdff dff_A_82FIWrjE3_0(.dout(w_dff_A_y4UVvr3y6_0),.din(w_dff_A_82FIWrjE3_0),.clk(gclk));
	jdff dff_A_y4UVvr3y6_0(.dout(w_dff_A_ya35myYx5_0),.din(w_dff_A_y4UVvr3y6_0),.clk(gclk));
	jdff dff_A_ya35myYx5_0(.dout(w_dff_A_Lz4R1lWK5_0),.din(w_dff_A_ya35myYx5_0),.clk(gclk));
	jdff dff_A_Lz4R1lWK5_0(.dout(w_dff_A_Zhq6baI88_0),.din(w_dff_A_Lz4R1lWK5_0),.clk(gclk));
	jdff dff_A_Zhq6baI88_0(.dout(w_dff_A_5LBMkHLK3_0),.din(w_dff_A_Zhq6baI88_0),.clk(gclk));
	jdff dff_A_5LBMkHLK3_0(.dout(w_dff_A_y1S8iZjm6_0),.din(w_dff_A_5LBMkHLK3_0),.clk(gclk));
	jdff dff_A_y1S8iZjm6_0(.dout(w_dff_A_0q7vflWe0_0),.din(w_dff_A_y1S8iZjm6_0),.clk(gclk));
	jdff dff_A_0q7vflWe0_0(.dout(w_dff_A_kvoyxFSh5_0),.din(w_dff_A_0q7vflWe0_0),.clk(gclk));
	jdff dff_A_kvoyxFSh5_0(.dout(w_dff_A_6rq2NHXN9_0),.din(w_dff_A_kvoyxFSh5_0),.clk(gclk));
	jdff dff_A_6rq2NHXN9_0(.dout(w_dff_A_N6H7OTw20_0),.din(w_dff_A_6rq2NHXN9_0),.clk(gclk));
	jdff dff_A_N6H7OTw20_0(.dout(w_dff_A_4s2LNkBy1_0),.din(w_dff_A_N6H7OTw20_0),.clk(gclk));
	jdff dff_A_4s2LNkBy1_0(.dout(w_dff_A_DBd6t99U2_0),.din(w_dff_A_4s2LNkBy1_0),.clk(gclk));
	jdff dff_A_DBd6t99U2_0(.dout(w_dff_A_TlhoMpTp2_0),.din(w_dff_A_DBd6t99U2_0),.clk(gclk));
	jdff dff_A_TlhoMpTp2_0(.dout(w_dff_A_sXCjoh2K5_0),.din(w_dff_A_TlhoMpTp2_0),.clk(gclk));
	jdff dff_A_sXCjoh2K5_0(.dout(w_dff_A_rVVTBUHX2_0),.din(w_dff_A_sXCjoh2K5_0),.clk(gclk));
	jdff dff_A_rVVTBUHX2_0(.dout(w_dff_A_enFI1pD69_0),.din(w_dff_A_rVVTBUHX2_0),.clk(gclk));
	jdff dff_A_enFI1pD69_0(.dout(w_dff_A_6kmL7lfO7_0),.din(w_dff_A_enFI1pD69_0),.clk(gclk));
	jdff dff_A_6kmL7lfO7_0(.dout(w_dff_A_uZ5zQV233_0),.din(w_dff_A_6kmL7lfO7_0),.clk(gclk));
	jdff dff_A_uZ5zQV233_0(.dout(w_dff_A_74mrreFB9_0),.din(w_dff_A_uZ5zQV233_0),.clk(gclk));
	jdff dff_A_74mrreFB9_0(.dout(w_dff_A_P60Qy7Dr8_0),.din(w_dff_A_74mrreFB9_0),.clk(gclk));
	jdff dff_A_P60Qy7Dr8_0(.dout(w_dff_A_tz9aYjWz2_0),.din(w_dff_A_P60Qy7Dr8_0),.clk(gclk));
	jdff dff_A_tz9aYjWz2_0(.dout(w_dff_A_VIvHBkx90_0),.din(w_dff_A_tz9aYjWz2_0),.clk(gclk));
	jdff dff_A_VIvHBkx90_0(.dout(w_dff_A_ZHWJkbpj3_0),.din(w_dff_A_VIvHBkx90_0),.clk(gclk));
	jdff dff_A_ZHWJkbpj3_0(.dout(w_dff_A_MFwOKpof3_0),.din(w_dff_A_ZHWJkbpj3_0),.clk(gclk));
	jdff dff_A_MFwOKpof3_0(.dout(w_dff_A_i5LCXn107_0),.din(w_dff_A_MFwOKpof3_0),.clk(gclk));
	jdff dff_A_i5LCXn107_0(.dout(w_dff_A_6RK1onP97_0),.din(w_dff_A_i5LCXn107_0),.clk(gclk));
	jdff dff_A_6RK1onP97_0(.dout(w_dff_A_EFtX4gxT3_0),.din(w_dff_A_6RK1onP97_0),.clk(gclk));
	jdff dff_A_EFtX4gxT3_0(.dout(w_dff_A_gBmXod542_0),.din(w_dff_A_EFtX4gxT3_0),.clk(gclk));
	jdff dff_A_gBmXod542_0(.dout(w_dff_A_qQ4ElGug8_0),.din(w_dff_A_gBmXod542_0),.clk(gclk));
	jdff dff_A_qQ4ElGug8_0(.dout(w_dff_A_2sqKCUKN9_0),.din(w_dff_A_qQ4ElGug8_0),.clk(gclk));
	jdff dff_A_2sqKCUKN9_0(.dout(w_dff_A_O333e3BQ6_0),.din(w_dff_A_2sqKCUKN9_0),.clk(gclk));
	jdff dff_A_O333e3BQ6_0(.dout(w_dff_A_itSpDTOm5_0),.din(w_dff_A_O333e3BQ6_0),.clk(gclk));
	jdff dff_A_itSpDTOm5_0(.dout(w_dff_A_snOHc84O4_0),.din(w_dff_A_itSpDTOm5_0),.clk(gclk));
	jdff dff_A_snOHc84O4_0(.dout(w_dff_A_SxJRLB578_0),.din(w_dff_A_snOHc84O4_0),.clk(gclk));
	jdff dff_A_SxJRLB578_0(.dout(w_dff_A_QfYySoUh0_0),.din(w_dff_A_SxJRLB578_0),.clk(gclk));
	jdff dff_A_QfYySoUh0_0(.dout(w_dff_A_UErrL4eL8_0),.din(w_dff_A_QfYySoUh0_0),.clk(gclk));
	jdff dff_A_UErrL4eL8_0(.dout(w_dff_A_ajGKrzye8_0),.din(w_dff_A_UErrL4eL8_0),.clk(gclk));
	jdff dff_A_ajGKrzye8_0(.dout(w_dff_A_7tJ5UrSc9_0),.din(w_dff_A_ajGKrzye8_0),.clk(gclk));
	jdff dff_A_7tJ5UrSc9_0(.dout(w_dff_A_dZzbELHd9_0),.din(w_dff_A_7tJ5UrSc9_0),.clk(gclk));
	jdff dff_A_dZzbELHd9_0(.dout(w_dff_A_HgeQCjLO0_0),.din(w_dff_A_dZzbELHd9_0),.clk(gclk));
	jdff dff_A_HgeQCjLO0_0(.dout(w_dff_A_7L0cfby70_0),.din(w_dff_A_HgeQCjLO0_0),.clk(gclk));
	jdff dff_A_7L0cfby70_0(.dout(w_dff_A_eHO7v2ZO2_0),.din(w_dff_A_7L0cfby70_0),.clk(gclk));
	jdff dff_A_eHO7v2ZO2_0(.dout(w_dff_A_yV0xkws93_0),.din(w_dff_A_eHO7v2ZO2_0),.clk(gclk));
	jdff dff_A_yV0xkws93_0(.dout(w_dff_A_mkQ40IJp6_0),.din(w_dff_A_yV0xkws93_0),.clk(gclk));
	jdff dff_A_mkQ40IJp6_0(.dout(w_dff_A_fJOoY3RV1_0),.din(w_dff_A_mkQ40IJp6_0),.clk(gclk));
	jdff dff_A_fJOoY3RV1_0(.dout(w_dff_A_sfQWWVT60_0),.din(w_dff_A_fJOoY3RV1_0),.clk(gclk));
	jdff dff_A_sfQWWVT60_0(.dout(w_dff_A_NDhZpc6m9_0),.din(w_dff_A_sfQWWVT60_0),.clk(gclk));
	jdff dff_A_NDhZpc6m9_0(.dout(w_dff_A_cWvrTatd2_0),.din(w_dff_A_NDhZpc6m9_0),.clk(gclk));
	jdff dff_A_cWvrTatd2_0(.dout(w_dff_A_7FniTJ6t0_0),.din(w_dff_A_cWvrTatd2_0),.clk(gclk));
	jdff dff_A_7FniTJ6t0_0(.dout(w_dff_A_G8Up5KFD1_0),.din(w_dff_A_7FniTJ6t0_0),.clk(gclk));
	jdff dff_A_G8Up5KFD1_0(.dout(w_dff_A_ZNGIY1Kc2_0),.din(w_dff_A_G8Up5KFD1_0),.clk(gclk));
	jdff dff_A_ZNGIY1Kc2_0(.dout(f72),.din(w_dff_A_ZNGIY1Kc2_0),.clk(gclk));
	jdff dff_A_EXeMsU4S3_2(.dout(w_dff_A_Zln0oU877_0),.din(w_dff_A_EXeMsU4S3_2),.clk(gclk));
	jdff dff_A_Zln0oU877_0(.dout(w_dff_A_ddoOc77z5_0),.din(w_dff_A_Zln0oU877_0),.clk(gclk));
	jdff dff_A_ddoOc77z5_0(.dout(w_dff_A_OeswcQRV0_0),.din(w_dff_A_ddoOc77z5_0),.clk(gclk));
	jdff dff_A_OeswcQRV0_0(.dout(w_dff_A_7bPWMjHM8_0),.din(w_dff_A_OeswcQRV0_0),.clk(gclk));
	jdff dff_A_7bPWMjHM8_0(.dout(w_dff_A_Q3UYzNZ84_0),.din(w_dff_A_7bPWMjHM8_0),.clk(gclk));
	jdff dff_A_Q3UYzNZ84_0(.dout(w_dff_A_UiloeydJ2_0),.din(w_dff_A_Q3UYzNZ84_0),.clk(gclk));
	jdff dff_A_UiloeydJ2_0(.dout(w_dff_A_OJk86uQq0_0),.din(w_dff_A_UiloeydJ2_0),.clk(gclk));
	jdff dff_A_OJk86uQq0_0(.dout(w_dff_A_2uAwSGJB2_0),.din(w_dff_A_OJk86uQq0_0),.clk(gclk));
	jdff dff_A_2uAwSGJB2_0(.dout(w_dff_A_P84pQi9B8_0),.din(w_dff_A_2uAwSGJB2_0),.clk(gclk));
	jdff dff_A_P84pQi9B8_0(.dout(w_dff_A_1v0ZCuPY3_0),.din(w_dff_A_P84pQi9B8_0),.clk(gclk));
	jdff dff_A_1v0ZCuPY3_0(.dout(w_dff_A_r4WMnlBu6_0),.din(w_dff_A_1v0ZCuPY3_0),.clk(gclk));
	jdff dff_A_r4WMnlBu6_0(.dout(w_dff_A_vdf4uaYD4_0),.din(w_dff_A_r4WMnlBu6_0),.clk(gclk));
	jdff dff_A_vdf4uaYD4_0(.dout(w_dff_A_2kPOqpwC0_0),.din(w_dff_A_vdf4uaYD4_0),.clk(gclk));
	jdff dff_A_2kPOqpwC0_0(.dout(w_dff_A_kJcnqBpd1_0),.din(w_dff_A_2kPOqpwC0_0),.clk(gclk));
	jdff dff_A_kJcnqBpd1_0(.dout(w_dff_A_hT9RjCqx5_0),.din(w_dff_A_kJcnqBpd1_0),.clk(gclk));
	jdff dff_A_hT9RjCqx5_0(.dout(w_dff_A_26C6OUBy8_0),.din(w_dff_A_hT9RjCqx5_0),.clk(gclk));
	jdff dff_A_26C6OUBy8_0(.dout(w_dff_A_rHv977LH6_0),.din(w_dff_A_26C6OUBy8_0),.clk(gclk));
	jdff dff_A_rHv977LH6_0(.dout(w_dff_A_8yzyMVC58_0),.din(w_dff_A_rHv977LH6_0),.clk(gclk));
	jdff dff_A_8yzyMVC58_0(.dout(w_dff_A_R0f9gUP06_0),.din(w_dff_A_8yzyMVC58_0),.clk(gclk));
	jdff dff_A_R0f9gUP06_0(.dout(w_dff_A_vpHkwVLa3_0),.din(w_dff_A_R0f9gUP06_0),.clk(gclk));
	jdff dff_A_vpHkwVLa3_0(.dout(w_dff_A_57Z0k43U5_0),.din(w_dff_A_vpHkwVLa3_0),.clk(gclk));
	jdff dff_A_57Z0k43U5_0(.dout(w_dff_A_AVXp5ds75_0),.din(w_dff_A_57Z0k43U5_0),.clk(gclk));
	jdff dff_A_AVXp5ds75_0(.dout(w_dff_A_UrXnx3686_0),.din(w_dff_A_AVXp5ds75_0),.clk(gclk));
	jdff dff_A_UrXnx3686_0(.dout(w_dff_A_vExjHH2k7_0),.din(w_dff_A_UrXnx3686_0),.clk(gclk));
	jdff dff_A_vExjHH2k7_0(.dout(w_dff_A_qIxMHUAc7_0),.din(w_dff_A_vExjHH2k7_0),.clk(gclk));
	jdff dff_A_qIxMHUAc7_0(.dout(w_dff_A_DzVIQta27_0),.din(w_dff_A_qIxMHUAc7_0),.clk(gclk));
	jdff dff_A_DzVIQta27_0(.dout(w_dff_A_ir2Cgy7G3_0),.din(w_dff_A_DzVIQta27_0),.clk(gclk));
	jdff dff_A_ir2Cgy7G3_0(.dout(w_dff_A_UTSAnnYM9_0),.din(w_dff_A_ir2Cgy7G3_0),.clk(gclk));
	jdff dff_A_UTSAnnYM9_0(.dout(w_dff_A_oV688GxJ2_0),.din(w_dff_A_UTSAnnYM9_0),.clk(gclk));
	jdff dff_A_oV688GxJ2_0(.dout(w_dff_A_CU9778F21_0),.din(w_dff_A_oV688GxJ2_0),.clk(gclk));
	jdff dff_A_CU9778F21_0(.dout(w_dff_A_y8nwg7Q93_0),.din(w_dff_A_CU9778F21_0),.clk(gclk));
	jdff dff_A_y8nwg7Q93_0(.dout(w_dff_A_OSuq24jR4_0),.din(w_dff_A_y8nwg7Q93_0),.clk(gclk));
	jdff dff_A_OSuq24jR4_0(.dout(w_dff_A_jGRYtIQz1_0),.din(w_dff_A_OSuq24jR4_0),.clk(gclk));
	jdff dff_A_jGRYtIQz1_0(.dout(w_dff_A_abtHvNhj2_0),.din(w_dff_A_jGRYtIQz1_0),.clk(gclk));
	jdff dff_A_abtHvNhj2_0(.dout(w_dff_A_8qJ5ZTYG0_0),.din(w_dff_A_abtHvNhj2_0),.clk(gclk));
	jdff dff_A_8qJ5ZTYG0_0(.dout(w_dff_A_Q9Atw7Ot1_0),.din(w_dff_A_8qJ5ZTYG0_0),.clk(gclk));
	jdff dff_A_Q9Atw7Ot1_0(.dout(w_dff_A_OzSRRr1u3_0),.din(w_dff_A_Q9Atw7Ot1_0),.clk(gclk));
	jdff dff_A_OzSRRr1u3_0(.dout(w_dff_A_MhGw1nBV0_0),.din(w_dff_A_OzSRRr1u3_0),.clk(gclk));
	jdff dff_A_MhGw1nBV0_0(.dout(w_dff_A_JKg0nXE20_0),.din(w_dff_A_MhGw1nBV0_0),.clk(gclk));
	jdff dff_A_JKg0nXE20_0(.dout(w_dff_A_ioolUZBx4_0),.din(w_dff_A_JKg0nXE20_0),.clk(gclk));
	jdff dff_A_ioolUZBx4_0(.dout(w_dff_A_FCmgRkDz2_0),.din(w_dff_A_ioolUZBx4_0),.clk(gclk));
	jdff dff_A_FCmgRkDz2_0(.dout(w_dff_A_VesbgQ9o3_0),.din(w_dff_A_FCmgRkDz2_0),.clk(gclk));
	jdff dff_A_VesbgQ9o3_0(.dout(w_dff_A_pIdCw4Fc9_0),.din(w_dff_A_VesbgQ9o3_0),.clk(gclk));
	jdff dff_A_pIdCw4Fc9_0(.dout(w_dff_A_BYQxwySx2_0),.din(w_dff_A_pIdCw4Fc9_0),.clk(gclk));
	jdff dff_A_BYQxwySx2_0(.dout(w_dff_A_pCp4hosc2_0),.din(w_dff_A_BYQxwySx2_0),.clk(gclk));
	jdff dff_A_pCp4hosc2_0(.dout(w_dff_A_fxe47mxL9_0),.din(w_dff_A_pCp4hosc2_0),.clk(gclk));
	jdff dff_A_fxe47mxL9_0(.dout(w_dff_A_E7txir177_0),.din(w_dff_A_fxe47mxL9_0),.clk(gclk));
	jdff dff_A_E7txir177_0(.dout(w_dff_A_qRv1pvkc8_0),.din(w_dff_A_E7txir177_0),.clk(gclk));
	jdff dff_A_qRv1pvkc8_0(.dout(w_dff_A_MHwU2F0q6_0),.din(w_dff_A_qRv1pvkc8_0),.clk(gclk));
	jdff dff_A_MHwU2F0q6_0(.dout(w_dff_A_Gkfme8RG4_0),.din(w_dff_A_MHwU2F0q6_0),.clk(gclk));
	jdff dff_A_Gkfme8RG4_0(.dout(w_dff_A_niN05KA07_0),.din(w_dff_A_Gkfme8RG4_0),.clk(gclk));
	jdff dff_A_niN05KA07_0(.dout(w_dff_A_YPqapSkP7_0),.din(w_dff_A_niN05KA07_0),.clk(gclk));
	jdff dff_A_YPqapSkP7_0(.dout(w_dff_A_6q3kG0Zq9_0),.din(w_dff_A_YPqapSkP7_0),.clk(gclk));
	jdff dff_A_6q3kG0Zq9_0(.dout(f73),.din(w_dff_A_6q3kG0Zq9_0),.clk(gclk));
	jdff dff_A_kBneCYEu8_2(.dout(w_dff_A_TjZ8A8ix1_0),.din(w_dff_A_kBneCYEu8_2),.clk(gclk));
	jdff dff_A_TjZ8A8ix1_0(.dout(w_dff_A_1CiS67vV3_0),.din(w_dff_A_TjZ8A8ix1_0),.clk(gclk));
	jdff dff_A_1CiS67vV3_0(.dout(w_dff_A_z3bUp2Zk4_0),.din(w_dff_A_1CiS67vV3_0),.clk(gclk));
	jdff dff_A_z3bUp2Zk4_0(.dout(w_dff_A_vak0KR2D1_0),.din(w_dff_A_z3bUp2Zk4_0),.clk(gclk));
	jdff dff_A_vak0KR2D1_0(.dout(w_dff_A_24VX1jx52_0),.din(w_dff_A_vak0KR2D1_0),.clk(gclk));
	jdff dff_A_24VX1jx52_0(.dout(w_dff_A_BBODrWsH3_0),.din(w_dff_A_24VX1jx52_0),.clk(gclk));
	jdff dff_A_BBODrWsH3_0(.dout(w_dff_A_QZFHM5En2_0),.din(w_dff_A_BBODrWsH3_0),.clk(gclk));
	jdff dff_A_QZFHM5En2_0(.dout(w_dff_A_Wqhg9N3S4_0),.din(w_dff_A_QZFHM5En2_0),.clk(gclk));
	jdff dff_A_Wqhg9N3S4_0(.dout(w_dff_A_vXutZw1S8_0),.din(w_dff_A_Wqhg9N3S4_0),.clk(gclk));
	jdff dff_A_vXutZw1S8_0(.dout(w_dff_A_iciuHiHn6_0),.din(w_dff_A_vXutZw1S8_0),.clk(gclk));
	jdff dff_A_iciuHiHn6_0(.dout(w_dff_A_XcqqFZXf3_0),.din(w_dff_A_iciuHiHn6_0),.clk(gclk));
	jdff dff_A_XcqqFZXf3_0(.dout(w_dff_A_VTwqFdWs4_0),.din(w_dff_A_XcqqFZXf3_0),.clk(gclk));
	jdff dff_A_VTwqFdWs4_0(.dout(w_dff_A_0cNmxHt89_0),.din(w_dff_A_VTwqFdWs4_0),.clk(gclk));
	jdff dff_A_0cNmxHt89_0(.dout(w_dff_A_MLzdOCKr7_0),.din(w_dff_A_0cNmxHt89_0),.clk(gclk));
	jdff dff_A_MLzdOCKr7_0(.dout(w_dff_A_fQHa6Clv4_0),.din(w_dff_A_MLzdOCKr7_0),.clk(gclk));
	jdff dff_A_fQHa6Clv4_0(.dout(w_dff_A_RsHvLwOe4_0),.din(w_dff_A_fQHa6Clv4_0),.clk(gclk));
	jdff dff_A_RsHvLwOe4_0(.dout(w_dff_A_8SA1rCrf5_0),.din(w_dff_A_RsHvLwOe4_0),.clk(gclk));
	jdff dff_A_8SA1rCrf5_0(.dout(w_dff_A_zp4Gajy60_0),.din(w_dff_A_8SA1rCrf5_0),.clk(gclk));
	jdff dff_A_zp4Gajy60_0(.dout(w_dff_A_ZuFX1YDI5_0),.din(w_dff_A_zp4Gajy60_0),.clk(gclk));
	jdff dff_A_ZuFX1YDI5_0(.dout(w_dff_A_kptl2weY5_0),.din(w_dff_A_ZuFX1YDI5_0),.clk(gclk));
	jdff dff_A_kptl2weY5_0(.dout(w_dff_A_pziyDUgK7_0),.din(w_dff_A_kptl2weY5_0),.clk(gclk));
	jdff dff_A_pziyDUgK7_0(.dout(w_dff_A_W0DkZNNM0_0),.din(w_dff_A_pziyDUgK7_0),.clk(gclk));
	jdff dff_A_W0DkZNNM0_0(.dout(w_dff_A_9EVxH0J33_0),.din(w_dff_A_W0DkZNNM0_0),.clk(gclk));
	jdff dff_A_9EVxH0J33_0(.dout(w_dff_A_KgcQRq7J0_0),.din(w_dff_A_9EVxH0J33_0),.clk(gclk));
	jdff dff_A_KgcQRq7J0_0(.dout(w_dff_A_ne4hKc6D9_0),.din(w_dff_A_KgcQRq7J0_0),.clk(gclk));
	jdff dff_A_ne4hKc6D9_0(.dout(w_dff_A_pUAhSRLv2_0),.din(w_dff_A_ne4hKc6D9_0),.clk(gclk));
	jdff dff_A_pUAhSRLv2_0(.dout(w_dff_A_kdHeE7md9_0),.din(w_dff_A_pUAhSRLv2_0),.clk(gclk));
	jdff dff_A_kdHeE7md9_0(.dout(w_dff_A_BnSrrkiE1_0),.din(w_dff_A_kdHeE7md9_0),.clk(gclk));
	jdff dff_A_BnSrrkiE1_0(.dout(w_dff_A_5oIOcmNt4_0),.din(w_dff_A_BnSrrkiE1_0),.clk(gclk));
	jdff dff_A_5oIOcmNt4_0(.dout(w_dff_A_soqyhzV73_0),.din(w_dff_A_5oIOcmNt4_0),.clk(gclk));
	jdff dff_A_soqyhzV73_0(.dout(w_dff_A_KOeJhbke1_0),.din(w_dff_A_soqyhzV73_0),.clk(gclk));
	jdff dff_A_KOeJhbke1_0(.dout(w_dff_A_e0HoVtt94_0),.din(w_dff_A_KOeJhbke1_0),.clk(gclk));
	jdff dff_A_e0HoVtt94_0(.dout(w_dff_A_THonSYaz8_0),.din(w_dff_A_e0HoVtt94_0),.clk(gclk));
	jdff dff_A_THonSYaz8_0(.dout(w_dff_A_kE2YiNZ35_0),.din(w_dff_A_THonSYaz8_0),.clk(gclk));
	jdff dff_A_kE2YiNZ35_0(.dout(w_dff_A_WgHD6dXx9_0),.din(w_dff_A_kE2YiNZ35_0),.clk(gclk));
	jdff dff_A_WgHD6dXx9_0(.dout(w_dff_A_jiVWknzQ8_0),.din(w_dff_A_WgHD6dXx9_0),.clk(gclk));
	jdff dff_A_jiVWknzQ8_0(.dout(w_dff_A_9xRPcLUh0_0),.din(w_dff_A_jiVWknzQ8_0),.clk(gclk));
	jdff dff_A_9xRPcLUh0_0(.dout(w_dff_A_eENqY71f0_0),.din(w_dff_A_9xRPcLUh0_0),.clk(gclk));
	jdff dff_A_eENqY71f0_0(.dout(w_dff_A_1nvxvxJw7_0),.din(w_dff_A_eENqY71f0_0),.clk(gclk));
	jdff dff_A_1nvxvxJw7_0(.dout(w_dff_A_myuGvPEX5_0),.din(w_dff_A_1nvxvxJw7_0),.clk(gclk));
	jdff dff_A_myuGvPEX5_0(.dout(w_dff_A_zZ8XX7Im6_0),.din(w_dff_A_myuGvPEX5_0),.clk(gclk));
	jdff dff_A_zZ8XX7Im6_0(.dout(w_dff_A_m9GsMBpB0_0),.din(w_dff_A_zZ8XX7Im6_0),.clk(gclk));
	jdff dff_A_m9GsMBpB0_0(.dout(w_dff_A_h6jeR5BS2_0),.din(w_dff_A_m9GsMBpB0_0),.clk(gclk));
	jdff dff_A_h6jeR5BS2_0(.dout(w_dff_A_JQXCwFgF8_0),.din(w_dff_A_h6jeR5BS2_0),.clk(gclk));
	jdff dff_A_JQXCwFgF8_0(.dout(w_dff_A_7TUpj4h75_0),.din(w_dff_A_JQXCwFgF8_0),.clk(gclk));
	jdff dff_A_7TUpj4h75_0(.dout(w_dff_A_CyI9Vjt95_0),.din(w_dff_A_7TUpj4h75_0),.clk(gclk));
	jdff dff_A_CyI9Vjt95_0(.dout(w_dff_A_1aMdhNC21_0),.din(w_dff_A_CyI9Vjt95_0),.clk(gclk));
	jdff dff_A_1aMdhNC21_0(.dout(w_dff_A_y3Sh4eqa6_0),.din(w_dff_A_1aMdhNC21_0),.clk(gclk));
	jdff dff_A_y3Sh4eqa6_0(.dout(w_dff_A_fFGGIFZt1_0),.din(w_dff_A_y3Sh4eqa6_0),.clk(gclk));
	jdff dff_A_fFGGIFZt1_0(.dout(w_dff_A_UTQRMyaE7_0),.din(w_dff_A_fFGGIFZt1_0),.clk(gclk));
	jdff dff_A_UTQRMyaE7_0(.dout(w_dff_A_tf7ayJ1u7_0),.din(w_dff_A_UTQRMyaE7_0),.clk(gclk));
	jdff dff_A_tf7ayJ1u7_0(.dout(w_dff_A_no3YE7WY7_0),.din(w_dff_A_tf7ayJ1u7_0),.clk(gclk));
	jdff dff_A_no3YE7WY7_0(.dout(f74),.din(w_dff_A_no3YE7WY7_0),.clk(gclk));
	jdff dff_A_50Y8hj8Y4_2(.dout(w_dff_A_380q8mam8_0),.din(w_dff_A_50Y8hj8Y4_2),.clk(gclk));
	jdff dff_A_380q8mam8_0(.dout(w_dff_A_X7oXyS1x2_0),.din(w_dff_A_380q8mam8_0),.clk(gclk));
	jdff dff_A_X7oXyS1x2_0(.dout(w_dff_A_wpkHACFW3_0),.din(w_dff_A_X7oXyS1x2_0),.clk(gclk));
	jdff dff_A_wpkHACFW3_0(.dout(w_dff_A_InvMEHLe4_0),.din(w_dff_A_wpkHACFW3_0),.clk(gclk));
	jdff dff_A_InvMEHLe4_0(.dout(w_dff_A_F5HCMXON9_0),.din(w_dff_A_InvMEHLe4_0),.clk(gclk));
	jdff dff_A_F5HCMXON9_0(.dout(w_dff_A_CfyqoSyP1_0),.din(w_dff_A_F5HCMXON9_0),.clk(gclk));
	jdff dff_A_CfyqoSyP1_0(.dout(w_dff_A_toM6jEcl8_0),.din(w_dff_A_CfyqoSyP1_0),.clk(gclk));
	jdff dff_A_toM6jEcl8_0(.dout(w_dff_A_pwGVKEoY9_0),.din(w_dff_A_toM6jEcl8_0),.clk(gclk));
	jdff dff_A_pwGVKEoY9_0(.dout(w_dff_A_DZHNMTCB6_0),.din(w_dff_A_pwGVKEoY9_0),.clk(gclk));
	jdff dff_A_DZHNMTCB6_0(.dout(w_dff_A_4O5YjEMr2_0),.din(w_dff_A_DZHNMTCB6_0),.clk(gclk));
	jdff dff_A_4O5YjEMr2_0(.dout(w_dff_A_l8rg3K4r0_0),.din(w_dff_A_4O5YjEMr2_0),.clk(gclk));
	jdff dff_A_l8rg3K4r0_0(.dout(w_dff_A_coYJSFtM3_0),.din(w_dff_A_l8rg3K4r0_0),.clk(gclk));
	jdff dff_A_coYJSFtM3_0(.dout(w_dff_A_QaFodfrU7_0),.din(w_dff_A_coYJSFtM3_0),.clk(gclk));
	jdff dff_A_QaFodfrU7_0(.dout(w_dff_A_6eLxX7186_0),.din(w_dff_A_QaFodfrU7_0),.clk(gclk));
	jdff dff_A_6eLxX7186_0(.dout(w_dff_A_JqWqSuk32_0),.din(w_dff_A_6eLxX7186_0),.clk(gclk));
	jdff dff_A_JqWqSuk32_0(.dout(w_dff_A_yhKe7tuk4_0),.din(w_dff_A_JqWqSuk32_0),.clk(gclk));
	jdff dff_A_yhKe7tuk4_0(.dout(w_dff_A_4lsRD3MB4_0),.din(w_dff_A_yhKe7tuk4_0),.clk(gclk));
	jdff dff_A_4lsRD3MB4_0(.dout(w_dff_A_xnRVGa5p6_0),.din(w_dff_A_4lsRD3MB4_0),.clk(gclk));
	jdff dff_A_xnRVGa5p6_0(.dout(w_dff_A_dE1dSX6n5_0),.din(w_dff_A_xnRVGa5p6_0),.clk(gclk));
	jdff dff_A_dE1dSX6n5_0(.dout(w_dff_A_wYYNfpNG8_0),.din(w_dff_A_dE1dSX6n5_0),.clk(gclk));
	jdff dff_A_wYYNfpNG8_0(.dout(w_dff_A_ogNIVGzk8_0),.din(w_dff_A_wYYNfpNG8_0),.clk(gclk));
	jdff dff_A_ogNIVGzk8_0(.dout(w_dff_A_4mpehFMg3_0),.din(w_dff_A_ogNIVGzk8_0),.clk(gclk));
	jdff dff_A_4mpehFMg3_0(.dout(w_dff_A_un4NtM2z2_0),.din(w_dff_A_4mpehFMg3_0),.clk(gclk));
	jdff dff_A_un4NtM2z2_0(.dout(w_dff_A_0XgpDvg60_0),.din(w_dff_A_un4NtM2z2_0),.clk(gclk));
	jdff dff_A_0XgpDvg60_0(.dout(w_dff_A_g1mL9q8a0_0),.din(w_dff_A_0XgpDvg60_0),.clk(gclk));
	jdff dff_A_g1mL9q8a0_0(.dout(w_dff_A_UuSyHXzk4_0),.din(w_dff_A_g1mL9q8a0_0),.clk(gclk));
	jdff dff_A_UuSyHXzk4_0(.dout(w_dff_A_kf3VfFNM8_0),.din(w_dff_A_UuSyHXzk4_0),.clk(gclk));
	jdff dff_A_kf3VfFNM8_0(.dout(w_dff_A_BAYqhi505_0),.din(w_dff_A_kf3VfFNM8_0),.clk(gclk));
	jdff dff_A_BAYqhi505_0(.dout(w_dff_A_qfmkJNyU5_0),.din(w_dff_A_BAYqhi505_0),.clk(gclk));
	jdff dff_A_qfmkJNyU5_0(.dout(w_dff_A_IsOkEG7z2_0),.din(w_dff_A_qfmkJNyU5_0),.clk(gclk));
	jdff dff_A_IsOkEG7z2_0(.dout(w_dff_A_7UcO0olk3_0),.din(w_dff_A_IsOkEG7z2_0),.clk(gclk));
	jdff dff_A_7UcO0olk3_0(.dout(w_dff_A_MC7xgw8y3_0),.din(w_dff_A_7UcO0olk3_0),.clk(gclk));
	jdff dff_A_MC7xgw8y3_0(.dout(w_dff_A_6ZozluVv2_0),.din(w_dff_A_MC7xgw8y3_0),.clk(gclk));
	jdff dff_A_6ZozluVv2_0(.dout(w_dff_A_NdlSg1HD2_0),.din(w_dff_A_6ZozluVv2_0),.clk(gclk));
	jdff dff_A_NdlSg1HD2_0(.dout(w_dff_A_mWpxkfQk3_0),.din(w_dff_A_NdlSg1HD2_0),.clk(gclk));
	jdff dff_A_mWpxkfQk3_0(.dout(w_dff_A_0DbrXdlQ5_0),.din(w_dff_A_mWpxkfQk3_0),.clk(gclk));
	jdff dff_A_0DbrXdlQ5_0(.dout(w_dff_A_LRVsfhoq9_0),.din(w_dff_A_0DbrXdlQ5_0),.clk(gclk));
	jdff dff_A_LRVsfhoq9_0(.dout(w_dff_A_2kNjDGHY6_0),.din(w_dff_A_LRVsfhoq9_0),.clk(gclk));
	jdff dff_A_2kNjDGHY6_0(.dout(w_dff_A_ED7W3lqk3_0),.din(w_dff_A_2kNjDGHY6_0),.clk(gclk));
	jdff dff_A_ED7W3lqk3_0(.dout(w_dff_A_5T9p8brr2_0),.din(w_dff_A_ED7W3lqk3_0),.clk(gclk));
	jdff dff_A_5T9p8brr2_0(.dout(w_dff_A_8XdNfzqJ0_0),.din(w_dff_A_5T9p8brr2_0),.clk(gclk));
	jdff dff_A_8XdNfzqJ0_0(.dout(w_dff_A_wnWDUmlG4_0),.din(w_dff_A_8XdNfzqJ0_0),.clk(gclk));
	jdff dff_A_wnWDUmlG4_0(.dout(w_dff_A_cflT37il6_0),.din(w_dff_A_wnWDUmlG4_0),.clk(gclk));
	jdff dff_A_cflT37il6_0(.dout(w_dff_A_RCc5bRBT7_0),.din(w_dff_A_cflT37il6_0),.clk(gclk));
	jdff dff_A_RCc5bRBT7_0(.dout(w_dff_A_cYHMH3aM1_0),.din(w_dff_A_RCc5bRBT7_0),.clk(gclk));
	jdff dff_A_cYHMH3aM1_0(.dout(w_dff_A_eeJVynR56_0),.din(w_dff_A_cYHMH3aM1_0),.clk(gclk));
	jdff dff_A_eeJVynR56_0(.dout(w_dff_A_tN2npZYH6_0),.din(w_dff_A_eeJVynR56_0),.clk(gclk));
	jdff dff_A_tN2npZYH6_0(.dout(w_dff_A_8uOQsRJz6_0),.din(w_dff_A_tN2npZYH6_0),.clk(gclk));
	jdff dff_A_8uOQsRJz6_0(.dout(w_dff_A_xcl1jDOn2_0),.din(w_dff_A_8uOQsRJz6_0),.clk(gclk));
	jdff dff_A_xcl1jDOn2_0(.dout(w_dff_A_kluZOFwr9_0),.din(w_dff_A_xcl1jDOn2_0),.clk(gclk));
	jdff dff_A_kluZOFwr9_0(.dout(w_dff_A_LNISbhLH8_0),.din(w_dff_A_kluZOFwr9_0),.clk(gclk));
	jdff dff_A_LNISbhLH8_0(.dout(f75),.din(w_dff_A_LNISbhLH8_0),.clk(gclk));
	jdff dff_A_uKcBLu2n9_2(.dout(w_dff_A_HvNlbdOs7_0),.din(w_dff_A_uKcBLu2n9_2),.clk(gclk));
	jdff dff_A_HvNlbdOs7_0(.dout(w_dff_A_uQeD9Zd16_0),.din(w_dff_A_HvNlbdOs7_0),.clk(gclk));
	jdff dff_A_uQeD9Zd16_0(.dout(w_dff_A_m9g9yRsp0_0),.din(w_dff_A_uQeD9Zd16_0),.clk(gclk));
	jdff dff_A_m9g9yRsp0_0(.dout(w_dff_A_YZtPaWrA2_0),.din(w_dff_A_m9g9yRsp0_0),.clk(gclk));
	jdff dff_A_YZtPaWrA2_0(.dout(w_dff_A_bXAxPrgJ7_0),.din(w_dff_A_YZtPaWrA2_0),.clk(gclk));
	jdff dff_A_bXAxPrgJ7_0(.dout(w_dff_A_QtZzEh6R8_0),.din(w_dff_A_bXAxPrgJ7_0),.clk(gclk));
	jdff dff_A_QtZzEh6R8_0(.dout(w_dff_A_nMPD83vr7_0),.din(w_dff_A_QtZzEh6R8_0),.clk(gclk));
	jdff dff_A_nMPD83vr7_0(.dout(w_dff_A_901p4X1c4_0),.din(w_dff_A_nMPD83vr7_0),.clk(gclk));
	jdff dff_A_901p4X1c4_0(.dout(w_dff_A_tNy2uyJd2_0),.din(w_dff_A_901p4X1c4_0),.clk(gclk));
	jdff dff_A_tNy2uyJd2_0(.dout(w_dff_A_Z8HE94be5_0),.din(w_dff_A_tNy2uyJd2_0),.clk(gclk));
	jdff dff_A_Z8HE94be5_0(.dout(w_dff_A_436MqNVQ4_0),.din(w_dff_A_Z8HE94be5_0),.clk(gclk));
	jdff dff_A_436MqNVQ4_0(.dout(w_dff_A_yBhTrM2j2_0),.din(w_dff_A_436MqNVQ4_0),.clk(gclk));
	jdff dff_A_yBhTrM2j2_0(.dout(w_dff_A_nVf6cY2P2_0),.din(w_dff_A_yBhTrM2j2_0),.clk(gclk));
	jdff dff_A_nVf6cY2P2_0(.dout(w_dff_A_fOnTduJx7_0),.din(w_dff_A_nVf6cY2P2_0),.clk(gclk));
	jdff dff_A_fOnTduJx7_0(.dout(w_dff_A_ZBjk75Cn0_0),.din(w_dff_A_fOnTduJx7_0),.clk(gclk));
	jdff dff_A_ZBjk75Cn0_0(.dout(w_dff_A_2Cz1N7jj6_0),.din(w_dff_A_ZBjk75Cn0_0),.clk(gclk));
	jdff dff_A_2Cz1N7jj6_0(.dout(w_dff_A_3198nwiY2_0),.din(w_dff_A_2Cz1N7jj6_0),.clk(gclk));
	jdff dff_A_3198nwiY2_0(.dout(w_dff_A_TwRnH3f17_0),.din(w_dff_A_3198nwiY2_0),.clk(gclk));
	jdff dff_A_TwRnH3f17_0(.dout(w_dff_A_439zFR8x0_0),.din(w_dff_A_TwRnH3f17_0),.clk(gclk));
	jdff dff_A_439zFR8x0_0(.dout(w_dff_A_8mnjl5YU9_0),.din(w_dff_A_439zFR8x0_0),.clk(gclk));
	jdff dff_A_8mnjl5YU9_0(.dout(w_dff_A_RzUwzywh2_0),.din(w_dff_A_8mnjl5YU9_0),.clk(gclk));
	jdff dff_A_RzUwzywh2_0(.dout(w_dff_A_HCsF6nf21_0),.din(w_dff_A_RzUwzywh2_0),.clk(gclk));
	jdff dff_A_HCsF6nf21_0(.dout(w_dff_A_jkqJqvUh4_0),.din(w_dff_A_HCsF6nf21_0),.clk(gclk));
	jdff dff_A_jkqJqvUh4_0(.dout(w_dff_A_jWjWDhNx5_0),.din(w_dff_A_jkqJqvUh4_0),.clk(gclk));
	jdff dff_A_jWjWDhNx5_0(.dout(w_dff_A_vVNBJofN9_0),.din(w_dff_A_jWjWDhNx5_0),.clk(gclk));
	jdff dff_A_vVNBJofN9_0(.dout(w_dff_A_LVqNfCzz6_0),.din(w_dff_A_vVNBJofN9_0),.clk(gclk));
	jdff dff_A_LVqNfCzz6_0(.dout(w_dff_A_I813dbL64_0),.din(w_dff_A_LVqNfCzz6_0),.clk(gclk));
	jdff dff_A_I813dbL64_0(.dout(w_dff_A_5zUbsZL49_0),.din(w_dff_A_I813dbL64_0),.clk(gclk));
	jdff dff_A_5zUbsZL49_0(.dout(w_dff_A_emKkbmS10_0),.din(w_dff_A_5zUbsZL49_0),.clk(gclk));
	jdff dff_A_emKkbmS10_0(.dout(w_dff_A_Bk4Yr6xp4_0),.din(w_dff_A_emKkbmS10_0),.clk(gclk));
	jdff dff_A_Bk4Yr6xp4_0(.dout(w_dff_A_FpDYd6Yp6_0),.din(w_dff_A_Bk4Yr6xp4_0),.clk(gclk));
	jdff dff_A_FpDYd6Yp6_0(.dout(w_dff_A_Iu8gJkor6_0),.din(w_dff_A_FpDYd6Yp6_0),.clk(gclk));
	jdff dff_A_Iu8gJkor6_0(.dout(w_dff_A_22N3g46E3_0),.din(w_dff_A_Iu8gJkor6_0),.clk(gclk));
	jdff dff_A_22N3g46E3_0(.dout(w_dff_A_oh8Sdo6k9_0),.din(w_dff_A_22N3g46E3_0),.clk(gclk));
	jdff dff_A_oh8Sdo6k9_0(.dout(w_dff_A_q6da7xD82_0),.din(w_dff_A_oh8Sdo6k9_0),.clk(gclk));
	jdff dff_A_q6da7xD82_0(.dout(w_dff_A_x6zoRZYk4_0),.din(w_dff_A_q6da7xD82_0),.clk(gclk));
	jdff dff_A_x6zoRZYk4_0(.dout(w_dff_A_qVpcj7jv5_0),.din(w_dff_A_x6zoRZYk4_0),.clk(gclk));
	jdff dff_A_qVpcj7jv5_0(.dout(w_dff_A_6WeRIl7A2_0),.din(w_dff_A_qVpcj7jv5_0),.clk(gclk));
	jdff dff_A_6WeRIl7A2_0(.dout(w_dff_A_1KnrDZgR5_0),.din(w_dff_A_6WeRIl7A2_0),.clk(gclk));
	jdff dff_A_1KnrDZgR5_0(.dout(w_dff_A_zLGRwzUQ5_0),.din(w_dff_A_1KnrDZgR5_0),.clk(gclk));
	jdff dff_A_zLGRwzUQ5_0(.dout(w_dff_A_jHVo2UKZ5_0),.din(w_dff_A_zLGRwzUQ5_0),.clk(gclk));
	jdff dff_A_jHVo2UKZ5_0(.dout(w_dff_A_m1zYb7NW7_0),.din(w_dff_A_jHVo2UKZ5_0),.clk(gclk));
	jdff dff_A_m1zYb7NW7_0(.dout(w_dff_A_9UOwby586_0),.din(w_dff_A_m1zYb7NW7_0),.clk(gclk));
	jdff dff_A_9UOwby586_0(.dout(w_dff_A_k0PgebVk0_0),.din(w_dff_A_9UOwby586_0),.clk(gclk));
	jdff dff_A_k0PgebVk0_0(.dout(w_dff_A_OfHSRyVS1_0),.din(w_dff_A_k0PgebVk0_0),.clk(gclk));
	jdff dff_A_OfHSRyVS1_0(.dout(w_dff_A_F4I6rUl25_0),.din(w_dff_A_OfHSRyVS1_0),.clk(gclk));
	jdff dff_A_F4I6rUl25_0(.dout(w_dff_A_xwxd4ajW3_0),.din(w_dff_A_F4I6rUl25_0),.clk(gclk));
	jdff dff_A_xwxd4ajW3_0(.dout(w_dff_A_XEhTiZOz8_0),.din(w_dff_A_xwxd4ajW3_0),.clk(gclk));
	jdff dff_A_XEhTiZOz8_0(.dout(w_dff_A_xENpLPdo8_0),.din(w_dff_A_XEhTiZOz8_0),.clk(gclk));
	jdff dff_A_xENpLPdo8_0(.dout(w_dff_A_mXdx3Ypa7_0),.din(w_dff_A_xENpLPdo8_0),.clk(gclk));
	jdff dff_A_mXdx3Ypa7_0(.dout(f76),.din(w_dff_A_mXdx3Ypa7_0),.clk(gclk));
	jdff dff_A_RlfpDKF12_2(.dout(w_dff_A_4DonYcxZ2_0),.din(w_dff_A_RlfpDKF12_2),.clk(gclk));
	jdff dff_A_4DonYcxZ2_0(.dout(w_dff_A_B8HDxOQy5_0),.din(w_dff_A_4DonYcxZ2_0),.clk(gclk));
	jdff dff_A_B8HDxOQy5_0(.dout(w_dff_A_vdCQwJgC2_0),.din(w_dff_A_B8HDxOQy5_0),.clk(gclk));
	jdff dff_A_vdCQwJgC2_0(.dout(w_dff_A_vA1ZdwEd9_0),.din(w_dff_A_vdCQwJgC2_0),.clk(gclk));
	jdff dff_A_vA1ZdwEd9_0(.dout(w_dff_A_ARC4LZsm0_0),.din(w_dff_A_vA1ZdwEd9_0),.clk(gclk));
	jdff dff_A_ARC4LZsm0_0(.dout(w_dff_A_mWnDcfIB9_0),.din(w_dff_A_ARC4LZsm0_0),.clk(gclk));
	jdff dff_A_mWnDcfIB9_0(.dout(w_dff_A_ypgRplGv0_0),.din(w_dff_A_mWnDcfIB9_0),.clk(gclk));
	jdff dff_A_ypgRplGv0_0(.dout(w_dff_A_lsYs4WQt0_0),.din(w_dff_A_ypgRplGv0_0),.clk(gclk));
	jdff dff_A_lsYs4WQt0_0(.dout(w_dff_A_nnz5RsiZ8_0),.din(w_dff_A_lsYs4WQt0_0),.clk(gclk));
	jdff dff_A_nnz5RsiZ8_0(.dout(w_dff_A_giFPkiTO9_0),.din(w_dff_A_nnz5RsiZ8_0),.clk(gclk));
	jdff dff_A_giFPkiTO9_0(.dout(w_dff_A_SXJ0q3Ks3_0),.din(w_dff_A_giFPkiTO9_0),.clk(gclk));
	jdff dff_A_SXJ0q3Ks3_0(.dout(w_dff_A_3LmmaxXn8_0),.din(w_dff_A_SXJ0q3Ks3_0),.clk(gclk));
	jdff dff_A_3LmmaxXn8_0(.dout(w_dff_A_LtTDJPZR2_0),.din(w_dff_A_3LmmaxXn8_0),.clk(gclk));
	jdff dff_A_LtTDJPZR2_0(.dout(w_dff_A_foT4pxeZ4_0),.din(w_dff_A_LtTDJPZR2_0),.clk(gclk));
	jdff dff_A_foT4pxeZ4_0(.dout(w_dff_A_53QzjAf81_0),.din(w_dff_A_foT4pxeZ4_0),.clk(gclk));
	jdff dff_A_53QzjAf81_0(.dout(w_dff_A_ATpHjgT78_0),.din(w_dff_A_53QzjAf81_0),.clk(gclk));
	jdff dff_A_ATpHjgT78_0(.dout(w_dff_A_e0VT6QzL4_0),.din(w_dff_A_ATpHjgT78_0),.clk(gclk));
	jdff dff_A_e0VT6QzL4_0(.dout(w_dff_A_TWdJP5VH8_0),.din(w_dff_A_e0VT6QzL4_0),.clk(gclk));
	jdff dff_A_TWdJP5VH8_0(.dout(w_dff_A_q6F8wKw01_0),.din(w_dff_A_TWdJP5VH8_0),.clk(gclk));
	jdff dff_A_q6F8wKw01_0(.dout(w_dff_A_SpF0upsw2_0),.din(w_dff_A_q6F8wKw01_0),.clk(gclk));
	jdff dff_A_SpF0upsw2_0(.dout(w_dff_A_YBnZHitN9_0),.din(w_dff_A_SpF0upsw2_0),.clk(gclk));
	jdff dff_A_YBnZHitN9_0(.dout(w_dff_A_jUQBAWXz9_0),.din(w_dff_A_YBnZHitN9_0),.clk(gclk));
	jdff dff_A_jUQBAWXz9_0(.dout(w_dff_A_ecF1bpiO2_0),.din(w_dff_A_jUQBAWXz9_0),.clk(gclk));
	jdff dff_A_ecF1bpiO2_0(.dout(w_dff_A_cwxLrvwG9_0),.din(w_dff_A_ecF1bpiO2_0),.clk(gclk));
	jdff dff_A_cwxLrvwG9_0(.dout(w_dff_A_3Kv7FAwT0_0),.din(w_dff_A_cwxLrvwG9_0),.clk(gclk));
	jdff dff_A_3Kv7FAwT0_0(.dout(w_dff_A_MBDL2fvX3_0),.din(w_dff_A_3Kv7FAwT0_0),.clk(gclk));
	jdff dff_A_MBDL2fvX3_0(.dout(w_dff_A_S8ebt1Q11_0),.din(w_dff_A_MBDL2fvX3_0),.clk(gclk));
	jdff dff_A_S8ebt1Q11_0(.dout(w_dff_A_8fdtYeUp9_0),.din(w_dff_A_S8ebt1Q11_0),.clk(gclk));
	jdff dff_A_8fdtYeUp9_0(.dout(w_dff_A_mjXGhLxS5_0),.din(w_dff_A_8fdtYeUp9_0),.clk(gclk));
	jdff dff_A_mjXGhLxS5_0(.dout(w_dff_A_cmY9OMeK1_0),.din(w_dff_A_mjXGhLxS5_0),.clk(gclk));
	jdff dff_A_cmY9OMeK1_0(.dout(w_dff_A_izxOmPK24_0),.din(w_dff_A_cmY9OMeK1_0),.clk(gclk));
	jdff dff_A_izxOmPK24_0(.dout(w_dff_A_VBE13euG9_0),.din(w_dff_A_izxOmPK24_0),.clk(gclk));
	jdff dff_A_VBE13euG9_0(.dout(w_dff_A_YmhU2R6U4_0),.din(w_dff_A_VBE13euG9_0),.clk(gclk));
	jdff dff_A_YmhU2R6U4_0(.dout(w_dff_A_uFiOsNo44_0),.din(w_dff_A_YmhU2R6U4_0),.clk(gclk));
	jdff dff_A_uFiOsNo44_0(.dout(w_dff_A_zRjKlspb3_0),.din(w_dff_A_uFiOsNo44_0),.clk(gclk));
	jdff dff_A_zRjKlspb3_0(.dout(w_dff_A_hFvNIyOM3_0),.din(w_dff_A_zRjKlspb3_0),.clk(gclk));
	jdff dff_A_hFvNIyOM3_0(.dout(w_dff_A_kduNNEDK6_0),.din(w_dff_A_hFvNIyOM3_0),.clk(gclk));
	jdff dff_A_kduNNEDK6_0(.dout(w_dff_A_wCA7ujOc8_0),.din(w_dff_A_kduNNEDK6_0),.clk(gclk));
	jdff dff_A_wCA7ujOc8_0(.dout(w_dff_A_XyI67h5D6_0),.din(w_dff_A_wCA7ujOc8_0),.clk(gclk));
	jdff dff_A_XyI67h5D6_0(.dout(w_dff_A_N1xKqrTB1_0),.din(w_dff_A_XyI67h5D6_0),.clk(gclk));
	jdff dff_A_N1xKqrTB1_0(.dout(w_dff_A_OaeHKZhR1_0),.din(w_dff_A_N1xKqrTB1_0),.clk(gclk));
	jdff dff_A_OaeHKZhR1_0(.dout(w_dff_A_VqOlsUEJ2_0),.din(w_dff_A_OaeHKZhR1_0),.clk(gclk));
	jdff dff_A_VqOlsUEJ2_0(.dout(w_dff_A_Wt42TrZY5_0),.din(w_dff_A_VqOlsUEJ2_0),.clk(gclk));
	jdff dff_A_Wt42TrZY5_0(.dout(w_dff_A_cD2vn7133_0),.din(w_dff_A_Wt42TrZY5_0),.clk(gclk));
	jdff dff_A_cD2vn7133_0(.dout(w_dff_A_kINq8yqh2_0),.din(w_dff_A_cD2vn7133_0),.clk(gclk));
	jdff dff_A_kINq8yqh2_0(.dout(w_dff_A_QSEBN0SL5_0),.din(w_dff_A_kINq8yqh2_0),.clk(gclk));
	jdff dff_A_QSEBN0SL5_0(.dout(w_dff_A_l8H9QYxj0_0),.din(w_dff_A_QSEBN0SL5_0),.clk(gclk));
	jdff dff_A_l8H9QYxj0_0(.dout(w_dff_A_XD0GEFeW7_0),.din(w_dff_A_l8H9QYxj0_0),.clk(gclk));
	jdff dff_A_XD0GEFeW7_0(.dout(w_dff_A_OxCjHqpa7_0),.din(w_dff_A_XD0GEFeW7_0),.clk(gclk));
	jdff dff_A_OxCjHqpa7_0(.dout(f77),.din(w_dff_A_OxCjHqpa7_0),.clk(gclk));
	jdff dff_A_yWmtd95Z9_2(.dout(w_dff_A_qkZtBiSq1_0),.din(w_dff_A_yWmtd95Z9_2),.clk(gclk));
	jdff dff_A_qkZtBiSq1_0(.dout(w_dff_A_tScFh3Kl2_0),.din(w_dff_A_qkZtBiSq1_0),.clk(gclk));
	jdff dff_A_tScFh3Kl2_0(.dout(w_dff_A_36M7cNzF5_0),.din(w_dff_A_tScFh3Kl2_0),.clk(gclk));
	jdff dff_A_36M7cNzF5_0(.dout(w_dff_A_CndEV1K92_0),.din(w_dff_A_36M7cNzF5_0),.clk(gclk));
	jdff dff_A_CndEV1K92_0(.dout(w_dff_A_0h25dN1D6_0),.din(w_dff_A_CndEV1K92_0),.clk(gclk));
	jdff dff_A_0h25dN1D6_0(.dout(w_dff_A_oHXhD8j22_0),.din(w_dff_A_0h25dN1D6_0),.clk(gclk));
	jdff dff_A_oHXhD8j22_0(.dout(w_dff_A_bHuRnmKC2_0),.din(w_dff_A_oHXhD8j22_0),.clk(gclk));
	jdff dff_A_bHuRnmKC2_0(.dout(w_dff_A_F3vpQvgn6_0),.din(w_dff_A_bHuRnmKC2_0),.clk(gclk));
	jdff dff_A_F3vpQvgn6_0(.dout(w_dff_A_mZHBLTom4_0),.din(w_dff_A_F3vpQvgn6_0),.clk(gclk));
	jdff dff_A_mZHBLTom4_0(.dout(w_dff_A_etzstDjs6_0),.din(w_dff_A_mZHBLTom4_0),.clk(gclk));
	jdff dff_A_etzstDjs6_0(.dout(w_dff_A_AyGB1ZTc0_0),.din(w_dff_A_etzstDjs6_0),.clk(gclk));
	jdff dff_A_AyGB1ZTc0_0(.dout(w_dff_A_SJUkpxY93_0),.din(w_dff_A_AyGB1ZTc0_0),.clk(gclk));
	jdff dff_A_SJUkpxY93_0(.dout(w_dff_A_mP6XtOfq4_0),.din(w_dff_A_SJUkpxY93_0),.clk(gclk));
	jdff dff_A_mP6XtOfq4_0(.dout(w_dff_A_zfvjm2bz1_0),.din(w_dff_A_mP6XtOfq4_0),.clk(gclk));
	jdff dff_A_zfvjm2bz1_0(.dout(w_dff_A_YPoHV4Kg3_0),.din(w_dff_A_zfvjm2bz1_0),.clk(gclk));
	jdff dff_A_YPoHV4Kg3_0(.dout(w_dff_A_PVCzV6Ho8_0),.din(w_dff_A_YPoHV4Kg3_0),.clk(gclk));
	jdff dff_A_PVCzV6Ho8_0(.dout(w_dff_A_WmuU9RFK7_0),.din(w_dff_A_PVCzV6Ho8_0),.clk(gclk));
	jdff dff_A_WmuU9RFK7_0(.dout(w_dff_A_pMmWgtmU4_0),.din(w_dff_A_WmuU9RFK7_0),.clk(gclk));
	jdff dff_A_pMmWgtmU4_0(.dout(w_dff_A_RdlQZcB12_0),.din(w_dff_A_pMmWgtmU4_0),.clk(gclk));
	jdff dff_A_RdlQZcB12_0(.dout(w_dff_A_ggR422Dh2_0),.din(w_dff_A_RdlQZcB12_0),.clk(gclk));
	jdff dff_A_ggR422Dh2_0(.dout(w_dff_A_ncWh2HX84_0),.din(w_dff_A_ggR422Dh2_0),.clk(gclk));
	jdff dff_A_ncWh2HX84_0(.dout(w_dff_A_l70S9Sxu5_0),.din(w_dff_A_ncWh2HX84_0),.clk(gclk));
	jdff dff_A_l70S9Sxu5_0(.dout(w_dff_A_23pVAkUT1_0),.din(w_dff_A_l70S9Sxu5_0),.clk(gclk));
	jdff dff_A_23pVAkUT1_0(.dout(w_dff_A_ib1426oH9_0),.din(w_dff_A_23pVAkUT1_0),.clk(gclk));
	jdff dff_A_ib1426oH9_0(.dout(w_dff_A_b1EAwoEw3_0),.din(w_dff_A_ib1426oH9_0),.clk(gclk));
	jdff dff_A_b1EAwoEw3_0(.dout(w_dff_A_2zek97ag8_0),.din(w_dff_A_b1EAwoEw3_0),.clk(gclk));
	jdff dff_A_2zek97ag8_0(.dout(w_dff_A_oWryYxg27_0),.din(w_dff_A_2zek97ag8_0),.clk(gclk));
	jdff dff_A_oWryYxg27_0(.dout(w_dff_A_AXf38r8r6_0),.din(w_dff_A_oWryYxg27_0),.clk(gclk));
	jdff dff_A_AXf38r8r6_0(.dout(w_dff_A_RQCD9r8D8_0),.din(w_dff_A_AXf38r8r6_0),.clk(gclk));
	jdff dff_A_RQCD9r8D8_0(.dout(w_dff_A_iy1CD8ki6_0),.din(w_dff_A_RQCD9r8D8_0),.clk(gclk));
	jdff dff_A_iy1CD8ki6_0(.dout(w_dff_A_BZ7rYHzE1_0),.din(w_dff_A_iy1CD8ki6_0),.clk(gclk));
	jdff dff_A_BZ7rYHzE1_0(.dout(w_dff_A_W74HFkOY5_0),.din(w_dff_A_BZ7rYHzE1_0),.clk(gclk));
	jdff dff_A_W74HFkOY5_0(.dout(w_dff_A_zdvoRqev6_0),.din(w_dff_A_W74HFkOY5_0),.clk(gclk));
	jdff dff_A_zdvoRqev6_0(.dout(w_dff_A_hOMlBEIg4_0),.din(w_dff_A_zdvoRqev6_0),.clk(gclk));
	jdff dff_A_hOMlBEIg4_0(.dout(w_dff_A_PziKTnu00_0),.din(w_dff_A_hOMlBEIg4_0),.clk(gclk));
	jdff dff_A_PziKTnu00_0(.dout(w_dff_A_NcUkuUVK3_0),.din(w_dff_A_PziKTnu00_0),.clk(gclk));
	jdff dff_A_NcUkuUVK3_0(.dout(w_dff_A_KIpAsP4F0_0),.din(w_dff_A_NcUkuUVK3_0),.clk(gclk));
	jdff dff_A_KIpAsP4F0_0(.dout(w_dff_A_1PBDSoX25_0),.din(w_dff_A_KIpAsP4F0_0),.clk(gclk));
	jdff dff_A_1PBDSoX25_0(.dout(w_dff_A_F8AbN9jj0_0),.din(w_dff_A_1PBDSoX25_0),.clk(gclk));
	jdff dff_A_F8AbN9jj0_0(.dout(w_dff_A_bCu22zD62_0),.din(w_dff_A_F8AbN9jj0_0),.clk(gclk));
	jdff dff_A_bCu22zD62_0(.dout(w_dff_A_7C6icvPk2_0),.din(w_dff_A_bCu22zD62_0),.clk(gclk));
	jdff dff_A_7C6icvPk2_0(.dout(w_dff_A_jMSl0l025_0),.din(w_dff_A_7C6icvPk2_0),.clk(gclk));
	jdff dff_A_jMSl0l025_0(.dout(w_dff_A_FVKZY5wV7_0),.din(w_dff_A_jMSl0l025_0),.clk(gclk));
	jdff dff_A_FVKZY5wV7_0(.dout(w_dff_A_x7UftJps5_0),.din(w_dff_A_FVKZY5wV7_0),.clk(gclk));
	jdff dff_A_x7UftJps5_0(.dout(w_dff_A_MjHkPadH7_0),.din(w_dff_A_x7UftJps5_0),.clk(gclk));
	jdff dff_A_MjHkPadH7_0(.dout(w_dff_A_mgVfQPcp4_0),.din(w_dff_A_MjHkPadH7_0),.clk(gclk));
	jdff dff_A_mgVfQPcp4_0(.dout(w_dff_A_L3MUWpVP2_0),.din(w_dff_A_mgVfQPcp4_0),.clk(gclk));
	jdff dff_A_L3MUWpVP2_0(.dout(w_dff_A_ESH7nihC7_0),.din(w_dff_A_L3MUWpVP2_0),.clk(gclk));
	jdff dff_A_ESH7nihC7_0(.dout(f78),.din(w_dff_A_ESH7nihC7_0),.clk(gclk));
	jdff dff_A_iULoKlkx1_2(.dout(w_dff_A_hRb1WDEa6_0),.din(w_dff_A_iULoKlkx1_2),.clk(gclk));
	jdff dff_A_hRb1WDEa6_0(.dout(w_dff_A_Lda5KRtg5_0),.din(w_dff_A_hRb1WDEa6_0),.clk(gclk));
	jdff dff_A_Lda5KRtg5_0(.dout(w_dff_A_bFIitHTF7_0),.din(w_dff_A_Lda5KRtg5_0),.clk(gclk));
	jdff dff_A_bFIitHTF7_0(.dout(w_dff_A_XeOhAS495_0),.din(w_dff_A_bFIitHTF7_0),.clk(gclk));
	jdff dff_A_XeOhAS495_0(.dout(w_dff_A_EIGSAZnU0_0),.din(w_dff_A_XeOhAS495_0),.clk(gclk));
	jdff dff_A_EIGSAZnU0_0(.dout(w_dff_A_suP6yMeK3_0),.din(w_dff_A_EIGSAZnU0_0),.clk(gclk));
	jdff dff_A_suP6yMeK3_0(.dout(w_dff_A_eVjXcTaJ5_0),.din(w_dff_A_suP6yMeK3_0),.clk(gclk));
	jdff dff_A_eVjXcTaJ5_0(.dout(w_dff_A_B2RowLKo8_0),.din(w_dff_A_eVjXcTaJ5_0),.clk(gclk));
	jdff dff_A_B2RowLKo8_0(.dout(w_dff_A_u5SecGSH2_0),.din(w_dff_A_B2RowLKo8_0),.clk(gclk));
	jdff dff_A_u5SecGSH2_0(.dout(w_dff_A_F8FMi8VD0_0),.din(w_dff_A_u5SecGSH2_0),.clk(gclk));
	jdff dff_A_F8FMi8VD0_0(.dout(w_dff_A_IuH4HrD66_0),.din(w_dff_A_F8FMi8VD0_0),.clk(gclk));
	jdff dff_A_IuH4HrD66_0(.dout(w_dff_A_MXfMiRkz0_0),.din(w_dff_A_IuH4HrD66_0),.clk(gclk));
	jdff dff_A_MXfMiRkz0_0(.dout(w_dff_A_KLf448jv9_0),.din(w_dff_A_MXfMiRkz0_0),.clk(gclk));
	jdff dff_A_KLf448jv9_0(.dout(w_dff_A_w2DZAeCL5_0),.din(w_dff_A_KLf448jv9_0),.clk(gclk));
	jdff dff_A_w2DZAeCL5_0(.dout(w_dff_A_qUQu7PYp3_0),.din(w_dff_A_w2DZAeCL5_0),.clk(gclk));
	jdff dff_A_qUQu7PYp3_0(.dout(w_dff_A_DW3tUMo90_0),.din(w_dff_A_qUQu7PYp3_0),.clk(gclk));
	jdff dff_A_DW3tUMo90_0(.dout(w_dff_A_ml40Ebtd9_0),.din(w_dff_A_DW3tUMo90_0),.clk(gclk));
	jdff dff_A_ml40Ebtd9_0(.dout(w_dff_A_2q0z7P6E9_0),.din(w_dff_A_ml40Ebtd9_0),.clk(gclk));
	jdff dff_A_2q0z7P6E9_0(.dout(w_dff_A_euZLH25e8_0),.din(w_dff_A_2q0z7P6E9_0),.clk(gclk));
	jdff dff_A_euZLH25e8_0(.dout(w_dff_A_PZ7SHKic2_0),.din(w_dff_A_euZLH25e8_0),.clk(gclk));
	jdff dff_A_PZ7SHKic2_0(.dout(w_dff_A_WJch9ZpO9_0),.din(w_dff_A_PZ7SHKic2_0),.clk(gclk));
	jdff dff_A_WJch9ZpO9_0(.dout(w_dff_A_quIVjniU2_0),.din(w_dff_A_WJch9ZpO9_0),.clk(gclk));
	jdff dff_A_quIVjniU2_0(.dout(w_dff_A_M7Q6Agcq9_0),.din(w_dff_A_quIVjniU2_0),.clk(gclk));
	jdff dff_A_M7Q6Agcq9_0(.dout(w_dff_A_7oMQAG7l5_0),.din(w_dff_A_M7Q6Agcq9_0),.clk(gclk));
	jdff dff_A_7oMQAG7l5_0(.dout(w_dff_A_dzsqJTU21_0),.din(w_dff_A_7oMQAG7l5_0),.clk(gclk));
	jdff dff_A_dzsqJTU21_0(.dout(w_dff_A_IkcQABtj1_0),.din(w_dff_A_dzsqJTU21_0),.clk(gclk));
	jdff dff_A_IkcQABtj1_0(.dout(w_dff_A_GPFCbRyC3_0),.din(w_dff_A_IkcQABtj1_0),.clk(gclk));
	jdff dff_A_GPFCbRyC3_0(.dout(w_dff_A_SX7vW9ct8_0),.din(w_dff_A_GPFCbRyC3_0),.clk(gclk));
	jdff dff_A_SX7vW9ct8_0(.dout(w_dff_A_0LazYeen7_0),.din(w_dff_A_SX7vW9ct8_0),.clk(gclk));
	jdff dff_A_0LazYeen7_0(.dout(w_dff_A_BoEdLu2e2_0),.din(w_dff_A_0LazYeen7_0),.clk(gclk));
	jdff dff_A_BoEdLu2e2_0(.dout(w_dff_A_r2SqBUtD8_0),.din(w_dff_A_BoEdLu2e2_0),.clk(gclk));
	jdff dff_A_r2SqBUtD8_0(.dout(w_dff_A_0k217cT47_0),.din(w_dff_A_r2SqBUtD8_0),.clk(gclk));
	jdff dff_A_0k217cT47_0(.dout(w_dff_A_jd6fyX7m2_0),.din(w_dff_A_0k217cT47_0),.clk(gclk));
	jdff dff_A_jd6fyX7m2_0(.dout(w_dff_A_oDXlhhnW8_0),.din(w_dff_A_jd6fyX7m2_0),.clk(gclk));
	jdff dff_A_oDXlhhnW8_0(.dout(w_dff_A_VzuZuzZi1_0),.din(w_dff_A_oDXlhhnW8_0),.clk(gclk));
	jdff dff_A_VzuZuzZi1_0(.dout(w_dff_A_fG4EvSUN6_0),.din(w_dff_A_VzuZuzZi1_0),.clk(gclk));
	jdff dff_A_fG4EvSUN6_0(.dout(w_dff_A_IJnyghi77_0),.din(w_dff_A_fG4EvSUN6_0),.clk(gclk));
	jdff dff_A_IJnyghi77_0(.dout(w_dff_A_rdCuDiAg3_0),.din(w_dff_A_IJnyghi77_0),.clk(gclk));
	jdff dff_A_rdCuDiAg3_0(.dout(w_dff_A_wUqX7ldH1_0),.din(w_dff_A_rdCuDiAg3_0),.clk(gclk));
	jdff dff_A_wUqX7ldH1_0(.dout(w_dff_A_q1rZZC0K4_0),.din(w_dff_A_wUqX7ldH1_0),.clk(gclk));
	jdff dff_A_q1rZZC0K4_0(.dout(w_dff_A_EHbPQLf29_0),.din(w_dff_A_q1rZZC0K4_0),.clk(gclk));
	jdff dff_A_EHbPQLf29_0(.dout(w_dff_A_oBp2Hrva8_0),.din(w_dff_A_EHbPQLf29_0),.clk(gclk));
	jdff dff_A_oBp2Hrva8_0(.dout(w_dff_A_0glMPIVS2_0),.din(w_dff_A_oBp2Hrva8_0),.clk(gclk));
	jdff dff_A_0glMPIVS2_0(.dout(w_dff_A_a96g5GQv4_0),.din(w_dff_A_0glMPIVS2_0),.clk(gclk));
	jdff dff_A_a96g5GQv4_0(.dout(w_dff_A_8rK7WVdA8_0),.din(w_dff_A_a96g5GQv4_0),.clk(gclk));
	jdff dff_A_8rK7WVdA8_0(.dout(w_dff_A_Td3y2RKm7_0),.din(w_dff_A_8rK7WVdA8_0),.clk(gclk));
	jdff dff_A_Td3y2RKm7_0(.dout(w_dff_A_8gHFPLMH2_0),.din(w_dff_A_Td3y2RKm7_0),.clk(gclk));
	jdff dff_A_8gHFPLMH2_0(.dout(f79),.din(w_dff_A_8gHFPLMH2_0),.clk(gclk));
	jdff dff_A_E95bjTHE6_2(.dout(w_dff_A_EkTlbwSF6_0),.din(w_dff_A_E95bjTHE6_2),.clk(gclk));
	jdff dff_A_EkTlbwSF6_0(.dout(w_dff_A_VJtmhJed3_0),.din(w_dff_A_EkTlbwSF6_0),.clk(gclk));
	jdff dff_A_VJtmhJed3_0(.dout(w_dff_A_ory6Rcro9_0),.din(w_dff_A_VJtmhJed3_0),.clk(gclk));
	jdff dff_A_ory6Rcro9_0(.dout(w_dff_A_789X5lqI1_0),.din(w_dff_A_ory6Rcro9_0),.clk(gclk));
	jdff dff_A_789X5lqI1_0(.dout(w_dff_A_AWe4MnpT8_0),.din(w_dff_A_789X5lqI1_0),.clk(gclk));
	jdff dff_A_AWe4MnpT8_0(.dout(w_dff_A_OFWlbXqg9_0),.din(w_dff_A_AWe4MnpT8_0),.clk(gclk));
	jdff dff_A_OFWlbXqg9_0(.dout(w_dff_A_1I04ukaw6_0),.din(w_dff_A_OFWlbXqg9_0),.clk(gclk));
	jdff dff_A_1I04ukaw6_0(.dout(w_dff_A_hjd4ZPIZ3_0),.din(w_dff_A_1I04ukaw6_0),.clk(gclk));
	jdff dff_A_hjd4ZPIZ3_0(.dout(w_dff_A_bPECUQSg4_0),.din(w_dff_A_hjd4ZPIZ3_0),.clk(gclk));
	jdff dff_A_bPECUQSg4_0(.dout(w_dff_A_tANPOkyx9_0),.din(w_dff_A_bPECUQSg4_0),.clk(gclk));
	jdff dff_A_tANPOkyx9_0(.dout(w_dff_A_5LxVsuub5_0),.din(w_dff_A_tANPOkyx9_0),.clk(gclk));
	jdff dff_A_5LxVsuub5_0(.dout(w_dff_A_734NZw6D6_0),.din(w_dff_A_5LxVsuub5_0),.clk(gclk));
	jdff dff_A_734NZw6D6_0(.dout(w_dff_A_GuJyUhbp0_0),.din(w_dff_A_734NZw6D6_0),.clk(gclk));
	jdff dff_A_GuJyUhbp0_0(.dout(w_dff_A_XJkQ9pqk1_0),.din(w_dff_A_GuJyUhbp0_0),.clk(gclk));
	jdff dff_A_XJkQ9pqk1_0(.dout(w_dff_A_EmnbvvHE2_0),.din(w_dff_A_XJkQ9pqk1_0),.clk(gclk));
	jdff dff_A_EmnbvvHE2_0(.dout(w_dff_A_X5g9KCer4_0),.din(w_dff_A_EmnbvvHE2_0),.clk(gclk));
	jdff dff_A_X5g9KCer4_0(.dout(w_dff_A_Q1MI5oLg1_0),.din(w_dff_A_X5g9KCer4_0),.clk(gclk));
	jdff dff_A_Q1MI5oLg1_0(.dout(w_dff_A_u5SGxHBw3_0),.din(w_dff_A_Q1MI5oLg1_0),.clk(gclk));
	jdff dff_A_u5SGxHBw3_0(.dout(w_dff_A_rrICQaGk4_0),.din(w_dff_A_u5SGxHBw3_0),.clk(gclk));
	jdff dff_A_rrICQaGk4_0(.dout(w_dff_A_pGcTZ0tE1_0),.din(w_dff_A_rrICQaGk4_0),.clk(gclk));
	jdff dff_A_pGcTZ0tE1_0(.dout(w_dff_A_7BWyScQ28_0),.din(w_dff_A_pGcTZ0tE1_0),.clk(gclk));
	jdff dff_A_7BWyScQ28_0(.dout(w_dff_A_O8l17WgZ1_0),.din(w_dff_A_7BWyScQ28_0),.clk(gclk));
	jdff dff_A_O8l17WgZ1_0(.dout(w_dff_A_153vyNHY4_0),.din(w_dff_A_O8l17WgZ1_0),.clk(gclk));
	jdff dff_A_153vyNHY4_0(.dout(w_dff_A_wmySegux3_0),.din(w_dff_A_153vyNHY4_0),.clk(gclk));
	jdff dff_A_wmySegux3_0(.dout(w_dff_A_HI40fgjV3_0),.din(w_dff_A_wmySegux3_0),.clk(gclk));
	jdff dff_A_HI40fgjV3_0(.dout(w_dff_A_1SrDlBC40_0),.din(w_dff_A_HI40fgjV3_0),.clk(gclk));
	jdff dff_A_1SrDlBC40_0(.dout(w_dff_A_IQzhHR6F4_0),.din(w_dff_A_1SrDlBC40_0),.clk(gclk));
	jdff dff_A_IQzhHR6F4_0(.dout(w_dff_A_BkzKRszD2_0),.din(w_dff_A_IQzhHR6F4_0),.clk(gclk));
	jdff dff_A_BkzKRszD2_0(.dout(w_dff_A_h04rrvJB1_0),.din(w_dff_A_BkzKRszD2_0),.clk(gclk));
	jdff dff_A_h04rrvJB1_0(.dout(w_dff_A_t0tkoMpx9_0),.din(w_dff_A_h04rrvJB1_0),.clk(gclk));
	jdff dff_A_t0tkoMpx9_0(.dout(w_dff_A_bZQhJkMe0_0),.din(w_dff_A_t0tkoMpx9_0),.clk(gclk));
	jdff dff_A_bZQhJkMe0_0(.dout(w_dff_A_zaiFWFK59_0),.din(w_dff_A_bZQhJkMe0_0),.clk(gclk));
	jdff dff_A_zaiFWFK59_0(.dout(w_dff_A_3GXMC9mH3_0),.din(w_dff_A_zaiFWFK59_0),.clk(gclk));
	jdff dff_A_3GXMC9mH3_0(.dout(w_dff_A_aiQTVfsj5_0),.din(w_dff_A_3GXMC9mH3_0),.clk(gclk));
	jdff dff_A_aiQTVfsj5_0(.dout(w_dff_A_fvxgQ0L95_0),.din(w_dff_A_aiQTVfsj5_0),.clk(gclk));
	jdff dff_A_fvxgQ0L95_0(.dout(w_dff_A_2IzbuGBO9_0),.din(w_dff_A_fvxgQ0L95_0),.clk(gclk));
	jdff dff_A_2IzbuGBO9_0(.dout(w_dff_A_gzYSSEkJ2_0),.din(w_dff_A_2IzbuGBO9_0),.clk(gclk));
	jdff dff_A_gzYSSEkJ2_0(.dout(w_dff_A_Y6FuboB72_0),.din(w_dff_A_gzYSSEkJ2_0),.clk(gclk));
	jdff dff_A_Y6FuboB72_0(.dout(w_dff_A_YLFp524t3_0),.din(w_dff_A_Y6FuboB72_0),.clk(gclk));
	jdff dff_A_YLFp524t3_0(.dout(w_dff_A_deaxy2T96_0),.din(w_dff_A_YLFp524t3_0),.clk(gclk));
	jdff dff_A_deaxy2T96_0(.dout(w_dff_A_peUlOvJM1_0),.din(w_dff_A_deaxy2T96_0),.clk(gclk));
	jdff dff_A_peUlOvJM1_0(.dout(w_dff_A_lB3oYaCR8_0),.din(w_dff_A_peUlOvJM1_0),.clk(gclk));
	jdff dff_A_lB3oYaCR8_0(.dout(w_dff_A_vWLF5Wq77_0),.din(w_dff_A_lB3oYaCR8_0),.clk(gclk));
	jdff dff_A_vWLF5Wq77_0(.dout(w_dff_A_zmnA5sqz5_0),.din(w_dff_A_vWLF5Wq77_0),.clk(gclk));
	jdff dff_A_zmnA5sqz5_0(.dout(w_dff_A_AZUNBJU43_0),.din(w_dff_A_zmnA5sqz5_0),.clk(gclk));
	jdff dff_A_AZUNBJU43_0(.dout(w_dff_A_JbtFcLIb4_0),.din(w_dff_A_AZUNBJU43_0),.clk(gclk));
	jdff dff_A_JbtFcLIb4_0(.dout(f80),.din(w_dff_A_JbtFcLIb4_0),.clk(gclk));
	jdff dff_A_5ajlcE7V4_2(.dout(w_dff_A_yrq8RRxb6_0),.din(w_dff_A_5ajlcE7V4_2),.clk(gclk));
	jdff dff_A_yrq8RRxb6_0(.dout(w_dff_A_SRMDKckD6_0),.din(w_dff_A_yrq8RRxb6_0),.clk(gclk));
	jdff dff_A_SRMDKckD6_0(.dout(w_dff_A_VrxVSJdl0_0),.din(w_dff_A_SRMDKckD6_0),.clk(gclk));
	jdff dff_A_VrxVSJdl0_0(.dout(w_dff_A_RlvhMH4m9_0),.din(w_dff_A_VrxVSJdl0_0),.clk(gclk));
	jdff dff_A_RlvhMH4m9_0(.dout(w_dff_A_10ixQL8w0_0),.din(w_dff_A_RlvhMH4m9_0),.clk(gclk));
	jdff dff_A_10ixQL8w0_0(.dout(w_dff_A_02uvXEfK9_0),.din(w_dff_A_10ixQL8w0_0),.clk(gclk));
	jdff dff_A_02uvXEfK9_0(.dout(w_dff_A_Y4iLZifS1_0),.din(w_dff_A_02uvXEfK9_0),.clk(gclk));
	jdff dff_A_Y4iLZifS1_0(.dout(w_dff_A_AKZN3ET33_0),.din(w_dff_A_Y4iLZifS1_0),.clk(gclk));
	jdff dff_A_AKZN3ET33_0(.dout(w_dff_A_L2vIkbfK1_0),.din(w_dff_A_AKZN3ET33_0),.clk(gclk));
	jdff dff_A_L2vIkbfK1_0(.dout(w_dff_A_AUzPE6SA3_0),.din(w_dff_A_L2vIkbfK1_0),.clk(gclk));
	jdff dff_A_AUzPE6SA3_0(.dout(w_dff_A_bGLFVMNg6_0),.din(w_dff_A_AUzPE6SA3_0),.clk(gclk));
	jdff dff_A_bGLFVMNg6_0(.dout(w_dff_A_ovTPSDu90_0),.din(w_dff_A_bGLFVMNg6_0),.clk(gclk));
	jdff dff_A_ovTPSDu90_0(.dout(w_dff_A_4jttJpBA9_0),.din(w_dff_A_ovTPSDu90_0),.clk(gclk));
	jdff dff_A_4jttJpBA9_0(.dout(w_dff_A_NDIwV7dc8_0),.din(w_dff_A_4jttJpBA9_0),.clk(gclk));
	jdff dff_A_NDIwV7dc8_0(.dout(w_dff_A_CZ6Mui0E3_0),.din(w_dff_A_NDIwV7dc8_0),.clk(gclk));
	jdff dff_A_CZ6Mui0E3_0(.dout(w_dff_A_Z3GL3A8L0_0),.din(w_dff_A_CZ6Mui0E3_0),.clk(gclk));
	jdff dff_A_Z3GL3A8L0_0(.dout(w_dff_A_1ojMFOxX6_0),.din(w_dff_A_Z3GL3A8L0_0),.clk(gclk));
	jdff dff_A_1ojMFOxX6_0(.dout(w_dff_A_CbEU7rhi9_0),.din(w_dff_A_1ojMFOxX6_0),.clk(gclk));
	jdff dff_A_CbEU7rhi9_0(.dout(w_dff_A_9v7iZBZt6_0),.din(w_dff_A_CbEU7rhi9_0),.clk(gclk));
	jdff dff_A_9v7iZBZt6_0(.dout(w_dff_A_ahTrYK8P6_0),.din(w_dff_A_9v7iZBZt6_0),.clk(gclk));
	jdff dff_A_ahTrYK8P6_0(.dout(w_dff_A_1ojEdrYW0_0),.din(w_dff_A_ahTrYK8P6_0),.clk(gclk));
	jdff dff_A_1ojEdrYW0_0(.dout(w_dff_A_eIiR2u5o9_0),.din(w_dff_A_1ojEdrYW0_0),.clk(gclk));
	jdff dff_A_eIiR2u5o9_0(.dout(w_dff_A_Z1HHw6HT0_0),.din(w_dff_A_eIiR2u5o9_0),.clk(gclk));
	jdff dff_A_Z1HHw6HT0_0(.dout(w_dff_A_0BLxCuJ03_0),.din(w_dff_A_Z1HHw6HT0_0),.clk(gclk));
	jdff dff_A_0BLxCuJ03_0(.dout(w_dff_A_2IaUoFT26_0),.din(w_dff_A_0BLxCuJ03_0),.clk(gclk));
	jdff dff_A_2IaUoFT26_0(.dout(w_dff_A_C1w00jop1_0),.din(w_dff_A_2IaUoFT26_0),.clk(gclk));
	jdff dff_A_C1w00jop1_0(.dout(w_dff_A_P0TcQm7r4_0),.din(w_dff_A_C1w00jop1_0),.clk(gclk));
	jdff dff_A_P0TcQm7r4_0(.dout(w_dff_A_MTh4EHZj9_0),.din(w_dff_A_P0TcQm7r4_0),.clk(gclk));
	jdff dff_A_MTh4EHZj9_0(.dout(w_dff_A_uNYNhFHg7_0),.din(w_dff_A_MTh4EHZj9_0),.clk(gclk));
	jdff dff_A_uNYNhFHg7_0(.dout(w_dff_A_8H2zzh131_0),.din(w_dff_A_uNYNhFHg7_0),.clk(gclk));
	jdff dff_A_8H2zzh131_0(.dout(w_dff_A_5HtWgcmt4_0),.din(w_dff_A_8H2zzh131_0),.clk(gclk));
	jdff dff_A_5HtWgcmt4_0(.dout(w_dff_A_KHt6XktR9_0),.din(w_dff_A_5HtWgcmt4_0),.clk(gclk));
	jdff dff_A_KHt6XktR9_0(.dout(w_dff_A_W1JBg2YO2_0),.din(w_dff_A_KHt6XktR9_0),.clk(gclk));
	jdff dff_A_W1JBg2YO2_0(.dout(w_dff_A_SCF40G4p1_0),.din(w_dff_A_W1JBg2YO2_0),.clk(gclk));
	jdff dff_A_SCF40G4p1_0(.dout(w_dff_A_Pmso16Wt4_0),.din(w_dff_A_SCF40G4p1_0),.clk(gclk));
	jdff dff_A_Pmso16Wt4_0(.dout(w_dff_A_iBITEoki8_0),.din(w_dff_A_Pmso16Wt4_0),.clk(gclk));
	jdff dff_A_iBITEoki8_0(.dout(w_dff_A_w9QRzCAq2_0),.din(w_dff_A_iBITEoki8_0),.clk(gclk));
	jdff dff_A_w9QRzCAq2_0(.dout(w_dff_A_AxUGuuMg0_0),.din(w_dff_A_w9QRzCAq2_0),.clk(gclk));
	jdff dff_A_AxUGuuMg0_0(.dout(w_dff_A_CeEVVqsP7_0),.din(w_dff_A_AxUGuuMg0_0),.clk(gclk));
	jdff dff_A_CeEVVqsP7_0(.dout(w_dff_A_JWbKkE1b5_0),.din(w_dff_A_CeEVVqsP7_0),.clk(gclk));
	jdff dff_A_JWbKkE1b5_0(.dout(w_dff_A_GY1PQSS14_0),.din(w_dff_A_JWbKkE1b5_0),.clk(gclk));
	jdff dff_A_GY1PQSS14_0(.dout(w_dff_A_peXopZp01_0),.din(w_dff_A_GY1PQSS14_0),.clk(gclk));
	jdff dff_A_peXopZp01_0(.dout(w_dff_A_CxEFWK3D9_0),.din(w_dff_A_peXopZp01_0),.clk(gclk));
	jdff dff_A_CxEFWK3D9_0(.dout(w_dff_A_ZXdXoEhP7_0),.din(w_dff_A_CxEFWK3D9_0),.clk(gclk));
	jdff dff_A_ZXdXoEhP7_0(.dout(w_dff_A_9DMIZN2c4_0),.din(w_dff_A_ZXdXoEhP7_0),.clk(gclk));
	jdff dff_A_9DMIZN2c4_0(.dout(f81),.din(w_dff_A_9DMIZN2c4_0),.clk(gclk));
	jdff dff_A_Xic2Adtu8_2(.dout(w_dff_A_ae3fN4sz7_0),.din(w_dff_A_Xic2Adtu8_2),.clk(gclk));
	jdff dff_A_ae3fN4sz7_0(.dout(w_dff_A_QH3nMiW09_0),.din(w_dff_A_ae3fN4sz7_0),.clk(gclk));
	jdff dff_A_QH3nMiW09_0(.dout(w_dff_A_8KTAWJsc8_0),.din(w_dff_A_QH3nMiW09_0),.clk(gclk));
	jdff dff_A_8KTAWJsc8_0(.dout(w_dff_A_pwhuY45Y9_0),.din(w_dff_A_8KTAWJsc8_0),.clk(gclk));
	jdff dff_A_pwhuY45Y9_0(.dout(w_dff_A_CTN0kwmC8_0),.din(w_dff_A_pwhuY45Y9_0),.clk(gclk));
	jdff dff_A_CTN0kwmC8_0(.dout(w_dff_A_puY2T0OV1_0),.din(w_dff_A_CTN0kwmC8_0),.clk(gclk));
	jdff dff_A_puY2T0OV1_0(.dout(w_dff_A_an8NgWan7_0),.din(w_dff_A_puY2T0OV1_0),.clk(gclk));
	jdff dff_A_an8NgWan7_0(.dout(w_dff_A_zX5ZeUkR1_0),.din(w_dff_A_an8NgWan7_0),.clk(gclk));
	jdff dff_A_zX5ZeUkR1_0(.dout(w_dff_A_E2iaVVUK0_0),.din(w_dff_A_zX5ZeUkR1_0),.clk(gclk));
	jdff dff_A_E2iaVVUK0_0(.dout(w_dff_A_ZuXgAFUx9_0),.din(w_dff_A_E2iaVVUK0_0),.clk(gclk));
	jdff dff_A_ZuXgAFUx9_0(.dout(w_dff_A_NGl7jE5l4_0),.din(w_dff_A_ZuXgAFUx9_0),.clk(gclk));
	jdff dff_A_NGl7jE5l4_0(.dout(w_dff_A_9gwTamw38_0),.din(w_dff_A_NGl7jE5l4_0),.clk(gclk));
	jdff dff_A_9gwTamw38_0(.dout(w_dff_A_j7WgJTx71_0),.din(w_dff_A_9gwTamw38_0),.clk(gclk));
	jdff dff_A_j7WgJTx71_0(.dout(w_dff_A_V65MCLsK6_0),.din(w_dff_A_j7WgJTx71_0),.clk(gclk));
	jdff dff_A_V65MCLsK6_0(.dout(w_dff_A_uSeQGyzD7_0),.din(w_dff_A_V65MCLsK6_0),.clk(gclk));
	jdff dff_A_uSeQGyzD7_0(.dout(w_dff_A_oLANuLxA6_0),.din(w_dff_A_uSeQGyzD7_0),.clk(gclk));
	jdff dff_A_oLANuLxA6_0(.dout(w_dff_A_kD0lhMUr7_0),.din(w_dff_A_oLANuLxA6_0),.clk(gclk));
	jdff dff_A_kD0lhMUr7_0(.dout(w_dff_A_psXX62it7_0),.din(w_dff_A_kD0lhMUr7_0),.clk(gclk));
	jdff dff_A_psXX62it7_0(.dout(w_dff_A_meDuEnw66_0),.din(w_dff_A_psXX62it7_0),.clk(gclk));
	jdff dff_A_meDuEnw66_0(.dout(w_dff_A_sLnJVsKA3_0),.din(w_dff_A_meDuEnw66_0),.clk(gclk));
	jdff dff_A_sLnJVsKA3_0(.dout(w_dff_A_QsLVnZK26_0),.din(w_dff_A_sLnJVsKA3_0),.clk(gclk));
	jdff dff_A_QsLVnZK26_0(.dout(w_dff_A_ZEWEmoHY3_0),.din(w_dff_A_QsLVnZK26_0),.clk(gclk));
	jdff dff_A_ZEWEmoHY3_0(.dout(w_dff_A_VkMBIxlN5_0),.din(w_dff_A_ZEWEmoHY3_0),.clk(gclk));
	jdff dff_A_VkMBIxlN5_0(.dout(w_dff_A_UNfluSTA0_0),.din(w_dff_A_VkMBIxlN5_0),.clk(gclk));
	jdff dff_A_UNfluSTA0_0(.dout(w_dff_A_qKZ87JSS6_0),.din(w_dff_A_UNfluSTA0_0),.clk(gclk));
	jdff dff_A_qKZ87JSS6_0(.dout(w_dff_A_3bZjeuQH4_0),.din(w_dff_A_qKZ87JSS6_0),.clk(gclk));
	jdff dff_A_3bZjeuQH4_0(.dout(w_dff_A_AWxnT9AG4_0),.din(w_dff_A_3bZjeuQH4_0),.clk(gclk));
	jdff dff_A_AWxnT9AG4_0(.dout(w_dff_A_6cvzohV45_0),.din(w_dff_A_AWxnT9AG4_0),.clk(gclk));
	jdff dff_A_6cvzohV45_0(.dout(w_dff_A_UsTjmVRQ3_0),.din(w_dff_A_6cvzohV45_0),.clk(gclk));
	jdff dff_A_UsTjmVRQ3_0(.dout(w_dff_A_rR8zS27X9_0),.din(w_dff_A_UsTjmVRQ3_0),.clk(gclk));
	jdff dff_A_rR8zS27X9_0(.dout(w_dff_A_4ZqyfDqN2_0),.din(w_dff_A_rR8zS27X9_0),.clk(gclk));
	jdff dff_A_4ZqyfDqN2_0(.dout(w_dff_A_O3GU8iZ41_0),.din(w_dff_A_4ZqyfDqN2_0),.clk(gclk));
	jdff dff_A_O3GU8iZ41_0(.dout(w_dff_A_99ZTIEvf8_0),.din(w_dff_A_O3GU8iZ41_0),.clk(gclk));
	jdff dff_A_99ZTIEvf8_0(.dout(w_dff_A_8B4xFIAQ8_0),.din(w_dff_A_99ZTIEvf8_0),.clk(gclk));
	jdff dff_A_8B4xFIAQ8_0(.dout(w_dff_A_JxyxPhpD7_0),.din(w_dff_A_8B4xFIAQ8_0),.clk(gclk));
	jdff dff_A_JxyxPhpD7_0(.dout(w_dff_A_r7pYV3yF9_0),.din(w_dff_A_JxyxPhpD7_0),.clk(gclk));
	jdff dff_A_r7pYV3yF9_0(.dout(w_dff_A_AbmCaJOa0_0),.din(w_dff_A_r7pYV3yF9_0),.clk(gclk));
	jdff dff_A_AbmCaJOa0_0(.dout(w_dff_A_uxrj627s5_0),.din(w_dff_A_AbmCaJOa0_0),.clk(gclk));
	jdff dff_A_uxrj627s5_0(.dout(w_dff_A_ezZdDTRe3_0),.din(w_dff_A_uxrj627s5_0),.clk(gclk));
	jdff dff_A_ezZdDTRe3_0(.dout(w_dff_A_fvd9W8f35_0),.din(w_dff_A_ezZdDTRe3_0),.clk(gclk));
	jdff dff_A_fvd9W8f35_0(.dout(w_dff_A_JZpUUvKC0_0),.din(w_dff_A_fvd9W8f35_0),.clk(gclk));
	jdff dff_A_JZpUUvKC0_0(.dout(w_dff_A_YNha8dyU4_0),.din(w_dff_A_JZpUUvKC0_0),.clk(gclk));
	jdff dff_A_YNha8dyU4_0(.dout(w_dff_A_MSYyxAlT7_0),.din(w_dff_A_YNha8dyU4_0),.clk(gclk));
	jdff dff_A_MSYyxAlT7_0(.dout(w_dff_A_nfprwjxH9_0),.din(w_dff_A_MSYyxAlT7_0),.clk(gclk));
	jdff dff_A_nfprwjxH9_0(.dout(f82),.din(w_dff_A_nfprwjxH9_0),.clk(gclk));
	jdff dff_A_4p69wJXZ0_2(.dout(w_dff_A_w6swdRjt0_0),.din(w_dff_A_4p69wJXZ0_2),.clk(gclk));
	jdff dff_A_w6swdRjt0_0(.dout(w_dff_A_DYyitRvE0_0),.din(w_dff_A_w6swdRjt0_0),.clk(gclk));
	jdff dff_A_DYyitRvE0_0(.dout(w_dff_A_kDoJtfHJ4_0),.din(w_dff_A_DYyitRvE0_0),.clk(gclk));
	jdff dff_A_kDoJtfHJ4_0(.dout(w_dff_A_hwk1w0Aw7_0),.din(w_dff_A_kDoJtfHJ4_0),.clk(gclk));
	jdff dff_A_hwk1w0Aw7_0(.dout(w_dff_A_WE2zlTBT3_0),.din(w_dff_A_hwk1w0Aw7_0),.clk(gclk));
	jdff dff_A_WE2zlTBT3_0(.dout(w_dff_A_pj09o6s77_0),.din(w_dff_A_WE2zlTBT3_0),.clk(gclk));
	jdff dff_A_pj09o6s77_0(.dout(w_dff_A_PhFsf0Zp3_0),.din(w_dff_A_pj09o6s77_0),.clk(gclk));
	jdff dff_A_PhFsf0Zp3_0(.dout(w_dff_A_QvzyRWzt3_0),.din(w_dff_A_PhFsf0Zp3_0),.clk(gclk));
	jdff dff_A_QvzyRWzt3_0(.dout(w_dff_A_4VF5fkN18_0),.din(w_dff_A_QvzyRWzt3_0),.clk(gclk));
	jdff dff_A_4VF5fkN18_0(.dout(w_dff_A_Z7Zqzz4r7_0),.din(w_dff_A_4VF5fkN18_0),.clk(gclk));
	jdff dff_A_Z7Zqzz4r7_0(.dout(w_dff_A_BCFbvDCh8_0),.din(w_dff_A_Z7Zqzz4r7_0),.clk(gclk));
	jdff dff_A_BCFbvDCh8_0(.dout(w_dff_A_2otiWYib1_0),.din(w_dff_A_BCFbvDCh8_0),.clk(gclk));
	jdff dff_A_2otiWYib1_0(.dout(w_dff_A_JotKQPNE3_0),.din(w_dff_A_2otiWYib1_0),.clk(gclk));
	jdff dff_A_JotKQPNE3_0(.dout(w_dff_A_r4M2cirP2_0),.din(w_dff_A_JotKQPNE3_0),.clk(gclk));
	jdff dff_A_r4M2cirP2_0(.dout(w_dff_A_GfUjDvhG3_0),.din(w_dff_A_r4M2cirP2_0),.clk(gclk));
	jdff dff_A_GfUjDvhG3_0(.dout(w_dff_A_9NAaC6I83_0),.din(w_dff_A_GfUjDvhG3_0),.clk(gclk));
	jdff dff_A_9NAaC6I83_0(.dout(w_dff_A_e32dyhpt2_0),.din(w_dff_A_9NAaC6I83_0),.clk(gclk));
	jdff dff_A_e32dyhpt2_0(.dout(w_dff_A_xZn3NlHG0_0),.din(w_dff_A_e32dyhpt2_0),.clk(gclk));
	jdff dff_A_xZn3NlHG0_0(.dout(w_dff_A_Em9QqonB7_0),.din(w_dff_A_xZn3NlHG0_0),.clk(gclk));
	jdff dff_A_Em9QqonB7_0(.dout(w_dff_A_fK589tDi0_0),.din(w_dff_A_Em9QqonB7_0),.clk(gclk));
	jdff dff_A_fK589tDi0_0(.dout(w_dff_A_gGxVkSsJ6_0),.din(w_dff_A_fK589tDi0_0),.clk(gclk));
	jdff dff_A_gGxVkSsJ6_0(.dout(w_dff_A_7dXuuxyI1_0),.din(w_dff_A_gGxVkSsJ6_0),.clk(gclk));
	jdff dff_A_7dXuuxyI1_0(.dout(w_dff_A_p0Pr2fSO0_0),.din(w_dff_A_7dXuuxyI1_0),.clk(gclk));
	jdff dff_A_p0Pr2fSO0_0(.dout(w_dff_A_AHH1acAs2_0),.din(w_dff_A_p0Pr2fSO0_0),.clk(gclk));
	jdff dff_A_AHH1acAs2_0(.dout(w_dff_A_0BETMRhT9_0),.din(w_dff_A_AHH1acAs2_0),.clk(gclk));
	jdff dff_A_0BETMRhT9_0(.dout(w_dff_A_tZHuPoOe4_0),.din(w_dff_A_0BETMRhT9_0),.clk(gclk));
	jdff dff_A_tZHuPoOe4_0(.dout(w_dff_A_RvQ9PZEn5_0),.din(w_dff_A_tZHuPoOe4_0),.clk(gclk));
	jdff dff_A_RvQ9PZEn5_0(.dout(w_dff_A_f1kVDeZt4_0),.din(w_dff_A_RvQ9PZEn5_0),.clk(gclk));
	jdff dff_A_f1kVDeZt4_0(.dout(w_dff_A_DSas78eH1_0),.din(w_dff_A_f1kVDeZt4_0),.clk(gclk));
	jdff dff_A_DSas78eH1_0(.dout(w_dff_A_2NUdOyvW2_0),.din(w_dff_A_DSas78eH1_0),.clk(gclk));
	jdff dff_A_2NUdOyvW2_0(.dout(w_dff_A_lD6CANcD9_0),.din(w_dff_A_2NUdOyvW2_0),.clk(gclk));
	jdff dff_A_lD6CANcD9_0(.dout(w_dff_A_0piiSHpC6_0),.din(w_dff_A_lD6CANcD9_0),.clk(gclk));
	jdff dff_A_0piiSHpC6_0(.dout(w_dff_A_1rj5URsD7_0),.din(w_dff_A_0piiSHpC6_0),.clk(gclk));
	jdff dff_A_1rj5URsD7_0(.dout(w_dff_A_hZ5QwYQ18_0),.din(w_dff_A_1rj5URsD7_0),.clk(gclk));
	jdff dff_A_hZ5QwYQ18_0(.dout(w_dff_A_0tirzuB48_0),.din(w_dff_A_hZ5QwYQ18_0),.clk(gclk));
	jdff dff_A_0tirzuB48_0(.dout(w_dff_A_tQuJ6dAA6_0),.din(w_dff_A_0tirzuB48_0),.clk(gclk));
	jdff dff_A_tQuJ6dAA6_0(.dout(w_dff_A_SNJKiRpp2_0),.din(w_dff_A_tQuJ6dAA6_0),.clk(gclk));
	jdff dff_A_SNJKiRpp2_0(.dout(w_dff_A_rdkxDQHx8_0),.din(w_dff_A_SNJKiRpp2_0),.clk(gclk));
	jdff dff_A_rdkxDQHx8_0(.dout(w_dff_A_ucC8WALG7_0),.din(w_dff_A_rdkxDQHx8_0),.clk(gclk));
	jdff dff_A_ucC8WALG7_0(.dout(w_dff_A_PWtwCDQG6_0),.din(w_dff_A_ucC8WALG7_0),.clk(gclk));
	jdff dff_A_PWtwCDQG6_0(.dout(w_dff_A_V9eJRzxA7_0),.din(w_dff_A_PWtwCDQG6_0),.clk(gclk));
	jdff dff_A_V9eJRzxA7_0(.dout(w_dff_A_Pvlm2YmH9_0),.din(w_dff_A_V9eJRzxA7_0),.clk(gclk));
	jdff dff_A_Pvlm2YmH9_0(.dout(w_dff_A_no2IkSJL9_0),.din(w_dff_A_Pvlm2YmH9_0),.clk(gclk));
	jdff dff_A_no2IkSJL9_0(.dout(f83),.din(w_dff_A_no2IkSJL9_0),.clk(gclk));
	jdff dff_A_BzE0H6ap0_2(.dout(w_dff_A_jqXYV3io5_0),.din(w_dff_A_BzE0H6ap0_2),.clk(gclk));
	jdff dff_A_jqXYV3io5_0(.dout(w_dff_A_iM3cI7Ek6_0),.din(w_dff_A_jqXYV3io5_0),.clk(gclk));
	jdff dff_A_iM3cI7Ek6_0(.dout(w_dff_A_iN6VqhOQ0_0),.din(w_dff_A_iM3cI7Ek6_0),.clk(gclk));
	jdff dff_A_iN6VqhOQ0_0(.dout(w_dff_A_k2dItjQP9_0),.din(w_dff_A_iN6VqhOQ0_0),.clk(gclk));
	jdff dff_A_k2dItjQP9_0(.dout(w_dff_A_5gdDEE0T4_0),.din(w_dff_A_k2dItjQP9_0),.clk(gclk));
	jdff dff_A_5gdDEE0T4_0(.dout(w_dff_A_8bikkJeO1_0),.din(w_dff_A_5gdDEE0T4_0),.clk(gclk));
	jdff dff_A_8bikkJeO1_0(.dout(w_dff_A_82vovMh69_0),.din(w_dff_A_8bikkJeO1_0),.clk(gclk));
	jdff dff_A_82vovMh69_0(.dout(w_dff_A_gxoAJqr45_0),.din(w_dff_A_82vovMh69_0),.clk(gclk));
	jdff dff_A_gxoAJqr45_0(.dout(w_dff_A_Sr6lQnSW3_0),.din(w_dff_A_gxoAJqr45_0),.clk(gclk));
	jdff dff_A_Sr6lQnSW3_0(.dout(w_dff_A_zGojD2vJ2_0),.din(w_dff_A_Sr6lQnSW3_0),.clk(gclk));
	jdff dff_A_zGojD2vJ2_0(.dout(w_dff_A_4CVwlnPI9_0),.din(w_dff_A_zGojD2vJ2_0),.clk(gclk));
	jdff dff_A_4CVwlnPI9_0(.dout(w_dff_A_tYwnkX7K0_0),.din(w_dff_A_4CVwlnPI9_0),.clk(gclk));
	jdff dff_A_tYwnkX7K0_0(.dout(w_dff_A_fbUEDZNy0_0),.din(w_dff_A_tYwnkX7K0_0),.clk(gclk));
	jdff dff_A_fbUEDZNy0_0(.dout(w_dff_A_pypTNgHF6_0),.din(w_dff_A_fbUEDZNy0_0),.clk(gclk));
	jdff dff_A_pypTNgHF6_0(.dout(w_dff_A_uP2eD7y00_0),.din(w_dff_A_pypTNgHF6_0),.clk(gclk));
	jdff dff_A_uP2eD7y00_0(.dout(w_dff_A_oqehDbgi8_0),.din(w_dff_A_uP2eD7y00_0),.clk(gclk));
	jdff dff_A_oqehDbgi8_0(.dout(w_dff_A_5woHGs6L2_0),.din(w_dff_A_oqehDbgi8_0),.clk(gclk));
	jdff dff_A_5woHGs6L2_0(.dout(w_dff_A_lKDEsdBe9_0),.din(w_dff_A_5woHGs6L2_0),.clk(gclk));
	jdff dff_A_lKDEsdBe9_0(.dout(w_dff_A_j3ETKEMN7_0),.din(w_dff_A_lKDEsdBe9_0),.clk(gclk));
	jdff dff_A_j3ETKEMN7_0(.dout(w_dff_A_36FGHFrT1_0),.din(w_dff_A_j3ETKEMN7_0),.clk(gclk));
	jdff dff_A_36FGHFrT1_0(.dout(w_dff_A_RBktoPcE9_0),.din(w_dff_A_36FGHFrT1_0),.clk(gclk));
	jdff dff_A_RBktoPcE9_0(.dout(w_dff_A_jP9anIDS5_0),.din(w_dff_A_RBktoPcE9_0),.clk(gclk));
	jdff dff_A_jP9anIDS5_0(.dout(w_dff_A_RA90Km4p2_0),.din(w_dff_A_jP9anIDS5_0),.clk(gclk));
	jdff dff_A_RA90Km4p2_0(.dout(w_dff_A_O9mtDMsS0_0),.din(w_dff_A_RA90Km4p2_0),.clk(gclk));
	jdff dff_A_O9mtDMsS0_0(.dout(w_dff_A_sIaRBHlt7_0),.din(w_dff_A_O9mtDMsS0_0),.clk(gclk));
	jdff dff_A_sIaRBHlt7_0(.dout(w_dff_A_KtB7i6bB7_0),.din(w_dff_A_sIaRBHlt7_0),.clk(gclk));
	jdff dff_A_KtB7i6bB7_0(.dout(w_dff_A_BktbEgcv8_0),.din(w_dff_A_KtB7i6bB7_0),.clk(gclk));
	jdff dff_A_BktbEgcv8_0(.dout(w_dff_A_gmnaJajv8_0),.din(w_dff_A_BktbEgcv8_0),.clk(gclk));
	jdff dff_A_gmnaJajv8_0(.dout(w_dff_A_X1nZomeb0_0),.din(w_dff_A_gmnaJajv8_0),.clk(gclk));
	jdff dff_A_X1nZomeb0_0(.dout(w_dff_A_dIw0KlYv2_0),.din(w_dff_A_X1nZomeb0_0),.clk(gclk));
	jdff dff_A_dIw0KlYv2_0(.dout(w_dff_A_LxkoDsqn5_0),.din(w_dff_A_dIw0KlYv2_0),.clk(gclk));
	jdff dff_A_LxkoDsqn5_0(.dout(w_dff_A_noRtGyXv7_0),.din(w_dff_A_LxkoDsqn5_0),.clk(gclk));
	jdff dff_A_noRtGyXv7_0(.dout(w_dff_A_43sNXuGm1_0),.din(w_dff_A_noRtGyXv7_0),.clk(gclk));
	jdff dff_A_43sNXuGm1_0(.dout(w_dff_A_6zOs2XEH1_0),.din(w_dff_A_43sNXuGm1_0),.clk(gclk));
	jdff dff_A_6zOs2XEH1_0(.dout(w_dff_A_OM6j7uCh3_0),.din(w_dff_A_6zOs2XEH1_0),.clk(gclk));
	jdff dff_A_OM6j7uCh3_0(.dout(w_dff_A_o1R1GBQb2_0),.din(w_dff_A_OM6j7uCh3_0),.clk(gclk));
	jdff dff_A_o1R1GBQb2_0(.dout(w_dff_A_XvBrxUTX9_0),.din(w_dff_A_o1R1GBQb2_0),.clk(gclk));
	jdff dff_A_XvBrxUTX9_0(.dout(w_dff_A_XSKLV1JD8_0),.din(w_dff_A_XvBrxUTX9_0),.clk(gclk));
	jdff dff_A_XSKLV1JD8_0(.dout(w_dff_A_AsBXM55u6_0),.din(w_dff_A_XSKLV1JD8_0),.clk(gclk));
	jdff dff_A_AsBXM55u6_0(.dout(w_dff_A_6HtQQHLd3_0),.din(w_dff_A_AsBXM55u6_0),.clk(gclk));
	jdff dff_A_6HtQQHLd3_0(.dout(w_dff_A_vY6mp8l88_0),.din(w_dff_A_6HtQQHLd3_0),.clk(gclk));
	jdff dff_A_vY6mp8l88_0(.dout(w_dff_A_yV6ELeiR1_0),.din(w_dff_A_vY6mp8l88_0),.clk(gclk));
	jdff dff_A_yV6ELeiR1_0(.dout(f84),.din(w_dff_A_yV6ELeiR1_0),.clk(gclk));
	jdff dff_A_TrXEhtji4_2(.dout(w_dff_A_mpLTf4219_0),.din(w_dff_A_TrXEhtji4_2),.clk(gclk));
	jdff dff_A_mpLTf4219_0(.dout(w_dff_A_TdqsOJT54_0),.din(w_dff_A_mpLTf4219_0),.clk(gclk));
	jdff dff_A_TdqsOJT54_0(.dout(w_dff_A_65dX4yMa8_0),.din(w_dff_A_TdqsOJT54_0),.clk(gclk));
	jdff dff_A_65dX4yMa8_0(.dout(w_dff_A_1ZBM88Ll0_0),.din(w_dff_A_65dX4yMa8_0),.clk(gclk));
	jdff dff_A_1ZBM88Ll0_0(.dout(w_dff_A_izqwe0jp3_0),.din(w_dff_A_1ZBM88Ll0_0),.clk(gclk));
	jdff dff_A_izqwe0jp3_0(.dout(w_dff_A_GIYMBYEK8_0),.din(w_dff_A_izqwe0jp3_0),.clk(gclk));
	jdff dff_A_GIYMBYEK8_0(.dout(w_dff_A_hS0PaYuw6_0),.din(w_dff_A_GIYMBYEK8_0),.clk(gclk));
	jdff dff_A_hS0PaYuw6_0(.dout(w_dff_A_0TknbbLh5_0),.din(w_dff_A_hS0PaYuw6_0),.clk(gclk));
	jdff dff_A_0TknbbLh5_0(.dout(w_dff_A_2fCd8o253_0),.din(w_dff_A_0TknbbLh5_0),.clk(gclk));
	jdff dff_A_2fCd8o253_0(.dout(w_dff_A_e8aMue1E6_0),.din(w_dff_A_2fCd8o253_0),.clk(gclk));
	jdff dff_A_e8aMue1E6_0(.dout(w_dff_A_6svRrmX85_0),.din(w_dff_A_e8aMue1E6_0),.clk(gclk));
	jdff dff_A_6svRrmX85_0(.dout(w_dff_A_7G0JMF6y4_0),.din(w_dff_A_6svRrmX85_0),.clk(gclk));
	jdff dff_A_7G0JMF6y4_0(.dout(w_dff_A_Zx36iGOO1_0),.din(w_dff_A_7G0JMF6y4_0),.clk(gclk));
	jdff dff_A_Zx36iGOO1_0(.dout(w_dff_A_LdHkQoIm5_0),.din(w_dff_A_Zx36iGOO1_0),.clk(gclk));
	jdff dff_A_LdHkQoIm5_0(.dout(w_dff_A_XF8NdbBB3_0),.din(w_dff_A_LdHkQoIm5_0),.clk(gclk));
	jdff dff_A_XF8NdbBB3_0(.dout(w_dff_A_m8NfSNeS9_0),.din(w_dff_A_XF8NdbBB3_0),.clk(gclk));
	jdff dff_A_m8NfSNeS9_0(.dout(w_dff_A_Lmimkaom8_0),.din(w_dff_A_m8NfSNeS9_0),.clk(gclk));
	jdff dff_A_Lmimkaom8_0(.dout(w_dff_A_o23dxbw04_0),.din(w_dff_A_Lmimkaom8_0),.clk(gclk));
	jdff dff_A_o23dxbw04_0(.dout(w_dff_A_WVIy7PyL2_0),.din(w_dff_A_o23dxbw04_0),.clk(gclk));
	jdff dff_A_WVIy7PyL2_0(.dout(w_dff_A_egOplusY3_0),.din(w_dff_A_WVIy7PyL2_0),.clk(gclk));
	jdff dff_A_egOplusY3_0(.dout(w_dff_A_RphwYfE68_0),.din(w_dff_A_egOplusY3_0),.clk(gclk));
	jdff dff_A_RphwYfE68_0(.dout(w_dff_A_kKuXQA7Z0_0),.din(w_dff_A_RphwYfE68_0),.clk(gclk));
	jdff dff_A_kKuXQA7Z0_0(.dout(w_dff_A_KhMiOUSE8_0),.din(w_dff_A_kKuXQA7Z0_0),.clk(gclk));
	jdff dff_A_KhMiOUSE8_0(.dout(w_dff_A_nQ3r0zES9_0),.din(w_dff_A_KhMiOUSE8_0),.clk(gclk));
	jdff dff_A_nQ3r0zES9_0(.dout(w_dff_A_fT2aOutz6_0),.din(w_dff_A_nQ3r0zES9_0),.clk(gclk));
	jdff dff_A_fT2aOutz6_0(.dout(w_dff_A_nfqndw8i1_0),.din(w_dff_A_fT2aOutz6_0),.clk(gclk));
	jdff dff_A_nfqndw8i1_0(.dout(w_dff_A_1IWjK4N52_0),.din(w_dff_A_nfqndw8i1_0),.clk(gclk));
	jdff dff_A_1IWjK4N52_0(.dout(w_dff_A_ssx3bLXm1_0),.din(w_dff_A_1IWjK4N52_0),.clk(gclk));
	jdff dff_A_ssx3bLXm1_0(.dout(w_dff_A_KtaWNVou5_0),.din(w_dff_A_ssx3bLXm1_0),.clk(gclk));
	jdff dff_A_KtaWNVou5_0(.dout(w_dff_A_Nx4XsKVS1_0),.din(w_dff_A_KtaWNVou5_0),.clk(gclk));
	jdff dff_A_Nx4XsKVS1_0(.dout(w_dff_A_bZe6fj7x7_0),.din(w_dff_A_Nx4XsKVS1_0),.clk(gclk));
	jdff dff_A_bZe6fj7x7_0(.dout(w_dff_A_P2tHqJUu4_0),.din(w_dff_A_bZe6fj7x7_0),.clk(gclk));
	jdff dff_A_P2tHqJUu4_0(.dout(w_dff_A_G27dZytw9_0),.din(w_dff_A_P2tHqJUu4_0),.clk(gclk));
	jdff dff_A_G27dZytw9_0(.dout(w_dff_A_rq0lcUhd8_0),.din(w_dff_A_G27dZytw9_0),.clk(gclk));
	jdff dff_A_rq0lcUhd8_0(.dout(w_dff_A_FNArPyWS6_0),.din(w_dff_A_rq0lcUhd8_0),.clk(gclk));
	jdff dff_A_FNArPyWS6_0(.dout(w_dff_A_sTBbMO137_0),.din(w_dff_A_FNArPyWS6_0),.clk(gclk));
	jdff dff_A_sTBbMO137_0(.dout(w_dff_A_FUmyjLvz8_0),.din(w_dff_A_sTBbMO137_0),.clk(gclk));
	jdff dff_A_FUmyjLvz8_0(.dout(w_dff_A_CVFYPaIh5_0),.din(w_dff_A_FUmyjLvz8_0),.clk(gclk));
	jdff dff_A_CVFYPaIh5_0(.dout(w_dff_A_wzfi7FZF1_0),.din(w_dff_A_CVFYPaIh5_0),.clk(gclk));
	jdff dff_A_wzfi7FZF1_0(.dout(w_dff_A_BfRZoENc7_0),.din(w_dff_A_wzfi7FZF1_0),.clk(gclk));
	jdff dff_A_BfRZoENc7_0(.dout(w_dff_A_cf7dJh6C1_0),.din(w_dff_A_BfRZoENc7_0),.clk(gclk));
	jdff dff_A_cf7dJh6C1_0(.dout(f85),.din(w_dff_A_cf7dJh6C1_0),.clk(gclk));
	jdff dff_A_HRCPkfMi4_2(.dout(w_dff_A_2rSjB1rj9_0),.din(w_dff_A_HRCPkfMi4_2),.clk(gclk));
	jdff dff_A_2rSjB1rj9_0(.dout(w_dff_A_iqMRMa617_0),.din(w_dff_A_2rSjB1rj9_0),.clk(gclk));
	jdff dff_A_iqMRMa617_0(.dout(w_dff_A_6Fm8woOG7_0),.din(w_dff_A_iqMRMa617_0),.clk(gclk));
	jdff dff_A_6Fm8woOG7_0(.dout(w_dff_A_1lyaeRjh6_0),.din(w_dff_A_6Fm8woOG7_0),.clk(gclk));
	jdff dff_A_1lyaeRjh6_0(.dout(w_dff_A_k0ULkyCV0_0),.din(w_dff_A_1lyaeRjh6_0),.clk(gclk));
	jdff dff_A_k0ULkyCV0_0(.dout(w_dff_A_Ehiqzdjb8_0),.din(w_dff_A_k0ULkyCV0_0),.clk(gclk));
	jdff dff_A_Ehiqzdjb8_0(.dout(w_dff_A_qirzyIXZ2_0),.din(w_dff_A_Ehiqzdjb8_0),.clk(gclk));
	jdff dff_A_qirzyIXZ2_0(.dout(w_dff_A_O4Pu32G29_0),.din(w_dff_A_qirzyIXZ2_0),.clk(gclk));
	jdff dff_A_O4Pu32G29_0(.dout(w_dff_A_gwExHQ2I9_0),.din(w_dff_A_O4Pu32G29_0),.clk(gclk));
	jdff dff_A_gwExHQ2I9_0(.dout(w_dff_A_JgJFqoPU0_0),.din(w_dff_A_gwExHQ2I9_0),.clk(gclk));
	jdff dff_A_JgJFqoPU0_0(.dout(w_dff_A_qXjWXTUg2_0),.din(w_dff_A_JgJFqoPU0_0),.clk(gclk));
	jdff dff_A_qXjWXTUg2_0(.dout(w_dff_A_ZQ9de3FM2_0),.din(w_dff_A_qXjWXTUg2_0),.clk(gclk));
	jdff dff_A_ZQ9de3FM2_0(.dout(w_dff_A_xXRfod5m7_0),.din(w_dff_A_ZQ9de3FM2_0),.clk(gclk));
	jdff dff_A_xXRfod5m7_0(.dout(w_dff_A_mQWgElrW4_0),.din(w_dff_A_xXRfod5m7_0),.clk(gclk));
	jdff dff_A_mQWgElrW4_0(.dout(w_dff_A_7HuCOhJ69_0),.din(w_dff_A_mQWgElrW4_0),.clk(gclk));
	jdff dff_A_7HuCOhJ69_0(.dout(w_dff_A_NP7LGG3o7_0),.din(w_dff_A_7HuCOhJ69_0),.clk(gclk));
	jdff dff_A_NP7LGG3o7_0(.dout(w_dff_A_l2hV5m1P4_0),.din(w_dff_A_NP7LGG3o7_0),.clk(gclk));
	jdff dff_A_l2hV5m1P4_0(.dout(w_dff_A_HfKafrgH8_0),.din(w_dff_A_l2hV5m1P4_0),.clk(gclk));
	jdff dff_A_HfKafrgH8_0(.dout(w_dff_A_Gtybz85Q5_0),.din(w_dff_A_HfKafrgH8_0),.clk(gclk));
	jdff dff_A_Gtybz85Q5_0(.dout(w_dff_A_s9rS4OiU4_0),.din(w_dff_A_Gtybz85Q5_0),.clk(gclk));
	jdff dff_A_s9rS4OiU4_0(.dout(w_dff_A_FDAwbgv15_0),.din(w_dff_A_s9rS4OiU4_0),.clk(gclk));
	jdff dff_A_FDAwbgv15_0(.dout(w_dff_A_Lc4MaL958_0),.din(w_dff_A_FDAwbgv15_0),.clk(gclk));
	jdff dff_A_Lc4MaL958_0(.dout(w_dff_A_lA7XbW9O8_0),.din(w_dff_A_Lc4MaL958_0),.clk(gclk));
	jdff dff_A_lA7XbW9O8_0(.dout(w_dff_A_nBj4Wp078_0),.din(w_dff_A_lA7XbW9O8_0),.clk(gclk));
	jdff dff_A_nBj4Wp078_0(.dout(w_dff_A_MujaL6on7_0),.din(w_dff_A_nBj4Wp078_0),.clk(gclk));
	jdff dff_A_MujaL6on7_0(.dout(w_dff_A_WQ6erECb2_0),.din(w_dff_A_MujaL6on7_0),.clk(gclk));
	jdff dff_A_WQ6erECb2_0(.dout(w_dff_A_Ga2QGedC7_0),.din(w_dff_A_WQ6erECb2_0),.clk(gclk));
	jdff dff_A_Ga2QGedC7_0(.dout(w_dff_A_k4aPPfJc9_0),.din(w_dff_A_Ga2QGedC7_0),.clk(gclk));
	jdff dff_A_k4aPPfJc9_0(.dout(w_dff_A_arGQulI27_0),.din(w_dff_A_k4aPPfJc9_0),.clk(gclk));
	jdff dff_A_arGQulI27_0(.dout(w_dff_A_5LKyl36z9_0),.din(w_dff_A_arGQulI27_0),.clk(gclk));
	jdff dff_A_5LKyl36z9_0(.dout(w_dff_A_3dajWwuL6_0),.din(w_dff_A_5LKyl36z9_0),.clk(gclk));
	jdff dff_A_3dajWwuL6_0(.dout(w_dff_A_y751QZU46_0),.din(w_dff_A_3dajWwuL6_0),.clk(gclk));
	jdff dff_A_y751QZU46_0(.dout(w_dff_A_uM1C7RSr4_0),.din(w_dff_A_y751QZU46_0),.clk(gclk));
	jdff dff_A_uM1C7RSr4_0(.dout(w_dff_A_piPDTxBJ9_0),.din(w_dff_A_uM1C7RSr4_0),.clk(gclk));
	jdff dff_A_piPDTxBJ9_0(.dout(w_dff_A_QaAUtGFn1_0),.din(w_dff_A_piPDTxBJ9_0),.clk(gclk));
	jdff dff_A_QaAUtGFn1_0(.dout(w_dff_A_YPwmxXCC7_0),.din(w_dff_A_QaAUtGFn1_0),.clk(gclk));
	jdff dff_A_YPwmxXCC7_0(.dout(w_dff_A_wTOgwcv32_0),.din(w_dff_A_YPwmxXCC7_0),.clk(gclk));
	jdff dff_A_wTOgwcv32_0(.dout(w_dff_A_qn030i954_0),.din(w_dff_A_wTOgwcv32_0),.clk(gclk));
	jdff dff_A_qn030i954_0(.dout(w_dff_A_4QHExuNR0_0),.din(w_dff_A_qn030i954_0),.clk(gclk));
	jdff dff_A_4QHExuNR0_0(.dout(w_dff_A_eTDEE6CM9_0),.din(w_dff_A_4QHExuNR0_0),.clk(gclk));
	jdff dff_A_eTDEE6CM9_0(.dout(f86),.din(w_dff_A_eTDEE6CM9_0),.clk(gclk));
	jdff dff_A_OCpaXqst8_2(.dout(w_dff_A_aL5mmWiS6_0),.din(w_dff_A_OCpaXqst8_2),.clk(gclk));
	jdff dff_A_aL5mmWiS6_0(.dout(w_dff_A_bH462nvr3_0),.din(w_dff_A_aL5mmWiS6_0),.clk(gclk));
	jdff dff_A_bH462nvr3_0(.dout(w_dff_A_JTtXoK2j6_0),.din(w_dff_A_bH462nvr3_0),.clk(gclk));
	jdff dff_A_JTtXoK2j6_0(.dout(w_dff_A_pJWDczQd6_0),.din(w_dff_A_JTtXoK2j6_0),.clk(gclk));
	jdff dff_A_pJWDczQd6_0(.dout(w_dff_A_eF43UynL5_0),.din(w_dff_A_pJWDczQd6_0),.clk(gclk));
	jdff dff_A_eF43UynL5_0(.dout(w_dff_A_2F4wQ4656_0),.din(w_dff_A_eF43UynL5_0),.clk(gclk));
	jdff dff_A_2F4wQ4656_0(.dout(w_dff_A_dodhWfV67_0),.din(w_dff_A_2F4wQ4656_0),.clk(gclk));
	jdff dff_A_dodhWfV67_0(.dout(w_dff_A_M85m3UCZ3_0),.din(w_dff_A_dodhWfV67_0),.clk(gclk));
	jdff dff_A_M85m3UCZ3_0(.dout(w_dff_A_k5mq6NGH2_0),.din(w_dff_A_M85m3UCZ3_0),.clk(gclk));
	jdff dff_A_k5mq6NGH2_0(.dout(w_dff_A_45qwoUnC1_0),.din(w_dff_A_k5mq6NGH2_0),.clk(gclk));
	jdff dff_A_45qwoUnC1_0(.dout(w_dff_A_Zm8yimOu9_0),.din(w_dff_A_45qwoUnC1_0),.clk(gclk));
	jdff dff_A_Zm8yimOu9_0(.dout(w_dff_A_FtVypjpd1_0),.din(w_dff_A_Zm8yimOu9_0),.clk(gclk));
	jdff dff_A_FtVypjpd1_0(.dout(w_dff_A_0NQCeKcb4_0),.din(w_dff_A_FtVypjpd1_0),.clk(gclk));
	jdff dff_A_0NQCeKcb4_0(.dout(w_dff_A_oyOid39a5_0),.din(w_dff_A_0NQCeKcb4_0),.clk(gclk));
	jdff dff_A_oyOid39a5_0(.dout(w_dff_A_YS9ywHnL6_0),.din(w_dff_A_oyOid39a5_0),.clk(gclk));
	jdff dff_A_YS9ywHnL6_0(.dout(w_dff_A_jpXggtwh9_0),.din(w_dff_A_YS9ywHnL6_0),.clk(gclk));
	jdff dff_A_jpXggtwh9_0(.dout(w_dff_A_dnUP1o4t7_0),.din(w_dff_A_jpXggtwh9_0),.clk(gclk));
	jdff dff_A_dnUP1o4t7_0(.dout(w_dff_A_VcZJVNcg1_0),.din(w_dff_A_dnUP1o4t7_0),.clk(gclk));
	jdff dff_A_VcZJVNcg1_0(.dout(w_dff_A_asYK8RaT8_0),.din(w_dff_A_VcZJVNcg1_0),.clk(gclk));
	jdff dff_A_asYK8RaT8_0(.dout(w_dff_A_g7nJLmRe3_0),.din(w_dff_A_asYK8RaT8_0),.clk(gclk));
	jdff dff_A_g7nJLmRe3_0(.dout(w_dff_A_zaoU9vPq4_0),.din(w_dff_A_g7nJLmRe3_0),.clk(gclk));
	jdff dff_A_zaoU9vPq4_0(.dout(w_dff_A_W5OoMSxm9_0),.din(w_dff_A_zaoU9vPq4_0),.clk(gclk));
	jdff dff_A_W5OoMSxm9_0(.dout(w_dff_A_5JaNrVKA2_0),.din(w_dff_A_W5OoMSxm9_0),.clk(gclk));
	jdff dff_A_5JaNrVKA2_0(.dout(w_dff_A_2gtmGbdx0_0),.din(w_dff_A_5JaNrVKA2_0),.clk(gclk));
	jdff dff_A_2gtmGbdx0_0(.dout(w_dff_A_0J3tUHCV0_0),.din(w_dff_A_2gtmGbdx0_0),.clk(gclk));
	jdff dff_A_0J3tUHCV0_0(.dout(w_dff_A_o2qh2RJa6_0),.din(w_dff_A_0J3tUHCV0_0),.clk(gclk));
	jdff dff_A_o2qh2RJa6_0(.dout(w_dff_A_BNOrYJj89_0),.din(w_dff_A_o2qh2RJa6_0),.clk(gclk));
	jdff dff_A_BNOrYJj89_0(.dout(w_dff_A_HUqCe9rY8_0),.din(w_dff_A_BNOrYJj89_0),.clk(gclk));
	jdff dff_A_HUqCe9rY8_0(.dout(w_dff_A_Au62QzpP0_0),.din(w_dff_A_HUqCe9rY8_0),.clk(gclk));
	jdff dff_A_Au62QzpP0_0(.dout(w_dff_A_nqEkH5jt7_0),.din(w_dff_A_Au62QzpP0_0),.clk(gclk));
	jdff dff_A_nqEkH5jt7_0(.dout(w_dff_A_md8dCJji6_0),.din(w_dff_A_nqEkH5jt7_0),.clk(gclk));
	jdff dff_A_md8dCJji6_0(.dout(w_dff_A_YPHI7fn75_0),.din(w_dff_A_md8dCJji6_0),.clk(gclk));
	jdff dff_A_YPHI7fn75_0(.dout(w_dff_A_hUAL0c5w9_0),.din(w_dff_A_YPHI7fn75_0),.clk(gclk));
	jdff dff_A_hUAL0c5w9_0(.dout(w_dff_A_yGXTXH4b5_0),.din(w_dff_A_hUAL0c5w9_0),.clk(gclk));
	jdff dff_A_yGXTXH4b5_0(.dout(w_dff_A_scTJkbhP1_0),.din(w_dff_A_yGXTXH4b5_0),.clk(gclk));
	jdff dff_A_scTJkbhP1_0(.dout(w_dff_A_kVrUBjav0_0),.din(w_dff_A_scTJkbhP1_0),.clk(gclk));
	jdff dff_A_kVrUBjav0_0(.dout(w_dff_A_ry5okceN1_0),.din(w_dff_A_kVrUBjav0_0),.clk(gclk));
	jdff dff_A_ry5okceN1_0(.dout(w_dff_A_TatD4bdV2_0),.din(w_dff_A_ry5okceN1_0),.clk(gclk));
	jdff dff_A_TatD4bdV2_0(.dout(w_dff_A_izocvOpF5_0),.din(w_dff_A_TatD4bdV2_0),.clk(gclk));
	jdff dff_A_izocvOpF5_0(.dout(f87),.din(w_dff_A_izocvOpF5_0),.clk(gclk));
	jdff dff_A_LDFLxawb9_2(.dout(w_dff_A_tHuYhkTX8_0),.din(w_dff_A_LDFLxawb9_2),.clk(gclk));
	jdff dff_A_tHuYhkTX8_0(.dout(w_dff_A_hLRD023M9_0),.din(w_dff_A_tHuYhkTX8_0),.clk(gclk));
	jdff dff_A_hLRD023M9_0(.dout(w_dff_A_s5yBq3Zu2_0),.din(w_dff_A_hLRD023M9_0),.clk(gclk));
	jdff dff_A_s5yBq3Zu2_0(.dout(w_dff_A_H28RLnpR3_0),.din(w_dff_A_s5yBq3Zu2_0),.clk(gclk));
	jdff dff_A_H28RLnpR3_0(.dout(w_dff_A_fHKYOYnC1_0),.din(w_dff_A_H28RLnpR3_0),.clk(gclk));
	jdff dff_A_fHKYOYnC1_0(.dout(w_dff_A_vASC2l875_0),.din(w_dff_A_fHKYOYnC1_0),.clk(gclk));
	jdff dff_A_vASC2l875_0(.dout(w_dff_A_GL1cxy0p6_0),.din(w_dff_A_vASC2l875_0),.clk(gclk));
	jdff dff_A_GL1cxy0p6_0(.dout(w_dff_A_4hgHlFrK8_0),.din(w_dff_A_GL1cxy0p6_0),.clk(gclk));
	jdff dff_A_4hgHlFrK8_0(.dout(w_dff_A_3V51jYAo2_0),.din(w_dff_A_4hgHlFrK8_0),.clk(gclk));
	jdff dff_A_3V51jYAo2_0(.dout(w_dff_A_nYbXU8e86_0),.din(w_dff_A_3V51jYAo2_0),.clk(gclk));
	jdff dff_A_nYbXU8e86_0(.dout(w_dff_A_MQ1dVrCQ4_0),.din(w_dff_A_nYbXU8e86_0),.clk(gclk));
	jdff dff_A_MQ1dVrCQ4_0(.dout(w_dff_A_hRaXDNNJ6_0),.din(w_dff_A_MQ1dVrCQ4_0),.clk(gclk));
	jdff dff_A_hRaXDNNJ6_0(.dout(w_dff_A_9f2K14Wl0_0),.din(w_dff_A_hRaXDNNJ6_0),.clk(gclk));
	jdff dff_A_9f2K14Wl0_0(.dout(w_dff_A_A0IN27wo8_0),.din(w_dff_A_9f2K14Wl0_0),.clk(gclk));
	jdff dff_A_A0IN27wo8_0(.dout(w_dff_A_YAtJlaxc2_0),.din(w_dff_A_A0IN27wo8_0),.clk(gclk));
	jdff dff_A_YAtJlaxc2_0(.dout(w_dff_A_ntlwEz2f3_0),.din(w_dff_A_YAtJlaxc2_0),.clk(gclk));
	jdff dff_A_ntlwEz2f3_0(.dout(w_dff_A_C4D9PtUC8_0),.din(w_dff_A_ntlwEz2f3_0),.clk(gclk));
	jdff dff_A_C4D9PtUC8_0(.dout(w_dff_A_kXJN3uGx6_0),.din(w_dff_A_C4D9PtUC8_0),.clk(gclk));
	jdff dff_A_kXJN3uGx6_0(.dout(w_dff_A_f2QHW6iK3_0),.din(w_dff_A_kXJN3uGx6_0),.clk(gclk));
	jdff dff_A_f2QHW6iK3_0(.dout(w_dff_A_bYB5QZVH1_0),.din(w_dff_A_f2QHW6iK3_0),.clk(gclk));
	jdff dff_A_bYB5QZVH1_0(.dout(w_dff_A_b5K3EeYA0_0),.din(w_dff_A_bYB5QZVH1_0),.clk(gclk));
	jdff dff_A_b5K3EeYA0_0(.dout(w_dff_A_LyHIUixr3_0),.din(w_dff_A_b5K3EeYA0_0),.clk(gclk));
	jdff dff_A_LyHIUixr3_0(.dout(w_dff_A_Q5eV4ttV0_0),.din(w_dff_A_LyHIUixr3_0),.clk(gclk));
	jdff dff_A_Q5eV4ttV0_0(.dout(w_dff_A_buEUpT5x9_0),.din(w_dff_A_Q5eV4ttV0_0),.clk(gclk));
	jdff dff_A_buEUpT5x9_0(.dout(w_dff_A_a9Cq3sRo7_0),.din(w_dff_A_buEUpT5x9_0),.clk(gclk));
	jdff dff_A_a9Cq3sRo7_0(.dout(w_dff_A_O24ThT117_0),.din(w_dff_A_a9Cq3sRo7_0),.clk(gclk));
	jdff dff_A_O24ThT117_0(.dout(w_dff_A_K18XR8Xr6_0),.din(w_dff_A_O24ThT117_0),.clk(gclk));
	jdff dff_A_K18XR8Xr6_0(.dout(w_dff_A_j2NTQjsH6_0),.din(w_dff_A_K18XR8Xr6_0),.clk(gclk));
	jdff dff_A_j2NTQjsH6_0(.dout(w_dff_A_WhluNXyf6_0),.din(w_dff_A_j2NTQjsH6_0),.clk(gclk));
	jdff dff_A_WhluNXyf6_0(.dout(w_dff_A_9xtWOCfE8_0),.din(w_dff_A_WhluNXyf6_0),.clk(gclk));
	jdff dff_A_9xtWOCfE8_0(.dout(w_dff_A_NvOBlU3t9_0),.din(w_dff_A_9xtWOCfE8_0),.clk(gclk));
	jdff dff_A_NvOBlU3t9_0(.dout(w_dff_A_dCFjroEQ9_0),.din(w_dff_A_NvOBlU3t9_0),.clk(gclk));
	jdff dff_A_dCFjroEQ9_0(.dout(w_dff_A_4Z7M4SiK4_0),.din(w_dff_A_dCFjroEQ9_0),.clk(gclk));
	jdff dff_A_4Z7M4SiK4_0(.dout(w_dff_A_AJCKv0OJ9_0),.din(w_dff_A_4Z7M4SiK4_0),.clk(gclk));
	jdff dff_A_AJCKv0OJ9_0(.dout(w_dff_A_D96b6KHj4_0),.din(w_dff_A_AJCKv0OJ9_0),.clk(gclk));
	jdff dff_A_D96b6KHj4_0(.dout(w_dff_A_QHQsfEFF3_0),.din(w_dff_A_D96b6KHj4_0),.clk(gclk));
	jdff dff_A_QHQsfEFF3_0(.dout(w_dff_A_A6Dz6kOs4_0),.din(w_dff_A_QHQsfEFF3_0),.clk(gclk));
	jdff dff_A_A6Dz6kOs4_0(.dout(w_dff_A_n1lhhwon3_0),.din(w_dff_A_A6Dz6kOs4_0),.clk(gclk));
	jdff dff_A_n1lhhwon3_0(.dout(f88),.din(w_dff_A_n1lhhwon3_0),.clk(gclk));
	jdff dff_A_6JucvmkC3_2(.dout(w_dff_A_r8Uz5tCr3_0),.din(w_dff_A_6JucvmkC3_2),.clk(gclk));
	jdff dff_A_r8Uz5tCr3_0(.dout(w_dff_A_y5A7ROmk9_0),.din(w_dff_A_r8Uz5tCr3_0),.clk(gclk));
	jdff dff_A_y5A7ROmk9_0(.dout(w_dff_A_q7qUTkmZ4_0),.din(w_dff_A_y5A7ROmk9_0),.clk(gclk));
	jdff dff_A_q7qUTkmZ4_0(.dout(w_dff_A_9Ba0qRj96_0),.din(w_dff_A_q7qUTkmZ4_0),.clk(gclk));
	jdff dff_A_9Ba0qRj96_0(.dout(w_dff_A_mBnU1qsY4_0),.din(w_dff_A_9Ba0qRj96_0),.clk(gclk));
	jdff dff_A_mBnU1qsY4_0(.dout(w_dff_A_bJgbDpJn3_0),.din(w_dff_A_mBnU1qsY4_0),.clk(gclk));
	jdff dff_A_bJgbDpJn3_0(.dout(w_dff_A_BbDa7xMc0_0),.din(w_dff_A_bJgbDpJn3_0),.clk(gclk));
	jdff dff_A_BbDa7xMc0_0(.dout(w_dff_A_wVRommd89_0),.din(w_dff_A_BbDa7xMc0_0),.clk(gclk));
	jdff dff_A_wVRommd89_0(.dout(w_dff_A_C6jrz7uf4_0),.din(w_dff_A_wVRommd89_0),.clk(gclk));
	jdff dff_A_C6jrz7uf4_0(.dout(w_dff_A_VTxTo4Xn0_0),.din(w_dff_A_C6jrz7uf4_0),.clk(gclk));
	jdff dff_A_VTxTo4Xn0_0(.dout(w_dff_A_909EZ1Vm2_0),.din(w_dff_A_VTxTo4Xn0_0),.clk(gclk));
	jdff dff_A_909EZ1Vm2_0(.dout(w_dff_A_hHV0onUZ0_0),.din(w_dff_A_909EZ1Vm2_0),.clk(gclk));
	jdff dff_A_hHV0onUZ0_0(.dout(w_dff_A_K7gMtYAm4_0),.din(w_dff_A_hHV0onUZ0_0),.clk(gclk));
	jdff dff_A_K7gMtYAm4_0(.dout(w_dff_A_CmsjPF7W1_0),.din(w_dff_A_K7gMtYAm4_0),.clk(gclk));
	jdff dff_A_CmsjPF7W1_0(.dout(w_dff_A_nSZOk3yf3_0),.din(w_dff_A_CmsjPF7W1_0),.clk(gclk));
	jdff dff_A_nSZOk3yf3_0(.dout(w_dff_A_UyjAO2PB8_0),.din(w_dff_A_nSZOk3yf3_0),.clk(gclk));
	jdff dff_A_UyjAO2PB8_0(.dout(w_dff_A_Q0WTtCKU1_0),.din(w_dff_A_UyjAO2PB8_0),.clk(gclk));
	jdff dff_A_Q0WTtCKU1_0(.dout(w_dff_A_gojJTxL90_0),.din(w_dff_A_Q0WTtCKU1_0),.clk(gclk));
	jdff dff_A_gojJTxL90_0(.dout(w_dff_A_nDKChvTu5_0),.din(w_dff_A_gojJTxL90_0),.clk(gclk));
	jdff dff_A_nDKChvTu5_0(.dout(w_dff_A_InsADXP52_0),.din(w_dff_A_nDKChvTu5_0),.clk(gclk));
	jdff dff_A_InsADXP52_0(.dout(w_dff_A_451P4qkv5_0),.din(w_dff_A_InsADXP52_0),.clk(gclk));
	jdff dff_A_451P4qkv5_0(.dout(w_dff_A_teEmgDa31_0),.din(w_dff_A_451P4qkv5_0),.clk(gclk));
	jdff dff_A_teEmgDa31_0(.dout(w_dff_A_hW8ZtUsF5_0),.din(w_dff_A_teEmgDa31_0),.clk(gclk));
	jdff dff_A_hW8ZtUsF5_0(.dout(w_dff_A_LCfGoxfb7_0),.din(w_dff_A_hW8ZtUsF5_0),.clk(gclk));
	jdff dff_A_LCfGoxfb7_0(.dout(w_dff_A_L0Hj4WZc1_0),.din(w_dff_A_LCfGoxfb7_0),.clk(gclk));
	jdff dff_A_L0Hj4WZc1_0(.dout(w_dff_A_gZ1R2zXt6_0),.din(w_dff_A_L0Hj4WZc1_0),.clk(gclk));
	jdff dff_A_gZ1R2zXt6_0(.dout(w_dff_A_x0XWrMoh0_0),.din(w_dff_A_gZ1R2zXt6_0),.clk(gclk));
	jdff dff_A_x0XWrMoh0_0(.dout(w_dff_A_ICDD4oHo3_0),.din(w_dff_A_x0XWrMoh0_0),.clk(gclk));
	jdff dff_A_ICDD4oHo3_0(.dout(w_dff_A_vmsaB1HH5_0),.din(w_dff_A_ICDD4oHo3_0),.clk(gclk));
	jdff dff_A_vmsaB1HH5_0(.dout(w_dff_A_9mqdupKU3_0),.din(w_dff_A_vmsaB1HH5_0),.clk(gclk));
	jdff dff_A_9mqdupKU3_0(.dout(w_dff_A_X0974R2u0_0),.din(w_dff_A_9mqdupKU3_0),.clk(gclk));
	jdff dff_A_X0974R2u0_0(.dout(w_dff_A_6CNYcLKx3_0),.din(w_dff_A_X0974R2u0_0),.clk(gclk));
	jdff dff_A_6CNYcLKx3_0(.dout(w_dff_A_NCqyXU4Z2_0),.din(w_dff_A_6CNYcLKx3_0),.clk(gclk));
	jdff dff_A_NCqyXU4Z2_0(.dout(w_dff_A_PUluDnQW3_0),.din(w_dff_A_NCqyXU4Z2_0),.clk(gclk));
	jdff dff_A_PUluDnQW3_0(.dout(w_dff_A_hQwWJGOh7_0),.din(w_dff_A_PUluDnQW3_0),.clk(gclk));
	jdff dff_A_hQwWJGOh7_0(.dout(w_dff_A_xXVYilAv6_0),.din(w_dff_A_hQwWJGOh7_0),.clk(gclk));
	jdff dff_A_xXVYilAv6_0(.dout(w_dff_A_kNbKvpbM7_0),.din(w_dff_A_xXVYilAv6_0),.clk(gclk));
	jdff dff_A_kNbKvpbM7_0(.dout(f89),.din(w_dff_A_kNbKvpbM7_0),.clk(gclk));
	jdff dff_A_7kDqg9E90_2(.dout(w_dff_A_w1v5wgod7_0),.din(w_dff_A_7kDqg9E90_2),.clk(gclk));
	jdff dff_A_w1v5wgod7_0(.dout(w_dff_A_mrqQ34YW0_0),.din(w_dff_A_w1v5wgod7_0),.clk(gclk));
	jdff dff_A_mrqQ34YW0_0(.dout(w_dff_A_peT6RoWX1_0),.din(w_dff_A_mrqQ34YW0_0),.clk(gclk));
	jdff dff_A_peT6RoWX1_0(.dout(w_dff_A_zrYxOMZs0_0),.din(w_dff_A_peT6RoWX1_0),.clk(gclk));
	jdff dff_A_zrYxOMZs0_0(.dout(w_dff_A_UIquMr658_0),.din(w_dff_A_zrYxOMZs0_0),.clk(gclk));
	jdff dff_A_UIquMr658_0(.dout(w_dff_A_dAcENKSM7_0),.din(w_dff_A_UIquMr658_0),.clk(gclk));
	jdff dff_A_dAcENKSM7_0(.dout(w_dff_A_6pyLv7aY9_0),.din(w_dff_A_dAcENKSM7_0),.clk(gclk));
	jdff dff_A_6pyLv7aY9_0(.dout(w_dff_A_4GRSAY1B4_0),.din(w_dff_A_6pyLv7aY9_0),.clk(gclk));
	jdff dff_A_4GRSAY1B4_0(.dout(w_dff_A_z7q2J3wv7_0),.din(w_dff_A_4GRSAY1B4_0),.clk(gclk));
	jdff dff_A_z7q2J3wv7_0(.dout(w_dff_A_Trh8OoQS0_0),.din(w_dff_A_z7q2J3wv7_0),.clk(gclk));
	jdff dff_A_Trh8OoQS0_0(.dout(w_dff_A_yF9MVNaO4_0),.din(w_dff_A_Trh8OoQS0_0),.clk(gclk));
	jdff dff_A_yF9MVNaO4_0(.dout(w_dff_A_arc6ByMn9_0),.din(w_dff_A_yF9MVNaO4_0),.clk(gclk));
	jdff dff_A_arc6ByMn9_0(.dout(w_dff_A_bq6j5ewq2_0),.din(w_dff_A_arc6ByMn9_0),.clk(gclk));
	jdff dff_A_bq6j5ewq2_0(.dout(w_dff_A_Yg9vO6lc4_0),.din(w_dff_A_bq6j5ewq2_0),.clk(gclk));
	jdff dff_A_Yg9vO6lc4_0(.dout(w_dff_A_L7wIM2tI9_0),.din(w_dff_A_Yg9vO6lc4_0),.clk(gclk));
	jdff dff_A_L7wIM2tI9_0(.dout(w_dff_A_megLYJw99_0),.din(w_dff_A_L7wIM2tI9_0),.clk(gclk));
	jdff dff_A_megLYJw99_0(.dout(w_dff_A_c3stksiv6_0),.din(w_dff_A_megLYJw99_0),.clk(gclk));
	jdff dff_A_c3stksiv6_0(.dout(w_dff_A_eioubO7q2_0),.din(w_dff_A_c3stksiv6_0),.clk(gclk));
	jdff dff_A_eioubO7q2_0(.dout(w_dff_A_iEdmvH551_0),.din(w_dff_A_eioubO7q2_0),.clk(gclk));
	jdff dff_A_iEdmvH551_0(.dout(w_dff_A_nltm93702_0),.din(w_dff_A_iEdmvH551_0),.clk(gclk));
	jdff dff_A_nltm93702_0(.dout(w_dff_A_P9jat2O28_0),.din(w_dff_A_nltm93702_0),.clk(gclk));
	jdff dff_A_P9jat2O28_0(.dout(w_dff_A_NpNc9lKT6_0),.din(w_dff_A_P9jat2O28_0),.clk(gclk));
	jdff dff_A_NpNc9lKT6_0(.dout(w_dff_A_lkLePOwx5_0),.din(w_dff_A_NpNc9lKT6_0),.clk(gclk));
	jdff dff_A_lkLePOwx5_0(.dout(w_dff_A_KtzlBNsZ5_0),.din(w_dff_A_lkLePOwx5_0),.clk(gclk));
	jdff dff_A_KtzlBNsZ5_0(.dout(w_dff_A_Ozaj3MJi7_0),.din(w_dff_A_KtzlBNsZ5_0),.clk(gclk));
	jdff dff_A_Ozaj3MJi7_0(.dout(w_dff_A_r3xfQC3E5_0),.din(w_dff_A_Ozaj3MJi7_0),.clk(gclk));
	jdff dff_A_r3xfQC3E5_0(.dout(w_dff_A_UELLSaGU0_0),.din(w_dff_A_r3xfQC3E5_0),.clk(gclk));
	jdff dff_A_UELLSaGU0_0(.dout(w_dff_A_ORLJKkOG4_0),.din(w_dff_A_UELLSaGU0_0),.clk(gclk));
	jdff dff_A_ORLJKkOG4_0(.dout(w_dff_A_HPk4UVUJ8_0),.din(w_dff_A_ORLJKkOG4_0),.clk(gclk));
	jdff dff_A_HPk4UVUJ8_0(.dout(w_dff_A_qrccpb3i0_0),.din(w_dff_A_HPk4UVUJ8_0),.clk(gclk));
	jdff dff_A_qrccpb3i0_0(.dout(w_dff_A_bvv7RRTT7_0),.din(w_dff_A_qrccpb3i0_0),.clk(gclk));
	jdff dff_A_bvv7RRTT7_0(.dout(w_dff_A_G6Ijt2045_0),.din(w_dff_A_bvv7RRTT7_0),.clk(gclk));
	jdff dff_A_G6Ijt2045_0(.dout(w_dff_A_ZZeqKtMi4_0),.din(w_dff_A_G6Ijt2045_0),.clk(gclk));
	jdff dff_A_ZZeqKtMi4_0(.dout(w_dff_A_s2C7haa13_0),.din(w_dff_A_ZZeqKtMi4_0),.clk(gclk));
	jdff dff_A_s2C7haa13_0(.dout(w_dff_A_oAeOVQOF6_0),.din(w_dff_A_s2C7haa13_0),.clk(gclk));
	jdff dff_A_oAeOVQOF6_0(.dout(w_dff_A_VDrkGpMV2_0),.din(w_dff_A_oAeOVQOF6_0),.clk(gclk));
	jdff dff_A_VDrkGpMV2_0(.dout(f90),.din(w_dff_A_VDrkGpMV2_0),.clk(gclk));
	jdff dff_A_oKzz53IO5_2(.dout(w_dff_A_lyJ8Fdoz1_0),.din(w_dff_A_oKzz53IO5_2),.clk(gclk));
	jdff dff_A_lyJ8Fdoz1_0(.dout(w_dff_A_1xJrJYEB8_0),.din(w_dff_A_lyJ8Fdoz1_0),.clk(gclk));
	jdff dff_A_1xJrJYEB8_0(.dout(w_dff_A_xyQ40gwT1_0),.din(w_dff_A_1xJrJYEB8_0),.clk(gclk));
	jdff dff_A_xyQ40gwT1_0(.dout(w_dff_A_aI10CsNS8_0),.din(w_dff_A_xyQ40gwT1_0),.clk(gclk));
	jdff dff_A_aI10CsNS8_0(.dout(w_dff_A_XWcZECy74_0),.din(w_dff_A_aI10CsNS8_0),.clk(gclk));
	jdff dff_A_XWcZECy74_0(.dout(w_dff_A_Cys1BEmO3_0),.din(w_dff_A_XWcZECy74_0),.clk(gclk));
	jdff dff_A_Cys1BEmO3_0(.dout(w_dff_A_yZiay1Ra5_0),.din(w_dff_A_Cys1BEmO3_0),.clk(gclk));
	jdff dff_A_yZiay1Ra5_0(.dout(w_dff_A_CQcn7UCA4_0),.din(w_dff_A_yZiay1Ra5_0),.clk(gclk));
	jdff dff_A_CQcn7UCA4_0(.dout(w_dff_A_RXthB2Mn2_0),.din(w_dff_A_CQcn7UCA4_0),.clk(gclk));
	jdff dff_A_RXthB2Mn2_0(.dout(w_dff_A_IJfONVh88_0),.din(w_dff_A_RXthB2Mn2_0),.clk(gclk));
	jdff dff_A_IJfONVh88_0(.dout(w_dff_A_IdEcnlQK2_0),.din(w_dff_A_IJfONVh88_0),.clk(gclk));
	jdff dff_A_IdEcnlQK2_0(.dout(w_dff_A_tRJZPFQj6_0),.din(w_dff_A_IdEcnlQK2_0),.clk(gclk));
	jdff dff_A_tRJZPFQj6_0(.dout(w_dff_A_1NU2Sj192_0),.din(w_dff_A_tRJZPFQj6_0),.clk(gclk));
	jdff dff_A_1NU2Sj192_0(.dout(w_dff_A_6NWdFAQ88_0),.din(w_dff_A_1NU2Sj192_0),.clk(gclk));
	jdff dff_A_6NWdFAQ88_0(.dout(w_dff_A_6VZCquiV0_0),.din(w_dff_A_6NWdFAQ88_0),.clk(gclk));
	jdff dff_A_6VZCquiV0_0(.dout(w_dff_A_2Atwsl1e8_0),.din(w_dff_A_6VZCquiV0_0),.clk(gclk));
	jdff dff_A_2Atwsl1e8_0(.dout(w_dff_A_h7JwT59k0_0),.din(w_dff_A_2Atwsl1e8_0),.clk(gclk));
	jdff dff_A_h7JwT59k0_0(.dout(w_dff_A_1eHLkgSZ4_0),.din(w_dff_A_h7JwT59k0_0),.clk(gclk));
	jdff dff_A_1eHLkgSZ4_0(.dout(w_dff_A_iKWKqtI07_0),.din(w_dff_A_1eHLkgSZ4_0),.clk(gclk));
	jdff dff_A_iKWKqtI07_0(.dout(w_dff_A_9jX8atez9_0),.din(w_dff_A_iKWKqtI07_0),.clk(gclk));
	jdff dff_A_9jX8atez9_0(.dout(w_dff_A_x99zwbsx6_0),.din(w_dff_A_9jX8atez9_0),.clk(gclk));
	jdff dff_A_x99zwbsx6_0(.dout(w_dff_A_XGMUizW88_0),.din(w_dff_A_x99zwbsx6_0),.clk(gclk));
	jdff dff_A_XGMUizW88_0(.dout(w_dff_A_NgRQ9sQv0_0),.din(w_dff_A_XGMUizW88_0),.clk(gclk));
	jdff dff_A_NgRQ9sQv0_0(.dout(w_dff_A_YdYiZ7AU3_0),.din(w_dff_A_NgRQ9sQv0_0),.clk(gclk));
	jdff dff_A_YdYiZ7AU3_0(.dout(w_dff_A_VJQGOMM76_0),.din(w_dff_A_YdYiZ7AU3_0),.clk(gclk));
	jdff dff_A_VJQGOMM76_0(.dout(w_dff_A_T7Z2gSsz2_0),.din(w_dff_A_VJQGOMM76_0),.clk(gclk));
	jdff dff_A_T7Z2gSsz2_0(.dout(w_dff_A_YTdbOB5J2_0),.din(w_dff_A_T7Z2gSsz2_0),.clk(gclk));
	jdff dff_A_YTdbOB5J2_0(.dout(w_dff_A_MRXlh1625_0),.din(w_dff_A_YTdbOB5J2_0),.clk(gclk));
	jdff dff_A_MRXlh1625_0(.dout(w_dff_A_dnbNaOuy9_0),.din(w_dff_A_MRXlh1625_0),.clk(gclk));
	jdff dff_A_dnbNaOuy9_0(.dout(w_dff_A_5193G9Ww8_0),.din(w_dff_A_dnbNaOuy9_0),.clk(gclk));
	jdff dff_A_5193G9Ww8_0(.dout(w_dff_A_5uSi0a8m7_0),.din(w_dff_A_5193G9Ww8_0),.clk(gclk));
	jdff dff_A_5uSi0a8m7_0(.dout(w_dff_A_SrWgg1V45_0),.din(w_dff_A_5uSi0a8m7_0),.clk(gclk));
	jdff dff_A_SrWgg1V45_0(.dout(w_dff_A_5J7euuBr6_0),.din(w_dff_A_SrWgg1V45_0),.clk(gclk));
	jdff dff_A_5J7euuBr6_0(.dout(w_dff_A_G5dtKGF12_0),.din(w_dff_A_5J7euuBr6_0),.clk(gclk));
	jdff dff_A_G5dtKGF12_0(.dout(w_dff_A_I4pNf0av5_0),.din(w_dff_A_G5dtKGF12_0),.clk(gclk));
	jdff dff_A_I4pNf0av5_0(.dout(f91),.din(w_dff_A_I4pNf0av5_0),.clk(gclk));
	jdff dff_A_AEzxCK512_2(.dout(w_dff_A_GG2qHrda8_0),.din(w_dff_A_AEzxCK512_2),.clk(gclk));
	jdff dff_A_GG2qHrda8_0(.dout(w_dff_A_HEMTRrbP5_0),.din(w_dff_A_GG2qHrda8_0),.clk(gclk));
	jdff dff_A_HEMTRrbP5_0(.dout(w_dff_A_pmoD3Ghc4_0),.din(w_dff_A_HEMTRrbP5_0),.clk(gclk));
	jdff dff_A_pmoD3Ghc4_0(.dout(w_dff_A_36qEBrI93_0),.din(w_dff_A_pmoD3Ghc4_0),.clk(gclk));
	jdff dff_A_36qEBrI93_0(.dout(w_dff_A_9zlPCw3b3_0),.din(w_dff_A_36qEBrI93_0),.clk(gclk));
	jdff dff_A_9zlPCw3b3_0(.dout(w_dff_A_DjsrlyfB3_0),.din(w_dff_A_9zlPCw3b3_0),.clk(gclk));
	jdff dff_A_DjsrlyfB3_0(.dout(w_dff_A_ZKoYZQew1_0),.din(w_dff_A_DjsrlyfB3_0),.clk(gclk));
	jdff dff_A_ZKoYZQew1_0(.dout(w_dff_A_O0lCVhFz5_0),.din(w_dff_A_ZKoYZQew1_0),.clk(gclk));
	jdff dff_A_O0lCVhFz5_0(.dout(w_dff_A_7ZLbmI1O3_0),.din(w_dff_A_O0lCVhFz5_0),.clk(gclk));
	jdff dff_A_7ZLbmI1O3_0(.dout(w_dff_A_2ZrH3l2z6_0),.din(w_dff_A_7ZLbmI1O3_0),.clk(gclk));
	jdff dff_A_2ZrH3l2z6_0(.dout(w_dff_A_y4bBXwF59_0),.din(w_dff_A_2ZrH3l2z6_0),.clk(gclk));
	jdff dff_A_y4bBXwF59_0(.dout(w_dff_A_5EqS5cp89_0),.din(w_dff_A_y4bBXwF59_0),.clk(gclk));
	jdff dff_A_5EqS5cp89_0(.dout(w_dff_A_pqyHQPTf7_0),.din(w_dff_A_5EqS5cp89_0),.clk(gclk));
	jdff dff_A_pqyHQPTf7_0(.dout(w_dff_A_ZGXGSGaI8_0),.din(w_dff_A_pqyHQPTf7_0),.clk(gclk));
	jdff dff_A_ZGXGSGaI8_0(.dout(w_dff_A_kk8aeY6D9_0),.din(w_dff_A_ZGXGSGaI8_0),.clk(gclk));
	jdff dff_A_kk8aeY6D9_0(.dout(w_dff_A_Ym6T1lWP5_0),.din(w_dff_A_kk8aeY6D9_0),.clk(gclk));
	jdff dff_A_Ym6T1lWP5_0(.dout(w_dff_A_GMReuTzS9_0),.din(w_dff_A_Ym6T1lWP5_0),.clk(gclk));
	jdff dff_A_GMReuTzS9_0(.dout(w_dff_A_xCHzNYns4_0),.din(w_dff_A_GMReuTzS9_0),.clk(gclk));
	jdff dff_A_xCHzNYns4_0(.dout(w_dff_A_Y0viZO0d2_0),.din(w_dff_A_xCHzNYns4_0),.clk(gclk));
	jdff dff_A_Y0viZO0d2_0(.dout(w_dff_A_PGTCaPkD5_0),.din(w_dff_A_Y0viZO0d2_0),.clk(gclk));
	jdff dff_A_PGTCaPkD5_0(.dout(w_dff_A_FR07CoQ79_0),.din(w_dff_A_PGTCaPkD5_0),.clk(gclk));
	jdff dff_A_FR07CoQ79_0(.dout(w_dff_A_tRN7QY4J8_0),.din(w_dff_A_FR07CoQ79_0),.clk(gclk));
	jdff dff_A_tRN7QY4J8_0(.dout(w_dff_A_sOqrwEUk5_0),.din(w_dff_A_tRN7QY4J8_0),.clk(gclk));
	jdff dff_A_sOqrwEUk5_0(.dout(w_dff_A_FEnRIYzi5_0),.din(w_dff_A_sOqrwEUk5_0),.clk(gclk));
	jdff dff_A_FEnRIYzi5_0(.dout(w_dff_A_gVW96HaF4_0),.din(w_dff_A_FEnRIYzi5_0),.clk(gclk));
	jdff dff_A_gVW96HaF4_0(.dout(w_dff_A_3VGk58dE0_0),.din(w_dff_A_gVW96HaF4_0),.clk(gclk));
	jdff dff_A_3VGk58dE0_0(.dout(w_dff_A_KSIjEYaI7_0),.din(w_dff_A_3VGk58dE0_0),.clk(gclk));
	jdff dff_A_KSIjEYaI7_0(.dout(w_dff_A_uAg23j1w9_0),.din(w_dff_A_KSIjEYaI7_0),.clk(gclk));
	jdff dff_A_uAg23j1w9_0(.dout(w_dff_A_4Q9byydA5_0),.din(w_dff_A_uAg23j1w9_0),.clk(gclk));
	jdff dff_A_4Q9byydA5_0(.dout(w_dff_A_2vk2danU6_0),.din(w_dff_A_4Q9byydA5_0),.clk(gclk));
	jdff dff_A_2vk2danU6_0(.dout(w_dff_A_xFJkBUed9_0),.din(w_dff_A_2vk2danU6_0),.clk(gclk));
	jdff dff_A_xFJkBUed9_0(.dout(w_dff_A_bTMQQsJo4_0),.din(w_dff_A_xFJkBUed9_0),.clk(gclk));
	jdff dff_A_bTMQQsJo4_0(.dout(w_dff_A_gfT7eHZK6_0),.din(w_dff_A_bTMQQsJo4_0),.clk(gclk));
	jdff dff_A_gfT7eHZK6_0(.dout(w_dff_A_ha7sRvCT7_0),.din(w_dff_A_gfT7eHZK6_0),.clk(gclk));
	jdff dff_A_ha7sRvCT7_0(.dout(f92),.din(w_dff_A_ha7sRvCT7_0),.clk(gclk));
	jdff dff_A_Er2L8DHW9_2(.dout(w_dff_A_s0FhXH485_0),.din(w_dff_A_Er2L8DHW9_2),.clk(gclk));
	jdff dff_A_s0FhXH485_0(.dout(w_dff_A_H3KxTAOp2_0),.din(w_dff_A_s0FhXH485_0),.clk(gclk));
	jdff dff_A_H3KxTAOp2_0(.dout(w_dff_A_q4vYkGNi5_0),.din(w_dff_A_H3KxTAOp2_0),.clk(gclk));
	jdff dff_A_q4vYkGNi5_0(.dout(w_dff_A_27hEjulX3_0),.din(w_dff_A_q4vYkGNi5_0),.clk(gclk));
	jdff dff_A_27hEjulX3_0(.dout(w_dff_A_tm4LvgA97_0),.din(w_dff_A_27hEjulX3_0),.clk(gclk));
	jdff dff_A_tm4LvgA97_0(.dout(w_dff_A_LcTWEY0y3_0),.din(w_dff_A_tm4LvgA97_0),.clk(gclk));
	jdff dff_A_LcTWEY0y3_0(.dout(w_dff_A_dhjZMPjj6_0),.din(w_dff_A_LcTWEY0y3_0),.clk(gclk));
	jdff dff_A_dhjZMPjj6_0(.dout(w_dff_A_nAhy8jg97_0),.din(w_dff_A_dhjZMPjj6_0),.clk(gclk));
	jdff dff_A_nAhy8jg97_0(.dout(w_dff_A_iZ0FBQ177_0),.din(w_dff_A_nAhy8jg97_0),.clk(gclk));
	jdff dff_A_iZ0FBQ177_0(.dout(w_dff_A_C74O2baP2_0),.din(w_dff_A_iZ0FBQ177_0),.clk(gclk));
	jdff dff_A_C74O2baP2_0(.dout(w_dff_A_gurycyko8_0),.din(w_dff_A_C74O2baP2_0),.clk(gclk));
	jdff dff_A_gurycyko8_0(.dout(w_dff_A_5hlrvbOy0_0),.din(w_dff_A_gurycyko8_0),.clk(gclk));
	jdff dff_A_5hlrvbOy0_0(.dout(w_dff_A_HLpD1Wbu2_0),.din(w_dff_A_5hlrvbOy0_0),.clk(gclk));
	jdff dff_A_HLpD1Wbu2_0(.dout(w_dff_A_wFI9jBks7_0),.din(w_dff_A_HLpD1Wbu2_0),.clk(gclk));
	jdff dff_A_wFI9jBks7_0(.dout(w_dff_A_jVyFTlLG6_0),.din(w_dff_A_wFI9jBks7_0),.clk(gclk));
	jdff dff_A_jVyFTlLG6_0(.dout(w_dff_A_mVbs1mQK4_0),.din(w_dff_A_jVyFTlLG6_0),.clk(gclk));
	jdff dff_A_mVbs1mQK4_0(.dout(w_dff_A_QlmCQiEH4_0),.din(w_dff_A_mVbs1mQK4_0),.clk(gclk));
	jdff dff_A_QlmCQiEH4_0(.dout(w_dff_A_L6KSNkEp9_0),.din(w_dff_A_QlmCQiEH4_0),.clk(gclk));
	jdff dff_A_L6KSNkEp9_0(.dout(w_dff_A_j7CXxbfw8_0),.din(w_dff_A_L6KSNkEp9_0),.clk(gclk));
	jdff dff_A_j7CXxbfw8_0(.dout(w_dff_A_ZtrqJAz43_0),.din(w_dff_A_j7CXxbfw8_0),.clk(gclk));
	jdff dff_A_ZtrqJAz43_0(.dout(w_dff_A_RsvUncEq5_0),.din(w_dff_A_ZtrqJAz43_0),.clk(gclk));
	jdff dff_A_RsvUncEq5_0(.dout(w_dff_A_0pkwwZBt8_0),.din(w_dff_A_RsvUncEq5_0),.clk(gclk));
	jdff dff_A_0pkwwZBt8_0(.dout(w_dff_A_VpJKZxxq4_0),.din(w_dff_A_0pkwwZBt8_0),.clk(gclk));
	jdff dff_A_VpJKZxxq4_0(.dout(w_dff_A_c7ULtHPb4_0),.din(w_dff_A_VpJKZxxq4_0),.clk(gclk));
	jdff dff_A_c7ULtHPb4_0(.dout(w_dff_A_J6zzYJr99_0),.din(w_dff_A_c7ULtHPb4_0),.clk(gclk));
	jdff dff_A_J6zzYJr99_0(.dout(w_dff_A_fEDCAqdp5_0),.din(w_dff_A_J6zzYJr99_0),.clk(gclk));
	jdff dff_A_fEDCAqdp5_0(.dout(w_dff_A_jJz3Byz79_0),.din(w_dff_A_fEDCAqdp5_0),.clk(gclk));
	jdff dff_A_jJz3Byz79_0(.dout(w_dff_A_6ccVvoid0_0),.din(w_dff_A_jJz3Byz79_0),.clk(gclk));
	jdff dff_A_6ccVvoid0_0(.dout(w_dff_A_xNjEQSO61_0),.din(w_dff_A_6ccVvoid0_0),.clk(gclk));
	jdff dff_A_xNjEQSO61_0(.dout(w_dff_A_uLE9o1bl6_0),.din(w_dff_A_xNjEQSO61_0),.clk(gclk));
	jdff dff_A_uLE9o1bl6_0(.dout(w_dff_A_OeLNR1lA4_0),.din(w_dff_A_uLE9o1bl6_0),.clk(gclk));
	jdff dff_A_OeLNR1lA4_0(.dout(w_dff_A_yQAACRrt1_0),.din(w_dff_A_OeLNR1lA4_0),.clk(gclk));
	jdff dff_A_yQAACRrt1_0(.dout(w_dff_A_GteC1O896_0),.din(w_dff_A_yQAACRrt1_0),.clk(gclk));
	jdff dff_A_GteC1O896_0(.dout(f93),.din(w_dff_A_GteC1O896_0),.clk(gclk));
	jdff dff_A_XtJDEDOj6_2(.dout(w_dff_A_OyFx5A880_0),.din(w_dff_A_XtJDEDOj6_2),.clk(gclk));
	jdff dff_A_OyFx5A880_0(.dout(w_dff_A_KOaYgp0D9_0),.din(w_dff_A_OyFx5A880_0),.clk(gclk));
	jdff dff_A_KOaYgp0D9_0(.dout(w_dff_A_nkgGLMtD9_0),.din(w_dff_A_KOaYgp0D9_0),.clk(gclk));
	jdff dff_A_nkgGLMtD9_0(.dout(w_dff_A_IaiFbMsq2_0),.din(w_dff_A_nkgGLMtD9_0),.clk(gclk));
	jdff dff_A_IaiFbMsq2_0(.dout(w_dff_A_hiH3E2K55_0),.din(w_dff_A_IaiFbMsq2_0),.clk(gclk));
	jdff dff_A_hiH3E2K55_0(.dout(w_dff_A_nFdgBBVX7_0),.din(w_dff_A_hiH3E2K55_0),.clk(gclk));
	jdff dff_A_nFdgBBVX7_0(.dout(w_dff_A_f7KippQH5_0),.din(w_dff_A_nFdgBBVX7_0),.clk(gclk));
	jdff dff_A_f7KippQH5_0(.dout(w_dff_A_jZCayZcU5_0),.din(w_dff_A_f7KippQH5_0),.clk(gclk));
	jdff dff_A_jZCayZcU5_0(.dout(w_dff_A_EnygtvhL5_0),.din(w_dff_A_jZCayZcU5_0),.clk(gclk));
	jdff dff_A_EnygtvhL5_0(.dout(w_dff_A_pTJ5ZJAZ3_0),.din(w_dff_A_EnygtvhL5_0),.clk(gclk));
	jdff dff_A_pTJ5ZJAZ3_0(.dout(w_dff_A_V6FZ53R40_0),.din(w_dff_A_pTJ5ZJAZ3_0),.clk(gclk));
	jdff dff_A_V6FZ53R40_0(.dout(w_dff_A_g6SGFTmx0_0),.din(w_dff_A_V6FZ53R40_0),.clk(gclk));
	jdff dff_A_g6SGFTmx0_0(.dout(w_dff_A_wv7Zd7jA2_0),.din(w_dff_A_g6SGFTmx0_0),.clk(gclk));
	jdff dff_A_wv7Zd7jA2_0(.dout(w_dff_A_0DkXz5Rp1_0),.din(w_dff_A_wv7Zd7jA2_0),.clk(gclk));
	jdff dff_A_0DkXz5Rp1_0(.dout(w_dff_A_R4ehAkps4_0),.din(w_dff_A_0DkXz5Rp1_0),.clk(gclk));
	jdff dff_A_R4ehAkps4_0(.dout(w_dff_A_wHPL78TD7_0),.din(w_dff_A_R4ehAkps4_0),.clk(gclk));
	jdff dff_A_wHPL78TD7_0(.dout(w_dff_A_wjbkuumn2_0),.din(w_dff_A_wHPL78TD7_0),.clk(gclk));
	jdff dff_A_wjbkuumn2_0(.dout(w_dff_A_87Lomuc35_0),.din(w_dff_A_wjbkuumn2_0),.clk(gclk));
	jdff dff_A_87Lomuc35_0(.dout(w_dff_A_TemNoxqc6_0),.din(w_dff_A_87Lomuc35_0),.clk(gclk));
	jdff dff_A_TemNoxqc6_0(.dout(w_dff_A_6feuHVrJ0_0),.din(w_dff_A_TemNoxqc6_0),.clk(gclk));
	jdff dff_A_6feuHVrJ0_0(.dout(w_dff_A_0G0vAa8i2_0),.din(w_dff_A_6feuHVrJ0_0),.clk(gclk));
	jdff dff_A_0G0vAa8i2_0(.dout(w_dff_A_AHCT5n9d5_0),.din(w_dff_A_0G0vAa8i2_0),.clk(gclk));
	jdff dff_A_AHCT5n9d5_0(.dout(w_dff_A_mTbdqkSx3_0),.din(w_dff_A_AHCT5n9d5_0),.clk(gclk));
	jdff dff_A_mTbdqkSx3_0(.dout(w_dff_A_nrZDo8Ng2_0),.din(w_dff_A_mTbdqkSx3_0),.clk(gclk));
	jdff dff_A_nrZDo8Ng2_0(.dout(w_dff_A_ftSEOCsG1_0),.din(w_dff_A_nrZDo8Ng2_0),.clk(gclk));
	jdff dff_A_ftSEOCsG1_0(.dout(w_dff_A_FNAR7OHg0_0),.din(w_dff_A_ftSEOCsG1_0),.clk(gclk));
	jdff dff_A_FNAR7OHg0_0(.dout(w_dff_A_i2sXLfoG6_0),.din(w_dff_A_FNAR7OHg0_0),.clk(gclk));
	jdff dff_A_i2sXLfoG6_0(.dout(w_dff_A_Ib8X9Dm93_0),.din(w_dff_A_i2sXLfoG6_0),.clk(gclk));
	jdff dff_A_Ib8X9Dm93_0(.dout(w_dff_A_4iLw99K71_0),.din(w_dff_A_Ib8X9Dm93_0),.clk(gclk));
	jdff dff_A_4iLw99K71_0(.dout(w_dff_A_HOt6GUvs5_0),.din(w_dff_A_4iLw99K71_0),.clk(gclk));
	jdff dff_A_HOt6GUvs5_0(.dout(w_dff_A_3NTiZ3Yi6_0),.din(w_dff_A_HOt6GUvs5_0),.clk(gclk));
	jdff dff_A_3NTiZ3Yi6_0(.dout(w_dff_A_RFD5YmZp0_0),.din(w_dff_A_3NTiZ3Yi6_0),.clk(gclk));
	jdff dff_A_RFD5YmZp0_0(.dout(f94),.din(w_dff_A_RFD5YmZp0_0),.clk(gclk));
	jdff dff_A_AMFRU9o10_2(.dout(w_dff_A_jIVhXD069_0),.din(w_dff_A_AMFRU9o10_2),.clk(gclk));
	jdff dff_A_jIVhXD069_0(.dout(w_dff_A_yTp6qN5W8_0),.din(w_dff_A_jIVhXD069_0),.clk(gclk));
	jdff dff_A_yTp6qN5W8_0(.dout(w_dff_A_1zUFLRwG2_0),.din(w_dff_A_yTp6qN5W8_0),.clk(gclk));
	jdff dff_A_1zUFLRwG2_0(.dout(w_dff_A_VwrrkvWe2_0),.din(w_dff_A_1zUFLRwG2_0),.clk(gclk));
	jdff dff_A_VwrrkvWe2_0(.dout(w_dff_A_sfB2jh6E7_0),.din(w_dff_A_VwrrkvWe2_0),.clk(gclk));
	jdff dff_A_sfB2jh6E7_0(.dout(w_dff_A_CBgQENVl6_0),.din(w_dff_A_sfB2jh6E7_0),.clk(gclk));
	jdff dff_A_CBgQENVl6_0(.dout(w_dff_A_5sg1HbME6_0),.din(w_dff_A_CBgQENVl6_0),.clk(gclk));
	jdff dff_A_5sg1HbME6_0(.dout(w_dff_A_x8ExOody9_0),.din(w_dff_A_5sg1HbME6_0),.clk(gclk));
	jdff dff_A_x8ExOody9_0(.dout(w_dff_A_21NfC90x9_0),.din(w_dff_A_x8ExOody9_0),.clk(gclk));
	jdff dff_A_21NfC90x9_0(.dout(w_dff_A_qfCcvu7Y4_0),.din(w_dff_A_21NfC90x9_0),.clk(gclk));
	jdff dff_A_qfCcvu7Y4_0(.dout(w_dff_A_c6jxBjna5_0),.din(w_dff_A_qfCcvu7Y4_0),.clk(gclk));
	jdff dff_A_c6jxBjna5_0(.dout(w_dff_A_iGWbQu3n5_0),.din(w_dff_A_c6jxBjna5_0),.clk(gclk));
	jdff dff_A_iGWbQu3n5_0(.dout(w_dff_A_FmNSV9Zc5_0),.din(w_dff_A_iGWbQu3n5_0),.clk(gclk));
	jdff dff_A_FmNSV9Zc5_0(.dout(w_dff_A_pzOzmHdQ2_0),.din(w_dff_A_FmNSV9Zc5_0),.clk(gclk));
	jdff dff_A_pzOzmHdQ2_0(.dout(w_dff_A_OEUCuBTl8_0),.din(w_dff_A_pzOzmHdQ2_0),.clk(gclk));
	jdff dff_A_OEUCuBTl8_0(.dout(w_dff_A_wkWBZRef1_0),.din(w_dff_A_OEUCuBTl8_0),.clk(gclk));
	jdff dff_A_wkWBZRef1_0(.dout(w_dff_A_Fdfb4myi2_0),.din(w_dff_A_wkWBZRef1_0),.clk(gclk));
	jdff dff_A_Fdfb4myi2_0(.dout(w_dff_A_xBzxjasY5_0),.din(w_dff_A_Fdfb4myi2_0),.clk(gclk));
	jdff dff_A_xBzxjasY5_0(.dout(w_dff_A_K9CmqhHe0_0),.din(w_dff_A_xBzxjasY5_0),.clk(gclk));
	jdff dff_A_K9CmqhHe0_0(.dout(w_dff_A_mVI6TKSg5_0),.din(w_dff_A_K9CmqhHe0_0),.clk(gclk));
	jdff dff_A_mVI6TKSg5_0(.dout(w_dff_A_REjKV5va8_0),.din(w_dff_A_mVI6TKSg5_0),.clk(gclk));
	jdff dff_A_REjKV5va8_0(.dout(w_dff_A_gIuKOqEl3_0),.din(w_dff_A_REjKV5va8_0),.clk(gclk));
	jdff dff_A_gIuKOqEl3_0(.dout(w_dff_A_Z2OHPcQM9_0),.din(w_dff_A_gIuKOqEl3_0),.clk(gclk));
	jdff dff_A_Z2OHPcQM9_0(.dout(w_dff_A_exWGyCCJ8_0),.din(w_dff_A_Z2OHPcQM9_0),.clk(gclk));
	jdff dff_A_exWGyCCJ8_0(.dout(w_dff_A_0CUD4K4l6_0),.din(w_dff_A_exWGyCCJ8_0),.clk(gclk));
	jdff dff_A_0CUD4K4l6_0(.dout(w_dff_A_Pb8O3KwZ2_0),.din(w_dff_A_0CUD4K4l6_0),.clk(gclk));
	jdff dff_A_Pb8O3KwZ2_0(.dout(w_dff_A_9bxlpSS61_0),.din(w_dff_A_Pb8O3KwZ2_0),.clk(gclk));
	jdff dff_A_9bxlpSS61_0(.dout(w_dff_A_CCJJUVgd2_0),.din(w_dff_A_9bxlpSS61_0),.clk(gclk));
	jdff dff_A_CCJJUVgd2_0(.dout(w_dff_A_2Xvt5aW23_0),.din(w_dff_A_CCJJUVgd2_0),.clk(gclk));
	jdff dff_A_2Xvt5aW23_0(.dout(w_dff_A_ZOVD3b5g5_0),.din(w_dff_A_2Xvt5aW23_0),.clk(gclk));
	jdff dff_A_ZOVD3b5g5_0(.dout(w_dff_A_TlgeE8eC6_0),.din(w_dff_A_ZOVD3b5g5_0),.clk(gclk));
	jdff dff_A_TlgeE8eC6_0(.dout(f95),.din(w_dff_A_TlgeE8eC6_0),.clk(gclk));
	jdff dff_A_4HZtpbSH1_2(.dout(w_dff_A_OzbBedJb7_0),.din(w_dff_A_4HZtpbSH1_2),.clk(gclk));
	jdff dff_A_OzbBedJb7_0(.dout(w_dff_A_1MTZhLHc1_0),.din(w_dff_A_OzbBedJb7_0),.clk(gclk));
	jdff dff_A_1MTZhLHc1_0(.dout(w_dff_A_ne1HhVGo4_0),.din(w_dff_A_1MTZhLHc1_0),.clk(gclk));
	jdff dff_A_ne1HhVGo4_0(.dout(w_dff_A_9qr5Z93a6_0),.din(w_dff_A_ne1HhVGo4_0),.clk(gclk));
	jdff dff_A_9qr5Z93a6_0(.dout(w_dff_A_RjQ5wP8l1_0),.din(w_dff_A_9qr5Z93a6_0),.clk(gclk));
	jdff dff_A_RjQ5wP8l1_0(.dout(w_dff_A_4wBtinSQ2_0),.din(w_dff_A_RjQ5wP8l1_0),.clk(gclk));
	jdff dff_A_4wBtinSQ2_0(.dout(w_dff_A_8OhVbW7t9_0),.din(w_dff_A_4wBtinSQ2_0),.clk(gclk));
	jdff dff_A_8OhVbW7t9_0(.dout(w_dff_A_x0TcEQ1t1_0),.din(w_dff_A_8OhVbW7t9_0),.clk(gclk));
	jdff dff_A_x0TcEQ1t1_0(.dout(w_dff_A_E17ZPpId0_0),.din(w_dff_A_x0TcEQ1t1_0),.clk(gclk));
	jdff dff_A_E17ZPpId0_0(.dout(w_dff_A_T6bTbsre6_0),.din(w_dff_A_E17ZPpId0_0),.clk(gclk));
	jdff dff_A_T6bTbsre6_0(.dout(w_dff_A_m5mqXB9Y0_0),.din(w_dff_A_T6bTbsre6_0),.clk(gclk));
	jdff dff_A_m5mqXB9Y0_0(.dout(w_dff_A_QtfUI3C00_0),.din(w_dff_A_m5mqXB9Y0_0),.clk(gclk));
	jdff dff_A_QtfUI3C00_0(.dout(w_dff_A_TF6lvV6v0_0),.din(w_dff_A_QtfUI3C00_0),.clk(gclk));
	jdff dff_A_TF6lvV6v0_0(.dout(w_dff_A_WUOT6sek2_0),.din(w_dff_A_TF6lvV6v0_0),.clk(gclk));
	jdff dff_A_WUOT6sek2_0(.dout(w_dff_A_Cvgxm6IG7_0),.din(w_dff_A_WUOT6sek2_0),.clk(gclk));
	jdff dff_A_Cvgxm6IG7_0(.dout(w_dff_A_lC7hgAga4_0),.din(w_dff_A_Cvgxm6IG7_0),.clk(gclk));
	jdff dff_A_lC7hgAga4_0(.dout(w_dff_A_dqssucrA4_0),.din(w_dff_A_lC7hgAga4_0),.clk(gclk));
	jdff dff_A_dqssucrA4_0(.dout(w_dff_A_h5Ade49L3_0),.din(w_dff_A_dqssucrA4_0),.clk(gclk));
	jdff dff_A_h5Ade49L3_0(.dout(w_dff_A_bllbTu639_0),.din(w_dff_A_h5Ade49L3_0),.clk(gclk));
	jdff dff_A_bllbTu639_0(.dout(w_dff_A_WPcbLUlv7_0),.din(w_dff_A_bllbTu639_0),.clk(gclk));
	jdff dff_A_WPcbLUlv7_0(.dout(w_dff_A_WezhJCRD5_0),.din(w_dff_A_WPcbLUlv7_0),.clk(gclk));
	jdff dff_A_WezhJCRD5_0(.dout(w_dff_A_TPZG4tmn1_0),.din(w_dff_A_WezhJCRD5_0),.clk(gclk));
	jdff dff_A_TPZG4tmn1_0(.dout(w_dff_A_AH40itoX9_0),.din(w_dff_A_TPZG4tmn1_0),.clk(gclk));
	jdff dff_A_AH40itoX9_0(.dout(w_dff_A_FbErS4Kj5_0),.din(w_dff_A_AH40itoX9_0),.clk(gclk));
	jdff dff_A_FbErS4Kj5_0(.dout(w_dff_A_oEym1vmV9_0),.din(w_dff_A_FbErS4Kj5_0),.clk(gclk));
	jdff dff_A_oEym1vmV9_0(.dout(w_dff_A_wOnsUkqY4_0),.din(w_dff_A_oEym1vmV9_0),.clk(gclk));
	jdff dff_A_wOnsUkqY4_0(.dout(w_dff_A_U8Ri4lTr6_0),.din(w_dff_A_wOnsUkqY4_0),.clk(gclk));
	jdff dff_A_U8Ri4lTr6_0(.dout(w_dff_A_5ToOps0K2_0),.din(w_dff_A_U8Ri4lTr6_0),.clk(gclk));
	jdff dff_A_5ToOps0K2_0(.dout(w_dff_A_A1O5LbtV9_0),.din(w_dff_A_5ToOps0K2_0),.clk(gclk));
	jdff dff_A_A1O5LbtV9_0(.dout(w_dff_A_5SZGfYla9_0),.din(w_dff_A_A1O5LbtV9_0),.clk(gclk));
	jdff dff_A_5SZGfYla9_0(.dout(f96),.din(w_dff_A_5SZGfYla9_0),.clk(gclk));
	jdff dff_A_LhBO705X1_2(.dout(w_dff_A_zEpGsihP7_0),.din(w_dff_A_LhBO705X1_2),.clk(gclk));
	jdff dff_A_zEpGsihP7_0(.dout(w_dff_A_WRML9YSR7_0),.din(w_dff_A_zEpGsihP7_0),.clk(gclk));
	jdff dff_A_WRML9YSR7_0(.dout(w_dff_A_EbMEZZh34_0),.din(w_dff_A_WRML9YSR7_0),.clk(gclk));
	jdff dff_A_EbMEZZh34_0(.dout(w_dff_A_Jv1ane812_0),.din(w_dff_A_EbMEZZh34_0),.clk(gclk));
	jdff dff_A_Jv1ane812_0(.dout(w_dff_A_0NHjkmcn2_0),.din(w_dff_A_Jv1ane812_0),.clk(gclk));
	jdff dff_A_0NHjkmcn2_0(.dout(w_dff_A_S8x0eCf48_0),.din(w_dff_A_0NHjkmcn2_0),.clk(gclk));
	jdff dff_A_S8x0eCf48_0(.dout(w_dff_A_m7EI7u6d7_0),.din(w_dff_A_S8x0eCf48_0),.clk(gclk));
	jdff dff_A_m7EI7u6d7_0(.dout(w_dff_A_0kqtpuMh4_0),.din(w_dff_A_m7EI7u6d7_0),.clk(gclk));
	jdff dff_A_0kqtpuMh4_0(.dout(w_dff_A_YOIchtsx3_0),.din(w_dff_A_0kqtpuMh4_0),.clk(gclk));
	jdff dff_A_YOIchtsx3_0(.dout(w_dff_A_RJ6aH9HW3_0),.din(w_dff_A_YOIchtsx3_0),.clk(gclk));
	jdff dff_A_RJ6aH9HW3_0(.dout(w_dff_A_ykMiWOmd7_0),.din(w_dff_A_RJ6aH9HW3_0),.clk(gclk));
	jdff dff_A_ykMiWOmd7_0(.dout(w_dff_A_r9vIpNX69_0),.din(w_dff_A_ykMiWOmd7_0),.clk(gclk));
	jdff dff_A_r9vIpNX69_0(.dout(w_dff_A_zdj4RMZp5_0),.din(w_dff_A_r9vIpNX69_0),.clk(gclk));
	jdff dff_A_zdj4RMZp5_0(.dout(w_dff_A_Uz5G1Hr18_0),.din(w_dff_A_zdj4RMZp5_0),.clk(gclk));
	jdff dff_A_Uz5G1Hr18_0(.dout(w_dff_A_BvBDuFQC5_0),.din(w_dff_A_Uz5G1Hr18_0),.clk(gclk));
	jdff dff_A_BvBDuFQC5_0(.dout(w_dff_A_H1k3tpQC5_0),.din(w_dff_A_BvBDuFQC5_0),.clk(gclk));
	jdff dff_A_H1k3tpQC5_0(.dout(w_dff_A_NR8wCoVQ3_0),.din(w_dff_A_H1k3tpQC5_0),.clk(gclk));
	jdff dff_A_NR8wCoVQ3_0(.dout(w_dff_A_SOJoO6kf2_0),.din(w_dff_A_NR8wCoVQ3_0),.clk(gclk));
	jdff dff_A_SOJoO6kf2_0(.dout(w_dff_A_w2pwQ2km1_0),.din(w_dff_A_SOJoO6kf2_0),.clk(gclk));
	jdff dff_A_w2pwQ2km1_0(.dout(w_dff_A_iKLN3hkd6_0),.din(w_dff_A_w2pwQ2km1_0),.clk(gclk));
	jdff dff_A_iKLN3hkd6_0(.dout(w_dff_A_oYLQsRHv3_0),.din(w_dff_A_iKLN3hkd6_0),.clk(gclk));
	jdff dff_A_oYLQsRHv3_0(.dout(w_dff_A_uL5O8sbb5_0),.din(w_dff_A_oYLQsRHv3_0),.clk(gclk));
	jdff dff_A_uL5O8sbb5_0(.dout(w_dff_A_Aurm1clF5_0),.din(w_dff_A_uL5O8sbb5_0),.clk(gclk));
	jdff dff_A_Aurm1clF5_0(.dout(w_dff_A_mUpL9pL13_0),.din(w_dff_A_Aurm1clF5_0),.clk(gclk));
	jdff dff_A_mUpL9pL13_0(.dout(w_dff_A_RrdZ3eil9_0),.din(w_dff_A_mUpL9pL13_0),.clk(gclk));
	jdff dff_A_RrdZ3eil9_0(.dout(w_dff_A_cseoMQNJ7_0),.din(w_dff_A_RrdZ3eil9_0),.clk(gclk));
	jdff dff_A_cseoMQNJ7_0(.dout(w_dff_A_tllxPUpK9_0),.din(w_dff_A_cseoMQNJ7_0),.clk(gclk));
	jdff dff_A_tllxPUpK9_0(.dout(w_dff_A_AWDRmoyb0_0),.din(w_dff_A_tllxPUpK9_0),.clk(gclk));
	jdff dff_A_AWDRmoyb0_0(.dout(w_dff_A_re7SjTjq8_0),.din(w_dff_A_AWDRmoyb0_0),.clk(gclk));
	jdff dff_A_re7SjTjq8_0(.dout(f97),.din(w_dff_A_re7SjTjq8_0),.clk(gclk));
	jdff dff_A_rQuWRbM25_2(.dout(w_dff_A_sAQW3IEU1_0),.din(w_dff_A_rQuWRbM25_2),.clk(gclk));
	jdff dff_A_sAQW3IEU1_0(.dout(w_dff_A_p3eE2AWL6_0),.din(w_dff_A_sAQW3IEU1_0),.clk(gclk));
	jdff dff_A_p3eE2AWL6_0(.dout(w_dff_A_BMLHg5pi6_0),.din(w_dff_A_p3eE2AWL6_0),.clk(gclk));
	jdff dff_A_BMLHg5pi6_0(.dout(w_dff_A_3LVBQ0Pl4_0),.din(w_dff_A_BMLHg5pi6_0),.clk(gclk));
	jdff dff_A_3LVBQ0Pl4_0(.dout(w_dff_A_Dotap0Un6_0),.din(w_dff_A_3LVBQ0Pl4_0),.clk(gclk));
	jdff dff_A_Dotap0Un6_0(.dout(w_dff_A_1AchSSIF2_0),.din(w_dff_A_Dotap0Un6_0),.clk(gclk));
	jdff dff_A_1AchSSIF2_0(.dout(w_dff_A_3f3b0Iid8_0),.din(w_dff_A_1AchSSIF2_0),.clk(gclk));
	jdff dff_A_3f3b0Iid8_0(.dout(w_dff_A_7QRDJune4_0),.din(w_dff_A_3f3b0Iid8_0),.clk(gclk));
	jdff dff_A_7QRDJune4_0(.dout(w_dff_A_82QO3kuO9_0),.din(w_dff_A_7QRDJune4_0),.clk(gclk));
	jdff dff_A_82QO3kuO9_0(.dout(w_dff_A_5NcD73wh4_0),.din(w_dff_A_82QO3kuO9_0),.clk(gclk));
	jdff dff_A_5NcD73wh4_0(.dout(w_dff_A_hY5JxQdx9_0),.din(w_dff_A_5NcD73wh4_0),.clk(gclk));
	jdff dff_A_hY5JxQdx9_0(.dout(w_dff_A_trFWKzSG7_0),.din(w_dff_A_hY5JxQdx9_0),.clk(gclk));
	jdff dff_A_trFWKzSG7_0(.dout(w_dff_A_TCrAfWY33_0),.din(w_dff_A_trFWKzSG7_0),.clk(gclk));
	jdff dff_A_TCrAfWY33_0(.dout(w_dff_A_Y5x0x0nm7_0),.din(w_dff_A_TCrAfWY33_0),.clk(gclk));
	jdff dff_A_Y5x0x0nm7_0(.dout(w_dff_A_QNGsPW584_0),.din(w_dff_A_Y5x0x0nm7_0),.clk(gclk));
	jdff dff_A_QNGsPW584_0(.dout(w_dff_A_LoSkd3Sz7_0),.din(w_dff_A_QNGsPW584_0),.clk(gclk));
	jdff dff_A_LoSkd3Sz7_0(.dout(w_dff_A_BWZex2k27_0),.din(w_dff_A_LoSkd3Sz7_0),.clk(gclk));
	jdff dff_A_BWZex2k27_0(.dout(w_dff_A_ho1eOfeC8_0),.din(w_dff_A_BWZex2k27_0),.clk(gclk));
	jdff dff_A_ho1eOfeC8_0(.dout(w_dff_A_qd6suzrS7_0),.din(w_dff_A_ho1eOfeC8_0),.clk(gclk));
	jdff dff_A_qd6suzrS7_0(.dout(w_dff_A_Jw6s70ey5_0),.din(w_dff_A_qd6suzrS7_0),.clk(gclk));
	jdff dff_A_Jw6s70ey5_0(.dout(w_dff_A_cDA7P9sQ0_0),.din(w_dff_A_Jw6s70ey5_0),.clk(gclk));
	jdff dff_A_cDA7P9sQ0_0(.dout(w_dff_A_ZUoVrhUy8_0),.din(w_dff_A_cDA7P9sQ0_0),.clk(gclk));
	jdff dff_A_ZUoVrhUy8_0(.dout(w_dff_A_WYcXydrp6_0),.din(w_dff_A_ZUoVrhUy8_0),.clk(gclk));
	jdff dff_A_WYcXydrp6_0(.dout(w_dff_A_UqF2f45e4_0),.din(w_dff_A_WYcXydrp6_0),.clk(gclk));
	jdff dff_A_UqF2f45e4_0(.dout(w_dff_A_052u7nYm7_0),.din(w_dff_A_UqF2f45e4_0),.clk(gclk));
	jdff dff_A_052u7nYm7_0(.dout(w_dff_A_m1kegvqW0_0),.din(w_dff_A_052u7nYm7_0),.clk(gclk));
	jdff dff_A_m1kegvqW0_0(.dout(w_dff_A_XYL7coZp0_0),.din(w_dff_A_m1kegvqW0_0),.clk(gclk));
	jdff dff_A_XYL7coZp0_0(.dout(w_dff_A_xdsG2och5_0),.din(w_dff_A_XYL7coZp0_0),.clk(gclk));
	jdff dff_A_xdsG2och5_0(.dout(f98),.din(w_dff_A_xdsG2och5_0),.clk(gclk));
	jdff dff_A_jth7tJDE4_2(.dout(w_dff_A_V1dGsCCM7_0),.din(w_dff_A_jth7tJDE4_2),.clk(gclk));
	jdff dff_A_V1dGsCCM7_0(.dout(w_dff_A_oqpsioch9_0),.din(w_dff_A_V1dGsCCM7_0),.clk(gclk));
	jdff dff_A_oqpsioch9_0(.dout(w_dff_A_FBvVIzWY2_0),.din(w_dff_A_oqpsioch9_0),.clk(gclk));
	jdff dff_A_FBvVIzWY2_0(.dout(w_dff_A_xbRA5X9p5_0),.din(w_dff_A_FBvVIzWY2_0),.clk(gclk));
	jdff dff_A_xbRA5X9p5_0(.dout(w_dff_A_Nm9K2iCn4_0),.din(w_dff_A_xbRA5X9p5_0),.clk(gclk));
	jdff dff_A_Nm9K2iCn4_0(.dout(w_dff_A_609eHOsQ7_0),.din(w_dff_A_Nm9K2iCn4_0),.clk(gclk));
	jdff dff_A_609eHOsQ7_0(.dout(w_dff_A_LmHUcl7l8_0),.din(w_dff_A_609eHOsQ7_0),.clk(gclk));
	jdff dff_A_LmHUcl7l8_0(.dout(w_dff_A_vR2hI2l76_0),.din(w_dff_A_LmHUcl7l8_0),.clk(gclk));
	jdff dff_A_vR2hI2l76_0(.dout(w_dff_A_SDchV6BP6_0),.din(w_dff_A_vR2hI2l76_0),.clk(gclk));
	jdff dff_A_SDchV6BP6_0(.dout(w_dff_A_4RXx2lW24_0),.din(w_dff_A_SDchV6BP6_0),.clk(gclk));
	jdff dff_A_4RXx2lW24_0(.dout(w_dff_A_XC6hkmqM3_0),.din(w_dff_A_4RXx2lW24_0),.clk(gclk));
	jdff dff_A_XC6hkmqM3_0(.dout(w_dff_A_DU5JkoUh6_0),.din(w_dff_A_XC6hkmqM3_0),.clk(gclk));
	jdff dff_A_DU5JkoUh6_0(.dout(w_dff_A_f7dD0e0w5_0),.din(w_dff_A_DU5JkoUh6_0),.clk(gclk));
	jdff dff_A_f7dD0e0w5_0(.dout(w_dff_A_kdfSSpBn7_0),.din(w_dff_A_f7dD0e0w5_0),.clk(gclk));
	jdff dff_A_kdfSSpBn7_0(.dout(w_dff_A_X07Dzd4B8_0),.din(w_dff_A_kdfSSpBn7_0),.clk(gclk));
	jdff dff_A_X07Dzd4B8_0(.dout(w_dff_A_TjyJTRN73_0),.din(w_dff_A_X07Dzd4B8_0),.clk(gclk));
	jdff dff_A_TjyJTRN73_0(.dout(w_dff_A_T9LIP4ij6_0),.din(w_dff_A_TjyJTRN73_0),.clk(gclk));
	jdff dff_A_T9LIP4ij6_0(.dout(w_dff_A_dCuIuUfN1_0),.din(w_dff_A_T9LIP4ij6_0),.clk(gclk));
	jdff dff_A_dCuIuUfN1_0(.dout(w_dff_A_2yIgaWsg8_0),.din(w_dff_A_dCuIuUfN1_0),.clk(gclk));
	jdff dff_A_2yIgaWsg8_0(.dout(w_dff_A_Ulvsk4vP0_0),.din(w_dff_A_2yIgaWsg8_0),.clk(gclk));
	jdff dff_A_Ulvsk4vP0_0(.dout(w_dff_A_iheEw9AN7_0),.din(w_dff_A_Ulvsk4vP0_0),.clk(gclk));
	jdff dff_A_iheEw9AN7_0(.dout(w_dff_A_63E4zvyf8_0),.din(w_dff_A_iheEw9AN7_0),.clk(gclk));
	jdff dff_A_63E4zvyf8_0(.dout(w_dff_A_vBRWUc9B3_0),.din(w_dff_A_63E4zvyf8_0),.clk(gclk));
	jdff dff_A_vBRWUc9B3_0(.dout(w_dff_A_XHOBbnYp9_0),.din(w_dff_A_vBRWUc9B3_0),.clk(gclk));
	jdff dff_A_XHOBbnYp9_0(.dout(w_dff_A_JQxkL62B2_0),.din(w_dff_A_XHOBbnYp9_0),.clk(gclk));
	jdff dff_A_JQxkL62B2_0(.dout(w_dff_A_lMcdKPRB3_0),.din(w_dff_A_JQxkL62B2_0),.clk(gclk));
	jdff dff_A_lMcdKPRB3_0(.dout(w_dff_A_slMcurW44_0),.din(w_dff_A_lMcdKPRB3_0),.clk(gclk));
	jdff dff_A_slMcurW44_0(.dout(f99),.din(w_dff_A_slMcurW44_0),.clk(gclk));
	jdff dff_A_vGnqaJJF9_2(.dout(w_dff_A_TUq5Ubjf5_0),.din(w_dff_A_vGnqaJJF9_2),.clk(gclk));
	jdff dff_A_TUq5Ubjf5_0(.dout(w_dff_A_EPglFiZF0_0),.din(w_dff_A_TUq5Ubjf5_0),.clk(gclk));
	jdff dff_A_EPglFiZF0_0(.dout(w_dff_A_27Pf443e7_0),.din(w_dff_A_EPglFiZF0_0),.clk(gclk));
	jdff dff_A_27Pf443e7_0(.dout(w_dff_A_CkokMeok2_0),.din(w_dff_A_27Pf443e7_0),.clk(gclk));
	jdff dff_A_CkokMeok2_0(.dout(w_dff_A_8zeaxkIn2_0),.din(w_dff_A_CkokMeok2_0),.clk(gclk));
	jdff dff_A_8zeaxkIn2_0(.dout(w_dff_A_u82QWup05_0),.din(w_dff_A_8zeaxkIn2_0),.clk(gclk));
	jdff dff_A_u82QWup05_0(.dout(w_dff_A_gYo2DAND4_0),.din(w_dff_A_u82QWup05_0),.clk(gclk));
	jdff dff_A_gYo2DAND4_0(.dout(w_dff_A_fW51Of138_0),.din(w_dff_A_gYo2DAND4_0),.clk(gclk));
	jdff dff_A_fW51Of138_0(.dout(w_dff_A_v4W7ykMc4_0),.din(w_dff_A_fW51Of138_0),.clk(gclk));
	jdff dff_A_v4W7ykMc4_0(.dout(w_dff_A_wZ7I0XZw5_0),.din(w_dff_A_v4W7ykMc4_0),.clk(gclk));
	jdff dff_A_wZ7I0XZw5_0(.dout(w_dff_A_slYO8GMn1_0),.din(w_dff_A_wZ7I0XZw5_0),.clk(gclk));
	jdff dff_A_slYO8GMn1_0(.dout(w_dff_A_Bw7GPftn7_0),.din(w_dff_A_slYO8GMn1_0),.clk(gclk));
	jdff dff_A_Bw7GPftn7_0(.dout(w_dff_A_UT8Tuj5l2_0),.din(w_dff_A_Bw7GPftn7_0),.clk(gclk));
	jdff dff_A_UT8Tuj5l2_0(.dout(w_dff_A_nGZowy1a8_0),.din(w_dff_A_UT8Tuj5l2_0),.clk(gclk));
	jdff dff_A_nGZowy1a8_0(.dout(w_dff_A_JlqjK21E7_0),.din(w_dff_A_nGZowy1a8_0),.clk(gclk));
	jdff dff_A_JlqjK21E7_0(.dout(w_dff_A_Tx7FWKCP1_0),.din(w_dff_A_JlqjK21E7_0),.clk(gclk));
	jdff dff_A_Tx7FWKCP1_0(.dout(w_dff_A_UZ2YTpHk2_0),.din(w_dff_A_Tx7FWKCP1_0),.clk(gclk));
	jdff dff_A_UZ2YTpHk2_0(.dout(w_dff_A_ZXyfIqhh9_0),.din(w_dff_A_UZ2YTpHk2_0),.clk(gclk));
	jdff dff_A_ZXyfIqhh9_0(.dout(w_dff_A_OKIpevN61_0),.din(w_dff_A_ZXyfIqhh9_0),.clk(gclk));
	jdff dff_A_OKIpevN61_0(.dout(w_dff_A_epiqUJjz6_0),.din(w_dff_A_OKIpevN61_0),.clk(gclk));
	jdff dff_A_epiqUJjz6_0(.dout(w_dff_A_ME0a4nPr3_0),.din(w_dff_A_epiqUJjz6_0),.clk(gclk));
	jdff dff_A_ME0a4nPr3_0(.dout(w_dff_A_zhnxk0Qq3_0),.din(w_dff_A_ME0a4nPr3_0),.clk(gclk));
	jdff dff_A_zhnxk0Qq3_0(.dout(w_dff_A_2cpCqytp7_0),.din(w_dff_A_zhnxk0Qq3_0),.clk(gclk));
	jdff dff_A_2cpCqytp7_0(.dout(w_dff_A_k487bRJE0_0),.din(w_dff_A_2cpCqytp7_0),.clk(gclk));
	jdff dff_A_k487bRJE0_0(.dout(w_dff_A_L5DA1Ew38_0),.din(w_dff_A_k487bRJE0_0),.clk(gclk));
	jdff dff_A_L5DA1Ew38_0(.dout(w_dff_A_ZN5Pv19v0_0),.din(w_dff_A_L5DA1Ew38_0),.clk(gclk));
	jdff dff_A_ZN5Pv19v0_0(.dout(f100),.din(w_dff_A_ZN5Pv19v0_0),.clk(gclk));
	jdff dff_A_Fj4n1Rkq2_2(.dout(w_dff_A_hXEtOOHJ7_0),.din(w_dff_A_Fj4n1Rkq2_2),.clk(gclk));
	jdff dff_A_hXEtOOHJ7_0(.dout(w_dff_A_zPYaZlJv0_0),.din(w_dff_A_hXEtOOHJ7_0),.clk(gclk));
	jdff dff_A_zPYaZlJv0_0(.dout(w_dff_A_lsstklFy5_0),.din(w_dff_A_zPYaZlJv0_0),.clk(gclk));
	jdff dff_A_lsstklFy5_0(.dout(w_dff_A_okMKNz337_0),.din(w_dff_A_lsstklFy5_0),.clk(gclk));
	jdff dff_A_okMKNz337_0(.dout(w_dff_A_1sX6YB4P5_0),.din(w_dff_A_okMKNz337_0),.clk(gclk));
	jdff dff_A_1sX6YB4P5_0(.dout(w_dff_A_VB2xGp2w5_0),.din(w_dff_A_1sX6YB4P5_0),.clk(gclk));
	jdff dff_A_VB2xGp2w5_0(.dout(w_dff_A_TB8mrGKu0_0),.din(w_dff_A_VB2xGp2w5_0),.clk(gclk));
	jdff dff_A_TB8mrGKu0_0(.dout(w_dff_A_6gMvx1hS4_0),.din(w_dff_A_TB8mrGKu0_0),.clk(gclk));
	jdff dff_A_6gMvx1hS4_0(.dout(w_dff_A_ntZFqKDd6_0),.din(w_dff_A_6gMvx1hS4_0),.clk(gclk));
	jdff dff_A_ntZFqKDd6_0(.dout(w_dff_A_7N4kp3X63_0),.din(w_dff_A_ntZFqKDd6_0),.clk(gclk));
	jdff dff_A_7N4kp3X63_0(.dout(w_dff_A_bqWsk6JH0_0),.din(w_dff_A_7N4kp3X63_0),.clk(gclk));
	jdff dff_A_bqWsk6JH0_0(.dout(w_dff_A_TYQY54Mp1_0),.din(w_dff_A_bqWsk6JH0_0),.clk(gclk));
	jdff dff_A_TYQY54Mp1_0(.dout(w_dff_A_BHPBXFJe8_0),.din(w_dff_A_TYQY54Mp1_0),.clk(gclk));
	jdff dff_A_BHPBXFJe8_0(.dout(w_dff_A_jQ0eDOjk2_0),.din(w_dff_A_BHPBXFJe8_0),.clk(gclk));
	jdff dff_A_jQ0eDOjk2_0(.dout(w_dff_A_IqT8IT6l2_0),.din(w_dff_A_jQ0eDOjk2_0),.clk(gclk));
	jdff dff_A_IqT8IT6l2_0(.dout(w_dff_A_cCgJvPcb8_0),.din(w_dff_A_IqT8IT6l2_0),.clk(gclk));
	jdff dff_A_cCgJvPcb8_0(.dout(w_dff_A_eovcZIHQ7_0),.din(w_dff_A_cCgJvPcb8_0),.clk(gclk));
	jdff dff_A_eovcZIHQ7_0(.dout(w_dff_A_zEDwgM0L5_0),.din(w_dff_A_eovcZIHQ7_0),.clk(gclk));
	jdff dff_A_zEDwgM0L5_0(.dout(w_dff_A_fsnrjpag8_0),.din(w_dff_A_zEDwgM0L5_0),.clk(gclk));
	jdff dff_A_fsnrjpag8_0(.dout(w_dff_A_ST5L3gf98_0),.din(w_dff_A_fsnrjpag8_0),.clk(gclk));
	jdff dff_A_ST5L3gf98_0(.dout(w_dff_A_opiUc1bh3_0),.din(w_dff_A_ST5L3gf98_0),.clk(gclk));
	jdff dff_A_opiUc1bh3_0(.dout(w_dff_A_xl2jBpz60_0),.din(w_dff_A_opiUc1bh3_0),.clk(gclk));
	jdff dff_A_xl2jBpz60_0(.dout(w_dff_A_EAyseYti3_0),.din(w_dff_A_xl2jBpz60_0),.clk(gclk));
	jdff dff_A_EAyseYti3_0(.dout(w_dff_A_k7kRvua23_0),.din(w_dff_A_EAyseYti3_0),.clk(gclk));
	jdff dff_A_k7kRvua23_0(.dout(w_dff_A_LEtvUaOA7_0),.din(w_dff_A_k7kRvua23_0),.clk(gclk));
	jdff dff_A_LEtvUaOA7_0(.dout(f101),.din(w_dff_A_LEtvUaOA7_0),.clk(gclk));
	jdff dff_A_P3vaBdYA9_2(.dout(w_dff_A_wgW0wQKP7_0),.din(w_dff_A_P3vaBdYA9_2),.clk(gclk));
	jdff dff_A_wgW0wQKP7_0(.dout(w_dff_A_TEShzEva1_0),.din(w_dff_A_wgW0wQKP7_0),.clk(gclk));
	jdff dff_A_TEShzEva1_0(.dout(w_dff_A_kWujKEim4_0),.din(w_dff_A_TEShzEva1_0),.clk(gclk));
	jdff dff_A_kWujKEim4_0(.dout(w_dff_A_VmhHHbww9_0),.din(w_dff_A_kWujKEim4_0),.clk(gclk));
	jdff dff_A_VmhHHbww9_0(.dout(w_dff_A_JCso0TM61_0),.din(w_dff_A_VmhHHbww9_0),.clk(gclk));
	jdff dff_A_JCso0TM61_0(.dout(w_dff_A_mlH8pfmY3_0),.din(w_dff_A_JCso0TM61_0),.clk(gclk));
	jdff dff_A_mlH8pfmY3_0(.dout(w_dff_A_y31upuPF3_0),.din(w_dff_A_mlH8pfmY3_0),.clk(gclk));
	jdff dff_A_y31upuPF3_0(.dout(w_dff_A_WQ5oT3ZY3_0),.din(w_dff_A_y31upuPF3_0),.clk(gclk));
	jdff dff_A_WQ5oT3ZY3_0(.dout(w_dff_A_Utd4LhlA5_0),.din(w_dff_A_WQ5oT3ZY3_0),.clk(gclk));
	jdff dff_A_Utd4LhlA5_0(.dout(w_dff_A_LUFoTsyR0_0),.din(w_dff_A_Utd4LhlA5_0),.clk(gclk));
	jdff dff_A_LUFoTsyR0_0(.dout(w_dff_A_7BlsdwCI3_0),.din(w_dff_A_LUFoTsyR0_0),.clk(gclk));
	jdff dff_A_7BlsdwCI3_0(.dout(w_dff_A_5JG3KtDt2_0),.din(w_dff_A_7BlsdwCI3_0),.clk(gclk));
	jdff dff_A_5JG3KtDt2_0(.dout(w_dff_A_RYwAcxiH3_0),.din(w_dff_A_5JG3KtDt2_0),.clk(gclk));
	jdff dff_A_RYwAcxiH3_0(.dout(w_dff_A_WpCQYC4I6_0),.din(w_dff_A_RYwAcxiH3_0),.clk(gclk));
	jdff dff_A_WpCQYC4I6_0(.dout(w_dff_A_fbgpJ23L3_0),.din(w_dff_A_WpCQYC4I6_0),.clk(gclk));
	jdff dff_A_fbgpJ23L3_0(.dout(w_dff_A_C0MY41l90_0),.din(w_dff_A_fbgpJ23L3_0),.clk(gclk));
	jdff dff_A_C0MY41l90_0(.dout(w_dff_A_dtC4Y41o0_0),.din(w_dff_A_C0MY41l90_0),.clk(gclk));
	jdff dff_A_dtC4Y41o0_0(.dout(w_dff_A_ztH5nZhI4_0),.din(w_dff_A_dtC4Y41o0_0),.clk(gclk));
	jdff dff_A_ztH5nZhI4_0(.dout(w_dff_A_XJ4vC2Ol1_0),.din(w_dff_A_ztH5nZhI4_0),.clk(gclk));
	jdff dff_A_XJ4vC2Ol1_0(.dout(w_dff_A_hTSzYaC67_0),.din(w_dff_A_XJ4vC2Ol1_0),.clk(gclk));
	jdff dff_A_hTSzYaC67_0(.dout(w_dff_A_NI4DIGyU8_0),.din(w_dff_A_hTSzYaC67_0),.clk(gclk));
	jdff dff_A_NI4DIGyU8_0(.dout(w_dff_A_7QVvKskS0_0),.din(w_dff_A_NI4DIGyU8_0),.clk(gclk));
	jdff dff_A_7QVvKskS0_0(.dout(w_dff_A_POMwUXZ06_0),.din(w_dff_A_7QVvKskS0_0),.clk(gclk));
	jdff dff_A_POMwUXZ06_0(.dout(w_dff_A_mGf3FJTz7_0),.din(w_dff_A_POMwUXZ06_0),.clk(gclk));
	jdff dff_A_mGf3FJTz7_0(.dout(f102),.din(w_dff_A_mGf3FJTz7_0),.clk(gclk));
	jdff dff_A_XMlybQoI8_2(.dout(w_dff_A_DnPGD6s15_0),.din(w_dff_A_XMlybQoI8_2),.clk(gclk));
	jdff dff_A_DnPGD6s15_0(.dout(w_dff_A_aLqdgAdc8_0),.din(w_dff_A_DnPGD6s15_0),.clk(gclk));
	jdff dff_A_aLqdgAdc8_0(.dout(w_dff_A_VsMcGbNA4_0),.din(w_dff_A_aLqdgAdc8_0),.clk(gclk));
	jdff dff_A_VsMcGbNA4_0(.dout(w_dff_A_RRDLnXg30_0),.din(w_dff_A_VsMcGbNA4_0),.clk(gclk));
	jdff dff_A_RRDLnXg30_0(.dout(w_dff_A_0RLeMwV01_0),.din(w_dff_A_RRDLnXg30_0),.clk(gclk));
	jdff dff_A_0RLeMwV01_0(.dout(w_dff_A_SplXach55_0),.din(w_dff_A_0RLeMwV01_0),.clk(gclk));
	jdff dff_A_SplXach55_0(.dout(w_dff_A_Rup4IS1v6_0),.din(w_dff_A_SplXach55_0),.clk(gclk));
	jdff dff_A_Rup4IS1v6_0(.dout(w_dff_A_DUpeHa601_0),.din(w_dff_A_Rup4IS1v6_0),.clk(gclk));
	jdff dff_A_DUpeHa601_0(.dout(w_dff_A_gGBdJpjh0_0),.din(w_dff_A_DUpeHa601_0),.clk(gclk));
	jdff dff_A_gGBdJpjh0_0(.dout(w_dff_A_Dq5ar8i42_0),.din(w_dff_A_gGBdJpjh0_0),.clk(gclk));
	jdff dff_A_Dq5ar8i42_0(.dout(w_dff_A_wlDihNJk4_0),.din(w_dff_A_Dq5ar8i42_0),.clk(gclk));
	jdff dff_A_wlDihNJk4_0(.dout(w_dff_A_qSm3hOd71_0),.din(w_dff_A_wlDihNJk4_0),.clk(gclk));
	jdff dff_A_qSm3hOd71_0(.dout(w_dff_A_nJg4aDGr2_0),.din(w_dff_A_qSm3hOd71_0),.clk(gclk));
	jdff dff_A_nJg4aDGr2_0(.dout(w_dff_A_TfuZ4JPa7_0),.din(w_dff_A_nJg4aDGr2_0),.clk(gclk));
	jdff dff_A_TfuZ4JPa7_0(.dout(w_dff_A_vxsUmO9G3_0),.din(w_dff_A_TfuZ4JPa7_0),.clk(gclk));
	jdff dff_A_vxsUmO9G3_0(.dout(w_dff_A_y60o0Nyw9_0),.din(w_dff_A_vxsUmO9G3_0),.clk(gclk));
	jdff dff_A_y60o0Nyw9_0(.dout(w_dff_A_keigOqtW6_0),.din(w_dff_A_y60o0Nyw9_0),.clk(gclk));
	jdff dff_A_keigOqtW6_0(.dout(w_dff_A_G2nbdawe5_0),.din(w_dff_A_keigOqtW6_0),.clk(gclk));
	jdff dff_A_G2nbdawe5_0(.dout(w_dff_A_y1NYJzuH5_0),.din(w_dff_A_G2nbdawe5_0),.clk(gclk));
	jdff dff_A_y1NYJzuH5_0(.dout(w_dff_A_N54wXrV99_0),.din(w_dff_A_y1NYJzuH5_0),.clk(gclk));
	jdff dff_A_N54wXrV99_0(.dout(w_dff_A_UFL3lFAj9_0),.din(w_dff_A_N54wXrV99_0),.clk(gclk));
	jdff dff_A_UFL3lFAj9_0(.dout(w_dff_A_MYRBxoZT7_0),.din(w_dff_A_UFL3lFAj9_0),.clk(gclk));
	jdff dff_A_MYRBxoZT7_0(.dout(w_dff_A_vcPCwn541_0),.din(w_dff_A_MYRBxoZT7_0),.clk(gclk));
	jdff dff_A_vcPCwn541_0(.dout(f103),.din(w_dff_A_vcPCwn541_0),.clk(gclk));
	jdff dff_A_5ieeOtHr7_2(.dout(w_dff_A_zoSumTK41_0),.din(w_dff_A_5ieeOtHr7_2),.clk(gclk));
	jdff dff_A_zoSumTK41_0(.dout(w_dff_A_djrT8tsr0_0),.din(w_dff_A_zoSumTK41_0),.clk(gclk));
	jdff dff_A_djrT8tsr0_0(.dout(w_dff_A_SW1g5nM00_0),.din(w_dff_A_djrT8tsr0_0),.clk(gclk));
	jdff dff_A_SW1g5nM00_0(.dout(w_dff_A_cMwlRTG65_0),.din(w_dff_A_SW1g5nM00_0),.clk(gclk));
	jdff dff_A_cMwlRTG65_0(.dout(w_dff_A_zzmi3HH02_0),.din(w_dff_A_cMwlRTG65_0),.clk(gclk));
	jdff dff_A_zzmi3HH02_0(.dout(w_dff_A_QMOoHHeL5_0),.din(w_dff_A_zzmi3HH02_0),.clk(gclk));
	jdff dff_A_QMOoHHeL5_0(.dout(w_dff_A_gLMsXJs80_0),.din(w_dff_A_QMOoHHeL5_0),.clk(gclk));
	jdff dff_A_gLMsXJs80_0(.dout(w_dff_A_d3b9AFFd2_0),.din(w_dff_A_gLMsXJs80_0),.clk(gclk));
	jdff dff_A_d3b9AFFd2_0(.dout(w_dff_A_MqDIMbQG9_0),.din(w_dff_A_d3b9AFFd2_0),.clk(gclk));
	jdff dff_A_MqDIMbQG9_0(.dout(w_dff_A_xLkATVKT3_0),.din(w_dff_A_MqDIMbQG9_0),.clk(gclk));
	jdff dff_A_xLkATVKT3_0(.dout(w_dff_A_iX2EXJGN3_0),.din(w_dff_A_xLkATVKT3_0),.clk(gclk));
	jdff dff_A_iX2EXJGN3_0(.dout(w_dff_A_4Hojidmt9_0),.din(w_dff_A_iX2EXJGN3_0),.clk(gclk));
	jdff dff_A_4Hojidmt9_0(.dout(w_dff_A_YiNWJ4kD9_0),.din(w_dff_A_4Hojidmt9_0),.clk(gclk));
	jdff dff_A_YiNWJ4kD9_0(.dout(w_dff_A_SxbIkGKd3_0),.din(w_dff_A_YiNWJ4kD9_0),.clk(gclk));
	jdff dff_A_SxbIkGKd3_0(.dout(w_dff_A_hFFa02gQ4_0),.din(w_dff_A_SxbIkGKd3_0),.clk(gclk));
	jdff dff_A_hFFa02gQ4_0(.dout(w_dff_A_4SZg7hkt0_0),.din(w_dff_A_hFFa02gQ4_0),.clk(gclk));
	jdff dff_A_4SZg7hkt0_0(.dout(w_dff_A_2YGmEzHA8_0),.din(w_dff_A_4SZg7hkt0_0),.clk(gclk));
	jdff dff_A_2YGmEzHA8_0(.dout(w_dff_A_fbLZO0UM7_0),.din(w_dff_A_2YGmEzHA8_0),.clk(gclk));
	jdff dff_A_fbLZO0UM7_0(.dout(w_dff_A_H8mMMVgf0_0),.din(w_dff_A_fbLZO0UM7_0),.clk(gclk));
	jdff dff_A_H8mMMVgf0_0(.dout(w_dff_A_pI0NoPbT6_0),.din(w_dff_A_H8mMMVgf0_0),.clk(gclk));
	jdff dff_A_pI0NoPbT6_0(.dout(w_dff_A_MRXsOHl51_0),.din(w_dff_A_pI0NoPbT6_0),.clk(gclk));
	jdff dff_A_MRXsOHl51_0(.dout(w_dff_A_dX5aVNW90_0),.din(w_dff_A_MRXsOHl51_0),.clk(gclk));
	jdff dff_A_dX5aVNW90_0(.dout(f104),.din(w_dff_A_dX5aVNW90_0),.clk(gclk));
	jdff dff_A_ZOM6W9LV4_2(.dout(w_dff_A_mIgwi5UL9_0),.din(w_dff_A_ZOM6W9LV4_2),.clk(gclk));
	jdff dff_A_mIgwi5UL9_0(.dout(w_dff_A_XFpw9E6u2_0),.din(w_dff_A_mIgwi5UL9_0),.clk(gclk));
	jdff dff_A_XFpw9E6u2_0(.dout(w_dff_A_NZF4uEZs0_0),.din(w_dff_A_XFpw9E6u2_0),.clk(gclk));
	jdff dff_A_NZF4uEZs0_0(.dout(w_dff_A_MYFDGeFq7_0),.din(w_dff_A_NZF4uEZs0_0),.clk(gclk));
	jdff dff_A_MYFDGeFq7_0(.dout(w_dff_A_0hvkPZNW7_0),.din(w_dff_A_MYFDGeFq7_0),.clk(gclk));
	jdff dff_A_0hvkPZNW7_0(.dout(w_dff_A_XyHIVfkr3_0),.din(w_dff_A_0hvkPZNW7_0),.clk(gclk));
	jdff dff_A_XyHIVfkr3_0(.dout(w_dff_A_cERMalAW1_0),.din(w_dff_A_XyHIVfkr3_0),.clk(gclk));
	jdff dff_A_cERMalAW1_0(.dout(w_dff_A_maQDEzpY8_0),.din(w_dff_A_cERMalAW1_0),.clk(gclk));
	jdff dff_A_maQDEzpY8_0(.dout(w_dff_A_CkOgGDVh6_0),.din(w_dff_A_maQDEzpY8_0),.clk(gclk));
	jdff dff_A_CkOgGDVh6_0(.dout(w_dff_A_hRrtdQzl4_0),.din(w_dff_A_CkOgGDVh6_0),.clk(gclk));
	jdff dff_A_hRrtdQzl4_0(.dout(w_dff_A_VhbgBBqp3_0),.din(w_dff_A_hRrtdQzl4_0),.clk(gclk));
	jdff dff_A_VhbgBBqp3_0(.dout(w_dff_A_kKmAAYk10_0),.din(w_dff_A_VhbgBBqp3_0),.clk(gclk));
	jdff dff_A_kKmAAYk10_0(.dout(w_dff_A_Rf5lOyIV9_0),.din(w_dff_A_kKmAAYk10_0),.clk(gclk));
	jdff dff_A_Rf5lOyIV9_0(.dout(w_dff_A_HeTMY7S33_0),.din(w_dff_A_Rf5lOyIV9_0),.clk(gclk));
	jdff dff_A_HeTMY7S33_0(.dout(w_dff_A_sMpvmZLb5_0),.din(w_dff_A_HeTMY7S33_0),.clk(gclk));
	jdff dff_A_sMpvmZLb5_0(.dout(w_dff_A_pBeQ16zq6_0),.din(w_dff_A_sMpvmZLb5_0),.clk(gclk));
	jdff dff_A_pBeQ16zq6_0(.dout(w_dff_A_k96B1frD7_0),.din(w_dff_A_pBeQ16zq6_0),.clk(gclk));
	jdff dff_A_k96B1frD7_0(.dout(w_dff_A_sKaCFLvi4_0),.din(w_dff_A_k96B1frD7_0),.clk(gclk));
	jdff dff_A_sKaCFLvi4_0(.dout(w_dff_A_JaihCoN39_0),.din(w_dff_A_sKaCFLvi4_0),.clk(gclk));
	jdff dff_A_JaihCoN39_0(.dout(w_dff_A_OERwHGfQ5_0),.din(w_dff_A_JaihCoN39_0),.clk(gclk));
	jdff dff_A_OERwHGfQ5_0(.dout(w_dff_A_6Yj68FtL3_0),.din(w_dff_A_OERwHGfQ5_0),.clk(gclk));
	jdff dff_A_6Yj68FtL3_0(.dout(f105),.din(w_dff_A_6Yj68FtL3_0),.clk(gclk));
	jdff dff_A_URhuMiJa9_2(.dout(w_dff_A_R5xOR7iw0_0),.din(w_dff_A_URhuMiJa9_2),.clk(gclk));
	jdff dff_A_R5xOR7iw0_0(.dout(w_dff_A_AcrXoWmU0_0),.din(w_dff_A_R5xOR7iw0_0),.clk(gclk));
	jdff dff_A_AcrXoWmU0_0(.dout(w_dff_A_WIV82wZ56_0),.din(w_dff_A_AcrXoWmU0_0),.clk(gclk));
	jdff dff_A_WIV82wZ56_0(.dout(w_dff_A_mql5OtEv4_0),.din(w_dff_A_WIV82wZ56_0),.clk(gclk));
	jdff dff_A_mql5OtEv4_0(.dout(w_dff_A_X14564wG4_0),.din(w_dff_A_mql5OtEv4_0),.clk(gclk));
	jdff dff_A_X14564wG4_0(.dout(w_dff_A_HRLznOIr3_0),.din(w_dff_A_X14564wG4_0),.clk(gclk));
	jdff dff_A_HRLznOIr3_0(.dout(w_dff_A_83FIooh79_0),.din(w_dff_A_HRLznOIr3_0),.clk(gclk));
	jdff dff_A_83FIooh79_0(.dout(w_dff_A_eYcdS94q2_0),.din(w_dff_A_83FIooh79_0),.clk(gclk));
	jdff dff_A_eYcdS94q2_0(.dout(w_dff_A_x0Qy0WX98_0),.din(w_dff_A_eYcdS94q2_0),.clk(gclk));
	jdff dff_A_x0Qy0WX98_0(.dout(w_dff_A_KyRbk5do0_0),.din(w_dff_A_x0Qy0WX98_0),.clk(gclk));
	jdff dff_A_KyRbk5do0_0(.dout(w_dff_A_gXpRIzGV1_0),.din(w_dff_A_KyRbk5do0_0),.clk(gclk));
	jdff dff_A_gXpRIzGV1_0(.dout(w_dff_A_uFwR1n136_0),.din(w_dff_A_gXpRIzGV1_0),.clk(gclk));
	jdff dff_A_uFwR1n136_0(.dout(w_dff_A_Au45byRy8_0),.din(w_dff_A_uFwR1n136_0),.clk(gclk));
	jdff dff_A_Au45byRy8_0(.dout(w_dff_A_J7dGG6DA3_0),.din(w_dff_A_Au45byRy8_0),.clk(gclk));
	jdff dff_A_J7dGG6DA3_0(.dout(w_dff_A_yzi3vWZX4_0),.din(w_dff_A_J7dGG6DA3_0),.clk(gclk));
	jdff dff_A_yzi3vWZX4_0(.dout(w_dff_A_HVvuYU7h3_0),.din(w_dff_A_yzi3vWZX4_0),.clk(gclk));
	jdff dff_A_HVvuYU7h3_0(.dout(w_dff_A_ZuuRcs2H9_0),.din(w_dff_A_HVvuYU7h3_0),.clk(gclk));
	jdff dff_A_ZuuRcs2H9_0(.dout(w_dff_A_HPNQdwgI4_0),.din(w_dff_A_ZuuRcs2H9_0),.clk(gclk));
	jdff dff_A_HPNQdwgI4_0(.dout(w_dff_A_1icJqdb29_0),.din(w_dff_A_HPNQdwgI4_0),.clk(gclk));
	jdff dff_A_1icJqdb29_0(.dout(w_dff_A_3Lo9b6G18_0),.din(w_dff_A_1icJqdb29_0),.clk(gclk));
	jdff dff_A_3Lo9b6G18_0(.dout(f106),.din(w_dff_A_3Lo9b6G18_0),.clk(gclk));
	jdff dff_A_cwkY2DxV9_2(.dout(w_dff_A_QvqEaHKG4_0),.din(w_dff_A_cwkY2DxV9_2),.clk(gclk));
	jdff dff_A_QvqEaHKG4_0(.dout(w_dff_A_EjyZ383l8_0),.din(w_dff_A_QvqEaHKG4_0),.clk(gclk));
	jdff dff_A_EjyZ383l8_0(.dout(w_dff_A_JVRc0Ru27_0),.din(w_dff_A_EjyZ383l8_0),.clk(gclk));
	jdff dff_A_JVRc0Ru27_0(.dout(w_dff_A_Wjpi3EFy3_0),.din(w_dff_A_JVRc0Ru27_0),.clk(gclk));
	jdff dff_A_Wjpi3EFy3_0(.dout(w_dff_A_svbN2EnZ7_0),.din(w_dff_A_Wjpi3EFy3_0),.clk(gclk));
	jdff dff_A_svbN2EnZ7_0(.dout(w_dff_A_uq6gKeGI7_0),.din(w_dff_A_svbN2EnZ7_0),.clk(gclk));
	jdff dff_A_uq6gKeGI7_0(.dout(w_dff_A_1NPtqsrc0_0),.din(w_dff_A_uq6gKeGI7_0),.clk(gclk));
	jdff dff_A_1NPtqsrc0_0(.dout(w_dff_A_Q0YMngAh6_0),.din(w_dff_A_1NPtqsrc0_0),.clk(gclk));
	jdff dff_A_Q0YMngAh6_0(.dout(w_dff_A_IeCXc6Qg3_0),.din(w_dff_A_Q0YMngAh6_0),.clk(gclk));
	jdff dff_A_IeCXc6Qg3_0(.dout(w_dff_A_64UkebS74_0),.din(w_dff_A_IeCXc6Qg3_0),.clk(gclk));
	jdff dff_A_64UkebS74_0(.dout(w_dff_A_d2IRJ8AP8_0),.din(w_dff_A_64UkebS74_0),.clk(gclk));
	jdff dff_A_d2IRJ8AP8_0(.dout(w_dff_A_nklNoIf45_0),.din(w_dff_A_d2IRJ8AP8_0),.clk(gclk));
	jdff dff_A_nklNoIf45_0(.dout(w_dff_A_DZ28DWka4_0),.din(w_dff_A_nklNoIf45_0),.clk(gclk));
	jdff dff_A_DZ28DWka4_0(.dout(w_dff_A_rdmNDJLK3_0),.din(w_dff_A_DZ28DWka4_0),.clk(gclk));
	jdff dff_A_rdmNDJLK3_0(.dout(w_dff_A_ySSQOess4_0),.din(w_dff_A_rdmNDJLK3_0),.clk(gclk));
	jdff dff_A_ySSQOess4_0(.dout(w_dff_A_7eqsieVT7_0),.din(w_dff_A_ySSQOess4_0),.clk(gclk));
	jdff dff_A_7eqsieVT7_0(.dout(w_dff_A_oGHixy531_0),.din(w_dff_A_7eqsieVT7_0),.clk(gclk));
	jdff dff_A_oGHixy531_0(.dout(w_dff_A_e0xhZWKO7_0),.din(w_dff_A_oGHixy531_0),.clk(gclk));
	jdff dff_A_e0xhZWKO7_0(.dout(w_dff_A_0TBOmsVl5_0),.din(w_dff_A_e0xhZWKO7_0),.clk(gclk));
	jdff dff_A_0TBOmsVl5_0(.dout(f107),.din(w_dff_A_0TBOmsVl5_0),.clk(gclk));
	jdff dff_A_aQI6d3Nn2_2(.dout(w_dff_A_AzNc77CQ7_0),.din(w_dff_A_aQI6d3Nn2_2),.clk(gclk));
	jdff dff_A_AzNc77CQ7_0(.dout(w_dff_A_LCM4Yejg9_0),.din(w_dff_A_AzNc77CQ7_0),.clk(gclk));
	jdff dff_A_LCM4Yejg9_0(.dout(w_dff_A_uIPLGUNv6_0),.din(w_dff_A_LCM4Yejg9_0),.clk(gclk));
	jdff dff_A_uIPLGUNv6_0(.dout(w_dff_A_YCe56c4y2_0),.din(w_dff_A_uIPLGUNv6_0),.clk(gclk));
	jdff dff_A_YCe56c4y2_0(.dout(w_dff_A_eLLA1vKa2_0),.din(w_dff_A_YCe56c4y2_0),.clk(gclk));
	jdff dff_A_eLLA1vKa2_0(.dout(w_dff_A_1uwtFH7b0_0),.din(w_dff_A_eLLA1vKa2_0),.clk(gclk));
	jdff dff_A_1uwtFH7b0_0(.dout(w_dff_A_zMgjeUZL0_0),.din(w_dff_A_1uwtFH7b0_0),.clk(gclk));
	jdff dff_A_zMgjeUZL0_0(.dout(w_dff_A_CMUE9ayB0_0),.din(w_dff_A_zMgjeUZL0_0),.clk(gclk));
	jdff dff_A_CMUE9ayB0_0(.dout(w_dff_A_ktuva36K9_0),.din(w_dff_A_CMUE9ayB0_0),.clk(gclk));
	jdff dff_A_ktuva36K9_0(.dout(w_dff_A_FyeagAyb5_0),.din(w_dff_A_ktuva36K9_0),.clk(gclk));
	jdff dff_A_FyeagAyb5_0(.dout(w_dff_A_9QuLYpSU7_0),.din(w_dff_A_FyeagAyb5_0),.clk(gclk));
	jdff dff_A_9QuLYpSU7_0(.dout(w_dff_A_I9774roP9_0),.din(w_dff_A_9QuLYpSU7_0),.clk(gclk));
	jdff dff_A_I9774roP9_0(.dout(w_dff_A_woYQbONg7_0),.din(w_dff_A_I9774roP9_0),.clk(gclk));
	jdff dff_A_woYQbONg7_0(.dout(w_dff_A_aW0JcCXM5_0),.din(w_dff_A_woYQbONg7_0),.clk(gclk));
	jdff dff_A_aW0JcCXM5_0(.dout(w_dff_A_7jZtU57U6_0),.din(w_dff_A_aW0JcCXM5_0),.clk(gclk));
	jdff dff_A_7jZtU57U6_0(.dout(w_dff_A_y0zwjRrI2_0),.din(w_dff_A_7jZtU57U6_0),.clk(gclk));
	jdff dff_A_y0zwjRrI2_0(.dout(w_dff_A_IDNxqPEX8_0),.din(w_dff_A_y0zwjRrI2_0),.clk(gclk));
	jdff dff_A_IDNxqPEX8_0(.dout(w_dff_A_QovH0nhy8_0),.din(w_dff_A_IDNxqPEX8_0),.clk(gclk));
	jdff dff_A_QovH0nhy8_0(.dout(f108),.din(w_dff_A_QovH0nhy8_0),.clk(gclk));
	jdff dff_A_6RAzsJrE3_2(.dout(w_dff_A_fcPJaCHr9_0),.din(w_dff_A_6RAzsJrE3_2),.clk(gclk));
	jdff dff_A_fcPJaCHr9_0(.dout(w_dff_A_Pt75JKha0_0),.din(w_dff_A_fcPJaCHr9_0),.clk(gclk));
	jdff dff_A_Pt75JKha0_0(.dout(w_dff_A_pDrdtPCf8_0),.din(w_dff_A_Pt75JKha0_0),.clk(gclk));
	jdff dff_A_pDrdtPCf8_0(.dout(w_dff_A_9sOSToaq3_0),.din(w_dff_A_pDrdtPCf8_0),.clk(gclk));
	jdff dff_A_9sOSToaq3_0(.dout(w_dff_A_tats9DAT7_0),.din(w_dff_A_9sOSToaq3_0),.clk(gclk));
	jdff dff_A_tats9DAT7_0(.dout(w_dff_A_xVMTakRC2_0),.din(w_dff_A_tats9DAT7_0),.clk(gclk));
	jdff dff_A_xVMTakRC2_0(.dout(w_dff_A_U5svZFhj4_0),.din(w_dff_A_xVMTakRC2_0),.clk(gclk));
	jdff dff_A_U5svZFhj4_0(.dout(w_dff_A_qYmj0XIQ6_0),.din(w_dff_A_U5svZFhj4_0),.clk(gclk));
	jdff dff_A_qYmj0XIQ6_0(.dout(w_dff_A_j4BASZgP3_0),.din(w_dff_A_qYmj0XIQ6_0),.clk(gclk));
	jdff dff_A_j4BASZgP3_0(.dout(w_dff_A_FtrYgpAU5_0),.din(w_dff_A_j4BASZgP3_0),.clk(gclk));
	jdff dff_A_FtrYgpAU5_0(.dout(w_dff_A_LssIE8tW7_0),.din(w_dff_A_FtrYgpAU5_0),.clk(gclk));
	jdff dff_A_LssIE8tW7_0(.dout(w_dff_A_D23S3ID22_0),.din(w_dff_A_LssIE8tW7_0),.clk(gclk));
	jdff dff_A_D23S3ID22_0(.dout(w_dff_A_6fgPjKce4_0),.din(w_dff_A_D23S3ID22_0),.clk(gclk));
	jdff dff_A_6fgPjKce4_0(.dout(w_dff_A_ZSQ4I4Ui4_0),.din(w_dff_A_6fgPjKce4_0),.clk(gclk));
	jdff dff_A_ZSQ4I4Ui4_0(.dout(w_dff_A_jY6jEer21_0),.din(w_dff_A_ZSQ4I4Ui4_0),.clk(gclk));
	jdff dff_A_jY6jEer21_0(.dout(w_dff_A_R2MXtO1e0_0),.din(w_dff_A_jY6jEer21_0),.clk(gclk));
	jdff dff_A_R2MXtO1e0_0(.dout(w_dff_A_apYP00tx6_0),.din(w_dff_A_R2MXtO1e0_0),.clk(gclk));
	jdff dff_A_apYP00tx6_0(.dout(f109),.din(w_dff_A_apYP00tx6_0),.clk(gclk));
	jdff dff_A_ukMTbJQ36_2(.dout(w_dff_A_wvEQ7hdg0_0),.din(w_dff_A_ukMTbJQ36_2),.clk(gclk));
	jdff dff_A_wvEQ7hdg0_0(.dout(w_dff_A_VU1EFMrT3_0),.din(w_dff_A_wvEQ7hdg0_0),.clk(gclk));
	jdff dff_A_VU1EFMrT3_0(.dout(w_dff_A_ZNqCzFb72_0),.din(w_dff_A_VU1EFMrT3_0),.clk(gclk));
	jdff dff_A_ZNqCzFb72_0(.dout(w_dff_A_83vQJNTY9_0),.din(w_dff_A_ZNqCzFb72_0),.clk(gclk));
	jdff dff_A_83vQJNTY9_0(.dout(w_dff_A_Mtznnj0x6_0),.din(w_dff_A_83vQJNTY9_0),.clk(gclk));
	jdff dff_A_Mtznnj0x6_0(.dout(w_dff_A_VFIf5r337_0),.din(w_dff_A_Mtznnj0x6_0),.clk(gclk));
	jdff dff_A_VFIf5r337_0(.dout(w_dff_A_yxJPLhbU3_0),.din(w_dff_A_VFIf5r337_0),.clk(gclk));
	jdff dff_A_yxJPLhbU3_0(.dout(w_dff_A_LKgLger15_0),.din(w_dff_A_yxJPLhbU3_0),.clk(gclk));
	jdff dff_A_LKgLger15_0(.dout(w_dff_A_poO4AJMA0_0),.din(w_dff_A_LKgLger15_0),.clk(gclk));
	jdff dff_A_poO4AJMA0_0(.dout(w_dff_A_8Tl9X62H9_0),.din(w_dff_A_poO4AJMA0_0),.clk(gclk));
	jdff dff_A_8Tl9X62H9_0(.dout(w_dff_A_4Abr1N4q3_0),.din(w_dff_A_8Tl9X62H9_0),.clk(gclk));
	jdff dff_A_4Abr1N4q3_0(.dout(w_dff_A_z9ixAAkq1_0),.din(w_dff_A_4Abr1N4q3_0),.clk(gclk));
	jdff dff_A_z9ixAAkq1_0(.dout(w_dff_A_ytJE0TKo5_0),.din(w_dff_A_z9ixAAkq1_0),.clk(gclk));
	jdff dff_A_ytJE0TKo5_0(.dout(w_dff_A_cmvhdiwe7_0),.din(w_dff_A_ytJE0TKo5_0),.clk(gclk));
	jdff dff_A_cmvhdiwe7_0(.dout(w_dff_A_bqz4TNf24_0),.din(w_dff_A_cmvhdiwe7_0),.clk(gclk));
	jdff dff_A_bqz4TNf24_0(.dout(w_dff_A_stwvBZNp3_0),.din(w_dff_A_bqz4TNf24_0),.clk(gclk));
	jdff dff_A_stwvBZNp3_0(.dout(f110),.din(w_dff_A_stwvBZNp3_0),.clk(gclk));
	jdff dff_A_kWw534XR3_2(.dout(w_dff_A_BidquCIy1_0),.din(w_dff_A_kWw534XR3_2),.clk(gclk));
	jdff dff_A_BidquCIy1_0(.dout(w_dff_A_VarZBo5k7_0),.din(w_dff_A_BidquCIy1_0),.clk(gclk));
	jdff dff_A_VarZBo5k7_0(.dout(w_dff_A_bKn9TE068_0),.din(w_dff_A_VarZBo5k7_0),.clk(gclk));
	jdff dff_A_bKn9TE068_0(.dout(w_dff_A_awMKTcC25_0),.din(w_dff_A_bKn9TE068_0),.clk(gclk));
	jdff dff_A_awMKTcC25_0(.dout(w_dff_A_dTG30o3B6_0),.din(w_dff_A_awMKTcC25_0),.clk(gclk));
	jdff dff_A_dTG30o3B6_0(.dout(w_dff_A_Ly0DCpf35_0),.din(w_dff_A_dTG30o3B6_0),.clk(gclk));
	jdff dff_A_Ly0DCpf35_0(.dout(w_dff_A_TcdsbM6c6_0),.din(w_dff_A_Ly0DCpf35_0),.clk(gclk));
	jdff dff_A_TcdsbM6c6_0(.dout(w_dff_A_lPHYUwfF7_0),.din(w_dff_A_TcdsbM6c6_0),.clk(gclk));
	jdff dff_A_lPHYUwfF7_0(.dout(w_dff_A_1C4UwDMw2_0),.din(w_dff_A_lPHYUwfF7_0),.clk(gclk));
	jdff dff_A_1C4UwDMw2_0(.dout(w_dff_A_wA3cx3SH3_0),.din(w_dff_A_1C4UwDMw2_0),.clk(gclk));
	jdff dff_A_wA3cx3SH3_0(.dout(w_dff_A_VYIjAtFW9_0),.din(w_dff_A_wA3cx3SH3_0),.clk(gclk));
	jdff dff_A_VYIjAtFW9_0(.dout(w_dff_A_7amHe4Bo5_0),.din(w_dff_A_VYIjAtFW9_0),.clk(gclk));
	jdff dff_A_7amHe4Bo5_0(.dout(w_dff_A_M6xb7lpj5_0),.din(w_dff_A_7amHe4Bo5_0),.clk(gclk));
	jdff dff_A_M6xb7lpj5_0(.dout(w_dff_A_tSKYmCYO7_0),.din(w_dff_A_M6xb7lpj5_0),.clk(gclk));
	jdff dff_A_tSKYmCYO7_0(.dout(w_dff_A_bHjWloGN6_0),.din(w_dff_A_tSKYmCYO7_0),.clk(gclk));
	jdff dff_A_bHjWloGN6_0(.dout(f111),.din(w_dff_A_bHjWloGN6_0),.clk(gclk));
	jdff dff_A_bne51yCD0_2(.dout(w_dff_A_WK6EJDtf0_0),.din(w_dff_A_bne51yCD0_2),.clk(gclk));
	jdff dff_A_WK6EJDtf0_0(.dout(w_dff_A_ClhUFvES4_0),.din(w_dff_A_WK6EJDtf0_0),.clk(gclk));
	jdff dff_A_ClhUFvES4_0(.dout(w_dff_A_zqNRi1lD4_0),.din(w_dff_A_ClhUFvES4_0),.clk(gclk));
	jdff dff_A_zqNRi1lD4_0(.dout(w_dff_A_FfOHGaCs6_0),.din(w_dff_A_zqNRi1lD4_0),.clk(gclk));
	jdff dff_A_FfOHGaCs6_0(.dout(w_dff_A_qvxSnGmK1_0),.din(w_dff_A_FfOHGaCs6_0),.clk(gclk));
	jdff dff_A_qvxSnGmK1_0(.dout(w_dff_A_BtXzz1kR5_0),.din(w_dff_A_qvxSnGmK1_0),.clk(gclk));
	jdff dff_A_BtXzz1kR5_0(.dout(w_dff_A_QIUA7GFY1_0),.din(w_dff_A_BtXzz1kR5_0),.clk(gclk));
	jdff dff_A_QIUA7GFY1_0(.dout(w_dff_A_jzqemet56_0),.din(w_dff_A_QIUA7GFY1_0),.clk(gclk));
	jdff dff_A_jzqemet56_0(.dout(w_dff_A_IBAGth7O9_0),.din(w_dff_A_jzqemet56_0),.clk(gclk));
	jdff dff_A_IBAGth7O9_0(.dout(w_dff_A_B095ri797_0),.din(w_dff_A_IBAGth7O9_0),.clk(gclk));
	jdff dff_A_B095ri797_0(.dout(w_dff_A_n2L41IjT2_0),.din(w_dff_A_B095ri797_0),.clk(gclk));
	jdff dff_A_n2L41IjT2_0(.dout(w_dff_A_XagthY0s2_0),.din(w_dff_A_n2L41IjT2_0),.clk(gclk));
	jdff dff_A_XagthY0s2_0(.dout(w_dff_A_Am07XMav3_0),.din(w_dff_A_XagthY0s2_0),.clk(gclk));
	jdff dff_A_Am07XMav3_0(.dout(w_dff_A_co00XfWT4_0),.din(w_dff_A_Am07XMav3_0),.clk(gclk));
	jdff dff_A_co00XfWT4_0(.dout(f112),.din(w_dff_A_co00XfWT4_0),.clk(gclk));
	jdff dff_A_3U7JlSNO5_2(.dout(w_dff_A_pnLvFod86_0),.din(w_dff_A_3U7JlSNO5_2),.clk(gclk));
	jdff dff_A_pnLvFod86_0(.dout(w_dff_A_aY6E5eNv5_0),.din(w_dff_A_pnLvFod86_0),.clk(gclk));
	jdff dff_A_aY6E5eNv5_0(.dout(w_dff_A_Y9gpwtXe4_0),.din(w_dff_A_aY6E5eNv5_0),.clk(gclk));
	jdff dff_A_Y9gpwtXe4_0(.dout(w_dff_A_azWlgLyn6_0),.din(w_dff_A_Y9gpwtXe4_0),.clk(gclk));
	jdff dff_A_azWlgLyn6_0(.dout(w_dff_A_Usu1l2Kb3_0),.din(w_dff_A_azWlgLyn6_0),.clk(gclk));
	jdff dff_A_Usu1l2Kb3_0(.dout(w_dff_A_WtFxGp7T6_0),.din(w_dff_A_Usu1l2Kb3_0),.clk(gclk));
	jdff dff_A_WtFxGp7T6_0(.dout(w_dff_A_AKHwbQAN1_0),.din(w_dff_A_WtFxGp7T6_0),.clk(gclk));
	jdff dff_A_AKHwbQAN1_0(.dout(w_dff_A_MfGW3Onq8_0),.din(w_dff_A_AKHwbQAN1_0),.clk(gclk));
	jdff dff_A_MfGW3Onq8_0(.dout(w_dff_A_C1MbJwYK1_0),.din(w_dff_A_MfGW3Onq8_0),.clk(gclk));
	jdff dff_A_C1MbJwYK1_0(.dout(w_dff_A_mBejUqLh8_0),.din(w_dff_A_C1MbJwYK1_0),.clk(gclk));
	jdff dff_A_mBejUqLh8_0(.dout(w_dff_A_7LEqFVeF4_0),.din(w_dff_A_mBejUqLh8_0),.clk(gclk));
	jdff dff_A_7LEqFVeF4_0(.dout(w_dff_A_deTQa9lE0_0),.din(w_dff_A_7LEqFVeF4_0),.clk(gclk));
	jdff dff_A_deTQa9lE0_0(.dout(w_dff_A_fKhiDbuw8_0),.din(w_dff_A_deTQa9lE0_0),.clk(gclk));
	jdff dff_A_fKhiDbuw8_0(.dout(f113),.din(w_dff_A_fKhiDbuw8_0),.clk(gclk));
	jdff dff_A_3VmB04UB2_2(.dout(w_dff_A_HaTQCZom3_0),.din(w_dff_A_3VmB04UB2_2),.clk(gclk));
	jdff dff_A_HaTQCZom3_0(.dout(w_dff_A_qzCNFlmB7_0),.din(w_dff_A_HaTQCZom3_0),.clk(gclk));
	jdff dff_A_qzCNFlmB7_0(.dout(w_dff_A_dcPacLFt4_0),.din(w_dff_A_qzCNFlmB7_0),.clk(gclk));
	jdff dff_A_dcPacLFt4_0(.dout(w_dff_A_HaXPQeVw0_0),.din(w_dff_A_dcPacLFt4_0),.clk(gclk));
	jdff dff_A_HaXPQeVw0_0(.dout(w_dff_A_QHBz4jk01_0),.din(w_dff_A_HaXPQeVw0_0),.clk(gclk));
	jdff dff_A_QHBz4jk01_0(.dout(w_dff_A_rR5VlmdJ0_0),.din(w_dff_A_QHBz4jk01_0),.clk(gclk));
	jdff dff_A_rR5VlmdJ0_0(.dout(w_dff_A_rkgx6CZI6_0),.din(w_dff_A_rR5VlmdJ0_0),.clk(gclk));
	jdff dff_A_rkgx6CZI6_0(.dout(w_dff_A_ZOBgwSoD9_0),.din(w_dff_A_rkgx6CZI6_0),.clk(gclk));
	jdff dff_A_ZOBgwSoD9_0(.dout(w_dff_A_qpir5nay3_0),.din(w_dff_A_ZOBgwSoD9_0),.clk(gclk));
	jdff dff_A_qpir5nay3_0(.dout(w_dff_A_o1t3YtAy4_0),.din(w_dff_A_qpir5nay3_0),.clk(gclk));
	jdff dff_A_o1t3YtAy4_0(.dout(w_dff_A_ejOVAiHG2_0),.din(w_dff_A_o1t3YtAy4_0),.clk(gclk));
	jdff dff_A_ejOVAiHG2_0(.dout(w_dff_A_7RRxYpKw9_0),.din(w_dff_A_ejOVAiHG2_0),.clk(gclk));
	jdff dff_A_7RRxYpKw9_0(.dout(f114),.din(w_dff_A_7RRxYpKw9_0),.clk(gclk));
	jdff dff_A_3bA8xD5P2_2(.dout(w_dff_A_vSSzQQdW7_0),.din(w_dff_A_3bA8xD5P2_2),.clk(gclk));
	jdff dff_A_vSSzQQdW7_0(.dout(w_dff_A_M2OmrYFS7_0),.din(w_dff_A_vSSzQQdW7_0),.clk(gclk));
	jdff dff_A_M2OmrYFS7_0(.dout(w_dff_A_cZL1uRaJ3_0),.din(w_dff_A_M2OmrYFS7_0),.clk(gclk));
	jdff dff_A_cZL1uRaJ3_0(.dout(w_dff_A_9yJbI2Ln9_0),.din(w_dff_A_cZL1uRaJ3_0),.clk(gclk));
	jdff dff_A_9yJbI2Ln9_0(.dout(w_dff_A_eSducORv0_0),.din(w_dff_A_9yJbI2Ln9_0),.clk(gclk));
	jdff dff_A_eSducORv0_0(.dout(w_dff_A_Pv6XwFBY6_0),.din(w_dff_A_eSducORv0_0),.clk(gclk));
	jdff dff_A_Pv6XwFBY6_0(.dout(w_dff_A_CLQlnbdo5_0),.din(w_dff_A_Pv6XwFBY6_0),.clk(gclk));
	jdff dff_A_CLQlnbdo5_0(.dout(w_dff_A_1oBmfopY1_0),.din(w_dff_A_CLQlnbdo5_0),.clk(gclk));
	jdff dff_A_1oBmfopY1_0(.dout(w_dff_A_FbUW3vO70_0),.din(w_dff_A_1oBmfopY1_0),.clk(gclk));
	jdff dff_A_FbUW3vO70_0(.dout(w_dff_A_p6zFibIm6_0),.din(w_dff_A_FbUW3vO70_0),.clk(gclk));
	jdff dff_A_p6zFibIm6_0(.dout(w_dff_A_8uaIeREO3_0),.din(w_dff_A_p6zFibIm6_0),.clk(gclk));
	jdff dff_A_8uaIeREO3_0(.dout(f115),.din(w_dff_A_8uaIeREO3_0),.clk(gclk));
	jdff dff_A_fKN0jFwO9_2(.dout(w_dff_A_7XAfmi9u6_0),.din(w_dff_A_fKN0jFwO9_2),.clk(gclk));
	jdff dff_A_7XAfmi9u6_0(.dout(w_dff_A_OlFkYmOn2_0),.din(w_dff_A_7XAfmi9u6_0),.clk(gclk));
	jdff dff_A_OlFkYmOn2_0(.dout(w_dff_A_KCwq0QBL8_0),.din(w_dff_A_OlFkYmOn2_0),.clk(gclk));
	jdff dff_A_KCwq0QBL8_0(.dout(w_dff_A_Iz7WlUZf0_0),.din(w_dff_A_KCwq0QBL8_0),.clk(gclk));
	jdff dff_A_Iz7WlUZf0_0(.dout(w_dff_A_WCk5HKwe4_0),.din(w_dff_A_Iz7WlUZf0_0),.clk(gclk));
	jdff dff_A_WCk5HKwe4_0(.dout(w_dff_A_Xv5Trcx60_0),.din(w_dff_A_WCk5HKwe4_0),.clk(gclk));
	jdff dff_A_Xv5Trcx60_0(.dout(w_dff_A_SBEmuX9o8_0),.din(w_dff_A_Xv5Trcx60_0),.clk(gclk));
	jdff dff_A_SBEmuX9o8_0(.dout(w_dff_A_8dYujpQX8_0),.din(w_dff_A_SBEmuX9o8_0),.clk(gclk));
	jdff dff_A_8dYujpQX8_0(.dout(w_dff_A_4mHypyvg4_0),.din(w_dff_A_8dYujpQX8_0),.clk(gclk));
	jdff dff_A_4mHypyvg4_0(.dout(w_dff_A_LBRWsrIM0_0),.din(w_dff_A_4mHypyvg4_0),.clk(gclk));
	jdff dff_A_LBRWsrIM0_0(.dout(f116),.din(w_dff_A_LBRWsrIM0_0),.clk(gclk));
	jdff dff_A_llLQJvtS3_2(.dout(w_dff_A_xrBJtCSZ0_0),.din(w_dff_A_llLQJvtS3_2),.clk(gclk));
	jdff dff_A_xrBJtCSZ0_0(.dout(w_dff_A_UK5NQipZ2_0),.din(w_dff_A_xrBJtCSZ0_0),.clk(gclk));
	jdff dff_A_UK5NQipZ2_0(.dout(w_dff_A_7JQOCkeH0_0),.din(w_dff_A_UK5NQipZ2_0),.clk(gclk));
	jdff dff_A_7JQOCkeH0_0(.dout(w_dff_A_okE5sMLk3_0),.din(w_dff_A_7JQOCkeH0_0),.clk(gclk));
	jdff dff_A_okE5sMLk3_0(.dout(w_dff_A_mYpIoqg69_0),.din(w_dff_A_okE5sMLk3_0),.clk(gclk));
	jdff dff_A_mYpIoqg69_0(.dout(w_dff_A_tCCFH3Xv7_0),.din(w_dff_A_mYpIoqg69_0),.clk(gclk));
	jdff dff_A_tCCFH3Xv7_0(.dout(w_dff_A_jPfqylYA2_0),.din(w_dff_A_tCCFH3Xv7_0),.clk(gclk));
	jdff dff_A_jPfqylYA2_0(.dout(w_dff_A_zBR8Aika4_0),.din(w_dff_A_jPfqylYA2_0),.clk(gclk));
	jdff dff_A_zBR8Aika4_0(.dout(w_dff_A_EcfhzWiX4_0),.din(w_dff_A_zBR8Aika4_0),.clk(gclk));
	jdff dff_A_EcfhzWiX4_0(.dout(f117),.din(w_dff_A_EcfhzWiX4_0),.clk(gclk));
	jdff dff_A_9UxeUz0e4_2(.dout(w_dff_A_ZTGYclPq4_0),.din(w_dff_A_9UxeUz0e4_2),.clk(gclk));
	jdff dff_A_ZTGYclPq4_0(.dout(w_dff_A_U7yMt1zL1_0),.din(w_dff_A_ZTGYclPq4_0),.clk(gclk));
	jdff dff_A_U7yMt1zL1_0(.dout(w_dff_A_7PxYVrBw0_0),.din(w_dff_A_U7yMt1zL1_0),.clk(gclk));
	jdff dff_A_7PxYVrBw0_0(.dout(w_dff_A_Ymx8UBmT3_0),.din(w_dff_A_7PxYVrBw0_0),.clk(gclk));
	jdff dff_A_Ymx8UBmT3_0(.dout(w_dff_A_yXYCHHPO8_0),.din(w_dff_A_Ymx8UBmT3_0),.clk(gclk));
	jdff dff_A_yXYCHHPO8_0(.dout(w_dff_A_JaAJ4YBp6_0),.din(w_dff_A_yXYCHHPO8_0),.clk(gclk));
	jdff dff_A_JaAJ4YBp6_0(.dout(w_dff_A_gL7u1HKB1_0),.din(w_dff_A_JaAJ4YBp6_0),.clk(gclk));
	jdff dff_A_gL7u1HKB1_0(.dout(w_dff_A_SaestAav7_0),.din(w_dff_A_gL7u1HKB1_0),.clk(gclk));
	jdff dff_A_SaestAav7_0(.dout(f118),.din(w_dff_A_SaestAav7_0),.clk(gclk));
	jdff dff_A_VEKg84Oy2_2(.dout(w_dff_A_tY6J68k74_0),.din(w_dff_A_VEKg84Oy2_2),.clk(gclk));
	jdff dff_A_tY6J68k74_0(.dout(w_dff_A_AasODOBE5_0),.din(w_dff_A_tY6J68k74_0),.clk(gclk));
	jdff dff_A_AasODOBE5_0(.dout(w_dff_A_7jrMCY5F3_0),.din(w_dff_A_AasODOBE5_0),.clk(gclk));
	jdff dff_A_7jrMCY5F3_0(.dout(w_dff_A_B81ZmGIY8_0),.din(w_dff_A_7jrMCY5F3_0),.clk(gclk));
	jdff dff_A_B81ZmGIY8_0(.dout(w_dff_A_lVdqU8uU9_0),.din(w_dff_A_B81ZmGIY8_0),.clk(gclk));
	jdff dff_A_lVdqU8uU9_0(.dout(w_dff_A_r4Mbs7zM4_0),.din(w_dff_A_lVdqU8uU9_0),.clk(gclk));
	jdff dff_A_r4Mbs7zM4_0(.dout(w_dff_A_16l6xVEV2_0),.din(w_dff_A_r4Mbs7zM4_0),.clk(gclk));
	jdff dff_A_16l6xVEV2_0(.dout(f119),.din(w_dff_A_16l6xVEV2_0),.clk(gclk));
	jdff dff_A_qLw4TMU81_2(.dout(w_dff_A_gQUcPB1M3_0),.din(w_dff_A_qLw4TMU81_2),.clk(gclk));
	jdff dff_A_gQUcPB1M3_0(.dout(w_dff_A_gXUcJs2c8_0),.din(w_dff_A_gQUcPB1M3_0),.clk(gclk));
	jdff dff_A_gXUcJs2c8_0(.dout(w_dff_A_wFBaKcoN0_0),.din(w_dff_A_gXUcJs2c8_0),.clk(gclk));
	jdff dff_A_wFBaKcoN0_0(.dout(w_dff_A_7ieWQnUJ4_0),.din(w_dff_A_wFBaKcoN0_0),.clk(gclk));
	jdff dff_A_7ieWQnUJ4_0(.dout(w_dff_A_YydnO40Y0_0),.din(w_dff_A_7ieWQnUJ4_0),.clk(gclk));
	jdff dff_A_YydnO40Y0_0(.dout(w_dff_A_l8FPsNhz8_0),.din(w_dff_A_YydnO40Y0_0),.clk(gclk));
	jdff dff_A_l8FPsNhz8_0(.dout(f120),.din(w_dff_A_l8FPsNhz8_0),.clk(gclk));
	jdff dff_A_72ECXwuX6_2(.dout(w_dff_A_6fdH6ibw7_0),.din(w_dff_A_72ECXwuX6_2),.clk(gclk));
	jdff dff_A_6fdH6ibw7_0(.dout(w_dff_A_V9DHNrXJ1_0),.din(w_dff_A_6fdH6ibw7_0),.clk(gclk));
	jdff dff_A_V9DHNrXJ1_0(.dout(w_dff_A_YAN9LuKi3_0),.din(w_dff_A_V9DHNrXJ1_0),.clk(gclk));
	jdff dff_A_YAN9LuKi3_0(.dout(w_dff_A_DIG7appW3_0),.din(w_dff_A_YAN9LuKi3_0),.clk(gclk));
	jdff dff_A_DIG7appW3_0(.dout(w_dff_A_l7fEUm0g5_0),.din(w_dff_A_DIG7appW3_0),.clk(gclk));
	jdff dff_A_l7fEUm0g5_0(.dout(f121),.din(w_dff_A_l7fEUm0g5_0),.clk(gclk));
	jdff dff_A_pUdZQfwk6_2(.dout(w_dff_A_SYV3Wbhr8_0),.din(w_dff_A_pUdZQfwk6_2),.clk(gclk));
	jdff dff_A_SYV3Wbhr8_0(.dout(w_dff_A_c3di3RzO0_0),.din(w_dff_A_SYV3Wbhr8_0),.clk(gclk));
	jdff dff_A_c3di3RzO0_0(.dout(w_dff_A_HlzORNQm3_0),.din(w_dff_A_c3di3RzO0_0),.clk(gclk));
	jdff dff_A_HlzORNQm3_0(.dout(w_dff_A_rPEjnIGK4_0),.din(w_dff_A_HlzORNQm3_0),.clk(gclk));
	jdff dff_A_rPEjnIGK4_0(.dout(f122),.din(w_dff_A_rPEjnIGK4_0),.clk(gclk));
	jdff dff_A_njEGwhT63_2(.dout(w_dff_A_nDWIoLhN5_0),.din(w_dff_A_njEGwhT63_2),.clk(gclk));
	jdff dff_A_nDWIoLhN5_0(.dout(w_dff_A_YOPuAJXX3_0),.din(w_dff_A_nDWIoLhN5_0),.clk(gclk));
	jdff dff_A_YOPuAJXX3_0(.dout(w_dff_A_YgokwFm35_0),.din(w_dff_A_YOPuAJXX3_0),.clk(gclk));
	jdff dff_A_YgokwFm35_0(.dout(f123),.din(w_dff_A_YgokwFm35_0),.clk(gclk));
	jdff dff_A_qPETohS16_2(.dout(w_dff_A_YWhCSTZH9_0),.din(w_dff_A_qPETohS16_2),.clk(gclk));
	jdff dff_A_YWhCSTZH9_0(.dout(w_dff_A_Xe9XK3yk0_0),.din(w_dff_A_YWhCSTZH9_0),.clk(gclk));
	jdff dff_A_Xe9XK3yk0_0(.dout(f124),.din(w_dff_A_Xe9XK3yk0_0),.clk(gclk));
	jdff dff_A_Dk9V03BL7_2(.dout(w_dff_A_QYfAqV0p5_0),.din(w_dff_A_Dk9V03BL7_2),.clk(gclk));
	jdff dff_A_QYfAqV0p5_0(.dout(f125),.din(w_dff_A_QYfAqV0p5_0),.clk(gclk));
	jdff dff_A_e8TKNRw88_2(.dout(f126),.din(w_dff_A_e8TKNRw88_2),.clk(gclk));
endmodule

