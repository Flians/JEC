/*

c1908:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 969
	jor: 87
	jand: 120

Summary:
	jxor: 78
	jspl: 105
	jspl3: 86
	jnot: 30
	jdff: 969
	jor: 87
	jand: 120
*/

module c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n173;
	wire n174;
	wire n175;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n201;
	wire n203;
	wire n204;
	wire n206;
	wire n207;
	wire n208;
	wire n210;
	wire n211;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n220;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n270;
	wire n271;
	wire n272;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n348;
	wire n349;
	wire n350;
	wire n352;
	wire n353;
	wire n354;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n369;
	wire n370;
	wire n371;
	wire[2:0] w_G101_0;
	wire[2:0] w_G104_0;
	wire[2:0] w_G107_0;
	wire[2:0] w_G110_0;
	wire[2:0] w_G113_0;
	wire[2:0] w_G116_0;
	wire[2:0] w_G119_0;
	wire[2:0] w_G122_0;
	wire[1:0] w_G122_1;
	wire[2:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[2:0] w_G131_0;
	wire[2:0] w_G134_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G140_0;
	wire[2:0] w_G143_0;
	wire[2:0] w_G146_0;
	wire[2:0] w_G210_0;
	wire[1:0] w_G214_0;
	wire[2:0] w_G217_0;
	wire[1:0] w_G221_0;
	wire[1:0] w_G224_0;
	wire[1:0] w_G227_0;
	wire[2:0] w_G234_0;
	wire[1:0] w_G234_1;
	wire[2:0] w_G237_0;
	wire[2:0] w_G469_0;
	wire[2:0] w_G472_0;
	wire[2:0] w_G475_0;
	wire[2:0] w_G478_0;
	wire[1:0] w_G898_0;
	wire[1:0] w_G900_0;
	wire[2:0] w_G902_0;
	wire[2:0] w_G902_1;
	wire[2:0] w_G902_2;
	wire[2:0] w_G902_3;
	wire[2:0] w_G952_0;
	wire[2:0] w_G953_0;
	wire[2:0] w_G953_1;
	wire[1:0] w_G953_2;
	wire[2:0] w_n58_0;
	wire[2:0] w_n58_1;
	wire[2:0] w_n58_2;
	wire[1:0] w_n63_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n71_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n74_0;
	wire[2:0] w_n76_0;
	wire[2:0] w_n76_1;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[2:0] w_n81_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[2:0] w_n92_0;
	wire[1:0] w_n92_1;
	wire[2:0] w_n93_0;
	wire[1:0] w_n93_1;
	wire[1:0] w_n94_0;
	wire[2:0] w_n95_0;
	wire[1:0] w_n95_1;
	wire[2:0] w_n96_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n102_0;
	wire[2:0] w_n103_0;
	wire[2:0] w_n103_1;
	wire[2:0] w_n103_2;
	wire[2:0] w_n103_3;
	wire[1:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n109_0;
	wire[1:0] w_n110_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n112_0;
	wire[1:0] w_n112_1;
	wire[2:0] w_n113_0;
	wire[1:0] w_n118_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[2:0] w_n122_0;
	wire[1:0] w_n122_1;
	wire[1:0] w_n124_0;
	wire[1:0] w_n126_0;
	wire[1:0] w_n127_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n130_1;
	wire[2:0] w_n131_0;
	wire[2:0] w_n131_1;
	wire[1:0] w_n139_0;
	wire[1:0] w_n140_0;
	wire[2:0] w_n141_0;
	wire[1:0] w_n141_1;
	wire[2:0] w_n151_0;
	wire[1:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[1:0] w_n153_1;
	wire[2:0] w_n154_0;
	wire[1:0] w_n154_1;
	wire[1:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n157_0;
	wire[2:0] w_n160_0;
	wire[2:0] w_n160_1;
	wire[2:0] w_n161_0;
	wire[1:0] w_n161_1;
	wire[1:0] w_n162_0;
	wire[2:0] w_n163_0;
	wire[1:0] w_n163_1;
	wire[1:0] w_n164_0;
	wire[2:0] w_n165_0;
	wire[1:0] w_n166_0;
	wire[2:0] w_n168_0;
	wire[1:0] w_n168_1;
	wire[1:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n171_0;
	wire[2:0] w_n173_0;
	wire[1:0] w_n173_1;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[2:0] w_n177_0;
	wire[1:0] w_n178_0;
	wire[1:0] w_n180_0;
	wire[2:0] w_n182_0;
	wire[2:0] w_n182_1;
	wire[2:0] w_n183_0;
	wire[1:0] w_n184_0;
	wire[1:0] w_n186_0;
	wire[1:0] w_n189_0;
	wire[2:0] w_n191_0;
	wire[2:0] w_n192_0;
	wire[2:0] w_n195_0;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[1:0] w_n198_0;
	wire[2:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n208_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n211_0;
	wire[2:0] w_n214_0;
	wire[2:0] w_n216_0;
	wire[1:0] w_n216_1;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n226_0;
	wire[2:0] w_n242_0;
	wire[2:0] w_n242_1;
	wire[2:0] w_n242_2;
	wire[1:0] w_n243_0;
	wire[1:0] w_n249_0;
	wire[2:0] w_n258_0;
	wire[2:0] w_n265_0;
	wire[2:0] w_n265_1;
	wire[1:0] w_n265_2;
	wire[1:0] w_n274_0;
	wire[2:0] w_n278_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n280_0;
	wire[2:0] w_n282_0;
	wire[1:0] w_n282_1;
	wire[1:0] w_n286_0;
	wire[2:0] w_n287_0;
	wire[1:0] w_n287_1;
	wire[1:0] w_n288_0;
	wire[2:0] w_n291_0;
	wire[1:0] w_n291_1;
	wire[1:0] w_n292_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n294_0;
	wire[1:0] w_n297_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n307_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n316_0;
	wire[2:0] w_n317_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n329_0;
	wire[1:0] w_n341_0;
	wire w_dff_B_gRoE5hj54_0;
	wire w_dff_B_217tmLfb0_0;
	wire w_dff_B_oHQ6x86A1_0;
	wire w_dff_B_4hfbee0s3_0;
	wire w_dff_B_xdFdkSUS6_0;
	wire w_dff_B_CRDpuNq14_0;
	wire w_dff_B_Wmu07nX56_0;
	wire w_dff_B_EOM0QiK69_0;
	wire w_dff_A_vZtyeN6G0_0;
	wire w_dff_A_qF97oLAq4_0;
	wire w_dff_B_yzKj40tv6_0;
	wire w_dff_B_289zX16p1_0;
	wire w_dff_B_GpDgQbzg3_0;
	wire w_dff_B_u34d1zbb2_0;
	wire w_dff_B_apkQf78x5_0;
	wire w_dff_B_8bptot6U4_1;
	wire w_dff_B_8jT7SjKR1_1;
	wire w_dff_B_m3WdSuYS8_1;
	wire w_dff_B_xoFZ9m0Q5_1;
	wire w_dff_B_5rdrazH21_1;
	wire w_dff_B_wrzresxM1_1;
	wire w_dff_B_B0PUDSaL1_1;
	wire w_dff_B_4Ubn4dbK3_1;
	wire w_dff_B_PbRPsO087_1;
	wire w_dff_B_iCce1xkd1_1;
	wire w_dff_B_KLJ5GnLK6_1;
	wire w_dff_B_5lrRqkCa5_1;
	wire w_dff_B_XZG5oczu4_0;
	wire w_dff_B_fScDFGmE2_0;
	wire w_dff_B_RbllD0ED1_0;
	wire w_dff_B_2bokdNiJ8_0;
	wire w_dff_B_SMY5Hzsc2_0;
	wire w_dff_B_PgBXu2QW0_0;
	wire w_dff_B_yleaMZuA9_0;
	wire w_dff_B_Zgj2cefF6_0;
	wire w_dff_B_0QkUNGRR8_0;
	wire w_dff_B_Q1dCM7WX8_0;
	wire w_dff_B_pPDCAFuE9_0;
	wire w_dff_B_IdsyYkH62_0;
	wire w_dff_B_eRpUBvpO3_0;
	wire w_dff_B_dZJonO2V5_0;
	wire w_dff_A_tghaUmpO5_1;
	wire w_dff_A_SPJlyURP8_1;
	wire w_dff_A_cakV6Asy8_1;
	wire w_dff_A_7k7rpdAV8_1;
	wire w_dff_A_fGqdGEo11_1;
	wire w_dff_A_jqUECqvU3_1;
	wire w_dff_A_kfHkVYdZ7_1;
	wire w_dff_A_wp6dSsHc0_1;
	wire w_dff_A_2e1PIBh61_1;
	wire w_dff_A_CltLlal05_1;
	wire w_dff_A_UDBtD4919_1;
	wire w_dff_A_753kcTCD8_1;
	wire w_dff_A_fcy4FWCD2_1;
	wire w_dff_A_bbOLXKZv3_1;
	wire w_dff_A_p6LfYgvw2_1;
	wire w_dff_A_mYKh4gra4_1;
	wire w_dff_A_XWPLXkbd7_1;
	wire w_dff_A_OvCn3US17_1;
	wire w_dff_A_tCsfNudJ3_1;
	wire w_dff_A_DVFHJ7Yf3_1;
	wire w_dff_A_geUV8zZN0_1;
	wire w_dff_A_hBhBAH5X3_1;
	wire w_dff_A_S0EBWjgW5_1;
	wire w_dff_A_kYJkkiDr6_1;
	wire w_dff_A_zJkIfS6s9_1;
	wire w_dff_A_qS4IVq449_1;
	wire w_dff_A_NLCYjfDY7_1;
	wire w_dff_A_Kb9lV6dn4_1;
	wire w_dff_A_EG8S5HFF4_1;
	wire w_dff_A_scQnXMZO7_1;
	wire w_dff_A_UA7Si7RF3_1;
	wire w_dff_A_qxF7e5cA0_1;
	wire w_dff_A_aMP8TxdD8_2;
	wire w_dff_A_RJpXreUj8_2;
	wire w_dff_A_SzIJBEkJ2_2;
	wire w_dff_A_iHdRgjGT8_2;
	wire w_dff_A_c60Amz7F7_2;
	wire w_dff_A_LawalTON3_2;
	wire w_dff_A_662gdWoi6_2;
	wire w_dff_A_y7T4zg6q8_2;
	wire w_dff_A_aU4dkGcP3_2;
	wire w_dff_A_TXnEezUI4_2;
	wire w_dff_A_BdKpp2w27_2;
	wire w_dff_A_VK7IZjKm2_2;
	wire w_dff_A_glg6sRqQ9_2;
	wire w_dff_A_Fr9tkfCD7_2;
	wire w_dff_A_50hE6mO46_2;
	wire w_dff_A_gipLDijG6_2;
	wire w_dff_A_eA2euOQv1_2;
	wire w_dff_A_5FhJvPGZ3_0;
	wire w_dff_A_2LxxnF2Y5_1;
	wire w_dff_B_oDFlLFrH6_1;
	wire w_dff_B_kkZGT5ex4_1;
	wire w_dff_B_xpkfFFE45_1;
	wire w_dff_B_jqqewpTn7_1;
	wire w_dff_B_K1oilr9n8_1;
	wire w_dff_B_ME0ctDw45_1;
	wire w_dff_B_2i56dJIx9_1;
	wire w_dff_B_k5H5qfgk9_1;
	wire w_dff_B_ca6pTKAa9_1;
	wire w_dff_B_Q4JEGFuY1_1;
	wire w_dff_B_AeyW46c71_1;
	wire w_dff_B_BJrzF2mA7_1;
	wire w_dff_B_bnANAjms4_0;
	wire w_dff_B_uViSEPFG6_0;
	wire w_dff_B_Tof3qMPu7_0;
	wire w_dff_B_1LrVve8r9_0;
	wire w_dff_B_NMgCGL556_0;
	wire w_dff_B_f95KTXUO2_0;
	wire w_dff_B_vlrt9UZ56_0;
	wire w_dff_B_xlvujJv19_0;
	wire w_dff_B_KVJyetJt7_0;
	wire w_dff_B_SM8ao1kl0_0;
	wire w_dff_B_fUpP4j4k8_0;
	wire w_dff_B_0q1XVR3r5_0;
	wire w_dff_B_LxmA6KS07_0;
	wire w_dff_B_CIDRaylk5_0;
	wire w_dff_B_YKHt5J0m8_1;
	wire w_dff_B_0LxZ9BDq7_1;
	wire w_dff_B_mg6vrPOX5_1;
	wire w_dff_B_50NgK2HR5_1;
	wire w_dff_B_sMOGxZUK7_2;
	wire w_dff_A_N5usaIeo9_1;
	wire w_dff_B_d1LbOOHB1_2;
	wire w_dff_A_mbPiTqZQ8_2;
	wire w_dff_A_mDT284LI8_2;
	wire w_dff_B_baiLUCyu9_3;
	wire w_dff_B_UvX1D9mq7_3;
	wire w_dff_B_CBkZFcZr1_0;
	wire w_dff_B_BlbbzFwu8_0;
	wire w_dff_B_fjvq7sK88_0;
	wire w_dff_B_8XGhWZXF1_0;
	wire w_dff_B_rl3VHiSm3_0;
	wire w_dff_B_Pcqve8FC6_0;
	wire w_dff_B_dlKiSWxK3_0;
	wire w_dff_B_cbHEKBl85_0;
	wire w_dff_B_YFxpDKCm0_0;
	wire w_dff_B_R1AXzCN50_0;
	wire w_dff_B_Hmziks3v6_0;
	wire w_dff_B_7zCrDNGV5_0;
	wire w_dff_B_asktv9BC0_0;
	wire w_dff_B_GOGYS8gI2_0;
	wire w_dff_B_7U5xAF7x3_0;
	wire w_dff_B_6iqi2rmt3_0;
	wire w_dff_B_G6eqx5cE5_0;
	wire w_dff_B_O3xIvpoG1_0;
	wire w_dff_B_jz97CtEX7_0;
	wire w_dff_B_vE5mbV9l5_0;
	wire w_dff_B_UjTeNUhL0_0;
	wire w_dff_B_brPlIuhZ1_0;
	wire w_dff_B_jMb14Fsk5_0;
	wire w_dff_B_QvNXZIlv1_0;
	wire w_dff_B_M1X8Cc2u7_0;
	wire w_dff_B_XytGs9et4_0;
	wire w_dff_B_WoMQU8Xr6_1;
	wire w_dff_B_ARLySCip4_1;
	wire w_dff_B_L52U40XV7_1;
	wire w_dff_A_92hYar444_1;
	wire w_dff_A_5ld2p0Q47_2;
	wire w_dff_A_p4wmA6dm0_1;
	wire w_dff_A_eXF0yj0D6_1;
	wire w_dff_A_jRuMaBaC7_1;
	wire w_dff_A_lWXx1Z5k6_2;
	wire w_dff_A_GlRQ3DSW3_1;
	wire w_dff_A_e4tCZxkY8_0;
	wire w_dff_A_cgR5SqR31_2;
	wire w_dff_A_ESH28Yld7_0;
	wire w_dff_A_IKnNahbU2_1;
	wire w_dff_B_mZMqktea3_2;
	wire w_dff_A_t0AN5XoL1_0;
	wire w_dff_A_b8HLrhFj1_2;
	wire w_dff_A_nT7IT46z9_0;
	wire w_dff_A_474pC7iS8_2;
	wire w_dff_B_vhhNAn034_3;
	wire w_dff_B_l6WeeIPA1_3;
	wire w_dff_A_WRKgB4gP3_1;
	wire w_dff_A_DGIu3rtn2_2;
	wire w_dff_B_3funJieQ8_0;
	wire w_dff_B_rHg0aR1x2_0;
	wire w_dff_B_xdvJCgyA3_0;
	wire w_dff_B_sChwiXBc3_0;
	wire w_dff_B_YghbJD1r6_0;
	wire w_dff_B_JTOIhjbR0_0;
	wire w_dff_B_whwpl6tL4_0;
	wire w_dff_B_WKEiH8V11_0;
	wire w_dff_B_RJolY06a7_0;
	wire w_dff_B_nDtIyK1b5_0;
	wire w_dff_B_CezhDRNi8_0;
	wire w_dff_B_lAgyn7Xj9_0;
	wire w_dff_B_8cIoaHl79_0;
	wire w_dff_B_M8qScDlO8_0;
	wire w_dff_B_rRqdFC7O3_0;
	wire w_dff_A_Ob9VAU6x7_1;
	wire w_dff_A_ysFF107H1_1;
	wire w_dff_A_Et1FL7JO8_1;
	wire w_dff_A_1Nrd7bdF7_1;
	wire w_dff_A_CSzVkNdn9_1;
	wire w_dff_A_6j4EvXZe3_1;
	wire w_dff_A_OLB7P6zY3_1;
	wire w_dff_A_ktdHEVxd8_1;
	wire w_dff_A_ZwYm77281_1;
	wire w_dff_A_X2QLLxGJ3_1;
	wire w_dff_A_4XJfn4QY0_1;
	wire w_dff_A_LSYqAxwU5_1;
	wire w_dff_A_9BVGgBsK6_1;
	wire w_dff_A_pVWF1xs27_1;
	wire w_dff_A_tjfRjIee7_1;
	wire w_dff_A_xqcT2hvA9_1;
	wire w_dff_A_Y0O5LEFn9_1;
	wire w_dff_A_BRjINC0z0_2;
	wire w_dff_A_4uYM1mso0_2;
	wire w_dff_A_VaBScGfd5_2;
	wire w_dff_A_YoVImA6k2_2;
	wire w_dff_A_kGodJQwH7_2;
	wire w_dff_A_goLhS2s04_2;
	wire w_dff_A_KrMuT1pJ3_2;
	wire w_dff_A_aAn6CQMd5_2;
	wire w_dff_A_PbAlEzDK4_2;
	wire w_dff_A_ToiQrkkz7_2;
	wire w_dff_A_JFEL1nUo3_2;
	wire w_dff_A_rclqD4ZQ2_2;
	wire w_dff_A_Gyoi4zx37_2;
	wire w_dff_A_rafw39099_2;
	wire w_dff_A_4y5XQRZL7_2;
	wire w_dff_A_22myod8p8_2;
	wire w_dff_A_pWNy4AKp6_2;
	wire w_dff_B_2X3F5Utf0_1;
	wire w_dff_B_JXxE9l7T2_1;
	wire w_dff_A_xEIhDbgd1_0;
	wire w_dff_A_C9ZSpTRT0_1;
	wire w_dff_A_DevZQJIz3_2;
	wire w_dff_A_LVBGMoP22_0;
	wire w_dff_A_QKfCqza18_2;
	wire w_dff_B_ujxpdS7E3_0;
	wire w_dff_B_NgPS3SEX2_0;
	wire w_dff_B_twwOpmxt5_0;
	wire w_dff_A_jo4ZeTVu3_1;
	wire w_dff_A_iSuFEqde4_0;
	wire w_dff_A_AVw7lWSl2_2;
	wire w_dff_A_Yxw5h3ar9_1;
	wire w_dff_A_ceuQN59g7_0;
	wire w_dff_A_kAaKGw3K8_0;
	wire w_dff_A_qupKCXvj3_0;
	wire w_dff_A_sTeTl9j90_2;
	wire w_dff_A_XUkfqiMS7_2;
	wire w_dff_A_wPdwgXWI3_2;
	wire w_dff_A_Kq7nAxjJ6_2;
	wire w_dff_A_LuAz3Zoz4_0;
	wire w_dff_A_j1v6xOuW7_1;
	wire w_dff_A_pL9aPxaf8_1;
	wire w_dff_A_NybkuwfE7_2;
	wire w_dff_A_YxtIsUQ09_0;
	wire w_dff_A_dG3pUUhf3_1;
	wire w_dff_B_TYA0jWKs3_2;
	wire w_dff_A_s5YjsonR8_1;
	wire w_dff_A_xQT8wLcD4_1;
	wire w_dff_A_wHFsuuiJ8_0;
	wire w_dff_B_2T9zAfDd3_2;
	wire w_dff_A_D3qXC8054_2;
	wire w_dff_A_wQssL4Lw9_2;
	wire w_dff_A_hoRXZfFF0_2;
	wire w_dff_A_GAFQXiQk6_2;
	wire w_dff_B_f6Q2iOXQ1_1;
	wire w_dff_B_789dvlrH7_1;
	wire w_dff_B_zoWnA3Sw9_1;
	wire w_dff_B_2JLpDrk81_1;
	wire w_dff_B_gbbLE1r79_1;
	wire w_dff_A_yfhcaq8P3_1;
	wire w_dff_A_a9FOPwLV5_1;
	wire w_dff_A_soEHyxz21_1;
	wire w_dff_A_yMjaBLlH6_2;
	wire w_dff_A_6gvA7Kvb2_0;
	wire w_dff_A_MX6iKdHZ7_1;
	wire w_dff_A_EZQQlWfd2_2;
	wire w_dff_B_yxV8UGaj6_1;
	wire w_dff_B_Y4OnDzFr3_1;
	wire w_dff_B_WJrPwGVT1_1;
	wire w_dff_B_IfHaIX4n4_1;
	wire w_dff_B_Lhkdwcf79_1;
	wire w_dff_A_KOS7OcBZ2_1;
	wire w_dff_A_FJ51mBDe1_0;
	wire w_dff_A_zhsHfnEm0_1;
	wire w_dff_B_uzR4OQuH0_1;
	wire w_dff_B_2RgNAlMZ2_1;
	wire w_dff_B_MWxUAb5E4_1;
	wire w_dff_B_C0kAeFOd6_1;
	wire w_dff_B_3kB9E9WJ2_1;
	wire w_dff_A_UYistIdV0_0;
	wire w_dff_A_0fWTY5xz5_0;
	wire w_dff_A_BjEMlTet3_0;
	wire w_dff_A_3AxcHWoe5_0;
	wire w_dff_A_YCztvHnA2_0;
	wire w_dff_A_DcxoOiIG4_0;
	wire w_dff_A_omNvXYFU5_0;
	wire w_dff_A_9RO2IyyX7_0;
	wire w_dff_A_Q8zLMNXk4_0;
	wire w_dff_A_MvPLNjpo1_0;
	wire w_dff_A_PNR7F9bp4_0;
	wire w_dff_A_7QDaXC2d3_0;
	wire w_dff_A_DCDL6rW75_0;
	wire w_dff_A_7WMoCQIU0_1;
	wire w_dff_A_gjbdkYIb0_0;
	wire w_dff_A_0zhemYdL4_0;
	wire w_dff_A_khodaI6M6_0;
	wire w_dff_A_Gv8l8Q3L8_0;
	wire w_dff_A_ag7Im9mg7_0;
	wire w_dff_A_b7e3vnuK8_0;
	wire w_dff_A_DWLzeQDI0_0;
	wire w_dff_A_M2CmPuwm5_0;
	wire w_dff_A_sXfm6t2m7_0;
	wire w_dff_A_H0R0gBJm9_0;
	wire w_dff_A_ihMVvcDN0_0;
	wire w_dff_A_Hf6EEOXC0_0;
	wire w_dff_A_pfFUrYvS8_0;
	wire w_dff_A_MFR2jh6Q4_0;
	wire w_dff_A_r7RVUuaW0_0;
	wire w_dff_A_hi8HOVFL6_0;
	wire w_dff_A_Tbf7fEPQ5_2;
	wire w_dff_A_sg68VMId5_2;
	wire w_dff_A_PFpzELJV4_2;
	wire w_dff_A_qyPaySJa3_2;
	wire w_dff_A_1FjSXV9z0_2;
	wire w_dff_A_yjGMR8qv0_2;
	wire w_dff_A_iPJCIki71_1;
	wire w_dff_A_viYe8xIr3_1;
	wire w_dff_A_IDXMZJm00_2;
	wire w_dff_A_bFIRqKpw9_2;
	wire w_dff_A_LFpjap0v7_1;
	wire w_dff_A_tQ6X6L0b4_1;
	wire w_dff_A_hj8rotjC3_1;
	wire w_dff_A_zW9L4dHS9_2;
	wire w_dff_A_S133haJG2_2;
	wire w_dff_A_23L3vLrA3_2;
	wire w_dff_A_ILbxSRX01_1;
	wire w_dff_A_u2vrMGRA8_1;
	wire w_dff_A_gwtCXaDD2_1;
	wire w_dff_A_2zVWGoBz7_1;
	wire w_dff_A_0hn9qmfX6_0;
	wire w_dff_A_Z9ohuSKm0_0;
	wire w_dff_A_dn9w75tJ3_0;
	wire w_dff_A_zyA0znkD5_0;
	wire w_dff_A_NrlRSbuI4_0;
	wire w_dff_A_igCyGVkT9_0;
	wire w_dff_A_lGXE1MWv3_0;
	wire w_dff_A_sDXGCA2C6_0;
	wire w_dff_A_zzUgZ3Vr9_0;
	wire w_dff_A_WXRgklfM4_0;
	wire w_dff_A_FEe6EmbO6_0;
	wire w_dff_A_V7pe8dpK8_0;
	wire w_dff_A_dOdQglT95_0;
	wire w_dff_B_dEj9vy825_1;
	wire w_dff_A_kSftgAv93_1;
	wire w_dff_B_gGE3uEGs4_0;
	wire w_dff_B_C21Cr2AB5_0;
	wire w_dff_A_jjWIrSHE2_0;
	wire w_dff_A_UANKoWfV5_1;
	wire w_dff_A_HTLSczVE8_1;
	wire w_dff_A_Big4gnsf9_2;
	wire w_dff_A_mPRuzlGc6_2;
	wire w_dff_B_hVsy3OE97_3;
	wire w_dff_B_836m1ysa9_3;
	wire w_dff_A_jcYedj8v0_0;
	wire w_dff_A_3xNgarSq0_0;
	wire w_dff_A_Sqme8lOR8_1;
	wire w_dff_A_VCwZPWoZ7_1;
	wire w_dff_A_E0i33Pnj3_1;
	wire w_dff_A_Pc05VXXJ3_1;
	wire w_dff_A_VVcpvPLv4_1;
	wire w_dff_A_YUuSe0jM1_2;
	wire w_dff_A_RINZHuL81_2;
	wire w_dff_A_d2xjLCcJ0_2;
	wire w_dff_A_Vk0unUv63_2;
	wire w_dff_A_s4HEiENx9_2;
	wire w_dff_A_akdZEYzP7_1;
	wire w_dff_A_LMQzXh8Y3_2;
	wire w_dff_B_9df6Tjnu5_3;
	wire w_dff_B_yQ6CoJCA8_1;
	wire w_dff_B_hbFeXRny0_1;
	wire w_dff_B_e8gTMXUE6_1;
	wire w_dff_B_DtM3fqRY8_1;
	wire w_dff_B_fW3ODDb64_1;
	wire w_dff_A_nTA8dc2J4_0;
	wire w_dff_A_arDw1qDP6_0;
	wire w_dff_A_KdvZQnOx3_0;
	wire w_dff_A_vLUjnDP74_0;
	wire w_dff_A_HRu0UsxV7_0;
	wire w_dff_A_NOTBondg0_0;
	wire w_dff_A_2Poa2mue9_0;
	wire w_dff_A_Ys8MZafy6_0;
	wire w_dff_A_Jf4H14860_0;
	wire w_dff_A_IxYExDvf8_0;
	wire w_dff_A_WcXlRiwk9_0;
	wire w_dff_A_j4eWW6fM7_0;
	wire w_dff_A_0hIR9ZAy8_0;
	wire w_dff_A_Kj646pdm1_0;
	wire w_dff_A_3vWj2P5T0_0;
	wire w_dff_A_ykrmFzzJ4_0;
	wire w_dff_A_J6uPRhhx5_0;
	wire w_dff_A_U9Pq5whE9_0;
	wire w_dff_A_0fKSYsEz7_0;
	wire w_dff_A_gbWYWOX61_0;
	wire w_dff_A_seO9mZAi9_0;
	wire w_dff_A_K6pOlWRz7_0;
	wire w_dff_A_RPYC76iM6_0;
	wire w_dff_A_X8nYf7Ib2_0;
	wire w_dff_A_WFEKeYOX3_0;
	wire w_dff_A_gORIwm874_0;
	wire w_dff_A_PZfsSMQf1_0;
	wire w_dff_A_OxcboRLa7_0;
	wire w_dff_A_lgVNsBUw3_1;
	wire w_dff_A_2igJotMc4_0;
	wire w_dff_A_b7ZsRcXM4_0;
	wire w_dff_A_qtC2uJTM6_0;
	wire w_dff_A_zUO6yFtc2_0;
	wire w_dff_A_XiNJVHv52_0;
	wire w_dff_A_kc67abS97_0;
	wire w_dff_A_SdbcqVAH1_0;
	wire w_dff_A_S7jz1DP98_0;
	wire w_dff_A_aDnl2Ive5_0;
	wire w_dff_A_C8nH7f4g9_0;
	wire w_dff_A_e09HX4jy3_0;
	wire w_dff_A_XYgP6YE56_2;
	wire w_dff_A_hek1xz6t0_2;
	wire w_dff_A_0ikeNFih7_1;
	wire w_dff_A_Sc72a3VD2_1;
	wire w_dff_A_JDwHL18b8_2;
	wire w_dff_A_t7DcwMMq3_2;
	wire w_dff_A_uoALZ0xa1_2;
	wire w_dff_A_cLJcyHSe6_2;
	wire w_dff_A_RIZzNKuy0_2;
	wire w_dff_A_tt3a3Kk34_2;
	wire w_dff_A_lLBd2Mlm2_2;
	wire w_dff_B_zfUoBTQh6_0;
	wire w_dff_A_vwNAnwBi9_0;
	wire w_dff_A_zvGreQTX8_0;
	wire w_dff_A_8Fnq0ajR2_0;
	wire w_dff_A_gWODHQOU4_0;
	wire w_dff_A_u1nqCuJj4_0;
	wire w_dff_A_r5jycrNU8_0;
	wire w_dff_A_B6ByFUkx9_0;
	wire w_dff_A_vApP2TkF9_0;
	wire w_dff_A_q2lv8LCn5_0;
	wire w_dff_A_XuHVOHfK9_0;
	wire w_dff_A_3q3QRkbk6_0;
	wire w_dff_A_LQSVngut4_0;
	wire w_dff_A_4bB5OuEG5_0;
	wire w_dff_A_smsN2Iox9_0;
	wire w_dff_A_HAwpuHLL6_0;
	wire w_dff_B_rSPAN7jr8_0;
	wire w_dff_B_Riq3223L9_0;
	wire w_dff_A_w6sVhHoO8_0;
	wire w_dff_A_wvDoVApv4_0;
	wire w_dff_A_RWSKkCu97_0;
	wire w_dff_A_sGIdZOwg1_0;
	wire w_dff_A_eMpst64i5_0;
	wire w_dff_A_uhr4LGSY7_0;
	wire w_dff_A_4fhJFv3b4_0;
	wire w_dff_A_MmjVKcDN1_0;
	wire w_dff_A_eqj3wAXU6_0;
	wire w_dff_A_aLnQ2UFa6_0;
	wire w_dff_A_dmY5xswP2_0;
	wire w_dff_B_j1EcKPlT8_0;
	wire w_dff_A_5SAgPiya6_0;
	wire w_dff_A_g4KXJQXo9_0;
	wire w_dff_A_VhUWGECe0_0;
	wire w_dff_A_qL334ohz8_0;
	wire w_dff_A_2lQI52uQ4_0;
	wire w_dff_A_4utpvD5Q7_0;
	wire w_dff_A_uto0gISE3_0;
	wire w_dff_A_lTh5TlsS4_0;
	wire w_dff_A_GbRVivJi6_0;
	wire w_dff_A_3C7b3KkZ9_0;
	wire w_dff_A_8ccLeRGo3_0;
	wire w_dff_A_pltr9Sy91_2;
	wire w_dff_A_KAFUf0ie5_0;
	wire w_dff_A_bMLvj4vK6_0;
	wire w_dff_A_isC4nyop5_0;
	wire w_dff_A_1OCK4Hfe3_0;
	wire w_dff_A_FpjEbNeu5_0;
	wire w_dff_A_w6UiwGWK1_0;
	wire w_dff_A_UDv47Jyb2_0;
	wire w_dff_A_tMBLsMwz9_0;
	wire w_dff_A_HcNUUNC09_0;
	wire w_dff_A_a9np6C7j6_0;
	wire w_dff_A_iU37nXPr2_0;
	wire w_dff_B_lRv8V3uU9_1;
	wire w_dff_A_CqMkEHCF9_0;
	wire w_dff_A_bCHLZywt4_0;
	wire w_dff_A_Xm3AFnP14_0;
	wire w_dff_A_ramVYyqn5_0;
	wire w_dff_A_JpljhAPX5_0;
	wire w_dff_A_oaRh1Isg0_0;
	wire w_dff_A_EWEC3qSB8_0;
	wire w_dff_A_vajKnaec8_0;
	wire w_dff_A_gNVfRazD7_2;
	wire w_dff_A_VLPQj9N95_2;
	wire w_dff_A_jjicVHTu2_2;
	wire w_dff_A_S5z7eyd04_2;
	wire w_dff_A_HtXn5sey4_0;
	wire w_dff_A_mGkVDPT69_0;
	wire w_dff_A_Rkt191pb6_0;
	wire w_dff_A_a3stNVrJ1_2;
	wire w_dff_A_howrrxnu0_2;
	wire w_dff_A_Xxkx8BNO7_2;
	wire w_dff_A_kUpEp3qm3_2;
	wire w_dff_A_66Ajoyz44_2;
	wire w_dff_A_MBSKY7wZ0_1;
	wire w_dff_A_wymmlnrp4_1;
	wire w_dff_A_dBSwxGuH5_1;
	wire w_dff_A_2Owppcnm8_1;
	wire w_dff_A_IdGG1rts0_2;
	wire w_dff_A_n5rbimli5_2;
	wire w_dff_A_UjNvUUNS2_2;
	wire w_dff_A_zRemNt128_2;
	wire w_dff_A_2aGJKbXC9_2;
	wire w_dff_A_2Rq2Fr4M0_2;
	wire w_dff_A_itdnHQhG9_2;
	wire w_dff_A_Glw0nwvI2_2;
	wire w_dff_A_rcqTukSG5_2;
	wire w_dff_A_5djuqVFR4_0;
	wire w_dff_A_0sMTgjXs1_1;
	wire w_dff_A_ydXUKeDR6_0;
	wire w_dff_A_BinbQrpY8_0;
	wire w_dff_A_sB64z77S3_0;
	wire w_dff_A_jX8b1f1s6_1;
	wire w_dff_A_Ba13vm6k1_1;
	wire w_dff_A_WObRkVXM3_1;
	wire w_dff_A_Lj6B4xWL1_1;
	wire w_dff_A_4rPayeat6_1;
	wire w_dff_A_4kxpTksh5_1;
	wire w_dff_A_OzW7DTnm7_1;
	wire w_dff_A_Urd1DreW0_1;
	wire w_dff_A_CLhc1APU4_1;
	wire w_dff_A_PzMxH0kn3_1;
	wire w_dff_A_gjLME5Nz6_1;
	wire w_dff_A_5z0D4Avc7_1;
	wire w_dff_B_WXB1PzWk1_1;
	wire w_dff_B_OR4AFcGl9_1;
	wire w_dff_A_ny44Yxjq1_0;
	wire w_dff_A_t6Aqb92A9_0;
	wire w_dff_A_gmemrK8c4_0;
	wire w_dff_A_MxtWWakH8_0;
	wire w_dff_A_sp8c4X9D8_0;
	wire w_dff_A_ZD9dmgdA5_0;
	wire w_dff_A_N7knh9kF0_0;
	wire w_dff_A_DnZ0gSkA9_0;
	wire w_dff_A_aikiDzSt6_0;
	wire w_dff_A_bCg3G5HH0_0;
	wire w_dff_A_kods908k3_0;
	wire w_dff_A_yHCBM2o71_2;
	wire w_dff_A_4gro4Qq16_1;
	wire w_dff_A_MndoQkpc4_1;
	wire w_dff_A_O82f2qgK5_0;
	wire w_dff_A_9hXodets6_0;
	wire w_dff_A_IzmLdrPM4_0;
	wire w_dff_A_s9eyQzU52_0;
	wire w_dff_A_ijYW7ftR5_0;
	wire w_dff_A_nStjOTmZ5_0;
	wire w_dff_A_oaq1eUE38_0;
	wire w_dff_A_g1TcIJRt4_0;
	wire w_dff_A_7LILtQ9H7_0;
	wire w_dff_A_LA6PbRAi6_0;
	wire w_dff_A_tHxKLm443_0;
	wire w_dff_A_ZiHncPfI6_0;
	wire w_dff_A_ej3pzEcr5_0;
	wire w_dff_A_SXTVyYmQ3_0;
	wire w_dff_A_wF4hsBQF2_1;
	wire w_dff_A_i1Hwubp30_0;
	wire w_dff_A_aAnerfct9_0;
	wire w_dff_A_PAoRkGDN0_0;
	wire w_dff_A_Clgrptpj1_0;
	wire w_dff_A_v6chAHij5_0;
	wire w_dff_A_GcOqCF9K8_0;
	wire w_dff_A_Nyy2vzIP0_0;
	wire w_dff_A_O6B0a1403_0;
	wire w_dff_A_SeSyZGcX5_0;
	wire w_dff_A_iijTPlN86_0;
	wire w_dff_A_C8994UPm7_0;
	wire w_dff_A_rlIJPHfN1_1;
	wire w_dff_A_WndBmvHt3_1;
	wire w_dff_A_ARiPaSY28_0;
	wire w_dff_A_paWH26mO8_0;
	wire w_dff_A_oWK3JBLm4_0;
	wire w_dff_A_ANKfPbG39_0;
	wire w_dff_A_Z1iiLFEb2_0;
	wire w_dff_A_0FPz1Bmz4_0;
	wire w_dff_A_t7erJs8e7_0;
	wire w_dff_A_b0unMr1B5_0;
	wire w_dff_A_QBTBEDr06_0;
	wire w_dff_A_lGqwmx6k0_0;
	wire w_dff_B_pJ00iYd30_3;
	wire w_dff_A_2LDcOgv21_0;
	wire w_dff_A_gh9SyJsA6_0;
	wire w_dff_A_m86lGQxw3_0;
	wire w_dff_A_W2V6DUtM6_0;
	wire w_dff_A_WbCUFWBT6_0;
	wire w_dff_A_HM7cNEzm5_0;
	wire w_dff_A_LfoBj8Ja6_0;
	wire w_dff_A_vnKd2LCA2_0;
	wire w_dff_A_joXP8Esh0_0;
	wire w_dff_A_rPloaFkw3_0;
	wire w_dff_A_W6A9ZwZM7_0;
	wire w_dff_A_Mv9PS05C3_0;
	wire w_dff_A_6NzcPmKd8_0;
	wire w_dff_A_oF6pixnn9_0;
	wire w_dff_A_OepuZN8N2_0;
	wire w_dff_A_GoTNuIH95_0;
	wire w_dff_A_48hznqgR6_0;
	wire w_dff_A_hOBl3brz2_0;
	wire w_dff_A_vR3vijAC3_0;
	wire w_dff_A_JGwUCmuH4_0;
	wire w_dff_A_k0YkS6im8_0;
	wire w_dff_A_XBXSzFWV5_0;
	wire w_dff_A_mfxrm3Sh9_1;
	wire w_dff_A_GcLArIWj5_1;
	wire w_dff_A_AOQreN4t6_1;
	wire w_dff_A_GY65gK7N7_1;
	wire w_dff_A_ViEKZQb18_1;
	wire w_dff_A_YleF7ISi4_1;
	wire w_dff_A_YB1Nc0QZ0_1;
	wire w_dff_A_mWR2PQIy1_0;
	wire w_dff_A_VA5asiY78_0;
	wire w_dff_A_4KNi1YVI9_0;
	wire w_dff_A_K63yS8ea1_0;
	wire w_dff_A_XWmNXPPX1_0;
	wire w_dff_A_IACZD6388_0;
	wire w_dff_A_GPJKNxuc2_0;
	wire w_dff_A_A6t5laxm8_0;
	wire w_dff_A_DaKDpKmx2_0;
	wire w_dff_A_JOsJ6Rhk9_0;
	wire w_dff_A_KtTzOYmK8_0;
	wire w_dff_A_pyKFEhQI8_0;
	wire w_dff_A_KdXWk3gy3_0;
	wire w_dff_B_Bh3sPweE9_1;
	wire w_dff_B_UKEKbcmb4_1;
	wire w_dff_B_idvopbrR7_0;
	wire w_dff_A_lFvFyPPR1_1;
	wire w_dff_A_94f2hsQR2_1;
	wire w_dff_A_xSqjmXpx4_1;
	wire w_dff_A_j74IhGhE7_1;
	wire w_dff_A_7kYhQ0L47_1;
	wire w_dff_A_ACEK8Yt05_1;
	wire w_dff_A_4UCi0tU26_1;
	wire w_dff_A_zKzwhAVR1_1;
	wire w_dff_A_zdaY5l260_1;
	wire w_dff_A_NGqv4ogJ5_1;
	wire w_dff_A_FcIi9Brt1_1;
	wire w_dff_A_zeEAMW488_1;
	wire w_dff_A_TJajhCmD7_0;
	wire w_dff_A_CdrawaRy0_0;
	wire w_dff_A_C71pwByx9_0;
	wire w_dff_A_KBo7VCKl8_0;
	wire w_dff_A_eUXjmOwR6_0;
	wire w_dff_A_tYURWBIx1_0;
	wire w_dff_A_1krbR3pj6_0;
	wire w_dff_A_lW37oSFs1_0;
	wire w_dff_A_q7vpDMdE7_0;
	wire w_dff_A_D3wF8aWo3_0;
	wire w_dff_A_hpithpsj5_0;
	wire w_dff_A_Jw8eBKCr2_0;
	wire w_dff_A_uNHBq4bp3_0;
	wire w_dff_A_vPwzDTcv7_0;
	wire w_dff_A_PYdrpQmU8_0;
	wire w_dff_A_pWbL2WTr1_0;
	wire w_dff_A_fwFKgR1q5_0;
	wire w_dff_A_2FkRzDyw3_0;
	wire w_dff_A_nwUITX0C1_0;
	wire w_dff_A_ID4Pk6ml7_0;
	wire w_dff_A_jahA2CPO7_0;
	wire w_dff_A_tILj3M467_0;
	wire w_dff_A_TWcZ3hlV8_1;
	wire w_dff_A_vqQHzyQy5_2;
	wire w_dff_A_sCiPDOfo6_2;
	wire w_dff_A_e1THIr3i3_1;
	wire w_dff_A_h6dGnH6u5_0;
	wire w_dff_A_SU1pPER50_0;
	wire w_dff_A_Fk427TdG1_0;
	wire w_dff_A_x7rPlRLu2_0;
	wire w_dff_A_fXlHFcYu6_0;
	wire w_dff_A_9W0pmyp47_0;
	wire w_dff_A_zxqiynyj6_0;
	wire w_dff_A_mDgN9ZgF7_0;
	wire w_dff_A_kL1Z1Pm95_0;
	wire w_dff_A_kV9f1zVT7_0;
	wire w_dff_A_qJlt3UJN2_0;
	wire w_dff_A_7ka7thog0_0;
	wire w_dff_A_2bIecY3Y3_0;
	wire w_dff_A_YFHk7fnc7_0;
	wire w_dff_A_Ej80MD9W3_2;
	wire w_dff_B_hO9y6Zfl1_3;
	wire w_dff_B_NMvSU6qi8_3;
	wire w_dff_A_Uyxa1jdV3_0;
	wire w_dff_A_zkrzFq9t3_0;
	wire w_dff_A_K9SZtQG15_0;
	wire w_dff_A_cAq71eL22_0;
	wire w_dff_A_DMctQkqj2_0;
	wire w_dff_A_5kjPYsut1_0;
	wire w_dff_A_EPv2wLsB0_0;
	wire w_dff_A_mUg58g8w7_0;
	wire w_dff_A_Lqr4g2Ii4_0;
	wire w_dff_A_acBnNSvq5_0;
	wire w_dff_A_54YWHNz46_0;
	wire w_dff_A_8zc6us4R5_1;
	wire w_dff_A_AORReWib9_0;
	wire w_dff_A_KyWQvPab6_0;
	wire w_dff_A_Rzh3Lz0I1_0;
	wire w_dff_A_pF1zcXhi4_0;
	wire w_dff_A_rl57237d4_0;
	wire w_dff_A_pZkQA3H45_0;
	wire w_dff_A_spANxOh15_0;
	wire w_dff_A_qKeaOSgV5_0;
	wire w_dff_A_8K7YSytW6_0;
	wire w_dff_A_iOz0fSRG1_0;
	wire w_dff_A_julECBpF0_0;
	wire w_dff_A_ZgKH4qLv2_0;
	wire w_dff_A_1dOdWFbt4_0;
	wire w_dff_A_RvvqsymX1_0;
	wire w_dff_A_hIegGQQ95_0;
	wire w_dff_A_8I6G7J8J1_0;
	wire w_dff_A_A0OAUl0l0_0;
	wire w_dff_A_zM1WbSZ23_0;
	wire w_dff_A_PCdON3043_0;
	wire w_dff_A_EYRc5Jg54_0;
	wire w_dff_A_kHr6qwOO9_0;
	wire w_dff_A_6fVrQNeK2_0;
	wire w_dff_A_Ceh9Y6RA4_1;
	wire w_dff_A_zs8FWjcf8_0;
	wire w_dff_A_V4m9vpmB8_0;
	wire w_dff_A_QaqVoQ6i3_0;
	wire w_dff_A_N1JBoeja7_0;
	wire w_dff_A_Yhai2ikW0_2;
	wire w_dff_A_FLDsYRoa1_2;
	wire w_dff_A_6IOIBCTc9_2;
	wire w_dff_A_mcU4tgIv0_2;
	wire w_dff_A_2c3QfiNY0_0;
	wire w_dff_A_tiODlU1F4_0;
	wire w_dff_A_hOHbir0a9_0;
	wire w_dff_A_PDjWm0sn2_0;
	wire w_dff_A_oeZgErjw3_0;
	wire w_dff_A_rDDXlFen1_0;
	wire w_dff_A_vsKFgpCk8_0;
	wire w_dff_A_VAUH35qY0_0;
	wire w_dff_A_vTG6tajw1_0;
	wire w_dff_A_ucS4E2g80_0;
	wire w_dff_A_Jb8hfndA9_0;
	wire w_dff_A_bEVz6YNV4_0;
	wire w_dff_A_VoKtbupI5_0;
	wire w_dff_A_pjFHUqEz0_0;
	wire w_dff_A_pIvRJMFZ7_0;
	wire w_dff_A_dzFctr5t1_0;
	wire w_dff_A_T4qmQgTn8_0;
	wire w_dff_A_fKDY7Nsc9_0;
	wire w_dff_A_M02w6KUf3_1;
	wire w_dff_A_72LYaYfb0_1;
	wire w_dff_A_y4VWZT022_1;
	wire w_dff_A_lm7bARAI1_1;
	wire w_dff_A_VctRwhUr7_1;
	wire w_dff_A_l0eGAroD5_1;
	wire w_dff_A_H8dpCByK6_1;
	wire w_dff_B_3KlfMBQA9_3;
	wire w_dff_B_8tesdH5w4_3;
	wire w_dff_B_EhBHDecs2_3;
	wire w_dff_B_uKTTEheB9_3;
	wire w_dff_B_zc3zs5xo6_3;
	wire w_dff_B_Zwqu0bqe7_3;
	wire w_dff_B_sJBTHqkT3_3;
	wire w_dff_B_8ar9O2Ie3_3;
	wire w_dff_B_xfDn2R9L6_3;
	wire w_dff_B_QOUfgPnZ1_3;
	wire w_dff_B_U7vSbnKH4_3;
	wire w_dff_B_DqelCsKJ1_3;
	wire w_dff_B_D4fHQvLF9_3;
	wire w_dff_B_yNpts7NY5_3;
	wire w_dff_B_S7LHnDBT9_3;
	wire w_dff_B_YCfBBzZ70_3;
	wire w_dff_A_lOKFUup95_0;
	wire w_dff_A_6IiluKjv0_0;
	wire w_dff_A_P78E6ndu2_0;
	wire w_dff_A_OO4BfbEG7_0;
	wire w_dff_A_xipyZCpr9_0;
	wire w_dff_A_ziVXBFSx5_0;
	wire w_dff_A_ZHuVen6B4_0;
	wire w_dff_A_zpFHcZRZ8_0;
	wire w_dff_A_q69mUsiW8_0;
	wire w_dff_A_ddiVUbg04_0;
	wire w_dff_A_rh9P2G2O0_0;
	wire w_dff_A_2A6pMAIZ8_0;
	wire w_dff_A_ynZYaNpE5_0;
	wire w_dff_A_ytvGwuEO0_0;
	wire w_dff_A_KXfeyVnS8_0;
	wire w_dff_A_Pm1Qpj9M2_1;
	wire w_dff_A_R0LuugEo0_1;
	wire w_dff_A_F2zpO55S0_1;
	wire w_dff_A_B43PHoVe5_1;
	wire w_dff_A_qGTl746B6_1;
	wire w_dff_A_UVsxiAya9_1;
	wire w_dff_A_Iv2EG6hp6_1;
	wire w_dff_A_COnjRR6S4_1;
	wire w_dff_A_MNLVDXSy7_1;
	wire w_dff_A_ZgTAUQXH8_1;
	wire w_dff_A_iaZIgbic2_1;
	wire w_dff_A_UGqxG0g45_1;
	wire w_dff_A_GgAyF5bf5_2;
	wire w_dff_A_gL2fNxA12_2;
	wire w_dff_A_9j5upJDu4_2;
	wire w_dff_A_ffBxmw9z8_2;
	wire w_dff_A_WVS9tnBF5_2;
	wire w_dff_A_t6SN8CFU6_2;
	wire w_dff_A_PgL2PPIp4_2;
	wire w_dff_A_ymkJJMVU8_2;
	wire w_dff_A_HcSQSjMQ5_2;
	wire w_dff_A_qHM1NRBl1_2;
	wire w_dff_A_oPrdO45e4_2;
	wire w_dff_A_55uuqk1i8_2;
	wire w_dff_A_l4P3fljX2_2;
	wire w_dff_A_e8jTiCF58_2;
	wire w_dff_A_hiFdIg9Q8_2;
	wire w_dff_A_B6LlEjr60_1;
	wire w_dff_A_6i0kJJaO8_1;
	wire w_dff_A_jDjCFC3n9_1;
	wire w_dff_A_DiTXsm7e1_1;
	wire w_dff_A_RjD8HaVJ3_1;
	wire w_dff_A_WAk2OABQ1_1;
	wire w_dff_A_lRkGRM7K0_1;
	wire w_dff_A_7YDbiEcs0_1;
	wire w_dff_A_2OnvTU1x7_1;
	wire w_dff_A_PXeVG97y2_1;
	wire w_dff_A_kTVJeEXa9_1;
	wire w_dff_A_6BJkxyXk5_1;
	wire w_dff_A_nmLjS0oG8_1;
	wire w_dff_A_QdnxJQn89_1;
	wire w_dff_A_xvDgcW3l1_1;
	wire w_dff_A_GJtCJ9al0_1;
	wire w_dff_A_SjzwPv5X2_2;
	wire w_dff_B_PjuaBNu04_3;
	wire w_dff_A_1HIeDp7r2_2;
	wire w_dff_A_dpSwxm545_0;
	wire w_dff_A_mbF8eUps7_0;
	wire w_dff_A_HxWVCLTv5_0;
	wire w_dff_A_g7FwyZWy5_0;
	wire w_dff_A_6FZWLiIJ4_0;
	wire w_dff_A_QwsrG7Az8_0;
	wire w_dff_A_Cxg7nzTV6_0;
	wire w_dff_A_jzkZ6mNp7_2;
	wire w_dff_A_MHUHYXTa4_0;
	wire w_dff_A_JswjQ0108_0;
	wire w_dff_A_0o8yrJiR2_0;
	wire w_dff_A_8x2BsPps5_0;
	wire w_dff_A_q9TbdOh14_0;
	wire w_dff_A_uS4mnpUH5_0;
	wire w_dff_A_s1Tj0OV23_0;
	wire w_dff_A_25G69Rjr9_2;
	wire w_dff_A_10Sdgrvs1_0;
	wire w_dff_A_FaslhWba5_0;
	wire w_dff_A_1DTnCy7r5_0;
	wire w_dff_A_1ELhKcnn8_0;
	wire w_dff_A_SMhhcGkr1_0;
	wire w_dff_A_iSJ9zS557_0;
	wire w_dff_A_KvuzvACb3_0;
	wire w_dff_A_z3wcJUFY4_2;
	wire w_dff_A_fMbK2QzZ0_0;
	wire w_dff_A_Wo1G8lMq3_0;
	wire w_dff_A_7CQajTHE1_0;
	wire w_dff_A_8lqg625L3_0;
	wire w_dff_A_saG0aem95_0;
	wire w_dff_A_LOMJq8wV4_0;
	wire w_dff_A_mHbDUKf35_0;
	wire w_dff_A_WlpV7S0I3_2;
	wire w_dff_A_VoTwe0xA1_0;
	wire w_dff_A_a5uXxZFv3_0;
	wire w_dff_A_QdCzHjlB6_0;
	wire w_dff_A_So69hqCf3_0;
	wire w_dff_A_MiPx4MOj1_0;
	wire w_dff_A_CdOhcoDh7_0;
	wire w_dff_A_0q5J7Jwn5_0;
	wire w_dff_A_WaS3U3aF1_2;
	wire w_dff_A_tGyO216O7_0;
	wire w_dff_A_eU4F72ku8_0;
	wire w_dff_A_0luz7jIX0_0;
	wire w_dff_A_iSjbBr9t4_0;
	wire w_dff_A_iF7uQ93P1_0;
	wire w_dff_A_NwXul5tS7_0;
	wire w_dff_A_jnawhvD27_0;
	wire w_dff_A_kpZMc0eW0_2;
	wire w_dff_A_3b77LA202_0;
	wire w_dff_A_JFjWkVH60_0;
	wire w_dff_A_MQIPxl8C9_0;
	wire w_dff_A_LNxAYDtE5_0;
	wire w_dff_A_JnVtZDyB7_0;
	wire w_dff_A_nlz9VTaX2_0;
	wire w_dff_A_APdtuPOw8_0;
	wire w_dff_A_f5o7qxak1_2;
	wire w_dff_A_8vuCgLM62_0;
	wire w_dff_A_Dscj6AP62_0;
	wire w_dff_A_lNCbob4Z0_0;
	wire w_dff_A_tztno8Af8_0;
	wire w_dff_A_AGXe5uzd6_0;
	wire w_dff_A_fGrWdj768_0;
	wire w_dff_A_VFoC8jf03_0;
	wire w_dff_A_bVp1TW5f3_2;
	wire w_dff_A_DI95F5hg9_0;
	wire w_dff_A_OrR0toCO2_0;
	wire w_dff_A_YVx5EXNo1_0;
	wire w_dff_A_fBBFJml14_0;
	wire w_dff_A_rhUCwuWP0_0;
	wire w_dff_A_j6SjAFiZ1_0;
	wire w_dff_A_SImkO0Rk1_0;
	wire w_dff_A_2vzslNSD5_2;
	wire w_dff_A_sI4UH3hQ0_0;
	wire w_dff_A_SwaiIOem2_0;
	wire w_dff_A_VP0tGqfs2_0;
	wire w_dff_A_KA9w5xpi9_0;
	wire w_dff_A_BxGNppwU5_0;
	wire w_dff_A_4nlB5erg5_0;
	wire w_dff_A_y5BuBXWP1_0;
	wire w_dff_A_UFllNdkx6_2;
	wire w_dff_A_ghEs7qxg9_0;
	wire w_dff_A_7HEJrJgE8_0;
	wire w_dff_A_cUoP0DwX9_0;
	wire w_dff_A_lKrS4BBf5_0;
	wire w_dff_A_00VubZMV4_0;
	wire w_dff_A_cB17GowC3_0;
	wire w_dff_A_Bsw4eSI67_2;
	wire w_dff_A_iD9eMV6H3_0;
	wire w_dff_A_YooGIYis9_0;
	wire w_dff_A_Edk6p6ct2_0;
	wire w_dff_A_lDy7wSU71_0;
	wire w_dff_A_sEFpQIxZ1_0;
	wire w_dff_A_KT6DvG4N0_0;
	wire w_dff_A_T53P2MVF1_0;
	wire w_dff_A_l3LCzSx29_2;
	wire w_dff_A_6KJFuvAg5_0;
	wire w_dff_A_pGn8BuzS1_0;
	wire w_dff_A_W7ei9MpB7_0;
	wire w_dff_A_Gkdd7hlu2_0;
	wire w_dff_A_2nmwoshl0_0;
	wire w_dff_A_X3HwRawM5_0;
	wire w_dff_A_4htbBja82_0;
	wire w_dff_A_dFpioPX11_2;
	wire w_dff_A_jGdEnVPo9_0;
	wire w_dff_A_9vTYiUYL5_0;
	wire w_dff_A_pkzt4W3q0_0;
	wire w_dff_A_FH4fhV2K5_0;
	wire w_dff_A_RU9wFu5j4_0;
	wire w_dff_A_zd3tJsmm7_0;
	wire w_dff_A_5tpsoEHB4_0;
	wire w_dff_A_OOU44twI0_2;
	wire w_dff_A_QH3hzpep6_0;
	wire w_dff_A_BzPxYXdQ6_0;
	wire w_dff_A_dAi5970u2_0;
	wire w_dff_A_eMIknfsY4_0;
	wire w_dff_A_8jaJ9J2g5_0;
	wire w_dff_A_LkUdZLky5_0;
	wire w_dff_A_MQSqB57S8_0;
	wire w_dff_A_eEjNbT6i5_2;
	wire w_dff_A_9FGrK7kQ6_0;
	wire w_dff_A_JhBvAJBs9_0;
	wire w_dff_A_naPF2VXU4_0;
	wire w_dff_A_ocj3SyfO2_0;
	wire w_dff_A_M9RFyUEd8_0;
	wire w_dff_A_AVJuVzmJ7_0;
	wire w_dff_A_0mD1Bjnm5_0;
	wire w_dff_A_2RADLT291_2;
	wire w_dff_A_pXp8UqB39_2;
	wire w_dff_A_NOz3iSZT9_0;
	wire w_dff_A_yveDk3Uy2_2;
	wire w_dff_A_2BecV9tE0_0;
	wire w_dff_A_o6nunRDk6_2;
	jnot g000(.din(w_G902_3[2]),.dout(n58),.clk(gclk));
	jnot g001(.din(w_G221_0[1]),.dout(n59),.clk(gclk));
	jnot g002(.din(w_G234_1[1]),.dout(n60),.clk(gclk));
	jor g003(.dina(w_G953_2[1]),.dinb(n60),.dout(n61),.clk(gclk));
	jor g004(.dina(n61),.dinb(w_dff_B_lRv8V3uU9_1),.dout(n62),.clk(gclk));
	jnot g005(.din(w_G110_0[2]),.dout(n63),.clk(gclk));
	jxor g006(.dina(w_G119_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_dff_B_j1EcKPlT8_0),.dinb(n62),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n66),.clk(gclk));
	jxor g009(.dina(w_n66_0[1]),.dinb(w_G146_0[2]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_G137_0[2]),.dinb(w_G128_0[2]),.dout(n68),.clk(gclk));
	jxor g011(.dina(w_dff_B_Riq3223L9_0),.dinb(w_n67_0[1]),.dout(n69),.clk(gclk));
	jxor g012(.dina(w_dff_B_rSPAN7jr8_0),.dinb(n65),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_0[1]),.dinb(w_n58_2[2]),.dout(n71),.clk(gclk));
	jand g014(.dina(w_n58_2[1]),.dinb(w_G234_1[0]),.dout(n72),.clk(gclk));
	jnot g015(.din(n72),.dout(n73),.clk(gclk));
	jand g016(.dina(w_n73_0[1]),.dinb(w_G217_0[2]),.dout(n74),.clk(gclk));
	jnot g017(.din(w_n74_0[1]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_dff_B_zfUoBTQh6_0),.dinb(w_n71_0[1]),.dout(n76),.clk(gclk));
	jxor g019(.dina(w_G143_0[2]),.dinb(w_G128_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_n77_0[1]),.dinb(w_G146_0[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(w_G137_0[1]),.dinb(w_G134_0[2]),.dout(n79),.clk(gclk));
	jxor g022(.dina(n79),.dinb(w_G131_0[2]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[2]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(n82),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_2[0]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[1]),.dinb(w_n58_2[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(w_n91_0[1]),.dinb(w_G472_0[2]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[1]),.dinb(w_n76_1[2]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[1]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_1[1]),.dout(n96),.clk(gclk));
	jnot g039(.din(w_G101_0[1]),.dout(n97),.clk(gclk));
	jxor g040(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n98),.clk(gclk));
	jxor g041(.dina(n98),.dinb(n97),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_n99_0[1]),.dinb(w_n84_0[0]),.dout(n100),.clk(gclk));
	jxor g043(.dina(w_G122_1[1]),.dinb(w_G110_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_dff_B_C21Cr2AB5_0),.dinb(n100),.dout(n102),.clk(gclk));
	jnot g045(.din(w_G953_1[2]),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n103_3[2]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n78_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_dEj9vy825_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n102_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[1]),.dinb(w_n58_1[2]),.dout(n108),.clk(gclk));
	jand g051(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n109),.clk(gclk));
	jxor g052(.dina(w_n109_0[1]),.dinb(w_n108_0[1]),.dout(n110),.clk(gclk));
	jand g053(.dina(w_n110_0[1]),.dinb(w_n96_0[2]),.dout(n111),.clk(gclk));
	jand g054(.dina(w_n73_0[0]),.dinb(w_G221_0[0]),.dout(n112),.clk(gclk));
	jnot g055(.din(w_n112_1[1]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n103_3[1]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(w_G140_0[1]),.dinb(w_n63_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n99_0[0]),.dout(n117),.clk(gclk));
	jxor g060(.dina(n117),.dinb(w_n81_0[1]),.dout(n118),.clk(gclk));
	jand g061(.dina(w_n118_0[1]),.dinb(w_n58_1[1]),.dout(n119),.clk(gclk));
	jxor g062(.dina(w_n119_0[1]),.dinb(w_G469_0[2]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n113_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_0[1]),.dinb(w_n111_0[1]),.dout(n122),.clk(gclk));
	jor g065(.dina(w_n103_3[0]),.dinb(w_G898_0[1]),.dout(n123),.clk(gclk));
	jnot g066(.din(n123),.dout(n124),.clk(gclk));
	jand g067(.dina(w_G237_0[0]),.dinb(w_G234_0[2]),.dout(n125),.clk(gclk));
	jnot g068(.din(n125),.dout(n126),.clk(gclk));
	jand g069(.dina(w_n126_0[1]),.dinb(w_G902_3[0]),.dout(n127),.clk(gclk));
	jand g070(.dina(w_n127_0[1]),.dinb(w_n124_0[1]),.dout(n128),.clk(gclk));
	jand g071(.dina(w_n126_0[0]),.dinb(w_G952_0[2]),.dout(n129),.clk(gclk));
	jand g072(.dina(n129),.dinb(w_n103_2[2]),.dout(n130),.clk(gclk));
	jor g073(.dina(w_n130_1[1]),.dinb(n128),.dout(n131),.clk(gclk));
	jnot g074(.din(w_G478_0[2]),.dout(n132),.clk(gclk));
	jxor g075(.dina(w_n77_0[0]),.dinb(w_G134_0[1]),.dout(n133),.clk(gclk));
	jand g076(.dina(w_n103_2[1]),.dinb(w_G234_0[1]),.dout(n134),.clk(gclk));
	jand g077(.dina(n134),.dinb(w_G217_0[1]),.dout(n135),.clk(gclk));
	jxor g078(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n136),.clk(gclk));
	jxor g079(.dina(n136),.dinb(w_G107_0[1]),.dout(n137),.clk(gclk));
	jxor g080(.dina(w_dff_B_idvopbrR7_0),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_dff_B_UKEKbcmb4_1),.dout(n139),.clk(gclk));
	jand g082(.dina(w_n139_0[1]),.dinb(w_n58_1[0]),.dout(n140),.clk(gclk));
	jxor g083(.dina(w_n140_0[1]),.dinb(w_dff_B_Lhkdwcf79_1),.dout(n141),.clk(gclk));
	jnot g084(.din(w_G475_0[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_G122_0[2]),.dinb(w_G113_0[1]),.dout(n143),.clk(gclk));
	jxor g086(.dina(n143),.dinb(w_G104_0[1]),.dout(n144),.clk(gclk));
	jnot g087(.din(w_G214_0[0]),.dout(n145),.clk(gclk));
	jor g088(.dina(w_n86_0[0]),.dinb(n145),.dout(n146),.clk(gclk));
	jnot g089(.din(w_G131_0[1]),.dout(n147),.clk(gclk));
	jxor g090(.dina(w_G143_0[1]),.dinb(n147),.dout(n148),.clk(gclk));
	jxor g091(.dina(n148),.dinb(n146),.dout(n149),.clk(gclk));
	jxor g092(.dina(n149),.dinb(w_n67_0[0]),.dout(n150),.clk(gclk));
	jxor g093(.dina(n150),.dinb(w_dff_B_OR4AFcGl9_1),.dout(n151),.clk(gclk));
	jand g094(.dina(w_n151_0[2]),.dinb(w_n58_0[2]),.dout(n152),.clk(gclk));
	jxor g095(.dina(w_n152_0[1]),.dinb(w_dff_B_gbbLE1r79_1),.dout(n153),.clk(gclk));
	jand g096(.dina(w_n153_1[1]),.dinb(w_n141_1[1]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n131_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[1]),.dinb(w_n122_1[1]),.dout(n156),.clk(gclk));
	jand g099(.dina(w_n156_0[1]),.dinb(w_n93_1[1]),.dout(n157),.clk(gclk));
	jxor g100(.dina(w_n157_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_1HIeDp7r2_2),.clk(gclk));
	jnot g101(.din(w_G472_0[1]),.dout(n159),.clk(gclk));
	jxor g102(.dina(w_n91_0[0]),.dinb(w_dff_B_fW3ODDb64_1),.dout(n160),.clk(gclk));
	jand g103(.dina(w_n160_1[2]),.dinb(w_n76_1[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_1[1]),.dinb(w_n122_1[0]),.dout(n162),.clk(gclk));
	jxor g105(.dina(w_n152_0[0]),.dinb(w_G475_0[1]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_1[1]),.dinb(w_n141_1[0]),.dout(n164),.clk(gclk));
	jand g107(.dina(w_n164_0[1]),.dinb(w_n131_1[1]),.dout(n165),.clk(gclk));
	jand g108(.dina(w_n165_0[2]),.dinb(w_n162_0[1]),.dout(n166),.clk(gclk));
	jxor g109(.dina(w_n166_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_jzkZ6mNp7_2),.clk(gclk));
	jxor g110(.dina(w_n140_0[0]),.dinb(w_G478_0[1]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n153_1[0]),.dinb(w_n168_1[1]),.dout(n169),.clk(gclk));
	jand g112(.dina(w_n169_0[1]),.dinb(w_n131_1[0]),.dout(n170),.clk(gclk));
	jand g113(.dina(w_n170_0[1]),.dinb(w_n162_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n171_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_25G69Rjr9_2),.clk(gclk));
	jxor g115(.dina(w_n74_0[0]),.dinb(w_n71_0[0]),.dout(n173),.clk(gclk));
	jand g116(.dina(w_n160_1[1]),.dinb(w_n173_1[1]),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n174_0[1]),.dinb(w_n156_0[0]),.dout(n175),.clk(gclk));
	jxor g118(.dina(w_n175_0[1]),.dinb(w_G110_0[0]),.dout(w_dff_A_z3wcJUFY4_2),.clk(gclk));
	jand g119(.dina(w_n92_1[0]),.dinb(w_n173_1[0]),.dout(n177),.clk(gclk));
	jand g120(.dina(w_n177_0[2]),.dinb(w_n122_0[2]),.dout(n178),.clk(gclk));
	jor g121(.dina(w_n103_2[0]),.dinb(w_G900_0[1]),.dout(n179),.clk(gclk));
	jnot g122(.din(n179),.dout(n180),.clk(gclk));
	jand g123(.dina(w_n180_0[1]),.dinb(w_n127_0[0]),.dout(n181),.clk(gclk));
	jor g124(.dina(n181),.dinb(w_n130_1[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(w_n182_1[2]),.dinb(w_n169_0[0]),.dout(n183),.clk(gclk));
	jand g126(.dina(w_n183_0[2]),.dinb(w_n178_0[1]),.dout(n184),.clk(gclk));
	jxor g127(.dina(w_n184_0[1]),.dinb(w_G128_0[0]),.dout(w_dff_A_WlpV7S0I3_2),.clk(gclk));
	jand g128(.dina(w_n163_1[0]),.dinb(w_n168_1[0]),.dout(n186),.clk(gclk));
	jand g129(.dina(w_n186_0[1]),.dinb(w_n93_1[0]),.dout(n187),.clk(gclk));
	jand g130(.dina(n187),.dinb(w_n182_1[1]),.dout(n188),.clk(gclk));
	jand g131(.dina(n188),.dinb(w_n122_0[1]),.dout(n189),.clk(gclk));
	jxor g132(.dina(w_n189_0[1]),.dinb(w_G143_0[0]),.dout(w_dff_A_WaS3U3aF1_2),.clk(gclk));
	jand g133(.dina(w_n182_1[0]),.dinb(w_n164_0[0]),.dout(n191),.clk(gclk));
	jand g134(.dina(w_n191_0[2]),.dinb(w_n178_0[0]),.dout(n192),.clk(gclk));
	jxor g135(.dina(w_n192_0[2]),.dinb(w_G146_0[0]),.dout(w_dff_A_kpZMc0eW0_2),.clk(gclk));
	jnot g136(.din(w_G469_0[1]),.dout(n194),.clk(gclk));
	jxor g137(.dina(w_n119_0[0]),.dinb(w_dff_B_3kB9E9WJ2_1),.dout(n195),.clk(gclk));
	jand g138(.dina(w_n195_0[2]),.dinb(w_n113_0[1]),.dout(n196),.clk(gclk));
	jand g139(.dina(n196),.dinb(w_n111_0[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n93_0[2]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_0[1]),.dinb(w_n165_0[1]),.dout(n199),.clk(gclk));
	jxor g142(.dina(w_n199_0[2]),.dinb(w_G113_0[0]),.dout(w_dff_A_f5o7qxak1_2),.clk(gclk));
	jand g143(.dina(w_n198_0[0]),.dinb(w_n170_0[0]),.dout(n201),.clk(gclk));
	jxor g144(.dina(w_n201_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_bVp1TW5f3_2),.clk(gclk));
	jand g145(.dina(w_n177_0[1]),.dinb(w_n155_0[0]),.dout(n203),.clk(gclk));
	jand g146(.dina(n203),.dinb(w_n197_1[0]),.dout(n204),.clk(gclk));
	jxor g147(.dina(w_n204_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_2vzslNSD5_2),.clk(gclk));
	jand g148(.dina(w_n197_0[2]),.dinb(w_n161_1[0]),.dout(n206),.clk(gclk));
	jand g149(.dina(w_n206_0[1]),.dinb(w_n131_0[2]),.dout(n207),.clk(gclk));
	jand g150(.dina(n207),.dinb(w_n186_0[0]),.dout(n208),.clk(gclk));
	jxor g151(.dina(w_n208_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_UFllNdkx6_2),.clk(gclk));
	jand g152(.dina(w_n191_0[1]),.dinb(w_n174_0[0]),.dout(n210),.clk(gclk));
	jand g153(.dina(w_n210_0[1]),.dinb(w_n197_0[1]),.dout(n211),.clk(gclk));
	jxor g154(.dina(w_n211_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_Bsw4eSI67_2),.clk(gclk));
	jnot g155(.din(w_n109_0[0]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_dff_B_twwOpmxt5_0),.dinb(w_n108_0[0]),.dout(n214),.clk(gclk));
	jand g157(.dina(w_n214_0[2]),.dinb(w_n96_0[1]),.dout(n215),.clk(gclk));
	jand g158(.dina(n215),.dinb(w_n121_0[0]),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_1[1]),.dinb(w_n93_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[1]),.dinb(w_n191_0[0]),.dout(n218),.clk(gclk));
	jxor g161(.dina(w_n218_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_l3LCzSx29_2),.clk(gclk));
	jand g162(.dina(w_n217_0[0]),.dinb(w_n183_0[1]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_dFpioPX11_2),.clk(gclk));
	jand g164(.dina(w_n177_0[0]),.dinb(w_n154_1[0]),.dout(n222),.clk(gclk));
	jand g165(.dina(n222),.dinb(w_n182_0[2]),.dout(n223),.clk(gclk));
	jand g166(.dina(n223),.dinb(w_n216_1[0]),.dout(n224),.clk(gclk));
	jxor g167(.dina(w_n224_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_OOU44twI0_2),.clk(gclk));
	jand g168(.dina(w_n216_0[2]),.dinb(w_n210_0[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_eEjNbT6i5_2),.clk(gclk));
	jor g170(.dina(w_n171_0[0]),.dinb(w_n157_0[0]),.dout(n228),.clk(gclk));
	jor g171(.dina(n228),.dinb(w_n166_0[0]),.dout(n229),.clk(gclk));
	jor g172(.dina(n229),.dinb(w_n208_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n204_0[0]),.dinb(w_n201_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(w_n175_0[0]),.dout(n232),.clk(gclk));
	jor g175(.dina(n232),.dinb(w_n199_0[1]),.dout(n233),.clk(gclk));
	jor g176(.dina(n233),.dinb(n230),.dout(n234),.clk(gclk));
	jor g177(.dina(w_n226_0[0]),.dinb(w_n224_0[0]),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(w_n192_0[1]),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n218_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n211_0[0]),.dinb(w_n189_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(w_n184_0[0]),.dout(n239),.clk(gclk));
	jor g182(.dina(n239),.dinb(w_dff_B_JXxE9l7T2_1),.dout(n240),.clk(gclk));
	jor g183(.dina(n240),.dinb(w_dff_B_2X3F5Utf0_1),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n234),.dout(n242),.clk(gclk));
	jand g185(.dina(w_n195_0[1]),.dinb(w_n214_0[1]),.dout(n243),.clk(gclk));
	jxor g186(.dina(w_n112_1[0]),.dinb(w_n95_1[0]),.dout(n244),.clk(gclk));
	jand g187(.dina(w_dff_B_apkQf78x5_0),.dinb(w_n243_0[1]),.dout(n245),.clk(gclk));
	jor g188(.dina(n245),.dinb(w_n216_0[1]),.dout(n246),.clk(gclk));
	jand g189(.dina(n246),.dinb(w_n161_0[2]),.dout(n247),.clk(gclk));
	jand g190(.dina(w_n113_0[0]),.dinb(w_n96_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_289zX16p1_0),.dinb(w_n243_0[0]),.dout(n249),.clk(gclk));
	jxor g192(.dina(w_n160_1[0]),.dinb(w_n76_1[0]),.dout(n250),.clk(gclk));
	jand g193(.dina(w_dff_B_EOM0QiK69_0),.dinb(w_n249_0[1]),.dout(n251),.clk(gclk));
	jor g194(.dina(n251),.dinb(w_n206_0[0]),.dout(n252),.clk(gclk));
	jor g195(.dina(n252),.dinb(n247),.dout(n253),.clk(gclk));
	jand g196(.dina(n253),.dinb(w_n154_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(n254),.dinb(w_n130_0[2]),.dout(n255),.clk(gclk));
	jor g198(.dina(w_dff_B_Wmu07nX56_0),.dinb(w_n242_2[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_G952_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(w_n153_0[2]),.dinb(w_n141_0[2]),.dout(n258),.clk(gclk));
	jor g201(.dina(w_n154_0[1]),.dinb(w_n130_0[1]),.dout(n259),.clk(gclk));
	jand g202(.dina(n259),.dinb(w_n258_0[2]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n161_0[1]),.dout(n261),.clk(gclk));
	jand g204(.dina(n261),.dinb(w_n249_0[0]),.dout(n262),.clk(gclk));
	jor g205(.dina(n262),.dinb(w_G953_1[1]),.dout(n263),.clk(gclk));
	jor g206(.dina(w_dff_B_xdFdkSUS6_0),.dinb(n257),.dout(w_dff_A_2RADLT291_2),.clk(gclk));
	jor g207(.dina(w_n103_1[2]),.dinb(w_G952_0[0]),.dout(n265),.clk(gclk));
	jand g208(.dina(w_n242_2[1]),.dinb(w_G210_0[0]),.dout(n266),.clk(gclk));
	jand g209(.dina(n266),.dinb(w_G902_2[2]),.dout(n267),.clk(gclk));
	jxor g210(.dina(n267),.dinb(w_n107_0[0]),.dout(n268),.clk(gclk));
	jand g211(.dina(n268),.dinb(w_n265_2[1]),.dout(G51),.clk(gclk));
	jand g212(.dina(w_n242_2[0]),.dinb(w_G469_0[0]),.dout(n270),.clk(gclk));
	jand g213(.dina(n270),.dinb(w_G902_2[1]),.dout(n271),.clk(gclk));
	jxor g214(.dina(n271),.dinb(w_n118_0[0]),.dout(n272),.clk(gclk));
	jand g215(.dina(n272),.dinb(w_n265_2[0]),.dout(G54),.clk(gclk));
	jand g216(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n274),.clk(gclk));
	jand g217(.dina(w_n274_0[1]),.dinb(w_n242_1[2]),.dout(n275),.clk(gclk));
	jor g218(.dina(n275),.dinb(w_n151_0[1]),.dout(n276),.clk(gclk));
	jnot g219(.din(w_n151_0[0]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n131_0[1]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n92_0[2]),.dinb(w_n173_0[2]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n214_0[0]),.dinb(w_n95_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n120_0[0]),.dinb(w_n112_0[2]),.dout(n281),.clk(gclk));
	jor g224(.dina(n281),.dinb(w_n280_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_1[1]),.dinb(w_n279_0[1]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n278_0[2]),.dout(n284),.clk(gclk));
	jor g227(.dina(n284),.dinb(w_n258_0[1]),.dout(n285),.clk(gclk));
	jor g228(.dina(w_n195_0[0]),.dinb(w_n112_0[1]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n280_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n279_0[0]),.dinb(w_n287_1[1]),.dout(n288),.clk(gclk));
	jnot g231(.din(w_n165_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(n289),.dinb(w_n288_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n160_0[2]),.dinb(w_n173_0[1]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n163_0[2]),.dinb(w_n168_0[2]),.dout(n292),.clk(gclk));
	jor g235(.dina(w_n292_0[1]),.dinb(w_n278_0[1]),.dout(n293),.clk(gclk));
	jor g236(.dina(w_n293_0[1]),.dinb(w_n287_1[0]),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n294_0[1]),.dinb(w_n291_1[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n163_0[1]),.dinb(w_n141_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(n296),.dinb(w_n278_0[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(w_n297_0[1]),.dinb(w_n288_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n295),.dout(n299),.clk(gclk));
	jand g242(.dina(n299),.dinb(w_dff_B_50NgK2HR5_1),.dout(n300),.clk(gclk));
	jand g243(.dina(n300),.dinb(w_dff_B_mg6vrPOX5_1),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n199_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n92_0[1]),.dinb(w_n76_0[2]),.dout(n303),.clk(gclk));
	jor g246(.dina(w_n303_0[1]),.dinb(w_n294_0[0]),.dout(n304),.clk(gclk));
	jor g247(.dina(w_n282_1[0]),.dinb(w_n291_1[0]),.dout(n305),.clk(gclk));
	jor g248(.dina(n305),.dinb(w_n297_0[0]),.dout(n306),.clk(gclk));
	jor g249(.dina(w_n160_0[1]),.dinb(w_n76_0[1]),.dout(n307),.clk(gclk));
	jor g250(.dina(w_n307_0[2]),.dinb(w_n293_0[0]),.dout(n308),.clk(gclk));
	jor g251(.dina(n308),.dinb(w_n282_0[2]),.dout(n309),.clk(gclk));
	jand g252(.dina(n309),.dinb(n306),.dout(n310),.clk(gclk));
	jand g253(.dina(n310),.dinb(w_dff_B_0LxZ9BDq7_1),.dout(n311),.clk(gclk));
	jand g254(.dina(n311),.dinb(w_dff_B_YKHt5J0m8_1),.dout(n312),.clk(gclk));
	jand g255(.dina(n312),.dinb(n301),.dout(n313),.clk(gclk));
	jnot g256(.din(w_n192_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n110_0[0]),.dinb(w_n95_0[1]),.dout(n315),.clk(gclk));
	jor g258(.dina(n315),.dinb(w_n286_0[0]),.dout(n316),.clk(gclk));
	jnot g259(.din(w_n182_0[1]),.dout(n317),.clk(gclk));
	jor g260(.dina(w_n307_0[1]),.dinb(w_n292_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(n318),.dinb(w_n317_0[2]),.dout(n319),.clk(gclk));
	jor g262(.dina(n319),.dinb(w_n316_0[2]),.dout(n320),.clk(gclk));
	jor g263(.dina(w_n153_0[1]),.dinb(w_n168_0[1]),.dout(n321),.clk(gclk));
	jor g264(.dina(w_n317_0[1]),.dinb(n321),.dout(n322),.clk(gclk));
	jor g265(.dina(w_n322_0[1]),.dinb(w_n303_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(w_n316_0[1]),.dinb(w_n323_0[1]),.dout(n324),.clk(gclk));
	jand g267(.dina(n324),.dinb(n320),.dout(n325),.clk(gclk));
	jand g268(.dina(n325),.dinb(n314),.dout(n326),.clk(gclk));
	jor g269(.dina(w_n316_0[0]),.dinb(w_n291_0[2]),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n327_0[1]),.dinb(w_n322_0[0]),.dout(n328),.clk(gclk));
	jnot g271(.din(w_n183_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(w_n327_0[0]),.dinb(w_n329_0[1]),.dout(n330),.clk(gclk));
	jand g273(.dina(n330),.dinb(n328),.dout(n331),.clk(gclk));
	jor g274(.dina(w_n307_0[0]),.dinb(w_n287_0[2]),.dout(n332),.clk(gclk));
	jor g275(.dina(w_n329_0[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jor g276(.dina(w_n258_0[0]),.dinb(w_n291_0[1]),.dout(n334),.clk(gclk));
	jor g277(.dina(n334),.dinb(w_n317_0[0]),.dout(n335),.clk(gclk));
	jor g278(.dina(n335),.dinb(w_n287_0[1]),.dout(n336),.clk(gclk));
	jor g279(.dina(w_n323_0[0]),.dinb(w_n282_0[1]),.dout(n337),.clk(gclk));
	jand g280(.dina(n337),.dinb(n336),.dout(n338),.clk(gclk));
	jand g281(.dina(n338),.dinb(w_dff_B_L52U40XV7_1),.dout(n339),.clk(gclk));
	jand g282(.dina(n339),.dinb(w_dff_B_ARLySCip4_1),.dout(n340),.clk(gclk));
	jand g283(.dina(n340),.dinb(w_dff_B_WoMQU8Xr6_1),.dout(n341),.clk(gclk));
	jand g284(.dina(w_n341_0[1]),.dinb(w_n313_0[1]),.dout(n342),.clk(gclk));
	jnot g285(.din(w_n274_0[0]),.dout(n343),.clk(gclk));
	jor g286(.dina(w_dff_B_dZJonO2V5_0),.dinb(n342),.dout(n344),.clk(gclk));
	jor g287(.dina(n344),.dinb(w_dff_B_5lrRqkCa5_1),.dout(n345),.clk(gclk));
	jand g288(.dina(n345),.dinb(w_n265_1[2]),.dout(n346),.clk(gclk));
	jand g289(.dina(n346),.dinb(w_dff_B_8bptot6U4_1),.dout(G60),.clk(gclk));
	jand g290(.dina(w_n242_1[1]),.dinb(w_G478_0[0]),.dout(n348),.clk(gclk));
	jand g291(.dina(n348),.dinb(w_G902_1[2]),.dout(n349),.clk(gclk));
	jxor g292(.dina(n349),.dinb(w_n139_0[0]),.dout(n350),.clk(gclk));
	jand g293(.dina(n350),.dinb(w_n265_1[1]),.dout(G63),.clk(gclk));
	jand g294(.dina(w_n242_1[0]),.dinb(w_G217_0[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_G902_1[1]),.dout(n353),.clk(gclk));
	jxor g296(.dina(n353),.dinb(w_n70_0[0]),.dout(n354),.clk(gclk));
	jand g297(.dina(n354),.dinb(w_n265_1[0]),.dout(G66),.clk(gclk));
	jor g298(.dina(w_n124_0[0]),.dinb(w_n102_0[0]),.dout(n356),.clk(gclk));
	jor g299(.dina(w_n313_0[0]),.dinb(w_G953_1[0]),.dout(n357),.clk(gclk));
	jand g300(.dina(w_G898_0[0]),.dinb(w_G224_0[0]),.dout(n358),.clk(gclk));
	jor g301(.dina(n358),.dinb(w_n103_1[1]),.dout(n359),.clk(gclk));
	jand g302(.dina(w_dff_B_CIDRaylk5_0),.dinb(n357),.dout(n360),.clk(gclk));
	jxor g303(.dina(n360),.dinb(w_dff_B_BJrzF2mA7_1),.dout(w_dff_A_pXp8UqB39_2),.clk(gclk));
	jor g304(.dina(w_n341_0[0]),.dinb(w_G953_0[2]),.dout(n362),.clk(gclk));
	jand g305(.dina(w_G900_0[0]),.dinb(w_G227_0[0]),.dout(n363),.clk(gclk));
	jor g306(.dina(n363),.dinb(w_n103_1[0]),.dout(n364),.clk(gclk));
	jand g307(.dina(w_dff_B_XytGs9et4_0),.dinb(n362),.dout(n365),.clk(gclk));
	jxor g308(.dina(w_n81_0[0]),.dinb(w_n66_0[0]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(w_n180_0[0]),.dout(n367),.clk(gclk));
	jxor g310(.dina(w_dff_B_7zCrDNGV5_0),.dinb(n365),.dout(w_dff_A_yveDk3Uy2_2),.clk(gclk));
	jand g311(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(w_dff_B_rRqdFC7O3_0),.dinb(w_n242_0[2]),.dout(n370),.clk(gclk));
	jxor g313(.dina(n370),.dinb(w_n90_0[0]),.dout(n371),.clk(gclk));
	jand g314(.dina(n371),.dinb(w_n265_0[2]),.dout(w_dff_A_o6nunRDk6_2),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_e09HX4jy3_0),.doutb(w_G101_0[1]),.doutc(w_dff_A_hek1xz6t0_2),.din(G101));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_XBXSzFWV5_0),.doutb(w_dff_A_mfxrm3Sh9_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_tILj3M467_0),.doutb(w_dff_A_TWcZ3hlV8_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_dff_A_iU37nXPr2_0),.doutb(w_G110_0[1]),.doutc(w_G110_0[2]),.din(G110));
	jspl3 jspl3_w_G113_0(.douta(w_dff_A_W6A9ZwZM7_0),.doutb(w_G113_0[1]),.doutc(w_G113_0[2]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_hpithpsj5_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_8ccLeRGo3_0),.doutb(w_G119_0[1]),.doutc(w_dff_A_pltr9Sy91_2),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_zeEAMW488_1),.doutc(w_G122_0[2]),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_G122_1[1]),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_C8994UPm7_0),.doutb(w_dff_A_WndBmvHt3_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_julECBpF0_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl3 jspl3_w_G131_0(.douta(w_dff_A_kods908k3_0),.doutb(w_G131_0[1]),.doutc(w_dff_A_yHCBM2o71_2),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_6fVrQNeK2_0),.doutb(w_dff_A_Ceh9Y6RA4_1),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_dmY5xswP2_0),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_SXTVyYmQ3_0),.doutb(w_dff_A_wF4hsBQF2_1),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_dff_A_54YWHNz46_0),.doutb(w_dff_A_8zc6us4R5_1),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_lGqwmx6k0_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(w_dff_B_pJ00iYd30_3));
	jspl3 jspl3_w_G210_0(.douta(w_dff_A_OxcboRLa7_0),.doutb(w_dff_A_lgVNsBUw3_1),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_dff_A_MndoQkpc4_1),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_dff_A_YFHk7fnc7_0),.doutb(w_G217_0[1]),.doutc(w_dff_A_Ej80MD9W3_2),.din(w_dff_B_NMvSU6qi8_3));
	jspl jspl_w_G221_0(.douta(w_dff_A_ramVYyqn5_0),.doutb(w_G221_0[1]),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_dff_A_kSftgAv93_1),.din(G224));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_dff_A_7WMoCQIU0_1),.din(G227));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_e1THIr3i3_1),.doutc(w_G234_0[2]),.din(G234));
	jspl jspl_w_G234_1(.douta(w_dff_A_CqMkEHCF9_0),.doutb(w_G234_1[1]),.din(w_G234_0[0]));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_dff_A_hi8HOVFL6_0),.doutb(w_G469_0[1]),.doutc(w_dff_A_yjGMR8qv0_2),.din(G469));
	jspl3 jspl3_w_G472_0(.douta(w_G472_0[0]),.doutb(w_G472_0[1]),.doutc(w_dff_A_lLBd2Mlm2_2),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_YB1Nc0QZ0_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_dff_A_fKDY7Nsc9_0),.doutb(w_dff_A_l0eGAroD5_1),.doutc(w_G478_0[2]),.din(G478));
	jspl jspl_w_G898_0(.douta(w_G898_0[0]),.doutb(w_dff_A_0sMTgjXs1_1),.din(G898));
	jspl jspl_w_G900_0(.douta(w_G900_0[0]),.doutb(w_dff_A_j1v6xOuW7_1),.din(G900));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_dff_A_Y0O5LEFn9_1),.doutc(w_dff_A_pWNy4AKp6_2),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_dff_A_qxF7e5cA0_1),.doutc(w_dff_A_eA2euOQv1_2),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_dff_A_tiODlU1F4_0),.doutb(w_G902_3[1]),.doutc(w_G902_3[2]),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_GJtCJ9al0_1),.doutc(w_dff_A_SjzwPv5X2_2),.din(w_dff_B_PjuaBNu04_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_G953_0[1]),.doutc(w_dff_A_hiFdIg9Q8_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_KXfeyVnS8_0),.doutb(w_dff_A_UGqxG0g45_1),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_G953_2(.douta(w_G953_2[0]),.doutb(w_dff_A_4gro4Qq16_1),.din(w_G953_0[1]));
	jspl3 jspl3_w_n58_0(.douta(w_dff_A_N1JBoeja7_0),.doutb(w_n58_0[1]),.doutc(w_dff_A_mcU4tgIv0_2),.din(n58));
	jspl3 jspl3_w_n58_1(.douta(w_n58_1[0]),.doutb(w_n58_1[1]),.doutc(w_n58_1[2]),.din(w_n58_0[0]));
	jspl3 jspl3_w_n58_2(.douta(w_dff_A_vajKnaec8_0),.doutb(w_n58_2[1]),.doutc(w_dff_A_S5z7eyd04_2),.din(w_n58_0[1]));
	jspl jspl_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n66_0(.douta(w_dff_A_IzmLdrPM4_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_dff_A_O82f2qgK5_0),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n70_0(.douta(w_dff_A_HAwpuHLL6_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n74_0(.douta(w_dff_A_zvGreQTX8_0),.doutb(w_n74_0[1]),.din(n74));
	jspl3 jspl3_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.doutc(w_n76_0[2]),.din(n76));
	jspl3 jspl3_w_n76_1(.douta(w_n76_1[0]),.doutb(w_n76_1[1]),.doutc(w_n76_1[2]),.din(w_n76_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_dff_A_Sc72a3VD2_1),.doutc(w_dff_A_JDwHL18b8_2),.din(n81));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_0ikeNFih7_1),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_dff_A_j4eWW6fM7_0),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_dff_A_soEHyxz21_1),.doutc(w_dff_A_yMjaBLlH6_2),.din(n93));
	jspl jspl_w_n93_1(.douta(w_n93_1[0]),.doutb(w_dff_A_a9FOPwLV5_1),.din(w_n93_0[0]));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_dff_A_VVcpvPLv4_1),.doutc(w_dff_A_s4HEiENx9_2),.din(n95));
	jspl jspl_w_n95_1(.douta(w_dff_A_3xNgarSq0_0),.doutb(w_n95_1[1]),.din(w_n95_0[0]));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_HTLSczVE8_1),.doutc(w_dff_A_mPRuzlGc6_2),.din(w_dff_B_836m1ysa9_3));
	jspl jspl_w_n99_0(.douta(w_dff_A_jjWIrSHE2_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n103_1(.douta(w_n103_1[0]),.doutb(w_n103_1[1]),.doutc(w_n103_1[2]),.din(w_n103_0[0]));
	jspl3 jspl3_w_n103_2(.douta(w_n103_2[0]),.doutb(w_n103_2[1]),.doutc(w_dff_A_sCiPDOfo6_2),.din(w_n103_0[1]));
	jspl3 jspl3_w_n103_3(.douta(w_n103_3[0]),.doutb(w_n103_3[1]),.doutc(w_n103_3[2]),.din(w_n103_0[2]));
	jspl jspl_w_n107_0(.douta(w_dff_A_dOdQglT95_0),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_dff_A_2zVWGoBz7_1),.din(n109));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_dff_A_hj8rotjC3_1),.doutc(w_dff_A_23L3vLrA3_2),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_viYe8xIr3_1),.doutc(w_dff_A_bFIRqKpw9_2),.din(n113));
	jspl jspl_w_n118_0(.douta(w_dff_A_DCDL6rW75_0),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_KOS7OcBZ2_1),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl jspl_w_n124_0(.douta(w_dff_A_5djuqVFR4_0),.doutb(w_n124_0[1]),.din(n124));
	jspl jspl_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_2Owppcnm8_1),.doutc(w_dff_A_rcqTukSG5_2),.din(n130));
	jspl jspl_w_n130_1(.douta(w_n130_1[0]),.doutb(w_n130_1[1]),.din(w_n130_0[0]));
	jspl3 jspl3_w_n131_0(.douta(w_dff_A_Rkt191pb6_0),.doutb(w_n131_0[1]),.doutc(w_dff_A_66Ajoyz44_2),.din(n131));
	jspl3 jspl3_w_n131_1(.douta(w_n131_1[0]),.doutb(w_n131_1[1]),.doutc(w_n131_1[2]),.din(w_n131_0[0]));
	jspl jspl_w_n139_0(.douta(w_dff_A_KdXWk3gy3_0),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_5z0D4Avc7_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl jspl_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_dff_A_GAFQXiQk6_2),.din(n154));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.doutc(w_n160_0[2]),.din(n160));
	jspl3 jspl3_w_n160_1(.douta(w_n160_1[0]),.doutb(w_n160_1[1]),.doutc(w_n160_1[2]),.din(w_n160_0[0]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_dff_A_akdZEYzP7_1),.doutc(w_dff_A_LMQzXh8Y3_2),.din(w_dff_B_9df6Tjnu5_3));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_MX6iKdHZ7_1),.doutc(w_dff_A_EZQQlWfd2_2),.din(n165));
	jspl jspl_w_n166_0(.douta(w_dff_A_6gvA7Kvb2_0),.doutb(w_n166_0[1]),.din(n166));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl jspl_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.din(w_n168_0[0]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(w_dff_B_2T9zAfDd3_2));
	jspl jspl_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.din(n171));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.din(w_n173_0[0]));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_dff_A_dG3pUUhf3_1),.din(w_dff_B_TYA0jWKs3_2));
	jspl jspl_w_n175_0(.douta(w_dff_A_YxtIsUQ09_0),.doutb(w_n175_0[1]),.din(n175));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_dff_A_pL9aPxaf8_1),.doutc(w_dff_A_NybkuwfE7_2),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_dff_A_LuAz3Zoz4_0),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n182_0(.douta(w_dff_A_qupKCXvj3_0),.doutb(w_n182_0[1]),.doutc(w_dff_A_Kq7nAxjJ6_2),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_dff_A_Yxw5h3ar9_1),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n183_0(.douta(w_n183_0[0]),.doutb(w_dff_A_C9ZSpTRT0_1),.doutc(w_dff_A_DevZQJIz3_2),.din(n183));
	jspl jspl_w_n184_0(.douta(w_dff_A_xEIhDbgd1_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n186_0(.douta(w_dff_A_sB64z77S3_0),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n191_0(.douta(w_dff_A_iSuFEqde4_0),.doutb(w_n191_0[1]),.doutc(w_dff_A_AVw7lWSl2_2),.din(n191));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_dff_A_jo4ZeTVu3_1),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.doutc(w_n195_0[2]),.din(n195));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_dff_A_zhsHfnEm0_1),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_wHFsuuiJ8_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_dff_A_xQT8wLcD4_1),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n208_0(.douta(w_dff_A_FJ51mBDe1_0),.doutb(w_n208_0[1]),.din(n208));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.din(n211));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_dff_A_QKfCqza18_2),.din(n216));
	jspl jspl_w_n216_1(.douta(w_dff_A_LVBGMoP22_0),.doutb(w_n216_1[1]),.din(w_n216_0[0]));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n242_1(.douta(w_n242_1[0]),.doutb(w_n242_1[1]),.doutc(w_n242_1[2]),.din(w_n242_0[0]));
	jspl3 jspl3_w_n242_2(.douta(w_n242_2[0]),.doutb(w_n242_2[1]),.doutc(w_n242_2[2]),.din(w_n242_0[1]));
	jspl jspl_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n249_0(.douta(w_dff_A_qF97oLAq4_0),.doutb(w_n249_0[1]),.din(n249));
	jspl3 jspl3_w_n258_0(.douta(w_n258_0[0]),.doutb(w_dff_A_jRuMaBaC7_1),.doutc(w_dff_A_lWXx1Z5k6_2),.din(n258));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_dff_A_H8dpCByK6_1),.doutc(w_n265_0[2]),.din(w_dff_B_YCfBBzZ70_3));
	jspl3 jspl3_w_n265_1(.douta(w_dff_A_5FhJvPGZ3_0),.doutb(w_dff_A_2LxxnF2Y5_1),.doutc(w_n265_1[2]),.din(w_n265_0[0]));
	jspl jspl_w_n265_2(.douta(w_n265_2[0]),.doutb(w_n265_2[1]),.din(w_n265_0[1]));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_p6LfYgvw2_1),.din(n274));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_dff_A_mDT284LI8_2),.din(w_dff_B_UvX1D9mq7_3));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_d1LbOOHB1_2));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_dff_A_92hYar444_1),.doutc(w_dff_A_5ld2p0Q47_2),.din(n282));
	jspl jspl_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.din(w_n282_0[0]));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(n286));
	jspl3 jspl3_w_n287_0(.douta(w_n287_0[0]),.doutb(w_dff_A_GlRQ3DSW3_1),.doutc(w_n287_0[2]),.din(n287));
	jspl jspl_w_n287_1(.douta(w_n287_1[0]),.doutb(w_n287_1[1]),.din(w_n287_0[0]));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl3 jspl3_w_n291_0(.douta(w_dff_A_e4tCZxkY8_0),.doutb(w_n291_0[1]),.doutc(w_dff_A_cgR5SqR31_2),.din(n291));
	jspl jspl_w_n291_1(.douta(w_n291_1[0]),.doutb(w_dff_A_N5usaIeo9_1),.din(w_n291_0[0]));
	jspl jspl_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.din(n292));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.din(n294));
	jspl jspl_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.din(w_dff_B_sMOGxZUK7_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_IKnNahbU2_1),.din(w_dff_B_mZMqktea3_2));
	jspl3 jspl3_w_n307_0(.douta(w_dff_A_t0AN5XoL1_0),.doutb(w_n307_0[1]),.doutc(w_dff_A_b8HLrhFj1_2),.din(n307));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n316_0(.douta(w_n316_0[0]),.doutb(w_dff_A_WRKgB4gP3_1),.doutc(w_dff_A_DGIu3rtn2_2),.din(n316));
	jspl3 jspl3_w_n317_0(.douta(w_dff_A_nT7IT46z9_0),.doutb(w_n317_0[1]),.doutc(w_dff_A_474pC7iS8_2),.din(w_dff_B_l6WeeIPA1_3));
	jspl jspl_w_n322_0(.douta(w_dff_A_ESH28Yld7_0),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n341_0(.douta(w_n341_0[0]),.doutb(w_n341_0[1]),.din(n341));
	jdff dff_B_gRoE5hj54_0(.din(n263),.dout(w_dff_B_gRoE5hj54_0),.clk(gclk));
	jdff dff_B_217tmLfb0_0(.din(w_dff_B_gRoE5hj54_0),.dout(w_dff_B_217tmLfb0_0),.clk(gclk));
	jdff dff_B_oHQ6x86A1_0(.din(w_dff_B_217tmLfb0_0),.dout(w_dff_B_oHQ6x86A1_0),.clk(gclk));
	jdff dff_B_4hfbee0s3_0(.din(w_dff_B_oHQ6x86A1_0),.dout(w_dff_B_4hfbee0s3_0),.clk(gclk));
	jdff dff_B_xdFdkSUS6_0(.din(w_dff_B_4hfbee0s3_0),.dout(w_dff_B_xdFdkSUS6_0),.clk(gclk));
	jdff dff_B_CRDpuNq14_0(.din(n255),.dout(w_dff_B_CRDpuNq14_0),.clk(gclk));
	jdff dff_B_Wmu07nX56_0(.din(w_dff_B_CRDpuNq14_0),.dout(w_dff_B_Wmu07nX56_0),.clk(gclk));
	jdff dff_B_EOM0QiK69_0(.din(n250),.dout(w_dff_B_EOM0QiK69_0),.clk(gclk));
	jdff dff_A_vZtyeN6G0_0(.dout(w_n249_0[0]),.din(w_dff_A_vZtyeN6G0_0),.clk(gclk));
	jdff dff_A_qF97oLAq4_0(.dout(w_dff_A_vZtyeN6G0_0),.din(w_dff_A_qF97oLAq4_0),.clk(gclk));
	jdff dff_B_yzKj40tv6_0(.din(n248),.dout(w_dff_B_yzKj40tv6_0),.clk(gclk));
	jdff dff_B_289zX16p1_0(.din(w_dff_B_yzKj40tv6_0),.dout(w_dff_B_289zX16p1_0),.clk(gclk));
	jdff dff_B_GpDgQbzg3_0(.din(n244),.dout(w_dff_B_GpDgQbzg3_0),.clk(gclk));
	jdff dff_B_u34d1zbb2_0(.din(w_dff_B_GpDgQbzg3_0),.dout(w_dff_B_u34d1zbb2_0),.clk(gclk));
	jdff dff_B_apkQf78x5_0(.din(w_dff_B_u34d1zbb2_0),.dout(w_dff_B_apkQf78x5_0),.clk(gclk));
	jdff dff_B_8bptot6U4_1(.din(n276),.dout(w_dff_B_8bptot6U4_1),.clk(gclk));
	jdff dff_B_8jT7SjKR1_1(.din(n277),.dout(w_dff_B_8jT7SjKR1_1),.clk(gclk));
	jdff dff_B_m3WdSuYS8_1(.din(w_dff_B_8jT7SjKR1_1),.dout(w_dff_B_m3WdSuYS8_1),.clk(gclk));
	jdff dff_B_xoFZ9m0Q5_1(.din(w_dff_B_m3WdSuYS8_1),.dout(w_dff_B_xoFZ9m0Q5_1),.clk(gclk));
	jdff dff_B_5rdrazH21_1(.din(w_dff_B_xoFZ9m0Q5_1),.dout(w_dff_B_5rdrazH21_1),.clk(gclk));
	jdff dff_B_wrzresxM1_1(.din(w_dff_B_5rdrazH21_1),.dout(w_dff_B_wrzresxM1_1),.clk(gclk));
	jdff dff_B_B0PUDSaL1_1(.din(w_dff_B_wrzresxM1_1),.dout(w_dff_B_B0PUDSaL1_1),.clk(gclk));
	jdff dff_B_4Ubn4dbK3_1(.din(w_dff_B_B0PUDSaL1_1),.dout(w_dff_B_4Ubn4dbK3_1),.clk(gclk));
	jdff dff_B_PbRPsO087_1(.din(w_dff_B_4Ubn4dbK3_1),.dout(w_dff_B_PbRPsO087_1),.clk(gclk));
	jdff dff_B_iCce1xkd1_1(.din(w_dff_B_PbRPsO087_1),.dout(w_dff_B_iCce1xkd1_1),.clk(gclk));
	jdff dff_B_KLJ5GnLK6_1(.din(w_dff_B_iCce1xkd1_1),.dout(w_dff_B_KLJ5GnLK6_1),.clk(gclk));
	jdff dff_B_5lrRqkCa5_1(.din(w_dff_B_KLJ5GnLK6_1),.dout(w_dff_B_5lrRqkCa5_1),.clk(gclk));
	jdff dff_B_XZG5oczu4_0(.din(n343),.dout(w_dff_B_XZG5oczu4_0),.clk(gclk));
	jdff dff_B_fScDFGmE2_0(.din(w_dff_B_XZG5oczu4_0),.dout(w_dff_B_fScDFGmE2_0),.clk(gclk));
	jdff dff_B_RbllD0ED1_0(.din(w_dff_B_fScDFGmE2_0),.dout(w_dff_B_RbllD0ED1_0),.clk(gclk));
	jdff dff_B_2bokdNiJ8_0(.din(w_dff_B_RbllD0ED1_0),.dout(w_dff_B_2bokdNiJ8_0),.clk(gclk));
	jdff dff_B_SMY5Hzsc2_0(.din(w_dff_B_2bokdNiJ8_0),.dout(w_dff_B_SMY5Hzsc2_0),.clk(gclk));
	jdff dff_B_PgBXu2QW0_0(.din(w_dff_B_SMY5Hzsc2_0),.dout(w_dff_B_PgBXu2QW0_0),.clk(gclk));
	jdff dff_B_yleaMZuA9_0(.din(w_dff_B_PgBXu2QW0_0),.dout(w_dff_B_yleaMZuA9_0),.clk(gclk));
	jdff dff_B_Zgj2cefF6_0(.din(w_dff_B_yleaMZuA9_0),.dout(w_dff_B_Zgj2cefF6_0),.clk(gclk));
	jdff dff_B_0QkUNGRR8_0(.din(w_dff_B_Zgj2cefF6_0),.dout(w_dff_B_0QkUNGRR8_0),.clk(gclk));
	jdff dff_B_Q1dCM7WX8_0(.din(w_dff_B_0QkUNGRR8_0),.dout(w_dff_B_Q1dCM7WX8_0),.clk(gclk));
	jdff dff_B_pPDCAFuE9_0(.din(w_dff_B_Q1dCM7WX8_0),.dout(w_dff_B_pPDCAFuE9_0),.clk(gclk));
	jdff dff_B_IdsyYkH62_0(.din(w_dff_B_pPDCAFuE9_0),.dout(w_dff_B_IdsyYkH62_0),.clk(gclk));
	jdff dff_B_eRpUBvpO3_0(.din(w_dff_B_IdsyYkH62_0),.dout(w_dff_B_eRpUBvpO3_0),.clk(gclk));
	jdff dff_B_dZJonO2V5_0(.din(w_dff_B_eRpUBvpO3_0),.dout(w_dff_B_dZJonO2V5_0),.clk(gclk));
	jdff dff_A_tghaUmpO5_1(.dout(w_n274_0[1]),.din(w_dff_A_tghaUmpO5_1),.clk(gclk));
	jdff dff_A_SPJlyURP8_1(.dout(w_dff_A_tghaUmpO5_1),.din(w_dff_A_SPJlyURP8_1),.clk(gclk));
	jdff dff_A_cakV6Asy8_1(.dout(w_dff_A_SPJlyURP8_1),.din(w_dff_A_cakV6Asy8_1),.clk(gclk));
	jdff dff_A_7k7rpdAV8_1(.dout(w_dff_A_cakV6Asy8_1),.din(w_dff_A_7k7rpdAV8_1),.clk(gclk));
	jdff dff_A_fGqdGEo11_1(.dout(w_dff_A_7k7rpdAV8_1),.din(w_dff_A_fGqdGEo11_1),.clk(gclk));
	jdff dff_A_jqUECqvU3_1(.dout(w_dff_A_fGqdGEo11_1),.din(w_dff_A_jqUECqvU3_1),.clk(gclk));
	jdff dff_A_kfHkVYdZ7_1(.dout(w_dff_A_jqUECqvU3_1),.din(w_dff_A_kfHkVYdZ7_1),.clk(gclk));
	jdff dff_A_wp6dSsHc0_1(.dout(w_dff_A_kfHkVYdZ7_1),.din(w_dff_A_wp6dSsHc0_1),.clk(gclk));
	jdff dff_A_2e1PIBh61_1(.dout(w_dff_A_wp6dSsHc0_1),.din(w_dff_A_2e1PIBh61_1),.clk(gclk));
	jdff dff_A_CltLlal05_1(.dout(w_dff_A_2e1PIBh61_1),.din(w_dff_A_CltLlal05_1),.clk(gclk));
	jdff dff_A_UDBtD4919_1(.dout(w_dff_A_CltLlal05_1),.din(w_dff_A_UDBtD4919_1),.clk(gclk));
	jdff dff_A_753kcTCD8_1(.dout(w_dff_A_UDBtD4919_1),.din(w_dff_A_753kcTCD8_1),.clk(gclk));
	jdff dff_A_fcy4FWCD2_1(.dout(w_dff_A_753kcTCD8_1),.din(w_dff_A_fcy4FWCD2_1),.clk(gclk));
	jdff dff_A_bbOLXKZv3_1(.dout(w_dff_A_fcy4FWCD2_1),.din(w_dff_A_bbOLXKZv3_1),.clk(gclk));
	jdff dff_A_p6LfYgvw2_1(.dout(w_dff_A_bbOLXKZv3_1),.din(w_dff_A_p6LfYgvw2_1),.clk(gclk));
	jdff dff_A_mYKh4gra4_1(.dout(w_G902_2[1]),.din(w_dff_A_mYKh4gra4_1),.clk(gclk));
	jdff dff_A_XWPLXkbd7_1(.dout(w_dff_A_mYKh4gra4_1),.din(w_dff_A_XWPLXkbd7_1),.clk(gclk));
	jdff dff_A_OvCn3US17_1(.dout(w_dff_A_XWPLXkbd7_1),.din(w_dff_A_OvCn3US17_1),.clk(gclk));
	jdff dff_A_tCsfNudJ3_1(.dout(w_dff_A_OvCn3US17_1),.din(w_dff_A_tCsfNudJ3_1),.clk(gclk));
	jdff dff_A_DVFHJ7Yf3_1(.dout(w_dff_A_tCsfNudJ3_1),.din(w_dff_A_DVFHJ7Yf3_1),.clk(gclk));
	jdff dff_A_geUV8zZN0_1(.dout(w_dff_A_DVFHJ7Yf3_1),.din(w_dff_A_geUV8zZN0_1),.clk(gclk));
	jdff dff_A_hBhBAH5X3_1(.dout(w_dff_A_geUV8zZN0_1),.din(w_dff_A_hBhBAH5X3_1),.clk(gclk));
	jdff dff_A_S0EBWjgW5_1(.dout(w_dff_A_hBhBAH5X3_1),.din(w_dff_A_S0EBWjgW5_1),.clk(gclk));
	jdff dff_A_kYJkkiDr6_1(.dout(w_dff_A_S0EBWjgW5_1),.din(w_dff_A_kYJkkiDr6_1),.clk(gclk));
	jdff dff_A_zJkIfS6s9_1(.dout(w_dff_A_kYJkkiDr6_1),.din(w_dff_A_zJkIfS6s9_1),.clk(gclk));
	jdff dff_A_qS4IVq449_1(.dout(w_dff_A_zJkIfS6s9_1),.din(w_dff_A_qS4IVq449_1),.clk(gclk));
	jdff dff_A_NLCYjfDY7_1(.dout(w_dff_A_qS4IVq449_1),.din(w_dff_A_NLCYjfDY7_1),.clk(gclk));
	jdff dff_A_Kb9lV6dn4_1(.dout(w_dff_A_NLCYjfDY7_1),.din(w_dff_A_Kb9lV6dn4_1),.clk(gclk));
	jdff dff_A_EG8S5HFF4_1(.dout(w_dff_A_Kb9lV6dn4_1),.din(w_dff_A_EG8S5HFF4_1),.clk(gclk));
	jdff dff_A_scQnXMZO7_1(.dout(w_dff_A_EG8S5HFF4_1),.din(w_dff_A_scQnXMZO7_1),.clk(gclk));
	jdff dff_A_UA7Si7RF3_1(.dout(w_dff_A_scQnXMZO7_1),.din(w_dff_A_UA7Si7RF3_1),.clk(gclk));
	jdff dff_A_qxF7e5cA0_1(.dout(w_dff_A_UA7Si7RF3_1),.din(w_dff_A_qxF7e5cA0_1),.clk(gclk));
	jdff dff_A_aMP8TxdD8_2(.dout(w_G902_2[2]),.din(w_dff_A_aMP8TxdD8_2),.clk(gclk));
	jdff dff_A_RJpXreUj8_2(.dout(w_dff_A_aMP8TxdD8_2),.din(w_dff_A_RJpXreUj8_2),.clk(gclk));
	jdff dff_A_SzIJBEkJ2_2(.dout(w_dff_A_RJpXreUj8_2),.din(w_dff_A_SzIJBEkJ2_2),.clk(gclk));
	jdff dff_A_iHdRgjGT8_2(.dout(w_dff_A_SzIJBEkJ2_2),.din(w_dff_A_iHdRgjGT8_2),.clk(gclk));
	jdff dff_A_c60Amz7F7_2(.dout(w_dff_A_iHdRgjGT8_2),.din(w_dff_A_c60Amz7F7_2),.clk(gclk));
	jdff dff_A_LawalTON3_2(.dout(w_dff_A_c60Amz7F7_2),.din(w_dff_A_LawalTON3_2),.clk(gclk));
	jdff dff_A_662gdWoi6_2(.dout(w_dff_A_LawalTON3_2),.din(w_dff_A_662gdWoi6_2),.clk(gclk));
	jdff dff_A_y7T4zg6q8_2(.dout(w_dff_A_662gdWoi6_2),.din(w_dff_A_y7T4zg6q8_2),.clk(gclk));
	jdff dff_A_aU4dkGcP3_2(.dout(w_dff_A_y7T4zg6q8_2),.din(w_dff_A_aU4dkGcP3_2),.clk(gclk));
	jdff dff_A_TXnEezUI4_2(.dout(w_dff_A_aU4dkGcP3_2),.din(w_dff_A_TXnEezUI4_2),.clk(gclk));
	jdff dff_A_BdKpp2w27_2(.dout(w_dff_A_TXnEezUI4_2),.din(w_dff_A_BdKpp2w27_2),.clk(gclk));
	jdff dff_A_VK7IZjKm2_2(.dout(w_dff_A_BdKpp2w27_2),.din(w_dff_A_VK7IZjKm2_2),.clk(gclk));
	jdff dff_A_glg6sRqQ9_2(.dout(w_dff_A_VK7IZjKm2_2),.din(w_dff_A_glg6sRqQ9_2),.clk(gclk));
	jdff dff_A_Fr9tkfCD7_2(.dout(w_dff_A_glg6sRqQ9_2),.din(w_dff_A_Fr9tkfCD7_2),.clk(gclk));
	jdff dff_A_50hE6mO46_2(.dout(w_dff_A_Fr9tkfCD7_2),.din(w_dff_A_50hE6mO46_2),.clk(gclk));
	jdff dff_A_gipLDijG6_2(.dout(w_dff_A_50hE6mO46_2),.din(w_dff_A_gipLDijG6_2),.clk(gclk));
	jdff dff_A_eA2euOQv1_2(.dout(w_dff_A_gipLDijG6_2),.din(w_dff_A_eA2euOQv1_2),.clk(gclk));
	jdff dff_A_5FhJvPGZ3_0(.dout(w_n265_1[0]),.din(w_dff_A_5FhJvPGZ3_0),.clk(gclk));
	jdff dff_A_2LxxnF2Y5_1(.dout(w_n265_1[1]),.din(w_dff_A_2LxxnF2Y5_1),.clk(gclk));
	jdff dff_B_oDFlLFrH6_1(.din(n356),.dout(w_dff_B_oDFlLFrH6_1),.clk(gclk));
	jdff dff_B_kkZGT5ex4_1(.din(w_dff_B_oDFlLFrH6_1),.dout(w_dff_B_kkZGT5ex4_1),.clk(gclk));
	jdff dff_B_xpkfFFE45_1(.din(w_dff_B_kkZGT5ex4_1),.dout(w_dff_B_xpkfFFE45_1),.clk(gclk));
	jdff dff_B_jqqewpTn7_1(.din(w_dff_B_xpkfFFE45_1),.dout(w_dff_B_jqqewpTn7_1),.clk(gclk));
	jdff dff_B_K1oilr9n8_1(.din(w_dff_B_jqqewpTn7_1),.dout(w_dff_B_K1oilr9n8_1),.clk(gclk));
	jdff dff_B_ME0ctDw45_1(.din(w_dff_B_K1oilr9n8_1),.dout(w_dff_B_ME0ctDw45_1),.clk(gclk));
	jdff dff_B_2i56dJIx9_1(.din(w_dff_B_ME0ctDw45_1),.dout(w_dff_B_2i56dJIx9_1),.clk(gclk));
	jdff dff_B_k5H5qfgk9_1(.din(w_dff_B_2i56dJIx9_1),.dout(w_dff_B_k5H5qfgk9_1),.clk(gclk));
	jdff dff_B_ca6pTKAa9_1(.din(w_dff_B_k5H5qfgk9_1),.dout(w_dff_B_ca6pTKAa9_1),.clk(gclk));
	jdff dff_B_Q4JEGFuY1_1(.din(w_dff_B_ca6pTKAa9_1),.dout(w_dff_B_Q4JEGFuY1_1),.clk(gclk));
	jdff dff_B_AeyW46c71_1(.din(w_dff_B_Q4JEGFuY1_1),.dout(w_dff_B_AeyW46c71_1),.clk(gclk));
	jdff dff_B_BJrzF2mA7_1(.din(w_dff_B_AeyW46c71_1),.dout(w_dff_B_BJrzF2mA7_1),.clk(gclk));
	jdff dff_B_bnANAjms4_0(.din(n359),.dout(w_dff_B_bnANAjms4_0),.clk(gclk));
	jdff dff_B_uViSEPFG6_0(.din(w_dff_B_bnANAjms4_0),.dout(w_dff_B_uViSEPFG6_0),.clk(gclk));
	jdff dff_B_Tof3qMPu7_0(.din(w_dff_B_uViSEPFG6_0),.dout(w_dff_B_Tof3qMPu7_0),.clk(gclk));
	jdff dff_B_1LrVve8r9_0(.din(w_dff_B_Tof3qMPu7_0),.dout(w_dff_B_1LrVve8r9_0),.clk(gclk));
	jdff dff_B_NMgCGL556_0(.din(w_dff_B_1LrVve8r9_0),.dout(w_dff_B_NMgCGL556_0),.clk(gclk));
	jdff dff_B_f95KTXUO2_0(.din(w_dff_B_NMgCGL556_0),.dout(w_dff_B_f95KTXUO2_0),.clk(gclk));
	jdff dff_B_vlrt9UZ56_0(.din(w_dff_B_f95KTXUO2_0),.dout(w_dff_B_vlrt9UZ56_0),.clk(gclk));
	jdff dff_B_xlvujJv19_0(.din(w_dff_B_vlrt9UZ56_0),.dout(w_dff_B_xlvujJv19_0),.clk(gclk));
	jdff dff_B_KVJyetJt7_0(.din(w_dff_B_xlvujJv19_0),.dout(w_dff_B_KVJyetJt7_0),.clk(gclk));
	jdff dff_B_SM8ao1kl0_0(.din(w_dff_B_KVJyetJt7_0),.dout(w_dff_B_SM8ao1kl0_0),.clk(gclk));
	jdff dff_B_fUpP4j4k8_0(.din(w_dff_B_SM8ao1kl0_0),.dout(w_dff_B_fUpP4j4k8_0),.clk(gclk));
	jdff dff_B_0q1XVR3r5_0(.din(w_dff_B_fUpP4j4k8_0),.dout(w_dff_B_0q1XVR3r5_0),.clk(gclk));
	jdff dff_B_LxmA6KS07_0(.din(w_dff_B_0q1XVR3r5_0),.dout(w_dff_B_LxmA6KS07_0),.clk(gclk));
	jdff dff_B_CIDRaylk5_0(.din(w_dff_B_LxmA6KS07_0),.dout(w_dff_B_CIDRaylk5_0),.clk(gclk));
	jdff dff_B_YKHt5J0m8_1(.din(n302),.dout(w_dff_B_YKHt5J0m8_1),.clk(gclk));
	jdff dff_B_0LxZ9BDq7_1(.din(n304),.dout(w_dff_B_0LxZ9BDq7_1),.clk(gclk));
	jdff dff_B_mg6vrPOX5_1(.din(n285),.dout(w_dff_B_mg6vrPOX5_1),.clk(gclk));
	jdff dff_B_50NgK2HR5_1(.din(n290),.dout(w_dff_B_50NgK2HR5_1),.clk(gclk));
	jdff dff_B_sMOGxZUK7_2(.din(n297),.dout(w_dff_B_sMOGxZUK7_2),.clk(gclk));
	jdff dff_A_N5usaIeo9_1(.dout(w_n291_1[1]),.din(w_dff_A_N5usaIeo9_1),.clk(gclk));
	jdff dff_B_d1LbOOHB1_2(.din(n279),.dout(w_dff_B_d1LbOOHB1_2),.clk(gclk));
	jdff dff_A_mbPiTqZQ8_2(.dout(w_n278_0[2]),.din(w_dff_A_mbPiTqZQ8_2),.clk(gclk));
	jdff dff_A_mDT284LI8_2(.dout(w_dff_A_mbPiTqZQ8_2),.din(w_dff_A_mDT284LI8_2),.clk(gclk));
	jdff dff_B_baiLUCyu9_3(.din(n278),.dout(w_dff_B_baiLUCyu9_3),.clk(gclk));
	jdff dff_B_UvX1D9mq7_3(.din(w_dff_B_baiLUCyu9_3),.dout(w_dff_B_UvX1D9mq7_3),.clk(gclk));
	jdff dff_B_CBkZFcZr1_0(.din(n367),.dout(w_dff_B_CBkZFcZr1_0),.clk(gclk));
	jdff dff_B_BlbbzFwu8_0(.din(w_dff_B_CBkZFcZr1_0),.dout(w_dff_B_BlbbzFwu8_0),.clk(gclk));
	jdff dff_B_fjvq7sK88_0(.din(w_dff_B_BlbbzFwu8_0),.dout(w_dff_B_fjvq7sK88_0),.clk(gclk));
	jdff dff_B_8XGhWZXF1_0(.din(w_dff_B_fjvq7sK88_0),.dout(w_dff_B_8XGhWZXF1_0),.clk(gclk));
	jdff dff_B_rl3VHiSm3_0(.din(w_dff_B_8XGhWZXF1_0),.dout(w_dff_B_rl3VHiSm3_0),.clk(gclk));
	jdff dff_B_Pcqve8FC6_0(.din(w_dff_B_rl3VHiSm3_0),.dout(w_dff_B_Pcqve8FC6_0),.clk(gclk));
	jdff dff_B_dlKiSWxK3_0(.din(w_dff_B_Pcqve8FC6_0),.dout(w_dff_B_dlKiSWxK3_0),.clk(gclk));
	jdff dff_B_cbHEKBl85_0(.din(w_dff_B_dlKiSWxK3_0),.dout(w_dff_B_cbHEKBl85_0),.clk(gclk));
	jdff dff_B_YFxpDKCm0_0(.din(w_dff_B_cbHEKBl85_0),.dout(w_dff_B_YFxpDKCm0_0),.clk(gclk));
	jdff dff_B_R1AXzCN50_0(.din(w_dff_B_YFxpDKCm0_0),.dout(w_dff_B_R1AXzCN50_0),.clk(gclk));
	jdff dff_B_Hmziks3v6_0(.din(w_dff_B_R1AXzCN50_0),.dout(w_dff_B_Hmziks3v6_0),.clk(gclk));
	jdff dff_B_7zCrDNGV5_0(.din(w_dff_B_Hmziks3v6_0),.dout(w_dff_B_7zCrDNGV5_0),.clk(gclk));
	jdff dff_B_asktv9BC0_0(.din(n364),.dout(w_dff_B_asktv9BC0_0),.clk(gclk));
	jdff dff_B_GOGYS8gI2_0(.din(w_dff_B_asktv9BC0_0),.dout(w_dff_B_GOGYS8gI2_0),.clk(gclk));
	jdff dff_B_7U5xAF7x3_0(.din(w_dff_B_GOGYS8gI2_0),.dout(w_dff_B_7U5xAF7x3_0),.clk(gclk));
	jdff dff_B_6iqi2rmt3_0(.din(w_dff_B_7U5xAF7x3_0),.dout(w_dff_B_6iqi2rmt3_0),.clk(gclk));
	jdff dff_B_G6eqx5cE5_0(.din(w_dff_B_6iqi2rmt3_0),.dout(w_dff_B_G6eqx5cE5_0),.clk(gclk));
	jdff dff_B_O3xIvpoG1_0(.din(w_dff_B_G6eqx5cE5_0),.dout(w_dff_B_O3xIvpoG1_0),.clk(gclk));
	jdff dff_B_jz97CtEX7_0(.din(w_dff_B_O3xIvpoG1_0),.dout(w_dff_B_jz97CtEX7_0),.clk(gclk));
	jdff dff_B_vE5mbV9l5_0(.din(w_dff_B_jz97CtEX7_0),.dout(w_dff_B_vE5mbV9l5_0),.clk(gclk));
	jdff dff_B_UjTeNUhL0_0(.din(w_dff_B_vE5mbV9l5_0),.dout(w_dff_B_UjTeNUhL0_0),.clk(gclk));
	jdff dff_B_brPlIuhZ1_0(.din(w_dff_B_UjTeNUhL0_0),.dout(w_dff_B_brPlIuhZ1_0),.clk(gclk));
	jdff dff_B_jMb14Fsk5_0(.din(w_dff_B_brPlIuhZ1_0),.dout(w_dff_B_jMb14Fsk5_0),.clk(gclk));
	jdff dff_B_QvNXZIlv1_0(.din(w_dff_B_jMb14Fsk5_0),.dout(w_dff_B_QvNXZIlv1_0),.clk(gclk));
	jdff dff_B_M1X8Cc2u7_0(.din(w_dff_B_QvNXZIlv1_0),.dout(w_dff_B_M1X8Cc2u7_0),.clk(gclk));
	jdff dff_B_XytGs9et4_0(.din(w_dff_B_M1X8Cc2u7_0),.dout(w_dff_B_XytGs9et4_0),.clk(gclk));
	jdff dff_B_WoMQU8Xr6_1(.din(n326),.dout(w_dff_B_WoMQU8Xr6_1),.clk(gclk));
	jdff dff_B_ARLySCip4_1(.din(n331),.dout(w_dff_B_ARLySCip4_1),.clk(gclk));
	jdff dff_B_L52U40XV7_1(.din(n333),.dout(w_dff_B_L52U40XV7_1),.clk(gclk));
	jdff dff_A_92hYar444_1(.dout(w_n282_0[1]),.din(w_dff_A_92hYar444_1),.clk(gclk));
	jdff dff_A_5ld2p0Q47_2(.dout(w_n282_0[2]),.din(w_dff_A_5ld2p0Q47_2),.clk(gclk));
	jdff dff_A_p4wmA6dm0_1(.dout(w_n258_0[1]),.din(w_dff_A_p4wmA6dm0_1),.clk(gclk));
	jdff dff_A_eXF0yj0D6_1(.dout(w_dff_A_p4wmA6dm0_1),.din(w_dff_A_eXF0yj0D6_1),.clk(gclk));
	jdff dff_A_jRuMaBaC7_1(.dout(w_dff_A_eXF0yj0D6_1),.din(w_dff_A_jRuMaBaC7_1),.clk(gclk));
	jdff dff_A_lWXx1Z5k6_2(.dout(w_n258_0[2]),.din(w_dff_A_lWXx1Z5k6_2),.clk(gclk));
	jdff dff_A_GlRQ3DSW3_1(.dout(w_n287_0[1]),.din(w_dff_A_GlRQ3DSW3_1),.clk(gclk));
	jdff dff_A_e4tCZxkY8_0(.dout(w_n291_0[0]),.din(w_dff_A_e4tCZxkY8_0),.clk(gclk));
	jdff dff_A_cgR5SqR31_2(.dout(w_n291_0[2]),.din(w_dff_A_cgR5SqR31_2),.clk(gclk));
	jdff dff_A_ESH28Yld7_0(.dout(w_n322_0[0]),.din(w_dff_A_ESH28Yld7_0),.clk(gclk));
	jdff dff_A_IKnNahbU2_1(.dout(w_n303_0[1]),.din(w_dff_A_IKnNahbU2_1),.clk(gclk));
	jdff dff_B_mZMqktea3_2(.din(n303),.dout(w_dff_B_mZMqktea3_2),.clk(gclk));
	jdff dff_A_t0AN5XoL1_0(.dout(w_n307_0[0]),.din(w_dff_A_t0AN5XoL1_0),.clk(gclk));
	jdff dff_A_b8HLrhFj1_2(.dout(w_n307_0[2]),.din(w_dff_A_b8HLrhFj1_2),.clk(gclk));
	jdff dff_A_nT7IT46z9_0(.dout(w_n317_0[0]),.din(w_dff_A_nT7IT46z9_0),.clk(gclk));
	jdff dff_A_474pC7iS8_2(.dout(w_n317_0[2]),.din(w_dff_A_474pC7iS8_2),.clk(gclk));
	jdff dff_B_vhhNAn034_3(.din(n317),.dout(w_dff_B_vhhNAn034_3),.clk(gclk));
	jdff dff_B_l6WeeIPA1_3(.din(w_dff_B_vhhNAn034_3),.dout(w_dff_B_l6WeeIPA1_3),.clk(gclk));
	jdff dff_A_WRKgB4gP3_1(.dout(w_n316_0[1]),.din(w_dff_A_WRKgB4gP3_1),.clk(gclk));
	jdff dff_A_DGIu3rtn2_2(.dout(w_n316_0[2]),.din(w_dff_A_DGIu3rtn2_2),.clk(gclk));
	jdff dff_B_3funJieQ8_0(.din(n369),.dout(w_dff_B_3funJieQ8_0),.clk(gclk));
	jdff dff_B_rHg0aR1x2_0(.din(w_dff_B_3funJieQ8_0),.dout(w_dff_B_rHg0aR1x2_0),.clk(gclk));
	jdff dff_B_xdvJCgyA3_0(.din(w_dff_B_rHg0aR1x2_0),.dout(w_dff_B_xdvJCgyA3_0),.clk(gclk));
	jdff dff_B_sChwiXBc3_0(.din(w_dff_B_xdvJCgyA3_0),.dout(w_dff_B_sChwiXBc3_0),.clk(gclk));
	jdff dff_B_YghbJD1r6_0(.din(w_dff_B_sChwiXBc3_0),.dout(w_dff_B_YghbJD1r6_0),.clk(gclk));
	jdff dff_B_JTOIhjbR0_0(.din(w_dff_B_YghbJD1r6_0),.dout(w_dff_B_JTOIhjbR0_0),.clk(gclk));
	jdff dff_B_whwpl6tL4_0(.din(w_dff_B_JTOIhjbR0_0),.dout(w_dff_B_whwpl6tL4_0),.clk(gclk));
	jdff dff_B_WKEiH8V11_0(.din(w_dff_B_whwpl6tL4_0),.dout(w_dff_B_WKEiH8V11_0),.clk(gclk));
	jdff dff_B_RJolY06a7_0(.din(w_dff_B_WKEiH8V11_0),.dout(w_dff_B_RJolY06a7_0),.clk(gclk));
	jdff dff_B_nDtIyK1b5_0(.din(w_dff_B_RJolY06a7_0),.dout(w_dff_B_nDtIyK1b5_0),.clk(gclk));
	jdff dff_B_CezhDRNi8_0(.din(w_dff_B_nDtIyK1b5_0),.dout(w_dff_B_CezhDRNi8_0),.clk(gclk));
	jdff dff_B_lAgyn7Xj9_0(.din(w_dff_B_CezhDRNi8_0),.dout(w_dff_B_lAgyn7Xj9_0),.clk(gclk));
	jdff dff_B_8cIoaHl79_0(.din(w_dff_B_lAgyn7Xj9_0),.dout(w_dff_B_8cIoaHl79_0),.clk(gclk));
	jdff dff_B_M8qScDlO8_0(.din(w_dff_B_8cIoaHl79_0),.dout(w_dff_B_M8qScDlO8_0),.clk(gclk));
	jdff dff_B_rRqdFC7O3_0(.din(w_dff_B_M8qScDlO8_0),.dout(w_dff_B_rRqdFC7O3_0),.clk(gclk));
	jdff dff_A_Ob9VAU6x7_1(.dout(w_G902_1[1]),.din(w_dff_A_Ob9VAU6x7_1),.clk(gclk));
	jdff dff_A_ysFF107H1_1(.dout(w_dff_A_Ob9VAU6x7_1),.din(w_dff_A_ysFF107H1_1),.clk(gclk));
	jdff dff_A_Et1FL7JO8_1(.dout(w_dff_A_ysFF107H1_1),.din(w_dff_A_Et1FL7JO8_1),.clk(gclk));
	jdff dff_A_1Nrd7bdF7_1(.dout(w_dff_A_Et1FL7JO8_1),.din(w_dff_A_1Nrd7bdF7_1),.clk(gclk));
	jdff dff_A_CSzVkNdn9_1(.dout(w_dff_A_1Nrd7bdF7_1),.din(w_dff_A_CSzVkNdn9_1),.clk(gclk));
	jdff dff_A_6j4EvXZe3_1(.dout(w_dff_A_CSzVkNdn9_1),.din(w_dff_A_6j4EvXZe3_1),.clk(gclk));
	jdff dff_A_OLB7P6zY3_1(.dout(w_dff_A_6j4EvXZe3_1),.din(w_dff_A_OLB7P6zY3_1),.clk(gclk));
	jdff dff_A_ktdHEVxd8_1(.dout(w_dff_A_OLB7P6zY3_1),.din(w_dff_A_ktdHEVxd8_1),.clk(gclk));
	jdff dff_A_ZwYm77281_1(.dout(w_dff_A_ktdHEVxd8_1),.din(w_dff_A_ZwYm77281_1),.clk(gclk));
	jdff dff_A_X2QLLxGJ3_1(.dout(w_dff_A_ZwYm77281_1),.din(w_dff_A_X2QLLxGJ3_1),.clk(gclk));
	jdff dff_A_4XJfn4QY0_1(.dout(w_dff_A_X2QLLxGJ3_1),.din(w_dff_A_4XJfn4QY0_1),.clk(gclk));
	jdff dff_A_LSYqAxwU5_1(.dout(w_dff_A_4XJfn4QY0_1),.din(w_dff_A_LSYqAxwU5_1),.clk(gclk));
	jdff dff_A_9BVGgBsK6_1(.dout(w_dff_A_LSYqAxwU5_1),.din(w_dff_A_9BVGgBsK6_1),.clk(gclk));
	jdff dff_A_pVWF1xs27_1(.dout(w_dff_A_9BVGgBsK6_1),.din(w_dff_A_pVWF1xs27_1),.clk(gclk));
	jdff dff_A_tjfRjIee7_1(.dout(w_dff_A_pVWF1xs27_1),.din(w_dff_A_tjfRjIee7_1),.clk(gclk));
	jdff dff_A_xqcT2hvA9_1(.dout(w_dff_A_tjfRjIee7_1),.din(w_dff_A_xqcT2hvA9_1),.clk(gclk));
	jdff dff_A_Y0O5LEFn9_1(.dout(w_dff_A_xqcT2hvA9_1),.din(w_dff_A_Y0O5LEFn9_1),.clk(gclk));
	jdff dff_A_BRjINC0z0_2(.dout(w_G902_1[2]),.din(w_dff_A_BRjINC0z0_2),.clk(gclk));
	jdff dff_A_4uYM1mso0_2(.dout(w_dff_A_BRjINC0z0_2),.din(w_dff_A_4uYM1mso0_2),.clk(gclk));
	jdff dff_A_VaBScGfd5_2(.dout(w_dff_A_4uYM1mso0_2),.din(w_dff_A_VaBScGfd5_2),.clk(gclk));
	jdff dff_A_YoVImA6k2_2(.dout(w_dff_A_VaBScGfd5_2),.din(w_dff_A_YoVImA6k2_2),.clk(gclk));
	jdff dff_A_kGodJQwH7_2(.dout(w_dff_A_YoVImA6k2_2),.din(w_dff_A_kGodJQwH7_2),.clk(gclk));
	jdff dff_A_goLhS2s04_2(.dout(w_dff_A_kGodJQwH7_2),.din(w_dff_A_goLhS2s04_2),.clk(gclk));
	jdff dff_A_KrMuT1pJ3_2(.dout(w_dff_A_goLhS2s04_2),.din(w_dff_A_KrMuT1pJ3_2),.clk(gclk));
	jdff dff_A_aAn6CQMd5_2(.dout(w_dff_A_KrMuT1pJ3_2),.din(w_dff_A_aAn6CQMd5_2),.clk(gclk));
	jdff dff_A_PbAlEzDK4_2(.dout(w_dff_A_aAn6CQMd5_2),.din(w_dff_A_PbAlEzDK4_2),.clk(gclk));
	jdff dff_A_ToiQrkkz7_2(.dout(w_dff_A_PbAlEzDK4_2),.din(w_dff_A_ToiQrkkz7_2),.clk(gclk));
	jdff dff_A_JFEL1nUo3_2(.dout(w_dff_A_ToiQrkkz7_2),.din(w_dff_A_JFEL1nUo3_2),.clk(gclk));
	jdff dff_A_rclqD4ZQ2_2(.dout(w_dff_A_JFEL1nUo3_2),.din(w_dff_A_rclqD4ZQ2_2),.clk(gclk));
	jdff dff_A_Gyoi4zx37_2(.dout(w_dff_A_rclqD4ZQ2_2),.din(w_dff_A_Gyoi4zx37_2),.clk(gclk));
	jdff dff_A_rafw39099_2(.dout(w_dff_A_Gyoi4zx37_2),.din(w_dff_A_rafw39099_2),.clk(gclk));
	jdff dff_A_4y5XQRZL7_2(.dout(w_dff_A_rafw39099_2),.din(w_dff_A_4y5XQRZL7_2),.clk(gclk));
	jdff dff_A_22myod8p8_2(.dout(w_dff_A_4y5XQRZL7_2),.din(w_dff_A_22myod8p8_2),.clk(gclk));
	jdff dff_A_pWNy4AKp6_2(.dout(w_dff_A_22myod8p8_2),.din(w_dff_A_pWNy4AKp6_2),.clk(gclk));
	jdff dff_B_2X3F5Utf0_1(.din(n236),.dout(w_dff_B_2X3F5Utf0_1),.clk(gclk));
	jdff dff_B_JXxE9l7T2_1(.din(n237),.dout(w_dff_B_JXxE9l7T2_1),.clk(gclk));
	jdff dff_A_xEIhDbgd1_0(.dout(w_n184_0[0]),.din(w_dff_A_xEIhDbgd1_0),.clk(gclk));
	jdff dff_A_C9ZSpTRT0_1(.dout(w_n183_0[1]),.din(w_dff_A_C9ZSpTRT0_1),.clk(gclk));
	jdff dff_A_DevZQJIz3_2(.dout(w_n183_0[2]),.din(w_dff_A_DevZQJIz3_2),.clk(gclk));
	jdff dff_A_LVBGMoP22_0(.dout(w_n216_1[0]),.din(w_dff_A_LVBGMoP22_0),.clk(gclk));
	jdff dff_A_QKfCqza18_2(.dout(w_n216_0[2]),.din(w_dff_A_QKfCqza18_2),.clk(gclk));
	jdff dff_B_ujxpdS7E3_0(.din(n213),.dout(w_dff_B_ujxpdS7E3_0),.clk(gclk));
	jdff dff_B_NgPS3SEX2_0(.din(w_dff_B_ujxpdS7E3_0),.dout(w_dff_B_NgPS3SEX2_0),.clk(gclk));
	jdff dff_B_twwOpmxt5_0(.din(w_dff_B_NgPS3SEX2_0),.dout(w_dff_B_twwOpmxt5_0),.clk(gclk));
	jdff dff_A_jo4ZeTVu3_1(.dout(w_n192_0[1]),.din(w_dff_A_jo4ZeTVu3_1),.clk(gclk));
	jdff dff_A_iSuFEqde4_0(.dout(w_n191_0[0]),.din(w_dff_A_iSuFEqde4_0),.clk(gclk));
	jdff dff_A_AVw7lWSl2_2(.dout(w_n191_0[2]),.din(w_dff_A_AVw7lWSl2_2),.clk(gclk));
	jdff dff_A_Yxw5h3ar9_1(.dout(w_n182_1[1]),.din(w_dff_A_Yxw5h3ar9_1),.clk(gclk));
	jdff dff_A_ceuQN59g7_0(.dout(w_n182_0[0]),.din(w_dff_A_ceuQN59g7_0),.clk(gclk));
	jdff dff_A_kAaKGw3K8_0(.dout(w_dff_A_ceuQN59g7_0),.din(w_dff_A_kAaKGw3K8_0),.clk(gclk));
	jdff dff_A_qupKCXvj3_0(.dout(w_dff_A_kAaKGw3K8_0),.din(w_dff_A_qupKCXvj3_0),.clk(gclk));
	jdff dff_A_sTeTl9j90_2(.dout(w_n182_0[2]),.din(w_dff_A_sTeTl9j90_2),.clk(gclk));
	jdff dff_A_XUkfqiMS7_2(.dout(w_dff_A_sTeTl9j90_2),.din(w_dff_A_XUkfqiMS7_2),.clk(gclk));
	jdff dff_A_wPdwgXWI3_2(.dout(w_dff_A_XUkfqiMS7_2),.din(w_dff_A_wPdwgXWI3_2),.clk(gclk));
	jdff dff_A_Kq7nAxjJ6_2(.dout(w_dff_A_wPdwgXWI3_2),.din(w_dff_A_Kq7nAxjJ6_2),.clk(gclk));
	jdff dff_A_LuAz3Zoz4_0(.dout(w_n180_0[0]),.din(w_dff_A_LuAz3Zoz4_0),.clk(gclk));
	jdff dff_A_j1v6xOuW7_1(.dout(w_G900_0[1]),.din(w_dff_A_j1v6xOuW7_1),.clk(gclk));
	jdff dff_A_pL9aPxaf8_1(.dout(w_n177_0[1]),.din(w_dff_A_pL9aPxaf8_1),.clk(gclk));
	jdff dff_A_NybkuwfE7_2(.dout(w_n177_0[2]),.din(w_dff_A_NybkuwfE7_2),.clk(gclk));
	jdff dff_A_YxtIsUQ09_0(.dout(w_n175_0[0]),.din(w_dff_A_YxtIsUQ09_0),.clk(gclk));
	jdff dff_A_dG3pUUhf3_1(.dout(w_n174_0[1]),.din(w_dff_A_dG3pUUhf3_1),.clk(gclk));
	jdff dff_B_TYA0jWKs3_2(.din(n174),.dout(w_dff_B_TYA0jWKs3_2),.clk(gclk));
	jdff dff_A_s5YjsonR8_1(.dout(w_n199_0[1]),.din(w_dff_A_s5YjsonR8_1),.clk(gclk));
	jdff dff_A_xQT8wLcD4_1(.dout(w_dff_A_s5YjsonR8_1),.din(w_dff_A_xQT8wLcD4_1),.clk(gclk));
	jdff dff_A_wHFsuuiJ8_0(.dout(w_n197_1[0]),.din(w_dff_A_wHFsuuiJ8_0),.clk(gclk));
	jdff dff_B_2T9zAfDd3_2(.din(n170),.dout(w_dff_B_2T9zAfDd3_2),.clk(gclk));
	jdff dff_A_D3qXC8054_2(.dout(w_n154_0[2]),.din(w_dff_A_D3qXC8054_2),.clk(gclk));
	jdff dff_A_wQssL4Lw9_2(.dout(w_dff_A_D3qXC8054_2),.din(w_dff_A_wQssL4Lw9_2),.clk(gclk));
	jdff dff_A_hoRXZfFF0_2(.dout(w_dff_A_wQssL4Lw9_2),.din(w_dff_A_hoRXZfFF0_2),.clk(gclk));
	jdff dff_A_GAFQXiQk6_2(.dout(w_dff_A_hoRXZfFF0_2),.din(w_dff_A_GAFQXiQk6_2),.clk(gclk));
	jdff dff_B_f6Q2iOXQ1_1(.din(n142),.dout(w_dff_B_f6Q2iOXQ1_1),.clk(gclk));
	jdff dff_B_789dvlrH7_1(.din(w_dff_B_f6Q2iOXQ1_1),.dout(w_dff_B_789dvlrH7_1),.clk(gclk));
	jdff dff_B_zoWnA3Sw9_1(.din(w_dff_B_789dvlrH7_1),.dout(w_dff_B_zoWnA3Sw9_1),.clk(gclk));
	jdff dff_B_2JLpDrk81_1(.din(w_dff_B_zoWnA3Sw9_1),.dout(w_dff_B_2JLpDrk81_1),.clk(gclk));
	jdff dff_B_gbbLE1r79_1(.din(w_dff_B_2JLpDrk81_1),.dout(w_dff_B_gbbLE1r79_1),.clk(gclk));
	jdff dff_A_yfhcaq8P3_1(.dout(w_n93_1[1]),.din(w_dff_A_yfhcaq8P3_1),.clk(gclk));
	jdff dff_A_a9FOPwLV5_1(.dout(w_dff_A_yfhcaq8P3_1),.din(w_dff_A_a9FOPwLV5_1),.clk(gclk));
	jdff dff_A_soEHyxz21_1(.dout(w_n93_0[1]),.din(w_dff_A_soEHyxz21_1),.clk(gclk));
	jdff dff_A_yMjaBLlH6_2(.dout(w_n93_0[2]),.din(w_dff_A_yMjaBLlH6_2),.clk(gclk));
	jdff dff_A_6gvA7Kvb2_0(.dout(w_n166_0[0]),.din(w_dff_A_6gvA7Kvb2_0),.clk(gclk));
	jdff dff_A_MX6iKdHZ7_1(.dout(w_n165_0[1]),.din(w_dff_A_MX6iKdHZ7_1),.clk(gclk));
	jdff dff_A_EZQQlWfd2_2(.dout(w_n165_0[2]),.din(w_dff_A_EZQQlWfd2_2),.clk(gclk));
	jdff dff_B_yxV8UGaj6_1(.din(n132),.dout(w_dff_B_yxV8UGaj6_1),.clk(gclk));
	jdff dff_B_Y4OnDzFr3_1(.din(w_dff_B_yxV8UGaj6_1),.dout(w_dff_B_Y4OnDzFr3_1),.clk(gclk));
	jdff dff_B_WJrPwGVT1_1(.din(w_dff_B_Y4OnDzFr3_1),.dout(w_dff_B_WJrPwGVT1_1),.clk(gclk));
	jdff dff_B_IfHaIX4n4_1(.din(w_dff_B_WJrPwGVT1_1),.dout(w_dff_B_IfHaIX4n4_1),.clk(gclk));
	jdff dff_B_Lhkdwcf79_1(.din(w_dff_B_IfHaIX4n4_1),.dout(w_dff_B_Lhkdwcf79_1),.clk(gclk));
	jdff dff_A_KOS7OcBZ2_1(.dout(w_n122_0[1]),.din(w_dff_A_KOS7OcBZ2_1),.clk(gclk));
	jdff dff_A_FJ51mBDe1_0(.dout(w_n208_0[0]),.din(w_dff_A_FJ51mBDe1_0),.clk(gclk));
	jdff dff_A_zhsHfnEm0_1(.dout(w_n197_0[1]),.din(w_dff_A_zhsHfnEm0_1),.clk(gclk));
	jdff dff_B_uzR4OQuH0_1(.din(n194),.dout(w_dff_B_uzR4OQuH0_1),.clk(gclk));
	jdff dff_B_2RgNAlMZ2_1(.din(w_dff_B_uzR4OQuH0_1),.dout(w_dff_B_2RgNAlMZ2_1),.clk(gclk));
	jdff dff_B_MWxUAb5E4_1(.din(w_dff_B_2RgNAlMZ2_1),.dout(w_dff_B_MWxUAb5E4_1),.clk(gclk));
	jdff dff_B_C0kAeFOd6_1(.din(w_dff_B_MWxUAb5E4_1),.dout(w_dff_B_C0kAeFOd6_1),.clk(gclk));
	jdff dff_B_3kB9E9WJ2_1(.din(w_dff_B_C0kAeFOd6_1),.dout(w_dff_B_3kB9E9WJ2_1),.clk(gclk));
	jdff dff_A_UYistIdV0_0(.dout(w_n118_0[0]),.din(w_dff_A_UYistIdV0_0),.clk(gclk));
	jdff dff_A_0fWTY5xz5_0(.dout(w_dff_A_UYistIdV0_0),.din(w_dff_A_0fWTY5xz5_0),.clk(gclk));
	jdff dff_A_BjEMlTet3_0(.dout(w_dff_A_0fWTY5xz5_0),.din(w_dff_A_BjEMlTet3_0),.clk(gclk));
	jdff dff_A_3AxcHWoe5_0(.dout(w_dff_A_BjEMlTet3_0),.din(w_dff_A_3AxcHWoe5_0),.clk(gclk));
	jdff dff_A_YCztvHnA2_0(.dout(w_dff_A_3AxcHWoe5_0),.din(w_dff_A_YCztvHnA2_0),.clk(gclk));
	jdff dff_A_DcxoOiIG4_0(.dout(w_dff_A_YCztvHnA2_0),.din(w_dff_A_DcxoOiIG4_0),.clk(gclk));
	jdff dff_A_omNvXYFU5_0(.dout(w_dff_A_DcxoOiIG4_0),.din(w_dff_A_omNvXYFU5_0),.clk(gclk));
	jdff dff_A_9RO2IyyX7_0(.dout(w_dff_A_omNvXYFU5_0),.din(w_dff_A_9RO2IyyX7_0),.clk(gclk));
	jdff dff_A_Q8zLMNXk4_0(.dout(w_dff_A_9RO2IyyX7_0),.din(w_dff_A_Q8zLMNXk4_0),.clk(gclk));
	jdff dff_A_MvPLNjpo1_0(.dout(w_dff_A_Q8zLMNXk4_0),.din(w_dff_A_MvPLNjpo1_0),.clk(gclk));
	jdff dff_A_PNR7F9bp4_0(.dout(w_dff_A_MvPLNjpo1_0),.din(w_dff_A_PNR7F9bp4_0),.clk(gclk));
	jdff dff_A_7QDaXC2d3_0(.dout(w_dff_A_PNR7F9bp4_0),.din(w_dff_A_7QDaXC2d3_0),.clk(gclk));
	jdff dff_A_DCDL6rW75_0(.dout(w_dff_A_7QDaXC2d3_0),.din(w_dff_A_DCDL6rW75_0),.clk(gclk));
	jdff dff_A_7WMoCQIU0_1(.dout(w_G227_0[1]),.din(w_dff_A_7WMoCQIU0_1),.clk(gclk));
	jdff dff_A_gjbdkYIb0_0(.dout(w_G469_0[0]),.din(w_dff_A_gjbdkYIb0_0),.clk(gclk));
	jdff dff_A_0zhemYdL4_0(.dout(w_dff_A_gjbdkYIb0_0),.din(w_dff_A_0zhemYdL4_0),.clk(gclk));
	jdff dff_A_khodaI6M6_0(.dout(w_dff_A_0zhemYdL4_0),.din(w_dff_A_khodaI6M6_0),.clk(gclk));
	jdff dff_A_Gv8l8Q3L8_0(.dout(w_dff_A_khodaI6M6_0),.din(w_dff_A_Gv8l8Q3L8_0),.clk(gclk));
	jdff dff_A_ag7Im9mg7_0(.dout(w_dff_A_Gv8l8Q3L8_0),.din(w_dff_A_ag7Im9mg7_0),.clk(gclk));
	jdff dff_A_b7e3vnuK8_0(.dout(w_dff_A_ag7Im9mg7_0),.din(w_dff_A_b7e3vnuK8_0),.clk(gclk));
	jdff dff_A_DWLzeQDI0_0(.dout(w_dff_A_b7e3vnuK8_0),.din(w_dff_A_DWLzeQDI0_0),.clk(gclk));
	jdff dff_A_M2CmPuwm5_0(.dout(w_dff_A_DWLzeQDI0_0),.din(w_dff_A_M2CmPuwm5_0),.clk(gclk));
	jdff dff_A_sXfm6t2m7_0(.dout(w_dff_A_M2CmPuwm5_0),.din(w_dff_A_sXfm6t2m7_0),.clk(gclk));
	jdff dff_A_H0R0gBJm9_0(.dout(w_dff_A_sXfm6t2m7_0),.din(w_dff_A_H0R0gBJm9_0),.clk(gclk));
	jdff dff_A_ihMVvcDN0_0(.dout(w_dff_A_H0R0gBJm9_0),.din(w_dff_A_ihMVvcDN0_0),.clk(gclk));
	jdff dff_A_Hf6EEOXC0_0(.dout(w_dff_A_ihMVvcDN0_0),.din(w_dff_A_Hf6EEOXC0_0),.clk(gclk));
	jdff dff_A_pfFUrYvS8_0(.dout(w_dff_A_Hf6EEOXC0_0),.din(w_dff_A_pfFUrYvS8_0),.clk(gclk));
	jdff dff_A_MFR2jh6Q4_0(.dout(w_dff_A_pfFUrYvS8_0),.din(w_dff_A_MFR2jh6Q4_0),.clk(gclk));
	jdff dff_A_r7RVUuaW0_0(.dout(w_dff_A_MFR2jh6Q4_0),.din(w_dff_A_r7RVUuaW0_0),.clk(gclk));
	jdff dff_A_hi8HOVFL6_0(.dout(w_dff_A_r7RVUuaW0_0),.din(w_dff_A_hi8HOVFL6_0),.clk(gclk));
	jdff dff_A_Tbf7fEPQ5_2(.dout(w_G469_0[2]),.din(w_dff_A_Tbf7fEPQ5_2),.clk(gclk));
	jdff dff_A_sg68VMId5_2(.dout(w_dff_A_Tbf7fEPQ5_2),.din(w_dff_A_sg68VMId5_2),.clk(gclk));
	jdff dff_A_PFpzELJV4_2(.dout(w_dff_A_sg68VMId5_2),.din(w_dff_A_PFpzELJV4_2),.clk(gclk));
	jdff dff_A_qyPaySJa3_2(.dout(w_dff_A_PFpzELJV4_2),.din(w_dff_A_qyPaySJa3_2),.clk(gclk));
	jdff dff_A_1FjSXV9z0_2(.dout(w_dff_A_qyPaySJa3_2),.din(w_dff_A_1FjSXV9z0_2),.clk(gclk));
	jdff dff_A_yjGMR8qv0_2(.dout(w_dff_A_1FjSXV9z0_2),.din(w_dff_A_yjGMR8qv0_2),.clk(gclk));
	jdff dff_A_iPJCIki71_1(.dout(w_n113_0[1]),.din(w_dff_A_iPJCIki71_1),.clk(gclk));
	jdff dff_A_viYe8xIr3_1(.dout(w_dff_A_iPJCIki71_1),.din(w_dff_A_viYe8xIr3_1),.clk(gclk));
	jdff dff_A_IDXMZJm00_2(.dout(w_n113_0[2]),.din(w_dff_A_IDXMZJm00_2),.clk(gclk));
	jdff dff_A_bFIRqKpw9_2(.dout(w_dff_A_IDXMZJm00_2),.din(w_dff_A_bFIRqKpw9_2),.clk(gclk));
	jdff dff_A_LFpjap0v7_1(.dout(w_n112_0[1]),.din(w_dff_A_LFpjap0v7_1),.clk(gclk));
	jdff dff_A_tQ6X6L0b4_1(.dout(w_dff_A_LFpjap0v7_1),.din(w_dff_A_tQ6X6L0b4_1),.clk(gclk));
	jdff dff_A_hj8rotjC3_1(.dout(w_dff_A_tQ6X6L0b4_1),.din(w_dff_A_hj8rotjC3_1),.clk(gclk));
	jdff dff_A_zW9L4dHS9_2(.dout(w_n112_0[2]),.din(w_dff_A_zW9L4dHS9_2),.clk(gclk));
	jdff dff_A_S133haJG2_2(.dout(w_dff_A_zW9L4dHS9_2),.din(w_dff_A_S133haJG2_2),.clk(gclk));
	jdff dff_A_23L3vLrA3_2(.dout(w_dff_A_S133haJG2_2),.din(w_dff_A_23L3vLrA3_2),.clk(gclk));
	jdff dff_A_ILbxSRX01_1(.dout(w_n109_0[1]),.din(w_dff_A_ILbxSRX01_1),.clk(gclk));
	jdff dff_A_u2vrMGRA8_1(.dout(w_dff_A_ILbxSRX01_1),.din(w_dff_A_u2vrMGRA8_1),.clk(gclk));
	jdff dff_A_gwtCXaDD2_1(.dout(w_dff_A_u2vrMGRA8_1),.din(w_dff_A_gwtCXaDD2_1),.clk(gclk));
	jdff dff_A_2zVWGoBz7_1(.dout(w_dff_A_gwtCXaDD2_1),.din(w_dff_A_2zVWGoBz7_1),.clk(gclk));
	jdff dff_A_0hn9qmfX6_0(.dout(w_n107_0[0]),.din(w_dff_A_0hn9qmfX6_0),.clk(gclk));
	jdff dff_A_Z9ohuSKm0_0(.dout(w_dff_A_0hn9qmfX6_0),.din(w_dff_A_Z9ohuSKm0_0),.clk(gclk));
	jdff dff_A_dn9w75tJ3_0(.dout(w_dff_A_Z9ohuSKm0_0),.din(w_dff_A_dn9w75tJ3_0),.clk(gclk));
	jdff dff_A_zyA0znkD5_0(.dout(w_dff_A_dn9w75tJ3_0),.din(w_dff_A_zyA0znkD5_0),.clk(gclk));
	jdff dff_A_NrlRSbuI4_0(.dout(w_dff_A_zyA0znkD5_0),.din(w_dff_A_NrlRSbuI4_0),.clk(gclk));
	jdff dff_A_igCyGVkT9_0(.dout(w_dff_A_NrlRSbuI4_0),.din(w_dff_A_igCyGVkT9_0),.clk(gclk));
	jdff dff_A_lGXE1MWv3_0(.dout(w_dff_A_igCyGVkT9_0),.din(w_dff_A_lGXE1MWv3_0),.clk(gclk));
	jdff dff_A_sDXGCA2C6_0(.dout(w_dff_A_lGXE1MWv3_0),.din(w_dff_A_sDXGCA2C6_0),.clk(gclk));
	jdff dff_A_zzUgZ3Vr9_0(.dout(w_dff_A_sDXGCA2C6_0),.din(w_dff_A_zzUgZ3Vr9_0),.clk(gclk));
	jdff dff_A_WXRgklfM4_0(.dout(w_dff_A_zzUgZ3Vr9_0),.din(w_dff_A_WXRgklfM4_0),.clk(gclk));
	jdff dff_A_FEe6EmbO6_0(.dout(w_dff_A_WXRgklfM4_0),.din(w_dff_A_FEe6EmbO6_0),.clk(gclk));
	jdff dff_A_V7pe8dpK8_0(.dout(w_dff_A_FEe6EmbO6_0),.din(w_dff_A_V7pe8dpK8_0),.clk(gclk));
	jdff dff_A_dOdQglT95_0(.dout(w_dff_A_V7pe8dpK8_0),.din(w_dff_A_dOdQglT95_0),.clk(gclk));
	jdff dff_B_dEj9vy825_1(.din(n104),.dout(w_dff_B_dEj9vy825_1),.clk(gclk));
	jdff dff_A_kSftgAv93_1(.dout(w_G224_0[1]),.din(w_dff_A_kSftgAv93_1),.clk(gclk));
	jdff dff_B_gGE3uEGs4_0(.din(n101),.dout(w_dff_B_gGE3uEGs4_0),.clk(gclk));
	jdff dff_B_C21Cr2AB5_0(.din(w_dff_B_gGE3uEGs4_0),.dout(w_dff_B_C21Cr2AB5_0),.clk(gclk));
	jdff dff_A_jjWIrSHE2_0(.dout(w_n99_0[0]),.din(w_dff_A_jjWIrSHE2_0),.clk(gclk));
	jdff dff_A_UANKoWfV5_1(.dout(w_n96_0[1]),.din(w_dff_A_UANKoWfV5_1),.clk(gclk));
	jdff dff_A_HTLSczVE8_1(.dout(w_dff_A_UANKoWfV5_1),.din(w_dff_A_HTLSczVE8_1),.clk(gclk));
	jdff dff_A_Big4gnsf9_2(.dout(w_n96_0[2]),.din(w_dff_A_Big4gnsf9_2),.clk(gclk));
	jdff dff_A_mPRuzlGc6_2(.dout(w_dff_A_Big4gnsf9_2),.din(w_dff_A_mPRuzlGc6_2),.clk(gclk));
	jdff dff_B_hVsy3OE97_3(.din(n96),.dout(w_dff_B_hVsy3OE97_3),.clk(gclk));
	jdff dff_B_836m1ysa9_3(.din(w_dff_B_hVsy3OE97_3),.dout(w_dff_B_836m1ysa9_3),.clk(gclk));
	jdff dff_A_jcYedj8v0_0(.dout(w_n95_1[0]),.din(w_dff_A_jcYedj8v0_0),.clk(gclk));
	jdff dff_A_3xNgarSq0_0(.dout(w_dff_A_jcYedj8v0_0),.din(w_dff_A_3xNgarSq0_0),.clk(gclk));
	jdff dff_A_Sqme8lOR8_1(.dout(w_n95_0[1]),.din(w_dff_A_Sqme8lOR8_1),.clk(gclk));
	jdff dff_A_VCwZPWoZ7_1(.dout(w_dff_A_Sqme8lOR8_1),.din(w_dff_A_VCwZPWoZ7_1),.clk(gclk));
	jdff dff_A_E0i33Pnj3_1(.dout(w_dff_A_VCwZPWoZ7_1),.din(w_dff_A_E0i33Pnj3_1),.clk(gclk));
	jdff dff_A_Pc05VXXJ3_1(.dout(w_dff_A_E0i33Pnj3_1),.din(w_dff_A_Pc05VXXJ3_1),.clk(gclk));
	jdff dff_A_VVcpvPLv4_1(.dout(w_dff_A_Pc05VXXJ3_1),.din(w_dff_A_VVcpvPLv4_1),.clk(gclk));
	jdff dff_A_YUuSe0jM1_2(.dout(w_n95_0[2]),.din(w_dff_A_YUuSe0jM1_2),.clk(gclk));
	jdff dff_A_RINZHuL81_2(.dout(w_dff_A_YUuSe0jM1_2),.din(w_dff_A_RINZHuL81_2),.clk(gclk));
	jdff dff_A_d2xjLCcJ0_2(.dout(w_dff_A_RINZHuL81_2),.din(w_dff_A_d2xjLCcJ0_2),.clk(gclk));
	jdff dff_A_Vk0unUv63_2(.dout(w_dff_A_d2xjLCcJ0_2),.din(w_dff_A_Vk0unUv63_2),.clk(gclk));
	jdff dff_A_s4HEiENx9_2(.dout(w_dff_A_Vk0unUv63_2),.din(w_dff_A_s4HEiENx9_2),.clk(gclk));
	jdff dff_A_akdZEYzP7_1(.dout(w_n161_0[1]),.din(w_dff_A_akdZEYzP7_1),.clk(gclk));
	jdff dff_A_LMQzXh8Y3_2(.dout(w_n161_0[2]),.din(w_dff_A_LMQzXh8Y3_2),.clk(gclk));
	jdff dff_B_9df6Tjnu5_3(.din(n161),.dout(w_dff_B_9df6Tjnu5_3),.clk(gclk));
	jdff dff_B_yQ6CoJCA8_1(.din(n159),.dout(w_dff_B_yQ6CoJCA8_1),.clk(gclk));
	jdff dff_B_hbFeXRny0_1(.din(w_dff_B_yQ6CoJCA8_1),.dout(w_dff_B_hbFeXRny0_1),.clk(gclk));
	jdff dff_B_e8gTMXUE6_1(.din(w_dff_B_hbFeXRny0_1),.dout(w_dff_B_e8gTMXUE6_1),.clk(gclk));
	jdff dff_B_DtM3fqRY8_1(.din(w_dff_B_e8gTMXUE6_1),.dout(w_dff_B_DtM3fqRY8_1),.clk(gclk));
	jdff dff_B_fW3ODDb64_1(.din(w_dff_B_DtM3fqRY8_1),.dout(w_dff_B_fW3ODDb64_1),.clk(gclk));
	jdff dff_A_nTA8dc2J4_0(.dout(w_n90_0[0]),.din(w_dff_A_nTA8dc2J4_0),.clk(gclk));
	jdff dff_A_arDw1qDP6_0(.dout(w_dff_A_nTA8dc2J4_0),.din(w_dff_A_arDw1qDP6_0),.clk(gclk));
	jdff dff_A_KdvZQnOx3_0(.dout(w_dff_A_arDw1qDP6_0),.din(w_dff_A_KdvZQnOx3_0),.clk(gclk));
	jdff dff_A_vLUjnDP74_0(.dout(w_dff_A_KdvZQnOx3_0),.din(w_dff_A_vLUjnDP74_0),.clk(gclk));
	jdff dff_A_HRu0UsxV7_0(.dout(w_dff_A_vLUjnDP74_0),.din(w_dff_A_HRu0UsxV7_0),.clk(gclk));
	jdff dff_A_NOTBondg0_0(.dout(w_dff_A_HRu0UsxV7_0),.din(w_dff_A_NOTBondg0_0),.clk(gclk));
	jdff dff_A_2Poa2mue9_0(.dout(w_dff_A_NOTBondg0_0),.din(w_dff_A_2Poa2mue9_0),.clk(gclk));
	jdff dff_A_Ys8MZafy6_0(.dout(w_dff_A_2Poa2mue9_0),.din(w_dff_A_Ys8MZafy6_0),.clk(gclk));
	jdff dff_A_Jf4H14860_0(.dout(w_dff_A_Ys8MZafy6_0),.din(w_dff_A_Jf4H14860_0),.clk(gclk));
	jdff dff_A_IxYExDvf8_0(.dout(w_dff_A_Jf4H14860_0),.din(w_dff_A_IxYExDvf8_0),.clk(gclk));
	jdff dff_A_WcXlRiwk9_0(.dout(w_dff_A_IxYExDvf8_0),.din(w_dff_A_WcXlRiwk9_0),.clk(gclk));
	jdff dff_A_j4eWW6fM7_0(.dout(w_dff_A_WcXlRiwk9_0),.din(w_dff_A_j4eWW6fM7_0),.clk(gclk));
	jdff dff_A_0hIR9ZAy8_0(.dout(w_G210_0[0]),.din(w_dff_A_0hIR9ZAy8_0),.clk(gclk));
	jdff dff_A_Kj646pdm1_0(.dout(w_dff_A_0hIR9ZAy8_0),.din(w_dff_A_Kj646pdm1_0),.clk(gclk));
	jdff dff_A_3vWj2P5T0_0(.dout(w_dff_A_Kj646pdm1_0),.din(w_dff_A_3vWj2P5T0_0),.clk(gclk));
	jdff dff_A_ykrmFzzJ4_0(.dout(w_dff_A_3vWj2P5T0_0),.din(w_dff_A_ykrmFzzJ4_0),.clk(gclk));
	jdff dff_A_J6uPRhhx5_0(.dout(w_dff_A_ykrmFzzJ4_0),.din(w_dff_A_J6uPRhhx5_0),.clk(gclk));
	jdff dff_A_U9Pq5whE9_0(.dout(w_dff_A_J6uPRhhx5_0),.din(w_dff_A_U9Pq5whE9_0),.clk(gclk));
	jdff dff_A_0fKSYsEz7_0(.dout(w_dff_A_U9Pq5whE9_0),.din(w_dff_A_0fKSYsEz7_0),.clk(gclk));
	jdff dff_A_gbWYWOX61_0(.dout(w_dff_A_0fKSYsEz7_0),.din(w_dff_A_gbWYWOX61_0),.clk(gclk));
	jdff dff_A_seO9mZAi9_0(.dout(w_dff_A_gbWYWOX61_0),.din(w_dff_A_seO9mZAi9_0),.clk(gclk));
	jdff dff_A_K6pOlWRz7_0(.dout(w_dff_A_seO9mZAi9_0),.din(w_dff_A_K6pOlWRz7_0),.clk(gclk));
	jdff dff_A_RPYC76iM6_0(.dout(w_dff_A_K6pOlWRz7_0),.din(w_dff_A_RPYC76iM6_0),.clk(gclk));
	jdff dff_A_X8nYf7Ib2_0(.dout(w_dff_A_RPYC76iM6_0),.din(w_dff_A_X8nYf7Ib2_0),.clk(gclk));
	jdff dff_A_WFEKeYOX3_0(.dout(w_dff_A_X8nYf7Ib2_0),.din(w_dff_A_WFEKeYOX3_0),.clk(gclk));
	jdff dff_A_gORIwm874_0(.dout(w_dff_A_WFEKeYOX3_0),.din(w_dff_A_gORIwm874_0),.clk(gclk));
	jdff dff_A_PZfsSMQf1_0(.dout(w_dff_A_gORIwm874_0),.din(w_dff_A_PZfsSMQf1_0),.clk(gclk));
	jdff dff_A_OxcboRLa7_0(.dout(w_dff_A_PZfsSMQf1_0),.din(w_dff_A_OxcboRLa7_0),.clk(gclk));
	jdff dff_A_lgVNsBUw3_1(.dout(w_G210_0[1]),.din(w_dff_A_lgVNsBUw3_1),.clk(gclk));
	jdff dff_A_2igJotMc4_0(.dout(w_G101_0[0]),.din(w_dff_A_2igJotMc4_0),.clk(gclk));
	jdff dff_A_b7ZsRcXM4_0(.dout(w_dff_A_2igJotMc4_0),.din(w_dff_A_b7ZsRcXM4_0),.clk(gclk));
	jdff dff_A_qtC2uJTM6_0(.dout(w_dff_A_b7ZsRcXM4_0),.din(w_dff_A_qtC2uJTM6_0),.clk(gclk));
	jdff dff_A_zUO6yFtc2_0(.dout(w_dff_A_qtC2uJTM6_0),.din(w_dff_A_zUO6yFtc2_0),.clk(gclk));
	jdff dff_A_XiNJVHv52_0(.dout(w_dff_A_zUO6yFtc2_0),.din(w_dff_A_XiNJVHv52_0),.clk(gclk));
	jdff dff_A_kc67abS97_0(.dout(w_dff_A_XiNJVHv52_0),.din(w_dff_A_kc67abS97_0),.clk(gclk));
	jdff dff_A_SdbcqVAH1_0(.dout(w_dff_A_kc67abS97_0),.din(w_dff_A_SdbcqVAH1_0),.clk(gclk));
	jdff dff_A_S7jz1DP98_0(.dout(w_dff_A_SdbcqVAH1_0),.din(w_dff_A_S7jz1DP98_0),.clk(gclk));
	jdff dff_A_aDnl2Ive5_0(.dout(w_dff_A_S7jz1DP98_0),.din(w_dff_A_aDnl2Ive5_0),.clk(gclk));
	jdff dff_A_C8nH7f4g9_0(.dout(w_dff_A_aDnl2Ive5_0),.din(w_dff_A_C8nH7f4g9_0),.clk(gclk));
	jdff dff_A_e09HX4jy3_0(.dout(w_dff_A_C8nH7f4g9_0),.din(w_dff_A_e09HX4jy3_0),.clk(gclk));
	jdff dff_A_XYgP6YE56_2(.dout(w_G101_0[2]),.din(w_dff_A_XYgP6YE56_2),.clk(gclk));
	jdff dff_A_hek1xz6t0_2(.dout(w_dff_A_XYgP6YE56_2),.din(w_dff_A_hek1xz6t0_2),.clk(gclk));
	jdff dff_A_0ikeNFih7_1(.dout(w_n84_0[1]),.din(w_dff_A_0ikeNFih7_1),.clk(gclk));
	jdff dff_A_Sc72a3VD2_1(.dout(w_n81_0[1]),.din(w_dff_A_Sc72a3VD2_1),.clk(gclk));
	jdff dff_A_JDwHL18b8_2(.dout(w_n81_0[2]),.din(w_dff_A_JDwHL18b8_2),.clk(gclk));
	jdff dff_A_t7DcwMMq3_2(.dout(w_G472_0[2]),.din(w_dff_A_t7DcwMMq3_2),.clk(gclk));
	jdff dff_A_uoALZ0xa1_2(.dout(w_dff_A_t7DcwMMq3_2),.din(w_dff_A_uoALZ0xa1_2),.clk(gclk));
	jdff dff_A_cLJcyHSe6_2(.dout(w_dff_A_uoALZ0xa1_2),.din(w_dff_A_cLJcyHSe6_2),.clk(gclk));
	jdff dff_A_RIZzNKuy0_2(.dout(w_dff_A_cLJcyHSe6_2),.din(w_dff_A_RIZzNKuy0_2),.clk(gclk));
	jdff dff_A_tt3a3Kk34_2(.dout(w_dff_A_RIZzNKuy0_2),.din(w_dff_A_tt3a3Kk34_2),.clk(gclk));
	jdff dff_A_lLBd2Mlm2_2(.dout(w_dff_A_tt3a3Kk34_2),.din(w_dff_A_lLBd2Mlm2_2),.clk(gclk));
	jdff dff_B_zfUoBTQh6_0(.din(n75),.dout(w_dff_B_zfUoBTQh6_0),.clk(gclk));
	jdff dff_A_vwNAnwBi9_0(.dout(w_n74_0[0]),.din(w_dff_A_vwNAnwBi9_0),.clk(gclk));
	jdff dff_A_zvGreQTX8_0(.dout(w_dff_A_vwNAnwBi9_0),.din(w_dff_A_zvGreQTX8_0),.clk(gclk));
	jdff dff_A_8Fnq0ajR2_0(.dout(w_n70_0[0]),.din(w_dff_A_8Fnq0ajR2_0),.clk(gclk));
	jdff dff_A_gWODHQOU4_0(.dout(w_dff_A_8Fnq0ajR2_0),.din(w_dff_A_gWODHQOU4_0),.clk(gclk));
	jdff dff_A_u1nqCuJj4_0(.dout(w_dff_A_gWODHQOU4_0),.din(w_dff_A_u1nqCuJj4_0),.clk(gclk));
	jdff dff_A_r5jycrNU8_0(.dout(w_dff_A_u1nqCuJj4_0),.din(w_dff_A_r5jycrNU8_0),.clk(gclk));
	jdff dff_A_B6ByFUkx9_0(.dout(w_dff_A_r5jycrNU8_0),.din(w_dff_A_B6ByFUkx9_0),.clk(gclk));
	jdff dff_A_vApP2TkF9_0(.dout(w_dff_A_B6ByFUkx9_0),.din(w_dff_A_vApP2TkF9_0),.clk(gclk));
	jdff dff_A_q2lv8LCn5_0(.dout(w_dff_A_vApP2TkF9_0),.din(w_dff_A_q2lv8LCn5_0),.clk(gclk));
	jdff dff_A_XuHVOHfK9_0(.dout(w_dff_A_q2lv8LCn5_0),.din(w_dff_A_XuHVOHfK9_0),.clk(gclk));
	jdff dff_A_3q3QRkbk6_0(.dout(w_dff_A_XuHVOHfK9_0),.din(w_dff_A_3q3QRkbk6_0),.clk(gclk));
	jdff dff_A_LQSVngut4_0(.dout(w_dff_A_3q3QRkbk6_0),.din(w_dff_A_LQSVngut4_0),.clk(gclk));
	jdff dff_A_4bB5OuEG5_0(.dout(w_dff_A_LQSVngut4_0),.din(w_dff_A_4bB5OuEG5_0),.clk(gclk));
	jdff dff_A_smsN2Iox9_0(.dout(w_dff_A_4bB5OuEG5_0),.din(w_dff_A_smsN2Iox9_0),.clk(gclk));
	jdff dff_A_HAwpuHLL6_0(.dout(w_dff_A_smsN2Iox9_0),.din(w_dff_A_HAwpuHLL6_0),.clk(gclk));
	jdff dff_B_rSPAN7jr8_0(.din(n69),.dout(w_dff_B_rSPAN7jr8_0),.clk(gclk));
	jdff dff_B_Riq3223L9_0(.din(n68),.dout(w_dff_B_Riq3223L9_0),.clk(gclk));
	jdff dff_A_w6sVhHoO8_0(.dout(w_G137_0[0]),.din(w_dff_A_w6sVhHoO8_0),.clk(gclk));
	jdff dff_A_wvDoVApv4_0(.dout(w_dff_A_w6sVhHoO8_0),.din(w_dff_A_wvDoVApv4_0),.clk(gclk));
	jdff dff_A_RWSKkCu97_0(.dout(w_dff_A_wvDoVApv4_0),.din(w_dff_A_RWSKkCu97_0),.clk(gclk));
	jdff dff_A_sGIdZOwg1_0(.dout(w_dff_A_RWSKkCu97_0),.din(w_dff_A_sGIdZOwg1_0),.clk(gclk));
	jdff dff_A_eMpst64i5_0(.dout(w_dff_A_sGIdZOwg1_0),.din(w_dff_A_eMpst64i5_0),.clk(gclk));
	jdff dff_A_uhr4LGSY7_0(.dout(w_dff_A_eMpst64i5_0),.din(w_dff_A_uhr4LGSY7_0),.clk(gclk));
	jdff dff_A_4fhJFv3b4_0(.dout(w_dff_A_uhr4LGSY7_0),.din(w_dff_A_4fhJFv3b4_0),.clk(gclk));
	jdff dff_A_MmjVKcDN1_0(.dout(w_dff_A_4fhJFv3b4_0),.din(w_dff_A_MmjVKcDN1_0),.clk(gclk));
	jdff dff_A_eqj3wAXU6_0(.dout(w_dff_A_MmjVKcDN1_0),.din(w_dff_A_eqj3wAXU6_0),.clk(gclk));
	jdff dff_A_aLnQ2UFa6_0(.dout(w_dff_A_eqj3wAXU6_0),.din(w_dff_A_aLnQ2UFa6_0),.clk(gclk));
	jdff dff_A_dmY5xswP2_0(.dout(w_dff_A_aLnQ2UFa6_0),.din(w_dff_A_dmY5xswP2_0),.clk(gclk));
	jdff dff_B_j1EcKPlT8_0(.din(n64),.dout(w_dff_B_j1EcKPlT8_0),.clk(gclk));
	jdff dff_A_5SAgPiya6_0(.dout(w_G119_0[0]),.din(w_dff_A_5SAgPiya6_0),.clk(gclk));
	jdff dff_A_g4KXJQXo9_0(.dout(w_dff_A_5SAgPiya6_0),.din(w_dff_A_g4KXJQXo9_0),.clk(gclk));
	jdff dff_A_VhUWGECe0_0(.dout(w_dff_A_g4KXJQXo9_0),.din(w_dff_A_VhUWGECe0_0),.clk(gclk));
	jdff dff_A_qL334ohz8_0(.dout(w_dff_A_VhUWGECe0_0),.din(w_dff_A_qL334ohz8_0),.clk(gclk));
	jdff dff_A_2lQI52uQ4_0(.dout(w_dff_A_qL334ohz8_0),.din(w_dff_A_2lQI52uQ4_0),.clk(gclk));
	jdff dff_A_4utpvD5Q7_0(.dout(w_dff_A_2lQI52uQ4_0),.din(w_dff_A_4utpvD5Q7_0),.clk(gclk));
	jdff dff_A_uto0gISE3_0(.dout(w_dff_A_4utpvD5Q7_0),.din(w_dff_A_uto0gISE3_0),.clk(gclk));
	jdff dff_A_lTh5TlsS4_0(.dout(w_dff_A_uto0gISE3_0),.din(w_dff_A_lTh5TlsS4_0),.clk(gclk));
	jdff dff_A_GbRVivJi6_0(.dout(w_dff_A_lTh5TlsS4_0),.din(w_dff_A_GbRVivJi6_0),.clk(gclk));
	jdff dff_A_3C7b3KkZ9_0(.dout(w_dff_A_GbRVivJi6_0),.din(w_dff_A_3C7b3KkZ9_0),.clk(gclk));
	jdff dff_A_8ccLeRGo3_0(.dout(w_dff_A_3C7b3KkZ9_0),.din(w_dff_A_8ccLeRGo3_0),.clk(gclk));
	jdff dff_A_pltr9Sy91_2(.dout(w_G119_0[2]),.din(w_dff_A_pltr9Sy91_2),.clk(gclk));
	jdff dff_A_KAFUf0ie5_0(.dout(w_G110_0[0]),.din(w_dff_A_KAFUf0ie5_0),.clk(gclk));
	jdff dff_A_bMLvj4vK6_0(.dout(w_dff_A_KAFUf0ie5_0),.din(w_dff_A_bMLvj4vK6_0),.clk(gclk));
	jdff dff_A_isC4nyop5_0(.dout(w_dff_A_bMLvj4vK6_0),.din(w_dff_A_isC4nyop5_0),.clk(gclk));
	jdff dff_A_1OCK4Hfe3_0(.dout(w_dff_A_isC4nyop5_0),.din(w_dff_A_1OCK4Hfe3_0),.clk(gclk));
	jdff dff_A_FpjEbNeu5_0(.dout(w_dff_A_1OCK4Hfe3_0),.din(w_dff_A_FpjEbNeu5_0),.clk(gclk));
	jdff dff_A_w6UiwGWK1_0(.dout(w_dff_A_FpjEbNeu5_0),.din(w_dff_A_w6UiwGWK1_0),.clk(gclk));
	jdff dff_A_UDv47Jyb2_0(.dout(w_dff_A_w6UiwGWK1_0),.din(w_dff_A_UDv47Jyb2_0),.clk(gclk));
	jdff dff_A_tMBLsMwz9_0(.dout(w_dff_A_UDv47Jyb2_0),.din(w_dff_A_tMBLsMwz9_0),.clk(gclk));
	jdff dff_A_HcNUUNC09_0(.dout(w_dff_A_tMBLsMwz9_0),.din(w_dff_A_HcNUUNC09_0),.clk(gclk));
	jdff dff_A_a9np6C7j6_0(.dout(w_dff_A_HcNUUNC09_0),.din(w_dff_A_a9np6C7j6_0),.clk(gclk));
	jdff dff_A_iU37nXPr2_0(.dout(w_dff_A_a9np6C7j6_0),.din(w_dff_A_iU37nXPr2_0),.clk(gclk));
	jdff dff_B_lRv8V3uU9_1(.din(n59),.dout(w_dff_B_lRv8V3uU9_1),.clk(gclk));
	jdff dff_A_CqMkEHCF9_0(.dout(w_G234_1[0]),.din(w_dff_A_CqMkEHCF9_0),.clk(gclk));
	jdff dff_A_bCHLZywt4_0(.dout(w_G221_0[0]),.din(w_dff_A_bCHLZywt4_0),.clk(gclk));
	jdff dff_A_Xm3AFnP14_0(.dout(w_dff_A_bCHLZywt4_0),.din(w_dff_A_Xm3AFnP14_0),.clk(gclk));
	jdff dff_A_ramVYyqn5_0(.dout(w_dff_A_Xm3AFnP14_0),.din(w_dff_A_ramVYyqn5_0),.clk(gclk));
	jdff dff_A_JpljhAPX5_0(.dout(w_n58_2[0]),.din(w_dff_A_JpljhAPX5_0),.clk(gclk));
	jdff dff_A_oaRh1Isg0_0(.dout(w_dff_A_JpljhAPX5_0),.din(w_dff_A_oaRh1Isg0_0),.clk(gclk));
	jdff dff_A_EWEC3qSB8_0(.dout(w_dff_A_oaRh1Isg0_0),.din(w_dff_A_EWEC3qSB8_0),.clk(gclk));
	jdff dff_A_vajKnaec8_0(.dout(w_dff_A_EWEC3qSB8_0),.din(w_dff_A_vajKnaec8_0),.clk(gclk));
	jdff dff_A_gNVfRazD7_2(.dout(w_n58_2[2]),.din(w_dff_A_gNVfRazD7_2),.clk(gclk));
	jdff dff_A_VLPQj9N95_2(.dout(w_dff_A_gNVfRazD7_2),.din(w_dff_A_VLPQj9N95_2),.clk(gclk));
	jdff dff_A_jjicVHTu2_2(.dout(w_dff_A_VLPQj9N95_2),.din(w_dff_A_jjicVHTu2_2),.clk(gclk));
	jdff dff_A_S5z7eyd04_2(.dout(w_dff_A_jjicVHTu2_2),.din(w_dff_A_S5z7eyd04_2),.clk(gclk));
	jdff dff_A_HtXn5sey4_0(.dout(w_n131_0[0]),.din(w_dff_A_HtXn5sey4_0),.clk(gclk));
	jdff dff_A_mGkVDPT69_0(.dout(w_dff_A_HtXn5sey4_0),.din(w_dff_A_mGkVDPT69_0),.clk(gclk));
	jdff dff_A_Rkt191pb6_0(.dout(w_dff_A_mGkVDPT69_0),.din(w_dff_A_Rkt191pb6_0),.clk(gclk));
	jdff dff_A_a3stNVrJ1_2(.dout(w_n131_0[2]),.din(w_dff_A_a3stNVrJ1_2),.clk(gclk));
	jdff dff_A_howrrxnu0_2(.dout(w_dff_A_a3stNVrJ1_2),.din(w_dff_A_howrrxnu0_2),.clk(gclk));
	jdff dff_A_Xxkx8BNO7_2(.dout(w_dff_A_howrrxnu0_2),.din(w_dff_A_Xxkx8BNO7_2),.clk(gclk));
	jdff dff_A_kUpEp3qm3_2(.dout(w_dff_A_Xxkx8BNO7_2),.din(w_dff_A_kUpEp3qm3_2),.clk(gclk));
	jdff dff_A_66Ajoyz44_2(.dout(w_dff_A_kUpEp3qm3_2),.din(w_dff_A_66Ajoyz44_2),.clk(gclk));
	jdff dff_A_MBSKY7wZ0_1(.dout(w_n130_0[1]),.din(w_dff_A_MBSKY7wZ0_1),.clk(gclk));
	jdff dff_A_wymmlnrp4_1(.dout(w_dff_A_MBSKY7wZ0_1),.din(w_dff_A_wymmlnrp4_1),.clk(gclk));
	jdff dff_A_dBSwxGuH5_1(.dout(w_dff_A_wymmlnrp4_1),.din(w_dff_A_dBSwxGuH5_1),.clk(gclk));
	jdff dff_A_2Owppcnm8_1(.dout(w_dff_A_dBSwxGuH5_1),.din(w_dff_A_2Owppcnm8_1),.clk(gclk));
	jdff dff_A_IdGG1rts0_2(.dout(w_n130_0[2]),.din(w_dff_A_IdGG1rts0_2),.clk(gclk));
	jdff dff_A_n5rbimli5_2(.dout(w_dff_A_IdGG1rts0_2),.din(w_dff_A_n5rbimli5_2),.clk(gclk));
	jdff dff_A_UjNvUUNS2_2(.dout(w_dff_A_n5rbimli5_2),.din(w_dff_A_UjNvUUNS2_2),.clk(gclk));
	jdff dff_A_zRemNt128_2(.dout(w_dff_A_UjNvUUNS2_2),.din(w_dff_A_zRemNt128_2),.clk(gclk));
	jdff dff_A_2aGJKbXC9_2(.dout(w_dff_A_zRemNt128_2),.din(w_dff_A_2aGJKbXC9_2),.clk(gclk));
	jdff dff_A_2Rq2Fr4M0_2(.dout(w_dff_A_2aGJKbXC9_2),.din(w_dff_A_2Rq2Fr4M0_2),.clk(gclk));
	jdff dff_A_itdnHQhG9_2(.dout(w_dff_A_2Rq2Fr4M0_2),.din(w_dff_A_itdnHQhG9_2),.clk(gclk));
	jdff dff_A_Glw0nwvI2_2(.dout(w_dff_A_itdnHQhG9_2),.din(w_dff_A_Glw0nwvI2_2),.clk(gclk));
	jdff dff_A_rcqTukSG5_2(.dout(w_dff_A_Glw0nwvI2_2),.din(w_dff_A_rcqTukSG5_2),.clk(gclk));
	jdff dff_A_5djuqVFR4_0(.dout(w_n124_0[0]),.din(w_dff_A_5djuqVFR4_0),.clk(gclk));
	jdff dff_A_0sMTgjXs1_1(.dout(w_G898_0[1]),.din(w_dff_A_0sMTgjXs1_1),.clk(gclk));
	jdff dff_A_ydXUKeDR6_0(.dout(w_n186_0[0]),.din(w_dff_A_ydXUKeDR6_0),.clk(gclk));
	jdff dff_A_BinbQrpY8_0(.dout(w_dff_A_ydXUKeDR6_0),.din(w_dff_A_BinbQrpY8_0),.clk(gclk));
	jdff dff_A_sB64z77S3_0(.dout(w_dff_A_BinbQrpY8_0),.din(w_dff_A_sB64z77S3_0),.clk(gclk));
	jdff dff_A_jX8b1f1s6_1(.dout(w_n151_0[1]),.din(w_dff_A_jX8b1f1s6_1),.clk(gclk));
	jdff dff_A_Ba13vm6k1_1(.dout(w_dff_A_jX8b1f1s6_1),.din(w_dff_A_Ba13vm6k1_1),.clk(gclk));
	jdff dff_A_WObRkVXM3_1(.dout(w_dff_A_Ba13vm6k1_1),.din(w_dff_A_WObRkVXM3_1),.clk(gclk));
	jdff dff_A_Lj6B4xWL1_1(.dout(w_dff_A_WObRkVXM3_1),.din(w_dff_A_Lj6B4xWL1_1),.clk(gclk));
	jdff dff_A_4rPayeat6_1(.dout(w_dff_A_Lj6B4xWL1_1),.din(w_dff_A_4rPayeat6_1),.clk(gclk));
	jdff dff_A_4kxpTksh5_1(.dout(w_dff_A_4rPayeat6_1),.din(w_dff_A_4kxpTksh5_1),.clk(gclk));
	jdff dff_A_OzW7DTnm7_1(.dout(w_dff_A_4kxpTksh5_1),.din(w_dff_A_OzW7DTnm7_1),.clk(gclk));
	jdff dff_A_Urd1DreW0_1(.dout(w_dff_A_OzW7DTnm7_1),.din(w_dff_A_Urd1DreW0_1),.clk(gclk));
	jdff dff_A_CLhc1APU4_1(.dout(w_dff_A_Urd1DreW0_1),.din(w_dff_A_CLhc1APU4_1),.clk(gclk));
	jdff dff_A_PzMxH0kn3_1(.dout(w_dff_A_CLhc1APU4_1),.din(w_dff_A_PzMxH0kn3_1),.clk(gclk));
	jdff dff_A_gjLME5Nz6_1(.dout(w_dff_A_PzMxH0kn3_1),.din(w_dff_A_gjLME5Nz6_1),.clk(gclk));
	jdff dff_A_5z0D4Avc7_1(.dout(w_dff_A_gjLME5Nz6_1),.din(w_dff_A_5z0D4Avc7_1),.clk(gclk));
	jdff dff_B_WXB1PzWk1_1(.din(n144),.dout(w_dff_B_WXB1PzWk1_1),.clk(gclk));
	jdff dff_B_OR4AFcGl9_1(.din(w_dff_B_WXB1PzWk1_1),.dout(w_dff_B_OR4AFcGl9_1),.clk(gclk));
	jdff dff_A_ny44Yxjq1_0(.dout(w_G131_0[0]),.din(w_dff_A_ny44Yxjq1_0),.clk(gclk));
	jdff dff_A_t6Aqb92A9_0(.dout(w_dff_A_ny44Yxjq1_0),.din(w_dff_A_t6Aqb92A9_0),.clk(gclk));
	jdff dff_A_gmemrK8c4_0(.dout(w_dff_A_t6Aqb92A9_0),.din(w_dff_A_gmemrK8c4_0),.clk(gclk));
	jdff dff_A_MxtWWakH8_0(.dout(w_dff_A_gmemrK8c4_0),.din(w_dff_A_MxtWWakH8_0),.clk(gclk));
	jdff dff_A_sp8c4X9D8_0(.dout(w_dff_A_MxtWWakH8_0),.din(w_dff_A_sp8c4X9D8_0),.clk(gclk));
	jdff dff_A_ZD9dmgdA5_0(.dout(w_dff_A_sp8c4X9D8_0),.din(w_dff_A_ZD9dmgdA5_0),.clk(gclk));
	jdff dff_A_N7knh9kF0_0(.dout(w_dff_A_ZD9dmgdA5_0),.din(w_dff_A_N7knh9kF0_0),.clk(gclk));
	jdff dff_A_DnZ0gSkA9_0(.dout(w_dff_A_N7knh9kF0_0),.din(w_dff_A_DnZ0gSkA9_0),.clk(gclk));
	jdff dff_A_aikiDzSt6_0(.dout(w_dff_A_DnZ0gSkA9_0),.din(w_dff_A_aikiDzSt6_0),.clk(gclk));
	jdff dff_A_bCg3G5HH0_0(.dout(w_dff_A_aikiDzSt6_0),.din(w_dff_A_bCg3G5HH0_0),.clk(gclk));
	jdff dff_A_kods908k3_0(.dout(w_dff_A_bCg3G5HH0_0),.din(w_dff_A_kods908k3_0),.clk(gclk));
	jdff dff_A_yHCBM2o71_2(.dout(w_G131_0[2]),.din(w_dff_A_yHCBM2o71_2),.clk(gclk));
	jdff dff_A_4gro4Qq16_1(.dout(w_G953_2[1]),.din(w_dff_A_4gro4Qq16_1),.clk(gclk));
	jdff dff_A_MndoQkpc4_1(.dout(w_G214_0[1]),.din(w_dff_A_MndoQkpc4_1),.clk(gclk));
	jdff dff_A_O82f2qgK5_0(.dout(w_n67_0[0]),.din(w_dff_A_O82f2qgK5_0),.clk(gclk));
	jdff dff_A_9hXodets6_0(.dout(w_n66_0[0]),.din(w_dff_A_9hXodets6_0),.clk(gclk));
	jdff dff_A_IzmLdrPM4_0(.dout(w_dff_A_9hXodets6_0),.din(w_dff_A_IzmLdrPM4_0),.clk(gclk));
	jdff dff_A_s9eyQzU52_0(.dout(w_G140_0[0]),.din(w_dff_A_s9eyQzU52_0),.clk(gclk));
	jdff dff_A_ijYW7ftR5_0(.dout(w_dff_A_s9eyQzU52_0),.din(w_dff_A_ijYW7ftR5_0),.clk(gclk));
	jdff dff_A_nStjOTmZ5_0(.dout(w_dff_A_ijYW7ftR5_0),.din(w_dff_A_nStjOTmZ5_0),.clk(gclk));
	jdff dff_A_oaq1eUE38_0(.dout(w_dff_A_nStjOTmZ5_0),.din(w_dff_A_oaq1eUE38_0),.clk(gclk));
	jdff dff_A_g1TcIJRt4_0(.dout(w_dff_A_oaq1eUE38_0),.din(w_dff_A_g1TcIJRt4_0),.clk(gclk));
	jdff dff_A_7LILtQ9H7_0(.dout(w_dff_A_g1TcIJRt4_0),.din(w_dff_A_7LILtQ9H7_0),.clk(gclk));
	jdff dff_A_LA6PbRAi6_0(.dout(w_dff_A_7LILtQ9H7_0),.din(w_dff_A_LA6PbRAi6_0),.clk(gclk));
	jdff dff_A_tHxKLm443_0(.dout(w_dff_A_LA6PbRAi6_0),.din(w_dff_A_tHxKLm443_0),.clk(gclk));
	jdff dff_A_ZiHncPfI6_0(.dout(w_dff_A_tHxKLm443_0),.din(w_dff_A_ZiHncPfI6_0),.clk(gclk));
	jdff dff_A_ej3pzEcr5_0(.dout(w_dff_A_ZiHncPfI6_0),.din(w_dff_A_ej3pzEcr5_0),.clk(gclk));
	jdff dff_A_SXTVyYmQ3_0(.dout(w_dff_A_ej3pzEcr5_0),.din(w_dff_A_SXTVyYmQ3_0),.clk(gclk));
	jdff dff_A_wF4hsBQF2_1(.dout(w_G140_0[1]),.din(w_dff_A_wF4hsBQF2_1),.clk(gclk));
	jdff dff_A_i1Hwubp30_0(.dout(w_G125_0[0]),.din(w_dff_A_i1Hwubp30_0),.clk(gclk));
	jdff dff_A_aAnerfct9_0(.dout(w_dff_A_i1Hwubp30_0),.din(w_dff_A_aAnerfct9_0),.clk(gclk));
	jdff dff_A_PAoRkGDN0_0(.dout(w_dff_A_aAnerfct9_0),.din(w_dff_A_PAoRkGDN0_0),.clk(gclk));
	jdff dff_A_Clgrptpj1_0(.dout(w_dff_A_PAoRkGDN0_0),.din(w_dff_A_Clgrptpj1_0),.clk(gclk));
	jdff dff_A_v6chAHij5_0(.dout(w_dff_A_Clgrptpj1_0),.din(w_dff_A_v6chAHij5_0),.clk(gclk));
	jdff dff_A_GcOqCF9K8_0(.dout(w_dff_A_v6chAHij5_0),.din(w_dff_A_GcOqCF9K8_0),.clk(gclk));
	jdff dff_A_Nyy2vzIP0_0(.dout(w_dff_A_GcOqCF9K8_0),.din(w_dff_A_Nyy2vzIP0_0),.clk(gclk));
	jdff dff_A_O6B0a1403_0(.dout(w_dff_A_Nyy2vzIP0_0),.din(w_dff_A_O6B0a1403_0),.clk(gclk));
	jdff dff_A_SeSyZGcX5_0(.dout(w_dff_A_O6B0a1403_0),.din(w_dff_A_SeSyZGcX5_0),.clk(gclk));
	jdff dff_A_iijTPlN86_0(.dout(w_dff_A_SeSyZGcX5_0),.din(w_dff_A_iijTPlN86_0),.clk(gclk));
	jdff dff_A_C8994UPm7_0(.dout(w_dff_A_iijTPlN86_0),.din(w_dff_A_C8994UPm7_0),.clk(gclk));
	jdff dff_A_rlIJPHfN1_1(.dout(w_G125_0[1]),.din(w_dff_A_rlIJPHfN1_1),.clk(gclk));
	jdff dff_A_WndBmvHt3_1(.dout(w_dff_A_rlIJPHfN1_1),.din(w_dff_A_WndBmvHt3_1),.clk(gclk));
	jdff dff_A_ARiPaSY28_0(.dout(w_G146_0[0]),.din(w_dff_A_ARiPaSY28_0),.clk(gclk));
	jdff dff_A_paWH26mO8_0(.dout(w_dff_A_ARiPaSY28_0),.din(w_dff_A_paWH26mO8_0),.clk(gclk));
	jdff dff_A_oWK3JBLm4_0(.dout(w_dff_A_paWH26mO8_0),.din(w_dff_A_oWK3JBLm4_0),.clk(gclk));
	jdff dff_A_ANKfPbG39_0(.dout(w_dff_A_oWK3JBLm4_0),.din(w_dff_A_ANKfPbG39_0),.clk(gclk));
	jdff dff_A_Z1iiLFEb2_0(.dout(w_dff_A_ANKfPbG39_0),.din(w_dff_A_Z1iiLFEb2_0),.clk(gclk));
	jdff dff_A_0FPz1Bmz4_0(.dout(w_dff_A_Z1iiLFEb2_0),.din(w_dff_A_0FPz1Bmz4_0),.clk(gclk));
	jdff dff_A_t7erJs8e7_0(.dout(w_dff_A_0FPz1Bmz4_0),.din(w_dff_A_t7erJs8e7_0),.clk(gclk));
	jdff dff_A_b0unMr1B5_0(.dout(w_dff_A_t7erJs8e7_0),.din(w_dff_A_b0unMr1B5_0),.clk(gclk));
	jdff dff_A_QBTBEDr06_0(.dout(w_dff_A_b0unMr1B5_0),.din(w_dff_A_QBTBEDr06_0),.clk(gclk));
	jdff dff_A_lGqwmx6k0_0(.dout(w_dff_A_QBTBEDr06_0),.din(w_dff_A_lGqwmx6k0_0),.clk(gclk));
	jdff dff_B_pJ00iYd30_3(.din(G146),.dout(w_dff_B_pJ00iYd30_3),.clk(gclk));
	jdff dff_A_2LDcOgv21_0(.dout(w_G113_0[0]),.din(w_dff_A_2LDcOgv21_0),.clk(gclk));
	jdff dff_A_gh9SyJsA6_0(.dout(w_dff_A_2LDcOgv21_0),.din(w_dff_A_gh9SyJsA6_0),.clk(gclk));
	jdff dff_A_m86lGQxw3_0(.dout(w_dff_A_gh9SyJsA6_0),.din(w_dff_A_m86lGQxw3_0),.clk(gclk));
	jdff dff_A_W2V6DUtM6_0(.dout(w_dff_A_m86lGQxw3_0),.din(w_dff_A_W2V6DUtM6_0),.clk(gclk));
	jdff dff_A_WbCUFWBT6_0(.dout(w_dff_A_W2V6DUtM6_0),.din(w_dff_A_WbCUFWBT6_0),.clk(gclk));
	jdff dff_A_HM7cNEzm5_0(.dout(w_dff_A_WbCUFWBT6_0),.din(w_dff_A_HM7cNEzm5_0),.clk(gclk));
	jdff dff_A_LfoBj8Ja6_0(.dout(w_dff_A_HM7cNEzm5_0),.din(w_dff_A_LfoBj8Ja6_0),.clk(gclk));
	jdff dff_A_vnKd2LCA2_0(.dout(w_dff_A_LfoBj8Ja6_0),.din(w_dff_A_vnKd2LCA2_0),.clk(gclk));
	jdff dff_A_joXP8Esh0_0(.dout(w_dff_A_vnKd2LCA2_0),.din(w_dff_A_joXP8Esh0_0),.clk(gclk));
	jdff dff_A_rPloaFkw3_0(.dout(w_dff_A_joXP8Esh0_0),.din(w_dff_A_rPloaFkw3_0),.clk(gclk));
	jdff dff_A_W6A9ZwZM7_0(.dout(w_dff_A_rPloaFkw3_0),.din(w_dff_A_W6A9ZwZM7_0),.clk(gclk));
	jdff dff_A_Mv9PS05C3_0(.dout(w_G104_0[0]),.din(w_dff_A_Mv9PS05C3_0),.clk(gclk));
	jdff dff_A_6NzcPmKd8_0(.dout(w_dff_A_Mv9PS05C3_0),.din(w_dff_A_6NzcPmKd8_0),.clk(gclk));
	jdff dff_A_oF6pixnn9_0(.dout(w_dff_A_6NzcPmKd8_0),.din(w_dff_A_oF6pixnn9_0),.clk(gclk));
	jdff dff_A_OepuZN8N2_0(.dout(w_dff_A_oF6pixnn9_0),.din(w_dff_A_OepuZN8N2_0),.clk(gclk));
	jdff dff_A_GoTNuIH95_0(.dout(w_dff_A_OepuZN8N2_0),.din(w_dff_A_GoTNuIH95_0),.clk(gclk));
	jdff dff_A_48hznqgR6_0(.dout(w_dff_A_GoTNuIH95_0),.din(w_dff_A_48hznqgR6_0),.clk(gclk));
	jdff dff_A_hOBl3brz2_0(.dout(w_dff_A_48hznqgR6_0),.din(w_dff_A_hOBl3brz2_0),.clk(gclk));
	jdff dff_A_vR3vijAC3_0(.dout(w_dff_A_hOBl3brz2_0),.din(w_dff_A_vR3vijAC3_0),.clk(gclk));
	jdff dff_A_JGwUCmuH4_0(.dout(w_dff_A_vR3vijAC3_0),.din(w_dff_A_JGwUCmuH4_0),.clk(gclk));
	jdff dff_A_k0YkS6im8_0(.dout(w_dff_A_JGwUCmuH4_0),.din(w_dff_A_k0YkS6im8_0),.clk(gclk));
	jdff dff_A_XBXSzFWV5_0(.dout(w_dff_A_k0YkS6im8_0),.din(w_dff_A_XBXSzFWV5_0),.clk(gclk));
	jdff dff_A_mfxrm3Sh9_1(.dout(w_G104_0[1]),.din(w_dff_A_mfxrm3Sh9_1),.clk(gclk));
	jdff dff_A_GcLArIWj5_1(.dout(w_G475_0[1]),.din(w_dff_A_GcLArIWj5_1),.clk(gclk));
	jdff dff_A_AOQreN4t6_1(.dout(w_dff_A_GcLArIWj5_1),.din(w_dff_A_AOQreN4t6_1),.clk(gclk));
	jdff dff_A_GY65gK7N7_1(.dout(w_dff_A_AOQreN4t6_1),.din(w_dff_A_GY65gK7N7_1),.clk(gclk));
	jdff dff_A_ViEKZQb18_1(.dout(w_dff_A_GY65gK7N7_1),.din(w_dff_A_ViEKZQb18_1),.clk(gclk));
	jdff dff_A_YleF7ISi4_1(.dout(w_dff_A_ViEKZQb18_1),.din(w_dff_A_YleF7ISi4_1),.clk(gclk));
	jdff dff_A_YB1Nc0QZ0_1(.dout(w_dff_A_YleF7ISi4_1),.din(w_dff_A_YB1Nc0QZ0_1),.clk(gclk));
	jdff dff_A_mWR2PQIy1_0(.dout(w_n139_0[0]),.din(w_dff_A_mWR2PQIy1_0),.clk(gclk));
	jdff dff_A_VA5asiY78_0(.dout(w_dff_A_mWR2PQIy1_0),.din(w_dff_A_VA5asiY78_0),.clk(gclk));
	jdff dff_A_4KNi1YVI9_0(.dout(w_dff_A_VA5asiY78_0),.din(w_dff_A_4KNi1YVI9_0),.clk(gclk));
	jdff dff_A_K63yS8ea1_0(.dout(w_dff_A_4KNi1YVI9_0),.din(w_dff_A_K63yS8ea1_0),.clk(gclk));
	jdff dff_A_XWmNXPPX1_0(.dout(w_dff_A_K63yS8ea1_0),.din(w_dff_A_XWmNXPPX1_0),.clk(gclk));
	jdff dff_A_IACZD6388_0(.dout(w_dff_A_XWmNXPPX1_0),.din(w_dff_A_IACZD6388_0),.clk(gclk));
	jdff dff_A_GPJKNxuc2_0(.dout(w_dff_A_IACZD6388_0),.din(w_dff_A_GPJKNxuc2_0),.clk(gclk));
	jdff dff_A_A6t5laxm8_0(.dout(w_dff_A_GPJKNxuc2_0),.din(w_dff_A_A6t5laxm8_0),.clk(gclk));
	jdff dff_A_DaKDpKmx2_0(.dout(w_dff_A_A6t5laxm8_0),.din(w_dff_A_DaKDpKmx2_0),.clk(gclk));
	jdff dff_A_JOsJ6Rhk9_0(.dout(w_dff_A_DaKDpKmx2_0),.din(w_dff_A_JOsJ6Rhk9_0),.clk(gclk));
	jdff dff_A_KtTzOYmK8_0(.dout(w_dff_A_JOsJ6Rhk9_0),.din(w_dff_A_KtTzOYmK8_0),.clk(gclk));
	jdff dff_A_pyKFEhQI8_0(.dout(w_dff_A_KtTzOYmK8_0),.din(w_dff_A_pyKFEhQI8_0),.clk(gclk));
	jdff dff_A_KdXWk3gy3_0(.dout(w_dff_A_pyKFEhQI8_0),.din(w_dff_A_KdXWk3gy3_0),.clk(gclk));
	jdff dff_B_Bh3sPweE9_1(.din(n133),.dout(w_dff_B_Bh3sPweE9_1),.clk(gclk));
	jdff dff_B_UKEKbcmb4_1(.din(w_dff_B_Bh3sPweE9_1),.dout(w_dff_B_UKEKbcmb4_1),.clk(gclk));
	jdff dff_B_idvopbrR7_0(.din(n137),.dout(w_dff_B_idvopbrR7_0),.clk(gclk));
	jdff dff_A_lFvFyPPR1_1(.dout(w_G122_0[1]),.din(w_dff_A_lFvFyPPR1_1),.clk(gclk));
	jdff dff_A_94f2hsQR2_1(.dout(w_dff_A_lFvFyPPR1_1),.din(w_dff_A_94f2hsQR2_1),.clk(gclk));
	jdff dff_A_xSqjmXpx4_1(.dout(w_dff_A_94f2hsQR2_1),.din(w_dff_A_xSqjmXpx4_1),.clk(gclk));
	jdff dff_A_j74IhGhE7_1(.dout(w_dff_A_xSqjmXpx4_1),.din(w_dff_A_j74IhGhE7_1),.clk(gclk));
	jdff dff_A_7kYhQ0L47_1(.dout(w_dff_A_j74IhGhE7_1),.din(w_dff_A_7kYhQ0L47_1),.clk(gclk));
	jdff dff_A_ACEK8Yt05_1(.dout(w_dff_A_7kYhQ0L47_1),.din(w_dff_A_ACEK8Yt05_1),.clk(gclk));
	jdff dff_A_4UCi0tU26_1(.dout(w_dff_A_ACEK8Yt05_1),.din(w_dff_A_4UCi0tU26_1),.clk(gclk));
	jdff dff_A_zKzwhAVR1_1(.dout(w_dff_A_4UCi0tU26_1),.din(w_dff_A_zKzwhAVR1_1),.clk(gclk));
	jdff dff_A_zdaY5l260_1(.dout(w_dff_A_zKzwhAVR1_1),.din(w_dff_A_zdaY5l260_1),.clk(gclk));
	jdff dff_A_NGqv4ogJ5_1(.dout(w_dff_A_zdaY5l260_1),.din(w_dff_A_NGqv4ogJ5_1),.clk(gclk));
	jdff dff_A_FcIi9Brt1_1(.dout(w_dff_A_NGqv4ogJ5_1),.din(w_dff_A_FcIi9Brt1_1),.clk(gclk));
	jdff dff_A_zeEAMW488_1(.dout(w_dff_A_FcIi9Brt1_1),.din(w_dff_A_zeEAMW488_1),.clk(gclk));
	jdff dff_A_TJajhCmD7_0(.dout(w_G116_0[0]),.din(w_dff_A_TJajhCmD7_0),.clk(gclk));
	jdff dff_A_CdrawaRy0_0(.dout(w_dff_A_TJajhCmD7_0),.din(w_dff_A_CdrawaRy0_0),.clk(gclk));
	jdff dff_A_C71pwByx9_0(.dout(w_dff_A_CdrawaRy0_0),.din(w_dff_A_C71pwByx9_0),.clk(gclk));
	jdff dff_A_KBo7VCKl8_0(.dout(w_dff_A_C71pwByx9_0),.din(w_dff_A_KBo7VCKl8_0),.clk(gclk));
	jdff dff_A_eUXjmOwR6_0(.dout(w_dff_A_KBo7VCKl8_0),.din(w_dff_A_eUXjmOwR6_0),.clk(gclk));
	jdff dff_A_tYURWBIx1_0(.dout(w_dff_A_eUXjmOwR6_0),.din(w_dff_A_tYURWBIx1_0),.clk(gclk));
	jdff dff_A_1krbR3pj6_0(.dout(w_dff_A_tYURWBIx1_0),.din(w_dff_A_1krbR3pj6_0),.clk(gclk));
	jdff dff_A_lW37oSFs1_0(.dout(w_dff_A_1krbR3pj6_0),.din(w_dff_A_lW37oSFs1_0),.clk(gclk));
	jdff dff_A_q7vpDMdE7_0(.dout(w_dff_A_lW37oSFs1_0),.din(w_dff_A_q7vpDMdE7_0),.clk(gclk));
	jdff dff_A_D3wF8aWo3_0(.dout(w_dff_A_q7vpDMdE7_0),.din(w_dff_A_D3wF8aWo3_0),.clk(gclk));
	jdff dff_A_hpithpsj5_0(.dout(w_dff_A_D3wF8aWo3_0),.din(w_dff_A_hpithpsj5_0),.clk(gclk));
	jdff dff_A_Jw8eBKCr2_0(.dout(w_G107_0[0]),.din(w_dff_A_Jw8eBKCr2_0),.clk(gclk));
	jdff dff_A_uNHBq4bp3_0(.dout(w_dff_A_Jw8eBKCr2_0),.din(w_dff_A_uNHBq4bp3_0),.clk(gclk));
	jdff dff_A_vPwzDTcv7_0(.dout(w_dff_A_uNHBq4bp3_0),.din(w_dff_A_vPwzDTcv7_0),.clk(gclk));
	jdff dff_A_PYdrpQmU8_0(.dout(w_dff_A_vPwzDTcv7_0),.din(w_dff_A_PYdrpQmU8_0),.clk(gclk));
	jdff dff_A_pWbL2WTr1_0(.dout(w_dff_A_PYdrpQmU8_0),.din(w_dff_A_pWbL2WTr1_0),.clk(gclk));
	jdff dff_A_fwFKgR1q5_0(.dout(w_dff_A_pWbL2WTr1_0),.din(w_dff_A_fwFKgR1q5_0),.clk(gclk));
	jdff dff_A_2FkRzDyw3_0(.dout(w_dff_A_fwFKgR1q5_0),.din(w_dff_A_2FkRzDyw3_0),.clk(gclk));
	jdff dff_A_nwUITX0C1_0(.dout(w_dff_A_2FkRzDyw3_0),.din(w_dff_A_nwUITX0C1_0),.clk(gclk));
	jdff dff_A_ID4Pk6ml7_0(.dout(w_dff_A_nwUITX0C1_0),.din(w_dff_A_ID4Pk6ml7_0),.clk(gclk));
	jdff dff_A_jahA2CPO7_0(.dout(w_dff_A_ID4Pk6ml7_0),.din(w_dff_A_jahA2CPO7_0),.clk(gclk));
	jdff dff_A_tILj3M467_0(.dout(w_dff_A_jahA2CPO7_0),.din(w_dff_A_tILj3M467_0),.clk(gclk));
	jdff dff_A_TWcZ3hlV8_1(.dout(w_G107_0[1]),.din(w_dff_A_TWcZ3hlV8_1),.clk(gclk));
	jdff dff_A_vqQHzyQy5_2(.dout(w_n103_2[2]),.din(w_dff_A_vqQHzyQy5_2),.clk(gclk));
	jdff dff_A_sCiPDOfo6_2(.dout(w_dff_A_vqQHzyQy5_2),.din(w_dff_A_sCiPDOfo6_2),.clk(gclk));
	jdff dff_A_e1THIr3i3_1(.dout(w_G234_0[1]),.din(w_dff_A_e1THIr3i3_1),.clk(gclk));
	jdff dff_A_h6dGnH6u5_0(.dout(w_G217_0[0]),.din(w_dff_A_h6dGnH6u5_0),.clk(gclk));
	jdff dff_A_SU1pPER50_0(.dout(w_dff_A_h6dGnH6u5_0),.din(w_dff_A_SU1pPER50_0),.clk(gclk));
	jdff dff_A_Fk427TdG1_0(.dout(w_dff_A_SU1pPER50_0),.din(w_dff_A_Fk427TdG1_0),.clk(gclk));
	jdff dff_A_x7rPlRLu2_0(.dout(w_dff_A_Fk427TdG1_0),.din(w_dff_A_x7rPlRLu2_0),.clk(gclk));
	jdff dff_A_fXlHFcYu6_0(.dout(w_dff_A_x7rPlRLu2_0),.din(w_dff_A_fXlHFcYu6_0),.clk(gclk));
	jdff dff_A_9W0pmyp47_0(.dout(w_dff_A_fXlHFcYu6_0),.din(w_dff_A_9W0pmyp47_0),.clk(gclk));
	jdff dff_A_zxqiynyj6_0(.dout(w_dff_A_9W0pmyp47_0),.din(w_dff_A_zxqiynyj6_0),.clk(gclk));
	jdff dff_A_mDgN9ZgF7_0(.dout(w_dff_A_zxqiynyj6_0),.din(w_dff_A_mDgN9ZgF7_0),.clk(gclk));
	jdff dff_A_kL1Z1Pm95_0(.dout(w_dff_A_mDgN9ZgF7_0),.din(w_dff_A_kL1Z1Pm95_0),.clk(gclk));
	jdff dff_A_kV9f1zVT7_0(.dout(w_dff_A_kL1Z1Pm95_0),.din(w_dff_A_kV9f1zVT7_0),.clk(gclk));
	jdff dff_A_qJlt3UJN2_0(.dout(w_dff_A_kV9f1zVT7_0),.din(w_dff_A_qJlt3UJN2_0),.clk(gclk));
	jdff dff_A_7ka7thog0_0(.dout(w_dff_A_qJlt3UJN2_0),.din(w_dff_A_7ka7thog0_0),.clk(gclk));
	jdff dff_A_2bIecY3Y3_0(.dout(w_dff_A_7ka7thog0_0),.din(w_dff_A_2bIecY3Y3_0),.clk(gclk));
	jdff dff_A_YFHk7fnc7_0(.dout(w_dff_A_2bIecY3Y3_0),.din(w_dff_A_YFHk7fnc7_0),.clk(gclk));
	jdff dff_A_Ej80MD9W3_2(.dout(w_G217_0[2]),.din(w_dff_A_Ej80MD9W3_2),.clk(gclk));
	jdff dff_B_hO9y6Zfl1_3(.din(G217),.dout(w_dff_B_hO9y6Zfl1_3),.clk(gclk));
	jdff dff_B_NMvSU6qi8_3(.din(w_dff_B_hO9y6Zfl1_3),.dout(w_dff_B_NMvSU6qi8_3),.clk(gclk));
	jdff dff_A_Uyxa1jdV3_0(.dout(w_G143_0[0]),.din(w_dff_A_Uyxa1jdV3_0),.clk(gclk));
	jdff dff_A_zkrzFq9t3_0(.dout(w_dff_A_Uyxa1jdV3_0),.din(w_dff_A_zkrzFq9t3_0),.clk(gclk));
	jdff dff_A_K9SZtQG15_0(.dout(w_dff_A_zkrzFq9t3_0),.din(w_dff_A_K9SZtQG15_0),.clk(gclk));
	jdff dff_A_cAq71eL22_0(.dout(w_dff_A_K9SZtQG15_0),.din(w_dff_A_cAq71eL22_0),.clk(gclk));
	jdff dff_A_DMctQkqj2_0(.dout(w_dff_A_cAq71eL22_0),.din(w_dff_A_DMctQkqj2_0),.clk(gclk));
	jdff dff_A_5kjPYsut1_0(.dout(w_dff_A_DMctQkqj2_0),.din(w_dff_A_5kjPYsut1_0),.clk(gclk));
	jdff dff_A_EPv2wLsB0_0(.dout(w_dff_A_5kjPYsut1_0),.din(w_dff_A_EPv2wLsB0_0),.clk(gclk));
	jdff dff_A_mUg58g8w7_0(.dout(w_dff_A_EPv2wLsB0_0),.din(w_dff_A_mUg58g8w7_0),.clk(gclk));
	jdff dff_A_Lqr4g2Ii4_0(.dout(w_dff_A_mUg58g8w7_0),.din(w_dff_A_Lqr4g2Ii4_0),.clk(gclk));
	jdff dff_A_acBnNSvq5_0(.dout(w_dff_A_Lqr4g2Ii4_0),.din(w_dff_A_acBnNSvq5_0),.clk(gclk));
	jdff dff_A_54YWHNz46_0(.dout(w_dff_A_acBnNSvq5_0),.din(w_dff_A_54YWHNz46_0),.clk(gclk));
	jdff dff_A_8zc6us4R5_1(.dout(w_G143_0[1]),.din(w_dff_A_8zc6us4R5_1),.clk(gclk));
	jdff dff_A_AORReWib9_0(.dout(w_G128_0[0]),.din(w_dff_A_AORReWib9_0),.clk(gclk));
	jdff dff_A_KyWQvPab6_0(.dout(w_dff_A_AORReWib9_0),.din(w_dff_A_KyWQvPab6_0),.clk(gclk));
	jdff dff_A_Rzh3Lz0I1_0(.dout(w_dff_A_KyWQvPab6_0),.din(w_dff_A_Rzh3Lz0I1_0),.clk(gclk));
	jdff dff_A_pF1zcXhi4_0(.dout(w_dff_A_Rzh3Lz0I1_0),.din(w_dff_A_pF1zcXhi4_0),.clk(gclk));
	jdff dff_A_rl57237d4_0(.dout(w_dff_A_pF1zcXhi4_0),.din(w_dff_A_rl57237d4_0),.clk(gclk));
	jdff dff_A_pZkQA3H45_0(.dout(w_dff_A_rl57237d4_0),.din(w_dff_A_pZkQA3H45_0),.clk(gclk));
	jdff dff_A_spANxOh15_0(.dout(w_dff_A_pZkQA3H45_0),.din(w_dff_A_spANxOh15_0),.clk(gclk));
	jdff dff_A_qKeaOSgV5_0(.dout(w_dff_A_spANxOh15_0),.din(w_dff_A_qKeaOSgV5_0),.clk(gclk));
	jdff dff_A_8K7YSytW6_0(.dout(w_dff_A_qKeaOSgV5_0),.din(w_dff_A_8K7YSytW6_0),.clk(gclk));
	jdff dff_A_iOz0fSRG1_0(.dout(w_dff_A_8K7YSytW6_0),.din(w_dff_A_iOz0fSRG1_0),.clk(gclk));
	jdff dff_A_julECBpF0_0(.dout(w_dff_A_iOz0fSRG1_0),.din(w_dff_A_julECBpF0_0),.clk(gclk));
	jdff dff_A_ZgKH4qLv2_0(.dout(w_G134_0[0]),.din(w_dff_A_ZgKH4qLv2_0),.clk(gclk));
	jdff dff_A_1dOdWFbt4_0(.dout(w_dff_A_ZgKH4qLv2_0),.din(w_dff_A_1dOdWFbt4_0),.clk(gclk));
	jdff dff_A_RvvqsymX1_0(.dout(w_dff_A_1dOdWFbt4_0),.din(w_dff_A_RvvqsymX1_0),.clk(gclk));
	jdff dff_A_hIegGQQ95_0(.dout(w_dff_A_RvvqsymX1_0),.din(w_dff_A_hIegGQQ95_0),.clk(gclk));
	jdff dff_A_8I6G7J8J1_0(.dout(w_dff_A_hIegGQQ95_0),.din(w_dff_A_8I6G7J8J1_0),.clk(gclk));
	jdff dff_A_A0OAUl0l0_0(.dout(w_dff_A_8I6G7J8J1_0),.din(w_dff_A_A0OAUl0l0_0),.clk(gclk));
	jdff dff_A_zM1WbSZ23_0(.dout(w_dff_A_A0OAUl0l0_0),.din(w_dff_A_zM1WbSZ23_0),.clk(gclk));
	jdff dff_A_PCdON3043_0(.dout(w_dff_A_zM1WbSZ23_0),.din(w_dff_A_PCdON3043_0),.clk(gclk));
	jdff dff_A_EYRc5Jg54_0(.dout(w_dff_A_PCdON3043_0),.din(w_dff_A_EYRc5Jg54_0),.clk(gclk));
	jdff dff_A_kHr6qwOO9_0(.dout(w_dff_A_EYRc5Jg54_0),.din(w_dff_A_kHr6qwOO9_0),.clk(gclk));
	jdff dff_A_6fVrQNeK2_0(.dout(w_dff_A_kHr6qwOO9_0),.din(w_dff_A_6fVrQNeK2_0),.clk(gclk));
	jdff dff_A_Ceh9Y6RA4_1(.dout(w_G134_0[1]),.din(w_dff_A_Ceh9Y6RA4_1),.clk(gclk));
	jdff dff_A_zs8FWjcf8_0(.dout(w_n58_0[0]),.din(w_dff_A_zs8FWjcf8_0),.clk(gclk));
	jdff dff_A_V4m9vpmB8_0(.dout(w_dff_A_zs8FWjcf8_0),.din(w_dff_A_V4m9vpmB8_0),.clk(gclk));
	jdff dff_A_QaqVoQ6i3_0(.dout(w_dff_A_V4m9vpmB8_0),.din(w_dff_A_QaqVoQ6i3_0),.clk(gclk));
	jdff dff_A_N1JBoeja7_0(.dout(w_dff_A_QaqVoQ6i3_0),.din(w_dff_A_N1JBoeja7_0),.clk(gclk));
	jdff dff_A_Yhai2ikW0_2(.dout(w_n58_0[2]),.din(w_dff_A_Yhai2ikW0_2),.clk(gclk));
	jdff dff_A_FLDsYRoa1_2(.dout(w_dff_A_Yhai2ikW0_2),.din(w_dff_A_FLDsYRoa1_2),.clk(gclk));
	jdff dff_A_6IOIBCTc9_2(.dout(w_dff_A_FLDsYRoa1_2),.din(w_dff_A_6IOIBCTc9_2),.clk(gclk));
	jdff dff_A_mcU4tgIv0_2(.dout(w_dff_A_6IOIBCTc9_2),.din(w_dff_A_mcU4tgIv0_2),.clk(gclk));
	jdff dff_A_2c3QfiNY0_0(.dout(w_G902_3[0]),.din(w_dff_A_2c3QfiNY0_0),.clk(gclk));
	jdff dff_A_tiODlU1F4_0(.dout(w_dff_A_2c3QfiNY0_0),.din(w_dff_A_tiODlU1F4_0),.clk(gclk));
	jdff dff_A_hOHbir0a9_0(.dout(w_G478_0[0]),.din(w_dff_A_hOHbir0a9_0),.clk(gclk));
	jdff dff_A_PDjWm0sn2_0(.dout(w_dff_A_hOHbir0a9_0),.din(w_dff_A_PDjWm0sn2_0),.clk(gclk));
	jdff dff_A_oeZgErjw3_0(.dout(w_dff_A_PDjWm0sn2_0),.din(w_dff_A_oeZgErjw3_0),.clk(gclk));
	jdff dff_A_rDDXlFen1_0(.dout(w_dff_A_oeZgErjw3_0),.din(w_dff_A_rDDXlFen1_0),.clk(gclk));
	jdff dff_A_vsKFgpCk8_0(.dout(w_dff_A_rDDXlFen1_0),.din(w_dff_A_vsKFgpCk8_0),.clk(gclk));
	jdff dff_A_VAUH35qY0_0(.dout(w_dff_A_vsKFgpCk8_0),.din(w_dff_A_VAUH35qY0_0),.clk(gclk));
	jdff dff_A_vTG6tajw1_0(.dout(w_dff_A_VAUH35qY0_0),.din(w_dff_A_vTG6tajw1_0),.clk(gclk));
	jdff dff_A_ucS4E2g80_0(.dout(w_dff_A_vTG6tajw1_0),.din(w_dff_A_ucS4E2g80_0),.clk(gclk));
	jdff dff_A_Jb8hfndA9_0(.dout(w_dff_A_ucS4E2g80_0),.din(w_dff_A_Jb8hfndA9_0),.clk(gclk));
	jdff dff_A_bEVz6YNV4_0(.dout(w_dff_A_Jb8hfndA9_0),.din(w_dff_A_bEVz6YNV4_0),.clk(gclk));
	jdff dff_A_VoKtbupI5_0(.dout(w_dff_A_bEVz6YNV4_0),.din(w_dff_A_VoKtbupI5_0),.clk(gclk));
	jdff dff_A_pjFHUqEz0_0(.dout(w_dff_A_VoKtbupI5_0),.din(w_dff_A_pjFHUqEz0_0),.clk(gclk));
	jdff dff_A_pIvRJMFZ7_0(.dout(w_dff_A_pjFHUqEz0_0),.din(w_dff_A_pIvRJMFZ7_0),.clk(gclk));
	jdff dff_A_dzFctr5t1_0(.dout(w_dff_A_pIvRJMFZ7_0),.din(w_dff_A_dzFctr5t1_0),.clk(gclk));
	jdff dff_A_T4qmQgTn8_0(.dout(w_dff_A_dzFctr5t1_0),.din(w_dff_A_T4qmQgTn8_0),.clk(gclk));
	jdff dff_A_fKDY7Nsc9_0(.dout(w_dff_A_T4qmQgTn8_0),.din(w_dff_A_fKDY7Nsc9_0),.clk(gclk));
	jdff dff_A_M02w6KUf3_1(.dout(w_G478_0[1]),.din(w_dff_A_M02w6KUf3_1),.clk(gclk));
	jdff dff_A_72LYaYfb0_1(.dout(w_dff_A_M02w6KUf3_1),.din(w_dff_A_72LYaYfb0_1),.clk(gclk));
	jdff dff_A_y4VWZT022_1(.dout(w_dff_A_72LYaYfb0_1),.din(w_dff_A_y4VWZT022_1),.clk(gclk));
	jdff dff_A_lm7bARAI1_1(.dout(w_dff_A_y4VWZT022_1),.din(w_dff_A_lm7bARAI1_1),.clk(gclk));
	jdff dff_A_VctRwhUr7_1(.dout(w_dff_A_lm7bARAI1_1),.din(w_dff_A_VctRwhUr7_1),.clk(gclk));
	jdff dff_A_l0eGAroD5_1(.dout(w_dff_A_VctRwhUr7_1),.din(w_dff_A_l0eGAroD5_1),.clk(gclk));
	jdff dff_A_H8dpCByK6_1(.dout(w_n265_0[1]),.din(w_dff_A_H8dpCByK6_1),.clk(gclk));
	jdff dff_B_3KlfMBQA9_3(.din(n265),.dout(w_dff_B_3KlfMBQA9_3),.clk(gclk));
	jdff dff_B_8tesdH5w4_3(.din(w_dff_B_3KlfMBQA9_3),.dout(w_dff_B_8tesdH5w4_3),.clk(gclk));
	jdff dff_B_EhBHDecs2_3(.din(w_dff_B_8tesdH5w4_3),.dout(w_dff_B_EhBHDecs2_3),.clk(gclk));
	jdff dff_B_uKTTEheB9_3(.din(w_dff_B_EhBHDecs2_3),.dout(w_dff_B_uKTTEheB9_3),.clk(gclk));
	jdff dff_B_zc3zs5xo6_3(.din(w_dff_B_uKTTEheB9_3),.dout(w_dff_B_zc3zs5xo6_3),.clk(gclk));
	jdff dff_B_Zwqu0bqe7_3(.din(w_dff_B_zc3zs5xo6_3),.dout(w_dff_B_Zwqu0bqe7_3),.clk(gclk));
	jdff dff_B_sJBTHqkT3_3(.din(w_dff_B_Zwqu0bqe7_3),.dout(w_dff_B_sJBTHqkT3_3),.clk(gclk));
	jdff dff_B_8ar9O2Ie3_3(.din(w_dff_B_sJBTHqkT3_3),.dout(w_dff_B_8ar9O2Ie3_3),.clk(gclk));
	jdff dff_B_xfDn2R9L6_3(.din(w_dff_B_8ar9O2Ie3_3),.dout(w_dff_B_xfDn2R9L6_3),.clk(gclk));
	jdff dff_B_QOUfgPnZ1_3(.din(w_dff_B_xfDn2R9L6_3),.dout(w_dff_B_QOUfgPnZ1_3),.clk(gclk));
	jdff dff_B_U7vSbnKH4_3(.din(w_dff_B_QOUfgPnZ1_3),.dout(w_dff_B_U7vSbnKH4_3),.clk(gclk));
	jdff dff_B_DqelCsKJ1_3(.din(w_dff_B_U7vSbnKH4_3),.dout(w_dff_B_DqelCsKJ1_3),.clk(gclk));
	jdff dff_B_D4fHQvLF9_3(.din(w_dff_B_DqelCsKJ1_3),.dout(w_dff_B_D4fHQvLF9_3),.clk(gclk));
	jdff dff_B_yNpts7NY5_3(.din(w_dff_B_D4fHQvLF9_3),.dout(w_dff_B_yNpts7NY5_3),.clk(gclk));
	jdff dff_B_S7LHnDBT9_3(.din(w_dff_B_yNpts7NY5_3),.dout(w_dff_B_S7LHnDBT9_3),.clk(gclk));
	jdff dff_B_YCfBBzZ70_3(.din(w_dff_B_S7LHnDBT9_3),.dout(w_dff_B_YCfBBzZ70_3),.clk(gclk));
	jdff dff_A_lOKFUup95_0(.dout(w_G953_1[0]),.din(w_dff_A_lOKFUup95_0),.clk(gclk));
	jdff dff_A_6IiluKjv0_0(.dout(w_dff_A_lOKFUup95_0),.din(w_dff_A_6IiluKjv0_0),.clk(gclk));
	jdff dff_A_P78E6ndu2_0(.dout(w_dff_A_6IiluKjv0_0),.din(w_dff_A_P78E6ndu2_0),.clk(gclk));
	jdff dff_A_OO4BfbEG7_0(.dout(w_dff_A_P78E6ndu2_0),.din(w_dff_A_OO4BfbEG7_0),.clk(gclk));
	jdff dff_A_xipyZCpr9_0(.dout(w_dff_A_OO4BfbEG7_0),.din(w_dff_A_xipyZCpr9_0),.clk(gclk));
	jdff dff_A_ziVXBFSx5_0(.dout(w_dff_A_xipyZCpr9_0),.din(w_dff_A_ziVXBFSx5_0),.clk(gclk));
	jdff dff_A_ZHuVen6B4_0(.dout(w_dff_A_ziVXBFSx5_0),.din(w_dff_A_ZHuVen6B4_0),.clk(gclk));
	jdff dff_A_zpFHcZRZ8_0(.dout(w_dff_A_ZHuVen6B4_0),.din(w_dff_A_zpFHcZRZ8_0),.clk(gclk));
	jdff dff_A_q69mUsiW8_0(.dout(w_dff_A_zpFHcZRZ8_0),.din(w_dff_A_q69mUsiW8_0),.clk(gclk));
	jdff dff_A_ddiVUbg04_0(.dout(w_dff_A_q69mUsiW8_0),.din(w_dff_A_ddiVUbg04_0),.clk(gclk));
	jdff dff_A_rh9P2G2O0_0(.dout(w_dff_A_ddiVUbg04_0),.din(w_dff_A_rh9P2G2O0_0),.clk(gclk));
	jdff dff_A_2A6pMAIZ8_0(.dout(w_dff_A_rh9P2G2O0_0),.din(w_dff_A_2A6pMAIZ8_0),.clk(gclk));
	jdff dff_A_ynZYaNpE5_0(.dout(w_dff_A_2A6pMAIZ8_0),.din(w_dff_A_ynZYaNpE5_0),.clk(gclk));
	jdff dff_A_ytvGwuEO0_0(.dout(w_dff_A_ynZYaNpE5_0),.din(w_dff_A_ytvGwuEO0_0),.clk(gclk));
	jdff dff_A_KXfeyVnS8_0(.dout(w_dff_A_ytvGwuEO0_0),.din(w_dff_A_KXfeyVnS8_0),.clk(gclk));
	jdff dff_A_Pm1Qpj9M2_1(.dout(w_G953_1[1]),.din(w_dff_A_Pm1Qpj9M2_1),.clk(gclk));
	jdff dff_A_R0LuugEo0_1(.dout(w_dff_A_Pm1Qpj9M2_1),.din(w_dff_A_R0LuugEo0_1),.clk(gclk));
	jdff dff_A_F2zpO55S0_1(.dout(w_dff_A_R0LuugEo0_1),.din(w_dff_A_F2zpO55S0_1),.clk(gclk));
	jdff dff_A_B43PHoVe5_1(.dout(w_dff_A_F2zpO55S0_1),.din(w_dff_A_B43PHoVe5_1),.clk(gclk));
	jdff dff_A_qGTl746B6_1(.dout(w_dff_A_B43PHoVe5_1),.din(w_dff_A_qGTl746B6_1),.clk(gclk));
	jdff dff_A_UVsxiAya9_1(.dout(w_dff_A_qGTl746B6_1),.din(w_dff_A_UVsxiAya9_1),.clk(gclk));
	jdff dff_A_Iv2EG6hp6_1(.dout(w_dff_A_UVsxiAya9_1),.din(w_dff_A_Iv2EG6hp6_1),.clk(gclk));
	jdff dff_A_COnjRR6S4_1(.dout(w_dff_A_Iv2EG6hp6_1),.din(w_dff_A_COnjRR6S4_1),.clk(gclk));
	jdff dff_A_MNLVDXSy7_1(.dout(w_dff_A_COnjRR6S4_1),.din(w_dff_A_MNLVDXSy7_1),.clk(gclk));
	jdff dff_A_ZgTAUQXH8_1(.dout(w_dff_A_MNLVDXSy7_1),.din(w_dff_A_ZgTAUQXH8_1),.clk(gclk));
	jdff dff_A_iaZIgbic2_1(.dout(w_dff_A_ZgTAUQXH8_1),.din(w_dff_A_iaZIgbic2_1),.clk(gclk));
	jdff dff_A_UGqxG0g45_1(.dout(w_dff_A_iaZIgbic2_1),.din(w_dff_A_UGqxG0g45_1),.clk(gclk));
	jdff dff_A_GgAyF5bf5_2(.dout(w_G953_0[2]),.din(w_dff_A_GgAyF5bf5_2),.clk(gclk));
	jdff dff_A_gL2fNxA12_2(.dout(w_dff_A_GgAyF5bf5_2),.din(w_dff_A_gL2fNxA12_2),.clk(gclk));
	jdff dff_A_9j5upJDu4_2(.dout(w_dff_A_gL2fNxA12_2),.din(w_dff_A_9j5upJDu4_2),.clk(gclk));
	jdff dff_A_ffBxmw9z8_2(.dout(w_dff_A_9j5upJDu4_2),.din(w_dff_A_ffBxmw9z8_2),.clk(gclk));
	jdff dff_A_WVS9tnBF5_2(.dout(w_dff_A_ffBxmw9z8_2),.din(w_dff_A_WVS9tnBF5_2),.clk(gclk));
	jdff dff_A_t6SN8CFU6_2(.dout(w_dff_A_WVS9tnBF5_2),.din(w_dff_A_t6SN8CFU6_2),.clk(gclk));
	jdff dff_A_PgL2PPIp4_2(.dout(w_dff_A_t6SN8CFU6_2),.din(w_dff_A_PgL2PPIp4_2),.clk(gclk));
	jdff dff_A_ymkJJMVU8_2(.dout(w_dff_A_PgL2PPIp4_2),.din(w_dff_A_ymkJJMVU8_2),.clk(gclk));
	jdff dff_A_HcSQSjMQ5_2(.dout(w_dff_A_ymkJJMVU8_2),.din(w_dff_A_HcSQSjMQ5_2),.clk(gclk));
	jdff dff_A_qHM1NRBl1_2(.dout(w_dff_A_HcSQSjMQ5_2),.din(w_dff_A_qHM1NRBl1_2),.clk(gclk));
	jdff dff_A_oPrdO45e4_2(.dout(w_dff_A_qHM1NRBl1_2),.din(w_dff_A_oPrdO45e4_2),.clk(gclk));
	jdff dff_A_55uuqk1i8_2(.dout(w_dff_A_oPrdO45e4_2),.din(w_dff_A_55uuqk1i8_2),.clk(gclk));
	jdff dff_A_l4P3fljX2_2(.dout(w_dff_A_55uuqk1i8_2),.din(w_dff_A_l4P3fljX2_2),.clk(gclk));
	jdff dff_A_e8jTiCF58_2(.dout(w_dff_A_l4P3fljX2_2),.din(w_dff_A_e8jTiCF58_2),.clk(gclk));
	jdff dff_A_hiFdIg9Q8_2(.dout(w_dff_A_e8jTiCF58_2),.din(w_dff_A_hiFdIg9Q8_2),.clk(gclk));
	jdff dff_A_B6LlEjr60_1(.dout(w_G952_0[1]),.din(w_dff_A_B6LlEjr60_1),.clk(gclk));
	jdff dff_A_6i0kJJaO8_1(.dout(w_dff_A_B6LlEjr60_1),.din(w_dff_A_6i0kJJaO8_1),.clk(gclk));
	jdff dff_A_jDjCFC3n9_1(.dout(w_dff_A_6i0kJJaO8_1),.din(w_dff_A_jDjCFC3n9_1),.clk(gclk));
	jdff dff_A_DiTXsm7e1_1(.dout(w_dff_A_jDjCFC3n9_1),.din(w_dff_A_DiTXsm7e1_1),.clk(gclk));
	jdff dff_A_RjD8HaVJ3_1(.dout(w_dff_A_DiTXsm7e1_1),.din(w_dff_A_RjD8HaVJ3_1),.clk(gclk));
	jdff dff_A_WAk2OABQ1_1(.dout(w_dff_A_RjD8HaVJ3_1),.din(w_dff_A_WAk2OABQ1_1),.clk(gclk));
	jdff dff_A_lRkGRM7K0_1(.dout(w_dff_A_WAk2OABQ1_1),.din(w_dff_A_lRkGRM7K0_1),.clk(gclk));
	jdff dff_A_7YDbiEcs0_1(.dout(w_dff_A_lRkGRM7K0_1),.din(w_dff_A_7YDbiEcs0_1),.clk(gclk));
	jdff dff_A_2OnvTU1x7_1(.dout(w_dff_A_7YDbiEcs0_1),.din(w_dff_A_2OnvTU1x7_1),.clk(gclk));
	jdff dff_A_PXeVG97y2_1(.dout(w_dff_A_2OnvTU1x7_1),.din(w_dff_A_PXeVG97y2_1),.clk(gclk));
	jdff dff_A_kTVJeEXa9_1(.dout(w_dff_A_PXeVG97y2_1),.din(w_dff_A_kTVJeEXa9_1),.clk(gclk));
	jdff dff_A_6BJkxyXk5_1(.dout(w_dff_A_kTVJeEXa9_1),.din(w_dff_A_6BJkxyXk5_1),.clk(gclk));
	jdff dff_A_nmLjS0oG8_1(.dout(w_dff_A_6BJkxyXk5_1),.din(w_dff_A_nmLjS0oG8_1),.clk(gclk));
	jdff dff_A_QdnxJQn89_1(.dout(w_dff_A_nmLjS0oG8_1),.din(w_dff_A_QdnxJQn89_1),.clk(gclk));
	jdff dff_A_xvDgcW3l1_1(.dout(w_dff_A_QdnxJQn89_1),.din(w_dff_A_xvDgcW3l1_1),.clk(gclk));
	jdff dff_A_GJtCJ9al0_1(.dout(w_dff_A_xvDgcW3l1_1),.din(w_dff_A_GJtCJ9al0_1),.clk(gclk));
	jdff dff_A_SjzwPv5X2_2(.dout(w_G952_0[2]),.din(w_dff_A_SjzwPv5X2_2),.clk(gclk));
	jdff dff_B_PjuaBNu04_3(.din(G952),.dout(w_dff_B_PjuaBNu04_3),.clk(gclk));
	jdff dff_A_1HIeDp7r2_2(.dout(w_dff_A_dpSwxm545_0),.din(w_dff_A_1HIeDp7r2_2),.clk(gclk));
	jdff dff_A_dpSwxm545_0(.dout(w_dff_A_mbF8eUps7_0),.din(w_dff_A_dpSwxm545_0),.clk(gclk));
	jdff dff_A_mbF8eUps7_0(.dout(w_dff_A_HxWVCLTv5_0),.din(w_dff_A_mbF8eUps7_0),.clk(gclk));
	jdff dff_A_HxWVCLTv5_0(.dout(w_dff_A_g7FwyZWy5_0),.din(w_dff_A_HxWVCLTv5_0),.clk(gclk));
	jdff dff_A_g7FwyZWy5_0(.dout(w_dff_A_6FZWLiIJ4_0),.din(w_dff_A_g7FwyZWy5_0),.clk(gclk));
	jdff dff_A_6FZWLiIJ4_0(.dout(w_dff_A_QwsrG7Az8_0),.din(w_dff_A_6FZWLiIJ4_0),.clk(gclk));
	jdff dff_A_QwsrG7Az8_0(.dout(w_dff_A_Cxg7nzTV6_0),.din(w_dff_A_QwsrG7Az8_0),.clk(gclk));
	jdff dff_A_Cxg7nzTV6_0(.dout(G3),.din(w_dff_A_Cxg7nzTV6_0),.clk(gclk));
	jdff dff_A_jzkZ6mNp7_2(.dout(w_dff_A_MHUHYXTa4_0),.din(w_dff_A_jzkZ6mNp7_2),.clk(gclk));
	jdff dff_A_MHUHYXTa4_0(.dout(w_dff_A_JswjQ0108_0),.din(w_dff_A_MHUHYXTa4_0),.clk(gclk));
	jdff dff_A_JswjQ0108_0(.dout(w_dff_A_0o8yrJiR2_0),.din(w_dff_A_JswjQ0108_0),.clk(gclk));
	jdff dff_A_0o8yrJiR2_0(.dout(w_dff_A_8x2BsPps5_0),.din(w_dff_A_0o8yrJiR2_0),.clk(gclk));
	jdff dff_A_8x2BsPps5_0(.dout(w_dff_A_q9TbdOh14_0),.din(w_dff_A_8x2BsPps5_0),.clk(gclk));
	jdff dff_A_q9TbdOh14_0(.dout(w_dff_A_uS4mnpUH5_0),.din(w_dff_A_q9TbdOh14_0),.clk(gclk));
	jdff dff_A_uS4mnpUH5_0(.dout(w_dff_A_s1Tj0OV23_0),.din(w_dff_A_uS4mnpUH5_0),.clk(gclk));
	jdff dff_A_s1Tj0OV23_0(.dout(G6),.din(w_dff_A_s1Tj0OV23_0),.clk(gclk));
	jdff dff_A_25G69Rjr9_2(.dout(w_dff_A_10Sdgrvs1_0),.din(w_dff_A_25G69Rjr9_2),.clk(gclk));
	jdff dff_A_10Sdgrvs1_0(.dout(w_dff_A_FaslhWba5_0),.din(w_dff_A_10Sdgrvs1_0),.clk(gclk));
	jdff dff_A_FaslhWba5_0(.dout(w_dff_A_1DTnCy7r5_0),.din(w_dff_A_FaslhWba5_0),.clk(gclk));
	jdff dff_A_1DTnCy7r5_0(.dout(w_dff_A_1ELhKcnn8_0),.din(w_dff_A_1DTnCy7r5_0),.clk(gclk));
	jdff dff_A_1ELhKcnn8_0(.dout(w_dff_A_SMhhcGkr1_0),.din(w_dff_A_1ELhKcnn8_0),.clk(gclk));
	jdff dff_A_SMhhcGkr1_0(.dout(w_dff_A_iSJ9zS557_0),.din(w_dff_A_SMhhcGkr1_0),.clk(gclk));
	jdff dff_A_iSJ9zS557_0(.dout(w_dff_A_KvuzvACb3_0),.din(w_dff_A_iSJ9zS557_0),.clk(gclk));
	jdff dff_A_KvuzvACb3_0(.dout(G9),.din(w_dff_A_KvuzvACb3_0),.clk(gclk));
	jdff dff_A_z3wcJUFY4_2(.dout(w_dff_A_fMbK2QzZ0_0),.din(w_dff_A_z3wcJUFY4_2),.clk(gclk));
	jdff dff_A_fMbK2QzZ0_0(.dout(w_dff_A_Wo1G8lMq3_0),.din(w_dff_A_fMbK2QzZ0_0),.clk(gclk));
	jdff dff_A_Wo1G8lMq3_0(.dout(w_dff_A_7CQajTHE1_0),.din(w_dff_A_Wo1G8lMq3_0),.clk(gclk));
	jdff dff_A_7CQajTHE1_0(.dout(w_dff_A_8lqg625L3_0),.din(w_dff_A_7CQajTHE1_0),.clk(gclk));
	jdff dff_A_8lqg625L3_0(.dout(w_dff_A_saG0aem95_0),.din(w_dff_A_8lqg625L3_0),.clk(gclk));
	jdff dff_A_saG0aem95_0(.dout(w_dff_A_LOMJq8wV4_0),.din(w_dff_A_saG0aem95_0),.clk(gclk));
	jdff dff_A_LOMJq8wV4_0(.dout(w_dff_A_mHbDUKf35_0),.din(w_dff_A_LOMJq8wV4_0),.clk(gclk));
	jdff dff_A_mHbDUKf35_0(.dout(G12),.din(w_dff_A_mHbDUKf35_0),.clk(gclk));
	jdff dff_A_WlpV7S0I3_2(.dout(w_dff_A_VoTwe0xA1_0),.din(w_dff_A_WlpV7S0I3_2),.clk(gclk));
	jdff dff_A_VoTwe0xA1_0(.dout(w_dff_A_a5uXxZFv3_0),.din(w_dff_A_VoTwe0xA1_0),.clk(gclk));
	jdff dff_A_a5uXxZFv3_0(.dout(w_dff_A_QdCzHjlB6_0),.din(w_dff_A_a5uXxZFv3_0),.clk(gclk));
	jdff dff_A_QdCzHjlB6_0(.dout(w_dff_A_So69hqCf3_0),.din(w_dff_A_QdCzHjlB6_0),.clk(gclk));
	jdff dff_A_So69hqCf3_0(.dout(w_dff_A_MiPx4MOj1_0),.din(w_dff_A_So69hqCf3_0),.clk(gclk));
	jdff dff_A_MiPx4MOj1_0(.dout(w_dff_A_CdOhcoDh7_0),.din(w_dff_A_MiPx4MOj1_0),.clk(gclk));
	jdff dff_A_CdOhcoDh7_0(.dout(w_dff_A_0q5J7Jwn5_0),.din(w_dff_A_CdOhcoDh7_0),.clk(gclk));
	jdff dff_A_0q5J7Jwn5_0(.dout(G30),.din(w_dff_A_0q5J7Jwn5_0),.clk(gclk));
	jdff dff_A_WaS3U3aF1_2(.dout(w_dff_A_tGyO216O7_0),.din(w_dff_A_WaS3U3aF1_2),.clk(gclk));
	jdff dff_A_tGyO216O7_0(.dout(w_dff_A_eU4F72ku8_0),.din(w_dff_A_tGyO216O7_0),.clk(gclk));
	jdff dff_A_eU4F72ku8_0(.dout(w_dff_A_0luz7jIX0_0),.din(w_dff_A_eU4F72ku8_0),.clk(gclk));
	jdff dff_A_0luz7jIX0_0(.dout(w_dff_A_iSjbBr9t4_0),.din(w_dff_A_0luz7jIX0_0),.clk(gclk));
	jdff dff_A_iSjbBr9t4_0(.dout(w_dff_A_iF7uQ93P1_0),.din(w_dff_A_iSjbBr9t4_0),.clk(gclk));
	jdff dff_A_iF7uQ93P1_0(.dout(w_dff_A_NwXul5tS7_0),.din(w_dff_A_iF7uQ93P1_0),.clk(gclk));
	jdff dff_A_NwXul5tS7_0(.dout(w_dff_A_jnawhvD27_0),.din(w_dff_A_NwXul5tS7_0),.clk(gclk));
	jdff dff_A_jnawhvD27_0(.dout(G45),.din(w_dff_A_jnawhvD27_0),.clk(gclk));
	jdff dff_A_kpZMc0eW0_2(.dout(w_dff_A_3b77LA202_0),.din(w_dff_A_kpZMc0eW0_2),.clk(gclk));
	jdff dff_A_3b77LA202_0(.dout(w_dff_A_JFjWkVH60_0),.din(w_dff_A_3b77LA202_0),.clk(gclk));
	jdff dff_A_JFjWkVH60_0(.dout(w_dff_A_MQIPxl8C9_0),.din(w_dff_A_JFjWkVH60_0),.clk(gclk));
	jdff dff_A_MQIPxl8C9_0(.dout(w_dff_A_LNxAYDtE5_0),.din(w_dff_A_MQIPxl8C9_0),.clk(gclk));
	jdff dff_A_LNxAYDtE5_0(.dout(w_dff_A_JnVtZDyB7_0),.din(w_dff_A_LNxAYDtE5_0),.clk(gclk));
	jdff dff_A_JnVtZDyB7_0(.dout(w_dff_A_nlz9VTaX2_0),.din(w_dff_A_JnVtZDyB7_0),.clk(gclk));
	jdff dff_A_nlz9VTaX2_0(.dout(w_dff_A_APdtuPOw8_0),.din(w_dff_A_nlz9VTaX2_0),.clk(gclk));
	jdff dff_A_APdtuPOw8_0(.dout(G48),.din(w_dff_A_APdtuPOw8_0),.clk(gclk));
	jdff dff_A_f5o7qxak1_2(.dout(w_dff_A_8vuCgLM62_0),.din(w_dff_A_f5o7qxak1_2),.clk(gclk));
	jdff dff_A_8vuCgLM62_0(.dout(w_dff_A_Dscj6AP62_0),.din(w_dff_A_8vuCgLM62_0),.clk(gclk));
	jdff dff_A_Dscj6AP62_0(.dout(w_dff_A_lNCbob4Z0_0),.din(w_dff_A_Dscj6AP62_0),.clk(gclk));
	jdff dff_A_lNCbob4Z0_0(.dout(w_dff_A_tztno8Af8_0),.din(w_dff_A_lNCbob4Z0_0),.clk(gclk));
	jdff dff_A_tztno8Af8_0(.dout(w_dff_A_AGXe5uzd6_0),.din(w_dff_A_tztno8Af8_0),.clk(gclk));
	jdff dff_A_AGXe5uzd6_0(.dout(w_dff_A_fGrWdj768_0),.din(w_dff_A_AGXe5uzd6_0),.clk(gclk));
	jdff dff_A_fGrWdj768_0(.dout(w_dff_A_VFoC8jf03_0),.din(w_dff_A_fGrWdj768_0),.clk(gclk));
	jdff dff_A_VFoC8jf03_0(.dout(G15),.din(w_dff_A_VFoC8jf03_0),.clk(gclk));
	jdff dff_A_bVp1TW5f3_2(.dout(w_dff_A_DI95F5hg9_0),.din(w_dff_A_bVp1TW5f3_2),.clk(gclk));
	jdff dff_A_DI95F5hg9_0(.dout(w_dff_A_OrR0toCO2_0),.din(w_dff_A_DI95F5hg9_0),.clk(gclk));
	jdff dff_A_OrR0toCO2_0(.dout(w_dff_A_YVx5EXNo1_0),.din(w_dff_A_OrR0toCO2_0),.clk(gclk));
	jdff dff_A_YVx5EXNo1_0(.dout(w_dff_A_fBBFJml14_0),.din(w_dff_A_YVx5EXNo1_0),.clk(gclk));
	jdff dff_A_fBBFJml14_0(.dout(w_dff_A_rhUCwuWP0_0),.din(w_dff_A_fBBFJml14_0),.clk(gclk));
	jdff dff_A_rhUCwuWP0_0(.dout(w_dff_A_j6SjAFiZ1_0),.din(w_dff_A_rhUCwuWP0_0),.clk(gclk));
	jdff dff_A_j6SjAFiZ1_0(.dout(w_dff_A_SImkO0Rk1_0),.din(w_dff_A_j6SjAFiZ1_0),.clk(gclk));
	jdff dff_A_SImkO0Rk1_0(.dout(G18),.din(w_dff_A_SImkO0Rk1_0),.clk(gclk));
	jdff dff_A_2vzslNSD5_2(.dout(w_dff_A_sI4UH3hQ0_0),.din(w_dff_A_2vzslNSD5_2),.clk(gclk));
	jdff dff_A_sI4UH3hQ0_0(.dout(w_dff_A_SwaiIOem2_0),.din(w_dff_A_sI4UH3hQ0_0),.clk(gclk));
	jdff dff_A_SwaiIOem2_0(.dout(w_dff_A_VP0tGqfs2_0),.din(w_dff_A_SwaiIOem2_0),.clk(gclk));
	jdff dff_A_VP0tGqfs2_0(.dout(w_dff_A_KA9w5xpi9_0),.din(w_dff_A_VP0tGqfs2_0),.clk(gclk));
	jdff dff_A_KA9w5xpi9_0(.dout(w_dff_A_BxGNppwU5_0),.din(w_dff_A_KA9w5xpi9_0),.clk(gclk));
	jdff dff_A_BxGNppwU5_0(.dout(w_dff_A_4nlB5erg5_0),.din(w_dff_A_BxGNppwU5_0),.clk(gclk));
	jdff dff_A_4nlB5erg5_0(.dout(w_dff_A_y5BuBXWP1_0),.din(w_dff_A_4nlB5erg5_0),.clk(gclk));
	jdff dff_A_y5BuBXWP1_0(.dout(G21),.din(w_dff_A_y5BuBXWP1_0),.clk(gclk));
	jdff dff_A_UFllNdkx6_2(.dout(w_dff_A_ghEs7qxg9_0),.din(w_dff_A_UFllNdkx6_2),.clk(gclk));
	jdff dff_A_ghEs7qxg9_0(.dout(w_dff_A_7HEJrJgE8_0),.din(w_dff_A_ghEs7qxg9_0),.clk(gclk));
	jdff dff_A_7HEJrJgE8_0(.dout(w_dff_A_cUoP0DwX9_0),.din(w_dff_A_7HEJrJgE8_0),.clk(gclk));
	jdff dff_A_cUoP0DwX9_0(.dout(w_dff_A_lKrS4BBf5_0),.din(w_dff_A_cUoP0DwX9_0),.clk(gclk));
	jdff dff_A_lKrS4BBf5_0(.dout(w_dff_A_00VubZMV4_0),.din(w_dff_A_lKrS4BBf5_0),.clk(gclk));
	jdff dff_A_00VubZMV4_0(.dout(w_dff_A_cB17GowC3_0),.din(w_dff_A_00VubZMV4_0),.clk(gclk));
	jdff dff_A_cB17GowC3_0(.dout(G24),.din(w_dff_A_cB17GowC3_0),.clk(gclk));
	jdff dff_A_Bsw4eSI67_2(.dout(w_dff_A_iD9eMV6H3_0),.din(w_dff_A_Bsw4eSI67_2),.clk(gclk));
	jdff dff_A_iD9eMV6H3_0(.dout(w_dff_A_YooGIYis9_0),.din(w_dff_A_iD9eMV6H3_0),.clk(gclk));
	jdff dff_A_YooGIYis9_0(.dout(w_dff_A_Edk6p6ct2_0),.din(w_dff_A_YooGIYis9_0),.clk(gclk));
	jdff dff_A_Edk6p6ct2_0(.dout(w_dff_A_lDy7wSU71_0),.din(w_dff_A_Edk6p6ct2_0),.clk(gclk));
	jdff dff_A_lDy7wSU71_0(.dout(w_dff_A_sEFpQIxZ1_0),.din(w_dff_A_lDy7wSU71_0),.clk(gclk));
	jdff dff_A_sEFpQIxZ1_0(.dout(w_dff_A_KT6DvG4N0_0),.din(w_dff_A_sEFpQIxZ1_0),.clk(gclk));
	jdff dff_A_KT6DvG4N0_0(.dout(w_dff_A_T53P2MVF1_0),.din(w_dff_A_KT6DvG4N0_0),.clk(gclk));
	jdff dff_A_T53P2MVF1_0(.dout(G27),.din(w_dff_A_T53P2MVF1_0),.clk(gclk));
	jdff dff_A_l3LCzSx29_2(.dout(w_dff_A_6KJFuvAg5_0),.din(w_dff_A_l3LCzSx29_2),.clk(gclk));
	jdff dff_A_6KJFuvAg5_0(.dout(w_dff_A_pGn8BuzS1_0),.din(w_dff_A_6KJFuvAg5_0),.clk(gclk));
	jdff dff_A_pGn8BuzS1_0(.dout(w_dff_A_W7ei9MpB7_0),.din(w_dff_A_pGn8BuzS1_0),.clk(gclk));
	jdff dff_A_W7ei9MpB7_0(.dout(w_dff_A_Gkdd7hlu2_0),.din(w_dff_A_W7ei9MpB7_0),.clk(gclk));
	jdff dff_A_Gkdd7hlu2_0(.dout(w_dff_A_2nmwoshl0_0),.din(w_dff_A_Gkdd7hlu2_0),.clk(gclk));
	jdff dff_A_2nmwoshl0_0(.dout(w_dff_A_X3HwRawM5_0),.din(w_dff_A_2nmwoshl0_0),.clk(gclk));
	jdff dff_A_X3HwRawM5_0(.dout(w_dff_A_4htbBja82_0),.din(w_dff_A_X3HwRawM5_0),.clk(gclk));
	jdff dff_A_4htbBja82_0(.dout(G33),.din(w_dff_A_4htbBja82_0),.clk(gclk));
	jdff dff_A_dFpioPX11_2(.dout(w_dff_A_jGdEnVPo9_0),.din(w_dff_A_dFpioPX11_2),.clk(gclk));
	jdff dff_A_jGdEnVPo9_0(.dout(w_dff_A_9vTYiUYL5_0),.din(w_dff_A_jGdEnVPo9_0),.clk(gclk));
	jdff dff_A_9vTYiUYL5_0(.dout(w_dff_A_pkzt4W3q0_0),.din(w_dff_A_9vTYiUYL5_0),.clk(gclk));
	jdff dff_A_pkzt4W3q0_0(.dout(w_dff_A_FH4fhV2K5_0),.din(w_dff_A_pkzt4W3q0_0),.clk(gclk));
	jdff dff_A_FH4fhV2K5_0(.dout(w_dff_A_RU9wFu5j4_0),.din(w_dff_A_FH4fhV2K5_0),.clk(gclk));
	jdff dff_A_RU9wFu5j4_0(.dout(w_dff_A_zd3tJsmm7_0),.din(w_dff_A_RU9wFu5j4_0),.clk(gclk));
	jdff dff_A_zd3tJsmm7_0(.dout(w_dff_A_5tpsoEHB4_0),.din(w_dff_A_zd3tJsmm7_0),.clk(gclk));
	jdff dff_A_5tpsoEHB4_0(.dout(G36),.din(w_dff_A_5tpsoEHB4_0),.clk(gclk));
	jdff dff_A_OOU44twI0_2(.dout(w_dff_A_QH3hzpep6_0),.din(w_dff_A_OOU44twI0_2),.clk(gclk));
	jdff dff_A_QH3hzpep6_0(.dout(w_dff_A_BzPxYXdQ6_0),.din(w_dff_A_QH3hzpep6_0),.clk(gclk));
	jdff dff_A_BzPxYXdQ6_0(.dout(w_dff_A_dAi5970u2_0),.din(w_dff_A_BzPxYXdQ6_0),.clk(gclk));
	jdff dff_A_dAi5970u2_0(.dout(w_dff_A_eMIknfsY4_0),.din(w_dff_A_dAi5970u2_0),.clk(gclk));
	jdff dff_A_eMIknfsY4_0(.dout(w_dff_A_8jaJ9J2g5_0),.din(w_dff_A_eMIknfsY4_0),.clk(gclk));
	jdff dff_A_8jaJ9J2g5_0(.dout(w_dff_A_LkUdZLky5_0),.din(w_dff_A_8jaJ9J2g5_0),.clk(gclk));
	jdff dff_A_LkUdZLky5_0(.dout(w_dff_A_MQSqB57S8_0),.din(w_dff_A_LkUdZLky5_0),.clk(gclk));
	jdff dff_A_MQSqB57S8_0(.dout(G39),.din(w_dff_A_MQSqB57S8_0),.clk(gclk));
	jdff dff_A_eEjNbT6i5_2(.dout(w_dff_A_9FGrK7kQ6_0),.din(w_dff_A_eEjNbT6i5_2),.clk(gclk));
	jdff dff_A_9FGrK7kQ6_0(.dout(w_dff_A_JhBvAJBs9_0),.din(w_dff_A_9FGrK7kQ6_0),.clk(gclk));
	jdff dff_A_JhBvAJBs9_0(.dout(w_dff_A_naPF2VXU4_0),.din(w_dff_A_JhBvAJBs9_0),.clk(gclk));
	jdff dff_A_naPF2VXU4_0(.dout(w_dff_A_ocj3SyfO2_0),.din(w_dff_A_naPF2VXU4_0),.clk(gclk));
	jdff dff_A_ocj3SyfO2_0(.dout(w_dff_A_M9RFyUEd8_0),.din(w_dff_A_ocj3SyfO2_0),.clk(gclk));
	jdff dff_A_M9RFyUEd8_0(.dout(w_dff_A_AVJuVzmJ7_0),.din(w_dff_A_M9RFyUEd8_0),.clk(gclk));
	jdff dff_A_AVJuVzmJ7_0(.dout(w_dff_A_0mD1Bjnm5_0),.din(w_dff_A_AVJuVzmJ7_0),.clk(gclk));
	jdff dff_A_0mD1Bjnm5_0(.dout(G42),.din(w_dff_A_0mD1Bjnm5_0),.clk(gclk));
	jdff dff_A_2RADLT291_2(.dout(G75),.din(w_dff_A_2RADLT291_2),.clk(gclk));
	jdff dff_A_pXp8UqB39_2(.dout(w_dff_A_NOz3iSZT9_0),.din(w_dff_A_pXp8UqB39_2),.clk(gclk));
	jdff dff_A_NOz3iSZT9_0(.dout(G69),.din(w_dff_A_NOz3iSZT9_0),.clk(gclk));
	jdff dff_A_yveDk3Uy2_2(.dout(w_dff_A_2BecV9tE0_0),.din(w_dff_A_yveDk3Uy2_2),.clk(gclk));
	jdff dff_A_2BecV9tE0_0(.dout(G72),.din(w_dff_A_2BecV9tE0_0),.clk(gclk));
	jdff dff_A_o6nunRDk6_2(.dout(G57),.din(w_dff_A_o6nunRDk6_2),.clk(gclk));
endmodule

