/*

top:
	jspl: 56
	jspl3: 248
	jnot: 8
	jdff: 11
	jand: 304

Summary:
	jspl: 56
	jspl3: 248
	jnot: 8
	jdff: 11
	jand: 304

The maximum logic level gap of any gate:
	top: 1
*/

module gf_decoder(gclk, count0, count1, count2, count3, count4, count5, count6, count7, selectp10, selectp11, selectp12, selectp13, selectp14, selectp15, selectp16, selectp17, selectp18, selectp19, selectp110, selectp111, selectp112, selectp113, selectp114, selectp115, selectp116, selectp117, selectp118, selectp119, selectp120, selectp121, selectp122, selectp123, selectp124, selectp125, selectp126, selectp127, selectp128, selectp129, selectp130, selectp131, selectp132, selectp133, selectp134, selectp135, selectp136, selectp137, selectp138, selectp139, selectp140, selectp141, selectp142, selectp143, selectp144, selectp145, selectp146, selectp147, selectp148, selectp149, selectp150, selectp151, selectp152, selectp153, selectp154, selectp155, selectp156, selectp157, selectp158, selectp159, selectp160, selectp161, selectp162, selectp163, selectp164, selectp165, selectp166, selectp167, selectp168, selectp169, selectp170, selectp171, selectp172, selectp173, selectp174, selectp175, selectp176, selectp177, selectp178, selectp179, selectp180, selectp181, selectp182, selectp183, selectp184, selectp185, selectp186, selectp187, selectp188, selectp189, selectp190, selectp191, selectp192, selectp193, selectp194, selectp195, selectp196, selectp197, selectp198, selectp199, selectp1100, selectp1101, selectp1102, selectp1103, selectp1104, selectp1105, selectp1106, selectp1107, selectp1108, selectp1109, selectp1110, selectp1111, selectp1112, selectp1113, selectp1114, selectp1115, selectp1116, selectp1117, selectp1118, selectp1119, selectp1120, selectp1121, selectp1122, selectp1123, selectp1124, selectp1125, selectp1126, selectp1127, selectp20, selectp21, selectp22, selectp23, selectp24, selectp25, selectp26, selectp27, selectp28, selectp29, selectp210, selectp211, selectp212, selectp213, selectp214, selectp215, selectp216, selectp217, selectp218, selectp219, selectp220, selectp221, selectp222, selectp223, selectp224, selectp225, selectp226, selectp227, selectp228, selectp229, selectp230, selectp231, selectp232, selectp233, selectp234, selectp235, selectp236, selectp237, selectp238, selectp239, selectp240, selectp241, selectp242, selectp243, selectp244, selectp245, selectp246, selectp247, selectp248, selectp249, selectp250, selectp251, selectp252, selectp253, selectp254, selectp255, selectp256, selectp257, selectp258, selectp259, selectp260, selectp261, selectp262, selectp263, selectp264, selectp265, selectp266, selectp267, selectp268, selectp269, selectp270, selectp271, selectp272, selectp273, selectp274, selectp275, selectp276, selectp277, selectp278, selectp279, selectp280, selectp281, selectp282, selectp283, selectp284, selectp285, selectp286, selectp287, selectp288, selectp289, selectp290, selectp291, selectp292, selectp293, selectp294, selectp295, selectp296, selectp297, selectp298, selectp299, selectp2100, selectp2101, selectp2102, selectp2103, selectp2104, selectp2105, selectp2106, selectp2107, selectp2108, selectp2109, selectp2110, selectp2111, selectp2112, selectp2113, selectp2114, selectp2115, selectp2116, selectp2117, selectp2118, selectp2119, selectp2120, selectp2121, selectp2122, selectp2123, selectp2124, selectp2125, selectp2126, selectp2127);
	input gclk;
	input count0;
	input count1;
	input count2;
	input count3;
	input count4;
	input count5;
	input count6;
	input count7;
	output selectp10;
	output selectp11;
	output selectp12;
	output selectp13;
	output selectp14;
	output selectp15;
	output selectp16;
	output selectp17;
	output selectp18;
	output selectp19;
	output selectp110;
	output selectp111;
	output selectp112;
	output selectp113;
	output selectp114;
	output selectp115;
	output selectp116;
	output selectp117;
	output selectp118;
	output selectp119;
	output selectp120;
	output selectp121;
	output selectp122;
	output selectp123;
	output selectp124;
	output selectp125;
	output selectp126;
	output selectp127;
	output selectp128;
	output selectp129;
	output selectp130;
	output selectp131;
	output selectp132;
	output selectp133;
	output selectp134;
	output selectp135;
	output selectp136;
	output selectp137;
	output selectp138;
	output selectp139;
	output selectp140;
	output selectp141;
	output selectp142;
	output selectp143;
	output selectp144;
	output selectp145;
	output selectp146;
	output selectp147;
	output selectp148;
	output selectp149;
	output selectp150;
	output selectp151;
	output selectp152;
	output selectp153;
	output selectp154;
	output selectp155;
	output selectp156;
	output selectp157;
	output selectp158;
	output selectp159;
	output selectp160;
	output selectp161;
	output selectp162;
	output selectp163;
	output selectp164;
	output selectp165;
	output selectp166;
	output selectp167;
	output selectp168;
	output selectp169;
	output selectp170;
	output selectp171;
	output selectp172;
	output selectp173;
	output selectp174;
	output selectp175;
	output selectp176;
	output selectp177;
	output selectp178;
	output selectp179;
	output selectp180;
	output selectp181;
	output selectp182;
	output selectp183;
	output selectp184;
	output selectp185;
	output selectp186;
	output selectp187;
	output selectp188;
	output selectp189;
	output selectp190;
	output selectp191;
	output selectp192;
	output selectp193;
	output selectp194;
	output selectp195;
	output selectp196;
	output selectp197;
	output selectp198;
	output selectp199;
	output selectp1100;
	output selectp1101;
	output selectp1102;
	output selectp1103;
	output selectp1104;
	output selectp1105;
	output selectp1106;
	output selectp1107;
	output selectp1108;
	output selectp1109;
	output selectp1110;
	output selectp1111;
	output selectp1112;
	output selectp1113;
	output selectp1114;
	output selectp1115;
	output selectp1116;
	output selectp1117;
	output selectp1118;
	output selectp1119;
	output selectp1120;
	output selectp1121;
	output selectp1122;
	output selectp1123;
	output selectp1124;
	output selectp1125;
	output selectp1126;
	output selectp1127;
	output selectp20;
	output selectp21;
	output selectp22;
	output selectp23;
	output selectp24;
	output selectp25;
	output selectp26;
	output selectp27;
	output selectp28;
	output selectp29;
	output selectp210;
	output selectp211;
	output selectp212;
	output selectp213;
	output selectp214;
	output selectp215;
	output selectp216;
	output selectp217;
	output selectp218;
	output selectp219;
	output selectp220;
	output selectp221;
	output selectp222;
	output selectp223;
	output selectp224;
	output selectp225;
	output selectp226;
	output selectp227;
	output selectp228;
	output selectp229;
	output selectp230;
	output selectp231;
	output selectp232;
	output selectp233;
	output selectp234;
	output selectp235;
	output selectp236;
	output selectp237;
	output selectp238;
	output selectp239;
	output selectp240;
	output selectp241;
	output selectp242;
	output selectp243;
	output selectp244;
	output selectp245;
	output selectp246;
	output selectp247;
	output selectp248;
	output selectp249;
	output selectp250;
	output selectp251;
	output selectp252;
	output selectp253;
	output selectp254;
	output selectp255;
	output selectp256;
	output selectp257;
	output selectp258;
	output selectp259;
	output selectp260;
	output selectp261;
	output selectp262;
	output selectp263;
	output selectp264;
	output selectp265;
	output selectp266;
	output selectp267;
	output selectp268;
	output selectp269;
	output selectp270;
	output selectp271;
	output selectp272;
	output selectp273;
	output selectp274;
	output selectp275;
	output selectp276;
	output selectp277;
	output selectp278;
	output selectp279;
	output selectp280;
	output selectp281;
	output selectp282;
	output selectp283;
	output selectp284;
	output selectp285;
	output selectp286;
	output selectp287;
	output selectp288;
	output selectp289;
	output selectp290;
	output selectp291;
	output selectp292;
	output selectp293;
	output selectp294;
	output selectp295;
	output selectp296;
	output selectp297;
	output selectp298;
	output selectp299;
	output selectp2100;
	output selectp2101;
	output selectp2102;
	output selectp2103;
	output selectp2104;
	output selectp2105;
	output selectp2106;
	output selectp2107;
	output selectp2108;
	output selectp2109;
	output selectp2110;
	output selectp2111;
	output selectp2112;
	output selectp2113;
	output selectp2114;
	output selectp2115;
	output selectp2116;
	output selectp2117;
	output selectp2118;
	output selectp2119;
	output selectp2120;
	output selectp2121;
	output selectp2122;
	output selectp2123;
	output selectp2124;
	output selectp2125;
	output selectp2126;
	output selectp2127;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n278;
	wire n279;
	wire n281;
	wire n282;
	wire n284;
	wire n286;
	wire n287;
	wire n289;
	wire n290;
	wire n292;
	wire n294;
	wire n296;
	wire n297;
	wire n299;
	wire n301;
	wire n302;
	wire n304;
	wire n306;
	wire n308;
	wire n310;
	wire n312;
	wire n314;
	wire n315;
	wire n332;
	wire n333;
	wire n350;
	wire n351;
	wire n368;
	wire n369;
	wire n386;
	wire n403;
	wire n420;
	wire n437;
	wire n438;
	wire n439;
	wire n456;
	wire n473;
	wire n490;
	wire n507;
	wire n508;
	wire n525;
	wire n542;
	wire n559;
	wire[2:0] w_count0_0;
	wire[2:0] w_count1_0;
	wire[2:0] w_count2_0;
	wire[2:0] w_count3_0;
	wire[2:0] w_count4_0;
	wire[2:0] w_count5_0;
	wire[2:0] w_count6_0;
	wire[2:0] w_count7_0;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[2:0] w_n266_0;
	wire[1:0] w_n266_1;
	wire[1:0] w_n267_0;
	wire[2:0] w_n268_0;
	wire[1:0] w_n268_1;
	wire[2:0] w_n269_0;
	wire[2:0] w_n269_1;
	wire[2:0] w_n269_2;
	wire[2:0] w_n269_3;
	wire[2:0] w_n269_4;
	wire[2:0] w_n269_5;
	wire[2:0] w_n269_6;
	wire[1:0] w_n269_7;
	wire[1:0] w_n270_0;
	wire[1:0] w_n271_0;
	wire[2:0] w_n272_0;
	wire[1:0] w_n272_1;
	wire[1:0] w_n273_0;
	wire[1:0] w_n274_0;
	wire[2:0] w_n275_0;
	wire[1:0] w_n275_1;
	wire[2:0] w_n276_0;
	wire[2:0] w_n276_1;
	wire[2:0] w_n276_2;
	wire[2:0] w_n276_3;
	wire[2:0] w_n276_4;
	wire[2:0] w_n276_5;
	wire[2:0] w_n276_6;
	wire[1:0] w_n276_7;
	wire[2:0] w_n278_0;
	wire[1:0] w_n278_1;
	wire[2:0] w_n279_0;
	wire[2:0] w_n279_1;
	wire[2:0] w_n279_2;
	wire[2:0] w_n279_3;
	wire[2:0] w_n279_4;
	wire[2:0] w_n279_5;
	wire[2:0] w_n279_6;
	wire[1:0] w_n279_7;
	wire[2:0] w_n281_0;
	wire[1:0] w_n281_1;
	wire[2:0] w_n282_0;
	wire[2:0] w_n282_1;
	wire[2:0] w_n282_2;
	wire[2:0] w_n282_3;
	wire[2:0] w_n282_4;
	wire[2:0] w_n282_5;
	wire[2:0] w_n282_6;
	wire[1:0] w_n282_7;
	wire[2:0] w_n284_0;
	wire[2:0] w_n284_1;
	wire[2:0] w_n284_2;
	wire[2:0] w_n284_3;
	wire[2:0] w_n284_4;
	wire[2:0] w_n284_5;
	wire[2:0] w_n284_6;
	wire[1:0] w_n284_7;
	wire[2:0] w_n286_0;
	wire[1:0] w_n286_1;
	wire[2:0] w_n287_0;
	wire[2:0] w_n287_1;
	wire[2:0] w_n287_2;
	wire[2:0] w_n287_3;
	wire[2:0] w_n287_4;
	wire[2:0] w_n287_5;
	wire[2:0] w_n287_6;
	wire[1:0] w_n287_7;
	wire[2:0] w_n289_0;
	wire[1:0] w_n289_1;
	wire[2:0] w_n290_0;
	wire[2:0] w_n290_1;
	wire[2:0] w_n290_2;
	wire[2:0] w_n290_3;
	wire[2:0] w_n290_4;
	wire[2:0] w_n290_5;
	wire[2:0] w_n290_6;
	wire[1:0] w_n290_7;
	wire[2:0] w_n292_0;
	wire[2:0] w_n292_1;
	wire[2:0] w_n292_2;
	wire[2:0] w_n292_3;
	wire[2:0] w_n292_4;
	wire[2:0] w_n292_5;
	wire[2:0] w_n292_6;
	wire[1:0] w_n292_7;
	wire[2:0] w_n294_0;
	wire[2:0] w_n294_1;
	wire[2:0] w_n294_2;
	wire[2:0] w_n294_3;
	wire[2:0] w_n294_4;
	wire[2:0] w_n294_5;
	wire[2:0] w_n294_6;
	wire[1:0] w_n294_7;
	wire[2:0] w_n296_0;
	wire[1:0] w_n296_1;
	wire[2:0] w_n297_0;
	wire[2:0] w_n297_1;
	wire[2:0] w_n297_2;
	wire[2:0] w_n297_3;
	wire[2:0] w_n297_4;
	wire[2:0] w_n297_5;
	wire[2:0] w_n297_6;
	wire[1:0] w_n297_7;
	wire[2:0] w_n299_0;
	wire[2:0] w_n299_1;
	wire[2:0] w_n299_2;
	wire[2:0] w_n299_3;
	wire[2:0] w_n299_4;
	wire[2:0] w_n299_5;
	wire[2:0] w_n299_6;
	wire[1:0] w_n299_7;
	wire[2:0] w_n301_0;
	wire[1:0] w_n301_1;
	wire[2:0] w_n302_0;
	wire[2:0] w_n302_1;
	wire[2:0] w_n302_2;
	wire[2:0] w_n302_3;
	wire[2:0] w_n302_4;
	wire[2:0] w_n302_5;
	wire[2:0] w_n302_6;
	wire[1:0] w_n302_7;
	wire[2:0] w_n304_0;
	wire[2:0] w_n304_1;
	wire[2:0] w_n304_2;
	wire[2:0] w_n304_3;
	wire[2:0] w_n304_4;
	wire[2:0] w_n304_5;
	wire[2:0] w_n304_6;
	wire[1:0] w_n304_7;
	wire[2:0] w_n306_0;
	wire[2:0] w_n306_1;
	wire[2:0] w_n306_2;
	wire[2:0] w_n306_3;
	wire[2:0] w_n306_4;
	wire[2:0] w_n306_5;
	wire[2:0] w_n306_6;
	wire[1:0] w_n306_7;
	wire[2:0] w_n308_0;
	wire[2:0] w_n308_1;
	wire[2:0] w_n308_2;
	wire[2:0] w_n308_3;
	wire[2:0] w_n308_4;
	wire[2:0] w_n308_5;
	wire[2:0] w_n308_6;
	wire[1:0] w_n308_7;
	wire[2:0] w_n310_0;
	wire[2:0] w_n310_1;
	wire[2:0] w_n310_2;
	wire[2:0] w_n310_3;
	wire[2:0] w_n310_4;
	wire[2:0] w_n310_5;
	wire[2:0] w_n310_6;
	wire[1:0] w_n310_7;
	wire[2:0] w_n312_0;
	wire[2:0] w_n312_1;
	wire[2:0] w_n312_2;
	wire[2:0] w_n312_3;
	wire[2:0] w_n312_4;
	wire[2:0] w_n312_5;
	wire[2:0] w_n312_6;
	wire[1:0] w_n312_7;
	wire[2:0] w_n314_0;
	wire[1:0] w_n314_1;
	wire[2:0] w_n315_0;
	wire[2:0] w_n315_1;
	wire[2:0] w_n315_2;
	wire[2:0] w_n315_3;
	wire[2:0] w_n315_4;
	wire[2:0] w_n315_5;
	wire[2:0] w_n315_6;
	wire[1:0] w_n315_7;
	wire[2:0] w_n332_0;
	wire[1:0] w_n332_1;
	wire[2:0] w_n333_0;
	wire[2:0] w_n333_1;
	wire[2:0] w_n333_2;
	wire[2:0] w_n333_3;
	wire[2:0] w_n333_4;
	wire[2:0] w_n333_5;
	wire[2:0] w_n333_6;
	wire[1:0] w_n333_7;
	wire[2:0] w_n350_0;
	wire[1:0] w_n350_1;
	wire[2:0] w_n351_0;
	wire[2:0] w_n351_1;
	wire[2:0] w_n351_2;
	wire[2:0] w_n351_3;
	wire[2:0] w_n351_4;
	wire[2:0] w_n351_5;
	wire[2:0] w_n351_6;
	wire[1:0] w_n351_7;
	wire[2:0] w_n368_0;
	wire[1:0] w_n368_1;
	wire[2:0] w_n369_0;
	wire[2:0] w_n369_1;
	wire[2:0] w_n369_2;
	wire[2:0] w_n369_3;
	wire[2:0] w_n369_4;
	wire[2:0] w_n369_5;
	wire[2:0] w_n369_6;
	wire[1:0] w_n369_7;
	wire[2:0] w_n386_0;
	wire[2:0] w_n386_1;
	wire[2:0] w_n386_2;
	wire[2:0] w_n386_3;
	wire[2:0] w_n386_4;
	wire[2:0] w_n386_5;
	wire[2:0] w_n386_6;
	wire[1:0] w_n386_7;
	wire[2:0] w_n403_0;
	wire[2:0] w_n403_1;
	wire[2:0] w_n403_2;
	wire[2:0] w_n403_3;
	wire[2:0] w_n403_4;
	wire[2:0] w_n403_5;
	wire[2:0] w_n403_6;
	wire[1:0] w_n403_7;
	wire[2:0] w_n420_0;
	wire[2:0] w_n420_1;
	wire[2:0] w_n420_2;
	wire[2:0] w_n420_3;
	wire[2:0] w_n420_4;
	wire[2:0] w_n420_5;
	wire[2:0] w_n420_6;
	wire[1:0] w_n420_7;
	wire[1:0] w_n437_0;
	wire[2:0] w_n438_0;
	wire[1:0] w_n438_1;
	wire[2:0] w_n439_0;
	wire[2:0] w_n439_1;
	wire[2:0] w_n439_2;
	wire[2:0] w_n439_3;
	wire[2:0] w_n439_4;
	wire[2:0] w_n439_5;
	wire[2:0] w_n439_6;
	wire[1:0] w_n439_7;
	wire[2:0] w_n456_0;
	wire[2:0] w_n456_1;
	wire[2:0] w_n456_2;
	wire[2:0] w_n456_3;
	wire[2:0] w_n456_4;
	wire[2:0] w_n456_5;
	wire[2:0] w_n456_6;
	wire[1:0] w_n456_7;
	wire[2:0] w_n473_0;
	wire[2:0] w_n473_1;
	wire[2:0] w_n473_2;
	wire[2:0] w_n473_3;
	wire[2:0] w_n473_4;
	wire[2:0] w_n473_5;
	wire[2:0] w_n473_6;
	wire[1:0] w_n473_7;
	wire[2:0] w_n490_0;
	wire[2:0] w_n490_1;
	wire[2:0] w_n490_2;
	wire[2:0] w_n490_3;
	wire[2:0] w_n490_4;
	wire[2:0] w_n490_5;
	wire[2:0] w_n490_6;
	wire[1:0] w_n490_7;
	wire[2:0] w_n507_0;
	wire[1:0] w_n507_1;
	wire[2:0] w_n508_0;
	wire[2:0] w_n508_1;
	wire[2:0] w_n508_2;
	wire[2:0] w_n508_3;
	wire[2:0] w_n508_4;
	wire[2:0] w_n508_5;
	wire[2:0] w_n508_6;
	wire[1:0] w_n508_7;
	wire[2:0] w_n525_0;
	wire[2:0] w_n525_1;
	wire[2:0] w_n525_2;
	wire[2:0] w_n525_3;
	wire[2:0] w_n525_4;
	wire[2:0] w_n525_5;
	wire[2:0] w_n525_6;
	wire[1:0] w_n525_7;
	wire[2:0] w_n542_0;
	wire[2:0] w_n542_1;
	wire[2:0] w_n542_2;
	wire[2:0] w_n542_3;
	wire[2:0] w_n542_4;
	wire[2:0] w_n542_5;
	wire[2:0] w_n542_6;
	wire[1:0] w_n542_7;
	wire[2:0] w_n559_0;
	wire[2:0] w_n559_1;
	wire[2:0] w_n559_2;
	wire[2:0] w_n559_3;
	wire[2:0] w_n559_4;
	wire[2:0] w_n559_5;
	wire[2:0] w_n559_6;
	wire[1:0] w_n559_7;
	wire w_dff_A_Gf2kgLWc7_0;
	wire w_dff_A_6pXnAQTl5_2;
	wire w_dff_A_qjAdWqQ03_0;
	wire w_dff_A_060PweF86_2;
	wire w_dff_A_x9tybVmZ8_1;
	wire w_dff_A_hXKPEsEE7_2;
	wire w_dff_A_Ly8npyZr5_0;
	wire w_dff_A_egJSvUHp6_2;
	wire w_dff_A_J4cuJkSl9_1;
	wire w_dff_A_hkly1Ioj9_2;
	wire w_dff_A_oBp7Jqop7_2;
	jnot g000(.din(w_count4_0[2]),.dout(n264),.clk(gclk));
	jnot g001(.din(w_count5_0[2]),.dout(n265),.clk(gclk));
	jand g002(.dina(w_n265_0[1]),.dinb(w_n264_0[1]),.dout(n266),.clk(gclk));
	jnot g003(.din(w_count6_0[2]),.dout(n267),.clk(gclk));
	jand g004(.dina(w_count7_0[2]),.dinb(w_n267_0[1]),.dout(n268),.clk(gclk));
	jand g005(.dina(w_n268_1[1]),.dinb(w_n266_1[1]),.dout(n269),.clk(gclk));
	jnot g006(.din(w_count0_0[2]),.dout(n270),.clk(gclk));
	jnot g007(.din(w_count2_0[2]),.dout(n271),.clk(gclk));
	jand g008(.dina(w_n271_0[1]),.dinb(w_n270_0[1]),.dout(n272),.clk(gclk));
	jnot g009(.din(w_count1_0[2]),.dout(n273),.clk(gclk));
	jnot g010(.din(w_count3_0[2]),.dout(n274),.clk(gclk));
	jand g011(.dina(w_n274_0[1]),.dinb(w_n273_0[1]),.dout(n275),.clk(gclk));
	jand g012(.dina(w_n275_1[1]),.dinb(w_n272_1[1]),.dout(n276),.clk(gclk));
	jand g013(.dina(w_n276_7[1]),.dinb(w_n269_7[1]),.dout(selectp10),.clk(gclk));
	jand g014(.dina(w_n271_0[0]),.dinb(w_count0_0[1]),.dout(n278),.clk(gclk));
	jand g015(.dina(w_n278_1[1]),.dinb(w_n275_1[0]),.dout(n279),.clk(gclk));
	jand g016(.dina(w_n279_7[1]),.dinb(w_n269_7[0]),.dout(selectp11),.clk(gclk));
	jand g017(.dina(w_n274_0[0]),.dinb(w_count1_0[1]),.dout(n281),.clk(gclk));
	jand g018(.dina(w_n281_1[1]),.dinb(w_n272_1[0]),.dout(n282),.clk(gclk));
	jand g019(.dina(w_n282_7[1]),.dinb(w_n269_6[2]),.dout(selectp12),.clk(gclk));
	jand g020(.dina(w_n281_1[0]),.dinb(w_n278_1[0]),.dout(n284),.clk(gclk));
	jand g021(.dina(w_n284_7[1]),.dinb(w_n269_6[1]),.dout(selectp13),.clk(gclk));
	jand g022(.dina(w_count2_0[1]),.dinb(w_n270_0[0]),.dout(n286),.clk(gclk));
	jand g023(.dina(w_n286_1[1]),.dinb(w_n275_0[2]),.dout(n287),.clk(gclk));
	jand g024(.dina(w_n287_7[1]),.dinb(w_n269_6[0]),.dout(selectp14),.clk(gclk));
	jand g025(.dina(w_count2_0[0]),.dinb(w_count0_0[0]),.dout(n289),.clk(gclk));
	jand g026(.dina(w_n289_1[1]),.dinb(w_n275_0[1]),.dout(n290),.clk(gclk));
	jand g027(.dina(w_n290_7[1]),.dinb(w_n269_5[2]),.dout(selectp15),.clk(gclk));
	jand g028(.dina(w_n286_1[0]),.dinb(w_n281_0[2]),.dout(n292),.clk(gclk));
	jand g029(.dina(w_n292_7[1]),.dinb(w_n269_5[1]),.dout(selectp16),.clk(gclk));
	jand g030(.dina(w_n289_1[0]),.dinb(w_n281_0[1]),.dout(n294),.clk(gclk));
	jand g031(.dina(w_n294_7[1]),.dinb(w_n269_5[0]),.dout(selectp17),.clk(gclk));
	jand g032(.dina(w_count3_0[1]),.dinb(w_n273_0[0]),.dout(n296),.clk(gclk));
	jand g033(.dina(w_n296_1[1]),.dinb(w_n272_0[2]),.dout(n297),.clk(gclk));
	jand g034(.dina(w_n297_7[1]),.dinb(w_n269_4[2]),.dout(selectp18),.clk(gclk));
	jand g035(.dina(w_n296_1[0]),.dinb(w_n278_0[2]),.dout(n299),.clk(gclk));
	jand g036(.dina(w_n299_7[1]),.dinb(w_n269_4[1]),.dout(selectp19),.clk(gclk));
	jand g037(.dina(w_count3_0[0]),.dinb(w_count1_0[0]),.dout(n301),.clk(gclk));
	jand g038(.dina(w_n301_1[1]),.dinb(w_n272_0[1]),.dout(n302),.clk(gclk));
	jand g039(.dina(w_n302_7[1]),.dinb(w_n269_4[0]),.dout(selectp110),.clk(gclk));
	jand g040(.dina(w_n301_1[0]),.dinb(w_n278_0[1]),.dout(n304),.clk(gclk));
	jand g041(.dina(w_n304_7[1]),.dinb(w_n269_3[2]),.dout(selectp111),.clk(gclk));
	jand g042(.dina(w_n296_0[2]),.dinb(w_n286_0[2]),.dout(n306),.clk(gclk));
	jand g043(.dina(w_n306_7[1]),.dinb(w_n269_3[1]),.dout(selectp112),.clk(gclk));
	jand g044(.dina(w_n296_0[1]),.dinb(w_n289_0[2]),.dout(n308),.clk(gclk));
	jand g045(.dina(w_n308_7[1]),.dinb(w_n269_3[0]),.dout(selectp113),.clk(gclk));
	jand g046(.dina(w_n301_0[2]),.dinb(w_n286_0[1]),.dout(n310),.clk(gclk));
	jand g047(.dina(w_n310_7[1]),.dinb(w_n269_2[2]),.dout(selectp114),.clk(gclk));
	jand g048(.dina(w_n301_0[1]),.dinb(w_n289_0[1]),.dout(n312),.clk(gclk));
	jand g049(.dina(w_n312_7[1]),.dinb(w_n269_2[1]),.dout(selectp115),.clk(gclk));
	jand g050(.dina(w_n265_0[0]),.dinb(w_count4_0[1]),.dout(n314),.clk(gclk));
	jand g051(.dina(w_n314_1[1]),.dinb(w_n268_1[0]),.dout(n315),.clk(gclk));
	jand g052(.dina(w_n315_7[1]),.dinb(w_n276_7[0]),.dout(selectp116),.clk(gclk));
	jand g053(.dina(w_n315_7[0]),.dinb(w_n279_7[0]),.dout(selectp117),.clk(gclk));
	jand g054(.dina(w_n315_6[2]),.dinb(w_n282_7[0]),.dout(selectp118),.clk(gclk));
	jand g055(.dina(w_n315_6[1]),.dinb(w_n284_7[0]),.dout(selectp119),.clk(gclk));
	jand g056(.dina(w_n315_6[0]),.dinb(w_n287_7[0]),.dout(selectp120),.clk(gclk));
	jand g057(.dina(w_n315_5[2]),.dinb(w_n290_7[0]),.dout(selectp121),.clk(gclk));
	jand g058(.dina(w_n315_5[1]),.dinb(w_n292_7[0]),.dout(selectp122),.clk(gclk));
	jand g059(.dina(w_n315_5[0]),.dinb(w_n294_7[0]),.dout(selectp123),.clk(gclk));
	jand g060(.dina(w_n315_4[2]),.dinb(w_n297_7[0]),.dout(selectp124),.clk(gclk));
	jand g061(.dina(w_n315_4[1]),.dinb(w_n299_7[0]),.dout(selectp125),.clk(gclk));
	jand g062(.dina(w_n315_4[0]),.dinb(w_n302_7[0]),.dout(selectp126),.clk(gclk));
	jand g063(.dina(w_n315_3[2]),.dinb(w_n304_7[0]),.dout(selectp127),.clk(gclk));
	jand g064(.dina(w_n315_3[1]),.dinb(w_n306_7[0]),.dout(selectp128),.clk(gclk));
	jand g065(.dina(w_n315_3[0]),.dinb(w_n308_7[0]),.dout(selectp129),.clk(gclk));
	jand g066(.dina(w_n315_2[2]),.dinb(w_n310_7[0]),.dout(selectp130),.clk(gclk));
	jand g067(.dina(w_n315_2[1]),.dinb(w_n312_7[0]),.dout(selectp131),.clk(gclk));
	jand g068(.dina(w_count5_0[1]),.dinb(w_n264_0[0]),.dout(n332),.clk(gclk));
	jand g069(.dina(w_n332_1[1]),.dinb(w_n268_0[2]),.dout(n333),.clk(gclk));
	jand g070(.dina(w_n333_7[1]),.dinb(w_n276_6[2]),.dout(selectp132),.clk(gclk));
	jand g071(.dina(w_n333_7[0]),.dinb(w_n279_6[2]),.dout(selectp133),.clk(gclk));
	jand g072(.dina(w_n333_6[2]),.dinb(w_n282_6[2]),.dout(selectp134),.clk(gclk));
	jand g073(.dina(w_n333_6[1]),.dinb(w_n284_6[2]),.dout(selectp135),.clk(gclk));
	jand g074(.dina(w_n333_6[0]),.dinb(w_n287_6[2]),.dout(selectp136),.clk(gclk));
	jand g075(.dina(w_n333_5[2]),.dinb(w_n290_6[2]),.dout(selectp137),.clk(gclk));
	jand g076(.dina(w_n333_5[1]),.dinb(w_n292_6[2]),.dout(selectp138),.clk(gclk));
	jand g077(.dina(w_n333_5[0]),.dinb(w_n294_6[2]),.dout(selectp139),.clk(gclk));
	jand g078(.dina(w_n333_4[2]),.dinb(w_n297_6[2]),.dout(selectp140),.clk(gclk));
	jand g079(.dina(w_n333_4[1]),.dinb(w_n299_6[2]),.dout(selectp141),.clk(gclk));
	jand g080(.dina(w_n333_4[0]),.dinb(w_n302_6[2]),.dout(selectp142),.clk(gclk));
	jand g081(.dina(w_n333_3[2]),.dinb(w_n304_6[2]),.dout(selectp143),.clk(gclk));
	jand g082(.dina(w_n333_3[1]),.dinb(w_n306_6[2]),.dout(selectp144),.clk(gclk));
	jand g083(.dina(w_n333_3[0]),.dinb(w_n308_6[2]),.dout(selectp145),.clk(gclk));
	jand g084(.dina(w_n333_2[2]),.dinb(w_n310_6[2]),.dout(selectp146),.clk(gclk));
	jand g085(.dina(w_n333_2[1]),.dinb(w_n312_6[2]),.dout(selectp147),.clk(gclk));
	jand g086(.dina(w_count5_0[0]),.dinb(w_count4_0[0]),.dout(n350),.clk(gclk));
	jand g087(.dina(w_n350_1[1]),.dinb(w_n268_0[1]),.dout(n351),.clk(gclk));
	jand g088(.dina(w_n351_7[1]),.dinb(w_n276_6[1]),.dout(selectp148),.clk(gclk));
	jand g089(.dina(w_n351_7[0]),.dinb(w_n279_6[1]),.dout(selectp149),.clk(gclk));
	jand g090(.dina(w_n351_6[2]),.dinb(w_n282_6[1]),.dout(selectp150),.clk(gclk));
	jand g091(.dina(w_n351_6[1]),.dinb(w_n284_6[1]),.dout(selectp151),.clk(gclk));
	jand g092(.dina(w_n351_6[0]),.dinb(w_n287_6[1]),.dout(selectp152),.clk(gclk));
	jand g093(.dina(w_n351_5[2]),.dinb(w_n290_6[1]),.dout(selectp153),.clk(gclk));
	jand g094(.dina(w_n351_5[1]),.dinb(w_n292_6[1]),.dout(selectp154),.clk(gclk));
	jand g095(.dina(w_n351_5[0]),.dinb(w_n294_6[1]),.dout(selectp155),.clk(gclk));
	jand g096(.dina(w_n351_4[2]),.dinb(w_n297_6[1]),.dout(selectp156),.clk(gclk));
	jand g097(.dina(w_n351_4[1]),.dinb(w_n299_6[1]),.dout(selectp157),.clk(gclk));
	jand g098(.dina(w_n351_4[0]),.dinb(w_n302_6[1]),.dout(selectp158),.clk(gclk));
	jand g099(.dina(w_n351_3[2]),.dinb(w_n304_6[1]),.dout(selectp159),.clk(gclk));
	jand g100(.dina(w_n351_3[1]),.dinb(w_n306_6[1]),.dout(selectp160),.clk(gclk));
	jand g101(.dina(w_n351_3[0]),.dinb(w_n308_6[1]),.dout(selectp161),.clk(gclk));
	jand g102(.dina(w_n351_2[2]),.dinb(w_n310_6[1]),.dout(selectp162),.clk(gclk));
	jand g103(.dina(w_n351_2[1]),.dinb(w_n312_6[1]),.dout(selectp163),.clk(gclk));
	jand g104(.dina(w_count7_0[1]),.dinb(w_count6_0[1]),.dout(n368),.clk(gclk));
	jand g105(.dina(w_n368_1[1]),.dinb(w_n266_1[0]),.dout(n369),.clk(gclk));
	jand g106(.dina(w_n369_7[1]),.dinb(w_n276_6[0]),.dout(selectp164),.clk(gclk));
	jand g107(.dina(w_n369_7[0]),.dinb(w_n279_6[0]),.dout(selectp165),.clk(gclk));
	jand g108(.dina(w_n369_6[2]),.dinb(w_n282_6[0]),.dout(selectp166),.clk(gclk));
	jand g109(.dina(w_n369_6[1]),.dinb(w_n284_6[0]),.dout(selectp167),.clk(gclk));
	jand g110(.dina(w_n369_6[0]),.dinb(w_n287_6[0]),.dout(selectp168),.clk(gclk));
	jand g111(.dina(w_n369_5[2]),.dinb(w_n290_6[0]),.dout(selectp169),.clk(gclk));
	jand g112(.dina(w_n369_5[1]),.dinb(w_n292_6[0]),.dout(selectp170),.clk(gclk));
	jand g113(.dina(w_n369_5[0]),.dinb(w_n294_6[0]),.dout(selectp171),.clk(gclk));
	jand g114(.dina(w_n369_4[2]),.dinb(w_n297_6[0]),.dout(selectp172),.clk(gclk));
	jand g115(.dina(w_n369_4[1]),.dinb(w_n299_6[0]),.dout(selectp173),.clk(gclk));
	jand g116(.dina(w_n369_4[0]),.dinb(w_n302_6[0]),.dout(selectp174),.clk(gclk));
	jand g117(.dina(w_n369_3[2]),.dinb(w_n304_6[0]),.dout(selectp175),.clk(gclk));
	jand g118(.dina(w_n369_3[1]),.dinb(w_n306_6[0]),.dout(selectp176),.clk(gclk));
	jand g119(.dina(w_n369_3[0]),.dinb(w_n308_6[0]),.dout(selectp177),.clk(gclk));
	jand g120(.dina(w_n369_2[2]),.dinb(w_n310_6[0]),.dout(selectp178),.clk(gclk));
	jand g121(.dina(w_n369_2[1]),.dinb(w_n312_6[0]),.dout(selectp179),.clk(gclk));
	jand g122(.dina(w_n368_1[0]),.dinb(w_n314_1[0]),.dout(n386),.clk(gclk));
	jand g123(.dina(w_n386_7[1]),.dinb(w_n276_5[2]),.dout(selectp180),.clk(gclk));
	jand g124(.dina(w_n386_7[0]),.dinb(w_n279_5[2]),.dout(selectp181),.clk(gclk));
	jand g125(.dina(w_n386_6[2]),.dinb(w_n282_5[2]),.dout(selectp182),.clk(gclk));
	jand g126(.dina(w_n386_6[1]),.dinb(w_n284_5[2]),.dout(selectp183),.clk(gclk));
	jand g127(.dina(w_n386_6[0]),.dinb(w_n287_5[2]),.dout(selectp184),.clk(gclk));
	jand g128(.dina(w_n386_5[2]),.dinb(w_n290_5[2]),.dout(selectp185),.clk(gclk));
	jand g129(.dina(w_n386_5[1]),.dinb(w_n292_5[2]),.dout(selectp186),.clk(gclk));
	jand g130(.dina(w_n386_5[0]),.dinb(w_n294_5[2]),.dout(selectp187),.clk(gclk));
	jand g131(.dina(w_n386_4[2]),.dinb(w_n297_5[2]),.dout(selectp188),.clk(gclk));
	jand g132(.dina(w_n386_4[1]),.dinb(w_n299_5[2]),.dout(selectp189),.clk(gclk));
	jand g133(.dina(w_n386_4[0]),.dinb(w_n302_5[2]),.dout(selectp190),.clk(gclk));
	jand g134(.dina(w_n386_3[2]),.dinb(w_n304_5[2]),.dout(selectp191),.clk(gclk));
	jand g135(.dina(w_n386_3[1]),.dinb(w_n306_5[2]),.dout(selectp192),.clk(gclk));
	jand g136(.dina(w_n386_3[0]),.dinb(w_n308_5[2]),.dout(selectp193),.clk(gclk));
	jand g137(.dina(w_n386_2[2]),.dinb(w_n310_5[2]),.dout(selectp194),.clk(gclk));
	jand g138(.dina(w_n386_2[1]),.dinb(w_n312_5[2]),.dout(selectp195),.clk(gclk));
	jand g139(.dina(w_n368_0[2]),.dinb(w_n332_1[0]),.dout(n403),.clk(gclk));
	jand g140(.dina(w_n403_7[1]),.dinb(w_n276_5[1]),.dout(selectp196),.clk(gclk));
	jand g141(.dina(w_n403_7[0]),.dinb(w_n279_5[1]),.dout(selectp197),.clk(gclk));
	jand g142(.dina(w_n403_6[2]),.dinb(w_n282_5[1]),.dout(selectp198),.clk(gclk));
	jand g143(.dina(w_n403_6[1]),.dinb(w_n284_5[1]),.dout(selectp199),.clk(gclk));
	jand g144(.dina(w_n403_6[0]),.dinb(w_n287_5[1]),.dout(selectp1100),.clk(gclk));
	jand g145(.dina(w_n403_5[2]),.dinb(w_n290_5[1]),.dout(selectp1101),.clk(gclk));
	jand g146(.dina(w_n403_5[1]),.dinb(w_n292_5[1]),.dout(selectp1102),.clk(gclk));
	jand g147(.dina(w_n403_5[0]),.dinb(w_n294_5[1]),.dout(selectp1103),.clk(gclk));
	jand g148(.dina(w_n403_4[2]),.dinb(w_n297_5[1]),.dout(selectp1104),.clk(gclk));
	jand g149(.dina(w_n403_4[1]),.dinb(w_n299_5[1]),.dout(selectp1105),.clk(gclk));
	jand g150(.dina(w_n403_4[0]),.dinb(w_n302_5[1]),.dout(selectp1106),.clk(gclk));
	jand g151(.dina(w_n403_3[2]),.dinb(w_n304_5[1]),.dout(selectp1107),.clk(gclk));
	jand g152(.dina(w_n403_3[1]),.dinb(w_n306_5[1]),.dout(selectp1108),.clk(gclk));
	jand g153(.dina(w_n403_3[0]),.dinb(w_n308_5[1]),.dout(selectp1109),.clk(gclk));
	jand g154(.dina(w_n403_2[2]),.dinb(w_n310_5[1]),.dout(selectp1110),.clk(gclk));
	jand g155(.dina(w_n403_2[1]),.dinb(w_n312_5[1]),.dout(selectp1111),.clk(gclk));
	jand g156(.dina(w_n368_0[1]),.dinb(w_n350_1[0]),.dout(n420),.clk(gclk));
	jand g157(.dina(w_n420_7[1]),.dinb(w_n276_5[0]),.dout(selectp1112),.clk(gclk));
	jand g158(.dina(w_n420_7[0]),.dinb(w_n279_5[0]),.dout(selectp1113),.clk(gclk));
	jand g159(.dina(w_n420_6[2]),.dinb(w_n282_5[0]),.dout(selectp1114),.clk(gclk));
	jand g160(.dina(w_n420_6[1]),.dinb(w_n284_5[0]),.dout(selectp1115),.clk(gclk));
	jand g161(.dina(w_n420_6[0]),.dinb(w_n287_5[0]),.dout(selectp1116),.clk(gclk));
	jand g162(.dina(w_n420_5[2]),.dinb(w_n290_5[0]),.dout(selectp1117),.clk(gclk));
	jand g163(.dina(w_n420_5[1]),.dinb(w_n292_5[0]),.dout(selectp1118),.clk(gclk));
	jand g164(.dina(w_n420_5[0]),.dinb(w_n294_5[0]),.dout(selectp1119),.clk(gclk));
	jand g165(.dina(w_n420_4[2]),.dinb(w_n297_5[0]),.dout(selectp1120),.clk(gclk));
	jand g166(.dina(w_n420_4[1]),.dinb(w_n299_5[0]),.dout(selectp1121),.clk(gclk));
	jand g167(.dina(w_n420_4[0]),.dinb(w_n302_5[0]),.dout(selectp1122),.clk(gclk));
	jand g168(.dina(w_n420_3[2]),.dinb(w_n304_5[0]),.dout(selectp1123),.clk(gclk));
	jand g169(.dina(w_n420_3[1]),.dinb(w_n306_5[0]),.dout(selectp1124),.clk(gclk));
	jand g170(.dina(w_n420_3[0]),.dinb(w_n308_5[0]),.dout(selectp1125),.clk(gclk));
	jand g171(.dina(w_n420_2[2]),.dinb(w_n310_5[0]),.dout(selectp1126),.clk(gclk));
	jand g172(.dina(w_n420_2[1]),.dinb(w_n312_5[0]),.dout(w_dff_A_oBp7Jqop7_2),.clk(gclk));
	jnot g173(.din(w_count7_0[0]),.dout(n437),.clk(gclk));
	jand g174(.dina(w_n437_0[1]),.dinb(w_n267_0[0]),.dout(n438),.clk(gclk));
	jand g175(.dina(w_n438_1[1]),.dinb(w_n266_0[2]),.dout(n439),.clk(gclk));
	jand g176(.dina(w_n439_7[1]),.dinb(w_n276_4[2]),.dout(selectp20),.clk(gclk));
	jand g177(.dina(w_n439_7[0]),.dinb(w_n279_4[2]),.dout(selectp21),.clk(gclk));
	jand g178(.dina(w_n439_6[2]),.dinb(w_n282_4[2]),.dout(selectp22),.clk(gclk));
	jand g179(.dina(w_n439_6[1]),.dinb(w_n284_4[2]),.dout(selectp23),.clk(gclk));
	jand g180(.dina(w_n439_6[0]),.dinb(w_n287_4[2]),.dout(selectp24),.clk(gclk));
	jand g181(.dina(w_n439_5[2]),.dinb(w_n290_4[2]),.dout(selectp25),.clk(gclk));
	jand g182(.dina(w_n439_5[1]),.dinb(w_n292_4[2]),.dout(selectp26),.clk(gclk));
	jand g183(.dina(w_n439_5[0]),.dinb(w_n294_4[2]),.dout(selectp27),.clk(gclk));
	jand g184(.dina(w_n439_4[2]),.dinb(w_n297_4[2]),.dout(selectp28),.clk(gclk));
	jand g185(.dina(w_n439_4[1]),.dinb(w_n299_4[2]),.dout(selectp29),.clk(gclk));
	jand g186(.dina(w_n439_4[0]),.dinb(w_n302_4[2]),.dout(selectp210),.clk(gclk));
	jand g187(.dina(w_n439_3[2]),.dinb(w_n304_4[2]),.dout(selectp211),.clk(gclk));
	jand g188(.dina(w_n439_3[1]),.dinb(w_n306_4[2]),.dout(selectp212),.clk(gclk));
	jand g189(.dina(w_n439_3[0]),.dinb(w_n308_4[2]),.dout(selectp213),.clk(gclk));
	jand g190(.dina(w_n439_2[2]),.dinb(w_n310_4[2]),.dout(selectp214),.clk(gclk));
	jand g191(.dina(w_n439_2[1]),.dinb(w_n312_4[2]),.dout(selectp215),.clk(gclk));
	jand g192(.dina(w_n438_1[0]),.dinb(w_n314_0[2]),.dout(n456),.clk(gclk));
	jand g193(.dina(w_n456_7[1]),.dinb(w_n276_4[1]),.dout(selectp216),.clk(gclk));
	jand g194(.dina(w_n456_7[0]),.dinb(w_n279_4[1]),.dout(selectp217),.clk(gclk));
	jand g195(.dina(w_n456_6[2]),.dinb(w_n282_4[1]),.dout(selectp218),.clk(gclk));
	jand g196(.dina(w_n456_6[1]),.dinb(w_n284_4[1]),.dout(selectp219),.clk(gclk));
	jand g197(.dina(w_n456_6[0]),.dinb(w_n287_4[1]),.dout(selectp220),.clk(gclk));
	jand g198(.dina(w_n456_5[2]),.dinb(w_n290_4[1]),.dout(selectp221),.clk(gclk));
	jand g199(.dina(w_n456_5[1]),.dinb(w_n292_4[1]),.dout(selectp222),.clk(gclk));
	jand g200(.dina(w_n456_5[0]),.dinb(w_n294_4[1]),.dout(selectp223),.clk(gclk));
	jand g201(.dina(w_n456_4[2]),.dinb(w_n297_4[1]),.dout(selectp224),.clk(gclk));
	jand g202(.dina(w_n456_4[1]),.dinb(w_n299_4[1]),.dout(selectp225),.clk(gclk));
	jand g203(.dina(w_n456_4[0]),.dinb(w_n302_4[1]),.dout(selectp226),.clk(gclk));
	jand g204(.dina(w_n456_3[2]),.dinb(w_n304_4[1]),.dout(selectp227),.clk(gclk));
	jand g205(.dina(w_n456_3[1]),.dinb(w_n306_4[1]),.dout(selectp228),.clk(gclk));
	jand g206(.dina(w_n456_3[0]),.dinb(w_n308_4[1]),.dout(selectp229),.clk(gclk));
	jand g207(.dina(w_n456_2[2]),.dinb(w_n310_4[1]),.dout(selectp230),.clk(gclk));
	jand g208(.dina(w_n456_2[1]),.dinb(w_n312_4[1]),.dout(selectp231),.clk(gclk));
	jand g209(.dina(w_n438_0[2]),.dinb(w_n332_0[2]),.dout(n473),.clk(gclk));
	jand g210(.dina(w_n473_7[1]),.dinb(w_n276_4[0]),.dout(selectp232),.clk(gclk));
	jand g211(.dina(w_n473_7[0]),.dinb(w_n279_4[0]),.dout(selectp233),.clk(gclk));
	jand g212(.dina(w_n473_6[2]),.dinb(w_n282_4[0]),.dout(selectp234),.clk(gclk));
	jand g213(.dina(w_n473_6[1]),.dinb(w_n284_4[0]),.dout(selectp235),.clk(gclk));
	jand g214(.dina(w_n473_6[0]),.dinb(w_n287_4[0]),.dout(selectp236),.clk(gclk));
	jand g215(.dina(w_n473_5[2]),.dinb(w_n290_4[0]),.dout(selectp237),.clk(gclk));
	jand g216(.dina(w_n473_5[1]),.dinb(w_n292_4[0]),.dout(selectp238),.clk(gclk));
	jand g217(.dina(w_n473_5[0]),.dinb(w_n294_4[0]),.dout(selectp239),.clk(gclk));
	jand g218(.dina(w_n473_4[2]),.dinb(w_n297_4[0]),.dout(selectp240),.clk(gclk));
	jand g219(.dina(w_n473_4[1]),.dinb(w_n299_4[0]),.dout(selectp241),.clk(gclk));
	jand g220(.dina(w_n473_4[0]),.dinb(w_n302_4[0]),.dout(selectp242),.clk(gclk));
	jand g221(.dina(w_n473_3[2]),.dinb(w_n304_4[0]),.dout(selectp243),.clk(gclk));
	jand g222(.dina(w_n473_3[1]),.dinb(w_n306_4[0]),.dout(selectp244),.clk(gclk));
	jand g223(.dina(w_n473_3[0]),.dinb(w_n308_4[0]),.dout(selectp245),.clk(gclk));
	jand g224(.dina(w_n473_2[2]),.dinb(w_n310_4[0]),.dout(selectp246),.clk(gclk));
	jand g225(.dina(w_n473_2[1]),.dinb(w_n312_4[0]),.dout(selectp247),.clk(gclk));
	jand g226(.dina(w_n438_0[1]),.dinb(w_n350_0[2]),.dout(n490),.clk(gclk));
	jand g227(.dina(w_n490_7[1]),.dinb(w_n276_3[2]),.dout(selectp248),.clk(gclk));
	jand g228(.dina(w_n490_7[0]),.dinb(w_n279_3[2]),.dout(selectp249),.clk(gclk));
	jand g229(.dina(w_n490_6[2]),.dinb(w_n282_3[2]),.dout(selectp250),.clk(gclk));
	jand g230(.dina(w_n490_6[1]),.dinb(w_n284_3[2]),.dout(selectp251),.clk(gclk));
	jand g231(.dina(w_n490_6[0]),.dinb(w_n287_3[2]),.dout(selectp252),.clk(gclk));
	jand g232(.dina(w_n490_5[2]),.dinb(w_n290_3[2]),.dout(selectp253),.clk(gclk));
	jand g233(.dina(w_n490_5[1]),.dinb(w_n292_3[2]),.dout(selectp254),.clk(gclk));
	jand g234(.dina(w_n490_5[0]),.dinb(w_n294_3[2]),.dout(selectp255),.clk(gclk));
	jand g235(.dina(w_n490_4[2]),.dinb(w_n297_3[2]),.dout(selectp256),.clk(gclk));
	jand g236(.dina(w_n490_4[1]),.dinb(w_n299_3[2]),.dout(selectp257),.clk(gclk));
	jand g237(.dina(w_n490_4[0]),.dinb(w_n302_3[2]),.dout(selectp258),.clk(gclk));
	jand g238(.dina(w_n490_3[2]),.dinb(w_n304_3[2]),.dout(selectp259),.clk(gclk));
	jand g239(.dina(w_n490_3[1]),.dinb(w_n306_3[2]),.dout(selectp260),.clk(gclk));
	jand g240(.dina(w_n490_3[0]),.dinb(w_n308_3[2]),.dout(selectp261),.clk(gclk));
	jand g241(.dina(w_n490_2[2]),.dinb(w_n310_3[2]),.dout(selectp262),.clk(gclk));
	jand g242(.dina(w_n490_2[1]),.dinb(w_n312_3[2]),.dout(selectp263),.clk(gclk));
	jand g243(.dina(w_n437_0[0]),.dinb(w_count6_0[0]),.dout(n507),.clk(gclk));
	jand g244(.dina(w_n507_1[1]),.dinb(w_n266_0[1]),.dout(n508),.clk(gclk));
	jand g245(.dina(w_n508_7[1]),.dinb(w_n276_3[1]),.dout(selectp264),.clk(gclk));
	jand g246(.dina(w_n508_7[0]),.dinb(w_n279_3[1]),.dout(selectp265),.clk(gclk));
	jand g247(.dina(w_n508_6[2]),.dinb(w_n282_3[1]),.dout(selectp266),.clk(gclk));
	jand g248(.dina(w_n508_6[1]),.dinb(w_n284_3[1]),.dout(selectp267),.clk(gclk));
	jand g249(.dina(w_n508_6[0]),.dinb(w_n287_3[1]),.dout(selectp268),.clk(gclk));
	jand g250(.dina(w_n508_5[2]),.dinb(w_n290_3[1]),.dout(selectp269),.clk(gclk));
	jand g251(.dina(w_n508_5[1]),.dinb(w_n292_3[1]),.dout(selectp270),.clk(gclk));
	jand g252(.dina(w_n508_5[0]),.dinb(w_n294_3[1]),.dout(selectp271),.clk(gclk));
	jand g253(.dina(w_n508_4[2]),.dinb(w_n297_3[1]),.dout(selectp272),.clk(gclk));
	jand g254(.dina(w_n508_4[1]),.dinb(w_n299_3[1]),.dout(selectp273),.clk(gclk));
	jand g255(.dina(w_n508_4[0]),.dinb(w_n302_3[1]),.dout(selectp274),.clk(gclk));
	jand g256(.dina(w_n508_3[2]),.dinb(w_n304_3[1]),.dout(selectp275),.clk(gclk));
	jand g257(.dina(w_n508_3[1]),.dinb(w_n306_3[1]),.dout(selectp276),.clk(gclk));
	jand g258(.dina(w_n508_3[0]),.dinb(w_n308_3[1]),.dout(selectp277),.clk(gclk));
	jand g259(.dina(w_n508_2[2]),.dinb(w_n310_3[1]),.dout(selectp278),.clk(gclk));
	jand g260(.dina(w_n508_2[1]),.dinb(w_n312_3[1]),.dout(selectp279),.clk(gclk));
	jand g261(.dina(w_n507_1[0]),.dinb(w_n314_0[1]),.dout(n525),.clk(gclk));
	jand g262(.dina(w_n525_7[1]),.dinb(w_n276_3[0]),.dout(selectp280),.clk(gclk));
	jand g263(.dina(w_n525_7[0]),.dinb(w_n279_3[0]),.dout(selectp281),.clk(gclk));
	jand g264(.dina(w_n525_6[2]),.dinb(w_n282_3[0]),.dout(selectp282),.clk(gclk));
	jand g265(.dina(w_n525_6[1]),.dinb(w_n284_3[0]),.dout(selectp283),.clk(gclk));
	jand g266(.dina(w_n525_6[0]),.dinb(w_n287_3[0]),.dout(selectp284),.clk(gclk));
	jand g267(.dina(w_n525_5[2]),.dinb(w_n290_3[0]),.dout(selectp285),.clk(gclk));
	jand g268(.dina(w_n525_5[1]),.dinb(w_n292_3[0]),.dout(selectp286),.clk(gclk));
	jand g269(.dina(w_n525_5[0]),.dinb(w_n294_3[0]),.dout(selectp287),.clk(gclk));
	jand g270(.dina(w_n525_4[2]),.dinb(w_n297_3[0]),.dout(selectp288),.clk(gclk));
	jand g271(.dina(w_n525_4[1]),.dinb(w_n299_3[0]),.dout(selectp289),.clk(gclk));
	jand g272(.dina(w_n525_4[0]),.dinb(w_n302_3[0]),.dout(selectp290),.clk(gclk));
	jand g273(.dina(w_n525_3[2]),.dinb(w_n304_3[0]),.dout(selectp291),.clk(gclk));
	jand g274(.dina(w_n525_3[1]),.dinb(w_n306_3[0]),.dout(selectp292),.clk(gclk));
	jand g275(.dina(w_n525_3[0]),.dinb(w_n308_3[0]),.dout(selectp293),.clk(gclk));
	jand g276(.dina(w_n525_2[2]),.dinb(w_n310_3[0]),.dout(selectp294),.clk(gclk));
	jand g277(.dina(w_n525_2[1]),.dinb(w_n312_3[0]),.dout(selectp295),.clk(gclk));
	jand g278(.dina(w_n507_0[2]),.dinb(w_n332_0[1]),.dout(n542),.clk(gclk));
	jand g279(.dina(w_n542_7[1]),.dinb(w_n276_2[2]),.dout(selectp296),.clk(gclk));
	jand g280(.dina(w_n542_7[0]),.dinb(w_n279_2[2]),.dout(selectp297),.clk(gclk));
	jand g281(.dina(w_n542_6[2]),.dinb(w_n282_2[2]),.dout(selectp298),.clk(gclk));
	jand g282(.dina(w_n542_6[1]),.dinb(w_n284_2[2]),.dout(selectp299),.clk(gclk));
	jand g283(.dina(w_n542_6[0]),.dinb(w_n287_2[2]),.dout(selectp2100),.clk(gclk));
	jand g284(.dina(w_n542_5[2]),.dinb(w_n290_2[2]),.dout(selectp2101),.clk(gclk));
	jand g285(.dina(w_n542_5[1]),.dinb(w_n292_2[2]),.dout(selectp2102),.clk(gclk));
	jand g286(.dina(w_n542_5[0]),.dinb(w_n294_2[2]),.dout(selectp2103),.clk(gclk));
	jand g287(.dina(w_n542_4[2]),.dinb(w_n297_2[2]),.dout(selectp2104),.clk(gclk));
	jand g288(.dina(w_n542_4[1]),.dinb(w_n299_2[2]),.dout(selectp2105),.clk(gclk));
	jand g289(.dina(w_n542_4[0]),.dinb(w_n302_2[2]),.dout(selectp2106),.clk(gclk));
	jand g290(.dina(w_n542_3[2]),.dinb(w_n304_2[2]),.dout(selectp2107),.clk(gclk));
	jand g291(.dina(w_n542_3[1]),.dinb(w_n306_2[2]),.dout(selectp2108),.clk(gclk));
	jand g292(.dina(w_n542_3[0]),.dinb(w_n308_2[2]),.dout(selectp2109),.clk(gclk));
	jand g293(.dina(w_n542_2[2]),.dinb(w_n310_2[2]),.dout(selectp2110),.clk(gclk));
	jand g294(.dina(w_n542_2[1]),.dinb(w_n312_2[2]),.dout(selectp2111),.clk(gclk));
	jand g295(.dina(w_n507_0[1]),.dinb(w_n350_0[1]),.dout(n559),.clk(gclk));
	jand g296(.dina(w_n559_7[1]),.dinb(w_n276_2[1]),.dout(selectp2112),.clk(gclk));
	jand g297(.dina(w_n559_7[0]),.dinb(w_n279_2[1]),.dout(selectp2113),.clk(gclk));
	jand g298(.dina(w_n559_6[2]),.dinb(w_n282_2[1]),.dout(selectp2114),.clk(gclk));
	jand g299(.dina(w_n559_6[1]),.dinb(w_n284_2[1]),.dout(selectp2115),.clk(gclk));
	jand g300(.dina(w_n559_6[0]),.dinb(w_n287_2[1]),.dout(selectp2116),.clk(gclk));
	jand g301(.dina(w_n559_5[2]),.dinb(w_n290_2[1]),.dout(selectp2117),.clk(gclk));
	jand g302(.dina(w_n559_5[1]),.dinb(w_n292_2[1]),.dout(selectp2118),.clk(gclk));
	jand g303(.dina(w_n559_5[0]),.dinb(w_n294_2[1]),.dout(selectp2119),.clk(gclk));
	jand g304(.dina(w_n559_4[2]),.dinb(w_n297_2[1]),.dout(selectp2120),.clk(gclk));
	jand g305(.dina(w_n559_4[1]),.dinb(w_n299_2[1]),.dout(selectp2121),.clk(gclk));
	jand g306(.dina(w_n559_4[0]),.dinb(w_n302_2[1]),.dout(selectp2122),.clk(gclk));
	jand g307(.dina(w_n559_3[2]),.dinb(w_n304_2[1]),.dout(selectp2123),.clk(gclk));
	jand g308(.dina(w_n559_3[1]),.dinb(w_n306_2[1]),.dout(selectp2124),.clk(gclk));
	jand g309(.dina(w_n559_3[0]),.dinb(w_n308_2[1]),.dout(selectp2125),.clk(gclk));
	jand g310(.dina(w_n559_2[2]),.dinb(w_n310_2[1]),.dout(selectp2126),.clk(gclk));
	jand g311(.dina(w_n559_2[1]),.dinb(w_n312_2[1]),.dout(selectp2127),.clk(gclk));
	jspl3 jspl3_w_count0_0(.douta(w_count0_0[0]),.doutb(w_count0_0[1]),.doutc(w_count0_0[2]),.din(count0));
	jspl3 jspl3_w_count1_0(.douta(w_count1_0[0]),.doutb(w_count1_0[1]),.doutc(w_count1_0[2]),.din(count1));
	jspl3 jspl3_w_count2_0(.douta(w_count2_0[0]),.doutb(w_count2_0[1]),.doutc(w_count2_0[2]),.din(count2));
	jspl3 jspl3_w_count3_0(.douta(w_count3_0[0]),.doutb(w_count3_0[1]),.doutc(w_count3_0[2]),.din(count3));
	jspl3 jspl3_w_count4_0(.douta(w_count4_0[0]),.doutb(w_count4_0[1]),.doutc(w_count4_0[2]),.din(count4));
	jspl3 jspl3_w_count5_0(.douta(w_count5_0[0]),.doutb(w_count5_0[1]),.doutc(w_count5_0[2]),.din(count5));
	jspl3 jspl3_w_count6_0(.douta(w_count6_0[0]),.doutb(w_count6_0[1]),.doutc(w_count6_0[2]),.din(count6));
	jspl3 jspl3_w_count7_0(.douta(w_count7_0[0]),.doutb(w_count7_0[1]),.doutc(w_count7_0[2]),.din(count7));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(n265));
	jspl3 jspl3_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.doutc(w_n266_0[2]),.din(n266));
	jspl jspl_w_n266_1(.douta(w_n266_1[0]),.doutb(w_n266_1[1]),.din(w_n266_0[0]));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.doutc(w_n268_0[2]),.din(n268));
	jspl jspl_w_n268_1(.douta(w_n268_1[0]),.doutb(w_n268_1[1]),.din(w_n268_0[0]));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl3 jspl3_w_n269_2(.douta(w_n269_2[0]),.doutb(w_n269_2[1]),.doutc(w_n269_2[2]),.din(w_n269_0[1]));
	jspl3 jspl3_w_n269_3(.douta(w_n269_3[0]),.doutb(w_n269_3[1]),.doutc(w_n269_3[2]),.din(w_n269_0[2]));
	jspl3 jspl3_w_n269_4(.douta(w_n269_4[0]),.doutb(w_n269_4[1]),.doutc(w_n269_4[2]),.din(w_n269_1[0]));
	jspl3 jspl3_w_n269_5(.douta(w_n269_5[0]),.doutb(w_n269_5[1]),.doutc(w_n269_5[2]),.din(w_n269_1[1]));
	jspl3 jspl3_w_n269_6(.douta(w_n269_6[0]),.doutb(w_n269_6[1]),.doutc(w_n269_6[2]),.din(w_n269_1[2]));
	jspl jspl_w_n269_7(.douta(w_n269_7[0]),.doutb(w_n269_7[1]),.din(w_n269_2[0]));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.din(n271));
	jspl3 jspl3_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.doutc(w_n272_0[2]),.din(n272));
	jspl jspl_w_n272_1(.douta(w_n272_1[0]),.doutb(w_n272_1[1]),.din(w_n272_0[0]));
	jspl jspl_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl3 jspl3_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.doutc(w_n275_0[2]),.din(n275));
	jspl jspl_w_n275_1(.douta(w_n275_1[0]),.doutb(w_n275_1[1]),.din(w_n275_0[0]));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(n276));
	jspl3 jspl3_w_n276_1(.douta(w_n276_1[0]),.doutb(w_n276_1[1]),.doutc(w_n276_1[2]),.din(w_n276_0[0]));
	jspl3 jspl3_w_n276_2(.douta(w_n276_2[0]),.doutb(w_n276_2[1]),.doutc(w_n276_2[2]),.din(w_n276_0[1]));
	jspl3 jspl3_w_n276_3(.douta(w_n276_3[0]),.doutb(w_n276_3[1]),.doutc(w_n276_3[2]),.din(w_n276_0[2]));
	jspl3 jspl3_w_n276_4(.douta(w_n276_4[0]),.doutb(w_n276_4[1]),.doutc(w_n276_4[2]),.din(w_n276_1[0]));
	jspl3 jspl3_w_n276_5(.douta(w_n276_5[0]),.doutb(w_n276_5[1]),.doutc(w_n276_5[2]),.din(w_n276_1[1]));
	jspl3 jspl3_w_n276_6(.douta(w_n276_6[0]),.doutb(w_n276_6[1]),.doutc(w_n276_6[2]),.din(w_n276_1[2]));
	jspl jspl_w_n276_7(.douta(w_n276_7[0]),.doutb(w_n276_7[1]),.din(w_n276_2[0]));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_n278_0[2]),.din(n278));
	jspl jspl_w_n278_1(.douta(w_n278_1[0]),.doutb(w_n278_1[1]),.din(w_n278_0[0]));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl3 jspl3_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.doutc(w_n279_1[2]),.din(w_n279_0[0]));
	jspl3 jspl3_w_n279_2(.douta(w_n279_2[0]),.doutb(w_n279_2[1]),.doutc(w_n279_2[2]),.din(w_n279_0[1]));
	jspl3 jspl3_w_n279_3(.douta(w_n279_3[0]),.doutb(w_n279_3[1]),.doutc(w_n279_3[2]),.din(w_n279_0[2]));
	jspl3 jspl3_w_n279_4(.douta(w_n279_4[0]),.doutb(w_n279_4[1]),.doutc(w_n279_4[2]),.din(w_n279_1[0]));
	jspl3 jspl3_w_n279_5(.douta(w_n279_5[0]),.doutb(w_n279_5[1]),.doutc(w_n279_5[2]),.din(w_n279_1[1]));
	jspl3 jspl3_w_n279_6(.douta(w_n279_6[0]),.doutb(w_n279_6[1]),.doutc(w_n279_6[2]),.din(w_n279_1[2]));
	jspl jspl_w_n279_7(.douta(w_n279_7[0]),.doutb(w_n279_7[1]),.din(w_n279_2[0]));
	jspl3 jspl3_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.doutc(w_n281_0[2]),.din(n281));
	jspl jspl_w_n281_1(.douta(w_n281_1[0]),.doutb(w_n281_1[1]),.din(w_n281_0[0]));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.doutc(w_n282_0[2]),.din(n282));
	jspl3 jspl3_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.doutc(w_n282_1[2]),.din(w_n282_0[0]));
	jspl3 jspl3_w_n282_2(.douta(w_n282_2[0]),.doutb(w_n282_2[1]),.doutc(w_n282_2[2]),.din(w_n282_0[1]));
	jspl3 jspl3_w_n282_3(.douta(w_n282_3[0]),.doutb(w_n282_3[1]),.doutc(w_n282_3[2]),.din(w_n282_0[2]));
	jspl3 jspl3_w_n282_4(.douta(w_n282_4[0]),.doutb(w_n282_4[1]),.doutc(w_n282_4[2]),.din(w_n282_1[0]));
	jspl3 jspl3_w_n282_5(.douta(w_n282_5[0]),.doutb(w_n282_5[1]),.doutc(w_n282_5[2]),.din(w_n282_1[1]));
	jspl3 jspl3_w_n282_6(.douta(w_n282_6[0]),.doutb(w_n282_6[1]),.doutc(w_n282_6[2]),.din(w_n282_1[2]));
	jspl jspl_w_n282_7(.douta(w_n282_7[0]),.doutb(w_n282_7[1]),.din(w_n282_2[0]));
	jspl3 jspl3_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.doutc(w_n284_0[2]),.din(n284));
	jspl3 jspl3_w_n284_1(.douta(w_n284_1[0]),.doutb(w_n284_1[1]),.doutc(w_n284_1[2]),.din(w_n284_0[0]));
	jspl3 jspl3_w_n284_2(.douta(w_n284_2[0]),.doutb(w_n284_2[1]),.doutc(w_n284_2[2]),.din(w_n284_0[1]));
	jspl3 jspl3_w_n284_3(.douta(w_n284_3[0]),.doutb(w_n284_3[1]),.doutc(w_n284_3[2]),.din(w_n284_0[2]));
	jspl3 jspl3_w_n284_4(.douta(w_n284_4[0]),.doutb(w_n284_4[1]),.doutc(w_n284_4[2]),.din(w_n284_1[0]));
	jspl3 jspl3_w_n284_5(.douta(w_n284_5[0]),.doutb(w_n284_5[1]),.doutc(w_n284_5[2]),.din(w_n284_1[1]));
	jspl3 jspl3_w_n284_6(.douta(w_n284_6[0]),.doutb(w_n284_6[1]),.doutc(w_n284_6[2]),.din(w_n284_1[2]));
	jspl jspl_w_n284_7(.douta(w_n284_7[0]),.doutb(w_n284_7[1]),.din(w_n284_2[0]));
	jspl3 jspl3_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.doutc(w_n286_0[2]),.din(n286));
	jspl jspl_w_n286_1(.douta(w_n286_1[0]),.doutb(w_n286_1[1]),.din(w_n286_0[0]));
	jspl3 jspl3_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.doutc(w_n287_0[2]),.din(n287));
	jspl3 jspl3_w_n287_1(.douta(w_n287_1[0]),.doutb(w_n287_1[1]),.doutc(w_n287_1[2]),.din(w_n287_0[0]));
	jspl3 jspl3_w_n287_2(.douta(w_n287_2[0]),.doutb(w_n287_2[1]),.doutc(w_n287_2[2]),.din(w_n287_0[1]));
	jspl3 jspl3_w_n287_3(.douta(w_n287_3[0]),.doutb(w_n287_3[1]),.doutc(w_n287_3[2]),.din(w_n287_0[2]));
	jspl3 jspl3_w_n287_4(.douta(w_n287_4[0]),.doutb(w_n287_4[1]),.doutc(w_n287_4[2]),.din(w_n287_1[0]));
	jspl3 jspl3_w_n287_5(.douta(w_n287_5[0]),.doutb(w_n287_5[1]),.doutc(w_n287_5[2]),.din(w_n287_1[1]));
	jspl3 jspl3_w_n287_6(.douta(w_n287_6[0]),.doutb(w_n287_6[1]),.doutc(w_n287_6[2]),.din(w_n287_1[2]));
	jspl jspl_w_n287_7(.douta(w_n287_7[0]),.doutb(w_n287_7[1]),.din(w_n287_2[0]));
	jspl3 jspl3_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.doutc(w_n289_0[2]),.din(n289));
	jspl jspl_w_n289_1(.douta(w_n289_1[0]),.doutb(w_n289_1[1]),.din(w_n289_0[0]));
	jspl3 jspl3_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(n290));
	jspl3 jspl3_w_n290_1(.douta(w_n290_1[0]),.doutb(w_n290_1[1]),.doutc(w_n290_1[2]),.din(w_n290_0[0]));
	jspl3 jspl3_w_n290_2(.douta(w_n290_2[0]),.doutb(w_n290_2[1]),.doutc(w_n290_2[2]),.din(w_n290_0[1]));
	jspl3 jspl3_w_n290_3(.douta(w_n290_3[0]),.doutb(w_n290_3[1]),.doutc(w_n290_3[2]),.din(w_n290_0[2]));
	jspl3 jspl3_w_n290_4(.douta(w_n290_4[0]),.doutb(w_n290_4[1]),.doutc(w_n290_4[2]),.din(w_n290_1[0]));
	jspl3 jspl3_w_n290_5(.douta(w_n290_5[0]),.doutb(w_n290_5[1]),.doutc(w_n290_5[2]),.din(w_n290_1[1]));
	jspl3 jspl3_w_n290_6(.douta(w_n290_6[0]),.doutb(w_n290_6[1]),.doutc(w_n290_6[2]),.din(w_n290_1[2]));
	jspl jspl_w_n290_7(.douta(w_n290_7[0]),.doutb(w_n290_7[1]),.din(w_n290_2[0]));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl3 jspl3_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.doutc(w_n292_1[2]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n292_2(.douta(w_n292_2[0]),.doutb(w_n292_2[1]),.doutc(w_n292_2[2]),.din(w_n292_0[1]));
	jspl3 jspl3_w_n292_3(.douta(w_n292_3[0]),.doutb(w_n292_3[1]),.doutc(w_n292_3[2]),.din(w_n292_0[2]));
	jspl3 jspl3_w_n292_4(.douta(w_n292_4[0]),.doutb(w_n292_4[1]),.doutc(w_n292_4[2]),.din(w_n292_1[0]));
	jspl3 jspl3_w_n292_5(.douta(w_n292_5[0]),.doutb(w_n292_5[1]),.doutc(w_n292_5[2]),.din(w_n292_1[1]));
	jspl3 jspl3_w_n292_6(.douta(w_n292_6[0]),.doutb(w_n292_6[1]),.doutc(w_n292_6[2]),.din(w_n292_1[2]));
	jspl jspl_w_n292_7(.douta(w_n292_7[0]),.doutb(w_n292_7[1]),.din(w_n292_2[0]));
	jspl3 jspl3_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.doutc(w_n294_0[2]),.din(n294));
	jspl3 jspl3_w_n294_1(.douta(w_n294_1[0]),.doutb(w_n294_1[1]),.doutc(w_n294_1[2]),.din(w_n294_0[0]));
	jspl3 jspl3_w_n294_2(.douta(w_n294_2[0]),.doutb(w_n294_2[1]),.doutc(w_n294_2[2]),.din(w_n294_0[1]));
	jspl3 jspl3_w_n294_3(.douta(w_n294_3[0]),.doutb(w_n294_3[1]),.doutc(w_n294_3[2]),.din(w_n294_0[2]));
	jspl3 jspl3_w_n294_4(.douta(w_n294_4[0]),.doutb(w_n294_4[1]),.doutc(w_n294_4[2]),.din(w_n294_1[0]));
	jspl3 jspl3_w_n294_5(.douta(w_n294_5[0]),.doutb(w_n294_5[1]),.doutc(w_n294_5[2]),.din(w_n294_1[1]));
	jspl3 jspl3_w_n294_6(.douta(w_n294_6[0]),.doutb(w_n294_6[1]),.doutc(w_n294_6[2]),.din(w_n294_1[2]));
	jspl jspl_w_n294_7(.douta(w_n294_7[0]),.doutb(w_n294_7[1]),.din(w_n294_2[0]));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n296_1(.douta(w_n296_1[0]),.doutb(w_n296_1[1]),.din(w_n296_0[0]));
	jspl3 jspl3_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.doutc(w_n297_0[2]),.din(n297));
	jspl3 jspl3_w_n297_1(.douta(w_n297_1[0]),.doutb(w_n297_1[1]),.doutc(w_n297_1[2]),.din(w_n297_0[0]));
	jspl3 jspl3_w_n297_2(.douta(w_n297_2[0]),.doutb(w_n297_2[1]),.doutc(w_n297_2[2]),.din(w_n297_0[1]));
	jspl3 jspl3_w_n297_3(.douta(w_n297_3[0]),.doutb(w_n297_3[1]),.doutc(w_n297_3[2]),.din(w_n297_0[2]));
	jspl3 jspl3_w_n297_4(.douta(w_n297_4[0]),.doutb(w_n297_4[1]),.doutc(w_n297_4[2]),.din(w_n297_1[0]));
	jspl3 jspl3_w_n297_5(.douta(w_n297_5[0]),.doutb(w_n297_5[1]),.doutc(w_n297_5[2]),.din(w_n297_1[1]));
	jspl3 jspl3_w_n297_6(.douta(w_n297_6[0]),.doutb(w_n297_6[1]),.doutc(w_n297_6[2]),.din(w_n297_1[2]));
	jspl jspl_w_n297_7(.douta(w_n297_7[0]),.doutb(w_n297_7[1]),.din(w_n297_2[0]));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl3 jspl3_w_n299_1(.douta(w_n299_1[0]),.doutb(w_n299_1[1]),.doutc(w_n299_1[2]),.din(w_n299_0[0]));
	jspl3 jspl3_w_n299_2(.douta(w_n299_2[0]),.doutb(w_n299_2[1]),.doutc(w_n299_2[2]),.din(w_n299_0[1]));
	jspl3 jspl3_w_n299_3(.douta(w_n299_3[0]),.doutb(w_n299_3[1]),.doutc(w_n299_3[2]),.din(w_n299_0[2]));
	jspl3 jspl3_w_n299_4(.douta(w_n299_4[0]),.doutb(w_n299_4[1]),.doutc(w_n299_4[2]),.din(w_n299_1[0]));
	jspl3 jspl3_w_n299_5(.douta(w_n299_5[0]),.doutb(w_n299_5[1]),.doutc(w_n299_5[2]),.din(w_n299_1[1]));
	jspl3 jspl3_w_n299_6(.douta(w_n299_6[0]),.doutb(w_n299_6[1]),.doutc(w_n299_6[2]),.din(w_n299_1[2]));
	jspl jspl_w_n299_7(.douta(w_n299_7[0]),.doutb(w_n299_7[1]),.din(w_n299_2[0]));
	jspl3 jspl3_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.doutc(w_n301_0[2]),.din(n301));
	jspl jspl_w_n301_1(.douta(w_n301_1[0]),.doutb(w_n301_1[1]),.din(w_n301_0[0]));
	jspl3 jspl3_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.doutc(w_n302_0[2]),.din(n302));
	jspl3 jspl3_w_n302_1(.douta(w_n302_1[0]),.doutb(w_n302_1[1]),.doutc(w_n302_1[2]),.din(w_n302_0[0]));
	jspl3 jspl3_w_n302_2(.douta(w_n302_2[0]),.doutb(w_n302_2[1]),.doutc(w_n302_2[2]),.din(w_n302_0[1]));
	jspl3 jspl3_w_n302_3(.douta(w_n302_3[0]),.doutb(w_n302_3[1]),.doutc(w_n302_3[2]),.din(w_n302_0[2]));
	jspl3 jspl3_w_n302_4(.douta(w_n302_4[0]),.doutb(w_n302_4[1]),.doutc(w_n302_4[2]),.din(w_n302_1[0]));
	jspl3 jspl3_w_n302_5(.douta(w_n302_5[0]),.doutb(w_n302_5[1]),.doutc(w_n302_5[2]),.din(w_n302_1[1]));
	jspl3 jspl3_w_n302_6(.douta(w_n302_6[0]),.doutb(w_n302_6[1]),.doutc(w_n302_6[2]),.din(w_n302_1[2]));
	jspl jspl_w_n302_7(.douta(w_n302_7[0]),.doutb(w_n302_7[1]),.din(w_n302_2[0]));
	jspl3 jspl3_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.doutc(w_n304_0[2]),.din(n304));
	jspl3 jspl3_w_n304_1(.douta(w_n304_1[0]),.doutb(w_n304_1[1]),.doutc(w_n304_1[2]),.din(w_n304_0[0]));
	jspl3 jspl3_w_n304_2(.douta(w_n304_2[0]),.doutb(w_n304_2[1]),.doutc(w_n304_2[2]),.din(w_n304_0[1]));
	jspl3 jspl3_w_n304_3(.douta(w_n304_3[0]),.doutb(w_n304_3[1]),.doutc(w_n304_3[2]),.din(w_n304_0[2]));
	jspl3 jspl3_w_n304_4(.douta(w_n304_4[0]),.doutb(w_n304_4[1]),.doutc(w_n304_4[2]),.din(w_n304_1[0]));
	jspl3 jspl3_w_n304_5(.douta(w_n304_5[0]),.doutb(w_n304_5[1]),.doutc(w_n304_5[2]),.din(w_n304_1[1]));
	jspl3 jspl3_w_n304_6(.douta(w_n304_6[0]),.doutb(w_n304_6[1]),.doutc(w_n304_6[2]),.din(w_n304_1[2]));
	jspl jspl_w_n304_7(.douta(w_n304_7[0]),.doutb(w_n304_7[1]),.din(w_n304_2[0]));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.doutc(w_n306_0[2]),.din(n306));
	jspl3 jspl3_w_n306_1(.douta(w_n306_1[0]),.doutb(w_n306_1[1]),.doutc(w_n306_1[2]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n306_2(.douta(w_n306_2[0]),.doutb(w_n306_2[1]),.doutc(w_n306_2[2]),.din(w_n306_0[1]));
	jspl3 jspl3_w_n306_3(.douta(w_n306_3[0]),.doutb(w_n306_3[1]),.doutc(w_n306_3[2]),.din(w_n306_0[2]));
	jspl3 jspl3_w_n306_4(.douta(w_n306_4[0]),.doutb(w_n306_4[1]),.doutc(w_n306_4[2]),.din(w_n306_1[0]));
	jspl3 jspl3_w_n306_5(.douta(w_n306_5[0]),.doutb(w_n306_5[1]),.doutc(w_n306_5[2]),.din(w_n306_1[1]));
	jspl3 jspl3_w_n306_6(.douta(w_n306_6[0]),.doutb(w_n306_6[1]),.doutc(w_n306_6[2]),.din(w_n306_1[2]));
	jspl jspl_w_n306_7(.douta(w_n306_7[0]),.doutb(w_n306_7[1]),.din(w_n306_2[0]));
	jspl3 jspl3_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.doutc(w_n308_0[2]),.din(n308));
	jspl3 jspl3_w_n308_1(.douta(w_n308_1[0]),.doutb(w_n308_1[1]),.doutc(w_n308_1[2]),.din(w_n308_0[0]));
	jspl3 jspl3_w_n308_2(.douta(w_n308_2[0]),.doutb(w_n308_2[1]),.doutc(w_n308_2[2]),.din(w_n308_0[1]));
	jspl3 jspl3_w_n308_3(.douta(w_n308_3[0]),.doutb(w_n308_3[1]),.doutc(w_n308_3[2]),.din(w_n308_0[2]));
	jspl3 jspl3_w_n308_4(.douta(w_n308_4[0]),.doutb(w_n308_4[1]),.doutc(w_n308_4[2]),.din(w_n308_1[0]));
	jspl3 jspl3_w_n308_5(.douta(w_n308_5[0]),.doutb(w_n308_5[1]),.doutc(w_n308_5[2]),.din(w_n308_1[1]));
	jspl3 jspl3_w_n308_6(.douta(w_n308_6[0]),.doutb(w_n308_6[1]),.doutc(w_n308_6[2]),.din(w_n308_1[2]));
	jspl jspl_w_n308_7(.douta(w_n308_7[0]),.doutb(w_n308_7[1]),.din(w_n308_2[0]));
	jspl3 jspl3_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.doutc(w_n310_0[2]),.din(n310));
	jspl3 jspl3_w_n310_1(.douta(w_n310_1[0]),.doutb(w_n310_1[1]),.doutc(w_n310_1[2]),.din(w_n310_0[0]));
	jspl3 jspl3_w_n310_2(.douta(w_n310_2[0]),.doutb(w_n310_2[1]),.doutc(w_n310_2[2]),.din(w_n310_0[1]));
	jspl3 jspl3_w_n310_3(.douta(w_n310_3[0]),.doutb(w_n310_3[1]),.doutc(w_n310_3[2]),.din(w_n310_0[2]));
	jspl3 jspl3_w_n310_4(.douta(w_n310_4[0]),.doutb(w_n310_4[1]),.doutc(w_n310_4[2]),.din(w_n310_1[0]));
	jspl3 jspl3_w_n310_5(.douta(w_n310_5[0]),.doutb(w_n310_5[1]),.doutc(w_n310_5[2]),.din(w_n310_1[1]));
	jspl3 jspl3_w_n310_6(.douta(w_n310_6[0]),.doutb(w_n310_6[1]),.doutc(w_n310_6[2]),.din(w_n310_1[2]));
	jspl jspl_w_n310_7(.douta(w_n310_7[0]),.doutb(w_n310_7[1]),.din(w_n310_2[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_dff_A_J4cuJkSl9_1),.doutc(w_dff_A_hkly1Ioj9_2),.din(n312));
	jspl3 jspl3_w_n312_1(.douta(w_dff_A_Ly8npyZr5_0),.doutb(w_n312_1[1]),.doutc(w_dff_A_egJSvUHp6_2),.din(w_n312_0[0]));
	jspl3 jspl3_w_n312_2(.douta(w_n312_2[0]),.doutb(w_n312_2[1]),.doutc(w_n312_2[2]),.din(w_n312_0[1]));
	jspl3 jspl3_w_n312_3(.douta(w_n312_3[0]),.doutb(w_n312_3[1]),.doutc(w_n312_3[2]),.din(w_n312_0[2]));
	jspl3 jspl3_w_n312_4(.douta(w_n312_4[0]),.doutb(w_n312_4[1]),.doutc(w_n312_4[2]),.din(w_n312_1[0]));
	jspl3 jspl3_w_n312_5(.douta(w_n312_5[0]),.doutb(w_dff_A_x9tybVmZ8_1),.doutc(w_dff_A_hXKPEsEE7_2),.din(w_n312_1[1]));
	jspl3 jspl3_w_n312_6(.douta(w_n312_6[0]),.doutb(w_n312_6[1]),.doutc(w_n312_6[2]),.din(w_n312_1[2]));
	jspl jspl_w_n312_7(.douta(w_n312_7[0]),.doutb(w_n312_7[1]),.din(w_n312_2[0]));
	jspl3 jspl3_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n314_1(.douta(w_n314_1[0]),.doutb(w_n314_1[1]),.din(w_n314_0[0]));
	jspl3 jspl3_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.doutc(w_n315_0[2]),.din(n315));
	jspl3 jspl3_w_n315_1(.douta(w_n315_1[0]),.doutb(w_n315_1[1]),.doutc(w_n315_1[2]),.din(w_n315_0[0]));
	jspl3 jspl3_w_n315_2(.douta(w_n315_2[0]),.doutb(w_n315_2[1]),.doutc(w_n315_2[2]),.din(w_n315_0[1]));
	jspl3 jspl3_w_n315_3(.douta(w_n315_3[0]),.doutb(w_n315_3[1]),.doutc(w_n315_3[2]),.din(w_n315_0[2]));
	jspl3 jspl3_w_n315_4(.douta(w_n315_4[0]),.doutb(w_n315_4[1]),.doutc(w_n315_4[2]),.din(w_n315_1[0]));
	jspl3 jspl3_w_n315_5(.douta(w_n315_5[0]),.doutb(w_n315_5[1]),.doutc(w_n315_5[2]),.din(w_n315_1[1]));
	jspl3 jspl3_w_n315_6(.douta(w_n315_6[0]),.doutb(w_n315_6[1]),.doutc(w_n315_6[2]),.din(w_n315_1[2]));
	jspl jspl_w_n315_7(.douta(w_n315_7[0]),.doutb(w_n315_7[1]),.din(w_n315_2[0]));
	jspl3 jspl3_w_n332_0(.douta(w_n332_0[0]),.doutb(w_n332_0[1]),.doutc(w_n332_0[2]),.din(n332));
	jspl jspl_w_n332_1(.douta(w_n332_1[0]),.doutb(w_n332_1[1]),.din(w_n332_0[0]));
	jspl3 jspl3_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.doutc(w_n333_0[2]),.din(n333));
	jspl3 jspl3_w_n333_1(.douta(w_n333_1[0]),.doutb(w_n333_1[1]),.doutc(w_n333_1[2]),.din(w_n333_0[0]));
	jspl3 jspl3_w_n333_2(.douta(w_n333_2[0]),.doutb(w_n333_2[1]),.doutc(w_n333_2[2]),.din(w_n333_0[1]));
	jspl3 jspl3_w_n333_3(.douta(w_n333_3[0]),.doutb(w_n333_3[1]),.doutc(w_n333_3[2]),.din(w_n333_0[2]));
	jspl3 jspl3_w_n333_4(.douta(w_n333_4[0]),.doutb(w_n333_4[1]),.doutc(w_n333_4[2]),.din(w_n333_1[0]));
	jspl3 jspl3_w_n333_5(.douta(w_n333_5[0]),.doutb(w_n333_5[1]),.doutc(w_n333_5[2]),.din(w_n333_1[1]));
	jspl3 jspl3_w_n333_6(.douta(w_n333_6[0]),.doutb(w_n333_6[1]),.doutc(w_n333_6[2]),.din(w_n333_1[2]));
	jspl jspl_w_n333_7(.douta(w_n333_7[0]),.doutb(w_n333_7[1]),.din(w_n333_2[0]));
	jspl3 jspl3_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.doutc(w_n350_0[2]),.din(n350));
	jspl jspl_w_n350_1(.douta(w_n350_1[0]),.doutb(w_n350_1[1]),.din(w_n350_0[0]));
	jspl3 jspl3_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.doutc(w_n351_0[2]),.din(n351));
	jspl3 jspl3_w_n351_1(.douta(w_n351_1[0]),.doutb(w_n351_1[1]),.doutc(w_n351_1[2]),.din(w_n351_0[0]));
	jspl3 jspl3_w_n351_2(.douta(w_n351_2[0]),.doutb(w_n351_2[1]),.doutc(w_n351_2[2]),.din(w_n351_0[1]));
	jspl3 jspl3_w_n351_3(.douta(w_n351_3[0]),.doutb(w_n351_3[1]),.doutc(w_n351_3[2]),.din(w_n351_0[2]));
	jspl3 jspl3_w_n351_4(.douta(w_n351_4[0]),.doutb(w_n351_4[1]),.doutc(w_n351_4[2]),.din(w_n351_1[0]));
	jspl3 jspl3_w_n351_5(.douta(w_n351_5[0]),.doutb(w_n351_5[1]),.doutc(w_n351_5[2]),.din(w_n351_1[1]));
	jspl3 jspl3_w_n351_6(.douta(w_n351_6[0]),.doutb(w_n351_6[1]),.doutc(w_n351_6[2]),.din(w_n351_1[2]));
	jspl jspl_w_n351_7(.douta(w_n351_7[0]),.doutb(w_n351_7[1]),.din(w_n351_2[0]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl jspl_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.doutc(w_n369_0[2]),.din(n369));
	jspl3 jspl3_w_n369_1(.douta(w_n369_1[0]),.doutb(w_n369_1[1]),.doutc(w_n369_1[2]),.din(w_n369_0[0]));
	jspl3 jspl3_w_n369_2(.douta(w_n369_2[0]),.doutb(w_n369_2[1]),.doutc(w_n369_2[2]),.din(w_n369_0[1]));
	jspl3 jspl3_w_n369_3(.douta(w_n369_3[0]),.doutb(w_n369_3[1]),.doutc(w_n369_3[2]),.din(w_n369_0[2]));
	jspl3 jspl3_w_n369_4(.douta(w_n369_4[0]),.doutb(w_n369_4[1]),.doutc(w_n369_4[2]),.din(w_n369_1[0]));
	jspl3 jspl3_w_n369_5(.douta(w_n369_5[0]),.doutb(w_n369_5[1]),.doutc(w_n369_5[2]),.din(w_n369_1[1]));
	jspl3 jspl3_w_n369_6(.douta(w_n369_6[0]),.doutb(w_n369_6[1]),.doutc(w_n369_6[2]),.din(w_n369_1[2]));
	jspl jspl_w_n369_7(.douta(w_n369_7[0]),.doutb(w_n369_7[1]),.din(w_n369_2[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.doutc(w_n386_1[2]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n386_2(.douta(w_n386_2[0]),.doutb(w_n386_2[1]),.doutc(w_n386_2[2]),.din(w_n386_0[1]));
	jspl3 jspl3_w_n386_3(.douta(w_n386_3[0]),.doutb(w_n386_3[1]),.doutc(w_n386_3[2]),.din(w_n386_0[2]));
	jspl3 jspl3_w_n386_4(.douta(w_n386_4[0]),.doutb(w_n386_4[1]),.doutc(w_n386_4[2]),.din(w_n386_1[0]));
	jspl3 jspl3_w_n386_5(.douta(w_n386_5[0]),.doutb(w_n386_5[1]),.doutc(w_n386_5[2]),.din(w_n386_1[1]));
	jspl3 jspl3_w_n386_6(.douta(w_n386_6[0]),.doutb(w_n386_6[1]),.doutc(w_n386_6[2]),.din(w_n386_1[2]));
	jspl jspl_w_n386_7(.douta(w_n386_7[0]),.doutb(w_n386_7[1]),.din(w_n386_2[0]));
	jspl3 jspl3_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.doutc(w_n403_0[2]),.din(n403));
	jspl3 jspl3_w_n403_1(.douta(w_n403_1[0]),.doutb(w_n403_1[1]),.doutc(w_n403_1[2]),.din(w_n403_0[0]));
	jspl3 jspl3_w_n403_2(.douta(w_n403_2[0]),.doutb(w_n403_2[1]),.doutc(w_n403_2[2]),.din(w_n403_0[1]));
	jspl3 jspl3_w_n403_3(.douta(w_n403_3[0]),.doutb(w_n403_3[1]),.doutc(w_n403_3[2]),.din(w_n403_0[2]));
	jspl3 jspl3_w_n403_4(.douta(w_n403_4[0]),.doutb(w_n403_4[1]),.doutc(w_n403_4[2]),.din(w_n403_1[0]));
	jspl3 jspl3_w_n403_5(.douta(w_n403_5[0]),.doutb(w_n403_5[1]),.doutc(w_n403_5[2]),.din(w_n403_1[1]));
	jspl3 jspl3_w_n403_6(.douta(w_n403_6[0]),.doutb(w_n403_6[1]),.doutc(w_n403_6[2]),.din(w_n403_1[2]));
	jspl jspl_w_n403_7(.douta(w_n403_7[0]),.doutb(w_n403_7[1]),.din(w_n403_2[0]));
	jspl3 jspl3_w_n420_0(.douta(w_dff_A_qjAdWqQ03_0),.doutb(w_n420_0[1]),.doutc(w_dff_A_060PweF86_2),.din(n420));
	jspl3 jspl3_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.doutc(w_n420_1[2]),.din(w_n420_0[0]));
	jspl3 jspl3_w_n420_2(.douta(w_dff_A_Gf2kgLWc7_0),.doutb(w_n420_2[1]),.doutc(w_dff_A_6pXnAQTl5_2),.din(w_n420_0[1]));
	jspl3 jspl3_w_n420_3(.douta(w_n420_3[0]),.doutb(w_n420_3[1]),.doutc(w_n420_3[2]),.din(w_n420_0[2]));
	jspl3 jspl3_w_n420_4(.douta(w_n420_4[0]),.doutb(w_n420_4[1]),.doutc(w_n420_4[2]),.din(w_n420_1[0]));
	jspl3 jspl3_w_n420_5(.douta(w_n420_5[0]),.doutb(w_n420_5[1]),.doutc(w_n420_5[2]),.din(w_n420_1[1]));
	jspl3 jspl3_w_n420_6(.douta(w_n420_6[0]),.doutb(w_n420_6[1]),.doutc(w_n420_6[2]),.din(w_n420_1[2]));
	jspl jspl_w_n420_7(.douta(w_n420_7[0]),.doutb(w_n420_7[1]),.din(w_n420_2[0]));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl3 jspl3_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.doutc(w_n438_0[2]),.din(n438));
	jspl jspl_w_n438_1(.douta(w_n438_1[0]),.doutb(w_n438_1[1]),.din(w_n438_0[0]));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl3 jspl3_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.doutc(w_n439_1[2]),.din(w_n439_0[0]));
	jspl3 jspl3_w_n439_2(.douta(w_n439_2[0]),.doutb(w_n439_2[1]),.doutc(w_n439_2[2]),.din(w_n439_0[1]));
	jspl3 jspl3_w_n439_3(.douta(w_n439_3[0]),.doutb(w_n439_3[1]),.doutc(w_n439_3[2]),.din(w_n439_0[2]));
	jspl3 jspl3_w_n439_4(.douta(w_n439_4[0]),.doutb(w_n439_4[1]),.doutc(w_n439_4[2]),.din(w_n439_1[0]));
	jspl3 jspl3_w_n439_5(.douta(w_n439_5[0]),.doutb(w_n439_5[1]),.doutc(w_n439_5[2]),.din(w_n439_1[1]));
	jspl3 jspl3_w_n439_6(.douta(w_n439_6[0]),.doutb(w_n439_6[1]),.doutc(w_n439_6[2]),.din(w_n439_1[2]));
	jspl jspl_w_n439_7(.douta(w_n439_7[0]),.doutb(w_n439_7[1]),.din(w_n439_2[0]));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.doutc(w_n456_0[2]),.din(n456));
	jspl3 jspl3_w_n456_1(.douta(w_n456_1[0]),.doutb(w_n456_1[1]),.doutc(w_n456_1[2]),.din(w_n456_0[0]));
	jspl3 jspl3_w_n456_2(.douta(w_n456_2[0]),.doutb(w_n456_2[1]),.doutc(w_n456_2[2]),.din(w_n456_0[1]));
	jspl3 jspl3_w_n456_3(.douta(w_n456_3[0]),.doutb(w_n456_3[1]),.doutc(w_n456_3[2]),.din(w_n456_0[2]));
	jspl3 jspl3_w_n456_4(.douta(w_n456_4[0]),.doutb(w_n456_4[1]),.doutc(w_n456_4[2]),.din(w_n456_1[0]));
	jspl3 jspl3_w_n456_5(.douta(w_n456_5[0]),.doutb(w_n456_5[1]),.doutc(w_n456_5[2]),.din(w_n456_1[1]));
	jspl3 jspl3_w_n456_6(.douta(w_n456_6[0]),.doutb(w_n456_6[1]),.doutc(w_n456_6[2]),.din(w_n456_1[2]));
	jspl jspl_w_n456_7(.douta(w_n456_7[0]),.doutb(w_n456_7[1]),.din(w_n456_2[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_n473_0[2]),.din(n473));
	jspl3 jspl3_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl3 jspl3_w_n473_2(.douta(w_n473_2[0]),.doutb(w_n473_2[1]),.doutc(w_n473_2[2]),.din(w_n473_0[1]));
	jspl3 jspl3_w_n473_3(.douta(w_n473_3[0]),.doutb(w_n473_3[1]),.doutc(w_n473_3[2]),.din(w_n473_0[2]));
	jspl3 jspl3_w_n473_4(.douta(w_n473_4[0]),.doutb(w_n473_4[1]),.doutc(w_n473_4[2]),.din(w_n473_1[0]));
	jspl3 jspl3_w_n473_5(.douta(w_n473_5[0]),.doutb(w_n473_5[1]),.doutc(w_n473_5[2]),.din(w_n473_1[1]));
	jspl3 jspl3_w_n473_6(.douta(w_n473_6[0]),.doutb(w_n473_6[1]),.doutc(w_n473_6[2]),.din(w_n473_1[2]));
	jspl jspl_w_n473_7(.douta(w_n473_7[0]),.doutb(w_n473_7[1]),.din(w_n473_2[0]));
	jspl3 jspl3_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.doutc(w_n490_0[2]),.din(n490));
	jspl3 jspl3_w_n490_1(.douta(w_n490_1[0]),.doutb(w_n490_1[1]),.doutc(w_n490_1[2]),.din(w_n490_0[0]));
	jspl3 jspl3_w_n490_2(.douta(w_n490_2[0]),.doutb(w_n490_2[1]),.doutc(w_n490_2[2]),.din(w_n490_0[1]));
	jspl3 jspl3_w_n490_3(.douta(w_n490_3[0]),.doutb(w_n490_3[1]),.doutc(w_n490_3[2]),.din(w_n490_0[2]));
	jspl3 jspl3_w_n490_4(.douta(w_n490_4[0]),.doutb(w_n490_4[1]),.doutc(w_n490_4[2]),.din(w_n490_1[0]));
	jspl3 jspl3_w_n490_5(.douta(w_n490_5[0]),.doutb(w_n490_5[1]),.doutc(w_n490_5[2]),.din(w_n490_1[1]));
	jspl3 jspl3_w_n490_6(.douta(w_n490_6[0]),.doutb(w_n490_6[1]),.doutc(w_n490_6[2]),.din(w_n490_1[2]));
	jspl jspl_w_n490_7(.douta(w_n490_7[0]),.doutb(w_n490_7[1]),.din(w_n490_2[0]));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.doutc(w_n508_0[2]),.din(n508));
	jspl3 jspl3_w_n508_1(.douta(w_n508_1[0]),.doutb(w_n508_1[1]),.doutc(w_n508_1[2]),.din(w_n508_0[0]));
	jspl3 jspl3_w_n508_2(.douta(w_n508_2[0]),.doutb(w_n508_2[1]),.doutc(w_n508_2[2]),.din(w_n508_0[1]));
	jspl3 jspl3_w_n508_3(.douta(w_n508_3[0]),.doutb(w_n508_3[1]),.doutc(w_n508_3[2]),.din(w_n508_0[2]));
	jspl3 jspl3_w_n508_4(.douta(w_n508_4[0]),.doutb(w_n508_4[1]),.doutc(w_n508_4[2]),.din(w_n508_1[0]));
	jspl3 jspl3_w_n508_5(.douta(w_n508_5[0]),.doutb(w_n508_5[1]),.doutc(w_n508_5[2]),.din(w_n508_1[1]));
	jspl3 jspl3_w_n508_6(.douta(w_n508_6[0]),.doutb(w_n508_6[1]),.doutc(w_n508_6[2]),.din(w_n508_1[2]));
	jspl jspl_w_n508_7(.douta(w_n508_7[0]),.doutb(w_n508_7[1]),.din(w_n508_2[0]));
	jspl3 jspl3_w_n525_0(.douta(w_n525_0[0]),.doutb(w_n525_0[1]),.doutc(w_n525_0[2]),.din(n525));
	jspl3 jspl3_w_n525_1(.douta(w_n525_1[0]),.doutb(w_n525_1[1]),.doutc(w_n525_1[2]),.din(w_n525_0[0]));
	jspl3 jspl3_w_n525_2(.douta(w_n525_2[0]),.doutb(w_n525_2[1]),.doutc(w_n525_2[2]),.din(w_n525_0[1]));
	jspl3 jspl3_w_n525_3(.douta(w_n525_3[0]),.doutb(w_n525_3[1]),.doutc(w_n525_3[2]),.din(w_n525_0[2]));
	jspl3 jspl3_w_n525_4(.douta(w_n525_4[0]),.doutb(w_n525_4[1]),.doutc(w_n525_4[2]),.din(w_n525_1[0]));
	jspl3 jspl3_w_n525_5(.douta(w_n525_5[0]),.doutb(w_n525_5[1]),.doutc(w_n525_5[2]),.din(w_n525_1[1]));
	jspl3 jspl3_w_n525_6(.douta(w_n525_6[0]),.doutb(w_n525_6[1]),.doutc(w_n525_6[2]),.din(w_n525_1[2]));
	jspl jspl_w_n525_7(.douta(w_n525_7[0]),.doutb(w_n525_7[1]),.din(w_n525_2[0]));
	jspl3 jspl3_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.doutc(w_n542_0[2]),.din(n542));
	jspl3 jspl3_w_n542_1(.douta(w_n542_1[0]),.doutb(w_n542_1[1]),.doutc(w_n542_1[2]),.din(w_n542_0[0]));
	jspl3 jspl3_w_n542_2(.douta(w_n542_2[0]),.doutb(w_n542_2[1]),.doutc(w_n542_2[2]),.din(w_n542_0[1]));
	jspl3 jspl3_w_n542_3(.douta(w_n542_3[0]),.doutb(w_n542_3[1]),.doutc(w_n542_3[2]),.din(w_n542_0[2]));
	jspl3 jspl3_w_n542_4(.douta(w_n542_4[0]),.doutb(w_n542_4[1]),.doutc(w_n542_4[2]),.din(w_n542_1[0]));
	jspl3 jspl3_w_n542_5(.douta(w_n542_5[0]),.doutb(w_n542_5[1]),.doutc(w_n542_5[2]),.din(w_n542_1[1]));
	jspl3 jspl3_w_n542_6(.douta(w_n542_6[0]),.doutb(w_n542_6[1]),.doutc(w_n542_6[2]),.din(w_n542_1[2]));
	jspl jspl_w_n542_7(.douta(w_n542_7[0]),.doutb(w_n542_7[1]),.din(w_n542_2[0]));
	jspl3 jspl3_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.doutc(w_n559_0[2]),.din(n559));
	jspl3 jspl3_w_n559_1(.douta(w_n559_1[0]),.doutb(w_n559_1[1]),.doutc(w_n559_1[2]),.din(w_n559_0[0]));
	jspl3 jspl3_w_n559_2(.douta(w_n559_2[0]),.doutb(w_n559_2[1]),.doutc(w_n559_2[2]),.din(w_n559_0[1]));
	jspl3 jspl3_w_n559_3(.douta(w_n559_3[0]),.doutb(w_n559_3[1]),.doutc(w_n559_3[2]),.din(w_n559_0[2]));
	jspl3 jspl3_w_n559_4(.douta(w_n559_4[0]),.doutb(w_n559_4[1]),.doutc(w_n559_4[2]),.din(w_n559_1[0]));
	jspl3 jspl3_w_n559_5(.douta(w_n559_5[0]),.doutb(w_n559_5[1]),.doutc(w_n559_5[2]),.din(w_n559_1[1]));
	jspl3 jspl3_w_n559_6(.douta(w_n559_6[0]),.doutb(w_n559_6[1]),.doutc(w_n559_6[2]),.din(w_n559_1[2]));
	jspl jspl_w_n559_7(.douta(w_n559_7[0]),.doutb(w_n559_7[1]),.din(w_n559_2[0]));
	jdff dff_A_Gf2kgLWc7_0(.dout(w_n420_2[0]),.din(w_dff_A_Gf2kgLWc7_0),.clk(gclk));
	jdff dff_A_6pXnAQTl5_2(.dout(w_n420_2[2]),.din(w_dff_A_6pXnAQTl5_2),.clk(gclk));
	jdff dff_A_qjAdWqQ03_0(.dout(w_n420_0[0]),.din(w_dff_A_qjAdWqQ03_0),.clk(gclk));
	jdff dff_A_060PweF86_2(.dout(w_n420_0[2]),.din(w_dff_A_060PweF86_2),.clk(gclk));
	jdff dff_A_x9tybVmZ8_1(.dout(w_n312_5[1]),.din(w_dff_A_x9tybVmZ8_1),.clk(gclk));
	jdff dff_A_hXKPEsEE7_2(.dout(w_n312_5[2]),.din(w_dff_A_hXKPEsEE7_2),.clk(gclk));
	jdff dff_A_Ly8npyZr5_0(.dout(w_n312_1[0]),.din(w_dff_A_Ly8npyZr5_0),.clk(gclk));
	jdff dff_A_egJSvUHp6_2(.dout(w_n312_1[2]),.din(w_dff_A_egJSvUHp6_2),.clk(gclk));
	jdff dff_A_J4cuJkSl9_1(.dout(w_n312_0[1]),.din(w_dff_A_J4cuJkSl9_1),.clk(gclk));
	jdff dff_A_hkly1Ioj9_2(.dout(w_n312_0[2]),.din(w_dff_A_hkly1Ioj9_2),.clk(gclk));
	jdff dff_A_oBp7Jqop7_2(.dout(selectp1127),.din(w_dff_A_oBp7Jqop7_2),.clk(gclk));
endmodule

