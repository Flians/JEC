/*

c3540:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 276
	jand: 535
	jor: 374

Summary:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jdff: 276
	jand: 535
	jor: 374

The maximum logic level gap of any gate:
	c3540: 26
*/

module rf_c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[2:0] w_G1_2;
	wire[1:0] w_G1_3;
	wire[2:0] w_G13_0;
	wire[1:0] w_G13_1;
	wire[2:0] w_G20_0;
	wire[2:0] w_G20_1;
	wire[2:0] w_G20_2;
	wire[2:0] w_G20_3;
	wire[2:0] w_G20_4;
	wire[2:0] w_G20_5;
	wire[2:0] w_G20_6;
	wire[1:0] w_G20_7;
	wire[2:0] w_G33_0;
	wire[2:0] w_G33_1;
	wire[2:0] w_G33_2;
	wire[2:0] w_G33_3;
	wire[2:0] w_G33_4;
	wire[2:0] w_G33_5;
	wire[2:0] w_G33_6;
	wire[2:0] w_G33_7;
	wire[2:0] w_G33_8;
	wire[2:0] w_G33_9;
	wire[2:0] w_G33_10;
	wire[2:0] w_G33_11;
	wire[2:0] w_G41_0;
	wire[1:0] w_G41_1;
	wire[2:0] w_G45_0;
	wire[2:0] w_G45_1;
	wire[2:0] w_G50_0;
	wire[2:0] w_G50_1;
	wire[2:0] w_G50_2;
	wire[2:0] w_G50_3;
	wire[2:0] w_G50_4;
	wire[2:0] w_G50_5;
	wire[2:0] w_G58_0;
	wire[2:0] w_G58_1;
	wire[2:0] w_G58_2;
	wire[2:0] w_G58_3;
	wire[2:0] w_G58_4;
	wire[1:0] w_G58_5;
	wire[2:0] w_G68_0;
	wire[2:0] w_G68_1;
	wire[2:0] w_G68_2;
	wire[2:0] w_G68_3;
	wire[2:0] w_G68_4;
	wire[1:0] w_G68_5;
	wire[2:0] w_G77_0;
	wire[2:0] w_G77_1;
	wire[2:0] w_G77_2;
	wire[2:0] w_G77_3;
	wire[2:0] w_G77_4;
	wire[1:0] w_G77_5;
	wire[2:0] w_G87_0;
	wire[2:0] w_G87_1;
	wire[2:0] w_G87_2;
	wire[2:0] w_G87_3;
	wire[2:0] w_G97_0;
	wire[2:0] w_G97_1;
	wire[2:0] w_G97_2;
	wire[2:0] w_G97_3;
	wire[2:0] w_G97_4;
	wire[1:0] w_G97_5;
	wire[2:0] w_G107_0;
	wire[2:0] w_G107_1;
	wire[2:0] w_G107_2;
	wire[2:0] w_G107_3;
	wire[2:0] w_G107_4;
	wire[1:0] w_G107_5;
	wire[2:0] w_G116_0;
	wire[2:0] w_G116_1;
	wire[2:0] w_G116_2;
	wire[2:0] w_G116_3;
	wire[2:0] w_G116_4;
	wire[1:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[2:0] w_G132_0;
	wire[1:0] w_G132_1;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G143_0;
	wire[2:0] w_G143_1;
	wire[1:0] w_G143_2;
	wire[2:0] w_G150_0;
	wire[2:0] w_G150_1;
	wire[2:0] w_G150_2;
	wire[1:0] w_G150_3;
	wire[2:0] w_G159_0;
	wire[2:0] w_G159_1;
	wire[2:0] w_G159_2;
	wire[2:0] w_G159_3;
	wire[2:0] w_G169_0;
	wire[1:0] w_G169_1;
	wire[2:0] w_G179_0;
	wire[2:0] w_G179_1;
	wire[2:0] w_G179_2;
	wire[2:0] w_G190_0;
	wire[2:0] w_G190_1;
	wire[2:0] w_G190_2;
	wire[2:0] w_G190_3;
	wire[1:0] w_G190_4;
	wire[2:0] w_G200_0;
	wire[2:0] w_G200_1;
	wire[2:0] w_G200_2;
	wire[2:0] w_G200_3;
	wire[2:0] w_G200_4;
	wire[2:0] w_G213_0;
	wire[1:0] w_G223_0;
	wire[2:0] w_G226_0;
	wire[1:0] w_G226_1;
	wire[2:0] w_G232_0;
	wire[2:0] w_G232_1;
	wire[2:0] w_G238_0;
	wire[2:0] w_G238_1;
	wire[2:0] w_G244_0;
	wire[2:0] w_G244_1;
	wire[2:0] w_G250_0;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[2:0] w_G264_0;
	wire[1:0] w_G264_1;
	wire[2:0] w_G270_0;
	wire[2:0] w_G274_0;
	wire[2:0] w_G283_0;
	wire[2:0] w_G283_1;
	wire[2:0] w_G283_2;
	wire[2:0] w_G283_3;
	wire[2:0] w_G294_0;
	wire[2:0] w_G294_1;
	wire[2:0] w_G294_2;
	wire[1:0] w_G294_3;
	wire[2:0] w_G303_0;
	wire[2:0] w_G303_1;
	wire[2:0] w_G303_2;
	wire[2:0] w_G311_0;
	wire[2:0] w_G311_1;
	wire[2:0] w_G317_0;
	wire[1:0] w_G317_1;
	wire[2:0] w_G322_0;
	wire[1:0] w_G326_0;
	wire[1:0] w_G330_0;
	wire[1:0] w_G343_0;
	wire[2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire[1:0] w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire[1:0] w_G387_0;
	wire G387_fa_;
	wire[2:0] w_n72_0;
	wire[1:0] w_n72_1;
	wire[2:0] w_n73_0;
	wire[2:0] w_n73_1;
	wire[2:0] w_n73_2;
	wire[2:0] w_n74_0;
	wire[1:0] w_n74_1;
	wire[2:0] w_n75_0;
	wire[1:0] w_n75_1;
	wire[1:0] w_n76_0;
	wire[1:0] w_n77_0;
	wire[2:0] w_n79_0;
	wire[2:0] w_n80_0;
	wire[1:0] w_n80_1;
	wire[2:0] w_n81_0;
	wire[2:0] w_n85_0;
	wire[1:0] w_n86_0;
	wire[2:0] w_n88_0;
	wire[1:0] w_n88_1;
	wire[2:0] w_n91_0;
	wire[2:0] w_n91_1;
	wire[1:0] w_n93_0;
	wire[2:0] w_n97_0;
	wire[2:0] w_n97_1;
	wire[1:0] w_n97_2;
	wire[2:0] w_n98_0;
	wire[2:0] w_n98_1;
	wire[1:0] w_n98_2;
	wire[2:0] w_n103_0;
	wire[2:0] w_n105_0;
	wire[2:0] w_n105_1;
	wire[1:0] w_n105_2;
	wire[1:0] w_n106_0;
	wire[2:0] w_n112_0;
	wire[2:0] w_n112_1;
	wire[2:0] w_n112_2;
	wire[2:0] w_n112_3;
	wire[2:0] w_n112_4;
	wire[2:0] w_n112_5;
	wire[2:0] w_n113_0;
	wire[2:0] w_n113_1;
	wire[2:0] w_n113_2;
	wire[1:0] w_n113_3;
	wire[2:0] w_n114_0;
	wire[2:0] w_n114_1;
	wire[2:0] w_n115_0;
	wire[1:0] w_n115_1;
	wire[1:0] w_n116_0;
	wire[2:0] w_n118_0;
	wire[2:0] w_n121_0;
	wire[2:0] w_n122_0;
	wire[1:0] w_n122_1;
	wire[2:0] w_n123_0;
	wire[2:0] w_n123_1;
	wire[1:0] w_n131_0;
	wire[1:0] w_n135_0;
	wire[2:0] w_n137_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n144_0;
	wire[2:0] w_n146_0;
	wire[2:0] w_n146_1;
	wire[2:0] w_n146_2;
	wire[2:0] w_n146_3;
	wire[2:0] w_n147_0;
	wire[2:0] w_n148_0;
	wire[2:0] w_n148_1;
	wire[2:0] w_n148_2;
	wire[2:0] w_n148_3;
	wire[2:0] w_n148_4;
	wire[2:0] w_n148_5;
	wire[2:0] w_n148_6;
	wire[2:0] w_n148_7;
	wire[2:0] w_n148_8;
	wire[2:0] w_n148_9;
	wire[2:0] w_n149_0;
	wire[2:0] w_n149_1;
	wire[1:0] w_n149_2;
	wire[2:0] w_n151_0;
	wire[2:0] w_n151_1;
	wire[2:0] w_n151_2;
	wire[2:0] w_n151_3;
	wire[2:0] w_n151_4;
	wire[2:0] w_n152_0;
	wire[2:0] w_n152_1;
	wire[2:0] w_n152_2;
	wire[1:0] w_n152_3;
	wire[1:0] w_n154_0;
	wire[2:0] w_n155_0;
	wire[2:0] w_n155_1;
	wire[2:0] w_n155_2;
	wire[1:0] w_n155_3;
	wire[2:0] w_n157_0;
	wire[2:0] w_n161_0;
	wire[1:0] w_n161_1;
	wire[2:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[2:0] w_n166_0;
	wire[2:0] w_n166_1;
	wire[2:0] w_n166_2;
	wire[1:0] w_n166_3;
	wire[2:0] w_n170_0;
	wire[1:0] w_n172_0;
	wire[2:0] w_n179_0;
	wire[2:0] w_n179_1;
	wire[1:0] w_n180_0;
	wire[2:0] w_n185_0;
	wire[2:0] w_n185_1;
	wire[2:0] w_n185_2;
	wire[2:0] w_n185_3;
	wire[2:0] w_n189_0;
	wire[2:0] w_n189_1;
	wire[1:0] w_n189_2;
	wire[2:0] w_n190_0;
	wire[2:0] w_n190_1;
	wire[2:0] w_n191_0;
	wire[1:0] w_n195_0;
	wire[2:0] w_n196_0;
	wire[2:0] w_n196_1;
	wire[2:0] w_n196_2;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[2:0] w_n199_0;
	wire[1:0] w_n199_1;
	wire[1:0] w_n201_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n206_0;
	wire[2:0] w_n210_0;
	wire[1:0] w_n213_0;
	wire[1:0] w_n214_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n219_0;
	wire[2:0] w_n221_0;
	wire[1:0] w_n228_0;
	wire[2:0] w_n229_0;
	wire[1:0] w_n230_0;
	wire[2:0] w_n231_0;
	wire[2:0] w_n234_0;
	wire[1:0] w_n241_0;
	wire[2:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[2:0] w_n246_0;
	wire[1:0] w_n246_1;
	wire[1:0] w_n249_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n257_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n262_0;
	wire[2:0] w_n269_0;
	wire[2:0] w_n269_1;
	wire[1:0] w_n270_0;
	wire[2:0] w_n271_0;
	wire[2:0] w_n271_1;
	wire[2:0] w_n274_0;
	wire[1:0] w_n278_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n281_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n288_1;
	wire[1:0] w_n296_0;
	wire[1:0] w_n298_0;
	wire[1:0] w_n300_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n312_0;
	wire[1:0] w_n312_1;
	wire[1:0] w_n315_0;
	wire[1:0] w_n320_0;
	wire[1:0] w_n324_0;
	wire[1:0] w_n328_0;
	wire[1:0] w_n334_0;
	wire[1:0] w_n339_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n346_1;
	wire[2:0] w_n355_0;
	wire[1:0] w_n355_1;
	wire[1:0] w_n362_0;
	wire[2:0] w_n367_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n374_0;
	wire[1:0] w_n381_0;
	wire[2:0] w_n382_0;
	wire[1:0] w_n382_1;
	wire[2:0] w_n385_0;
	wire[1:0] w_n385_1;
	wire[2:0] w_n387_0;
	wire[1:0] w_n387_1;
	wire[1:0] w_n390_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n404_0;
	wire[1:0] w_n405_0;
	wire[2:0] w_n407_0;
	wire[2:0] w_n407_1;
	wire[1:0] w_n407_2;
	wire[1:0] w_n412_0;
	wire[2:0] w_n420_0;
	wire[1:0] w_n420_1;
	wire[2:0] w_n425_0;
	wire[2:0] w_n425_1;
	wire[1:0] w_n426_0;
	wire[1:0] w_n430_0;
	wire[2:0] w_n436_0;
	wire[2:0] w_n439_0;
	wire[1:0] w_n439_1;
	wire[1:0] w_n445_0;
	wire[1:0] w_n446_0;
	wire[2:0] w_n455_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n474_0;
	wire[1:0] w_n475_0;
	wire[1:0] w_n478_0;
	wire[1:0] w_n479_0;
	wire[1:0] w_n483_0;
	wire[1:0] w_n484_0;
	wire[2:0] w_n492_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n508_0;
	wire[1:0] w_n511_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n516_0;
	wire[1:0] w_n517_0;
	wire[2:0] w_n519_0;
	wire[2:0] w_n519_1;
	wire[1:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n528_0;
	wire[1:0] w_n532_0;
	wire[1:0] w_n534_0;
	wire[2:0] w_n536_0;
	wire[1:0] w_n539_0;
	wire[1:0] w_n541_0;
	wire[2:0] w_n542_0;
	wire[1:0] w_n543_0;
	wire[2:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[2:0] w_n552_0;
	wire[1:0] w_n552_1;
	wire[2:0] w_n553_0;
	wire[2:0] w_n553_1;
	wire[2:0] w_n553_2;
	wire[2:0] w_n554_0;
	wire[2:0] w_n554_1;
	wire[2:0] w_n554_2;
	wire[2:0] w_n554_3;
	wire[1:0] w_n556_0;
	wire[1:0] w_n557_0;
	wire[2:0] w_n561_0;
	wire[2:0] w_n563_0;
	wire[1:0] w_n564_0;
	wire[1:0] w_n565_0;
	wire[1:0] w_n567_0;
	wire[2:0] w_n571_0;
	wire[2:0] w_n572_0;
	wire[2:0] w_n573_0;
	wire[2:0] w_n576_0;
	wire[1:0] w_n576_1;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[2:0] w_n589_0;
	wire[2:0] w_n589_1;
	wire[2:0] w_n591_0;
	wire[1:0] w_n591_1;
	wire[2:0] w_n592_0;
	wire[2:0] w_n592_1;
	wire[1:0] w_n592_2;
	wire[2:0] w_n593_0;
	wire[1:0] w_n602_0;
	wire[2:0] w_n603_0;
	wire[2:0] w_n603_1;
	wire[1:0] w_n603_2;
	wire[2:0] w_n604_0;
	wire[2:0] w_n604_1;
	wire[1:0] w_n604_2;
	wire[2:0] w_n605_0;
	wire[2:0] w_n605_1;
	wire[2:0] w_n608_0;
	wire[2:0] w_n608_1;
	wire[2:0] w_n612_0;
	wire[2:0] w_n612_1;
	wire[2:0] w_n612_2;
	wire[2:0] w_n612_3;
	wire[1:0] w_n612_4;
	wire[2:0] w_n613_0;
	wire[1:0] w_n613_1;
	wire[1:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[2:0] w_n617_0;
	wire[2:0] w_n617_1;
	wire[2:0] w_n617_2;
	wire[2:0] w_n617_3;
	wire[2:0] w_n617_4;
	wire[2:0] w_n617_5;
	wire[1:0] w_n617_6;
	wire[1:0] w_n619_0;
	wire[1:0] w_n622_0;
	wire[2:0] w_n623_0;
	wire[2:0] w_n623_1;
	wire[2:0] w_n623_2;
	wire[2:0] w_n623_3;
	wire[2:0] w_n623_4;
	wire[1:0] w_n623_5;
	wire[1:0] w_n626_0;
	wire[2:0] w_n627_0;
	wire[2:0] w_n627_1;
	wire[2:0] w_n627_2;
	wire[2:0] w_n627_3;
	wire[2:0] w_n627_4;
	wire[2:0] w_n627_5;
	wire[2:0] w_n627_6;
	wire[1:0] w_n627_7;
	wire[2:0] w_n631_0;
	wire[2:0] w_n631_1;
	wire[2:0] w_n631_2;
	wire[2:0] w_n631_3;
	wire[2:0] w_n631_4;
	wire[2:0] w_n631_5;
	wire[2:0] w_n631_6;
	wire[1:0] w_n631_7;
	wire[2:0] w_n634_0;
	wire[2:0] w_n634_1;
	wire[2:0] w_n634_2;
	wire[2:0] w_n634_3;
	wire[1:0] w_n634_4;
	wire[2:0] w_n636_0;
	wire[2:0] w_n636_1;
	wire[2:0] w_n636_2;
	wire[2:0] w_n636_3;
	wire[2:0] w_n636_4;
	wire[2:0] w_n636_5;
	wire[2:0] w_n636_6;
	wire[1:0] w_n636_7;
	wire[1:0] w_n639_0;
	wire[2:0] w_n640_0;
	wire[2:0] w_n640_1;
	wire[2:0] w_n640_2;
	wire[2:0] w_n640_3;
	wire[2:0] w_n640_4;
	wire[2:0] w_n640_5;
	wire[2:0] w_n640_6;
	wire[1:0] w_n640_7;
	wire[2:0] w_n642_0;
	wire[2:0] w_n642_1;
	wire[2:0] w_n642_2;
	wire[2:0] w_n642_3;
	wire[2:0] w_n642_4;
	wire[2:0] w_n642_5;
	wire[2:0] w_n642_6;
	wire[1:0] w_n642_7;
	wire[1:0] w_n654_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n661_0;
	wire[2:0] w_n672_0;
	wire[1:0] w_n672_1;
	wire[2:0] w_n675_0;
	wire[1:0] w_n676_0;
	wire[1:0] w_n680_0;
	wire[1:0] w_n692_0;
	wire[2:0] w_n696_0;
	wire[2:0] w_n696_1;
	wire[1:0] w_n717_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n743_0;
	wire[1:0] w_n743_1;
	wire[1:0] w_n750_0;
	wire[1:0] w_n754_0;
	wire[2:0] w_n758_0;
	wire[1:0] w_n758_1;
	wire[1:0] w_n759_0;
	wire[1:0] w_n760_0;
	wire[2:0] w_n764_0;
	wire[2:0] w_n764_1;
	wire[1:0] w_n769_0;
	wire[2:0] w_n771_0;
	wire[1:0] w_n779_0;
	wire[1:0] w_n797_0;
	wire[1:0] w_n801_0;
	wire[1:0] w_n816_0;
	wire[1:0] w_n823_0;
	wire[1:0] w_n825_0;
	wire[2:0] w_n853_0;
	wire[2:0] w_n855_0;
	wire[2:0] w_n861_0;
	wire[1:0] w_n861_1;
	wire[1:0] w_n863_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n899_0;
	wire[1:0] w_n909_0;
	wire[2:0] w_n937_0;
	wire[1:0] w_n940_0;
	wire[1:0] w_n962_0;
	wire[2:0] w_n988_0;
	wire[1:0] w_n990_0;
	wire[2:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[2:0] w_n994_0;
	wire[2:0] w_n996_0;
	wire[1:0] w_n999_0;
	wire[2:0] w_n1001_0;
	wire[2:0] w_n1002_0;
	wire[1:0] w_n1003_0;
	wire[2:0] w_n1049_0;
	wire[1:0] w_n1052_0;
	wire[1:0] w_n1057_0;
	wire[1:0] w_n1059_0;
	wire[1:0] w_n1088_0;
	wire[2:0] w_n1114_0;
	wire[2:0] w_n1162_0;
	wire[1:0] w_n1164_0;
	wire[1:0] w_n1172_0;
	wire[1:0] w_n1175_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1184_0;
	wire[1:0] w_n1187_0;
	wire w_dff_B_M2bk8CTR9_1;
	wire w_dff_B_L5K1pX3c9_1;
	wire w_dff_B_tdIYQyy51_0;
	wire w_dff_B_hLperUKE3_0;
	wire w_dff_B_eTKitgFn8_0;
	wire w_dff_B_YXcrKEAJ2_0;
	wire w_dff_B_39kMmzie6_0;
	wire w_dff_B_cbUMfDkb0_0;
	wire w_dff_B_dFj2zYCq7_0;
	wire w_dff_B_lVRXuHPs2_0;
	wire w_dff_B_BEtrxYBi6_0;
	wire w_dff_B_emsRcblk9_0;
	wire w_dff_B_MbNWeus15_0;
	wire w_dff_B_RM9HVZop1_0;
	wire w_dff_B_4chH4i9T0_0;
	wire w_dff_B_9PPINYUl7_0;
	wire w_dff_B_J5SzWb9M1_0;
	wire w_dff_B_A9nccNNq1_0;
	wire w_dff_B_8MfOWSig9_0;
	wire w_dff_B_A4TviHsX6_0;
	wire w_dff_B_YMeEVwok3_0;
	wire w_dff_B_MCk3Ssc73_0;
	wire w_dff_B_QiudUgjP3_0;
	wire w_dff_B_KYiqwOBi3_0;
	wire w_dff_B_Irm9ncJQ4_0;
	wire w_dff_B_JQkHdphv9_0;
	wire w_dff_B_bDJtiRpV7_0;
	wire w_dff_B_qZMCsC4o3_0;
	wire w_dff_B_gaRAddgQ5_0;
	wire w_dff_A_JD9tOuMB5_0;
	wire w_dff_B_DTvBXyOK4_1;
	wire w_dff_B_eHuJ3Zsg4_1;
	wire w_dff_A_RftdTNmm0_1;
	wire w_dff_B_5PKNBKz49_1;
	wire w_dff_B_iCS2njBI1_1;
	wire w_dff_B_Xbn8CJNi1_1;
	wire w_dff_B_NFbYal1R0_1;
	wire w_dff_B_kzVggnsM9_1;
	wire w_dff_A_EeJc0YC55_0;
	wire w_dff_A_ZQmF1xtq7_0;
	wire w_dff_A_qaUH8K5X8_1;
	wire w_dff_A_4C8JbJYO9_0;
	wire w_dff_A_VmTMOllq2_0;
	wire w_dff_A_ZMqnxzvf1_0;
	wire w_dff_B_B8lF4AdG4_0;
	wire w_dff_B_K7Mb3bCB7_0;
	wire w_dff_B_jdHu0q5J0_0;
	wire w_dff_B_Q5u8Ir0H9_0;
	wire w_dff_B_9CjI7fM78_1;
	wire w_dff_B_Y0HyG9oT8_1;
	wire w_dff_A_Y8dPIE7f0_1;
	wire w_dff_A_HGPx0bsZ1_0;
	wire w_dff_A_mWJJ95QE5_0;
	wire w_dff_A_eHaXs8ak3_2;
	wire w_dff_A_BDdeUnCZ1_0;
	wire w_dff_A_OWxnm4cp3_0;
	wire w_dff_A_RNsFj8bQ7_0;
	wire w_dff_A_ET1kx94Z1_0;
	wire w_dff_A_BBwZ4xyJ9_0;
	wire w_dff_A_RX6J1BbH9_0;
	wire w_dff_A_pMt8nEKh0_0;
	wire w_dff_A_ycarUudx2_0;
	wire w_dff_A_kL1Ia3kA9_0;
	wire w_dff_A_wAuMb2Va8_0;
	wire w_dff_A_MQ1551cG6_0;
	wire w_dff_A_v8W7uE694_0;
	wire w_dff_A_9seO9t8D3_0;
	wire w_dff_A_TUygGutm7_0;
	wire w_dff_A_p43BVdkF8_0;
	wire w_dff_A_i0lg6pko8_0;
	wire w_dff_A_AwYQKIbY0_0;
	wire w_dff_A_z00g9Up74_0;
	wire w_dff_A_rTC27Ujv9_0;
	wire w_dff_A_ZuYHJo5F0_0;
	wire w_dff_A_XRgZIweo0_0;
	wire w_dff_A_4iFfzkXn1_0;
	wire w_dff_A_8v7uQRFZ6_0;
	wire w_dff_A_PVrdWs1m7_0;
	wire w_dff_A_cyNhmvic6_1;
	wire w_dff_A_ya2Aiw553_0;
	wire w_dff_A_6Z7j5pSM8_0;
	wire w_dff_A_DKHdOct33_0;
	wire w_dff_A_iFlNSgwe4_0;
	wire w_dff_A_5vnT0x4x4_0;
	wire w_dff_A_Fwm8XYaE1_0;
	wire w_dff_A_rKoB023L2_0;
	wire w_dff_A_MDXAVeua5_0;
	wire w_dff_A_DBa16L9l0_0;
	wire w_dff_A_0fwKqOTm2_0;
	wire w_dff_A_w45RH9sP7_0;
	wire w_dff_A_T55bB0ag8_0;
	wire w_dff_A_Gn435XAr0_0;
	wire w_dff_A_y1rFtMDE7_0;
	wire w_dff_A_sQMFf0Uv6_0;
	wire w_dff_A_y1V3Up6c1_0;
	wire w_dff_A_gx07RHvg3_0;
	wire w_dff_A_lDM1FK4F9_0;
	wire w_dff_A_buWJidtA9_0;
	wire w_dff_A_xSd0AmbU7_0;
	wire w_dff_A_Ua7qVgcQ1_0;
	wire w_dff_A_UDg6dnwl5_0;
	wire w_dff_A_MaMy1aGw3_0;
	wire w_dff_A_6n9RzDAU9_2;
	wire w_dff_A_iNSP9uw25_0;
	wire w_dff_A_CBPNOo2U9_0;
	wire w_dff_A_JvvWstK53_0;
	wire w_dff_A_nzgTBldx3_0;
	wire w_dff_A_T9L7FZvb1_0;
	wire w_dff_A_xYQy2Xfl7_0;
	wire w_dff_A_RFKNx8NZ0_0;
	wire w_dff_A_f9us52zi7_0;
	wire w_dff_A_T9oJ1gxD2_0;
	wire w_dff_A_dBa4KbTK0_0;
	wire w_dff_A_MfeAzOyP9_0;
	wire w_dff_A_vkpN7A7S9_0;
	wire w_dff_A_9FzQSQQg7_0;
	wire w_dff_A_vDuzeeR05_0;
	wire w_dff_A_PZ8IaZCk7_0;
	wire w_dff_A_eCwCsQfR5_0;
	wire w_dff_A_SoS4AyFT1_0;
	wire w_dff_A_mtE2qBZj4_0;
	wire w_dff_A_L3dAmn8P4_0;
	wire w_dff_A_NF138Mhz6_0;
	wire w_dff_A_x8w3OkNr6_2;
	wire w_dff_A_t3WM7HnJ4_0;
	wire w_dff_A_fmUKup6j7_0;
	wire w_dff_A_Iib65AKQ2_0;
	wire w_dff_A_PH8Lw6Nm5_0;
	wire w_dff_A_nQlaNGRY6_0;
	wire w_dff_A_tBFinChI6_0;
	wire w_dff_A_SnGa4QSV0_0;
	wire w_dff_A_Z7a0zdQI7_0;
	wire w_dff_A_JKlPqns47_0;
	wire w_dff_A_NPlDhGk86_0;
	wire w_dff_A_Z5CYrWyN0_0;
	wire w_dff_A_o63knkld1_0;
	wire w_dff_A_OeGHYLmr5_0;
	wire w_dff_A_EVSH4rOi8_0;
	wire w_dff_A_WG0SuF1k2_0;
	wire w_dff_A_4pK8wCXV0_0;
	wire w_dff_A_e7ox6w9F9_0;
	wire w_dff_A_Z0c9FQ7z3_0;
	wire w_dff_A_mPX9ATHL6_0;
	wire w_dff_A_hc8aJAzE8_0;
	wire w_dff_A_g5PN8qbD9_0;
	wire w_dff_A_S97nMcH87_0;
	wire w_dff_A_2CuGPe2C3_0;
	wire w_dff_A_MMM98mI96_2;
	wire w_dff_A_YrGIIctL5_0;
	wire w_dff_A_orUO2Ost2_0;
	wire w_dff_A_YdwBZwp39_0;
	wire w_dff_A_OZFTCYku7_0;
	wire w_dff_A_cssR2C1c8_0;
	wire w_dff_A_FfGxyauN6_0;
	wire w_dff_A_53HRLule7_0;
	wire w_dff_A_o12pm6UI9_0;
	wire w_dff_A_PqmNOBEM2_0;
	wire w_dff_A_ThQHPZvC2_0;
	wire w_dff_A_ko0gb4Uk0_0;
	wire w_dff_A_SSBgdHsN2_0;
	wire w_dff_A_NkCpB6At9_0;
	wire w_dff_A_I3XUg78F4_0;
	wire w_dff_A_csKpg7Vr3_0;
	wire w_dff_A_8PAszGGU4_0;
	wire w_dff_A_69Tfxs4k6_0;
	wire w_dff_A_AG6pyT1G1_0;
	wire w_dff_A_XrDOxc951_0;
	wire w_dff_A_qOIsBatc1_0;
	wire w_dff_A_zxLaVc240_0;
	wire w_dff_A_CwuYsNzx1_0;
	wire w_dff_A_rBcBKz039_0;
	wire w_dff_A_pVqNiwPA5_2;
	wire w_dff_A_TPRssbmc8_0;
	wire w_dff_A_s5w8MOP58_0;
	wire w_dff_A_ImsFZWhO1_0;
	wire w_dff_A_qMgARpnT2_0;
	wire w_dff_A_eTu77bM78_0;
	wire w_dff_A_011DCSol9_0;
	wire w_dff_A_gx0RmkDW7_0;
	wire w_dff_A_EOnlBFNd4_0;
	wire w_dff_A_1BfvGWRs3_0;
	wire w_dff_A_OPG2z6hB5_0;
	wire w_dff_A_6vdob3ul3_0;
	wire w_dff_A_pfdSVIcz9_0;
	wire w_dff_A_O4NSYRy27_0;
	wire w_dff_A_m84hN0bh5_2;
	wire w_dff_A_6UGpNuVA1_0;
	wire w_dff_A_dM8FEHoY5_0;
	wire w_dff_A_ZPtrLbS69_0;
	wire w_dff_A_uF27NlyY1_0;
	wire w_dff_A_ALf8UQqd3_0;
	wire w_dff_A_U65q1uSE1_0;
	wire w_dff_A_BRMIDGBu3_0;
	wire w_dff_A_qlaIbqXv0_0;
	wire w_dff_A_EDn6K2rB2_0;
	wire w_dff_A_dV9SLUXR1_0;
	wire w_dff_A_zAvXALRF6_0;
	wire w_dff_A_m8XhH8tq7_2;
	wire w_dff_A_m9IwkISh1_0;
	wire w_dff_A_qzfDZh0X6_0;
	wire w_dff_A_cm4dQeg76_0;
	wire w_dff_A_hksdxLHH8_0;
	wire w_dff_A_hzpk3Q5F4_0;
	wire w_dff_A_OSBCI5aM6_0;
	wire w_dff_A_qMmPkybN2_0;
	wire w_dff_A_c020QNlg6_0;
	wire w_dff_A_roHWtaR75_0;
	wire w_dff_A_5113JSsV7_0;
	wire w_dff_A_suxkJc9W4_2;
	wire w_dff_A_Z8JREjjN9_0;
	wire w_dff_A_7pgYwA4l1_0;
	wire w_dff_A_0FQj6WAO3_0;
	wire w_dff_A_ofbc0hAk3_0;
	wire w_dff_A_76SFJWpT8_0;
	wire w_dff_A_3yh6VbIy4_0;
	wire w_dff_A_YA1W9wn41_0;
	wire w_dff_A_OJoT2UhP0_0;
	wire w_dff_A_lgEufWyi0_0;
	wire w_dff_A_FH1rm7wP5_0;
	wire w_dff_A_QVGVQfYK5_2;
	wire w_dff_A_pO225CQ91_0;
	wire w_dff_A_pM3r58Os8_0;
	wire w_dff_A_XQxYVzmv4_0;
	wire w_dff_A_ZkoGnkeN7_0;
	wire w_dff_A_8yzMmy9m2_0;
	wire w_dff_A_37tdttyl5_0;
	wire w_dff_A_TBeJSWGG1_0;
	wire w_dff_A_5THm0ccg7_0;
	wire w_dff_A_3mqd2LSB1_0;
	wire w_dff_A_TTs0Ebo48_0;
	wire w_dff_A_CAs6wypP0_1;
	wire w_dff_A_04yIwS3a1_0;
	wire w_dff_A_xjM1qNsL6_0;
	wire w_dff_A_Y0gcCkcp8_0;
	wire w_dff_A_RDkaEOis8_0;
	wire w_dff_A_Z6Sxk4LA1_0;
	wire w_dff_A_zSE96s8W0_0;
	wire w_dff_A_J1Db1Fso2_0;
	wire w_dff_A_8Faaqfu06_2;
	wire w_dff_A_fgvTXq5c7_0;
	wire w_dff_A_SqT9QFom1_0;
	wire w_dff_A_VQjg5Bf97_0;
	wire w_dff_A_uvV2URYd5_0;
	wire w_dff_A_iCSTSP0S7_2;
	wire w_dff_A_pbvNBtfW3_0;
	wire w_dff_A_j05d5K929_0;
	wire w_dff_A_CYRV8SvA9_0;
	wire w_dff_A_RTDFHfRV3_0;
	wire w_dff_A_QIL9dh5f4_1;
	wire w_dff_A_Pc7m9k791_0;
	wire w_dff_A_uwKuCJ2R9_0;
	wire w_dff_A_Z3X71WYa8_0;
	wire w_dff_A_tzjOiDPM2_0;
	wire w_dff_A_TX9cKArf8_0;
	wire w_dff_A_yJeu9qUG8_0;
	wire w_dff_A_C8WizjaC4_1;
	wire w_dff_A_W8ZDHHB99_0;
	wire w_dff_A_zxDUn9Pe6_0;
	wire w_dff_A_jF25fous3_0;
	wire w_dff_A_cWd8y1Eo7_0;
	wire w_dff_A_x6MFrcXs1_0;
	wire w_dff_A_4BLq7DIM7_1;
	wire w_dff_A_L9dsrKyh3_0;
	wire w_dff_A_a5H6vCKM6_0;
	wire w_dff_A_eJfTlNBL5_0;
	wire w_dff_A_mUQgB1iF3_0;
	wire w_dff_A_Kdmz1GUI9_1;
	wire w_dff_A_uVGAMC2O8_0;
	wire w_dff_A_rTlkI1I64_0;
	wire w_dff_A_3TPEWlaZ5_1;
	wire w_dff_A_OpvJBNVA6_0;
	wire w_dff_A_wVG6D6Ml7_0;
	wire w_dff_A_PVlWremV5_0;
	wire w_dff_A_5wTVWcMF7_0;
	wire w_dff_A_snNc0Gbh4_1;
	wire w_dff_A_Znbnrzrt0_2;
	jnot g0000(.din(w_G77_5[1]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[1]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[1]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_1[1]),.dinb(w_n74_1[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[1]),.dout(w_dff_A_eHaXs8ak3_2),.clk(gclk));
	jnot g0007(.din(w_G97_5[1]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G107_5[1]),.dout(n80),.clk(gclk));
	jand g0009(.dina(w_n80_1[1]),.dinb(w_n79_0[2]),.dout(n81),.clk(gclk));
	jnot g0010(.din(w_n81_0[2]),.dout(n82),.clk(gclk));
	jand g0011(.dina(n82),.dinb(w_G87_3[2]),.dout(n83),.clk(gclk));
	jnot g0012(.din(n83),.dout(G355_fa_),.clk(gclk));
	jand g0013(.dina(w_G20_7[1]),.dinb(w_G1_3[1]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G226_1[1]),.dout(n86),.clk(gclk));
	jor g0015(.dina(w_n86_0[1]),.dinb(w_n73_2[1]),.dout(n87),.clk(gclk));
	jnot g0016(.din(w_G264_1[1]),.dout(n88),.clk(gclk));
	jor g0017(.dina(w_n88_1[1]),.dinb(w_n80_1[0]),.dout(n89),.clk(gclk));
	jand g0018(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jnot g0019(.din(w_G257_1[2]),.dout(n91),.clk(gclk));
	jor g0020(.dina(w_n91_1[2]),.dinb(w_n79_0[1]),.dout(n92),.clk(gclk));
	jnot g0021(.din(w_G238_1[2]),.dout(n93),.clk(gclk));
	jor g0022(.dina(w_n93_0[1]),.dinb(w_n75_1[0]),.dout(n94),.clk(gclk));
	jand g0023(.dina(n94),.dinb(n92),.dout(n95),.clk(gclk));
	jand g0024(.dina(n95),.dinb(n90),.dout(n96),.clk(gclk));
	jnot g0025(.din(w_G87_3[1]),.dout(n97),.clk(gclk));
	jnot g0026(.din(w_G250_0[2]),.dout(n98),.clk(gclk));
	jor g0027(.dina(w_n98_2[1]),.dinb(w_n97_2[1]),.dout(n99),.clk(gclk));
	jnot g0028(.din(w_G232_1[2]),.dout(n100),.clk(gclk));
	jor g0029(.dina(n100),.dinb(w_n74_1[0]),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(n99),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G244_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(w_n103_0[2]),.dinb(w_n72_1[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_4[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(w_n106_0[1]),.dinb(w_n105_2[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jand g0037(.dina(n108),.dinb(n102),.dout(n109),.clk(gclk));
	jand g0038(.dina(n109),.dinb(n96),.dout(n110),.clk(gclk));
	jor g0039(.dina(n110),.dinb(w_n85_0[2]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_G20_7[0]),.dout(n112),.clk(gclk));
	jnot g0041(.din(w_G1_3[0]),.dout(n113),.clk(gclk));
	jnot g0042(.din(w_G13_1[1]),.dout(n114),.clk(gclk));
	jor g0043(.dina(w_n114_1[2]),.dinb(w_n113_3[1]),.dout(n115),.clk(gclk));
	jor g0044(.dina(w_n115_1[1]),.dinb(w_n112_5[2]),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jor g0048(.dina(n119),.dinb(w_n116_0[1]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n114_1[1]),.dinb(w_G1_2[2]),.dout(n121),.clk(gclk));
	jand g0050(.dina(w_n121_0[2]),.dinb(w_G20_6[2]),.dout(n122),.clk(gclk));
	jnot g0051(.din(w_n122_1[1]),.dout(n123),.clk(gclk));
	jand g0052(.dina(w_n88_1[0]),.dinb(w_n91_1[1]),.dout(n124),.clk(gclk));
	jor g0053(.dina(n124),.dinb(w_n98_2[0]),.dout(n125),.clk(gclk));
	jor g0054(.dina(n125),.dinb(w_n123_1[2]),.dout(n126),.clk(gclk));
	jand g0055(.dina(n126),.dinb(n120),.dout(n127),.clk(gclk));
	jand g0056(.dina(n127),.dinb(w_dff_B_M2bk8CTR9_1),.dout(w_dff_A_6n9RzDAU9_2),.clk(gclk));
	jxor g0057(.dina(w_G270_0[1]),.dinb(w_G264_1[0]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_G257_1[1]),.dinb(w_n98_1[2]),.dout(n130),.clk(gclk));
	jxor g0059(.dina(n130),.dinb(n129),.dout(n131),.clk(gclk));
	jnot g0060(.din(w_n131_0[1]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G244_1[1]),.dinb(w_G238_1[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(w_G232_1[1]),.dinb(w_n86_0[0]),.dout(n134),.clk(gclk));
	jxor g0063(.dina(n134),.dinb(n133),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_n135_0[1]),.dinb(n132),.dout(w_dff_A_x8w3OkNr6_2),.clk(gclk));
	jxor g0065(.dina(w_G68_5[0]),.dinb(w_G58_5[0]),.dout(n137),.clk(gclk));
	jnot g0066(.din(w_n137_0[2]),.dout(n138),.clk(gclk));
	jxor g0067(.dina(w_G77_5[0]),.dinb(w_G50_5[0]),.dout(n139),.clk(gclk));
	jxor g0068(.dina(n139),.dinb(n138),.dout(n140),.clk(gclk));
	jnot g0069(.din(w_n140_0[1]),.dout(n141),.clk(gclk));
	jxor g0070(.dina(w_G116_4[1]),.dinb(w_G107_5[0]),.dout(n142),.clk(gclk));
	jxor g0071(.dina(w_G97_5[0]),.dinb(w_n97_2[0]),.dout(n143),.clk(gclk));
	jxor g0072(.dina(n143),.dinb(n142),.dout(n144),.clk(gclk));
	jxor g0073(.dina(w_n144_0[1]),.dinb(n141),.dout(w_dff_A_MMM98mI96_2),.clk(gclk));
	jnot g0074(.din(w_G169_1[1]),.dout(n146),.clk(gclk));
	jand g0075(.dina(w_G13_1[0]),.dinb(w_G1_2[1]),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_G33_11[2]),.dout(n148),.clk(gclk));
	jnot g0077(.din(w_G41_1[1]),.dout(n149),.clk(gclk));
	jor g0078(.dina(w_n149_2[1]),.dinb(w_n148_9[2]),.dout(n150),.clk(gclk));
	jand g0079(.dina(n150),.dinb(w_n147_0[2]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G1698_0[2]),.dinb(w_n148_9[1]),.dout(n152),.clk(gclk));
	jand g0081(.dina(w_n152_3[1]),.dinb(w_G244_1[0]),.dout(n153),.clk(gclk));
	jnot g0082(.din(w_G1698_0[1]),.dout(n154),.clk(gclk));
	jand g0083(.dina(w_n154_0[1]),.dinb(w_n148_9[0]),.dout(n155),.clk(gclk));
	jand g0084(.dina(w_n155_3[1]),.dinb(w_G238_1[0]),.dout(n156),.clk(gclk));
	jand g0085(.dina(w_G116_4[0]),.dinb(w_G33_11[1]),.dout(n157),.clk(gclk));
	jor g0086(.dina(w_n157_0[2]),.dinb(n156),.dout(n158),.clk(gclk));
	jor g0087(.dina(n158),.dinb(n153),.dout(n159),.clk(gclk));
	jand g0088(.dina(n159),.dinb(w_n151_4[2]),.dout(n160),.clk(gclk));
	jnot g0089(.din(w_G45_1[2]),.dout(n161),.clk(gclk));
	jor g0090(.dina(w_n161_1[1]),.dinb(w_G1_2[0]),.dout(n162),.clk(gclk));
	jand g0091(.dina(w_n162_0[2]),.dinb(w_n98_1[1]),.dout(n163),.clk(gclk));
	jnot g0092(.din(w_n163_0[1]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_G41_1[0]),.dinb(w_G33_11[0]),.dout(n165),.clk(gclk));
	jor g0094(.dina(n165),.dinb(w_n115_1[0]),.dout(n166),.clk(gclk));
	jor g0095(.dina(w_n162_0[1]),.dinb(w_G274_0[2]),.dout(n167),.clk(gclk));
	jand g0096(.dina(n167),.dinb(w_n166_3[1]),.dout(n168),.clk(gclk));
	jand g0097(.dina(n168),.dinb(n164),.dout(n169),.clk(gclk));
	jor g0098(.dina(n169),.dinb(n160),.dout(n170),.clk(gclk));
	jand g0099(.dina(w_n170_0[2]),.dinb(w_n146_3[2]),.dout(n171),.clk(gclk));
	jand g0100(.dina(w_G97_4[2]),.dinb(w_G33_10[2]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G68_4[2]),.dinb(w_n148_8[2]),.dout(n173),.clk(gclk));
	jor g0102(.dina(n173),.dinb(w_G20_6[1]),.dout(n174),.clk(gclk));
	jor g0103(.dina(n174),.dinb(w_n172_0[1]),.dout(n175),.clk(gclk));
	jnot g0104(.din(n175),.dout(n176),.clk(gclk));
	jor g0105(.dina(w_n112_5[1]),.dinb(w_n113_3[0]),.dout(n177),.clk(gclk));
	jor g0106(.dina(n177),.dinb(w_n148_8[1]),.dout(n178),.clk(gclk));
	jand g0107(.dina(n178),.dinb(w_n115_0[2]),.dout(n179),.clk(gclk));
	jand g0108(.dina(w_n81_0[1]),.dinb(w_n97_1[2]),.dout(n180),.clk(gclk));
	jand g0109(.dina(w_n180_0[1]),.dinb(w_G20_6[0]),.dout(n181),.clk(gclk));
	jor g0110(.dina(n181),.dinb(w_n179_1[2]),.dout(n182),.clk(gclk));
	jor g0111(.dina(n182),.dinb(n176),.dout(n183),.clk(gclk));
	jand g0112(.dina(w_G20_5[2]),.dinb(w_n113_2[2]),.dout(n184),.clk(gclk));
	jand g0113(.dina(n184),.dinb(w_G13_0[2]),.dout(n185),.clk(gclk));
	jand g0114(.dina(w_n185_3[2]),.dinb(w_n97_1[1]),.dout(n186),.clk(gclk));
	jnot g0115(.din(n186),.dout(n187),.clk(gclk));
	jand g0116(.dina(w_n85_0[1]),.dinb(w_G33_10[1]),.dout(n188),.clk(gclk));
	jor g0117(.dina(n188),.dinb(w_n147_0[1]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n185_3[1]),.dinb(w_n189_2[1]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_G33_10[0]),.dinb(w_n113_2[1]),.dout(n191),.clk(gclk));
	jor g0120(.dina(w_n191_0[2]),.dinb(w_n97_1[0]),.dout(n192),.clk(gclk));
	jor g0121(.dina(n192),.dinb(w_n190_1[2]),.dout(n193),.clk(gclk));
	jand g0122(.dina(n193),.dinb(n187),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(n183),.dout(n195),.clk(gclk));
	jnot g0124(.din(w_G179_2[2]),.dout(n196),.clk(gclk));
	jor g0125(.dina(w_n154_0[0]),.dinb(w_G33_9[2]),.dout(n197),.clk(gclk));
	jor g0126(.dina(w_n197_1[1]),.dinb(w_n103_0[1]),.dout(n198),.clk(gclk));
	jor g0127(.dina(w_G1698_0[0]),.dinb(w_G33_9[1]),.dout(n199),.clk(gclk));
	jor g0128(.dina(w_n199_1[1]),.dinb(w_n93_0[0]),.dout(n200),.clk(gclk));
	jnot g0129(.din(w_n157_0[1]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n201_0[1]),.dinb(n200),.dout(n202),.clk(gclk));
	jand g0131(.dina(n202),.dinb(n198),.dout(n203),.clk(gclk));
	jor g0132(.dina(n203),.dinb(w_n166_3[0]),.dout(n204),.clk(gclk));
	jnot g0133(.din(w_G274_0[1]),.dout(n205),.clk(gclk));
	jand g0134(.dina(w_G45_1[1]),.dinb(w_n113_2[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(w_n206_0[1]),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jor g0136(.dina(n207),.dinb(w_n151_4[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n163_0[0]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(n204),.dout(n210),.clk(gclk));
	jand g0139(.dina(w_n210_0[2]),.dinb(w_n196_2[2]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n195_0[1]),.dout(n212),.clk(gclk));
	jor g0141(.dina(n212),.dinb(n171),.dout(n213),.clk(gclk));
	jnot g0142(.din(w_n195_0[0]),.dout(n214),.clk(gclk));
	jand g0143(.dina(w_n210_0[1]),.dinb(w_G190_4[1]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n170_0[1]),.dinb(w_G200_4[2]),.dout(n216),.clk(gclk));
	jor g0145(.dina(n216),.dinb(n215),.dout(n217),.clk(gclk));
	jor g0146(.dina(n217),.dinb(w_n214_0[1]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_n218_0[1]),.dinb(w_n213_0[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(w_n197_1[0]),.dinb(w_n98_1[0]),.dout(n220),.clk(gclk));
	jand g0149(.dina(w_G283_3[2]),.dinb(w_G33_9[0]),.dout(n221),.clk(gclk));
	jnot g0150(.din(w_n221_0[2]),.dout(n222),.clk(gclk));
	jor g0151(.dina(w_n199_1[0]),.dinb(w_n103_0[0]),.dout(n223),.clk(gclk));
	jand g0152(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jand g0153(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jor g0154(.dina(n225),.dinb(w_n166_2[2]),.dout(n226),.clk(gclk));
	jor g0155(.dina(w_n151_4[0]),.dinb(w_n205_0[0]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n162_0[0]),.dinb(w_G41_0[2]),.dout(n228),.clk(gclk));
	jor g0157(.dina(w_n228_0[1]),.dinb(n227),.dout(n229),.clk(gclk));
	jand g0158(.dina(w_n206_0[0]),.dinb(w_n149_2[0]),.dout(n230),.clk(gclk));
	jor g0159(.dina(w_n230_0[1]),.dinb(w_n151_3[2]),.dout(n231),.clk(gclk));
	jor g0160(.dina(w_n231_0[2]),.dinb(w_n91_1[0]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[2]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(n226),.dout(n234),.clk(gclk));
	jor g0163(.dina(w_n234_0[2]),.dinb(w_n146_3[1]),.dout(n235),.clk(gclk));
	jand g0164(.dina(w_n152_3[0]),.dinb(w_G250_0[1]),.dout(n236),.clk(gclk));
	jand g0165(.dina(w_n155_3[0]),.dinb(w_G244_0[2]),.dout(n237),.clk(gclk));
	jor g0166(.dina(n237),.dinb(w_n221_0[1]),.dout(n238),.clk(gclk));
	jor g0167(.dina(n238),.dinb(n236),.dout(n239),.clk(gclk));
	jand g0168(.dina(n239),.dinb(w_n151_3[1]),.dout(n240),.clk(gclk));
	jand g0169(.dina(w_n166_2[1]),.dinb(w_G274_0[0]),.dout(n241),.clk(gclk));
	jand g0170(.dina(w_n230_0[0]),.dinb(w_n241_0[1]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n228_0[0]),.dinb(w_n166_2[0]),.dout(n243),.clk(gclk));
	jand g0172(.dina(w_n243_0[2]),.dinb(w_G257_1[0]),.dout(n244),.clk(gclk));
	jor g0173(.dina(n244),.dinb(w_n242_0[2]),.dout(n245),.clk(gclk));
	jor g0174(.dina(n245),.dinb(n240),.dout(n246),.clk(gclk));
	jor g0175(.dina(w_n246_1[1]),.dinb(w_n196_2[1]),.dout(n247),.clk(gclk));
	jand g0176(.dina(n247),.dinb(n235),.dout(n248),.clk(gclk));
	jand g0177(.dina(w_G107_4[2]),.dinb(w_G33_8[2]),.dout(n249),.clk(gclk));
	jand g0178(.dina(w_G77_4[2]),.dinb(w_n148_8[0]),.dout(n250),.clk(gclk));
	jor g0179(.dina(n250),.dinb(w_G20_5[1]),.dout(n251),.clk(gclk));
	jor g0180(.dina(n251),.dinb(w_n249_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(w_G107_4[1]),.dinb(w_G97_4[1]),.dout(n253),.clk(gclk));
	jor g0182(.dina(n253),.dinb(w_n112_5[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(w_n81_0[0]),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_0[1]),.dinb(n252),.dout(n256),.clk(gclk));
	jand g0185(.dina(n256),.dinb(w_n189_2[0]),.dout(n257),.clk(gclk));
	jnot g0186(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g0187(.dina(w_n185_3[0]),.dinb(w_n79_0[0]),.dout(n259),.clk(gclk));
	jnot g0188(.din(w_n259_0[1]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n191_0[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_n261_0[1]),.dinb(w_G97_4[0]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[1]),.dout(n263),.clk(gclk));
	jor g0192(.dina(n263),.dinb(w_n190_1[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(n260),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(n258),.dout(n266),.clk(gclk));
	jor g0195(.dina(n266),.dinb(n248),.dout(n267),.clk(gclk));
	jand g0196(.dina(w_n246_1[0]),.dinb(w_G200_4[1]),.dout(n268),.clk(gclk));
	jor g0197(.dina(w_n112_4[2]),.dinb(w_G1_1[2]),.dout(n269),.clk(gclk));
	jor g0198(.dina(w_n269_1[2]),.dinb(w_n114_1[0]),.dout(n270),.clk(gclk));
	jand g0199(.dina(w_n270_0[1]),.dinb(w_n179_1[1]),.dout(n271),.clk(gclk));
	jand g0200(.dina(w_n262_0[0]),.dinb(w_n271_1[2]),.dout(n272),.clk(gclk));
	jor g0201(.dina(n272),.dinb(w_n259_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n257_0[0]),.dout(n274),.clk(gclk));
	jand g0203(.dina(w_n234_0[1]),.dinb(w_G190_4[0]),.dout(n275),.clk(gclk));
	jor g0204(.dina(n275),.dinb(w_n274_0[2]),.dout(n276),.clk(gclk));
	jor g0205(.dina(n276),.dinb(n268),.dout(n277),.clk(gclk));
	jand g0206(.dina(n277),.dinb(n267),.dout(n278),.clk(gclk));
	jand g0207(.dina(w_n278_0[1]),.dinb(w_n219_0[1]),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n152_2[2]),.dinb(w_G264_0[2]),.dout(n280),.clk(gclk));
	jand g0209(.dina(w_G303_2[2]),.dinb(w_G33_8[1]),.dout(n281),.clk(gclk));
	jand g0210(.dina(w_n155_2[2]),.dinb(w_G257_0[2]),.dout(n282),.clk(gclk));
	jor g0211(.dina(n282),.dinb(w_n281_0[1]),.dout(n283),.clk(gclk));
	jor g0212(.dina(n283),.dinb(n280),.dout(n284),.clk(gclk));
	jand g0213(.dina(n284),.dinb(w_n151_3[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_n243_0[1]),.dinb(w_G270_0[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_n242_0[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(n285),.dout(n288),.clk(gclk));
	jand g0217(.dina(w_n288_1[1]),.dinb(w_n146_3[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(w_G97_3[2]),.dinb(w_n148_7[2]),.dout(n290),.clk(gclk));
	jor g0219(.dina(n290),.dinb(w_G20_5[0]),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(w_n221_0[0]),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n105_2[0]),.dinb(w_G20_4[2]),.dout(n293),.clk(gclk));
	jnot g0222(.din(n293),.dout(n294),.clk(gclk));
	jand g0223(.dina(n294),.dinb(w_n189_1[2]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(n292),.dout(n296),.clk(gclk));
	jnot g0225(.din(w_n296_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(w_n185_2[2]),.dinb(w_n105_1[2]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n191_0[0]),.dinb(w_n105_1[1]),.dout(n300),.clk(gclk));
	jor g0229(.dina(w_n300_0[1]),.dinb(w_n190_1[0]),.dout(n301),.clk(gclk));
	jand g0230(.dina(n301),.dinb(n299),.dout(n302),.clk(gclk));
	jand g0231(.dina(n302),.dinb(n297),.dout(n303),.clk(gclk));
	jor g0232(.dina(w_n197_0[2]),.dinb(w_n88_0[2]),.dout(n304),.clk(gclk));
	jnot g0233(.din(w_n281_0[0]),.dout(n305),.clk(gclk));
	jor g0234(.dina(w_n199_0[2]),.dinb(w_n91_0[2]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(n305),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n304),.dout(n308),.clk(gclk));
	jor g0237(.dina(n308),.dinb(w_n166_1[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n231_0[1]),.dinb(w_n106_0[0]),.dout(n310),.clk(gclk));
	jand g0239(.dina(n310),.dinb(w_n229_0[1]),.dout(n311),.clk(gclk));
	jand g0240(.dina(n311),.dinb(n309),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_1[1]),.dinb(w_n196_2[0]),.dout(n313),.clk(gclk));
	jor g0242(.dina(n313),.dinb(w_n303_0[1]),.dout(n314),.clk(gclk));
	jor g0243(.dina(n314),.dinb(n289),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_n288_1[0]),.dinb(w_G200_4[0]),.dout(n316),.clk(gclk));
	jnot g0245(.din(w_n300_0[0]),.dout(n317),.clk(gclk));
	jand g0246(.dina(n317),.dinb(w_n271_1[1]),.dout(n318),.clk(gclk));
	jor g0247(.dina(n318),.dinb(w_n298_0[0]),.dout(n319),.clk(gclk));
	jor g0248(.dina(n319),.dinb(w_n296_0[0]),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n312_1[0]),.dinb(w_G190_3[2]),.dout(n321),.clk(gclk));
	jor g0250(.dina(n321),.dinb(w_n320_0[1]),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(n316),.dout(n323),.clk(gclk));
	jand g0252(.dina(n323),.dinb(w_n315_0[1]),.dout(n324),.clk(gclk));
	jor g0253(.dina(w_n97_0[2]),.dinb(w_G33_8[0]),.dout(n325),.clk(gclk));
	jand g0254(.dina(n325),.dinb(w_n112_4[1]),.dout(n326),.clk(gclk));
	jand g0255(.dina(n326),.dinb(w_n201_0[0]),.dout(n327),.clk(gclk));
	jor g0256(.dina(n327),.dinb(w_n179_1[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(w_n328_0[1]),.dinb(w_G20_4[1]),.dout(n329),.clk(gclk));
	jand g0258(.dina(n329),.dinb(w_G107_4[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n328_0[0]),.dinb(w_n270_0[0]),.dout(n331),.clk(gclk));
	jor g0260(.dina(n331),.dinb(n330),.dout(n332),.clk(gclk));
	jand g0261(.dina(w_n261_0[0]),.dinb(w_G107_3[2]),.dout(n333),.clk(gclk));
	jand g0262(.dina(n333),.dinb(w_n271_1[0]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jand g0264(.dina(n335),.dinb(n332),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n197_0[1]),.dinb(w_n91_0[1]),.dout(n337),.clk(gclk));
	jor g0266(.dina(w_n199_0[1]),.dinb(w_n98_0[2]),.dout(n338),.clk(gclk));
	jand g0267(.dina(w_G294_3[1]),.dinb(w_G33_7[2]),.dout(n339),.clk(gclk));
	jnot g0268(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jand g0269(.dina(n340),.dinb(n338),.dout(n341),.clk(gclk));
	jand g0270(.dina(n341),.dinb(n337),.dout(n342),.clk(gclk));
	jor g0271(.dina(n342),.dinb(w_n166_1[1]),.dout(n343),.clk(gclk));
	jor g0272(.dina(w_n231_0[0]),.dinb(w_n88_0[1]),.dout(n344),.clk(gclk));
	jand g0273(.dina(n344),.dinb(w_n229_0[0]),.dout(n345),.clk(gclk));
	jand g0274(.dina(n345),.dinb(n343),.dout(n346),.clk(gclk));
	jand g0275(.dina(w_n346_1[1]),.dinb(w_n196_1[2]),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n152_2[1]),.dinb(w_G257_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n155_2[1]),.dinb(w_G250_0[0]),.dout(n349),.clk(gclk));
	jor g0278(.dina(w_n339_0[0]),.dinb(n349),.dout(n350),.clk(gclk));
	jor g0279(.dina(n350),.dinb(n348),.dout(n351),.clk(gclk));
	jand g0280(.dina(n351),.dinb(w_n151_2[2]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n243_0[0]),.dinb(w_G264_0[1]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_n242_0[0]),.dout(n354),.clk(gclk));
	jor g0283(.dina(n354),.dinb(n352),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_1[1]),.dinb(w_n146_2[2]),.dout(n356),.clk(gclk));
	jor g0285(.dina(n356),.dinb(n347),.dout(n357),.clk(gclk));
	jor g0286(.dina(n357),.dinb(n336),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_G87_3[0]),.dinb(w_n148_7[1]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_G20_4[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(w_n157_0[0]),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n189_1[1]),.dout(n362),.clk(gclk));
	jand g0291(.dina(w_n362_0[1]),.dinb(w_n112_4[0]),.dout(n363),.clk(gclk));
	jor g0292(.dina(n363),.dinb(w_n80_0[2]),.dout(n364),.clk(gclk));
	jor g0293(.dina(w_n362_0[0]),.dinb(w_n185_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(n365),.dinb(n364),.dout(n366),.clk(gclk));
	jor g0295(.dina(w_n334_0[0]),.dinb(n366),.dout(n367),.clk(gclk));
	jor g0296(.dina(w_n355_1[0]),.dinb(w_G190_3[1]),.dout(n368),.clk(gclk));
	jor g0297(.dina(w_n346_1[0]),.dinb(w_G200_3[2]),.dout(n369),.clk(gclk));
	jand g0298(.dina(n369),.dinb(n368),.dout(n370),.clk(gclk));
	jor g0299(.dina(n370),.dinb(w_n367_0[2]),.dout(n371),.clk(gclk));
	jand g0300(.dina(w_n371_0[1]),.dinb(n358),.dout(n372),.clk(gclk));
	jand g0301(.dina(w_n372_0[1]),.dinb(w_n324_0[1]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n279_0[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n155_2[0]),.dinb(w_G232_1[0]),.dout(n375),.clk(gclk));
	jand g0304(.dina(w_n152_2[0]),.dinb(w_G238_0[2]),.dout(n376),.clk(gclk));
	jor g0305(.dina(n376),.dinb(w_n249_0[0]),.dout(n377),.clk(gclk));
	jor g0306(.dina(n377),.dinb(n375),.dout(n378),.clk(gclk));
	jand g0307(.dina(n378),.dinb(w_n151_2[1]),.dout(n379),.clk(gclk));
	jand g0308(.dina(w_n161_1[0]),.dinb(w_n149_1[2]),.dout(n380),.clk(gclk));
	jor g0309(.dina(n380),.dinb(w_G1_1[1]),.dout(n381),.clk(gclk));
	jand g0310(.dina(w_n381_0[1]),.dinb(w_n166_1[0]),.dout(n382),.clk(gclk));
	jand g0311(.dina(w_n382_1[1]),.dinb(w_G244_0[1]),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n381_0[0]),.dout(n384),.clk(gclk));
	jand g0313(.dina(n384),.dinb(w_n241_0[0]),.dout(n385),.clk(gclk));
	jor g0314(.dina(w_n385_1[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n379),.dout(n387),.clk(gclk));
	jand g0316(.dina(w_n387_1[1]),.dinb(w_n146_2[1]),.dout(n388),.clk(gclk));
	jnot g0317(.din(n388),.dout(n389),.clk(gclk));
	jand g0318(.dina(w_G87_2[2]),.dinb(w_G33_7[1]),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_G58_4[2]),.dinb(w_n148_7[0]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_G20_3[2]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(w_n390_0[1]),.dout(n393),.clk(gclk));
	jor g0322(.dina(w_G77_4[1]),.dinb(w_n112_3[2]),.dout(n394),.clk(gclk));
	jand g0323(.dina(n394),.dinb(w_n189_1[0]),.dout(n395),.clk(gclk));
	jand g0324(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0325(.dina(w_n185_2[0]),.dinb(w_n72_0[2]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n269_1[1]),.dinb(w_G77_4[0]),.dout(n398),.clk(gclk));
	jand g0327(.dina(n398),.dinb(w_n271_0[2]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(n397),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(n396),.dout(n401),.clk(gclk));
	jor g0330(.dina(w_n387_1[0]),.dinb(w_G179_2[1]),.dout(n402),.clk(gclk));
	jand g0331(.dina(n402),.dinb(w_n401_0[2]),.dout(n403),.clk(gclk));
	jand g0332(.dina(n403),.dinb(n389),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jand g0334(.dina(w_n387_0[2]),.dinb(w_G200_3[1]),.dout(n406),.clk(gclk));
	jnot g0335(.din(w_G190_3[0]),.dout(n407),.clk(gclk));
	jor g0336(.dina(w_n387_0[1]),.dinb(w_n407_2[1]),.dout(n408),.clk(gclk));
	jnot g0337(.din(n408),.dout(n409),.clk(gclk));
	jor g0338(.dina(n409),.dinb(w_n401_0[1]),.dout(n410),.clk(gclk));
	jor g0339(.dina(n410),.dinb(n406),.dout(n411),.clk(gclk));
	jand g0340(.dina(n411),.dinb(w_n405_0[1]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_n155_1[2]),.dinb(w_G226_1[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n152_1[2]),.dinb(w_G232_0[2]),.dout(n414),.clk(gclk));
	jor g0343(.dina(n414),.dinb(w_n172_0[0]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(n413),.dout(n416),.clk(gclk));
	jand g0345(.dina(n416),.dinb(w_n151_2[0]),.dout(n417),.clk(gclk));
	jand g0346(.dina(w_n382_1[0]),.dinb(w_G238_0[1]),.dout(n418),.clk(gclk));
	jor g0347(.dina(n418),.dinb(w_n385_1[0]),.dout(n419),.clk(gclk));
	jor g0348(.dina(n419),.dinb(n417),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n420_1[1]),.dinb(w_n146_2[0]),.dout(n421),.clk(gclk));
	jnot g0350(.din(n421),.dout(n422),.clk(gclk));
	jand g0351(.dina(w_n269_1[0]),.dinb(w_G68_4[1]),.dout(n423),.clk(gclk));
	jand g0352(.dina(n423),.dinb(w_n271_0[1]),.dout(n424),.clk(gclk));
	jand g0353(.dina(w_n148_6[2]),.dinb(w_n114_0[2]),.dout(n425),.clk(gclk));
	jnot g0354(.din(w_n425_1[2]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n426_0[1]),.dinb(w_n85_0[0]),.dout(n427),.clk(gclk));
	jor g0356(.dina(n427),.dinb(w_n185_1[2]),.dout(n428),.clk(gclk));
	jand g0357(.dina(n428),.dinb(w_n75_0[2]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_G77_3[2]),.dinb(w_G33_7[0]),.dout(n430),.clk(gclk));
	jand g0359(.dina(w_G50_4[2]),.dinb(w_n148_6[1]),.dout(n431),.clk(gclk));
	jor g0360(.dina(n431),.dinb(w_n430_0[1]),.dout(n432),.clk(gclk));
	jand g0361(.dina(n432),.dinb(w_n112_3[1]),.dout(n433),.clk(gclk));
	jand g0362(.dina(n433),.dinb(w_n189_0[2]),.dout(n434),.clk(gclk));
	jor g0363(.dina(n434),.dinb(n429),.dout(n435),.clk(gclk));
	jor g0364(.dina(n435),.dinb(n424),.dout(n436),.clk(gclk));
	jor g0365(.dina(w_n420_1[0]),.dinb(w_G179_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n436_0[2]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(n422),.dout(n439),.clk(gclk));
	jnot g0368(.din(w_n439_1[1]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_n420_0[2]),.dinb(w_G200_3[0]),.dout(n441),.clk(gclk));
	jor g0370(.dina(w_n420_0[1]),.dinb(w_n407_2[0]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(n443),.dinb(w_n436_0[1]),.dout(n444),.clk(gclk));
	jor g0373(.dina(n444),.dinb(n441),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(n440),.dout(n446),.clk(gclk));
	jand g0375(.dina(w_n446_0[1]),.dinb(w_n412_0[1]),.dout(n447),.clk(gclk));
	jand g0376(.dina(w_n152_1[1]),.dinb(w_G223_0[1]),.dout(n448),.clk(gclk));
	jand g0377(.dina(w_n155_1[1]),.dinb(G222),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n430_0[0]),.dout(n450),.clk(gclk));
	jor g0379(.dina(n450),.dinb(n448),.dout(n451),.clk(gclk));
	jand g0380(.dina(n451),.dinb(w_n151_1[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n382_0[2]),.dinb(w_G226_0[2]),.dout(n453),.clk(gclk));
	jor g0382(.dina(n453),.dinb(w_n385_0[2]),.dout(n454),.clk(gclk));
	jor g0383(.dina(n454),.dinb(n452),.dout(n455),.clk(gclk));
	jand g0384(.dina(w_n455_0[2]),.dinb(w_n146_1[2]),.dout(n456),.clk(gclk));
	jand g0385(.dina(w_n269_0[2]),.dinb(w_G50_4[1]),.dout(n457),.clk(gclk));
	jnot g0386(.din(n457),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n190_0[2]),.dout(n459),.clk(gclk));
	jor g0388(.dina(w_n77_0[0]),.dinb(w_n112_3[0]),.dout(n460),.clk(gclk));
	jnot g0389(.din(w_G150_3[1]),.dout(n461),.clk(gclk));
	jand g0390(.dina(w_n148_6[0]),.dinb(w_n112_2[2]),.dout(n462),.clk(gclk));
	jnot g0391(.din(w_n462_0[2]),.dout(n463),.clk(gclk));
	jor g0392(.dina(n463),.dinb(n461),.dout(n464),.clk(gclk));
	jand g0393(.dina(w_G33_6[2]),.dinb(w_n112_2[1]),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n465_0[1]),.dinb(w_G58_4[1]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jand g0396(.dina(n467),.dinb(n464),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(n460),.dout(n469),.clk(gclk));
	jor g0398(.dina(n469),.dinb(w_n179_0[2]),.dout(n470),.clk(gclk));
	jand g0399(.dina(w_n185_1[1]),.dinb(w_n73_2[0]),.dout(n471),.clk(gclk));
	jnot g0400(.din(n471),.dout(n472),.clk(gclk));
	jand g0401(.dina(n472),.dinb(n470),.dout(n473),.clk(gclk));
	jand g0402(.dina(n473),.dinb(n459),.dout(n474),.clk(gclk));
	jnot g0403(.din(w_n455_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n475_0[1]),.dinb(w_n196_1[1]),.dout(n476),.clk(gclk));
	jor g0405(.dina(n476),.dinb(w_n474_0[1]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(n456),.dout(n478),.clk(gclk));
	jnot g0407(.din(w_n474_0[0]),.dout(n479),.clk(gclk));
	jand g0408(.dina(w_n475_0[0]),.dinb(w_G190_2[2]),.dout(n480),.clk(gclk));
	jand g0409(.dina(w_n455_0[0]),.dinb(w_G200_2[2]),.dout(n481),.clk(gclk));
	jor g0410(.dina(n481),.dinb(n480),.dout(n482),.clk(gclk));
	jor g0411(.dina(n482),.dinb(w_n479_0[1]),.dout(n483),.clk(gclk));
	jand g0412(.dina(w_n483_0[1]),.dinb(w_n478_0[1]),.dout(n484),.clk(gclk));
	jand g0413(.dina(w_n152_1[0]),.dinb(w_G226_0[1]),.dout(n485),.clk(gclk));
	jand g0414(.dina(w_n155_1[0]),.dinb(w_G223_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(w_n390_0[0]),.dout(n487),.clk(gclk));
	jor g0416(.dina(n487),.dinb(n485),.dout(n488),.clk(gclk));
	jand g0417(.dina(n488),.dinb(w_n151_1[1]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n382_0[1]),.dinb(w_G232_0[1]),.dout(n490),.clk(gclk));
	jor g0419(.dina(n490),.dinb(w_n385_0[1]),.dout(n491),.clk(gclk));
	jor g0420(.dina(n491),.dinb(n489),.dout(n492),.clk(gclk));
	jand g0421(.dina(w_n492_0[2]),.dinb(w_n146_1[1]),.dout(n493),.clk(gclk));
	jand g0422(.dina(w_n269_0[1]),.dinb(w_G58_4[0]),.dout(n494),.clk(gclk));
	jnot g0423(.din(n494),.dout(n495),.clk(gclk));
	jor g0424(.dina(n495),.dinb(w_n190_0[1]),.dout(n496),.clk(gclk));
	jor g0425(.dina(w_n137_0[1]),.dinb(w_n112_2[0]),.dout(n497),.clk(gclk));
	jand g0426(.dina(w_n462_0[1]),.dinb(w_G159_3[2]),.dout(n498),.clk(gclk));
	jand g0427(.dina(w_n465_0[0]),.dinb(w_G68_4[0]),.dout(n499),.clk(gclk));
	jor g0428(.dina(n499),.dinb(n498),.dout(n500),.clk(gclk));
	jnot g0429(.din(n500),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(n497),.dout(n502),.clk(gclk));
	jor g0431(.dina(n502),.dinb(w_n179_0[1]),.dout(n503),.clk(gclk));
	jand g0432(.dina(w_n185_1[0]),.dinb(w_n74_0[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(n504),.dout(n505),.clk(gclk));
	jand g0434(.dina(n505),.dinb(n503),.dout(n506),.clk(gclk));
	jand g0435(.dina(n506),.dinb(n496),.dout(n507),.clk(gclk));
	jnot g0436(.din(w_n492_0[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(w_n508_0[1]),.dinb(w_n196_1[0]),.dout(n509),.clk(gclk));
	jor g0438(.dina(n509),.dinb(w_n507_0[1]),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(n493),.dout(n511),.clk(gclk));
	jnot g0440(.din(w_n507_0[0]),.dout(n512),.clk(gclk));
	jand g0441(.dina(w_n508_0[0]),.dinb(w_G190_2[1]),.dout(n513),.clk(gclk));
	jand g0442(.dina(w_n492_0[0]),.dinb(w_G200_2[1]),.dout(n514),.clk(gclk));
	jor g0443(.dina(n514),.dinb(n513),.dout(n515),.clk(gclk));
	jor g0444(.dina(n515),.dinb(w_n512_0[1]),.dout(n516),.clk(gclk));
	jand g0445(.dina(w_n516_0[1]),.dinb(w_n511_0[1]),.dout(n517),.clk(gclk));
	jand g0446(.dina(w_n517_0[1]),.dinb(w_n484_0[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(n447),.dout(n519),.clk(gclk));
	jand g0448(.dina(w_n519_1[2]),.dinb(w_n374_0[1]),.dout(w_dff_A_pVqNiwPA5_2),.clk(gclk));
	jor g0449(.dina(w_n355_0[2]),.dinb(w_G179_1[2]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n346_0[2]),.dinb(w_G169_1[0]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(n521),.dout(n523),.clk(gclk));
	jand g0452(.dina(w_n523_0[1]),.dinb(w_n367_0[1]),.dout(n524),.clk(gclk));
	jor g0453(.dina(w_n312_0[2]),.dinb(w_G169_0[2]),.dout(n525),.clk(gclk));
	jor g0454(.dina(w_n288_0[2]),.dinb(w_G179_1[1]),.dout(n526),.clk(gclk));
	jand g0455(.dina(n526),.dinb(w_n320_0[0]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(n525),.dout(n528),.clk(gclk));
	jand g0457(.dina(w_n371_0[0]),.dinb(w_n528_0[1]),.dout(n529),.clk(gclk));
	jor g0458(.dina(n529),.dinb(w_n524_0[1]),.dout(n530),.clk(gclk));
	jand g0459(.dina(n530),.dinb(w_n279_0[0]),.dout(n531),.clk(gclk));
	jnot g0460(.din(w_n213_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(w_n246_0[2]),.dinb(w_G169_0[1]),.dout(n533),.clk(gclk));
	jand g0462(.dina(w_n234_0[0]),.dinb(w_G179_1[0]),.dout(n534),.clk(gclk));
	jor g0463(.dina(w_n534_0[1]),.dinb(n533),.dout(n535),.clk(gclk));
	jand g0464(.dina(w_n274_0[1]),.dinb(n535),.dout(n536),.clk(gclk));
	jand g0465(.dina(w_n536_0[2]),.dinb(w_n218_0[0]),.dout(n537),.clk(gclk));
	jor g0466(.dina(n537),.dinb(w_n532_0[1]),.dout(n538),.clk(gclk));
	jor g0467(.dina(n538),.dinb(n531),.dout(n539),.clk(gclk));
	jand g0468(.dina(w_n539_0[1]),.dinb(w_n519_1[1]),.dout(n540),.clk(gclk));
	jnot g0469(.din(w_n478_0[0]),.dout(n541),.clk(gclk));
	jnot g0470(.din(w_n511_0[0]),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n439_1[0]),.dinb(w_n404_0[1]),.dout(n543),.clk(gclk));
	jand g0472(.dina(w_n543_0[1]),.dinb(w_n445_0[0]),.dout(n544),.clk(gclk));
	jor g0473(.dina(n544),.dinb(w_n542_0[2]),.dout(n545),.clk(gclk));
	jand g0474(.dina(n545),.dinb(w_n516_0[0]),.dout(n546),.clk(gclk));
	jor g0475(.dina(n546),.dinb(w_n541_0[1]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n483_0[0]),.dout(n548),.clk(gclk));
	jor g0477(.dina(w_n548_0[2]),.dinb(w_dff_B_L5K1pX3c9_1),.dout(w_dff_A_m84hN0bh5_2),.clk(gclk));
	jand g0478(.dina(w_n112_1[2]),.dinb(w_G13_0[1]),.dout(n550),.clk(gclk));
	jand g0479(.dina(w_G213_0[2]),.dinb(w_n113_1[2]),.dout(n551),.clk(gclk));
	jand g0480(.dina(n551),.dinb(w_n550_0[1]),.dout(n552),.clk(gclk));
	jand g0481(.dina(w_n552_1[1]),.dinb(w_G343_0[1]),.dout(n553),.clk(gclk));
	jnot g0482(.din(w_n553_2[2]),.dout(n554),.clk(gclk));
	jand g0483(.dina(w_n554_3[2]),.dinb(w_n524_0[0]),.dout(n555),.clk(gclk));
	jand g0484(.dina(w_n554_3[1]),.dinb(w_n528_0[0]),.dout(n556),.clk(gclk));
	jand g0485(.dina(w_n553_2[1]),.dinb(w_n367_0[0]),.dout(n557),.clk(gclk));
	jnot g0486(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(w_n372_0[0]),.dout(n559),.clk(gclk));
	jand g0488(.dina(w_n557_0[0]),.dinb(w_n523_0[0]),.dout(n560),.clk(gclk));
	jor g0489(.dina(n560),.dinb(n559),.dout(n561),.clk(gclk));
	jand g0490(.dina(w_n561_0[2]),.dinb(w_n556_0[1]),.dout(n562),.clk(gclk));
	jor g0491(.dina(n562),.dinb(n555),.dout(n563),.clk(gclk));
	jnot g0492(.din(w_n561_0[1]),.dout(n564),.clk(gclk));
	jnot g0493(.din(w_G330_0[1]),.dout(n565),.clk(gclk));
	jnot g0494(.din(w_n324_0[0]),.dout(n566),.clk(gclk));
	jor g0495(.dina(w_n554_3[0]),.dinb(w_n303_0[0]),.dout(n567),.clk(gclk));
	jnot g0496(.din(w_n567_0[1]),.dout(n568),.clk(gclk));
	jor g0497(.dina(n568),.dinb(n566),.dout(n569),.clk(gclk));
	jor g0498(.dina(w_n567_0[0]),.dinb(w_n315_0[0]),.dout(n570),.clk(gclk));
	jand g0499(.dina(n570),.dinb(n569),.dout(n571),.clk(gclk));
	jor g0500(.dina(w_n571_0[2]),.dinb(w_n565_0[1]),.dout(n572),.clk(gclk));
	jor g0501(.dina(w_n572_0[2]),.dinb(w_n564_0[1]),.dout(n573),.clk(gclk));
	jnot g0502(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jor g0503(.dina(n574),.dinb(w_n563_0[2]),.dout(w_dff_A_m8XhH8tq7_2),.clk(gclk));
	jand g0504(.dina(w_n554_2[2]),.dinb(w_n539_0[0]),.dout(n576),.clk(gclk));
	jor g0505(.dina(w_n553_2[0]),.dinb(w_n374_0[0]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n346_0[1]),.dinb(w_n210_0[0]),.dout(n578),.clk(gclk));
	jand g0507(.dina(n578),.dinb(w_n312_0[1]),.dout(n579),.clk(gclk));
	jand g0508(.dina(n579),.dinb(w_n534_0[0]),.dout(n580),.clk(gclk));
	jand g0509(.dina(w_n288_0[1]),.dinb(w_n196_0[2]),.dout(n581),.clk(gclk));
	jand g0510(.dina(w_n355_0[1]),.dinb(w_n246_0[1]),.dout(n582),.clk(gclk));
	jand g0511(.dina(n582),.dinb(w_n170_0[0]),.dout(n583),.clk(gclk));
	jand g0512(.dina(n583),.dinb(n581),.dout(n584),.clk(gclk));
	jor g0513(.dina(n584),.dinb(w_n554_2[1]),.dout(n585),.clk(gclk));
	jor g0514(.dina(n585),.dinb(n580),.dout(n586),.clk(gclk));
	jand g0515(.dina(n586),.dinb(w_G330_0[0]),.dout(n587),.clk(gclk));
	jand g0516(.dina(n587),.dinb(n577),.dout(n588),.clk(gclk));
	jor g0517(.dina(w_n588_1[1]),.dinb(w_n576_1[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(w_n589_1[2]),.dinb(w_n113_1[1]),.dout(n590),.clk(gclk));
	jand g0519(.dina(w_n122_1[0]),.dinb(w_n149_1[1]),.dout(n591),.clk(gclk));
	jnot g0520(.din(w_n591_1[1]),.dout(n592),.clk(gclk));
	jand g0521(.dina(w_n180_0[0]),.dinb(w_n105_1[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(w_n593_0[2]),.dinb(w_G1_1[0]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n592_2[1]),.dout(n595),.clk(gclk));
	jand g0524(.dina(w_n591_1[0]),.dinb(w_n118_0[1]),.dout(n596),.clk(gclk));
	jor g0525(.dina(n596),.dinb(n595),.dout(n597),.clk(gclk));
	jor g0526(.dina(w_dff_B_emsRcblk9_0),.dinb(n590),.dout(w_dff_A_suxkJc9W4_2),.clk(gclk));
	jand g0527(.dina(w_n571_0[1]),.dinb(w_n565_0[0]),.dout(n599),.clk(gclk));
	jnot g0528(.din(n599),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n550_0[0]),.dinb(w_G45_1[0]),.dout(n601),.clk(gclk));
	jor g0530(.dina(n601),.dinb(w_n113_1[0]),.dout(n602),.clk(gclk));
	jnot g0531(.din(w_n602_0[1]),.dout(n603),.clk(gclk));
	jand g0532(.dina(w_n603_2[1]),.dinb(w_n592_2[0]),.dout(n604),.clk(gclk));
	jnot g0533(.din(w_n604_2[1]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_1[2]),.dinb(w_n572_0[1]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(n600),.dout(n607),.clk(gclk));
	jand g0536(.dina(w_n462_0[0]),.dinb(w_n114_0[1]),.dout(n608),.clk(gclk));
	jand g0537(.dina(w_n608_1[2]),.dinb(w_n571_0[0]),.dout(n609),.clk(gclk));
	jnot g0538(.din(n609),.dout(n610),.clk(gclk));
	jand g0539(.dina(w_n146_1[0]),.dinb(w_G20_3[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n115_0[1]),.dout(n612),.clk(gclk));
	jand g0541(.dina(w_G179_0[2]),.dinb(w_G20_3[0]),.dout(n613),.clk(gclk));
	jnot g0542(.din(w_n613_1[1]),.dout(n614),.clk(gclk));
	jand g0543(.dina(w_G200_2[0]),.dinb(w_G20_2[2]),.dout(n615),.clk(gclk));
	jand g0544(.dina(w_n615_0[1]),.dinb(n614),.dout(n616),.clk(gclk));
	jand g0545(.dina(w_n616_0[1]),.dinb(w_G190_2[0]),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n617_6[1]),.dinb(w_G303_2[1]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n407_1[2]),.dinb(w_G20_2[1]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[1]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n615_0[0]),.dinb(w_n613_1[0]),.dout(n621),.clk(gclk));
	jnot g0550(.din(n621),.dout(n622),.clk(gclk));
	jand g0551(.dina(w_n622_0[1]),.dinb(n620),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_n623_5[1]),.dinb(w_G294_3[0]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_G200_1[2]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_n613_0[2]),.dinb(n625),.dout(n626),.clk(gclk));
	jand g0555(.dina(w_n626_0[1]),.dinb(w_G190_1[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(w_n627_7[1]),.dinb(w_G322_0[2]),.dout(n628),.clk(gclk));
	jor g0557(.dina(n628),.dinb(n624),.dout(n629),.clk(gclk));
	jor g0558(.dina(n629),.dinb(n618),.dout(n630),.clk(gclk));
	jand g0559(.dina(w_n622_0[0]),.dinb(w_n619_0[0]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n631_7[1]),.dinb(G329),.dout(n632),.clk(gclk));
	jor g0561(.dina(n632),.dinb(w_n148_5[2]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n616_0[0]),.dinb(w_n407_1[1]),.dout(n634),.clk(gclk));
	jand g0563(.dina(w_n634_4[1]),.dinb(w_G283_3[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_n626_0[0]),.dinb(w_n407_1[0]),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n636_7[1]),.dinb(w_G311_1[2]),.dout(n637),.clk(gclk));
	jor g0566(.dina(n637),.dinb(n635),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n613_0[1]),.dinb(w_G200_1[1]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n639_0[1]),.dinb(w_G190_1[1]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G326_0[1]),.dout(n641),.clk(gclk));
	jand g0570(.dina(w_n639_0[0]),.dinb(w_n407_0[2]),.dout(n642),.clk(gclk));
	jand g0571(.dina(w_n642_7[1]),.dinb(w_G317_1[1]),.dout(n643),.clk(gclk));
	jor g0572(.dina(n643),.dinb(n641),.dout(n644),.clk(gclk));
	jor g0573(.dina(n644),.dinb(n638),.dout(n645),.clk(gclk));
	jor g0574(.dina(n645),.dinb(n633),.dout(n646),.clk(gclk));
	jor g0575(.dina(n646),.dinb(n630),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n631_7[0]),.dinb(w_G159_3[1]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n640_7[0]),.dinb(w_G50_4[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n642_7[0]),.dinb(w_G68_3[2]),.dout(n650),.clk(gclk));
	jor g0579(.dina(n650),.dinb(n649),.dout(n651),.clk(gclk));
	jor g0580(.dina(n651),.dinb(n648),.dout(n652),.clk(gclk));
	jnot g0581(.din(n652),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n617_6[0]),.dinb(w_G87_2[1]),.dout(n654),.clk(gclk));
	jnot g0583(.din(w_n654_0[1]),.dout(n655),.clk(gclk));
	jand g0584(.dina(n655),.dinb(w_n148_5[1]),.dout(n656),.clk(gclk));
	jand g0585(.dina(w_n634_4[0]),.dinb(w_G107_3[1]),.dout(n657),.clk(gclk));
	jand g0586(.dina(w_n636_7[0]),.dinb(w_G77_3[1]),.dout(n658),.clk(gclk));
	jor g0587(.dina(n658),.dinb(w_n657_0[1]),.dout(n659),.clk(gclk));
	jand g0588(.dina(w_n627_7[0]),.dinb(w_G58_3[2]),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n623_5[0]),.dinb(w_G97_3[1]),.dout(n661),.clk(gclk));
	jor g0590(.dina(w_n661_0[1]),.dinb(n660),.dout(n662),.clk(gclk));
	jor g0591(.dina(n662),.dinb(n659),.dout(n663),.clk(gclk));
	jnot g0592(.din(n663),.dout(n664),.clk(gclk));
	jand g0593(.dina(n664),.dinb(n656),.dout(n665),.clk(gclk));
	jand g0594(.dina(n665),.dinb(n653),.dout(n666),.clk(gclk));
	jnot g0595(.din(n666),.dout(n667),.clk(gclk));
	jand g0596(.dina(n667),.dinb(n647),.dout(n668),.clk(gclk));
	jor g0597(.dina(n668),.dinb(w_n612_4[1]),.dout(n669),.clk(gclk));
	jnot g0598(.din(w_n608_1[1]),.dout(n670),.clk(gclk));
	jand g0599(.dina(w_n612_4[0]),.dinb(n670),.dout(n671),.clk(gclk));
	jnot g0600(.din(n671),.dout(n672),.clk(gclk));
	jand g0601(.dina(w_n140_0[0]),.dinb(w_G45_0[2]),.dout(n673),.clk(gclk));
	jand g0602(.dina(w_n118_0[0]),.dinb(w_n161_0[2]),.dout(n674),.clk(gclk));
	jand g0603(.dina(w_n122_0[2]),.dinb(w_G33_6[1]),.dout(n675),.clk(gclk));
	jnot g0604(.din(w_n675_0[2]),.dout(n676),.clk(gclk));
	jor g0605(.dina(w_n676_0[1]),.dinb(n674),.dout(n677),.clk(gclk));
	jor g0606(.dina(n677),.dinb(n673),.dout(n678),.clk(gclk));
	jand g0607(.dina(w_n123_1[1]),.dinb(w_n105_0[2]),.dout(n679),.clk(gclk));
	jand g0608(.dina(w_n122_0[1]),.dinb(w_n148_5[0]),.dout(n680),.clk(gclk));
	jand g0609(.dina(w_n680_0[1]),.dinb(w_G355_0),.dout(n681),.clk(gclk));
	jor g0610(.dina(n681),.dinb(w_dff_B_Y0HyG9oT8_1),.dout(n682),.clk(gclk));
	jnot g0611(.din(n682),.dout(n683),.clk(gclk));
	jand g0612(.dina(n683),.dinb(w_dff_B_9CjI7fM78_1),.dout(n684),.clk(gclk));
	jor g0613(.dina(n684),.dinb(w_n672_1[1]),.dout(n685),.clk(gclk));
	jand g0614(.dina(n685),.dinb(w_n604_2[0]),.dout(n686),.clk(gclk));
	jand g0615(.dina(w_dff_B_Q5u8Ir0H9_0),.dinb(n669),.dout(n687),.clk(gclk));
	jand g0616(.dina(w_dff_B_K7Mb3bCB7_0),.dinb(n610),.dout(n688),.clk(gclk));
	jor g0617(.dina(n688),.dinb(n607),.dout(G396_fa_),.clk(gclk));
	jnot g0618(.din(w_n588_1[0]),.dout(n690),.clk(gclk));
	jnot g0619(.din(w_n401_0[0]),.dout(n691),.clk(gclk));
	jor g0620(.dina(w_n554_2[0]),.dinb(n691),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_n412_0[0]),.dout(n693),.clk(gclk));
	jor g0622(.dina(w_n692_0[0]),.dinb(w_n405_0[0]),.dout(n694),.clk(gclk));
	jnot g0623(.din(n694),.dout(n695),.clk(gclk));
	jor g0624(.dina(n695),.dinb(n693),.dout(n696),.clk(gclk));
	jxor g0625(.dina(w_n696_1[2]),.dinb(w_n576_1[0]),.dout(n697),.clk(gclk));
	jnot g0626(.din(n697),.dout(n698),.clk(gclk));
	jand g0627(.dina(n698),.dinb(n690),.dout(n699),.clk(gclk));
	jor g0628(.dina(w_n991_0[2]),.dinb(w_n604_1[2]),.dout(n701),.clk(gclk));
	jor g0629(.dina(n701),.dinb(n699),.dout(n702),.clk(gclk));
	jnot g0630(.din(w_n696_1[1]),.dout(n703),.clk(gclk));
	jand g0631(.dina(n703),.dinb(w_n425_1[1]),.dout(n704),.clk(gclk));
	jnot g0632(.din(n704),.dout(n705),.clk(gclk));
	jand g0633(.dina(w_n631_6[2]),.dinb(w_G132_1[1]),.dout(n706),.clk(gclk));
	jand g0634(.dina(w_n623_4[2]),.dinb(w_G58_3[1]),.dout(n707),.clk(gclk));
	jand g0635(.dina(w_n642_6[2]),.dinb(w_G150_3[0]),.dout(n708),.clk(gclk));
	jor g0636(.dina(n708),.dinb(n707),.dout(n709),.clk(gclk));
	jor g0637(.dina(n709),.dinb(n706),.dout(n710),.clk(gclk));
	jand g0638(.dina(w_n617_5[2]),.dinb(w_G50_3[2]),.dout(n711),.clk(gclk));
	jor g0639(.dina(n711),.dinb(w_G33_6[0]),.dout(n712),.clk(gclk));
	jand g0640(.dina(w_n636_6[2]),.dinb(w_G159_3[0]),.dout(n713),.clk(gclk));
	jand g0641(.dina(w_n627_6[2]),.dinb(w_G143_2[1]),.dout(n714),.clk(gclk));
	jor g0642(.dina(n714),.dinb(n713),.dout(n715),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G137_1[2]),.dout(n716),.clk(gclk));
	jand g0644(.dina(w_n634_3[2]),.dinb(w_G68_3[1]),.dout(n717),.clk(gclk));
	jor g0645(.dina(w_n717_0[1]),.dinb(n716),.dout(n718),.clk(gclk));
	jor g0646(.dina(n718),.dinb(n715),.dout(n719),.clk(gclk));
	jor g0647(.dina(n719),.dinb(n712),.dout(n720),.clk(gclk));
	jor g0648(.dina(n720),.dinb(n710),.dout(n721),.clk(gclk));
	jand g0649(.dina(w_n631_6[1]),.dinb(w_G311_1[1]),.dout(n722),.clk(gclk));
	jand g0650(.dina(w_n617_5[1]),.dinb(w_G107_3[0]),.dout(n723),.clk(gclk));
	jand g0651(.dina(w_n642_6[1]),.dinb(w_G283_3[0]),.dout(n724),.clk(gclk));
	jor g0652(.dina(n724),.dinb(n723),.dout(n725),.clk(gclk));
	jor g0653(.dina(n725),.dinb(n722),.dout(n726),.clk(gclk));
	jnot g0654(.din(n726),.dout(n727),.clk(gclk));
	jand g0655(.dina(w_n634_3[1]),.dinb(w_G87_2[0]),.dout(n728),.clk(gclk));
	jnot g0656(.din(w_n728_0[1]),.dout(n729),.clk(gclk));
	jand g0657(.dina(n729),.dinb(w_G33_5[2]),.dout(n730),.clk(gclk));
	jand g0658(.dina(w_n636_6[1]),.dinb(w_G116_3[2]),.dout(n731),.clk(gclk));
	jand g0659(.dina(w_n627_6[1]),.dinb(w_G294_2[2]),.dout(n732),.clk(gclk));
	jor g0660(.dina(n732),.dinb(n731),.dout(n733),.clk(gclk));
	jand g0661(.dina(w_n640_6[1]),.dinb(w_G303_2[0]),.dout(n734),.clk(gclk));
	jor g0662(.dina(n734),.dinb(w_n661_0[0]),.dout(n735),.clk(gclk));
	jor g0663(.dina(n735),.dinb(n733),.dout(n736),.clk(gclk));
	jnot g0664(.din(n736),.dout(n737),.clk(gclk));
	jand g0665(.dina(n737),.dinb(n730),.dout(n738),.clk(gclk));
	jand g0666(.dina(n738),.dinb(n727),.dout(n739),.clk(gclk));
	jnot g0667(.din(n739),.dout(n740),.clk(gclk));
	jand g0668(.dina(n740),.dinb(n721),.dout(n741),.clk(gclk));
	jor g0669(.dina(n741),.dinb(w_n612_3[2]),.dout(n742),.clk(gclk));
	jand g0670(.dina(w_n612_3[1]),.dinb(w_n426_0[0]),.dout(n743),.clk(gclk));
	jand g0671(.dina(w_n743_1[1]),.dinb(w_n72_0[1]),.dout(n744),.clk(gclk));
	jor g0672(.dina(n744),.dinb(w_n605_1[1]),.dout(n745),.clk(gclk));
	jnot g0673(.din(n745),.dout(n746),.clk(gclk));
	jand g0674(.dina(n746),.dinb(n742),.dout(n747),.clk(gclk));
	jand g0675(.dina(n747),.dinb(n705),.dout(n748),.clk(gclk));
	jnot g0676(.din(n748),.dout(n749),.clk(gclk));
	jand g0677(.dina(n749),.dinb(n702),.dout(n750),.clk(gclk));
	jnot g0678(.din(w_n750_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0679(.din(w_n552_1[0]),.dout(n752),.clk(gclk));
	jand g0680(.dina(n752),.dinb(w_n542_0[1]),.dout(n753),.clk(gclk));
	jand g0681(.dina(w_n552_0[2]),.dinb(w_n512_0[0]),.dout(n754),.clk(gclk));
	jnot g0682(.din(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0683(.dina(n755),.dinb(w_n517_0[0]),.dout(n756),.clk(gclk));
	jand g0684(.dina(w_n754_0[0]),.dinb(w_n542_0[0]),.dout(n757),.clk(gclk));
	jor g0685(.dina(n757),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0686(.dina(w_n696_1[0]),.dinb(w_n576_0[2]),.dout(n759),.clk(gclk));
	jand g0687(.dina(w_n553_1[2]),.dinb(w_n436_0[0]),.dout(n760),.clk(gclk));
	jnot g0688(.din(w_n760_0[1]),.dout(n761),.clk(gclk));
	jand g0689(.dina(n761),.dinb(w_n446_0[0]),.dout(n762),.clk(gclk));
	jand g0690(.dina(w_n760_0[0]),.dinb(w_n439_0[2]),.dout(n763),.clk(gclk));
	jor g0691(.dina(n763),.dinb(n762),.dout(n764),.clk(gclk));
	jand g0692(.dina(w_n764_1[2]),.dinb(w_n759_0[1]),.dout(n765),.clk(gclk));
	jor g0693(.dina(w_n764_1[1]),.dinb(w_n439_0[1]),.dout(n766),.clk(gclk));
	jand g0694(.dina(w_n554_1[2]),.dinb(w_n543_0[0]),.dout(n767),.clk(gclk));
	jand g0695(.dina(n767),.dinb(n766),.dout(n768),.clk(gclk));
	jor g0696(.dina(n768),.dinb(n765),.dout(n769),.clk(gclk));
	jand g0697(.dina(w_n769_0[1]),.dinb(w_n758_1[1]),.dout(n770),.clk(gclk));
	jor g0698(.dina(n770),.dinb(n753),.dout(n771),.clk(gclk));
	jnot g0699(.din(w_n771_0[2]),.dout(n772),.clk(gclk));
	jand g0700(.dina(w_n576_0[1]),.dinb(w_n519_1[0]),.dout(n773),.clk(gclk));
	jor g0701(.dina(n773),.dinb(w_n548_0[1]),.dout(n774),.clk(gclk));
	jand g0702(.dina(w_n764_1[0]),.dinb(w_n696_0[2]),.dout(n775),.clk(gclk));
	jand g0703(.dina(n775),.dinb(w_n758_1[0]),.dout(n776),.clk(gclk));
	jxor g0704(.dina(n776),.dinb(w_n519_0[2]),.dout(n777),.clk(gclk));
	jand g0705(.dina(n777),.dinb(w_n588_0[2]),.dout(n778),.clk(gclk));
	jxor g0706(.dina(n778),.dinb(n774),.dout(n779),.clk(gclk));
	jnot g0707(.din(w_n779_0[1]),.dout(n780),.clk(gclk));
	jor g0708(.dina(n780),.dinb(n772),.dout(n781),.clk(gclk));
	jor g0709(.dina(w_n779_0[0]),.dinb(w_n771_0[1]),.dout(n782),.clk(gclk));
	jnot g0710(.din(w_n121_0[1]),.dout(n783),.clk(gclk));
	jand g0711(.dina(n783),.dinb(w_n116_0[0]),.dout(n784),.clk(gclk));
	jand g0712(.dina(n784),.dinb(n782),.dout(n785),.clk(gclk));
	jand g0713(.dina(n785),.dinb(n781),.dout(n786),.clk(gclk));
	jand g0714(.dina(w_G77_3[0]),.dinb(w_G50_3[1]),.dout(n787),.clk(gclk));
	jand g0715(.dina(n787),.dinb(w_n137_0[0]),.dout(n788),.clk(gclk));
	jand g0716(.dina(w_G68_3[0]),.dinb(w_n73_1[2]),.dout(n789),.clk(gclk));
	jor g0717(.dina(n789),.dinb(n788),.dout(n790),.clk(gclk));
	jand g0718(.dina(n790),.dinb(w_n121_0[0]),.dout(n791),.clk(gclk));
	jnot g0719(.din(w_n255_0[0]),.dout(n792),.clk(gclk));
	jand g0720(.dina(w_n147_0[0]),.dinb(w_G116_3[1]),.dout(n793),.clk(gclk));
	jand g0721(.dina(n793),.dinb(n792),.dout(n794),.clk(gclk));
	jor g0722(.dina(n794),.dinb(n791),.dout(n795),.clk(gclk));
	jor g0723(.dina(w_dff_B_gaRAddgQ5_0),.dinb(n786),.dout(w_dff_A_8Faaqfu06_2),.clk(gclk));
	jand g0724(.dina(w_n553_1[1]),.dinb(w_n214_0[0]),.dout(n797),.clk(gclk));
	jnot g0725(.din(w_n797_0[1]),.dout(n798),.clk(gclk));
	jand g0726(.dina(n798),.dinb(w_n219_0[0]),.dout(n799),.clk(gclk));
	jand g0727(.dina(w_n797_0[0]),.dinb(w_n532_0[0]),.dout(n800),.clk(gclk));
	jor g0728(.dina(n800),.dinb(n799),.dout(n801),.clk(gclk));
	jnot g0729(.din(w_n801_0[1]),.dout(n802),.clk(gclk));
	jand g0730(.dina(n802),.dinb(w_n608_1[0]),.dout(n803),.clk(gclk));
	jnot g0731(.din(n803),.dout(n804),.clk(gclk));
	jand g0732(.dina(w_n631_6[0]),.dinb(w_G317_1[0]),.dout(n805),.clk(gclk));
	jand g0733(.dina(w_n623_4[1]),.dinb(w_G107_2[2]),.dout(n806),.clk(gclk));
	jand g0734(.dina(w_n642_6[0]),.dinb(w_G294_2[1]),.dout(n807),.clk(gclk));
	jor g0735(.dina(n807),.dinb(n806),.dout(n808),.clk(gclk));
	jor g0736(.dina(n808),.dinb(n805),.dout(n809),.clk(gclk));
	jand g0737(.dina(w_n617_5[0]),.dinb(w_G116_3[0]),.dout(n810),.clk(gclk));
	jor g0738(.dina(n810),.dinb(w_n148_4[2]),.dout(n811),.clk(gclk));
	jand g0739(.dina(w_n636_6[0]),.dinb(w_G283_2[2]),.dout(n812),.clk(gclk));
	jand g0740(.dina(w_n627_6[0]),.dinb(w_G303_1[2]),.dout(n813),.clk(gclk));
	jor g0741(.dina(n813),.dinb(n812),.dout(n814),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G311_1[0]),.dout(n815),.clk(gclk));
	jand g0743(.dina(w_n634_3[0]),.dinb(w_G97_3[0]),.dout(n816),.clk(gclk));
	jor g0744(.dina(w_n816_0[1]),.dinb(n815),.dout(n817),.clk(gclk));
	jor g0745(.dina(n817),.dinb(n814),.dout(n818),.clk(gclk));
	jor g0746(.dina(n818),.dinb(n811),.dout(n819),.clk(gclk));
	jor g0747(.dina(n819),.dinb(n809),.dout(n820),.clk(gclk));
	jand g0748(.dina(w_n631_5[2]),.dinb(w_G137_1[1]),.dout(n821),.clk(gclk));
	jnot g0749(.din(n821),.dout(n822),.clk(gclk));
	jand g0750(.dina(w_n623_4[0]),.dinb(w_G68_2[2]),.dout(n823),.clk(gclk));
	jnot g0751(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jand g0752(.dina(w_n634_2[2]),.dinb(w_G77_2[2]),.dout(n825),.clk(gclk));
	jnot g0753(.din(w_n825_0[1]),.dout(n826),.clk(gclk));
	jand g0754(.dina(n826),.dinb(n824),.dout(n827),.clk(gclk));
	jand g0755(.dina(n827),.dinb(n822),.dout(n828),.clk(gclk));
	jand g0756(.dina(w_n642_5[2]),.dinb(w_G159_2[2]),.dout(n829),.clk(gclk));
	jor g0757(.dina(n829),.dinb(w_G33_5[1]),.dout(n830),.clk(gclk));
	jand g0758(.dina(w_n640_5[2]),.dinb(w_G143_2[0]),.dout(n831),.clk(gclk));
	jand g0759(.dina(w_n627_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jor g0760(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jand g0761(.dina(w_n636_5[2]),.dinb(w_G50_3[0]),.dout(n834),.clk(gclk));
	jand g0762(.dina(w_n617_4[2]),.dinb(w_G58_3[0]),.dout(n835),.clk(gclk));
	jor g0763(.dina(n835),.dinb(n834),.dout(n836),.clk(gclk));
	jor g0764(.dina(n836),.dinb(n833),.dout(n837),.clk(gclk));
	jor g0765(.dina(n837),.dinb(n830),.dout(n838),.clk(gclk));
	jnot g0766(.din(n838),.dout(n839),.clk(gclk));
	jand g0767(.dina(n839),.dinb(n828),.dout(n840),.clk(gclk));
	jnot g0768(.din(n840),.dout(n841),.clk(gclk));
	jand g0769(.dina(n841),.dinb(n820),.dout(n842),.clk(gclk));
	jor g0770(.dina(n842),.dinb(w_n612_3[0]),.dout(n843),.clk(gclk));
	jand g0771(.dina(w_n675_0[1]),.dinb(w_n131_0[0]),.dout(n844),.clk(gclk));
	jand g0772(.dina(w_n123_1[0]),.dinb(w_G87_1[2]),.dout(n845),.clk(gclk));
	jor g0773(.dina(n845),.dinb(w_n672_1[0]),.dout(n846),.clk(gclk));
	jor g0774(.dina(n846),.dinb(n844),.dout(n847),.clk(gclk));
	jand g0775(.dina(n847),.dinb(w_n604_1[1]),.dout(n848),.clk(gclk));
	jand g0776(.dina(n848),.dinb(n843),.dout(n849),.clk(gclk));
	jand g0777(.dina(n849),.dinb(n804),.dout(n850),.clk(gclk));
	jnot g0778(.din(w_n589_1[1]),.dout(n851),.clk(gclk));
	jxor g0779(.dina(w_n561_0[0]),.dinb(w_n556_0[0]),.dout(n852),.clk(gclk));
	jxor g0780(.dina(n852),.dinb(w_n572_0[0]),.dout(n853),.clk(gclk));
	jnot g0781(.din(w_n853_0[2]),.dout(n854),.clk(gclk));
	jand g0782(.dina(n854),.dinb(n851),.dout(n855),.clk(gclk));
	jnot g0783(.din(w_n278_0[0]),.dout(n856),.clk(gclk));
	jand g0784(.dina(w_n553_1[0]),.dinb(w_n274_0[0]),.dout(n857),.clk(gclk));
	jor g0785(.dina(n857),.dinb(n856),.dout(n858),.clk(gclk));
	jand g0786(.dina(w_n553_0[2]),.dinb(w_n536_0[1]),.dout(n859),.clk(gclk));
	jnot g0787(.din(n859),.dout(n860),.clk(gclk));
	jand g0788(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jxor g0789(.dina(w_n861_1[1]),.dinb(w_n573_0[1]),.dout(n862),.clk(gclk));
	jxor g0790(.dina(n862),.dinb(w_n563_0[1]),.dout(n863),.clk(gclk));
	jand g0791(.dina(w_n863_0[1]),.dinb(w_n855_0[2]),.dout(n864),.clk(gclk));
	jor g0792(.dina(w_n864_0[1]),.dinb(w_n589_1[0]),.dout(n865),.clk(gclk));
	jand g0793(.dina(n865),.dinb(w_n591_0[2]),.dout(n866),.clk(gclk));
	jor g0794(.dina(n866),.dinb(w_n602_0[0]),.dout(n867),.clk(gclk));
	jand g0795(.dina(w_n554_1[1]),.dinb(w_n536_0[0]),.dout(n868),.clk(gclk));
	jnot g0796(.din(w_n861_1[0]),.dout(n869),.clk(gclk));
	jand g0797(.dina(n869),.dinb(w_n563_0[0]),.dout(n870),.clk(gclk));
	jor g0798(.dina(n870),.dinb(n868),.dout(n871),.clk(gclk));
	jor g0799(.dina(w_n861_0[2]),.dinb(w_n573_0[0]),.dout(n872),.clk(gclk));
	jxor g0800(.dina(n872),.dinb(w_n801_0[0]),.dout(n873),.clk(gclk));
	jxor g0801(.dina(n873),.dinb(n871),.dout(n874),.clk(gclk));
	jnot g0802(.din(n874),.dout(n875),.clk(gclk));
	jand g0803(.dina(n875),.dinb(n867),.dout(n876),.clk(gclk));
	jor g0804(.dina(n876),.dinb(n850),.dout(G387_fa_),.clk(gclk));
	jand g0805(.dina(w_n853_0[1]),.dinb(w_n589_0[2]),.dout(n878),.clk(gclk));
	jor g0806(.dina(w_n855_0[1]),.dinb(w_n592_1[2]),.dout(n879),.clk(gclk));
	jor g0807(.dina(n879),.dinb(n878),.dout(n880),.clk(gclk));
	jor g0808(.dina(w_n853_0[0]),.dinb(w_n603_2[0]),.dout(n881),.clk(gclk));
	jand g0809(.dina(w_n608_0[2]),.dinb(w_n564_0[0]),.dout(n882),.clk(gclk));
	jand g0810(.dina(w_n631_5[1]),.dinb(w_G326_0[0]),.dout(n883),.clk(gclk));
	jand g0811(.dina(w_n623_3[2]),.dinb(w_G283_2[1]),.dout(n884),.clk(gclk));
	jand g0812(.dina(w_n627_5[1]),.dinb(w_G317_0[2]),.dout(n885),.clk(gclk));
	jor g0813(.dina(n885),.dinb(n884),.dout(n886),.clk(gclk));
	jor g0814(.dina(n886),.dinb(n883),.dout(n887),.clk(gclk));
	jand g0815(.dina(w_n617_4[1]),.dinb(w_G294_2[0]),.dout(n888),.clk(gclk));
	jor g0816(.dina(n888),.dinb(w_n148_4[1]),.dout(n889),.clk(gclk));
	jand g0817(.dina(w_n634_2[1]),.dinb(w_G116_2[2]),.dout(n890),.clk(gclk));
	jand g0818(.dina(w_n636_5[1]),.dinb(w_G303_1[1]),.dout(n891),.clk(gclk));
	jor g0819(.dina(n891),.dinb(n890),.dout(n892),.clk(gclk));
	jand g0820(.dina(w_n640_5[1]),.dinb(w_G322_0[1]),.dout(n893),.clk(gclk));
	jand g0821(.dina(w_n642_5[1]),.dinb(w_G311_0[2]),.dout(n894),.clk(gclk));
	jor g0822(.dina(n894),.dinb(n893),.dout(n895),.clk(gclk));
	jor g0823(.dina(n895),.dinb(n892),.dout(n896),.clk(gclk));
	jor g0824(.dina(n896),.dinb(n889),.dout(n897),.clk(gclk));
	jor g0825(.dina(n897),.dinb(n887),.dout(n898),.clk(gclk));
	jand g0826(.dina(w_n623_3[1]),.dinb(w_G87_1[1]),.dout(n899),.clk(gclk));
	jand g0827(.dina(w_n642_5[0]),.dinb(w_G58_2[2]),.dout(n900),.clk(gclk));
	jor g0828(.dina(n900),.dinb(w_n816_0[0]),.dout(n901),.clk(gclk));
	jor g0829(.dina(n901),.dinb(w_n899_0[1]),.dout(n902),.clk(gclk));
	jand g0830(.dina(w_n631_5[0]),.dinb(w_G150_2[1]),.dout(n903),.clk(gclk));
	jor g0831(.dina(n903),.dinb(w_G33_5[0]),.dout(n904),.clk(gclk));
	jand g0832(.dina(w_n640_5[0]),.dinb(w_G159_2[1]),.dout(n905),.clk(gclk));
	jand g0833(.dina(w_n636_5[0]),.dinb(w_G68_2[1]),.dout(n906),.clk(gclk));
	jor g0834(.dina(n906),.dinb(n905),.dout(n907),.clk(gclk));
	jand g0835(.dina(w_n627_5[0]),.dinb(w_G50_2[2]),.dout(n908),.clk(gclk));
	jand g0836(.dina(w_n617_4[0]),.dinb(w_G77_2[1]),.dout(n909),.clk(gclk));
	jor g0837(.dina(w_n909_0[1]),.dinb(n908),.dout(n910),.clk(gclk));
	jor g0838(.dina(n910),.dinb(n907),.dout(n911),.clk(gclk));
	jor g0839(.dina(n911),.dinb(n904),.dout(n912),.clk(gclk));
	jor g0840(.dina(n912),.dinb(n902),.dout(n913),.clk(gclk));
	jand g0841(.dina(n913),.dinb(n898),.dout(n914),.clk(gclk));
	jor g0842(.dina(n914),.dinb(w_n612_2[2]),.dout(n915),.clk(gclk));
	jand g0843(.dina(w_n135_0[0]),.dinb(w_G45_0[1]),.dout(n916),.clk(gclk));
	jand g0844(.dina(w_G77_2[0]),.dinb(w_G68_2[0]),.dout(n917),.clk(gclk));
	jnot g0845(.din(n917),.dout(n918),.clk(gclk));
	jand g0846(.dina(w_G58_2[1]),.dinb(w_n161_0[1]),.dout(n919),.clk(gclk));
	jand g0847(.dina(n919),.dinb(w_n73_1[1]),.dout(n920),.clk(gclk));
	jand g0848(.dina(n920),.dinb(n918),.dout(n921),.clk(gclk));
	jand g0849(.dina(n921),.dinb(w_n593_0[1]),.dout(n922),.clk(gclk));
	jor g0850(.dina(n922),.dinb(w_n676_0[0]),.dout(n923),.clk(gclk));
	jor g0851(.dina(n923),.dinb(n916),.dout(n924),.clk(gclk));
	jand g0852(.dina(w_n123_0[2]),.dinb(w_n80_0[1]),.dout(n925),.clk(gclk));
	jnot g0853(.din(w_n593_0[0]),.dout(n926),.clk(gclk));
	jand g0854(.dina(w_n680_0[0]),.dinb(n926),.dout(n927),.clk(gclk));
	jor g0855(.dina(n927),.dinb(n925),.dout(n928),.clk(gclk));
	jnot g0856(.din(n928),.dout(n929),.clk(gclk));
	jand g0857(.dina(n929),.dinb(n924),.dout(n930),.clk(gclk));
	jor g0858(.dina(n930),.dinb(w_n672_0[2]),.dout(n931),.clk(gclk));
	jand g0859(.dina(n931),.dinb(w_n604_1[0]),.dout(n932),.clk(gclk));
	jand g0860(.dina(n932),.dinb(n915),.dout(n933),.clk(gclk));
	jnot g0861(.din(n933),.dout(n934),.clk(gclk));
	jor g0862(.dina(n934),.dinb(n882),.dout(n935),.clk(gclk));
	jand g0863(.dina(n935),.dinb(n881),.dout(n936),.clk(gclk));
	jand g0864(.dina(n936),.dinb(n880),.dout(n937),.clk(gclk));
	jnot g0865(.din(w_n937_0[2]),.dout(w_dff_A_QIL9dh5f4_1),.clk(gclk));
	jnot g0866(.din(w_n855_0[0]),.dout(n939),.clk(gclk));
	jnot g0867(.din(w_n863_0[0]),.dout(n940),.clk(gclk));
	jand g0868(.dina(w_n940_0[1]),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0869(.dina(w_n864_0[0]),.dinb(w_n592_1[1]),.dout(n942),.clk(gclk));
	jor g0870(.dina(n942),.dinb(n941),.dout(n943),.clk(gclk));
	jor g0871(.dina(w_n940_0[0]),.dinb(w_n603_1[2]),.dout(n944),.clk(gclk));
	jand g0872(.dina(w_n861_0[1]),.dinb(w_n608_0[1]),.dout(n945),.clk(gclk));
	jnot g0873(.din(n945),.dout(n946),.clk(gclk));
	jand g0874(.dina(w_n623_3[0]),.dinb(w_G116_2[1]),.dout(n947),.clk(gclk));
	jand g0875(.dina(w_n617_3[2]),.dinb(w_G283_2[0]),.dout(n948),.clk(gclk));
	jand g0876(.dina(w_n642_4[2]),.dinb(w_G303_1[0]),.dout(n949),.clk(gclk));
	jor g0877(.dina(n949),.dinb(n948),.dout(n950),.clk(gclk));
	jor g0878(.dina(n950),.dinb(n947),.dout(n951),.clk(gclk));
	jand g0879(.dina(w_n631_4[2]),.dinb(w_G322_0[0]),.dout(n952),.clk(gclk));
	jor g0880(.dina(n952),.dinb(w_n148_4[0]),.dout(n953),.clk(gclk));
	jand g0881(.dina(w_n636_4[2]),.dinb(w_G294_1[2]),.dout(n954),.clk(gclk));
	jand g0882(.dina(w_n627_4[2]),.dinb(w_G311_0[1]),.dout(n955),.clk(gclk));
	jor g0883(.dina(n955),.dinb(n954),.dout(n956),.clk(gclk));
	jand g0884(.dina(w_n640_4[2]),.dinb(w_G317_0[1]),.dout(n957),.clk(gclk));
	jor g0885(.dina(n957),.dinb(w_n657_0[0]),.dout(n958),.clk(gclk));
	jor g0886(.dina(n958),.dinb(n956),.dout(n959),.clk(gclk));
	jor g0887(.dina(n959),.dinb(n953),.dout(n960),.clk(gclk));
	jor g0888(.dina(n960),.dinb(n951),.dout(n961),.clk(gclk));
	jand g0889(.dina(w_n623_2[2]),.dinb(w_G77_1[2]),.dout(n962),.clk(gclk));
	jand g0890(.dina(w_n617_3[1]),.dinb(w_G68_1[2]),.dout(n963),.clk(gclk));
	jand g0891(.dina(w_n642_4[1]),.dinb(w_G50_2[1]),.dout(n964),.clk(gclk));
	jor g0892(.dina(n964),.dinb(n963),.dout(n965),.clk(gclk));
	jor g0893(.dina(n965),.dinb(w_n962_0[1]),.dout(n966),.clk(gclk));
	jand g0894(.dina(w_n631_4[1]),.dinb(w_G143_1[2]),.dout(n967),.clk(gclk));
	jor g0895(.dina(n967),.dinb(w_G33_4[2]),.dout(n968),.clk(gclk));
	jand g0896(.dina(w_n636_4[1]),.dinb(w_G58_2[0]),.dout(n969),.clk(gclk));
	jand g0897(.dina(w_n627_4[1]),.dinb(w_G159_2[0]),.dout(n970),.clk(gclk));
	jor g0898(.dina(n970),.dinb(n969),.dout(n971),.clk(gclk));
	jand g0899(.dina(w_n640_4[1]),.dinb(w_G150_2[0]),.dout(n972),.clk(gclk));
	jor g0900(.dina(n972),.dinb(w_n728_0[0]),.dout(n973),.clk(gclk));
	jor g0901(.dina(n973),.dinb(n971),.dout(n974),.clk(gclk));
	jor g0902(.dina(n974),.dinb(n968),.dout(n975),.clk(gclk));
	jor g0903(.dina(n975),.dinb(n966),.dout(n976),.clk(gclk));
	jand g0904(.dina(n976),.dinb(n961),.dout(n977),.clk(gclk));
	jor g0905(.dina(n977),.dinb(w_n612_2[1]),.dout(n978),.clk(gclk));
	jand g0906(.dina(w_n675_0[0]),.dinb(w_n144_0[0]),.dout(n979),.clk(gclk));
	jand g0907(.dina(w_n123_0[1]),.dinb(w_G97_2[2]),.dout(n980),.clk(gclk));
	jor g0908(.dina(n980),.dinb(w_n672_0[1]),.dout(n981),.clk(gclk));
	jor g0909(.dina(n981),.dinb(n979),.dout(n982),.clk(gclk));
	jand g0910(.dina(n982),.dinb(w_n604_0[2]),.dout(n983),.clk(gclk));
	jand g0911(.dina(n983),.dinb(n978),.dout(n984),.clk(gclk));
	jand g0912(.dina(n984),.dinb(n946),.dout(n985),.clk(gclk));
	jnot g0913(.din(n985),.dout(n986),.clk(gclk));
	jand g0914(.dina(n986),.dinb(n944),.dout(n987),.clk(gclk));
	jand g0915(.dina(n987),.dinb(n943),.dout(n988),.clk(gclk));
	jnot g0916(.din(w_n988_0[2]),.dout(w_dff_A_C8WizjaC4_1),.clk(gclk));
	jnot g0917(.din(w_n758_0[2]),.dout(n990),.clk(gclk));
	jand g0918(.dina(w_n696_0[1]),.dinb(w_n588_0[1]),.dout(n991),.clk(gclk));
	jand g0919(.dina(w_n991_0[1]),.dinb(w_n764_0[2]),.dout(n992),.clk(gclk));
	jxor g0920(.dina(w_n992_0[1]),.dinb(w_n990_0[1]),.dout(n993),.clk(gclk));
	jxor g0921(.dina(n993),.dinb(w_n769_0[0]),.dout(n994),.clk(gclk));
	jand g0922(.dina(w_n589_0[1]),.dinb(w_n519_0[1]),.dout(n995),.clk(gclk));
	jor g0923(.dina(n995),.dinb(w_n548_0[0]),.dout(n996),.clk(gclk));
	jand g0924(.dina(w_n554_1[0]),.dinb(w_n404_0[0]),.dout(n997),.clk(gclk));
	jor g0925(.dina(n997),.dinb(w_n759_0[0]),.dout(n998),.clk(gclk));
	jnot g0926(.din(w_n764_0[1]),.dout(n999),.clk(gclk));
	jxor g0927(.dina(w_n991_0[0]),.dinb(w_n999_0[1]),.dout(n1000),.clk(gclk));
	jxor g0928(.dina(n1000),.dinb(n998),.dout(n1001),.clk(gclk));
	jor g0929(.dina(w_n1001_0[2]),.dinb(w_n996_0[2]),.dout(n1002),.clk(gclk));
	jor g0930(.dina(w_n1002_0[2]),.dinb(w_n994_0[2]),.dout(n1003),.clk(gclk));
	jnot g0931(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0932(.dina(w_n1002_0[1]),.dinb(w_n994_0[1]),.dout(n1005),.clk(gclk));
	jor g0933(.dina(n1005),.dinb(w_n592_1[0]),.dout(n1006),.clk(gclk));
	jor g0934(.dina(n1006),.dinb(n1004),.dout(n1007),.clk(gclk));
	jor g0935(.dina(w_n994_0[0]),.dinb(w_n603_1[1]),.dout(n1008),.clk(gclk));
	jand g0936(.dina(w_n990_0[0]),.dinb(w_n425_1[0]),.dout(n1009),.clk(gclk));
	jnot g0937(.din(n1009),.dout(n1010),.clk(gclk));
	jand g0938(.dina(w_n631_4[0]),.dinb(w_G125_0[1]),.dout(n1011),.clk(gclk));
	jand g0939(.dina(w_n623_2[1]),.dinb(w_G159_1[2]),.dout(n1012),.clk(gclk));
	jand g0940(.dina(w_n642_4[0]),.dinb(w_G137_1[0]),.dout(n1013),.clk(gclk));
	jor g0941(.dina(n1013),.dinb(n1012),.dout(n1014),.clk(gclk));
	jor g0942(.dina(n1014),.dinb(n1011),.dout(n1015),.clk(gclk));
	jand g0943(.dina(w_n617_3[0]),.dinb(w_G150_1[2]),.dout(n1016),.clk(gclk));
	jor g0944(.dina(n1016),.dinb(w_G33_4[1]),.dout(n1017),.clk(gclk));
	jand g0945(.dina(w_n636_4[0]),.dinb(w_G143_1[1]),.dout(n1018),.clk(gclk));
	jand g0946(.dina(w_n627_4[0]),.dinb(w_G132_1[0]),.dout(n1019),.clk(gclk));
	jor g0947(.dina(n1019),.dinb(n1018),.dout(n1020),.clk(gclk));
	jand g0948(.dina(w_n640_4[0]),.dinb(w_G128_0[2]),.dout(n1021),.clk(gclk));
	jand g0949(.dina(w_n634_2[0]),.dinb(w_G50_2[0]),.dout(n1022),.clk(gclk));
	jor g0950(.dina(n1022),.dinb(n1021),.dout(n1023),.clk(gclk));
	jor g0951(.dina(n1023),.dinb(n1020),.dout(n1024),.clk(gclk));
	jor g0952(.dina(n1024),.dinb(n1017),.dout(n1025),.clk(gclk));
	jor g0953(.dina(n1025),.dinb(n1015),.dout(n1026),.clk(gclk));
	jand g0954(.dina(w_n631_3[2]),.dinb(w_G294_1[1]),.dout(n1027),.clk(gclk));
	jand g0955(.dina(w_n642_3[2]),.dinb(w_G107_2[1]),.dout(n1028),.clk(gclk));
	jor g0956(.dina(n1028),.dinb(w_n962_0[0]),.dout(n1029),.clk(gclk));
	jor g0957(.dina(n1029),.dinb(n1027),.dout(n1030),.clk(gclk));
	jand g0958(.dina(w_n640_3[2]),.dinb(w_G283_1[2]),.dout(n1031),.clk(gclk));
	jor g0959(.dina(n1031),.dinb(w_n148_3[2]),.dout(n1032),.clk(gclk));
	jand g0960(.dina(w_n636_3[2]),.dinb(w_G97_2[1]),.dout(n1033),.clk(gclk));
	jand g0961(.dina(w_n627_3[2]),.dinb(w_G116_2[0]),.dout(n1034),.clk(gclk));
	jor g0962(.dina(n1034),.dinb(n1033),.dout(n1035),.clk(gclk));
	jor g0963(.dina(w_n717_0[0]),.dinb(w_n654_0[0]),.dout(n1036),.clk(gclk));
	jor g0964(.dina(n1036),.dinb(n1035),.dout(n1037),.clk(gclk));
	jor g0965(.dina(n1037),.dinb(n1032),.dout(n1038),.clk(gclk));
	jor g0966(.dina(n1038),.dinb(n1030),.dout(n1039),.clk(gclk));
	jand g0967(.dina(n1039),.dinb(n1026),.dout(n1040),.clk(gclk));
	jor g0968(.dina(n1040),.dinb(w_n612_2[0]),.dout(n1041),.clk(gclk));
	jand g0969(.dina(w_n743_1[0]),.dinb(w_n74_0[1]),.dout(n1042),.clk(gclk));
	jor g0970(.dina(n1042),.dinb(w_n605_1[0]),.dout(n1043),.clk(gclk));
	jnot g0971(.din(n1043),.dout(n1044),.clk(gclk));
	jand g0972(.dina(n1044),.dinb(n1041),.dout(n1045),.clk(gclk));
	jand g0973(.dina(n1045),.dinb(n1010),.dout(n1046),.clk(gclk));
	jnot g0974(.din(n1046),.dout(n1047),.clk(gclk));
	jand g0975(.dina(n1047),.dinb(n1008),.dout(n1048),.clk(gclk));
	jand g0976(.dina(n1048),.dinb(n1007),.dout(n1049),.clk(gclk));
	jnot g0977(.din(w_n1049_0[2]),.dout(w_dff_A_4BLq7DIM7_1),.clk(gclk));
	jand g0978(.dina(w_n992_0[0]),.dinb(w_n758_0[1]),.dout(n1051),.clk(gclk));
	jand g0979(.dina(w_n552_0[1]),.dinb(w_n479_0[0]),.dout(n1052),.clk(gclk));
	jnot g0980(.din(w_n1052_0[1]),.dout(n1053),.clk(gclk));
	jand g0981(.dina(n1053),.dinb(w_n484_0[0]),.dout(n1054),.clk(gclk));
	jand g0982(.dina(w_n1052_0[0]),.dinb(w_n541_0[0]),.dout(n1055),.clk(gclk));
	jor g0983(.dina(n1055),.dinb(n1054),.dout(n1056),.clk(gclk));
	jnot g0984(.din(n1056),.dout(n1057),.clk(gclk));
	jxor g0985(.dina(w_n1057_0[1]),.dinb(w_n771_0[0]),.dout(n1058),.clk(gclk));
	jxor g0986(.dina(n1058),.dinb(n1051),.dout(n1059),.clk(gclk));
	jor g0987(.dina(w_n1059_0[1]),.dinb(w_n603_1[0]),.dout(n1060),.clk(gclk));
	jnot g0988(.din(w_n996_0[1]),.dout(n1061),.clk(gclk));
	jand g0989(.dina(w_n1003_0[0]),.dinb(n1061),.dout(n1062),.clk(gclk));
	jor g0990(.dina(n1062),.dinb(w_n592_0[2]),.dout(n1063),.clk(gclk));
	jor g0991(.dina(n1063),.dinb(w_n1059_0[0]),.dout(n1064),.clk(gclk));
	jand g0992(.dina(w_n1057_0[0]),.dinb(w_n425_0[2]),.dout(n1065),.clk(gclk));
	jnot g0993(.din(w_n612_1[2]),.dout(n1066),.clk(gclk));
	jand g0994(.dina(w_n642_3[1]),.dinb(w_G132_0[2]),.dout(n1067),.clk(gclk));
	jand g0995(.dina(w_n627_3[1]),.dinb(w_G128_0[1]),.dout(n1068),.clk(gclk));
	jand g0996(.dina(w_n636_3[1]),.dinb(w_G137_0[2]),.dout(n1069),.clk(gclk));
	jor g0997(.dina(n1069),.dinb(n1068),.dout(n1070),.clk(gclk));
	jor g0998(.dina(n1070),.dinb(n1067),.dout(n1071),.clk(gclk));
	jnot g0999(.din(n1071),.dout(n1072),.clk(gclk));
	jand g1000(.dina(w_n623_2[0]),.dinb(w_G150_1[1]),.dout(n1073),.clk(gclk));
	jnot g1001(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1002(.dina(w_n149_1[0]),.dinb(w_n148_3[1]),.dout(n1075),.clk(gclk));
	jand g1003(.dina(n1075),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_G125_0[0]),.dout(n1077),.clk(gclk));
	jand g1005(.dina(w_n617_2[2]),.dinb(w_G143_1[0]),.dout(n1078),.clk(gclk));
	jor g1006(.dina(n1078),.dinb(n1077),.dout(n1079),.clk(gclk));
	jand g1007(.dina(w_n631_3[1]),.dinb(G124),.dout(n1080),.clk(gclk));
	jand g1008(.dina(w_n634_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jor g1009(.dina(n1081),.dinb(n1080),.dout(n1082),.clk(gclk));
	jor g1010(.dina(n1082),.dinb(n1079),.dout(n1083),.clk(gclk));
	jnot g1011(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1012(.dina(n1084),.dinb(n1076),.dout(n1085),.clk(gclk));
	jand g1013(.dina(n1085),.dinb(n1072),.dout(n1086),.clk(gclk));
	jand g1014(.dina(w_n627_3[0]),.dinb(w_G107_2[0]),.dout(n1087),.clk(gclk));
	jand g1015(.dina(w_n634_1[1]),.dinb(w_G58_1[2]),.dout(n1088),.clk(gclk));
	jand g1016(.dina(w_n636_3[0]),.dinb(w_G87_1[0]),.dout(n1089),.clk(gclk));
	jor g1017(.dina(n1089),.dinb(w_n1088_0[1]),.dout(n1090),.clk(gclk));
	jor g1018(.dina(n1090),.dinb(n1087),.dout(n1091),.clk(gclk));
	jnot g1019(.din(n1091),.dout(n1092),.clk(gclk));
	jand g1020(.dina(w_n642_3[0]),.dinb(w_G97_2[0]),.dout(n1093),.clk(gclk));
	jnot g1021(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1022(.dina(w_n149_0[2]),.dinb(w_G33_4[0]),.dout(n1095),.clk(gclk));
	jand g1023(.dina(n1095),.dinb(n1094),.dout(n1096),.clk(gclk));
	jand g1024(.dina(w_n631_3[0]),.dinb(w_G283_1[1]),.dout(n1097),.clk(gclk));
	jor g1025(.dina(n1097),.dinb(w_n823_0[0]),.dout(n1098),.clk(gclk));
	jand g1026(.dina(w_n640_3[0]),.dinb(w_G116_1[2]),.dout(n1099),.clk(gclk));
	jor g1027(.dina(n1099),.dinb(w_n909_0[0]),.dout(n1100),.clk(gclk));
	jor g1028(.dina(n1100),.dinb(n1098),.dout(n1101),.clk(gclk));
	jnot g1029(.din(n1101),.dout(n1102),.clk(gclk));
	jand g1030(.dina(n1102),.dinb(n1096),.dout(n1103),.clk(gclk));
	jand g1031(.dina(n1103),.dinb(n1092),.dout(n1104),.clk(gclk));
	jand g1032(.dina(w_n73_1[0]),.dinb(w_G41_0[1]),.dout(n1105),.clk(gclk));
	jor g1033(.dina(n1105),.dinb(n1104),.dout(n1106),.clk(gclk));
	jor g1034(.dina(n1106),.dinb(n1086),.dout(n1107),.clk(gclk));
	jand g1035(.dina(n1107),.dinb(n1066),.dout(n1108),.clk(gclk));
	jand g1036(.dina(w_n743_0[2]),.dinb(w_n73_0[2]),.dout(n1109),.clk(gclk));
	jor g1037(.dina(n1109),.dinb(w_n605_0[2]),.dout(n1110),.clk(gclk));
	jor g1038(.dina(n1110),.dinb(n1108),.dout(n1111),.clk(gclk));
	jor g1039(.dina(n1111),.dinb(n1065),.dout(n1112),.clk(gclk));
	jand g1040(.dina(n1112),.dinb(n1064),.dout(n1113),.clk(gclk));
	jand g1041(.dina(n1113),.dinb(n1060),.dout(n1114),.clk(gclk));
	jnot g1042(.din(w_n1114_0[2]),.dout(w_dff_A_Kdmz1GUI9_1),.clk(gclk));
	jand g1043(.dina(w_n1001_0[1]),.dinb(w_n996_0[0]),.dout(n1116),.clk(gclk));
	jnot g1044(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1045(.dina(w_n1002_0[0]),.dinb(w_n591_0[1]),.dout(n1118),.clk(gclk));
	jand g1046(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jnot g1047(.din(n1119),.dout(n1120),.clk(gclk));
	jor g1048(.dina(w_n1001_0[0]),.dinb(w_n603_0[2]),.dout(n1121),.clk(gclk));
	jand g1049(.dina(w_n999_0[0]),.dinb(w_n425_0[1]),.dout(n1122),.clk(gclk));
	jnot g1050(.din(n1122),.dout(n1123),.clk(gclk));
	jand g1051(.dina(w_n623_1[2]),.dinb(w_G50_1[2]),.dout(n1124),.clk(gclk));
	jand g1052(.dina(w_n617_2[1]),.dinb(w_G159_1[0]),.dout(n1125),.clk(gclk));
	jand g1053(.dina(w_n642_2[2]),.dinb(w_G143_0[2]),.dout(n1126),.clk(gclk));
	jor g1054(.dina(n1126),.dinb(n1125),.dout(n1127),.clk(gclk));
	jor g1055(.dina(n1127),.dinb(n1124),.dout(n1128),.clk(gclk));
	jand g1056(.dina(w_n631_2[2]),.dinb(w_G128_0[0]),.dout(n1129),.clk(gclk));
	jor g1057(.dina(n1129),.dinb(w_G33_3[2]),.dout(n1130),.clk(gclk));
	jand g1058(.dina(w_n636_2[2]),.dinb(w_G150_1[0]),.dout(n1131),.clk(gclk));
	jand g1059(.dina(w_n627_2[2]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jor g1060(.dina(n1132),.dinb(n1131),.dout(n1133),.clk(gclk));
	jand g1061(.dina(w_n640_2[2]),.dinb(w_G132_0[1]),.dout(n1134),.clk(gclk));
	jor g1062(.dina(n1134),.dinb(w_n1088_0[0]),.dout(n1135),.clk(gclk));
	jor g1063(.dina(n1135),.dinb(n1133),.dout(n1136),.clk(gclk));
	jor g1064(.dina(n1136),.dinb(n1130),.dout(n1137),.clk(gclk));
	jor g1065(.dina(n1137),.dinb(n1128),.dout(n1138),.clk(gclk));
	jand g1066(.dina(w_n617_2[0]),.dinb(w_G97_1[2]),.dout(n1139),.clk(gclk));
	jand g1067(.dina(w_n640_2[1]),.dinb(w_G294_1[0]),.dout(n1140),.clk(gclk));
	jand g1068(.dina(w_n642_2[1]),.dinb(w_G116_1[1]),.dout(n1141),.clk(gclk));
	jor g1069(.dina(n1141),.dinb(n1140),.dout(n1142),.clk(gclk));
	jor g1070(.dina(n1142),.dinb(n1139),.dout(n1143),.clk(gclk));
	jand g1071(.dina(w_n631_2[1]),.dinb(w_G303_0[2]),.dout(n1144),.clk(gclk));
	jor g1072(.dina(n1144),.dinb(w_n148_3[0]),.dout(n1145),.clk(gclk));
	jand g1073(.dina(w_n636_2[1]),.dinb(w_G107_1[2]),.dout(n1146),.clk(gclk));
	jand g1074(.dina(w_n627_2[1]),.dinb(w_G283_1[0]),.dout(n1147),.clk(gclk));
	jor g1075(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jor g1076(.dina(w_n899_0[0]),.dinb(w_n825_0[0]),.dout(n1149),.clk(gclk));
	jor g1077(.dina(n1149),.dinb(n1148),.dout(n1150),.clk(gclk));
	jor g1078(.dina(n1150),.dinb(n1145),.dout(n1151),.clk(gclk));
	jor g1079(.dina(n1151),.dinb(n1143),.dout(n1152),.clk(gclk));
	jand g1080(.dina(n1152),.dinb(n1138),.dout(n1153),.clk(gclk));
	jor g1081(.dina(n1153),.dinb(w_n612_1[1]),.dout(n1154),.clk(gclk));
	jand g1082(.dina(w_n743_0[1]),.dinb(w_n75_0[1]),.dout(n1155),.clk(gclk));
	jor g1083(.dina(n1155),.dinb(w_n605_0[1]),.dout(n1156),.clk(gclk));
	jnot g1084(.din(n1156),.dout(n1157),.clk(gclk));
	jand g1085(.dina(n1157),.dinb(n1154),.dout(n1158),.clk(gclk));
	jand g1086(.dina(n1158),.dinb(n1123),.dout(n1159),.clk(gclk));
	jnot g1087(.din(n1159),.dout(n1160),.clk(gclk));
	jand g1088(.dina(n1160),.dinb(n1121),.dout(n1161),.clk(gclk));
	jand g1089(.dina(n1161),.dinb(n1120),.dout(n1162),.clk(gclk));
	jnot g1090(.din(w_n1162_0[2]),.dout(w_dff_A_3TPEWlaZ5_1),.clk(gclk));
	jand g1091(.dina(w_n1114_0[1]),.dinb(w_n1049_0[1]),.dout(n1164),.clk(gclk));
	jnot g1092(.din(w_G387_0[1]),.dout(n1165),.clk(gclk));
	jnot g1093(.din(w_G396_0[1]),.dout(n1166),.clk(gclk));
	jand g1094(.dina(w_n937_0[1]),.dinb(w_dff_B_eHuJ3Zsg4_1),.dout(n1167),.clk(gclk));
	jand g1095(.dina(n1167),.dinb(w_n750_0[0]),.dout(n1168),.clk(gclk));
	jand g1096(.dina(n1168),.dinb(w_n988_0[1]),.dout(n1169),.clk(gclk));
	jand g1097(.dina(n1169),.dinb(w_n1162_0[1]),.dout(n1170),.clk(gclk));
	jand g1098(.dina(n1170),.dinb(n1165),.dout(n1171),.clk(gclk));
	jand g1099(.dina(n1171),.dinb(w_n1164_0[1]),.dout(n1172),.clk(gclk));
	jnot g1100(.din(w_n1172_0[1]),.dout(w_dff_A_snNc0Gbh4_1),.clk(gclk));
	jnot g1101(.din(w_G213_0[1]),.dout(n1174),.clk(gclk));
	jnot g1102(.din(w_G343_0[0]),.dout(n1175),.clk(gclk));
	jand g1103(.dina(w_n1164_0[0]),.dinb(w_n1175_0[1]),.dout(n1176),.clk(gclk));
	jor g1104(.dina(n1176),.dinb(n1174),.dout(n1177),.clk(gclk));
	jor g1105(.dina(n1177),.dinb(w_n1172_0[0]),.dout(G409),.clk(gclk));
	jxor g1106(.dina(w_n1162_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1107(.dina(w_n937_0[0]),.dinb(w_G396_0[0]),.dout(n1180),.clk(gclk));
	jxor g1108(.dina(w_n988_0[0]),.dinb(w_G387_0[0]),.dout(n1181),.clk(gclk));
	jxor g1109(.dina(n1181),.dinb(w_dff_B_kzVggnsM9_1),.dout(n1182),.clk(gclk));
	jxor g1110(.dina(n1182),.dinb(w_dff_B_iCS2njBI1_1),.dout(n1183),.clk(gclk));
	jand g1111(.dina(w_n1175_0[0]),.dinb(w_G213_0[0]),.dout(n1184),.clk(gclk));
	jnot g1112(.din(w_n1184_0[1]),.dout(n1185),.clk(gclk));
	jor g1113(.dina(n1185),.dinb(G2897),.dout(n1186),.clk(gclk));
	jxor g1114(.dina(w_n1114_0[0]),.dinb(w_n1049_0[0]),.dout(n1187),.clk(gclk));
	jor g1115(.dina(w_n1187_0[1]),.dinb(w_n1184_0[0]),.dout(n1188),.clk(gclk));
	jand g1116(.dina(n1188),.dinb(n1186),.dout(n1189),.clk(gclk));
	jxor g1117(.dina(n1189),.dinb(w_n1183_0[1]),.dout(G405),.clk(gclk));
	jxor g1118(.dina(w_n1187_0[0]),.dinb(w_n1183_0[0]),.dout(w_dff_A_Znbnrzrt0_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.doutc(w_G1_2[2]),.din(w_G1_0[1]));
	jspl jspl_w_G1_3(.douta(w_G1_3[0]),.doutb(w_G1_3[1]),.din(w_G1_0[2]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_G13_0[1]),.doutc(w_G13_0[2]),.din(G13));
	jspl jspl_w_G13_1(.douta(w_G13_1[0]),.doutb(w_G13_1[1]),.din(w_G13_0[0]));
	jspl3 jspl3_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_G20_1[0]),.doutb(w_G20_1[1]),.doutc(w_G20_1[2]),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_G20_2[1]),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_G20_3[1]),.doutc(w_G20_3[2]),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_G20_4[0]),.doutb(w_G20_4[1]),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_G20_5[0]),.doutb(w_G20_5[1]),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_G20_6[0]),.doutb(w_G20_6[1]),.doutc(w_G20_6[2]),.din(w_G20_1[2]));
	jspl jspl_w_G20_7(.douta(w_G20_7[0]),.doutb(w_G20_7[1]),.din(w_G20_2[0]));
	jspl3 jspl3_w_G33_0(.douta(w_G33_0[0]),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_G33_1[0]),.doutb(w_G33_1[1]),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_G33_3[2]),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_G33_4[1]),.doutc(w_G33_4[2]),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_G33_5[0]),.doutb(w_G33_5[1]),.doutc(w_G33_5[2]),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_G33_6[0]),.doutb(w_G33_6[1]),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_G33_8[0]),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_G33_9[0]),.doutb(w_G33_9[1]),.doutc(w_G33_9[2]),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_G33_10[0]),.doutb(w_G33_10[1]),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.doutc(w_G41_0[2]),.din(G41));
	jspl jspl_w_G41_1(.douta(w_G41_1[0]),.doutb(w_G41_1[1]),.din(w_G41_0[0]));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_G45_0[1]),.doutc(w_G45_0[2]),.din(G45));
	jspl3 jspl3_w_G45_1(.douta(w_G45_1[0]),.doutb(w_G45_1[1]),.doutc(w_G45_1[2]),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_G50_0[1]),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_G50_1[0]),.doutb(w_G50_1[1]),.doutc(w_G50_1[2]),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_G50_2[0]),.doutb(w_G50_2[1]),.doutc(w_G50_2[2]),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_G50_3[0]),.doutb(w_G50_3[1]),.doutc(w_G50_3[2]),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_G50_4[0]),.doutb(w_G50_4[1]),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_G50_5[1]),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_G58_0[1]),.doutc(w_G58_0[2]),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_G58_1[0]),.doutb(w_G58_1[1]),.doutc(w_G58_1[2]),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_G58_2[0]),.doutb(w_G58_2[1]),.doutc(w_G58_2[2]),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_G58_3[0]),.doutb(w_G58_3[1]),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_G58_4[0]),.doutb(w_G58_4[1]),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl jspl_w_G58_5(.douta(w_G58_5[0]),.doutb(w_G58_5[1]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_G68_0[2]),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_G68_1[0]),.doutb(w_G68_1[1]),.doutc(w_G68_1[2]),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_G68_2[1]),.doutc(w_G68_2[2]),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_G68_3[1]),.doutc(w_G68_3[2]),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_G68_4[0]),.doutb(w_G68_4[1]),.doutc(w_G68_4[2]),.din(w_G68_1[0]));
	jspl jspl_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_G77_0[1]),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_G77_1[0]),.doutb(w_G77_1[1]),.doutc(w_G77_1[2]),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_G77_2[0]),.doutb(w_G77_2[1]),.doutc(w_G77_2[2]),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_G77_3[0]),.doutb(w_G77_3[1]),.doutc(w_G77_3[2]),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_G77_4[0]),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl jspl_w_G77_5(.douta(w_G77_5[0]),.doutb(w_G77_5[1]),.din(w_G77_1[1]));
	jspl3 jspl3_w_G87_0(.douta(w_G87_0[0]),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_G87_1[1]),.doutc(w_G87_1[2]),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_G87_2[0]),.doutb(w_G87_2[1]),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_G87_3[0]),.doutb(w_G87_3[1]),.doutc(w_G87_3[2]),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_G97_0[1]),.doutc(w_G97_0[2]),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_G97_1[2]),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_G97_2[2]),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_G97_3[0]),.doutb(w_G97_3[1]),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_G97_4[0]),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl jspl_w_G97_5(.douta(w_G97_5[0]),.doutb(w_G97_5[1]),.din(w_G97_1[1]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_G107_1[2]),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_G107_2[2]),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_G107_3[0]),.doutb(w_G107_3[1]),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl3 jspl3_w_G107_4(.douta(w_G107_4[0]),.doutb(w_G107_4[1]),.doutc(w_G107_4[2]),.din(w_G107_1[0]));
	jspl jspl_w_G107_5(.douta(w_G107_5[0]),.doutb(w_G107_5[1]),.din(w_G107_1[1]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_G116_1[1]),.doutc(w_G116_1[2]),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_G116_2[1]),.doutc(w_G116_2[2]),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_G116_3[0]),.doutb(w_G116_3[1]),.doutc(w_G116_3[2]),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_G116_4[0]),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_G125_0[1]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(G132));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_G132_1[1]),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_G137_1[1]),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.doutc(w_G143_1[2]),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_G150_0[0]),.doutb(w_G150_0[1]),.doutc(w_G150_0[2]),.din(G150));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_G150_1[1]),.doutc(w_G150_1[2]),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_G150_2[1]),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_G150_3[0]),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_G159_0[0]),.doutb(w_G159_0[1]),.doutc(w_G159_0[2]),.din(G159));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_G159_3[0]),.doutb(w_G159_3[1]),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_G169_0[0]),.doutb(w_G169_0[1]),.doutc(w_G169_0[2]),.din(G169));
	jspl jspl_w_G169_1(.douta(w_G169_1[0]),.doutb(w_G169_1[1]),.din(w_G169_0[0]));
	jspl3 jspl3_w_G179_0(.douta(w_G179_0[0]),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_G179_2[0]),.doutb(w_G179_2[1]),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_G190_0[0]),.doutb(w_G190_0[1]),.doutc(w_G190_0[2]),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_G190_1[0]),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_G190_2[1]),.doutc(w_G190_2[2]),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_G190_3[1]),.doutc(w_G190_3[2]),.din(w_G190_0[2]));
	jspl jspl_w_G190_4(.douta(w_G190_4[0]),.doutb(w_G190_4[1]),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_G200_0[2]),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_G200_1[0]),.doutb(w_G200_1[1]),.doutc(w_G200_1[2]),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_G200_2[1]),.doutc(w_G200_2[2]),.din(w_G200_0[1]));
	jspl3 jspl3_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.doutc(w_G200_3[2]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G200_4(.douta(w_G200_4[0]),.doutb(w_G200_4[1]),.doutc(w_G200_4[2]),.din(w_G200_1[0]));
	jspl3 jspl3_w_G213_0(.douta(w_G213_0[0]),.doutb(w_G213_0[1]),.doutc(w_G213_0[2]),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(G223));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl jspl_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_G232_0[1]),.doutc(w_G232_0[2]),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_G232_1[0]),.doutb(w_G232_1[1]),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_G238_0[1]),.doutc(w_G238_0[2]),.din(G238));
	jspl3 jspl3_w_G238_1(.douta(w_G238_1[0]),.doutb(w_G238_1[1]),.doutc(w_G238_1[2]),.din(w_G238_0[0]));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_G244_0[1]),.doutc(w_G244_0[2]),.din(G244));
	jspl3 jspl3_w_G244_1(.douta(w_G244_1[0]),.doutb(w_G244_1[1]),.doutc(w_G244_1[2]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_G250_0[0]),.doutb(w_G250_0[1]),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_G264_0[0]),.doutb(w_G264_0[1]),.doutc(w_G264_0[2]),.din(G264));
	jspl jspl_w_G264_1(.douta(w_G264_1[0]),.doutb(w_G264_1[1]),.din(w_G264_0[0]));
	jspl3 jspl3_w_G270_0(.douta(w_G270_0[0]),.doutb(w_G270_0[1]),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_G274_0[0]),.doutb(w_G274_0[1]),.doutc(w_G274_0[2]),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_G283_0[0]),.doutb(w_G283_0[1]),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_G283_1[1]),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_G283_2[0]),.doutb(w_G283_2[1]),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_G283_3[0]),.doutb(w_G283_3[1]),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_G294_0[0]),.doutb(w_G294_0[1]),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_G294_1[1]),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_G294_2[0]),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_G294_3[0]),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_G303_0[0]),.doutb(w_G303_0[1]),.doutc(w_G303_0[2]),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_G303_2[0]),.doutb(w_G303_2[1]),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(G311));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_G311_1[1]),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(G317));
	jspl jspl_w_G317_1(.douta(w_G317_1[0]),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_G322_0[0]),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(G322));
	jspl jspl_w_G326_0(.douta(w_G326_0[0]),.doutb(w_G326_0[1]),.din(G326));
	jspl jspl_w_G330_0(.douta(w_G330_0[0]),.doutb(w_G330_0[1]),.din(G330));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_G343_0[1]),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_G1698_0[2]),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_G355_0),.doutb(w_dff_A_cyNhmvic6_1),.din(G355_fa_));
	jspl3 jspl3_w_G396_0(.douta(w_dff_A_ZMqnxzvf1_0),.doutb(w_G396_0[1]),.doutc(w_dff_A_QVGVQfYK5_2),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_mWJJ95QE5_0),.doutb(w_dff_A_CAs6wypP0_1),.din(G384_fa_));
	jspl3 jspl3_w_G387_0(.douta(w_G387_0[0]),.doutb(w_G387_0[1]),.doutc(w_dff_A_iCSTSP0S7_2),.din(G387_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_n72_0[1]),.doutc(w_n72_0[2]),.din(n72));
	jspl jspl_w_n72_1(.douta(w_n72_1[0]),.doutb(w_n72_1[1]),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_n73_0[2]),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_n73_1[1]),.doutc(w_n73_1[2]),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_n73_2[0]),.doutb(w_n73_2[1]),.doutc(w_n73_2[2]),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.doutc(w_n75_0[2]),.din(n75));
	jspl jspl_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.din(w_n75_0[0]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl jspl_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.doutc(w_n85_0[2]),.din(n85));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.doutc(w_n88_0[2]),.din(n88));
	jspl jspl_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.din(w_n88_0[0]));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_n91_1[0]),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl3 jspl3_w_n97_1(.douta(w_n97_1[0]),.doutb(w_n97_1[1]),.doutc(w_n97_1[2]),.din(w_n97_0[0]));
	jspl jspl_w_n97_2(.douta(w_n97_2[0]),.doutb(w_n97_2[1]),.din(w_n97_0[1]));
	jspl3 jspl3_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.doutc(w_n98_0[2]),.din(n98));
	jspl3 jspl3_w_n98_1(.douta(w_n98_1[0]),.doutb(w_n98_1[1]),.doutc(w_n98_1[2]),.din(w_n98_0[0]));
	jspl jspl_w_n98_2(.douta(w_n98_2[0]),.doutb(w_n98_2[1]),.din(w_n98_0[1]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n105_0(.douta(w_n105_0[0]),.doutb(w_n105_0[1]),.doutc(w_n105_0[2]),.din(n105));
	jspl3 jspl3_w_n105_1(.douta(w_n105_1[0]),.doutb(w_n105_1[1]),.doutc(w_n105_1[2]),.din(w_n105_0[0]));
	jspl jspl_w_n105_2(.douta(w_n105_2[0]),.doutb(w_n105_2[1]),.din(w_n105_0[1]));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl3 jspl3_w_n112_3(.douta(w_n112_3[0]),.doutb(w_n112_3[1]),.doutc(w_n112_3[2]),.din(w_n112_0[2]));
	jspl3 jspl3_w_n112_4(.douta(w_n112_4[0]),.doutb(w_n112_4[1]),.doutc(w_n112_4[2]),.din(w_n112_1[0]));
	jspl3 jspl3_w_n112_5(.douta(w_n112_5[0]),.doutb(w_n112_5[1]),.doutc(w_n112_5[2]),.din(w_n112_1[1]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl3 jspl3_w_n113_1(.douta(w_n113_1[0]),.doutb(w_n113_1[1]),.doutc(w_n113_1[2]),.din(w_n113_0[0]));
	jspl3 jspl3_w_n113_2(.douta(w_n113_2[0]),.doutb(w_n113_2[1]),.doutc(w_n113_2[2]),.din(w_n113_0[1]));
	jspl jspl_w_n113_3(.douta(w_n113_3[0]),.doutb(w_n113_3[1]),.din(w_n113_0[2]));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl3 jspl3_w_n114_1(.douta(w_n114_1[0]),.doutb(w_n114_1[1]),.doutc(w_n114_1[2]),.din(w_n114_0[0]));
	jspl3 jspl3_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.doutc(w_n115_0[2]),.din(n115));
	jspl jspl_w_n115_1(.douta(w_n115_1[0]),.doutb(w_n115_1[1]),.din(w_n115_0[0]));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.din(n116));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl3 jspl3_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.doutc(w_n123_1[2]),.din(w_n123_0[0]));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.din(n135));
	jspl3 jspl3_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.doutc(w_n137_0[2]),.din(n137));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(n144));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.doutc(w_n146_0[2]),.din(n146));
	jspl3 jspl3_w_n146_1(.douta(w_n146_1[0]),.doutb(w_n146_1[1]),.doutc(w_n146_1[2]),.din(w_n146_0[0]));
	jspl3 jspl3_w_n146_2(.douta(w_n146_2[0]),.doutb(w_n146_2[1]),.doutc(w_n146_2[2]),.din(w_n146_0[1]));
	jspl3 jspl3_w_n146_3(.douta(w_n146_3[0]),.doutb(w_n146_3[1]),.doutc(w_n146_3[2]),.din(w_n146_0[2]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.doutc(w_n148_1[2]),.din(w_n148_0[0]));
	jspl3 jspl3_w_n148_2(.douta(w_n148_2[0]),.doutb(w_n148_2[1]),.doutc(w_n148_2[2]),.din(w_n148_0[1]));
	jspl3 jspl3_w_n148_3(.douta(w_n148_3[0]),.doutb(w_n148_3[1]),.doutc(w_n148_3[2]),.din(w_n148_0[2]));
	jspl3 jspl3_w_n148_4(.douta(w_n148_4[0]),.doutb(w_n148_4[1]),.doutc(w_n148_4[2]),.din(w_n148_1[0]));
	jspl3 jspl3_w_n148_5(.douta(w_n148_5[0]),.doutb(w_n148_5[1]),.doutc(w_n148_5[2]),.din(w_n148_1[1]));
	jspl3 jspl3_w_n148_6(.douta(w_n148_6[0]),.doutb(w_n148_6[1]),.doutc(w_n148_6[2]),.din(w_n148_1[2]));
	jspl3 jspl3_w_n148_7(.douta(w_n148_7[0]),.doutb(w_n148_7[1]),.doutc(w_n148_7[2]),.din(w_n148_2[0]));
	jspl3 jspl3_w_n148_8(.douta(w_n148_8[0]),.doutb(w_n148_8[1]),.doutc(w_n148_8[2]),.din(w_n148_2[1]));
	jspl3 jspl3_w_n148_9(.douta(w_n148_9[0]),.doutb(w_n148_9[1]),.doutc(w_n148_9[2]),.din(w_n148_2[2]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_n149_2[0]),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_n151_1[1]),.doutc(w_n151_1[2]),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_n151_3[0]),.doutb(w_n151_3[1]),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_n151_4[1]),.doutc(w_n151_4[2]),.din(w_n151_1[0]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n152_1(.douta(w_n152_1[0]),.doutb(w_n152_1[1]),.doutc(w_n152_1[2]),.din(w_n152_0[0]));
	jspl3 jspl3_w_n152_2(.douta(w_n152_2[0]),.doutb(w_n152_2[1]),.doutc(w_n152_2[2]),.din(w_n152_0[1]));
	jspl jspl_w_n152_3(.douta(w_n152_3[0]),.doutb(w_n152_3[1]),.din(w_n152_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n155_2(.douta(w_n155_2[0]),.doutb(w_n155_2[1]),.doutc(w_n155_2[2]),.din(w_n155_0[1]));
	jspl jspl_w_n155_3(.douta(w_n155_3[0]),.doutb(w_n155_3[1]),.din(w_n155_0[2]));
	jspl3 jspl3_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.doutc(w_n157_0[2]),.din(n157));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.doutc(w_n166_1[2]),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_n166_2[2]),.din(w_n166_0[1]));
	jspl jspl_w_n166_3(.douta(w_n166_3[0]),.doutb(w_n166_3[1]),.din(w_n166_0[2]));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.doutc(w_n179_0[2]),.din(n179));
	jspl3 jspl3_w_n179_1(.douta(w_n179_1[0]),.doutb(w_n179_1[1]),.doutc(w_n179_1[2]),.din(w_n179_0[0]));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_n185_1[2]),.din(w_n185_0[0]));
	jspl3 jspl3_w_n185_2(.douta(w_n185_2[0]),.doutb(w_n185_2[1]),.doutc(w_n185_2[2]),.din(w_n185_0[1]));
	jspl3 jspl3_w_n185_3(.douta(w_n185_3[0]),.doutb(w_n185_3[1]),.doutc(w_n185_3[2]),.din(w_n185_0[2]));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_n189_0[2]),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_n189_1[1]),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl jspl_w_n189_2(.douta(w_n189_2[0]),.doutb(w_n189_2[1]),.din(w_n189_0[1]));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl3 jspl3_w_n190_1(.douta(w_n190_1[0]),.doutb(w_n190_1[1]),.doutc(w_n190_1[2]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl3 jspl3_w_n196_1(.douta(w_n196_1[0]),.doutb(w_n196_1[1]),.doutc(w_n196_1[2]),.din(w_n196_0[0]));
	jspl3 jspl3_w_n196_2(.douta(w_n196_2[0]),.doutb(w_n196_2[1]),.doutc(w_n196_2[2]),.din(w_n196_0[1]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n199_1(.douta(w_n199_1[0]),.doutb(w_n199_1[1]),.din(w_n199_0[0]));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.doutc(w_n210_0[2]),.din(n210));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.din(n214));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl3 jspl3_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.doutc(w_n221_0[2]),.din(n221));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(n229));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.din(w_n246_0[0]));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.doutc(w_n274_0[2]),.din(n274));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.din(n281));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.din(w_n288_0[0]));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(n300));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_n339_0[1]),.din(n339));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl jspl_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.din(w_n355_0[0]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.doutc(w_n382_0[2]),.din(n382));
	jspl jspl_w_n382_1(.douta(w_n382_1[0]),.doutb(w_n382_1[1]),.din(w_n382_0[0]));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl jspl_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.doutc(w_n407_0[2]),.din(n407));
	jspl3 jspl3_w_n407_1(.douta(w_n407_1[0]),.doutb(w_n407_1[1]),.doutc(w_n407_1[2]),.din(w_n407_0[0]));
	jspl jspl_w_n407_2(.douta(w_n407_2[0]),.doutb(w_n407_2[1]),.din(w_n407_0[1]));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl3 jspl3_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jspl jspl_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.din(w_n420_0[0]));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n425_1(.douta(w_n425_1[0]),.doutb(w_n425_1[1]),.doutc(w_n425_1[2]),.din(w_n425_0[0]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.din(w_n439_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl3 jspl3_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.doutc(w_n455_0[2]),.din(n455));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.din(n475));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.doutc(w_n492_0[2]),.din(n492));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.doutc(w_n519_0[2]),.din(n519));
	jspl3 jspl3_w_n519_1(.douta(w_n519_1[0]),.doutb(w_n519_1[1]),.doutc(w_n519_1[2]),.din(w_n519_0[0]));
	jspl jspl_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.doutc(w_n536_0[2]),.din(n536));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl3 jspl3_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.doutc(w_n542_0[2]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.doutc(w_n548_0[2]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.doutc(w_n552_0[2]),.din(n552));
	jspl jspl_w_n552_1(.douta(w_n552_1[0]),.doutb(w_n552_1[1]),.din(w_n552_0[0]));
	jspl3 jspl3_w_n553_0(.douta(w_n553_0[0]),.doutb(w_n553_0[1]),.doutc(w_n553_0[2]),.din(n553));
	jspl3 jspl3_w_n553_1(.douta(w_n553_1[0]),.doutb(w_n553_1[1]),.doutc(w_n553_1[2]),.din(w_n553_0[0]));
	jspl3 jspl3_w_n553_2(.douta(w_n553_2[0]),.doutb(w_n553_2[1]),.doutc(w_n553_2[2]),.din(w_n553_0[1]));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.doutc(w_n554_0[2]),.din(n554));
	jspl3 jspl3_w_n554_1(.douta(w_n554_1[0]),.doutb(w_n554_1[1]),.doutc(w_n554_1[2]),.din(w_n554_0[0]));
	jspl3 jspl3_w_n554_2(.douta(w_n554_2[0]),.doutb(w_n554_2[1]),.doutc(w_n554_2[2]),.din(w_n554_0[1]));
	jspl3 jspl3_w_n554_3(.douta(w_n554_3[0]),.doutb(w_n554_3[1]),.doutc(w_n554_3[2]),.din(w_n554_0[2]));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(n556));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.doutc(w_n563_0[2]),.din(n563));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(n567));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n576_1(.douta(w_n576_1[0]),.doutb(w_n576_1[1]),.din(w_n576_0[0]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl3 jspl3_w_n589_1(.douta(w_n589_1[0]),.doutb(w_n589_1[1]),.doutc(w_n589_1[2]),.din(w_n589_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.doutc(w_n592_0[2]),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_n592_1[0]),.doutb(w_n592_1[1]),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl jspl_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.din(w_n592_0[1]));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl3 jspl3_w_n603_1(.douta(w_n603_1[0]),.doutb(w_n603_1[1]),.doutc(w_n603_1[2]),.din(w_n603_0[0]));
	jspl jspl_w_n603_2(.douta(w_n603_2[0]),.doutb(w_n603_2[1]),.din(w_n603_0[1]));
	jspl3 jspl3_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_n604_1[0]),.doutb(w_n604_1[1]),.doutc(w_n604_1[2]),.din(w_n604_0[0]));
	jspl jspl_w_n604_2(.douta(w_n604_2[0]),.doutb(w_n604_2[1]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_n605_1[2]),.din(w_n605_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.doutc(w_n608_0[2]),.din(n608));
	jspl3 jspl3_w_n608_1(.douta(w_n608_1[0]),.doutb(w_n608_1[1]),.doutc(w_n608_1[2]),.din(w_n608_0[0]));
	jspl3 jspl3_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.doutc(w_n612_0[2]),.din(n612));
	jspl3 jspl3_w_n612_1(.douta(w_n612_1[0]),.doutb(w_n612_1[1]),.doutc(w_n612_1[2]),.din(w_n612_0[0]));
	jspl3 jspl3_w_n612_2(.douta(w_n612_2[0]),.doutb(w_n612_2[1]),.doutc(w_n612_2[2]),.din(w_n612_0[1]));
	jspl3 jspl3_w_n612_3(.douta(w_n612_3[0]),.doutb(w_n612_3[1]),.doutc(w_n612_3[2]),.din(w_n612_0[2]));
	jspl jspl_w_n612_4(.douta(w_n612_4[0]),.doutb(w_n612_4[1]),.din(w_n612_1[0]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl jspl_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.din(w_n613_0[0]));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl3 jspl3_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.doutc(w_n617_1[2]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n617_2(.douta(w_n617_2[0]),.doutb(w_n617_2[1]),.doutc(w_n617_2[2]),.din(w_n617_0[1]));
	jspl3 jspl3_w_n617_3(.douta(w_n617_3[0]),.doutb(w_n617_3[1]),.doutc(w_n617_3[2]),.din(w_n617_0[2]));
	jspl3 jspl3_w_n617_4(.douta(w_n617_4[0]),.doutb(w_n617_4[1]),.doutc(w_n617_4[2]),.din(w_n617_1[0]));
	jspl3 jspl3_w_n617_5(.douta(w_n617_5[0]),.doutb(w_n617_5[1]),.doutc(w_n617_5[2]),.din(w_n617_1[1]));
	jspl jspl_w_n617_6(.douta(w_n617_6[0]),.doutb(w_n617_6[1]),.din(w_n617_1[2]));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.doutc(w_n623_0[2]),.din(n623));
	jspl3 jspl3_w_n623_1(.douta(w_n623_1[0]),.doutb(w_n623_1[1]),.doutc(w_n623_1[2]),.din(w_n623_0[0]));
	jspl3 jspl3_w_n623_2(.douta(w_n623_2[0]),.doutb(w_n623_2[1]),.doutc(w_n623_2[2]),.din(w_n623_0[1]));
	jspl3 jspl3_w_n623_3(.douta(w_n623_3[0]),.doutb(w_n623_3[1]),.doutc(w_n623_3[2]),.din(w_n623_0[2]));
	jspl3 jspl3_w_n623_4(.douta(w_n623_4[0]),.doutb(w_n623_4[1]),.doutc(w_n623_4[2]),.din(w_n623_1[0]));
	jspl jspl_w_n623_5(.douta(w_n623_5[0]),.doutb(w_n623_5[1]),.din(w_n623_1[1]));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl3 jspl3_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.doutc(w_n627_1[2]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n627_2(.douta(w_n627_2[0]),.doutb(w_n627_2[1]),.doutc(w_n627_2[2]),.din(w_n627_0[1]));
	jspl3 jspl3_w_n627_3(.douta(w_n627_3[0]),.doutb(w_n627_3[1]),.doutc(w_n627_3[2]),.din(w_n627_0[2]));
	jspl3 jspl3_w_n627_4(.douta(w_n627_4[0]),.doutb(w_n627_4[1]),.doutc(w_n627_4[2]),.din(w_n627_1[0]));
	jspl3 jspl3_w_n627_5(.douta(w_n627_5[0]),.doutb(w_n627_5[1]),.doutc(w_n627_5[2]),.din(w_n627_1[1]));
	jspl3 jspl3_w_n627_6(.douta(w_n627_6[0]),.doutb(w_n627_6[1]),.doutc(w_n627_6[2]),.din(w_n627_1[2]));
	jspl jspl_w_n627_7(.douta(w_n627_7[0]),.doutb(w_n627_7[1]),.din(w_n627_2[0]));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n631_1(.douta(w_n631_1[0]),.doutb(w_n631_1[1]),.doutc(w_n631_1[2]),.din(w_n631_0[0]));
	jspl3 jspl3_w_n631_2(.douta(w_n631_2[0]),.doutb(w_n631_2[1]),.doutc(w_n631_2[2]),.din(w_n631_0[1]));
	jspl3 jspl3_w_n631_3(.douta(w_n631_3[0]),.doutb(w_n631_3[1]),.doutc(w_n631_3[2]),.din(w_n631_0[2]));
	jspl3 jspl3_w_n631_4(.douta(w_n631_4[0]),.doutb(w_n631_4[1]),.doutc(w_n631_4[2]),.din(w_n631_1[0]));
	jspl3 jspl3_w_n631_5(.douta(w_n631_5[0]),.doutb(w_n631_5[1]),.doutc(w_n631_5[2]),.din(w_n631_1[1]));
	jspl3 jspl3_w_n631_6(.douta(w_n631_6[0]),.doutb(w_n631_6[1]),.doutc(w_n631_6[2]),.din(w_n631_1[2]));
	jspl jspl_w_n631_7(.douta(w_n631_7[0]),.doutb(w_n631_7[1]),.din(w_n631_2[0]));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n634_1(.douta(w_n634_1[0]),.doutb(w_n634_1[1]),.doutc(w_n634_1[2]),.din(w_n634_0[0]));
	jspl3 jspl3_w_n634_2(.douta(w_n634_2[0]),.doutb(w_n634_2[1]),.doutc(w_n634_2[2]),.din(w_n634_0[1]));
	jspl3 jspl3_w_n634_3(.douta(w_n634_3[0]),.doutb(w_n634_3[1]),.doutc(w_n634_3[2]),.din(w_n634_0[2]));
	jspl jspl_w_n634_4(.douta(w_n634_4[0]),.doutb(w_n634_4[1]),.din(w_n634_1[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n636_1(.douta(w_n636_1[0]),.doutb(w_n636_1[1]),.doutc(w_n636_1[2]),.din(w_n636_0[0]));
	jspl3 jspl3_w_n636_2(.douta(w_n636_2[0]),.doutb(w_n636_2[1]),.doutc(w_n636_2[2]),.din(w_n636_0[1]));
	jspl3 jspl3_w_n636_3(.douta(w_n636_3[0]),.doutb(w_n636_3[1]),.doutc(w_n636_3[2]),.din(w_n636_0[2]));
	jspl3 jspl3_w_n636_4(.douta(w_n636_4[0]),.doutb(w_n636_4[1]),.doutc(w_n636_4[2]),.din(w_n636_1[0]));
	jspl3 jspl3_w_n636_5(.douta(w_n636_5[0]),.doutb(w_n636_5[1]),.doutc(w_n636_5[2]),.din(w_n636_1[1]));
	jspl3 jspl3_w_n636_6(.douta(w_n636_6[0]),.doutb(w_n636_6[1]),.doutc(w_n636_6[2]),.din(w_n636_1[2]));
	jspl jspl_w_n636_7(.douta(w_n636_7[0]),.doutb(w_n636_7[1]),.din(w_n636_2[0]));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl3 jspl3_w_n642_1(.douta(w_n642_1[0]),.doutb(w_n642_1[1]),.doutc(w_n642_1[2]),.din(w_n642_0[0]));
	jspl3 jspl3_w_n642_2(.douta(w_n642_2[0]),.doutb(w_n642_2[1]),.doutc(w_n642_2[2]),.din(w_n642_0[1]));
	jspl3 jspl3_w_n642_3(.douta(w_n642_3[0]),.doutb(w_n642_3[1]),.doutc(w_n642_3[2]),.din(w_n642_0[2]));
	jspl3 jspl3_w_n642_4(.douta(w_n642_4[0]),.doutb(w_n642_4[1]),.doutc(w_n642_4[2]),.din(w_n642_1[0]));
	jspl3 jspl3_w_n642_5(.douta(w_n642_5[0]),.doutb(w_n642_5[1]),.doutc(w_n642_5[2]),.din(w_n642_1[1]));
	jspl3 jspl3_w_n642_6(.douta(w_n642_6[0]),.doutb(w_n642_6[1]),.doutc(w_n642_6[2]),.din(w_n642_1[2]));
	jspl jspl_w_n642_7(.douta(w_n642_7[0]),.doutb(w_n642_7[1]),.din(w_n642_2[0]));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_n672_0[2]),.din(n672));
	jspl jspl_w_n672_1(.douta(w_n672_1[0]),.doutb(w_n672_1[1]),.din(w_n672_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.doutc(w_n696_0[2]),.din(n696));
	jspl3 jspl3_w_n696_1(.douta(w_n696_1[0]),.doutb(w_n696_1[1]),.doutc(w_n696_1[2]),.din(w_n696_0[0]));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl jspl_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.din(w_n743_0[0]));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_n758_1[1]),.din(w_n758_0[0]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_n764_0[2]),.din(n764));
	jspl3 jspl3_w_n764_1(.douta(w_n764_1[0]),.doutb(w_n764_1[1]),.doutc(w_n764_1[2]),.din(w_n764_0[0]));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.doutc(w_n853_0[2]),.din(n853));
	jspl3 jspl3_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl3 jspl3_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.doutc(w_n861_0[2]),.din(n861));
	jspl jspl_w_n861_1(.douta(w_n861_1[0]),.doutb(w_n861_1[1]),.din(w_n861_0[0]));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.din(n940));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl3 jspl3_w_n988_0(.douta(w_dff_A_ZQmF1xtq7_0),.doutb(w_dff_A_qaUH8K5X8_1),.doutc(w_n988_0[2]),.din(n988));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(n990));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl3 jspl3_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.doutc(w_n1001_0[2]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.doutc(w_n1002_0[2]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl3 jspl3_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.doutc(w_n1049_0[2]),.din(n1049));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_dff_A_Y8dPIE7f0_1),.doutc(w_n1162_0[2]),.din(n1162));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1172_0(.douta(w_dff_A_JD9tOuMB5_0),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(n1175));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_dff_A_RftdTNmm0_1),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(n1184));
	jspl jspl_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.din(n1187));
	jdff dff_B_M2bk8CTR9_1(.din(n111),.dout(w_dff_B_M2bk8CTR9_1),.clk(gclk));
	jdff dff_B_L5K1pX3c9_1(.din(n540),.dout(w_dff_B_L5K1pX3c9_1),.clk(gclk));
	jdff dff_B_tdIYQyy51_0(.din(n597),.dout(w_dff_B_tdIYQyy51_0),.clk(gclk));
	jdff dff_B_hLperUKE3_0(.din(w_dff_B_tdIYQyy51_0),.dout(w_dff_B_hLperUKE3_0),.clk(gclk));
	jdff dff_B_eTKitgFn8_0(.din(w_dff_B_hLperUKE3_0),.dout(w_dff_B_eTKitgFn8_0),.clk(gclk));
	jdff dff_B_YXcrKEAJ2_0(.din(w_dff_B_eTKitgFn8_0),.dout(w_dff_B_YXcrKEAJ2_0),.clk(gclk));
	jdff dff_B_39kMmzie6_0(.din(w_dff_B_YXcrKEAJ2_0),.dout(w_dff_B_39kMmzie6_0),.clk(gclk));
	jdff dff_B_cbUMfDkb0_0(.din(w_dff_B_39kMmzie6_0),.dout(w_dff_B_cbUMfDkb0_0),.clk(gclk));
	jdff dff_B_dFj2zYCq7_0(.din(w_dff_B_cbUMfDkb0_0),.dout(w_dff_B_dFj2zYCq7_0),.clk(gclk));
	jdff dff_B_lVRXuHPs2_0(.din(w_dff_B_dFj2zYCq7_0),.dout(w_dff_B_lVRXuHPs2_0),.clk(gclk));
	jdff dff_B_BEtrxYBi6_0(.din(w_dff_B_lVRXuHPs2_0),.dout(w_dff_B_BEtrxYBi6_0),.clk(gclk));
	jdff dff_B_emsRcblk9_0(.din(w_dff_B_BEtrxYBi6_0),.dout(w_dff_B_emsRcblk9_0),.clk(gclk));
	jdff dff_B_MbNWeus15_0(.din(n795),.dout(w_dff_B_MbNWeus15_0),.clk(gclk));
	jdff dff_B_RM9HVZop1_0(.din(w_dff_B_MbNWeus15_0),.dout(w_dff_B_RM9HVZop1_0),.clk(gclk));
	jdff dff_B_4chH4i9T0_0(.din(w_dff_B_RM9HVZop1_0),.dout(w_dff_B_4chH4i9T0_0),.clk(gclk));
	jdff dff_B_9PPINYUl7_0(.din(w_dff_B_4chH4i9T0_0),.dout(w_dff_B_9PPINYUl7_0),.clk(gclk));
	jdff dff_B_J5SzWb9M1_0(.din(w_dff_B_9PPINYUl7_0),.dout(w_dff_B_J5SzWb9M1_0),.clk(gclk));
	jdff dff_B_A9nccNNq1_0(.din(w_dff_B_J5SzWb9M1_0),.dout(w_dff_B_A9nccNNq1_0),.clk(gclk));
	jdff dff_B_8MfOWSig9_0(.din(w_dff_B_A9nccNNq1_0),.dout(w_dff_B_8MfOWSig9_0),.clk(gclk));
	jdff dff_B_A4TviHsX6_0(.din(w_dff_B_8MfOWSig9_0),.dout(w_dff_B_A4TviHsX6_0),.clk(gclk));
	jdff dff_B_YMeEVwok3_0(.din(w_dff_B_A4TviHsX6_0),.dout(w_dff_B_YMeEVwok3_0),.clk(gclk));
	jdff dff_B_MCk3Ssc73_0(.din(w_dff_B_YMeEVwok3_0),.dout(w_dff_B_MCk3Ssc73_0),.clk(gclk));
	jdff dff_B_QiudUgjP3_0(.din(w_dff_B_MCk3Ssc73_0),.dout(w_dff_B_QiudUgjP3_0),.clk(gclk));
	jdff dff_B_KYiqwOBi3_0(.din(w_dff_B_QiudUgjP3_0),.dout(w_dff_B_KYiqwOBi3_0),.clk(gclk));
	jdff dff_B_Irm9ncJQ4_0(.din(w_dff_B_KYiqwOBi3_0),.dout(w_dff_B_Irm9ncJQ4_0),.clk(gclk));
	jdff dff_B_JQkHdphv9_0(.din(w_dff_B_Irm9ncJQ4_0),.dout(w_dff_B_JQkHdphv9_0),.clk(gclk));
	jdff dff_B_bDJtiRpV7_0(.din(w_dff_B_JQkHdphv9_0),.dout(w_dff_B_bDJtiRpV7_0),.clk(gclk));
	jdff dff_B_qZMCsC4o3_0(.din(w_dff_B_bDJtiRpV7_0),.dout(w_dff_B_qZMCsC4o3_0),.clk(gclk));
	jdff dff_B_gaRAddgQ5_0(.din(w_dff_B_qZMCsC4o3_0),.dout(w_dff_B_gaRAddgQ5_0),.clk(gclk));
	jdff dff_A_JD9tOuMB5_0(.dout(w_n1172_0[0]),.din(w_dff_A_JD9tOuMB5_0),.clk(gclk));
	jdff dff_B_DTvBXyOK4_1(.din(n1166),.dout(w_dff_B_DTvBXyOK4_1),.clk(gclk));
	jdff dff_B_eHuJ3Zsg4_1(.din(w_dff_B_DTvBXyOK4_1),.dout(w_dff_B_eHuJ3Zsg4_1),.clk(gclk));
	jdff dff_A_RftdTNmm0_1(.dout(w_n1183_0[1]),.din(w_dff_A_RftdTNmm0_1),.clk(gclk));
	jdff dff_B_5PKNBKz49_1(.din(n1179),.dout(w_dff_B_5PKNBKz49_1),.clk(gclk));
	jdff dff_B_iCS2njBI1_1(.din(w_dff_B_5PKNBKz49_1),.dout(w_dff_B_iCS2njBI1_1),.clk(gclk));
	jdff dff_B_Xbn8CJNi1_1(.din(n1180),.dout(w_dff_B_Xbn8CJNi1_1),.clk(gclk));
	jdff dff_B_NFbYal1R0_1(.din(w_dff_B_Xbn8CJNi1_1),.dout(w_dff_B_NFbYal1R0_1),.clk(gclk));
	jdff dff_B_kzVggnsM9_1(.din(w_dff_B_NFbYal1R0_1),.dout(w_dff_B_kzVggnsM9_1),.clk(gclk));
	jdff dff_A_EeJc0YC55_0(.dout(w_n988_0[0]),.din(w_dff_A_EeJc0YC55_0),.clk(gclk));
	jdff dff_A_ZQmF1xtq7_0(.dout(w_dff_A_EeJc0YC55_0),.din(w_dff_A_ZQmF1xtq7_0),.clk(gclk));
	jdff dff_A_qaUH8K5X8_1(.dout(w_n988_0[1]),.din(w_dff_A_qaUH8K5X8_1),.clk(gclk));
	jdff dff_A_4C8JbJYO9_0(.dout(w_G396_0[0]),.din(w_dff_A_4C8JbJYO9_0),.clk(gclk));
	jdff dff_A_VmTMOllq2_0(.dout(w_dff_A_4C8JbJYO9_0),.din(w_dff_A_VmTMOllq2_0),.clk(gclk));
	jdff dff_A_ZMqnxzvf1_0(.dout(w_dff_A_VmTMOllq2_0),.din(w_dff_A_ZMqnxzvf1_0),.clk(gclk));
	jdff dff_B_B8lF4AdG4_0(.din(n687),.dout(w_dff_B_B8lF4AdG4_0),.clk(gclk));
	jdff dff_B_K7Mb3bCB7_0(.din(w_dff_B_B8lF4AdG4_0),.dout(w_dff_B_K7Mb3bCB7_0),.clk(gclk));
	jdff dff_B_jdHu0q5J0_0(.din(n686),.dout(w_dff_B_jdHu0q5J0_0),.clk(gclk));
	jdff dff_B_Q5u8Ir0H9_0(.din(w_dff_B_jdHu0q5J0_0),.dout(w_dff_B_Q5u8Ir0H9_0),.clk(gclk));
	jdff dff_B_9CjI7fM78_1(.din(n678),.dout(w_dff_B_9CjI7fM78_1),.clk(gclk));
	jdff dff_B_Y0HyG9oT8_1(.din(n679),.dout(w_dff_B_Y0HyG9oT8_1),.clk(gclk));
	jdff dff_A_Y8dPIE7f0_1(.dout(w_n1162_0[1]),.din(w_dff_A_Y8dPIE7f0_1),.clk(gclk));
	jdff dff_A_HGPx0bsZ1_0(.dout(w_G384_0),.din(w_dff_A_HGPx0bsZ1_0),.clk(gclk));
	jdff dff_A_mWJJ95QE5_0(.dout(w_dff_A_HGPx0bsZ1_0),.din(w_dff_A_mWJJ95QE5_0),.clk(gclk));
	jdff dff_A_eHaXs8ak3_2(.dout(w_dff_A_BDdeUnCZ1_0),.din(w_dff_A_eHaXs8ak3_2),.clk(gclk));
	jdff dff_A_BDdeUnCZ1_0(.dout(w_dff_A_OWxnm4cp3_0),.din(w_dff_A_BDdeUnCZ1_0),.clk(gclk));
	jdff dff_A_OWxnm4cp3_0(.dout(w_dff_A_RNsFj8bQ7_0),.din(w_dff_A_OWxnm4cp3_0),.clk(gclk));
	jdff dff_A_RNsFj8bQ7_0(.dout(w_dff_A_ET1kx94Z1_0),.din(w_dff_A_RNsFj8bQ7_0),.clk(gclk));
	jdff dff_A_ET1kx94Z1_0(.dout(w_dff_A_BBwZ4xyJ9_0),.din(w_dff_A_ET1kx94Z1_0),.clk(gclk));
	jdff dff_A_BBwZ4xyJ9_0(.dout(w_dff_A_RX6J1BbH9_0),.din(w_dff_A_BBwZ4xyJ9_0),.clk(gclk));
	jdff dff_A_RX6J1BbH9_0(.dout(w_dff_A_pMt8nEKh0_0),.din(w_dff_A_RX6J1BbH9_0),.clk(gclk));
	jdff dff_A_pMt8nEKh0_0(.dout(w_dff_A_ycarUudx2_0),.din(w_dff_A_pMt8nEKh0_0),.clk(gclk));
	jdff dff_A_ycarUudx2_0(.dout(w_dff_A_kL1Ia3kA9_0),.din(w_dff_A_ycarUudx2_0),.clk(gclk));
	jdff dff_A_kL1Ia3kA9_0(.dout(w_dff_A_wAuMb2Va8_0),.din(w_dff_A_kL1Ia3kA9_0),.clk(gclk));
	jdff dff_A_wAuMb2Va8_0(.dout(w_dff_A_MQ1551cG6_0),.din(w_dff_A_wAuMb2Va8_0),.clk(gclk));
	jdff dff_A_MQ1551cG6_0(.dout(w_dff_A_v8W7uE694_0),.din(w_dff_A_MQ1551cG6_0),.clk(gclk));
	jdff dff_A_v8W7uE694_0(.dout(w_dff_A_9seO9t8D3_0),.din(w_dff_A_v8W7uE694_0),.clk(gclk));
	jdff dff_A_9seO9t8D3_0(.dout(w_dff_A_TUygGutm7_0),.din(w_dff_A_9seO9t8D3_0),.clk(gclk));
	jdff dff_A_TUygGutm7_0(.dout(w_dff_A_p43BVdkF8_0),.din(w_dff_A_TUygGutm7_0),.clk(gclk));
	jdff dff_A_p43BVdkF8_0(.dout(w_dff_A_i0lg6pko8_0),.din(w_dff_A_p43BVdkF8_0),.clk(gclk));
	jdff dff_A_i0lg6pko8_0(.dout(w_dff_A_AwYQKIbY0_0),.din(w_dff_A_i0lg6pko8_0),.clk(gclk));
	jdff dff_A_AwYQKIbY0_0(.dout(w_dff_A_z00g9Up74_0),.din(w_dff_A_AwYQKIbY0_0),.clk(gclk));
	jdff dff_A_z00g9Up74_0(.dout(w_dff_A_rTC27Ujv9_0),.din(w_dff_A_z00g9Up74_0),.clk(gclk));
	jdff dff_A_rTC27Ujv9_0(.dout(w_dff_A_ZuYHJo5F0_0),.din(w_dff_A_rTC27Ujv9_0),.clk(gclk));
	jdff dff_A_ZuYHJo5F0_0(.dout(w_dff_A_XRgZIweo0_0),.din(w_dff_A_ZuYHJo5F0_0),.clk(gclk));
	jdff dff_A_XRgZIweo0_0(.dout(w_dff_A_4iFfzkXn1_0),.din(w_dff_A_XRgZIweo0_0),.clk(gclk));
	jdff dff_A_4iFfzkXn1_0(.dout(w_dff_A_8v7uQRFZ6_0),.din(w_dff_A_4iFfzkXn1_0),.clk(gclk));
	jdff dff_A_8v7uQRFZ6_0(.dout(w_dff_A_PVrdWs1m7_0),.din(w_dff_A_8v7uQRFZ6_0),.clk(gclk));
	jdff dff_A_PVrdWs1m7_0(.dout(G353),.din(w_dff_A_PVrdWs1m7_0),.clk(gclk));
	jdff dff_A_cyNhmvic6_1(.dout(w_dff_A_ya2Aiw553_0),.din(w_dff_A_cyNhmvic6_1),.clk(gclk));
	jdff dff_A_ya2Aiw553_0(.dout(w_dff_A_6Z7j5pSM8_0),.din(w_dff_A_ya2Aiw553_0),.clk(gclk));
	jdff dff_A_6Z7j5pSM8_0(.dout(w_dff_A_DKHdOct33_0),.din(w_dff_A_6Z7j5pSM8_0),.clk(gclk));
	jdff dff_A_DKHdOct33_0(.dout(w_dff_A_iFlNSgwe4_0),.din(w_dff_A_DKHdOct33_0),.clk(gclk));
	jdff dff_A_iFlNSgwe4_0(.dout(w_dff_A_5vnT0x4x4_0),.din(w_dff_A_iFlNSgwe4_0),.clk(gclk));
	jdff dff_A_5vnT0x4x4_0(.dout(w_dff_A_Fwm8XYaE1_0),.din(w_dff_A_5vnT0x4x4_0),.clk(gclk));
	jdff dff_A_Fwm8XYaE1_0(.dout(w_dff_A_rKoB023L2_0),.din(w_dff_A_Fwm8XYaE1_0),.clk(gclk));
	jdff dff_A_rKoB023L2_0(.dout(w_dff_A_MDXAVeua5_0),.din(w_dff_A_rKoB023L2_0),.clk(gclk));
	jdff dff_A_MDXAVeua5_0(.dout(w_dff_A_DBa16L9l0_0),.din(w_dff_A_MDXAVeua5_0),.clk(gclk));
	jdff dff_A_DBa16L9l0_0(.dout(w_dff_A_0fwKqOTm2_0),.din(w_dff_A_DBa16L9l0_0),.clk(gclk));
	jdff dff_A_0fwKqOTm2_0(.dout(w_dff_A_w45RH9sP7_0),.din(w_dff_A_0fwKqOTm2_0),.clk(gclk));
	jdff dff_A_w45RH9sP7_0(.dout(w_dff_A_T55bB0ag8_0),.din(w_dff_A_w45RH9sP7_0),.clk(gclk));
	jdff dff_A_T55bB0ag8_0(.dout(w_dff_A_Gn435XAr0_0),.din(w_dff_A_T55bB0ag8_0),.clk(gclk));
	jdff dff_A_Gn435XAr0_0(.dout(w_dff_A_y1rFtMDE7_0),.din(w_dff_A_Gn435XAr0_0),.clk(gclk));
	jdff dff_A_y1rFtMDE7_0(.dout(w_dff_A_sQMFf0Uv6_0),.din(w_dff_A_y1rFtMDE7_0),.clk(gclk));
	jdff dff_A_sQMFf0Uv6_0(.dout(w_dff_A_y1V3Up6c1_0),.din(w_dff_A_sQMFf0Uv6_0),.clk(gclk));
	jdff dff_A_y1V3Up6c1_0(.dout(w_dff_A_gx07RHvg3_0),.din(w_dff_A_y1V3Up6c1_0),.clk(gclk));
	jdff dff_A_gx07RHvg3_0(.dout(w_dff_A_lDM1FK4F9_0),.din(w_dff_A_gx07RHvg3_0),.clk(gclk));
	jdff dff_A_lDM1FK4F9_0(.dout(w_dff_A_buWJidtA9_0),.din(w_dff_A_lDM1FK4F9_0),.clk(gclk));
	jdff dff_A_buWJidtA9_0(.dout(w_dff_A_xSd0AmbU7_0),.din(w_dff_A_buWJidtA9_0),.clk(gclk));
	jdff dff_A_xSd0AmbU7_0(.dout(w_dff_A_Ua7qVgcQ1_0),.din(w_dff_A_xSd0AmbU7_0),.clk(gclk));
	jdff dff_A_Ua7qVgcQ1_0(.dout(w_dff_A_UDg6dnwl5_0),.din(w_dff_A_Ua7qVgcQ1_0),.clk(gclk));
	jdff dff_A_UDg6dnwl5_0(.dout(w_dff_A_MaMy1aGw3_0),.din(w_dff_A_UDg6dnwl5_0),.clk(gclk));
	jdff dff_A_MaMy1aGw3_0(.dout(G355),.din(w_dff_A_MaMy1aGw3_0),.clk(gclk));
	jdff dff_A_6n9RzDAU9_2(.dout(w_dff_A_iNSP9uw25_0),.din(w_dff_A_6n9RzDAU9_2),.clk(gclk));
	jdff dff_A_iNSP9uw25_0(.dout(w_dff_A_CBPNOo2U9_0),.din(w_dff_A_iNSP9uw25_0),.clk(gclk));
	jdff dff_A_CBPNOo2U9_0(.dout(w_dff_A_JvvWstK53_0),.din(w_dff_A_CBPNOo2U9_0),.clk(gclk));
	jdff dff_A_JvvWstK53_0(.dout(w_dff_A_nzgTBldx3_0),.din(w_dff_A_JvvWstK53_0),.clk(gclk));
	jdff dff_A_nzgTBldx3_0(.dout(w_dff_A_T9L7FZvb1_0),.din(w_dff_A_nzgTBldx3_0),.clk(gclk));
	jdff dff_A_T9L7FZvb1_0(.dout(w_dff_A_xYQy2Xfl7_0),.din(w_dff_A_T9L7FZvb1_0),.clk(gclk));
	jdff dff_A_xYQy2Xfl7_0(.dout(w_dff_A_RFKNx8NZ0_0),.din(w_dff_A_xYQy2Xfl7_0),.clk(gclk));
	jdff dff_A_RFKNx8NZ0_0(.dout(w_dff_A_f9us52zi7_0),.din(w_dff_A_RFKNx8NZ0_0),.clk(gclk));
	jdff dff_A_f9us52zi7_0(.dout(w_dff_A_T9oJ1gxD2_0),.din(w_dff_A_f9us52zi7_0),.clk(gclk));
	jdff dff_A_T9oJ1gxD2_0(.dout(w_dff_A_dBa4KbTK0_0),.din(w_dff_A_T9oJ1gxD2_0),.clk(gclk));
	jdff dff_A_dBa4KbTK0_0(.dout(w_dff_A_MfeAzOyP9_0),.din(w_dff_A_dBa4KbTK0_0),.clk(gclk));
	jdff dff_A_MfeAzOyP9_0(.dout(w_dff_A_vkpN7A7S9_0),.din(w_dff_A_MfeAzOyP9_0),.clk(gclk));
	jdff dff_A_vkpN7A7S9_0(.dout(w_dff_A_9FzQSQQg7_0),.din(w_dff_A_vkpN7A7S9_0),.clk(gclk));
	jdff dff_A_9FzQSQQg7_0(.dout(w_dff_A_vDuzeeR05_0),.din(w_dff_A_9FzQSQQg7_0),.clk(gclk));
	jdff dff_A_vDuzeeR05_0(.dout(w_dff_A_PZ8IaZCk7_0),.din(w_dff_A_vDuzeeR05_0),.clk(gclk));
	jdff dff_A_PZ8IaZCk7_0(.dout(w_dff_A_eCwCsQfR5_0),.din(w_dff_A_PZ8IaZCk7_0),.clk(gclk));
	jdff dff_A_eCwCsQfR5_0(.dout(w_dff_A_SoS4AyFT1_0),.din(w_dff_A_eCwCsQfR5_0),.clk(gclk));
	jdff dff_A_SoS4AyFT1_0(.dout(w_dff_A_mtE2qBZj4_0),.din(w_dff_A_SoS4AyFT1_0),.clk(gclk));
	jdff dff_A_mtE2qBZj4_0(.dout(w_dff_A_L3dAmn8P4_0),.din(w_dff_A_mtE2qBZj4_0),.clk(gclk));
	jdff dff_A_L3dAmn8P4_0(.dout(w_dff_A_NF138Mhz6_0),.din(w_dff_A_L3dAmn8P4_0),.clk(gclk));
	jdff dff_A_NF138Mhz6_0(.dout(G361),.din(w_dff_A_NF138Mhz6_0),.clk(gclk));
	jdff dff_A_x8w3OkNr6_2(.dout(w_dff_A_t3WM7HnJ4_0),.din(w_dff_A_x8w3OkNr6_2),.clk(gclk));
	jdff dff_A_t3WM7HnJ4_0(.dout(w_dff_A_fmUKup6j7_0),.din(w_dff_A_t3WM7HnJ4_0),.clk(gclk));
	jdff dff_A_fmUKup6j7_0(.dout(w_dff_A_Iib65AKQ2_0),.din(w_dff_A_fmUKup6j7_0),.clk(gclk));
	jdff dff_A_Iib65AKQ2_0(.dout(w_dff_A_PH8Lw6Nm5_0),.din(w_dff_A_Iib65AKQ2_0),.clk(gclk));
	jdff dff_A_PH8Lw6Nm5_0(.dout(w_dff_A_nQlaNGRY6_0),.din(w_dff_A_PH8Lw6Nm5_0),.clk(gclk));
	jdff dff_A_nQlaNGRY6_0(.dout(w_dff_A_tBFinChI6_0),.din(w_dff_A_nQlaNGRY6_0),.clk(gclk));
	jdff dff_A_tBFinChI6_0(.dout(w_dff_A_SnGa4QSV0_0),.din(w_dff_A_tBFinChI6_0),.clk(gclk));
	jdff dff_A_SnGa4QSV0_0(.dout(w_dff_A_Z7a0zdQI7_0),.din(w_dff_A_SnGa4QSV0_0),.clk(gclk));
	jdff dff_A_Z7a0zdQI7_0(.dout(w_dff_A_JKlPqns47_0),.din(w_dff_A_Z7a0zdQI7_0),.clk(gclk));
	jdff dff_A_JKlPqns47_0(.dout(w_dff_A_NPlDhGk86_0),.din(w_dff_A_JKlPqns47_0),.clk(gclk));
	jdff dff_A_NPlDhGk86_0(.dout(w_dff_A_Z5CYrWyN0_0),.din(w_dff_A_NPlDhGk86_0),.clk(gclk));
	jdff dff_A_Z5CYrWyN0_0(.dout(w_dff_A_o63knkld1_0),.din(w_dff_A_Z5CYrWyN0_0),.clk(gclk));
	jdff dff_A_o63knkld1_0(.dout(w_dff_A_OeGHYLmr5_0),.din(w_dff_A_o63knkld1_0),.clk(gclk));
	jdff dff_A_OeGHYLmr5_0(.dout(w_dff_A_EVSH4rOi8_0),.din(w_dff_A_OeGHYLmr5_0),.clk(gclk));
	jdff dff_A_EVSH4rOi8_0(.dout(w_dff_A_WG0SuF1k2_0),.din(w_dff_A_EVSH4rOi8_0),.clk(gclk));
	jdff dff_A_WG0SuF1k2_0(.dout(w_dff_A_4pK8wCXV0_0),.din(w_dff_A_WG0SuF1k2_0),.clk(gclk));
	jdff dff_A_4pK8wCXV0_0(.dout(w_dff_A_e7ox6w9F9_0),.din(w_dff_A_4pK8wCXV0_0),.clk(gclk));
	jdff dff_A_e7ox6w9F9_0(.dout(w_dff_A_Z0c9FQ7z3_0),.din(w_dff_A_e7ox6w9F9_0),.clk(gclk));
	jdff dff_A_Z0c9FQ7z3_0(.dout(w_dff_A_mPX9ATHL6_0),.din(w_dff_A_Z0c9FQ7z3_0),.clk(gclk));
	jdff dff_A_mPX9ATHL6_0(.dout(w_dff_A_hc8aJAzE8_0),.din(w_dff_A_mPX9ATHL6_0),.clk(gclk));
	jdff dff_A_hc8aJAzE8_0(.dout(w_dff_A_g5PN8qbD9_0),.din(w_dff_A_hc8aJAzE8_0),.clk(gclk));
	jdff dff_A_g5PN8qbD9_0(.dout(w_dff_A_S97nMcH87_0),.din(w_dff_A_g5PN8qbD9_0),.clk(gclk));
	jdff dff_A_S97nMcH87_0(.dout(w_dff_A_2CuGPe2C3_0),.din(w_dff_A_S97nMcH87_0),.clk(gclk));
	jdff dff_A_2CuGPe2C3_0(.dout(G358),.din(w_dff_A_2CuGPe2C3_0),.clk(gclk));
	jdff dff_A_MMM98mI96_2(.dout(w_dff_A_YrGIIctL5_0),.din(w_dff_A_MMM98mI96_2),.clk(gclk));
	jdff dff_A_YrGIIctL5_0(.dout(w_dff_A_orUO2Ost2_0),.din(w_dff_A_YrGIIctL5_0),.clk(gclk));
	jdff dff_A_orUO2Ost2_0(.dout(w_dff_A_YdwBZwp39_0),.din(w_dff_A_orUO2Ost2_0),.clk(gclk));
	jdff dff_A_YdwBZwp39_0(.dout(w_dff_A_OZFTCYku7_0),.din(w_dff_A_YdwBZwp39_0),.clk(gclk));
	jdff dff_A_OZFTCYku7_0(.dout(w_dff_A_cssR2C1c8_0),.din(w_dff_A_OZFTCYku7_0),.clk(gclk));
	jdff dff_A_cssR2C1c8_0(.dout(w_dff_A_FfGxyauN6_0),.din(w_dff_A_cssR2C1c8_0),.clk(gclk));
	jdff dff_A_FfGxyauN6_0(.dout(w_dff_A_53HRLule7_0),.din(w_dff_A_FfGxyauN6_0),.clk(gclk));
	jdff dff_A_53HRLule7_0(.dout(w_dff_A_o12pm6UI9_0),.din(w_dff_A_53HRLule7_0),.clk(gclk));
	jdff dff_A_o12pm6UI9_0(.dout(w_dff_A_PqmNOBEM2_0),.din(w_dff_A_o12pm6UI9_0),.clk(gclk));
	jdff dff_A_PqmNOBEM2_0(.dout(w_dff_A_ThQHPZvC2_0),.din(w_dff_A_PqmNOBEM2_0),.clk(gclk));
	jdff dff_A_ThQHPZvC2_0(.dout(w_dff_A_ko0gb4Uk0_0),.din(w_dff_A_ThQHPZvC2_0),.clk(gclk));
	jdff dff_A_ko0gb4Uk0_0(.dout(w_dff_A_SSBgdHsN2_0),.din(w_dff_A_ko0gb4Uk0_0),.clk(gclk));
	jdff dff_A_SSBgdHsN2_0(.dout(w_dff_A_NkCpB6At9_0),.din(w_dff_A_SSBgdHsN2_0),.clk(gclk));
	jdff dff_A_NkCpB6At9_0(.dout(w_dff_A_I3XUg78F4_0),.din(w_dff_A_NkCpB6At9_0),.clk(gclk));
	jdff dff_A_I3XUg78F4_0(.dout(w_dff_A_csKpg7Vr3_0),.din(w_dff_A_I3XUg78F4_0),.clk(gclk));
	jdff dff_A_csKpg7Vr3_0(.dout(w_dff_A_8PAszGGU4_0),.din(w_dff_A_csKpg7Vr3_0),.clk(gclk));
	jdff dff_A_8PAszGGU4_0(.dout(w_dff_A_69Tfxs4k6_0),.din(w_dff_A_8PAszGGU4_0),.clk(gclk));
	jdff dff_A_69Tfxs4k6_0(.dout(w_dff_A_AG6pyT1G1_0),.din(w_dff_A_69Tfxs4k6_0),.clk(gclk));
	jdff dff_A_AG6pyT1G1_0(.dout(w_dff_A_XrDOxc951_0),.din(w_dff_A_AG6pyT1G1_0),.clk(gclk));
	jdff dff_A_XrDOxc951_0(.dout(w_dff_A_qOIsBatc1_0),.din(w_dff_A_XrDOxc951_0),.clk(gclk));
	jdff dff_A_qOIsBatc1_0(.dout(w_dff_A_zxLaVc240_0),.din(w_dff_A_qOIsBatc1_0),.clk(gclk));
	jdff dff_A_zxLaVc240_0(.dout(w_dff_A_CwuYsNzx1_0),.din(w_dff_A_zxLaVc240_0),.clk(gclk));
	jdff dff_A_CwuYsNzx1_0(.dout(w_dff_A_rBcBKz039_0),.din(w_dff_A_CwuYsNzx1_0),.clk(gclk));
	jdff dff_A_rBcBKz039_0(.dout(G351),.din(w_dff_A_rBcBKz039_0),.clk(gclk));
	jdff dff_A_pVqNiwPA5_2(.dout(w_dff_A_TPRssbmc8_0),.din(w_dff_A_pVqNiwPA5_2),.clk(gclk));
	jdff dff_A_TPRssbmc8_0(.dout(w_dff_A_s5w8MOP58_0),.din(w_dff_A_TPRssbmc8_0),.clk(gclk));
	jdff dff_A_s5w8MOP58_0(.dout(w_dff_A_ImsFZWhO1_0),.din(w_dff_A_s5w8MOP58_0),.clk(gclk));
	jdff dff_A_ImsFZWhO1_0(.dout(w_dff_A_qMgARpnT2_0),.din(w_dff_A_ImsFZWhO1_0),.clk(gclk));
	jdff dff_A_qMgARpnT2_0(.dout(w_dff_A_eTu77bM78_0),.din(w_dff_A_qMgARpnT2_0),.clk(gclk));
	jdff dff_A_eTu77bM78_0(.dout(w_dff_A_011DCSol9_0),.din(w_dff_A_eTu77bM78_0),.clk(gclk));
	jdff dff_A_011DCSol9_0(.dout(w_dff_A_gx0RmkDW7_0),.din(w_dff_A_011DCSol9_0),.clk(gclk));
	jdff dff_A_gx0RmkDW7_0(.dout(w_dff_A_EOnlBFNd4_0),.din(w_dff_A_gx0RmkDW7_0),.clk(gclk));
	jdff dff_A_EOnlBFNd4_0(.dout(w_dff_A_1BfvGWRs3_0),.din(w_dff_A_EOnlBFNd4_0),.clk(gclk));
	jdff dff_A_1BfvGWRs3_0(.dout(w_dff_A_OPG2z6hB5_0),.din(w_dff_A_1BfvGWRs3_0),.clk(gclk));
	jdff dff_A_OPG2z6hB5_0(.dout(w_dff_A_6vdob3ul3_0),.din(w_dff_A_OPG2z6hB5_0),.clk(gclk));
	jdff dff_A_6vdob3ul3_0(.dout(w_dff_A_pfdSVIcz9_0),.din(w_dff_A_6vdob3ul3_0),.clk(gclk));
	jdff dff_A_pfdSVIcz9_0(.dout(w_dff_A_O4NSYRy27_0),.din(w_dff_A_pfdSVIcz9_0),.clk(gclk));
	jdff dff_A_O4NSYRy27_0(.dout(G372),.din(w_dff_A_O4NSYRy27_0),.clk(gclk));
	jdff dff_A_m84hN0bh5_2(.dout(w_dff_A_6UGpNuVA1_0),.din(w_dff_A_m84hN0bh5_2),.clk(gclk));
	jdff dff_A_6UGpNuVA1_0(.dout(w_dff_A_dM8FEHoY5_0),.din(w_dff_A_6UGpNuVA1_0),.clk(gclk));
	jdff dff_A_dM8FEHoY5_0(.dout(w_dff_A_ZPtrLbS69_0),.din(w_dff_A_dM8FEHoY5_0),.clk(gclk));
	jdff dff_A_ZPtrLbS69_0(.dout(w_dff_A_uF27NlyY1_0),.din(w_dff_A_ZPtrLbS69_0),.clk(gclk));
	jdff dff_A_uF27NlyY1_0(.dout(w_dff_A_ALf8UQqd3_0),.din(w_dff_A_uF27NlyY1_0),.clk(gclk));
	jdff dff_A_ALf8UQqd3_0(.dout(w_dff_A_U65q1uSE1_0),.din(w_dff_A_ALf8UQqd3_0),.clk(gclk));
	jdff dff_A_U65q1uSE1_0(.dout(w_dff_A_BRMIDGBu3_0),.din(w_dff_A_U65q1uSE1_0),.clk(gclk));
	jdff dff_A_BRMIDGBu3_0(.dout(w_dff_A_qlaIbqXv0_0),.din(w_dff_A_BRMIDGBu3_0),.clk(gclk));
	jdff dff_A_qlaIbqXv0_0(.dout(w_dff_A_EDn6K2rB2_0),.din(w_dff_A_qlaIbqXv0_0),.clk(gclk));
	jdff dff_A_EDn6K2rB2_0(.dout(w_dff_A_dV9SLUXR1_0),.din(w_dff_A_EDn6K2rB2_0),.clk(gclk));
	jdff dff_A_dV9SLUXR1_0(.dout(w_dff_A_zAvXALRF6_0),.din(w_dff_A_dV9SLUXR1_0),.clk(gclk));
	jdff dff_A_zAvXALRF6_0(.dout(G369),.din(w_dff_A_zAvXALRF6_0),.clk(gclk));
	jdff dff_A_m8XhH8tq7_2(.dout(w_dff_A_m9IwkISh1_0),.din(w_dff_A_m8XhH8tq7_2),.clk(gclk));
	jdff dff_A_m9IwkISh1_0(.dout(w_dff_A_qzfDZh0X6_0),.din(w_dff_A_m9IwkISh1_0),.clk(gclk));
	jdff dff_A_qzfDZh0X6_0(.dout(w_dff_A_cm4dQeg76_0),.din(w_dff_A_qzfDZh0X6_0),.clk(gclk));
	jdff dff_A_cm4dQeg76_0(.dout(w_dff_A_hksdxLHH8_0),.din(w_dff_A_cm4dQeg76_0),.clk(gclk));
	jdff dff_A_hksdxLHH8_0(.dout(w_dff_A_hzpk3Q5F4_0),.din(w_dff_A_hksdxLHH8_0),.clk(gclk));
	jdff dff_A_hzpk3Q5F4_0(.dout(w_dff_A_OSBCI5aM6_0),.din(w_dff_A_hzpk3Q5F4_0),.clk(gclk));
	jdff dff_A_OSBCI5aM6_0(.dout(w_dff_A_qMmPkybN2_0),.din(w_dff_A_OSBCI5aM6_0),.clk(gclk));
	jdff dff_A_qMmPkybN2_0(.dout(w_dff_A_c020QNlg6_0),.din(w_dff_A_qMmPkybN2_0),.clk(gclk));
	jdff dff_A_c020QNlg6_0(.dout(w_dff_A_roHWtaR75_0),.din(w_dff_A_c020QNlg6_0),.clk(gclk));
	jdff dff_A_roHWtaR75_0(.dout(w_dff_A_5113JSsV7_0),.din(w_dff_A_roHWtaR75_0),.clk(gclk));
	jdff dff_A_5113JSsV7_0(.dout(G399),.din(w_dff_A_5113JSsV7_0),.clk(gclk));
	jdff dff_A_suxkJc9W4_2(.dout(w_dff_A_Z8JREjjN9_0),.din(w_dff_A_suxkJc9W4_2),.clk(gclk));
	jdff dff_A_Z8JREjjN9_0(.dout(w_dff_A_7pgYwA4l1_0),.din(w_dff_A_Z8JREjjN9_0),.clk(gclk));
	jdff dff_A_7pgYwA4l1_0(.dout(w_dff_A_0FQj6WAO3_0),.din(w_dff_A_7pgYwA4l1_0),.clk(gclk));
	jdff dff_A_0FQj6WAO3_0(.dout(w_dff_A_ofbc0hAk3_0),.din(w_dff_A_0FQj6WAO3_0),.clk(gclk));
	jdff dff_A_ofbc0hAk3_0(.dout(w_dff_A_76SFJWpT8_0),.din(w_dff_A_ofbc0hAk3_0),.clk(gclk));
	jdff dff_A_76SFJWpT8_0(.dout(w_dff_A_3yh6VbIy4_0),.din(w_dff_A_76SFJWpT8_0),.clk(gclk));
	jdff dff_A_3yh6VbIy4_0(.dout(w_dff_A_YA1W9wn41_0),.din(w_dff_A_3yh6VbIy4_0),.clk(gclk));
	jdff dff_A_YA1W9wn41_0(.dout(w_dff_A_OJoT2UhP0_0),.din(w_dff_A_YA1W9wn41_0),.clk(gclk));
	jdff dff_A_OJoT2UhP0_0(.dout(w_dff_A_lgEufWyi0_0),.din(w_dff_A_OJoT2UhP0_0),.clk(gclk));
	jdff dff_A_lgEufWyi0_0(.dout(w_dff_A_FH1rm7wP5_0),.din(w_dff_A_lgEufWyi0_0),.clk(gclk));
	jdff dff_A_FH1rm7wP5_0(.dout(G364),.din(w_dff_A_FH1rm7wP5_0),.clk(gclk));
	jdff dff_A_QVGVQfYK5_2(.dout(w_dff_A_pO225CQ91_0),.din(w_dff_A_QVGVQfYK5_2),.clk(gclk));
	jdff dff_A_pO225CQ91_0(.dout(w_dff_A_pM3r58Os8_0),.din(w_dff_A_pO225CQ91_0),.clk(gclk));
	jdff dff_A_pM3r58Os8_0(.dout(w_dff_A_XQxYVzmv4_0),.din(w_dff_A_pM3r58Os8_0),.clk(gclk));
	jdff dff_A_XQxYVzmv4_0(.dout(w_dff_A_ZkoGnkeN7_0),.din(w_dff_A_XQxYVzmv4_0),.clk(gclk));
	jdff dff_A_ZkoGnkeN7_0(.dout(w_dff_A_8yzMmy9m2_0),.din(w_dff_A_ZkoGnkeN7_0),.clk(gclk));
	jdff dff_A_8yzMmy9m2_0(.dout(w_dff_A_37tdttyl5_0),.din(w_dff_A_8yzMmy9m2_0),.clk(gclk));
	jdff dff_A_37tdttyl5_0(.dout(w_dff_A_TBeJSWGG1_0),.din(w_dff_A_37tdttyl5_0),.clk(gclk));
	jdff dff_A_TBeJSWGG1_0(.dout(w_dff_A_5THm0ccg7_0),.din(w_dff_A_TBeJSWGG1_0),.clk(gclk));
	jdff dff_A_5THm0ccg7_0(.dout(w_dff_A_3mqd2LSB1_0),.din(w_dff_A_5THm0ccg7_0),.clk(gclk));
	jdff dff_A_3mqd2LSB1_0(.dout(w_dff_A_TTs0Ebo48_0),.din(w_dff_A_3mqd2LSB1_0),.clk(gclk));
	jdff dff_A_TTs0Ebo48_0(.dout(G396),.din(w_dff_A_TTs0Ebo48_0),.clk(gclk));
	jdff dff_A_CAs6wypP0_1(.dout(w_dff_A_04yIwS3a1_0),.din(w_dff_A_CAs6wypP0_1),.clk(gclk));
	jdff dff_A_04yIwS3a1_0(.dout(w_dff_A_xjM1qNsL6_0),.din(w_dff_A_04yIwS3a1_0),.clk(gclk));
	jdff dff_A_xjM1qNsL6_0(.dout(w_dff_A_Y0gcCkcp8_0),.din(w_dff_A_xjM1qNsL6_0),.clk(gclk));
	jdff dff_A_Y0gcCkcp8_0(.dout(w_dff_A_RDkaEOis8_0),.din(w_dff_A_Y0gcCkcp8_0),.clk(gclk));
	jdff dff_A_RDkaEOis8_0(.dout(w_dff_A_Z6Sxk4LA1_0),.din(w_dff_A_RDkaEOis8_0),.clk(gclk));
	jdff dff_A_Z6Sxk4LA1_0(.dout(w_dff_A_zSE96s8W0_0),.din(w_dff_A_Z6Sxk4LA1_0),.clk(gclk));
	jdff dff_A_zSE96s8W0_0(.dout(w_dff_A_J1Db1Fso2_0),.din(w_dff_A_zSE96s8W0_0),.clk(gclk));
	jdff dff_A_J1Db1Fso2_0(.dout(G384),.din(w_dff_A_J1Db1Fso2_0),.clk(gclk));
	jdff dff_A_8Faaqfu06_2(.dout(w_dff_A_fgvTXq5c7_0),.din(w_dff_A_8Faaqfu06_2),.clk(gclk));
	jdff dff_A_fgvTXq5c7_0(.dout(w_dff_A_SqT9QFom1_0),.din(w_dff_A_fgvTXq5c7_0),.clk(gclk));
	jdff dff_A_SqT9QFom1_0(.dout(w_dff_A_VQjg5Bf97_0),.din(w_dff_A_SqT9QFom1_0),.clk(gclk));
	jdff dff_A_VQjg5Bf97_0(.dout(w_dff_A_uvV2URYd5_0),.din(w_dff_A_VQjg5Bf97_0),.clk(gclk));
	jdff dff_A_uvV2URYd5_0(.dout(G367),.din(w_dff_A_uvV2URYd5_0),.clk(gclk));
	jdff dff_A_iCSTSP0S7_2(.dout(w_dff_A_pbvNBtfW3_0),.din(w_dff_A_iCSTSP0S7_2),.clk(gclk));
	jdff dff_A_pbvNBtfW3_0(.dout(w_dff_A_j05d5K929_0),.din(w_dff_A_pbvNBtfW3_0),.clk(gclk));
	jdff dff_A_j05d5K929_0(.dout(w_dff_A_CYRV8SvA9_0),.din(w_dff_A_j05d5K929_0),.clk(gclk));
	jdff dff_A_CYRV8SvA9_0(.dout(w_dff_A_RTDFHfRV3_0),.din(w_dff_A_CYRV8SvA9_0),.clk(gclk));
	jdff dff_A_RTDFHfRV3_0(.dout(G387),.din(w_dff_A_RTDFHfRV3_0),.clk(gclk));
	jdff dff_A_QIL9dh5f4_1(.dout(w_dff_A_Pc7m9k791_0),.din(w_dff_A_QIL9dh5f4_1),.clk(gclk));
	jdff dff_A_Pc7m9k791_0(.dout(w_dff_A_uwKuCJ2R9_0),.din(w_dff_A_Pc7m9k791_0),.clk(gclk));
	jdff dff_A_uwKuCJ2R9_0(.dout(w_dff_A_Z3X71WYa8_0),.din(w_dff_A_uwKuCJ2R9_0),.clk(gclk));
	jdff dff_A_Z3X71WYa8_0(.dout(w_dff_A_tzjOiDPM2_0),.din(w_dff_A_Z3X71WYa8_0),.clk(gclk));
	jdff dff_A_tzjOiDPM2_0(.dout(w_dff_A_TX9cKArf8_0),.din(w_dff_A_tzjOiDPM2_0),.clk(gclk));
	jdff dff_A_TX9cKArf8_0(.dout(w_dff_A_yJeu9qUG8_0),.din(w_dff_A_TX9cKArf8_0),.clk(gclk));
	jdff dff_A_yJeu9qUG8_0(.dout(G393),.din(w_dff_A_yJeu9qUG8_0),.clk(gclk));
	jdff dff_A_C8WizjaC4_1(.dout(w_dff_A_W8ZDHHB99_0),.din(w_dff_A_C8WizjaC4_1),.clk(gclk));
	jdff dff_A_W8ZDHHB99_0(.dout(w_dff_A_zxDUn9Pe6_0),.din(w_dff_A_W8ZDHHB99_0),.clk(gclk));
	jdff dff_A_zxDUn9Pe6_0(.dout(w_dff_A_jF25fous3_0),.din(w_dff_A_zxDUn9Pe6_0),.clk(gclk));
	jdff dff_A_jF25fous3_0(.dout(w_dff_A_cWd8y1Eo7_0),.din(w_dff_A_jF25fous3_0),.clk(gclk));
	jdff dff_A_cWd8y1Eo7_0(.dout(w_dff_A_x6MFrcXs1_0),.din(w_dff_A_cWd8y1Eo7_0),.clk(gclk));
	jdff dff_A_x6MFrcXs1_0(.dout(G390),.din(w_dff_A_x6MFrcXs1_0),.clk(gclk));
	jdff dff_A_4BLq7DIM7_1(.dout(w_dff_A_L9dsrKyh3_0),.din(w_dff_A_4BLq7DIM7_1),.clk(gclk));
	jdff dff_A_L9dsrKyh3_0(.dout(w_dff_A_a5H6vCKM6_0),.din(w_dff_A_L9dsrKyh3_0),.clk(gclk));
	jdff dff_A_a5H6vCKM6_0(.dout(w_dff_A_eJfTlNBL5_0),.din(w_dff_A_a5H6vCKM6_0),.clk(gclk));
	jdff dff_A_eJfTlNBL5_0(.dout(w_dff_A_mUQgB1iF3_0),.din(w_dff_A_eJfTlNBL5_0),.clk(gclk));
	jdff dff_A_mUQgB1iF3_0(.dout(G378),.din(w_dff_A_mUQgB1iF3_0),.clk(gclk));
	jdff dff_A_Kdmz1GUI9_1(.dout(w_dff_A_uVGAMC2O8_0),.din(w_dff_A_Kdmz1GUI9_1),.clk(gclk));
	jdff dff_A_uVGAMC2O8_0(.dout(w_dff_A_rTlkI1I64_0),.din(w_dff_A_uVGAMC2O8_0),.clk(gclk));
	jdff dff_A_rTlkI1I64_0(.dout(G375),.din(w_dff_A_rTlkI1I64_0),.clk(gclk));
	jdff dff_A_3TPEWlaZ5_1(.dout(w_dff_A_OpvJBNVA6_0),.din(w_dff_A_3TPEWlaZ5_1),.clk(gclk));
	jdff dff_A_OpvJBNVA6_0(.dout(w_dff_A_wVG6D6Ml7_0),.din(w_dff_A_OpvJBNVA6_0),.clk(gclk));
	jdff dff_A_wVG6D6Ml7_0(.dout(w_dff_A_PVlWremV5_0),.din(w_dff_A_wVG6D6Ml7_0),.clk(gclk));
	jdff dff_A_PVlWremV5_0(.dout(w_dff_A_5wTVWcMF7_0),.din(w_dff_A_PVlWremV5_0),.clk(gclk));
	jdff dff_A_5wTVWcMF7_0(.dout(G381),.din(w_dff_A_5wTVWcMF7_0),.clk(gclk));
	jdff dff_A_snNc0Gbh4_1(.dout(G407),.din(w_dff_A_snNc0Gbh4_1),.clk(gclk));
	jdff dff_A_Znbnrzrt0_2(.dout(G402),.din(w_dff_A_Znbnrzrt0_2),.clk(gclk));
endmodule

