/*
rf_c5315:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 4692
	jand: 605
	jor: 419

Summary:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 4692
	jand: 605
	jor: 419

The maximum logic level gap of any gate:
	rf_c5315: 21
*/

module rf_c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1157;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G4_0;
	wire [1:0] w_G4_1;
	wire [1:0] w_G11_0;
	wire [1:0] w_G14_0;
	wire [1:0] w_G17_0;
	wire [1:0] w_G20_0;
	wire [1:0] w_G37_0;
	wire [1:0] w_G40_0;
	wire [1:0] w_G43_0;
	wire [1:0] w_G46_0;
	wire [1:0] w_G49_0;
	wire [1:0] w_G54_0;
	wire [1:0] w_G61_0;
	wire [1:0] w_G64_0;
	wire [1:0] w_G67_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G73_0;
	wire [1:0] w_G76_0;
	wire [1:0] w_G91_0;
	wire [1:0] w_G100_0;
	wire [1:0] w_G103_0;
	wire [1:0] w_G106_0;
	wire [1:0] w_G109_0;
	wire [1:0] w_G123_0;
	wire [1:0] w_G132_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G137_2;
	wire [2:0] w_G137_3;
	wire [2:0] w_G137_4;
	wire [2:0] w_G137_5;
	wire [2:0] w_G137_6;
	wire [2:0] w_G137_7;
	wire [2:0] w_G137_8;
	wire [1:0] w_G137_9;
	wire [2:0] w_G141_0;
	wire [2:0] w_G141_1;
	wire [2:0] w_G141_2;
	wire [1:0] w_G146_0;
	wire [1:0] w_G149_0;
	wire [1:0] w_G152_0;
	wire [1:0] w_G155_0;
	wire [1:0] w_G158_0;
	wire [1:0] w_G161_0;
	wire [1:0] w_G164_0;
	wire [1:0] w_G167_0;
	wire [1:0] w_G170_0;
	wire [1:0] w_G173_0;
	wire [1:0] w_G182_0;
	wire [1:0] w_G185_0;
	wire [1:0] w_G188_0;
	wire [1:0] w_G191_0;
	wire [1:0] w_G194_0;
	wire [1:0] w_G197_0;
	wire [1:0] w_G200_0;
	wire [1:0] w_G203_0;
	wire [2:0] w_G206_0;
	wire [2:0] w_G210_0;
	wire [2:0] w_G210_1;
	wire [2:0] w_G210_2;
	wire [2:0] w_G218_0;
	wire [2:0] w_G218_1;
	wire [2:0] w_G218_2;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [2:0] w_G226_2;
	wire [2:0] w_G234_0;
	wire [2:0] w_G234_1;
	wire [1:0] w_G234_2;
	wire [2:0] w_G242_0;
	wire [2:0] w_G242_1;
	wire [1:0] w_G245_0;
	wire [2:0] w_G248_0;
	wire [2:0] w_G248_1;
	wire [2:0] w_G248_2;
	wire [2:0] w_G248_3;
	wire [2:0] w_G248_4;
	wire [1:0] w_G248_5;
	wire [2:0] w_G251_0;
	wire [2:0] w_G251_1;
	wire [2:0] w_G251_2;
	wire [2:0] w_G251_3;
	wire [2:0] w_G251_4;
	wire [2:0] w_G254_0;
	wire [2:0] w_G254_1;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G257_2;
	wire [2:0] w_G265_0;
	wire [2:0] w_G265_1;
	wire [1:0] w_G265_2;
	wire [2:0] w_G273_0;
	wire [2:0] w_G273_1;
	wire [2:0] w_G273_2;
	wire [1:0] w_G280_0;
	wire [2:0] w_G281_0;
	wire [2:0] w_G281_1;
	wire [1:0] w_G281_2;
	wire [1:0] w_G289_0;
	wire [2:0] w_G293_0;
	wire [2:0] w_G299_0;
	wire [2:0] w_G302_0;
	wire [2:0] w_G308_0;
	wire [2:0] w_G308_1;
	wire [2:0] w_G316_0;
	wire [2:0] w_G316_1;
	wire [2:0] w_G324_0;
	wire [2:0] w_G324_1;
	wire [1:0] w_G331_0;
	wire [2:0] w_G332_0;
	wire [2:0] w_G332_1;
	wire [2:0] w_G332_2;
	wire [2:0] w_G332_3;
	wire [2:0] w_G332_4;
	wire [2:0] w_G335_0;
	wire [2:0] w_G335_1;
	wire [2:0] w_G335_2;
	wire [2:0] w_G335_3;
	wire [1:0] w_G335_4;
	wire [2:0] w_G341_0;
	wire [2:0] w_G341_1;
	wire [2:0] w_G341_2;
	wire [1:0] w_G348_0;
	wire [2:0] w_G351_0;
	wire [2:0] w_G351_1;
	wire [2:0] w_G351_2;
	wire [1:0] w_G358_0;
	wire [2:0] w_G361_0;
	wire [1:0] w_G369_0;
	wire [2:0] w_G374_0;
	wire [2:0] w_G389_0;
	wire [2:0] w_G400_0;
	wire [1:0] w_G400_1;
	wire [2:0] w_G411_0;
	wire [2:0] w_G422_0;
	wire [2:0] w_G422_1;
	wire [1:0] w_G422_2;
	wire [2:0] w_G435_0;
	wire [2:0] w_G435_1;
	wire [2:0] w_G446_0;
	wire [2:0] w_G446_1;
	wire [2:0] w_G457_0;
	wire [2:0] w_G457_1;
	wire [1:0] w_G457_2;
	wire [2:0] w_G468_0;
	wire [2:0] w_G468_1;
	wire [2:0] w_G479_0;
	wire [1:0] w_G479_1;
	wire [2:0] w_G490_0;
	wire [2:0] w_G490_1;
	wire [2:0] w_G503_0;
	wire [2:0] w_G503_1;
	wire [2:0] w_G514_0;
	wire [1:0] w_G514_1;
	wire [2:0] w_G523_0;
	wire [1:0] w_G523_1;
	wire [2:0] w_G534_0;
	wire [2:0] w_G534_1;
	wire [2:0] w_G545_0;
	wire [2:0] w_G549_0;
	wire [1:0] w_G552_0;
	wire [1:0] w_G559_0;
	wire [1:0] w_G562_0;
	wire [2:0] w_G1497_0;
	wire [2:0] w_G1689_0;
	wire [2:0] w_G1690_0;
	wire [2:0] w_G1691_0;
	wire [2:0] w_G1694_0;
	wire [2:0] w_G2174_0;
	wire [2:0] w_G2358_0;
	wire [2:0] w_G2358_1;
	wire [2:0] w_G2358_2;
	wire [1:0] w_G3173_0;
	wire [2:0] w_G3546_0;
	wire [2:0] w_G3546_1;
	wire [2:0] w_G3546_2;
	wire [2:0] w_G3546_3;
	wire [2:0] w_G3546_4;
	wire [1:0] w_G3546_5;
	wire [2:0] w_G3548_0;
	wire [2:0] w_G3548_1;
	wire [2:0] w_G3548_2;
	wire [2:0] w_G3548_3;
	wire [2:0] w_G3548_4;
	wire [1:0] w_G3552_0;
	wire [1:0] w_G3717_0;
	wire [2:0] w_G3724_0;
	wire [2:0] w_G4087_0;
	wire [2:0] w_G4088_0;
	wire [2:0] w_G4089_0;
	wire [2:0] w_G4090_0;
	wire [2:0] w_G4091_0;
	wire [2:0] w_G4091_1;
	wire [2:0] w_G4091_2;
	wire [2:0] w_G4092_0;
	wire [2:0] w_G4092_1;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G600_0;
	wire G600_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G611_0;
	wire G611_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire [2:0] w_G809_0;
	wire [2:0] w_G809_1;
	wire [2:0] w_G809_2;
	wire [1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G1000_0;
	wire G1000_fa_;
	wire w_G826_0;
	wire G826_fa_;
	wire w_G828_0;
	wire G828_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G867_0;
	wire G867_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [2:0] w_n326_0;
	wire [2:0] w_n326_1;
	wire [1:0] w_n326_2;
	wire [1:0] w_n333_0;
	wire [1:0] w_n336_0;
	wire [1:0] w_n360_0;
	wire [1:0] w_n362_0;
	wire [2:0] w_n366_0;
	wire [2:0] w_n366_1;
	wire [2:0] w_n366_2;
	wire [2:0] w_n366_3;
	wire [2:0] w_n366_4;
	wire [2:0] w_n368_0;
	wire [2:0] w_n368_1;
	wire [2:0] w_n368_2;
	wire [2:0] w_n368_3;
	wire [2:0] w_n368_4;
	wire [1:0] w_n368_5;
	wire [2:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n385_0;
	wire [2:0] w_n385_1;
	wire [2:0] w_n386_0;
	wire [2:0] w_n386_1;
	wire [2:0] w_n386_2;
	wire [2:0] w_n386_3;
	wire [2:0] w_n386_4;
	wire [2:0] w_n388_0;
	wire [2:0] w_n388_1;
	wire [2:0] w_n389_0;
	wire [2:0] w_n389_1;
	wire [2:0] w_n389_2;
	wire [2:0] w_n389_3;
	wire [2:0] w_n389_4;
	wire [1:0] w_n397_0;
	wire [2:0] w_n398_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n402_0;
	wire [2:0] w_n402_1;
	wire [1:0] w_n402_2;
	wire [1:0] w_n403_0;
	wire [2:0] w_n405_0;
	wire [2:0] w_n405_1;
	wire [1:0] w_n405_2;
	wire [1:0] w_n407_0;
	wire [1:0] w_n408_0;
	wire [2:0] w_n410_0;
	wire [1:0] w_n410_1;
	wire [1:0] w_n414_0;
	wire [1:0] w_n416_0;
	wire [2:0] w_n419_0;
	wire [2:0] w_n424_0;
	wire [2:0] w_n424_1;
	wire [1:0] w_n424_2;
	wire [1:0] w_n426_0;
	wire [1:0] w_n434_0;
	wire [2:0] w_n435_0;
	wire [2:0] w_n435_1;
	wire [2:0] w_n437_0;
	wire [2:0] w_n437_1;
	wire [1:0] w_n445_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n449_1;
	wire [2:0] w_n451_0;
	wire [1:0] w_n451_1;
	wire [1:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [1:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [1:0] w_n471_1;
	wire [2:0] w_n473_0;
	wire [2:0] w_n473_1;
	wire [1:0] w_n481_0;
	wire [2:0] w_n484_0;
	wire [1:0] w_n484_1;
	wire [2:0] w_n486_0;
	wire [1:0] w_n486_1;
	wire [1:0] w_n494_0;
	wire [2:0] w_n495_0;
	wire [2:0] w_n495_1;
	wire [2:0] w_n497_0;
	wire [1:0] w_n497_1;
	wire [1:0] w_n505_0;
	wire [2:0] w_n507_0;
	wire [1:0] w_n507_1;
	wire [1:0] w_n509_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n518_0;
	wire [1:0] w_n518_1;
	wire [2:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [1:0] w_n530_1;
	wire [1:0] w_n532_0;
	wire [1:0] w_n540_0;
	wire [2:0] w_n541_0;
	wire [1:0] w_n541_1;
	wire [1:0] w_n543_0;
	wire [1:0] w_n551_0;
	wire [2:0] w_n556_0;
	wire [2:0] w_n556_1;
	wire [2:0] w_n556_2;
	wire [2:0] w_n556_3;
	wire [2:0] w_n556_4;
	wire [1:0] w_n556_5;
	wire [2:0] w_n560_0;
	wire [1:0] w_n560_1;
	wire [2:0] w_n561_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n567_0;
	wire [1:0] w_n567_1;
	wire [1:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [2:0] w_n571_0;
	wire [1:0] w_n571_1;
	wire [2:0] w_n572_0;
	wire [2:0] w_n574_0;
	wire [2:0] w_n577_0;
	wire [2:0] w_n578_0;
	wire [2:0] w_n582_0;
	wire [1:0] w_n582_1;
	wire [2:0] w_n583_0;
	wire [1:0] w_n583_1;
	wire [1:0] w_n585_0;
	wire [2:0] w_n587_0;
	wire [1:0] w_n587_1;
	wire [2:0] w_n590_0;
	wire [1:0] w_n590_1;
	wire [1:0] w_n591_0;
	wire [2:0] w_n595_0;
	wire [1:0] w_n595_1;
	wire [2:0] w_n596_0;
	wire [2:0] w_n600_0;
	wire [1:0] w_n600_1;
	wire [1:0] w_n601_0;
	wire [2:0] w_n604_0;
	wire [2:0] w_n605_0;
	wire [2:0] w_n605_1;
	wire [2:0] w_n605_2;
	wire [2:0] w_n607_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n609_1;
	wire [2:0] w_n609_2;
	wire [2:0] w_n609_3;
	wire [2:0] w_n609_4;
	wire [2:0] w_n609_5;
	wire [2:0] w_n613_0;
	wire [2:0] w_n614_0;
	wire [2:0] w_n614_1;
	wire [1:0] w_n614_2;
	wire [2:0] w_n617_0;
	wire [1:0] w_n617_1;
	wire [2:0] w_n618_0;
	wire [1:0] w_n618_1;
	wire [2:0] w_n621_0;
	wire [2:0] w_n621_1;
	wire [1:0] w_n621_2;
	wire [2:0] w_n622_0;
	wire [1:0] w_n622_1;
	wire [1:0] w_n623_0;
	wire [2:0] w_n624_0;
	wire [2:0] w_n624_1;
	wire [2:0] w_n625_0;
	wire [2:0] w_n628_0;
	wire [2:0] w_n629_0;
	wire [1:0] w_n631_0;
	wire [2:0] w_n633_0;
	wire [1:0] w_n633_1;
	wire [2:0] w_n636_0;
	wire [1:0] w_n636_1;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [1:0] w_n641_0;
	wire [1:0] w_n642_0;
	wire [2:0] w_n645_0;
	wire [2:0] w_n646_0;
	wire [2:0] w_n649_0;
	wire [1:0] w_n649_1;
	wire [1:0] w_n650_0;
	wire [2:0] w_n651_0;
	wire [1:0] w_n651_1;
	wire [1:0] w_n652_0;
	wire [1:0] w_n661_0;
	wire [1:0] w_n671_0;
	wire [1:0] w_n677_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n679_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n681_0;
	wire [2:0] w_n681_1;
	wire [1:0] w_n681_2;
	wire [1:0] w_n682_0;
	wire [2:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [2:0] w_n691_0;
	wire [2:0] w_n693_0;
	wire [2:0] w_n696_0;
	wire [1:0] w_n697_0;
	wire [1:0] w_n700_0;
	wire [1:0] w_n702_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n705_0;
	wire [1:0] w_n706_0;
	wire [2:0] w_n707_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n716_0;
	wire [2:0] w_n717_0;
	wire [1:0] w_n720_0;
	wire [2:0] w_n721_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n726_0;
	wire [2:0] w_n727_0;
	wire [2:0] w_n729_0;
	wire [1:0] w_n729_1;
	wire [2:0] w_n732_0;
	wire [1:0] w_n733_0;
	wire [1:0] w_n735_0;
	wire [1:0] w_n736_0;
	wire [2:0] w_n739_0;
	wire [1:0] w_n739_1;
	wire [1:0] w_n740_0;
	wire [1:0] w_n741_0;
	wire [1:0] w_n742_0;
	wire [2:0] w_n744_0;
	wire [2:0] w_n744_1;
	wire [2:0] w_n746_0;
	wire [2:0] w_n746_1;
	wire [2:0] w_n747_0;
	wire [2:0] w_n747_1;
	wire [2:0] w_n747_2;
	wire [2:0] w_n747_3;
	wire [2:0] w_n748_0;
	wire [2:0] w_n748_1;
	wire [2:0] w_n748_2;
	wire [2:0] w_n748_3;
	wire [1:0] w_n748_4;
	wire [2:0] w_n750_0;
	wire [1:0] w_n750_1;
	wire [2:0] w_n751_0;
	wire [2:0] w_n751_1;
	wire [1:0] w_n751_2;
	wire [2:0] w_n753_0;
	wire [2:0] w_n753_1;
	wire [2:0] w_n753_2;
	wire [2:0] w_n753_3;
	wire [2:0] w_n753_4;
	wire [2:0] w_n753_5;
	wire [2:0] w_n753_6;
	wire [2:0] w_n753_7;
	wire [1:0] w_n753_8;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n761_0;
	wire [2:0] w_n765_0;
	wire [2:0] w_n765_1;
	wire [2:0] w_n765_2;
	wire [2:0] w_n765_3;
	wire [2:0] w_n765_4;
	wire [2:0] w_n765_5;
	wire [1:0] w_n771_0;
	wire [1:0] w_n779_0;
	wire [2:0] w_n781_0;
	wire [2:0] w_n783_0;
	wire [1:0] w_n783_1;
	wire [1:0] w_n786_0;
	wire [1:0] w_n787_0;
	wire [2:0] w_n789_0;
	wire [2:0] w_n791_0;
	wire [1:0] w_n791_1;
	wire [1:0] w_n792_0;
	wire [2:0] w_n793_0;
	wire [2:0] w_n793_1;
	wire [2:0] w_n793_2;
	wire [2:0] w_n793_3;
	wire [1:0] w_n793_4;
	wire [2:0] w_n795_0;
	wire [1:0] w_n795_1;
	wire [1:0] w_n796_0;
	wire [2:0] w_n797_0;
	wire [2:0] w_n797_1;
	wire [2:0] w_n797_2;
	wire [2:0] w_n797_3;
	wire [1:0] w_n797_4;
	wire [2:0] w_n799_0;
	wire [2:0] w_n799_1;
	wire [2:0] w_n799_2;
	wire [2:0] w_n799_3;
	wire [1:0] w_n799_4;
	wire [2:0] w_n801_0;
	wire [2:0] w_n801_1;
	wire [2:0] w_n801_2;
	wire [2:0] w_n801_3;
	wire [1:0] w_n801_4;
	wire [2:0] w_n806_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n821_0;
	wire [2:0] w_n828_0;
	wire [1:0] w_n829_0;
	wire [1:0] w_n832_0;
	wire [1:0] w_n839_0;
	wire [2:0] w_n840_0;
	wire [2:0] w_n840_1;
	wire [2:0] w_n840_2;
	wire [2:0] w_n840_3;
	wire [1:0] w_n840_4;
	wire [1:0] w_n842_0;
	wire [2:0] w_n843_0;
	wire [2:0] w_n843_1;
	wire [2:0] w_n843_2;
	wire [2:0] w_n843_3;
	wire [1:0] w_n843_4;
	wire [2:0] w_n845_0;
	wire [2:0] w_n845_1;
	wire [2:0] w_n845_2;
	wire [2:0] w_n845_3;
	wire [1:0] w_n845_4;
	wire [2:0] w_n847_0;
	wire [2:0] w_n847_1;
	wire [2:0] w_n847_2;
	wire [2:0] w_n847_3;
	wire [1:0] w_n847_4;
	wire [1:0] w_n853_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n856_0;
	wire [1:0] w_n857_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n862_0;
	wire [1:0] w_n869_0;
	wire [1:0] w_n877_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n892_0;
	wire [1:0] w_n914_0;
	wire [1:0] w_n928_0;
	wire [2:0] w_n930_0;
	wire [1:0] w_n932_0;
	wire [2:0] w_n936_0;
	wire [1:0] w_n938_0;
	wire [1:0] w_n941_0;
	wire [1:0] w_n943_0;
	wire [1:0] w_n944_0;
	wire [1:0] w_n946_0;
	wire [2:0] w_n948_0;
	wire [1:0] w_n953_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n968_0;
	wire [1:0] w_n971_0;
	wire [1:0] w_n972_0;
	wire [1:0] w_n973_0;
	wire [1:0] w_n984_0;
	wire [2:0] w_n985_0;
	wire [2:0] w_n985_1;
	wire [2:0] w_n985_2;
	wire [2:0] w_n985_3;
	wire [1:0] w_n985_4;
	wire [1:0] w_n987_0;
	wire [2:0] w_n988_0;
	wire [2:0] w_n988_1;
	wire [2:0] w_n988_2;
	wire [2:0] w_n988_3;
	wire [1:0] w_n988_4;
	wire [2:0] w_n990_0;
	wire [2:0] w_n990_1;
	wire [2:0] w_n990_2;
	wire [2:0] w_n990_3;
	wire [1:0] w_n990_4;
	wire [2:0] w_n992_0;
	wire [2:0] w_n992_1;
	wire [2:0] w_n992_2;
	wire [2:0] w_n992_3;
	wire [1:0] w_n992_4;
	wire [1:0] w_n998_0;
	wire [2:0] w_n999_0;
	wire [2:0] w_n999_1;
	wire [2:0] w_n999_2;
	wire [2:0] w_n999_3;
	wire [1:0] w_n999_4;
	wire [1:0] w_n1001_0;
	wire [2:0] w_n1002_0;
	wire [2:0] w_n1002_1;
	wire [2:0] w_n1002_2;
	wire [2:0] w_n1002_3;
	wire [1:0] w_n1002_4;
	wire [2:0] w_n1004_0;
	wire [2:0] w_n1004_1;
	wire [2:0] w_n1004_2;
	wire [2:0] w_n1004_3;
	wire [1:0] w_n1004_4;
	wire [2:0] w_n1006_0;
	wire [2:0] w_n1006_1;
	wire [2:0] w_n1006_2;
	wire [2:0] w_n1006_3;
	wire [1:0] w_n1006_4;
	wire [2:0] w_n1012_0;
	wire [1:0] w_n1012_1;
	wire [2:0] w_n1014_0;
	wire [1:0] w_n1014_1;
	wire [2:0] w_n1021_0;
	wire [1:0] w_n1021_1;
	wire [2:0] w_n1023_0;
	wire [1:0] w_n1023_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1032_0;
	wire [1:0] w_n1032_1;
	wire [2:0] w_n1039_0;
	wire [1:0] w_n1039_1;
	wire [2:0] w_n1041_0;
	wire [1:0] w_n1041_1;
	wire [1:0] w_n1142_0;
	wire [1:0] w_n1151_0;
	wire [2:0] w_n1163_0;
	wire [2:0] w_n1163_1;
	wire [2:0] w_n1197_0;
	wire [2:0] w_n1197_1;
	wire [2:0] w_n1205_0;
	wire [2:0] w_n1205_1;
	wire [2:0] w_n1235_0;
	wire [1:0] w_n1235_1;
	wire [2:0] w_n1242_0;
	wire [1:0] w_n1242_1;
	wire [2:0] w_n1244_0;
	wire [1:0] w_n1244_1;
	wire [2:0] w_n1251_0;
	wire [1:0] w_n1251_1;
	wire [2:0] w_n1253_0;
	wire [1:0] w_n1253_1;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1383_0;
	wire [1:0] w_n1391_0;
	wire [1:0] w_n1394_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1399_0;
	wire [1:0] w_n1409_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1411_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1434_0;
	wire [1:0] w_n1438_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1452_0;
	wire [1:0] w_n1494_0;
	wire [1:0] w_n1533_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1553_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1568_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1597_0;
	wire [2:0] w_n1601_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1609_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1624_0;
	wire [1:0] w_n1629_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1634_0;
	wire w_dff_B_XssIjf5V0_1;
	wire w_dff_B_Dal5NXoy4_0;
	wire w_dff_B_Mca1lwmy8_1;
	wire w_dff_B_Fm0mRtxx3_1;
	wire w_dff_B_D7BgWf7S7_2;
	wire w_dff_B_S57yGqN83_1;
	wire w_dff_B_fnTBsdyL9_1;
	wire w_dff_B_IrVW51x29_0;
	wire w_dff_B_KSZfTLzP9_1;
	wire w_dff_B_ODt69OBG6_1;
	wire w_dff_B_TiA3PYaH3_0;
	wire w_dff_B_Jfk8n5Ey8_1;
	wire w_dff_A_WQWmgh6x2_0;
	wire w_dff_A_gygGVr8w1_0;
	wire w_dff_A_fB1lmueH0_0;
	wire w_dff_A_NRmMTPDk0_0;
	wire w_dff_A_AFxMaLQZ3_1;
	wire w_dff_A_9EmKaLaE6_1;
	wire w_dff_A_yAeXsPl21_1;
	wire w_dff_A_9tMO6vDT1_1;
	wire w_dff_B_Gkskymn36_1;
	wire w_dff_B_p9XI6owv5_0;
	wire w_dff_B_cVsNJJHb0_1;
	wire w_dff_B_JmCqyBqc5_1;
	wire w_dff_B_aSvu7Tg51_0;
	wire w_dff_B_dEkF10QY7_1;
	wire w_dff_A_ZMRpH7Cm0_0;
	wire w_dff_A_bt1O9L7I5_1;
	wire w_dff_A_J13aWE4G7_1;
	wire w_dff_A_tFnwf5qe7_1;
	wire w_dff_A_HybsOoa34_1;
	wire w_dff_A_8SuW07jG0_1;
	wire w_dff_A_ihCZD1qn1_2;
	wire w_dff_A_zVDY3vDk9_2;
	wire w_dff_A_MJuLq9HB7_2;
	wire w_dff_A_a5cZcJOE8_2;
	wire w_dff_B_WsR53Ip04_1;
	wire w_dff_B_3CzV9Jej8_1;
	wire w_dff_B_Nz0flp8Q2_0;
	wire w_dff_B_pkjSE7L20_1;
	wire w_dff_B_kW56YRH88_1;
	wire w_dff_B_Ly8y0O7P7_2;
	wire w_dff_B_HmIOfsGO3_2;
	wire w_dff_B_DEkXRBgq2_2;
	wire w_dff_B_giZSAE6j8_2;
	wire w_dff_B_8PzF9dIk4_1;
	wire w_dff_B_ED7Z7xQZ9_1;
	wire w_dff_B_2WzSiiHc7_1;
	wire w_dff_B_7XrR9Fu38_1;
	wire w_dff_B_ip7ldRLj3_1;
	wire w_dff_B_ZcvBg8Sc2_1;
	wire w_dff_B_fnflHZ8W5_1;
	wire w_dff_A_hrZEm7iI5_1;
	wire w_dff_A_bispfRPv1_1;
	wire w_dff_B_vZrKh8sv0_3;
	wire w_dff_B_yYpi79nI5_3;
	wire w_dff_B_NxnJO8Er8_3;
	wire w_dff_B_AeDOD12Z9_0;
	wire w_dff_B_whth4iwK4_2;
	wire w_dff_B_5CtWqWG32_2;
	wire w_dff_B_f5WSunBa1_2;
	wire w_dff_B_YGtMakNp9_2;
	wire w_dff_B_2SZsCcUg8_2;
	wire w_dff_A_Z33aOacp4_0;
	wire w_dff_A_QHGVysha6_0;
	wire w_dff_A_vT0gjAMZ6_0;
	wire w_dff_A_JAk0xbai5_0;
	wire w_dff_A_IN0CntKv1_0;
	wire w_dff_A_KZ6qEmH77_0;
	wire w_dff_B_PhzMjzHb8_0;
	wire w_dff_B_fBDCGOM50_0;
	wire w_dff_B_rGxtK9wi5_0;
	wire w_dff_B_ph7LqdJY4_0;
	wire w_dff_B_3ewiIPnx2_0;
	wire w_dff_B_viMLJl540_0;
	wire w_dff_B_b35jbf2Z3_0;
	wire w_dff_B_zpGI0mAt6_0;
	wire w_dff_B_nQPXoJiJ7_0;
	wire w_dff_B_rgBzz1bG1_0;
	wire w_dff_B_U2olVBQR0_0;
	wire w_dff_B_yMh7HUE44_0;
	wire w_dff_B_MZhMwQa67_2;
	wire w_dff_B_5X48FtVM3_2;
	wire w_dff_B_CChcr1BA4_2;
	wire w_dff_B_bXABOWnN9_0;
	wire w_dff_B_W2wYqFAe1_0;
	wire w_dff_B_KaCYtSDu2_0;
	wire w_dff_B_IrpWIMHD3_1;
	wire w_dff_B_EhSDyr2c9_1;
	wire w_dff_B_InlKldaq1_1;
	wire w_dff_B_3wJGaPeF1_1;
	wire w_dff_B_WESzWxWL2_0;
	wire w_dff_B_mSFnHuVU1_0;
	wire w_dff_B_mAUt7xJU8_0;
	wire w_dff_B_tjDkCpYo4_0;
	wire w_dff_B_wAe7Cz920_0;
	wire w_dff_B_DEajMSUz6_0;
	wire w_dff_B_99g6zTEi2_0;
	wire w_dff_B_1qYgqFH83_0;
	wire w_dff_B_RAli3rd30_0;
	wire w_dff_B_0MqjEfGd0_0;
	wire w_dff_B_8OjgUUdK4_0;
	wire w_dff_B_yzSYTJWf6_0;
	wire w_dff_B_R7asPy7h5_0;
	wire w_dff_B_M9SHpA5H4_0;
	wire w_dff_B_fSRNsPI46_0;
	wire w_dff_B_XV3u2wTd0_0;
	wire w_dff_B_avY0gwYw0_0;
	wire w_dff_B_6TjWitqE6_0;
	wire w_dff_B_E8Ow1mSb0_2;
	wire w_dff_B_mg0MgxRV1_2;
	wire w_dff_B_uQNPPLHu0_2;
	wire w_dff_B_wwrx8AHY9_1;
	wire w_dff_B_B227RsBo4_0;
	wire w_dff_B_xFtzP4mP1_1;
	wire w_dff_B_QRg1MG1I3_1;
	wire w_dff_B_CzAGbBpC4_0;
	wire w_dff_B_33JdFQzd1_0;
	wire w_dff_B_plweYquy5_1;
	wire w_dff_B_gUgiBgL93_1;
	wire w_dff_B_qPKMQyte9_0;
	wire w_dff_B_KjOV1hzk1_1;
	wire w_dff_B_47TbZlIf2_0;
	wire w_dff_B_4FPXO9oq2_0;
	wire w_dff_B_9do6CGYe5_0;
	wire w_dff_B_DK7afoQR6_0;
	wire w_dff_B_FWWB7Nqj3_0;
	wire w_dff_B_PEUGs7Ix9_0;
	wire w_dff_B_CygcLcqT8_0;
	wire w_dff_B_piNr54hs0_0;
	wire w_dff_B_JYeiFR921_0;
	wire w_dff_B_Rv5YJH7z6_0;
	wire w_dff_B_vn7svMmu9_0;
	wire w_dff_B_BAeuSWTx6_0;
	wire w_dff_B_ztWLRg0X4_0;
	wire w_dff_B_Ww6v3SSi1_0;
	wire w_dff_A_q3zLCPm63_0;
	wire w_dff_A_A48mdAmP4_0;
	wire w_dff_A_LvF52s4v5_0;
	wire w_dff_A_a47M2xaZ7_0;
	wire w_dff_A_ZgPCGr6Y6_0;
	wire w_dff_A_fcQliiep9_0;
	wire w_dff_A_DrEaSfxY2_0;
	wire w_dff_A_3dQy5vFe3_0;
	wire w_dff_A_xq15hH6Z1_0;
	wire w_dff_A_cvnKx47M1_0;
	wire w_dff_A_Uwkh47Si4_0;
	wire w_dff_A_sJx77pRG2_0;
	wire w_dff_A_VC7dsWwV8_0;
	wire w_dff_A_m61YsGgv0_0;
	wire w_dff_A_pDba1ues0_0;
	wire w_dff_B_4QTYj42L0_0;
	wire w_dff_B_CYoRH7bO6_0;
	wire w_dff_B_8sSrWfTZ6_0;
	wire w_dff_B_8w1o0Pwi9_0;
	wire w_dff_B_bvSipQJx4_0;
	wire w_dff_B_c7m6rXMD7_0;
	wire w_dff_B_m58G5xzA9_0;
	wire w_dff_B_4fJtjy4U4_0;
	wire w_dff_B_CDytwPxH1_0;
	wire w_dff_B_rwa9BTLw4_0;
	wire w_dff_B_gz8CIbCF7_0;
	wire w_dff_B_jHgqreCB4_0;
	wire w_dff_B_QIFUOnRh2_0;
	wire w_dff_B_syxrlt572_0;
	wire w_dff_B_ZkBOZRCt1_0;
	wire w_dff_B_Kmqbff6M7_0;
	wire w_dff_B_blFGw6jZ5_0;
	wire w_dff_B_e5WHWo593_0;
	wire w_dff_B_7ZzqMHBu9_0;
	wire w_dff_B_XbiAhNVy0_0;
	wire w_dff_B_P6BvjMBa8_0;
	wire w_dff_B_45NXoFSz2_0;
	wire w_dff_B_gOnz1Z622_0;
	wire w_dff_B_zng9M7Sd3_0;
	wire w_dff_B_KQnOpBxn5_0;
	wire w_dff_B_fvPzOQNK9_0;
	wire w_dff_B_KLoCxCNO9_0;
	wire w_dff_B_5xcSTM5P5_0;
	wire w_dff_B_fdVVnm3y2_0;
	wire w_dff_B_KEyaKCrz6_0;
	wire w_dff_B_MDnUbVep0_0;
	wire w_dff_B_zRMVweWr4_0;
	wire w_dff_B_04HM0IyZ8_0;
	wire w_dff_A_Oc0bOI7p6_1;
	wire w_dff_A_Y9bywIRN2_1;
	wire w_dff_A_ZwpPDw3o7_2;
	wire w_dff_A_5SOsB5WF6_2;
	wire w_dff_A_8pRe6LkT2_2;
	wire w_dff_A_rTCJRv862_2;
	wire w_dff_A_8LEd86GY1_1;
	wire w_dff_A_eHXEDivT4_2;
	wire w_dff_A_kG0CDKnq1_2;
	wire w_dff_B_lpijphA11_0;
	wire w_dff_B_GYqsEJOj8_0;
	wire w_dff_B_i6JhRNwU6_0;
	wire w_dff_B_gmAs5Kix2_0;
	wire w_dff_B_jBIxtsFT1_0;
	wire w_dff_B_7CYsb0fn5_0;
	wire w_dff_B_WgB243ov3_0;
	wire w_dff_B_VRcPIPAr5_0;
	wire w_dff_B_0IPoP4RU7_0;
	wire w_dff_B_gq8X0Bec3_0;
	wire w_dff_B_CLUWGzWf2_0;
	wire w_dff_B_J9GBjOcs0_0;
	wire w_dff_B_IqO4jrNW8_0;
	wire w_dff_B_JUusCXk67_0;
	wire w_dff_B_S7J5IsmI3_2;
	wire w_dff_B_Rli16P8U4_2;
	wire w_dff_B_dxC1OtnG9_2;
	wire w_dff_A_H9e2wXoZ0_0;
	wire w_dff_A_4VNwIuYC1_0;
	wire w_dff_A_mhPKSX9G0_0;
	wire w_dff_A_00N8qH0f4_0;
	wire w_dff_A_6Rxdd2bt0_0;
	wire w_dff_A_P2fmNh136_0;
	wire w_dff_A_7Ey6VMuo4_0;
	wire w_dff_A_rBWeQVvN4_0;
	wire w_dff_A_wE6aJrTb1_0;
	wire w_dff_A_h3x6bsEl5_0;
	wire w_dff_A_sgNgf0vX6_0;
	wire w_dff_A_waHlxvN38_0;
	wire w_dff_A_pamI7Pxv1_0;
	wire w_dff_A_6f9epyeH3_0;
	wire w_dff_A_2YFHNRle2_0;
	wire w_dff_B_tm7n7pgN3_0;
	wire w_dff_B_spxeXEEB7_0;
	wire w_dff_B_B0H0h72i4_0;
	wire w_dff_B_StLHkQiI3_0;
	wire w_dff_B_3PaLHpKP9_0;
	wire w_dff_B_euwC8bRQ4_0;
	wire w_dff_B_PJQewawI0_0;
	wire w_dff_B_DDX5Fy4I6_0;
	wire w_dff_B_NqcF3pch4_0;
	wire w_dff_B_Je3HVV2R8_0;
	wire w_dff_B_e9AgWHTM3_0;
	wire w_dff_B_bMwGzXBW6_0;
	wire w_dff_B_ntYLpOYK3_2;
	wire w_dff_B_K85BdsWi9_2;
	wire w_dff_B_l3xCiwCo2_2;
	wire w_dff_B_XCDHoueb2_0;
	wire w_dff_B_TErgr8ko2_0;
	wire w_dff_B_unBvVqnu6_0;
	wire w_dff_B_D9SjgIIo7_0;
	wire w_dff_B_ajTPpUqU0_0;
	wire w_dff_B_hQ1ZOIEw6_0;
	wire w_dff_B_sgHFWcFo8_0;
	wire w_dff_B_JyGP5icQ1_0;
	wire w_dff_B_u5lrbKGc5_0;
	wire w_dff_B_TKf1DxH57_0;
	wire w_dff_B_NwksgsXy5_0;
	wire w_dff_B_JPVxV5JX3_2;
	wire w_dff_B_41uG2RLG8_2;
	wire w_dff_B_SAJzS6I19_2;
	wire w_dff_B_DMJtnIM71_0;
	wire w_dff_B_nyxe27eH1_0;
	wire w_dff_B_J3jcYmM34_0;
	wire w_dff_B_O7THjFWr7_0;
	wire w_dff_B_GaElTtFk0_0;
	wire w_dff_B_dIDC2yNE2_0;
	wire w_dff_B_Mb9koHU65_0;
	wire w_dff_B_NBwEMJkl1_0;
	wire w_dff_B_QKeZNlHr6_0;
	wire w_dff_B_TZ3jdvfl1_0;
	wire w_dff_B_gGqDyEHP8_2;
	wire w_dff_B_tFN5R1Mz9_2;
	wire w_dff_B_dmDgtYiK5_2;
	wire w_dff_A_P2xNaJpc5_1;
	wire w_dff_A_np2aySLL9_1;
	wire w_dff_A_wHs9jq1k8_2;
	wire w_dff_A_4OVrbwy44_2;
	wire w_dff_A_oxwMc8g02_2;
	wire w_dff_A_ILrysShD0_2;
	wire w_dff_A_2SUQv1QZ1_1;
	wire w_dff_A_1WNx31T11_2;
	wire w_dff_A_GSoiYBCs5_2;
	wire w_dff_B_XTnXtpgM8_0;
	wire w_dff_B_gtS9rtlA1_0;
	wire w_dff_B_a4nihD729_0;
	wire w_dff_B_Xh8RYayb9_0;
	wire w_dff_B_mCRNHctH2_0;
	wire w_dff_B_x8zkF9130_0;
	wire w_dff_B_vn3QLHjX3_0;
	wire w_dff_B_KW5161zW1_0;
	wire w_dff_B_kcz1biqD4_0;
	wire w_dff_B_GB4tiu9b0_0;
	wire w_dff_B_ay1FvGnp2_0;
	wire w_dff_B_DhAD15Lh7_0;
	wire w_dff_B_W3ZZw4Cn9_0;
	wire w_dff_B_WjCWHaAT4_0;
	wire w_dff_A_BxdxAuTy3_0;
	wire w_dff_A_QRetefqs5_0;
	wire w_dff_A_0rMw0z2f3_0;
	wire w_dff_A_fMXsBj9m6_0;
	wire w_dff_A_MmLzWgdh3_0;
	wire w_dff_A_noo8JoPT4_0;
	wire w_dff_A_LzgFPlqJ2_0;
	wire w_dff_A_gHzBM0LF5_0;
	wire w_dff_A_EysPXUwI6_0;
	wire w_dff_A_AyI6GO7f7_0;
	wire w_dff_A_guqWhoe00_0;
	wire w_dff_A_YiYShXeA3_0;
	wire w_dff_A_KRV72M3l8_0;
	wire w_dff_A_KyShtKWw0_0;
	wire w_dff_A_p7tmQuyS8_0;
	wire w_dff_B_FHdlhyxr5_0;
	wire w_dff_B_P6gQ9s1P0_0;
	wire w_dff_B_T3z170Uf8_0;
	wire w_dff_B_gq0Tum2J9_0;
	wire w_dff_B_oBnIaTDD1_0;
	wire w_dff_B_TWbyM5508_0;
	wire w_dff_B_nXtGAaXD7_0;
	wire w_dff_B_uSdc2ox50_0;
	wire w_dff_B_W18ARSSY5_0;
	wire w_dff_B_UroukBto2_0;
	wire w_dff_B_EoeafYTF2_0;
	wire w_dff_B_KlIGP9566_0;
	wire w_dff_B_K7rIN2yn3_0;
	wire w_dff_B_62J7ihQl9_0;
	wire w_dff_B_1v5WwXJz9_0;
	wire w_dff_B_bxUHRyXk9_0;
	wire w_dff_B_kriV0NXd8_0;
	wire w_dff_B_c7xR3tpJ3_0;
	wire w_dff_B_3E2BngQZ8_0;
	wire w_dff_B_D7JximM67_0;
	wire w_dff_B_0aRS2stc2_0;
	wire w_dff_A_1BC24AqY8_0;
	wire w_dff_A_gko4YKyK2_2;
	wire w_dff_A_px96T8OU9_2;
	wire w_dff_A_E9gPA6Lu8_2;
	wire w_dff_A_e6UNA8IQ6_2;
	wire w_dff_B_BprNyinQ4_0;
	wire w_dff_B_OS5ZA7bL9_0;
	wire w_dff_B_VEjMUxYL5_0;
	wire w_dff_B_no1Xjybo0_0;
	wire w_dff_B_EmVfzZRj6_0;
	wire w_dff_B_1KUHvEMk1_0;
	wire w_dff_B_x8V8CaWD3_0;
	wire w_dff_B_u5SYxqAU4_0;
	wire w_dff_B_JaNqa41D0_0;
	wire w_dff_B_soNc0u147_0;
	wire w_dff_B_5qbHPi520_0;
	wire w_dff_B_xkoqWe9W8_0;
	wire w_dff_A_DyrteZ6p1_0;
	wire w_dff_A_HppuP6Js1_0;
	wire w_dff_A_DDViaX6f7_0;
	wire w_dff_A_dpyfnwzd8_0;
	wire w_dff_A_atiftQfm6_1;
	wire w_dff_A_SSmOGXFU7_1;
	wire w_dff_A_qNjLDCVg7_0;
	wire w_dff_A_fCAycZkA0_0;
	wire w_dff_A_cN4ywjen3_1;
	wire w_dff_B_OgIeoO6B4_0;
	wire w_dff_B_En1prRs44_0;
	wire w_dff_B_fwlSjpo56_0;
	wire w_dff_B_upMTLFBi1_0;
	wire w_dff_B_QNvj0gwz1_0;
	wire w_dff_B_ZhMkt2bJ3_0;
	wire w_dff_B_9dOWhQTQ3_0;
	wire w_dff_B_zThJXWQv4_0;
	wire w_dff_B_vl0nWUn87_0;
	wire w_dff_B_8NuyTHxS8_0;
	wire w_dff_B_KanJafkY3_0;
	wire w_dff_B_70WijCaP4_0;
	wire w_dff_B_GzcXBlx84_0;
	wire w_dff_B_5KDeyqNZ2_0;
	wire w_dff_B_JcnLwAmB3_2;
	wire w_dff_B_XcbrhrKy6_2;
	wire w_dff_B_YbWxK6xW4_2;
	wire w_dff_A_9eKJdbRh4_0;
	wire w_dff_A_sLqpRWvs9_0;
	wire w_dff_A_GgBhcmtO9_0;
	wire w_dff_A_47zHNPzp2_0;
	wire w_dff_A_deeyw11t2_0;
	wire w_dff_A_6Vi4GMIZ8_0;
	wire w_dff_A_kMyjH4IQ1_0;
	wire w_dff_B_ZpKwYiag7_0;
	wire w_dff_B_AP3B4fjv9_0;
	wire w_dff_B_BOcGSZIL7_0;
	wire w_dff_B_RgcqJiYQ9_0;
	wire w_dff_B_COUyQcJW3_0;
	wire w_dff_B_6PCInH3y0_0;
	wire w_dff_B_eKL3llTz4_0;
	wire w_dff_B_FDZowcrK5_0;
	wire w_dff_B_MC7EYT0u1_1;
	wire w_dff_B_TXDqdpuD8_1;
	wire w_dff_B_6x1nUjZV6_0;
	wire w_dff_B_9iNE9XXP0_1;
	wire w_dff_A_RR97Thn17_0;
	wire w_dff_A_7nm7N9su5_0;
	wire w_dff_A_3MCc1XmU7_0;
	wire w_dff_A_waTVUbUa8_0;
	wire w_dff_A_Rr2iFJ0p9_0;
	wire w_dff_A_exPsBILN4_0;
	wire w_dff_A_mLONIbjn9_0;
	wire w_dff_A_a9Qm4DtW7_0;
	wire w_dff_B_fq9rhGuf4_0;
	wire w_dff_B_PuyzAVSH1_0;
	wire w_dff_B_8mQ0XSkc9_0;
	wire w_dff_B_R7YEhzvu4_0;
	wire w_dff_B_PR0izhPs7_0;
	wire w_dff_B_ULeG9tiY5_0;
	wire w_dff_B_Vk0JY3u23_0;
	wire w_dff_B_94rHWRBM0_0;
	wire w_dff_B_1cLKOKWl7_0;
	wire w_dff_B_WUOp7OYO9_0;
	wire w_dff_B_M89nhxxV1_1;
	wire w_dff_B_Pvx58Jyu8_1;
	wire w_dff_B_FGBLF5RG1_0;
	wire w_dff_B_4NDoHUfP4_1;
	wire w_dff_B_iNlZN9jk3_1;
	wire w_dff_B_5zist2W43_1;
	wire w_dff_B_EmjnAZEq6_1;
	wire w_dff_B_pHWzAP7Y9_1;
	wire w_dff_B_AuHxWxW40_1;
	wire w_dff_B_73bDIewy7_1;
	wire w_dff_B_IomaU9x00_0;
	wire w_dff_B_b8GBKIl80_0;
	wire w_dff_B_CNjIMwUF5_0;
	wire w_dff_B_iljtuNsl0_0;
	wire w_dff_B_OKBLelgK2_0;
	wire w_dff_B_aOxlDQ062_0;
	wire w_dff_B_yOorlP4o7_0;
	wire w_dff_B_PZcdhNna8_0;
	wire w_dff_B_wahLog2R8_0;
	wire w_dff_B_Dria40VK9_0;
	wire w_dff_B_rhmpJRnq2_2;
	wire w_dff_B_Kcwo7PKd4_2;
	wire w_dff_B_oPu1wzDG3_2;
	wire w_dff_B_wTdfFCYR9_0;
	wire w_dff_B_Dplxahew3_0;
	wire w_dff_B_0cZsRaBs4_1;
	wire w_dff_B_UlMVrDl49_1;
	wire w_dff_A_y5ATf2KU7_1;
	wire w_dff_B_hpRNacob3_0;
	wire w_dff_B_ME1rjpGW3_1;
	wire w_dff_A_zE2BDkb14_0;
	wire w_dff_B_1cDh0C0P1_0;
	wire w_dff_B_e6H0owVM2_0;
	wire w_dff_B_XV6f11p15_0;
	wire w_dff_B_i7cpOCT88_0;
	wire w_dff_B_2NrrkCob0_0;
	wire w_dff_B_WEhjN6ji8_0;
	wire w_dff_B_HkCz8Ird5_1;
	wire w_dff_B_mEvSGX876_1;
	wire w_dff_B_NznqOe2n0_0;
	wire w_dff_B_9BFouGyv7_1;
	wire w_dff_B_90uOtjj17_0;
	wire w_dff_A_Ovfi9hOb9_1;
	wire w_dff_A_g0BHYwOQ1_1;
	wire w_dff_A_973G9RMs0_1;
	wire w_dff_A_Dg47uAWB2_1;
	wire w_dff_A_MA2pURe37_2;
	wire w_dff_A_srnJSoTh0_2;
	wire w_dff_A_Rt3k4Nc34_0;
	wire w_dff_A_UZDXURbz1_0;
	wire w_dff_A_kZc9yHur4_0;
	wire w_dff_A_rYHWvkE08_0;
	wire w_dff_A_fGYOpEif8_1;
	wire w_dff_A_AHSc45R73_1;
	wire w_dff_A_hKm7mnYD0_1;
	wire w_dff_A_E3CF4CRp0_1;
	wire w_dff_B_joGhvehh8_0;
	wire w_dff_B_reDfHA2s8_0;
	wire w_dff_B_3ZpPZ9th1_0;
	wire w_dff_B_zi3z1JL30_0;
	wire w_dff_B_MY3JNuaJ7_0;
	wire w_dff_B_PFdWbYIz0_0;
	wire w_dff_B_CgAU9tAa9_0;
	wire w_dff_B_SIQJrTRL8_0;
	wire w_dff_B_t6ibS3ha3_0;
	wire w_dff_B_q1U8qdc83_0;
	wire w_dff_B_htxaFz5i3_0;
	wire w_dff_B_Jwib4FT85_2;
	wire w_dff_B_nx8Dlb4J8_2;
	wire w_dff_B_tyClrbYL5_2;
	wire w_dff_B_qGUnuodJ7_0;
	wire w_dff_B_folb1ScY3_0;
	wire w_dff_B_ItJBMpig6_0;
	wire w_dff_B_qQWnhljy2_0;
	wire w_dff_B_PgOv85E25_1;
	wire w_dff_B_oO4A8jg59_1;
	wire w_dff_B_90sOMuAW5_0;
	wire w_dff_B_AHuoukWT8_1;
	wire w_dff_A_wy6D8lKC3_0;
	wire w_dff_A_SKuI1rEA3_0;
	wire w_dff_A_aaSUKXGg5_0;
	wire w_dff_A_sW34QoFa6_0;
	wire w_dff_A_J2Ts6Yvv4_0;
	wire w_dff_A_9oh8lctW9_0;
	wire w_dff_B_Y7QT4HVk9_0;
	wire w_dff_B_V597U4Y40_0;
	wire w_dff_B_FUXuW4ch9_0;
	wire w_dff_B_xfw8lBFP9_0;
	wire w_dff_B_UWRP0Y5A5_0;
	wire w_dff_B_u9EAxGG46_0;
	wire w_dff_B_Y8q27l6j4_0;
	wire w_dff_B_cytzVKcL3_1;
	wire w_dff_B_A0F7fsOW6_1;
	wire w_dff_A_8VKltBBU2_1;
	wire w_dff_B_YwJWY0nX7_0;
	wire w_dff_B_v0xWcDdw6_1;
	wire w_dff_B_ZNFHKvU31_0;
	wire w_dff_B_6hklEctc2_0;
	wire w_dff_B_DuHVaRYy5_0;
	wire w_dff_B_WS8OTYFr8_0;
	wire w_dff_B_hLJV7IoA7_0;
	wire w_dff_B_lgFfUvub0_0;
	wire w_dff_B_PhJv75Xw4_0;
	wire w_dff_B_wPp1weZE4_0;
	wire w_dff_B_hUShEWNF6_0;
	wire w_dff_B_y8teBY6p8_0;
	wire w_dff_B_tntgAJsr9_0;
	wire w_dff_B_1vcrToXD2_0;
	wire w_dff_B_Yql3Al7D3_2;
	wire w_dff_B_eeyDiJgY2_2;
	wire w_dff_B_uqpvHaIJ6_2;
	wire w_dff_A_B0n1OQAi3_0;
	wire w_dff_A_63pvQg8h8_0;
	wire w_dff_A_BN4vH3IG5_0;
	wire w_dff_A_6mb7RBXC1_0;
	wire w_dff_A_64erkCvW5_1;
	wire w_dff_A_BCAe3P7R0_1;
	wire w_dff_B_S2Or8NpQ2_0;
	wire w_dff_B_AGGj8wiS0_0;
	wire w_dff_B_BAfeW1eF9_0;
	wire w_dff_B_35uPWueG1_0;
	wire w_dff_B_yl3JbdgC0_0;
	wire w_dff_B_J1JxYypK8_0;
	wire w_dff_B_AEPhoVEA0_1;
	wire w_dff_B_eRjeDWEg4_1;
	wire w_dff_B_Zz6Hvt2A8_0;
	wire w_dff_B_33ZGEYC72_1;
	wire w_dff_B_6NNxzr0W7_1;
	wire w_dff_B_8cbz5lvv5_1;
	wire w_dff_B_bjNjYMa54_1;
	wire w_dff_B_ltmbQhDK8_1;
	wire w_dff_A_hd1Eoys54_2;
	wire w_dff_A_GZRNoypF2_2;
	wire w_dff_A_4CavtIdX3_2;
	wire w_dff_A_wV0klqvI2_2;
	wire w_dff_B_Kk0V9Pnr3_3;
	wire w_dff_B_4K1igsW85_3;
	wire w_dff_A_sS2V6STz4_1;
	wire w_dff_A_sHOXtqEZ9_1;
	wire w_dff_A_PUPh2Q1J9_2;
	wire w_dff_A_bpcWVSnb9_2;
	wire w_dff_A_w1Xm0ZBY8_2;
	wire w_dff_A_p1fNNdqi8_2;
	wire w_dff_A_5Ni3oU0t8_0;
	wire w_dff_A_i86dQOnh2_0;
	wire w_dff_A_QwZ9RiFX5_1;
	wire w_dff_B_0iCX4q2L4_0;
	wire w_dff_B_1IUmLE8N8_0;
	wire w_dff_B_5MhM0mvX9_0;
	wire w_dff_B_PIIXsSd08_0;
	wire w_dff_B_yRUs2IVr8_0;
	wire w_dff_B_fZP1RiSL2_0;
	wire w_dff_B_EcPTGb4R5_0;
	wire w_dff_B_wCO12kb00_0;
	wire w_dff_B_CXvXgtDY2_1;
	wire w_dff_B_QJsdoiVI0_1;
	wire w_dff_B_twvL3bjd5_0;
	wire w_dff_B_XnnT7VXe0_1;
	wire w_dff_B_orm6dmTT0_0;
	wire w_dff_A_S3A9iaE13_0;
	wire w_dff_A_krEBoHMt1_0;
	wire w_dff_A_zbBOPd4Q6_0;
	wire w_dff_A_SL3qSCfQ3_0;
	wire w_dff_B_rZlufikp0_0;
	wire w_dff_B_Z8QgmcpH3_0;
	wire w_dff_B_Sx6bZPfX9_0;
	wire w_dff_B_tURWSTxm3_0;
	wire w_dff_B_EJIcXACC0_0;
	wire w_dff_B_RLQnn9YY0_0;
	wire w_dff_B_R1vwRNSd9_0;
	wire w_dff_B_KkfVonDU0_0;
	wire w_dff_B_UydwmAn19_0;
	wire w_dff_B_KFyg94CR6_0;
	wire w_dff_B_aieW1T711_0;
	wire w_dff_B_w7QhIpOV3_0;
	wire w_dff_B_JFohs4FV4_1;
	wire w_dff_B_b8ZWHRwQ6_1;
	wire w_dff_B_i6tiRbtz5_1;
	wire w_dff_B_azQH0x1a7_1;
	wire w_dff_B_FsbrXkvc7_1;
	wire w_dff_B_n1caYDXs8_1;
	wire w_dff_B_jOuKGlAG2_0;
	wire w_dff_B_XofCy3am5_0;
	wire w_dff_B_aYYrDuJW6_0;
	wire w_dff_B_PBruMV9M2_0;
	wire w_dff_B_HpBSRuLH3_0;
	wire w_dff_B_5aYLOKsi5_0;
	wire w_dff_B_tIFftIpk1_0;
	wire w_dff_B_zNJNcfz89_0;
	wire w_dff_B_ICcObu3u6_0;
	wire w_dff_B_MojCcEFQ2_0;
	wire w_dff_B_1z8FhPUv6_0;
	wire w_dff_B_Jp3qyDQ02_0;
	wire w_dff_B_5nfTkvUg1_0;
	wire w_dff_B_7N6eNxPt9_0;
	wire w_dff_B_MWWNPNaA3_0;
	wire w_dff_B_FMrwp04V2_0;
	wire w_dff_B_J0YdLulo1_1;
	wire w_dff_A_K6SzOKp15_0;
	wire w_dff_A_qeirXqOk5_0;
	wire w_dff_A_osSimo5V6_0;
	wire w_dff_A_aKgV9xIY9_0;
	wire w_dff_A_sGtT0UpU5_0;
	wire w_dff_A_wtCkzWpC0_0;
	wire w_dff_A_d2klbvkf6_0;
	wire w_dff_A_j4F8Q4Q48_0;
	wire w_dff_A_KupFvMek0_0;
	wire w_dff_A_YMQddjrZ0_0;
	wire w_dff_A_neHuwbZB1_0;
	wire w_dff_A_vCMXz4iL1_0;
	wire w_dff_A_bkx6wXmx2_2;
	wire w_dff_A_INHrCEno2_2;
	wire w_dff_A_yAzh50XK3_2;
	wire w_dff_A_fRLBZb3v8_2;
	wire w_dff_A_HVpc9jXd3_2;
	wire w_dff_A_URkEzGnw4_2;
	wire w_dff_A_DBvuUKK06_2;
	wire w_dff_A_8RgLcLau1_2;
	wire w_dff_A_T83pYknB7_2;
	wire w_dff_A_8zQhIFMF0_2;
	wire w_dff_A_GIzrlDgr3_2;
	wire w_dff_A_bbsteKd83_2;
	wire w_dff_A_9wEnWf2n6_2;
	wire w_dff_A_007DtaO53_2;
	wire w_dff_A_afgfJBNd1_2;
	wire w_dff_A_awaVXosT6_2;
	wire w_dff_A_NZxTyMrq2_2;
	wire w_dff_A_Y3km0hto5_2;
	wire w_dff_A_CyhbJpPf8_0;
	wire w_dff_A_mp7Tnzcw8_0;
	wire w_dff_A_gsfJ6xKn8_0;
	wire w_dff_A_O9AgyIXz0_0;
	wire w_dff_A_oOM8QH7N3_0;
	wire w_dff_A_GoffM0QW2_0;
	wire w_dff_A_YEkxEUIG5_0;
	wire w_dff_A_yt364Pk02_0;
	wire w_dff_A_ALYqXm6s4_0;
	wire w_dff_A_YzTymrLW3_0;
	wire w_dff_A_zzsJyB2j0_0;
	wire w_dff_A_ZG2Bd2je4_0;
	wire w_dff_A_de4oxTsm6_0;
	wire w_dff_B_eXbFNvuK9_2;
	wire w_dff_B_PQ2AeFZf3_2;
	wire w_dff_B_i0Dq756B2_2;
	wire w_dff_B_9S8cjbQD0_1;
	wire w_dff_B_U0OOsFzQ1_0;
	wire w_dff_B_Fk7TrJzz6_0;
	wire w_dff_B_NHXjAi4F9_0;
	wire w_dff_A_66KJWVwp8_0;
	wire w_dff_B_UFlG5cKM3_1;
	wire w_dff_A_AS70YKql5_0;
	wire w_dff_B_QE8FytI96_1;
	wire w_dff_B_FhiAzXBB6_1;
	wire w_dff_B_g1TD5Row9_1;
	wire w_dff_B_JEPeCu9J0_1;
	wire w_dff_B_ZG2jwuz38_0;
	wire w_dff_B_zQ4MytPc7_1;
	wire w_dff_B_jyM7J1ZV9_0;
	wire w_dff_A_7RobHvig9_0;
	wire w_dff_A_jNOtSQy00_0;
	wire w_dff_A_3vlUtqyv9_0;
	wire w_dff_A_XwwuUsln0_0;
	wire w_dff_B_MvjSQb1U2_0;
	wire w_dff_A_9cjRjcFv5_0;
	wire w_dff_B_Ut5Bnd300_0;
	wire w_dff_B_bhGgs7uv5_0;
	wire w_dff_B_UFJ4mJEx3_0;
	wire w_dff_B_z9LDfLam6_0;
	wire w_dff_B_pi18C67K0_0;
	wire w_dff_B_58hRtFy36_0;
	wire w_dff_B_s7n5lhpd8_0;
	wire w_dff_B_dtPFA2SD7_0;
	wire w_dff_B_9bPkADha1_0;
	wire w_dff_B_Yh1o87DF4_0;
	wire w_dff_B_q9XTkk1d1_0;
	wire w_dff_B_GU6O5mJw0_0;
	wire w_dff_B_QNxPHZKg8_0;
	wire w_dff_B_Wc5IvLvh3_0;
	wire w_dff_B_FlTFRELI9_0;
	wire w_dff_B_aEuozjhT5_0;
	wire w_dff_B_I2ermMkl7_0;
	wire w_dff_B_2C2LaIa98_0;
	wire w_dff_B_K8TlxGVZ4_0;
	wire w_dff_B_vTLCDkIb0_0;
	wire w_dff_B_Gpl903cN2_0;
	wire w_dff_B_OtsaWbz08_0;
	wire w_dff_B_ZhQRZYta7_0;
	wire w_dff_B_ofde5ZOi0_0;
	wire w_dff_B_b4G56N331_0;
	wire w_dff_B_uPHCEmRC4_0;
	wire w_dff_B_F12qWcb15_0;
	wire w_dff_B_nU5g4WdW9_0;
	wire w_dff_B_X5lc8ERA2_0;
	wire w_dff_B_E4BG8Ayw5_0;
	wire w_dff_B_IOi2av3N4_0;
	wire w_dff_B_DZcULegl0_0;
	wire w_dff_B_Qx7oNdWy9_0;
	wire w_dff_B_0ztLduFz5_0;
	wire w_dff_B_nsPRMNxz1_0;
	wire w_dff_B_Ih13jZBk8_0;
	wire w_dff_B_skpGvuxw4_2;
	wire w_dff_B_G5rMUXF48_2;
	wire w_dff_B_pc46jYw56_2;
	wire w_dff_B_xiEtWRdJ3_0;
	wire w_dff_B_0QXWl8xb1_0;
	wire w_dff_B_axFCVXAq9_0;
	wire w_dff_B_q14bpZdM0_0;
	wire w_dff_B_xKfuQ16J7_0;
	wire w_dff_B_XW5a9qpS3_0;
	wire w_dff_B_qoNtuyfN5_0;
	wire w_dff_B_lo5eZZYj4_0;
	wire w_dff_B_wR7cML9x6_0;
	wire w_dff_B_rw2nfGOk0_0;
	wire w_dff_B_sZjXSQc00_0;
	wire w_dff_B_1MYmZ2Hh8_0;
	wire w_dff_B_vZJ4MQiT0_0;
	wire w_dff_B_zU4wzDf07_0;
	wire w_dff_B_2rdPzQxt5_0;
	wire w_dff_B_wsrvTRFU1_0;
	wire w_dff_B_bKng4ZYj7_0;
	wire w_dff_B_7sDRp8Pe6_0;
	wire w_dff_B_jcLLwElZ8_0;
	wire w_dff_B_X3W3I4CG0_0;
	wire w_dff_B_bxdHV3Tb7_0;
	wire w_dff_B_Y7YCJUoX5_0;
	wire w_dff_B_qlpAoWjL2_0;
	wire w_dff_B_7MN0tEj44_0;
	wire w_dff_B_xl0qGUAI6_0;
	wire w_dff_B_rM0t2XlX6_0;
	wire w_dff_B_FAavZQ1G2_0;
	wire w_dff_B_4j68Ncvl4_0;
	wire w_dff_B_vwzFit9Q6_0;
	wire w_dff_B_Hj7tOlfS8_0;
	wire w_dff_B_nBFTz95a8_0;
	wire w_dff_B_CiOblOqN6_0;
	wire w_dff_B_bOm6xuOr3_0;
	wire w_dff_B_uwUSbe004_0;
	wire w_dff_A_dkRHlgvt0_2;
	wire w_dff_A_ZgzYrzSU2_2;
	wire w_dff_B_qYJGFmw80_0;
	wire w_dff_B_0xGmt1ef9_0;
	wire w_dff_B_WlUJvoLS4_0;
	wire w_dff_B_lRZuuHgY9_0;
	wire w_dff_B_f1jKh4Xk8_0;
	wire w_dff_B_hnUKu0HQ6_0;
	wire w_dff_B_jFCmLIkr3_0;
	wire w_dff_B_zEnMY9dx2_0;
	wire w_dff_B_Tg6LPpdP0_0;
	wire w_dff_B_gP81Hn0u5_0;
	wire w_dff_B_o0wuvb1b9_0;
	wire w_dff_B_IIGwLfn26_0;
	wire w_dff_B_ohzHHHUB2_0;
	wire w_dff_B_q77aGSrk7_0;
	wire w_dff_B_t94d85kX8_0;
	wire w_dff_B_5jWzyvJG7_0;
	wire w_dff_B_NypKMHDv5_0;
	wire w_dff_B_PoebvJ2P8_0;
	wire w_dff_B_8fRSbgka8_0;
	wire w_dff_B_UmrBnTNH2_0;
	wire w_dff_B_v9cFAZLn5_0;
	wire w_dff_B_zqDTnKjs4_0;
	wire w_dff_B_4vle1Qcn3_0;
	wire w_dff_B_k16y28oq0_0;
	wire w_dff_B_uv1yIhmW3_0;
	wire w_dff_B_2jKjYMzD8_0;
	wire w_dff_B_ywD1xsZl0_0;
	wire w_dff_B_Z0ns3pPN8_0;
	wire w_dff_B_g4KtRWBn3_0;
	wire w_dff_B_1DRwYKOB2_0;
	wire w_dff_B_77g5Gz7d0_0;
	wire w_dff_B_LhUW3Ydi0_0;
	wire w_dff_B_Izl0K9OX4_0;
	wire w_dff_B_zwPJdQEF4_2;
	wire w_dff_B_eXvMRe1b0_2;
	wire w_dff_B_SYbYFckq7_2;
	wire w_dff_B_8a1wdmuh6_0;
	wire w_dff_B_LcHVNjN99_0;
	wire w_dff_B_18MsEnw70_0;
	wire w_dff_B_HVS95MvC7_0;
	wire w_dff_B_GGddtJoi9_0;
	wire w_dff_B_fal9RzBR4_0;
	wire w_dff_B_L6FrlyfN6_0;
	wire w_dff_B_OxoekeWa1_0;
	wire w_dff_B_2Kc6ThxV7_0;
	wire w_dff_B_YI2taczn0_0;
	wire w_dff_B_Fj3NFwt24_0;
	wire w_dff_B_uNgBiU0g9_0;
	wire w_dff_B_vRurAE3o3_0;
	wire w_dff_B_UrgNl8Ee5_0;
	wire w_dff_B_OftxRVgy5_0;
	wire w_dff_B_aiw9eHOp9_0;
	wire w_dff_B_jlLPp9Vx4_0;
	wire w_dff_B_mOQjkljC0_2;
	wire w_dff_B_zoqcHgRF3_2;
	wire w_dff_B_0gLVztIc0_2;
	wire w_dff_A_YZB8mdmT1_2;
	wire w_dff_A_WCC2ZLwE1_2;
	wire w_dff_B_pBf9AXCt4_0;
	wire w_dff_B_yMNdH2HB6_0;
	wire w_dff_B_hjkvwDCd0_0;
	wire w_dff_B_AcGrsj9n5_0;
	wire w_dff_B_xrmpRsv10_0;
	wire w_dff_B_3dgRN1Um7_0;
	wire w_dff_B_mWlX1zib4_0;
	wire w_dff_B_XBWApV9K6_0;
	wire w_dff_B_QfUT9LvJ3_0;
	wire w_dff_B_ciLEGZ418_0;
	wire w_dff_B_AlFxUvzv6_0;
	wire w_dff_B_HeI2mYQu0_0;
	wire w_dff_B_MziJslA06_0;
	wire w_dff_B_VVs6pJHk9_0;
	wire w_dff_B_pcFZ3uXV4_0;
	wire w_dff_B_vi4xFXql7_0;
	wire w_dff_B_cQ9zOYqq2_2;
	wire w_dff_B_QWTeqsKZ6_2;
	wire w_dff_B_jN6unUfh7_2;
	wire w_dff_B_Ow9FdZNy8_0;
	wire w_dff_B_YGPUoZBU2_0;
	wire w_dff_B_rNED4cpP6_0;
	wire w_dff_B_ttIkTcL76_0;
	wire w_dff_B_83KDtTui9_0;
	wire w_dff_B_hUY0udmf3_0;
	wire w_dff_B_hEznpjwG7_0;
	wire w_dff_B_wcQSsuKc3_0;
	wire w_dff_B_RcKiMlGo0_0;
	wire w_dff_B_7EqxGuFx2_0;
	wire w_dff_B_v6JDwg0L9_0;
	wire w_dff_B_OKspzJNu7_0;
	wire w_dff_B_APgepRj83_0;
	wire w_dff_B_NgUwY59h6_0;
	wire w_dff_B_bdxp7AcU3_0;
	wire w_dff_B_fis0PEsW9_0;
	wire w_dff_A_y1kofuVU5_0;
	wire w_dff_A_bZhs7fic4_0;
	wire w_dff_A_H5oXzNSF8_0;
	wire w_dff_A_H3FSjW8n1_0;
	wire w_dff_A_ZlmiawB56_0;
	wire w_dff_A_qp4LGAap9_1;
	wire w_dff_B_agRsUJDf4_0;
	wire w_dff_B_ZKwsOfHf5_0;
	wire w_dff_B_V3uCsFml0_0;
	wire w_dff_B_SQHPePvO3_0;
	wire w_dff_B_TDWBnvTb7_0;
	wire w_dff_B_xr8B8iLi1_0;
	wire w_dff_B_12MprNB32_0;
	wire w_dff_B_5aEKSf3m8_0;
	wire w_dff_B_RkBc9UVD7_0;
	wire w_dff_B_3hqkoWtI1_0;
	wire w_dff_B_sIJUYtiF0_0;
	wire w_dff_B_6nGtx7Bc5_0;
	wire w_dff_B_7UyEt8Gt1_0;
	wire w_dff_B_wjNWKAFj7_0;
	wire w_dff_B_EBRwlS4T6_0;
	wire w_dff_B_V85onpWG4_0;
	wire w_dff_B_294IO92r3_0;
	wire w_dff_B_d0YDtxRG3_0;
	wire w_dff_B_LAXbZkme6_0;
	wire w_dff_B_wMMrjdzF3_0;
	wire w_dff_B_Tv3AhgpP7_0;
	wire w_dff_B_cbFc7pic9_0;
	wire w_dff_B_8GxulXDB4_0;
	wire w_dff_B_dM2C0V3V7_0;
	wire w_dff_B_g5vUnsM18_0;
	wire w_dff_B_KOhDaaUz2_0;
	wire w_dff_B_O3LfvDXL3_0;
	wire w_dff_B_xyw0L8UL6_0;
	wire w_dff_B_AAfTTh1A4_0;
	wire w_dff_B_ViAWt65H6_0;
	wire w_dff_B_MkvfGRyR6_0;
	wire w_dff_B_cssxxx1u9_0;
	wire w_dff_B_C1YjVtUI7_0;
	wire w_dff_B_FfSLbWuY1_0;
	wire w_dff_A_7OW5y9l72_0;
	wire w_dff_A_l4jMXvw94_1;
	wire w_dff_A_PHBE6jlE2_0;
	wire w_dff_A_o45GCSCM4_1;
	wire w_dff_B_gVdEtFX19_0;
	wire w_dff_B_Ba0686lj8_0;
	wire w_dff_B_qsfq8MbL0_0;
	wire w_dff_B_KfOZ8Leu1_0;
	wire w_dff_B_vj1MW3nq9_0;
	wire w_dff_B_uS61SSR74_0;
	wire w_dff_B_C9ky7vOl1_0;
	wire w_dff_B_R2CeI2Jc3_0;
	wire w_dff_B_kMat4lox3_0;
	wire w_dff_B_Rdg9HmST9_0;
	wire w_dff_B_JhlFtZgN5_0;
	wire w_dff_B_3CmVi0QK0_0;
	wire w_dff_B_yBsCen7m0_0;
	wire w_dff_B_V5ZrAPuN6_0;
	wire w_dff_B_xyVYWRYK9_0;
	wire w_dff_B_s55vGzNJ3_0;
	wire w_dff_B_UhZT5YK20_0;
	wire w_dff_B_KImXdIga2_0;
	wire w_dff_A_RQQIh7vn0_0;
	wire w_dff_B_ZmFCOJy13_0;
	wire w_dff_B_JbI7LX1H9_0;
	wire w_dff_B_LMESYq2w5_0;
	wire w_dff_B_8hAu5rcr9_0;
	wire w_dff_B_a35Fo7iV8_0;
	wire w_dff_B_t3yeZgE34_0;
	wire w_dff_B_4xMKYaLx1_0;
	wire w_dff_B_7PEwpT1r2_0;
	wire w_dff_B_zu2voKMB9_0;
	wire w_dff_B_QUWFna4i9_0;
	wire w_dff_B_5Bds0IZW2_0;
	wire w_dff_B_CIdUXag39_0;
	wire w_dff_B_vmB6lXpv2_0;
	wire w_dff_B_SWDiZyBP0_0;
	wire w_dff_B_ccTWhB2x9_0;
	wire w_dff_B_OKMz4WVo9_0;
	wire w_dff_B_SGUhAMb97_2;
	wire w_dff_B_IFxkz3Y08_2;
	wire w_dff_B_mLxJD7f59_2;
	wire w_dff_B_I9S9Xa0x6_0;
	wire w_dff_B_TEtLmidp4_0;
	wire w_dff_B_96xzDBIs6_0;
	wire w_dff_B_LHpPA1Wf7_0;
	wire w_dff_B_cFYJGVhW7_0;
	wire w_dff_B_RMXQNnOq9_0;
	wire w_dff_B_L4qQWu689_0;
	wire w_dff_B_kmG4DrdP9_0;
	wire w_dff_B_AQUBKamq2_0;
	wire w_dff_B_E1ByTHYL4_0;
	wire w_dff_B_62huH6Nq1_0;
	wire w_dff_B_3epKLyCT9_1;
	wire w_dff_B_tYfQVzEI9_1;
	wire w_dff_B_17aiqjGc4_0;
	wire w_dff_B_dSejLMxx2_0;
	wire w_dff_B_nek2bSjm6_0;
	wire w_dff_B_IX8EgRQH2_0;
	wire w_dff_B_xbHkbq0I8_0;
	wire w_dff_B_UnPCY6Db0_0;
	wire w_dff_B_dihwUXjS5_0;
	wire w_dff_B_gCnKLI5i2_0;
	wire w_dff_B_9CBb133i7_0;
	wire w_dff_B_jGhB8Mmf3_0;
	wire w_dff_B_p23c7erm3_0;
	wire w_dff_B_kWzdq82a2_0;
	wire w_dff_B_0TVAYJPD2_1;
	wire w_dff_B_AKDvo7Ba7_1;
	wire w_dff_B_2wflkQor3_0;
	wire w_dff_B_YdcdSCpG9_1;
	wire w_dff_B_09Q8taF07_0;
	wire w_dff_B_zEuw58Vs5_0;
	wire w_dff_B_qtFTJ7YN5_0;
	wire w_dff_B_0rmgxtLS1_0;
	wire w_dff_B_dYrKAl9E6_0;
	wire w_dff_B_EJQTvFzO7_0;
	wire w_dff_B_BiTMPZqi6_0;
	wire w_dff_B_dqkJ1ncm3_0;
	wire w_dff_B_fmMG05vF3_0;
	wire w_dff_B_AtuYmRCA6_0;
	wire w_dff_B_IFHSWs6i4_0;
	wire w_dff_B_d8G8CC2Z5_0;
	wire w_dff_B_aj8h4fjM8_0;
	wire w_dff_B_GURgKlrr4_0;
	wire w_dff_B_qCbrYods6_0;
	wire w_dff_B_lXYnlb5b3_0;
	wire w_dff_B_SAWpM6fQ5_0;
	wire w_dff_B_MAJmmH5t1_2;
	wire w_dff_B_50RCKjQP1_2;
	wire w_dff_B_cFW4n59S5_2;
	wire w_dff_B_LIqQJyqB7_0;
	wire w_dff_B_154GA88v8_0;
	wire w_dff_B_scoLKQWQ0_0;
	wire w_dff_B_H5TTfpr02_0;
	wire w_dff_B_WVwjElLV1_0;
	wire w_dff_B_r8tieEPh9_0;
	wire w_dff_B_xGpnWdoj3_0;
	wire w_dff_B_fKnP5ZTG4_0;
	wire w_dff_B_zpKo9Ccc5_0;
	wire w_dff_B_vJHcfLve3_0;
	wire w_dff_B_3J5EAi6i6_0;
	wire w_dff_B_1QghGSTZ5_0;
	wire w_dff_B_odjM5rvn3_1;
	wire w_dff_B_h2p3nyxB3_1;
	wire w_dff_A_sUW6gcWQ9_1;
	wire w_dff_B_quMq9nbg5_1;
	wire w_dff_B_sQCErxne2_1;
	wire w_dff_B_4EsNKvRA1_1;
	wire w_dff_B_l8XGactB8_1;
	wire w_dff_B_xlzh8Ftl9_1;
	wire w_dff_B_c0G0nXkd0_1;
	wire w_dff_B_kZeNUo0G9_1;
	wire w_dff_B_3nxzTJoj7_1;
	wire w_dff_B_kOVmyXKi0_1;
	wire w_dff_B_udGqIPxm7_1;
	wire w_dff_B_IMe2uchO1_0;
	wire w_dff_B_ZReIIt4W8_0;
	wire w_dff_B_gw0ZtexQ4_0;
	wire w_dff_B_7sCawKEX8_0;
	wire w_dff_B_8Ui3d48h8_0;
	wire w_dff_B_mSSl9zLJ1_0;
	wire w_dff_B_sNTc23mc7_0;
	wire w_dff_B_9oJ52C180_0;
	wire w_dff_B_MqaT0KJJ5_0;
	wire w_dff_B_AQXaAoau3_0;
	wire w_dff_B_xAXaJ5Ik2_0;
	wire w_dff_B_pxnY8ccd7_0;
	wire w_dff_B_7PZywBut2_0;
	wire w_dff_B_Nj5vdTif5_1;
	wire w_dff_B_StV1voEx0_1;
	wire w_dff_B_gG2uUQz25_0;
	wire w_dff_B_ETgeSkvN4_1;
	wire w_dff_B_ixPsF8PX5_1;
	wire w_dff_B_4qSErFbZ5_1;
	wire w_dff_B_55kHWLt07_1;
	wire w_dff_B_PdoLO2ui9_1;
	wire w_dff_B_Uo6Ck4sD7_1;
	wire w_dff_B_Us86aFVR4_1;
	wire w_dff_B_mXczXv536_1;
	wire w_dff_B_sf9LzMDB0_1;
	wire w_dff_B_c7gxiID30_1;
	wire w_dff_B_TffRr9w90_1;
	wire w_dff_B_3c94yB1b0_1;
	wire w_dff_B_fpTMEgEi4_1;
	wire w_dff_B_eeznKk6L0_1;
	wire w_dff_B_ConUEDM16_1;
	wire w_dff_B_qsOYPMWr4_1;
	wire w_dff_B_VbZ4XuZP0_1;
	wire w_dff_B_P1WrViCA7_1;
	wire w_dff_B_iBWYpPYu7_1;
	wire w_dff_B_e5HQDqVp5_1;
	wire w_dff_A_sAzoij892_1;
	wire w_dff_A_6FYOdVxK6_1;
	wire w_dff_A_zNPmARhV5_1;
	wire w_dff_A_77DusoA61_1;
	wire w_dff_A_aLhqdgZU3_1;
	wire w_dff_A_Vgr5vevl1_1;
	wire w_dff_A_vb2M1OE24_1;
	wire w_dff_A_Ck6oxcC35_1;
	wire w_dff_A_RBGRznVJ7_1;
	wire w_dff_A_zeRLM1kf4_1;
	wire w_dff_A_BmECUsk12_1;
	wire w_dff_A_Gu5nNEwY7_1;
	wire w_dff_A_FBNMLUe16_1;
	wire w_dff_A_nDfkBzeK5_2;
	wire w_dff_A_9RebKp3i9_2;
	wire w_dff_A_gNbujCMb7_2;
	wire w_dff_A_aLH5F6Tt6_2;
	wire w_dff_A_Pimr12Am7_2;
	wire w_dff_A_ElQe45RG5_2;
	wire w_dff_A_2s2YT0uI2_2;
	wire w_dff_A_btSBnyTP2_2;
	wire w_dff_A_BPkgQXW11_2;
	wire w_dff_A_SQAQH26V5_2;
	wire w_dff_A_iNS2XPFK1_2;
	wire w_dff_A_L5frsO004_2;
	wire w_dff_B_9pLJ2O540_0;
	wire w_dff_B_cPWzW0kk4_0;
	wire w_dff_B_Xe9zhxh66_0;
	wire w_dff_B_7iguyQVm5_0;
	wire w_dff_B_RNLWmLJJ1_0;
	wire w_dff_B_RHF8iTjG5_0;
	wire w_dff_B_pQW52dv74_0;
	wire w_dff_B_7y1vDWQp2_0;
	wire w_dff_B_5vVcP5lv2_0;
	wire w_dff_B_Bm4FV72o3_0;
	wire w_dff_B_j0If32eX7_0;
	wire w_dff_B_CjZodt2l6_0;
	wire w_dff_B_DLpxs9L61_0;
	wire w_dff_B_yqIm284c6_0;
	wire w_dff_B_Bbjyg1EH7_0;
	wire w_dff_B_RyyWYobz7_0;
	wire w_dff_B_powhZxEO6_0;
	wire w_dff_B_TvkVAIn21_2;
	wire w_dff_B_14vpiaKB5_2;
	wire w_dff_B_7lMbWqIo5_2;
	wire w_dff_B_B84uG7bX8_0;
	wire w_dff_B_QjU99fHA3_0;
	wire w_dff_B_ucHpOF5h4_0;
	wire w_dff_B_Ym1Q9bcb1_0;
	wire w_dff_B_ncHijzMR4_0;
	wire w_dff_B_y0ZkcAHI7_0;
	wire w_dff_B_pY4kvoBt2_0;
	wire w_dff_B_TvlAC35e3_0;
	wire w_dff_B_Mlmerch91_0;
	wire w_dff_B_pehWNw4f6_0;
	wire w_dff_B_KrP1yuHQ9_0;
	wire w_dff_B_marBBmw55_0;
	wire w_dff_B_HXk0kOAM5_1;
	wire w_dff_B_uKr8CYGs6_1;
	wire w_dff_A_aeevJOVS0_0;
	wire w_dff_A_vEyg9jp74_0;
	wire w_dff_A_X6QMuLAm1_0;
	wire w_dff_A_q9i9WFuA3_0;
	wire w_dff_A_SBknElrP1_2;
	wire w_dff_A_YlD1YxIp1_2;
	wire w_dff_A_H1qLvIgG7_1;
	wire w_dff_A_xsOeO7oV5_1;
	wire w_dff_A_ylCN2lH88_1;
	wire w_dff_A_8yOW4PUZ0_1;
	wire w_dff_A_y7CO8UH03_1;
	wire w_dff_A_qzHdiVqZ7_1;
	wire w_dff_A_EnI1yzei1_1;
	wire w_dff_A_UQoh7LGe2_1;
	wire w_dff_A_wOf1Cfte0_2;
	wire w_dff_A_N3h0DbEd0_2;
	wire w_dff_A_wRFxOKzz0_2;
	wire w_dff_A_a3B1miSq9_2;
	wire w_dff_B_qXzrlhWH2_3;
	wire w_dff_A_qNY8BP3v7_0;
	wire w_dff_A_UXajs5TU9_0;
	wire w_dff_A_aPAD6atK6_0;
	wire w_dff_A_WBxupp7Q1_0;
	wire w_dff_A_n4a7JNKr9_0;
	wire w_dff_A_sTj0VN4c4_0;
	wire w_dff_A_e0JYmab19_0;
	wire w_dff_A_wDe8DPcc0_0;
	wire w_dff_A_SqI2yV546_1;
	wire w_dff_A_3Vi918I32_1;
	wire w_dff_A_gU6XlNYE1_1;
	wire w_dff_A_H5bf7n1u2_0;
	wire w_dff_A_ITNR949C7_1;
	wire w_dff_B_S9J7nqW47_0;
	wire w_dff_B_qSC0jK4B7_0;
	wire w_dff_B_74MEXcp64_0;
	wire w_dff_B_XNwsMo0y7_0;
	wire w_dff_B_yNmVYCKB9_0;
	wire w_dff_B_9U6ylI2J2_0;
	wire w_dff_B_XdZik20e3_0;
	wire w_dff_B_vMziX8uU1_0;
	wire w_dff_B_r7ZKzvHx2_0;
	wire w_dff_B_9DeFJJmY7_0;
	wire w_dff_B_WPzhHrAb9_0;
	wire w_dff_B_PqJq7Mgt4_0;
	wire w_dff_B_XGAPpf743_0;
	wire w_dff_B_Nm4EO94P3_1;
	wire w_dff_B_vNPPy6ed3_1;
	wire w_dff_B_jFICK1UL1_3;
	wire w_dff_B_rUp8ULsw4_3;
	wire w_dff_A_BsgYYTw75_1;
	wire w_dff_B_Bb8vETym4_0;
	wire w_dff_B_GertBESm2_3;
	wire w_dff_B_SCzYglrG4_1;
	wire w_dff_A_fYU173FL6_0;
	wire w_dff_A_tjHVlKCN6_1;
	wire w_dff_A_383ZEy6I1_0;
	wire w_dff_A_ju5dP4BX9_1;
	wire w_dff_A_y0ZRGQTF0_0;
	wire w_dff_A_sKZThTtb6_0;
	wire w_dff_A_q4R3ZE6d8_0;
	wire w_dff_A_ZCPtQnaG6_0;
	wire w_dff_A_so03MYB81_0;
	wire w_dff_A_a9J6yTKK2_1;
	wire w_dff_A_ZJQjY5Xt2_1;
	wire w_dff_A_9IoQ8PG53_1;
	wire w_dff_A_HjS9J4X52_1;
	wire w_dff_A_Fl8KFQKn2_1;
	wire w_dff_A_2NRd1JdT9_1;
	wire w_dff_B_n7cutjcq9_0;
	wire w_dff_B_yptsFa2p8_0;
	wire w_dff_B_JRsmjG7t2_0;
	wire w_dff_B_dZSZV8M57_0;
	wire w_dff_B_BSzS8LU70_0;
	wire w_dff_B_JVHhIBho1_0;
	wire w_dff_B_plbfaqeX3_0;
	wire w_dff_B_7eWOYkPS2_0;
	wire w_dff_B_gKVHduvz1_0;
	wire w_dff_B_JV9dXuVZ5_0;
	wire w_dff_B_jeGq64yM1_0;
	wire w_dff_B_9pGaziJu7_0;
	wire w_dff_B_aV5fYulz2_0;
	wire w_dff_B_sLKrHYsW7_0;
	wire w_dff_B_quMSMqcC0_0;
	wire w_dff_B_ZUaMsc4b2_0;
	wire w_dff_B_AM3vBMxa2_0;
	wire w_dff_B_nXPPc2nM8_0;
	wire w_dff_B_wnoB62px8_2;
	wire w_dff_B_tpfWh4pm0_2;
	wire w_dff_B_YXrldbBk9_2;
	wire w_dff_B_7FRchA6w4_0;
	wire w_dff_B_4RhB5ZPW2_0;
	wire w_dff_B_7D0ylB5Q9_0;
	wire w_dff_B_rEAdzYBT9_0;
	wire w_dff_B_AhbaE4kP1_0;
	wire w_dff_B_u1HQjpXg7_0;
	wire w_dff_B_bmMGZWz43_0;
	wire w_dff_B_IQ4cwdyf5_0;
	wire w_dff_B_3Of4yyyn8_0;
	wire w_dff_B_ZRG9BTvk1_0;
	wire w_dff_B_WMfun7bd3_0;
	wire w_dff_B_aH6Nh85K3_0;
	wire w_dff_B_BWNbPEii0_0;
	wire w_dff_B_BKEKWhze3_1;
	wire w_dff_B_FE6uwSmS0_1;
	wire w_dff_A_7EUgJjEv4_1;
	wire w_dff_A_BrrDWsJJ5_0;
	wire w_dff_B_k7ccmGjA3_2;
	wire w_dff_B_BCyhDCpA1_0;
	wire w_dff_B_JbPk5Cbw3_0;
	wire w_dff_B_t0QenPJK3_0;
	wire w_dff_B_enuUWqnO6_0;
	wire w_dff_A_FMfDTZPu3_0;
	wire w_dff_A_mAXDZyS17_0;
	wire w_dff_A_d7HrMQip3_0;
	wire w_dff_A_6B2gmyQI5_0;
	wire w_dff_A_lCuEXdLn1_0;
	wire w_dff_A_LqY3TKdd0_0;
	wire w_dff_A_jq7VWQt19_0;
	wire w_dff_A_vpdtxn4N0_0;
	wire w_dff_A_hGTaNu9B9_0;
	wire w_dff_A_G8LGNIc74_0;
	wire w_dff_A_cDwjwPSq8_0;
	wire w_dff_A_NB5iNk0F7_0;
	wire w_dff_A_1J23STzd1_0;
	wire w_dff_A_sIKpZPM87_0;
	wire w_dff_A_xo8iiHrd0_0;
	wire w_dff_A_fqc6Redu2_0;
	wire w_dff_A_8apAwvBr9_0;
	wire w_dff_A_Myua4Nl51_0;
	wire w_dff_A_XOvFG1JA5_0;
	wire w_dff_A_Zh3Fzkn12_0;
	wire w_dff_A_4cCoBgTJ8_1;
	wire w_dff_A_q30IOs7B4_1;
	wire w_dff_A_0YA5gX3L0_1;
	wire w_dff_A_tA6W320N7_1;
	wire w_dff_A_G7C3MKLi5_1;
	wire w_dff_A_mibvx99g4_1;
	wire w_dff_A_B163nOEO9_1;
	wire w_dff_A_B6nQ4l5Q2_1;
	wire w_dff_A_uvpUTQee1_1;
	wire w_dff_B_QB6mvxpj1_0;
	wire w_dff_B_bXm5ay248_0;
	wire w_dff_B_A0CdZTO27_0;
	wire w_dff_B_DMr4WauW9_0;
	wire w_dff_B_inQ3U82g4_0;
	wire w_dff_B_aYmgZKAm5_0;
	wire w_dff_B_KElNYV6G7_0;
	wire w_dff_B_DBi65DCa4_0;
	wire w_dff_B_VY6FUyUR8_0;
	wire w_dff_B_U2snLKEJ8_0;
	wire w_dff_B_NxDyucTm8_0;
	wire w_dff_B_5R5KWFjg0_0;
	wire w_dff_B_JUKEnXWI7_0;
	wire w_dff_B_lhXixDxu4_0;
	wire w_dff_B_2j8GxOw91_0;
	wire w_dff_B_20Y1p8ix0_0;
	wire w_dff_B_P1l3ehr71_1;
	wire w_dff_B_9G85qHLp6_1;
	wire w_dff_A_frt58SoM2_0;
	wire w_dff_A_OYaMXLGe7_2;
	wire w_dff_A_YKKmtzwo8_2;
	wire w_dff_A_LGVtW3Qv9_2;
	wire w_dff_A_PvOiRHAm7_2;
	wire w_dff_B_V0ZC5LCV6_1;
	wire w_dff_B_F36k1EPQ8_1;
	wire w_dff_B_zTMLTtux5_1;
	wire w_dff_B_4RvYDFRq3_1;
	wire w_dff_B_Uw8cvXCJ3_1;
	wire w_dff_B_KyJLUTO75_1;
	wire w_dff_B_thd4XTy23_1;
	wire w_dff_B_TG5KVz8b0_1;
	wire w_dff_B_Jbi5ZFtY8_1;
	wire w_dff_B_ErAA75Sg3_1;
	wire w_dff_B_2xvbEX6b6_1;
	wire w_dff_B_rBz9tB1n5_1;
	wire w_dff_B_xo2Xg6bR2_1;
	wire w_dff_B_2TknPHmb6_1;
	wire w_dff_B_4BqlQqfc9_1;
	wire w_dff_B_5knzVkgt4_1;
	wire w_dff_B_nyszu3Qx9_1;
	wire w_dff_B_PSye6bXg7_1;
	wire w_dff_B_yZEvMHkQ1_0;
	wire w_dff_A_bDtXZSfF2_1;
	wire w_dff_A_aZsRZRzc4_1;
	wire w_dff_A_m6tBuxuy5_1;
	wire w_dff_A_LyJqcdhE2_1;
	wire w_dff_A_XQ85SI904_1;
	wire w_dff_A_KUzeLFZw3_1;
	wire w_dff_B_nm6Aqo8B0_3;
	wire w_dff_B_iP6ndz3S4_3;
	wire w_dff_B_CpQk12DH3_3;
	wire w_dff_B_3zTcJTIs9_3;
	wire w_dff_B_hPJG0ldp5_2;
	wire w_dff_B_GP2YH0ms9_2;
	wire w_dff_B_mWMwWwPY5_2;
	wire w_dff_B_vwcFlwia3_2;
	wire w_dff_B_QYKlooOo9_2;
	wire w_dff_B_eTDh0uSx2_2;
	wire w_dff_B_VN8rMfKo1_2;
	wire w_dff_B_RbRQ8xPU8_2;
	wire w_dff_B_MVJDqufb2_2;
	wire w_dff_A_HLAl1M521_1;
	wire w_dff_A_xFXK0hL58_1;
	wire w_dff_A_VoHkmlRv2_1;
	wire w_dff_A_PssrBKtE0_2;
	wire w_dff_A_uE9d4O748_2;
	wire w_dff_A_ZDayzo5r4_2;
	wire w_dff_A_PRChFjBw1_2;
	wire w_dff_A_05wwoAWZ0_0;
	wire w_dff_A_CeJleYnU5_0;
	wire w_dff_A_KzdNH0DK9_0;
	wire w_dff_A_oieLvGfZ1_0;
	wire w_dff_A_0FC9zjOJ3_0;
	wire w_dff_A_h5iRJ6oW1_0;
	wire w_dff_A_rCFMe4uN1_0;
	wire w_dff_A_PKfuQANw6_0;
	wire w_dff_A_oKPUfezU1_0;
	wire w_dff_A_UXYtXNr46_0;
	wire w_dff_A_dhsvvXga0_0;
	wire w_dff_A_W1gUI3au0_0;
	wire w_dff_A_LoCCPFDQ2_0;
	wire w_dff_A_njKGqq1g9_1;
	wire w_dff_A_bzzNAAMX7_1;
	wire w_dff_A_DeQWqwRF8_1;
	wire w_dff_A_Hulc4xtm9_1;
	wire w_dff_A_vtSH9Vbn1_1;
	wire w_dff_A_NWZp0gGh3_1;
	wire w_dff_A_Xu5BlIp72_1;
	wire w_dff_B_hWyTCKRT3_1;
	wire w_dff_B_VDLvyCjj0_1;
	wire w_dff_B_sbds70jh7_1;
	wire w_dff_B_xVKvmOMW7_1;
	wire w_dff_B_NAl70N4K8_1;
	wire w_dff_B_5xB1GOzx7_1;
	wire w_dff_B_AoYBY6MI2_1;
	wire w_dff_B_TtEPmjQ46_1;
	wire w_dff_B_clzf3T6G8_1;
	wire w_dff_B_cFeYhvnw4_1;
	wire w_dff_B_CJ9UndW83_1;
	wire w_dff_B_N5MmGJLS4_1;
	wire w_dff_B_8DsBHhks9_1;
	wire w_dff_B_guLETHEL6_1;
	wire w_dff_B_RO1PxrYt8_1;
	wire w_dff_B_NlmNpPso8_1;
	wire w_dff_B_uTZn3X140_1;
	wire w_dff_B_O590Tvgi3_1;
	wire w_dff_B_pt4Np9lk0_1;
	wire w_dff_B_2fu0Yukz0_1;
	wire w_dff_B_XKFhEpvU7_1;
	wire w_dff_B_X16GS3k32_1;
	wire w_dff_B_lEZqV0FP4_1;
	wire w_dff_B_d00V3A903_1;
	wire w_dff_B_SiQpf2OB4_1;
	wire w_dff_B_37Wt5caT1_1;
	wire w_dff_B_isjrsp5R5_1;
	wire w_dff_B_3Szipj2D7_1;
	wire w_dff_B_2ltHrkJs4_1;
	wire w_dff_B_nZ2gg8PF1_1;
	wire w_dff_B_AxlY0AT22_1;
	wire w_dff_B_sqUS6HAx9_1;
	wire w_dff_B_xiX3QdBV9_1;
	wire w_dff_B_JpiBi7vB6_1;
	wire w_dff_B_LESUyLpb0_1;
	wire w_dff_B_9zXaKAsG7_1;
	wire w_dff_B_BYPKNXFo4_1;
	wire w_dff_B_bUlMydrC4_1;
	wire w_dff_B_Oyc7erkj0_0;
	wire w_dff_B_3UQXGzYe1_0;
	wire w_dff_B_p9iI1GCm6_0;
	wire w_dff_B_Fv8oce7b2_0;
	wire w_dff_B_xfdXn3gh8_0;
	wire w_dff_B_24RTbt2l6_0;
	wire w_dff_B_T5QHiW5g4_0;
	wire w_dff_B_XUHRBrMY2_0;
	wire w_dff_B_rM8hLnGy8_0;
	wire w_dff_B_8nFpynAk6_0;
	wire w_dff_B_6O0TcsTE8_0;
	wire w_dff_B_1ERHSp2e2_0;
	wire w_dff_B_KgQ5RStM5_0;
	wire w_dff_B_iQkfhazn3_0;
	wire w_dff_B_YxjzLB4X2_0;
	wire w_dff_B_A6trlIz93_0;
	wire w_dff_B_7CFLzJwE9_0;
	wire w_dff_B_Acos7NPE2_0;
	wire w_dff_B_pn9fF3NJ2_0;
	wire w_dff_B_zVkRJpEp9_0;
	wire w_dff_A_gDFl44Nf8_1;
	wire w_dff_A_QK4tJ5KJ2_1;
	wire w_dff_A_WTFoR4Xs3_1;
	wire w_dff_A_WnvQZK9R1_1;
	wire w_dff_A_YYBwUoaC1_1;
	wire w_dff_A_Vv1X4RK16_1;
	wire w_dff_A_6t5wCJPH9_1;
	wire w_dff_A_nloeYeZH8_1;
	wire w_dff_A_Zb1Np2Q13_1;
	wire w_dff_A_hOA9568S6_1;
	wire w_dff_A_iywbZGbf1_1;
	wire w_dff_A_TgEIV9iS0_1;
	wire w_dff_A_y3HvpBwO3_1;
	wire w_dff_A_wr4dtUjX9_1;
	wire w_dff_A_rKVaqn901_2;
	wire w_dff_A_ldK5lY4G6_2;
	wire w_dff_A_681pEa5P3_2;
	wire w_dff_A_XDMjJR8f2_2;
	wire w_dff_A_SwdNfqQS8_2;
	wire w_dff_A_1IUCxP8Q5_2;
	wire w_dff_A_SjRh2TnK2_2;
	wire w_dff_A_wffqRqnD2_2;
	wire w_dff_A_9b4ItQma5_2;
	wire w_dff_A_AJGiieCM9_2;
	wire w_dff_A_Zxi2yntb3_1;
	wire w_dff_A_iW9kNU8j2_1;
	wire w_dff_A_P6fUHoeO5_1;
	wire w_dff_A_YyMhI7br9_1;
	wire w_dff_A_hFiRqPYe5_1;
	wire w_dff_A_9yNuijDT7_1;
	wire w_dff_A_J9s8QZEi9_1;
	wire w_dff_A_5fop84UG1_1;
	wire w_dff_A_ZFi2FESZ2_1;
	wire w_dff_A_oRQ7d04F4_1;
	wire w_dff_A_MsSSaf845_1;
	wire w_dff_A_dsfKY5Mi9_2;
	wire w_dff_B_Jj9PwHD67_3;
	wire w_dff_B_4yw7WmsD5_3;
	wire w_dff_B_z3NZq9r76_3;
	wire w_dff_B_i40G09E43_3;
	wire w_dff_B_BWtFMQnv4_3;
	wire w_dff_B_XABObqKV1_3;
	wire w_dff_A_09hrrOSP0_1;
	wire w_dff_A_ICxSbAIE1_1;
	wire w_dff_A_4bNrqtOu9_1;
	wire w_dff_A_56k5cqEv8_1;
	wire w_dff_A_zei0RHmK3_1;
	wire w_dff_A_rmTAStox6_1;
	wire w_dff_A_LIfvZvJn4_1;
	wire w_dff_A_AoZXPVz36_1;
	wire w_dff_A_6wYzzrQc6_1;
	wire w_dff_A_GJPIIFRs0_1;
	wire w_dff_A_d3nwqLTE2_1;
	wire w_dff_A_AhPdWlgx8_1;
	wire w_dff_A_qeOascDE5_1;
	wire w_dff_A_xjWfmCDl7_1;
	wire w_dff_A_y0oRANoW6_2;
	wire w_dff_A_Kzu7LfBS5_2;
	wire w_dff_A_ePmZYUO09_2;
	wire w_dff_A_6XrdGx970_2;
	wire w_dff_A_9HOSXcbI1_2;
	wire w_dff_A_v7rzEFQq9_2;
	wire w_dff_A_kSD2nT7G3_2;
	wire w_dff_A_taAU0pJb7_2;
	wire w_dff_A_bktD94j34_2;
	wire w_dff_A_S5eA9kuy6_2;
	wire w_dff_A_ODzzS0E23_1;
	wire w_dff_A_NB3Sle5t5_1;
	wire w_dff_A_4yarnEib1_1;
	wire w_dff_A_mzgCjKZS7_1;
	wire w_dff_A_a1MPQaHw2_1;
	wire w_dff_A_vcICGs300_1;
	wire w_dff_A_A7zNrVPA7_1;
	wire w_dff_A_VzlFDMJE1_1;
	wire w_dff_A_60iMxWrC7_1;
	wire w_dff_A_NlNYudBi9_1;
	wire w_dff_A_rbDetDgH9_1;
	wire w_dff_A_SX3MLxt72_2;
	wire w_dff_A_02duTM8P5_2;
	wire w_dff_A_x3tz2ruC5_2;
	wire w_dff_A_4S0qJLoI6_2;
	wire w_dff_B_zmntCGcZ5_3;
	wire w_dff_B_hc2jIxY07_3;
	wire w_dff_B_F7pcUx834_3;
	wire w_dff_B_SwKN3pzG4_3;
	wire w_dff_B_tAHh98pf8_3;
	wire w_dff_B_YW0PqZyk2_3;
	wire w_dff_B_dFN2gYon5_3;
	wire w_dff_A_Ts5zBysZ3_2;
	wire w_dff_A_Jh1PO9Ub9_1;
	wire w_dff_B_zaTCGnqh1_0;
	wire w_dff_B_PAWhwoeG8_0;
	wire w_dff_B_PfRReHWk3_0;
	wire w_dff_B_11Gsk3zY7_0;
	wire w_dff_B_QYWkJchj3_0;
	wire w_dff_B_3vcKBv499_0;
	wire w_dff_B_R3xUY0fx2_0;
	wire w_dff_B_F1YHIbtk3_0;
	wire w_dff_B_MGpcTcz82_0;
	wire w_dff_B_wlON81Hb1_0;
	wire w_dff_B_9LPqMGjj0_0;
	wire w_dff_B_BGfBg8vY1_0;
	wire w_dff_B_eT7K70c91_0;
	wire w_dff_B_1vmN5luf3_0;
	wire w_dff_B_5KAjjyVv9_0;
	wire w_dff_B_08wO1yN45_0;
	wire w_dff_B_IkqgK7uJ3_0;
	wire w_dff_B_Qrk93bQG4_0;
	wire w_dff_B_vy2zsUTI4_0;
	wire w_dff_B_Iw1JI7LE5_0;
	wire w_dff_B_tjMC8laf8_2;
	wire w_dff_B_R6qd8A5o3_2;
	wire w_dff_B_UE8GuEbX6_2;
	wire w_dff_A_Bw91KRzU6_1;
	wire w_dff_A_mFSizQAB5_1;
	wire w_dff_A_Tcv2PsEN5_1;
	wire w_dff_A_U4ln5SHA2_1;
	wire w_dff_A_2Gept2Jo6_1;
	wire w_dff_A_KYNLNk6S2_1;
	wire w_dff_A_UIvSCv7u3_1;
	wire w_dff_A_0f3R6dKC7_1;
	wire w_dff_A_rTCv7y8G5_1;
	wire w_dff_A_NXzMwWYT0_1;
	wire w_dff_A_7Wvx59Ze7_1;
	wire w_dff_A_eF1kCpAo5_1;
	wire w_dff_A_QMvxRlkL1_1;
	wire w_dff_A_WGJbEyxO9_1;
	wire w_dff_A_mVjjwKGe3_2;
	wire w_dff_A_QV4le3QW2_2;
	wire w_dff_A_OpxzFyJB1_2;
	wire w_dff_A_77LzJhx87_2;
	wire w_dff_A_fTlAtfnV2_2;
	wire w_dff_A_XB4NSBmK9_2;
	wire w_dff_A_juotzPK26_2;
	wire w_dff_A_IZVpXalT3_2;
	wire w_dff_A_xS6GkIMI7_2;
	wire w_dff_A_Hwmo3KAh3_2;
	wire w_dff_A_49N5uduP5_1;
	wire w_dff_A_7HfHjDa84_1;
	wire w_dff_A_HXCNTPbk8_1;
	wire w_dff_A_cQmn4lFP1_1;
	wire w_dff_A_pNvcG4Z20_1;
	wire w_dff_A_yZz1gfvG6_1;
	wire w_dff_A_cv2rVsIN5_1;
	wire w_dff_A_4uWKlkDW5_1;
	wire w_dff_A_kPq7nZkf0_1;
	wire w_dff_A_oo9ebvOe3_1;
	wire w_dff_A_kk7zswMP6_1;
	wire w_dff_A_ETtXIzyY5_2;
	wire w_dff_B_HS0SdTZg8_3;
	wire w_dff_B_mhtNTZ0c1_3;
	wire w_dff_B_TbCKI1Rc8_3;
	wire w_dff_B_E5kYmR2p0_3;
	wire w_dff_B_QUibiwm78_3;
	wire w_dff_B_YNwcWui00_3;
	wire w_dff_A_lQRkkn7L6_1;
	wire w_dff_A_A0rPgeOt2_1;
	wire w_dff_A_cVR335jI7_1;
	wire w_dff_A_ffNL8TsJ5_1;
	wire w_dff_A_bxRoYoQg0_1;
	wire w_dff_A_A4WVKjca8_1;
	wire w_dff_A_8ZmzrnB93_1;
	wire w_dff_A_trCIINZ53_1;
	wire w_dff_A_RmHbgeXA6_1;
	wire w_dff_A_muBslIKH4_1;
	wire w_dff_A_DU33Q8n40_1;
	wire w_dff_A_kkTUnA3w1_1;
	wire w_dff_A_u8b5jmpL2_1;
	wire w_dff_A_nLzfCQsM7_1;
	wire w_dff_A_VWpPITbl1_2;
	wire w_dff_A_VriCAyT59_2;
	wire w_dff_A_9veWSEuW6_2;
	wire w_dff_A_ESY4zw8P7_2;
	wire w_dff_A_WrvQyqRj9_2;
	wire w_dff_A_34mx983w1_2;
	wire w_dff_A_sj5abWxI0_2;
	wire w_dff_A_3ZL6epNk0_2;
	wire w_dff_A_ETkTuboE4_2;
	wire w_dff_A_8wZX448Z7_2;
	wire w_dff_A_xWdDvhNX3_1;
	wire w_dff_A_sgeRwZNV6_1;
	wire w_dff_A_yd8p5ipB7_1;
	wire w_dff_A_TXkCGyfc9_1;
	wire w_dff_A_fbiWGzUq3_1;
	wire w_dff_A_1ysmOmuF8_1;
	wire w_dff_A_MNw5UL0q4_1;
	wire w_dff_A_XN9drVBE1_1;
	wire w_dff_A_FOjqyKUo7_1;
	wire w_dff_A_2QcyE6Bd0_1;
	wire w_dff_A_Yw8dhu3K1_1;
	wire w_dff_A_MPqETHIJ7_2;
	wire w_dff_A_MgUL0Bl02_2;
	wire w_dff_A_2s3zZm4n4_2;
	wire w_dff_A_1eiEKxGE0_2;
	wire w_dff_B_d13xtpX31_3;
	wire w_dff_B_46qk7RXw5_3;
	wire w_dff_B_wGWUR7wr4_3;
	wire w_dff_B_bByIaimR9_3;
	wire w_dff_B_7dhOLKPu5_3;
	wire w_dff_B_rXjKCc991_3;
	wire w_dff_B_ybEFOdHf6_3;
	wire w_dff_A_4CRskux41_1;
	wire w_dff_A_SGVINllK6_2;
	wire w_dff_B_WDSJg6To0_1;
	wire w_dff_B_W0VuoQNR9_0;
	wire w_dff_B_SJ2s7CJX8_0;
	wire w_dff_B_H8iMtuMh1_0;
	wire w_dff_B_0PYhF4O05_0;
	wire w_dff_B_iEFiicFC9_0;
	wire w_dff_B_0qwySIf04_0;
	wire w_dff_B_nODTLu8j8_0;
	wire w_dff_B_hwZ2QBFM2_0;
	wire w_dff_B_cq9WxawO3_0;
	wire w_dff_B_guJLuw7V8_0;
	wire w_dff_B_ap0gar116_0;
	wire w_dff_B_ze3dQJQJ8_0;
	wire w_dff_B_N72LmPrQ6_0;
	wire w_dff_B_MivFnubg2_0;
	wire w_dff_B_eEimXZ8n5_0;
	wire w_dff_B_8hT4PvgW8_0;
	wire w_dff_B_vLSC3Jhc8_0;
	wire w_dff_B_0HFVwDKA1_0;
	wire w_dff_B_fNWvu0Ba5_1;
	wire w_dff_B_Y8Kz8GFj8_1;
	wire w_dff_B_SycmWz7h0_1;
	wire w_dff_B_77Z1O1pc6_1;
	wire w_dff_B_SLkzalUW6_1;
	wire w_dff_B_WmxQRnwC7_1;
	wire w_dff_B_Mq51PVmM5_1;
	wire w_dff_B_SHf0hWt57_1;
	wire w_dff_B_4eLVmgno8_1;
	wire w_dff_B_ZJJK44hD6_1;
	wire w_dff_B_OZcxFgxD3_1;
	wire w_dff_B_S8tdATFH8_1;
	wire w_dff_B_RE3od9HI0_1;
	wire w_dff_B_ipm9Ljwo2_1;
	wire w_dff_B_pq6E21WS5_1;
	wire w_dff_B_SZKGjNZO4_1;
	wire w_dff_B_f9O6MNGd0_1;
	wire w_dff_B_Y58RtSJ29_1;
	wire w_dff_B_wotfyTJE5_1;
	wire w_dff_B_lU0gpBps2_1;
	wire w_dff_A_iHELKUG08_0;
	wire w_dff_A_JLMDq7te7_0;
	wire w_dff_A_XlXlueqR2_0;
	wire w_dff_A_C65bxzey1_0;
	wire w_dff_A_jwdxQDeC6_0;
	wire w_dff_A_RS3E63ZZ8_0;
	wire w_dff_A_zaEMJS5y1_2;
	wire w_dff_A_f1Ac9L4z1_2;
	wire w_dff_A_4Q7Rqo8r2_2;
	wire w_dff_A_5S8BuSF53_2;
	wire w_dff_A_n2SQzVNL3_2;
	wire w_dff_A_KeYBZipT4_2;
	wire w_dff_A_RMdziKXA7_2;
	wire w_dff_A_xs8At4Ad5_2;
	wire w_dff_A_ssuHvV1x9_2;
	wire w_dff_A_YEuyJf9P2_2;
	wire w_dff_A_eZyDpLQi3_2;
	wire w_dff_A_3d2wZlUO0_2;
	wire w_dff_A_XBNuIOju5_2;
	wire w_dff_A_wXEszY9E9_2;
	wire w_dff_A_Y4SC1a0I0_2;
	wire w_dff_A_QLIc4odz2_2;
	wire w_dff_A_IkYQX1ya8_2;
	wire w_dff_A_WcX8CP5O4_2;
	wire w_dff_A_eXFg4IlW1_1;
	wire w_dff_A_ScsDh4u38_1;
	wire w_dff_A_xhc8N4CO3_1;
	wire w_dff_A_V8lgoi8O3_1;
	wire w_dff_A_rqzMa1as8_1;
	wire w_dff_A_vKmt0qfj2_1;
	wire w_dff_A_SBDi12mP8_1;
	wire w_dff_A_0n4bZYXa1_1;
	wire w_dff_A_wQW1a9xD2_1;
	wire w_dff_A_gu81xreD1_1;
	wire w_dff_A_OxxtIKWa9_1;
	wire w_dff_A_3Vgv66q52_1;
	wire w_dff_A_qB07bLz41_1;
	wire w_dff_A_JNnxzt9i4_1;
	wire w_dff_A_SnYGJwgI1_1;
	wire w_dff_A_q74Muz0Z9_1;
	wire w_dff_A_FmQcAuyX1_2;
	wire w_dff_A_bVDZBFzy6_2;
	wire w_dff_A_BJg2IT4b6_2;
	wire w_dff_A_PMsPWmz07_2;
	wire w_dff_A_JVDka3Zi9_2;
	wire w_dff_A_pmBhRDCS4_2;
	wire w_dff_A_srwLQ5c40_2;
	wire w_dff_B_ADl4x1I67_1;
	wire w_dff_B_YIkN63ix3_1;
	wire w_dff_B_02i94erj1_1;
	wire w_dff_B_1RqGvp9P5_1;
	wire w_dff_B_0ZkJsJOg0_1;
	wire w_dff_B_xbZwIeDv3_1;
	wire w_dff_B_CCf1sQqX0_1;
	wire w_dff_B_7i3JhJil5_1;
	wire w_dff_B_WdTnOeSQ7_1;
	wire w_dff_B_ZILFCqnK7_1;
	wire w_dff_B_s0jOnRZr4_1;
	wire w_dff_B_T0AZJEkz9_1;
	wire w_dff_B_H9PfolCh3_1;
	wire w_dff_B_IFzlGp5n3_1;
	wire w_dff_B_4dMFw2le9_1;
	wire w_dff_B_N973HRmS5_1;
	wire w_dff_B_gag6sJdH4_1;
	wire w_dff_B_ZhBvSANF8_1;
	wire w_dff_B_2TT89mhw0_1;
	wire w_dff_A_KaS8Gjmp7_0;
	wire w_dff_A_YDSjYdWi1_0;
	wire w_dff_A_6sNleYyk2_0;
	wire w_dff_A_QeuITl8g9_0;
	wire w_dff_A_uopNGU9Q9_0;
	wire w_dff_A_A64mu9WC9_0;
	wire w_dff_A_Nky4KSlY5_0;
	wire w_dff_A_YXbuRvEe6_2;
	wire w_dff_A_E8b3whZb0_2;
	wire w_dff_A_Z6sV74iU8_2;
	wire w_dff_A_ygwnds2u5_2;
	wire w_dff_A_BkgepQIr4_2;
	wire w_dff_A_EDUFbXmI6_2;
	wire w_dff_A_Fqya9Ppc7_2;
	wire w_dff_A_bvgAqDQA7_2;
	wire w_dff_A_yYPMmlIl2_2;
	wire w_dff_A_Yp2IxehB0_2;
	wire w_dff_A_Gi0yjUwF7_2;
	wire w_dff_A_7LVqeWkA3_2;
	wire w_dff_A_OsZUJQAV4_2;
	wire w_dff_A_Vf9Gdczv3_2;
	wire w_dff_A_LHry1Kob6_2;
	wire w_dff_A_yj4xZaDO9_2;
	wire w_dff_A_qDdl9PUa3_2;
	wire w_dff_A_Gx3srTJB5_2;
	wire w_dff_A_9vZJQ24L1_2;
	wire w_dff_A_SzmOzkWV1_1;
	wire w_dff_A_EawolTbo1_1;
	wire w_dff_A_c5kw5qj53_1;
	wire w_dff_A_CySUXMTS8_1;
	wire w_dff_A_0FhMjHqI6_1;
	wire w_dff_A_VUbQvf5T2_1;
	wire w_dff_A_KRZJpQur7_1;
	wire w_dff_A_VewggG2H4_1;
	wire w_dff_A_6QfcUjhk5_1;
	wire w_dff_A_qno6efzJ4_1;
	wire w_dff_A_foLlheHq1_1;
	wire w_dff_A_QOzIT3WG2_1;
	wire w_dff_A_DSCTJOUl1_1;
	wire w_dff_A_uKVMB4oG5_1;
	wire w_dff_A_4G2HRrGl2_1;
	wire w_dff_A_EoNtu0H00_1;
	wire w_dff_A_RFQeJ0rj8_1;
	wire w_dff_A_MN9hvVqO9_2;
	wire w_dff_A_zY7AvL4P7_2;
	wire w_dff_A_5tARJulS1_2;
	wire w_dff_A_iqPyKJ4v2_2;
	wire w_dff_A_HPm1gUJ59_2;
	wire w_dff_A_DF7xBQUR0_2;
	wire w_dff_A_KtPzDrIM2_2;
	wire w_dff_A_dwSHW1VY7_2;
	wire w_dff_A_TZqrMTYV7_2;
	wire w_dff_A_nShUj1GO1_2;
	wire w_dff_A_XlHVV9RA6_2;
	wire w_dff_A_kWN7fJzX1_1;
	wire w_dff_A_shACUS9a7_2;
	wire w_dff_B_kO1xlF5h5_1;
	wire w_dff_B_LfIV5xTx3_0;
	wire w_dff_B_UiMih9lw6_0;
	wire w_dff_B_bmXPNjKx8_0;
	wire w_dff_B_0XCAjgoC6_0;
	wire w_dff_B_7mLXmI0j0_0;
	wire w_dff_B_zibivfLm9_0;
	wire w_dff_B_rDNdzLCw9_0;
	wire w_dff_B_aCpFc6yW1_0;
	wire w_dff_B_xG6T76pF6_0;
	wire w_dff_B_6ARhtCrO9_0;
	wire w_dff_B_nLYEia8J2_0;
	wire w_dff_B_sMYYjckc0_0;
	wire w_dff_B_lpK4u32E2_0;
	wire w_dff_B_Q6TBJCfg7_0;
	wire w_dff_B_DenSSNA57_0;
	wire w_dff_B_i1VLYggP1_0;
	wire w_dff_B_7zETgrhx6_0;
	wire w_dff_B_sUjayH6W6_0;
	wire w_dff_B_pjxcf6tk2_1;
	wire w_dff_B_fnBqcRVL1_2;
	wire w_dff_B_9ka1Ae2n2_2;
	wire w_dff_B_uXGqDPoi2_2;
	wire w_dff_B_5nRWFFqr8_1;
	wire w_dff_B_BSIomkER9_1;
	wire w_dff_B_mRgcY9Nb7_1;
	wire w_dff_B_nCoNP1I53_1;
	wire w_dff_B_jSEeUeMY0_1;
	wire w_dff_B_DNB5IOhH3_1;
	wire w_dff_B_jcYqNVaM4_1;
	wire w_dff_B_bsWaEmUV7_1;
	wire w_dff_B_nvfFrwUp2_1;
	wire w_dff_B_oQwCSowM1_1;
	wire w_dff_B_H4yjJnyj3_1;
	wire w_dff_B_q7zrlhNy5_1;
	wire w_dff_B_IYsRfYYL9_1;
	wire w_dff_B_GTWJnPbN0_1;
	wire w_dff_B_3YKgXkRR4_1;
	wire w_dff_B_whtlgsNr0_1;
	wire w_dff_B_iOwKKTv57_1;
	wire w_dff_B_Gt6abUR49_1;
	wire w_dff_B_QQQYwGwz9_1;
	wire w_dff_B_nSyVskDI9_0;
	wire w_dff_B_8wF03YzM8_0;
	wire w_dff_B_aPuqufsa5_0;
	wire w_dff_B_8VUeNZon6_0;
	wire w_dff_B_yHoVVJiQ8_0;
	wire w_dff_B_WfVGL2fU4_0;
	wire w_dff_B_GY4ZbLlM0_0;
	wire w_dff_B_ITN3cMfV3_0;
	wire w_dff_B_HrHYRHr98_0;
	wire w_dff_B_cBe28yCV4_0;
	wire w_dff_B_XUgYyT8M9_0;
	wire w_dff_B_R9gTmzsv8_0;
	wire w_dff_B_AWCXUrGL8_0;
	wire w_dff_B_zvaA5D1N9_0;
	wire w_dff_B_g8Zkx60P2_0;
	wire w_dff_B_5MZ4CJjg4_0;
	wire w_dff_B_6rYAchRu8_0;
	wire w_dff_B_U9I6NSKP4_0;
	wire w_dff_B_VkqJ4JdF2_0;
	wire w_dff_A_2qNBQAAz1_1;
	wire w_dff_A_KXq6F43g4_1;
	wire w_dff_A_M7eigc2J0_1;
	wire w_dff_A_mE0bREcL4_1;
	wire w_dff_A_e3XV9LNK4_1;
	wire w_dff_A_vxnwc74m0_1;
	wire w_dff_A_WlQMOzsc4_1;
	wire w_dff_A_q6RkgbSP8_1;
	wire w_dff_A_XhfRU2u52_1;
	wire w_dff_A_0V4Iu1L22_1;
	wire w_dff_A_Y90mAvUv5_1;
	wire w_dff_A_1iWUyKb64_1;
	wire w_dff_A_stdcJoPf5_1;
	wire w_dff_A_4erDwzrp7_1;
	wire w_dff_A_H93Uu6Zn8_1;
	wire w_dff_A_pR8iYj328_1;
	wire w_dff_A_EAQwzC245_1;
	wire w_dff_A_cKvkMZMF8_1;
	wire w_dff_A_a0wee1C72_1;
	wire w_dff_A_lOfGrWq38_1;
	wire w_dff_B_EiferPjr7_1;
	wire w_dff_B_LEYSzV9g6_1;
	wire w_dff_B_WDjFJlta3_1;
	wire w_dff_B_A5UV8FbO1_1;
	wire w_dff_B_vPNP0QHB0_1;
	wire w_dff_B_srRKSC302_1;
	wire w_dff_A_uP4cssC57_1;
	wire w_dff_B_zLvkXYvw7_1;
	wire w_dff_B_Ctzvl1pv9_1;
	wire w_dff_B_ccoYs86D7_1;
	wire w_dff_B_fAtLgESn2_1;
	wire w_dff_B_h2h6XhD24_1;
	wire w_dff_B_78h5uKli9_1;
	wire w_dff_B_y4lPWIZM9_1;
	wire w_dff_B_Ycw62p2G9_1;
	wire w_dff_B_OKGcimLH4_1;
	wire w_dff_B_T5OrYCv76_1;
	wire w_dff_B_B8p0AihC4_0;
	wire w_dff_B_rYpnkdck4_0;
	wire w_dff_A_DAnZjvDa5_1;
	wire w_dff_A_RU3PesLf9_1;
	wire w_dff_A_i4tnNOao0_1;
	wire w_dff_B_JlEetKWX5_0;
	wire w_dff_B_93VvCCoL9_1;
	wire w_dff_B_fBAZfIPF1_1;
	wire w_dff_B_CmMYRjGy6_1;
	wire w_dff_B_k8wkP7V45_1;
	wire w_dff_B_l5805JJW3_1;
	wire w_dff_B_qtoGbi9Q3_1;
	wire w_dff_B_DvW9Xmlr0_1;
	wire w_dff_B_mn2IDOe53_1;
	wire w_dff_B_ImFpiWwF0_1;
	wire w_dff_B_6ADLqYUy0_1;
	wire w_dff_B_8lN77ZZV8_1;
	wire w_dff_B_E8bw2Xc02_1;
	wire w_dff_B_5hVWzVVv8_1;
	wire w_dff_B_xPpdEmg91_1;
	wire w_dff_B_hahaZNaU7_1;
	wire w_dff_B_m1reyT1g6_1;
	wire w_dff_B_DZsrSaJC9_1;
	wire w_dff_B_5XddWEBp3_0;
	wire w_dff_A_HcOHyT6M2_0;
	wire w_dff_A_X51ckPEc8_0;
	wire w_dff_A_dwyuefgZ4_0;
	wire w_dff_B_41D4gjXK6_1;
	wire w_dff_A_q39Y62Qo9_1;
	wire w_dff_A_7U8dAIfM4_0;
	wire w_dff_A_Dj08AoB85_0;
	wire w_dff_A_3BqQ1vZL7_0;
	wire w_dff_A_GRkkIbkc5_0;
	wire w_dff_A_yFlhvwaL7_0;
	wire w_dff_A_vMZcvEne7_2;
	wire w_dff_A_v8ccX43L2_2;
	wire w_dff_A_6R0eBoST5_2;
	wire w_dff_A_43kEHPEg7_2;
	wire w_dff_A_7VdfCcrB8_2;
	wire w_dff_A_SfMgCxe87_2;
	wire w_dff_A_J6xtzue03_1;
	wire w_dff_A_exhrGTRb2_1;
	wire w_dff_A_U8cEK5rx7_1;
	wire w_dff_A_bsDESXrn1_1;
	wire w_dff_A_Llzfcz2D6_1;
	wire w_dff_A_9p8FwHgm0_1;
	wire w_dff_A_oFlFmqrn6_2;
	wire w_dff_A_VZ74eUt02_2;
	wire w_dff_B_3haLFshg7_2;
	wire w_dff_B_YNCr1ghA7_2;
	wire w_dff_B_H8r2rb7a7_2;
	wire w_dff_B_qSk3uBpR2_2;
	wire w_dff_B_kx3bsKHd9_2;
	wire w_dff_B_5c34sflw2_2;
	wire w_dff_B_YU7MduXM0_2;
	wire w_dff_B_PlWYkjCq5_2;
	wire w_dff_B_G0r8g5BP1_2;
	wire w_dff_A_p02ZZeyY1_1;
	wire w_dff_A_PiutBOKW9_1;
	wire w_dff_A_fo7ty2Ig3_1;
	wire w_dff_A_vi7fcVaA1_1;
	wire w_dff_A_qyJST7g97_1;
	wire w_dff_A_T9XOHi6A6_1;
	wire w_dff_A_FmJG8Dnv8_1;
	wire w_dff_A_19NKEVfM8_1;
	wire w_dff_A_zsOTnmHl7_1;
	wire w_dff_A_8mvt0AeL9_1;
	wire w_dff_A_ZHVBNmEb4_1;
	wire w_dff_A_oxz4LApm0_1;
	wire w_dff_A_2vLDGwbn1_1;
	wire w_dff_A_YybsqF5R9_1;
	wire w_dff_A_lDwR0oxZ1_2;
	wire w_dff_A_83I4TDbd0_0;
	wire w_dff_A_VhoHiYwh2_0;
	wire w_dff_A_XEg2A39h3_0;
	wire w_dff_A_1MjHR3At8_0;
	wire w_dff_A_FKyPYXmF7_0;
	wire w_dff_A_CRdPderv7_0;
	wire w_dff_A_nQxZ6Apw4_0;
	wire w_dff_A_bInQ2ewd0_0;
	wire w_dff_A_8aOzhEPB5_0;
	wire w_dff_A_9i10deTR1_0;
	wire w_dff_A_yQLIJlPF6_0;
	wire w_dff_A_07bBmpDT9_0;
	wire w_dff_B_jKVjrq5X9_1;
	wire w_dff_B_fhLSiVLT7_0;
	wire w_dff_B_E6HVoo1T4_0;
	wire w_dff_B_TQRLK7av2_0;
	wire w_dff_B_0jfqp2Sr6_0;
	wire w_dff_A_A7pyJF0q2_1;
	wire w_dff_A_GIQAnLri7_1;
	wire w_dff_A_c2uT18W97_1;
	wire w_dff_A_h1JDWaJA3_1;
	wire w_dff_A_qkS26nqD6_1;
	wire w_dff_B_M8L1t6OB9_2;
	wire w_dff_B_sCZfvn0t7_2;
	wire w_dff_B_Ki3Mc9955_2;
	wire w_dff_B_p2gEwM9Z5_2;
	wire w_dff_B_qYv6NP3V6_2;
	wire w_dff_B_246mbD024_0;
	wire w_dff_B_IKKyRrnr9_0;
	wire w_dff_B_S1s3UIPE3_1;
	wire w_dff_B_dh32HErn3_1;
	wire w_dff_B_Q5aEoJqx2_1;
	wire w_dff_A_qLi9mKAP9_1;
	wire w_dff_A_i29xRiPG6_1;
	wire w_dff_A_MmFNpZCS8_1;
	wire w_dff_A_HmG6Z6ho0_2;
	wire w_dff_A_2gdmoAsn9_2;
	wire w_dff_A_6tH0pIWo0_2;
	wire w_dff_A_RMtnfA0Q2_2;
	wire w_dff_A_Cx4XFVwu0_2;
	wire w_dff_A_ppNgcQAy5_2;
	wire w_dff_A_uonOlQ6T0_2;
	wire w_dff_B_5M9btRQs8_3;
	wire w_dff_A_l8vT5vQK1_0;
	wire w_dff_A_VNLyh4yD4_0;
	wire w_dff_A_t9r41Nco3_0;
	wire w_dff_A_vw1ZzAog0_0;
	wire w_dff_A_kLsYy4kh4_0;
	wire w_dff_A_rhwnmWmK9_0;
	wire w_dff_A_ohl3pi0p0_0;
	wire w_dff_A_nXyAlhw77_0;
	wire w_dff_A_KnkyxPvf7_0;
	wire w_dff_B_1KEajjX92_1;
	wire w_dff_A_kUQDiRdJ1_1;
	wire w_dff_A_JlBhJpDg0_0;
	wire w_dff_A_d4qRLEDP4_0;
	wire w_dff_A_a3SyjLHw4_0;
	wire w_dff_A_sutFpcGy7_0;
	wire w_dff_A_uCbpn1v40_0;
	wire w_dff_A_D8G3IhyY8_0;
	wire w_dff_A_ye3YonQl8_0;
	wire w_dff_A_wNlLgMxG5_0;
	wire w_dff_A_yKP8tZG88_0;
	wire w_dff_A_OuggQ7wO4_2;
	wire w_dff_A_xoIC4ohq8_2;
	wire w_dff_A_cPVSayx24_2;
	wire w_dff_A_LSHlXkhS6_2;
	wire w_dff_A_FIgmJxWn2_2;
	wire w_dff_A_MlFFv0D18_2;
	wire w_dff_B_5BaMNZE13_0;
	wire w_dff_B_d9S4yyXW1_1;
	wire w_dff_A_Ah5jx5xq6_0;
	wire w_dff_A_5FaKLTAu6_0;
	wire w_dff_A_hdHaghVi9_0;
	wire w_dff_A_7y3fmF6K9_0;
	wire w_dff_A_KMCz86P61_0;
	wire w_dff_A_ZHwX3Y8X3_0;
	wire w_dff_A_T63qrX6K1_0;
	wire w_dff_A_EgHcgpFC8_0;
	wire w_dff_A_mB80jkcS5_0;
	wire w_dff_A_zpxvzAgL6_0;
	wire w_dff_A_OwxKxIKB0_0;
	wire w_dff_A_RZPL5dbr7_0;
	wire w_dff_A_mdWYaNkU6_0;
	wire w_dff_B_kjeHPyV10_0;
	wire w_dff_B_Ku26dCwl2_1;
	wire w_dff_A_7qnZTphL5_1;
	wire w_dff_A_BkVAH2ZV8_2;
	wire w_dff_A_vwcKKIkE5_2;
	wire w_dff_A_VRwsdY0y4_2;
	wire w_dff_A_A3OPp8uX3_2;
	wire w_dff_A_azJ1Cwza1_2;
	wire w_dff_A_6qlwNx9c4_2;
	wire w_dff_A_BeDjNIWs3_2;
	wire w_dff_A_sp6qozvR2_2;
	wire w_dff_A_tAJIxZZM3_2;
	wire w_dff_A_zHqaBtl11_2;
	wire w_dff_A_m2MJmds47_2;
	wire w_dff_B_y2tM4x287_1;
	wire w_dff_B_9MSpMEdm3_1;
	wire w_dff_B_l1rPpzD15_0;
	wire w_dff_B_QJtKWBiP2_0;
	wire w_dff_B_bavSCnqv8_0;
	wire w_dff_A_607vqbmS9_0;
	wire w_dff_A_0bob9csf8_0;
	wire w_dff_A_HIdUAKGh5_0;
	wire w_dff_A_nmDxEz0M2_1;
	wire w_dff_A_YPqa7FE77_1;
	wire w_dff_A_ArazxxYs6_1;
	wire w_dff_A_y078HFsd3_1;
	wire w_dff_B_VrYukKn71_0;
	wire w_dff_A_PGqWpFTY3_0;
	wire w_dff_A_ye7KwXvM9_2;
	wire w_dff_A_rPjvbile5_0;
	wire w_dff_B_rkiHOKfh7_0;
	wire w_dff_A_7yrUm62o8_0;
	wire w_dff_A_zm4lqhY66_0;
	wire w_dff_A_5Xz5M9m92_0;
	wire w_dff_A_ekf3WwRm4_0;
	wire w_dff_A_pqviEFAC5_0;
	wire w_dff_A_rjfCWH7v3_0;
	wire w_dff_A_JZRfTq6S6_0;
	wire w_dff_A_IBfCtatM8_0;
	wire w_dff_A_tO8jjP8l6_0;
	wire w_dff_A_5bV9BeUp6_0;
	wire w_dff_A_2PvgxPFn8_0;
	wire w_dff_A_J7IMqfUf0_2;
	wire w_dff_A_eqOLkfew4_2;
	wire w_dff_A_bYIpvWPS6_2;
	wire w_dff_A_G1x36azM6_2;
	wire w_dff_A_CNIbL2NR6_2;
	wire w_dff_A_wKjQFHTu1_2;
	wire w_dff_A_ESHT4cdV3_2;
	wire w_dff_A_yp2Uiusj4_2;
	wire w_dff_B_JGqAcsRr8_1;
	wire w_dff_B_GHUFqe1f3_1;
	wire w_dff_B_fulIQZQl7_1;
	wire w_dff_B_9sooi4Uc8_1;
	wire w_dff_B_8kjyRUHx5_1;
	wire w_dff_B_UwWcPl1b7_1;
	wire w_dff_B_SLHDcqRL3_1;
	wire w_dff_B_t1eZh6es9_1;
	wire w_dff_B_b1MTaIZk2_1;
	wire w_dff_B_LeAwGtZq7_1;
	wire w_dff_B_boRSAyMn0_1;
	wire w_dff_B_WFuUAlZN4_1;
	wire w_dff_B_znUCkEJB4_1;
	wire w_dff_B_W4dZU0oB8_1;
	wire w_dff_B_J8ZZvl7V7_1;
	wire w_dff_A_jDdGjmD57_0;
	wire w_dff_A_IFsxbyU17_0;
	wire w_dff_A_9v7IrxGW5_1;
	wire w_dff_A_xwNgPe5F2_1;
	wire w_dff_A_QfJbN9cG1_1;
	wire w_dff_A_fZ1P4Zf60_1;
	wire w_dff_A_c6KmzTiU9_1;
	wire w_dff_A_BlrkuVzQ3_1;
	wire w_dff_A_JD0BOWzY6_0;
	wire w_dff_A_tNKKSYbO1_0;
	wire w_dff_A_UvZHh7uC5_1;
	wire w_dff_A_6QtFNhGn3_1;
	wire w_dff_A_bRFzw5NC2_1;
	wire w_dff_A_HKufdfLD0_1;
	wire w_dff_A_tGhsZud05_2;
	wire w_dff_A_CKr4KLtG9_2;
	wire w_dff_A_IcUKXp9b7_0;
	wire w_dff_A_IDL7tBGd6_0;
	wire w_dff_A_n0fgwF552_0;
	wire w_dff_A_S9nwTBvd1_1;
	wire w_dff_A_289YKKsd7_0;
	wire w_dff_A_5nV0ELg97_2;
	wire w_dff_A_gHKJPNrq2_0;
	wire w_dff_A_tX71DhYN1_0;
	wire w_dff_A_vjaJejNG5_0;
	wire w_dff_A_JWom5X3a3_0;
	wire w_dff_A_2HCW811z8_1;
	wire w_dff_A_MGTmNajW1_1;
	wire w_dff_A_O8HdHmMk5_2;
	wire w_dff_A_e2wFTsdm5_2;
	wire w_dff_A_sDamZIWu9_2;
	wire w_dff_A_HBGiEuX35_2;
	wire w_dff_B_rYGqbmNG0_1;
	wire w_dff_A_LT5SgMpK3_0;
	wire w_dff_A_TWNRPvyV2_2;
	wire w_dff_A_7Eb9Jmja7_1;
	wire w_dff_A_dWzcPerA0_0;
	wire w_dff_A_CaI8okV65_0;
	wire w_dff_A_3PmkaxBr7_0;
	wire w_dff_A_Sg7RcbN19_0;
	wire w_dff_A_rjwvY9S35_0;
	wire w_dff_A_ydPM95mj5_0;
	wire w_dff_A_2zAA9Umb0_0;
	wire w_dff_B_SQxsLgcW7_1;
	wire w_dff_B_fwDQ9fKU8_1;
	wire w_dff_A_u6mEIkBT1_1;
	wire w_dff_A_YprWSQXl2_1;
	wire w_dff_A_UQf0Whvu4_1;
	wire w_dff_A_8JQLu9eK9_1;
	wire w_dff_A_MkKKhlk65_1;
	wire w_dff_A_u5EHQxMO5_1;
	wire w_dff_A_LNrO9Vr24_1;
	wire w_dff_A_dRdZwZm91_1;
	wire w_dff_A_sUXL1Gpm1_1;
	wire w_dff_A_PSud7I7X4_1;
	wire w_dff_A_2nGnnnYf9_1;
	wire w_dff_A_nArJsp985_1;
	wire w_dff_A_h6TM1nLb0_1;
	wire w_dff_A_jl11dvRb3_1;
	wire w_dff_A_BuIuQJ7E7_1;
	wire w_dff_A_mlFn4RIz5_1;
	wire w_dff_A_mJUPKJal7_1;
	wire w_dff_A_kLbvHeRq5_1;
	wire w_dff_A_WWz6kItk5_2;
	wire w_dff_A_yoTy8XiB6_2;
	wire w_dff_A_FO2LjoWX8_2;
	wire w_dff_A_jRCz178b5_2;
	wire w_dff_A_H3iU3qlg3_2;
	wire w_dff_A_iDrou3bl9_2;
	wire w_dff_A_DVM9SFrA2_2;
	wire w_dff_A_bD7SVp1N3_2;
	wire w_dff_A_fxY25Nyx7_2;
	wire w_dff_A_m8eHBqdZ6_2;
	wire w_dff_A_vJ2Onia90_0;
	wire w_dff_A_fOBNq5Es2_0;
	wire w_dff_B_khmYPcgz9_1;
	wire w_dff_B_Cn27TpIJ0_1;
	wire w_dff_B_rhIZik0W9_1;
	wire w_dff_B_kRJT3wse7_1;
	wire w_dff_A_7Lv7AdWl5_1;
	wire w_dff_A_ddU9OMzw0_0;
	wire w_dff_A_VW1wU9Xh5_0;
	wire w_dff_A_wK71iNMU8_0;
	wire w_dff_A_t8pGFjp86_0;
	wire w_dff_A_MIQ1Y4FX5_1;
	wire w_dff_A_THHCLd8W5_1;
	wire w_dff_A_uvjxOwaX1_1;
	wire w_dff_A_C7If0JOz7_2;
	wire w_dff_A_y0LvTvBl1_2;
	wire w_dff_A_TIFXSPOy5_2;
	wire w_dff_A_Pru7XwWy6_2;
	wire w_dff_A_2TCoX7101_1;
	wire w_dff_A_o35FUYa91_1;
	wire w_dff_B_j3XPcoFH2_1;
	wire w_dff_B_5XAEIhWx1_1;
	wire w_dff_A_x1spk4jM5_2;
	wire w_dff_B_Q4dSipxa8_3;
	wire w_dff_A_5nmcFANn6_0;
	wire w_dff_A_gEgy98RR2_0;
	wire w_dff_A_hFq9wJpJ8_0;
	wire w_dff_A_5qhikpfe9_1;
	wire w_dff_B_aWUAzN4U2_1;
	wire w_dff_A_kJ1VNvQG9_1;
	wire w_dff_A_cvrUomGe6_1;
	wire w_dff_A_1OY5sP727_1;
	wire w_dff_A_VidaYrBB3_2;
	wire w_dff_A_xiyzJKe73_2;
	wire w_dff_A_0pFK2Ner1_2;
	wire w_dff_A_OglsVBYO9_0;
	wire w_dff_A_Rtj5CWw78_2;
	wire w_dff_A_6st0OpoW4_1;
	wire w_dff_A_FlZ0ONBZ3_2;
	wire w_dff_A_rhNxgrBE4_2;
	wire w_dff_A_iMsQLFAt3_1;
	wire w_dff_B_TBo6RMLm5_1;
	wire w_dff_B_Ywm0ecfJ3_1;
	wire w_dff_B_lAeKIlEP8_1;
	wire w_dff_B_Nsmg6kdC0_1;
	wire w_dff_B_HrGeroVV9_1;
	wire w_dff_A_T7u7M1HZ3_0;
	wire w_dff_A_TiknX4FY5_0;
	wire w_dff_A_4rgexoVy5_0;
	wire w_dff_A_FWhTANMH7_1;
	wire w_dff_A_sGs16ISw7_1;
	wire w_dff_A_yhl7EdmH5_1;
	wire w_dff_A_gzcDVFSt0_1;
	wire w_dff_A_eREKj2st1_1;
	wire w_dff_A_LAxhXHmZ7_2;
	wire w_dff_A_fTEYH5MJ3_2;
	wire w_dff_A_4J7QjujL1_2;
	wire w_dff_A_msxUPXKl5_0;
	wire w_dff_B_DYaX8Hgu3_1;
	wire w_dff_B_Ad7FIs4t6_1;
	wire w_dff_A_HqRQQ5Dw3_0;
	wire w_dff_A_v2PmSzza2_0;
	wire w_dff_A_RvHiWXFc7_0;
	wire w_dff_A_V2gQG1eZ7_0;
	wire w_dff_A_MvzDF7Oj4_0;
	wire w_dff_A_C5PijlUF7_1;
	wire w_dff_A_GTBQ4FCe4_1;
	wire w_dff_A_1kxmuCHH2_1;
	wire w_dff_A_DtmHDySL8_2;
	wire w_dff_A_swKeyPw01_2;
	wire w_dff_A_5hM7wWQg4_2;
	wire w_dff_A_77KRC1lc4_0;
	wire w_dff_A_4NWISi2H3_0;
	wire w_dff_A_j41D3iUL7_1;
	wire w_dff_A_9RxrP5xD1_0;
	wire w_dff_A_USqn9juS4_2;
	wire w_dff_A_rU5hIRg20_1;
	wire w_dff_B_a2v8VoHg4_1;
	wire w_dff_B_nc06qPDF0_1;
	wire w_dff_A_X8JEPTvo8_0;
	wire w_dff_A_SLhPDG6J2_2;
	wire w_dff_A_rVsBUueX2_2;
	wire w_dff_A_QGecVUIb6_0;
	wire w_dff_A_92YtTzxb0_1;
	wire w_dff_A_6KjX17et2_1;
	wire w_dff_A_6PiK53K50_1;
	wire w_dff_A_RDUmUsws8_2;
	wire w_dff_A_zDMoByYg7_2;
	wire w_dff_A_bcnZ5QXg4_1;
	wire w_dff_A_8Kvxk1sW7_2;
	wire w_dff_A_aze7x1926_2;
	wire w_dff_A_pFPTIqm75_2;
	wire w_dff_A_uZpT0iYG7_2;
	wire w_dff_A_hvkmYb9T5_2;
	wire w_dff_A_W4QeQyRj1_2;
	wire w_dff_A_yBmEkHR52_2;
	wire w_dff_A_ph5qFrFO9_2;
	wire w_dff_A_q9xs8aBf7_2;
	wire w_dff_A_IW8s2snX7_2;
	wire w_dff_A_rxs8mDsb4_2;
	wire w_dff_A_xCoe0Yxo1_2;
	wire w_dff_A_NLKlnGtd4_0;
	wire w_dff_A_HYLUqFkp4_0;
	wire w_dff_A_GYLgjmw42_0;
	wire w_dff_A_nm9NQ2Pf3_0;
	wire w_dff_A_EfLg9am28_0;
	wire w_dff_A_LW7Mt9wV8_0;
	wire w_dff_A_7eioFKEk0_2;
	wire w_dff_A_ZuuYbSaV3_2;
	wire w_dff_A_h1nyXclN6_2;
	wire w_dff_A_fdlHF7ir3_2;
	wire w_dff_A_HZ5IFSO28_2;
	wire w_dff_A_KF45V0xS4_2;
	wire w_dff_A_bISymSaK6_2;
	wire w_dff_A_taQFjGuE7_2;
	wire w_dff_A_Voo3CxCM6_2;
	wire w_dff_A_ND6PrY139_2;
	wire w_dff_A_Z9p8ucLv1_2;
	wire w_dff_A_AIgbrBNr3_2;
	wire w_dff_A_xLgZBadQ1_2;
	wire w_dff_A_RW3szw4Z4_2;
	wire w_dff_A_IjIs24Tj0_2;
	wire w_dff_A_kW6BxD995_2;
	wire w_dff_A_Ytz3WvXx7_2;
	wire w_dff_A_IDxTqGVC1_2;
	wire w_dff_A_Deyg2NPH8_1;
	wire w_dff_A_RMquG1VH5_1;
	wire w_dff_A_qAkVl2KR2_1;
	wire w_dff_A_S8Q5VEb37_1;
	wire w_dff_A_iGo2aX4h1_1;
	wire w_dff_A_QldryrM18_1;
	wire w_dff_A_OmHXET6u8_1;
	wire w_dff_A_afAF2FrS8_1;
	wire w_dff_A_zWIkN5RY2_1;
	wire w_dff_A_2CqVssKs0_1;
	wire w_dff_A_JreCyYxF9_1;
	wire w_dff_A_wYxPPXOo4_1;
	wire w_dff_A_7aE8ig800_1;
	wire w_dff_A_TH0PPm387_1;
	wire w_dff_A_zOfvnnl55_1;
	wire w_dff_A_32D0wbyv8_1;
	wire w_dff_A_wsDP1bJN1_2;
	wire w_dff_A_QRo3H8Pp1_2;
	wire w_dff_A_jk0adFD75_2;
	wire w_dff_A_FaY6W2PO3_2;
	wire w_dff_A_xchrOceB9_2;
	wire w_dff_A_SA6K04Ui8_2;
	wire w_dff_A_wXW4sHwz1_2;
	wire w_dff_B_D0CWybsJ3_1;
	wire w_dff_B_E9pVTg2h6_1;
	wire w_dff_B_gYfskHur3_1;
	wire w_dff_B_iYhTyRRk3_1;
	wire w_dff_B_Wik5T94l9_1;
	wire w_dff_B_f7yEEDOe6_1;
	wire w_dff_B_YNReeq394_1;
	wire w_dff_B_266Bsybs0_1;
	wire w_dff_B_U7qNGUDw4_1;
	wire w_dff_B_w8H034wv6_1;
	wire w_dff_B_obFN7baq1_1;
	wire w_dff_B_KqzyrakD9_1;
	wire w_dff_B_qhIFKDUt1_1;
	wire w_dff_B_403AIYZk7_1;
	wire w_dff_B_on9cbfOZ0_1;
	wire w_dff_B_AvbfHbsE0_1;
	wire w_dff_B_3cmqoIzR5_1;
	wire w_dff_B_BhU5I1SB5_1;
	wire w_dff_B_y6t5PHBq2_1;
	wire w_dff_B_m9RvD3KT2_0;
	wire w_dff_B_bAjPbLHg5_0;
	wire w_dff_B_t283aIEp3_0;
	wire w_dff_B_07k7FyeT2_0;
	wire w_dff_B_K80B8jMO0_0;
	wire w_dff_B_rThIxeqp0_0;
	wire w_dff_B_kbljello1_0;
	wire w_dff_B_sqNmiUWR4_0;
	wire w_dff_B_oeJrBfkf2_0;
	wire w_dff_B_dj564phh1_0;
	wire w_dff_B_eg3XnDXj7_0;
	wire w_dff_B_ruonKnZQ4_0;
	wire w_dff_B_jZD2Stwo6_0;
	wire w_dff_B_sb0Pk6hN5_0;
	wire w_dff_B_55jthq2E1_0;
	wire w_dff_B_qSjIQnq75_0;
	wire w_dff_B_ZCNmBO4p3_0;
	wire w_dff_B_bcAW2MU46_0;
	wire w_dff_B_CczamCeA6_0;
	wire w_dff_B_y6eSBI4b3_1;
	wire w_dff_B_cybQlxok1_1;
	wire w_dff_B_71f4yUDK4_1;
	wire w_dff_B_cMGm7CZg8_1;
	wire w_dff_B_5OhrnJ7w7_1;
	wire w_dff_B_cEHmt6JV6_1;
	wire w_dff_B_SSdPyBsD3_1;
	wire w_dff_B_JxnJFHBJ9_1;
	wire w_dff_B_voDq9m3C7_0;
	wire w_dff_B_OBkh3hor7_0;
	wire w_dff_B_Y0KUzQp49_1;
	wire w_dff_B_fDgFNn5p1_0;
	wire w_dff_B_HmHRIsmj7_0;
	wire w_dff_B_13uFmaH52_0;
	wire w_dff_B_8LDZHcFf0_0;
	wire w_dff_B_oHymJl9Z4_1;
	wire w_dff_B_p0OjHqQ14_1;
	wire w_dff_B_Oo98Fwqg2_1;
	wire w_dff_B_hvQyuDWe6_1;
	wire w_dff_B_kfga65Hg1_1;
	wire w_dff_B_oKx2tdWk3_1;
	wire w_dff_B_s6FttiPF9_1;
	wire w_dff_B_BK8bDYqc8_1;
	wire w_dff_B_NRoWvbCT3_1;
	wire w_dff_B_zJkuUrqE1_1;
	wire w_dff_B_CPYGXWMg6_1;
	wire w_dff_B_gm7OfTpl8_1;
	wire w_dff_B_KRgvwtkw4_1;
	wire w_dff_B_TWtG4G4Q2_1;
	wire w_dff_B_m5YzHZ2X8_1;
	wire w_dff_B_WWxDy1XO9_1;
	wire w_dff_B_ZEHe0Y898_1;
	wire w_dff_B_NyEhML011_1;
	wire w_dff_B_8v8wTRNY5_1;
	wire w_dff_B_PtQ18N2B6_1;
	wire w_dff_B_XIfNXhkf4_1;
	wire w_dff_B_GIHZRyBw4_1;
	wire w_dff_B_LvevyD0u7_1;
	wire w_dff_A_hEsPBp8w3_0;
	wire w_dff_A_1lupsNG66_1;
	wire w_dff_B_MtLqDPHt3_2;
	wire w_dff_B_Br1j1YCb7_2;
	wire w_dff_B_jurjrizg7_2;
	wire w_dff_B_kllcc4En5_2;
	wire w_dff_A_QxLJaRx41_0;
	wire w_dff_A_9O4EolNm4_0;
	wire w_dff_A_srsVW9Af9_0;
	wire w_dff_A_j8tzyT2m1_0;
	wire w_dff_A_jHm2wTS61_1;
	wire w_dff_A_zKmaTsBv8_1;
	wire w_dff_B_fiDJVqRi0_1;
	wire w_dff_B_9mibG71Y7_0;
	wire w_dff_B_IJNya5Rl8_1;
	wire w_dff_A_ikduT0UA6_0;
	wire w_dff_A_i0edykUa5_0;
	wire w_dff_B_LOnslHMK5_2;
	wire w_dff_B_KrP6ACxw1_2;
	wire w_dff_B_tMwK3bNH7_2;
	wire w_dff_B_JjpdH9y39_2;
	wire w_dff_B_bsSRZaF56_2;
	wire w_dff_B_bK8R2NEB5_2;
	wire w_dff_B_3kGxsvzi2_0;
	wire w_dff_B_IknBggBW4_0;
	wire w_dff_B_wrBjtwS76_0;
	wire w_dff_B_CCqndtHG8_0;
	wire w_dff_B_7ohlDYPp9_0;
	wire w_dff_B_e0AiH9RI4_0;
	wire w_dff_B_SCPpuGLX7_0;
	wire w_dff_B_3TEKFXjF7_0;
	wire w_dff_A_BSIOabYs3_2;
	wire w_dff_A_y1EzK1zt2_2;
	wire w_dff_A_wJ97G8MC0_2;
	wire w_dff_A_aKdImrnP2_2;
	wire w_dff_A_SsmDP4dU2_2;
	wire w_dff_A_l3KMi0Lf5_2;
	wire w_dff_A_YPhObIO37_2;
	wire w_dff_A_jWiQ0e9t3_2;
	wire w_dff_A_YYDdGiXM6_2;
	wire w_dff_A_aTQiV29g7_2;
	wire w_dff_A_jLfgwm3B2_2;
	wire w_dff_A_vtSVt5Ke4_2;
	wire w_dff_A_oxQIZz4S9_1;
	wire w_dff_A_GKLhhMUB8_1;
	wire w_dff_A_rrWg23Ee9_1;
	wire w_dff_A_ogIfQWlc6_1;
	wire w_dff_A_1syFJ1BI3_1;
	wire w_dff_A_wopdOaqf6_1;
	wire w_dff_A_Zw8N9znH7_1;
	wire w_dff_A_vvnwE0dB6_1;
	wire w_dff_A_JiOFjd856_1;
	wire w_dff_A_YA3kvibd3_2;
	wire w_dff_A_lcrB65fP0_2;
	wire w_dff_A_Dnw3qxl19_2;
	wire w_dff_A_HhCA1haI8_2;
	wire w_dff_A_myzx6miw8_2;
	wire w_dff_A_SuTsqUUz7_2;
	wire w_dff_A_lTS9xalW3_2;
	wire w_dff_A_xzbAIfva8_2;
	wire w_dff_A_DcNViKZO3_2;
	wire w_dff_B_8w9SjXgu8_3;
	wire w_dff_B_cNCEHzcg0_3;
	wire w_dff_A_QPJrCzQ94_1;
	wire w_dff_A_uQWcp82E3_1;
	wire w_dff_A_HcWZaaDr7_1;
	wire w_dff_A_RabxUM5u6_0;
	wire w_dff_B_LWfr27by0_1;
	wire w_dff_B_zHdUCnVa4_1;
	wire w_dff_B_0rl6XDgm3_0;
	wire w_dff_B_PV5733b09_1;
	wire w_dff_B_yJUIuqCl3_2;
	wire w_dff_A_d2qPCzLc6_0;
	wire w_dff_B_IrYITDwn2_0;
	wire w_dff_B_I4f65N7O1_1;
	wire w_dff_A_BSGd3JMX3_1;
	wire w_dff_A_3ESHHXks4_1;
	wire w_dff_A_cwv6t5gy6_1;
	wire w_dff_A_m14ZmyXb3_1;
	wire w_dff_A_SkQ9pSQd8_1;
	wire w_dff_A_jEfh31XR7_1;
	wire w_dff_A_mLPZdrPX1_1;
	wire w_dff_A_ifObSwrm4_1;
	wire w_dff_A_pCOCpnTh6_1;
	wire w_dff_B_jqKCjf4A8_2;
	wire w_dff_B_JLAvMhPP4_2;
	wire w_dff_B_tHW24P2b1_2;
	wire w_dff_A_0flIumw26_0;
	wire w_dff_A_NFa9gf9t3_0;
	wire w_dff_A_PfRuB1eH7_0;
	wire w_dff_A_S5K49NIm7_0;
	wire w_dff_A_09eiEXdN9_0;
	wire w_dff_B_p3feOSO34_1;
	wire w_dff_B_WCFRpAvJ0_1;
	wire w_dff_B_6kfQng679_0;
	wire w_dff_A_ZUHGbJNA8_0;
	wire w_dff_B_CbaEUmP63_0;
	wire w_dff_B_SDAncjIu4_0;
	wire w_dff_A_7dpqGCjC5_0;
	wire w_dff_A_x5NtLHI71_0;
	wire w_dff_A_bnNVtO9w5_0;
	wire w_dff_A_63KvYAOB7_0;
	wire w_dff_A_BPpn6oSc2_0;
	wire w_dff_A_JRHCN90s7_0;
	wire w_dff_A_EXbfzPrL4_0;
	wire w_dff_A_P8xOK5uz1_1;
	wire w_dff_A_uK6OIkPM0_1;
	wire w_dff_A_wIlEuhuF7_1;
	wire w_dff_A_9WJodyuM8_1;
	wire w_dff_A_IwN1l2Xb1_0;
	wire w_dff_A_fMctWRTU0_0;
	wire w_dff_A_92dWOa9m5_0;
	wire w_dff_A_zTGz7cTw7_0;
	wire w_dff_A_mMMU0x3m6_0;
	wire w_dff_A_YLbN2nBA3_0;
	wire w_dff_B_Q17ELFLL2_2;
	wire w_dff_B_f1SPZpZX8_2;
	wire w_dff_A_LT7SfRtI1_0;
	wire w_dff_A_QeGAPcQN6_1;
	wire w_dff_A_TYKPX5VY6_1;
	wire w_dff_A_Q094VyXA8_1;
	wire w_dff_A_ZrUszQjG6_0;
	wire w_dff_A_5X3yEdkl6_0;
	wire w_dff_A_GrRXcfIM7_0;
	wire w_dff_A_Bb9lsqzh5_0;
	wire w_dff_A_kEMwIXIn5_0;
	wire w_dff_A_0Fa8os3z7_0;
	wire w_dff_A_FS4Kxid42_0;
	wire w_dff_A_oWUaqytK7_0;
	wire w_dff_A_dG2Mjsc11_0;
	wire w_dff_A_eSrgxN3W7_0;
	wire w_dff_A_OYUQNdxS0_0;
	wire w_dff_A_JqaM0uqn6_0;
	wire w_dff_A_JIsGZ0Ow2_2;
	wire w_dff_A_UsYkc8JY3_2;
	wire w_dff_A_bFLN5keE7_2;
	wire w_dff_A_2PVSg64j2_2;
	wire w_dff_A_kdVLLeTI5_2;
	wire w_dff_A_t9pvmhFv2_2;
	wire w_dff_A_PU2cSZfk8_2;
	wire w_dff_A_pMmppbiq0_2;
	wire w_dff_A_er9MN6VG4_2;
	wire w_dff_A_EWHZ9Osq4_2;
	wire w_dff_B_oq0Ywofd2_1;
	wire w_dff_B_gZDI64Ns3_1;
	wire w_dff_B_7T1LkwOg9_1;
	wire w_dff_B_ahsHh9Ol7_1;
	wire w_dff_B_CbbG04359_1;
	wire w_dff_B_bOYmoYFs5_1;
	wire w_dff_B_Xz7zCVNm5_1;
	wire w_dff_B_9hso8GXL7_1;
	wire w_dff_B_1PaqHFXG2_1;
	wire w_dff_A_8v12xvBk6_1;
	wire w_dff_A_JOLCGD738_0;
	wire w_dff_A_NiKCeGge1_0;
	wire w_dff_A_hVs7x4Xo4_1;
	wire w_dff_A_qTLdxIJi4_1;
	wire w_dff_A_ssmlvYDc9_1;
	wire w_dff_A_EvD6p0zS9_1;
	wire w_dff_A_VD5hiWkc2_2;
	wire w_dff_A_4yccVk0V6_2;
	wire w_dff_A_9prX5OOG0_2;
	wire w_dff_A_SU22FOku6_1;
	wire w_dff_A_dIXvuexv7_1;
	wire w_dff_A_iqc2tmVP1_0;
	wire w_dff_A_pe5x4dCf1_0;
	wire w_dff_A_CZu92rYw1_0;
	wire w_dff_A_Vpom8c187_1;
	wire w_dff_B_97Od1iLj9_2;
	wire w_dff_A_rdwYEB797_0;
	wire w_dff_A_BUnEjW585_1;
	wire w_dff_A_EeOODEu20_1;
	wire w_dff_A_LoROC9dG1_1;
	wire w_dff_A_6jdQc28D4_1;
	wire w_dff_A_cdBdRrEJ6_1;
	wire w_dff_B_c5b0SisU2_1;
	wire w_dff_B_OdDnxJVz1_1;
	wire w_dff_B_nYHrPa6X7_2;
	wire w_dff_B_NCF2avyc2_2;
	wire w_dff_B_70esU5vR8_2;
	wire w_dff_B_8sWR1LZ04_2;
	wire w_dff_B_MNvJXFBW1_2;
	wire w_dff_B_rABvzCqa6_2;
	wire w_dff_B_piFvOyF13_2;
	wire w_dff_B_FvrOhXZl9_2;
	wire w_dff_B_BIDd6ZH78_2;
	wire w_dff_B_4ofr7wj29_2;
	wire w_dff_A_fAbKqvX35_2;
	wire w_dff_A_OQaTlxtk6_2;
	wire w_dff_A_uMBcqh5w8_2;
	wire w_dff_A_96EIOfti0_2;
	wire w_dff_A_OVx7vuIf6_2;
	wire w_dff_A_3W9nTXQe8_1;
	wire w_dff_A_CZc7oxpZ0_1;
	wire w_dff_A_p16N9eAf4_1;
	wire w_dff_A_IRvJ5n7H9_1;
	wire w_dff_A_mRHePuIw5_1;
	wire w_dff_A_ZM6t2rqF7_1;
	wire w_dff_A_nLtBEqxt1_1;
	wire w_dff_B_y2DrAnYB0_0;
	wire w_dff_A_X5VE5Rn87_0;
	wire w_dff_B_ex8iQiFj3_1;
	wire w_dff_A_I48WH7cW8_0;
	wire w_dff_A_xwueaaXp8_0;
	wire w_dff_A_3XYAaoiY3_1;
	wire w_dff_A_BBMmeLKm0_1;
	wire w_dff_A_rEbBXL8M5_1;
	wire w_dff_A_gq866Uyx9_1;
	wire w_dff_A_iFiqIPSR9_1;
	wire w_dff_A_pTzrZNO72_1;
	wire w_dff_A_habZwT1r8_1;
	wire w_dff_A_hLTnTAOU5_1;
	wire w_dff_A_huzUM75a1_1;
	wire w_dff_A_wi0ZbLkl6_1;
	wire w_dff_A_n8KaUCZM2_1;
	wire w_dff_A_3kVqWks17_1;
	wire w_dff_A_rc6cyPT01_1;
	wire w_dff_A_nJ2td3iY0_1;
	wire w_dff_A_Gt3ZoqjV6_1;
	wire w_dff_A_K7sE6wq35_1;
	wire w_dff_B_7O06H6yB2_0;
	wire w_dff_B_oSc3NJlp1_1;
	wire w_dff_A_Y0C5iHwL0_0;
	wire w_dff_A_6CHDTV882_2;
	wire w_dff_A_SJM3llbf3_1;
	wire w_dff_A_u8JSnDQi1_1;
	wire w_dff_A_il7T7hol3_1;
	wire w_dff_A_IV7T04QO9_1;
	wire w_dff_A_NgP28wni9_1;
	wire w_dff_A_cuQLzaUW8_1;
	wire w_dff_A_bmyElyw24_1;
	wire w_dff_A_2ljb2NLh7_1;
	wire w_dff_A_1pPdm0Gj8_1;
	wire w_dff_A_830R7nnO7_1;
	wire w_dff_A_HWW4jZFn9_1;
	wire w_dff_A_nFQtPAcr9_1;
	wire w_dff_A_8s4z32cf7_1;
	wire w_dff_A_zfGaarHY9_1;
	wire w_dff_A_EdWZtHnH2_1;
	wire w_dff_A_zQQQTv6k9_1;
	wire w_dff_A_vGWoQ90w7_1;
	wire w_dff_A_HAUkrzKr3_2;
	wire w_dff_A_U6v1aeNf5_2;
	wire w_dff_A_G3jFXJA17_2;
	wire w_dff_A_n6Sv8eHr5_2;
	wire w_dff_A_uuHG5Q250_2;
	wire w_dff_A_Ru9HNxHt3_2;
	wire w_dff_A_uAOJH08I9_2;
	wire w_dff_A_NYquPSHS8_2;
	wire w_dff_A_5GaXf1406_2;
	wire w_dff_A_pMnAPbPy2_2;
	wire w_dff_A_fUn5nLBT4_2;
	wire w_dff_A_s5nuRzJv2_2;
	wire w_dff_A_VThthqik6_2;
	wire w_dff_A_zxu4Y6xJ2_2;
	wire w_dff_A_2vUuaBgp4_2;
	wire w_dff_A_wnUidp9P8_2;
	wire w_dff_A_GkHTtTX37_2;
	wire w_dff_A_9KWaRm4D7_2;
	wire w_dff_A_gV6NFZlV5_2;
	wire w_dff_A_vaajNmmr9_2;
	wire w_dff_A_xCnhGROG9_2;
	wire w_dff_A_ydaMKyjA1_2;
	wire w_dff_A_COWnrVOF2_2;
	wire w_dff_A_0n8QOOed6_2;
	wire w_dff_A_QMHeXJpH0_2;
	wire w_dff_A_2K3aXCom4_2;
	wire w_dff_A_mDT9zZ7v2_2;
	wire w_dff_B_otbjf07u4_2;
	wire w_dff_B_m1R52wP16_1;
	wire w_dff_B_AJTqV7fd2_1;
	wire w_dff_A_1YbHecmV2_0;
	wire w_dff_A_posRy3dw0_2;
	wire w_dff_A_8RSXgteW1_2;
	wire w_dff_A_d064H4t07_0;
	wire w_dff_A_Zw8gwf5R7_0;
	wire w_dff_A_6BR4DVNt6_1;
	wire w_dff_A_HlJL891t2_1;
	wire w_dff_A_rbLJ0fbJ2_2;
	wire w_dff_B_YIiBl1PT1_1;
	wire w_dff_B_pwRFMlrp9_1;
	wire w_dff_A_VieoZLRK7_2;
	wire w_dff_A_yQsZz6LY3_2;
	wire w_dff_B_c5M0faWB5_3;
	wire w_dff_B_s5CmWdDh1_1;
	wire w_dff_A_KFQivGam9_1;
	wire w_dff_A_PP7ffUZ67_0;
	wire w_dff_A_ntbxNQMz8_0;
	wire w_dff_A_G0yvkdsE8_1;
	wire w_dff_A_0vmrnqG67_0;
	wire w_dff_B_8WJiVgDg4_1;
	wire w_dff_B_dA7S9O0q4_1;
	wire w_dff_A_yzVfqSoE5_0;
	wire w_dff_A_XPcdGorN6_2;
	wire w_dff_A_C9wiUB3i5_2;
	wire w_dff_A_SQiowSOU1_0;
	wire w_dff_A_KwfjedKL4_1;
	wire w_dff_A_LR4UwY9l0_1;
	wire w_dff_A_ttdzmNqI7_2;
	wire w_dff_A_rSBlSYSC0_2;
	wire w_dff_A_bodr78eO0_2;
	wire w_dff_A_GHf1WuLw3_0;
	wire w_dff_A_e3JIbNxC8_2;
	wire w_dff_B_F7dSwWAA2_1;
	wire w_dff_B_t4xIJt4T5_1;
	wire w_dff_A_CQDvDQIN0_0;
	wire w_dff_A_KbGIdVt48_2;
	wire w_dff_A_53wdL9Ic4_2;
	wire w_dff_A_ZMRooXgA5_0;
	wire w_dff_A_jk4Zfurw9_0;
	wire w_dff_A_rrQKLtgY1_1;
	wire w_dff_A_zwQWhkLL1_0;
	wire w_dff_A_Z2ld8Ms42_2;
	wire w_dff_B_CggUUJyJ9_1;
	wire w_dff_B_McPhVsr13_1;
	wire w_dff_B_M2BfNANf4_1;
	wire w_dff_B_xqQZZMkN9_1;
	wire w_dff_A_2Fos1n793_1;
	wire w_dff_A_K1sSTTDM4_1;
	wire w_dff_A_PpQBE0k26_0;
	wire w_dff_A_ikHJwaSR6_0;
	wire w_dff_A_5utZaRT63_0;
	wire w_dff_A_kIlLJhno4_0;
	wire w_dff_A_uzNAGVgL4_2;
	wire w_dff_A_NIHaGDVF2_2;
	wire w_dff_A_Wvhep0ki2_1;
	wire w_dff_A_W0Bp2O9F7_2;
	wire w_dff_B_drKLrYsS4_1;
	wire w_dff_B_p5kmLarl3_1;
	wire w_dff_B_juMTaES87_2;
	wire w_dff_A_FCoTUeF00_0;
	wire w_dff_A_X5buWeyf0_0;
	wire w_dff_A_P62yhVsH3_0;
	wire w_dff_A_6D3Di4A10_1;
	wire w_dff_B_rzADqUVV1_1;
	wire w_dff_A_sblDCa1a4_1;
	wire w_dff_A_8XrAwFnq4_1;
	wire w_dff_A_IcWadWZz6_1;
	wire w_dff_A_u3XK0Zs11_2;
	wire w_dff_A_KoCm3FHP7_2;
	wire w_dff_A_KNLrAf8K1_2;
	wire w_dff_A_9a9Fd7d06_0;
	wire w_dff_B_vP9uQ1Iv3_1;
	wire w_dff_B_Z0Onc9aE6_1;
	wire w_dff_B_E0EfueVk5_2;
	wire w_dff_A_dTobYgT19_0;
	wire w_dff_B_PS8UhcAt3_1;
	wire w_dff_A_8jIdLr0h7_1;
	wire w_dff_A_Hs8KFHmw9_0;
	wire w_dff_A_bi0OmC4g3_0;
	wire w_dff_A_dQHbuo6n9_0;
	wire w_dff_A_1yF74THA3_2;
	wire w_dff_A_TPUCpvG71_2;
	wire w_dff_A_g05iV4qr9_1;
	wire w_dff_A_umsvQfiS2_2;
	wire w_dff_A_K6d3lJfk5_1;
	wire w_dff_A_CwMNRSJ39_2;
	wire w_dff_A_6CZxVukQ2_0;
	wire w_dff_B_J4fIGD0M8_1;
	wire w_dff_B_jPvxMSUl7_1;
	wire w_dff_A_a3DYy5kJ1_0;
	wire w_dff_A_WDwUZNW40_0;
	wire w_dff_A_JOkU9xyp2_0;
	wire w_dff_A_5RAOQJeX5_0;
	wire w_dff_A_RDfsVM6X2_1;
	wire w_dff_A_PjIXy07J6_1;
	wire w_dff_A_L84Mh0M65_1;
	wire w_dff_A_1SfBBiXl2_1;
	wire w_dff_A_WTBqrzoc1_1;
	wire w_dff_A_G6lbEGdA0_1;
	wire w_dff_A_pJCGRX3l2_2;
	wire w_dff_A_WL2r15fE7_2;
	wire w_dff_A_yGjiDEl32_2;
	wire w_dff_A_jWocplEn0_2;
	wire w_dff_A_4WsIfzAC9_0;
	wire w_dff_B_PzdBPeFS4_1;
	wire w_dff_B_ESW2Jyin8_1;
	wire w_dff_A_cQwm38V27_0;
	wire w_dff_A_Q5zt9qC28_1;
	wire w_dff_A_HpUvt8bN7_1;
	wire w_dff_A_L1bi1yru6_2;
	wire w_dff_A_iVswdcIQ0_2;
	wire w_dff_A_zsQn6rAz9_1;
	wire w_dff_A_6xE1kp3C5_1;
	wire w_dff_A_yPEI7Z7s6_1;
	wire w_dff_A_IxdqBATw2_1;
	wire w_dff_A_CvTLzAgQ6_2;
	wire w_dff_A_145FCC1R1_0;
	wire w_dff_A_E0jDH5bB5_0;
	wire w_dff_A_9326LpdF4_0;
	wire w_dff_A_BKERlw5H5_0;
	wire w_dff_A_93DnRBLx5_1;
	wire w_dff_A_6JXrWEu75_1;
	wire w_dff_A_fxjrjCh67_1;
	wire w_dff_A_jKyhf4HO5_2;
	wire w_dff_A_3rQhbg9g1_2;
	wire w_dff_A_1AEaBP9I6_2;
	wire w_dff_A_93tWPI9q8_2;
	wire w_dff_A_xBie47Qk2_1;
	wire w_dff_A_EmzcZY9t8_2;
	wire w_dff_A_y5HQIe6X9_0;
	wire w_dff_A_5gdKQzfI4_2;
	wire w_dff_A_MYR8O7PY4_0;
	wire w_dff_A_tBnMUCjT0_0;
	wire w_dff_A_ca1oavqp1_0;
	wire w_dff_A_gnnwhmDU5_0;
	wire w_dff_A_mzXovG4n0_0;
	wire w_dff_A_0hup6JtJ1_0;
	wire w_dff_A_s8Cwsbp59_0;
	wire w_dff_A_9J9gV7LA9_0;
	wire w_dff_A_UMSDBrGl4_0;
	wire w_dff_A_vPrnZUAq7_0;
	wire w_dff_A_c9obuGxY8_0;
	wire w_dff_A_zdrI3PDS9_1;
	wire w_dff_A_BoMi0olI2_0;
	wire w_dff_A_nvTaLphW4_0;
	wire w_dff_A_QsJjPFXN5_0;
	wire w_dff_A_j3O89ShG0_0;
	wire w_dff_A_S0vDBA0J9_0;
	wire w_dff_A_iW9HFaD08_0;
	wire w_dff_A_rrccWHtp0_0;
	wire w_dff_A_Ikjyje7n8_2;
	wire w_dff_A_TOXxie9F4_2;
	wire w_dff_A_apl4wpDY6_2;
	wire w_dff_A_WaRh8NRP3_2;
	wire w_dff_A_fYJv7fYP2_2;
	wire w_dff_A_lIlX7Wn50_2;
	wire w_dff_A_LJliNtAy7_2;
	wire w_dff_A_1bp8sStG3_2;
	wire w_dff_A_3DLSZKbP5_2;
	wire w_dff_A_mYHbTfFD9_2;
	wire w_dff_A_szsVc30w8_2;
	wire w_dff_A_F3pXSx5e6_2;
	wire w_dff_A_MUqtxYMl0_2;
	wire w_dff_A_WcsDrtic9_2;
	wire w_dff_A_IvX1SISW3_2;
	wire w_dff_A_lAQC2soE4_2;
	wire w_dff_A_tRXZgcD47_2;
	wire w_dff_A_ZKRb0Opf1_2;
	wire w_dff_A_A9I8q0GE3_2;
	wire w_dff_A_ppyogrIt4_1;
	wire w_dff_A_8b3QS6fT7_1;
	wire w_dff_A_uJdOCJWZ0_1;
	wire w_dff_A_Ie5jSKVK5_1;
	wire w_dff_A_b6C8S39j3_1;
	wire w_dff_A_ciBTzmfd6_1;
	wire w_dff_A_7wqJ9Bsa1_1;
	wire w_dff_A_VVDAx3uY1_1;
	wire w_dff_A_AD2tdsOF8_1;
	wire w_dff_A_4Xvbbywf5_1;
	wire w_dff_A_quyEqx870_1;
	wire w_dff_A_SJc8o4by1_1;
	wire w_dff_A_M7vcgRzt2_1;
	wire w_dff_A_oqBQk2bZ4_1;
	wire w_dff_A_jXWACblp2_1;
	wire w_dff_A_I0qaYEYe2_1;
	wire w_dff_A_YkaaOJ3u5_1;
	wire w_dff_A_kmY6zEzX4_2;
	wire w_dff_A_YSXjvyKU1_2;
	wire w_dff_A_WtJarjZg2_2;
	wire w_dff_A_puxkd1286_2;
	wire w_dff_A_LBmRRY814_2;
	wire w_dff_A_VQwgBGOY4_2;
	wire w_dff_A_Dhp9Osxv4_2;
	wire w_dff_A_i7mXiXBc4_2;
	wire w_dff_A_pal6TTlv8_2;
	wire w_dff_A_c6gSTUhR6_2;
	wire w_dff_A_KgaFGU7S5_2;
	wire w_dff_A_UygF6HbI1_1;
	wire w_dff_A_T9Chpajb1_2;
	wire w_dff_B_7NAwkOja3_2;
	wire w_dff_B_RNOSPl9T2_2;
	wire w_dff_B_E8goaBHO6_2;
	wire w_dff_B_kD7A8Gu39_2;
	wire w_dff_B_5VSnKx8E3_2;
	wire w_dff_B_4MJXGFq35_2;
	wire w_dff_B_IgrxV5K80_2;
	wire w_dff_B_SQ4edi7L6_2;
	wire w_dff_B_XO2G3nyv7_2;
	wire w_dff_B_qrXm9Kl65_2;
	wire w_dff_B_0BJ2ic2B4_2;
	wire w_dff_B_W6OUSo1Y4_2;
	wire w_dff_B_ZCsYp7Y29_2;
	wire w_dff_B_myZIM1NK6_2;
	wire w_dff_B_vet7eIdY0_2;
	wire w_dff_B_xwoFjAZC4_2;
	wire w_dff_B_265D6Uep9_2;
	wire w_dff_B_ZbQa7PCp5_2;
	wire w_dff_B_tzjSzFk76_2;
	wire w_dff_B_J7FJ6BEE5_2;
	wire w_dff_B_FNrz4wUl8_2;
	wire w_dff_B_6IqE0GFm7_2;
	wire w_dff_B_jW1C4NRR4_2;
	wire w_dff_B_XDizpPKl7_2;
	wire w_dff_A_PxRY2uzP1_2;
	wire w_dff_A_RDqLBym93_2;
	wire w_dff_A_SsyNtHW39_2;
	wire w_dff_A_5fuBd4Rc0_2;
	wire w_dff_A_2a4lBvd87_2;
	wire w_dff_A_lj9TLTIy0_2;
	wire w_dff_A_0VuRgy847_2;
	wire w_dff_A_YrtCm23Q6_2;
	wire w_dff_A_WAFqwUEP9_2;
	wire w_dff_A_LD2TpBWz4_2;
	wire w_dff_A_k2vTd8Xu7_2;
	wire w_dff_A_KA52KHCR6_2;
	wire w_dff_A_NGxsdPAI3_2;
	wire w_dff_A_UaBDrsHk9_2;
	wire w_dff_A_Sz8mgOhv0_2;
	wire w_dff_A_dUYkmnTs3_2;
	wire w_dff_A_FGNPx9p15_2;
	wire w_dff_A_i4GR8iVn4_2;
	wire w_dff_A_DUw5Epjj0_2;
	wire w_dff_A_hhI9bfnN0_2;
	wire w_dff_A_zy1gQ3ov1_2;
	wire w_dff_A_Uyj3YvV44_2;
	wire w_dff_A_LoVGMRWh5_2;
	wire w_dff_A_fuRUgZwW6_0;
	wire w_dff_A_pHqyWyMF6_0;
	wire w_dff_A_BA92vPRz0_0;
	wire w_dff_A_bhah2Hxn6_0;
	wire w_dff_A_sKt9M6kK5_0;
	wire w_dff_A_q9h7freb6_0;
	wire w_dff_A_e9Y3whVb1_0;
	wire w_dff_A_SscALKln3_0;
	wire w_dff_A_mv9Qe9hZ8_0;
	wire w_dff_A_5RacaMh79_0;
	wire w_dff_A_OhqbPePe9_0;
	wire w_dff_A_yfeF5XSX1_0;
	wire w_dff_A_hhoDlKC51_0;
	wire w_dff_A_cag0b5qf4_0;
	wire w_dff_A_PasI4ITh8_0;
	wire w_dff_A_Y7lYWyOM7_0;
	wire w_dff_A_hyar6FWU7_1;
	wire w_dff_A_L5vcJehQ6_1;
	wire w_dff_A_OCY1RXdO1_1;
	wire w_dff_A_jRZYI5ML9_1;
	wire w_dff_A_fN4BFm7N2_1;
	wire w_dff_A_KRs8Gbmq9_1;
	wire w_dff_A_tgGPUvU04_1;
	wire w_dff_A_4elJ960V5_1;
	wire w_dff_A_SxVrNxLb4_1;
	wire w_dff_A_QQuo31aY2_1;
	wire w_dff_A_qfPzuRhQ3_1;
	wire w_dff_A_cb5G565l2_1;
	wire w_dff_A_3RHCVIMc4_0;
	wire w_dff_A_ISAWvOxo3_0;
	wire w_dff_A_9Y9yy8zR4_0;
	wire w_dff_A_3irR0KP65_0;
	wire w_dff_A_JhPOMwGL6_0;
	wire w_dff_A_hYbRxPIL1_0;
	wire w_dff_A_mSDgAZtS5_0;
	wire w_dff_A_1nelbSrb4_0;
	wire w_dff_A_y309zFKo4_0;
	wire w_dff_A_B5kI9FwV9_0;
	wire w_dff_A_ny7ajQjk6_0;
	wire w_dff_A_AJE5QduK8_0;
	wire w_dff_A_t07HMYYV8_0;
	wire w_dff_A_Vn6bD5F74_0;
	wire w_dff_A_sQKv8hqb0_0;
	wire w_dff_A_XFJScwnh8_0;
	wire w_dff_A_PLWBdEet3_0;
	wire w_dff_A_xeKRPcYs3_0;
	wire w_dff_A_p16RC3072_0;
	wire w_dff_A_oizumvxp6_0;
	wire w_dff_A_0HHe19PL3_0;
	wire w_dff_A_AstgGGaD1_0;
	wire w_dff_A_pCLflLim8_0;
	wire w_dff_A_4HYNfnur1_0;
	wire w_dff_A_HUppY1yx4_1;
	wire w_dff_A_JkxxEBys7_0;
	wire w_dff_A_q0n3POXW3_0;
	wire w_dff_A_cehktUxD0_0;
	wire w_dff_A_M44KfxPO4_0;
	wire w_dff_A_5bBBem6b8_0;
	wire w_dff_A_GPrB7LAM2_0;
	wire w_dff_A_TGBFibZw6_0;
	wire w_dff_A_apRmpxY45_0;
	wire w_dff_A_T89OFW921_0;
	wire w_dff_A_8yYH2IQ27_0;
	wire w_dff_A_R4kJCjqO1_0;
	wire w_dff_A_q9P3EMcU5_0;
	wire w_dff_A_PCp7I8GM7_0;
	wire w_dff_A_VsAtRIEU7_0;
	wire w_dff_A_hIBPr7HU2_0;
	wire w_dff_A_0c2WevMi6_0;
	wire w_dff_A_x2swy0xC4_0;
	wire w_dff_A_Q5s0T84Y1_0;
	wire w_dff_A_SZdqoSlS9_0;
	wire w_dff_A_Ih4eRD3R7_0;
	wire w_dff_A_ViwAE7JN3_0;
	wire w_dff_A_wIcM7nXD6_0;
	wire w_dff_A_gR3xRhPa6_0;
	wire w_dff_A_s7fIBDsj0_0;
	wire w_dff_A_bgbfZxUg8_1;
	wire w_dff_A_3iukpOH64_0;
	wire w_dff_A_N2tLGc6e0_0;
	wire w_dff_A_382wXYrB6_0;
	wire w_dff_A_wognC2Q89_0;
	wire w_dff_A_DmT4I2r63_0;
	wire w_dff_A_AQZkrOwm2_0;
	wire w_dff_A_UTpaR8fz6_0;
	wire w_dff_A_wrgdHrHz8_0;
	wire w_dff_A_HdUoc6hb0_0;
	wire w_dff_A_Zwd2PX9a0_0;
	wire w_dff_A_2BwNehvp7_0;
	wire w_dff_A_0h2tkLmC1_0;
	wire w_dff_A_iXK43Zs41_0;
	wire w_dff_A_OmLbW4Iy4_0;
	wire w_dff_A_HubVTvWd0_0;
	wire w_dff_A_KxWanDai5_0;
	wire w_dff_A_hIH32iKu8_0;
	wire w_dff_A_4PpY3odB6_0;
	wire w_dff_A_qb9watoE0_0;
	wire w_dff_A_DDikxFB50_0;
	wire w_dff_A_0HXgrLo47_0;
	wire w_dff_A_ioyeN63Z6_0;
	wire w_dff_A_JN965QCk0_0;
	wire w_dff_A_a7Abiasf0_0;
	wire w_dff_A_xnuHcXtR9_1;
	wire w_dff_A_Spw7PSBT8_0;
	wire w_dff_A_Xd0gO3jg3_0;
	wire w_dff_A_dYJW6aHA3_0;
	wire w_dff_A_wyOinnPZ9_0;
	wire w_dff_A_FAJL4wXN9_0;
	wire w_dff_A_UqfFpiUn5_0;
	wire w_dff_A_waGytCvG3_0;
	wire w_dff_A_d59ubn9F1_0;
	wire w_dff_A_NaNrlEHF1_0;
	wire w_dff_A_seAYEsp76_0;
	wire w_dff_A_T1823c4M5_0;
	wire w_dff_A_PHux2mT88_0;
	wire w_dff_A_GkeuVsPt3_0;
	wire w_dff_A_LXypeAx94_0;
	wire w_dff_A_He3iXIhu0_0;
	wire w_dff_A_dhrAaJGI9_0;
	wire w_dff_A_5jo1I6l73_0;
	wire w_dff_A_iVV58X7c6_0;
	wire w_dff_A_WSa20qeo2_0;
	wire w_dff_A_xkFAl7Fg1_0;
	wire w_dff_A_9CD5bB7k9_0;
	wire w_dff_A_JVyna9ul2_0;
	wire w_dff_A_RPmdp4rG3_0;
	wire w_dff_A_S8O1fbJY7_0;
	wire w_dff_A_ywNt4EiO1_1;
	wire w_dff_A_VVNM3nxk7_0;
	wire w_dff_A_mmjtDoSM2_0;
	wire w_dff_A_b2Sh4jsb2_0;
	wire w_dff_A_6hYJGPOL7_0;
	wire w_dff_A_5umprcy05_0;
	wire w_dff_A_D5UXYMnK7_0;
	wire w_dff_A_bMwFVns33_0;
	wire w_dff_A_40wmxGgT3_0;
	wire w_dff_A_fgKMQkj48_0;
	wire w_dff_A_0ZQxhR5e9_0;
	wire w_dff_A_8dPtbYpI0_0;
	wire w_dff_A_Fq3HN0CL1_0;
	wire w_dff_A_Bd05Wsy23_0;
	wire w_dff_A_ALM58iN24_0;
	wire w_dff_A_6t3ZeJx36_0;
	wire w_dff_A_g3hPaqWW1_0;
	wire w_dff_A_vz1QgAqq4_0;
	wire w_dff_A_klPbOt779_0;
	wire w_dff_A_XQsxFS3V8_0;
	wire w_dff_A_iP1vrYH23_0;
	wire w_dff_A_koqwoAFO7_0;
	wire w_dff_A_LkXpchdi4_0;
	wire w_dff_A_IOYig3dL4_0;
	wire w_dff_A_RiPmO5jO7_0;
	wire w_dff_A_wEbXZwDn0_1;
	wire w_dff_A_HSvLcFhP5_0;
	wire w_dff_A_BCZSTrqm4_0;
	wire w_dff_A_311DW8Cb4_0;
	wire w_dff_A_EM8T03Ww0_0;
	wire w_dff_A_7mfxGjPM5_0;
	wire w_dff_A_yGoa4VFG3_0;
	wire w_dff_A_BCLyTzPz5_0;
	wire w_dff_A_dSxoOqCP5_0;
	wire w_dff_A_AaFa3NAg8_0;
	wire w_dff_A_onjYlMBl9_0;
	wire w_dff_A_XfTgz1Vg6_0;
	wire w_dff_A_JncHxJWa5_0;
	wire w_dff_A_1g6dkrv70_0;
	wire w_dff_A_Yvh6AOlh0_0;
	wire w_dff_A_aSNyovvN8_0;
	wire w_dff_A_Ev5iRoSw1_0;
	wire w_dff_A_ENUbs8W56_0;
	wire w_dff_A_Wuoudu227_0;
	wire w_dff_A_rJulTKrw4_0;
	wire w_dff_A_gOIlfFh00_0;
	wire w_dff_A_NwZT58qA1_0;
	wire w_dff_A_shR6BZ6X7_0;
	wire w_dff_A_YY9zUnjr2_0;
	wire w_dff_A_jrqvbr3c8_0;
	wire w_dff_A_XBKdFEY12_1;
	wire w_dff_A_W3blJKaT6_0;
	wire w_dff_A_m5lxHlBy9_0;
	wire w_dff_A_hDxQ0zxn9_0;
	wire w_dff_A_Hlx88qOv2_0;
	wire w_dff_A_SRZmYHN44_0;
	wire w_dff_A_j8WvfXCf3_0;
	wire w_dff_A_hGPvJOyA4_0;
	wire w_dff_A_1CGvhTYl6_0;
	wire w_dff_A_y4T2JSsi1_0;
	wire w_dff_A_ghNw8vfW5_0;
	wire w_dff_A_lQLqOei06_0;
	wire w_dff_A_3un9PmG75_0;
	wire w_dff_A_U8ZpNnbz5_0;
	wire w_dff_A_CQI7aj3O9_0;
	wire w_dff_A_PymAOf9O4_0;
	wire w_dff_A_WFBKwnf95_0;
	wire w_dff_A_bUgXr9FK0_0;
	wire w_dff_A_5ga8yakY1_0;
	wire w_dff_A_jyezGBJM0_0;
	wire w_dff_A_ADE6YPIK2_0;
	wire w_dff_A_ZMSHaKc78_0;
	wire w_dff_A_StMOIgqG7_0;
	wire w_dff_A_VVPO2BMh9_0;
	wire w_dff_A_oe8Go6Nb7_0;
	wire w_dff_A_5UiApBuf0_1;
	wire w_dff_A_ZOfNn9lZ0_0;
	wire w_dff_A_pCIAjKVy3_0;
	wire w_dff_A_lfRHEVvT8_0;
	wire w_dff_A_CCsFULqC1_0;
	wire w_dff_A_q26Ia2Vz8_0;
	wire w_dff_A_txdgd2aV0_0;
	wire w_dff_A_Tqyn0PGs2_0;
	wire w_dff_A_PupEY9tU4_0;
	wire w_dff_A_GulXQyOr1_0;
	wire w_dff_A_VwJ7xpip8_0;
	wire w_dff_A_JiNepxSR2_0;
	wire w_dff_A_fdfoUjCQ8_0;
	wire w_dff_A_evjQ1GOQ6_0;
	wire w_dff_A_Ai2LZgHB2_0;
	wire w_dff_A_qkThCd3n6_0;
	wire w_dff_A_wP7OkQIs7_0;
	wire w_dff_A_0gh7OFPG4_0;
	wire w_dff_A_Bc87HXuD6_0;
	wire w_dff_A_IXJSGref9_0;
	wire w_dff_A_3RJ4Z2zp8_0;
	wire w_dff_A_nZsYqJsJ8_0;
	wire w_dff_A_jmvhyzkZ3_0;
	wire w_dff_A_TZvXZ9uQ0_0;
	wire w_dff_A_uHLArAq26_0;
	wire w_dff_A_lAjJ6ntN2_1;
	wire w_dff_A_gX4l8LdO0_0;
	wire w_dff_A_Ez6ANdeV7_0;
	wire w_dff_A_0KZsZlnI4_0;
	wire w_dff_A_dLJb00FY5_0;
	wire w_dff_A_UJcq1LMn1_0;
	wire w_dff_A_lD83Iwof9_0;
	wire w_dff_A_Nx1kym4p3_0;
	wire w_dff_A_QavivzIi6_0;
	wire w_dff_A_2t2VTaDi9_0;
	wire w_dff_A_CDtK9NDC3_0;
	wire w_dff_A_MJ9UoudK5_0;
	wire w_dff_A_btQjM91A6_0;
	wire w_dff_A_ncjZG1842_0;
	wire w_dff_A_BTtIqM3W0_0;
	wire w_dff_A_YPsrmVI95_0;
	wire w_dff_A_efGUEy068_0;
	wire w_dff_A_XMI3Hs1t2_0;
	wire w_dff_A_43dXQUqv6_0;
	wire w_dff_A_c6UIM3pj6_0;
	wire w_dff_A_t6VnbjB46_0;
	wire w_dff_A_saPPbtAo1_0;
	wire w_dff_A_woxLorAt1_0;
	wire w_dff_A_xC83BlN51_0;
	wire w_dff_A_yFnvOrBl4_0;
	wire w_dff_A_0HHr3PS48_1;
	wire w_dff_A_Qmt1iINc8_0;
	wire w_dff_A_aEUtmnu55_0;
	wire w_dff_A_68hFG8kh9_0;
	wire w_dff_A_i1ZtKfQ55_0;
	wire w_dff_A_02bHml4r6_0;
	wire w_dff_A_1D89T5S51_0;
	wire w_dff_A_1eccpagy6_0;
	wire w_dff_A_69nOebat5_0;
	wire w_dff_A_NrxZeAKF7_0;
	wire w_dff_A_DhUKxEso9_0;
	wire w_dff_A_IhPRGPGP1_0;
	wire w_dff_A_RqErZqyq3_0;
	wire w_dff_A_mvELn8jo3_0;
	wire w_dff_A_XLzwTO640_0;
	wire w_dff_A_WbG5VX9j6_0;
	wire w_dff_A_PcQC7G1V9_0;
	wire w_dff_A_yXkrA4Gj0_0;
	wire w_dff_A_lg24CHzt4_0;
	wire w_dff_A_U4yiVyUN6_0;
	wire w_dff_A_IuxKDhvs7_0;
	wire w_dff_A_uJSbDNmw2_0;
	wire w_dff_A_9D16R5mB7_0;
	wire w_dff_A_nqZkEy4U6_0;
	wire w_dff_A_ALW4vH0j8_0;
	wire w_dff_A_pVw4klAf8_1;
	wire w_dff_A_QLZW3LF36_0;
	wire w_dff_A_U6fvBceE8_0;
	wire w_dff_A_j2UNdXJB2_0;
	wire w_dff_A_mhqfB2Nq4_0;
	wire w_dff_A_lvme9Jct0_0;
	wire w_dff_A_jJFicvkV8_0;
	wire w_dff_A_6YMLwFrZ2_0;
	wire w_dff_A_ja7oAzQ41_0;
	wire w_dff_A_nGvgUjE06_0;
	wire w_dff_A_24EAdmNA6_0;
	wire w_dff_A_GZdqD08q0_0;
	wire w_dff_A_4VY4z9Pt4_0;
	wire w_dff_A_il4hTyVm3_0;
	wire w_dff_A_ZEhDEe0d7_0;
	wire w_dff_A_RST6M91K4_0;
	wire w_dff_A_NxDDcVaf2_0;
	wire w_dff_A_dvmq6JXW8_0;
	wire w_dff_A_NQkEYQCw9_0;
	wire w_dff_A_BKhPLSCs0_0;
	wire w_dff_A_JPzGiUwV2_0;
	wire w_dff_A_l2wvO4NR9_0;
	wire w_dff_A_W2E9JpJS4_0;
	wire w_dff_A_YI2X50pv5_0;
	wire w_dff_A_XqTn1v4h0_0;
	wire w_dff_A_Kl1VYOge1_1;
	wire w_dff_A_B3EwKRTa9_0;
	wire w_dff_A_rbVVryLn6_0;
	wire w_dff_A_c6k24Z1B1_0;
	wire w_dff_A_2SynLc0q1_0;
	wire w_dff_A_O3rLhcNa3_0;
	wire w_dff_A_YFCZmZn02_0;
	wire w_dff_A_DE6c4i8X6_0;
	wire w_dff_A_NeIydeCE1_0;
	wire w_dff_A_2Gutarxx1_0;
	wire w_dff_A_NuPQ2fAM5_0;
	wire w_dff_A_GwN5urio6_0;
	wire w_dff_A_k0m57NFn4_0;
	wire w_dff_A_MRZmuARF4_0;
	wire w_dff_A_veRZFaGf5_0;
	wire w_dff_A_EXIBH7FF2_0;
	wire w_dff_A_AtIWkV7A8_0;
	wire w_dff_A_TFfMWMZO1_0;
	wire w_dff_A_iLXbjr3R9_0;
	wire w_dff_A_d4aptmOa9_0;
	wire w_dff_A_q2MZOYAs3_0;
	wire w_dff_A_KMZPdXSE5_0;
	wire w_dff_A_BbSM9Wij0_0;
	wire w_dff_A_hlhQvUvX2_0;
	wire w_dff_A_6NRR88zZ4_0;
	wire w_dff_A_xWfJIjhY9_2;
	wire w_dff_A_W4QEECt23_0;
	wire w_dff_A_MXJCNFNP1_0;
	wire w_dff_A_cSP4Twnl9_0;
	wire w_dff_A_iXMe5Czr1_0;
	wire w_dff_A_xFIVFouJ1_0;
	wire w_dff_A_0gMiaVB54_0;
	wire w_dff_A_9jo7rlqd1_0;
	wire w_dff_A_3JCQ8Gq22_0;
	wire w_dff_A_Ax7jbXJF4_0;
	wire w_dff_A_nFmYb7tG1_0;
	wire w_dff_A_6VGXosrO9_0;
	wire w_dff_A_R0wUTnBv8_0;
	wire w_dff_A_qw6D6rlu2_0;
	wire w_dff_A_OioMYsVH6_0;
	wire w_dff_A_Pfcmgsu95_0;
	wire w_dff_A_i8mtKWq51_0;
	wire w_dff_A_IsSgKvSD1_0;
	wire w_dff_A_uzhGcz4w8_0;
	wire w_dff_A_HsMeHz2e6_0;
	wire w_dff_A_n5iaUi1I4_0;
	wire w_dff_A_TXXm7fNr1_0;
	wire w_dff_A_r6nBd33b4_0;
	wire w_dff_A_7eHj7Vmb0_0;
	wire w_dff_A_aMOluZcQ8_0;
	wire w_dff_A_DKH03zRr9_1;
	wire w_dff_A_V9Dl4hlm9_0;
	wire w_dff_A_ZevjiADK7_0;
	wire w_dff_A_YH5oIzoM3_0;
	wire w_dff_A_TYuXSnAM2_0;
	wire w_dff_A_ubolZQDz4_0;
	wire w_dff_A_J1c3ZeLx1_0;
	wire w_dff_A_OCHDOgu56_0;
	wire w_dff_A_wU3Gi6uw6_0;
	wire w_dff_A_5z0GlFRk3_0;
	wire w_dff_A_ISNGNLqq6_0;
	wire w_dff_A_itNXrn802_0;
	wire w_dff_A_Cjtrg6io1_0;
	wire w_dff_A_xtaWXGfw8_0;
	wire w_dff_A_SugRY9d51_0;
	wire w_dff_A_fXetze8D1_0;
	wire w_dff_A_PoTC19mg5_0;
	wire w_dff_A_dOIkIvFI4_0;
	wire w_dff_A_qYYjo8Di4_0;
	wire w_dff_A_50UqEfcW1_0;
	wire w_dff_A_enR1XClG3_0;
	wire w_dff_A_9S2mwn7J5_0;
	wire w_dff_A_RpaTGwKC1_0;
	wire w_dff_A_lo72eVtF8_0;
	wire w_dff_A_0TcMbMkW1_0;
	wire w_dff_A_C4E6I9xm8_1;
	wire w_dff_A_J3wecKfl8_0;
	wire w_dff_A_PVdshIEX2_0;
	wire w_dff_A_9tqw22TR0_0;
	wire w_dff_A_o3O10GqH6_0;
	wire w_dff_A_VKsIspZl5_0;
	wire w_dff_A_w7nMf7iq6_0;
	wire w_dff_A_gD03OdNp1_0;
	wire w_dff_A_pWObaypn4_0;
	wire w_dff_A_JhTP2HUO8_0;
	wire w_dff_A_vNHZzIe48_0;
	wire w_dff_A_LcUEyZrV4_0;
	wire w_dff_A_tb1jacsR7_0;
	wire w_dff_A_KIy3WwXd8_0;
	wire w_dff_A_K1ZQVDtw3_0;
	wire w_dff_A_JprNTZPk2_0;
	wire w_dff_A_QObp4Vzv6_0;
	wire w_dff_A_uFxb5Z0a8_0;
	wire w_dff_A_mfr59jnh5_0;
	wire w_dff_A_hmAAue0G0_0;
	wire w_dff_A_KhmX7SqM9_0;
	wire w_dff_A_82TbgnjM3_0;
	wire w_dff_A_qur3YhbT2_0;
	wire w_dff_A_PgAh9jYo8_0;
	wire w_dff_A_vJqoAf853_0;
	wire w_dff_A_IneqafsU3_1;
	wire w_dff_A_bdp2HV5j4_0;
	wire w_dff_A_ZMxhpMte3_0;
	wire w_dff_A_T24lEb8t1_0;
	wire w_dff_A_zDmCoZu30_0;
	wire w_dff_A_woHPVkCV7_0;
	wire w_dff_A_s6T66enI5_0;
	wire w_dff_A_60S9acg72_0;
	wire w_dff_A_IsYTu06N0_0;
	wire w_dff_A_CDoPbfqB5_0;
	wire w_dff_A_wB8aa1u45_0;
	wire w_dff_A_SpKjj8Rh2_0;
	wire w_dff_A_FiJF7Unv8_0;
	wire w_dff_A_PUkP4kX68_0;
	wire w_dff_A_HpCYed7l8_0;
	wire w_dff_A_HP3KpLfy3_0;
	wire w_dff_A_utArNpwp5_0;
	wire w_dff_A_nn2F6oWB8_0;
	wire w_dff_A_wFixckNx2_0;
	wire w_dff_A_DcnDZqoU9_0;
	wire w_dff_A_fnWcAW433_0;
	wire w_dff_A_j6BIrdjI5_0;
	wire w_dff_A_zF1ysYqI0_0;
	wire w_dff_A_JSZIW3jV1_0;
	wire w_dff_A_kfRy5ahu9_0;
	wire w_dff_A_1xSfMYMt0_1;
	wire w_dff_A_9LKRB3f68_0;
	wire w_dff_A_gc0i5aTx3_0;
	wire w_dff_A_ZnFsmU7S4_0;
	wire w_dff_A_LXhdFnde2_0;
	wire w_dff_A_OK9feKSz0_0;
	wire w_dff_A_teOyDpbz2_0;
	wire w_dff_A_P1SAHPB60_0;
	wire w_dff_A_agHq9Vxe8_0;
	wire w_dff_A_W6mCaI3z2_0;
	wire w_dff_A_8vAThO435_0;
	wire w_dff_A_eP8CBvWY0_0;
	wire w_dff_A_lJPviwf89_0;
	wire w_dff_A_KQClxOC20_0;
	wire w_dff_A_xYtiwiq53_0;
	wire w_dff_A_jROIc4bY6_0;
	wire w_dff_A_V1qaUMme6_0;
	wire w_dff_A_jAtJSnBV4_0;
	wire w_dff_A_Q4j7EZNm1_0;
	wire w_dff_A_dGN7hzBT7_0;
	wire w_dff_A_hR5xHatP1_0;
	wire w_dff_A_FszJodIF2_0;
	wire w_dff_A_mAvnTKmL2_0;
	wire w_dff_A_S6IQxkHY2_0;
	wire w_dff_A_aqqtuCRt9_0;
	wire w_dff_A_ZCfZqptZ2_2;
	wire w_dff_A_AkxK3PXr7_0;
	wire w_dff_A_j94OQCS04_0;
	wire w_dff_A_cQBw3GLb0_0;
	wire w_dff_A_ysenTGml1_0;
	wire w_dff_A_AxYT9JZM0_0;
	wire w_dff_A_hKYqQDsu7_0;
	wire w_dff_A_1r1Xn5aR6_0;
	wire w_dff_A_q78m1Ni15_0;
	wire w_dff_A_FOJ9xqi72_0;
	wire w_dff_A_oWZFgUY55_0;
	wire w_dff_A_Zct95VyD4_0;
	wire w_dff_A_Yl725GGn9_0;
	wire w_dff_A_4vRX5qte9_0;
	wire w_dff_A_TzdtOuMs7_0;
	wire w_dff_A_ZsjCNNIt6_0;
	wire w_dff_A_sNtzgHPm3_0;
	wire w_dff_A_W3L6Sddn7_0;
	wire w_dff_A_UAHvOLWt6_0;
	wire w_dff_A_J7uiRwTk6_0;
	wire w_dff_A_l6pT0S5f5_0;
	wire w_dff_A_yXpblTTG0_0;
	wire w_dff_A_uS9K5RRB1_0;
	wire w_dff_A_Xtw3kVUu5_0;
	wire w_dff_A_dlMMGcj04_0;
	wire w_dff_A_85EWI87F1_2;
	wire w_dff_A_wUlp3ZHb7_0;
	wire w_dff_A_CtFMHTU65_0;
	wire w_dff_A_VRHQM1D97_0;
	wire w_dff_A_vuJDotK36_0;
	wire w_dff_A_smtJ0N6p1_0;
	wire w_dff_A_nVzTU1wv0_0;
	wire w_dff_A_vgYyKTxe5_0;
	wire w_dff_A_CbaKDPNt4_0;
	wire w_dff_A_NJXZjmGw5_0;
	wire w_dff_A_U8hkgIES8_0;
	wire w_dff_A_aCh7I36M3_0;
	wire w_dff_A_gVs8XcDN0_0;
	wire w_dff_A_zkZJzAKK1_0;
	wire w_dff_A_2EEfBfON7_0;
	wire w_dff_A_m8vJpnEV2_0;
	wire w_dff_A_uUKXjEl93_0;
	wire w_dff_A_RAsSNRWz7_0;
	wire w_dff_A_NTzsG20u9_0;
	wire w_dff_A_H8wcQRyh4_0;
	wire w_dff_A_L6kVtjQ69_0;
	wire w_dff_A_RRt0yPzE5_0;
	wire w_dff_A_7o8UcTC54_0;
	wire w_dff_A_0ncU4kYV4_0;
	wire w_dff_A_wbIT1XPG9_2;
	wire w_dff_A_vgwIbBju5_0;
	wire w_dff_A_bkFvrZ5J3_0;
	wire w_dff_A_xRcw8JG86_0;
	wire w_dff_A_kbBSzTe02_0;
	wire w_dff_A_7bH0luB35_0;
	wire w_dff_A_zHxniMfJ0_0;
	wire w_dff_A_GXJk6YgY3_0;
	wire w_dff_A_DklyxYxz6_0;
	wire w_dff_A_5J3lHr7j0_0;
	wire w_dff_A_gkAYmFWb4_0;
	wire w_dff_A_Z9izDOnl8_0;
	wire w_dff_A_2UoyOGkc1_0;
	wire w_dff_A_besySP5H1_0;
	wire w_dff_A_T1cYBKAv7_0;
	wire w_dff_A_DWjNw2ar2_0;
	wire w_dff_A_yiRhqAu64_0;
	wire w_dff_A_3s9vnMc08_0;
	wire w_dff_A_1XzhlFWJ2_0;
	wire w_dff_A_wSKLq0gu0_0;
	wire w_dff_A_BCZp0mBa3_0;
	wire w_dff_A_uApHQBbg7_0;
	wire w_dff_A_es2KX2yR9_0;
	wire w_dff_A_frJMrqSo1_0;
	wire w_dff_A_baaaIop22_1;
	wire w_dff_A_qHT3LPmz5_0;
	wire w_dff_A_zMglTbSo5_0;
	wire w_dff_A_h9dnR1xR0_0;
	wire w_dff_A_Wb0DyuPT7_0;
	wire w_dff_A_rn7xnLiI9_0;
	wire w_dff_A_gpoeS98b4_0;
	wire w_dff_A_cJHceGsL9_0;
	wire w_dff_A_u3soHglQ8_0;
	wire w_dff_A_XrlUDqrv8_0;
	wire w_dff_A_3yjouAZG0_0;
	wire w_dff_A_jwnGBlz66_0;
	wire w_dff_A_NqnhHSnG4_0;
	wire w_dff_A_ZzH1PtJZ5_0;
	wire w_dff_A_x7LHgaJv8_0;
	wire w_dff_A_VZvGSK4Y3_0;
	wire w_dff_A_TYHC74x96_0;
	wire w_dff_A_23nFjEDI6_0;
	wire w_dff_A_ET4TfNhs6_0;
	wire w_dff_A_yMhm8xQV2_0;
	wire w_dff_A_Pco2ROqo6_0;
	wire w_dff_A_pv6D1KCd8_0;
	wire w_dff_A_WHxedDe84_0;
	wire w_dff_A_Q52y1VST8_0;
	wire w_dff_A_0NtsHe4k0_1;
	wire w_dff_A_z8SEhmuw8_0;
	wire w_dff_A_0JW3qpPK1_0;
	wire w_dff_A_uZQRpj9u4_0;
	wire w_dff_A_UOWIhbIO6_0;
	wire w_dff_A_fcI1VUiZ9_0;
	wire w_dff_A_BWbThhkX9_0;
	wire w_dff_A_4qtfWl6m2_0;
	wire w_dff_A_UIUiWn8S4_0;
	wire w_dff_A_fvWGtN4H3_0;
	wire w_dff_A_VgWcOzhL8_0;
	wire w_dff_A_8VCmIRiZ1_0;
	wire w_dff_A_aiG5mRhr7_0;
	wire w_dff_A_rnff7rdv9_0;
	wire w_dff_A_C5fA222u1_0;
	wire w_dff_A_in6rFIyp5_0;
	wire w_dff_A_xHmOpUZn8_0;
	wire w_dff_A_ZO8cscaM6_0;
	wire w_dff_A_N8nSplsF6_0;
	wire w_dff_A_22FwJYlc0_0;
	wire w_dff_A_xbtWDrRh7_0;
	wire w_dff_A_JzC9FgC18_0;
	wire w_dff_A_DhTOD46w3_0;
	wire w_dff_A_0lLBpF6k3_0;
	wire w_dff_A_910Pao2f1_0;
	wire w_dff_A_U6IqrDOA3_1;
	wire w_dff_A_JFuCtzja3_0;
	wire w_dff_A_gBl0FTYb2_0;
	wire w_dff_A_1U6gpGID3_0;
	wire w_dff_A_tzfrMzca0_0;
	wire w_dff_A_7nS1bCmI1_0;
	wire w_dff_A_TxHYNhcK3_0;
	wire w_dff_A_6joH87FZ8_0;
	wire w_dff_A_Q1vsS2BU7_0;
	wire w_dff_A_1lOXF1qY7_0;
	wire w_dff_A_QxvhYoBx7_0;
	wire w_dff_A_SLCOGf525_0;
	wire w_dff_A_4roXJf559_0;
	wire w_dff_A_r1zjsBTd8_0;
	wire w_dff_A_CLtav2Qi1_0;
	wire w_dff_A_WF6cgsK41_0;
	wire w_dff_A_dJChjvxg0_0;
	wire w_dff_A_8ofXVN961_0;
	wire w_dff_A_2WY6iaes8_0;
	wire w_dff_A_PhvR06020_0;
	wire w_dff_A_gZnyTgn10_0;
	wire w_dff_A_OovXxVAL4_0;
	wire w_dff_A_XeYo21uv6_0;
	wire w_dff_A_EoG4hnUo0_0;
	wire w_dff_A_Xe6emeEV6_0;
	wire w_dff_A_NmT0XjCB0_1;
	wire w_dff_A_RZMcr9ml7_0;
	wire w_dff_A_n5rXPReW6_0;
	wire w_dff_A_ixu9Ajnm3_0;
	wire w_dff_A_uawdFRIq5_0;
	wire w_dff_A_97KL3mNg1_0;
	wire w_dff_A_pms3kupZ5_0;
	wire w_dff_A_TRzUWzqA9_0;
	wire w_dff_A_4GOOIoBm5_0;
	wire w_dff_A_ILzC5j1Y5_0;
	wire w_dff_A_2KgoG5uF9_0;
	wire w_dff_A_rCHZvA3y5_0;
	wire w_dff_A_Q8wagKWl2_0;
	wire w_dff_A_vlO09x095_0;
	wire w_dff_A_hHuvKOIz6_0;
	wire w_dff_A_3HceagY58_0;
	wire w_dff_A_SlaJdS6O3_0;
	wire w_dff_A_Z0wJn0BU4_0;
	wire w_dff_A_PMJ4zAW60_0;
	wire w_dff_A_0ZzEXFnr9_0;
	wire w_dff_A_MVqRmjUv6_0;
	wire w_dff_A_iNYzOTkj1_0;
	wire w_dff_A_zC9HvHJF1_0;
	wire w_dff_A_yEObtYBs5_0;
	wire w_dff_A_2jxIV3B49_0;
	wire w_dff_A_FwI0aGbj2_1;
	wire w_dff_A_XHPaJRCE4_0;
	wire w_dff_A_Mhc8ZdV60_0;
	wire w_dff_A_InkJaXhL9_0;
	wire w_dff_A_3k09P2nw0_0;
	wire w_dff_A_ndQSjTAy5_0;
	wire w_dff_A_z4Vz3Q9U8_0;
	wire w_dff_A_MolwkUZP4_0;
	wire w_dff_A_lMu4vz877_0;
	wire w_dff_A_1xNYFVuB7_0;
	wire w_dff_A_92MBFYl93_0;
	wire w_dff_A_A1R43ry02_0;
	wire w_dff_A_mi3U7mX09_0;
	wire w_dff_A_J4z8VsmN4_0;
	wire w_dff_A_cALNuMci9_0;
	wire w_dff_A_tHyB8OW05_0;
	wire w_dff_A_cjPvDO8B7_0;
	wire w_dff_A_1vUF3bQz3_0;
	wire w_dff_A_OwwzloIQ9_0;
	wire w_dff_A_YYP46nOo1_0;
	wire w_dff_A_SuKMQElZ8_0;
	wire w_dff_A_SeUcB0pi6_0;
	wire w_dff_A_TSnMP6gk0_0;
	wire w_dff_A_mIPC2zON9_0;
	wire w_dff_A_9Ueuxn9R0_0;
	wire w_dff_A_IM6ysSsv4_1;
	wire w_dff_A_zY63OBZr1_0;
	wire w_dff_A_ktX1edDQ1_0;
	wire w_dff_A_QJZkZGhW5_0;
	wire w_dff_A_WAeZpLlO6_0;
	wire w_dff_A_A7bdGS0l1_0;
	wire w_dff_A_XlA4f5kQ4_0;
	wire w_dff_A_e4AlmKNp9_0;
	wire w_dff_A_aKQt76y24_0;
	wire w_dff_A_a3EsAeRB6_0;
	wire w_dff_A_PoGMbfkG8_0;
	wire w_dff_A_QJOSBcQ79_0;
	wire w_dff_A_qh2QGmt83_0;
	wire w_dff_A_tPJmWqXF3_0;
	wire w_dff_A_6j2Kddnx8_0;
	wire w_dff_A_VJkgFuuW7_0;
	wire w_dff_A_NmESWnZK6_0;
	wire w_dff_A_SHBUuRdc2_0;
	wire w_dff_A_JV1R3ej42_0;
	wire w_dff_A_7uLaISER7_0;
	wire w_dff_A_Gl01ovTA0_0;
	wire w_dff_A_c9eWRvHJ3_0;
	wire w_dff_A_2zS9LLHd5_0;
	wire w_dff_A_q7TqjPED9_0;
	wire w_dff_A_r9Ba313H0_0;
	wire w_dff_A_ELUGCjOB6_1;
	wire w_dff_A_nCOVKXJW4_0;
	wire w_dff_A_gDFQfVk81_0;
	wire w_dff_A_x1x58NKi6_0;
	wire w_dff_A_DADGKog67_0;
	wire w_dff_A_s3y8BDx91_0;
	wire w_dff_A_adgIwvf93_0;
	wire w_dff_A_uQ4JskQk3_0;
	wire w_dff_A_DdINJAaW6_0;
	wire w_dff_A_3n3LtgKK4_0;
	wire w_dff_A_6ZgYHm3y4_0;
	wire w_dff_A_mBmZXUZ80_0;
	wire w_dff_A_rsAcAc5H9_0;
	wire w_dff_A_XtXrAGbu0_0;
	wire w_dff_A_tyukI0qE2_0;
	wire w_dff_A_DsSsIf3L7_0;
	wire w_dff_A_qHLc86ct6_0;
	wire w_dff_A_shdq50ZH0_0;
	wire w_dff_A_j5IFX4Zg0_0;
	wire w_dff_A_vCy38a642_0;
	wire w_dff_A_VD7wn6bm6_0;
	wire w_dff_A_TJXtEoKU1_0;
	wire w_dff_A_JO5766qF6_0;
	wire w_dff_A_4rNpAa2X8_0;
	wire w_dff_A_Z42TPgXx5_0;
	wire w_dff_A_keD9V7g93_2;
	wire w_dff_A_6No7jZ3l5_0;
	wire w_dff_A_YwCOvnJB1_0;
	wire w_dff_A_e2Zwj5m62_0;
	wire w_dff_A_jj23SIgP4_0;
	wire w_dff_A_IpvWiYMh2_0;
	wire w_dff_A_RRAU7Feh9_0;
	wire w_dff_A_Rs4lQiv80_0;
	wire w_dff_A_TaIA0Syt7_0;
	wire w_dff_A_Xl2iu4F66_0;
	wire w_dff_A_vTMnpaNz6_0;
	wire w_dff_A_D9yertSl6_0;
	wire w_dff_A_Yb8R0NBp9_0;
	wire w_dff_A_zoiV8HqI0_0;
	wire w_dff_A_frH1zcVH3_0;
	wire w_dff_A_jlSvN7Gi6_0;
	wire w_dff_A_l2yUoy9h5_0;
	wire w_dff_A_zoYPNHe88_0;
	wire w_dff_A_bwEjAIaO7_0;
	wire w_dff_A_w7sR6eES9_0;
	wire w_dff_A_AsVarqsG3_0;
	wire w_dff_A_uJzgPcEF4_0;
	wire w_dff_A_PeVg3iqd4_0;
	wire w_dff_A_x86FEGCI7_2;
	wire w_dff_A_QZa27yH73_0;
	wire w_dff_A_b9fGvEec6_0;
	wire w_dff_A_iGk5muXF6_0;
	wire w_dff_A_Gh3424E94_0;
	wire w_dff_A_LCebUzlT4_0;
	wire w_dff_A_PxdHmspX4_0;
	wire w_dff_A_TivC2nGk7_0;
	wire w_dff_A_u9Lazg1R2_0;
	wire w_dff_A_Vsi66rb35_0;
	wire w_dff_A_Z1fiM0vR6_0;
	wire w_dff_A_3NZ0yDjb3_0;
	wire w_dff_A_6SUEWyFS5_0;
	wire w_dff_A_YSCxAza49_0;
	wire w_dff_A_BlGFREtI4_0;
	wire w_dff_A_s5FtIMzv5_0;
	wire w_dff_A_00AvwFTZ2_0;
	wire w_dff_A_hhMxq2Tc8_0;
	wire w_dff_A_fMEkWrrV5_0;
	wire w_dff_A_rkNNEXs64_0;
	wire w_dff_A_aOJlDXK89_0;
	wire w_dff_A_vS5vbLYA1_0;
	wire w_dff_A_KofkMd3a9_0;
	wire w_dff_A_0g7TGgoS7_0;
	wire w_dff_A_YeaIpaov7_1;
	wire w_dff_A_jiXK9IhC9_0;
	wire w_dff_A_0iaZKLE90_0;
	wire w_dff_A_o39kVAQT8_0;
	wire w_dff_A_BtRLGDEP0_0;
	wire w_dff_A_99i7LAPF7_0;
	wire w_dff_A_57O3sZWL4_0;
	wire w_dff_A_xlNFVysj3_0;
	wire w_dff_A_XrLXivbj2_0;
	wire w_dff_A_L6iGirEZ7_0;
	wire w_dff_A_2JxubHvP6_0;
	wire w_dff_A_BZKSH1bR1_0;
	wire w_dff_A_o1MoDGsA2_0;
	wire w_dff_A_MkJoJj2e9_0;
	wire w_dff_A_948uc08y8_0;
	wire w_dff_A_zRXXoYv12_0;
	wire w_dff_A_Z9DbpMDw3_0;
	wire w_dff_A_wFCG80GU4_0;
	wire w_dff_A_aygIYzC69_0;
	wire w_dff_A_xwJ2ZW0q4_0;
	wire w_dff_A_KwXllmL38_0;
	wire w_dff_A_Ebnw4n3T0_0;
	wire w_dff_A_GLVGhJ037_0;
	wire w_dff_A_jcMUFEnB7_0;
	wire w_dff_A_TvHVLmIo4_0;
	wire w_dff_A_SpO2BMhM3_1;
	wire w_dff_A_jCo04NMI5_0;
	wire w_dff_A_47nucgNw2_0;
	wire w_dff_A_kWzdgH5L4_0;
	wire w_dff_A_UqajSPWh9_0;
	wire w_dff_A_JKzZdKFE9_0;
	wire w_dff_A_jJba68X70_0;
	wire w_dff_A_4GlW8KNG1_0;
	wire w_dff_A_uFgZRCcw0_0;
	wire w_dff_A_X5fIxnN13_0;
	wire w_dff_A_UXfhf2CA5_0;
	wire w_dff_A_nRP8m8mD1_0;
	wire w_dff_A_aiFZ5ciw2_0;
	wire w_dff_A_qHkjQACn7_0;
	wire w_dff_A_qjEkwSO13_0;
	wire w_dff_A_s81eWuvH7_0;
	wire w_dff_A_Mw9uFUtC9_0;
	wire w_dff_A_8PszQ2VZ8_0;
	wire w_dff_A_kQXK6ufu9_0;
	wire w_dff_A_03d5zdZt4_0;
	wire w_dff_A_meMuVMTn9_0;
	wire w_dff_A_4VSEAS7z3_0;
	wire w_dff_A_OhWZ7Kp21_0;
	wire w_dff_A_L5bNWsc53_0;
	wire w_dff_A_OtBO3pev2_0;
	wire w_dff_A_abVhkHvY7_1;
	wire w_dff_A_V85JZFxw4_0;
	wire w_dff_A_d3Gpi8Jc0_0;
	wire w_dff_A_jcmEfclu4_0;
	wire w_dff_A_Yb6Nbclj0_0;
	wire w_dff_A_R1AK6bSL6_0;
	wire w_dff_A_R8FvGvkB6_0;
	wire w_dff_A_kcFAIxA96_0;
	wire w_dff_A_qZIX0z0i8_0;
	wire w_dff_A_famX9DUw0_0;
	wire w_dff_A_gNC84Z308_0;
	wire w_dff_A_ofIv66Zj4_0;
	wire w_dff_A_w6uY1qWn7_0;
	wire w_dff_A_6LpPMPaN4_0;
	wire w_dff_A_xEfkJmnA8_0;
	wire w_dff_A_8G9h2CEO0_0;
	wire w_dff_A_XKpVDc3B3_0;
	wire w_dff_A_ebKE19mp1_0;
	wire w_dff_A_lBxUdizI1_0;
	wire w_dff_A_XRZtbF221_0;
	wire w_dff_A_FUWpOhri7_0;
	wire w_dff_A_eOzo2qa53_0;
	wire w_dff_A_jznu23Zk0_0;
	wire w_dff_A_9YXdI7EP2_0;
	wire w_dff_A_ML9mQqH98_0;
	wire w_dff_A_qpWbjoOy4_1;
	wire w_dff_A_oaFPvoaF5_0;
	wire w_dff_A_TrKS8yWm2_0;
	wire w_dff_A_E4VJRHTl3_0;
	wire w_dff_A_mXSY4zYP5_0;
	wire w_dff_A_w9A5TP2H2_0;
	wire w_dff_A_VlZUHRa21_0;
	wire w_dff_A_IvtZ7P7g1_0;
	wire w_dff_A_BfS3k26j9_0;
	wire w_dff_A_JOfFvtra7_0;
	wire w_dff_A_KvfZLhqi5_0;
	wire w_dff_A_9y1c4S6c9_0;
	wire w_dff_A_ZojNuHXZ5_0;
	wire w_dff_A_xpH9CXJM5_0;
	wire w_dff_A_fKaLlKz50_0;
	wire w_dff_A_6MgvSZpQ6_0;
	wire w_dff_A_AqsUbGqI2_0;
	wire w_dff_A_sHrKWhtn6_0;
	wire w_dff_A_k4QmlshR7_0;
	wire w_dff_A_ptLqqP2h2_0;
	wire w_dff_A_TiUNK2D95_0;
	wire w_dff_A_uKi4mG2o3_0;
	wire w_dff_A_EstgPHQC2_0;
	wire w_dff_A_TkpcScS52_0;
	wire w_dff_A_wsNhdpVO8_0;
	wire w_dff_A_lD6XExhc7_1;
	wire w_dff_A_Jl4ZNpnA1_0;
	wire w_dff_A_YRcS2ikS6_0;
	wire w_dff_A_c9n10fjS4_0;
	wire w_dff_A_QTjUCbq50_0;
	wire w_dff_A_XMibHe3f4_0;
	wire w_dff_A_Hgy08DiC8_0;
	wire w_dff_A_ty6mWJ6Y6_0;
	wire w_dff_A_NcpEUnwM2_0;
	wire w_dff_A_zHy5uA2U5_0;
	wire w_dff_A_k6LFJOLP7_0;
	wire w_dff_A_GQGhDm5G4_0;
	wire w_dff_A_iiw7dC0S9_0;
	wire w_dff_A_pGv4YvHQ3_0;
	wire w_dff_A_ReWdVeme4_0;
	wire w_dff_A_IDiLCvME8_0;
	wire w_dff_A_ATyGnFjX3_0;
	wire w_dff_A_FsvZQZ7i2_0;
	wire w_dff_A_RsX6UkSY0_0;
	wire w_dff_A_EsQzUZc85_0;
	wire w_dff_A_brVQAggx3_0;
	wire w_dff_A_cwqWPGr07_0;
	wire w_dff_A_dVrG7hGV7_0;
	wire w_dff_A_FrYoED5t0_0;
	wire w_dff_A_TpleHrMc4_0;
	wire w_dff_A_4e4EIA5N1_1;
	wire w_dff_A_NNj3eLVc1_0;
	wire w_dff_A_3HlQ2bnD6_0;
	wire w_dff_A_K0APsira4_0;
	wire w_dff_A_5mirhI067_0;
	wire w_dff_A_SgChimeS9_0;
	wire w_dff_A_I7tJAHJo4_0;
	wire w_dff_A_jEORaBQ79_0;
	wire w_dff_A_981HW88k6_0;
	wire w_dff_A_rAG8wnC35_0;
	wire w_dff_A_yEMSOdVg2_0;
	wire w_dff_A_7H2nFOht3_0;
	wire w_dff_A_0fRBeq0C1_0;
	wire w_dff_A_8X4qeEpt1_0;
	wire w_dff_A_ja6OvJz09_0;
	wire w_dff_A_FpJLk7TL0_0;
	wire w_dff_A_LzWbjckA9_0;
	wire w_dff_A_s9R8RfWi8_0;
	wire w_dff_A_pqgIY3NN1_0;
	wire w_dff_A_26dtetRk3_0;
	wire w_dff_A_h3Zg1kjR9_0;
	wire w_dff_A_EtvJhjP99_0;
	wire w_dff_A_yiqcB09d7_0;
	wire w_dff_A_iCRYLmRz2_0;
	wire w_dff_A_Uhx4mFUf4_0;
	wire w_dff_A_5DKWnxSc5_2;
	wire w_dff_A_xVQWH6Tr1_0;
	wire w_dff_A_uI2A11gr1_0;
	wire w_dff_A_xr7y9Smy1_0;
	wire w_dff_A_E4DmUa6Y8_0;
	wire w_dff_A_KCPLWmcP4_0;
	wire w_dff_A_6WVWdltR0_0;
	wire w_dff_A_ahA86vOb6_0;
	wire w_dff_A_6KcVJOQL8_0;
	wire w_dff_A_oIjlbJoV5_0;
	wire w_dff_A_x57fBEvW9_0;
	wire w_dff_A_YwmGE3Am3_0;
	wire w_dff_A_pd1p2vGz2_0;
	wire w_dff_A_nKTgTCH18_0;
	wire w_dff_A_QP5hFykY0_0;
	wire w_dff_A_WeoXHbwr4_0;
	wire w_dff_A_Ydk4Ner15_0;
	wire w_dff_A_uI1fL5E10_0;
	wire w_dff_A_NhiN46YI3_0;
	wire w_dff_A_BvVZYSyB5_0;
	wire w_dff_A_CPpuDR8l0_0;
	wire w_dff_A_2AJPeBJv2_0;
	wire w_dff_A_CXKw5YL30_2;
	wire w_dff_A_sN8DakQO6_0;
	wire w_dff_A_JcOoUIoU0_0;
	wire w_dff_A_AMQ9nWoi5_0;
	wire w_dff_A_ffv8D3iP0_0;
	wire w_dff_A_NLkBdWcm3_0;
	wire w_dff_A_rkUBQDy35_0;
	wire w_dff_A_gYFtotOP3_0;
	wire w_dff_A_WHcSynkR0_0;
	wire w_dff_A_lBDItlpU6_0;
	wire w_dff_A_07oRUG598_0;
	wire w_dff_A_luXZfeUs5_0;
	wire w_dff_A_zVtXFOHs9_0;
	wire w_dff_A_WGsCsiRH9_0;
	wire w_dff_A_NweTt4l64_0;
	wire w_dff_A_if2qgv0H6_0;
	wire w_dff_A_wAsJxjbj2_0;
	wire w_dff_A_9xIy5x3z4_0;
	wire w_dff_A_6JOjYtxb7_0;
	wire w_dff_A_cRKkT0PC0_0;
	wire w_dff_A_aItKAicj2_0;
	wire w_dff_A_wTQCLBXD0_0;
	wire w_dff_A_TR3QSKJ91_2;
	wire w_dff_A_RkLtvXpE6_0;
	wire w_dff_A_z0TMj8TG3_0;
	wire w_dff_A_64wFIkQ95_0;
	wire w_dff_A_puWSMKTF7_0;
	wire w_dff_A_dk9tfpKv2_0;
	wire w_dff_A_8tTZc8Kw2_0;
	wire w_dff_A_Xevm6M2H3_0;
	wire w_dff_A_FyPeZUxw6_0;
	wire w_dff_A_9aTbQNIu4_0;
	wire w_dff_A_nzxuVn7x7_0;
	wire w_dff_A_gLUPRY4w4_0;
	wire w_dff_A_PBKA6CSE2_0;
	wire w_dff_A_40L5QOHL3_0;
	wire w_dff_A_VDZx6CGd6_0;
	wire w_dff_A_wr4CqXl23_0;
	wire w_dff_A_TjeCiBd20_0;
	wire w_dff_A_jh06xNKB8_0;
	wire w_dff_A_xpbmMFm96_0;
	wire w_dff_A_3X92xAxM1_0;
	wire w_dff_A_3aVTff5Z7_0;
	wire w_dff_A_wISkywuW2_0;
	wire w_dff_A_9yC0VVfO7_2;
	wire w_dff_A_jFXPlW4o6_0;
	wire w_dff_A_xJpXaXBX8_0;
	wire w_dff_A_5kSP9aBD0_0;
	wire w_dff_A_zNTpmbIP0_0;
	wire w_dff_A_a2AJYJZY2_0;
	wire w_dff_A_S7QEW4ah1_0;
	wire w_dff_A_9NJzThi50_0;
	wire w_dff_A_ilQaAq009_0;
	wire w_dff_A_I6OnOS4L9_0;
	wire w_dff_A_Kqfm5GjQ8_0;
	wire w_dff_A_DQQxTDK83_0;
	wire w_dff_A_2z7dsrkQ1_0;
	wire w_dff_A_7xiub2BF7_0;
	wire w_dff_A_pj51po7o9_0;
	wire w_dff_A_jekEyZBi1_0;
	wire w_dff_A_1mn3SqOD2_0;
	wire w_dff_A_A90jU8Hx4_0;
	wire w_dff_A_NS9tbqK98_0;
	wire w_dff_A_TGZ9z4nW7_0;
	wire w_dff_A_ymbLtiM65_0;
	wire w_dff_A_D3s1irdO4_0;
	wire w_dff_A_lQWDjGuG1_0;
	wire w_dff_A_rizW0C430_2;
	wire w_dff_A_KgAAbwuH8_0;
	wire w_dff_A_7nnuyk1Q2_0;
	wire w_dff_A_vYgPw98P2_0;
	wire w_dff_A_GiHiMhTQ7_0;
	wire w_dff_A_AUqkSgAN4_0;
	wire w_dff_A_aDDEqaYT7_0;
	wire w_dff_A_wChBvq3p6_0;
	wire w_dff_A_vJm1Pm654_0;
	wire w_dff_A_MQroQ7IC1_0;
	wire w_dff_A_GiyvZx260_0;
	wire w_dff_A_jcrhMJgS8_0;
	wire w_dff_A_gs4gCJG75_0;
	wire w_dff_A_43PrkEhK8_0;
	wire w_dff_A_blgBBLO64_0;
	wire w_dff_A_Mn3y9pAO6_0;
	wire w_dff_A_OmwUq7pT7_0;
	wire w_dff_A_wTIzYJdY3_0;
	wire w_dff_A_X6fMt0Zj0_0;
	wire w_dff_A_kU02qcPQ1_0;
	wire w_dff_A_adtuXUxE0_0;
	wire w_dff_A_elugQIR87_2;
	wire w_dff_A_vjOvb3W06_0;
	wire w_dff_A_f7oJb32k4_0;
	wire w_dff_A_cGLVsDBl2_0;
	wire w_dff_A_LAicCfTh9_0;
	wire w_dff_A_zPpsueOZ2_0;
	wire w_dff_A_ncAURSH36_0;
	wire w_dff_A_kCSS4AZq0_0;
	wire w_dff_A_NYHD2jE67_0;
	wire w_dff_A_oYi4of0D3_0;
	wire w_dff_A_Hb4ytExg0_0;
	wire w_dff_A_mhiIvyDJ5_0;
	wire w_dff_A_GMirbeNl4_0;
	wire w_dff_A_6PHqUvff5_0;
	wire w_dff_A_NhBUSYdt2_0;
	wire w_dff_A_njyrBR860_0;
	wire w_dff_A_0fI8E1tn5_0;
	wire w_dff_A_LjAQVpdm0_0;
	wire w_dff_A_hOjv7GI27_0;
	wire w_dff_A_fvRySZuu8_0;
	wire w_dff_A_FrydKVP70_0;
	wire w_dff_A_FaokHENP3_2;
	wire w_dff_A_0QcR0jCY9_0;
	wire w_dff_A_fkXPbOey1_0;
	wire w_dff_A_FBlijyyz1_0;
	wire w_dff_A_oaAOkGXK3_0;
	wire w_dff_A_K7S56rVT4_0;
	wire w_dff_A_KCQuRw3E0_0;
	wire w_dff_A_fgZNn9MB6_0;
	wire w_dff_A_TbSvztVd9_0;
	wire w_dff_A_S7lPsxhh1_0;
	wire w_dff_A_xOKC3ko35_0;
	wire w_dff_A_d3Ip3zeE9_0;
	wire w_dff_A_64YrB5C19_0;
	wire w_dff_A_iSOwSdHN7_0;
	wire w_dff_A_n29ScSW67_0;
	wire w_dff_A_xQwsdKbI5_0;
	wire w_dff_A_XqEADTOL7_0;
	wire w_dff_A_QXQ2Bv1S2_0;
	wire w_dff_A_ao6Jk5qP6_0;
	wire w_dff_A_xTYZkzUF4_0;
	wire w_dff_A_K4tG1aVx5_0;
	wire w_dff_A_xsbWQ4I27_2;
	wire w_dff_A_ZmxnlbO75_0;
	wire w_dff_A_pGGRNlkO6_0;
	wire w_dff_A_vT2fL17A8_0;
	wire w_dff_A_HyQ7vQWy2_0;
	wire w_dff_A_gUlXqVgu7_0;
	wire w_dff_A_mFipyJM54_0;
	wire w_dff_A_vnhY7zrE0_0;
	wire w_dff_A_zvh8j5m56_0;
	wire w_dff_A_NX87CFfs2_0;
	wire w_dff_A_bMeo0Xii2_0;
	wire w_dff_A_0gDixBLJ5_0;
	wire w_dff_A_ShcqrH7E4_0;
	wire w_dff_A_uXKUj2lM3_0;
	wire w_dff_A_ayzisLxe1_0;
	wire w_dff_A_B7C4cCNj4_0;
	wire w_dff_A_VyHL6giX3_0;
	wire w_dff_A_p7En6qza1_0;
	wire w_dff_A_wlaTIjaE6_0;
	wire w_dff_A_ASPWIk2T1_0;
	wire w_dff_A_6SUGHeB62_0;
	wire w_dff_A_BEb53Iaq1_2;
	wire w_dff_A_oloWKfMa0_0;
	wire w_dff_A_pqD3GZ3g8_0;
	wire w_dff_A_EYGuIKep0_0;
	wire w_dff_A_9LMeRw9x6_0;
	wire w_dff_A_deNX8pML9_0;
	wire w_dff_A_MxDtdVQe0_0;
	wire w_dff_A_nl4mcWAu4_0;
	wire w_dff_A_ewEv8Ybp9_0;
	wire w_dff_A_U6aBBlE37_0;
	wire w_dff_A_sgeIN7sc3_0;
	wire w_dff_A_P1ICeaaJ8_0;
	wire w_dff_A_QA7VTbku3_0;
	wire w_dff_A_sgG74Gx40_0;
	wire w_dff_A_CUgQ3iz31_0;
	wire w_dff_A_aJMDk6zR2_0;
	wire w_dff_A_SUtsIFMm6_0;
	wire w_dff_A_j4efVi3O6_2;
	wire w_dff_A_Yq0pu1wW0_0;
	wire w_dff_A_GOBiuBFn1_0;
	wire w_dff_A_WbbPGbyL9_0;
	wire w_dff_A_QUDDyT3N6_0;
	wire w_dff_A_SRlVGceg3_0;
	wire w_dff_A_uALdLlXS3_0;
	wire w_dff_A_5DWrPsbL7_0;
	wire w_dff_A_TJ8wjj571_0;
	wire w_dff_A_g4gbUWNR7_0;
	wire w_dff_A_awoE7okF8_0;
	wire w_dff_A_lUxuw5nY6_0;
	wire w_dff_A_HON1Q2SL5_0;
	wire w_dff_A_VA68RU7z1_0;
	wire w_dff_A_iT40JmC66_0;
	wire w_dff_A_U5oLsT2f1_0;
	wire w_dff_A_I4bktKWu6_0;
	wire w_dff_A_4Xgg3Wdu6_2;
	wire w_dff_A_1M4z8uvC6_0;
	wire w_dff_A_5FiHU8d02_0;
	wire w_dff_A_tjm3Ww215_0;
	wire w_dff_A_71ej5SFX2_0;
	wire w_dff_A_TkQReInG0_0;
	wire w_dff_A_3Nz5jTUP4_0;
	wire w_dff_A_GuaHMZHy1_0;
	wire w_dff_A_G3Nt3byh6_0;
	wire w_dff_A_CJkqSmBs2_0;
	wire w_dff_A_MN2Ias6m6_0;
	wire w_dff_A_aWeCwI952_0;
	wire w_dff_A_KD0XfKV14_0;
	wire w_dff_A_IiaX7pO55_0;
	wire w_dff_A_LnHzd7tf5_0;
	wire w_dff_A_n3GGxwow0_2;
	wire w_dff_A_BC4hp5hS2_0;
	wire w_dff_A_8Tk9dvqi4_0;
	wire w_dff_A_35g2JW3m8_0;
	wire w_dff_A_HCgQiUjK2_0;
	wire w_dff_A_wzBljx7g8_0;
	wire w_dff_A_t0eXidmG0_0;
	wire w_dff_A_Vz2gVHAS2_0;
	wire w_dff_A_igQvbAAg2_0;
	wire w_dff_A_dNQgYKEB7_0;
	wire w_dff_A_HZi5PSZl0_0;
	wire w_dff_A_Y3j9diA04_0;
	wire w_dff_A_tSL6M70X7_0;
	wire w_dff_A_KL55QyXJ1_0;
	wire w_dff_A_Svx5lZzP2_0;
	wire w_dff_A_58pnp1Fr3_0;
	wire w_dff_A_Qysn4twB7_0;
	wire w_dff_A_QmKqJRIv2_2;
	wire w_dff_A_qkdo91Fi2_0;
	wire w_dff_A_OGCZ5huo7_0;
	wire w_dff_A_5UvpBk0r5_0;
	wire w_dff_A_x0JF5A1q7_0;
	wire w_dff_A_QL1opl1b8_0;
	wire w_dff_A_3OlaC27m3_0;
	wire w_dff_A_vVvcsjH78_0;
	wire w_dff_A_6eBH2sMQ8_0;
	wire w_dff_A_0fdM7YKm5_0;
	wire w_dff_A_iDGcRBmp4_0;
	wire w_dff_A_jEyBLj9Q6_0;
	wire w_dff_A_pU8QpZRt2_0;
	wire w_dff_A_yW1sngvI9_0;
	wire w_dff_A_j1vu3Yto4_0;
	wire w_dff_A_zMkrSvUF8_0;
	wire w_dff_A_silvTFXx7_0;
	wire w_dff_A_t4OEWpbI4_2;
	wire w_dff_A_XSGwYZJ66_0;
	wire w_dff_A_qKUKWfzu2_0;
	wire w_dff_A_qxukhu7v4_0;
	wire w_dff_A_qBLwA6M94_0;
	wire w_dff_A_JG0L87Ww6_0;
	wire w_dff_A_2E0x3VZI3_0;
	wire w_dff_A_fuXWis3a2_0;
	wire w_dff_A_0ReWyaKS8_0;
	wire w_dff_A_fKGZCOfD7_0;
	wire w_dff_A_PF4yy7YQ5_0;
	wire w_dff_A_EPhcu3l71_0;
	wire w_dff_A_84XnLP5F1_0;
	wire w_dff_A_DW0i6k8X9_0;
	wire w_dff_A_Vto4TfUX5_0;
	wire w_dff_A_8MThqmXy2_1;
	wire w_dff_A_DifVr3Om1_0;
	wire w_dff_A_Ng0oECXB3_0;
	wire w_dff_A_l0AW4AGy0_0;
	wire w_dff_A_mmWYF7Z63_0;
	wire w_dff_A_G1z6TzYy4_0;
	wire w_dff_A_z7M6r6dH6_0;
	wire w_dff_A_ttc7DjDN3_0;
	wire w_dff_A_njPV4DTd3_0;
	wire w_dff_A_JqmkJdmq5_0;
	wire w_dff_A_2tof4Dml2_0;
	wire w_dff_A_QK0QUSLo3_0;
	wire w_dff_A_W8pZpPQW0_0;
	wire w_dff_A_hwvb23Lb6_0;
	wire w_dff_A_7ZzzLzVy7_0;
	wire w_dff_A_Y9LsZRIZ3_0;
	wire w_dff_A_R3Bi5i7L2_0;
	wire w_dff_A_dJA0b8xC9_0;
	wire w_dff_A_Ez533ZU05_0;
	wire w_dff_A_yP86I3PT5_0;
	wire w_dff_A_pheM8mO71_0;
	wire w_dff_A_FM7ga7ou8_1;
	wire w_dff_A_liYurLTQ9_0;
	wire w_dff_A_n80DzAQ95_0;
	wire w_dff_A_TkSX4e669_0;
	wire w_dff_A_V1PAS0K72_0;
	wire w_dff_A_86hg12ZQ9_0;
	wire w_dff_A_zseMmEC93_0;
	wire w_dff_A_bYF9qzDW2_0;
	wire w_dff_A_ZRANlNYg9_0;
	wire w_dff_A_IK7n4Vwj6_0;
	wire w_dff_A_ttrUmXIN0_0;
	wire w_dff_A_UkrFsFir7_0;
	wire w_dff_A_NHS2pa075_0;
	wire w_dff_A_dxCAVoLL3_0;
	wire w_dff_A_Q1qsc3s55_0;
	wire w_dff_A_4e1Us7Ku2_0;
	wire w_dff_A_hfWDkREK5_0;
	wire w_dff_A_iqOjJnuo3_0;
	wire w_dff_A_ntWxwqQK1_0;
	wire w_dff_A_2xFGmuuI8_0;
	wire w_dff_A_JRAIqznC6_0;
	wire w_dff_A_x5Bdeqtt8_2;
	wire w_dff_A_hPhp5Y865_0;
	wire w_dff_A_b14ek91s8_0;
	wire w_dff_A_ZfCVIXFP5_0;
	wire w_dff_A_zGLOD5nD8_0;
	wire w_dff_A_ANbg6Wwm2_0;
	wire w_dff_A_rG5dGwXV3_0;
	wire w_dff_A_yI5iJGLK9_0;
	wire w_dff_A_g6nfOlMj9_0;
	wire w_dff_A_DemqSCnw7_0;
	wire w_dff_A_VCVhWC6d6_0;
	wire w_dff_A_7iGFQniU7_0;
	wire w_dff_A_dUvFZuI17_2;
	wire w_dff_A_XDTo9of91_0;
	wire w_dff_A_k3CyBxZC2_0;
	wire w_dff_A_n1DUMr9q9_0;
	wire w_dff_A_1TzUogFk7_0;
	wire w_dff_A_1lDnUSeg9_0;
	wire w_dff_A_mGNG4H3s8_0;
	wire w_dff_A_Y6F9dhiL1_0;
	wire w_dff_A_3Br8LzRX7_0;
	wire w_dff_A_g7JJJbif9_0;
	wire w_dff_A_9YmxPRjd2_0;
	wire w_dff_A_dVFojz512_0;
	wire w_dff_A_KD56kTfy9_2;
	wire w_dff_A_d4narGFS4_0;
	wire w_dff_A_R5rS28be5_0;
	wire w_dff_A_a4yXc90U1_0;
	wire w_dff_A_x4bT6BTj0_0;
	wire w_dff_A_XVnWRPNy5_0;
	wire w_dff_A_8vHnto142_0;
	wire w_dff_A_NkyevxkC1_0;
	wire w_dff_A_i7NRLqUr7_0;
	wire w_dff_A_PkvviMUt2_0;
	wire w_dff_A_YmyiEMt48_0;
	wire w_dff_A_YsqjyaXh4_0;
	wire w_dff_A_Cy9lkNbV7_2;
	wire w_dff_A_NhrnOveV2_0;
	wire w_dff_A_7Yvj5zxD4_0;
	wire w_dff_A_X3xuNiyw9_0;
	wire w_dff_A_Qvyp2K459_0;
	wire w_dff_A_c7vrLhPU0_0;
	wire w_dff_A_sUSzQodi5_0;
	wire w_dff_A_uPhWfkZE8_0;
	wire w_dff_A_2NiPPrNn4_0;
	wire w_dff_A_XryDxHHc7_0;
	wire w_dff_A_b0E8rjz12_0;
	wire w_dff_A_cZ9PTVaY6_0;
	wire w_dff_A_snZJi9ST6_1;
	wire w_dff_A_aq8I2DKO3_0;
	wire w_dff_A_7cy1O96o3_0;
	wire w_dff_A_IOaltbKl6_0;
	wire w_dff_A_EMmGKFik4_0;
	wire w_dff_A_nz9wzjG16_0;
	wire w_dff_A_X8V0nYfi7_0;
	wire w_dff_A_TajhmYGg3_0;
	wire w_dff_A_Y0a6UnnT6_0;
	wire w_dff_A_ao25x0TM2_0;
	wire w_dff_A_yASrjxQ85_0;
	wire w_dff_A_7qI3Ea5C9_0;
	wire w_dff_A_9tdBiNxn1_0;
	wire w_dff_A_4pz3WHHu2_0;
	wire w_dff_A_q7fYNNpk5_0;
	wire w_dff_A_VFHKjjf15_0;
	wire w_dff_A_iRbCYIBv5_0;
	wire w_dff_A_NoqhdNf00_0;
	wire w_dff_A_DEjCMjYR1_0;
	wire w_dff_A_NU9RSijT7_1;
	wire w_dff_A_Ep3zLD1i4_0;
	wire w_dff_A_Ybo5zWwy2_0;
	wire w_dff_A_isKRucTK0_0;
	wire w_dff_A_QAWQtNTc2_0;
	wire w_dff_A_Uw61XWbZ4_0;
	wire w_dff_A_2OaVpKAG8_0;
	wire w_dff_A_E8YSR3hE2_0;
	wire w_dff_A_1vQVqcdV0_0;
	wire w_dff_A_E420atvZ0_0;
	wire w_dff_A_lO8HBcVh6_0;
	wire w_dff_A_CC1DrSrT2_0;
	wire w_dff_A_kkH6UtBj1_0;
	wire w_dff_A_vOZGE8vc3_0;
	wire w_dff_A_lqf1ogiV1_0;
	wire w_dff_A_k1dgeqFz8_0;
	wire w_dff_A_0NMOQF9m1_0;
	wire w_dff_A_wVNaNbx41_0;
	wire w_dff_A_ZXolT0V26_1;
	wire w_dff_A_ZZq4kYo64_0;
	wire w_dff_A_kldSVPQ84_0;
	wire w_dff_A_kqFFAjy18_0;
	wire w_dff_A_df8MVVbc5_0;
	wire w_dff_A_gjHY7BFg2_0;
	wire w_dff_A_N1YpechW1_0;
	wire w_dff_A_Xs2t9kTr4_0;
	wire w_dff_A_JN19R1lq1_0;
	wire w_dff_A_v9VaeYR98_0;
	wire w_dff_A_2WGcBnbR7_0;
	wire w_dff_A_ipFZ34Lt1_0;
	wire w_dff_A_iTZPwjIH7_0;
	wire w_dff_A_kXYckNTh4_0;
	wire w_dff_A_gww8E7655_0;
	wire w_dff_A_oOE0Yfsj3_0;
	wire w_dff_A_ya5AUVCw8_0;
	wire w_dff_A_hTLAoxsz8_0;
	wire w_dff_A_ThmdqykU8_1;
	wire w_dff_A_dh5p1ikk2_0;
	wire w_dff_A_pEqBSy1B5_0;
	wire w_dff_A_vGTJbVse1_0;
	wire w_dff_A_MhaL0zvK2_0;
	wire w_dff_A_3tpwft3G5_0;
	wire w_dff_A_VkYGSsx51_0;
	wire w_dff_A_ZHMTSP3i6_2;
	wire w_dff_A_V4EC7Dd53_0;
	wire w_dff_A_aYgdNbkN9_0;
	wire w_dff_A_UNBiD9eu9_0;
	wire w_dff_A_9oNu4w210_0;
	wire w_dff_A_h3ZyZ3hk0_0;
	wire w_dff_A_umIRhdYr8_0;
	wire w_dff_A_cKv4AR9w0_0;
	wire w_dff_A_jMxXD8LX8_0;
	wire w_dff_A_7d04FC6Z1_0;
	wire w_dff_A_CQB6sj5B2_0;
	wire w_dff_A_VvWL19su1_0;
	wire w_dff_A_UOiucRSY6_0;
	wire w_dff_A_br8hVELs5_0;
	wire w_dff_A_IbBxoM2o5_0;
	wire w_dff_A_wR17c80c2_1;
	wire w_dff_A_XfJEjMF64_0;
	wire w_dff_A_og1H0ZN97_0;
	wire w_dff_A_SM2wA2Wy3_0;
	wire w_dff_A_MUGDUylO6_0;
	wire w_dff_A_bBuWOqqy7_0;
	wire w_dff_A_c2vFd4CO8_0;
	wire w_dff_A_PSykAM4I7_0;
	wire w_dff_A_bkq4kN653_0;
	wire w_dff_A_rB5l1Dxt4_0;
	wire w_dff_A_7WDLAm422_0;
	wire w_dff_A_FdOzntpk3_0;
	wire w_dff_A_5Xx6TgKH7_1;
	wire w_dff_A_lMOqQ0rS8_0;
	wire w_dff_A_t7z3xsnm6_0;
	wire w_dff_A_OetBEDxM9_0;
	wire w_dff_A_icOXVjl64_0;
	wire w_dff_A_shiYJbDp9_0;
	wire w_dff_A_rAXf54PX9_0;
	wire w_dff_A_Jg4vQ9HV2_0;
	wire w_dff_A_WcamD9mg6_0;
	wire w_dff_A_JuZhTEyw5_0;
	wire w_dff_A_goRRc3wp5_0;
	wire w_dff_A_DDmMEMTW2_0;
	wire w_dff_A_8MZY8CUr4_0;
	wire w_dff_A_AA3ph8CU2_0;
	wire w_dff_A_qqGvtkqc6_1;
	wire w_dff_A_qGoG3T8h0_0;
	wire w_dff_A_Ii5ZwzAM5_0;
	wire w_dff_A_ybg4YFsM6_0;
	wire w_dff_A_PWBe3cmi9_0;
	wire w_dff_A_9jv2sYF36_0;
	wire w_dff_A_18j6Fyyx0_0;
	wire w_dff_A_389TtBxd9_0;
	wire w_dff_A_2IXg8DsH0_0;
	wire w_dff_A_oXW4n89S0_0;
	wire w_dff_A_LqJlf77v3_0;
	wire w_dff_A_SBVJSIm32_0;
	wire w_dff_A_0ulM0GLY8_0;
	wire w_dff_A_jPf8QPi70_0;
	wire w_dff_A_NzPM8eWl4_0;
	wire w_dff_A_r7DH87ma9_0;
	wire w_dff_A_7O2wzkaw1_2;
	wire w_dff_A_ilQmmqJD0_0;
	wire w_dff_A_IYtFxu9W0_0;
	wire w_dff_A_e2k2DRdl7_0;
	wire w_dff_A_WeGYUlUa8_0;
	wire w_dff_A_cr3jm7j96_0;
	wire w_dff_A_WFMfEKIz5_0;
	wire w_dff_A_6Etd3qUY3_0;
	wire w_dff_A_BHu1VUKb9_0;
	wire w_dff_A_yykVMFx44_0;
	wire w_dff_A_rarOqqIw2_0;
	wire w_dff_A_h2U5pKVg1_0;
	wire w_dff_A_pbVMcsM92_0;
	wire w_dff_A_MuzgbhDl3_0;
	wire w_dff_A_1jIKfZT23_0;
	wire w_dff_A_N7LHGUu06_1;
	wire w_dff_A_Uqa9WElK9_0;
	wire w_dff_A_drEy0vdf7_0;
	wire w_dff_A_vCOILdJZ5_0;
	wire w_dff_A_RV1WwCaw6_0;
	wire w_dff_A_ISZ4NYmR7_0;
	wire w_dff_A_Hpj30Ax63_0;
	wire w_dff_A_mFOiPj4c2_0;
	wire w_dff_A_ppkBLltQ7_0;
	wire w_dff_A_dPMgjU3R7_0;
	wire w_dff_A_Z21vggDg8_1;
	wire w_dff_A_c64wwYKJ4_0;
	wire w_dff_A_ypNE6hvh7_0;
	wire w_dff_A_CvZYO3aI0_0;
	wire w_dff_A_g94nGanx7_0;
	wire w_dff_A_p1vJkx1M8_0;
	wire w_dff_A_A7pY0dpX1_0;
	wire w_dff_A_hYyeh1fV6_0;
	wire w_dff_A_ZAVSQPGH8_0;
	wire w_dff_A_p11MuTuQ9_0;
	wire w_dff_A_PZOjwCQ04_0;
	wire w_dff_A_hq6ePeyd7_0;
	wire w_dff_A_5zsUPBA47_1;
	wire w_dff_A_VYoBtlWz3_0;
	wire w_dff_A_RkhlHoH04_0;
	wire w_dff_A_m9DOy8Tk0_0;
	wire w_dff_A_U50f7xEO2_0;
	wire w_dff_A_pgJa7A665_0;
	wire w_dff_A_93DO8Yf21_0;
	wire w_dff_A_jwa96Fl75_0;
	wire w_dff_A_HnAfBtkG4_0;
	wire w_dff_A_Fulb2dLV5_0;
	wire w_dff_A_Zp2sodSg8_0;
	wire w_dff_A_6hDRUkCX4_0;
	wire w_dff_A_Q01r9AYR6_0;
	wire w_dff_A_M2r8JevI0_1;
	wire w_dff_A_4NKiSx5A2_0;
	wire w_dff_A_VWi6s1Jw2_0;
	wire w_dff_A_podGFzGD8_0;
	wire w_dff_A_dBpxepUG6_0;
	wire w_dff_A_k5ZtWuAc5_0;
	wire w_dff_A_ODIXZ89F6_0;
	wire w_dff_A_JAenVpx02_0;
	wire w_dff_A_IHvtxObP5_0;
	wire w_dff_A_bMf3h5LL5_0;
	wire w_dff_A_b4ooQjrS2_0;
	wire w_dff_A_gUT7qUu26_0;
	wire w_dff_A_ufoCXX3U0_0;
	wire w_dff_A_3QUBX8Qt3_0;
	wire w_dff_A_rsHUFwPC0_1;
	wire w_dff_A_T9asdqcq4_0;
	wire w_dff_A_ixcoWCSO2_0;
	wire w_dff_A_PtOWfpMy2_0;
	wire w_dff_A_DBRdP60S9_0;
	wire w_dff_A_Yc6tf6mU9_0;
	wire w_dff_A_tMCRbGHo2_0;
	wire w_dff_A_rz5qe9ya3_0;
	wire w_dff_A_x6hpU3qV9_0;
	wire w_dff_A_CAcrCyCy6_0;
	wire w_dff_A_UlofxvGN3_0;
	wire w_dff_A_MB8Gfrb67_0;
	wire w_dff_A_TmORDFHX5_0;
	wire w_dff_A_3d3sMt6m5_0;
	wire w_dff_A_PUJJon1W6_0;
	wire w_dff_A_Gz5Kq3nn1_0;
	wire w_dff_A_xJCTIBfG9_0;
	wire w_dff_A_vxWk0kuz4_1;
	wire w_dff_A_lol7tGyc9_0;
	wire w_dff_A_iKEkTV5t6_0;
	wire w_dff_A_o0iOlF0S9_0;
	wire w_dff_A_txTUDvuk0_0;
	wire w_dff_A_gpSSDnqP8_0;
	wire w_dff_A_gKKBMyGH2_0;
	wire w_dff_A_ujXf7ey06_0;
	wire w_dff_A_qdLImWtr9_0;
	wire w_dff_A_a52EhNS14_0;
	wire w_dff_A_C11h4Fyo7_0;
	wire w_dff_A_z4QWg72y8_0;
	wire w_dff_A_18nj1Z018_0;
	wire w_dff_A_P057rDQ20_0;
	wire w_dff_A_lqnMz7y54_0;
	wire w_dff_A_TscTtr5T5_0;
	wire w_dff_A_WFluOpEp0_0;
	wire w_dff_A_v6IyGWyY9_0;
	wire w_dff_A_UkYV04p32_0;
	wire w_dff_A_ZwVSUgu01_2;
	wire w_dff_A_cx4CKnL32_0;
	wire w_dff_A_PlH2NXOH3_0;
	wire w_dff_A_XoYOnOg67_0;
	wire w_dff_A_51s5SvMF4_0;
	wire w_dff_A_aPAHZ5LL4_2;
	wire w_dff_A_1nQkdxS48_0;
	wire w_dff_A_SYXW0W7J6_0;
	wire w_dff_A_JNkxd2Je5_0;
	wire w_dff_A_1sFFBQuW9_0;
	wire w_dff_A_UbtI2DGo5_0;
	wire w_dff_A_G63HbYJb4_0;
	wire w_dff_A_FqGrfaly0_0;
	wire w_dff_A_BjvcmaIf8_2;
	wire w_dff_A_O1uS5i5W7_0;
	wire w_dff_A_Iyon78Eh2_0;
	wire w_dff_A_PSu94Fp34_0;
	wire w_dff_A_FJ6BLk6H5_0;
	wire w_dff_A_t8fnELcm5_0;
	wire w_dff_A_Qy9pUNkj4_0;
	wire w_dff_A_yw6LOFQ46_0;
	wire w_dff_A_wvNU9kS00_0;
	wire w_dff_A_1sDO05d45_0;
	wire w_dff_A_gF1yE8Rg5_0;
	wire w_dff_A_Y8i03vy06_0;
	wire w_dff_A_ONibe0tZ3_0;
	wire w_dff_A_jjXailx57_0;
	wire w_dff_A_T2PMMgd24_2;
	wire w_dff_A_mZ8pUlFz5_0;
	wire w_dff_A_TNXH6GIs1_0;
	wire w_dff_A_1ej4X1Vz2_0;
	wire w_dff_A_KkGM2XdS9_0;
	wire w_dff_A_I4WTF1c89_0;
	wire w_dff_A_8IpmZLyl1_0;
	wire w_dff_A_ncsfzng79_0;
	wire w_dff_A_I7zMWBsM7_0;
	wire w_dff_A_dHBnbEgv2_0;
	wire w_dff_A_7dbf1h419_0;
	wire w_dff_A_fTI4crZ25_0;
	wire w_dff_A_3h2XP5c53_0;
	wire w_dff_A_MjH02BQJ1_0;
	wire w_dff_A_xNgk3bJf2_2;
	wire w_dff_A_W2BFYOlt5_0;
	wire w_dff_A_s48iNXK05_0;
	wire w_dff_A_bKoO846w1_0;
	wire w_dff_A_VhQuBeBX9_0;
	wire w_dff_A_pP2OPXy75_0;
	wire w_dff_A_UcorWion6_0;
	wire w_dff_A_g0IwlMxo1_2;
	wire w_dff_A_lwtRUbdz2_0;
	wire w_dff_A_M8Yz6tkD9_0;
	wire w_dff_A_jeVaUGCm4_0;
	wire w_dff_A_ADLXexMg5_0;
	wire w_dff_A_Ec8wgNHe0_0;
	wire w_dff_A_q1ZP4Ju71_0;
	wire w_dff_A_CWPC1Hao1_0;
	wire w_dff_A_E9glpBty5_0;
	wire w_dff_A_m9mvQOBB9_2;
	wire w_dff_A_ksAJL9kY7_0;
	wire w_dff_A_1Y3wWmRJ0_0;
	wire w_dff_A_aPagkDPs1_0;
	wire w_dff_A_QWdDj9Qn7_0;
	wire w_dff_A_njL2hrF09_0;
	wire w_dff_A_xDSaxUyy4_0;
	wire w_dff_A_ltxeGomy7_0;
	wire w_dff_A_2YYotMmc5_0;
	wire w_dff_A_yHFZUxf10_0;
	wire w_dff_A_V5IgNeJF5_2;
	wire w_dff_A_WpKOQMgU6_0;
	wire w_dff_A_Q4LeZp0o5_0;
	wire w_dff_A_FvOsX6rh2_0;
	wire w_dff_A_7BkNzJCb6_0;
	wire w_dff_A_BJ3sBhf47_0;
	wire w_dff_A_eEZWHRGO0_0;
	wire w_dff_A_bC9aoJ696_0;
	wire w_dff_A_XblsMeDR1_0;
	wire w_dff_A_EuGEL2YL8_0;
	wire w_dff_A_psBQKyDZ2_0;
	wire w_dff_A_cPQHNv5B9_2;
	wire w_dff_A_Ex4eapIB2_0;
	wire w_dff_A_CDNEXem76_0;
	wire w_dff_A_j2MpnEKC7_0;
	wire w_dff_A_ccbMY84v3_0;
	wire w_dff_A_jIVTXgdV8_0;
	wire w_dff_A_HNL4anZJ1_0;
	wire w_dff_A_oRgwlr2S2_2;
	wire w_dff_A_uz6TL8Fv8_0;
	wire w_dff_A_SU6dX10N2_0;
	wire w_dff_A_e658WdM31_0;
	wire w_dff_A_pGhyNCH50_0;
	wire w_dff_A_WJQibS2G0_0;
	wire w_dff_A_HUolGx9D6_0;
	wire w_dff_A_ICfuHqFr6_0;
	wire w_dff_A_P7pf4Vfe9_0;
	wire w_dff_A_7sYsf6TN1_2;
	wire w_dff_A_vNqj2az50_0;
	wire w_dff_A_WyJvKw7E0_0;
	wire w_dff_A_7onYI73d0_0;
	wire w_dff_A_IqxEx9ys7_0;
	wire w_dff_A_XDTDN5YN7_0;
	wire w_dff_A_8xqp0GbX0_0;
	wire w_dff_A_7cTf1T4i3_0;
	wire w_dff_A_AGcDh32s5_0;
	wire w_dff_A_NQrAO3Rv3_0;
	wire w_dff_A_axuI5cBD5_2;
	wire w_dff_A_6qTWw12u7_0;
	wire w_dff_A_nlQVr92Q0_0;
	wire w_dff_A_r8CcTp2v1_0;
	wire w_dff_A_FiW4QVMn3_0;
	wire w_dff_A_1Zb7RLc86_0;
	wire w_dff_A_OUTDsZUk6_0;
	wire w_dff_A_89UOq2Qy0_0;
	wire w_dff_A_l9nTWXBB3_0;
	wire w_dff_A_CYnA1xGP9_0;
	wire w_dff_A_aQZEqZ2H8_0;
	wire w_dff_A_6rpt8BSf5_2;
	wire w_dff_A_z17Rcdpv0_0;
	wire w_dff_A_KyNOtPHU3_0;
	wire w_dff_A_yawDQFw12_0;
	wire w_dff_A_cSrNiilW2_0;
	wire w_dff_A_utYL87sS2_0;
	wire w_dff_A_8re8Z0rV0_2;
	wire w_dff_A_GRR10IgP0_0;
	wire w_dff_A_cJNFi75R8_0;
	wire w_dff_A_ndU0ew5q3_0;
	wire w_dff_A_5tssc9dj5_0;
	wire w_dff_A_6Ux2QBei0_0;
	wire w_dff_A_cW0sIP7H9_0;
	wire w_dff_A_yZQ2yunU8_0;
	wire w_dff_A_inf7Of335_0;
	wire w_dff_A_pTC26Tiz3_0;
	wire w_dff_A_3hWNAct47_2;
	wire w_dff_A_vRwhH48E3_0;
	wire w_dff_A_Cy3dTs2N4_0;
	wire w_dff_A_CdPWBX9T4_0;
	wire w_dff_A_pNUKCvzA0_0;
	wire w_dff_A_yJUKYI1N5_0;
	wire w_dff_A_T2bI25Oj5_0;
	wire w_dff_A_zsBSBdfK1_0;
	wire w_dff_A_NK31XUtu1_0;
	wire w_dff_A_BCHA1aqF8_2;
	wire w_dff_A_4tbiLbgq2_0;
	wire w_dff_A_0rAlDyUm2_0;
	wire w_dff_A_ZpX5zIOT4_0;
	wire w_dff_A_EAuFQQyb3_0;
	wire w_dff_A_F4PkPkyH6_0;
	wire w_dff_A_c9VTKL0p0_0;
	wire w_dff_A_4ZYvl2q66_0;
	wire w_dff_A_Dt6jwWtM8_2;
	wire w_dff_A_X8y2MPUc5_0;
	wire w_dff_A_01xYAUnS3_0;
	wire w_dff_A_HRPcuduB5_0;
	wire w_dff_A_Wbt5YpQd5_0;
	wire w_dff_A_t38XyCSz3_0;
	wire w_dff_A_MqQBwMxU9_2;
	wire w_dff_A_8PyI6sKE1_0;
	wire w_dff_A_KosG7yld5_0;
	wire w_dff_A_Ei7LzMha6_0;
	wire w_dff_A_I4j4iM1L0_0;
	wire w_dff_A_LhURLAYy2_0;
	wire w_dff_A_H303VnPt9_0;
	wire w_dff_A_Pgb2sB8L8_0;
	wire w_dff_A_jOZEJrWW1_0;
	wire w_dff_A_RYqammxv7_0;
	wire w_dff_A_AX6UZEQe8_2;
	wire w_dff_A_JGwoNHNd1_0;
	wire w_dff_A_DLSBcTjB7_0;
	wire w_dff_A_60WASzlJ6_0;
	wire w_dff_A_5DR4MYjN6_0;
	wire w_dff_A_1fEYA2CO0_0;
	wire w_dff_A_VEesDnjg3_0;
	wire w_dff_A_w0wt9ylw3_0;
	wire w_dff_A_74UZtK6D7_0;
	wire w_dff_A_pI4UzbjX7_2;
	wire w_dff_A_PD7GVt7w3_0;
	wire w_dff_A_VIbBDNCn6_0;
	wire w_dff_A_W0P9SmEA4_0;
	wire w_dff_A_Ny37ee9D9_0;
	wire w_dff_A_q0FWV8NW2_0;
	wire w_dff_A_ShpImyfo3_0;
	wire w_dff_A_NbP1wXAe0_0;
	wire w_dff_A_PL0nReCd3_2;
	wire w_dff_A_u6EqJ3Cf5_0;
	wire w_dff_A_irnvtUxB4_0;
	wire w_dff_A_Nmyz9r8A8_0;
	wire w_dff_A_0pY5zyR49_0;
	wire w_dff_A_wjwk8NfH6_2;
	wire w_dff_A_xgw7p0Rd0_0;
	wire w_dff_A_2MfCMQnB8_0;
	wire w_dff_A_osVvMOyj5_0;
	wire w_dff_A_pWQMjWgi5_0;
	wire w_dff_A_MgBElAsh9_0;
	wire w_dff_A_Fc2CDHyE3_0;
	wire w_dff_A_KEmcbVxm3_0;
	wire w_dff_A_r5dLtpmm2_0;
	wire w_dff_A_H9l19U0M7_1;
	wire w_dff_A_sXU9p2Em6_0;
	wire w_dff_A_s63tS9o31_0;
	wire w_dff_A_ll0iwTxF4_0;
	wire w_dff_A_BS2SFMqn9_0;
	wire w_dff_A_G7R4DQMb4_1;
	wire w_dff_A_YL4vOG652_0;
	wire w_dff_A_bDH0qyyM4_0;
	wire w_dff_A_wEHEWSJm2_0;
	wire w_dff_A_SjK7TBBe2_0;
	wire w_dff_A_AR8ckWXU8_0;
	wire w_dff_A_ju0hEPEo9_0;
	wire w_dff_A_5aEQ9g5v0_0;
	wire w_dff_A_Bmlo6mAl5_1;
	wire w_dff_A_U8enSGN17_0;
	wire w_dff_A_AZMS5jDx8_0;
	wire w_dff_A_XlDDOS1I0_0;
	wire w_dff_A_EC7USFKY8_0;
	wire w_dff_A_QdSxRkTV5_0;
	wire w_dff_A_IPO3asO77_0;
	wire w_dff_A_IEdhuDou6_0;
	wire w_dff_A_FIVSn6jT5_1;
	wire w_dff_A_Qi12p23v0_0;
	wire w_dff_A_nTf3kGoq3_0;
	wire w_dff_A_aqjkUbL88_0;
	wire w_dff_A_eJEjRJto9_0;
	wire w_dff_A_hqvWELcf9_0;
	wire w_dff_A_oW4Mql2N5_0;
	wire w_dff_A_CGCd2iDo0_0;
	wire w_dff_A_vkIbfGlh2_0;
	wire w_dff_A_kppvDxAs8_2;
	wire w_dff_A_CJc1MQX59_0;
	wire w_dff_A_NHzDBLZ10_0;
	wire w_dff_A_0kZnrD8X5_0;
	wire w_dff_A_FQcx36GC3_0;
	wire w_dff_A_7HfiSwIN0_0;
	wire w_dff_A_K4h0biQT9_0;
	wire w_dff_A_OIHn8raU3_0;
	wire w_dff_A_zwbI27Zl7_0;
	wire w_dff_A_qiqBJ46L3_0;
	wire w_dff_A_JuBUJKWv1_0;
	wire w_dff_A_a2gz8XBV4_0;
	wire w_dff_A_fBGxTbSY1_0;
	wire w_dff_A_vLnah9Nh3_0;
	wire w_dff_A_zEGDd7WI3_0;
	wire w_dff_A_G2xREmvo6_0;
	wire w_dff_A_Db0Se1s10_1;
	wire w_dff_A_0yPptQX48_0;
	wire w_dff_A_ve4s6jcr8_0;
	wire w_dff_A_ybX7Iq9q0_0;
	wire w_dff_A_Xvirj3x92_1;
	wire w_dff_A_9HLefwsM7_0;
	wire w_dff_A_ZKR4KOu15_0;
	wire w_dff_A_1vfEAqKj1_0;
	wire w_dff_A_UTqRB3JZ8_0;
	wire w_dff_A_0gsqbsOX9_1;
	wire w_dff_A_2MU3zQs79_0;
	wire w_dff_A_8YV8pcFe0_0;
	wire w_dff_A_clG1kHoL9_0;
	wire w_dff_A_DN5dca3V1_0;
	wire w_dff_A_0s4VnOCC6_0;
	wire w_dff_A_2JE9l8j69_0;
	wire w_dff_A_Y9DXbQ481_1;
	wire w_dff_A_kyD7zK7U1_0;
	wire w_dff_A_1rSdnZCe4_0;
	wire w_dff_A_xdEoz0CS8_0;
	wire w_dff_A_3jeAbU1w5_0;
	wire w_dff_A_NjzqUsoA9_0;
	wire w_dff_A_6yUTm2Ws8_0;
	wire w_dff_A_rCo1GP2Y6_0;
	wire w_dff_A_UTwmXiJV5_2;
	wire w_dff_A_TXy3L1NG6_0;
	wire w_dff_A_fWRL19Y44_0;
	wire w_dff_A_cpxnTtkT7_2;
	wire w_dff_A_DkB9eyZc1_0;
	wire w_dff_A_vkSUaR3g5_0;
	wire w_dff_A_zT3XBVAo1_2;
	wire w_dff_A_DUQ5RHt73_0;
	wire w_dff_A_3mGJs6Ph6_0;
	wire w_dff_A_Wh7K7oZ84_0;
	wire w_dff_A_8UD0c5Ru2_2;
	wire w_dff_A_tWlDItD29_0;
	wire w_dff_A_AqPdayHI6_0;
	wire w_dff_A_nF3iWpjD1_0;
	wire w_dff_A_PIldz9RX9_2;
	wire w_dff_A_sD9RiPX72_0;
	wire w_dff_A_WO8lGLWg1_0;
	wire w_dff_A_u65Zf4pJ9_0;
	wire w_dff_A_EWnvNPoH7_0;
	wire w_dff_A_zLFP5pWE0_2;
	wire w_dff_A_ngOjbvSY8_0;
	wire w_dff_A_YB3NsWiX5_0;
	wire w_dff_A_4jrRbgWU5_0;
	wire w_dff_A_Jc6Rpzbn3_2;
	wire w_dff_A_USWGTGjs0_0;
	wire w_dff_A_AYIiujB36_0;
	wire w_dff_A_2oSbqiNS6_0;
	wire w_dff_A_W3LY4oTh8_2;
	wire w_dff_A_p4Z6OHCa9_0;
	wire w_dff_A_Uh9DHK8c5_0;
	wire w_dff_A_mtX3FGsz2_0;
	wire w_dff_A_TCsuykfJ9_0;
	wire w_dff_A_FMg1FwX22_2;
	wire w_dff_A_oMhcGBxd0_0;
	wire w_dff_A_DlsGPHEV0_0;
	wire w_dff_A_R2caKM6X3_0;
	wire w_dff_A_1QlhlnXk4_2;
	wire w_dff_A_0phmmXY59_0;
	wire w_dff_A_9HeNAnN46_0;
	wire w_dff_A_yqoRBsWS7_2;
	wire w_dff_A_HJOc8wDx5_0;
	wire w_dff_A_wNH9s7Zb0_0;
	wire w_dff_A_GDUy23aV8_2;
	wire w_dff_A_3cv1kEqb2_0;
	wire w_dff_A_Koy1Jatt2_2;
	wire w_dff_A_2UHCS21P1_0;
	wire w_dff_A_gmRVeP8O9_0;
	wire w_dff_A_TAD277UN8_0;
	wire w_dff_A_pBwC6pVv9_2;
	wire w_dff_A_uRcD19pB1_0;
	wire w_dff_A_gRXC4Tr85_0;
	wire w_dff_A_R1XS5Ihe0_2;
	wire w_dff_A_gk80YyZu3_0;
	wire w_dff_A_tBzr0fGn3_0;
	wire w_dff_A_8T6yUygj4_2;
	wire w_dff_A_83ihCwOD9_0;
	wire w_dff_A_SURhQcVE9_2;
	wire w_dff_A_5JQSpGdh3_0;
	wire w_dff_A_IphPcu077_0;
	wire w_dff_A_pNCoGSMR1_0;
	wire w_dff_A_uG8smKgl3_2;
	wire w_dff_A_YDRa4Cqv9_0;
	wire w_dff_A_Gb01iVMQ7_0;
	wire w_dff_A_B66RrRug7_0;
	wire w_dff_A_jKaG1UkO8_2;
	wire w_dff_A_1hgo6KA25_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_xnuHcXtR9_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(G366),.dout(G600_fa_),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_5UiApBuf0_1),.clk(gclk));
	jdff g0005(.din(G338),.dout(G611_fa_),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_xWfJIjhY9_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_DKH03zRr9_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_C4E6I9xm8_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_IneqafsU3_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_1xSfMYMt0_1),.clk(gclk));
	jor g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_ZCfZqptZ2_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_XssIjf5V0_1),.dout(w_dff_A_85EWI87F1_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_Dal5NXoy4_0),.dinb(w_n316_0[1]),.dout(w_dff_A_wbIT1XPG9_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_baaaIop22_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_Mca1lwmy8_1),.dout(w_dff_A_keD9V7g93_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_Fm0mRtxx3_1),.dout(w_dff_A_5DKWnxSc5_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_CXKw5YL30_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_S57yGqN83_1),.dout(w_dff_A_9yC0VVfO7_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_KSZfTLzP9_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_IrVW51x29_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_fnTBsdyL9_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_rizW0C430_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_Jfk8n5Ey8_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_TiA3PYaH3_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_ODt69OBG6_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_elugQIR87_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_cVsNJJHb0_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_p9XI6owv5_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_Gkskymn36_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_FaokHENP3_2),.clk(gclk));
	jand g0054(.dina(w_n326_0[2]),.dinb(w_dff_B_dEkF10QY7_1),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_G2358_0[2]),.dinb(G80),.dout(n356),.clk(gclk));
	jor g0056(.dina(w_dff_B_aSvu7Tg51_0),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_JmCqyBqc5_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_xsbWQ4I27_2),.clk(gclk));
	jnot g0059(.din(w_G308_1[2]),.dout(n360),.clk(gclk));
	jand g0060(.dina(w_n360_0[1]),.dinb(w_G251_4[2]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G479_1[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(w_G308_1[1]),.dinb(w_G248_5[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_n362_0[1]),.dout(n364),.clk(gclk));
	jor g0064(.dina(n364),.dinb(n361),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G254_1[2]),.dout(n366),.clk(gclk));
	jand g0066(.dina(w_n360_0[0]),.dinb(w_n366_4[2]),.dout(n367),.clk(gclk));
	jnot g0067(.din(w_G242_1[2]),.dout(n368),.clk(gclk));
	jand g0068(.dina(w_G308_1[0]),.dinb(w_n368_5[1]),.dout(n369),.clk(gclk));
	jor g0069(.dina(n369),.dinb(w_G479_1[0]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(w_dff_B_Ad7FIs4t6_1),.dout(n371),.clk(gclk));
	jand g0071(.dina(n371),.dinb(w_dff_B_DYaX8Hgu3_1),.dout(n372),.clk(gclk));
	jnot g0072(.din(w_G316_1[2]),.dout(n373),.clk(gclk));
	jand g0073(.dina(w_n373_0[1]),.dinb(w_G251_4[1]),.dout(n374),.clk(gclk));
	jnot g0074(.din(w_G490_1[2]),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_G316_1[1]),.dinb(w_G248_5[0]),.dout(n376),.clk(gclk));
	jor g0076(.dina(n376),.dinb(n375),.dout(n377),.clk(gclk));
	jor g0077(.dina(n377),.dinb(n374),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n373_0[0]),.dinb(w_n366_4[1]),.dout(n379),.clk(gclk));
	jand g0079(.dina(w_G316_1[0]),.dinb(w_n368_5[0]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_G490_1[1]),.dout(n381),.clk(gclk));
	jor g0081(.dina(n381),.dinb(w_dff_B_HrGeroVV9_1),.dout(n382),.clk(gclk));
	jand g0082(.dina(n382),.dinb(w_dff_B_Nsmg6kdC0_1),.dout(n383),.clk(gclk));
	jand g0083(.dina(w_n383_0[2]),.dinb(w_n372_0[2]),.dout(n384),.clk(gclk));
	jnot g0084(.din(w_G351_2[2]),.dout(n385),.clk(gclk));
	jnot g0085(.din(G3550),.dout(n386),.clk(gclk));
	jand g0086(.dina(w_n386_4[2]),.dinb(w_n385_1[2]),.dout(n387),.clk(gclk));
	jnot g0087(.din(w_G534_1[2]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G3552_0[1]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n389_4[2]),.dinb(w_G351_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n388_1[2]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(w_dff_B_ME1rjpGW3_1),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3548_4[2]),.dinb(w_n385_1[1]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3546_5[1]),.dinb(w_G351_2[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_G534_1[1]),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0096(.dina(w_dff_B_hpRNacob3_0),.dinb(n392),.dout(n397),.clk(gclk));
	jnot g0097(.din(w_G293_0[2]),.dout(n398),.clk(gclk));
	jand g0098(.dina(w_n398_0[2]),.dinb(w_n366_4[0]),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G293_0[1]),.dinb(w_n368_4[2]),.dout(n400),.clk(gclk));
	jor g0100(.dina(n400),.dinb(n399),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G251_4[0]),.dout(n402),.clk(gclk));
	jnot g0102(.din(w_G302_0[2]),.dout(n403),.clk(gclk));
	jand g0103(.dina(w_n403_0[1]),.dinb(w_n402_2[1]),.dout(n404),.clk(gclk));
	jnot g0104(.din(w_G248_4[2]),.dout(n405),.clk(gclk));
	jand g0105(.dina(w_G302_0[1]),.dinb(w_n405_2[1]),.dout(n406),.clk(gclk));
	jor g0106(.dina(n406),.dinb(n404),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_n407_0[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_n408_0[1]),.dinb(w_n401_0[2]),.dout(n409),.clk(gclk));
	jnot g0109(.din(w_G514_1[1]),.dout(n410),.clk(gclk));
	jnot g0110(.din(w_G3546_5[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(w_n410_1[1]),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G3552_0[0]),.dinb(w_G514_1[0]),.dout(n413),.clk(gclk));
	jor g0113(.dina(w_dff_B_Zz6Hvt2A8_0),.dinb(n412),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_n414_0[1]),.dout(n415),.clk(gclk));
	jnot g0115(.din(w_G361_0[2]),.dout(n416),.clk(gclk));
	jand g0116(.dina(w_n416_0[1]),.dinb(w_n402_2[0]),.dout(n417),.clk(gclk));
	jand g0117(.dina(w_G361_0[1]),.dinb(w_n405_2[0]),.dout(n418),.clk(gclk));
	jor g0118(.dina(n418),.dinb(n417),.dout(n419),.clk(gclk));
	jnot g0119(.din(w_n419_0[2]),.dout(n420),.clk(gclk));
	jand g0120(.dina(n420),.dinb(n415),.dout(n421),.clk(gclk));
	jand g0121(.dina(n421),.dinb(n409),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(w_n397_0[1]),.dout(n423),.clk(gclk));
	jnot g0123(.din(w_G324_1[2]),.dout(n424),.clk(gclk));
	jand g0124(.dina(w_n386_4[1]),.dinb(w_n424_2[1]),.dout(n425),.clk(gclk));
	jnot g0125(.din(w_G503_1[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_n389_4[1]),.dinb(w_G324_1[1]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(w_n426_0[1]),.dout(n428),.clk(gclk));
	jor g0128(.dina(n428),.dinb(w_dff_B_9iNE9XXP0_1),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_G3548_4[1]),.dinb(w_n424_2[0]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G3546_4[2]),.dinb(w_G324_1[0]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(w_G503_1[1]),.dout(n432),.clk(gclk));
	jor g0132(.dina(n432),.dinb(n430),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_dff_B_6x1nUjZV6_0),.dinb(n429),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G341_2[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n386_4[0]),.dinb(w_n435_1[2]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G523_1[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n389_4[0]),.dinb(w_G341_2[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_1[2]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(w_dff_B_AHuoukWT8_1),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3548_4[0]),.dinb(w_n435_1[1]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3546_4[1]),.dinb(w_G341_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_G523_1[0]),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(n441),.dout(n444),.clk(gclk));
	jand g0144(.dina(w_dff_B_90sOMuAW5_0),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(w_n434_0[1]),.dout(n446),.clk(gclk));
	jand g0146(.dina(w_dff_B_Nz0flp8Q2_0),.dinb(n423),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(w_dff_B_3CzV9Jej8_1),.dout(w_dff_A_BEb53Iaq1_2),.clk(gclk));
	jnot g0148(.din(w_G265_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n386_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G400_1[1]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n389_3[2]),.dinb(w_G265_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_1[1]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(w_dff_B_v0xWcDdw6_1),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3546_4[0]),.dinb(w_G265_1[2]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_G400_1[0]),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(n455),.dout(n458),.clk(gclk));
	jand g0158(.dina(w_dff_B_YwJWY0nX7_0),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n386_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n389_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(w_dff_B_4NDoHUfP4_1),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_G435_1[1]),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(n466),.dout(n469),.clk(gclk));
	jand g0169(.dina(w_dff_B_FGBLF5RG1_0),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G257_2[2]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n386_3[0]),.dinb(w_n471_1[1]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G389_0[2]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n389_3[0]),.dinb(w_G257_2[1]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[2]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(w_dff_B_XnnT7VXe0_1),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3548_3[0]),.dinb(w_n471_1[0]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3546_3[1]),.dinb(w_G257_2[0]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_G389_0[1]),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(n477),.dout(n480),.clk(gclk));
	jand g0180(.dina(w_dff_B_twvL3bjd5_0),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jand g0182(.dina(n482),.dinb(w_n459_0[1]),.dout(n483),.clk(gclk));
	jnot g0183(.din(w_G273_2[2]),.dout(n484),.clk(gclk));
	jand g0184(.dina(w_n386_2[2]),.dinb(w_n484_1[1]),.dout(n485),.clk(gclk));
	jnot g0185(.din(w_G411_0[2]),.dout(n486),.clk(gclk));
	jand g0186(.dina(w_n389_2[2]),.dinb(w_G273_2[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_n486_1[1]),.dout(n488),.clk(gclk));
	jor g0188(.dina(n488),.dinb(w_dff_B_9BFouGyv7_1),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n484_1[0]),.dout(n490),.clk(gclk));
	jand g0190(.dina(w_G3546_3[0]),.dinb(w_G273_2[0]),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G411_0[1]),.dout(n492),.clk(gclk));
	jor g0192(.dina(n492),.dinb(n490),.dout(n493),.clk(gclk));
	jand g0193(.dina(w_dff_B_NznqOe2n0_0),.dinb(n489),.dout(n494),.clk(gclk));
	jnot g0194(.din(w_G281_2[1]),.dout(n495),.clk(gclk));
	jand g0195(.dina(w_n386_2[1]),.dinb(w_n495_1[2]),.dout(n496),.clk(gclk));
	jnot g0196(.din(w_G374_0[2]),.dout(n497),.clk(gclk));
	jand g0197(.dina(w_n389_2[1]),.dinb(w_G281_2[0]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_n497_1[1]),.dout(n499),.clk(gclk));
	jor g0199(.dina(n499),.dinb(w_dff_B_KjOV1hzk1_1),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n495_1[1]),.dout(n501),.clk(gclk));
	jand g0201(.dina(w_G3546_2[2]),.dinb(w_G281_1[2]),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G374_0[1]),.dout(n503),.clk(gclk));
	jor g0203(.dina(n503),.dinb(n501),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_dff_B_qPKMQyte9_0),.dinb(n500),.dout(n505),.clk(gclk));
	jand g0205(.dina(w_n505_0[1]),.dinb(w_n494_0[1]),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[2]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n386_2[0]),.dinb(w_n507_1[1]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n389_2[0]),.dinb(w_G218_2[1]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[1]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(w_dff_B_ETgeSkvN4_1),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3548_2[0]),.dinb(w_n507_1[0]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3546_2[1]),.dinb(w_G218_2[0]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_G468_1[1]),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(n513),.dout(n516),.clk(gclk));
	jand g0216(.dina(w_dff_B_gG2uUQz25_0),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G206_0[2]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_G251_3[2]),.dinb(w_n518_1[1]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G446_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_G248_4[1]),.dinb(w_G206_0[1]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(n520),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(n519),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_n366_3[2]),.dinb(w_n518_1[0]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_n368_4[1]),.dinb(w_G206_0[0]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_G446_1[1]),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_dff_B_jPvxMSUl7_1),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(w_dff_B_J4fIGD0M8_1),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[2]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G226_2[2]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n386_1[2]),.dinb(w_n530_1[1]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G422_2[1]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n389_1[2]),.dinb(w_G226_2[1]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_0[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(w_dff_B_YdcdSCpG9_1),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3548_1[2]),.dinb(w_n530_1[0]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3546_2[0]),.dinb(w_G226_2[0]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_G422_2[0]),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(n536),.dout(n539),.clk(gclk));
	jand g0239(.dina(w_dff_B_2wflkQor3_0),.dinb(n535),.dout(n540),.clk(gclk));
	jnot g0240(.din(w_G210_2[2]),.dout(n541),.clk(gclk));
	jand g0241(.dina(w_n386_1[1]),.dinb(w_n541_1[1]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G457_2[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_n389_1[1]),.dinb(w_G210_2[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_n543_0[1]),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(w_dff_B_SCzYglrG4_1),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_G3548_1[1]),.dinb(w_n541_1[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_G3546_1[2]),.dinb(w_G210_2[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(w_G457_2[0]),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(n547),.dout(n550),.clk(gclk));
	jand g0250(.dina(w_dff_B_Bb8vETym4_0),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[1]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(w_dff_B_kW56YRH88_1),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_dff_B_pkjSE7L20_1),.dout(w_dff_A_j4efVi3O6_2),.clk(gclk));
	jnot g0255(.din(w_G335_4[1]),.dout(n556),.clk(gclk));
	jor g0256(.dina(w_n556_5[1]),.dinb(w_dff_B_OdDnxJVz1_1),.dout(n557),.clk(gclk));
	jand g0257(.dina(w_n556_5[0]),.dinb(w_n460_1[0]),.dout(n558),.clk(gclk));
	jnot g0258(.din(n558),.dout(n559),.clk(gclk));
	jand g0259(.dina(n559),.dinb(w_dff_B_c5b0SisU2_1),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_1[1]),.dinb(w_G435_1[0]),.dout(n561),.clk(gclk));
	jnot g0261(.din(w_n561_0[2]),.dout(n562),.clk(gclk));
	jnot g0262(.din(G288),.dout(n563),.clk(gclk));
	jand g0263(.dina(w_G335_4[0]),.dinb(n563),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n556_4[2]),.dinb(w_n495_1[0]),.dout(n565),.clk(gclk));
	jor g0265(.dina(n565),.dinb(n564),.dout(n566),.clk(gclk));
	jxor g0266(.dina(w_n566_0[2]),.dinb(w_n497_1[0]),.dout(n567),.clk(gclk));
	jor g0267(.dina(w_n556_4[1]),.dinb(w_G280_0[1]),.dout(n568),.clk(gclk));
	jor g0268(.dina(w_G335_3[2]),.dinb(w_G273_1[2]),.dout(n569),.clk(gclk));
	jand g0269(.dina(w_n569_0[1]),.dinb(n568),.dout(n570),.clk(gclk));
	jxor g0270(.dina(w_n570_0[1]),.dinb(w_n486_1[0]),.dout(n571),.clk(gclk));
	jnot g0271(.din(w_n571_1[1]),.dout(n572),.clk(gclk));
	jand g0272(.dina(w_n572_0[2]),.dinb(w_n567_1[1]),.dout(n573),.clk(gclk));
	jnot g0273(.din(n573),.dout(n574),.clk(gclk));
	jor g0274(.dina(w_n556_4[0]),.dinb(w_dff_B_ex8iQiFj3_1),.dout(n575),.clk(gclk));
	jor g0275(.dina(w_G335_3[1]),.dinb(w_G257_1[2]),.dout(n576),.clk(gclk));
	jand g0276(.dina(w_dff_B_y2DrAnYB0_0),.dinb(n575),.dout(n577),.clk(gclk));
	jxor g0277(.dina(w_n577_0[2]),.dinb(w_n473_1[1]),.dout(n578),.clk(gclk));
	jnot g0278(.din(G272),.dout(n579),.clk(gclk));
	jand g0279(.dina(w_G335_3[0]),.dinb(n579),.dout(n580),.clk(gclk));
	jand g0280(.dina(w_n556_3[2]),.dinb(w_n449_1[0]),.dout(n581),.clk(gclk));
	jor g0281(.dina(n581),.dinb(n580),.dout(n582),.clk(gclk));
	jxor g0282(.dina(w_n582_1[1]),.dinb(w_G400_0[2]),.dout(n583),.clk(gclk));
	jor g0283(.dina(w_n583_1[1]),.dinb(w_n578_0[2]),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_dff_B_SDAncjIu4_0),.dinb(w_n574_0[2]),.dout(n585),.clk(gclk));
	jor g0285(.dina(w_n585_0[1]),.dinb(w_n562_0[1]),.dout(n586),.clk(gclk));
	jnot g0286(.din(n586),.dout(n587),.clk(gclk));
	jor g0287(.dina(w_n556_3[1]),.dinb(w_dff_B_oSc3NJlp1_1),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_2[2]),.dinb(w_G210_1[2]),.dout(n589),.clk(gclk));
	jand g0289(.dina(w_dff_B_7O06H6yB2_0),.dinb(n588),.dout(n590),.clk(gclk));
	jxor g0290(.dina(w_n590_1[1]),.dinb(w_G457_1[2]),.dout(n591),.clk(gclk));
	jor g0291(.dina(w_n556_3[0]),.dinb(w_dff_B_WCFRpAvJ0_1),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_2[2]),.dinb(w_n518_0[2]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jand g0294(.dina(n594),.dinb(w_dff_B_p3feOSO34_1),.dout(n595),.clk(gclk));
	jxor g0295(.dina(w_n595_1[1]),.dinb(w_G446_1[0]),.dout(n596),.clk(gclk));
	jand g0296(.dina(w_n596_0[2]),.dinb(w_n591_0[1]),.dout(n597),.clk(gclk));
	jor g0297(.dina(w_n556_2[1]),.dinb(w_dff_B_PV5733b09_1),.dout(n598),.clk(gclk));
	jor g0298(.dina(w_G335_2[1]),.dinb(w_G226_1[2]),.dout(n599),.clk(gclk));
	jand g0299(.dina(w_dff_B_0rl6XDgm3_0),.dinb(n598),.dout(n600),.clk(gclk));
	jxor g0300(.dina(w_n600_1[1]),.dinb(w_G422_1[2]),.dout(n601),.clk(gclk));
	jor g0301(.dina(w_n556_2[0]),.dinb(w_dff_B_I4f65N7O1_1),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_G335_2[0]),.dinb(w_G218_1[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_dff_B_IrYITDwn2_0),.dinb(n602),.dout(n604),.clk(gclk));
	jxor g0304(.dina(w_n604_0[2]),.dinb(w_G468_1[0]),.dout(n605),.clk(gclk));
	jand g0305(.dina(w_n605_2[2]),.dinb(w_n601_0[1]),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_AeDOD12Z9_0),.dinb(n597),.dout(n607),.clk(gclk));
	jand g0307(.dina(w_n607_0[2]),.dinb(w_n587_1[1]),.dout(w_dff_A_4Xgg3Wdu6_2),.clk(gclk));
	jnot g0308(.din(w_G332_4[2]),.dout(n609),.clk(gclk));
	jor g0309(.dina(w_n609_5[2]),.dinb(w_G331_0[1]),.dout(n610),.clk(gclk));
	jand g0310(.dina(w_n609_5[1]),.dinb(w_n424_1[2]),.dout(n611),.clk(gclk));
	jnot g0311(.din(n611),.dout(n612),.clk(gclk));
	jand g0312(.dina(n612),.dinb(w_dff_B_rYGqbmNG0_1),.dout(n613),.clk(gclk));
	jxor g0313(.dina(w_n613_0[2]),.dinb(w_G503_1[0]),.dout(n614),.clk(gclk));
	jor g0314(.dina(w_G358_0[0]),.dinb(w_n609_5[0]),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_G351_1[2]),.dinb(w_G332_4[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(w_dff_B_rkiHOKfh7_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_n388_1[1]),.dout(n618),.clk(gclk));
	jand g0318(.dina(w_G600_0),.dinb(w_G332_4[0]),.dout(n619),.clk(gclk));
	jand g0319(.dina(w_n416_0[0]),.dinb(w_n609_4[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(n620),.dinb(n619),.dout(n621),.clk(gclk));
	jnot g0321(.din(w_n621_2[1]),.dout(n622),.clk(gclk));
	jor g0322(.dina(w_n622_1[1]),.dinb(w_n618_1[1]),.dout(n623),.clk(gclk));
	jand g0323(.dina(w_G611_0),.dinb(w_G332_3[2]),.dout(n624),.clk(gclk));
	jxor g0324(.dina(w_n624_1[2]),.dinb(w_G514_0[2]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G348_0[0]),.dinb(w_n609_4[1]),.dout(n626),.clk(gclk));
	jor g0326(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n627),.clk(gclk));
	jand g0327(.dina(w_dff_B_VrYukKn71_0),.dinb(n626),.dout(n628),.clk(gclk));
	jxor g0328(.dina(w_n628_0[2]),.dinb(w_n437_1[1]),.dout(n629),.clk(gclk));
	jor g0329(.dina(w_n629_0[2]),.dinb(w_n625_0[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(w_n623_0[1]),.dout(n631),.clk(gclk));
	jnot g0331(.din(w_n631_0[1]),.dout(n632),.clk(gclk));
	jand g0332(.dina(n632),.dinb(w_n614_2[1]),.dout(n633),.clk(gclk));
	jand g0333(.dina(w_G332_3[0]),.dinb(w_G593_0),.dout(n634),.clk(gclk));
	jand g0334(.dina(w_n609_4[0]),.dinb(w_n398_0[1]),.dout(n635),.clk(gclk));
	jor g0335(.dina(n635),.dinb(n634),.dout(n636),.clk(gclk));
	jor g0336(.dina(w_n609_3[2]),.dinb(w_dff_B_9MSpMEdm3_1),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n609_3[1]),.dinb(w_n403_0[0]),.dout(n638),.clk(gclk));
	jnot g0338(.din(n638),.dout(n639),.clk(gclk));
	jand g0339(.dina(n639),.dinb(w_dff_B_y2tM4x287_1),.dout(n640),.clk(gclk));
	jnot g0340(.din(w_n640_1[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n641_0[1]),.dinb(w_n636_1[1]),.dout(n642),.clk(gclk));
	jor g0342(.dina(w_n609_3[0]),.dinb(w_dff_B_Ku26dCwl2_1),.dout(n643),.clk(gclk));
	jor g0343(.dina(w_G332_2[2]),.dinb(w_G308_0[2]),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_dff_B_kjeHPyV10_0),.dinb(n643),.dout(n645),.clk(gclk));
	jxor g0345(.dina(w_n645_0[2]),.dinb(w_G479_0[2]),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n609_2[2]),.dinb(w_dff_B_d9S4yyXW1_1),.dout(n647),.clk(gclk));
	jor g0347(.dina(w_G332_2[1]),.dinb(w_G316_0[2]),.dout(n648),.clk(gclk));
	jand g0348(.dina(w_dff_B_5BaMNZE13_0),.dinb(n647),.dout(n649),.clk(gclk));
	jxor g0349(.dina(w_n649_1[1]),.dinb(w_G490_1[0]),.dout(n650),.clk(gclk));
	jand g0350(.dina(w_n650_0[1]),.dinb(w_n646_0[2]),.dout(n651),.clk(gclk));
	jand g0351(.dina(w_n651_1[1]),.dinb(w_n642_0[1]),.dout(n652),.clk(gclk));
	jand g0352(.dina(w_n652_0[1]),.dinb(w_n633_1[1]),.dout(w_dff_A_n3GGxwow0_2),.clk(gclk));
	jxor g0353(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n654),.clk(gclk));
	jxor g0354(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n655),.clk(gclk));
	jxor g0355(.dina(n655),.dinb(n654),.dout(n656),.clk(gclk));
	jxor g0356(.dina(w_G369_0[1]),.dinb(w_G361_0[0]),.dout(n657),.clk(gclk));
	jxor g0357(.dina(n657),.dinb(w_n424_1[1]),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_G302_0[0]),.dinb(w_n398_0[0]),.dout(n659),.clk(gclk));
	jxor g0359(.dina(n659),.dinb(n658),.dout(n660),.clk(gclk));
	jxor g0360(.dina(n660),.dinb(w_dff_B_UFlG5cKM3_1),.dout(n661),.clk(gclk));
	jnot g0361(.din(w_n661_0[1]),.dout(w_dff_A_8MThqmXy2_1),.clk(gclk));
	jxor g0362(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G273_1[1]),.dinb(w_G265_1[1]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(n667),.dinb(n666),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_G210_1[1]),.dinb(w_n518_0[1]),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n668),.dout(n670),.clk(gclk));
	jxor g0370(.dina(n670),.dinb(w_dff_B_QE8FytI96_1),.dout(n671),.clk(gclk));
	jnot g0371(.din(w_n671_0[1]),.dout(w_dff_A_FM7ga7ou8_1),.clk(gclk));
	jnot g0372(.din(w_n560_1[0]),.dout(n673),.clk(gclk));
	jand g0373(.dina(n673),.dinb(w_n462_0[1]),.dout(n674),.clk(gclk));
	jnot g0374(.din(n674),.dout(n675),.clk(gclk));
	jand g0375(.dina(w_n560_0[2]),.dinb(w_G435_0[2]),.dout(n676),.clk(gclk));
	jnot g0376(.din(w_n577_0[1]),.dout(n677),.clk(gclk));
	jand g0377(.dina(w_n677_0[1]),.dinb(w_n473_1[0]),.dout(n678),.clk(gclk));
	jor g0378(.dina(w_n677_0[0]),.dinb(w_n473_0[2]),.dout(n679),.clk(gclk));
	jand g0379(.dina(w_n582_1[0]),.dinb(w_n451_1[0]),.dout(n680),.clk(gclk));
	jor g0380(.dina(w_n566_0[1]),.dinb(w_n497_0[2]),.dout(n681),.clk(gclk));
	jor g0381(.dina(w_n571_1[0]),.dinb(w_n681_2[1]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_G280_0[0]),.dout(n683),.clk(gclk));
	jand g0383(.dina(w_G335_1[2]),.dinb(n683),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n569_0[0]),.dout(n685),.clk(gclk));
	jor g0385(.dina(n685),.dinb(n684),.dout(n686),.clk(gclk));
	jor g0386(.dina(n686),.dinb(w_n486_0[2]),.dout(n687),.clk(gclk));
	jor g0387(.dina(w_n582_0[2]),.dinb(w_n451_0[2]),.dout(n688),.clk(gclk));
	jand g0388(.dina(n688),.dinb(w_n687_0[2]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n682_0[1]),.dout(n690),.clk(gclk));
	jor g0390(.dina(n690),.dinb(w_n680_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n691_0[2]),.dinb(w_n679_0[1]),.dout(n692),.clk(gclk));
	jor g0392(.dina(n692),.dinb(w_n678_0[1]),.dout(n693),.clk(gclk));
	jnot g0393(.din(w_n693_0[2]),.dout(n694),.clk(gclk));
	jor g0394(.dina(n694),.dinb(w_dff_B_1PaqHFXG2_1),.dout(n695),.clk(gclk));
	jand g0395(.dina(n695),.dinb(w_dff_B_ahsHh9Ol7_1),.dout(n696),.clk(gclk));
	jand g0396(.dina(w_n696_0[2]),.dinb(w_n607_0[1]),.dout(n697),.clk(gclk));
	jand g0397(.dina(w_n595_1[0]),.dinb(w_G446_0[2]),.dout(n698),.clk(gclk));
	jor g0398(.dina(w_n595_0[2]),.dinb(w_G446_0[1]),.dout(n699),.clk(gclk));
	jor g0399(.dina(w_n590_1[0]),.dinb(w_G457_1[1]),.dout(n700),.clk(gclk));
	jand g0400(.dina(w_n590_0[2]),.dinb(w_G457_1[0]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n604_0[1]),.dinb(w_G468_0[2]),.dout(n702),.clk(gclk));
	jand g0402(.dina(w_n600_1[0]),.dinb(w_G422_1[1]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n605_2[1]),.dinb(w_n703_0[2]),.dout(n704),.clk(gclk));
	jor g0404(.dina(n704),.dinb(w_n702_0[1]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n705_0[1]),.dinb(w_dff_B_zHdUCnVa4_1),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n706_0[1]),.dinb(w_n700_0[1]),.dout(n707),.clk(gclk));
	jand g0407(.dina(w_n707_0[2]),.dinb(w_dff_B_fnflHZ8W5_1),.dout(n708),.clk(gclk));
	jor g0408(.dina(n708),.dinb(w_dff_B_7XrR9Fu38_1),.dout(n709),.clk(gclk));
	jor g0409(.dina(w_n709_0[1]),.dinb(w_n697_0[1]),.dout(w_dff_A_x5Bdeqtt8_2),.clk(gclk));
	jand g0410(.dina(w_n613_0[1]),.dinb(w_G503_0[2]),.dout(n711),.clk(gclk));
	jor g0411(.dina(w_n624_1[1]),.dinb(w_n410_1[0]),.dout(n712),.clk(gclk));
	jand g0412(.dina(w_n624_1[0]),.dinb(w_n410_0[2]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_G599_0),.dinb(w_G332_2[0]),.dout(n714),.clk(gclk));
	jand g0414(.dina(w_n435_1[0]),.dinb(w_n609_2[1]),.dout(n715),.clk(gclk));
	jor g0415(.dina(n715),.dinb(n714),.dout(n716),.clk(gclk));
	jand g0416(.dina(w_n716_0[1]),.dinb(w_n437_1[0]),.dout(n717),.clk(gclk));
	jand g0417(.dina(w_G612_0),.dinb(w_G332_1[2]),.dout(n718),.clk(gclk));
	jand g0418(.dina(w_n385_1[0]),.dinb(w_n609_2[0]),.dout(n719),.clk(gclk));
	jor g0419(.dina(n719),.dinb(n718),.dout(n720),.clk(gclk));
	jand g0420(.dina(w_n720_0[1]),.dinb(w_n388_1[0]),.dout(n721),.clk(gclk));
	jor g0421(.dina(w_n621_2[0]),.dinb(w_n721_0[2]),.dout(n722),.clk(gclk));
	jor g0422(.dina(w_n720_0[0]),.dinb(w_n388_0[2]),.dout(n723),.clk(gclk));
	jor g0423(.dina(w_n716_0[0]),.dinb(w_n437_0[2]),.dout(n724),.clk(gclk));
	jand g0424(.dina(n724),.dinb(w_n723_0[1]),.dout(n725),.clk(gclk));
	jand g0425(.dina(n725),.dinb(n722),.dout(n726),.clk(gclk));
	jor g0426(.dina(w_n726_0[1]),.dinb(w_n717_0[2]),.dout(n727),.clk(gclk));
	jor g0427(.dina(w_n727_0[2]),.dinb(w_dff_B_J8ZZvl7V7_1),.dout(n728),.clk(gclk));
	jand g0428(.dina(n728),.dinb(w_dff_B_boRSAyMn0_1),.dout(n729),.clk(gclk));
	jnot g0429(.din(w_n729_1[1]),.dout(n730),.clk(gclk));
	jand g0430(.dina(n730),.dinb(w_n614_2[0]),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_dff_B_UwWcPl1b7_1),.dout(n732),.clk(gclk));
	jand g0432(.dina(w_n732_0[2]),.dinb(w_n651_1[0]),.dout(n733),.clk(gclk));
	jnot g0433(.din(w_n642_0[0]),.dout(n734),.clk(gclk));
	jnot g0434(.din(w_n645_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[1]),.dinb(w_n362_0[0]),.dout(n736),.clk(gclk));
	jnot g0436(.din(w_n736_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n645_0[0]),.dinb(w_G479_0[1]),.dout(n738),.clk(gclk));
	jand g0438(.dina(w_n649_1[0]),.dinb(w_G490_0[2]),.dout(n739),.clk(gclk));
	jor g0439(.dina(w_n739_1[1]),.dinb(n738),.dout(n740),.clk(gclk));
	jand g0440(.dina(w_n740_0[1]),.dinb(n737),.dout(n741),.clk(gclk));
	jor g0441(.dina(w_n741_0[1]),.dinb(n734),.dout(n742),.clk(gclk));
	jor g0442(.dina(w_n742_0[1]),.dinb(w_n733_0[1]),.dout(w_dff_A_dUvFZuI17_2),.clk(gclk));
	jnot g0443(.din(w_G54_0[1]),.dout(n744),.clk(gclk));
	jxor g0444(.dina(w_n621_1[2]),.dinb(w_n744_1[2]),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_G4092_1[2]),.dout(n746),.clk(gclk));
	jand g0446(.dina(w_n746_1[2]),.dinb(w_G4091_2[2]),.dout(n747),.clk(gclk));
	jnot g0447(.din(w_n747_3[2]),.dout(n748),.clk(gclk));
	jor g0448(.dina(w_n748_4[1]),.dinb(n745),.dout(n749),.clk(gclk));
	jnot g0449(.din(w_G4091_2[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n746_1[1]),.dinb(w_n750_1[1]),.dout(n751),.clk(gclk));
	jand g0451(.dina(w_n751_2[1]),.dinb(w_n419_0[1]),.dout(n752),.clk(gclk));
	jand g0452(.dina(w_G4092_1[1]),.dinb(w_n750_1[0]),.dout(n753),.clk(gclk));
	jand g0453(.dina(w_n753_8[1]),.dinb(w_dff_B_QRg1MG1I3_1),.dout(n754),.clk(gclk));
	jor g0454(.dina(w_dff_B_B227RsBo4_0),.dinb(n752),.dout(n755),.clk(gclk));
	jnot g0455(.din(n755),.dout(n756),.clk(gclk));
	jand g0456(.dina(n756),.dinb(w_dff_B_wwrx8AHY9_1),.dout(G822_fa_),.clk(gclk));
	jnot g0457(.din(w_n618_1[0]),.dout(n758),.clk(gclk));
	jand g0458(.dina(w_n621_1[1]),.dinb(w_n744_1[1]),.dout(n759),.clk(gclk));
	jnot g0459(.din(w_n759_0[1]),.dout(n760),.clk(gclk));
	jand g0460(.dina(w_n760_0[1]),.dinb(n758),.dout(n761),.clk(gclk));
	jand g0461(.dina(w_n759_0[0]),.dinb(w_n618_0[2]),.dout(n762),.clk(gclk));
	jor g0462(.dina(n762),.dinb(w_n748_4[0]),.dout(n763),.clk(gclk));
	jor g0463(.dina(n763),.dinb(w_n761_0[1]),.dout(n764),.clk(gclk));
	jnot g0464(.din(w_n751_2[0]),.dout(n765),.clk(gclk));
	jor g0465(.dina(w_n765_5[2]),.dinb(w_n397_0[0]),.dout(n766),.clk(gclk));
	jand g0466(.dina(w_n753_8[0]),.dinb(w_dff_B_UlMVrDl49_1),.dout(n767),.clk(gclk));
	jnot g0467(.din(n767),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_dff_B_Dplxahew3_0),.dinb(n766),.dout(n769),.clk(gclk));
	jand g0469(.dina(n769),.dinb(n764),.dout(G838_fa_),.clk(gclk));
	jxor g0470(.dina(w_n567_1[0]),.dinb(w_G4_1[1]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n771_0[1]),.dinb(w_n747_3[1]),.dout(n772),.clk(gclk));
	jnot g0472(.din(n772),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_n765_5[1]),.dinb(w_n505_0[0]),.dout(n774),.clk(gclk));
	jand g0474(.dina(w_n753_7[2]),.dinb(w_dff_B_gUgiBgL93_1),.dout(n775),.clk(gclk));
	jnot g0475(.din(n775),.dout(n776),.clk(gclk));
	jand g0476(.dina(w_dff_B_33JdFQzd1_0),.dinb(n774),.dout(n777),.clk(gclk));
	jand g0477(.dina(n777),.dinb(n773),.dout(G861_fa_),.clk(gclk));
	jnot g0478(.din(w_n636_1[0]),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n633_1[0]),.dinb(w_G54_0[0]),.dout(n780),.clk(gclk));
	jor g0480(.dina(w_dff_B_enuUWqnO6_0),.dinb(w_n732_0[1]),.dout(n781),.clk(gclk));
	jand g0481(.dina(w_n781_0[2]),.dinb(w_n651_0[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(n782),.dinb(w_n741_0[0]),.dout(n783),.clk(gclk));
	jnot g0483(.din(w_n783_1[1]),.dout(n784),.clk(gclk));
	jor g0484(.dina(n784),.dinb(w_n779_0[1]),.dout(n785),.clk(gclk));
	jxor g0485(.dina(w_n640_1[1]),.dinb(w_n779_0[0]),.dout(n786),.clk(gclk));
	jnot g0486(.din(w_n786_0[1]),.dout(n787),.clk(gclk));
	jor g0487(.dina(w_n787_0[1]),.dinb(w_n783_1[0]),.dout(n788),.clk(gclk));
	jand g0488(.dina(w_dff_B_BCyhDCpA1_0),.dinb(n785),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n789_0[2]),.dout(w_dff_A_ThmdqykU8_1),.clk(gclk));
	jnot g0490(.din(w_G861_0),.dout(n791),.clk(gclk));
	jnot g0491(.din(w_G4087_0[2]),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_G4088_0[2]),.dinb(w_n792_0[1]),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n793_4[1]),.dinb(w_n791_1[1]),.dout(n794),.clk(gclk));
	jnot g0494(.din(w_G822_0),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_G4088_0[1]),.dout(n796),.clk(gclk));
	jand g0496(.dina(w_n796_0[1]),.dinb(w_n792_0[0]),.dout(n797),.clk(gclk));
	jand g0497(.dina(w_n797_4[1]),.dinb(w_n795_1[1]),.dout(n798),.clk(gclk));
	jand g0498(.dina(w_n796_0[0]),.dinb(w_G4087_0[1]),.dout(n799),.clk(gclk));
	jand g0499(.dina(w_n799_4[1]),.dinb(w_G11_0[1]),.dout(n800),.clk(gclk));
	jand g0500(.dina(w_G4088_0[0]),.dinb(w_G4087_0[0]),.dout(n801),.clk(gclk));
	jand g0501(.dina(w_n801_4[1]),.dinb(w_G61_0[1]),.dout(n802),.clk(gclk));
	jor g0502(.dina(w_dff_B_viMLJl540_0),.dinb(n800),.dout(n803),.clk(gclk));
	jor g0503(.dina(w_dff_B_3ewiIPnx2_0),.dinb(n798),.dout(n804),.clk(gclk));
	jor g0504(.dina(n804),.dinb(n794),.dout(w_dff_A_ZHMTSP3i6_2),.clk(gclk));
	jand g0505(.dina(w_n729_1[0]),.dinb(w_n631_0[0]),.dout(n806),.clk(gclk));
	jand g0506(.dina(w_n729_0[2]),.dinb(w_n744_1[0]),.dout(n807),.clk(gclk));
	jor g0507(.dina(n807),.dinb(w_n806_0[2]),.dout(n808),.clk(gclk));
	jxor g0508(.dina(n808),.dinb(w_n614_1[2]),.dout(n809),.clk(gclk));
	jor g0509(.dina(w_n809_0[1]),.dinb(w_n748_3[2]),.dout(n810),.clk(gclk));
	jor g0510(.dina(w_n765_5[0]),.dinb(w_n434_0[0]),.dout(n811),.clk(gclk));
	jand g0511(.dina(w_n753_7[1]),.dinb(w_dff_B_TXDqdpuD8_1),.dout(n812),.clk(gclk));
	jnot g0512(.din(n812),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_dff_B_FDZowcrK5_0),.dinb(n811),.dout(n814),.clk(gclk));
	jand g0514(.dina(w_dff_B_6PCInH3y0_0),.dinb(n810),.dout(G832_fa_),.clk(gclk));
	jnot g0515(.din(w_n625_0[1]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n727_0[1]),.dinb(w_n744_0[2]),.dout(n817),.clk(gclk));
	jand g0517(.dina(w_n726_0[0]),.dinb(w_n623_0[0]),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n717_0[1]),.dout(n819),.clk(gclk));
	jor g0519(.dina(w_n819_0[1]),.dinb(n817),.dout(n820),.clk(gclk));
	jxor g0520(.dina(n820),.dinb(w_dff_B_ltmbQhDK8_1),.dout(n821),.clk(gclk));
	jor g0521(.dina(w_n821_0[1]),.dinb(w_n748_3[1]),.dout(n822),.clk(gclk));
	jand g0522(.dina(w_n751_1[2]),.dinb(w_n414_0[0]),.dout(n823),.clk(gclk));
	jand g0523(.dina(w_n753_7[0]),.dinb(w_dff_B_eRjeDWEg4_1),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_dff_B_J1JxYypK8_0),.dinb(n823),.dout(n825),.clk(gclk));
	jnot g0525(.din(n825),.dout(n826),.clk(gclk));
	jand g0526(.dina(w_dff_B_yl3JbdgC0_0),.dinb(n822),.dout(G834_fa_),.clk(gclk));
	jor g0527(.dina(w_n617_1[0]),.dinb(w_G534_1[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n617_0[2]),.dinb(w_G534_0[2]),.dout(n829),.clk(gclk));
	jor g0529(.dina(w_n760_0[0]),.dinb(w_n829_0[1]),.dout(n830),.clk(gclk));
	jand g0530(.dina(n830),.dinb(w_n828_0[2]),.dout(n831),.clk(gclk));
	jxor g0531(.dina(n831),.dinb(w_n629_0[1]),.dout(n832),.clk(gclk));
	jor g0532(.dina(w_n832_0[1]),.dinb(w_n748_3[0]),.dout(n833),.clk(gclk));
	jor g0533(.dina(w_n765_4[2]),.dinb(w_n445_0[0]),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n753_6[2]),.dinb(w_dff_B_oO4A8jg59_1),.dout(n835),.clk(gclk));
	jnot g0535(.din(n835),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_dff_B_qQWnhljy2_0),.dinb(n834),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_dff_B_folb1ScY3_0),.dinb(n833),.dout(G836_fa_),.clk(gclk));
	jnot g0538(.din(w_G4090_0[2]),.dout(n839),.clk(gclk));
	jand g0539(.dina(w_n839_0[1]),.dinb(w_G4089_0[2]),.dout(n840),.clk(gclk));
	jand g0540(.dina(w_n840_4[1]),.dinb(w_n791_1[0]),.dout(n841),.clk(gclk));
	jnot g0541(.din(w_G4089_0[1]),.dout(n842),.clk(gclk));
	jand g0542(.dina(w_n839_0[0]),.dinb(w_n842_0[1]),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n843_4[1]),.dinb(w_n795_1[0]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_G4090_0[1]),.dinb(w_n842_0[0]),.dout(n845),.clk(gclk));
	jand g0545(.dina(w_n845_4[1]),.dinb(w_G11_0[0]),.dout(n846),.clk(gclk));
	jand g0546(.dina(w_G4090_0[0]),.dinb(w_G4089_0[0]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_4[1]),.dinb(w_G61_0[0]),.dout(n848),.clk(gclk));
	jor g0548(.dina(w_dff_B_yMh7HUE44_0),.dinb(n846),.dout(n849),.clk(gclk));
	jor g0549(.dina(w_dff_B_U2olVBQR0_0),.dinb(n844),.dout(n850),.clk(gclk));
	jor g0550(.dina(n850),.dinb(n841),.dout(w_dff_A_7O2wzkaw1_2),.clk(gclk));
	jnot g0551(.din(w_n678_0[0]),.dout(n852),.clk(gclk));
	jnot g0552(.din(w_n679_0[0]),.dout(n853),.clk(gclk));
	jor g0553(.dina(w_n583_1[0]),.dinb(w_n574_0[1]),.dout(n854),.clk(gclk));
	jand g0554(.dina(n854),.dinb(w_n691_0[1]),.dout(n855),.clk(gclk));
	jnot g0555(.din(w_n855_0[1]),.dout(n856),.clk(gclk));
	jnot g0556(.din(w_n691_0[0]),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n857_0[1]),.dinb(w_G4_1[0]),.dout(n858),.clk(gclk));
	jand g0558(.dina(w_dff_B_orm6dmTT0_0),.dinb(w_n856_0[1]),.dout(n859),.clk(gclk));
	jor g0559(.dina(w_n859_0[1]),.dinb(w_n853_0[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(w_dff_B_73bDIewy7_1),.dout(n861),.clk(gclk));
	jxor g0561(.dina(n861),.dinb(w_n562_0[0]),.dout(n862),.clk(gclk));
	jor g0562(.dina(w_n862_0[1]),.dinb(w_n748_2[2]),.dout(n863),.clk(gclk));
	jor g0563(.dina(w_n765_4[1]),.dinb(w_n470_0[0]),.dout(n864),.clk(gclk));
	jand g0564(.dina(w_n753_6[1]),.dinb(w_dff_B_Pvx58Jyu8_1),.dout(n865),.clk(gclk));
	jnot g0565(.din(n865),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_dff_B_WUOp7OYO9_0),.dinb(n864),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_dff_B_94rHWRBM0_0),.dinb(n863),.dout(G871_fa_),.clk(gclk));
	jxor g0568(.dina(w_n859_0[0]),.dinb(w_n578_0[1]),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_n869_0[1]),.dinb(w_n748_2[1]),.dout(n870),.clk(gclk));
	jor g0570(.dina(w_n765_4[0]),.dinb(w_n481_0[0]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n753_6[0]),.dinb(w_dff_B_QJsdoiVI0_1),.dout(n872),.clk(gclk));
	jnot g0572(.din(n872),.dout(n873),.clk(gclk));
	jand g0573(.dina(w_dff_B_wCO12kb00_0),.dinb(n871),.dout(n874),.clk(gclk));
	jand g0574(.dina(w_dff_B_fZP1RiSL2_0),.dinb(n870),.dout(G873_fa_),.clk(gclk));
	jand g0575(.dina(w_n567_0[2]),.dinb(w_G4_0[2]),.dout(n876),.clk(gclk));
	jnot g0576(.din(n876),.dout(n877),.clk(gclk));
	jand g0577(.dina(w_n877_0[1]),.dinb(w_n681_2[0]),.dout(n878),.clk(gclk));
	jor g0578(.dina(n878),.dinb(w_n571_0[2]),.dout(n879),.clk(gclk));
	jand g0579(.dina(w_n879_0[1]),.dinb(w_n687_0[1]),.dout(n880),.clk(gclk));
	jxor g0580(.dina(n880),.dinb(w_n583_0[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n881_0[1]),.dinb(w_n747_3[0]),.dout(n882),.clk(gclk));
	jnot g0582(.din(n882),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_n765_3[2]),.dinb(w_n459_0[0]),.dout(n884),.clk(gclk));
	jand g0584(.dina(w_n753_5[2]),.dinb(w_dff_B_A0F7fsOW6_1),.dout(n885),.clk(gclk));
	jnot g0585(.din(n885),.dout(n886),.clk(gclk));
	jand g0586(.dina(w_dff_B_Y8q27l6j4_0),.dinb(n884),.dout(n887),.clk(gclk));
	jand g0587(.dina(w_dff_B_UWRP0Y5A5_0),.dinb(n883),.dout(G875_fa_),.clk(gclk));
	jand g0588(.dina(w_n571_0[1]),.dinb(w_n681_1[2]),.dout(n889),.clk(gclk));
	jand g0589(.dina(w_dff_B_90uOtjj17_0),.dinb(w_n877_0[0]),.dout(n890),.clk(gclk));
	jnot g0590(.din(n890),.dout(n891),.clk(gclk));
	jand g0591(.dina(n891),.dinb(w_n879_0[0]),.dout(n892),.clk(gclk));
	jand g0592(.dina(w_n892_0[1]),.dinb(w_n747_2[2]),.dout(n893),.clk(gclk));
	jnot g0593(.din(n893),.dout(n894),.clk(gclk));
	jor g0594(.dina(w_n765_3[1]),.dinb(w_n494_0[0]),.dout(n895),.clk(gclk));
	jand g0595(.dina(w_n753_5[1]),.dinb(w_dff_B_mEvSGX876_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jand g0597(.dina(w_dff_B_WEhjN6ji8_0),.dinb(n895),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_dff_B_i7cpOCT88_0),.dinb(n894),.dout(G877_fa_),.clk(gclk));
	jxor g0599(.dina(w_n649_0[2]),.dinb(w_n735_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_n786_0[0]),.dout(n901),.clk(gclk));
	jxor g0601(.dina(n901),.dinb(w_n621_1[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_G369_0[0]),.dinb(w_n609_1[2]),.dout(n903),.clk(gclk));
	jand g0603(.dina(G372),.dinb(w_G332_1[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(w_dff_B_jyM7J1ZV9_0),.dinb(n903),.dout(n905),.clk(gclk));
	jxor g0605(.dina(n905),.dinb(w_n617_0[1]),.dout(n906),.clk(gclk));
	jxor g0606(.dina(n906),.dinb(w_n628_0[1]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_G331_0[0]),.dout(n908),.clk(gclk));
	jand g0608(.dina(w_n624_0[2]),.dinb(w_dff_B_zQ4MytPc7_1),.dout(n909),.clk(gclk));
	jnot g0609(.din(w_n624_0[1]),.dout(n910),.clk(gclk));
	jand g0610(.dina(w_dff_B_ZG2jwuz38_0),.dinb(w_n613_0[0]),.dout(n911),.clk(gclk));
	jor g0611(.dina(n911),.dinb(w_dff_B_JEPeCu9J0_1),.dout(n912),.clk(gclk));
	jxor g0612(.dina(n912),.dinb(w_dff_B_FhiAzXBB6_1),.dout(n913),.clk(gclk));
	jxor g0613(.dina(n913),.dinb(n902),.dout(n914),.clk(gclk));
	jnot g0614(.din(w_n914_0[1]),.dout(w_dff_A_rsHUFwPC0_1),.clk(gclk));
	jxor g0615(.dina(w_n577_0[0]),.dinb(w_n566_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n582_0[1]),.dinb(w_n570_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_n590_0[1]),.dout(n919),.clk(gclk));
	jand g0619(.dina(w_n556_1[2]),.dinb(w_G289_0[0]),.dout(n920),.clk(gclk));
	jand g0620(.dina(w_G335_1[1]),.dinb(G292),.dout(n921),.clk(gclk));
	jor g0621(.dina(w_dff_B_MvjSQb1U2_0),.dinb(n920),.dout(n922),.clk(gclk));
	jxor g0622(.dina(n922),.dinb(w_n600_0[2]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(n923),.dinb(w_n560_0[1]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n604_0[0]),.dinb(w_n595_0[1]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jxor g0626(.dina(n926),.dinb(n919),.dout(G1000_fa_),.clk(gclk));
	jnot g0627(.din(w_n596_0[1]),.dout(n928),.clk(gclk));
	jnot g0628(.din(w_n707_0[1]),.dout(n929),.clk(gclk));
	jnot g0629(.din(w_n700_0[0]),.dout(n930),.clk(gclk));
	jnot g0630(.din(w_n605_2[0]),.dout(n931),.clk(gclk));
	jnot g0631(.din(w_n601_0[0]),.dout(n932),.clk(gclk));
	jnot g0632(.din(w_n696_0[1]),.dout(n933),.clk(gclk));
	jand g0633(.dina(w_n587_1[0]),.dinb(w_G4_0[1]),.dout(n934),.clk(gclk));
	jnot g0634(.din(n934),.dout(n935),.clk(gclk));
	jand g0635(.dina(w_dff_B_yZEvMHkQ1_0),.dinb(n933),.dout(n936),.clk(gclk));
	jor g0636(.dina(w_n936_0[2]),.dinb(w_n932_0[1]),.dout(n937),.clk(gclk));
	jor g0637(.dina(n937),.dinb(w_dff_B_PSye6bXg7_1),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n938_0[1]),.dinb(w_n930_0[2]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_dff_B_TG5KVz8b0_1),.dout(n940),.clk(gclk));
	jxor g0640(.dina(n940),.dinb(w_n928_0[1]),.dout(n941),.clk(gclk));
	jnot g0641(.din(w_n941_0[1]),.dout(n942),.clk(gclk));
	jnot g0642(.din(w_n591_0[0]),.dout(n943),.clk(gclk));
	jnot g0643(.din(w_n705_0[0]),.dout(n944),.clk(gclk));
	jand g0644(.dina(w_n938_0[0]),.dinb(w_n944_0[1]),.dout(n945),.clk(gclk));
	jxor g0645(.dina(n945),.dinb(w_n943_0[1]),.dout(n946),.clk(gclk));
	jnot g0646(.din(w_n946_0[1]),.dout(n947),.clk(gclk));
	jor g0647(.dina(w_n600_0[1]),.dinb(w_G422_1[0]),.dout(n948),.clk(gclk));
	jnot g0648(.din(w_n948_0[2]),.dout(n949),.clk(gclk));
	jnot g0649(.din(w_n703_0[1]),.dout(n950),.clk(gclk));
	jand g0650(.dina(w_n936_0[1]),.dinb(w_dff_B_e5HQDqVp5_1),.dout(n951),.clk(gclk));
	jor g0651(.dina(n951),.dinb(w_dff_B_TffRr9w90_1),.dout(n952),.clk(gclk));
	jxor g0652(.dina(n952),.dinb(w_n605_1[2]),.dout(n953),.clk(gclk));
	jxor g0653(.dina(w_n936_0[0]),.dinb(w_n932_0[0]),.dout(n954),.clk(gclk));
	jnot g0654(.din(w_n954_0[1]),.dout(n955),.clk(gclk));
	jnot g0655(.din(w_n881_0[0]),.dout(n956),.clk(gclk));
	jnot g0656(.din(w_n771_0[0]),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n892_0[0]),.dout(n958),.clk(gclk));
	jand g0658(.dina(n958),.dinb(w_dff_B_3wJGaPeF1_1),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(n956),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n869_0[0]),.dout(n961),.clk(gclk));
	jand g0661(.dina(w_dff_B_KaCYtSDu2_0),.dinb(w_n862_0[0]),.dout(n962),.clk(gclk));
	jand g0662(.dina(w_dff_B_W2wYqFAe1_0),.dinb(n955),.dout(n963),.clk(gclk));
	jand g0663(.dina(n963),.dinb(w_n953_0[1]),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_dff_B_bXABOWnN9_0),.dinb(n947),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(n942),.dout(w_dff_A_ZwVSUgu01_2),.clk(gclk));
	jnot g0666(.din(w_n646_0[1]),.dout(n967),.clk(gclk));
	jor g0667(.dina(w_n649_0[1]),.dinb(w_G490_0[1]),.dout(n968),.clk(gclk));
	jor g0668(.dina(w_n781_0[1]),.dinb(w_n739_1[0]),.dout(n969),.clk(gclk));
	jand g0669(.dina(n969),.dinb(w_n968_0[1]),.dout(n970),.clk(gclk));
	jxor g0670(.dina(n970),.dinb(w_dff_B_udGqIPxm7_1),.dout(n971),.clk(gclk));
	jxor g0671(.dina(w_n783_0[2]),.dinb(w_n640_1[0]),.dout(n972),.clk(gclk));
	jxor g0672(.dina(w_n781_0[0]),.dinb(w_n650_0[0]),.dout(n973),.clk(gclk));
	jnot g0673(.din(w_n973_0[1]),.dout(n974),.clk(gclk));
	jor g0674(.dina(w_n621_0[2]),.dinb(w_n744_0[1]),.dout(n975),.clk(gclk));
	jand g0675(.dina(n975),.dinb(w_n636_0[2]),.dout(n976),.clk(gclk));
	jand g0676(.dina(w_dff_B_DEajMSUz6_0),.dinb(w_n761_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_dff_B_wAe7Cz920_0),.dinb(w_n832_0[0]),.dout(n978),.clk(gclk));
	jand g0678(.dina(w_dff_B_tjDkCpYo4_0),.dinb(w_n821_0[0]),.dout(n979),.clk(gclk));
	jand g0679(.dina(w_dff_B_mAUt7xJU8_0),.dinb(w_n809_0[0]),.dout(n980),.clk(gclk));
	jand g0680(.dina(w_dff_B_mSFnHuVU1_0),.dinb(n974),.dout(n981),.clk(gclk));
	jand g0681(.dina(n981),.dinb(w_n972_0[1]),.dout(n982),.clk(gclk));
	jand g0682(.dina(n982),.dinb(w_n971_0[1]),.dout(w_dff_A_aPAHZ5LL4_2),.clk(gclk));
	jnot g0683(.din(w_G1690_0[2]),.dout(n984),.clk(gclk));
	jand g0684(.dina(w_n984_0[1]),.dinb(w_G1689_0[2]),.dout(n985),.clk(gclk));
	jand g0685(.dina(w_n985_4[1]),.dinb(w_n791_0[2]),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_G1689_0[1]),.dout(n987),.clk(gclk));
	jand g0687(.dina(w_n984_0[0]),.dinb(w_n987_0[1]),.dout(n988),.clk(gclk));
	jand g0688(.dina(w_n988_4[1]),.dinb(w_n795_0[2]),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_G1690_0[1]),.dinb(w_n987_0[0]),.dout(n990),.clk(gclk));
	jand g0690(.dina(w_n990_4[1]),.dinb(w_G182_0[1]),.dout(n991),.clk(gclk));
	jand g0691(.dina(w_G1690_0[0]),.dinb(w_G1689_0[0]),.dout(n992),.clk(gclk));
	jand g0692(.dina(w_n992_4[1]),.dinb(w_G185_0[1]),.dout(n993),.clk(gclk));
	jor g0693(.dina(w_dff_B_yzSYTJWf6_0),.dinb(n991),.dout(n994),.clk(gclk));
	jor g0694(.dina(w_dff_B_8OjgUUdK4_0),.dinb(n989),.dout(n995),.clk(gclk));
	jor g0695(.dina(n995),.dinb(n986),.dout(n996),.clk(gclk));
	jand g0696(.dina(n996),.dinb(w_G137_9[1]),.dout(w_dff_A_BjvcmaIf8_2),.clk(gclk));
	jnot g0697(.din(w_G1694_0[2]),.dout(n998),.clk(gclk));
	jand g0698(.dina(w_n998_0[1]),.dinb(w_G1691_0[2]),.dout(n999),.clk(gclk));
	jand g0699(.dina(w_n999_4[1]),.dinb(w_n791_0[1]),.dout(n1000),.clk(gclk));
	jnot g0700(.din(w_G1691_0[1]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_n998_0[0]),.dinb(w_n1001_0[1]),.dout(n1002),.clk(gclk));
	jand g0702(.dina(w_n1002_4[1]),.dinb(w_n795_0[1]),.dout(n1003),.clk(gclk));
	jand g0703(.dina(w_G1694_0[1]),.dinb(w_n1001_0[0]),.dout(n1004),.clk(gclk));
	jand g0704(.dina(w_n1004_4[1]),.dinb(w_G182_0[0]),.dout(n1005),.clk(gclk));
	jand g0705(.dina(w_G1694_0[0]),.dinb(w_G1691_0[0]),.dout(n1006),.clk(gclk));
	jand g0706(.dina(w_n1006_4[1]),.dinb(w_G185_0[0]),.dout(n1007),.clk(gclk));
	jor g0707(.dina(w_dff_B_6TjWitqE6_0),.dinb(n1005),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_dff_B_avY0gwYw0_0),.dinb(n1003),.dout(n1009),.clk(gclk));
	jor g0709(.dina(n1009),.dinb(n1000),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_G137_9[0]),.dout(w_dff_A_T2PMMgd24_2),.clk(gclk));
	jnot g0711(.din(w_G871_0),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_1[1]),.dinb(w_n793_4[0]),.dout(n1013),.clk(gclk));
	jnot g0713(.din(w_G832_0),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_1[1]),.dinb(w_n797_4[0]),.dout(n1015),.clk(gclk));
	jand g0715(.dina(w_n799_4[0]),.dinb(w_G43_0[1]),.dout(n1016),.clk(gclk));
	jand g0716(.dina(w_n801_4[0]),.dinb(w_G37_0[1]),.dout(n1017),.clk(gclk));
	jor g0717(.dina(w_dff_B_Ww6v3SSi1_0),.dinb(n1016),.dout(n1018),.clk(gclk));
	jor g0718(.dina(w_dff_B_ztWLRg0X4_0),.dinb(n1015),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_dff_B_47TbZlIf2_0),.dinb(n1013),.dout(w_dff_A_xNgk3bJf2_2),.clk(gclk));
	jnot g0720(.din(w_G873_0),.dout(n1021),.clk(gclk));
	jand g0721(.dina(w_n1021_1[1]),.dinb(w_n793_3[2]),.dout(n1022),.clk(gclk));
	jnot g0722(.din(w_G834_0),.dout(n1023),.clk(gclk));
	jand g0723(.dina(w_n1023_1[1]),.dinb(w_n797_3[2]),.dout(n1024),.clk(gclk));
	jand g0724(.dina(w_n799_3[2]),.dinb(w_G76_0[1]),.dout(n1025),.clk(gclk));
	jand g0725(.dina(w_n801_3[2]),.dinb(w_G20_0[1]),.dout(n1026),.clk(gclk));
	jor g0726(.dina(w_dff_B_jHgqreCB4_0),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0727(.dina(w_dff_B_gz8CIbCF7_0),.dinb(n1024),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_4QTYj42L0_0),.dinb(n1022),.dout(w_dff_A_g0IwlMxo1_2),.clk(gclk));
	jnot g0729(.din(w_G875_0),.dout(n1030),.clk(gclk));
	jand g0730(.dina(w_n1030_1[1]),.dinb(w_n793_3[1]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G836_0),.dout(n1032),.clk(gclk));
	jand g0732(.dina(w_n1032_1[1]),.dinb(w_n797_3[1]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(w_n799_3[1]),.dinb(w_G73_0[1]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(w_n801_3[1]),.dinb(w_G17_0[1]),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_dff_B_gOnz1Z622_0),.dinb(n1034),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_dff_B_45NXoFSz2_0),.dinb(n1033),.dout(n1037),.clk(gclk));
	jor g0737(.dina(w_dff_B_syxrlt572_0),.dinb(n1031),.dout(w_dff_A_m9mvQOBB9_2),.clk(gclk));
	jnot g0738(.din(w_G877_0),.dout(n1039),.clk(gclk));
	jand g0739(.dina(w_n1039_1[1]),.dinb(w_n793_3[0]),.dout(n1040),.clk(gclk));
	jnot g0740(.din(w_G838_0),.dout(n1041),.clk(gclk));
	jand g0741(.dina(w_n797_3[0]),.dinb(w_n1041_1[1]),.dout(n1042),.clk(gclk));
	jand g0742(.dina(w_n799_3[0]),.dinb(w_G67_0[1]),.dout(n1043),.clk(gclk));
	jand g0743(.dina(w_n801_3[0]),.dinb(w_G70_0[1]),.dout(n1044),.clk(gclk));
	jor g0744(.dina(w_dff_B_04HM0IyZ8_0),.dinb(n1043),.dout(n1045),.clk(gclk));
	jor g0745(.dina(w_dff_B_zRMVweWr4_0),.dinb(n1042),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_dff_B_fvPzOQNK9_0),.dinb(n1040),.dout(w_dff_A_V5IgNeJF5_2),.clk(gclk));
	jand g0747(.dina(w_n1012_1[0]),.dinb(w_n840_4[0]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(w_n843_4[0]),.dinb(w_n1014_1[0]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(w_n845_4[0]),.dinb(w_G43_0[0]),.dout(n1050),.clk(gclk));
	jand g0750(.dina(w_n847_4[0]),.dinb(w_G37_0[0]),.dout(n1051),.clk(gclk));
	jor g0751(.dina(w_dff_B_JUusCXk67_0),.dinb(n1050),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_dff_B_IqO4jrNW8_0),.dinb(n1049),.dout(n1053),.clk(gclk));
	jor g0753(.dina(w_dff_B_lpijphA11_0),.dinb(n1048),.dout(w_dff_A_cPQHNv5B9_2),.clk(gclk));
	jand g0754(.dina(w_n1021_1[0]),.dinb(w_n840_3[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(w_n843_3[2]),.dinb(w_n1023_1[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(w_n845_3[2]),.dinb(w_G76_0[0]),.dout(n1057),.clk(gclk));
	jand g0757(.dina(w_n847_3[2]),.dinb(w_G20_0[0]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_dff_B_bMwGzXBW6_0),.dinb(n1057),.dout(n1059),.clk(gclk));
	jor g0759(.dina(w_dff_B_e9AgWHTM3_0),.dinb(n1056),.dout(n1060),.clk(gclk));
	jor g0760(.dina(w_dff_B_tm7n7pgN3_0),.dinb(n1055),.dout(w_dff_A_oRgwlr2S2_2),.clk(gclk));
	jand g0761(.dina(w_n1030_1[0]),.dinb(w_n840_3[1]),.dout(n1062),.clk(gclk));
	jand g0762(.dina(w_n843_3[1]),.dinb(w_n1032_1[0]),.dout(n1063),.clk(gclk));
	jand g0763(.dina(w_n845_3[1]),.dinb(w_G73_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(w_n847_3[1]),.dinb(w_G17_0[0]),.dout(n1065),.clk(gclk));
	jor g0765(.dina(w_dff_B_NwksgsXy5_0),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_dff_B_TKf1DxH57_0),.dinb(n1063),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_dff_B_TErgr8ko2_0),.dinb(n1062),.dout(w_dff_A_7sYsf6TN1_2),.clk(gclk));
	jand g0768(.dina(w_n1039_1[0]),.dinb(w_n840_3[0]),.dout(n1069),.clk(gclk));
	jand g0769(.dina(w_n843_3[0]),.dinb(w_n1041_1[0]),.dout(n1070),.clk(gclk));
	jand g0770(.dina(w_n845_3[0]),.dinb(w_G67_0[0]),.dout(n1071),.clk(gclk));
	jand g0771(.dina(w_n847_3[0]),.dinb(w_G70_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_dff_B_TZ3jdvfl1_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0773(.dina(w_dff_B_QKeZNlHr6_0),.dinb(n1070),.dout(n1074),.clk(gclk));
	jor g0774(.dina(w_dff_B_J3jcYmM34_0),.dinb(n1069),.dout(w_dff_A_axuI5cBD5_2),.clk(gclk));
	jand g0775(.dina(w_n985_4[0]),.dinb(w_n1012_0[2]),.dout(n1076),.clk(gclk));
	jand g0776(.dina(w_n988_4[0]),.dinb(w_n1014_0[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_n990_4[0]),.dinb(w_G200_0[1]),.dout(n1078),.clk(gclk));
	jand g0778(.dina(w_n992_4[0]),.dinb(w_G170_0[1]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(w_dff_B_WjCWHaAT4_0),.dinb(n1078),.dout(n1080),.clk(gclk));
	jor g0780(.dina(w_dff_B_W3ZZw4Cn9_0),.dinb(n1077),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_dff_B_XTnXtpgM8_0),.dinb(n1076),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G137_8[2]),.dout(w_dff_A_6rpt8BSf5_2),.clk(gclk));
	jand g0783(.dina(w_n985_3[2]),.dinb(w_n1039_0[2]),.dout(n1084),.clk(gclk));
	jand g0784(.dina(w_n988_3[2]),.dinb(w_n1041_0[2]),.dout(n1085),.clk(gclk));
	jand g0785(.dina(w_n990_3[2]),.dinb(w_G188_0[1]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(w_n992_3[2]),.dinb(w_G158_0[1]),.dout(n1087),.clk(gclk));
	jor g0787(.dina(w_dff_B_UroukBto2_0),.dinb(n1086),.dout(n1088),.clk(gclk));
	jor g0788(.dina(w_dff_B_W18ARSSY5_0),.dinb(n1085),.dout(n1089),.clk(gclk));
	jor g0789(.dina(w_dff_B_T3z170Uf8_0),.dinb(n1084),.dout(n1090),.clk(gclk));
	jand g0790(.dina(n1090),.dinb(w_G137_8[1]),.dout(w_dff_A_8re8Z0rV0_2),.clk(gclk));
	jand g0791(.dina(w_n985_3[1]),.dinb(w_n1030_0[2]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(w_n988_3[1]),.dinb(w_n1032_0[2]),.dout(n1093),.clk(gclk));
	jand g0793(.dina(w_n990_3[1]),.dinb(w_G155_0[1]),.dout(n1094),.clk(gclk));
	jand g0794(.dina(w_n992_3[1]),.dinb(w_G152_0[1]),.dout(n1095),.clk(gclk));
	jor g0795(.dina(w_dff_B_0aRS2stc2_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jor g0796(.dina(w_dff_B_D7JximM67_0),.dinb(n1093),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_KlIGP9566_0),.dinb(n1092),.dout(n1098),.clk(gclk));
	jand g0798(.dina(n1098),.dinb(w_G137_8[0]),.dout(w_dff_A_3hWNAct47_2),.clk(gclk));
	jand g0799(.dina(w_n985_3[0]),.dinb(w_n1021_0[2]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(w_n988_3[0]),.dinb(w_n1023_0[2]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(w_n990_3[0]),.dinb(w_G149_0[1]),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n992_3[0]),.dinb(w_G146_0[1]),.dout(n1103),.clk(gclk));
	jor g0803(.dina(w_dff_B_xkoqWe9W8_0),.dinb(n1102),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_5qbHPi520_0),.dinb(n1101),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_BprNyinQ4_0),.dinb(n1100),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_7[2]),.dout(w_dff_A_BCHA1aqF8_2),.clk(gclk));
	jand g0807(.dina(w_n999_4[0]),.dinb(w_n1012_0[1]),.dout(n1108),.clk(gclk));
	jand g0808(.dina(w_n1002_4[0]),.dinb(w_n1014_0[1]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(w_n1004_4[0]),.dinb(w_G200_0[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_n1006_4[0]),.dinb(w_G170_0[0]),.dout(n1111),.clk(gclk));
	jor g0811(.dina(w_dff_B_5KDeyqNZ2_0),.dinb(n1110),.dout(n1112),.clk(gclk));
	jor g0812(.dina(w_dff_B_GzcXBlx84_0),.dinb(n1109),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_OgIeoO6B4_0),.dinb(n1108),.dout(n1114),.clk(gclk));
	jand g0814(.dina(n1114),.dinb(w_G137_7[1]),.dout(w_dff_A_Dt6jwWtM8_2),.clk(gclk));
	jand g0815(.dina(w_n999_3[2]),.dinb(w_n1039_0[1]),.dout(n1116),.clk(gclk));
	jand g0816(.dina(w_n1002_3[2]),.dinb(w_n1041_0[1]),.dout(n1117),.clk(gclk));
	jand g0817(.dina(w_n1004_3[2]),.dinb(w_G188_0[0]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(w_n1006_3[2]),.dinb(w_G158_0[0]),.dout(n1119),.clk(gclk));
	jor g0819(.dina(w_dff_B_Dria40VK9_0),.dinb(n1118),.dout(n1120),.clk(gclk));
	jor g0820(.dina(w_dff_B_wahLog2R8_0),.dinb(n1117),.dout(n1121),.clk(gclk));
	jor g0821(.dina(w_dff_B_CNjIMwUF5_0),.dinb(n1116),.dout(n1122),.clk(gclk));
	jand g0822(.dina(n1122),.dinb(w_G137_7[0]),.dout(w_dff_A_MqQBwMxU9_2),.clk(gclk));
	jand g0823(.dina(w_n999_3[1]),.dinb(w_n1030_0[1]),.dout(n1124),.clk(gclk));
	jand g0824(.dina(w_n1002_3[1]),.dinb(w_n1032_0[1]),.dout(n1125),.clk(gclk));
	jand g0825(.dina(w_n1004_3[1]),.dinb(w_G155_0[0]),.dout(n1126),.clk(gclk));
	jand g0826(.dina(w_n1006_3[1]),.dinb(w_G152_0[0]),.dout(n1127),.clk(gclk));
	jor g0827(.dina(w_dff_B_htxaFz5i3_0),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g0828(.dina(w_dff_B_q1U8qdc83_0),.dinb(n1125),.dout(n1129),.clk(gclk));
	jor g0829(.dina(w_dff_B_reDfHA2s8_0),.dinb(n1124),.dout(n1130),.clk(gclk));
	jand g0830(.dina(n1130),.dinb(w_G137_6[2]),.dout(w_dff_A_AX6UZEQe8_2),.clk(gclk));
	jand g0831(.dina(w_n999_3[0]),.dinb(w_n1021_0[1]),.dout(n1132),.clk(gclk));
	jand g0832(.dina(w_n1002_3[0]),.dinb(w_n1023_0[1]),.dout(n1133),.clk(gclk));
	jand g0833(.dina(w_n1004_3[0]),.dinb(w_G149_0[0]),.dout(n1134),.clk(gclk));
	jand g0834(.dina(w_n1006_3[0]),.dinb(w_G146_0[0]),.dout(n1135),.clk(gclk));
	jor g0835(.dina(w_dff_B_1vcrToXD2_0),.dinb(n1134),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_dff_B_tntgAJsr9_0),.dinb(n1133),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_dff_B_ZNFHKvU31_0),.dinb(n1132),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(w_G137_6[1]),.dout(w_dff_A_pI4UzbjX7_2),.clk(gclk));
	jand g0839(.dina(w_n789_0[1]),.dinb(w_G3724_0[2]),.dout(n1140),.clk(gclk));
	jnot g0840(.din(w_G3717_0[1]),.dout(n1141),.clk(gclk));
	jnot g0841(.din(w_G3724_0[1]),.dout(n1142),.clk(gclk));
	jand g0842(.dina(w_n1142_0[1]),.dinb(w_G123_0[1]),.dout(n1143),.clk(gclk));
	jor g0843(.dina(n1143),.dinb(w_dff_B_J0YdLulo1_1),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_dff_B_FMrwp04V2_0),.dinb(n1140),.dout(n1145),.clk(gclk));
	jnot g0845(.din(G135),.dout(n1146),.clk(gclk));
	jnot g0846(.din(G4115),.dout(n1147),.clk(gclk));
	jor g0847(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jxor g0848(.dina(w_n636_0[1]),.dinb(w_G132_0[1]),.dout(n1149),.clk(gclk));
	jand g0849(.dina(n1149),.dinb(w_G3724_0[0]),.dout(n1150),.clk(gclk));
	jnot g0850(.din(w_n401_0[1]),.dout(n1151),.clk(gclk));
	jand g0851(.dina(w_n1151_0[1]),.dinb(w_n1142_0[0]),.dout(n1152),.clk(gclk));
	jor g0852(.dina(n1152),.dinb(w_G3717_0[0]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(n1153),.dinb(w_dff_B_n1caYDXs8_1),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_dff_B_FsbrXkvc7_1),.dout(n1155),.clk(gclk));
	jand g0855(.dina(w_dff_B_w7QhIpOV3_0),.dinb(n1145),.dout(w_dff_A_PL0nReCd3_2),.clk(gclk));
	jor g0856(.dina(w_n783_0[1]),.dinb(w_n640_0[2]),.dout(n1157),.clk(gclk));
	jxor g0857(.dina(n1157),.dinb(w_G132_0[0]),.dout(w_dff_A_wjwk8NfH6_2),.clk(gclk));
	jand g0858(.dina(w_n789_0[0]),.dinb(w_n747_2[1]),.dout(n1159),.clk(gclk));
	jand g0859(.dina(w_n753_5[0]),.dinb(w_G123_0[0]),.dout(n1160),.clk(gclk));
	jand g0860(.dina(w_n751_1[1]),.dinb(w_n1151_0[0]),.dout(n1161),.clk(gclk));
	jor g0861(.dina(n1161),.dinb(w_dff_B_FE6uwSmS0_1),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_dff_B_BWNbPEii0_0),.dinb(n1159),.dout(n1163),.clk(gclk));
	jnot g0863(.din(w_n1163_1[2]),.dout(w_dff_A_H9l19U0M7_1),.clk(gclk));
	jor g0864(.dina(w_n972_0[0]),.dinb(w_n748_2[0]),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n751_1[0]),.dinb(w_n407_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n753_4[2]),.dinb(w_dff_B_uKr8CYGs6_1),.dout(n1167),.clk(gclk));
	jor g0867(.dina(w_dff_B_marBBmw55_0),.dinb(n1166),.dout(n1168),.clk(gclk));
	jnot g0868(.din(n1168),.dout(n1169),.clk(gclk));
	jand g0869(.dina(w_dff_B_KrP1yuHQ9_0),.dinb(n1165),.dout(G826_fa_),.clk(gclk));
	jor g0870(.dina(w_n971_0[0]),.dinb(w_n748_1[2]),.dout(n1171),.clk(gclk));
	jor g0871(.dina(w_n765_3[0]),.dinb(w_n372_0[1]),.dout(n1172),.clk(gclk));
	jand g0872(.dina(w_n753_4[1]),.dinb(w_dff_B_h2p3nyxB3_1),.dout(n1173),.clk(gclk));
	jnot g0873(.din(n1173),.dout(n1174),.clk(gclk));
	jand g0874(.dina(w_dff_B_1QghGSTZ5_0),.dinb(n1172),.dout(n1175),.clk(gclk));
	jand g0875(.dina(w_dff_B_vJHcfLve3_0),.dinb(n1171),.dout(G828_fa_),.clk(gclk));
	jand g0876(.dina(w_n973_0[0]),.dinb(w_n747_2[0]),.dout(n1177),.clk(gclk));
	jnot g0877(.din(n1177),.dout(n1178),.clk(gclk));
	jor g0878(.dina(w_n765_2[2]),.dinb(w_n383_0[1]),.dout(n1179),.clk(gclk));
	jand g0879(.dina(w_n753_4[0]),.dinb(w_dff_B_tYfQVzEI9_1),.dout(n1180),.clk(gclk));
	jnot g0880(.din(n1180),.dout(n1181),.clk(gclk));
	jand g0881(.dina(w_dff_B_62huH6Nq1_0),.dinb(n1179),.dout(n1182),.clk(gclk));
	jand g0882(.dina(w_dff_B_AQUBKamq2_0),.dinb(n1178),.dout(G830_fa_),.clk(gclk));
	jnot g0883(.din(w_G1000_0),.dout(n1184),.clk(gclk));
	jand g0884(.dina(w_G559_0[0]),.dinb(w_G245_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(n1185),.dinb(w_n318_0[0]),.dout(n1186),.clk(gclk));
	jand g0886(.dina(n1186),.dinb(w_G601_0),.dout(n1187),.clk(gclk));
	jand g0887(.dina(w_dff_B_NHXjAi4F9_0),.dinb(w_n661_0[0]),.dout(n1188),.clk(gclk));
	jand g0888(.dina(n1188),.dinb(w_n671_0[0]),.dout(n1189),.clk(gclk));
	jand g0889(.dina(w_dff_B_Fk7TrJzz6_0),.dinb(w_n914_0[0]),.dout(n1190),.clk(gclk));
	jand g0890(.dina(n1190),.dinb(w_dff_B_9S8cjbQD0_1),.dout(w_dff_A_kppvDxAs8_2),.clk(gclk));
	jand g0891(.dina(w_n941_0[0]),.dinb(w_n747_1[2]),.dout(n1192),.clk(gclk));
	jnot g0892(.din(w_n528_0[1]),.dout(n1193),.clk(gclk));
	jand g0893(.dina(w_n751_0[2]),.dinb(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_n753_3[2]),.dinb(w_dff_B_9G85qHLp6_1),.dout(n1195),.clk(gclk));
	jor g0895(.dina(w_dff_B_20Y1p8ix0_0),.dinb(n1194),.dout(n1196),.clk(gclk));
	jor g0896(.dina(w_dff_B_5R5KWFjg0_0),.dinb(n1192),.dout(n1197),.clk(gclk));
	jnot g0897(.din(w_n1197_1[2]),.dout(w_dff_A_Db0Se1s10_1),.clk(gclk));
	jand g0898(.dina(w_n946_0[0]),.dinb(w_n747_1[1]),.dout(n1199),.clk(gclk));
	jor g0899(.dina(w_n765_2[1]),.dinb(w_n551_0[0]),.dout(n1200),.clk(gclk));
	jand g0900(.dina(w_n753_3[1]),.dinb(w_dff_B_vNPPy6ed3_1),.dout(n1201),.clk(gclk));
	jnot g0901(.din(n1201),.dout(n1202),.clk(gclk));
	jand g0902(.dina(w_dff_B_XGAPpf743_0),.dinb(n1200),.dout(n1203),.clk(gclk));
	jnot g0903(.din(n1203),.dout(n1204),.clk(gclk));
	jor g0904(.dina(w_dff_B_WPzhHrAb9_0),.dinb(n1199),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_Xvirj3x92_1),.clk(gclk));
	jor g0906(.dina(w_n953_0[0]),.dinb(w_n748_1[1]),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n765_2[0]),.dinb(w_n517_0[0]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n753_3[0]),.dinb(w_dff_B_StV1voEx0_1),.dout(n1209),.clk(gclk));
	jnot g0909(.din(n1209),.dout(n1210),.clk(gclk));
	jand g0910(.dina(w_dff_B_7PZywBut2_0),.dinb(n1208),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_xAXaJ5Ik2_0),.dinb(n1207),.dout(G867_fa_),.clk(gclk));
	jand g0912(.dina(w_n954_0[0]),.dinb(w_n747_1[0]),.dout(n1213),.clk(gclk));
	jnot g0913(.din(n1213),.dout(n1214),.clk(gclk));
	jor g0914(.dina(w_n765_1[2]),.dinb(w_n540_0[0]),.dout(n1215),.clk(gclk));
	jand g0915(.dina(w_n753_2[2]),.dinb(w_dff_B_AKDvo7Ba7_1),.dout(n1216),.clk(gclk));
	jnot g0916(.din(n1216),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_dff_B_kWzdq82a2_0),.dinb(n1215),.dout(n1218),.clk(gclk));
	jand g0918(.dina(w_dff_B_jGhB8Mmf3_0),.dinb(n1214),.dout(G869_fa_),.clk(gclk));
	jand g0919(.dina(w_n1197_1[1]),.dinb(w_n840_2[2]),.dout(n1220),.clk(gclk));
	jand g0920(.dina(w_n1163_1[1]),.dinb(w_n843_2[2]),.dout(n1221),.clk(gclk));
	jand g0921(.dina(w_n845_2[2]),.dinb(w_G109_0[1]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_n847_2[2]),.dinb(w_G106_0[1]),.dout(n1223),.clk(gclk));
	jor g0923(.dina(w_dff_B_2C2LaIa98_0),.dinb(n1222),.dout(n1224),.clk(gclk));
	jor g0924(.dina(w_dff_B_I2ermMkl7_0),.dinb(n1221),.dout(n1225),.clk(gclk));
	jor g0925(.dina(n1225),.dinb(n1220),.dout(w_dff_A_UTwmXiJV5_2),.clk(gclk));
	jand g0926(.dina(w_n1197_1[0]),.dinb(w_n793_2[2]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_n1163_1[0]),.dinb(w_n797_2[2]),.dout(n1228),.clk(gclk));
	jand g0928(.dina(w_n799_2[2]),.dinb(w_G109_0[0]),.dout(n1229),.clk(gclk));
	jand g0929(.dina(w_n801_2[2]),.dinb(w_G106_0[0]),.dout(n1230),.clk(gclk));
	jor g0930(.dina(w_dff_B_Ih13jZBk8_0),.dinb(n1229),.dout(n1231),.clk(gclk));
	jor g0931(.dina(w_dff_B_nsPRMNxz1_0),.dinb(n1228),.dout(n1232),.clk(gclk));
	jor g0932(.dina(n1232),.dinb(n1227),.dout(w_dff_A_cpxnTtkT7_2),.clk(gclk));
	jand g0933(.dina(w_n1205_1[1]),.dinb(w_n793_2[1]),.dout(n1234),.clk(gclk));
	jnot g0934(.din(w_G826_0),.dout(n1235),.clk(gclk));
	jand g0935(.dina(w_n1235_1[1]),.dinb(w_n797_2[1]),.dout(n1236),.clk(gclk));
	jand g0936(.dina(w_n799_2[1]),.dinb(w_G46_0[1]),.dout(n1237),.clk(gclk));
	jand g0937(.dina(w_n801_2[1]),.dinb(w_G49_0[1]),.dout(n1238),.clk(gclk));
	jor g0938(.dina(w_dff_B_bKng4ZYj7_0),.dinb(n1237),.dout(n1239),.clk(gclk));
	jor g0939(.dina(w_dff_B_wsrvTRFU1_0),.dinb(n1236),.dout(n1240),.clk(gclk));
	jor g0940(.dina(n1240),.dinb(n1234),.dout(w_dff_A_zT3XBVAo1_2),.clk(gclk));
	jnot g0941(.din(w_G867_0),.dout(n1242),.clk(gclk));
	jand g0942(.dina(w_n1242_1[1]),.dinb(w_n793_2[0]),.dout(n1243),.clk(gclk));
	jnot g0943(.din(w_G828_0),.dout(n1244),.clk(gclk));
	jand g0944(.dina(w_n1244_1[1]),.dinb(w_n797_2[0]),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n799_2[0]),.dinb(w_G100_0[1]),.dout(n1246),.clk(gclk));
	jand g0946(.dina(w_n801_2[0]),.dinb(w_G103_0[1]),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_dff_B_uwUSbe004_0),.dinb(n1246),.dout(n1248),.clk(gclk));
	jor g0948(.dina(w_dff_B_bOm6xuOr3_0),.dinb(n1245),.dout(n1249),.clk(gclk));
	jor g0949(.dina(n1249),.dinb(n1243),.dout(w_dff_A_8UD0c5Ru2_2),.clk(gclk));
	jnot g0950(.din(w_G869_0),.dout(n1251),.clk(gclk));
	jand g0951(.dina(w_n1251_1[1]),.dinb(w_n793_1[2]),.dout(n1252),.clk(gclk));
	jnot g0952(.din(w_G830_0),.dout(n1253),.clk(gclk));
	jand g0953(.dina(w_n1253_1[1]),.dinb(w_n797_1[2]),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n799_1[2]),.dinb(w_G91_0[1]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n801_1[2]),.dinb(w_G40_0[1]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(w_dff_B_5jWzyvJG7_0),.dinb(n1255),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_t94d85kX8_0),.dinb(n1254),.dout(n1258),.clk(gclk));
	jor g0958(.dina(n1258),.dinb(n1252),.dout(w_dff_A_PIldz9RX9_2),.clk(gclk));
	jand g0959(.dina(w_n1205_1[0]),.dinb(w_n840_2[1]),.dout(n1260),.clk(gclk));
	jand g0960(.dina(w_n1235_1[0]),.dinb(w_n843_2[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(w_n845_2[1]),.dinb(w_G46_0[0]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(w_n847_2[1]),.dinb(w_G49_0[0]),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_dff_B_Izl0K9OX4_0),.dinb(n1262),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_dff_B_LhUW3Ydi0_0),.dinb(n1261),.dout(n1265),.clk(gclk));
	jor g0965(.dina(n1265),.dinb(n1260),.dout(w_dff_A_zLFP5pWE0_2),.clk(gclk));
	jand g0966(.dina(w_n1242_1[0]),.dinb(w_n840_2[0]),.dout(n1267),.clk(gclk));
	jand g0967(.dina(w_n1244_1[0]),.dinb(w_n843_2[0]),.dout(n1268),.clk(gclk));
	jand g0968(.dina(w_n845_2[0]),.dinb(w_G100_0[0]),.dout(n1269),.clk(gclk));
	jand g0969(.dina(w_n847_2[0]),.dinb(w_G103_0[0]),.dout(n1270),.clk(gclk));
	jor g0970(.dina(w_dff_B_jlLPp9Vx4_0),.dinb(n1269),.dout(n1271),.clk(gclk));
	jor g0971(.dina(w_dff_B_aiw9eHOp9_0),.dinb(n1268),.dout(n1272),.clk(gclk));
	jor g0972(.dina(n1272),.dinb(n1267),.dout(w_dff_A_Jc6Rpzbn3_2),.clk(gclk));
	jand g0973(.dina(w_n1251_1[0]),.dinb(w_n840_1[2]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(w_n1253_1[0]),.dinb(w_n843_1[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(w_n845_1[2]),.dinb(w_G91_0[0]),.dout(n1276),.clk(gclk));
	jand g0976(.dina(w_n847_1[2]),.dinb(w_G40_0[0]),.dout(n1277),.clk(gclk));
	jor g0977(.dina(w_dff_B_vi4xFXql7_0),.dinb(n1276),.dout(n1278),.clk(gclk));
	jor g0978(.dina(w_dff_B_pcFZ3uXV4_0),.dinb(n1275),.dout(n1279),.clk(gclk));
	jor g0979(.dina(n1279),.dinb(n1274),.dout(w_dff_A_W3LY4oTh8_2),.clk(gclk));
	jand g0980(.dina(w_n1251_0[2]),.dinb(w_n985_2[2]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(w_n1253_0[2]),.dinb(w_n988_2[2]),.dout(n1282),.clk(gclk));
	jand g0982(.dina(w_n990_2[2]),.dinb(w_G203_0[1]),.dout(n1283),.clk(gclk));
	jand g0983(.dina(w_n992_2[2]),.dinb(w_G173_0[1]),.dout(n1284),.clk(gclk));
	jor g0984(.dina(w_dff_B_fis0PEsW9_0),.dinb(n1283),.dout(n1285),.clk(gclk));
	jor g0985(.dina(w_dff_B_bdxp7AcU3_0),.dinb(n1282),.dout(n1286),.clk(gclk));
	jor g0986(.dina(n1286),.dinb(n1281),.dout(n1287),.clk(gclk));
	jand g0987(.dina(n1287),.dinb(w_G137_6[0]),.dout(w_dff_A_FMg1FwX22_2),.clk(gclk));
	jand g0988(.dina(w_n1242_0[2]),.dinb(w_n985_2[1]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(w_n1244_0[2]),.dinb(w_n988_2[1]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(w_n990_2[1]),.dinb(w_G197_0[1]),.dout(n1291),.clk(gclk));
	jand g0991(.dina(w_n992_2[1]),.dinb(w_G167_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_dff_B_294IO92r3_0),.dinb(n1291),.dout(n1293),.clk(gclk));
	jor g0993(.dina(w_dff_B_V85onpWG4_0),.dinb(n1290),.dout(n1294),.clk(gclk));
	jor g0994(.dina(n1294),.dinb(n1289),.dout(n1295),.clk(gclk));
	jand g0995(.dina(n1295),.dinb(w_G137_5[2]),.dout(w_dff_A_1QlhlnXk4_2),.clk(gclk));
	jand g0996(.dina(w_n1205_0[2]),.dinb(w_n985_2[0]),.dout(n1297),.clk(gclk));
	jand g0997(.dina(w_n1235_0[2]),.dinb(w_n988_2[0]),.dout(n1298),.clk(gclk));
	jand g0998(.dina(w_n990_2[0]),.dinb(w_G194_0[1]),.dout(n1299),.clk(gclk));
	jand g0999(.dina(w_n992_2[0]),.dinb(w_G164_0[1]),.dout(n1300),.clk(gclk));
	jor g1000(.dina(w_dff_B_FfSLbWuY1_0),.dinb(n1299),.dout(n1301),.clk(gclk));
	jor g1001(.dina(w_dff_B_C1YjVtUI7_0),.dinb(n1298),.dout(n1302),.clk(gclk));
	jor g1002(.dina(n1302),.dinb(n1297),.dout(n1303),.clk(gclk));
	jand g1003(.dina(n1303),.dinb(w_G137_5[1]),.dout(w_dff_A_yqoRBsWS7_2),.clk(gclk));
	jand g1004(.dina(w_n1197_0[2]),.dinb(w_n985_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(w_n1163_0[2]),.dinb(w_n988_1[2]),.dout(n1306),.clk(gclk));
	jand g1006(.dina(w_n990_1[2]),.dinb(w_G191_0[1]),.dout(n1307),.clk(gclk));
	jand g1007(.dina(w_n992_1[2]),.dinb(w_G161_0[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_dff_B_KImXdIga2_0),.dinb(n1307),.dout(n1309),.clk(gclk));
	jor g1009(.dina(w_dff_B_UhZT5YK20_0),.dinb(n1306),.dout(n1310),.clk(gclk));
	jor g1010(.dina(n1310),.dinb(n1305),.dout(n1311),.clk(gclk));
	jand g1011(.dina(n1311),.dinb(w_G137_5[0]),.dout(w_dff_A_GDUy23aV8_2),.clk(gclk));
	jand g1012(.dina(w_n1251_0[1]),.dinb(w_n999_2[2]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(w_n1253_0[1]),.dinb(w_n1002_2[2]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(w_n1004_2[2]),.dinb(w_G203_0[0]),.dout(n1315),.clk(gclk));
	jand g1015(.dina(w_n1006_2[2]),.dinb(w_G173_0[0]),.dout(n1316),.clk(gclk));
	jor g1016(.dina(w_dff_B_OKMz4WVo9_0),.dinb(n1315),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_dff_B_ccTWhB2x9_0),.dinb(n1314),.dout(n1318),.clk(gclk));
	jor g1018(.dina(n1318),.dinb(n1313),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_G137_4[2]),.dout(w_dff_A_Koy1Jatt2_2),.clk(gclk));
	jand g1020(.dina(w_n1242_0[1]),.dinb(w_n999_2[1]),.dout(n1321),.clk(gclk));
	jand g1021(.dina(w_n1244_0[1]),.dinb(w_n1002_2[1]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(w_n1004_2[1]),.dinb(w_G197_0[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(w_n1006_2[1]),.dinb(w_G167_0[0]),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_SAWpM6fQ5_0),.dinb(n1323),.dout(n1325),.clk(gclk));
	jor g1025(.dina(w_dff_B_lXYnlb5b3_0),.dinb(n1322),.dout(n1326),.clk(gclk));
	jor g1026(.dina(n1326),.dinb(n1321),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_G137_4[1]),.dout(w_dff_A_pBwC6pVv9_2),.clk(gclk));
	jand g1028(.dina(w_n1205_0[1]),.dinb(w_n999_2[0]),.dout(n1329),.clk(gclk));
	jand g1029(.dina(w_n1235_0[1]),.dinb(w_n1002_2[0]),.dout(n1330),.clk(gclk));
	jand g1030(.dina(w_n1004_2[0]),.dinb(w_G194_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(w_n1006_2[0]),.dinb(w_G164_0[0]),.dout(n1332),.clk(gclk));
	jor g1032(.dina(w_dff_B_powhZxEO6_0),.dinb(n1331),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_RyyWYobz7_0),.dinb(n1330),.dout(n1334),.clk(gclk));
	jor g1034(.dina(n1334),.dinb(n1329),.dout(n1335),.clk(gclk));
	jand g1035(.dina(n1335),.dinb(w_G137_4[0]),.dout(w_dff_A_R1XS5Ihe0_2),.clk(gclk));
	jand g1036(.dina(w_n1197_0[1]),.dinb(w_n999_1[2]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(w_n1163_0[1]),.dinb(w_n1002_1[2]),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n1004_1[2]),.dinb(w_G191_0[0]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n1006_1[2]),.dinb(w_G161_0[0]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(w_dff_B_nXPPc2nM8_0),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_AM3vBMxa2_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jor g1042(.dina(n1342),.dinb(n1337),.dout(n1343),.clk(gclk));
	jand g1043(.dina(n1343),.dinb(w_G137_3[2]),.dout(w_dff_A_8T6yUygj4_2),.clk(gclk));
	jor g1044(.dina(w_G4091_2[0]),.dinb(G120),.dout(n1345),.clk(gclk));
	jand g1045(.dina(w_n435_0[2]),.dinb(w_G251_3[1]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1347),.clk(gclk));
	jor g1047(.dina(n1347),.dinb(w_n437_0[1]),.dout(n1348),.clk(gclk));
	jor g1048(.dina(n1348),.dinb(n1346),.dout(n1349),.clk(gclk));
	jand g1049(.dina(w_n435_0[1]),.dinb(w_n366_3[1]),.dout(n1350),.clk(gclk));
	jand g1050(.dina(w_G341_0[2]),.dinb(w_n368_4[0]),.dout(n1351),.clk(gclk));
	jor g1051(.dina(n1351),.dinb(w_G523_0[2]),.dout(n1352),.clk(gclk));
	jor g1052(.dina(n1352),.dinb(w_dff_B_nc06qPDF0_1),.dout(n1353),.clk(gclk));
	jand g1053(.dina(n1353),.dinb(w_dff_B_a2v8VoHg4_1),.dout(n1354),.clk(gclk));
	jxor g1054(.dina(w_n408_0[0]),.dinb(w_n401_0[0]),.dout(n1355),.clk(gclk));
	jxor g1055(.dina(w_n383_0[0]),.dinb(w_n372_0[0]),.dout(n1356),.clk(gclk));
	jxor g1056(.dina(n1356),.dinb(w_dff_B_lAeKIlEP8_1),.dout(n1357),.clk(gclk));
	jxor g1057(.dina(n1357),.dinb(w_dff_B_Ywm0ecfJ3_1),.dout(n1358),.clk(gclk));
	jnot g1058(.din(w_n1358_0[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(w_n410_0[1]),.dinb(w_G248_3[2]),.dout(n1360),.clk(gclk));
	jor g1060(.dina(w_G514_0[1]),.dinb(w_n368_3[2]),.dout(n1361),.clk(gclk));
	jand g1061(.dina(n1361),.dinb(n1360),.dout(n1362),.clk(gclk));
	jxor g1062(.dina(n1362),.dinb(w_n419_0[0]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_G351_1[0]),.dinb(w_n402_1[2]),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n385_0[2]),.dinb(w_n405_1[2]),.dout(n1365),.clk(gclk));
	jand g1065(.dina(n1365),.dinb(w_G534_0[1]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_aWUAzN4U2_1),.dout(n1367),.clk(gclk));
	jor g1067(.dina(w_G351_0[2]),.dinb(w_G254_1[1]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(w_n385_0[1]),.dinb(w_G242_1[1]),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_n388_0[1]),.dout(n1370),.clk(gclk));
	jand g1070(.dina(n1370),.dinb(w_dff_B_5XAEIhWx1_1),.dout(n1371),.clk(gclk));
	jor g1071(.dina(n1371),.dinb(n1367),.dout(n1372),.clk(gclk));
	jand g1072(.dina(w_n424_1[0]),.dinb(w_G251_3[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(w_G324_0[2]),.dinb(w_G248_3[1]),.dout(n1374),.clk(gclk));
	jor g1074(.dina(n1374),.dinb(w_n426_0[0]),.dout(n1375),.clk(gclk));
	jor g1075(.dina(n1375),.dinb(n1373),.dout(n1376),.clk(gclk));
	jand g1076(.dina(w_n424_0[2]),.dinb(w_n366_3[0]),.dout(n1377),.clk(gclk));
	jand g1077(.dina(w_G324_0[1]),.dinb(w_n368_3[1]),.dout(n1378),.clk(gclk));
	jor g1078(.dina(n1378),.dinb(w_G503_0[1]),.dout(n1379),.clk(gclk));
	jor g1079(.dina(n1379),.dinb(w_dff_B_kRJT3wse7_1),.dout(n1380),.clk(gclk));
	jand g1080(.dina(n1380),.dinb(w_dff_B_rhIZik0W9_1),.dout(n1381),.clk(gclk));
	jxor g1081(.dina(n1381),.dinb(n1372),.dout(n1382),.clk(gclk));
	jxor g1082(.dina(n1382),.dinb(w_dff_B_Cn27TpIJ0_1),.dout(n1383),.clk(gclk));
	jnot g1083(.din(w_n1383_0[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(w_n1383_0[0]),.dinb(n1359),.dout(n1385),.clk(gclk));
	jor g1085(.dina(n1385),.dinb(w_G4091_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1345),.dinb(w_n746_1[0]),.dout(n1388),.clk(gclk));
	jand g1087(.dina(n1384),.dinb(w_n1358_0[0]),.dout(n1389),.clk(gclk));
	jor g1088(.dina(n1386),.dinb(w_dff_B_fwDQ9fKU8_1),.dout(n1390),.clk(gclk));
	jand g1089(.dina(n1390),.dinb(w_n746_0[2]),.dout(n1391),.clk(gclk));
	jnot g1090(.din(w_n1391_0[1]),.dout(n1392),.clk(gclk));
	jand g1091(.dina(w_n633_0[2]),.dinb(w_G2174_0[2]),.dout(n1393),.clk(gclk));
	jor g1092(.dina(w_dff_B_bavSCnqv8_0),.dinb(w_n732_0[0]),.dout(n1394),.clk(gclk));
	jand g1093(.dina(w_n736_0[0]),.dinb(w_n640_0[1]),.dout(n1395),.clk(gclk));
	jor g1094(.dina(w_n740_0[0]),.dinb(w_n641_0[0]),.dout(n1396),.clk(gclk));
	jand g1095(.dina(n1396),.dinb(w_n646_0[0]),.dout(n1397),.clk(gclk));
	jor g1096(.dina(n1397),.dinb(w_dff_B_1KEajjX92_1),.dout(n1398),.clk(gclk));
	jnot g1097(.din(w_n1398_0[1]),.dout(n1399),.clk(gclk));
	jand g1098(.dina(w_n1399_0[1]),.dinb(w_n739_0[2]),.dout(n1400),.clk(gclk));
	jnot g1099(.din(w_n739_0[1]),.dout(n1401),.clk(gclk));
	jand g1100(.dina(w_n1398_0[0]),.dinb(w_dff_B_Q5aEoJqx2_1),.dout(n1402),.clk(gclk));
	jor g1101(.dina(n1402),.dinb(w_n651_0[1]),.dout(n1403),.clk(gclk));
	jor g1102(.dina(n1403),.dinb(n1400),.dout(n1404),.clk(gclk));
	jand g1103(.dina(w_dff_B_IKKyRrnr9_0),.dinb(w_n1394_0[1]),.dout(n1405),.clk(gclk));
	jnot g1104(.din(w_n1394_0[0]),.dout(n1406),.clk(gclk));
	jxor g1105(.dina(w_n1399_0[0]),.dinb(w_n968_0[0]),.dout(n1407),.clk(gclk));
	jand g1106(.dina(w_dff_B_0jfqp2Sr6_0),.dinb(n1406),.dout(n1408),.clk(gclk));
	jor g1107(.dina(n1408),.dinb(w_dff_B_jKVjrq5X9_1),.dout(n1409),.clk(gclk));
	jnot g1108(.din(w_n1409_0[1]),.dout(n1410),.clk(gclk));
	jxor g1109(.dina(w_n629_0[0]),.dinb(w_n625_0[0]),.dout(n1411),.clk(gclk));
	jnot g1110(.din(w_n1411_0[1]),.dout(n1412),.clk(gclk));
	jxor g1111(.dina(w_n806_0[1]),.dinb(w_n828_0[1]),.dout(n1413),.clk(gclk));
	jnot g1112(.din(w_n614_1[1]),.dout(n1414),.clk(gclk));
	jnot g1113(.din(w_n717_0[0]),.dout(n1415),.clk(gclk));
	jand g1114(.dina(w_n622_1[0]),.dinb(w_n828_0[0]),.dout(n1416),.clk(gclk));
	jand g1115(.dina(w_n628_0[0]),.dinb(w_G523_0[1]),.dout(n1417),.clk(gclk));
	jor g1116(.dina(n1417),.dinb(w_n829_0[0]),.dout(n1418),.clk(gclk));
	jor g1117(.dina(n1418),.dinb(n1416),.dout(n1419),.clk(gclk));
	jand g1118(.dina(n1419),.dinb(w_dff_B_41D4gjXK6_1),.dout(n1420),.clk(gclk));
	jxor g1119(.dina(w_n622_0[2]),.dinb(w_n618_0[1]),.dout(n1421),.clk(gclk));
	jnot g1120(.din(w_n1421_0[1]),.dout(n1422),.clk(gclk));
	jor g1121(.dina(w_dff_B_5XddWEBp3_0),.dinb(n1420),.dout(n1423),.clk(gclk));
	jor g1122(.dina(w_n1421_0[0]),.dinb(w_n819_0[0]),.dout(n1424),.clk(gclk));
	jand g1123(.dina(n1424),.dinb(w_dff_B_DZsrSaJC9_1),.dout(n1425),.clk(gclk));
	jxor g1124(.dina(w_n1425_0[1]),.dinb(w_dff_B_m1reyT1g6_1),.dout(n1426),.clk(gclk));
	jand g1125(.dina(n1426),.dinb(n1413),.dout(n1427),.clk(gclk));
	jnot g1126(.din(w_G2174_0[1]),.dout(n1428),.clk(gclk));
	jxor g1127(.dina(w_n806_0[0]),.dinb(w_n721_0[1]),.dout(n1429),.clk(gclk));
	jxor g1128(.dina(w_n1425_0[0]),.dinb(w_n614_1[0]),.dout(n1430),.clk(gclk));
	jand g1129(.dina(n1430),.dinb(n1429),.dout(n1431),.clk(gclk));
	jor g1130(.dina(n1431),.dinb(w_dff_B_E8bw2Xc02_1),.dout(n1432),.clk(gclk));
	jor g1131(.dina(n1432),.dinb(w_dff_B_93VvCCoL9_1),.dout(n1433),.clk(gclk));
	jxor g1132(.dina(w_n729_0[1]),.dinb(w_n614_0[2]),.dout(n1434),.clk(gclk));
	jnot g1133(.din(w_n1434_0[1]),.dout(n1435),.clk(gclk));
	jor g1134(.dina(w_n622_0[1]),.dinb(w_n721_0[0]),.dout(n1436),.clk(gclk));
	jand g1135(.dina(n1436),.dinb(w_n723_0[0]),.dout(n1437),.clk(gclk));
	jxor g1136(.dina(w_dff_B_JlEetKWX5_0),.dinb(w_n727_0[0]),.dout(n1438),.clk(gclk));
	jand g1137(.dina(w_n1438_0[1]),.dinb(n1435),.dout(n1439),.clk(gclk));
	jnot g1138(.din(w_n1438_0[0]),.dout(n1440),.clk(gclk));
	jand g1139(.dina(w_dff_B_rYpnkdck4_0),.dinb(w_n1434_0[0]),.dout(n1441),.clk(gclk));
	jor g1140(.dina(n1441),.dinb(w_G2174_0[0]),.dout(n1442),.clk(gclk));
	jor g1141(.dina(n1442),.dinb(n1439),.dout(n1443),.clk(gclk));
	jand g1142(.dina(w_dff_B_B8p0AihC4_0),.dinb(n1433),.dout(n1444),.clk(gclk));
	jxor g1143(.dina(n1444),.dinb(w_n787_0[0]),.dout(n1445),.clk(gclk));
	jxor g1144(.dina(w_n1445_0[1]),.dinb(w_dff_B_T5OrYCv76_1),.dout(n1446),.clk(gclk));
	jor g1145(.dina(w_n1446_0[1]),.dinb(w_n1410_0[1]),.dout(n1447),.clk(gclk));
	jxor g1146(.dina(w_n1445_0[0]),.dinb(w_n1411_0[0]),.dout(n1448),.clk(gclk));
	jor g1147(.dina(n1448),.dinb(w_n1409_0[0]),.dout(n1449),.clk(gclk));
	jand g1148(.dina(n1449),.dinb(w_G4091_1[1]),.dout(n1450),.clk(gclk));
	jand g1149(.dina(n1450),.dinb(w_n1447_0[1]),.dout(n1451),.clk(gclk));
	jor g1150(.dina(n1451),.dinb(w_dff_B_srRKSC302_1),.dout(n1452),.clk(gclk));
	jand g1151(.dina(w_n1452_0[1]),.dinb(w_dff_B_pt4Np9lk0_1),.dout(w_dff_A_SURhQcVE9_2),.clk(gclk));
	jor g1152(.dina(w_G4091_1[0]),.dinb(G118),.dout(n1454),.clk(gclk));
	jand g1153(.dina(w_G251_2[2]),.dinb(w_n460_0[2]),.dout(n1455),.clk(gclk));
	jand g1154(.dina(w_G248_3[0]),.dinb(w_G234_1[0]),.dout(n1456),.clk(gclk));
	jor g1155(.dina(n1456),.dinb(w_n462_0[0]),.dout(n1457),.clk(gclk));
	jor g1156(.dina(n1457),.dinb(n1455),.dout(n1458),.clk(gclk));
	jand g1157(.dina(w_n366_2[2]),.dinb(w_n460_0[1]),.dout(n1459),.clk(gclk));
	jand g1158(.dina(w_n368_3[0]),.dinb(w_G234_0[2]),.dout(n1460),.clk(gclk));
	jor g1159(.dina(n1460),.dinb(w_G435_0[1]),.dout(n1461),.clk(gclk));
	jor g1160(.dina(n1461),.dinb(w_dff_B_ESW2Jyin8_1),.dout(n1462),.clk(gclk));
	jand g1161(.dina(n1462),.dinb(w_dff_B_PzdBPeFS4_1),.dout(n1463),.clk(gclk));
	jor g1162(.dina(w_n402_1[1]),.dinb(w_G226_1[0]),.dout(n1464),.clk(gclk));
	jor g1163(.dina(w_n405_1[1]),.dinb(w_n530_0[2]),.dout(n1465),.clk(gclk));
	jand g1164(.dina(n1465),.dinb(w_G422_0[2]),.dout(n1466),.clk(gclk));
	jand g1165(.dina(n1466),.dinb(w_dff_B_PS8UhcAt3_1),.dout(n1467),.clk(gclk));
	jor g1166(.dina(w_G254_1[0]),.dinb(w_G226_0[2]),.dout(n1468),.clk(gclk));
	jor g1167(.dina(w_G242_1[0]),.dinb(w_n530_0[1]),.dout(n1469),.clk(gclk));
	jand g1168(.dina(n1469),.dinb(w_n532_0[0]),.dout(n1470),.clk(gclk));
	jand g1169(.dina(n1470),.dinb(w_dff_B_Z0Onc9aE6_1),.dout(n1471),.clk(gclk));
	jor g1170(.dina(n1471),.dinb(n1467),.dout(n1472),.clk(gclk));
	jxor g1171(.dina(n1472),.dinb(w_n528_0[0]),.dout(n1473),.clk(gclk));
	jor g1172(.dina(w_n402_1[0]),.dinb(w_G218_1[0]),.dout(n1474),.clk(gclk));
	jor g1173(.dina(w_n405_1[0]),.dinb(w_n507_0[2]),.dout(n1475),.clk(gclk));
	jand g1174(.dina(n1475),.dinb(w_G468_0[1]),.dout(n1476),.clk(gclk));
	jand g1175(.dina(n1476),.dinb(w_dff_B_rzADqUVV1_1),.dout(n1477),.clk(gclk));
	jor g1176(.dina(w_G254_0[2]),.dinb(w_G218_0[2]),.dout(n1478),.clk(gclk));
	jor g1177(.dina(w_G242_0[2]),.dinb(w_n507_0[1]),.dout(n1479),.clk(gclk));
	jand g1178(.dina(n1479),.dinb(w_n509_0[0]),.dout(n1480),.clk(gclk));
	jand g1179(.dina(n1480),.dinb(w_dff_B_p5kmLarl3_1),.dout(n1481),.clk(gclk));
	jor g1180(.dina(n1481),.dinb(n1477),.dout(n1482),.clk(gclk));
	jand g1181(.dina(w_G251_2[1]),.dinb(w_n541_0[2]),.dout(n1483),.clk(gclk));
	jand g1182(.dina(w_G248_2[2]),.dinb(w_G210_1[0]),.dout(n1484),.clk(gclk));
	jor g1183(.dina(n1484),.dinb(w_n543_0[0]),.dout(n1485),.clk(gclk));
	jor g1184(.dina(n1485),.dinb(n1483),.dout(n1486),.clk(gclk));
	jand g1185(.dina(w_n366_2[1]),.dinb(w_n541_0[1]),.dout(n1487),.clk(gclk));
	jand g1186(.dina(w_n368_2[2]),.dinb(w_G210_0[2]),.dout(n1488),.clk(gclk));
	jor g1187(.dina(n1488),.dinb(w_G457_0[2]),.dout(n1489),.clk(gclk));
	jor g1188(.dina(n1489),.dinb(w_dff_B_xqQZZMkN9_1),.dout(n1490),.clk(gclk));
	jand g1189(.dina(n1490),.dinb(w_dff_B_M2BfNANf4_1),.dout(n1491),.clk(gclk));
	jxor g1190(.dina(n1491),.dinb(n1482),.dout(n1492),.clk(gclk));
	jxor g1191(.dina(n1492),.dinb(n1473),.dout(n1493),.clk(gclk));
	jxor g1192(.dina(n1493),.dinb(w_dff_B_McPhVsr13_1),.dout(n1494),.clk(gclk));
	jand g1193(.dina(w_n495_0[2]),.dinb(w_G251_2[0]),.dout(n1495),.clk(gclk));
	jand g1194(.dina(w_G281_1[0]),.dinb(w_G248_2[1]),.dout(n1496),.clk(gclk));
	jor g1195(.dina(n1496),.dinb(w_n497_0[1]),.dout(n1497),.clk(gclk));
	jor g1196(.dina(n1497),.dinb(n1495),.dout(n1498),.clk(gclk));
	jand g1197(.dina(w_n495_0[1]),.dinb(w_n366_2[0]),.dout(n1499),.clk(gclk));
	jand g1198(.dina(w_G281_0[2]),.dinb(w_n368_2[1]),.dout(n1500),.clk(gclk));
	jor g1199(.dina(n1500),.dinb(w_G374_0[0]),.dout(n1501),.clk(gclk));
	jor g1200(.dina(n1501),.dinb(w_dff_B_t4xIJt4T5_1),.dout(n1502),.clk(gclk));
	jand g1201(.dina(n1502),.dinb(w_dff_B_F7dSwWAA2_1),.dout(n1503),.clk(gclk));
	jand g1202(.dina(w_n449_0[2]),.dinb(w_G251_1[2]),.dout(n1504),.clk(gclk));
	jand g1203(.dina(w_G265_1[0]),.dinb(w_G248_2[0]),.dout(n1505),.clk(gclk));
	jor g1204(.dina(n1505),.dinb(w_n451_0[1]),.dout(n1506),.clk(gclk));
	jor g1205(.dina(n1506),.dinb(n1504),.dout(n1507),.clk(gclk));
	jand g1206(.dina(w_n449_0[1]),.dinb(w_n366_1[2]),.dout(n1508),.clk(gclk));
	jand g1207(.dina(w_G265_0[2]),.dinb(w_n368_2[0]),.dout(n1509),.clk(gclk));
	jor g1208(.dina(n1509),.dinb(w_G400_0[1]),.dout(n1510),.clk(gclk));
	jor g1209(.dina(n1510),.dinb(w_dff_B_dA7S9O0q4_1),.dout(n1511),.clk(gclk));
	jand g1210(.dina(n1511),.dinb(w_dff_B_8WJiVgDg4_1),.dout(n1512),.clk(gclk));
	jxor g1211(.dina(n1512),.dinb(n1503),.dout(n1513),.clk(gclk));
	jor g1212(.dina(w_G257_1[0]),.dinb(w_n402_0[2]),.dout(n1514),.clk(gclk));
	jor g1213(.dina(w_n471_0[2]),.dinb(w_n405_0[2]),.dout(n1515),.clk(gclk));
	jand g1214(.dina(n1515),.dinb(w_G389_0[0]),.dout(n1516),.clk(gclk));
	jand g1215(.dina(n1516),.dinb(w_dff_B_s5CmWdDh1_1),.dout(n1517),.clk(gclk));
	jor g1216(.dina(w_G257_0[2]),.dinb(w_G254_0[1]),.dout(n1518),.clk(gclk));
	jor g1217(.dina(w_n471_0[1]),.dinb(w_G242_0[1]),.dout(n1519),.clk(gclk));
	jand g1218(.dina(n1519),.dinb(w_n473_0[1]),.dout(n1520),.clk(gclk));
	jand g1219(.dina(n1520),.dinb(w_dff_B_pwRFMlrp9_1),.dout(n1521),.clk(gclk));
	jor g1220(.dina(n1521),.dinb(n1517),.dout(n1522),.clk(gclk));
	jand g1221(.dina(w_n484_0[2]),.dinb(w_G251_1[1]),.dout(n1523),.clk(gclk));
	jand g1222(.dina(w_G273_1[0]),.dinb(w_G248_1[2]),.dout(n1524),.clk(gclk));
	jor g1223(.dina(n1524),.dinb(w_n486_0[1]),.dout(n1525),.clk(gclk));
	jor g1224(.dina(n1525),.dinb(n1523),.dout(n1526),.clk(gclk));
	jand g1225(.dina(w_n484_0[1]),.dinb(w_n366_1[1]),.dout(n1527),.clk(gclk));
	jand g1226(.dina(w_G273_0[2]),.dinb(w_n368_1[2]),.dout(n1528),.clk(gclk));
	jor g1227(.dina(n1528),.dinb(w_G411_0[0]),.dout(n1529),.clk(gclk));
	jor g1228(.dina(n1529),.dinb(w_dff_B_AJTqV7fd2_1),.dout(n1530),.clk(gclk));
	jand g1229(.dina(n1530),.dinb(w_dff_B_m1R52wP16_1),.dout(n1531),.clk(gclk));
	jxor g1230(.dina(n1531),.dinb(n1522),.dout(n1532),.clk(gclk));
	jxor g1231(.dina(n1532),.dinb(n1513),.dout(n1533),.clk(gclk));
	jand g1232(.dina(w_n1533_0[1]),.dinb(w_n1494_0[1]),.dout(n1534),.clk(gclk));
	jnot g1233(.din(n1534),.dout(n1535),.clk(gclk));
	jor g1234(.dina(w_n1533_0[0]),.dinb(w_n1494_0[0]),.dout(n1536),.clk(gclk));
	jand g1235(.dina(n1536),.dinb(w_n750_0[2]),.dout(n1537),.clk(gclk));
	jand g1236(.dina(n1537),.dinb(n1535),.dout(n1538),.clk(gclk));
	jor g1237(.dina(n1454),.dinb(w_n746_0[1]),.dout(n1539),.clk(gclk));
	jor g1238(.dina(n1538),.dinb(w_G4092_1[0]),.dout(n1540),.clk(gclk));
	jxor g1239(.dina(w_n583_0[1]),.dinb(w_n578_0[0]),.dout(n1541),.clk(gclk));
	jxor g1240(.dina(n1541),.dinb(w_n943_0[0]),.dout(n1542),.clk(gclk));
	jnot g1241(.din(n1542),.dout(n1543),.clk(gclk));
	jand g1242(.dina(w_n587_0[2]),.dinb(w_G1497_0[2]),.dout(n1544),.clk(gclk));
	jor g1243(.dina(w_dff_B_6kfQng679_0),.dinb(w_n696_0[0]),.dout(n1545),.clk(gclk));
	jnot g1244(.din(w_n1545_0[1]),.dout(n1546),.clk(gclk));
	jor g1245(.dina(w_n944_0[0]),.dinb(w_n930_0[1]),.dout(n1547),.clk(gclk));
	jand g1246(.dina(n1547),.dinb(w_n706_0[0]),.dout(n1548),.clk(gclk));
	jxor g1247(.dina(n1548),.dinb(w_n928_0[0]),.dout(n1549),.clk(gclk));
	jxor g1248(.dina(w_n605_1[1]),.dinb(w_n948_0[1]),.dout(n1550),.clk(gclk));
	jxor g1249(.dina(w_dff_B_3TEKFXjF7_0),.dinb(n1549),.dout(n1551),.clk(gclk));
	jand g1250(.dina(w_dff_B_wrBjtwS76_0),.dinb(n1546),.dout(n1552),.clk(gclk));
	jxor g1251(.dina(w_n605_1[0]),.dinb(w_n703_0[0]),.dout(n1553),.clk(gclk));
	jand g1252(.dina(w_n605_0[2]),.dinb(w_n948_0[0]),.dout(n1554),.clk(gclk));
	jor g1253(.dina(n1554),.dinb(w_n702_0[0]),.dout(n1555),.clk(gclk));
	jnot g1254(.din(w_n1555_0[1]),.dout(n1556),.clk(gclk));
	jor g1255(.dina(n1556),.dinb(w_n930_0[0]),.dout(n1557),.clk(gclk));
	jor g1256(.dina(w_n1555_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1257(.dina(n1558),.dinb(w_dff_B_IJNya5Rl8_1),.dout(n1559),.clk(gclk));
	jxor g1258(.dina(n1559),.dinb(w_n596_0[0]),.dout(n1560),.clk(gclk));
	jand g1259(.dina(w_n1560_0[1]),.dinb(w_n1553_0[1]),.dout(n1561),.clk(gclk));
	jnot g1260(.din(n1561),.dout(n1562),.clk(gclk));
	jor g1261(.dina(w_n1560_0[0]),.dinb(w_n1553_0[0]),.dout(n1563),.clk(gclk));
	jand g1262(.dina(w_dff_B_9mibG71Y7_0),.dinb(w_n1545_0[0]),.dout(n1564),.clk(gclk));
	jand g1263(.dina(n1564),.dinb(w_dff_B_fiDJVqRi0_1),.dout(n1565),.clk(gclk));
	jor g1264(.dina(n1565),.dinb(n1552),.dout(n1566),.clk(gclk));
	jnot g1265(.din(w_G1497_0[1]),.dout(n1567),.clk(gclk));
	jand g1266(.dina(w_n682_0[0]),.dinb(w_n687_0[0]),.dout(n1568),.clk(gclk));
	jand g1267(.dina(w_n1568_0[1]),.dinb(w_n574_0[0]),.dout(n1569),.clk(gclk));
	jxor g1268(.dina(n1569),.dinb(w_n561_0[1]),.dout(n1570),.clk(gclk));
	jxor g1269(.dina(w_n572_0[1]),.dinb(w_n681_1[1]),.dout(n1571),.clk(gclk));
	jor g1270(.dina(w_n856_0[0]),.dinb(w_n853_0[0]),.dout(n1572),.clk(gclk));
	jand g1271(.dina(w_n693_0[1]),.dinb(w_n585_0[0]),.dout(n1573),.clk(gclk));
	jor g1272(.dina(n1573),.dinb(w_n855_0[0]),.dout(n1574),.clk(gclk));
	jand g1273(.dina(n1574),.dinb(n1572),.dout(n1575),.clk(gclk));
	jxor g1274(.dina(n1575),.dinb(w_dff_B_LvevyD0u7_1),.dout(n1576),.clk(gclk));
	jxor g1275(.dina(n1576),.dinb(w_dff_B_ZEHe0Y898_1),.dout(n1577),.clk(gclk));
	jor g1276(.dina(n1577),.dinb(w_dff_B_KRgvwtkw4_1),.dout(n1578),.clk(gclk));
	jxor g1277(.dina(w_n693_0[0]),.dinb(w_n572_0[0]),.dout(n1579),.clk(gclk));
	jor g1278(.dina(w_n857_0[0]),.dinb(w_n681_1[0]),.dout(n1580),.clk(gclk));
	jnot g1279(.din(w_n681_0[2]),.dout(n1581),.clk(gclk));
	jor g1280(.dina(w_n680_0[0]),.dinb(n1581),.dout(n1582),.clk(gclk));
	jor g1281(.dina(n1582),.dinb(w_n689_0[0]),.dout(n1583),.clk(gclk));
	jxor g1282(.dina(n1583),.dinb(w_n567_0[1]),.dout(n1584),.clk(gclk));
	jand g1283(.dina(w_dff_B_8LDZHcFf0_0),.dinb(n1580),.dout(n1585),.clk(gclk));
	jxor g1284(.dina(w_n1568_0[0]),.dinb(w_n561_0[0]),.dout(n1586),.clk(gclk));
	jxor g1285(.dina(w_dff_B_13uFmaH52_0),.dinb(n1585),.dout(n1587),.clk(gclk));
	jxor g1286(.dina(n1587),.dinb(w_dff_B_Y0KUzQp49_1),.dout(n1588),.clk(gclk));
	jor g1287(.dina(n1588),.dinb(w_G1497_0[0]),.dout(n1589),.clk(gclk));
	jand g1288(.dina(w_dff_B_OBkh3hor7_0),.dinb(n1578),.dout(n1590),.clk(gclk));
	jxor g1289(.dina(n1590),.dinb(n1566),.dout(n1591),.clk(gclk));
	jand g1290(.dina(w_n1591_0[1]),.dinb(w_n1543_0[1]),.dout(n1592),.clk(gclk));
	jnot g1291(.din(n1592),.dout(n1593),.clk(gclk));
	jor g1292(.dina(w_n1591_0[0]),.dinb(w_n1543_0[0]),.dout(n1594),.clk(gclk));
	jand g1293(.dina(n1594),.dinb(w_G4091_0[2]),.dout(n1595),.clk(gclk));
	jand g1294(.dina(n1595),.dinb(n1593),.dout(n1596),.clk(gclk));
	jor g1295(.dina(n1596),.dinb(w_dff_B_JxnJFHBJ9_1),.dout(n1597),.clk(gclk));
	jand g1296(.dina(w_n1597_0[1]),.dinb(w_dff_B_bUlMydrC4_1),.dout(w_dff_A_uG8smKgl3_2),.clk(gclk));
	jand g1297(.dina(w_G4092_0[2]),.dinb(G97),.dout(n1599),.clk(gclk));
	jnot g1298(.din(n1599),.dout(n1600),.clk(gclk));
	jand g1299(.dina(w_dff_B_CczamCeA6_0),.dinb(w_n1597_0[0]),.dout(n1601),.clk(gclk));
	jnot g1300(.din(w_n1601_0[2]),.dout(n1602),.clk(gclk));
	jand g1301(.dina(w_n1602_0[1]),.dinb(w_n793_1[1]),.dout(n1603),.clk(gclk));
	jnot g1302(.din(w_n1447_0[0]),.dout(n1604),.clk(gclk));
	jand g1303(.dina(w_n1446_0[0]),.dinb(w_n1410_0[0]),.dout(n1605),.clk(gclk));
	jor g1304(.dina(n1605),.dinb(w_n750_0[1]),.dout(n1606),.clk(gclk));
	jor g1305(.dina(n1606),.dinb(n1604),.dout(n1607),.clk(gclk));
	jand g1306(.dina(n1607),.dinb(w_n1391_0[0]),.dout(n1608),.clk(gclk));
	jand g1307(.dina(w_G4092_0[1]),.dinb(G94),.dout(n1609),.clk(gclk));
	jor g1308(.dina(w_n1609_0[1]),.dinb(n1608),.dout(n1610),.clk(gclk));
	jand g1309(.dina(w_n1610_0[1]),.dinb(w_n797_1[1]),.dout(n1611),.clk(gclk));
	jand g1310(.dina(w_n799_1[1]),.dinb(w_G14_0[1]),.dout(n1612),.clk(gclk));
	jand g1311(.dina(w_n801_1[1]),.dinb(w_G64_0[1]),.dout(n1613),.clk(gclk));
	jor g1312(.dina(w_dff_B_zVkRJpEp9_0),.dinb(n1612),.dout(n1614),.clk(gclk));
	jor g1313(.dina(w_dff_B_pn9fF3NJ2_0),.dinb(n1611),.dout(n1615),.clk(gclk));
	jor g1314(.dina(n1615),.dinb(n1603),.dout(w_dff_A_jKaG1UkO8_2),.clk(gclk));
	jand g1315(.dina(w_n1602_0[0]),.dinb(w_n840_1[1]),.dout(n1617),.clk(gclk));
	jand g1316(.dina(w_n1610_0[0]),.dinb(w_n843_1[1]),.dout(n1618),.clk(gclk));
	jand g1317(.dina(w_n845_1[1]),.dinb(w_G14_0[0]),.dout(n1619),.clk(gclk));
	jand g1318(.dina(w_n847_1[1]),.dinb(w_G64_0[0]),.dout(n1620),.clk(gclk));
	jor g1319(.dina(w_dff_B_Iw1JI7LE5_0),.dinb(n1619),.dout(n1621),.clk(gclk));
	jor g1320(.dina(w_dff_B_vy2zsUTI4_0),.dinb(n1618),.dout(n1622),.clk(gclk));
	jor g1321(.dina(n1622),.dinb(n1617),.dout(w_dff_A_1hgo6KA25_2),.clk(gclk));
	jnot g1322(.din(w_G137_3[1]),.dout(n1624),.clk(gclk));
	jnot g1323(.din(w_n985_1[1]),.dout(n1625),.clk(gclk));
	jor g1324(.dina(w_n1601_0[1]),.dinb(w_dff_B_2TT89mhw0_1),.dout(n1626),.clk(gclk));
	jnot g1325(.din(w_n988_1[1]),.dout(n1627),.clk(gclk));
	jnot g1326(.din(w_n1609_0[0]),.dout(n1628),.clk(gclk));
	jand g1327(.dina(w_dff_B_VkqJ4JdF2_0),.dinb(w_n1452_0[0]),.dout(n1629),.clk(gclk));
	jor g1328(.dina(w_n1629_0[1]),.dinb(w_dff_B_lU0gpBps2_1),.dout(n1630),.clk(gclk));
	jnot g1329(.din(G179),.dout(n1631),.clk(gclk));
	jnot g1330(.din(w_n992_1[1]),.dout(n1632),.clk(gclk));
	jor g1331(.dina(n1632),.dinb(w_n1631_0[1]),.dout(n1633),.clk(gclk));
	jnot g1332(.din(G176),.dout(n1634),.clk(gclk));
	jnot g1333(.din(w_n990_1[1]),.dout(n1635),.clk(gclk));
	jor g1334(.dina(n1635),.dinb(w_n1634_0[1]),.dout(n1636),.clk(gclk));
	jand g1335(.dina(n1636),.dinb(w_dff_B_fNWvu0Ba5_1),.dout(n1637),.clk(gclk));
	jand g1336(.dina(w_dff_B_0HFVwDKA1_0),.dinb(n1630),.dout(n1638),.clk(gclk));
	jand g1337(.dina(n1638),.dinb(w_dff_B_WDSJg6To0_1),.dout(n1639),.clk(gclk));
	jor g1338(.dina(n1639),.dinb(w_n1624_0[1]),.dout(G658),.clk(gclk));
	jnot g1339(.din(w_n999_1[1]),.dout(n1641),.clk(gclk));
	jor g1340(.dina(w_n1601_0[0]),.dinb(w_dff_B_y6t5PHBq2_1),.dout(n1642),.clk(gclk));
	jnot g1341(.din(w_n1002_1[1]),.dout(n1643),.clk(gclk));
	jor g1342(.dina(w_n1629_0[0]),.dinb(w_dff_B_QQQYwGwz9_1),.dout(n1644),.clk(gclk));
	jnot g1343(.din(w_n1006_1[1]),.dout(n1645),.clk(gclk));
	jor g1344(.dina(n1645),.dinb(w_n1631_0[0]),.dout(n1646),.clk(gclk));
	jnot g1345(.din(w_n1004_1[1]),.dout(n1647),.clk(gclk));
	jor g1346(.dina(n1647),.dinb(w_n1634_0[0]),.dout(n1648),.clk(gclk));
	jand g1347(.dina(n1648),.dinb(w_dff_B_pjxcf6tk2_1),.dout(n1649),.clk(gclk));
	jand g1348(.dina(w_dff_B_sUjayH6W6_0),.dinb(n1644),.dout(n1650),.clk(gclk));
	jand g1349(.dina(n1650),.dinb(w_dff_B_kO1xlF5h5_1),.dout(n1651),.clk(gclk));
	jor g1350(.dina(n1651),.dinb(w_n1624_0[0]),.dout(G690),.clk(gclk));
	jdff g1351(.din(w_G141_1[0]),.dout(w_dff_A_cb5G565l2_1),.clk(gclk));
	jdff g1352(.din(w_G293_0[0]),.dout(w_dff_A_HUppY1yx4_1),.clk(gclk));
	jdff g1353(.din(w_G3173_0[0]),.dout(w_dff_A_bgbfZxUg8_1),.clk(gclk));
	jnot g1354(.din(w_G545_0[1]),.dout(w_dff_A_lAjJ6ntN2_1),.clk(gclk));
	jnot g1355(.din(w_G545_0[0]),.dout(w_dff_A_0HHr3PS48_1),.clk(gclk));
	jdff g1356(.din(w_G137_3[0]),.dout(w_dff_A_0NtsHe4k0_1),.clk(gclk));
	jdff g1357(.din(w_G141_0[2]),.dout(w_dff_A_U6IqrDOA3_1),.clk(gclk));
	jdff g1358(.din(w_G1_2[0]),.dout(w_dff_A_NmT0XjCB0_1),.clk(gclk));
	jdff g1359(.din(w_G549_0[1]),.dout(w_dff_A_FwI0aGbj2_1),.clk(gclk));
	jdff g1360(.din(w_G299_0[1]),.dout(w_dff_A_IM6ysSsv4_1),.clk(gclk));
	jnot g1361(.din(w_G549_0[0]),.dout(w_dff_A_ELUGCjOB6_1),.clk(gclk));
	jdff g1362(.din(w_G1_1[2]),.dout(w_dff_A_YeaIpaov7_1),.clk(gclk));
	jdff g1363(.din(w_G1_1[1]),.dout(w_dff_A_SpO2BMhM3_1),.clk(gclk));
	jdff g1364(.din(w_G1_1[0]),.dout(w_dff_A_abVhkHvY7_1),.clk(gclk));
	jdff g1365(.din(w_G1_0[2]),.dout(w_dff_A_qpWbjoOy4_1),.clk(gclk));
	jdff g1366(.din(w_G299_0[0]),.dout(w_dff_A_lD6XExhc7_1),.clk(gclk));
	jor g1367(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_TR3QSKJ91_2),.clk(gclk));
	jand g1368(.dina(w_n652_0[0]),.dinb(w_n633_0[1]),.dout(w_dff_A_QmKqJRIv2_2),.clk(gclk));
	jand g1369(.dina(w_n607_0[0]),.dinb(w_n587_0[1]),.dout(w_dff_A_t4OEWpbI4_2),.clk(gclk));
	jor g1370(.dina(w_n709_0[0]),.dinb(w_n697_0[0]),.dout(w_dff_A_KD56kTfy9_2),.clk(gclk));
	jor g1371(.dina(w_n742_0[0]),.dinb(w_n733_0[0]),.dout(w_dff_A_Cy9lkNbV7_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_KUzeLFZw3_1),.doutc(w_G4_0[2]),.din(w_dff_B_3zTcJTIs9_3));
	jspl jspl_w_G4_1(.douta(w_dff_A_SL3qSCfQ3_0),.doutb(w_G4_1[1]),.din(w_G4_0[0]));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(w_dff_B_CChcr1BA4_2));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(w_dff_B_UE8GuEbX6_2));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_JPVxV5JX3_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_ntYLpOYK3_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_S7J5IsmI3_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_cQ9zOYqq2_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(w_dff_B_dxC1OtnG9_2));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(w_dff_B_SYbYFckq7_2));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_zwPJdQEF4_2));
	jspl jspl_w_G54_0(.douta(w_dff_A_vpdtxn4N0_0),.doutb(w_G54_0[1]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_MZhMwQa67_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_tjMC8laf8_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(w_dff_B_dmDgtYiK5_2));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_gGqDyEHP8_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(w_dff_B_SAJzS6I19_2));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(w_dff_B_l3xCiwCo2_2));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(w_dff_B_jN6unUfh7_2));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(w_dff_B_0gLVztIc0_2));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_mOQjkljC0_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_skpGvuxw4_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(w_dff_B_pc46jYw56_2));
	jspl jspl_w_G123_0(.douta(w_dff_A_BrrDWsJJ5_0),.doutb(w_G123_0[1]),.din(w_dff_B_k7ccmGjA3_2));
	jspl jspl_w_G132_0(.douta(w_dff_A_de4oxTsm6_0),.doutb(w_G132_0[1]),.din(w_dff_B_i0Dq756B2_2));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_Y7lYWyOM7_0),.doutb(w_dff_A_qfPzuRhQ3_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_so03MYB81_0),.doutb(w_dff_A_2NRd1JdT9_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_rYHWvkE08_0),.doutb(w_dff_A_E3CF4CRp0_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_LoVGMRWh5_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_383ZEy6I1_0),.doutb(w_dff_A_ju5dP4BX9_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_RQQIh7vn0_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_ZlmiawB56_0),.doutb(w_dff_A_qp4LGAap9_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_Dg47uAWB2_1),.doutc(w_dff_A_srnJSoTh0_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_dff_A_1BC24AqY8_0),.doutb(w_G137_8[1]),.doutc(w_dff_A_e6UNA8IQ6_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_8SuW07jG0_1),.doutc(w_dff_A_a5cZcJOE8_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_NRmMTPDk0_0),.doutb(w_dff_A_9tMO6vDT1_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_Yql3Al7D3_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_uqpvHaIJ6_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_Jwib4FT85_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_tyClrbYL5_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_rhmpJRnq2_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_wnoB62px8_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_TvkVAIn21_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_MAJmmH5t1_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_JcnLwAmB3_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_SGUhAMb97_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_uQNPPLHu0_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_E8Ow1mSb0_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_oPu1wzDG3_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_YXrldbBk9_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_7lMbWqIo5_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_cFW4n59S5_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_YbWxK6xW4_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_mLxJD7f59_2));
	jspl3 jspl3_w_G206_0(.douta(w_dff_A_4WsIfzAC9_0),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_W0Bp2O9F7_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_dff_A_2Fos1n793_1),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl3 jspl3_w_G210_2(.douta(w_G210_2[0]),.doutb(w_dff_A_Wvhep0ki2_1),.doutc(w_G210_2[2]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_9a9Fd7d06_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl3 jspl3_w_G218_2(.douta(w_G218_2[0]),.doutb(w_dff_A_sblDCa1a4_1),.doutc(w_G218_2[2]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_6CZxVukQ2_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G226_2(.douta(w_G226_2[0]),.doutb(w_dff_A_8jIdLr0h7_1),.doutc(w_G226_2[2]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_5gdKQzfI4_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_y5HQIe6X9_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_HpUvt8bN7_1),.doutc(w_dff_A_L1bi1yru6_2),.din(G242));
	jspl3 jspl3_w_G242_1(.douta(w_dff_A_cQwm38V27_0),.doutb(w_dff_A_Q5zt9qC28_1),.doutc(w_G242_1[2]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_G245_0[0]),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_iVswdcIQ0_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl jspl_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_xBie47Qk2_1),.doutc(w_dff_A_EmzcZY9t8_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_G251_1[0]),.doutb(w_dff_A_K6d3lJfk5_1),.doutc(w_dff_A_CwMNRSJ39_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_dff_A_g05iV4qr9_1),.doutc(w_dff_A_umsvQfiS2_2),.din(w_G251_1[0]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl3 jspl3_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.doutc(w_G254_1[2]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_0vmrnqG67_0),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G257_2(.douta(w_G257_2[0]),.doutb(w_dff_A_KFQivGam9_1),.doutc(w_G257_2[2]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_e3JIbNxC8_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_G265_1[1]),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl jspl_w_G265_2(.douta(w_dff_A_GHf1WuLw3_0),.doutb(w_G265_2[1]),.din(w_G265_0[1]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_rbLJ0fbJ2_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_G273_1[1]),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl3 jspl3_w_G273_2(.douta(w_G273_2[0]),.doutb(w_dff_A_HlJL891t2_1),.doutc(w_G273_2[2]),.din(w_G273_0[1]));
	jspl jspl_w_G280_0(.douta(w_G280_0[0]),.doutb(w_dff_A_dIXvuexv7_1),.din(G280));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_Z2ld8Ms42_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_zwQWhkLL1_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_dff_A_9cjRjcFv5_0),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_rU5hIRg20_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_4NWISi2H3_0),.doutb(w_dff_A_j41D3iUL7_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_77KRC1lc4_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_G316_0[2]),.din(G316));
	jspl3 jspl3_w_G316_1(.douta(w_dff_A_msxUPXKl5_0),.doutb(w_G316_1[1]),.doutc(w_G316_1[2]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_dff_A_o35FUYa91_1),.doutc(w_G324_0[2]),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_2TCoX7101_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_7Eb9Jmja7_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_G332_1[1]),.doutc(w_dff_A_TWNRPvyV2_2),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_IDL7tBGd6_0),.doutb(w_G332_2[1]),.doutc(w_G332_2[2]),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_dff_A_289YKKsd7_0),.doutb(w_G332_3[1]),.doutc(w_dff_A_5nV0ELg97_2),.din(w_G332_0[2]));
	jspl3 jspl3_w_G332_4(.douta(w_dff_A_LT5SgMpK3_0),.doutb(w_G332_4[1]),.doutc(w_G332_4[2]),.din(w_G332_1[0]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl3 jspl3_w_G335_1(.douta(w_G335_1[0]),.doutb(w_G335_1[1]),.doutc(w_dff_A_6CHDTV882_2),.din(w_G335_0[0]));
	jspl3 jspl3_w_G335_2(.douta(w_G335_2[0]),.doutb(w_G335_2[1]),.doutc(w_G335_2[2]),.din(w_G335_0[1]));
	jspl3 jspl3_w_G335_3(.douta(w_dff_A_X5VE5Rn87_0),.doutb(w_G335_3[1]),.doutc(w_G335_3[2]),.din(w_G335_0[2]));
	jspl jspl_w_G335_4(.douta(w_dff_A_Y0C5iHwL0_0),.doutb(w_G335_4[1]),.din(w_G335_1[0]));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_8Kvxk1sW7_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_bcnZ5QXg4_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_IcUKXp9b7_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_G351_0[2]),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_dff_A_OglsVBYO9_0),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_kJ1VNvQG9_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_JD0BOWzY6_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_dff_A_iMsQLFAt3_1),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G369_0(.douta(w_dff_A_7RobHvig9_0),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_dff_A_jk4Zfurw9_0),.doutb(w_dff_A_rrQKLtgY1_1),.doutc(w_G374_0[2]),.din(G374));
	jspl3 jspl3_w_G389_0(.douta(w_dff_A_ntbxNQMz8_0),.doutb(w_dff_A_G0yvkdsE8_1),.doutc(w_G389_0[2]),.din(G389));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_LR4UwY9l0_1),.doutc(w_dff_A_bodr78eO0_2),.din(G400));
	jspl jspl_w_G400_1(.douta(w_dff_A_SQiowSOU1_0),.doutb(w_G400_1[1]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_Zw8gwf5R7_0),.doutb(w_dff_A_6BR4DVNt6_1),.doutc(w_G411_0[2]),.din(G411));
	jspl3 jspl3_w_G422_0(.douta(w_dff_A_dQHbuo6n9_0),.doutb(w_G422_0[1]),.doutc(w_dff_A_TPUCpvG71_2),.din(G422));
	jspl3 jspl3_w_G422_1(.douta(w_G422_1[0]),.doutb(w_G422_1[1]),.doutc(w_G422_1[2]),.din(w_G422_0[0]));
	jspl jspl_w_G422_2(.douta(w_dff_A_dTobYgT19_0),.doutb(w_G422_2[1]),.din(w_G422_0[1]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_fxjrjCh67_1),.doutc(w_dff_A_93tWPI9q8_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_BKERlw5H5_0),.doutb(w_dff_A_93DnRBLx5_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_G6lbEGdA0_1),.doutc(w_dff_A_jWocplEn0_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_5RAOQJeX5_0),.doutb(w_dff_A_PjIXy07J6_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_dff_A_kIlLJhno4_0),.doutb(w_G457_0[1]),.doutc(w_dff_A_NIHaGDVF2_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_G457_1[0]),.doutb(w_G457_1[1]),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl jspl_w_G457_2(.douta(w_dff_A_PpQBE0k26_0),.doutb(w_G457_2[1]),.din(w_G457_0[1]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_IcWadWZz6_1),.doutc(w_dff_A_KNLrAf8K1_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_P62yhVsH3_0),.doutb(w_dff_A_6D3Di4A10_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_G479_0[0]),.doutb(w_dff_A_1kxmuCHH2_1),.doutc(w_dff_A_5hM7wWQg4_2),.din(G479));
	jspl jspl_w_G479_1(.douta(w_dff_A_MvzDF7Oj4_0),.doutb(w_G479_1[1]),.din(w_G479_0[0]));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_eREKj2st1_1),.doutc(w_dff_A_4J7QjujL1_2),.din(G490));
	jspl3 jspl3_w_G490_1(.douta(w_dff_A_4rgexoVy5_0),.doutb(w_dff_A_sGs16ISw7_1),.doutc(w_G490_1[2]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_G503_0[0]),.doutb(w_dff_A_uvjxOwaX1_1),.doutc(w_dff_A_Pru7XwWy6_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_dff_A_t8pGFjp86_0),.doutb(w_dff_A_MIQ1Y4FX5_1),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl3 jspl3_w_G514_0(.douta(w_G514_0[0]),.doutb(w_dff_A_6st0OpoW4_1),.doutc(w_dff_A_rhNxgrBE4_2),.din(G514));
	jspl jspl_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.din(w_G514_0[0]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_6PiK53K50_1),.doutc(w_dff_A_zDMoByYg7_2),.din(G523));
	jspl jspl_w_G523_1(.douta(w_dff_A_QGecVUIb6_0),.doutb(w_G523_1[1]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_G534_0[0]),.doutb(w_dff_A_1OY5sP727_1),.doutc(w_dff_A_0pFK2Ner1_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_dff_A_hFq9wJpJ8_0),.doutb(w_dff_A_5qhikpfe9_1),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_G559_0[0]),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_JqaM0uqn6_0),.doutb(w_G1497_0[1]),.doutc(w_dff_A_EWHZ9Osq4_2),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_G1689_0[1]),.doutc(w_dff_A_shACUS9a7_2),.din(G1689));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_kWN7fJzX1_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_G1691_0[1]),.doutc(w_dff_A_T9Chpajb1_2),.din(G1691));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_UygF6HbI1_1),.doutc(w_G1694_0[2]),.din(G1694));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_2PvgxPFn8_0),.doutb(w_G2174_0[1]),.doutc(w_dff_A_yp2Uiusj4_2),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_ZMRpH7Cm0_0),.doutb(w_dff_A_bt1O9L7I5_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_GertBESm2_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_j4F8Q4Q48_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_dff_A_vCMXz4iL1_0),.doutb(w_G3724_0[1]),.doutc(w_dff_A_Y3km0hto5_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_Jh1PO9Ub9_1),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_dff_A_Ts5zBysZ3_2),.din(G4088));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_dff_A_SGVINllK6_2),.din(G4089));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_4CRskux41_1),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_G4091_0[1]),.doutc(w_dff_A_mDT9zZ7v2_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_G4091_1[0]),.doutb(w_dff_A_kLbvHeRq5_1),.doutc(w_dff_A_m8eHBqdZ6_2),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_G4091_2[0]),.doutb(w_G4091_2[1]),.doutc(w_dff_A_5GaXf1406_2),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_G4092_0[1]),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_c9obuGxY8_0),.doutb(w_dff_A_zdrI3PDS9_1),.doutc(w_G4092_1[2]),.din(w_G4092_0[0]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_ywNt4EiO1_1),.din(G599_fa_));
	jspl jspl_w_G600_0(.douta(w_G600_0),.doutb(w_dff_A_wEbXZwDn0_1),.din(G600_fa_));
	jspl jspl_w_G601_0(.douta(w_dff_A_66KJWVwp8_0),.doutb(w_dff_A_XBKdFEY12_1),.din(G601_fa_));
	jspl jspl_w_G611_0(.douta(w_G611_0),.doutb(w_dff_A_pVw4klAf8_1),.din(G611_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_Kl1VYOge1_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_x86FEGCI7_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_4e4EIA5N1_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_snZJi9ST6_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_NU9RSijT7_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_ZXolT0V26_1),.din(G861_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_wR17c80c2_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_5Xx6TgKH7_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_qqGvtkqc6_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_N7LHGUu06_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_Z21vggDg8_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_5zsUPBA47_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_M2r8JevI0_1),.din(G877_fa_));
	jspl jspl_w_G1000_0(.douta(w_G1000_0),.doutb(w_dff_A_vxWk0kuz4_1),.din(G1000_fa_));
	jspl jspl_w_G826_0(.douta(w_G826_0),.doutb(w_dff_A_G7R4DQMb4_1),.din(G826_fa_));
	jspl jspl_w_G828_0(.douta(w_G828_0),.doutb(w_dff_A_Bmlo6mAl5_1),.din(G828_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_FIVSn6jT5_1),.din(G830_fa_));
	jspl jspl_w_G867_0(.douta(w_G867_0),.doutb(w_dff_A_0gsqbsOX9_1),.din(G867_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_Y9DXbQ481_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_D7BgWf7S7_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_dff_A_RvHiWXFc7_0),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n366_2(.douta(w_n366_2[0]),.doutb(w_n366_2[1]),.doutc(w_n366_2[2]),.din(w_n366_0[1]));
	jspl3 jspl3_w_n366_3(.douta(w_n366_3[0]),.doutb(w_n366_3[1]),.doutc(w_n366_3[2]),.din(w_n366_0[2]));
	jspl3 jspl3_w_n366_4(.douta(w_n366_4[0]),.doutb(w_n366_4[1]),.doutc(w_n366_4[2]),.din(w_n366_1[0]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl3 jspl3_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.doutc(w_n368_1[2]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n368_2(.douta(w_n368_2[0]),.doutb(w_n368_2[1]),.doutc(w_n368_2[2]),.din(w_n368_0[1]));
	jspl3 jspl3_w_n368_3(.douta(w_n368_3[0]),.doutb(w_n368_3[1]),.doutc(w_n368_3[2]),.din(w_n368_0[2]));
	jspl3 jspl3_w_n368_4(.douta(w_n368_4[0]),.doutb(w_n368_4[1]),.doutc(w_n368_4[2]),.din(w_n368_1[0]));
	jspl jspl_w_n368_5(.douta(w_n368_5[0]),.doutb(w_n368_5[1]),.din(w_n368_1[1]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl3 jspl3_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.doutc(w_n385_1[2]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.doutc(w_n386_1[2]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n386_2(.douta(w_n386_2[0]),.doutb(w_n386_2[1]),.doutc(w_n386_2[2]),.din(w_n386_0[1]));
	jspl3 jspl3_w_n386_3(.douta(w_n386_3[0]),.doutb(w_n386_3[1]),.doutc(w_n386_3[2]),.din(w_n386_0[2]));
	jspl3 jspl3_w_n386_4(.douta(w_n386_4[0]),.doutb(w_n386_4[1]),.doutc(w_n386_4[2]),.din(w_n386_1[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_dff_A_x1spk4jM5_2),.din(w_dff_B_Q4dSipxa8_3));
	jspl3 jspl3_w_n388_1(.douta(w_dff_A_tNKKSYbO1_0),.doutb(w_dff_A_UvZHh7uC5_1),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl3 jspl3_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.doutc(w_n389_1[2]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n389_2(.douta(w_n389_2[0]),.doutb(w_n389_2[1]),.doutc(w_n389_2[2]),.din(w_n389_0[1]));
	jspl3 jspl3_w_n389_3(.douta(w_n389_3[0]),.doutb(w_n389_3[1]),.doutc(w_n389_3[2]),.din(w_n389_0[2]));
	jspl3 jspl3_w_n389_4(.douta(w_n389_4[0]),.doutb(w_n389_4[1]),.doutc(w_n389_4[2]),.din(w_n389_1[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_dff_A_y5ATf2KU7_1),.din(n397));
	jspl3 jspl3_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.doutc(w_n398_0[2]),.din(n398));
	jspl3 jspl3_w_n401_0(.douta(w_dff_A_9RxrP5xD1_0),.doutb(w_n401_0[1]),.doutc(w_dff_A_USqn9juS4_2),.din(n401));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.doutc(w_n402_1[2]),.din(w_n402_0[0]));
	jspl jspl_w_n402_2(.douta(w_n402_2[0]),.doutb(w_n402_2[1]),.din(w_n402_0[1]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n405_1(.douta(w_n405_1[0]),.doutb(w_n405_1[1]),.doutc(w_n405_1[2]),.din(w_n405_0[0]));
	jspl jspl_w_n405_2(.douta(w_n405_2[0]),.doutb(w_n405_2[1]),.din(w_n405_0[1]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_dff_A_Rtj5CWw78_2),.din(n410));
	jspl jspl_w_n410_1(.douta(w_dff_A_gHKJPNrq2_0),.doutb(w_n410_1[1]),.din(w_n410_0[0]));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(n416));
	jspl3 jspl3_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.doutc(w_n419_0[2]),.din(n419));
	jspl3 jspl3_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.doutc(w_n424_0[2]),.din(n424));
	jspl3 jspl3_w_n424_1(.douta(w_n424_1[0]),.doutb(w_n424_1[1]),.doutc(w_n424_1[2]),.din(w_n424_0[0]));
	jspl jspl_w_n424_2(.douta(w_n424_2[0]),.doutb(w_n424_2[1]),.din(w_n424_0[1]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_dff_A_7Lv7AdWl5_1),.din(n426));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl3 jspl3_w_n437_0(.douta(w_dff_A_X8JEPTvo8_0),.doutb(w_n437_0[1]),.doutc(w_dff_A_rVsBUueX2_2),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_dff_A_n0fgwF552_0),.doutb(w_dff_A_S9nwTBvd1_1),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_dff_A_yzVfqSoE5_0),.doutb(w_n451_0[1]),.doutc(w_dff_A_C9wiUB3i5_2),.din(n451));
	jspl jspl_w_n451_1(.douta(w_dff_A_rdwYEB797_0),.doutb(w_n451_1[1]),.din(w_n451_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_8VKltBBU2_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_IxdqBATw2_1),.doutc(w_dff_A_CvTLzAgQ6_2),.din(n462));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_dff_A_yQsZz6LY3_2),.din(w_dff_B_c5M0faWB5_3));
	jspl3 jspl3_w_n473_1(.douta(w_dff_A_xwueaaXp8_0),.doutb(w_dff_A_3XYAaoiY3_1),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.doutc(w_n484_0[2]),.din(n484));
	jspl jspl_w_n484_1(.douta(w_n484_1[0]),.doutb(w_n484_1[1]),.din(w_n484_0[0]));
	jspl3 jspl3_w_n486_0(.douta(w_dff_A_1YbHecmV2_0),.doutb(w_n486_0[1]),.doutc(w_dff_A_8RSXgteW1_2),.din(n486));
	jspl jspl_w_n486_1(.douta(w_dff_A_iqc2tmVP1_0),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl3 jspl3_w_n495_1(.douta(w_n495_1[0]),.doutb(w_n495_1[1]),.doutc(w_n495_1[2]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n497_0(.douta(w_dff_A_CQDvDQIN0_0),.doutb(w_n497_0[1]),.doutc(w_dff_A_53wdL9Ic4_2),.din(n497));
	jspl jspl_w_n497_1(.douta(w_dff_A_IwN1l2Xb1_0),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_juMTaES87_2));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl jspl_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl jspl_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_E0EfueVk5_2));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl3 jspl3_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.doutc(w_n541_0[2]),.din(n541));
	jspl jspl_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.din(w_n541_0[0]));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_dff_A_K1sSTTDM4_1),.din(n543));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl jspl_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl jspl_w_n560_1(.douta(w_n560_1[0]),.doutb(w_n560_1[1]),.din(w_n560_0[0]));
	jspl3 jspl3_w_n561_0(.douta(w_dff_A_LT7SfRtI1_0),.doutb(w_dff_A_Q094VyXA8_1),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n562_0(.douta(w_dff_A_YLbN2nBA3_0),.doutb(w_n562_0[1]),.din(w_dff_B_f1SPZpZX8_2));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_dff_A_9WJodyuM8_1),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_dff_A_P8xOK5uz1_1),.din(w_n567_0[0]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_dff_A_SU22FOku6_1),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_dff_A_9prX5OOG0_2),.din(n571));
	jspl jspl_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.din(w_n571_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_dff_A_EXbfzPrL4_0),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_dff_A_nLtBEqxt1_1),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.doutc(w_n582_0[2]),.din(n582));
	jspl jspl_w_n582_1(.douta(w_n582_1[0]),.doutb(w_n582_1[1]),.din(w_n582_0[0]));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_dff_A_OVx7vuIf6_2),.din(n583));
	jspl jspl_w_n583_1(.douta(w_dff_A_bnNVtO9w5_0),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl jspl_w_n585_0(.douta(w_dff_A_ZUHGbJNA8_0),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl jspl_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_dff_A_K7sE6wq35_1),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.din(w_n590_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_nJ2td3iY0_1),.din(n591));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl jspl_w_n595_1(.douta(w_n595_1[0]),.doutb(w_n595_1[1]),.din(w_n595_0[0]));
	jspl3 jspl3_w_n596_0(.douta(w_dff_A_09eiEXdN9_0),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl jspl_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.din(w_n600_0[0]));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_d2qPCzLc6_0),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_vtSVt5Ke4_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n605_2(.douta(w_n605_2[0]),.doutb(w_n605_2[1]),.doutc(w_n605_2[2]),.din(w_n605_0[1]));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_dff_A_bispfRPv1_1),.doutc(w_n607_0[2]),.din(w_dff_B_NxnJO8Er8_3));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.doutc(w_n609_1[2]),.din(w_n609_0[0]));
	jspl3 jspl3_w_n609_2(.douta(w_n609_2[0]),.doutb(w_n609_2[1]),.doutc(w_n609_2[2]),.din(w_n609_0[1]));
	jspl3 jspl3_w_n609_3(.douta(w_n609_3[0]),.doutb(w_n609_3[1]),.doutc(w_n609_3[2]),.din(w_n609_0[2]));
	jspl3 jspl3_w_n609_4(.douta(w_n609_4[0]),.doutb(w_n609_4[1]),.doutc(w_n609_4[2]),.din(w_n609_1[0]));
	jspl3 jspl3_w_n609_5(.douta(w_n609_5[0]),.doutb(w_n609_5[1]),.doutc(w_n609_5[2]),.din(w_n609_1[1]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_dff_A_MGTmNajW1_1),.doutc(w_dff_A_HBGiEuX35_2),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_dff_A_yFlhvwaL7_0),.doutb(w_n614_1[1]),.doutc(w_dff_A_SfMgCxe87_2),.din(w_n614_0[0]));
	jspl jspl_w_n614_2(.douta(w_dff_A_JWom5X3a3_0),.doutb(w_n614_2[1]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n618_1(.douta(w_n618_1[0]),.doutb(w_n618_1[1]),.din(w_n618_0[0]));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n621_1(.douta(w_dff_A_XwwuUsln0_0),.doutb(w_n621_1[1]),.doutc(w_n621_1[2]),.din(w_n621_0[0]));
	jspl jspl_w_n621_2(.douta(w_dff_A_IFsxbyU17_0),.doutb(w_n621_2[1]),.din(w_n621_0[1]));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl jspl_w_n623_0(.douta(w_dff_A_rPjvbile5_0),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl3 jspl3_w_n624_1(.douta(w_n624_1[0]),.doutb(w_n624_1[1]),.doutc(w_n624_1[2]),.din(w_n624_0[0]));
	jspl3 jspl3_w_n625_0(.douta(w_dff_A_PGqWpFTY3_0),.doutb(w_n625_0[1]),.doutc(w_dff_A_ye7KwXvM9_2),.din(n625));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_dff_A_y078HFsd3_1),.doutc(w_n628_0[2]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_dff_A_ArazxxYs6_1),.doutc(w_n629_0[2]),.din(n629));
	jspl jspl_w_n631_0(.douta(w_dff_A_HIdUAKGh5_0),.doutb(w_n631_0[1]),.din(n631));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl jspl_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_dff_A_lDwR0oxZ1_2),.din(n636));
	jspl jspl_w_n636_1(.douta(w_n636_1[0]),.doutb(w_dff_A_YybsqF5R9_1),.din(w_n636_0[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_dff_A_7qnZTphL5_1),.doutc(w_dff_A_m2MJmds47_2),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_dff_A_OwxKxIKB0_0),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl3 jspl3_w_n646_0(.douta(w_dff_A_mdWYaNkU6_0),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.doutc(w_dff_A_MlFFv0D18_2),.din(n649));
	jspl jspl_w_n649_1(.douta(w_n649_1[0]),.doutb(w_n649_1[1]),.din(w_n649_0[0]));
	jspl jspl_w_n650_0(.douta(w_dff_A_KnkyxPvf7_0),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_dff_A_MmFNpZCS8_1),.doutc(w_dff_A_uonOlQ6T0_2),.din(w_dff_B_5M9btRQs8_3));
	jspl jspl_w_n651_1(.douta(w_dff_A_KZ6qEmH77_0),.doutb(w_n651_1[1]),.din(w_n651_0[0]));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_Ly8y0O7P7_2));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n671_0(.douta(w_dff_A_AS70YKql5_0),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_dff_A_cdBdRrEJ6_1),.din(n678));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_dff_A_EeOODEu20_1),.din(n679));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_dff_A_Vpom8c187_1),.din(w_dff_B_97Od1iLj9_2));
	jspl3 jspl3_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.doutc(w_n681_0[2]),.din(n681));
	jspl3 jspl3_w_n681_1(.douta(w_dff_A_j8tzyT2m1_0),.doutb(w_dff_A_jHm2wTS61_1),.doutc(w_n681_1[2]),.din(w_n681_0[0]));
	jspl jspl_w_n681_2(.douta(w_dff_A_CZu92rYw1_0),.doutb(w_n681_2[1]),.din(w_n681_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl3 jspl3_w_n687_0(.douta(w_dff_A_NiKCeGge1_0),.doutb(w_dff_A_EvD6p0zS9_1),.doutc(w_n687_0[2]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_dff_A_JOLCGD738_0),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_dff_A_8v12xvBk6_1),.doutc(w_n691_0[2]),.din(n691));
	jspl3 jspl3_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.doutc(w_n693_0[2]),.din(n693));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.doutc(w_n696_0[2]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_dff_A_HcWZaaDr7_1),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(w_dff_B_yJUIuqCl3_2));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_dff_A_RabxUM5u6_0),.doutb(w_n706_0[1]),.din(n706));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_giZSAE6j8_2));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_HKufdfLD0_1),.doutc(w_dff_A_CKr4KLtG9_2),.din(n717));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl3 jspl3_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_BlrkuVzQ3_1),.doutc(w_n721_0[2]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_dff_A_jDdGjmD57_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl3 jspl3_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.doutc(w_dff_A_FIgmJxWn2_2),.din(n739));
	jspl jspl_w_n739_1(.douta(w_dff_A_yKP8tZG88_0),.doutb(w_n739_1[1]),.din(w_n739_0[0]));
	jspl jspl_w_n740_0(.douta(w_n740_0[0]),.doutb(w_dff_A_kUQDiRdJ1_1),.din(n740));
	jspl jspl_w_n741_0(.douta(w_dff_A_xo8iiHrd0_0),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_2SZsCcUg8_2));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_dff_A_wV0klqvI2_2),.din(w_dff_B_4K1igsW85_3));
	jspl3 jspl3_w_n744_1(.douta(w_dff_A_9oh8lctW9_0),.doutb(w_n744_1[1]),.doutc(w_n744_1[2]),.din(w_n744_0[0]));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_dff_A_xCoe0Yxo1_2),.din(n746));
	jspl3 jspl3_w_n746_1(.douta(w_n746_1[0]),.doutb(w_n746_1[1]),.doutc(w_n746_1[2]),.din(w_n746_0[0]));
	jspl3 jspl3_w_n747_0(.douta(w_dff_A_LoCCPFDQ2_0),.doutb(w_dff_A_Xu5BlIp72_1),.doutc(w_n747_0[2]),.din(n747));
	jspl3 jspl3_w_n747_1(.douta(w_n747_1[0]),.doutb(w_dff_A_VoHkmlRv2_1),.doutc(w_dff_A_PRChFjBw1_2),.din(w_n747_0[0]));
	jspl3 jspl3_w_n747_2(.douta(w_dff_A_Zh3Fzkn12_0),.doutb(w_dff_A_uvpUTQee1_1),.doutc(w_n747_2[2]),.din(w_n747_0[1]));
	jspl3 jspl3_w_n747_3(.douta(w_dff_A_wDe8DPcc0_0),.doutb(w_dff_A_gU6XlNYE1_1),.doutc(w_n747_3[2]),.din(w_n747_0[2]));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_dff_A_UQoh7LGe2_1),.doutc(w_dff_A_a3B1miSq9_2),.din(w_dff_B_qXzrlhWH2_3));
	jspl3 jspl3_w_n748_1(.douta(w_n748_1[0]),.doutb(w_dff_A_FBNMLUe16_1),.doutc(w_dff_A_L5frsO004_2),.din(w_n748_0[0]));
	jspl3 jspl3_w_n748_2(.douta(w_dff_A_q9i9WFuA3_0),.doutb(w_n748_2[1]),.doutc(w_dff_A_YlD1YxIp1_2),.din(w_n748_0[1]));
	jspl3 jspl3_w_n748_3(.douta(w_n748_3[0]),.doutb(w_dff_A_sHOXtqEZ9_1),.doutc(w_dff_A_p1fNNdqi8_2),.din(w_n748_0[2]));
	jspl jspl_w_n748_4(.douta(w_dff_A_zE2BDkb14_0),.doutb(w_n748_4[1]),.din(w_n748_1[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_dff_A_vGWoQ90w7_1),.doutc(w_dff_A_NYquPSHS8_2),.din(n750));
	jspl jspl_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n751_0(.douta(w_dff_A_frt58SoM2_0),.doutb(w_n751_0[1]),.doutc(w_dff_A_PvOiRHAm7_2),.din(n751));
	jspl3 jspl3_w_n751_1(.douta(w_n751_1[0]),.doutb(w_dff_A_7EUgJjEv4_1),.doutc(w_n751_1[2]),.din(w_n751_0[0]));
	jspl jspl_w_n751_2(.douta(w_n751_2[0]),.doutb(w_dff_A_BsgYYTw75_1),.din(w_n751_0[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl3 jspl3_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.doutc(w_n753_1[2]),.din(w_n753_0[0]));
	jspl3 jspl3_w_n753_2(.douta(w_n753_2[0]),.doutb(w_n753_2[1]),.doutc(w_n753_2[2]),.din(w_n753_0[1]));
	jspl3 jspl3_w_n753_3(.douta(w_n753_3[0]),.doutb(w_n753_3[1]),.doutc(w_n753_3[2]),.din(w_n753_0[2]));
	jspl3 jspl3_w_n753_4(.douta(w_n753_4[0]),.doutb(w_n753_4[1]),.doutc(w_n753_4[2]),.din(w_n753_1[0]));
	jspl3 jspl3_w_n753_5(.douta(w_n753_5[0]),.doutb(w_n753_5[1]),.doutc(w_n753_5[2]),.din(w_n753_1[1]));
	jspl3 jspl3_w_n753_6(.douta(w_n753_6[0]),.doutb(w_n753_6[1]),.doutc(w_n753_6[2]),.din(w_n753_1[2]));
	jspl3 jspl3_w_n753_7(.douta(w_n753_7[0]),.doutb(w_n753_7[1]),.doutc(w_n753_7[2]),.din(w_n753_2[0]));
	jspl jspl_w_n753_8(.douta(w_n753_8[0]),.doutb(w_n753_8[1]),.din(w_n753_2[1]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl3 jspl3_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.doutc(w_n765_0[2]),.din(w_dff_B_rUp8ULsw4_3));
	jspl3 jspl3_w_n765_1(.douta(w_n765_1[0]),.doutb(w_n765_1[1]),.doutc(w_n765_1[2]),.din(w_n765_0[0]));
	jspl3 jspl3_w_n765_2(.douta(w_n765_2[0]),.doutb(w_n765_2[1]),.doutc(w_n765_2[2]),.din(w_n765_0[1]));
	jspl3 jspl3_w_n765_3(.douta(w_n765_3[0]),.doutb(w_n765_3[1]),.doutc(w_n765_3[2]),.din(w_n765_0[2]));
	jspl3 jspl3_w_n765_4(.douta(w_n765_4[0]),.doutb(w_n765_4[1]),.doutc(w_n765_4[2]),.din(w_n765_1[0]));
	jspl3 jspl3_w_n765_5(.douta(w_n765_5[0]),.doutb(w_n765_5[1]),.doutc(w_n765_5[2]),.din(w_n765_1[1]));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_dff_A_oxz4LApm0_1),.din(n779));
	jspl3 jspl3_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.doutc(w_n781_0[2]),.din(n781));
	jspl3 jspl3_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.doutc(w_n783_0[2]),.din(n783));
	jspl jspl_w_n783_1(.douta(w_n783_1[0]),.doutb(w_n783_1[1]),.din(w_n783_0[0]));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_G0r8g5BP1_2));
	jspl3 jspl3_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.doutc(w_n789_0[2]),.din(n789));
	jspl3 jspl3_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.doutc(w_n791_0[2]),.din(n791));
	jspl jspl_w_n791_1(.douta(w_n791_1[0]),.doutb(w_n791_1[1]),.din(w_n791_0[0]));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_dff_A_rbDetDgH9_1),.doutc(w_dff_A_4S0qJLoI6_2),.din(w_dff_B_dFN2gYon5_3));
	jspl3 jspl3_w_n793_1(.douta(w_n793_1[0]),.doutb(w_dff_A_xjWfmCDl7_1),.doutc(w_dff_A_S5eA9kuy6_2),.din(w_n793_0[0]));
	jspl3 jspl3_w_n793_2(.douta(w_n793_2[0]),.doutb(w_n793_2[1]),.doutc(w_dff_A_ZgzYrzSU2_2),.din(w_n793_0[1]));
	jspl3 jspl3_w_n793_3(.douta(w_n793_3[0]),.doutb(w_dff_A_8LEd86GY1_1),.doutc(w_dff_A_kG0CDKnq1_2),.din(w_n793_0[2]));
	jspl jspl_w_n793_4(.douta(w_dff_A_pDba1ues0_0),.doutb(w_n793_4[1]),.din(w_n793_1[0]));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_dff_A_MsSSaf845_1),.doutc(w_dff_A_dsfKY5Mi9_2),.din(w_dff_B_XABObqKV1_3));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_dff_A_wr4dtUjX9_1),.doutc(w_dff_A_AJGiieCM9_2),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_dff_A_dkRHlgvt0_2),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_n797_3[0]),.doutb(w_dff_A_Y9bywIRN2_1),.doutc(w_dff_A_rTCJRv862_2),.din(w_n797_0[2]));
	jspl jspl_w_n797_4(.douta(w_dff_A_DrEaSfxY2_0),.doutb(w_n797_4[1]),.din(w_n797_1[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.doutc(w_n799_1[2]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n799_2(.douta(w_n799_2[0]),.doutb(w_n799_2[1]),.doutc(w_n799_2[2]),.din(w_n799_0[1]));
	jspl3 jspl3_w_n799_3(.douta(w_n799_3[0]),.doutb(w_n799_3[1]),.doutc(w_n799_3[2]),.din(w_n799_0[2]));
	jspl jspl_w_n799_4(.douta(w_n799_4[0]),.doutb(w_n799_4[1]),.din(w_n799_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl3 jspl3_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.doutc(w_n801_1[2]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n801_2(.douta(w_n801_2[0]),.doutb(w_n801_2[1]),.doutc(w_n801_2[2]),.din(w_n801_0[1]));
	jspl3 jspl3_w_n801_3(.douta(w_n801_3[0]),.doutb(w_n801_3[1]),.doutc(w_n801_3[2]),.din(w_n801_0[2]));
	jspl jspl_w_n801_4(.douta(w_n801_4[0]),.doutb(w_n801_4[1]),.din(w_n801_1[0]));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl3 jspl3_w_n828_0(.douta(w_n828_0[0]),.doutb(w_dff_A_9p8FwHgm0_1),.doutc(w_dff_A_VZ74eUt02_2),.din(n828));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_dff_A_q39Y62Qo9_1),.din(n829));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl3 jspl3_w_n840_0(.douta(w_n840_0[0]),.doutb(w_dff_A_Yw8dhu3K1_1),.doutc(w_dff_A_1eiEKxGE0_2),.din(w_dff_B_ybEFOdHf6_3));
	jspl3 jspl3_w_n840_1(.douta(w_n840_1[0]),.doutb(w_dff_A_nLzfCQsM7_1),.doutc(w_dff_A_8wZX448Z7_2),.din(w_n840_0[0]));
	jspl3 jspl3_w_n840_2(.douta(w_n840_2[0]),.doutb(w_n840_2[1]),.doutc(w_dff_A_WCC2ZLwE1_2),.din(w_n840_0[1]));
	jspl3 jspl3_w_n840_3(.douta(w_n840_3[0]),.doutb(w_dff_A_2SUQv1QZ1_1),.doutc(w_dff_A_GSoiYBCs5_2),.din(w_n840_0[2]));
	jspl jspl_w_n840_4(.douta(w_dff_A_2YFHNRle2_0),.doutb(w_n840_4[1]),.din(w_n840_1[0]));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_dff_A_kk7zswMP6_1),.doutc(w_dff_A_ETtXIzyY5_2),.din(w_dff_B_YNwcWui00_3));
	jspl3 jspl3_w_n843_1(.douta(w_n843_1[0]),.doutb(w_dff_A_WGJbEyxO9_1),.doutc(w_dff_A_Hwmo3KAh3_2),.din(w_n843_0[0]));
	jspl3 jspl3_w_n843_2(.douta(w_n843_2[0]),.doutb(w_n843_2[1]),.doutc(w_dff_A_YZB8mdmT1_2),.din(w_n843_0[1]));
	jspl3 jspl3_w_n843_3(.douta(w_n843_3[0]),.doutb(w_dff_A_np2aySLL9_1),.doutc(w_dff_A_ILrysShD0_2),.din(w_n843_0[2]));
	jspl jspl_w_n843_4(.douta(w_dff_A_7Ey6VMuo4_0),.doutb(w_n843_4[1]),.din(w_n843_1[0]));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl3 jspl3_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.doutc(w_n845_1[2]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n845_2(.douta(w_n845_2[0]),.doutb(w_n845_2[1]),.doutc(w_n845_2[2]),.din(w_n845_0[1]));
	jspl3 jspl3_w_n845_3(.douta(w_n845_3[0]),.doutb(w_n845_3[1]),.doutc(w_n845_3[2]),.din(w_n845_0[2]));
	jspl jspl_w_n845_4(.douta(w_n845_4[0]),.doutb(w_n845_4[1]),.din(w_n845_1[0]));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl3 jspl3_w_n847_1(.douta(w_n847_1[0]),.doutb(w_n847_1[1]),.doutc(w_n847_1[2]),.din(w_n847_0[0]));
	jspl3 jspl3_w_n847_2(.douta(w_n847_2[0]),.doutb(w_n847_2[1]),.doutc(w_n847_2[2]),.din(w_n847_0[1]));
	jspl3 jspl3_w_n847_3(.douta(w_n847_3[0]),.doutb(w_n847_3[1]),.doutc(w_n847_3[2]),.din(w_n847_0[2]));
	jspl jspl_w_n847_4(.douta(w_n847_4[0]),.doutb(w_n847_4[1]),.din(w_n847_1[0]));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_dff_A_1lupsNG66_1),.din(w_dff_B_kllcc4En5_2));
	jspl jspl_w_n855_0(.douta(w_dff_A_hEsPBp8w3_0),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n928_0(.douta(w_n928_0[0]),.doutb(w_dff_A_pCOCpnTh6_1),.din(w_dff_B_tHW24P2b1_2));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_dff_A_DcNViKZO3_2),.din(w_dff_B_cNCEHzcg0_3));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(w_dff_B_MVJDqufb2_2));
	jspl3 jspl3_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.doutc(w_n936_0[2]),.din(n936));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_dff_A_rc6cyPT01_1),.din(n943));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_dff_A_JiOFjd856_1),.din(n944));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl3 jspl3_w_n948_0(.douta(w_n948_0[0]),.doutb(w_n948_0[1]),.doutc(w_n948_0[2]),.din(n948));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_dff_A_qkS26nqD6_1),.din(w_dff_B_qYv6NP3V6_2));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_dff_A_sUW6gcWQ9_1),.din(n971));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl3 jspl3_w_n985_0(.douta(w_n985_0[0]),.doutb(w_dff_A_RFQeJ0rj8_1),.doutc(w_dff_A_XlHVV9RA6_2),.din(n985));
	jspl3 jspl3_w_n985_1(.douta(w_dff_A_Nky4KSlY5_0),.doutb(w_n985_1[1]),.doutc(w_dff_A_9vZJQ24L1_2),.din(w_n985_0[0]));
	jspl3 jspl3_w_n985_2(.douta(w_dff_A_PHBE6jlE2_0),.doutb(w_dff_A_o45GCSCM4_1),.doutc(w_n985_2[2]),.din(w_n985_0[1]));
	jspl3 jspl3_w_n985_3(.douta(w_dff_A_fCAycZkA0_0),.doutb(w_dff_A_cN4ywjen3_1),.doutc(w_n985_3[2]),.din(w_n985_0[2]));
	jspl jspl_w_n985_4(.douta(w_dff_A_p7tmQuyS8_0),.doutb(w_n985_4[1]),.din(w_n985_1[0]));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_dff_A_q74Muz0Z9_1),.doutc(w_dff_A_srwLQ5c40_2),.din(n988));
	jspl3 jspl3_w_n988_1(.douta(w_dff_A_RS3E63ZZ8_0),.doutb(w_n988_1[1]),.doutc(w_dff_A_WcX8CP5O4_2),.din(w_n988_0[0]));
	jspl3 jspl3_w_n988_2(.douta(w_dff_A_7OW5y9l72_0),.doutb(w_dff_A_l4jMXvw94_1),.doutc(w_n988_2[2]),.din(w_n988_0[1]));
	jspl3 jspl3_w_n988_3(.douta(w_dff_A_dpyfnwzd8_0),.doutb(w_dff_A_SSmOGXFU7_1),.doutc(w_n988_3[2]),.din(w_n988_0[2]));
	jspl jspl_w_n988_4(.douta(w_dff_A_LzgFPlqJ2_0),.doutb(w_n988_4[1]),.din(w_n988_1[0]));
	jspl3 jspl3_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.doutc(w_n990_0[2]),.din(n990));
	jspl3 jspl3_w_n990_1(.douta(w_n990_1[0]),.doutb(w_n990_1[1]),.doutc(w_n990_1[2]),.din(w_n990_0[0]));
	jspl3 jspl3_w_n990_2(.douta(w_n990_2[0]),.doutb(w_n990_2[1]),.doutc(w_n990_2[2]),.din(w_n990_0[1]));
	jspl3 jspl3_w_n990_3(.douta(w_n990_3[0]),.doutb(w_n990_3[1]),.doutc(w_n990_3[2]),.din(w_n990_0[2]));
	jspl jspl_w_n990_4(.douta(w_n990_4[0]),.doutb(w_n990_4[1]),.din(w_n990_1[0]));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n992_2(.douta(w_n992_2[0]),.doutb(w_n992_2[1]),.doutc(w_n992_2[2]),.din(w_n992_0[1]));
	jspl3 jspl3_w_n992_3(.douta(w_n992_3[0]),.doutb(w_n992_3[1]),.doutc(w_n992_3[2]),.din(w_n992_0[2]));
	jspl jspl_w_n992_4(.douta(w_n992_4[0]),.doutb(w_n992_4[1]),.din(w_n992_1[0]));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_YkaaOJ3u5_1),.doutc(w_dff_A_KgaFGU7S5_2),.din(n999));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_rrccWHtp0_0),.doutb(w_n999_1[1]),.doutc(w_dff_A_A9I8q0GE3_2),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_fYU173FL6_0),.doutb(w_dff_A_tjHVlKCN6_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_i86dQOnh2_0),.doutb(w_dff_A_QwZ9RiFX5_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl jspl_w_n999_4(.douta(w_dff_A_a9Qm4DtW7_0),.doutb(w_n999_4[1]),.din(w_n999_1[0]));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_dff_A_32D0wbyv8_1),.doutc(w_dff_A_wXW4sHwz1_2),.din(n1002));
	jspl3 jspl3_w_n1002_1(.douta(w_dff_A_LW7Mt9wV8_0),.doutb(w_n1002_1[1]),.doutc(w_dff_A_IDxTqGVC1_2),.din(w_n1002_0[0]));
	jspl3 jspl3_w_n1002_2(.douta(w_dff_A_H5bf7n1u2_0),.doutb(w_dff_A_ITNR949C7_1),.doutc(w_n1002_2[2]),.din(w_n1002_0[1]));
	jspl3 jspl3_w_n1002_3(.douta(w_dff_A_6mb7RBXC1_0),.doutb(w_dff_A_BCAe3P7R0_1),.doutc(w_n1002_3[2]),.din(w_n1002_0[2]));
	jspl jspl_w_n1002_4(.douta(w_dff_A_kMyjH4IQ1_0),.doutb(w_n1002_4[1]),.din(w_n1002_1[0]));
	jspl3 jspl3_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.doutc(w_n1004_0[2]),.din(n1004));
	jspl3 jspl3_w_n1004_1(.douta(w_n1004_1[0]),.doutb(w_n1004_1[1]),.doutc(w_n1004_1[2]),.din(w_n1004_0[0]));
	jspl3 jspl3_w_n1004_2(.douta(w_n1004_2[0]),.doutb(w_n1004_2[1]),.doutc(w_n1004_2[2]),.din(w_n1004_0[1]));
	jspl3 jspl3_w_n1004_3(.douta(w_n1004_3[0]),.doutb(w_n1004_3[1]),.doutc(w_n1004_3[2]),.din(w_n1004_0[2]));
	jspl jspl_w_n1004_4(.douta(w_n1004_4[0]),.doutb(w_n1004_4[1]),.din(w_n1004_1[0]));
	jspl3 jspl3_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.doutc(w_n1006_0[2]),.din(n1006));
	jspl3 jspl3_w_n1006_1(.douta(w_n1006_1[0]),.doutb(w_n1006_1[1]),.doutc(w_n1006_1[2]),.din(w_n1006_0[0]));
	jspl3 jspl3_w_n1006_2(.douta(w_n1006_2[0]),.doutb(w_n1006_2[1]),.doutc(w_n1006_2[2]),.din(w_n1006_0[1]));
	jspl3 jspl3_w_n1006_3(.douta(w_n1006_3[0]),.doutb(w_n1006_3[1]),.doutc(w_n1006_3[2]),.din(w_n1006_0[2]));
	jspl jspl_w_n1006_4(.douta(w_n1006_4[0]),.doutb(w_n1006_4[1]),.din(w_n1006_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl jspl_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.doutc(w_n1023_0[2]),.din(n1023));
	jspl jspl_w_n1023_1(.douta(w_n1023_1[0]),.doutb(w_n1023_1[1]),.din(w_n1023_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl jspl_w_n1039_1(.douta(w_n1039_1[0]),.doutb(w_n1039_1[1]),.din(w_n1039_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl jspl_w_n1142_0(.douta(w_dff_A_osSimo5V6_0),.doutb(w_n1142_0[1]),.din(n1142));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl3 jspl3_w_n1163_1(.douta(w_n1163_1[0]),.doutb(w_n1163_1[1]),.doutc(w_n1163_1[2]),.din(w_n1163_0[0]));
	jspl3 jspl3_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.doutc(w_n1197_0[2]),.din(n1197));
	jspl3 jspl3_w_n1197_1(.douta(w_n1197_1[0]),.doutb(w_n1197_1[1]),.doutc(w_n1197_1[2]),.din(w_n1197_0[0]));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.doutc(w_n1235_0[2]),.din(n1235));
	jspl jspl_w_n1235_1(.douta(w_n1235_1[0]),.doutb(w_n1235_1[1]),.din(w_n1235_0[0]));
	jspl3 jspl3_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.doutc(w_n1242_0[2]),.din(n1242));
	jspl jspl_w_n1242_1(.douta(w_n1242_1[0]),.doutb(w_n1242_1[1]),.din(w_n1242_0[0]));
	jspl3 jspl3_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.doutc(w_n1244_0[2]),.din(n1244));
	jspl jspl_w_n1244_1(.douta(w_n1244_1[0]),.doutb(w_n1244_1[1]),.din(w_n1244_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl jspl_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1253_1(.douta(w_n1253_1[0]),.doutb(w_n1253_1[1]),.din(w_n1253_0[0]));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1383_0(.douta(w_dff_A_fOBNq5Es2_0),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1391_0(.douta(w_dff_A_2zAA9Umb0_0),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1409_0(.douta(w_dff_A_07bBmpDT9_0),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1411_0(.douta(w_dff_A_yQLIJlPF6_0),.doutb(w_n1411_0[1]),.din(n1411));
	jspl jspl_w_n1421_0(.douta(w_dff_A_dwyuefgZ4_0),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_dff_A_i4tnNOao0_1),.din(n1438));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_dff_A_uP4cssC57_1),.din(n1447));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(n1494));
	jspl jspl_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.din(w_dff_B_otbjf07u4_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(w_dff_B_4ofr7wj29_2));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_bK8R2NEB5_2));
	jspl jspl_w_n1555_0(.douta(w_dff_A_i0edykUa5_0),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_dff_A_zKmaTsBv8_1),.din(n1568));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl3 jspl3_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.doutc(w_n1601_0[2]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_dff_A_lOfGrWq38_1),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(w_dff_B_XDizpPKl7_2));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(w_dff_B_uXGqDPoi2_2));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(w_dff_B_9ka1Ae2n2_2));
	jdff dff_B_XssIjf5V0_1(.din(G136),.dout(w_dff_B_XssIjf5V0_1),.clk(gclk));
	jdff dff_B_Dal5NXoy4_0(.din(G2824),.dout(w_dff_B_Dal5NXoy4_0),.clk(gclk));
	jdff dff_B_Mca1lwmy8_1(.din(n320),.dout(w_dff_B_Mca1lwmy8_1),.clk(gclk));
	jdff dff_B_Fm0mRtxx3_1(.din(n327),.dout(w_dff_B_Fm0mRtxx3_1),.clk(gclk));
	jdff dff_B_D7BgWf7S7_2(.din(n333),.dout(w_dff_B_D7BgWf7S7_2),.clk(gclk));
	jdff dff_B_S57yGqN83_1(.din(n338),.dout(w_dff_B_S57yGqN83_1),.clk(gclk));
	jdff dff_B_fnTBsdyL9_1(.din(n340),.dout(w_dff_B_fnTBsdyL9_1),.clk(gclk));
	jdff dff_B_IrVW51x29_0(.din(n341),.dout(w_dff_B_IrVW51x29_0),.clk(gclk));
	jdff dff_B_KSZfTLzP9_1(.din(G24),.dout(w_dff_B_KSZfTLzP9_1),.clk(gclk));
	jdff dff_B_ODt69OBG6_1(.din(n345),.dout(w_dff_B_ODt69OBG6_1),.clk(gclk));
	jdff dff_B_TiA3PYaH3_0(.din(n346),.dout(w_dff_B_TiA3PYaH3_0),.clk(gclk));
	jdff dff_B_Jfk8n5Ey8_1(.din(G26),.dout(w_dff_B_Jfk8n5Ey8_1),.clk(gclk));
	jdff dff_A_WQWmgh6x2_0(.dout(w_G141_2[0]),.din(w_dff_A_WQWmgh6x2_0),.clk(gclk));
	jdff dff_A_gygGVr8w1_0(.dout(w_dff_A_WQWmgh6x2_0),.din(w_dff_A_gygGVr8w1_0),.clk(gclk));
	jdff dff_A_fB1lmueH0_0(.dout(w_dff_A_gygGVr8w1_0),.din(w_dff_A_fB1lmueH0_0),.clk(gclk));
	jdff dff_A_NRmMTPDk0_0(.dout(w_dff_A_fB1lmueH0_0),.din(w_dff_A_NRmMTPDk0_0),.clk(gclk));
	jdff dff_A_AFxMaLQZ3_1(.dout(w_G141_2[1]),.din(w_dff_A_AFxMaLQZ3_1),.clk(gclk));
	jdff dff_A_9EmKaLaE6_1(.dout(w_dff_A_AFxMaLQZ3_1),.din(w_dff_A_9EmKaLaE6_1),.clk(gclk));
	jdff dff_A_yAeXsPl21_1(.dout(w_dff_A_9EmKaLaE6_1),.din(w_dff_A_yAeXsPl21_1),.clk(gclk));
	jdff dff_A_9tMO6vDT1_1(.dout(w_dff_A_yAeXsPl21_1),.din(w_dff_A_9tMO6vDT1_1),.clk(gclk));
	jdff dff_B_Gkskymn36_1(.din(n350),.dout(w_dff_B_Gkskymn36_1),.clk(gclk));
	jdff dff_B_p9XI6owv5_0(.din(n351),.dout(w_dff_B_p9XI6owv5_0),.clk(gclk));
	jdff dff_B_cVsNJJHb0_1(.din(G79),.dout(w_dff_B_cVsNJJHb0_1),.clk(gclk));
	jdff dff_B_JmCqyBqc5_1(.din(n355),.dout(w_dff_B_JmCqyBqc5_1),.clk(gclk));
	jdff dff_B_aSvu7Tg51_0(.din(n356),.dout(w_dff_B_aSvu7Tg51_0),.clk(gclk));
	jdff dff_B_dEkF10QY7_1(.din(G82),.dout(w_dff_B_dEkF10QY7_1),.clk(gclk));
	jdff dff_A_ZMRpH7Cm0_0(.dout(w_G2358_2[0]),.din(w_dff_A_ZMRpH7Cm0_0),.clk(gclk));
	jdff dff_A_bt1O9L7I5_1(.dout(w_G2358_2[1]),.din(w_dff_A_bt1O9L7I5_1),.clk(gclk));
	jdff dff_A_J13aWE4G7_1(.dout(w_G141_1[1]),.din(w_dff_A_J13aWE4G7_1),.clk(gclk));
	jdff dff_A_tFnwf5qe7_1(.dout(w_dff_A_J13aWE4G7_1),.din(w_dff_A_tFnwf5qe7_1),.clk(gclk));
	jdff dff_A_HybsOoa34_1(.dout(w_dff_A_tFnwf5qe7_1),.din(w_dff_A_HybsOoa34_1),.clk(gclk));
	jdff dff_A_8SuW07jG0_1(.dout(w_dff_A_HybsOoa34_1),.din(w_dff_A_8SuW07jG0_1),.clk(gclk));
	jdff dff_A_ihCZD1qn1_2(.dout(w_G141_1[2]),.din(w_dff_A_ihCZD1qn1_2),.clk(gclk));
	jdff dff_A_zVDY3vDk9_2(.dout(w_dff_A_ihCZD1qn1_2),.din(w_dff_A_zVDY3vDk9_2),.clk(gclk));
	jdff dff_A_MJuLq9HB7_2(.dout(w_dff_A_zVDY3vDk9_2),.din(w_dff_A_MJuLq9HB7_2),.clk(gclk));
	jdff dff_A_a5cZcJOE8_2(.dout(w_dff_A_MJuLq9HB7_2),.din(w_dff_A_a5cZcJOE8_2),.clk(gclk));
	jdff dff_B_WsR53Ip04_1(.din(n384),.dout(w_dff_B_WsR53Ip04_1),.clk(gclk));
	jdff dff_B_3CzV9Jej8_1(.din(w_dff_B_WsR53Ip04_1),.dout(w_dff_B_3CzV9Jej8_1),.clk(gclk));
	jdff dff_B_Nz0flp8Q2_0(.din(n446),.dout(w_dff_B_Nz0flp8Q2_0),.clk(gclk));
	jdff dff_B_pkjSE7L20_1(.din(n483),.dout(w_dff_B_pkjSE7L20_1),.clk(gclk));
	jdff dff_B_kW56YRH88_1(.din(n506),.dout(w_dff_B_kW56YRH88_1),.clk(gclk));
	jdff dff_B_Ly8y0O7P7_2(.din(n652),.dout(w_dff_B_Ly8y0O7P7_2),.clk(gclk));
	jdff dff_B_HmIOfsGO3_2(.din(n709),.dout(w_dff_B_HmIOfsGO3_2),.clk(gclk));
	jdff dff_B_DEkXRBgq2_2(.din(w_dff_B_HmIOfsGO3_2),.dout(w_dff_B_DEkXRBgq2_2),.clk(gclk));
	jdff dff_B_giZSAE6j8_2(.din(w_dff_B_DEkXRBgq2_2),.dout(w_dff_B_giZSAE6j8_2),.clk(gclk));
	jdff dff_B_8PzF9dIk4_1(.din(n698),.dout(w_dff_B_8PzF9dIk4_1),.clk(gclk));
	jdff dff_B_ED7Z7xQZ9_1(.din(w_dff_B_8PzF9dIk4_1),.dout(w_dff_B_ED7Z7xQZ9_1),.clk(gclk));
	jdff dff_B_2WzSiiHc7_1(.din(w_dff_B_ED7Z7xQZ9_1),.dout(w_dff_B_2WzSiiHc7_1),.clk(gclk));
	jdff dff_B_7XrR9Fu38_1(.din(w_dff_B_2WzSiiHc7_1),.dout(w_dff_B_7XrR9Fu38_1),.clk(gclk));
	jdff dff_B_ip7ldRLj3_1(.din(n699),.dout(w_dff_B_ip7ldRLj3_1),.clk(gclk));
	jdff dff_B_ZcvBg8Sc2_1(.din(w_dff_B_ip7ldRLj3_1),.dout(w_dff_B_ZcvBg8Sc2_1),.clk(gclk));
	jdff dff_B_fnflHZ8W5_1(.din(w_dff_B_ZcvBg8Sc2_1),.dout(w_dff_B_fnflHZ8W5_1),.clk(gclk));
	jdff dff_A_hrZEm7iI5_1(.dout(w_n607_0[1]),.din(w_dff_A_hrZEm7iI5_1),.clk(gclk));
	jdff dff_A_bispfRPv1_1(.dout(w_dff_A_hrZEm7iI5_1),.din(w_dff_A_bispfRPv1_1),.clk(gclk));
	jdff dff_B_vZrKh8sv0_3(.din(n607),.dout(w_dff_B_vZrKh8sv0_3),.clk(gclk));
	jdff dff_B_yYpi79nI5_3(.din(w_dff_B_vZrKh8sv0_3),.dout(w_dff_B_yYpi79nI5_3),.clk(gclk));
	jdff dff_B_NxnJO8Er8_3(.din(w_dff_B_yYpi79nI5_3),.dout(w_dff_B_NxnJO8Er8_3),.clk(gclk));
	jdff dff_B_AeDOD12Z9_0(.din(n606),.dout(w_dff_B_AeDOD12Z9_0),.clk(gclk));
	jdff dff_B_whth4iwK4_2(.din(n742),.dout(w_dff_B_whth4iwK4_2),.clk(gclk));
	jdff dff_B_5CtWqWG32_2(.din(w_dff_B_whth4iwK4_2),.dout(w_dff_B_5CtWqWG32_2),.clk(gclk));
	jdff dff_B_f5WSunBa1_2(.din(w_dff_B_5CtWqWG32_2),.dout(w_dff_B_f5WSunBa1_2),.clk(gclk));
	jdff dff_B_YGtMakNp9_2(.din(w_dff_B_f5WSunBa1_2),.dout(w_dff_B_YGtMakNp9_2),.clk(gclk));
	jdff dff_B_2SZsCcUg8_2(.din(w_dff_B_YGtMakNp9_2),.dout(w_dff_B_2SZsCcUg8_2),.clk(gclk));
	jdff dff_A_Z33aOacp4_0(.dout(w_n651_1[0]),.din(w_dff_A_Z33aOacp4_0),.clk(gclk));
	jdff dff_A_QHGVysha6_0(.dout(w_dff_A_Z33aOacp4_0),.din(w_dff_A_QHGVysha6_0),.clk(gclk));
	jdff dff_A_vT0gjAMZ6_0(.dout(w_dff_A_QHGVysha6_0),.din(w_dff_A_vT0gjAMZ6_0),.clk(gclk));
	jdff dff_A_JAk0xbai5_0(.dout(w_dff_A_vT0gjAMZ6_0),.din(w_dff_A_JAk0xbai5_0),.clk(gclk));
	jdff dff_A_IN0CntKv1_0(.dout(w_dff_A_JAk0xbai5_0),.din(w_dff_A_IN0CntKv1_0),.clk(gclk));
	jdff dff_A_KZ6qEmH77_0(.dout(w_dff_A_IN0CntKv1_0),.din(w_dff_A_KZ6qEmH77_0),.clk(gclk));
	jdff dff_B_PhzMjzHb8_0(.din(n803),.dout(w_dff_B_PhzMjzHb8_0),.clk(gclk));
	jdff dff_B_fBDCGOM50_0(.din(w_dff_B_PhzMjzHb8_0),.dout(w_dff_B_fBDCGOM50_0),.clk(gclk));
	jdff dff_B_rGxtK9wi5_0(.din(w_dff_B_fBDCGOM50_0),.dout(w_dff_B_rGxtK9wi5_0),.clk(gclk));
	jdff dff_B_ph7LqdJY4_0(.din(w_dff_B_rGxtK9wi5_0),.dout(w_dff_B_ph7LqdJY4_0),.clk(gclk));
	jdff dff_B_3ewiIPnx2_0(.din(w_dff_B_ph7LqdJY4_0),.dout(w_dff_B_3ewiIPnx2_0),.clk(gclk));
	jdff dff_B_viMLJl540_0(.din(n802),.dout(w_dff_B_viMLJl540_0),.clk(gclk));
	jdff dff_B_b35jbf2Z3_0(.din(n849),.dout(w_dff_B_b35jbf2Z3_0),.clk(gclk));
	jdff dff_B_zpGI0mAt6_0(.din(w_dff_B_b35jbf2Z3_0),.dout(w_dff_B_zpGI0mAt6_0),.clk(gclk));
	jdff dff_B_nQPXoJiJ7_0(.din(w_dff_B_zpGI0mAt6_0),.dout(w_dff_B_nQPXoJiJ7_0),.clk(gclk));
	jdff dff_B_rgBzz1bG1_0(.din(w_dff_B_nQPXoJiJ7_0),.dout(w_dff_B_rgBzz1bG1_0),.clk(gclk));
	jdff dff_B_U2olVBQR0_0(.din(w_dff_B_rgBzz1bG1_0),.dout(w_dff_B_U2olVBQR0_0),.clk(gclk));
	jdff dff_B_yMh7HUE44_0(.din(n848),.dout(w_dff_B_yMh7HUE44_0),.clk(gclk));
	jdff dff_B_MZhMwQa67_2(.din(G61),.dout(w_dff_B_MZhMwQa67_2),.clk(gclk));
	jdff dff_B_5X48FtVM3_2(.din(G11),.dout(w_dff_B_5X48FtVM3_2),.clk(gclk));
	jdff dff_B_CChcr1BA4_2(.din(w_dff_B_5X48FtVM3_2),.dout(w_dff_B_CChcr1BA4_2),.clk(gclk));
	jdff dff_B_bXABOWnN9_0(.din(n964),.dout(w_dff_B_bXABOWnN9_0),.clk(gclk));
	jdff dff_B_W2wYqFAe1_0(.din(n962),.dout(w_dff_B_W2wYqFAe1_0),.clk(gclk));
	jdff dff_B_KaCYtSDu2_0(.din(n961),.dout(w_dff_B_KaCYtSDu2_0),.clk(gclk));
	jdff dff_B_IrpWIMHD3_1(.din(n957),.dout(w_dff_B_IrpWIMHD3_1),.clk(gclk));
	jdff dff_B_EhSDyr2c9_1(.din(w_dff_B_IrpWIMHD3_1),.dout(w_dff_B_EhSDyr2c9_1),.clk(gclk));
	jdff dff_B_InlKldaq1_1(.din(w_dff_B_EhSDyr2c9_1),.dout(w_dff_B_InlKldaq1_1),.clk(gclk));
	jdff dff_B_3wJGaPeF1_1(.din(w_dff_B_InlKldaq1_1),.dout(w_dff_B_3wJGaPeF1_1),.clk(gclk));
	jdff dff_B_WESzWxWL2_0(.din(n980),.dout(w_dff_B_WESzWxWL2_0),.clk(gclk));
	jdff dff_B_mSFnHuVU1_0(.din(w_dff_B_WESzWxWL2_0),.dout(w_dff_B_mSFnHuVU1_0),.clk(gclk));
	jdff dff_B_mAUt7xJU8_0(.din(n979),.dout(w_dff_B_mAUt7xJU8_0),.clk(gclk));
	jdff dff_B_tjDkCpYo4_0(.din(n978),.dout(w_dff_B_tjDkCpYo4_0),.clk(gclk));
	jdff dff_B_wAe7Cz920_0(.din(n977),.dout(w_dff_B_wAe7Cz920_0),.clk(gclk));
	jdff dff_B_DEajMSUz6_0(.din(n976),.dout(w_dff_B_DEajMSUz6_0),.clk(gclk));
	jdff dff_B_99g6zTEi2_0(.din(n994),.dout(w_dff_B_99g6zTEi2_0),.clk(gclk));
	jdff dff_B_1qYgqFH83_0(.din(w_dff_B_99g6zTEi2_0),.dout(w_dff_B_1qYgqFH83_0),.clk(gclk));
	jdff dff_B_RAli3rd30_0(.din(w_dff_B_1qYgqFH83_0),.dout(w_dff_B_RAli3rd30_0),.clk(gclk));
	jdff dff_B_0MqjEfGd0_0(.din(w_dff_B_RAli3rd30_0),.dout(w_dff_B_0MqjEfGd0_0),.clk(gclk));
	jdff dff_B_8OjgUUdK4_0(.din(w_dff_B_0MqjEfGd0_0),.dout(w_dff_B_8OjgUUdK4_0),.clk(gclk));
	jdff dff_B_yzSYTJWf6_0(.din(n993),.dout(w_dff_B_yzSYTJWf6_0),.clk(gclk));
	jdff dff_B_R7asPy7h5_0(.din(n1008),.dout(w_dff_B_R7asPy7h5_0),.clk(gclk));
	jdff dff_B_M9SHpA5H4_0(.din(w_dff_B_R7asPy7h5_0),.dout(w_dff_B_M9SHpA5H4_0),.clk(gclk));
	jdff dff_B_fSRNsPI46_0(.din(w_dff_B_M9SHpA5H4_0),.dout(w_dff_B_fSRNsPI46_0),.clk(gclk));
	jdff dff_B_XV3u2wTd0_0(.din(w_dff_B_fSRNsPI46_0),.dout(w_dff_B_XV3u2wTd0_0),.clk(gclk));
	jdff dff_B_avY0gwYw0_0(.din(w_dff_B_XV3u2wTd0_0),.dout(w_dff_B_avY0gwYw0_0),.clk(gclk));
	jdff dff_B_6TjWitqE6_0(.din(n1007),.dout(w_dff_B_6TjWitqE6_0),.clk(gclk));
	jdff dff_B_E8Ow1mSb0_2(.din(G185),.dout(w_dff_B_E8Ow1mSb0_2),.clk(gclk));
	jdff dff_B_mg0MgxRV1_2(.din(G182),.dout(w_dff_B_mg0MgxRV1_2),.clk(gclk));
	jdff dff_B_uQNPPLHu0_2(.din(w_dff_B_mg0MgxRV1_2),.dout(w_dff_B_uQNPPLHu0_2),.clk(gclk));
	jdff dff_B_wwrx8AHY9_1(.din(n749),.dout(w_dff_B_wwrx8AHY9_1),.clk(gclk));
	jdff dff_B_B227RsBo4_0(.din(n754),.dout(w_dff_B_B227RsBo4_0),.clk(gclk));
	jdff dff_B_xFtzP4mP1_1(.din(G131),.dout(w_dff_B_xFtzP4mP1_1),.clk(gclk));
	jdff dff_B_QRg1MG1I3_1(.din(w_dff_B_xFtzP4mP1_1),.dout(w_dff_B_QRg1MG1I3_1),.clk(gclk));
	jdff dff_B_CzAGbBpC4_0(.din(n776),.dout(w_dff_B_CzAGbBpC4_0),.clk(gclk));
	jdff dff_B_33JdFQzd1_0(.din(w_dff_B_CzAGbBpC4_0),.dout(w_dff_B_33JdFQzd1_0),.clk(gclk));
	jdff dff_B_plweYquy5_1(.din(G117),.dout(w_dff_B_plweYquy5_1),.clk(gclk));
	jdff dff_B_gUgiBgL93_1(.din(w_dff_B_plweYquy5_1),.dout(w_dff_B_gUgiBgL93_1),.clk(gclk));
	jdff dff_B_qPKMQyte9_0(.din(n504),.dout(w_dff_B_qPKMQyte9_0),.clk(gclk));
	jdff dff_B_KjOV1hzk1_1(.din(n496),.dout(w_dff_B_KjOV1hzk1_1),.clk(gclk));
	jdff dff_B_47TbZlIf2_0(.din(n1019),.dout(w_dff_B_47TbZlIf2_0),.clk(gclk));
	jdff dff_B_4FPXO9oq2_0(.din(n1018),.dout(w_dff_B_4FPXO9oq2_0),.clk(gclk));
	jdff dff_B_9do6CGYe5_0(.din(w_dff_B_4FPXO9oq2_0),.dout(w_dff_B_9do6CGYe5_0),.clk(gclk));
	jdff dff_B_DK7afoQR6_0(.din(w_dff_B_9do6CGYe5_0),.dout(w_dff_B_DK7afoQR6_0),.clk(gclk));
	jdff dff_B_FWWB7Nqj3_0(.din(w_dff_B_DK7afoQR6_0),.dout(w_dff_B_FWWB7Nqj3_0),.clk(gclk));
	jdff dff_B_PEUGs7Ix9_0(.din(w_dff_B_FWWB7Nqj3_0),.dout(w_dff_B_PEUGs7Ix9_0),.clk(gclk));
	jdff dff_B_CygcLcqT8_0(.din(w_dff_B_PEUGs7Ix9_0),.dout(w_dff_B_CygcLcqT8_0),.clk(gclk));
	jdff dff_B_piNr54hs0_0(.din(w_dff_B_CygcLcqT8_0),.dout(w_dff_B_piNr54hs0_0),.clk(gclk));
	jdff dff_B_JYeiFR921_0(.din(w_dff_B_piNr54hs0_0),.dout(w_dff_B_JYeiFR921_0),.clk(gclk));
	jdff dff_B_Rv5YJH7z6_0(.din(w_dff_B_JYeiFR921_0),.dout(w_dff_B_Rv5YJH7z6_0),.clk(gclk));
	jdff dff_B_vn7svMmu9_0(.din(w_dff_B_Rv5YJH7z6_0),.dout(w_dff_B_vn7svMmu9_0),.clk(gclk));
	jdff dff_B_BAeuSWTx6_0(.din(w_dff_B_vn7svMmu9_0),.dout(w_dff_B_BAeuSWTx6_0),.clk(gclk));
	jdff dff_B_ztWLRg0X4_0(.din(w_dff_B_BAeuSWTx6_0),.dout(w_dff_B_ztWLRg0X4_0),.clk(gclk));
	jdff dff_B_Ww6v3SSi1_0(.din(n1017),.dout(w_dff_B_Ww6v3SSi1_0),.clk(gclk));
	jdff dff_A_q3zLCPm63_0(.dout(w_n797_4[0]),.din(w_dff_A_q3zLCPm63_0),.clk(gclk));
	jdff dff_A_A48mdAmP4_0(.dout(w_dff_A_q3zLCPm63_0),.din(w_dff_A_A48mdAmP4_0),.clk(gclk));
	jdff dff_A_LvF52s4v5_0(.dout(w_dff_A_A48mdAmP4_0),.din(w_dff_A_LvF52s4v5_0),.clk(gclk));
	jdff dff_A_a47M2xaZ7_0(.dout(w_dff_A_LvF52s4v5_0),.din(w_dff_A_a47M2xaZ7_0),.clk(gclk));
	jdff dff_A_ZgPCGr6Y6_0(.dout(w_dff_A_a47M2xaZ7_0),.din(w_dff_A_ZgPCGr6Y6_0),.clk(gclk));
	jdff dff_A_fcQliiep9_0(.dout(w_dff_A_ZgPCGr6Y6_0),.din(w_dff_A_fcQliiep9_0),.clk(gclk));
	jdff dff_A_DrEaSfxY2_0(.dout(w_dff_A_fcQliiep9_0),.din(w_dff_A_DrEaSfxY2_0),.clk(gclk));
	jdff dff_A_3dQy5vFe3_0(.dout(w_n793_4[0]),.din(w_dff_A_3dQy5vFe3_0),.clk(gclk));
	jdff dff_A_xq15hH6Z1_0(.dout(w_dff_A_3dQy5vFe3_0),.din(w_dff_A_xq15hH6Z1_0),.clk(gclk));
	jdff dff_A_cvnKx47M1_0(.dout(w_dff_A_xq15hH6Z1_0),.din(w_dff_A_cvnKx47M1_0),.clk(gclk));
	jdff dff_A_Uwkh47Si4_0(.dout(w_dff_A_cvnKx47M1_0),.din(w_dff_A_Uwkh47Si4_0),.clk(gclk));
	jdff dff_A_sJx77pRG2_0(.dout(w_dff_A_Uwkh47Si4_0),.din(w_dff_A_sJx77pRG2_0),.clk(gclk));
	jdff dff_A_VC7dsWwV8_0(.dout(w_dff_A_sJx77pRG2_0),.din(w_dff_A_VC7dsWwV8_0),.clk(gclk));
	jdff dff_A_m61YsGgv0_0(.dout(w_dff_A_VC7dsWwV8_0),.din(w_dff_A_m61YsGgv0_0),.clk(gclk));
	jdff dff_A_pDba1ues0_0(.dout(w_dff_A_m61YsGgv0_0),.din(w_dff_A_pDba1ues0_0),.clk(gclk));
	jdff dff_B_4QTYj42L0_0(.din(n1028),.dout(w_dff_B_4QTYj42L0_0),.clk(gclk));
	jdff dff_B_CYoRH7bO6_0(.din(n1027),.dout(w_dff_B_CYoRH7bO6_0),.clk(gclk));
	jdff dff_B_8sSrWfTZ6_0(.din(w_dff_B_CYoRH7bO6_0),.dout(w_dff_B_8sSrWfTZ6_0),.clk(gclk));
	jdff dff_B_8w1o0Pwi9_0(.din(w_dff_B_8sSrWfTZ6_0),.dout(w_dff_B_8w1o0Pwi9_0),.clk(gclk));
	jdff dff_B_bvSipQJx4_0(.din(w_dff_B_8w1o0Pwi9_0),.dout(w_dff_B_bvSipQJx4_0),.clk(gclk));
	jdff dff_B_c7m6rXMD7_0(.din(w_dff_B_bvSipQJx4_0),.dout(w_dff_B_c7m6rXMD7_0),.clk(gclk));
	jdff dff_B_m58G5xzA9_0(.din(w_dff_B_c7m6rXMD7_0),.dout(w_dff_B_m58G5xzA9_0),.clk(gclk));
	jdff dff_B_4fJtjy4U4_0(.din(w_dff_B_m58G5xzA9_0),.dout(w_dff_B_4fJtjy4U4_0),.clk(gclk));
	jdff dff_B_CDytwPxH1_0(.din(w_dff_B_4fJtjy4U4_0),.dout(w_dff_B_CDytwPxH1_0),.clk(gclk));
	jdff dff_B_rwa9BTLw4_0(.din(w_dff_B_CDytwPxH1_0),.dout(w_dff_B_rwa9BTLw4_0),.clk(gclk));
	jdff dff_B_gz8CIbCF7_0(.din(w_dff_B_rwa9BTLw4_0),.dout(w_dff_B_gz8CIbCF7_0),.clk(gclk));
	jdff dff_B_jHgqreCB4_0(.din(n1026),.dout(w_dff_B_jHgqreCB4_0),.clk(gclk));
	jdff dff_B_QIFUOnRh2_0(.din(n1037),.dout(w_dff_B_QIFUOnRh2_0),.clk(gclk));
	jdff dff_B_syxrlt572_0(.din(w_dff_B_QIFUOnRh2_0),.dout(w_dff_B_syxrlt572_0),.clk(gclk));
	jdff dff_B_ZkBOZRCt1_0(.din(n1036),.dout(w_dff_B_ZkBOZRCt1_0),.clk(gclk));
	jdff dff_B_Kmqbff6M7_0(.din(w_dff_B_ZkBOZRCt1_0),.dout(w_dff_B_Kmqbff6M7_0),.clk(gclk));
	jdff dff_B_blFGw6jZ5_0(.din(w_dff_B_Kmqbff6M7_0),.dout(w_dff_B_blFGw6jZ5_0),.clk(gclk));
	jdff dff_B_e5WHWo593_0(.din(w_dff_B_blFGw6jZ5_0),.dout(w_dff_B_e5WHWo593_0),.clk(gclk));
	jdff dff_B_7ZzqMHBu9_0(.din(w_dff_B_e5WHWo593_0),.dout(w_dff_B_7ZzqMHBu9_0),.clk(gclk));
	jdff dff_B_XbiAhNVy0_0(.din(w_dff_B_7ZzqMHBu9_0),.dout(w_dff_B_XbiAhNVy0_0),.clk(gclk));
	jdff dff_B_P6BvjMBa8_0(.din(w_dff_B_XbiAhNVy0_0),.dout(w_dff_B_P6BvjMBa8_0),.clk(gclk));
	jdff dff_B_45NXoFSz2_0(.din(w_dff_B_P6BvjMBa8_0),.dout(w_dff_B_45NXoFSz2_0),.clk(gclk));
	jdff dff_B_gOnz1Z622_0(.din(n1035),.dout(w_dff_B_gOnz1Z622_0),.clk(gclk));
	jdff dff_B_zng9M7Sd3_0(.din(n1046),.dout(w_dff_B_zng9M7Sd3_0),.clk(gclk));
	jdff dff_B_KQnOpBxn5_0(.din(w_dff_B_zng9M7Sd3_0),.dout(w_dff_B_KQnOpBxn5_0),.clk(gclk));
	jdff dff_B_fvPzOQNK9_0(.din(w_dff_B_KQnOpBxn5_0),.dout(w_dff_B_fvPzOQNK9_0),.clk(gclk));
	jdff dff_B_KLoCxCNO9_0(.din(n1045),.dout(w_dff_B_KLoCxCNO9_0),.clk(gclk));
	jdff dff_B_5xcSTM5P5_0(.din(w_dff_B_KLoCxCNO9_0),.dout(w_dff_B_5xcSTM5P5_0),.clk(gclk));
	jdff dff_B_fdVVnm3y2_0(.din(w_dff_B_5xcSTM5P5_0),.dout(w_dff_B_fdVVnm3y2_0),.clk(gclk));
	jdff dff_B_KEyaKCrz6_0(.din(w_dff_B_fdVVnm3y2_0),.dout(w_dff_B_KEyaKCrz6_0),.clk(gclk));
	jdff dff_B_MDnUbVep0_0(.din(w_dff_B_KEyaKCrz6_0),.dout(w_dff_B_MDnUbVep0_0),.clk(gclk));
	jdff dff_B_zRMVweWr4_0(.din(w_dff_B_MDnUbVep0_0),.dout(w_dff_B_zRMVweWr4_0),.clk(gclk));
	jdff dff_B_04HM0IyZ8_0(.din(n1044),.dout(w_dff_B_04HM0IyZ8_0),.clk(gclk));
	jdff dff_A_Oc0bOI7p6_1(.dout(w_n797_3[1]),.din(w_dff_A_Oc0bOI7p6_1),.clk(gclk));
	jdff dff_A_Y9bywIRN2_1(.dout(w_dff_A_Oc0bOI7p6_1),.din(w_dff_A_Y9bywIRN2_1),.clk(gclk));
	jdff dff_A_ZwpPDw3o7_2(.dout(w_n797_3[2]),.din(w_dff_A_ZwpPDw3o7_2),.clk(gclk));
	jdff dff_A_5SOsB5WF6_2(.dout(w_dff_A_ZwpPDw3o7_2),.din(w_dff_A_5SOsB5WF6_2),.clk(gclk));
	jdff dff_A_8pRe6LkT2_2(.dout(w_dff_A_5SOsB5WF6_2),.din(w_dff_A_8pRe6LkT2_2),.clk(gclk));
	jdff dff_A_rTCJRv862_2(.dout(w_dff_A_8pRe6LkT2_2),.din(w_dff_A_rTCJRv862_2),.clk(gclk));
	jdff dff_A_8LEd86GY1_1(.dout(w_n793_3[1]),.din(w_dff_A_8LEd86GY1_1),.clk(gclk));
	jdff dff_A_eHXEDivT4_2(.dout(w_n793_3[2]),.din(w_dff_A_eHXEDivT4_2),.clk(gclk));
	jdff dff_A_kG0CDKnq1_2(.dout(w_dff_A_eHXEDivT4_2),.din(w_dff_A_kG0CDKnq1_2),.clk(gclk));
	jdff dff_B_lpijphA11_0(.din(n1053),.dout(w_dff_B_lpijphA11_0),.clk(gclk));
	jdff dff_B_GYqsEJOj8_0(.din(n1052),.dout(w_dff_B_GYqsEJOj8_0),.clk(gclk));
	jdff dff_B_i6JhRNwU6_0(.din(w_dff_B_GYqsEJOj8_0),.dout(w_dff_B_i6JhRNwU6_0),.clk(gclk));
	jdff dff_B_gmAs5Kix2_0(.din(w_dff_B_i6JhRNwU6_0),.dout(w_dff_B_gmAs5Kix2_0),.clk(gclk));
	jdff dff_B_jBIxtsFT1_0(.din(w_dff_B_gmAs5Kix2_0),.dout(w_dff_B_jBIxtsFT1_0),.clk(gclk));
	jdff dff_B_7CYsb0fn5_0(.din(w_dff_B_jBIxtsFT1_0),.dout(w_dff_B_7CYsb0fn5_0),.clk(gclk));
	jdff dff_B_WgB243ov3_0(.din(w_dff_B_7CYsb0fn5_0),.dout(w_dff_B_WgB243ov3_0),.clk(gclk));
	jdff dff_B_VRcPIPAr5_0(.din(w_dff_B_WgB243ov3_0),.dout(w_dff_B_VRcPIPAr5_0),.clk(gclk));
	jdff dff_B_0IPoP4RU7_0(.din(w_dff_B_VRcPIPAr5_0),.dout(w_dff_B_0IPoP4RU7_0),.clk(gclk));
	jdff dff_B_gq8X0Bec3_0(.din(w_dff_B_0IPoP4RU7_0),.dout(w_dff_B_gq8X0Bec3_0),.clk(gclk));
	jdff dff_B_CLUWGzWf2_0(.din(w_dff_B_gq8X0Bec3_0),.dout(w_dff_B_CLUWGzWf2_0),.clk(gclk));
	jdff dff_B_J9GBjOcs0_0(.din(w_dff_B_CLUWGzWf2_0),.dout(w_dff_B_J9GBjOcs0_0),.clk(gclk));
	jdff dff_B_IqO4jrNW8_0(.din(w_dff_B_J9GBjOcs0_0),.dout(w_dff_B_IqO4jrNW8_0),.clk(gclk));
	jdff dff_B_JUusCXk67_0(.din(n1051),.dout(w_dff_B_JUusCXk67_0),.clk(gclk));
	jdff dff_B_S7J5IsmI3_2(.din(G37),.dout(w_dff_B_S7J5IsmI3_2),.clk(gclk));
	jdff dff_B_Rli16P8U4_2(.din(G43),.dout(w_dff_B_Rli16P8U4_2),.clk(gclk));
	jdff dff_B_dxC1OtnG9_2(.din(w_dff_B_Rli16P8U4_2),.dout(w_dff_B_dxC1OtnG9_2),.clk(gclk));
	jdff dff_A_H9e2wXoZ0_0(.dout(w_n843_4[0]),.din(w_dff_A_H9e2wXoZ0_0),.clk(gclk));
	jdff dff_A_4VNwIuYC1_0(.dout(w_dff_A_H9e2wXoZ0_0),.din(w_dff_A_4VNwIuYC1_0),.clk(gclk));
	jdff dff_A_mhPKSX9G0_0(.dout(w_dff_A_4VNwIuYC1_0),.din(w_dff_A_mhPKSX9G0_0),.clk(gclk));
	jdff dff_A_00N8qH0f4_0(.dout(w_dff_A_mhPKSX9G0_0),.din(w_dff_A_00N8qH0f4_0),.clk(gclk));
	jdff dff_A_6Rxdd2bt0_0(.dout(w_dff_A_00N8qH0f4_0),.din(w_dff_A_6Rxdd2bt0_0),.clk(gclk));
	jdff dff_A_P2fmNh136_0(.dout(w_dff_A_6Rxdd2bt0_0),.din(w_dff_A_P2fmNh136_0),.clk(gclk));
	jdff dff_A_7Ey6VMuo4_0(.dout(w_dff_A_P2fmNh136_0),.din(w_dff_A_7Ey6VMuo4_0),.clk(gclk));
	jdff dff_A_rBWeQVvN4_0(.dout(w_n840_4[0]),.din(w_dff_A_rBWeQVvN4_0),.clk(gclk));
	jdff dff_A_wE6aJrTb1_0(.dout(w_dff_A_rBWeQVvN4_0),.din(w_dff_A_wE6aJrTb1_0),.clk(gclk));
	jdff dff_A_h3x6bsEl5_0(.dout(w_dff_A_wE6aJrTb1_0),.din(w_dff_A_h3x6bsEl5_0),.clk(gclk));
	jdff dff_A_sgNgf0vX6_0(.dout(w_dff_A_h3x6bsEl5_0),.din(w_dff_A_sgNgf0vX6_0),.clk(gclk));
	jdff dff_A_waHlxvN38_0(.dout(w_dff_A_sgNgf0vX6_0),.din(w_dff_A_waHlxvN38_0),.clk(gclk));
	jdff dff_A_pamI7Pxv1_0(.dout(w_dff_A_waHlxvN38_0),.din(w_dff_A_pamI7Pxv1_0),.clk(gclk));
	jdff dff_A_6f9epyeH3_0(.dout(w_dff_A_pamI7Pxv1_0),.din(w_dff_A_6f9epyeH3_0),.clk(gclk));
	jdff dff_A_2YFHNRle2_0(.dout(w_dff_A_6f9epyeH3_0),.din(w_dff_A_2YFHNRle2_0),.clk(gclk));
	jdff dff_B_tm7n7pgN3_0(.din(n1060),.dout(w_dff_B_tm7n7pgN3_0),.clk(gclk));
	jdff dff_B_spxeXEEB7_0(.din(n1059),.dout(w_dff_B_spxeXEEB7_0),.clk(gclk));
	jdff dff_B_B0H0h72i4_0(.din(w_dff_B_spxeXEEB7_0),.dout(w_dff_B_B0H0h72i4_0),.clk(gclk));
	jdff dff_B_StLHkQiI3_0(.din(w_dff_B_B0H0h72i4_0),.dout(w_dff_B_StLHkQiI3_0),.clk(gclk));
	jdff dff_B_3PaLHpKP9_0(.din(w_dff_B_StLHkQiI3_0),.dout(w_dff_B_3PaLHpKP9_0),.clk(gclk));
	jdff dff_B_euwC8bRQ4_0(.din(w_dff_B_3PaLHpKP9_0),.dout(w_dff_B_euwC8bRQ4_0),.clk(gclk));
	jdff dff_B_PJQewawI0_0(.din(w_dff_B_euwC8bRQ4_0),.dout(w_dff_B_PJQewawI0_0),.clk(gclk));
	jdff dff_B_DDX5Fy4I6_0(.din(w_dff_B_PJQewawI0_0),.dout(w_dff_B_DDX5Fy4I6_0),.clk(gclk));
	jdff dff_B_NqcF3pch4_0(.din(w_dff_B_DDX5Fy4I6_0),.dout(w_dff_B_NqcF3pch4_0),.clk(gclk));
	jdff dff_B_Je3HVV2R8_0(.din(w_dff_B_NqcF3pch4_0),.dout(w_dff_B_Je3HVV2R8_0),.clk(gclk));
	jdff dff_B_e9AgWHTM3_0(.din(w_dff_B_Je3HVV2R8_0),.dout(w_dff_B_e9AgWHTM3_0),.clk(gclk));
	jdff dff_B_bMwGzXBW6_0(.din(n1058),.dout(w_dff_B_bMwGzXBW6_0),.clk(gclk));
	jdff dff_B_ntYLpOYK3_2(.din(G20),.dout(w_dff_B_ntYLpOYK3_2),.clk(gclk));
	jdff dff_B_K85BdsWi9_2(.din(G76),.dout(w_dff_B_K85BdsWi9_2),.clk(gclk));
	jdff dff_B_l3xCiwCo2_2(.din(w_dff_B_K85BdsWi9_2),.dout(w_dff_B_l3xCiwCo2_2),.clk(gclk));
	jdff dff_B_XCDHoueb2_0(.din(n1067),.dout(w_dff_B_XCDHoueb2_0),.clk(gclk));
	jdff dff_B_TErgr8ko2_0(.din(w_dff_B_XCDHoueb2_0),.dout(w_dff_B_TErgr8ko2_0),.clk(gclk));
	jdff dff_B_unBvVqnu6_0(.din(n1066),.dout(w_dff_B_unBvVqnu6_0),.clk(gclk));
	jdff dff_B_D9SjgIIo7_0(.din(w_dff_B_unBvVqnu6_0),.dout(w_dff_B_D9SjgIIo7_0),.clk(gclk));
	jdff dff_B_ajTPpUqU0_0(.din(w_dff_B_D9SjgIIo7_0),.dout(w_dff_B_ajTPpUqU0_0),.clk(gclk));
	jdff dff_B_hQ1ZOIEw6_0(.din(w_dff_B_ajTPpUqU0_0),.dout(w_dff_B_hQ1ZOIEw6_0),.clk(gclk));
	jdff dff_B_sgHFWcFo8_0(.din(w_dff_B_hQ1ZOIEw6_0),.dout(w_dff_B_sgHFWcFo8_0),.clk(gclk));
	jdff dff_B_JyGP5icQ1_0(.din(w_dff_B_sgHFWcFo8_0),.dout(w_dff_B_JyGP5icQ1_0),.clk(gclk));
	jdff dff_B_u5lrbKGc5_0(.din(w_dff_B_JyGP5icQ1_0),.dout(w_dff_B_u5lrbKGc5_0),.clk(gclk));
	jdff dff_B_TKf1DxH57_0(.din(w_dff_B_u5lrbKGc5_0),.dout(w_dff_B_TKf1DxH57_0),.clk(gclk));
	jdff dff_B_NwksgsXy5_0(.din(n1065),.dout(w_dff_B_NwksgsXy5_0),.clk(gclk));
	jdff dff_B_JPVxV5JX3_2(.din(G17),.dout(w_dff_B_JPVxV5JX3_2),.clk(gclk));
	jdff dff_B_41uG2RLG8_2(.din(G73),.dout(w_dff_B_41uG2RLG8_2),.clk(gclk));
	jdff dff_B_SAJzS6I19_2(.din(w_dff_B_41uG2RLG8_2),.dout(w_dff_B_SAJzS6I19_2),.clk(gclk));
	jdff dff_B_DMJtnIM71_0(.din(n1074),.dout(w_dff_B_DMJtnIM71_0),.clk(gclk));
	jdff dff_B_nyxe27eH1_0(.din(w_dff_B_DMJtnIM71_0),.dout(w_dff_B_nyxe27eH1_0),.clk(gclk));
	jdff dff_B_J3jcYmM34_0(.din(w_dff_B_nyxe27eH1_0),.dout(w_dff_B_J3jcYmM34_0),.clk(gclk));
	jdff dff_B_O7THjFWr7_0(.din(n1073),.dout(w_dff_B_O7THjFWr7_0),.clk(gclk));
	jdff dff_B_GaElTtFk0_0(.din(w_dff_B_O7THjFWr7_0),.dout(w_dff_B_GaElTtFk0_0),.clk(gclk));
	jdff dff_B_dIDC2yNE2_0(.din(w_dff_B_GaElTtFk0_0),.dout(w_dff_B_dIDC2yNE2_0),.clk(gclk));
	jdff dff_B_Mb9koHU65_0(.din(w_dff_B_dIDC2yNE2_0),.dout(w_dff_B_Mb9koHU65_0),.clk(gclk));
	jdff dff_B_NBwEMJkl1_0(.din(w_dff_B_Mb9koHU65_0),.dout(w_dff_B_NBwEMJkl1_0),.clk(gclk));
	jdff dff_B_QKeZNlHr6_0(.din(w_dff_B_NBwEMJkl1_0),.dout(w_dff_B_QKeZNlHr6_0),.clk(gclk));
	jdff dff_B_TZ3jdvfl1_0(.din(n1072),.dout(w_dff_B_TZ3jdvfl1_0),.clk(gclk));
	jdff dff_B_gGqDyEHP8_2(.din(G70),.dout(w_dff_B_gGqDyEHP8_2),.clk(gclk));
	jdff dff_B_tFN5R1Mz9_2(.din(G67),.dout(w_dff_B_tFN5R1Mz9_2),.clk(gclk));
	jdff dff_B_dmDgtYiK5_2(.din(w_dff_B_tFN5R1Mz9_2),.dout(w_dff_B_dmDgtYiK5_2),.clk(gclk));
	jdff dff_A_P2xNaJpc5_1(.dout(w_n843_3[1]),.din(w_dff_A_P2xNaJpc5_1),.clk(gclk));
	jdff dff_A_np2aySLL9_1(.dout(w_dff_A_P2xNaJpc5_1),.din(w_dff_A_np2aySLL9_1),.clk(gclk));
	jdff dff_A_wHs9jq1k8_2(.dout(w_n843_3[2]),.din(w_dff_A_wHs9jq1k8_2),.clk(gclk));
	jdff dff_A_4OVrbwy44_2(.dout(w_dff_A_wHs9jq1k8_2),.din(w_dff_A_4OVrbwy44_2),.clk(gclk));
	jdff dff_A_oxwMc8g02_2(.dout(w_dff_A_4OVrbwy44_2),.din(w_dff_A_oxwMc8g02_2),.clk(gclk));
	jdff dff_A_ILrysShD0_2(.dout(w_dff_A_oxwMc8g02_2),.din(w_dff_A_ILrysShD0_2),.clk(gclk));
	jdff dff_A_2SUQv1QZ1_1(.dout(w_n840_3[1]),.din(w_dff_A_2SUQv1QZ1_1),.clk(gclk));
	jdff dff_A_1WNx31T11_2(.dout(w_n840_3[2]),.din(w_dff_A_1WNx31T11_2),.clk(gclk));
	jdff dff_A_GSoiYBCs5_2(.dout(w_dff_A_1WNx31T11_2),.din(w_dff_A_GSoiYBCs5_2),.clk(gclk));
	jdff dff_B_XTnXtpgM8_0(.din(n1081),.dout(w_dff_B_XTnXtpgM8_0),.clk(gclk));
	jdff dff_B_gtS9rtlA1_0(.din(n1080),.dout(w_dff_B_gtS9rtlA1_0),.clk(gclk));
	jdff dff_B_a4nihD729_0(.din(w_dff_B_gtS9rtlA1_0),.dout(w_dff_B_a4nihD729_0),.clk(gclk));
	jdff dff_B_Xh8RYayb9_0(.din(w_dff_B_a4nihD729_0),.dout(w_dff_B_Xh8RYayb9_0),.clk(gclk));
	jdff dff_B_mCRNHctH2_0(.din(w_dff_B_Xh8RYayb9_0),.dout(w_dff_B_mCRNHctH2_0),.clk(gclk));
	jdff dff_B_x8zkF9130_0(.din(w_dff_B_mCRNHctH2_0),.dout(w_dff_B_x8zkF9130_0),.clk(gclk));
	jdff dff_B_vn3QLHjX3_0(.din(w_dff_B_x8zkF9130_0),.dout(w_dff_B_vn3QLHjX3_0),.clk(gclk));
	jdff dff_B_KW5161zW1_0(.din(w_dff_B_vn3QLHjX3_0),.dout(w_dff_B_KW5161zW1_0),.clk(gclk));
	jdff dff_B_kcz1biqD4_0(.din(w_dff_B_KW5161zW1_0),.dout(w_dff_B_kcz1biqD4_0),.clk(gclk));
	jdff dff_B_GB4tiu9b0_0(.din(w_dff_B_kcz1biqD4_0),.dout(w_dff_B_GB4tiu9b0_0),.clk(gclk));
	jdff dff_B_ay1FvGnp2_0(.din(w_dff_B_GB4tiu9b0_0),.dout(w_dff_B_ay1FvGnp2_0),.clk(gclk));
	jdff dff_B_DhAD15Lh7_0(.din(w_dff_B_ay1FvGnp2_0),.dout(w_dff_B_DhAD15Lh7_0),.clk(gclk));
	jdff dff_B_W3ZZw4Cn9_0(.din(w_dff_B_DhAD15Lh7_0),.dout(w_dff_B_W3ZZw4Cn9_0),.clk(gclk));
	jdff dff_B_WjCWHaAT4_0(.din(n1079),.dout(w_dff_B_WjCWHaAT4_0),.clk(gclk));
	jdff dff_A_BxdxAuTy3_0(.dout(w_n988_4[0]),.din(w_dff_A_BxdxAuTy3_0),.clk(gclk));
	jdff dff_A_QRetefqs5_0(.dout(w_dff_A_BxdxAuTy3_0),.din(w_dff_A_QRetefqs5_0),.clk(gclk));
	jdff dff_A_0rMw0z2f3_0(.dout(w_dff_A_QRetefqs5_0),.din(w_dff_A_0rMw0z2f3_0),.clk(gclk));
	jdff dff_A_fMXsBj9m6_0(.dout(w_dff_A_0rMw0z2f3_0),.din(w_dff_A_fMXsBj9m6_0),.clk(gclk));
	jdff dff_A_MmLzWgdh3_0(.dout(w_dff_A_fMXsBj9m6_0),.din(w_dff_A_MmLzWgdh3_0),.clk(gclk));
	jdff dff_A_noo8JoPT4_0(.dout(w_dff_A_MmLzWgdh3_0),.din(w_dff_A_noo8JoPT4_0),.clk(gclk));
	jdff dff_A_LzgFPlqJ2_0(.dout(w_dff_A_noo8JoPT4_0),.din(w_dff_A_LzgFPlqJ2_0),.clk(gclk));
	jdff dff_A_gHzBM0LF5_0(.dout(w_n985_4[0]),.din(w_dff_A_gHzBM0LF5_0),.clk(gclk));
	jdff dff_A_EysPXUwI6_0(.dout(w_dff_A_gHzBM0LF5_0),.din(w_dff_A_EysPXUwI6_0),.clk(gclk));
	jdff dff_A_AyI6GO7f7_0(.dout(w_dff_A_EysPXUwI6_0),.din(w_dff_A_AyI6GO7f7_0),.clk(gclk));
	jdff dff_A_guqWhoe00_0(.dout(w_dff_A_AyI6GO7f7_0),.din(w_dff_A_guqWhoe00_0),.clk(gclk));
	jdff dff_A_YiYShXeA3_0(.dout(w_dff_A_guqWhoe00_0),.din(w_dff_A_YiYShXeA3_0),.clk(gclk));
	jdff dff_A_KRV72M3l8_0(.dout(w_dff_A_YiYShXeA3_0),.din(w_dff_A_KRV72M3l8_0),.clk(gclk));
	jdff dff_A_KyShtKWw0_0(.dout(w_dff_A_KRV72M3l8_0),.din(w_dff_A_KyShtKWw0_0),.clk(gclk));
	jdff dff_A_p7tmQuyS8_0(.dout(w_dff_A_KyShtKWw0_0),.din(w_dff_A_p7tmQuyS8_0),.clk(gclk));
	jdff dff_B_FHdlhyxr5_0(.din(n1089),.dout(w_dff_B_FHdlhyxr5_0),.clk(gclk));
	jdff dff_B_P6gQ9s1P0_0(.din(w_dff_B_FHdlhyxr5_0),.dout(w_dff_B_P6gQ9s1P0_0),.clk(gclk));
	jdff dff_B_T3z170Uf8_0(.din(w_dff_B_P6gQ9s1P0_0),.dout(w_dff_B_T3z170Uf8_0),.clk(gclk));
	jdff dff_B_gq0Tum2J9_0(.din(n1088),.dout(w_dff_B_gq0Tum2J9_0),.clk(gclk));
	jdff dff_B_oBnIaTDD1_0(.din(w_dff_B_gq0Tum2J9_0),.dout(w_dff_B_oBnIaTDD1_0),.clk(gclk));
	jdff dff_B_TWbyM5508_0(.din(w_dff_B_oBnIaTDD1_0),.dout(w_dff_B_TWbyM5508_0),.clk(gclk));
	jdff dff_B_nXtGAaXD7_0(.din(w_dff_B_TWbyM5508_0),.dout(w_dff_B_nXtGAaXD7_0),.clk(gclk));
	jdff dff_B_uSdc2ox50_0(.din(w_dff_B_nXtGAaXD7_0),.dout(w_dff_B_uSdc2ox50_0),.clk(gclk));
	jdff dff_B_W18ARSSY5_0(.din(w_dff_B_uSdc2ox50_0),.dout(w_dff_B_W18ARSSY5_0),.clk(gclk));
	jdff dff_B_UroukBto2_0(.din(n1087),.dout(w_dff_B_UroukBto2_0),.clk(gclk));
	jdff dff_B_EoeafYTF2_0(.din(n1097),.dout(w_dff_B_EoeafYTF2_0),.clk(gclk));
	jdff dff_B_KlIGP9566_0(.din(w_dff_B_EoeafYTF2_0),.dout(w_dff_B_KlIGP9566_0),.clk(gclk));
	jdff dff_B_K7rIN2yn3_0(.din(n1096),.dout(w_dff_B_K7rIN2yn3_0),.clk(gclk));
	jdff dff_B_62J7ihQl9_0(.din(w_dff_B_K7rIN2yn3_0),.dout(w_dff_B_62J7ihQl9_0),.clk(gclk));
	jdff dff_B_1v5WwXJz9_0(.din(w_dff_B_62J7ihQl9_0),.dout(w_dff_B_1v5WwXJz9_0),.clk(gclk));
	jdff dff_B_bxUHRyXk9_0(.din(w_dff_B_1v5WwXJz9_0),.dout(w_dff_B_bxUHRyXk9_0),.clk(gclk));
	jdff dff_B_kriV0NXd8_0(.din(w_dff_B_bxUHRyXk9_0),.dout(w_dff_B_kriV0NXd8_0),.clk(gclk));
	jdff dff_B_c7xR3tpJ3_0(.din(w_dff_B_kriV0NXd8_0),.dout(w_dff_B_c7xR3tpJ3_0),.clk(gclk));
	jdff dff_B_3E2BngQZ8_0(.din(w_dff_B_c7xR3tpJ3_0),.dout(w_dff_B_3E2BngQZ8_0),.clk(gclk));
	jdff dff_B_D7JximM67_0(.din(w_dff_B_3E2BngQZ8_0),.dout(w_dff_B_D7JximM67_0),.clk(gclk));
	jdff dff_B_0aRS2stc2_0(.din(n1095),.dout(w_dff_B_0aRS2stc2_0),.clk(gclk));
	jdff dff_A_1BC24AqY8_0(.dout(w_G137_8[0]),.din(w_dff_A_1BC24AqY8_0),.clk(gclk));
	jdff dff_A_gko4YKyK2_2(.dout(w_G137_8[2]),.din(w_dff_A_gko4YKyK2_2),.clk(gclk));
	jdff dff_A_px96T8OU9_2(.dout(w_dff_A_gko4YKyK2_2),.din(w_dff_A_px96T8OU9_2),.clk(gclk));
	jdff dff_A_E9gPA6Lu8_2(.dout(w_dff_A_px96T8OU9_2),.din(w_dff_A_E9gPA6Lu8_2),.clk(gclk));
	jdff dff_A_e6UNA8IQ6_2(.dout(w_dff_A_E9gPA6Lu8_2),.din(w_dff_A_e6UNA8IQ6_2),.clk(gclk));
	jdff dff_B_BprNyinQ4_0(.din(n1105),.dout(w_dff_B_BprNyinQ4_0),.clk(gclk));
	jdff dff_B_OS5ZA7bL9_0(.din(n1104),.dout(w_dff_B_OS5ZA7bL9_0),.clk(gclk));
	jdff dff_B_VEjMUxYL5_0(.din(w_dff_B_OS5ZA7bL9_0),.dout(w_dff_B_VEjMUxYL5_0),.clk(gclk));
	jdff dff_B_no1Xjybo0_0(.din(w_dff_B_VEjMUxYL5_0),.dout(w_dff_B_no1Xjybo0_0),.clk(gclk));
	jdff dff_B_EmVfzZRj6_0(.din(w_dff_B_no1Xjybo0_0),.dout(w_dff_B_EmVfzZRj6_0),.clk(gclk));
	jdff dff_B_1KUHvEMk1_0(.din(w_dff_B_EmVfzZRj6_0),.dout(w_dff_B_1KUHvEMk1_0),.clk(gclk));
	jdff dff_B_x8V8CaWD3_0(.din(w_dff_B_1KUHvEMk1_0),.dout(w_dff_B_x8V8CaWD3_0),.clk(gclk));
	jdff dff_B_u5SYxqAU4_0(.din(w_dff_B_x8V8CaWD3_0),.dout(w_dff_B_u5SYxqAU4_0),.clk(gclk));
	jdff dff_B_JaNqa41D0_0(.din(w_dff_B_u5SYxqAU4_0),.dout(w_dff_B_JaNqa41D0_0),.clk(gclk));
	jdff dff_B_soNc0u147_0(.din(w_dff_B_JaNqa41D0_0),.dout(w_dff_B_soNc0u147_0),.clk(gclk));
	jdff dff_B_5qbHPi520_0(.din(w_dff_B_soNc0u147_0),.dout(w_dff_B_5qbHPi520_0),.clk(gclk));
	jdff dff_B_xkoqWe9W8_0(.din(n1103),.dout(w_dff_B_xkoqWe9W8_0),.clk(gclk));
	jdff dff_A_DyrteZ6p1_0(.dout(w_n988_3[0]),.din(w_dff_A_DyrteZ6p1_0),.clk(gclk));
	jdff dff_A_HppuP6Js1_0(.dout(w_dff_A_DyrteZ6p1_0),.din(w_dff_A_HppuP6Js1_0),.clk(gclk));
	jdff dff_A_DDViaX6f7_0(.dout(w_dff_A_HppuP6Js1_0),.din(w_dff_A_DDViaX6f7_0),.clk(gclk));
	jdff dff_A_dpyfnwzd8_0(.dout(w_dff_A_DDViaX6f7_0),.din(w_dff_A_dpyfnwzd8_0),.clk(gclk));
	jdff dff_A_atiftQfm6_1(.dout(w_n988_3[1]),.din(w_dff_A_atiftQfm6_1),.clk(gclk));
	jdff dff_A_SSmOGXFU7_1(.dout(w_dff_A_atiftQfm6_1),.din(w_dff_A_SSmOGXFU7_1),.clk(gclk));
	jdff dff_A_qNjLDCVg7_0(.dout(w_n985_3[0]),.din(w_dff_A_qNjLDCVg7_0),.clk(gclk));
	jdff dff_A_fCAycZkA0_0(.dout(w_dff_A_qNjLDCVg7_0),.din(w_dff_A_fCAycZkA0_0),.clk(gclk));
	jdff dff_A_cN4ywjen3_1(.dout(w_n985_3[1]),.din(w_dff_A_cN4ywjen3_1),.clk(gclk));
	jdff dff_B_OgIeoO6B4_0(.din(n1113),.dout(w_dff_B_OgIeoO6B4_0),.clk(gclk));
	jdff dff_B_En1prRs44_0(.din(n1112),.dout(w_dff_B_En1prRs44_0),.clk(gclk));
	jdff dff_B_fwlSjpo56_0(.din(w_dff_B_En1prRs44_0),.dout(w_dff_B_fwlSjpo56_0),.clk(gclk));
	jdff dff_B_upMTLFBi1_0(.din(w_dff_B_fwlSjpo56_0),.dout(w_dff_B_upMTLFBi1_0),.clk(gclk));
	jdff dff_B_QNvj0gwz1_0(.din(w_dff_B_upMTLFBi1_0),.dout(w_dff_B_QNvj0gwz1_0),.clk(gclk));
	jdff dff_B_ZhMkt2bJ3_0(.din(w_dff_B_QNvj0gwz1_0),.dout(w_dff_B_ZhMkt2bJ3_0),.clk(gclk));
	jdff dff_B_9dOWhQTQ3_0(.din(w_dff_B_ZhMkt2bJ3_0),.dout(w_dff_B_9dOWhQTQ3_0),.clk(gclk));
	jdff dff_B_zThJXWQv4_0(.din(w_dff_B_9dOWhQTQ3_0),.dout(w_dff_B_zThJXWQv4_0),.clk(gclk));
	jdff dff_B_vl0nWUn87_0(.din(w_dff_B_zThJXWQv4_0),.dout(w_dff_B_vl0nWUn87_0),.clk(gclk));
	jdff dff_B_8NuyTHxS8_0(.din(w_dff_B_vl0nWUn87_0),.dout(w_dff_B_8NuyTHxS8_0),.clk(gclk));
	jdff dff_B_KanJafkY3_0(.din(w_dff_B_8NuyTHxS8_0),.dout(w_dff_B_KanJafkY3_0),.clk(gclk));
	jdff dff_B_70WijCaP4_0(.din(w_dff_B_KanJafkY3_0),.dout(w_dff_B_70WijCaP4_0),.clk(gclk));
	jdff dff_B_GzcXBlx84_0(.din(w_dff_B_70WijCaP4_0),.dout(w_dff_B_GzcXBlx84_0),.clk(gclk));
	jdff dff_B_5KDeyqNZ2_0(.din(n1111),.dout(w_dff_B_5KDeyqNZ2_0),.clk(gclk));
	jdff dff_B_JcnLwAmB3_2(.din(G170),.dout(w_dff_B_JcnLwAmB3_2),.clk(gclk));
	jdff dff_B_XcbrhrKy6_2(.din(G200),.dout(w_dff_B_XcbrhrKy6_2),.clk(gclk));
	jdff dff_B_YbWxK6xW4_2(.din(w_dff_B_XcbrhrKy6_2),.dout(w_dff_B_YbWxK6xW4_2),.clk(gclk));
	jdff dff_A_9eKJdbRh4_0(.dout(w_n1002_4[0]),.din(w_dff_A_9eKJdbRh4_0),.clk(gclk));
	jdff dff_A_sLqpRWvs9_0(.dout(w_dff_A_9eKJdbRh4_0),.din(w_dff_A_sLqpRWvs9_0),.clk(gclk));
	jdff dff_A_GgBhcmtO9_0(.dout(w_dff_A_sLqpRWvs9_0),.din(w_dff_A_GgBhcmtO9_0),.clk(gclk));
	jdff dff_A_47zHNPzp2_0(.dout(w_dff_A_GgBhcmtO9_0),.din(w_dff_A_47zHNPzp2_0),.clk(gclk));
	jdff dff_A_deeyw11t2_0(.dout(w_dff_A_47zHNPzp2_0),.din(w_dff_A_deeyw11t2_0),.clk(gclk));
	jdff dff_A_6Vi4GMIZ8_0(.dout(w_dff_A_deeyw11t2_0),.din(w_dff_A_6Vi4GMIZ8_0),.clk(gclk));
	jdff dff_A_kMyjH4IQ1_0(.dout(w_dff_A_6Vi4GMIZ8_0),.din(w_dff_A_kMyjH4IQ1_0),.clk(gclk));
	jdff dff_B_ZpKwYiag7_0(.din(n814),.dout(w_dff_B_ZpKwYiag7_0),.clk(gclk));
	jdff dff_B_AP3B4fjv9_0(.din(w_dff_B_ZpKwYiag7_0),.dout(w_dff_B_AP3B4fjv9_0),.clk(gclk));
	jdff dff_B_BOcGSZIL7_0(.din(w_dff_B_AP3B4fjv9_0),.dout(w_dff_B_BOcGSZIL7_0),.clk(gclk));
	jdff dff_B_RgcqJiYQ9_0(.din(w_dff_B_BOcGSZIL7_0),.dout(w_dff_B_RgcqJiYQ9_0),.clk(gclk));
	jdff dff_B_COUyQcJW3_0(.din(w_dff_B_RgcqJiYQ9_0),.dout(w_dff_B_COUyQcJW3_0),.clk(gclk));
	jdff dff_B_6PCInH3y0_0(.din(w_dff_B_COUyQcJW3_0),.dout(w_dff_B_6PCInH3y0_0),.clk(gclk));
	jdff dff_B_eKL3llTz4_0(.din(n813),.dout(w_dff_B_eKL3llTz4_0),.clk(gclk));
	jdff dff_B_FDZowcrK5_0(.din(w_dff_B_eKL3llTz4_0),.dout(w_dff_B_FDZowcrK5_0),.clk(gclk));
	jdff dff_B_MC7EYT0u1_1(.din(G52),.dout(w_dff_B_MC7EYT0u1_1),.clk(gclk));
	jdff dff_B_TXDqdpuD8_1(.din(w_dff_B_MC7EYT0u1_1),.dout(w_dff_B_TXDqdpuD8_1),.clk(gclk));
	jdff dff_B_6x1nUjZV6_0(.din(n433),.dout(w_dff_B_6x1nUjZV6_0),.clk(gclk));
	jdff dff_B_9iNE9XXP0_1(.din(n425),.dout(w_dff_B_9iNE9XXP0_1),.clk(gclk));
	jdff dff_A_RR97Thn17_0(.dout(w_n999_4[0]),.din(w_dff_A_RR97Thn17_0),.clk(gclk));
	jdff dff_A_7nm7N9su5_0(.dout(w_dff_A_RR97Thn17_0),.din(w_dff_A_7nm7N9su5_0),.clk(gclk));
	jdff dff_A_3MCc1XmU7_0(.dout(w_dff_A_7nm7N9su5_0),.din(w_dff_A_3MCc1XmU7_0),.clk(gclk));
	jdff dff_A_waTVUbUa8_0(.dout(w_dff_A_3MCc1XmU7_0),.din(w_dff_A_waTVUbUa8_0),.clk(gclk));
	jdff dff_A_Rr2iFJ0p9_0(.dout(w_dff_A_waTVUbUa8_0),.din(w_dff_A_Rr2iFJ0p9_0),.clk(gclk));
	jdff dff_A_exPsBILN4_0(.dout(w_dff_A_Rr2iFJ0p9_0),.din(w_dff_A_exPsBILN4_0),.clk(gclk));
	jdff dff_A_mLONIbjn9_0(.dout(w_dff_A_exPsBILN4_0),.din(w_dff_A_mLONIbjn9_0),.clk(gclk));
	jdff dff_A_a9Qm4DtW7_0(.dout(w_dff_A_mLONIbjn9_0),.din(w_dff_A_a9Qm4DtW7_0),.clk(gclk));
	jdff dff_B_fq9rhGuf4_0(.din(n867),.dout(w_dff_B_fq9rhGuf4_0),.clk(gclk));
	jdff dff_B_PuyzAVSH1_0(.din(w_dff_B_fq9rhGuf4_0),.dout(w_dff_B_PuyzAVSH1_0),.clk(gclk));
	jdff dff_B_8mQ0XSkc9_0(.din(w_dff_B_PuyzAVSH1_0),.dout(w_dff_B_8mQ0XSkc9_0),.clk(gclk));
	jdff dff_B_R7YEhzvu4_0(.din(w_dff_B_8mQ0XSkc9_0),.dout(w_dff_B_R7YEhzvu4_0),.clk(gclk));
	jdff dff_B_PR0izhPs7_0(.din(w_dff_B_R7YEhzvu4_0),.dout(w_dff_B_PR0izhPs7_0),.clk(gclk));
	jdff dff_B_ULeG9tiY5_0(.din(w_dff_B_PR0izhPs7_0),.dout(w_dff_B_ULeG9tiY5_0),.clk(gclk));
	jdff dff_B_Vk0JY3u23_0(.din(w_dff_B_ULeG9tiY5_0),.dout(w_dff_B_Vk0JY3u23_0),.clk(gclk));
	jdff dff_B_94rHWRBM0_0(.din(w_dff_B_Vk0JY3u23_0),.dout(w_dff_B_94rHWRBM0_0),.clk(gclk));
	jdff dff_B_1cLKOKWl7_0(.din(n866),.dout(w_dff_B_1cLKOKWl7_0),.clk(gclk));
	jdff dff_B_WUOp7OYO9_0(.din(w_dff_B_1cLKOKWl7_0),.dout(w_dff_B_WUOp7OYO9_0),.clk(gclk));
	jdff dff_B_M89nhxxV1_1(.din(G122),.dout(w_dff_B_M89nhxxV1_1),.clk(gclk));
	jdff dff_B_Pvx58Jyu8_1(.din(w_dff_B_M89nhxxV1_1),.dout(w_dff_B_Pvx58Jyu8_1),.clk(gclk));
	jdff dff_B_FGBLF5RG1_0(.din(n469),.dout(w_dff_B_FGBLF5RG1_0),.clk(gclk));
	jdff dff_B_4NDoHUfP4_1(.din(n461),.dout(w_dff_B_4NDoHUfP4_1),.clk(gclk));
	jdff dff_B_iNlZN9jk3_1(.din(n852),.dout(w_dff_B_iNlZN9jk3_1),.clk(gclk));
	jdff dff_B_5zist2W43_1(.din(w_dff_B_iNlZN9jk3_1),.dout(w_dff_B_5zist2W43_1),.clk(gclk));
	jdff dff_B_EmjnAZEq6_1(.din(w_dff_B_5zist2W43_1),.dout(w_dff_B_EmjnAZEq6_1),.clk(gclk));
	jdff dff_B_pHWzAP7Y9_1(.din(w_dff_B_EmjnAZEq6_1),.dout(w_dff_B_pHWzAP7Y9_1),.clk(gclk));
	jdff dff_B_AuHxWxW40_1(.din(w_dff_B_pHWzAP7Y9_1),.dout(w_dff_B_AuHxWxW40_1),.clk(gclk));
	jdff dff_B_73bDIewy7_1(.din(w_dff_B_AuHxWxW40_1),.dout(w_dff_B_73bDIewy7_1),.clk(gclk));
	jdff dff_B_IomaU9x00_0(.din(n1121),.dout(w_dff_B_IomaU9x00_0),.clk(gclk));
	jdff dff_B_b8GBKIl80_0(.din(w_dff_B_IomaU9x00_0),.dout(w_dff_B_b8GBKIl80_0),.clk(gclk));
	jdff dff_B_CNjIMwUF5_0(.din(w_dff_B_b8GBKIl80_0),.dout(w_dff_B_CNjIMwUF5_0),.clk(gclk));
	jdff dff_B_iljtuNsl0_0(.din(n1120),.dout(w_dff_B_iljtuNsl0_0),.clk(gclk));
	jdff dff_B_OKBLelgK2_0(.din(w_dff_B_iljtuNsl0_0),.dout(w_dff_B_OKBLelgK2_0),.clk(gclk));
	jdff dff_B_aOxlDQ062_0(.din(w_dff_B_OKBLelgK2_0),.dout(w_dff_B_aOxlDQ062_0),.clk(gclk));
	jdff dff_B_yOorlP4o7_0(.din(w_dff_B_aOxlDQ062_0),.dout(w_dff_B_yOorlP4o7_0),.clk(gclk));
	jdff dff_B_PZcdhNna8_0(.din(w_dff_B_yOorlP4o7_0),.dout(w_dff_B_PZcdhNna8_0),.clk(gclk));
	jdff dff_B_wahLog2R8_0(.din(w_dff_B_PZcdhNna8_0),.dout(w_dff_B_wahLog2R8_0),.clk(gclk));
	jdff dff_B_Dria40VK9_0(.din(n1119),.dout(w_dff_B_Dria40VK9_0),.clk(gclk));
	jdff dff_B_rhmpJRnq2_2(.din(G158),.dout(w_dff_B_rhmpJRnq2_2),.clk(gclk));
	jdff dff_B_Kcwo7PKd4_2(.din(G188),.dout(w_dff_B_Kcwo7PKd4_2),.clk(gclk));
	jdff dff_B_oPu1wzDG3_2(.din(w_dff_B_Kcwo7PKd4_2),.dout(w_dff_B_oPu1wzDG3_2),.clk(gclk));
	jdff dff_B_wTdfFCYR9_0(.din(n768),.dout(w_dff_B_wTdfFCYR9_0),.clk(gclk));
	jdff dff_B_Dplxahew3_0(.din(w_dff_B_wTdfFCYR9_0),.dout(w_dff_B_Dplxahew3_0),.clk(gclk));
	jdff dff_B_0cZsRaBs4_1(.din(G129),.dout(w_dff_B_0cZsRaBs4_1),.clk(gclk));
	jdff dff_B_UlMVrDl49_1(.din(w_dff_B_0cZsRaBs4_1),.dout(w_dff_B_UlMVrDl49_1),.clk(gclk));
	jdff dff_A_y5ATf2KU7_1(.dout(w_n397_0[1]),.din(w_dff_A_y5ATf2KU7_1),.clk(gclk));
	jdff dff_B_hpRNacob3_0(.din(n396),.dout(w_dff_B_hpRNacob3_0),.clk(gclk));
	jdff dff_B_ME1rjpGW3_1(.din(n387),.dout(w_dff_B_ME1rjpGW3_1),.clk(gclk));
	jdff dff_A_zE2BDkb14_0(.dout(w_n748_4[0]),.din(w_dff_A_zE2BDkb14_0),.clk(gclk));
	jdff dff_B_1cDh0C0P1_0(.din(n898),.dout(w_dff_B_1cDh0C0P1_0),.clk(gclk));
	jdff dff_B_e6H0owVM2_0(.din(w_dff_B_1cDh0C0P1_0),.dout(w_dff_B_e6H0owVM2_0),.clk(gclk));
	jdff dff_B_XV6f11p15_0(.din(w_dff_B_e6H0owVM2_0),.dout(w_dff_B_XV6f11p15_0),.clk(gclk));
	jdff dff_B_i7cpOCT88_0(.din(w_dff_B_XV6f11p15_0),.dout(w_dff_B_i7cpOCT88_0),.clk(gclk));
	jdff dff_B_2NrrkCob0_0(.din(n897),.dout(w_dff_B_2NrrkCob0_0),.clk(gclk));
	jdff dff_B_WEhjN6ji8_0(.din(w_dff_B_2NrrkCob0_0),.dout(w_dff_B_WEhjN6ji8_0),.clk(gclk));
	jdff dff_B_HkCz8Ird5_1(.din(G126),.dout(w_dff_B_HkCz8Ird5_1),.clk(gclk));
	jdff dff_B_mEvSGX876_1(.din(w_dff_B_HkCz8Ird5_1),.dout(w_dff_B_mEvSGX876_1),.clk(gclk));
	jdff dff_B_NznqOe2n0_0(.din(n493),.dout(w_dff_B_NznqOe2n0_0),.clk(gclk));
	jdff dff_B_9BFouGyv7_1(.din(n485),.dout(w_dff_B_9BFouGyv7_1),.clk(gclk));
	jdff dff_B_90uOtjj17_0(.din(n889),.dout(w_dff_B_90uOtjj17_0),.clk(gclk));
	jdff dff_A_Ovfi9hOb9_1(.dout(w_G137_7[1]),.din(w_dff_A_Ovfi9hOb9_1),.clk(gclk));
	jdff dff_A_g0BHYwOQ1_1(.dout(w_dff_A_Ovfi9hOb9_1),.din(w_dff_A_g0BHYwOQ1_1),.clk(gclk));
	jdff dff_A_973G9RMs0_1(.dout(w_dff_A_g0BHYwOQ1_1),.din(w_dff_A_973G9RMs0_1),.clk(gclk));
	jdff dff_A_Dg47uAWB2_1(.dout(w_dff_A_973G9RMs0_1),.din(w_dff_A_Dg47uAWB2_1),.clk(gclk));
	jdff dff_A_MA2pURe37_2(.dout(w_G137_7[2]),.din(w_dff_A_MA2pURe37_2),.clk(gclk));
	jdff dff_A_srnJSoTh0_2(.dout(w_dff_A_MA2pURe37_2),.din(w_dff_A_srnJSoTh0_2),.clk(gclk));
	jdff dff_A_Rt3k4Nc34_0(.dout(w_G137_2[0]),.din(w_dff_A_Rt3k4Nc34_0),.clk(gclk));
	jdff dff_A_UZDXURbz1_0(.dout(w_dff_A_Rt3k4Nc34_0),.din(w_dff_A_UZDXURbz1_0),.clk(gclk));
	jdff dff_A_kZc9yHur4_0(.dout(w_dff_A_UZDXURbz1_0),.din(w_dff_A_kZc9yHur4_0),.clk(gclk));
	jdff dff_A_rYHWvkE08_0(.dout(w_dff_A_kZc9yHur4_0),.din(w_dff_A_rYHWvkE08_0),.clk(gclk));
	jdff dff_A_fGYOpEif8_1(.dout(w_G137_2[1]),.din(w_dff_A_fGYOpEif8_1),.clk(gclk));
	jdff dff_A_AHSc45R73_1(.dout(w_dff_A_fGYOpEif8_1),.din(w_dff_A_AHSc45R73_1),.clk(gclk));
	jdff dff_A_hKm7mnYD0_1(.dout(w_dff_A_AHSc45R73_1),.din(w_dff_A_hKm7mnYD0_1),.clk(gclk));
	jdff dff_A_E3CF4CRp0_1(.dout(w_dff_A_hKm7mnYD0_1),.din(w_dff_A_E3CF4CRp0_1),.clk(gclk));
	jdff dff_B_joGhvehh8_0(.din(n1129),.dout(w_dff_B_joGhvehh8_0),.clk(gclk));
	jdff dff_B_reDfHA2s8_0(.din(w_dff_B_joGhvehh8_0),.dout(w_dff_B_reDfHA2s8_0),.clk(gclk));
	jdff dff_B_3ZpPZ9th1_0(.din(n1128),.dout(w_dff_B_3ZpPZ9th1_0),.clk(gclk));
	jdff dff_B_zi3z1JL30_0(.din(w_dff_B_3ZpPZ9th1_0),.dout(w_dff_B_zi3z1JL30_0),.clk(gclk));
	jdff dff_B_MY3JNuaJ7_0(.din(w_dff_B_zi3z1JL30_0),.dout(w_dff_B_MY3JNuaJ7_0),.clk(gclk));
	jdff dff_B_PFdWbYIz0_0(.din(w_dff_B_MY3JNuaJ7_0),.dout(w_dff_B_PFdWbYIz0_0),.clk(gclk));
	jdff dff_B_CgAU9tAa9_0(.din(w_dff_B_PFdWbYIz0_0),.dout(w_dff_B_CgAU9tAa9_0),.clk(gclk));
	jdff dff_B_SIQJrTRL8_0(.din(w_dff_B_CgAU9tAa9_0),.dout(w_dff_B_SIQJrTRL8_0),.clk(gclk));
	jdff dff_B_t6ibS3ha3_0(.din(w_dff_B_SIQJrTRL8_0),.dout(w_dff_B_t6ibS3ha3_0),.clk(gclk));
	jdff dff_B_q1U8qdc83_0(.din(w_dff_B_t6ibS3ha3_0),.dout(w_dff_B_q1U8qdc83_0),.clk(gclk));
	jdff dff_B_htxaFz5i3_0(.din(n1127),.dout(w_dff_B_htxaFz5i3_0),.clk(gclk));
	jdff dff_B_Jwib4FT85_2(.din(G152),.dout(w_dff_B_Jwib4FT85_2),.clk(gclk));
	jdff dff_B_nx8Dlb4J8_2(.din(G155),.dout(w_dff_B_nx8Dlb4J8_2),.clk(gclk));
	jdff dff_B_tyClrbYL5_2(.din(w_dff_B_nx8Dlb4J8_2),.dout(w_dff_B_tyClrbYL5_2),.clk(gclk));
	jdff dff_B_qGUnuodJ7_0(.din(n837),.dout(w_dff_B_qGUnuodJ7_0),.clk(gclk));
	jdff dff_B_folb1ScY3_0(.din(w_dff_B_qGUnuodJ7_0),.dout(w_dff_B_folb1ScY3_0),.clk(gclk));
	jdff dff_B_ItJBMpig6_0(.din(n836),.dout(w_dff_B_ItJBMpig6_0),.clk(gclk));
	jdff dff_B_qQWnhljy2_0(.din(w_dff_B_ItJBMpig6_0),.dout(w_dff_B_qQWnhljy2_0),.clk(gclk));
	jdff dff_B_PgOv85E25_1(.din(G119),.dout(w_dff_B_PgOv85E25_1),.clk(gclk));
	jdff dff_B_oO4A8jg59_1(.din(w_dff_B_PgOv85E25_1),.dout(w_dff_B_oO4A8jg59_1),.clk(gclk));
	jdff dff_B_90sOMuAW5_0(.din(n444),.dout(w_dff_B_90sOMuAW5_0),.clk(gclk));
	jdff dff_B_AHuoukWT8_1(.din(n436),.dout(w_dff_B_AHuoukWT8_1),.clk(gclk));
	jdff dff_A_wy6D8lKC3_0(.dout(w_n744_1[0]),.din(w_dff_A_wy6D8lKC3_0),.clk(gclk));
	jdff dff_A_SKuI1rEA3_0(.dout(w_dff_A_wy6D8lKC3_0),.din(w_dff_A_SKuI1rEA3_0),.clk(gclk));
	jdff dff_A_aaSUKXGg5_0(.dout(w_dff_A_SKuI1rEA3_0),.din(w_dff_A_aaSUKXGg5_0),.clk(gclk));
	jdff dff_A_sW34QoFa6_0(.dout(w_dff_A_aaSUKXGg5_0),.din(w_dff_A_sW34QoFa6_0),.clk(gclk));
	jdff dff_A_J2Ts6Yvv4_0(.dout(w_dff_A_sW34QoFa6_0),.din(w_dff_A_J2Ts6Yvv4_0),.clk(gclk));
	jdff dff_A_9oh8lctW9_0(.dout(w_dff_A_J2Ts6Yvv4_0),.din(w_dff_A_9oh8lctW9_0),.clk(gclk));
	jdff dff_B_Y7QT4HVk9_0(.din(n887),.dout(w_dff_B_Y7QT4HVk9_0),.clk(gclk));
	jdff dff_B_V597U4Y40_0(.din(w_dff_B_Y7QT4HVk9_0),.dout(w_dff_B_V597U4Y40_0),.clk(gclk));
	jdff dff_B_FUXuW4ch9_0(.din(w_dff_B_V597U4Y40_0),.dout(w_dff_B_FUXuW4ch9_0),.clk(gclk));
	jdff dff_B_xfw8lBFP9_0(.din(w_dff_B_FUXuW4ch9_0),.dout(w_dff_B_xfw8lBFP9_0),.clk(gclk));
	jdff dff_B_UWRP0Y5A5_0(.din(w_dff_B_xfw8lBFP9_0),.dout(w_dff_B_UWRP0Y5A5_0),.clk(gclk));
	jdff dff_B_u9EAxGG46_0(.din(n886),.dout(w_dff_B_u9EAxGG46_0),.clk(gclk));
	jdff dff_B_Y8q27l6j4_0(.din(w_dff_B_u9EAxGG46_0),.dout(w_dff_B_Y8q27l6j4_0),.clk(gclk));
	jdff dff_B_cytzVKcL3_1(.din(G127),.dout(w_dff_B_cytzVKcL3_1),.clk(gclk));
	jdff dff_B_A0F7fsOW6_1(.din(w_dff_B_cytzVKcL3_1),.dout(w_dff_B_A0F7fsOW6_1),.clk(gclk));
	jdff dff_A_8VKltBBU2_1(.dout(w_n459_0[1]),.din(w_dff_A_8VKltBBU2_1),.clk(gclk));
	jdff dff_B_YwJWY0nX7_0(.din(n458),.dout(w_dff_B_YwJWY0nX7_0),.clk(gclk));
	jdff dff_B_v0xWcDdw6_1(.din(n450),.dout(w_dff_B_v0xWcDdw6_1),.clk(gclk));
	jdff dff_B_ZNFHKvU31_0(.din(n1137),.dout(w_dff_B_ZNFHKvU31_0),.clk(gclk));
	jdff dff_B_6hklEctc2_0(.din(n1136),.dout(w_dff_B_6hklEctc2_0),.clk(gclk));
	jdff dff_B_DuHVaRYy5_0(.din(w_dff_B_6hklEctc2_0),.dout(w_dff_B_DuHVaRYy5_0),.clk(gclk));
	jdff dff_B_WS8OTYFr8_0(.din(w_dff_B_DuHVaRYy5_0),.dout(w_dff_B_WS8OTYFr8_0),.clk(gclk));
	jdff dff_B_hLJV7IoA7_0(.din(w_dff_B_WS8OTYFr8_0),.dout(w_dff_B_hLJV7IoA7_0),.clk(gclk));
	jdff dff_B_lgFfUvub0_0(.din(w_dff_B_hLJV7IoA7_0),.dout(w_dff_B_lgFfUvub0_0),.clk(gclk));
	jdff dff_B_PhJv75Xw4_0(.din(w_dff_B_lgFfUvub0_0),.dout(w_dff_B_PhJv75Xw4_0),.clk(gclk));
	jdff dff_B_wPp1weZE4_0(.din(w_dff_B_PhJv75Xw4_0),.dout(w_dff_B_wPp1weZE4_0),.clk(gclk));
	jdff dff_B_hUShEWNF6_0(.din(w_dff_B_wPp1weZE4_0),.dout(w_dff_B_hUShEWNF6_0),.clk(gclk));
	jdff dff_B_y8teBY6p8_0(.din(w_dff_B_hUShEWNF6_0),.dout(w_dff_B_y8teBY6p8_0),.clk(gclk));
	jdff dff_B_tntgAJsr9_0(.din(w_dff_B_y8teBY6p8_0),.dout(w_dff_B_tntgAJsr9_0),.clk(gclk));
	jdff dff_B_1vcrToXD2_0(.din(n1135),.dout(w_dff_B_1vcrToXD2_0),.clk(gclk));
	jdff dff_B_Yql3Al7D3_2(.din(G146),.dout(w_dff_B_Yql3Al7D3_2),.clk(gclk));
	jdff dff_B_eeyDiJgY2_2(.din(G149),.dout(w_dff_B_eeyDiJgY2_2),.clk(gclk));
	jdff dff_B_uqpvHaIJ6_2(.din(w_dff_B_eeyDiJgY2_2),.dout(w_dff_B_uqpvHaIJ6_2),.clk(gclk));
	jdff dff_A_B0n1OQAi3_0(.dout(w_n1002_3[0]),.din(w_dff_A_B0n1OQAi3_0),.clk(gclk));
	jdff dff_A_63pvQg8h8_0(.dout(w_dff_A_B0n1OQAi3_0),.din(w_dff_A_63pvQg8h8_0),.clk(gclk));
	jdff dff_A_BN4vH3IG5_0(.dout(w_dff_A_63pvQg8h8_0),.din(w_dff_A_BN4vH3IG5_0),.clk(gclk));
	jdff dff_A_6mb7RBXC1_0(.dout(w_dff_A_BN4vH3IG5_0),.din(w_dff_A_6mb7RBXC1_0),.clk(gclk));
	jdff dff_A_64erkCvW5_1(.dout(w_n1002_3[1]),.din(w_dff_A_64erkCvW5_1),.clk(gclk));
	jdff dff_A_BCAe3P7R0_1(.dout(w_dff_A_64erkCvW5_1),.din(w_dff_A_BCAe3P7R0_1),.clk(gclk));
	jdff dff_B_S2Or8NpQ2_0(.din(n826),.dout(w_dff_B_S2Or8NpQ2_0),.clk(gclk));
	jdff dff_B_AGGj8wiS0_0(.din(w_dff_B_S2Or8NpQ2_0),.dout(w_dff_B_AGGj8wiS0_0),.clk(gclk));
	jdff dff_B_BAfeW1eF9_0(.din(w_dff_B_AGGj8wiS0_0),.dout(w_dff_B_BAfeW1eF9_0),.clk(gclk));
	jdff dff_B_35uPWueG1_0(.din(w_dff_B_BAfeW1eF9_0),.dout(w_dff_B_35uPWueG1_0),.clk(gclk));
	jdff dff_B_yl3JbdgC0_0(.din(w_dff_B_35uPWueG1_0),.dout(w_dff_B_yl3JbdgC0_0),.clk(gclk));
	jdff dff_B_J1JxYypK8_0(.din(n824),.dout(w_dff_B_J1JxYypK8_0),.clk(gclk));
	jdff dff_B_AEPhoVEA0_1(.din(G130),.dout(w_dff_B_AEPhoVEA0_1),.clk(gclk));
	jdff dff_B_eRjeDWEg4_1(.din(w_dff_B_AEPhoVEA0_1),.dout(w_dff_B_eRjeDWEg4_1),.clk(gclk));
	jdff dff_B_Zz6Hvt2A8_0(.din(n413),.dout(w_dff_B_Zz6Hvt2A8_0),.clk(gclk));
	jdff dff_B_33ZGEYC72_1(.din(n816),.dout(w_dff_B_33ZGEYC72_1),.clk(gclk));
	jdff dff_B_6NNxzr0W7_1(.din(w_dff_B_33ZGEYC72_1),.dout(w_dff_B_6NNxzr0W7_1),.clk(gclk));
	jdff dff_B_8cbz5lvv5_1(.din(w_dff_B_6NNxzr0W7_1),.dout(w_dff_B_8cbz5lvv5_1),.clk(gclk));
	jdff dff_B_bjNjYMa54_1(.din(w_dff_B_8cbz5lvv5_1),.dout(w_dff_B_bjNjYMa54_1),.clk(gclk));
	jdff dff_B_ltmbQhDK8_1(.din(w_dff_B_bjNjYMa54_1),.dout(w_dff_B_ltmbQhDK8_1),.clk(gclk));
	jdff dff_A_hd1Eoys54_2(.dout(w_n744_0[2]),.din(w_dff_A_hd1Eoys54_2),.clk(gclk));
	jdff dff_A_GZRNoypF2_2(.dout(w_dff_A_hd1Eoys54_2),.din(w_dff_A_GZRNoypF2_2),.clk(gclk));
	jdff dff_A_4CavtIdX3_2(.dout(w_dff_A_GZRNoypF2_2),.din(w_dff_A_4CavtIdX3_2),.clk(gclk));
	jdff dff_A_wV0klqvI2_2(.dout(w_dff_A_4CavtIdX3_2),.din(w_dff_A_wV0klqvI2_2),.clk(gclk));
	jdff dff_B_Kk0V9Pnr3_3(.din(n744),.dout(w_dff_B_Kk0V9Pnr3_3),.clk(gclk));
	jdff dff_B_4K1igsW85_3(.din(w_dff_B_Kk0V9Pnr3_3),.dout(w_dff_B_4K1igsW85_3),.clk(gclk));
	jdff dff_A_sS2V6STz4_1(.dout(w_n748_3[1]),.din(w_dff_A_sS2V6STz4_1),.clk(gclk));
	jdff dff_A_sHOXtqEZ9_1(.dout(w_dff_A_sS2V6STz4_1),.din(w_dff_A_sHOXtqEZ9_1),.clk(gclk));
	jdff dff_A_PUPh2Q1J9_2(.dout(w_n748_3[2]),.din(w_dff_A_PUPh2Q1J9_2),.clk(gclk));
	jdff dff_A_bpcWVSnb9_2(.dout(w_dff_A_PUPh2Q1J9_2),.din(w_dff_A_bpcWVSnb9_2),.clk(gclk));
	jdff dff_A_w1Xm0ZBY8_2(.dout(w_dff_A_bpcWVSnb9_2),.din(w_dff_A_w1Xm0ZBY8_2),.clk(gclk));
	jdff dff_A_p1fNNdqi8_2(.dout(w_dff_A_w1Xm0ZBY8_2),.din(w_dff_A_p1fNNdqi8_2),.clk(gclk));
	jdff dff_A_5Ni3oU0t8_0(.dout(w_n999_3[0]),.din(w_dff_A_5Ni3oU0t8_0),.clk(gclk));
	jdff dff_A_i86dQOnh2_0(.dout(w_dff_A_5Ni3oU0t8_0),.din(w_dff_A_i86dQOnh2_0),.clk(gclk));
	jdff dff_A_QwZ9RiFX5_1(.dout(w_n999_3[1]),.din(w_dff_A_QwZ9RiFX5_1),.clk(gclk));
	jdff dff_B_0iCX4q2L4_0(.din(n874),.dout(w_dff_B_0iCX4q2L4_0),.clk(gclk));
	jdff dff_B_1IUmLE8N8_0(.din(w_dff_B_0iCX4q2L4_0),.dout(w_dff_B_1IUmLE8N8_0),.clk(gclk));
	jdff dff_B_5MhM0mvX9_0(.din(w_dff_B_1IUmLE8N8_0),.dout(w_dff_B_5MhM0mvX9_0),.clk(gclk));
	jdff dff_B_PIIXsSd08_0(.din(w_dff_B_5MhM0mvX9_0),.dout(w_dff_B_PIIXsSd08_0),.clk(gclk));
	jdff dff_B_yRUs2IVr8_0(.din(w_dff_B_PIIXsSd08_0),.dout(w_dff_B_yRUs2IVr8_0),.clk(gclk));
	jdff dff_B_fZP1RiSL2_0(.din(w_dff_B_yRUs2IVr8_0),.dout(w_dff_B_fZP1RiSL2_0),.clk(gclk));
	jdff dff_B_EcPTGb4R5_0(.din(n873),.dout(w_dff_B_EcPTGb4R5_0),.clk(gclk));
	jdff dff_B_wCO12kb00_0(.din(w_dff_B_EcPTGb4R5_0),.dout(w_dff_B_wCO12kb00_0),.clk(gclk));
	jdff dff_B_CXvXgtDY2_1(.din(G128),.dout(w_dff_B_CXvXgtDY2_1),.clk(gclk));
	jdff dff_B_QJsdoiVI0_1(.din(w_dff_B_CXvXgtDY2_1),.dout(w_dff_B_QJsdoiVI0_1),.clk(gclk));
	jdff dff_B_twvL3bjd5_0(.din(n480),.dout(w_dff_B_twvL3bjd5_0),.clk(gclk));
	jdff dff_B_XnnT7VXe0_1(.din(n472),.dout(w_dff_B_XnnT7VXe0_1),.clk(gclk));
	jdff dff_B_orm6dmTT0_0(.din(n858),.dout(w_dff_B_orm6dmTT0_0),.clk(gclk));
	jdff dff_A_S3A9iaE13_0(.dout(w_G4_1[0]),.din(w_dff_A_S3A9iaE13_0),.clk(gclk));
	jdff dff_A_krEBoHMt1_0(.dout(w_dff_A_S3A9iaE13_0),.din(w_dff_A_krEBoHMt1_0),.clk(gclk));
	jdff dff_A_zbBOPd4Q6_0(.dout(w_dff_A_krEBoHMt1_0),.din(w_dff_A_zbBOPd4Q6_0),.clk(gclk));
	jdff dff_A_SL3qSCfQ3_0(.dout(w_dff_A_zbBOPd4Q6_0),.din(w_dff_A_SL3qSCfQ3_0),.clk(gclk));
	jdff dff_B_rZlufikp0_0(.din(n1155),.dout(w_dff_B_rZlufikp0_0),.clk(gclk));
	jdff dff_B_Z8QgmcpH3_0(.din(w_dff_B_rZlufikp0_0),.dout(w_dff_B_Z8QgmcpH3_0),.clk(gclk));
	jdff dff_B_Sx6bZPfX9_0(.din(w_dff_B_Z8QgmcpH3_0),.dout(w_dff_B_Sx6bZPfX9_0),.clk(gclk));
	jdff dff_B_tURWSTxm3_0(.din(w_dff_B_Sx6bZPfX9_0),.dout(w_dff_B_tURWSTxm3_0),.clk(gclk));
	jdff dff_B_EJIcXACC0_0(.din(w_dff_B_tURWSTxm3_0),.dout(w_dff_B_EJIcXACC0_0),.clk(gclk));
	jdff dff_B_RLQnn9YY0_0(.din(w_dff_B_EJIcXACC0_0),.dout(w_dff_B_RLQnn9YY0_0),.clk(gclk));
	jdff dff_B_R1vwRNSd9_0(.din(w_dff_B_RLQnn9YY0_0),.dout(w_dff_B_R1vwRNSd9_0),.clk(gclk));
	jdff dff_B_KkfVonDU0_0(.din(w_dff_B_R1vwRNSd9_0),.dout(w_dff_B_KkfVonDU0_0),.clk(gclk));
	jdff dff_B_UydwmAn19_0(.din(w_dff_B_KkfVonDU0_0),.dout(w_dff_B_UydwmAn19_0),.clk(gclk));
	jdff dff_B_KFyg94CR6_0(.din(w_dff_B_UydwmAn19_0),.dout(w_dff_B_KFyg94CR6_0),.clk(gclk));
	jdff dff_B_aieW1T711_0(.din(w_dff_B_KFyg94CR6_0),.dout(w_dff_B_aieW1T711_0),.clk(gclk));
	jdff dff_B_w7QhIpOV3_0(.din(w_dff_B_aieW1T711_0),.dout(w_dff_B_w7QhIpOV3_0),.clk(gclk));
	jdff dff_B_JFohs4FV4_1(.din(n1148),.dout(w_dff_B_JFohs4FV4_1),.clk(gclk));
	jdff dff_B_b8ZWHRwQ6_1(.din(w_dff_B_JFohs4FV4_1),.dout(w_dff_B_b8ZWHRwQ6_1),.clk(gclk));
	jdff dff_B_i6tiRbtz5_1(.din(w_dff_B_b8ZWHRwQ6_1),.dout(w_dff_B_i6tiRbtz5_1),.clk(gclk));
	jdff dff_B_azQH0x1a7_1(.din(w_dff_B_i6tiRbtz5_1),.dout(w_dff_B_azQH0x1a7_1),.clk(gclk));
	jdff dff_B_FsbrXkvc7_1(.din(w_dff_B_azQH0x1a7_1),.dout(w_dff_B_FsbrXkvc7_1),.clk(gclk));
	jdff dff_B_n1caYDXs8_1(.din(n1150),.dout(w_dff_B_n1caYDXs8_1),.clk(gclk));
	jdff dff_B_jOuKGlAG2_0(.din(n1144),.dout(w_dff_B_jOuKGlAG2_0),.clk(gclk));
	jdff dff_B_XofCy3am5_0(.din(w_dff_B_jOuKGlAG2_0),.dout(w_dff_B_XofCy3am5_0),.clk(gclk));
	jdff dff_B_aYYrDuJW6_0(.din(w_dff_B_XofCy3am5_0),.dout(w_dff_B_aYYrDuJW6_0),.clk(gclk));
	jdff dff_B_PBruMV9M2_0(.din(w_dff_B_aYYrDuJW6_0),.dout(w_dff_B_PBruMV9M2_0),.clk(gclk));
	jdff dff_B_HpBSRuLH3_0(.din(w_dff_B_PBruMV9M2_0),.dout(w_dff_B_HpBSRuLH3_0),.clk(gclk));
	jdff dff_B_5aYLOKsi5_0(.din(w_dff_B_HpBSRuLH3_0),.dout(w_dff_B_5aYLOKsi5_0),.clk(gclk));
	jdff dff_B_tIFftIpk1_0(.din(w_dff_B_5aYLOKsi5_0),.dout(w_dff_B_tIFftIpk1_0),.clk(gclk));
	jdff dff_B_zNJNcfz89_0(.din(w_dff_B_tIFftIpk1_0),.dout(w_dff_B_zNJNcfz89_0),.clk(gclk));
	jdff dff_B_ICcObu3u6_0(.din(w_dff_B_zNJNcfz89_0),.dout(w_dff_B_ICcObu3u6_0),.clk(gclk));
	jdff dff_B_MojCcEFQ2_0(.din(w_dff_B_ICcObu3u6_0),.dout(w_dff_B_MojCcEFQ2_0),.clk(gclk));
	jdff dff_B_1z8FhPUv6_0(.din(w_dff_B_MojCcEFQ2_0),.dout(w_dff_B_1z8FhPUv6_0),.clk(gclk));
	jdff dff_B_Jp3qyDQ02_0(.din(w_dff_B_1z8FhPUv6_0),.dout(w_dff_B_Jp3qyDQ02_0),.clk(gclk));
	jdff dff_B_5nfTkvUg1_0(.din(w_dff_B_Jp3qyDQ02_0),.dout(w_dff_B_5nfTkvUg1_0),.clk(gclk));
	jdff dff_B_7N6eNxPt9_0(.din(w_dff_B_5nfTkvUg1_0),.dout(w_dff_B_7N6eNxPt9_0),.clk(gclk));
	jdff dff_B_MWWNPNaA3_0(.din(w_dff_B_7N6eNxPt9_0),.dout(w_dff_B_MWWNPNaA3_0),.clk(gclk));
	jdff dff_B_FMrwp04V2_0(.din(w_dff_B_MWWNPNaA3_0),.dout(w_dff_B_FMrwp04V2_0),.clk(gclk));
	jdff dff_B_J0YdLulo1_1(.din(n1141),.dout(w_dff_B_J0YdLulo1_1),.clk(gclk));
	jdff dff_A_K6SzOKp15_0(.dout(w_n1142_0[0]),.din(w_dff_A_K6SzOKp15_0),.clk(gclk));
	jdff dff_A_qeirXqOk5_0(.dout(w_dff_A_K6SzOKp15_0),.din(w_dff_A_qeirXqOk5_0),.clk(gclk));
	jdff dff_A_osSimo5V6_0(.dout(w_dff_A_qeirXqOk5_0),.din(w_dff_A_osSimo5V6_0),.clk(gclk));
	jdff dff_A_aKgV9xIY9_0(.dout(w_G3717_0[0]),.din(w_dff_A_aKgV9xIY9_0),.clk(gclk));
	jdff dff_A_sGtT0UpU5_0(.dout(w_dff_A_aKgV9xIY9_0),.din(w_dff_A_sGtT0UpU5_0),.clk(gclk));
	jdff dff_A_wtCkzWpC0_0(.dout(w_dff_A_sGtT0UpU5_0),.din(w_dff_A_wtCkzWpC0_0),.clk(gclk));
	jdff dff_A_d2klbvkf6_0(.dout(w_dff_A_wtCkzWpC0_0),.din(w_dff_A_d2klbvkf6_0),.clk(gclk));
	jdff dff_A_j4F8Q4Q48_0(.dout(w_dff_A_d2klbvkf6_0),.din(w_dff_A_j4F8Q4Q48_0),.clk(gclk));
	jdff dff_A_KupFvMek0_0(.dout(w_G3724_0[0]),.din(w_dff_A_KupFvMek0_0),.clk(gclk));
	jdff dff_A_YMQddjrZ0_0(.dout(w_dff_A_KupFvMek0_0),.din(w_dff_A_YMQddjrZ0_0),.clk(gclk));
	jdff dff_A_neHuwbZB1_0(.dout(w_dff_A_YMQddjrZ0_0),.din(w_dff_A_neHuwbZB1_0),.clk(gclk));
	jdff dff_A_vCMXz4iL1_0(.dout(w_dff_A_neHuwbZB1_0),.din(w_dff_A_vCMXz4iL1_0),.clk(gclk));
	jdff dff_A_bkx6wXmx2_2(.dout(w_G3724_0[2]),.din(w_dff_A_bkx6wXmx2_2),.clk(gclk));
	jdff dff_A_INHrCEno2_2(.dout(w_dff_A_bkx6wXmx2_2),.din(w_dff_A_INHrCEno2_2),.clk(gclk));
	jdff dff_A_yAzh50XK3_2(.dout(w_dff_A_INHrCEno2_2),.din(w_dff_A_yAzh50XK3_2),.clk(gclk));
	jdff dff_A_fRLBZb3v8_2(.dout(w_dff_A_yAzh50XK3_2),.din(w_dff_A_fRLBZb3v8_2),.clk(gclk));
	jdff dff_A_HVpc9jXd3_2(.dout(w_dff_A_fRLBZb3v8_2),.din(w_dff_A_HVpc9jXd3_2),.clk(gclk));
	jdff dff_A_URkEzGnw4_2(.dout(w_dff_A_HVpc9jXd3_2),.din(w_dff_A_URkEzGnw4_2),.clk(gclk));
	jdff dff_A_DBvuUKK06_2(.dout(w_dff_A_URkEzGnw4_2),.din(w_dff_A_DBvuUKK06_2),.clk(gclk));
	jdff dff_A_8RgLcLau1_2(.dout(w_dff_A_DBvuUKK06_2),.din(w_dff_A_8RgLcLau1_2),.clk(gclk));
	jdff dff_A_T83pYknB7_2(.dout(w_dff_A_8RgLcLau1_2),.din(w_dff_A_T83pYknB7_2),.clk(gclk));
	jdff dff_A_8zQhIFMF0_2(.dout(w_dff_A_T83pYknB7_2),.din(w_dff_A_8zQhIFMF0_2),.clk(gclk));
	jdff dff_A_GIzrlDgr3_2(.dout(w_dff_A_8zQhIFMF0_2),.din(w_dff_A_GIzrlDgr3_2),.clk(gclk));
	jdff dff_A_bbsteKd83_2(.dout(w_dff_A_GIzrlDgr3_2),.din(w_dff_A_bbsteKd83_2),.clk(gclk));
	jdff dff_A_9wEnWf2n6_2(.dout(w_dff_A_bbsteKd83_2),.din(w_dff_A_9wEnWf2n6_2),.clk(gclk));
	jdff dff_A_007DtaO53_2(.dout(w_dff_A_9wEnWf2n6_2),.din(w_dff_A_007DtaO53_2),.clk(gclk));
	jdff dff_A_afgfJBNd1_2(.dout(w_dff_A_007DtaO53_2),.din(w_dff_A_afgfJBNd1_2),.clk(gclk));
	jdff dff_A_awaVXosT6_2(.dout(w_dff_A_afgfJBNd1_2),.din(w_dff_A_awaVXosT6_2),.clk(gclk));
	jdff dff_A_NZxTyMrq2_2(.dout(w_dff_A_awaVXosT6_2),.din(w_dff_A_NZxTyMrq2_2),.clk(gclk));
	jdff dff_A_Y3km0hto5_2(.dout(w_dff_A_NZxTyMrq2_2),.din(w_dff_A_Y3km0hto5_2),.clk(gclk));
	jdff dff_A_CyhbJpPf8_0(.dout(w_G132_0[0]),.din(w_dff_A_CyhbJpPf8_0),.clk(gclk));
	jdff dff_A_mp7Tnzcw8_0(.dout(w_dff_A_CyhbJpPf8_0),.din(w_dff_A_mp7Tnzcw8_0),.clk(gclk));
	jdff dff_A_gsfJ6xKn8_0(.dout(w_dff_A_mp7Tnzcw8_0),.din(w_dff_A_gsfJ6xKn8_0),.clk(gclk));
	jdff dff_A_O9AgyIXz0_0(.dout(w_dff_A_gsfJ6xKn8_0),.din(w_dff_A_O9AgyIXz0_0),.clk(gclk));
	jdff dff_A_oOM8QH7N3_0(.dout(w_dff_A_O9AgyIXz0_0),.din(w_dff_A_oOM8QH7N3_0),.clk(gclk));
	jdff dff_A_GoffM0QW2_0(.dout(w_dff_A_oOM8QH7N3_0),.din(w_dff_A_GoffM0QW2_0),.clk(gclk));
	jdff dff_A_YEkxEUIG5_0(.dout(w_dff_A_GoffM0QW2_0),.din(w_dff_A_YEkxEUIG5_0),.clk(gclk));
	jdff dff_A_yt364Pk02_0(.dout(w_dff_A_YEkxEUIG5_0),.din(w_dff_A_yt364Pk02_0),.clk(gclk));
	jdff dff_A_ALYqXm6s4_0(.dout(w_dff_A_yt364Pk02_0),.din(w_dff_A_ALYqXm6s4_0),.clk(gclk));
	jdff dff_A_YzTymrLW3_0(.dout(w_dff_A_ALYqXm6s4_0),.din(w_dff_A_YzTymrLW3_0),.clk(gclk));
	jdff dff_A_zzsJyB2j0_0(.dout(w_dff_A_YzTymrLW3_0),.din(w_dff_A_zzsJyB2j0_0),.clk(gclk));
	jdff dff_A_ZG2Bd2je4_0(.dout(w_dff_A_zzsJyB2j0_0),.din(w_dff_A_ZG2Bd2je4_0),.clk(gclk));
	jdff dff_A_de4oxTsm6_0(.dout(w_dff_A_ZG2Bd2je4_0),.din(w_dff_A_de4oxTsm6_0),.clk(gclk));
	jdff dff_B_eXbFNvuK9_2(.din(G132),.dout(w_dff_B_eXbFNvuK9_2),.clk(gclk));
	jdff dff_B_PQ2AeFZf3_2(.din(w_dff_B_eXbFNvuK9_2),.dout(w_dff_B_PQ2AeFZf3_2),.clk(gclk));
	jdff dff_B_i0Dq756B2_2(.din(w_dff_B_PQ2AeFZf3_2),.dout(w_dff_B_i0Dq756B2_2),.clk(gclk));
	jdff dff_B_9S8cjbQD0_1(.din(n1184),.dout(w_dff_B_9S8cjbQD0_1),.clk(gclk));
	jdff dff_B_U0OOsFzQ1_0(.din(n1189),.dout(w_dff_B_U0OOsFzQ1_0),.clk(gclk));
	jdff dff_B_Fk7TrJzz6_0(.din(w_dff_B_U0OOsFzQ1_0),.dout(w_dff_B_Fk7TrJzz6_0),.clk(gclk));
	jdff dff_B_NHXjAi4F9_0(.din(n1187),.dout(w_dff_B_NHXjAi4F9_0),.clk(gclk));
	jdff dff_A_66KJWVwp8_0(.dout(w_G601_0),.din(w_dff_A_66KJWVwp8_0),.clk(gclk));
	jdff dff_B_UFlG5cKM3_1(.din(n656),.dout(w_dff_B_UFlG5cKM3_1),.clk(gclk));
	jdff dff_A_AS70YKql5_0(.dout(w_n671_0[0]),.din(w_dff_A_AS70YKql5_0),.clk(gclk));
	jdff dff_B_QE8FytI96_1(.din(n665),.dout(w_dff_B_QE8FytI96_1),.clk(gclk));
	jdff dff_B_FhiAzXBB6_1(.din(n907),.dout(w_dff_B_FhiAzXBB6_1),.clk(gclk));
	jdff dff_B_g1TD5Row9_1(.din(n909),.dout(w_dff_B_g1TD5Row9_1),.clk(gclk));
	jdff dff_B_JEPeCu9J0_1(.din(w_dff_B_g1TD5Row9_1),.dout(w_dff_B_JEPeCu9J0_1),.clk(gclk));
	jdff dff_B_ZG2jwuz38_0(.din(n910),.dout(w_dff_B_ZG2jwuz38_0),.clk(gclk));
	jdff dff_B_zQ4MytPc7_1(.din(n908),.dout(w_dff_B_zQ4MytPc7_1),.clk(gclk));
	jdff dff_B_jyM7J1ZV9_0(.din(n904),.dout(w_dff_B_jyM7J1ZV9_0),.clk(gclk));
	jdff dff_A_7RobHvig9_0(.dout(w_G369_0[0]),.din(w_dff_A_7RobHvig9_0),.clk(gclk));
	jdff dff_A_jNOtSQy00_0(.dout(w_n621_1[0]),.din(w_dff_A_jNOtSQy00_0),.clk(gclk));
	jdff dff_A_3vlUtqyv9_0(.dout(w_dff_A_jNOtSQy00_0),.din(w_dff_A_3vlUtqyv9_0),.clk(gclk));
	jdff dff_A_XwwuUsln0_0(.dout(w_dff_A_3vlUtqyv9_0),.din(w_dff_A_XwwuUsln0_0),.clk(gclk));
	jdff dff_B_MvjSQb1U2_0(.din(n921),.dout(w_dff_B_MvjSQb1U2_0),.clk(gclk));
	jdff dff_A_9cjRjcFv5_0(.dout(w_G289_0[0]),.din(w_dff_A_9cjRjcFv5_0),.clk(gclk));
	jdff dff_B_Ut5Bnd300_0(.din(n1224),.dout(w_dff_B_Ut5Bnd300_0),.clk(gclk));
	jdff dff_B_bhGgs7uv5_0(.din(w_dff_B_Ut5Bnd300_0),.dout(w_dff_B_bhGgs7uv5_0),.clk(gclk));
	jdff dff_B_UFJ4mJEx3_0(.din(w_dff_B_bhGgs7uv5_0),.dout(w_dff_B_UFJ4mJEx3_0),.clk(gclk));
	jdff dff_B_z9LDfLam6_0(.din(w_dff_B_UFJ4mJEx3_0),.dout(w_dff_B_z9LDfLam6_0),.clk(gclk));
	jdff dff_B_pi18C67K0_0(.din(w_dff_B_z9LDfLam6_0),.dout(w_dff_B_pi18C67K0_0),.clk(gclk));
	jdff dff_B_58hRtFy36_0(.din(w_dff_B_pi18C67K0_0),.dout(w_dff_B_58hRtFy36_0),.clk(gclk));
	jdff dff_B_s7n5lhpd8_0(.din(w_dff_B_58hRtFy36_0),.dout(w_dff_B_s7n5lhpd8_0),.clk(gclk));
	jdff dff_B_dtPFA2SD7_0(.din(w_dff_B_s7n5lhpd8_0),.dout(w_dff_B_dtPFA2SD7_0),.clk(gclk));
	jdff dff_B_9bPkADha1_0(.din(w_dff_B_dtPFA2SD7_0),.dout(w_dff_B_9bPkADha1_0),.clk(gclk));
	jdff dff_B_Yh1o87DF4_0(.din(w_dff_B_9bPkADha1_0),.dout(w_dff_B_Yh1o87DF4_0),.clk(gclk));
	jdff dff_B_q9XTkk1d1_0(.din(w_dff_B_Yh1o87DF4_0),.dout(w_dff_B_q9XTkk1d1_0),.clk(gclk));
	jdff dff_B_GU6O5mJw0_0(.din(w_dff_B_q9XTkk1d1_0),.dout(w_dff_B_GU6O5mJw0_0),.clk(gclk));
	jdff dff_B_QNxPHZKg8_0(.din(w_dff_B_GU6O5mJw0_0),.dout(w_dff_B_QNxPHZKg8_0),.clk(gclk));
	jdff dff_B_Wc5IvLvh3_0(.din(w_dff_B_QNxPHZKg8_0),.dout(w_dff_B_Wc5IvLvh3_0),.clk(gclk));
	jdff dff_B_FlTFRELI9_0(.din(w_dff_B_Wc5IvLvh3_0),.dout(w_dff_B_FlTFRELI9_0),.clk(gclk));
	jdff dff_B_aEuozjhT5_0(.din(w_dff_B_FlTFRELI9_0),.dout(w_dff_B_aEuozjhT5_0),.clk(gclk));
	jdff dff_B_I2ermMkl7_0(.din(w_dff_B_aEuozjhT5_0),.dout(w_dff_B_I2ermMkl7_0),.clk(gclk));
	jdff dff_B_2C2LaIa98_0(.din(n1223),.dout(w_dff_B_2C2LaIa98_0),.clk(gclk));
	jdff dff_B_K8TlxGVZ4_0(.din(n1231),.dout(w_dff_B_K8TlxGVZ4_0),.clk(gclk));
	jdff dff_B_vTLCDkIb0_0(.din(w_dff_B_K8TlxGVZ4_0),.dout(w_dff_B_vTLCDkIb0_0),.clk(gclk));
	jdff dff_B_Gpl903cN2_0(.din(w_dff_B_vTLCDkIb0_0),.dout(w_dff_B_Gpl903cN2_0),.clk(gclk));
	jdff dff_B_OtsaWbz08_0(.din(w_dff_B_Gpl903cN2_0),.dout(w_dff_B_OtsaWbz08_0),.clk(gclk));
	jdff dff_B_ZhQRZYta7_0(.din(w_dff_B_OtsaWbz08_0),.dout(w_dff_B_ZhQRZYta7_0),.clk(gclk));
	jdff dff_B_ofde5ZOi0_0(.din(w_dff_B_ZhQRZYta7_0),.dout(w_dff_B_ofde5ZOi0_0),.clk(gclk));
	jdff dff_B_b4G56N331_0(.din(w_dff_B_ofde5ZOi0_0),.dout(w_dff_B_b4G56N331_0),.clk(gclk));
	jdff dff_B_uPHCEmRC4_0(.din(w_dff_B_b4G56N331_0),.dout(w_dff_B_uPHCEmRC4_0),.clk(gclk));
	jdff dff_B_F12qWcb15_0(.din(w_dff_B_uPHCEmRC4_0),.dout(w_dff_B_F12qWcb15_0),.clk(gclk));
	jdff dff_B_nU5g4WdW9_0(.din(w_dff_B_F12qWcb15_0),.dout(w_dff_B_nU5g4WdW9_0),.clk(gclk));
	jdff dff_B_X5lc8ERA2_0(.din(w_dff_B_nU5g4WdW9_0),.dout(w_dff_B_X5lc8ERA2_0),.clk(gclk));
	jdff dff_B_E4BG8Ayw5_0(.din(w_dff_B_X5lc8ERA2_0),.dout(w_dff_B_E4BG8Ayw5_0),.clk(gclk));
	jdff dff_B_IOi2av3N4_0(.din(w_dff_B_E4BG8Ayw5_0),.dout(w_dff_B_IOi2av3N4_0),.clk(gclk));
	jdff dff_B_DZcULegl0_0(.din(w_dff_B_IOi2av3N4_0),.dout(w_dff_B_DZcULegl0_0),.clk(gclk));
	jdff dff_B_Qx7oNdWy9_0(.din(w_dff_B_DZcULegl0_0),.dout(w_dff_B_Qx7oNdWy9_0),.clk(gclk));
	jdff dff_B_0ztLduFz5_0(.din(w_dff_B_Qx7oNdWy9_0),.dout(w_dff_B_0ztLduFz5_0),.clk(gclk));
	jdff dff_B_nsPRMNxz1_0(.din(w_dff_B_0ztLduFz5_0),.dout(w_dff_B_nsPRMNxz1_0),.clk(gclk));
	jdff dff_B_Ih13jZBk8_0(.din(n1230),.dout(w_dff_B_Ih13jZBk8_0),.clk(gclk));
	jdff dff_B_skpGvuxw4_2(.din(G106),.dout(w_dff_B_skpGvuxw4_2),.clk(gclk));
	jdff dff_B_G5rMUXF48_2(.din(G109),.dout(w_dff_B_G5rMUXF48_2),.clk(gclk));
	jdff dff_B_pc46jYw56_2(.din(w_dff_B_G5rMUXF48_2),.dout(w_dff_B_pc46jYw56_2),.clk(gclk));
	jdff dff_B_xiEtWRdJ3_0(.din(n1239),.dout(w_dff_B_xiEtWRdJ3_0),.clk(gclk));
	jdff dff_B_0QXWl8xb1_0(.din(w_dff_B_xiEtWRdJ3_0),.dout(w_dff_B_0QXWl8xb1_0),.clk(gclk));
	jdff dff_B_axFCVXAq9_0(.din(w_dff_B_0QXWl8xb1_0),.dout(w_dff_B_axFCVXAq9_0),.clk(gclk));
	jdff dff_B_q14bpZdM0_0(.din(w_dff_B_axFCVXAq9_0),.dout(w_dff_B_q14bpZdM0_0),.clk(gclk));
	jdff dff_B_xKfuQ16J7_0(.din(w_dff_B_q14bpZdM0_0),.dout(w_dff_B_xKfuQ16J7_0),.clk(gclk));
	jdff dff_B_XW5a9qpS3_0(.din(w_dff_B_xKfuQ16J7_0),.dout(w_dff_B_XW5a9qpS3_0),.clk(gclk));
	jdff dff_B_qoNtuyfN5_0(.din(w_dff_B_XW5a9qpS3_0),.dout(w_dff_B_qoNtuyfN5_0),.clk(gclk));
	jdff dff_B_lo5eZZYj4_0(.din(w_dff_B_qoNtuyfN5_0),.dout(w_dff_B_lo5eZZYj4_0),.clk(gclk));
	jdff dff_B_wR7cML9x6_0(.din(w_dff_B_lo5eZZYj4_0),.dout(w_dff_B_wR7cML9x6_0),.clk(gclk));
	jdff dff_B_rw2nfGOk0_0(.din(w_dff_B_wR7cML9x6_0),.dout(w_dff_B_rw2nfGOk0_0),.clk(gclk));
	jdff dff_B_sZjXSQc00_0(.din(w_dff_B_rw2nfGOk0_0),.dout(w_dff_B_sZjXSQc00_0),.clk(gclk));
	jdff dff_B_1MYmZ2Hh8_0(.din(w_dff_B_sZjXSQc00_0),.dout(w_dff_B_1MYmZ2Hh8_0),.clk(gclk));
	jdff dff_B_vZJ4MQiT0_0(.din(w_dff_B_1MYmZ2Hh8_0),.dout(w_dff_B_vZJ4MQiT0_0),.clk(gclk));
	jdff dff_B_zU4wzDf07_0(.din(w_dff_B_vZJ4MQiT0_0),.dout(w_dff_B_zU4wzDf07_0),.clk(gclk));
	jdff dff_B_2rdPzQxt5_0(.din(w_dff_B_zU4wzDf07_0),.dout(w_dff_B_2rdPzQxt5_0),.clk(gclk));
	jdff dff_B_wsrvTRFU1_0(.din(w_dff_B_2rdPzQxt5_0),.dout(w_dff_B_wsrvTRFU1_0),.clk(gclk));
	jdff dff_B_bKng4ZYj7_0(.din(n1238),.dout(w_dff_B_bKng4ZYj7_0),.clk(gclk));
	jdff dff_B_7sDRp8Pe6_0(.din(n1248),.dout(w_dff_B_7sDRp8Pe6_0),.clk(gclk));
	jdff dff_B_jcLLwElZ8_0(.din(w_dff_B_7sDRp8Pe6_0),.dout(w_dff_B_jcLLwElZ8_0),.clk(gclk));
	jdff dff_B_X3W3I4CG0_0(.din(w_dff_B_jcLLwElZ8_0),.dout(w_dff_B_X3W3I4CG0_0),.clk(gclk));
	jdff dff_B_bxdHV3Tb7_0(.din(w_dff_B_X3W3I4CG0_0),.dout(w_dff_B_bxdHV3Tb7_0),.clk(gclk));
	jdff dff_B_Y7YCJUoX5_0(.din(w_dff_B_bxdHV3Tb7_0),.dout(w_dff_B_Y7YCJUoX5_0),.clk(gclk));
	jdff dff_B_qlpAoWjL2_0(.din(w_dff_B_Y7YCJUoX5_0),.dout(w_dff_B_qlpAoWjL2_0),.clk(gclk));
	jdff dff_B_7MN0tEj44_0(.din(w_dff_B_qlpAoWjL2_0),.dout(w_dff_B_7MN0tEj44_0),.clk(gclk));
	jdff dff_B_xl0qGUAI6_0(.din(w_dff_B_7MN0tEj44_0),.dout(w_dff_B_xl0qGUAI6_0),.clk(gclk));
	jdff dff_B_rM0t2XlX6_0(.din(w_dff_B_xl0qGUAI6_0),.dout(w_dff_B_rM0t2XlX6_0),.clk(gclk));
	jdff dff_B_FAavZQ1G2_0(.din(w_dff_B_rM0t2XlX6_0),.dout(w_dff_B_FAavZQ1G2_0),.clk(gclk));
	jdff dff_B_4j68Ncvl4_0(.din(w_dff_B_FAavZQ1G2_0),.dout(w_dff_B_4j68Ncvl4_0),.clk(gclk));
	jdff dff_B_vwzFit9Q6_0(.din(w_dff_B_4j68Ncvl4_0),.dout(w_dff_B_vwzFit9Q6_0),.clk(gclk));
	jdff dff_B_Hj7tOlfS8_0(.din(w_dff_B_vwzFit9Q6_0),.dout(w_dff_B_Hj7tOlfS8_0),.clk(gclk));
	jdff dff_B_nBFTz95a8_0(.din(w_dff_B_Hj7tOlfS8_0),.dout(w_dff_B_nBFTz95a8_0),.clk(gclk));
	jdff dff_B_CiOblOqN6_0(.din(w_dff_B_nBFTz95a8_0),.dout(w_dff_B_CiOblOqN6_0),.clk(gclk));
	jdff dff_B_bOm6xuOr3_0(.din(w_dff_B_CiOblOqN6_0),.dout(w_dff_B_bOm6xuOr3_0),.clk(gclk));
	jdff dff_B_uwUSbe004_0(.din(n1247),.dout(w_dff_B_uwUSbe004_0),.clk(gclk));
	jdff dff_A_dkRHlgvt0_2(.dout(w_n797_2[2]),.din(w_dff_A_dkRHlgvt0_2),.clk(gclk));
	jdff dff_A_ZgzYrzSU2_2(.dout(w_n793_2[2]),.din(w_dff_A_ZgzYrzSU2_2),.clk(gclk));
	jdff dff_B_qYJGFmw80_0(.din(n1257),.dout(w_dff_B_qYJGFmw80_0),.clk(gclk));
	jdff dff_B_0xGmt1ef9_0(.din(w_dff_B_qYJGFmw80_0),.dout(w_dff_B_0xGmt1ef9_0),.clk(gclk));
	jdff dff_B_WlUJvoLS4_0(.din(w_dff_B_0xGmt1ef9_0),.dout(w_dff_B_WlUJvoLS4_0),.clk(gclk));
	jdff dff_B_lRZuuHgY9_0(.din(w_dff_B_WlUJvoLS4_0),.dout(w_dff_B_lRZuuHgY9_0),.clk(gclk));
	jdff dff_B_f1jKh4Xk8_0(.din(w_dff_B_lRZuuHgY9_0),.dout(w_dff_B_f1jKh4Xk8_0),.clk(gclk));
	jdff dff_B_hnUKu0HQ6_0(.din(w_dff_B_f1jKh4Xk8_0),.dout(w_dff_B_hnUKu0HQ6_0),.clk(gclk));
	jdff dff_B_jFCmLIkr3_0(.din(w_dff_B_hnUKu0HQ6_0),.dout(w_dff_B_jFCmLIkr3_0),.clk(gclk));
	jdff dff_B_zEnMY9dx2_0(.din(w_dff_B_jFCmLIkr3_0),.dout(w_dff_B_zEnMY9dx2_0),.clk(gclk));
	jdff dff_B_Tg6LPpdP0_0(.din(w_dff_B_zEnMY9dx2_0),.dout(w_dff_B_Tg6LPpdP0_0),.clk(gclk));
	jdff dff_B_gP81Hn0u5_0(.din(w_dff_B_Tg6LPpdP0_0),.dout(w_dff_B_gP81Hn0u5_0),.clk(gclk));
	jdff dff_B_o0wuvb1b9_0(.din(w_dff_B_gP81Hn0u5_0),.dout(w_dff_B_o0wuvb1b9_0),.clk(gclk));
	jdff dff_B_IIGwLfn26_0(.din(w_dff_B_o0wuvb1b9_0),.dout(w_dff_B_IIGwLfn26_0),.clk(gclk));
	jdff dff_B_ohzHHHUB2_0(.din(w_dff_B_IIGwLfn26_0),.dout(w_dff_B_ohzHHHUB2_0),.clk(gclk));
	jdff dff_B_q77aGSrk7_0(.din(w_dff_B_ohzHHHUB2_0),.dout(w_dff_B_q77aGSrk7_0),.clk(gclk));
	jdff dff_B_t94d85kX8_0(.din(w_dff_B_q77aGSrk7_0),.dout(w_dff_B_t94d85kX8_0),.clk(gclk));
	jdff dff_B_5jWzyvJG7_0(.din(n1256),.dout(w_dff_B_5jWzyvJG7_0),.clk(gclk));
	jdff dff_B_NypKMHDv5_0(.din(n1264),.dout(w_dff_B_NypKMHDv5_0),.clk(gclk));
	jdff dff_B_PoebvJ2P8_0(.din(w_dff_B_NypKMHDv5_0),.dout(w_dff_B_PoebvJ2P8_0),.clk(gclk));
	jdff dff_B_8fRSbgka8_0(.din(w_dff_B_PoebvJ2P8_0),.dout(w_dff_B_8fRSbgka8_0),.clk(gclk));
	jdff dff_B_UmrBnTNH2_0(.din(w_dff_B_8fRSbgka8_0),.dout(w_dff_B_UmrBnTNH2_0),.clk(gclk));
	jdff dff_B_v9cFAZLn5_0(.din(w_dff_B_UmrBnTNH2_0),.dout(w_dff_B_v9cFAZLn5_0),.clk(gclk));
	jdff dff_B_zqDTnKjs4_0(.din(w_dff_B_v9cFAZLn5_0),.dout(w_dff_B_zqDTnKjs4_0),.clk(gclk));
	jdff dff_B_4vle1Qcn3_0(.din(w_dff_B_zqDTnKjs4_0),.dout(w_dff_B_4vle1Qcn3_0),.clk(gclk));
	jdff dff_B_k16y28oq0_0(.din(w_dff_B_4vle1Qcn3_0),.dout(w_dff_B_k16y28oq0_0),.clk(gclk));
	jdff dff_B_uv1yIhmW3_0(.din(w_dff_B_k16y28oq0_0),.dout(w_dff_B_uv1yIhmW3_0),.clk(gclk));
	jdff dff_B_2jKjYMzD8_0(.din(w_dff_B_uv1yIhmW3_0),.dout(w_dff_B_2jKjYMzD8_0),.clk(gclk));
	jdff dff_B_ywD1xsZl0_0(.din(w_dff_B_2jKjYMzD8_0),.dout(w_dff_B_ywD1xsZl0_0),.clk(gclk));
	jdff dff_B_Z0ns3pPN8_0(.din(w_dff_B_ywD1xsZl0_0),.dout(w_dff_B_Z0ns3pPN8_0),.clk(gclk));
	jdff dff_B_g4KtRWBn3_0(.din(w_dff_B_Z0ns3pPN8_0),.dout(w_dff_B_g4KtRWBn3_0),.clk(gclk));
	jdff dff_B_1DRwYKOB2_0(.din(w_dff_B_g4KtRWBn3_0),.dout(w_dff_B_1DRwYKOB2_0),.clk(gclk));
	jdff dff_B_77g5Gz7d0_0(.din(w_dff_B_1DRwYKOB2_0),.dout(w_dff_B_77g5Gz7d0_0),.clk(gclk));
	jdff dff_B_LhUW3Ydi0_0(.din(w_dff_B_77g5Gz7d0_0),.dout(w_dff_B_LhUW3Ydi0_0),.clk(gclk));
	jdff dff_B_Izl0K9OX4_0(.din(n1263),.dout(w_dff_B_Izl0K9OX4_0),.clk(gclk));
	jdff dff_B_zwPJdQEF4_2(.din(G49),.dout(w_dff_B_zwPJdQEF4_2),.clk(gclk));
	jdff dff_B_eXvMRe1b0_2(.din(G46),.dout(w_dff_B_eXvMRe1b0_2),.clk(gclk));
	jdff dff_B_SYbYFckq7_2(.din(w_dff_B_eXvMRe1b0_2),.dout(w_dff_B_SYbYFckq7_2),.clk(gclk));
	jdff dff_B_8a1wdmuh6_0(.din(n1271),.dout(w_dff_B_8a1wdmuh6_0),.clk(gclk));
	jdff dff_B_LcHVNjN99_0(.din(w_dff_B_8a1wdmuh6_0),.dout(w_dff_B_LcHVNjN99_0),.clk(gclk));
	jdff dff_B_18MsEnw70_0(.din(w_dff_B_LcHVNjN99_0),.dout(w_dff_B_18MsEnw70_0),.clk(gclk));
	jdff dff_B_HVS95MvC7_0(.din(w_dff_B_18MsEnw70_0),.dout(w_dff_B_HVS95MvC7_0),.clk(gclk));
	jdff dff_B_GGddtJoi9_0(.din(w_dff_B_HVS95MvC7_0),.dout(w_dff_B_GGddtJoi9_0),.clk(gclk));
	jdff dff_B_fal9RzBR4_0(.din(w_dff_B_GGddtJoi9_0),.dout(w_dff_B_fal9RzBR4_0),.clk(gclk));
	jdff dff_B_L6FrlyfN6_0(.din(w_dff_B_fal9RzBR4_0),.dout(w_dff_B_L6FrlyfN6_0),.clk(gclk));
	jdff dff_B_OxoekeWa1_0(.din(w_dff_B_L6FrlyfN6_0),.dout(w_dff_B_OxoekeWa1_0),.clk(gclk));
	jdff dff_B_2Kc6ThxV7_0(.din(w_dff_B_OxoekeWa1_0),.dout(w_dff_B_2Kc6ThxV7_0),.clk(gclk));
	jdff dff_B_YI2taczn0_0(.din(w_dff_B_2Kc6ThxV7_0),.dout(w_dff_B_YI2taczn0_0),.clk(gclk));
	jdff dff_B_Fj3NFwt24_0(.din(w_dff_B_YI2taczn0_0),.dout(w_dff_B_Fj3NFwt24_0),.clk(gclk));
	jdff dff_B_uNgBiU0g9_0(.din(w_dff_B_Fj3NFwt24_0),.dout(w_dff_B_uNgBiU0g9_0),.clk(gclk));
	jdff dff_B_vRurAE3o3_0(.din(w_dff_B_uNgBiU0g9_0),.dout(w_dff_B_vRurAE3o3_0),.clk(gclk));
	jdff dff_B_UrgNl8Ee5_0(.din(w_dff_B_vRurAE3o3_0),.dout(w_dff_B_UrgNl8Ee5_0),.clk(gclk));
	jdff dff_B_OftxRVgy5_0(.din(w_dff_B_UrgNl8Ee5_0),.dout(w_dff_B_OftxRVgy5_0),.clk(gclk));
	jdff dff_B_aiw9eHOp9_0(.din(w_dff_B_OftxRVgy5_0),.dout(w_dff_B_aiw9eHOp9_0),.clk(gclk));
	jdff dff_B_jlLPp9Vx4_0(.din(n1270),.dout(w_dff_B_jlLPp9Vx4_0),.clk(gclk));
	jdff dff_B_mOQjkljC0_2(.din(G103),.dout(w_dff_B_mOQjkljC0_2),.clk(gclk));
	jdff dff_B_zoqcHgRF3_2(.din(G100),.dout(w_dff_B_zoqcHgRF3_2),.clk(gclk));
	jdff dff_B_0gLVztIc0_2(.din(w_dff_B_zoqcHgRF3_2),.dout(w_dff_B_0gLVztIc0_2),.clk(gclk));
	jdff dff_A_YZB8mdmT1_2(.dout(w_n843_2[2]),.din(w_dff_A_YZB8mdmT1_2),.clk(gclk));
	jdff dff_A_WCC2ZLwE1_2(.dout(w_n840_2[2]),.din(w_dff_A_WCC2ZLwE1_2),.clk(gclk));
	jdff dff_B_pBf9AXCt4_0(.din(n1278),.dout(w_dff_B_pBf9AXCt4_0),.clk(gclk));
	jdff dff_B_yMNdH2HB6_0(.din(w_dff_B_pBf9AXCt4_0),.dout(w_dff_B_yMNdH2HB6_0),.clk(gclk));
	jdff dff_B_hjkvwDCd0_0(.din(w_dff_B_yMNdH2HB6_0),.dout(w_dff_B_hjkvwDCd0_0),.clk(gclk));
	jdff dff_B_AcGrsj9n5_0(.din(w_dff_B_hjkvwDCd0_0),.dout(w_dff_B_AcGrsj9n5_0),.clk(gclk));
	jdff dff_B_xrmpRsv10_0(.din(w_dff_B_AcGrsj9n5_0),.dout(w_dff_B_xrmpRsv10_0),.clk(gclk));
	jdff dff_B_3dgRN1Um7_0(.din(w_dff_B_xrmpRsv10_0),.dout(w_dff_B_3dgRN1Um7_0),.clk(gclk));
	jdff dff_B_mWlX1zib4_0(.din(w_dff_B_3dgRN1Um7_0),.dout(w_dff_B_mWlX1zib4_0),.clk(gclk));
	jdff dff_B_XBWApV9K6_0(.din(w_dff_B_mWlX1zib4_0),.dout(w_dff_B_XBWApV9K6_0),.clk(gclk));
	jdff dff_B_QfUT9LvJ3_0(.din(w_dff_B_XBWApV9K6_0),.dout(w_dff_B_QfUT9LvJ3_0),.clk(gclk));
	jdff dff_B_ciLEGZ418_0(.din(w_dff_B_QfUT9LvJ3_0),.dout(w_dff_B_ciLEGZ418_0),.clk(gclk));
	jdff dff_B_AlFxUvzv6_0(.din(w_dff_B_ciLEGZ418_0),.dout(w_dff_B_AlFxUvzv6_0),.clk(gclk));
	jdff dff_B_HeI2mYQu0_0(.din(w_dff_B_AlFxUvzv6_0),.dout(w_dff_B_HeI2mYQu0_0),.clk(gclk));
	jdff dff_B_MziJslA06_0(.din(w_dff_B_HeI2mYQu0_0),.dout(w_dff_B_MziJslA06_0),.clk(gclk));
	jdff dff_B_VVs6pJHk9_0(.din(w_dff_B_MziJslA06_0),.dout(w_dff_B_VVs6pJHk9_0),.clk(gclk));
	jdff dff_B_pcFZ3uXV4_0(.din(w_dff_B_VVs6pJHk9_0),.dout(w_dff_B_pcFZ3uXV4_0),.clk(gclk));
	jdff dff_B_vi4xFXql7_0(.din(n1277),.dout(w_dff_B_vi4xFXql7_0),.clk(gclk));
	jdff dff_B_cQ9zOYqq2_2(.din(G40),.dout(w_dff_B_cQ9zOYqq2_2),.clk(gclk));
	jdff dff_B_QWTeqsKZ6_2(.din(G91),.dout(w_dff_B_QWTeqsKZ6_2),.clk(gclk));
	jdff dff_B_jN6unUfh7_2(.din(w_dff_B_QWTeqsKZ6_2),.dout(w_dff_B_jN6unUfh7_2),.clk(gclk));
	jdff dff_B_Ow9FdZNy8_0(.din(n1285),.dout(w_dff_B_Ow9FdZNy8_0),.clk(gclk));
	jdff dff_B_YGPUoZBU2_0(.din(w_dff_B_Ow9FdZNy8_0),.dout(w_dff_B_YGPUoZBU2_0),.clk(gclk));
	jdff dff_B_rNED4cpP6_0(.din(w_dff_B_YGPUoZBU2_0),.dout(w_dff_B_rNED4cpP6_0),.clk(gclk));
	jdff dff_B_ttIkTcL76_0(.din(w_dff_B_rNED4cpP6_0),.dout(w_dff_B_ttIkTcL76_0),.clk(gclk));
	jdff dff_B_83KDtTui9_0(.din(w_dff_B_ttIkTcL76_0),.dout(w_dff_B_83KDtTui9_0),.clk(gclk));
	jdff dff_B_hUY0udmf3_0(.din(w_dff_B_83KDtTui9_0),.dout(w_dff_B_hUY0udmf3_0),.clk(gclk));
	jdff dff_B_hEznpjwG7_0(.din(w_dff_B_hUY0udmf3_0),.dout(w_dff_B_hEznpjwG7_0),.clk(gclk));
	jdff dff_B_wcQSsuKc3_0(.din(w_dff_B_hEznpjwG7_0),.dout(w_dff_B_wcQSsuKc3_0),.clk(gclk));
	jdff dff_B_RcKiMlGo0_0(.din(w_dff_B_wcQSsuKc3_0),.dout(w_dff_B_RcKiMlGo0_0),.clk(gclk));
	jdff dff_B_7EqxGuFx2_0(.din(w_dff_B_RcKiMlGo0_0),.dout(w_dff_B_7EqxGuFx2_0),.clk(gclk));
	jdff dff_B_v6JDwg0L9_0(.din(w_dff_B_7EqxGuFx2_0),.dout(w_dff_B_v6JDwg0L9_0),.clk(gclk));
	jdff dff_B_OKspzJNu7_0(.din(w_dff_B_v6JDwg0L9_0),.dout(w_dff_B_OKspzJNu7_0),.clk(gclk));
	jdff dff_B_APgepRj83_0(.din(w_dff_B_OKspzJNu7_0),.dout(w_dff_B_APgepRj83_0),.clk(gclk));
	jdff dff_B_NgUwY59h6_0(.din(w_dff_B_APgepRj83_0),.dout(w_dff_B_NgUwY59h6_0),.clk(gclk));
	jdff dff_B_bdxp7AcU3_0(.din(w_dff_B_NgUwY59h6_0),.dout(w_dff_B_bdxp7AcU3_0),.clk(gclk));
	jdff dff_B_fis0PEsW9_0(.din(n1284),.dout(w_dff_B_fis0PEsW9_0),.clk(gclk));
	jdff dff_A_y1kofuVU5_0(.dout(w_G137_6[0]),.din(w_dff_A_y1kofuVU5_0),.clk(gclk));
	jdff dff_A_bZhs7fic4_0(.dout(w_dff_A_y1kofuVU5_0),.din(w_dff_A_bZhs7fic4_0),.clk(gclk));
	jdff dff_A_H5oXzNSF8_0(.dout(w_dff_A_bZhs7fic4_0),.din(w_dff_A_H5oXzNSF8_0),.clk(gclk));
	jdff dff_A_H3FSjW8n1_0(.dout(w_dff_A_H5oXzNSF8_0),.din(w_dff_A_H3FSjW8n1_0),.clk(gclk));
	jdff dff_A_ZlmiawB56_0(.dout(w_dff_A_H3FSjW8n1_0),.din(w_dff_A_ZlmiawB56_0),.clk(gclk));
	jdff dff_A_qp4LGAap9_1(.dout(w_G137_6[1]),.din(w_dff_A_qp4LGAap9_1),.clk(gclk));
	jdff dff_B_agRsUJDf4_0(.din(n1293),.dout(w_dff_B_agRsUJDf4_0),.clk(gclk));
	jdff dff_B_ZKwsOfHf5_0(.din(w_dff_B_agRsUJDf4_0),.dout(w_dff_B_ZKwsOfHf5_0),.clk(gclk));
	jdff dff_B_V3uCsFml0_0(.din(w_dff_B_ZKwsOfHf5_0),.dout(w_dff_B_V3uCsFml0_0),.clk(gclk));
	jdff dff_B_SQHPePvO3_0(.din(w_dff_B_V3uCsFml0_0),.dout(w_dff_B_SQHPePvO3_0),.clk(gclk));
	jdff dff_B_TDWBnvTb7_0(.din(w_dff_B_SQHPePvO3_0),.dout(w_dff_B_TDWBnvTb7_0),.clk(gclk));
	jdff dff_B_xr8B8iLi1_0(.din(w_dff_B_TDWBnvTb7_0),.dout(w_dff_B_xr8B8iLi1_0),.clk(gclk));
	jdff dff_B_12MprNB32_0(.din(w_dff_B_xr8B8iLi1_0),.dout(w_dff_B_12MprNB32_0),.clk(gclk));
	jdff dff_B_5aEKSf3m8_0(.din(w_dff_B_12MprNB32_0),.dout(w_dff_B_5aEKSf3m8_0),.clk(gclk));
	jdff dff_B_RkBc9UVD7_0(.din(w_dff_B_5aEKSf3m8_0),.dout(w_dff_B_RkBc9UVD7_0),.clk(gclk));
	jdff dff_B_3hqkoWtI1_0(.din(w_dff_B_RkBc9UVD7_0),.dout(w_dff_B_3hqkoWtI1_0),.clk(gclk));
	jdff dff_B_sIJUYtiF0_0(.din(w_dff_B_3hqkoWtI1_0),.dout(w_dff_B_sIJUYtiF0_0),.clk(gclk));
	jdff dff_B_6nGtx7Bc5_0(.din(w_dff_B_sIJUYtiF0_0),.dout(w_dff_B_6nGtx7Bc5_0),.clk(gclk));
	jdff dff_B_7UyEt8Gt1_0(.din(w_dff_B_6nGtx7Bc5_0),.dout(w_dff_B_7UyEt8Gt1_0),.clk(gclk));
	jdff dff_B_wjNWKAFj7_0(.din(w_dff_B_7UyEt8Gt1_0),.dout(w_dff_B_wjNWKAFj7_0),.clk(gclk));
	jdff dff_B_EBRwlS4T6_0(.din(w_dff_B_wjNWKAFj7_0),.dout(w_dff_B_EBRwlS4T6_0),.clk(gclk));
	jdff dff_B_V85onpWG4_0(.din(w_dff_B_EBRwlS4T6_0),.dout(w_dff_B_V85onpWG4_0),.clk(gclk));
	jdff dff_B_294IO92r3_0(.din(n1292),.dout(w_dff_B_294IO92r3_0),.clk(gclk));
	jdff dff_B_d0YDtxRG3_0(.din(n1301),.dout(w_dff_B_d0YDtxRG3_0),.clk(gclk));
	jdff dff_B_LAXbZkme6_0(.din(w_dff_B_d0YDtxRG3_0),.dout(w_dff_B_LAXbZkme6_0),.clk(gclk));
	jdff dff_B_wMMrjdzF3_0(.din(w_dff_B_LAXbZkme6_0),.dout(w_dff_B_wMMrjdzF3_0),.clk(gclk));
	jdff dff_B_Tv3AhgpP7_0(.din(w_dff_B_wMMrjdzF3_0),.dout(w_dff_B_Tv3AhgpP7_0),.clk(gclk));
	jdff dff_B_cbFc7pic9_0(.din(w_dff_B_Tv3AhgpP7_0),.dout(w_dff_B_cbFc7pic9_0),.clk(gclk));
	jdff dff_B_8GxulXDB4_0(.din(w_dff_B_cbFc7pic9_0),.dout(w_dff_B_8GxulXDB4_0),.clk(gclk));
	jdff dff_B_dM2C0V3V7_0(.din(w_dff_B_8GxulXDB4_0),.dout(w_dff_B_dM2C0V3V7_0),.clk(gclk));
	jdff dff_B_g5vUnsM18_0(.din(w_dff_B_dM2C0V3V7_0),.dout(w_dff_B_g5vUnsM18_0),.clk(gclk));
	jdff dff_B_KOhDaaUz2_0(.din(w_dff_B_g5vUnsM18_0),.dout(w_dff_B_KOhDaaUz2_0),.clk(gclk));
	jdff dff_B_O3LfvDXL3_0(.din(w_dff_B_KOhDaaUz2_0),.dout(w_dff_B_O3LfvDXL3_0),.clk(gclk));
	jdff dff_B_xyw0L8UL6_0(.din(w_dff_B_O3LfvDXL3_0),.dout(w_dff_B_xyw0L8UL6_0),.clk(gclk));
	jdff dff_B_AAfTTh1A4_0(.din(w_dff_B_xyw0L8UL6_0),.dout(w_dff_B_AAfTTh1A4_0),.clk(gclk));
	jdff dff_B_ViAWt65H6_0(.din(w_dff_B_AAfTTh1A4_0),.dout(w_dff_B_ViAWt65H6_0),.clk(gclk));
	jdff dff_B_MkvfGRyR6_0(.din(w_dff_B_ViAWt65H6_0),.dout(w_dff_B_MkvfGRyR6_0),.clk(gclk));
	jdff dff_B_cssxxx1u9_0(.din(w_dff_B_MkvfGRyR6_0),.dout(w_dff_B_cssxxx1u9_0),.clk(gclk));
	jdff dff_B_C1YjVtUI7_0(.din(w_dff_B_cssxxx1u9_0),.dout(w_dff_B_C1YjVtUI7_0),.clk(gclk));
	jdff dff_B_FfSLbWuY1_0(.din(n1300),.dout(w_dff_B_FfSLbWuY1_0),.clk(gclk));
	jdff dff_A_7OW5y9l72_0(.dout(w_n988_2[0]),.din(w_dff_A_7OW5y9l72_0),.clk(gclk));
	jdff dff_A_l4jMXvw94_1(.dout(w_n988_2[1]),.din(w_dff_A_l4jMXvw94_1),.clk(gclk));
	jdff dff_A_PHBE6jlE2_0(.dout(w_n985_2[0]),.din(w_dff_A_PHBE6jlE2_0),.clk(gclk));
	jdff dff_A_o45GCSCM4_1(.dout(w_n985_2[1]),.din(w_dff_A_o45GCSCM4_1),.clk(gclk));
	jdff dff_B_gVdEtFX19_0(.din(n1309),.dout(w_dff_B_gVdEtFX19_0),.clk(gclk));
	jdff dff_B_Ba0686lj8_0(.din(w_dff_B_gVdEtFX19_0),.dout(w_dff_B_Ba0686lj8_0),.clk(gclk));
	jdff dff_B_qsfq8MbL0_0(.din(w_dff_B_Ba0686lj8_0),.dout(w_dff_B_qsfq8MbL0_0),.clk(gclk));
	jdff dff_B_KfOZ8Leu1_0(.din(w_dff_B_qsfq8MbL0_0),.dout(w_dff_B_KfOZ8Leu1_0),.clk(gclk));
	jdff dff_B_vj1MW3nq9_0(.din(w_dff_B_KfOZ8Leu1_0),.dout(w_dff_B_vj1MW3nq9_0),.clk(gclk));
	jdff dff_B_uS61SSR74_0(.din(w_dff_B_vj1MW3nq9_0),.dout(w_dff_B_uS61SSR74_0),.clk(gclk));
	jdff dff_B_C9ky7vOl1_0(.din(w_dff_B_uS61SSR74_0),.dout(w_dff_B_C9ky7vOl1_0),.clk(gclk));
	jdff dff_B_R2CeI2Jc3_0(.din(w_dff_B_C9ky7vOl1_0),.dout(w_dff_B_R2CeI2Jc3_0),.clk(gclk));
	jdff dff_B_kMat4lox3_0(.din(w_dff_B_R2CeI2Jc3_0),.dout(w_dff_B_kMat4lox3_0),.clk(gclk));
	jdff dff_B_Rdg9HmST9_0(.din(w_dff_B_kMat4lox3_0),.dout(w_dff_B_Rdg9HmST9_0),.clk(gclk));
	jdff dff_B_JhlFtZgN5_0(.din(w_dff_B_Rdg9HmST9_0),.dout(w_dff_B_JhlFtZgN5_0),.clk(gclk));
	jdff dff_B_3CmVi0QK0_0(.din(w_dff_B_JhlFtZgN5_0),.dout(w_dff_B_3CmVi0QK0_0),.clk(gclk));
	jdff dff_B_yBsCen7m0_0(.din(w_dff_B_3CmVi0QK0_0),.dout(w_dff_B_yBsCen7m0_0),.clk(gclk));
	jdff dff_B_V5ZrAPuN6_0(.din(w_dff_B_yBsCen7m0_0),.dout(w_dff_B_V5ZrAPuN6_0),.clk(gclk));
	jdff dff_B_xyVYWRYK9_0(.din(w_dff_B_V5ZrAPuN6_0),.dout(w_dff_B_xyVYWRYK9_0),.clk(gclk));
	jdff dff_B_s55vGzNJ3_0(.din(w_dff_B_xyVYWRYK9_0),.dout(w_dff_B_s55vGzNJ3_0),.clk(gclk));
	jdff dff_B_UhZT5YK20_0(.din(w_dff_B_s55vGzNJ3_0),.dout(w_dff_B_UhZT5YK20_0),.clk(gclk));
	jdff dff_B_KImXdIga2_0(.din(n1308),.dout(w_dff_B_KImXdIga2_0),.clk(gclk));
	jdff dff_A_RQQIh7vn0_0(.dout(w_G137_5[0]),.din(w_dff_A_RQQIh7vn0_0),.clk(gclk));
	jdff dff_B_ZmFCOJy13_0(.din(n1317),.dout(w_dff_B_ZmFCOJy13_0),.clk(gclk));
	jdff dff_B_JbI7LX1H9_0(.din(w_dff_B_ZmFCOJy13_0),.dout(w_dff_B_JbI7LX1H9_0),.clk(gclk));
	jdff dff_B_LMESYq2w5_0(.din(w_dff_B_JbI7LX1H9_0),.dout(w_dff_B_LMESYq2w5_0),.clk(gclk));
	jdff dff_B_8hAu5rcr9_0(.din(w_dff_B_LMESYq2w5_0),.dout(w_dff_B_8hAu5rcr9_0),.clk(gclk));
	jdff dff_B_a35Fo7iV8_0(.din(w_dff_B_8hAu5rcr9_0),.dout(w_dff_B_a35Fo7iV8_0),.clk(gclk));
	jdff dff_B_t3yeZgE34_0(.din(w_dff_B_a35Fo7iV8_0),.dout(w_dff_B_t3yeZgE34_0),.clk(gclk));
	jdff dff_B_4xMKYaLx1_0(.din(w_dff_B_t3yeZgE34_0),.dout(w_dff_B_4xMKYaLx1_0),.clk(gclk));
	jdff dff_B_7PEwpT1r2_0(.din(w_dff_B_4xMKYaLx1_0),.dout(w_dff_B_7PEwpT1r2_0),.clk(gclk));
	jdff dff_B_zu2voKMB9_0(.din(w_dff_B_7PEwpT1r2_0),.dout(w_dff_B_zu2voKMB9_0),.clk(gclk));
	jdff dff_B_QUWFna4i9_0(.din(w_dff_B_zu2voKMB9_0),.dout(w_dff_B_QUWFna4i9_0),.clk(gclk));
	jdff dff_B_5Bds0IZW2_0(.din(w_dff_B_QUWFna4i9_0),.dout(w_dff_B_5Bds0IZW2_0),.clk(gclk));
	jdff dff_B_CIdUXag39_0(.din(w_dff_B_5Bds0IZW2_0),.dout(w_dff_B_CIdUXag39_0),.clk(gclk));
	jdff dff_B_vmB6lXpv2_0(.din(w_dff_B_CIdUXag39_0),.dout(w_dff_B_vmB6lXpv2_0),.clk(gclk));
	jdff dff_B_SWDiZyBP0_0(.din(w_dff_B_vmB6lXpv2_0),.dout(w_dff_B_SWDiZyBP0_0),.clk(gclk));
	jdff dff_B_ccTWhB2x9_0(.din(w_dff_B_SWDiZyBP0_0),.dout(w_dff_B_ccTWhB2x9_0),.clk(gclk));
	jdff dff_B_OKMz4WVo9_0(.din(n1316),.dout(w_dff_B_OKMz4WVo9_0),.clk(gclk));
	jdff dff_B_SGUhAMb97_2(.din(G173),.dout(w_dff_B_SGUhAMb97_2),.clk(gclk));
	jdff dff_B_IFxkz3Y08_2(.din(G203),.dout(w_dff_B_IFxkz3Y08_2),.clk(gclk));
	jdff dff_B_mLxJD7f59_2(.din(w_dff_B_IFxkz3Y08_2),.dout(w_dff_B_mLxJD7f59_2),.clk(gclk));
	jdff dff_B_I9S9Xa0x6_0(.din(n1182),.dout(w_dff_B_I9S9Xa0x6_0),.clk(gclk));
	jdff dff_B_TEtLmidp4_0(.din(w_dff_B_I9S9Xa0x6_0),.dout(w_dff_B_TEtLmidp4_0),.clk(gclk));
	jdff dff_B_96xzDBIs6_0(.din(w_dff_B_TEtLmidp4_0),.dout(w_dff_B_96xzDBIs6_0),.clk(gclk));
	jdff dff_B_LHpPA1Wf7_0(.din(w_dff_B_96xzDBIs6_0),.dout(w_dff_B_LHpPA1Wf7_0),.clk(gclk));
	jdff dff_B_cFYJGVhW7_0(.din(w_dff_B_LHpPA1Wf7_0),.dout(w_dff_B_cFYJGVhW7_0),.clk(gclk));
	jdff dff_B_RMXQNnOq9_0(.din(w_dff_B_cFYJGVhW7_0),.dout(w_dff_B_RMXQNnOq9_0),.clk(gclk));
	jdff dff_B_L4qQWu689_0(.din(w_dff_B_RMXQNnOq9_0),.dout(w_dff_B_L4qQWu689_0),.clk(gclk));
	jdff dff_B_kmG4DrdP9_0(.din(w_dff_B_L4qQWu689_0),.dout(w_dff_B_kmG4DrdP9_0),.clk(gclk));
	jdff dff_B_AQUBKamq2_0(.din(w_dff_B_kmG4DrdP9_0),.dout(w_dff_B_AQUBKamq2_0),.clk(gclk));
	jdff dff_B_E1ByTHYL4_0(.din(n1181),.dout(w_dff_B_E1ByTHYL4_0),.clk(gclk));
	jdff dff_B_62huH6Nq1_0(.din(w_dff_B_E1ByTHYL4_0),.dout(w_dff_B_62huH6Nq1_0),.clk(gclk));
	jdff dff_B_3epKLyCT9_1(.din(G112),.dout(w_dff_B_3epKLyCT9_1),.clk(gclk));
	jdff dff_B_tYfQVzEI9_1(.din(w_dff_B_3epKLyCT9_1),.dout(w_dff_B_tYfQVzEI9_1),.clk(gclk));
	jdff dff_B_17aiqjGc4_0(.din(n1218),.dout(w_dff_B_17aiqjGc4_0),.clk(gclk));
	jdff dff_B_dSejLMxx2_0(.din(w_dff_B_17aiqjGc4_0),.dout(w_dff_B_dSejLMxx2_0),.clk(gclk));
	jdff dff_B_nek2bSjm6_0(.din(w_dff_B_dSejLMxx2_0),.dout(w_dff_B_nek2bSjm6_0),.clk(gclk));
	jdff dff_B_IX8EgRQH2_0(.din(w_dff_B_nek2bSjm6_0),.dout(w_dff_B_IX8EgRQH2_0),.clk(gclk));
	jdff dff_B_xbHkbq0I8_0(.din(w_dff_B_IX8EgRQH2_0),.dout(w_dff_B_xbHkbq0I8_0),.clk(gclk));
	jdff dff_B_UnPCY6Db0_0(.din(w_dff_B_xbHkbq0I8_0),.dout(w_dff_B_UnPCY6Db0_0),.clk(gclk));
	jdff dff_B_dihwUXjS5_0(.din(w_dff_B_UnPCY6Db0_0),.dout(w_dff_B_dihwUXjS5_0),.clk(gclk));
	jdff dff_B_gCnKLI5i2_0(.din(w_dff_B_dihwUXjS5_0),.dout(w_dff_B_gCnKLI5i2_0),.clk(gclk));
	jdff dff_B_9CBb133i7_0(.din(w_dff_B_gCnKLI5i2_0),.dout(w_dff_B_9CBb133i7_0),.clk(gclk));
	jdff dff_B_jGhB8Mmf3_0(.din(w_dff_B_9CBb133i7_0),.dout(w_dff_B_jGhB8Mmf3_0),.clk(gclk));
	jdff dff_B_p23c7erm3_0(.din(n1217),.dout(w_dff_B_p23c7erm3_0),.clk(gclk));
	jdff dff_B_kWzdq82a2_0(.din(w_dff_B_p23c7erm3_0),.dout(w_dff_B_kWzdq82a2_0),.clk(gclk));
	jdff dff_B_0TVAYJPD2_1(.din(G113),.dout(w_dff_B_0TVAYJPD2_1),.clk(gclk));
	jdff dff_B_AKDvo7Ba7_1(.din(w_dff_B_0TVAYJPD2_1),.dout(w_dff_B_AKDvo7Ba7_1),.clk(gclk));
	jdff dff_B_2wflkQor3_0(.din(n539),.dout(w_dff_B_2wflkQor3_0),.clk(gclk));
	jdff dff_B_YdcdSCpG9_1(.din(n531),.dout(w_dff_B_YdcdSCpG9_1),.clk(gclk));
	jdff dff_B_09Q8taF07_0(.din(n1325),.dout(w_dff_B_09Q8taF07_0),.clk(gclk));
	jdff dff_B_zEuw58Vs5_0(.din(w_dff_B_09Q8taF07_0),.dout(w_dff_B_zEuw58Vs5_0),.clk(gclk));
	jdff dff_B_qtFTJ7YN5_0(.din(w_dff_B_zEuw58Vs5_0),.dout(w_dff_B_qtFTJ7YN5_0),.clk(gclk));
	jdff dff_B_0rmgxtLS1_0(.din(w_dff_B_qtFTJ7YN5_0),.dout(w_dff_B_0rmgxtLS1_0),.clk(gclk));
	jdff dff_B_dYrKAl9E6_0(.din(w_dff_B_0rmgxtLS1_0),.dout(w_dff_B_dYrKAl9E6_0),.clk(gclk));
	jdff dff_B_EJQTvFzO7_0(.din(w_dff_B_dYrKAl9E6_0),.dout(w_dff_B_EJQTvFzO7_0),.clk(gclk));
	jdff dff_B_BiTMPZqi6_0(.din(w_dff_B_EJQTvFzO7_0),.dout(w_dff_B_BiTMPZqi6_0),.clk(gclk));
	jdff dff_B_dqkJ1ncm3_0(.din(w_dff_B_BiTMPZqi6_0),.dout(w_dff_B_dqkJ1ncm3_0),.clk(gclk));
	jdff dff_B_fmMG05vF3_0(.din(w_dff_B_dqkJ1ncm3_0),.dout(w_dff_B_fmMG05vF3_0),.clk(gclk));
	jdff dff_B_AtuYmRCA6_0(.din(w_dff_B_fmMG05vF3_0),.dout(w_dff_B_AtuYmRCA6_0),.clk(gclk));
	jdff dff_B_IFHSWs6i4_0(.din(w_dff_B_AtuYmRCA6_0),.dout(w_dff_B_IFHSWs6i4_0),.clk(gclk));
	jdff dff_B_d8G8CC2Z5_0(.din(w_dff_B_IFHSWs6i4_0),.dout(w_dff_B_d8G8CC2Z5_0),.clk(gclk));
	jdff dff_B_aj8h4fjM8_0(.din(w_dff_B_d8G8CC2Z5_0),.dout(w_dff_B_aj8h4fjM8_0),.clk(gclk));
	jdff dff_B_GURgKlrr4_0(.din(w_dff_B_aj8h4fjM8_0),.dout(w_dff_B_GURgKlrr4_0),.clk(gclk));
	jdff dff_B_qCbrYods6_0(.din(w_dff_B_GURgKlrr4_0),.dout(w_dff_B_qCbrYods6_0),.clk(gclk));
	jdff dff_B_lXYnlb5b3_0(.din(w_dff_B_qCbrYods6_0),.dout(w_dff_B_lXYnlb5b3_0),.clk(gclk));
	jdff dff_B_SAWpM6fQ5_0(.din(n1324),.dout(w_dff_B_SAWpM6fQ5_0),.clk(gclk));
	jdff dff_B_MAJmmH5t1_2(.din(G167),.dout(w_dff_B_MAJmmH5t1_2),.clk(gclk));
	jdff dff_B_50RCKjQP1_2(.din(G197),.dout(w_dff_B_50RCKjQP1_2),.clk(gclk));
	jdff dff_B_cFW4n59S5_2(.din(w_dff_B_50RCKjQP1_2),.dout(w_dff_B_cFW4n59S5_2),.clk(gclk));
	jdff dff_B_LIqQJyqB7_0(.din(n1175),.dout(w_dff_B_LIqQJyqB7_0),.clk(gclk));
	jdff dff_B_154GA88v8_0(.din(w_dff_B_LIqQJyqB7_0),.dout(w_dff_B_154GA88v8_0),.clk(gclk));
	jdff dff_B_scoLKQWQ0_0(.din(w_dff_B_154GA88v8_0),.dout(w_dff_B_scoLKQWQ0_0),.clk(gclk));
	jdff dff_B_H5TTfpr02_0(.din(w_dff_B_scoLKQWQ0_0),.dout(w_dff_B_H5TTfpr02_0),.clk(gclk));
	jdff dff_B_WVwjElLV1_0(.din(w_dff_B_H5TTfpr02_0),.dout(w_dff_B_WVwjElLV1_0),.clk(gclk));
	jdff dff_B_r8tieEPh9_0(.din(w_dff_B_WVwjElLV1_0),.dout(w_dff_B_r8tieEPh9_0),.clk(gclk));
	jdff dff_B_xGpnWdoj3_0(.din(w_dff_B_r8tieEPh9_0),.dout(w_dff_B_xGpnWdoj3_0),.clk(gclk));
	jdff dff_B_fKnP5ZTG4_0(.din(w_dff_B_xGpnWdoj3_0),.dout(w_dff_B_fKnP5ZTG4_0),.clk(gclk));
	jdff dff_B_zpKo9Ccc5_0(.din(w_dff_B_fKnP5ZTG4_0),.dout(w_dff_B_zpKo9Ccc5_0),.clk(gclk));
	jdff dff_B_vJHcfLve3_0(.din(w_dff_B_zpKo9Ccc5_0),.dout(w_dff_B_vJHcfLve3_0),.clk(gclk));
	jdff dff_B_3J5EAi6i6_0(.din(n1174),.dout(w_dff_B_3J5EAi6i6_0),.clk(gclk));
	jdff dff_B_1QghGSTZ5_0(.din(w_dff_B_3J5EAi6i6_0),.dout(w_dff_B_1QghGSTZ5_0),.clk(gclk));
	jdff dff_B_odjM5rvn3_1(.din(G116),.dout(w_dff_B_odjM5rvn3_1),.clk(gclk));
	jdff dff_B_h2p3nyxB3_1(.din(w_dff_B_odjM5rvn3_1),.dout(w_dff_B_h2p3nyxB3_1),.clk(gclk));
	jdff dff_A_sUW6gcWQ9_1(.dout(w_n971_0[1]),.din(w_dff_A_sUW6gcWQ9_1),.clk(gclk));
	jdff dff_B_quMq9nbg5_1(.din(n967),.dout(w_dff_B_quMq9nbg5_1),.clk(gclk));
	jdff dff_B_sQCErxne2_1(.din(w_dff_B_quMq9nbg5_1),.dout(w_dff_B_sQCErxne2_1),.clk(gclk));
	jdff dff_B_4EsNKvRA1_1(.din(w_dff_B_sQCErxne2_1),.dout(w_dff_B_4EsNKvRA1_1),.clk(gclk));
	jdff dff_B_l8XGactB8_1(.din(w_dff_B_4EsNKvRA1_1),.dout(w_dff_B_l8XGactB8_1),.clk(gclk));
	jdff dff_B_xlzh8Ftl9_1(.din(w_dff_B_l8XGactB8_1),.dout(w_dff_B_xlzh8Ftl9_1),.clk(gclk));
	jdff dff_B_c0G0nXkd0_1(.din(w_dff_B_xlzh8Ftl9_1),.dout(w_dff_B_c0G0nXkd0_1),.clk(gclk));
	jdff dff_B_kZeNUo0G9_1(.din(w_dff_B_c0G0nXkd0_1),.dout(w_dff_B_kZeNUo0G9_1),.clk(gclk));
	jdff dff_B_3nxzTJoj7_1(.din(w_dff_B_kZeNUo0G9_1),.dout(w_dff_B_3nxzTJoj7_1),.clk(gclk));
	jdff dff_B_kOVmyXKi0_1(.din(w_dff_B_3nxzTJoj7_1),.dout(w_dff_B_kOVmyXKi0_1),.clk(gclk));
	jdff dff_B_udGqIPxm7_1(.din(w_dff_B_kOVmyXKi0_1),.dout(w_dff_B_udGqIPxm7_1),.clk(gclk));
	jdff dff_B_IMe2uchO1_0(.din(n1211),.dout(w_dff_B_IMe2uchO1_0),.clk(gclk));
	jdff dff_B_ZReIIt4W8_0(.din(w_dff_B_IMe2uchO1_0),.dout(w_dff_B_ZReIIt4W8_0),.clk(gclk));
	jdff dff_B_gw0ZtexQ4_0(.din(w_dff_B_ZReIIt4W8_0),.dout(w_dff_B_gw0ZtexQ4_0),.clk(gclk));
	jdff dff_B_7sCawKEX8_0(.din(w_dff_B_gw0ZtexQ4_0),.dout(w_dff_B_7sCawKEX8_0),.clk(gclk));
	jdff dff_B_8Ui3d48h8_0(.din(w_dff_B_7sCawKEX8_0),.dout(w_dff_B_8Ui3d48h8_0),.clk(gclk));
	jdff dff_B_mSSl9zLJ1_0(.din(w_dff_B_8Ui3d48h8_0),.dout(w_dff_B_mSSl9zLJ1_0),.clk(gclk));
	jdff dff_B_sNTc23mc7_0(.din(w_dff_B_mSSl9zLJ1_0),.dout(w_dff_B_sNTc23mc7_0),.clk(gclk));
	jdff dff_B_9oJ52C180_0(.din(w_dff_B_sNTc23mc7_0),.dout(w_dff_B_9oJ52C180_0),.clk(gclk));
	jdff dff_B_MqaT0KJJ5_0(.din(w_dff_B_9oJ52C180_0),.dout(w_dff_B_MqaT0KJJ5_0),.clk(gclk));
	jdff dff_B_AQXaAoau3_0(.din(w_dff_B_MqaT0KJJ5_0),.dout(w_dff_B_AQXaAoau3_0),.clk(gclk));
	jdff dff_B_xAXaJ5Ik2_0(.din(w_dff_B_AQXaAoau3_0),.dout(w_dff_B_xAXaJ5Ik2_0),.clk(gclk));
	jdff dff_B_pxnY8ccd7_0(.din(n1210),.dout(w_dff_B_pxnY8ccd7_0),.clk(gclk));
	jdff dff_B_7PZywBut2_0(.din(w_dff_B_pxnY8ccd7_0),.dout(w_dff_B_7PZywBut2_0),.clk(gclk));
	jdff dff_B_Nj5vdTif5_1(.din(G53),.dout(w_dff_B_Nj5vdTif5_1),.clk(gclk));
	jdff dff_B_StV1voEx0_1(.din(w_dff_B_Nj5vdTif5_1),.dout(w_dff_B_StV1voEx0_1),.clk(gclk));
	jdff dff_B_gG2uUQz25_0(.din(n516),.dout(w_dff_B_gG2uUQz25_0),.clk(gclk));
	jdff dff_B_ETgeSkvN4_1(.din(n508),.dout(w_dff_B_ETgeSkvN4_1),.clk(gclk));
	jdff dff_B_ixPsF8PX5_1(.din(n949),.dout(w_dff_B_ixPsF8PX5_1),.clk(gclk));
	jdff dff_B_4qSErFbZ5_1(.din(w_dff_B_ixPsF8PX5_1),.dout(w_dff_B_4qSErFbZ5_1),.clk(gclk));
	jdff dff_B_55kHWLt07_1(.din(w_dff_B_4qSErFbZ5_1),.dout(w_dff_B_55kHWLt07_1),.clk(gclk));
	jdff dff_B_PdoLO2ui9_1(.din(w_dff_B_55kHWLt07_1),.dout(w_dff_B_PdoLO2ui9_1),.clk(gclk));
	jdff dff_B_Uo6Ck4sD7_1(.din(w_dff_B_PdoLO2ui9_1),.dout(w_dff_B_Uo6Ck4sD7_1),.clk(gclk));
	jdff dff_B_Us86aFVR4_1(.din(w_dff_B_Uo6Ck4sD7_1),.dout(w_dff_B_Us86aFVR4_1),.clk(gclk));
	jdff dff_B_mXczXv536_1(.din(w_dff_B_Us86aFVR4_1),.dout(w_dff_B_mXczXv536_1),.clk(gclk));
	jdff dff_B_sf9LzMDB0_1(.din(w_dff_B_mXczXv536_1),.dout(w_dff_B_sf9LzMDB0_1),.clk(gclk));
	jdff dff_B_c7gxiID30_1(.din(w_dff_B_sf9LzMDB0_1),.dout(w_dff_B_c7gxiID30_1),.clk(gclk));
	jdff dff_B_TffRr9w90_1(.din(w_dff_B_c7gxiID30_1),.dout(w_dff_B_TffRr9w90_1),.clk(gclk));
	jdff dff_B_3c94yB1b0_1(.din(n950),.dout(w_dff_B_3c94yB1b0_1),.clk(gclk));
	jdff dff_B_fpTMEgEi4_1(.din(w_dff_B_3c94yB1b0_1),.dout(w_dff_B_fpTMEgEi4_1),.clk(gclk));
	jdff dff_B_eeznKk6L0_1(.din(w_dff_B_fpTMEgEi4_1),.dout(w_dff_B_eeznKk6L0_1),.clk(gclk));
	jdff dff_B_ConUEDM16_1(.din(w_dff_B_eeznKk6L0_1),.dout(w_dff_B_ConUEDM16_1),.clk(gclk));
	jdff dff_B_qsOYPMWr4_1(.din(w_dff_B_ConUEDM16_1),.dout(w_dff_B_qsOYPMWr4_1),.clk(gclk));
	jdff dff_B_VbZ4XuZP0_1(.din(w_dff_B_qsOYPMWr4_1),.dout(w_dff_B_VbZ4XuZP0_1),.clk(gclk));
	jdff dff_B_P1WrViCA7_1(.din(w_dff_B_VbZ4XuZP0_1),.dout(w_dff_B_P1WrViCA7_1),.clk(gclk));
	jdff dff_B_iBWYpPYu7_1(.din(w_dff_B_P1WrViCA7_1),.dout(w_dff_B_iBWYpPYu7_1),.clk(gclk));
	jdff dff_B_e5HQDqVp5_1(.din(w_dff_B_iBWYpPYu7_1),.dout(w_dff_B_e5HQDqVp5_1),.clk(gclk));
	jdff dff_A_sAzoij892_1(.dout(w_n748_1[1]),.din(w_dff_A_sAzoij892_1),.clk(gclk));
	jdff dff_A_6FYOdVxK6_1(.dout(w_dff_A_sAzoij892_1),.din(w_dff_A_6FYOdVxK6_1),.clk(gclk));
	jdff dff_A_zNPmARhV5_1(.dout(w_dff_A_6FYOdVxK6_1),.din(w_dff_A_zNPmARhV5_1),.clk(gclk));
	jdff dff_A_77DusoA61_1(.dout(w_dff_A_zNPmARhV5_1),.din(w_dff_A_77DusoA61_1),.clk(gclk));
	jdff dff_A_aLhqdgZU3_1(.dout(w_dff_A_77DusoA61_1),.din(w_dff_A_aLhqdgZU3_1),.clk(gclk));
	jdff dff_A_Vgr5vevl1_1(.dout(w_dff_A_aLhqdgZU3_1),.din(w_dff_A_Vgr5vevl1_1),.clk(gclk));
	jdff dff_A_vb2M1OE24_1(.dout(w_dff_A_Vgr5vevl1_1),.din(w_dff_A_vb2M1OE24_1),.clk(gclk));
	jdff dff_A_Ck6oxcC35_1(.dout(w_dff_A_vb2M1OE24_1),.din(w_dff_A_Ck6oxcC35_1),.clk(gclk));
	jdff dff_A_RBGRznVJ7_1(.dout(w_dff_A_Ck6oxcC35_1),.din(w_dff_A_RBGRznVJ7_1),.clk(gclk));
	jdff dff_A_zeRLM1kf4_1(.dout(w_dff_A_RBGRznVJ7_1),.din(w_dff_A_zeRLM1kf4_1),.clk(gclk));
	jdff dff_A_BmECUsk12_1(.dout(w_dff_A_zeRLM1kf4_1),.din(w_dff_A_BmECUsk12_1),.clk(gclk));
	jdff dff_A_Gu5nNEwY7_1(.dout(w_dff_A_BmECUsk12_1),.din(w_dff_A_Gu5nNEwY7_1),.clk(gclk));
	jdff dff_A_FBNMLUe16_1(.dout(w_dff_A_Gu5nNEwY7_1),.din(w_dff_A_FBNMLUe16_1),.clk(gclk));
	jdff dff_A_nDfkBzeK5_2(.dout(w_n748_1[2]),.din(w_dff_A_nDfkBzeK5_2),.clk(gclk));
	jdff dff_A_9RebKp3i9_2(.dout(w_dff_A_nDfkBzeK5_2),.din(w_dff_A_9RebKp3i9_2),.clk(gclk));
	jdff dff_A_gNbujCMb7_2(.dout(w_dff_A_9RebKp3i9_2),.din(w_dff_A_gNbujCMb7_2),.clk(gclk));
	jdff dff_A_aLH5F6Tt6_2(.dout(w_dff_A_gNbujCMb7_2),.din(w_dff_A_aLH5F6Tt6_2),.clk(gclk));
	jdff dff_A_Pimr12Am7_2(.dout(w_dff_A_aLH5F6Tt6_2),.din(w_dff_A_Pimr12Am7_2),.clk(gclk));
	jdff dff_A_ElQe45RG5_2(.dout(w_dff_A_Pimr12Am7_2),.din(w_dff_A_ElQe45RG5_2),.clk(gclk));
	jdff dff_A_2s2YT0uI2_2(.dout(w_dff_A_ElQe45RG5_2),.din(w_dff_A_2s2YT0uI2_2),.clk(gclk));
	jdff dff_A_btSBnyTP2_2(.dout(w_dff_A_2s2YT0uI2_2),.din(w_dff_A_btSBnyTP2_2),.clk(gclk));
	jdff dff_A_BPkgQXW11_2(.dout(w_dff_A_btSBnyTP2_2),.din(w_dff_A_BPkgQXW11_2),.clk(gclk));
	jdff dff_A_SQAQH26V5_2(.dout(w_dff_A_BPkgQXW11_2),.din(w_dff_A_SQAQH26V5_2),.clk(gclk));
	jdff dff_A_iNS2XPFK1_2(.dout(w_dff_A_SQAQH26V5_2),.din(w_dff_A_iNS2XPFK1_2),.clk(gclk));
	jdff dff_A_L5frsO004_2(.dout(w_dff_A_iNS2XPFK1_2),.din(w_dff_A_L5frsO004_2),.clk(gclk));
	jdff dff_B_9pLJ2O540_0(.din(n1333),.dout(w_dff_B_9pLJ2O540_0),.clk(gclk));
	jdff dff_B_cPWzW0kk4_0(.din(w_dff_B_9pLJ2O540_0),.dout(w_dff_B_cPWzW0kk4_0),.clk(gclk));
	jdff dff_B_Xe9zhxh66_0(.din(w_dff_B_cPWzW0kk4_0),.dout(w_dff_B_Xe9zhxh66_0),.clk(gclk));
	jdff dff_B_7iguyQVm5_0(.din(w_dff_B_Xe9zhxh66_0),.dout(w_dff_B_7iguyQVm5_0),.clk(gclk));
	jdff dff_B_RNLWmLJJ1_0(.din(w_dff_B_7iguyQVm5_0),.dout(w_dff_B_RNLWmLJJ1_0),.clk(gclk));
	jdff dff_B_RHF8iTjG5_0(.din(w_dff_B_RNLWmLJJ1_0),.dout(w_dff_B_RHF8iTjG5_0),.clk(gclk));
	jdff dff_B_pQW52dv74_0(.din(w_dff_B_RHF8iTjG5_0),.dout(w_dff_B_pQW52dv74_0),.clk(gclk));
	jdff dff_B_7y1vDWQp2_0(.din(w_dff_B_pQW52dv74_0),.dout(w_dff_B_7y1vDWQp2_0),.clk(gclk));
	jdff dff_B_5vVcP5lv2_0(.din(w_dff_B_7y1vDWQp2_0),.dout(w_dff_B_5vVcP5lv2_0),.clk(gclk));
	jdff dff_B_Bm4FV72o3_0(.din(w_dff_B_5vVcP5lv2_0),.dout(w_dff_B_Bm4FV72o3_0),.clk(gclk));
	jdff dff_B_j0If32eX7_0(.din(w_dff_B_Bm4FV72o3_0),.dout(w_dff_B_j0If32eX7_0),.clk(gclk));
	jdff dff_B_CjZodt2l6_0(.din(w_dff_B_j0If32eX7_0),.dout(w_dff_B_CjZodt2l6_0),.clk(gclk));
	jdff dff_B_DLpxs9L61_0(.din(w_dff_B_CjZodt2l6_0),.dout(w_dff_B_DLpxs9L61_0),.clk(gclk));
	jdff dff_B_yqIm284c6_0(.din(w_dff_B_DLpxs9L61_0),.dout(w_dff_B_yqIm284c6_0),.clk(gclk));
	jdff dff_B_Bbjyg1EH7_0(.din(w_dff_B_yqIm284c6_0),.dout(w_dff_B_Bbjyg1EH7_0),.clk(gclk));
	jdff dff_B_RyyWYobz7_0(.din(w_dff_B_Bbjyg1EH7_0),.dout(w_dff_B_RyyWYobz7_0),.clk(gclk));
	jdff dff_B_powhZxEO6_0(.din(n1332),.dout(w_dff_B_powhZxEO6_0),.clk(gclk));
	jdff dff_B_TvkVAIn21_2(.din(G164),.dout(w_dff_B_TvkVAIn21_2),.clk(gclk));
	jdff dff_B_14vpiaKB5_2(.din(G194),.dout(w_dff_B_14vpiaKB5_2),.clk(gclk));
	jdff dff_B_7lMbWqIo5_2(.din(w_dff_B_14vpiaKB5_2),.dout(w_dff_B_7lMbWqIo5_2),.clk(gclk));
	jdff dff_B_B84uG7bX8_0(.din(n1169),.dout(w_dff_B_B84uG7bX8_0),.clk(gclk));
	jdff dff_B_QjU99fHA3_0(.din(w_dff_B_B84uG7bX8_0),.dout(w_dff_B_QjU99fHA3_0),.clk(gclk));
	jdff dff_B_ucHpOF5h4_0(.din(w_dff_B_QjU99fHA3_0),.dout(w_dff_B_ucHpOF5h4_0),.clk(gclk));
	jdff dff_B_Ym1Q9bcb1_0(.din(w_dff_B_ucHpOF5h4_0),.dout(w_dff_B_Ym1Q9bcb1_0),.clk(gclk));
	jdff dff_B_ncHijzMR4_0(.din(w_dff_B_Ym1Q9bcb1_0),.dout(w_dff_B_ncHijzMR4_0),.clk(gclk));
	jdff dff_B_y0ZkcAHI7_0(.din(w_dff_B_ncHijzMR4_0),.dout(w_dff_B_y0ZkcAHI7_0),.clk(gclk));
	jdff dff_B_pY4kvoBt2_0(.din(w_dff_B_y0ZkcAHI7_0),.dout(w_dff_B_pY4kvoBt2_0),.clk(gclk));
	jdff dff_B_TvlAC35e3_0(.din(w_dff_B_pY4kvoBt2_0),.dout(w_dff_B_TvlAC35e3_0),.clk(gclk));
	jdff dff_B_Mlmerch91_0(.din(w_dff_B_TvlAC35e3_0),.dout(w_dff_B_Mlmerch91_0),.clk(gclk));
	jdff dff_B_pehWNw4f6_0(.din(w_dff_B_Mlmerch91_0),.dout(w_dff_B_pehWNw4f6_0),.clk(gclk));
	jdff dff_B_KrP1yuHQ9_0(.din(w_dff_B_pehWNw4f6_0),.dout(w_dff_B_KrP1yuHQ9_0),.clk(gclk));
	jdff dff_B_marBBmw55_0(.din(n1167),.dout(w_dff_B_marBBmw55_0),.clk(gclk));
	jdff dff_B_HXk0kOAM5_1(.din(G121),.dout(w_dff_B_HXk0kOAM5_1),.clk(gclk));
	jdff dff_B_uKr8CYGs6_1(.din(w_dff_B_HXk0kOAM5_1),.dout(w_dff_B_uKr8CYGs6_1),.clk(gclk));
	jdff dff_A_aeevJOVS0_0(.dout(w_n748_2[0]),.din(w_dff_A_aeevJOVS0_0),.clk(gclk));
	jdff dff_A_vEyg9jp74_0(.dout(w_dff_A_aeevJOVS0_0),.din(w_dff_A_vEyg9jp74_0),.clk(gclk));
	jdff dff_A_X6QMuLAm1_0(.dout(w_dff_A_vEyg9jp74_0),.din(w_dff_A_X6QMuLAm1_0),.clk(gclk));
	jdff dff_A_q9i9WFuA3_0(.dout(w_dff_A_X6QMuLAm1_0),.din(w_dff_A_q9i9WFuA3_0),.clk(gclk));
	jdff dff_A_SBknElrP1_2(.dout(w_n748_2[2]),.din(w_dff_A_SBknElrP1_2),.clk(gclk));
	jdff dff_A_YlD1YxIp1_2(.dout(w_dff_A_SBknElrP1_2),.din(w_dff_A_YlD1YxIp1_2),.clk(gclk));
	jdff dff_A_H1qLvIgG7_1(.dout(w_n748_0[1]),.din(w_dff_A_H1qLvIgG7_1),.clk(gclk));
	jdff dff_A_xsOeO7oV5_1(.dout(w_dff_A_H1qLvIgG7_1),.din(w_dff_A_xsOeO7oV5_1),.clk(gclk));
	jdff dff_A_ylCN2lH88_1(.dout(w_dff_A_xsOeO7oV5_1),.din(w_dff_A_ylCN2lH88_1),.clk(gclk));
	jdff dff_A_8yOW4PUZ0_1(.dout(w_dff_A_ylCN2lH88_1),.din(w_dff_A_8yOW4PUZ0_1),.clk(gclk));
	jdff dff_A_y7CO8UH03_1(.dout(w_dff_A_8yOW4PUZ0_1),.din(w_dff_A_y7CO8UH03_1),.clk(gclk));
	jdff dff_A_qzHdiVqZ7_1(.dout(w_dff_A_y7CO8UH03_1),.din(w_dff_A_qzHdiVqZ7_1),.clk(gclk));
	jdff dff_A_EnI1yzei1_1(.dout(w_dff_A_qzHdiVqZ7_1),.din(w_dff_A_EnI1yzei1_1),.clk(gclk));
	jdff dff_A_UQoh7LGe2_1(.dout(w_dff_A_EnI1yzei1_1),.din(w_dff_A_UQoh7LGe2_1),.clk(gclk));
	jdff dff_A_wOf1Cfte0_2(.dout(w_n748_0[2]),.din(w_dff_A_wOf1Cfte0_2),.clk(gclk));
	jdff dff_A_N3h0DbEd0_2(.dout(w_dff_A_wOf1Cfte0_2),.din(w_dff_A_N3h0DbEd0_2),.clk(gclk));
	jdff dff_A_wRFxOKzz0_2(.dout(w_dff_A_N3h0DbEd0_2),.din(w_dff_A_wRFxOKzz0_2),.clk(gclk));
	jdff dff_A_a3B1miSq9_2(.dout(w_dff_A_wRFxOKzz0_2),.din(w_dff_A_a3B1miSq9_2),.clk(gclk));
	jdff dff_B_qXzrlhWH2_3(.din(n748),.dout(w_dff_B_qXzrlhWH2_3),.clk(gclk));
	jdff dff_A_qNY8BP3v7_0(.dout(w_n747_3[0]),.din(w_dff_A_qNY8BP3v7_0),.clk(gclk));
	jdff dff_A_UXajs5TU9_0(.dout(w_dff_A_qNY8BP3v7_0),.din(w_dff_A_UXajs5TU9_0),.clk(gclk));
	jdff dff_A_aPAD6atK6_0(.dout(w_dff_A_UXajs5TU9_0),.din(w_dff_A_aPAD6atK6_0),.clk(gclk));
	jdff dff_A_WBxupp7Q1_0(.dout(w_dff_A_aPAD6atK6_0),.din(w_dff_A_WBxupp7Q1_0),.clk(gclk));
	jdff dff_A_n4a7JNKr9_0(.dout(w_dff_A_WBxupp7Q1_0),.din(w_dff_A_n4a7JNKr9_0),.clk(gclk));
	jdff dff_A_sTj0VN4c4_0(.dout(w_dff_A_n4a7JNKr9_0),.din(w_dff_A_sTj0VN4c4_0),.clk(gclk));
	jdff dff_A_e0JYmab19_0(.dout(w_dff_A_sTj0VN4c4_0),.din(w_dff_A_e0JYmab19_0),.clk(gclk));
	jdff dff_A_wDe8DPcc0_0(.dout(w_dff_A_e0JYmab19_0),.din(w_dff_A_wDe8DPcc0_0),.clk(gclk));
	jdff dff_A_SqI2yV546_1(.dout(w_n747_3[1]),.din(w_dff_A_SqI2yV546_1),.clk(gclk));
	jdff dff_A_3Vi918I32_1(.dout(w_dff_A_SqI2yV546_1),.din(w_dff_A_3Vi918I32_1),.clk(gclk));
	jdff dff_A_gU6XlNYE1_1(.dout(w_dff_A_3Vi918I32_1),.din(w_dff_A_gU6XlNYE1_1),.clk(gclk));
	jdff dff_A_H5bf7n1u2_0(.dout(w_n1002_2[0]),.din(w_dff_A_H5bf7n1u2_0),.clk(gclk));
	jdff dff_A_ITNR949C7_1(.dout(w_n1002_2[1]),.din(w_dff_A_ITNR949C7_1),.clk(gclk));
	jdff dff_B_S9J7nqW47_0(.din(n1204),.dout(w_dff_B_S9J7nqW47_0),.clk(gclk));
	jdff dff_B_qSC0jK4B7_0(.din(w_dff_B_S9J7nqW47_0),.dout(w_dff_B_qSC0jK4B7_0),.clk(gclk));
	jdff dff_B_74MEXcp64_0(.din(w_dff_B_qSC0jK4B7_0),.dout(w_dff_B_74MEXcp64_0),.clk(gclk));
	jdff dff_B_XNwsMo0y7_0(.din(w_dff_B_74MEXcp64_0),.dout(w_dff_B_XNwsMo0y7_0),.clk(gclk));
	jdff dff_B_yNmVYCKB9_0(.din(w_dff_B_XNwsMo0y7_0),.dout(w_dff_B_yNmVYCKB9_0),.clk(gclk));
	jdff dff_B_9U6ylI2J2_0(.din(w_dff_B_yNmVYCKB9_0),.dout(w_dff_B_9U6ylI2J2_0),.clk(gclk));
	jdff dff_B_XdZik20e3_0(.din(w_dff_B_9U6ylI2J2_0),.dout(w_dff_B_XdZik20e3_0),.clk(gclk));
	jdff dff_B_vMziX8uU1_0(.din(w_dff_B_XdZik20e3_0),.dout(w_dff_B_vMziX8uU1_0),.clk(gclk));
	jdff dff_B_r7ZKzvHx2_0(.din(w_dff_B_vMziX8uU1_0),.dout(w_dff_B_r7ZKzvHx2_0),.clk(gclk));
	jdff dff_B_9DeFJJmY7_0(.din(w_dff_B_r7ZKzvHx2_0),.dout(w_dff_B_9DeFJJmY7_0),.clk(gclk));
	jdff dff_B_WPzhHrAb9_0(.din(w_dff_B_9DeFJJmY7_0),.dout(w_dff_B_WPzhHrAb9_0),.clk(gclk));
	jdff dff_B_PqJq7Mgt4_0(.din(n1202),.dout(w_dff_B_PqJq7Mgt4_0),.clk(gclk));
	jdff dff_B_XGAPpf743_0(.din(w_dff_B_PqJq7Mgt4_0),.dout(w_dff_B_XGAPpf743_0),.clk(gclk));
	jdff dff_B_Nm4EO94P3_1(.din(G114),.dout(w_dff_B_Nm4EO94P3_1),.clk(gclk));
	jdff dff_B_vNPPy6ed3_1(.din(w_dff_B_Nm4EO94P3_1),.dout(w_dff_B_vNPPy6ed3_1),.clk(gclk));
	jdff dff_B_jFICK1UL1_3(.din(n765),.dout(w_dff_B_jFICK1UL1_3),.clk(gclk));
	jdff dff_B_rUp8ULsw4_3(.din(w_dff_B_jFICK1UL1_3),.dout(w_dff_B_rUp8ULsw4_3),.clk(gclk));
	jdff dff_A_BsgYYTw75_1(.dout(w_n751_2[1]),.din(w_dff_A_BsgYYTw75_1),.clk(gclk));
	jdff dff_B_Bb8vETym4_0(.din(n550),.dout(w_dff_B_Bb8vETym4_0),.clk(gclk));
	jdff dff_B_GertBESm2_3(.din(G3548),.dout(w_dff_B_GertBESm2_3),.clk(gclk));
	jdff dff_B_SCzYglrG4_1(.din(n542),.dout(w_dff_B_SCzYglrG4_1),.clk(gclk));
	jdff dff_A_fYU173FL6_0(.dout(w_n999_2[0]),.din(w_dff_A_fYU173FL6_0),.clk(gclk));
	jdff dff_A_tjHVlKCN6_1(.dout(w_n999_2[1]),.din(w_dff_A_tjHVlKCN6_1),.clk(gclk));
	jdff dff_A_383ZEy6I1_0(.dout(w_G137_4[0]),.din(w_dff_A_383ZEy6I1_0),.clk(gclk));
	jdff dff_A_ju5dP4BX9_1(.dout(w_G137_4[1]),.din(w_dff_A_ju5dP4BX9_1),.clk(gclk));
	jdff dff_A_y0ZRGQTF0_0(.dout(w_G137_1[0]),.din(w_dff_A_y0ZRGQTF0_0),.clk(gclk));
	jdff dff_A_sKZThTtb6_0(.dout(w_dff_A_y0ZRGQTF0_0),.din(w_dff_A_sKZThTtb6_0),.clk(gclk));
	jdff dff_A_q4R3ZE6d8_0(.dout(w_dff_A_sKZThTtb6_0),.din(w_dff_A_q4R3ZE6d8_0),.clk(gclk));
	jdff dff_A_ZCPtQnaG6_0(.dout(w_dff_A_q4R3ZE6d8_0),.din(w_dff_A_ZCPtQnaG6_0),.clk(gclk));
	jdff dff_A_so03MYB81_0(.dout(w_dff_A_ZCPtQnaG6_0),.din(w_dff_A_so03MYB81_0),.clk(gclk));
	jdff dff_A_a9J6yTKK2_1(.dout(w_G137_1[1]),.din(w_dff_A_a9J6yTKK2_1),.clk(gclk));
	jdff dff_A_ZJQjY5Xt2_1(.dout(w_dff_A_a9J6yTKK2_1),.din(w_dff_A_ZJQjY5Xt2_1),.clk(gclk));
	jdff dff_A_9IoQ8PG53_1(.dout(w_dff_A_ZJQjY5Xt2_1),.din(w_dff_A_9IoQ8PG53_1),.clk(gclk));
	jdff dff_A_HjS9J4X52_1(.dout(w_dff_A_9IoQ8PG53_1),.din(w_dff_A_HjS9J4X52_1),.clk(gclk));
	jdff dff_A_Fl8KFQKn2_1(.dout(w_dff_A_HjS9J4X52_1),.din(w_dff_A_Fl8KFQKn2_1),.clk(gclk));
	jdff dff_A_2NRd1JdT9_1(.dout(w_dff_A_Fl8KFQKn2_1),.din(w_dff_A_2NRd1JdT9_1),.clk(gclk));
	jdff dff_B_n7cutjcq9_0(.din(n1341),.dout(w_dff_B_n7cutjcq9_0),.clk(gclk));
	jdff dff_B_yptsFa2p8_0(.din(w_dff_B_n7cutjcq9_0),.dout(w_dff_B_yptsFa2p8_0),.clk(gclk));
	jdff dff_B_JRsmjG7t2_0(.din(w_dff_B_yptsFa2p8_0),.dout(w_dff_B_JRsmjG7t2_0),.clk(gclk));
	jdff dff_B_dZSZV8M57_0(.din(w_dff_B_JRsmjG7t2_0),.dout(w_dff_B_dZSZV8M57_0),.clk(gclk));
	jdff dff_B_BSzS8LU70_0(.din(w_dff_B_dZSZV8M57_0),.dout(w_dff_B_BSzS8LU70_0),.clk(gclk));
	jdff dff_B_JVHhIBho1_0(.din(w_dff_B_BSzS8LU70_0),.dout(w_dff_B_JVHhIBho1_0),.clk(gclk));
	jdff dff_B_plbfaqeX3_0(.din(w_dff_B_JVHhIBho1_0),.dout(w_dff_B_plbfaqeX3_0),.clk(gclk));
	jdff dff_B_7eWOYkPS2_0(.din(w_dff_B_plbfaqeX3_0),.dout(w_dff_B_7eWOYkPS2_0),.clk(gclk));
	jdff dff_B_gKVHduvz1_0(.din(w_dff_B_7eWOYkPS2_0),.dout(w_dff_B_gKVHduvz1_0),.clk(gclk));
	jdff dff_B_JV9dXuVZ5_0(.din(w_dff_B_gKVHduvz1_0),.dout(w_dff_B_JV9dXuVZ5_0),.clk(gclk));
	jdff dff_B_jeGq64yM1_0(.din(w_dff_B_JV9dXuVZ5_0),.dout(w_dff_B_jeGq64yM1_0),.clk(gclk));
	jdff dff_B_9pGaziJu7_0(.din(w_dff_B_jeGq64yM1_0),.dout(w_dff_B_9pGaziJu7_0),.clk(gclk));
	jdff dff_B_aV5fYulz2_0(.din(w_dff_B_9pGaziJu7_0),.dout(w_dff_B_aV5fYulz2_0),.clk(gclk));
	jdff dff_B_sLKrHYsW7_0(.din(w_dff_B_aV5fYulz2_0),.dout(w_dff_B_sLKrHYsW7_0),.clk(gclk));
	jdff dff_B_quMSMqcC0_0(.din(w_dff_B_sLKrHYsW7_0),.dout(w_dff_B_quMSMqcC0_0),.clk(gclk));
	jdff dff_B_ZUaMsc4b2_0(.din(w_dff_B_quMSMqcC0_0),.dout(w_dff_B_ZUaMsc4b2_0),.clk(gclk));
	jdff dff_B_AM3vBMxa2_0(.din(w_dff_B_ZUaMsc4b2_0),.dout(w_dff_B_AM3vBMxa2_0),.clk(gclk));
	jdff dff_B_nXPPc2nM8_0(.din(n1340),.dout(w_dff_B_nXPPc2nM8_0),.clk(gclk));
	jdff dff_B_wnoB62px8_2(.din(G161),.dout(w_dff_B_wnoB62px8_2),.clk(gclk));
	jdff dff_B_tpfWh4pm0_2(.din(G191),.dout(w_dff_B_tpfWh4pm0_2),.clk(gclk));
	jdff dff_B_YXrldbBk9_2(.din(w_dff_B_tpfWh4pm0_2),.dout(w_dff_B_YXrldbBk9_2),.clk(gclk));
	jdff dff_B_7FRchA6w4_0(.din(n1162),.dout(w_dff_B_7FRchA6w4_0),.clk(gclk));
	jdff dff_B_4RhB5ZPW2_0(.din(w_dff_B_7FRchA6w4_0),.dout(w_dff_B_4RhB5ZPW2_0),.clk(gclk));
	jdff dff_B_7D0ylB5Q9_0(.din(w_dff_B_4RhB5ZPW2_0),.dout(w_dff_B_7D0ylB5Q9_0),.clk(gclk));
	jdff dff_B_rEAdzYBT9_0(.din(w_dff_B_7D0ylB5Q9_0),.dout(w_dff_B_rEAdzYBT9_0),.clk(gclk));
	jdff dff_B_AhbaE4kP1_0(.din(w_dff_B_rEAdzYBT9_0),.dout(w_dff_B_AhbaE4kP1_0),.clk(gclk));
	jdff dff_B_u1HQjpXg7_0(.din(w_dff_B_AhbaE4kP1_0),.dout(w_dff_B_u1HQjpXg7_0),.clk(gclk));
	jdff dff_B_bmMGZWz43_0(.din(w_dff_B_u1HQjpXg7_0),.dout(w_dff_B_bmMGZWz43_0),.clk(gclk));
	jdff dff_B_IQ4cwdyf5_0(.din(w_dff_B_bmMGZWz43_0),.dout(w_dff_B_IQ4cwdyf5_0),.clk(gclk));
	jdff dff_B_3Of4yyyn8_0(.din(w_dff_B_IQ4cwdyf5_0),.dout(w_dff_B_3Of4yyyn8_0),.clk(gclk));
	jdff dff_B_ZRG9BTvk1_0(.din(w_dff_B_3Of4yyyn8_0),.dout(w_dff_B_ZRG9BTvk1_0),.clk(gclk));
	jdff dff_B_WMfun7bd3_0(.din(w_dff_B_ZRG9BTvk1_0),.dout(w_dff_B_WMfun7bd3_0),.clk(gclk));
	jdff dff_B_aH6Nh85K3_0(.din(w_dff_B_WMfun7bd3_0),.dout(w_dff_B_aH6Nh85K3_0),.clk(gclk));
	jdff dff_B_BWNbPEii0_0(.din(w_dff_B_aH6Nh85K3_0),.dout(w_dff_B_BWNbPEii0_0),.clk(gclk));
	jdff dff_B_BKEKWhze3_1(.din(n1160),.dout(w_dff_B_BKEKWhze3_1),.clk(gclk));
	jdff dff_B_FE6uwSmS0_1(.din(w_dff_B_BKEKWhze3_1),.dout(w_dff_B_FE6uwSmS0_1),.clk(gclk));
	jdff dff_A_7EUgJjEv4_1(.dout(w_n751_1[1]),.din(w_dff_A_7EUgJjEv4_1),.clk(gclk));
	jdff dff_A_BrrDWsJJ5_0(.dout(w_G123_0[0]),.din(w_dff_A_BrrDWsJJ5_0),.clk(gclk));
	jdff dff_B_k7ccmGjA3_2(.din(G123),.dout(w_dff_B_k7ccmGjA3_2),.clk(gclk));
	jdff dff_B_BCyhDCpA1_0(.din(n788),.dout(w_dff_B_BCyhDCpA1_0),.clk(gclk));
	jdff dff_B_JbPk5Cbw3_0(.din(n780),.dout(w_dff_B_JbPk5Cbw3_0),.clk(gclk));
	jdff dff_B_t0QenPJK3_0(.din(w_dff_B_JbPk5Cbw3_0),.dout(w_dff_B_t0QenPJK3_0),.clk(gclk));
	jdff dff_B_enuUWqnO6_0(.din(w_dff_B_t0QenPJK3_0),.dout(w_dff_B_enuUWqnO6_0),.clk(gclk));
	jdff dff_A_FMfDTZPu3_0(.dout(w_G54_0[0]),.din(w_dff_A_FMfDTZPu3_0),.clk(gclk));
	jdff dff_A_mAXDZyS17_0(.dout(w_dff_A_FMfDTZPu3_0),.din(w_dff_A_mAXDZyS17_0),.clk(gclk));
	jdff dff_A_d7HrMQip3_0(.dout(w_dff_A_mAXDZyS17_0),.din(w_dff_A_d7HrMQip3_0),.clk(gclk));
	jdff dff_A_6B2gmyQI5_0(.dout(w_dff_A_d7HrMQip3_0),.din(w_dff_A_6B2gmyQI5_0),.clk(gclk));
	jdff dff_A_lCuEXdLn1_0(.dout(w_dff_A_6B2gmyQI5_0),.din(w_dff_A_lCuEXdLn1_0),.clk(gclk));
	jdff dff_A_LqY3TKdd0_0(.dout(w_dff_A_lCuEXdLn1_0),.din(w_dff_A_LqY3TKdd0_0),.clk(gclk));
	jdff dff_A_jq7VWQt19_0(.dout(w_dff_A_LqY3TKdd0_0),.din(w_dff_A_jq7VWQt19_0),.clk(gclk));
	jdff dff_A_vpdtxn4N0_0(.dout(w_dff_A_jq7VWQt19_0),.din(w_dff_A_vpdtxn4N0_0),.clk(gclk));
	jdff dff_A_hGTaNu9B9_0(.dout(w_n741_0[0]),.din(w_dff_A_hGTaNu9B9_0),.clk(gclk));
	jdff dff_A_G8LGNIc74_0(.dout(w_dff_A_hGTaNu9B9_0),.din(w_dff_A_G8LGNIc74_0),.clk(gclk));
	jdff dff_A_cDwjwPSq8_0(.dout(w_dff_A_G8LGNIc74_0),.din(w_dff_A_cDwjwPSq8_0),.clk(gclk));
	jdff dff_A_NB5iNk0F7_0(.dout(w_dff_A_cDwjwPSq8_0),.din(w_dff_A_NB5iNk0F7_0),.clk(gclk));
	jdff dff_A_1J23STzd1_0(.dout(w_dff_A_NB5iNk0F7_0),.din(w_dff_A_1J23STzd1_0),.clk(gclk));
	jdff dff_A_sIKpZPM87_0(.dout(w_dff_A_1J23STzd1_0),.din(w_dff_A_sIKpZPM87_0),.clk(gclk));
	jdff dff_A_xo8iiHrd0_0(.dout(w_dff_A_sIKpZPM87_0),.din(w_dff_A_xo8iiHrd0_0),.clk(gclk));
	jdff dff_A_fqc6Redu2_0(.dout(w_n747_2[0]),.din(w_dff_A_fqc6Redu2_0),.clk(gclk));
	jdff dff_A_8apAwvBr9_0(.dout(w_dff_A_fqc6Redu2_0),.din(w_dff_A_8apAwvBr9_0),.clk(gclk));
	jdff dff_A_Myua4Nl51_0(.dout(w_dff_A_8apAwvBr9_0),.din(w_dff_A_Myua4Nl51_0),.clk(gclk));
	jdff dff_A_XOvFG1JA5_0(.dout(w_dff_A_Myua4Nl51_0),.din(w_dff_A_XOvFG1JA5_0),.clk(gclk));
	jdff dff_A_Zh3Fzkn12_0(.dout(w_dff_A_XOvFG1JA5_0),.din(w_dff_A_Zh3Fzkn12_0),.clk(gclk));
	jdff dff_A_4cCoBgTJ8_1(.dout(w_n747_2[1]),.din(w_dff_A_4cCoBgTJ8_1),.clk(gclk));
	jdff dff_A_q30IOs7B4_1(.dout(w_dff_A_4cCoBgTJ8_1),.din(w_dff_A_q30IOs7B4_1),.clk(gclk));
	jdff dff_A_0YA5gX3L0_1(.dout(w_dff_A_q30IOs7B4_1),.din(w_dff_A_0YA5gX3L0_1),.clk(gclk));
	jdff dff_A_tA6W320N7_1(.dout(w_dff_A_0YA5gX3L0_1),.din(w_dff_A_tA6W320N7_1),.clk(gclk));
	jdff dff_A_G7C3MKLi5_1(.dout(w_dff_A_tA6W320N7_1),.din(w_dff_A_G7C3MKLi5_1),.clk(gclk));
	jdff dff_A_mibvx99g4_1(.dout(w_dff_A_G7C3MKLi5_1),.din(w_dff_A_mibvx99g4_1),.clk(gclk));
	jdff dff_A_B163nOEO9_1(.dout(w_dff_A_mibvx99g4_1),.din(w_dff_A_B163nOEO9_1),.clk(gclk));
	jdff dff_A_B6nQ4l5Q2_1(.dout(w_dff_A_B163nOEO9_1),.din(w_dff_A_B6nQ4l5Q2_1),.clk(gclk));
	jdff dff_A_uvpUTQee1_1(.dout(w_dff_A_B6nQ4l5Q2_1),.din(w_dff_A_uvpUTQee1_1),.clk(gclk));
	jdff dff_B_QB6mvxpj1_0(.din(n1196),.dout(w_dff_B_QB6mvxpj1_0),.clk(gclk));
	jdff dff_B_bXm5ay248_0(.din(w_dff_B_QB6mvxpj1_0),.dout(w_dff_B_bXm5ay248_0),.clk(gclk));
	jdff dff_B_A0CdZTO27_0(.din(w_dff_B_bXm5ay248_0),.dout(w_dff_B_A0CdZTO27_0),.clk(gclk));
	jdff dff_B_DMr4WauW9_0(.din(w_dff_B_A0CdZTO27_0),.dout(w_dff_B_DMr4WauW9_0),.clk(gclk));
	jdff dff_B_inQ3U82g4_0(.din(w_dff_B_DMr4WauW9_0),.dout(w_dff_B_inQ3U82g4_0),.clk(gclk));
	jdff dff_B_aYmgZKAm5_0(.din(w_dff_B_inQ3U82g4_0),.dout(w_dff_B_aYmgZKAm5_0),.clk(gclk));
	jdff dff_B_KElNYV6G7_0(.din(w_dff_B_aYmgZKAm5_0),.dout(w_dff_B_KElNYV6G7_0),.clk(gclk));
	jdff dff_B_DBi65DCa4_0(.din(w_dff_B_KElNYV6G7_0),.dout(w_dff_B_DBi65DCa4_0),.clk(gclk));
	jdff dff_B_VY6FUyUR8_0(.din(w_dff_B_DBi65DCa4_0),.dout(w_dff_B_VY6FUyUR8_0),.clk(gclk));
	jdff dff_B_U2snLKEJ8_0(.din(w_dff_B_VY6FUyUR8_0),.dout(w_dff_B_U2snLKEJ8_0),.clk(gclk));
	jdff dff_B_NxDyucTm8_0(.din(w_dff_B_U2snLKEJ8_0),.dout(w_dff_B_NxDyucTm8_0),.clk(gclk));
	jdff dff_B_5R5KWFjg0_0(.din(w_dff_B_NxDyucTm8_0),.dout(w_dff_B_5R5KWFjg0_0),.clk(gclk));
	jdff dff_B_JUKEnXWI7_0(.din(n1195),.dout(w_dff_B_JUKEnXWI7_0),.clk(gclk));
	jdff dff_B_lhXixDxu4_0(.din(w_dff_B_JUKEnXWI7_0),.dout(w_dff_B_lhXixDxu4_0),.clk(gclk));
	jdff dff_B_2j8GxOw91_0(.din(w_dff_B_lhXixDxu4_0),.dout(w_dff_B_2j8GxOw91_0),.clk(gclk));
	jdff dff_B_20Y1p8ix0_0(.din(w_dff_B_2j8GxOw91_0),.dout(w_dff_B_20Y1p8ix0_0),.clk(gclk));
	jdff dff_B_P1l3ehr71_1(.din(G115),.dout(w_dff_B_P1l3ehr71_1),.clk(gclk));
	jdff dff_B_9G85qHLp6_1(.din(w_dff_B_P1l3ehr71_1),.dout(w_dff_B_9G85qHLp6_1),.clk(gclk));
	jdff dff_A_frt58SoM2_0(.dout(w_n751_0[0]),.din(w_dff_A_frt58SoM2_0),.clk(gclk));
	jdff dff_A_OYaMXLGe7_2(.dout(w_n751_0[2]),.din(w_dff_A_OYaMXLGe7_2),.clk(gclk));
	jdff dff_A_YKKmtzwo8_2(.dout(w_dff_A_OYaMXLGe7_2),.din(w_dff_A_YKKmtzwo8_2),.clk(gclk));
	jdff dff_A_LGVtW3Qv9_2(.dout(w_dff_A_YKKmtzwo8_2),.din(w_dff_A_LGVtW3Qv9_2),.clk(gclk));
	jdff dff_A_PvOiRHAm7_2(.dout(w_dff_A_LGVtW3Qv9_2),.din(w_dff_A_PvOiRHAm7_2),.clk(gclk));
	jdff dff_B_V0ZC5LCV6_1(.din(n929),.dout(w_dff_B_V0ZC5LCV6_1),.clk(gclk));
	jdff dff_B_F36k1EPQ8_1(.din(w_dff_B_V0ZC5LCV6_1),.dout(w_dff_B_F36k1EPQ8_1),.clk(gclk));
	jdff dff_B_zTMLTtux5_1(.din(w_dff_B_F36k1EPQ8_1),.dout(w_dff_B_zTMLTtux5_1),.clk(gclk));
	jdff dff_B_4RvYDFRq3_1(.din(w_dff_B_zTMLTtux5_1),.dout(w_dff_B_4RvYDFRq3_1),.clk(gclk));
	jdff dff_B_Uw8cvXCJ3_1(.din(w_dff_B_4RvYDFRq3_1),.dout(w_dff_B_Uw8cvXCJ3_1),.clk(gclk));
	jdff dff_B_KyJLUTO75_1(.din(w_dff_B_Uw8cvXCJ3_1),.dout(w_dff_B_KyJLUTO75_1),.clk(gclk));
	jdff dff_B_thd4XTy23_1(.din(w_dff_B_KyJLUTO75_1),.dout(w_dff_B_thd4XTy23_1),.clk(gclk));
	jdff dff_B_TG5KVz8b0_1(.din(w_dff_B_thd4XTy23_1),.dout(w_dff_B_TG5KVz8b0_1),.clk(gclk));
	jdff dff_B_Jbi5ZFtY8_1(.din(n931),.dout(w_dff_B_Jbi5ZFtY8_1),.clk(gclk));
	jdff dff_B_ErAA75Sg3_1(.din(w_dff_B_Jbi5ZFtY8_1),.dout(w_dff_B_ErAA75Sg3_1),.clk(gclk));
	jdff dff_B_2xvbEX6b6_1(.din(w_dff_B_ErAA75Sg3_1),.dout(w_dff_B_2xvbEX6b6_1),.clk(gclk));
	jdff dff_B_rBz9tB1n5_1(.din(w_dff_B_2xvbEX6b6_1),.dout(w_dff_B_rBz9tB1n5_1),.clk(gclk));
	jdff dff_B_xo2Xg6bR2_1(.din(w_dff_B_rBz9tB1n5_1),.dout(w_dff_B_xo2Xg6bR2_1),.clk(gclk));
	jdff dff_B_2TknPHmb6_1(.din(w_dff_B_xo2Xg6bR2_1),.dout(w_dff_B_2TknPHmb6_1),.clk(gclk));
	jdff dff_B_4BqlQqfc9_1(.din(w_dff_B_2TknPHmb6_1),.dout(w_dff_B_4BqlQqfc9_1),.clk(gclk));
	jdff dff_B_5knzVkgt4_1(.din(w_dff_B_4BqlQqfc9_1),.dout(w_dff_B_5knzVkgt4_1),.clk(gclk));
	jdff dff_B_nyszu3Qx9_1(.din(w_dff_B_5knzVkgt4_1),.dout(w_dff_B_nyszu3Qx9_1),.clk(gclk));
	jdff dff_B_PSye6bXg7_1(.din(w_dff_B_nyszu3Qx9_1),.dout(w_dff_B_PSye6bXg7_1),.clk(gclk));
	jdff dff_B_yZEvMHkQ1_0(.din(n935),.dout(w_dff_B_yZEvMHkQ1_0),.clk(gclk));
	jdff dff_A_bDtXZSfF2_1(.dout(w_G4_0[1]),.din(w_dff_A_bDtXZSfF2_1),.clk(gclk));
	jdff dff_A_aZsRZRzc4_1(.dout(w_dff_A_bDtXZSfF2_1),.din(w_dff_A_aZsRZRzc4_1),.clk(gclk));
	jdff dff_A_m6tBuxuy5_1(.dout(w_dff_A_aZsRZRzc4_1),.din(w_dff_A_m6tBuxuy5_1),.clk(gclk));
	jdff dff_A_LyJqcdhE2_1(.dout(w_dff_A_m6tBuxuy5_1),.din(w_dff_A_LyJqcdhE2_1),.clk(gclk));
	jdff dff_A_XQ85SI904_1(.dout(w_dff_A_LyJqcdhE2_1),.din(w_dff_A_XQ85SI904_1),.clk(gclk));
	jdff dff_A_KUzeLFZw3_1(.dout(w_dff_A_XQ85SI904_1),.din(w_dff_A_KUzeLFZw3_1),.clk(gclk));
	jdff dff_B_nm6Aqo8B0_3(.din(G4),.dout(w_dff_B_nm6Aqo8B0_3),.clk(gclk));
	jdff dff_B_iP6ndz3S4_3(.din(w_dff_B_nm6Aqo8B0_3),.dout(w_dff_B_iP6ndz3S4_3),.clk(gclk));
	jdff dff_B_CpQk12DH3_3(.din(w_dff_B_iP6ndz3S4_3),.dout(w_dff_B_CpQk12DH3_3),.clk(gclk));
	jdff dff_B_3zTcJTIs9_3(.din(w_dff_B_CpQk12DH3_3),.dout(w_dff_B_3zTcJTIs9_3),.clk(gclk));
	jdff dff_B_hPJG0ldp5_2(.din(n932),.dout(w_dff_B_hPJG0ldp5_2),.clk(gclk));
	jdff dff_B_GP2YH0ms9_2(.din(w_dff_B_hPJG0ldp5_2),.dout(w_dff_B_GP2YH0ms9_2),.clk(gclk));
	jdff dff_B_mWMwWwPY5_2(.din(w_dff_B_GP2YH0ms9_2),.dout(w_dff_B_mWMwWwPY5_2),.clk(gclk));
	jdff dff_B_vwcFlwia3_2(.din(w_dff_B_mWMwWwPY5_2),.dout(w_dff_B_vwcFlwia3_2),.clk(gclk));
	jdff dff_B_QYKlooOo9_2(.din(w_dff_B_vwcFlwia3_2),.dout(w_dff_B_QYKlooOo9_2),.clk(gclk));
	jdff dff_B_eTDh0uSx2_2(.din(w_dff_B_QYKlooOo9_2),.dout(w_dff_B_eTDh0uSx2_2),.clk(gclk));
	jdff dff_B_VN8rMfKo1_2(.din(w_dff_B_eTDh0uSx2_2),.dout(w_dff_B_VN8rMfKo1_2),.clk(gclk));
	jdff dff_B_RbRQ8xPU8_2(.din(w_dff_B_VN8rMfKo1_2),.dout(w_dff_B_RbRQ8xPU8_2),.clk(gclk));
	jdff dff_B_MVJDqufb2_2(.din(w_dff_B_RbRQ8xPU8_2),.dout(w_dff_B_MVJDqufb2_2),.clk(gclk));
	jdff dff_A_HLAl1M521_1(.dout(w_n747_1[1]),.din(w_dff_A_HLAl1M521_1),.clk(gclk));
	jdff dff_A_xFXK0hL58_1(.dout(w_dff_A_HLAl1M521_1),.din(w_dff_A_xFXK0hL58_1),.clk(gclk));
	jdff dff_A_VoHkmlRv2_1(.dout(w_dff_A_xFXK0hL58_1),.din(w_dff_A_VoHkmlRv2_1),.clk(gclk));
	jdff dff_A_PssrBKtE0_2(.dout(w_n747_1[2]),.din(w_dff_A_PssrBKtE0_2),.clk(gclk));
	jdff dff_A_uE9d4O748_2(.dout(w_dff_A_PssrBKtE0_2),.din(w_dff_A_uE9d4O748_2),.clk(gclk));
	jdff dff_A_ZDayzo5r4_2(.dout(w_dff_A_uE9d4O748_2),.din(w_dff_A_ZDayzo5r4_2),.clk(gclk));
	jdff dff_A_PRChFjBw1_2(.dout(w_dff_A_ZDayzo5r4_2),.din(w_dff_A_PRChFjBw1_2),.clk(gclk));
	jdff dff_A_05wwoAWZ0_0(.dout(w_n747_0[0]),.din(w_dff_A_05wwoAWZ0_0),.clk(gclk));
	jdff dff_A_CeJleYnU5_0(.dout(w_dff_A_05wwoAWZ0_0),.din(w_dff_A_CeJleYnU5_0),.clk(gclk));
	jdff dff_A_KzdNH0DK9_0(.dout(w_dff_A_CeJleYnU5_0),.din(w_dff_A_KzdNH0DK9_0),.clk(gclk));
	jdff dff_A_oieLvGfZ1_0(.dout(w_dff_A_KzdNH0DK9_0),.din(w_dff_A_oieLvGfZ1_0),.clk(gclk));
	jdff dff_A_0FC9zjOJ3_0(.dout(w_dff_A_oieLvGfZ1_0),.din(w_dff_A_0FC9zjOJ3_0),.clk(gclk));
	jdff dff_A_h5iRJ6oW1_0(.dout(w_dff_A_0FC9zjOJ3_0),.din(w_dff_A_h5iRJ6oW1_0),.clk(gclk));
	jdff dff_A_rCFMe4uN1_0(.dout(w_dff_A_h5iRJ6oW1_0),.din(w_dff_A_rCFMe4uN1_0),.clk(gclk));
	jdff dff_A_PKfuQANw6_0(.dout(w_dff_A_rCFMe4uN1_0),.din(w_dff_A_PKfuQANw6_0),.clk(gclk));
	jdff dff_A_oKPUfezU1_0(.dout(w_dff_A_PKfuQANw6_0),.din(w_dff_A_oKPUfezU1_0),.clk(gclk));
	jdff dff_A_UXYtXNr46_0(.dout(w_dff_A_oKPUfezU1_0),.din(w_dff_A_UXYtXNr46_0),.clk(gclk));
	jdff dff_A_dhsvvXga0_0(.dout(w_dff_A_UXYtXNr46_0),.din(w_dff_A_dhsvvXga0_0),.clk(gclk));
	jdff dff_A_W1gUI3au0_0(.dout(w_dff_A_dhsvvXga0_0),.din(w_dff_A_W1gUI3au0_0),.clk(gclk));
	jdff dff_A_LoCCPFDQ2_0(.dout(w_dff_A_W1gUI3au0_0),.din(w_dff_A_LoCCPFDQ2_0),.clk(gclk));
	jdff dff_A_njKGqq1g9_1(.dout(w_n747_0[1]),.din(w_dff_A_njKGqq1g9_1),.clk(gclk));
	jdff dff_A_bzzNAAMX7_1(.dout(w_dff_A_njKGqq1g9_1),.din(w_dff_A_bzzNAAMX7_1),.clk(gclk));
	jdff dff_A_DeQWqwRF8_1(.dout(w_dff_A_bzzNAAMX7_1),.din(w_dff_A_DeQWqwRF8_1),.clk(gclk));
	jdff dff_A_Hulc4xtm9_1(.dout(w_dff_A_DeQWqwRF8_1),.din(w_dff_A_Hulc4xtm9_1),.clk(gclk));
	jdff dff_A_vtSH9Vbn1_1(.dout(w_dff_A_Hulc4xtm9_1),.din(w_dff_A_vtSH9Vbn1_1),.clk(gclk));
	jdff dff_A_NWZp0gGh3_1(.dout(w_dff_A_vtSH9Vbn1_1),.din(w_dff_A_NWZp0gGh3_1),.clk(gclk));
	jdff dff_A_Xu5BlIp72_1(.dout(w_dff_A_NWZp0gGh3_1),.din(w_dff_A_Xu5BlIp72_1),.clk(gclk));
	jdff dff_B_hWyTCKRT3_1(.din(n1388),.dout(w_dff_B_hWyTCKRT3_1),.clk(gclk));
	jdff dff_B_VDLvyCjj0_1(.din(w_dff_B_hWyTCKRT3_1),.dout(w_dff_B_VDLvyCjj0_1),.clk(gclk));
	jdff dff_B_sbds70jh7_1(.din(w_dff_B_VDLvyCjj0_1),.dout(w_dff_B_sbds70jh7_1),.clk(gclk));
	jdff dff_B_xVKvmOMW7_1(.din(w_dff_B_sbds70jh7_1),.dout(w_dff_B_xVKvmOMW7_1),.clk(gclk));
	jdff dff_B_NAl70N4K8_1(.din(w_dff_B_xVKvmOMW7_1),.dout(w_dff_B_NAl70N4K8_1),.clk(gclk));
	jdff dff_B_5xB1GOzx7_1(.din(w_dff_B_NAl70N4K8_1),.dout(w_dff_B_5xB1GOzx7_1),.clk(gclk));
	jdff dff_B_AoYBY6MI2_1(.din(w_dff_B_5xB1GOzx7_1),.dout(w_dff_B_AoYBY6MI2_1),.clk(gclk));
	jdff dff_B_TtEPmjQ46_1(.din(w_dff_B_AoYBY6MI2_1),.dout(w_dff_B_TtEPmjQ46_1),.clk(gclk));
	jdff dff_B_clzf3T6G8_1(.din(w_dff_B_TtEPmjQ46_1),.dout(w_dff_B_clzf3T6G8_1),.clk(gclk));
	jdff dff_B_cFeYhvnw4_1(.din(w_dff_B_clzf3T6G8_1),.dout(w_dff_B_cFeYhvnw4_1),.clk(gclk));
	jdff dff_B_CJ9UndW83_1(.din(w_dff_B_cFeYhvnw4_1),.dout(w_dff_B_CJ9UndW83_1),.clk(gclk));
	jdff dff_B_N5MmGJLS4_1(.din(w_dff_B_CJ9UndW83_1),.dout(w_dff_B_N5MmGJLS4_1),.clk(gclk));
	jdff dff_B_8DsBHhks9_1(.din(w_dff_B_N5MmGJLS4_1),.dout(w_dff_B_8DsBHhks9_1),.clk(gclk));
	jdff dff_B_guLETHEL6_1(.din(w_dff_B_8DsBHhks9_1),.dout(w_dff_B_guLETHEL6_1),.clk(gclk));
	jdff dff_B_RO1PxrYt8_1(.din(w_dff_B_guLETHEL6_1),.dout(w_dff_B_RO1PxrYt8_1),.clk(gclk));
	jdff dff_B_NlmNpPso8_1(.din(w_dff_B_RO1PxrYt8_1),.dout(w_dff_B_NlmNpPso8_1),.clk(gclk));
	jdff dff_B_uTZn3X140_1(.din(w_dff_B_NlmNpPso8_1),.dout(w_dff_B_uTZn3X140_1),.clk(gclk));
	jdff dff_B_O590Tvgi3_1(.din(w_dff_B_uTZn3X140_1),.dout(w_dff_B_O590Tvgi3_1),.clk(gclk));
	jdff dff_B_pt4Np9lk0_1(.din(w_dff_B_O590Tvgi3_1),.dout(w_dff_B_pt4Np9lk0_1),.clk(gclk));
	jdff dff_B_2fu0Yukz0_1(.din(n1539),.dout(w_dff_B_2fu0Yukz0_1),.clk(gclk));
	jdff dff_B_XKFhEpvU7_1(.din(w_dff_B_2fu0Yukz0_1),.dout(w_dff_B_XKFhEpvU7_1),.clk(gclk));
	jdff dff_B_X16GS3k32_1(.din(w_dff_B_XKFhEpvU7_1),.dout(w_dff_B_X16GS3k32_1),.clk(gclk));
	jdff dff_B_lEZqV0FP4_1(.din(w_dff_B_X16GS3k32_1),.dout(w_dff_B_lEZqV0FP4_1),.clk(gclk));
	jdff dff_B_d00V3A903_1(.din(w_dff_B_lEZqV0FP4_1),.dout(w_dff_B_d00V3A903_1),.clk(gclk));
	jdff dff_B_SiQpf2OB4_1(.din(w_dff_B_d00V3A903_1),.dout(w_dff_B_SiQpf2OB4_1),.clk(gclk));
	jdff dff_B_37Wt5caT1_1(.din(w_dff_B_SiQpf2OB4_1),.dout(w_dff_B_37Wt5caT1_1),.clk(gclk));
	jdff dff_B_isjrsp5R5_1(.din(w_dff_B_37Wt5caT1_1),.dout(w_dff_B_isjrsp5R5_1),.clk(gclk));
	jdff dff_B_3Szipj2D7_1(.din(w_dff_B_isjrsp5R5_1),.dout(w_dff_B_3Szipj2D7_1),.clk(gclk));
	jdff dff_B_2ltHrkJs4_1(.din(w_dff_B_3Szipj2D7_1),.dout(w_dff_B_2ltHrkJs4_1),.clk(gclk));
	jdff dff_B_nZ2gg8PF1_1(.din(w_dff_B_2ltHrkJs4_1),.dout(w_dff_B_nZ2gg8PF1_1),.clk(gclk));
	jdff dff_B_AxlY0AT22_1(.din(w_dff_B_nZ2gg8PF1_1),.dout(w_dff_B_AxlY0AT22_1),.clk(gclk));
	jdff dff_B_sqUS6HAx9_1(.din(w_dff_B_AxlY0AT22_1),.dout(w_dff_B_sqUS6HAx9_1),.clk(gclk));
	jdff dff_B_xiX3QdBV9_1(.din(w_dff_B_sqUS6HAx9_1),.dout(w_dff_B_xiX3QdBV9_1),.clk(gclk));
	jdff dff_B_JpiBi7vB6_1(.din(w_dff_B_xiX3QdBV9_1),.dout(w_dff_B_JpiBi7vB6_1),.clk(gclk));
	jdff dff_B_LESUyLpb0_1(.din(w_dff_B_JpiBi7vB6_1),.dout(w_dff_B_LESUyLpb0_1),.clk(gclk));
	jdff dff_B_9zXaKAsG7_1(.din(w_dff_B_LESUyLpb0_1),.dout(w_dff_B_9zXaKAsG7_1),.clk(gclk));
	jdff dff_B_BYPKNXFo4_1(.din(w_dff_B_9zXaKAsG7_1),.dout(w_dff_B_BYPKNXFo4_1),.clk(gclk));
	jdff dff_B_bUlMydrC4_1(.din(w_dff_B_BYPKNXFo4_1),.dout(w_dff_B_bUlMydrC4_1),.clk(gclk));
	jdff dff_B_Oyc7erkj0_0(.din(n1614),.dout(w_dff_B_Oyc7erkj0_0),.clk(gclk));
	jdff dff_B_3UQXGzYe1_0(.din(w_dff_B_Oyc7erkj0_0),.dout(w_dff_B_3UQXGzYe1_0),.clk(gclk));
	jdff dff_B_p9iI1GCm6_0(.din(w_dff_B_3UQXGzYe1_0),.dout(w_dff_B_p9iI1GCm6_0),.clk(gclk));
	jdff dff_B_Fv8oce7b2_0(.din(w_dff_B_p9iI1GCm6_0),.dout(w_dff_B_Fv8oce7b2_0),.clk(gclk));
	jdff dff_B_xfdXn3gh8_0(.din(w_dff_B_Fv8oce7b2_0),.dout(w_dff_B_xfdXn3gh8_0),.clk(gclk));
	jdff dff_B_24RTbt2l6_0(.din(w_dff_B_xfdXn3gh8_0),.dout(w_dff_B_24RTbt2l6_0),.clk(gclk));
	jdff dff_B_T5QHiW5g4_0(.din(w_dff_B_24RTbt2l6_0),.dout(w_dff_B_T5QHiW5g4_0),.clk(gclk));
	jdff dff_B_XUHRBrMY2_0(.din(w_dff_B_T5QHiW5g4_0),.dout(w_dff_B_XUHRBrMY2_0),.clk(gclk));
	jdff dff_B_rM8hLnGy8_0(.din(w_dff_B_XUHRBrMY2_0),.dout(w_dff_B_rM8hLnGy8_0),.clk(gclk));
	jdff dff_B_8nFpynAk6_0(.din(w_dff_B_rM8hLnGy8_0),.dout(w_dff_B_8nFpynAk6_0),.clk(gclk));
	jdff dff_B_6O0TcsTE8_0(.din(w_dff_B_8nFpynAk6_0),.dout(w_dff_B_6O0TcsTE8_0),.clk(gclk));
	jdff dff_B_1ERHSp2e2_0(.din(w_dff_B_6O0TcsTE8_0),.dout(w_dff_B_1ERHSp2e2_0),.clk(gclk));
	jdff dff_B_KgQ5RStM5_0(.din(w_dff_B_1ERHSp2e2_0),.dout(w_dff_B_KgQ5RStM5_0),.clk(gclk));
	jdff dff_B_iQkfhazn3_0(.din(w_dff_B_KgQ5RStM5_0),.dout(w_dff_B_iQkfhazn3_0),.clk(gclk));
	jdff dff_B_YxjzLB4X2_0(.din(w_dff_B_iQkfhazn3_0),.dout(w_dff_B_YxjzLB4X2_0),.clk(gclk));
	jdff dff_B_A6trlIz93_0(.din(w_dff_B_YxjzLB4X2_0),.dout(w_dff_B_A6trlIz93_0),.clk(gclk));
	jdff dff_B_7CFLzJwE9_0(.din(w_dff_B_A6trlIz93_0),.dout(w_dff_B_7CFLzJwE9_0),.clk(gclk));
	jdff dff_B_Acos7NPE2_0(.din(w_dff_B_7CFLzJwE9_0),.dout(w_dff_B_Acos7NPE2_0),.clk(gclk));
	jdff dff_B_pn9fF3NJ2_0(.din(w_dff_B_Acos7NPE2_0),.dout(w_dff_B_pn9fF3NJ2_0),.clk(gclk));
	jdff dff_B_zVkRJpEp9_0(.din(n1613),.dout(w_dff_B_zVkRJpEp9_0),.clk(gclk));
	jdff dff_A_gDFl44Nf8_1(.dout(w_n797_1[1]),.din(w_dff_A_gDFl44Nf8_1),.clk(gclk));
	jdff dff_A_QK4tJ5KJ2_1(.dout(w_dff_A_gDFl44Nf8_1),.din(w_dff_A_QK4tJ5KJ2_1),.clk(gclk));
	jdff dff_A_WTFoR4Xs3_1(.dout(w_dff_A_QK4tJ5KJ2_1),.din(w_dff_A_WTFoR4Xs3_1),.clk(gclk));
	jdff dff_A_WnvQZK9R1_1(.dout(w_dff_A_WTFoR4Xs3_1),.din(w_dff_A_WnvQZK9R1_1),.clk(gclk));
	jdff dff_A_YYBwUoaC1_1(.dout(w_dff_A_WnvQZK9R1_1),.din(w_dff_A_YYBwUoaC1_1),.clk(gclk));
	jdff dff_A_Vv1X4RK16_1(.dout(w_dff_A_YYBwUoaC1_1),.din(w_dff_A_Vv1X4RK16_1),.clk(gclk));
	jdff dff_A_6t5wCJPH9_1(.dout(w_dff_A_Vv1X4RK16_1),.din(w_dff_A_6t5wCJPH9_1),.clk(gclk));
	jdff dff_A_nloeYeZH8_1(.dout(w_dff_A_6t5wCJPH9_1),.din(w_dff_A_nloeYeZH8_1),.clk(gclk));
	jdff dff_A_Zb1Np2Q13_1(.dout(w_dff_A_nloeYeZH8_1),.din(w_dff_A_Zb1Np2Q13_1),.clk(gclk));
	jdff dff_A_hOA9568S6_1(.dout(w_dff_A_Zb1Np2Q13_1),.din(w_dff_A_hOA9568S6_1),.clk(gclk));
	jdff dff_A_iywbZGbf1_1(.dout(w_dff_A_hOA9568S6_1),.din(w_dff_A_iywbZGbf1_1),.clk(gclk));
	jdff dff_A_TgEIV9iS0_1(.dout(w_dff_A_iywbZGbf1_1),.din(w_dff_A_TgEIV9iS0_1),.clk(gclk));
	jdff dff_A_y3HvpBwO3_1(.dout(w_dff_A_TgEIV9iS0_1),.din(w_dff_A_y3HvpBwO3_1),.clk(gclk));
	jdff dff_A_wr4dtUjX9_1(.dout(w_dff_A_y3HvpBwO3_1),.din(w_dff_A_wr4dtUjX9_1),.clk(gclk));
	jdff dff_A_rKVaqn901_2(.dout(w_n797_1[2]),.din(w_dff_A_rKVaqn901_2),.clk(gclk));
	jdff dff_A_ldK5lY4G6_2(.dout(w_dff_A_rKVaqn901_2),.din(w_dff_A_ldK5lY4G6_2),.clk(gclk));
	jdff dff_A_681pEa5P3_2(.dout(w_dff_A_ldK5lY4G6_2),.din(w_dff_A_681pEa5P3_2),.clk(gclk));
	jdff dff_A_XDMjJR8f2_2(.dout(w_dff_A_681pEa5P3_2),.din(w_dff_A_XDMjJR8f2_2),.clk(gclk));
	jdff dff_A_SwdNfqQS8_2(.dout(w_dff_A_XDMjJR8f2_2),.din(w_dff_A_SwdNfqQS8_2),.clk(gclk));
	jdff dff_A_1IUCxP8Q5_2(.dout(w_dff_A_SwdNfqQS8_2),.din(w_dff_A_1IUCxP8Q5_2),.clk(gclk));
	jdff dff_A_SjRh2TnK2_2(.dout(w_dff_A_1IUCxP8Q5_2),.din(w_dff_A_SjRh2TnK2_2),.clk(gclk));
	jdff dff_A_wffqRqnD2_2(.dout(w_dff_A_SjRh2TnK2_2),.din(w_dff_A_wffqRqnD2_2),.clk(gclk));
	jdff dff_A_9b4ItQma5_2(.dout(w_dff_A_wffqRqnD2_2),.din(w_dff_A_9b4ItQma5_2),.clk(gclk));
	jdff dff_A_AJGiieCM9_2(.dout(w_dff_A_9b4ItQma5_2),.din(w_dff_A_AJGiieCM9_2),.clk(gclk));
	jdff dff_A_Zxi2yntb3_1(.dout(w_n797_0[1]),.din(w_dff_A_Zxi2yntb3_1),.clk(gclk));
	jdff dff_A_iW9kNU8j2_1(.dout(w_dff_A_Zxi2yntb3_1),.din(w_dff_A_iW9kNU8j2_1),.clk(gclk));
	jdff dff_A_P6fUHoeO5_1(.dout(w_dff_A_iW9kNU8j2_1),.din(w_dff_A_P6fUHoeO5_1),.clk(gclk));
	jdff dff_A_YyMhI7br9_1(.dout(w_dff_A_P6fUHoeO5_1),.din(w_dff_A_YyMhI7br9_1),.clk(gclk));
	jdff dff_A_hFiRqPYe5_1(.dout(w_dff_A_YyMhI7br9_1),.din(w_dff_A_hFiRqPYe5_1),.clk(gclk));
	jdff dff_A_9yNuijDT7_1(.dout(w_dff_A_hFiRqPYe5_1),.din(w_dff_A_9yNuijDT7_1),.clk(gclk));
	jdff dff_A_J9s8QZEi9_1(.dout(w_dff_A_9yNuijDT7_1),.din(w_dff_A_J9s8QZEi9_1),.clk(gclk));
	jdff dff_A_5fop84UG1_1(.dout(w_dff_A_J9s8QZEi9_1),.din(w_dff_A_5fop84UG1_1),.clk(gclk));
	jdff dff_A_ZFi2FESZ2_1(.dout(w_dff_A_5fop84UG1_1),.din(w_dff_A_ZFi2FESZ2_1),.clk(gclk));
	jdff dff_A_oRQ7d04F4_1(.dout(w_dff_A_ZFi2FESZ2_1),.din(w_dff_A_oRQ7d04F4_1),.clk(gclk));
	jdff dff_A_MsSSaf845_1(.dout(w_dff_A_oRQ7d04F4_1),.din(w_dff_A_MsSSaf845_1),.clk(gclk));
	jdff dff_A_dsfKY5Mi9_2(.dout(w_n797_0[2]),.din(w_dff_A_dsfKY5Mi9_2),.clk(gclk));
	jdff dff_B_Jj9PwHD67_3(.din(n797),.dout(w_dff_B_Jj9PwHD67_3),.clk(gclk));
	jdff dff_B_4yw7WmsD5_3(.din(w_dff_B_Jj9PwHD67_3),.dout(w_dff_B_4yw7WmsD5_3),.clk(gclk));
	jdff dff_B_z3NZq9r76_3(.din(w_dff_B_4yw7WmsD5_3),.dout(w_dff_B_z3NZq9r76_3),.clk(gclk));
	jdff dff_B_i40G09E43_3(.din(w_dff_B_z3NZq9r76_3),.dout(w_dff_B_i40G09E43_3),.clk(gclk));
	jdff dff_B_BWtFMQnv4_3(.din(w_dff_B_i40G09E43_3),.dout(w_dff_B_BWtFMQnv4_3),.clk(gclk));
	jdff dff_B_XABObqKV1_3(.din(w_dff_B_BWtFMQnv4_3),.dout(w_dff_B_XABObqKV1_3),.clk(gclk));
	jdff dff_A_09hrrOSP0_1(.dout(w_n793_1[1]),.din(w_dff_A_09hrrOSP0_1),.clk(gclk));
	jdff dff_A_ICxSbAIE1_1(.dout(w_dff_A_09hrrOSP0_1),.din(w_dff_A_ICxSbAIE1_1),.clk(gclk));
	jdff dff_A_4bNrqtOu9_1(.dout(w_dff_A_ICxSbAIE1_1),.din(w_dff_A_4bNrqtOu9_1),.clk(gclk));
	jdff dff_A_56k5cqEv8_1(.dout(w_dff_A_4bNrqtOu9_1),.din(w_dff_A_56k5cqEv8_1),.clk(gclk));
	jdff dff_A_zei0RHmK3_1(.dout(w_dff_A_56k5cqEv8_1),.din(w_dff_A_zei0RHmK3_1),.clk(gclk));
	jdff dff_A_rmTAStox6_1(.dout(w_dff_A_zei0RHmK3_1),.din(w_dff_A_rmTAStox6_1),.clk(gclk));
	jdff dff_A_LIfvZvJn4_1(.dout(w_dff_A_rmTAStox6_1),.din(w_dff_A_LIfvZvJn4_1),.clk(gclk));
	jdff dff_A_AoZXPVz36_1(.dout(w_dff_A_LIfvZvJn4_1),.din(w_dff_A_AoZXPVz36_1),.clk(gclk));
	jdff dff_A_6wYzzrQc6_1(.dout(w_dff_A_AoZXPVz36_1),.din(w_dff_A_6wYzzrQc6_1),.clk(gclk));
	jdff dff_A_GJPIIFRs0_1(.dout(w_dff_A_6wYzzrQc6_1),.din(w_dff_A_GJPIIFRs0_1),.clk(gclk));
	jdff dff_A_d3nwqLTE2_1(.dout(w_dff_A_GJPIIFRs0_1),.din(w_dff_A_d3nwqLTE2_1),.clk(gclk));
	jdff dff_A_AhPdWlgx8_1(.dout(w_dff_A_d3nwqLTE2_1),.din(w_dff_A_AhPdWlgx8_1),.clk(gclk));
	jdff dff_A_qeOascDE5_1(.dout(w_dff_A_AhPdWlgx8_1),.din(w_dff_A_qeOascDE5_1),.clk(gclk));
	jdff dff_A_xjWfmCDl7_1(.dout(w_dff_A_qeOascDE5_1),.din(w_dff_A_xjWfmCDl7_1),.clk(gclk));
	jdff dff_A_y0oRANoW6_2(.dout(w_n793_1[2]),.din(w_dff_A_y0oRANoW6_2),.clk(gclk));
	jdff dff_A_Kzu7LfBS5_2(.dout(w_dff_A_y0oRANoW6_2),.din(w_dff_A_Kzu7LfBS5_2),.clk(gclk));
	jdff dff_A_ePmZYUO09_2(.dout(w_dff_A_Kzu7LfBS5_2),.din(w_dff_A_ePmZYUO09_2),.clk(gclk));
	jdff dff_A_6XrdGx970_2(.dout(w_dff_A_ePmZYUO09_2),.din(w_dff_A_6XrdGx970_2),.clk(gclk));
	jdff dff_A_9HOSXcbI1_2(.dout(w_dff_A_6XrdGx970_2),.din(w_dff_A_9HOSXcbI1_2),.clk(gclk));
	jdff dff_A_v7rzEFQq9_2(.dout(w_dff_A_9HOSXcbI1_2),.din(w_dff_A_v7rzEFQq9_2),.clk(gclk));
	jdff dff_A_kSD2nT7G3_2(.dout(w_dff_A_v7rzEFQq9_2),.din(w_dff_A_kSD2nT7G3_2),.clk(gclk));
	jdff dff_A_taAU0pJb7_2(.dout(w_dff_A_kSD2nT7G3_2),.din(w_dff_A_taAU0pJb7_2),.clk(gclk));
	jdff dff_A_bktD94j34_2(.dout(w_dff_A_taAU0pJb7_2),.din(w_dff_A_bktD94j34_2),.clk(gclk));
	jdff dff_A_S5eA9kuy6_2(.dout(w_dff_A_bktD94j34_2),.din(w_dff_A_S5eA9kuy6_2),.clk(gclk));
	jdff dff_A_ODzzS0E23_1(.dout(w_n793_0[1]),.din(w_dff_A_ODzzS0E23_1),.clk(gclk));
	jdff dff_A_NB3Sle5t5_1(.dout(w_dff_A_ODzzS0E23_1),.din(w_dff_A_NB3Sle5t5_1),.clk(gclk));
	jdff dff_A_4yarnEib1_1(.dout(w_dff_A_NB3Sle5t5_1),.din(w_dff_A_4yarnEib1_1),.clk(gclk));
	jdff dff_A_mzgCjKZS7_1(.dout(w_dff_A_4yarnEib1_1),.din(w_dff_A_mzgCjKZS7_1),.clk(gclk));
	jdff dff_A_a1MPQaHw2_1(.dout(w_dff_A_mzgCjKZS7_1),.din(w_dff_A_a1MPQaHw2_1),.clk(gclk));
	jdff dff_A_vcICGs300_1(.dout(w_dff_A_a1MPQaHw2_1),.din(w_dff_A_vcICGs300_1),.clk(gclk));
	jdff dff_A_A7zNrVPA7_1(.dout(w_dff_A_vcICGs300_1),.din(w_dff_A_A7zNrVPA7_1),.clk(gclk));
	jdff dff_A_VzlFDMJE1_1(.dout(w_dff_A_A7zNrVPA7_1),.din(w_dff_A_VzlFDMJE1_1),.clk(gclk));
	jdff dff_A_60iMxWrC7_1(.dout(w_dff_A_VzlFDMJE1_1),.din(w_dff_A_60iMxWrC7_1),.clk(gclk));
	jdff dff_A_NlNYudBi9_1(.dout(w_dff_A_60iMxWrC7_1),.din(w_dff_A_NlNYudBi9_1),.clk(gclk));
	jdff dff_A_rbDetDgH9_1(.dout(w_dff_A_NlNYudBi9_1),.din(w_dff_A_rbDetDgH9_1),.clk(gclk));
	jdff dff_A_SX3MLxt72_2(.dout(w_n793_0[2]),.din(w_dff_A_SX3MLxt72_2),.clk(gclk));
	jdff dff_A_02duTM8P5_2(.dout(w_dff_A_SX3MLxt72_2),.din(w_dff_A_02duTM8P5_2),.clk(gclk));
	jdff dff_A_x3tz2ruC5_2(.dout(w_dff_A_02duTM8P5_2),.din(w_dff_A_x3tz2ruC5_2),.clk(gclk));
	jdff dff_A_4S0qJLoI6_2(.dout(w_dff_A_x3tz2ruC5_2),.din(w_dff_A_4S0qJLoI6_2),.clk(gclk));
	jdff dff_B_zmntCGcZ5_3(.din(n793),.dout(w_dff_B_zmntCGcZ5_3),.clk(gclk));
	jdff dff_B_hc2jIxY07_3(.din(w_dff_B_zmntCGcZ5_3),.dout(w_dff_B_hc2jIxY07_3),.clk(gclk));
	jdff dff_B_F7pcUx834_3(.din(w_dff_B_hc2jIxY07_3),.dout(w_dff_B_F7pcUx834_3),.clk(gclk));
	jdff dff_B_SwKN3pzG4_3(.din(w_dff_B_F7pcUx834_3),.dout(w_dff_B_SwKN3pzG4_3),.clk(gclk));
	jdff dff_B_tAHh98pf8_3(.din(w_dff_B_SwKN3pzG4_3),.dout(w_dff_B_tAHh98pf8_3),.clk(gclk));
	jdff dff_B_YW0PqZyk2_3(.din(w_dff_B_tAHh98pf8_3),.dout(w_dff_B_YW0PqZyk2_3),.clk(gclk));
	jdff dff_B_dFN2gYon5_3(.din(w_dff_B_YW0PqZyk2_3),.dout(w_dff_B_dFN2gYon5_3),.clk(gclk));
	jdff dff_A_Ts5zBysZ3_2(.dout(w_G4088_0[2]),.din(w_dff_A_Ts5zBysZ3_2),.clk(gclk));
	jdff dff_A_Jh1PO9Ub9_1(.dout(w_G4087_0[1]),.din(w_dff_A_Jh1PO9Ub9_1),.clk(gclk));
	jdff dff_B_zaTCGnqh1_0(.din(n1621),.dout(w_dff_B_zaTCGnqh1_0),.clk(gclk));
	jdff dff_B_PAWhwoeG8_0(.din(w_dff_B_zaTCGnqh1_0),.dout(w_dff_B_PAWhwoeG8_0),.clk(gclk));
	jdff dff_B_PfRReHWk3_0(.din(w_dff_B_PAWhwoeG8_0),.dout(w_dff_B_PfRReHWk3_0),.clk(gclk));
	jdff dff_B_11Gsk3zY7_0(.din(w_dff_B_PfRReHWk3_0),.dout(w_dff_B_11Gsk3zY7_0),.clk(gclk));
	jdff dff_B_QYWkJchj3_0(.din(w_dff_B_11Gsk3zY7_0),.dout(w_dff_B_QYWkJchj3_0),.clk(gclk));
	jdff dff_B_3vcKBv499_0(.din(w_dff_B_QYWkJchj3_0),.dout(w_dff_B_3vcKBv499_0),.clk(gclk));
	jdff dff_B_R3xUY0fx2_0(.din(w_dff_B_3vcKBv499_0),.dout(w_dff_B_R3xUY0fx2_0),.clk(gclk));
	jdff dff_B_F1YHIbtk3_0(.din(w_dff_B_R3xUY0fx2_0),.dout(w_dff_B_F1YHIbtk3_0),.clk(gclk));
	jdff dff_B_MGpcTcz82_0(.din(w_dff_B_F1YHIbtk3_0),.dout(w_dff_B_MGpcTcz82_0),.clk(gclk));
	jdff dff_B_wlON81Hb1_0(.din(w_dff_B_MGpcTcz82_0),.dout(w_dff_B_wlON81Hb1_0),.clk(gclk));
	jdff dff_B_9LPqMGjj0_0(.din(w_dff_B_wlON81Hb1_0),.dout(w_dff_B_9LPqMGjj0_0),.clk(gclk));
	jdff dff_B_BGfBg8vY1_0(.din(w_dff_B_9LPqMGjj0_0),.dout(w_dff_B_BGfBg8vY1_0),.clk(gclk));
	jdff dff_B_eT7K70c91_0(.din(w_dff_B_BGfBg8vY1_0),.dout(w_dff_B_eT7K70c91_0),.clk(gclk));
	jdff dff_B_1vmN5luf3_0(.din(w_dff_B_eT7K70c91_0),.dout(w_dff_B_1vmN5luf3_0),.clk(gclk));
	jdff dff_B_5KAjjyVv9_0(.din(w_dff_B_1vmN5luf3_0),.dout(w_dff_B_5KAjjyVv9_0),.clk(gclk));
	jdff dff_B_08wO1yN45_0(.din(w_dff_B_5KAjjyVv9_0),.dout(w_dff_B_08wO1yN45_0),.clk(gclk));
	jdff dff_B_IkqgK7uJ3_0(.din(w_dff_B_08wO1yN45_0),.dout(w_dff_B_IkqgK7uJ3_0),.clk(gclk));
	jdff dff_B_Qrk93bQG4_0(.din(w_dff_B_IkqgK7uJ3_0),.dout(w_dff_B_Qrk93bQG4_0),.clk(gclk));
	jdff dff_B_vy2zsUTI4_0(.din(w_dff_B_Qrk93bQG4_0),.dout(w_dff_B_vy2zsUTI4_0),.clk(gclk));
	jdff dff_B_Iw1JI7LE5_0(.din(n1620),.dout(w_dff_B_Iw1JI7LE5_0),.clk(gclk));
	jdff dff_B_tjMC8laf8_2(.din(G64),.dout(w_dff_B_tjMC8laf8_2),.clk(gclk));
	jdff dff_B_R6qd8A5o3_2(.din(G14),.dout(w_dff_B_R6qd8A5o3_2),.clk(gclk));
	jdff dff_B_UE8GuEbX6_2(.din(w_dff_B_R6qd8A5o3_2),.dout(w_dff_B_UE8GuEbX6_2),.clk(gclk));
	jdff dff_A_Bw91KRzU6_1(.dout(w_n843_1[1]),.din(w_dff_A_Bw91KRzU6_1),.clk(gclk));
	jdff dff_A_mFSizQAB5_1(.dout(w_dff_A_Bw91KRzU6_1),.din(w_dff_A_mFSizQAB5_1),.clk(gclk));
	jdff dff_A_Tcv2PsEN5_1(.dout(w_dff_A_mFSizQAB5_1),.din(w_dff_A_Tcv2PsEN5_1),.clk(gclk));
	jdff dff_A_U4ln5SHA2_1(.dout(w_dff_A_Tcv2PsEN5_1),.din(w_dff_A_U4ln5SHA2_1),.clk(gclk));
	jdff dff_A_2Gept2Jo6_1(.dout(w_dff_A_U4ln5SHA2_1),.din(w_dff_A_2Gept2Jo6_1),.clk(gclk));
	jdff dff_A_KYNLNk6S2_1(.dout(w_dff_A_2Gept2Jo6_1),.din(w_dff_A_KYNLNk6S2_1),.clk(gclk));
	jdff dff_A_UIvSCv7u3_1(.dout(w_dff_A_KYNLNk6S2_1),.din(w_dff_A_UIvSCv7u3_1),.clk(gclk));
	jdff dff_A_0f3R6dKC7_1(.dout(w_dff_A_UIvSCv7u3_1),.din(w_dff_A_0f3R6dKC7_1),.clk(gclk));
	jdff dff_A_rTCv7y8G5_1(.dout(w_dff_A_0f3R6dKC7_1),.din(w_dff_A_rTCv7y8G5_1),.clk(gclk));
	jdff dff_A_NXzMwWYT0_1(.dout(w_dff_A_rTCv7y8G5_1),.din(w_dff_A_NXzMwWYT0_1),.clk(gclk));
	jdff dff_A_7Wvx59Ze7_1(.dout(w_dff_A_NXzMwWYT0_1),.din(w_dff_A_7Wvx59Ze7_1),.clk(gclk));
	jdff dff_A_eF1kCpAo5_1(.dout(w_dff_A_7Wvx59Ze7_1),.din(w_dff_A_eF1kCpAo5_1),.clk(gclk));
	jdff dff_A_QMvxRlkL1_1(.dout(w_dff_A_eF1kCpAo5_1),.din(w_dff_A_QMvxRlkL1_1),.clk(gclk));
	jdff dff_A_WGJbEyxO9_1(.dout(w_dff_A_QMvxRlkL1_1),.din(w_dff_A_WGJbEyxO9_1),.clk(gclk));
	jdff dff_A_mVjjwKGe3_2(.dout(w_n843_1[2]),.din(w_dff_A_mVjjwKGe3_2),.clk(gclk));
	jdff dff_A_QV4le3QW2_2(.dout(w_dff_A_mVjjwKGe3_2),.din(w_dff_A_QV4le3QW2_2),.clk(gclk));
	jdff dff_A_OpxzFyJB1_2(.dout(w_dff_A_QV4le3QW2_2),.din(w_dff_A_OpxzFyJB1_2),.clk(gclk));
	jdff dff_A_77LzJhx87_2(.dout(w_dff_A_OpxzFyJB1_2),.din(w_dff_A_77LzJhx87_2),.clk(gclk));
	jdff dff_A_fTlAtfnV2_2(.dout(w_dff_A_77LzJhx87_2),.din(w_dff_A_fTlAtfnV2_2),.clk(gclk));
	jdff dff_A_XB4NSBmK9_2(.dout(w_dff_A_fTlAtfnV2_2),.din(w_dff_A_XB4NSBmK9_2),.clk(gclk));
	jdff dff_A_juotzPK26_2(.dout(w_dff_A_XB4NSBmK9_2),.din(w_dff_A_juotzPK26_2),.clk(gclk));
	jdff dff_A_IZVpXalT3_2(.dout(w_dff_A_juotzPK26_2),.din(w_dff_A_IZVpXalT3_2),.clk(gclk));
	jdff dff_A_xS6GkIMI7_2(.dout(w_dff_A_IZVpXalT3_2),.din(w_dff_A_xS6GkIMI7_2),.clk(gclk));
	jdff dff_A_Hwmo3KAh3_2(.dout(w_dff_A_xS6GkIMI7_2),.din(w_dff_A_Hwmo3KAh3_2),.clk(gclk));
	jdff dff_A_49N5uduP5_1(.dout(w_n843_0[1]),.din(w_dff_A_49N5uduP5_1),.clk(gclk));
	jdff dff_A_7HfHjDa84_1(.dout(w_dff_A_49N5uduP5_1),.din(w_dff_A_7HfHjDa84_1),.clk(gclk));
	jdff dff_A_HXCNTPbk8_1(.dout(w_dff_A_7HfHjDa84_1),.din(w_dff_A_HXCNTPbk8_1),.clk(gclk));
	jdff dff_A_cQmn4lFP1_1(.dout(w_dff_A_HXCNTPbk8_1),.din(w_dff_A_cQmn4lFP1_1),.clk(gclk));
	jdff dff_A_pNvcG4Z20_1(.dout(w_dff_A_cQmn4lFP1_1),.din(w_dff_A_pNvcG4Z20_1),.clk(gclk));
	jdff dff_A_yZz1gfvG6_1(.dout(w_dff_A_pNvcG4Z20_1),.din(w_dff_A_yZz1gfvG6_1),.clk(gclk));
	jdff dff_A_cv2rVsIN5_1(.dout(w_dff_A_yZz1gfvG6_1),.din(w_dff_A_cv2rVsIN5_1),.clk(gclk));
	jdff dff_A_4uWKlkDW5_1(.dout(w_dff_A_cv2rVsIN5_1),.din(w_dff_A_4uWKlkDW5_1),.clk(gclk));
	jdff dff_A_kPq7nZkf0_1(.dout(w_dff_A_4uWKlkDW5_1),.din(w_dff_A_kPq7nZkf0_1),.clk(gclk));
	jdff dff_A_oo9ebvOe3_1(.dout(w_dff_A_kPq7nZkf0_1),.din(w_dff_A_oo9ebvOe3_1),.clk(gclk));
	jdff dff_A_kk7zswMP6_1(.dout(w_dff_A_oo9ebvOe3_1),.din(w_dff_A_kk7zswMP6_1),.clk(gclk));
	jdff dff_A_ETtXIzyY5_2(.dout(w_n843_0[2]),.din(w_dff_A_ETtXIzyY5_2),.clk(gclk));
	jdff dff_B_HS0SdTZg8_3(.din(n843),.dout(w_dff_B_HS0SdTZg8_3),.clk(gclk));
	jdff dff_B_mhtNTZ0c1_3(.din(w_dff_B_HS0SdTZg8_3),.dout(w_dff_B_mhtNTZ0c1_3),.clk(gclk));
	jdff dff_B_TbCKI1Rc8_3(.din(w_dff_B_mhtNTZ0c1_3),.dout(w_dff_B_TbCKI1Rc8_3),.clk(gclk));
	jdff dff_B_E5kYmR2p0_3(.din(w_dff_B_TbCKI1Rc8_3),.dout(w_dff_B_E5kYmR2p0_3),.clk(gclk));
	jdff dff_B_QUibiwm78_3(.din(w_dff_B_E5kYmR2p0_3),.dout(w_dff_B_QUibiwm78_3),.clk(gclk));
	jdff dff_B_YNwcWui00_3(.din(w_dff_B_QUibiwm78_3),.dout(w_dff_B_YNwcWui00_3),.clk(gclk));
	jdff dff_A_lQRkkn7L6_1(.dout(w_n840_1[1]),.din(w_dff_A_lQRkkn7L6_1),.clk(gclk));
	jdff dff_A_A0rPgeOt2_1(.dout(w_dff_A_lQRkkn7L6_1),.din(w_dff_A_A0rPgeOt2_1),.clk(gclk));
	jdff dff_A_cVR335jI7_1(.dout(w_dff_A_A0rPgeOt2_1),.din(w_dff_A_cVR335jI7_1),.clk(gclk));
	jdff dff_A_ffNL8TsJ5_1(.dout(w_dff_A_cVR335jI7_1),.din(w_dff_A_ffNL8TsJ5_1),.clk(gclk));
	jdff dff_A_bxRoYoQg0_1(.dout(w_dff_A_ffNL8TsJ5_1),.din(w_dff_A_bxRoYoQg0_1),.clk(gclk));
	jdff dff_A_A4WVKjca8_1(.dout(w_dff_A_bxRoYoQg0_1),.din(w_dff_A_A4WVKjca8_1),.clk(gclk));
	jdff dff_A_8ZmzrnB93_1(.dout(w_dff_A_A4WVKjca8_1),.din(w_dff_A_8ZmzrnB93_1),.clk(gclk));
	jdff dff_A_trCIINZ53_1(.dout(w_dff_A_8ZmzrnB93_1),.din(w_dff_A_trCIINZ53_1),.clk(gclk));
	jdff dff_A_RmHbgeXA6_1(.dout(w_dff_A_trCIINZ53_1),.din(w_dff_A_RmHbgeXA6_1),.clk(gclk));
	jdff dff_A_muBslIKH4_1(.dout(w_dff_A_RmHbgeXA6_1),.din(w_dff_A_muBslIKH4_1),.clk(gclk));
	jdff dff_A_DU33Q8n40_1(.dout(w_dff_A_muBslIKH4_1),.din(w_dff_A_DU33Q8n40_1),.clk(gclk));
	jdff dff_A_kkTUnA3w1_1(.dout(w_dff_A_DU33Q8n40_1),.din(w_dff_A_kkTUnA3w1_1),.clk(gclk));
	jdff dff_A_u8b5jmpL2_1(.dout(w_dff_A_kkTUnA3w1_1),.din(w_dff_A_u8b5jmpL2_1),.clk(gclk));
	jdff dff_A_nLzfCQsM7_1(.dout(w_dff_A_u8b5jmpL2_1),.din(w_dff_A_nLzfCQsM7_1),.clk(gclk));
	jdff dff_A_VWpPITbl1_2(.dout(w_n840_1[2]),.din(w_dff_A_VWpPITbl1_2),.clk(gclk));
	jdff dff_A_VriCAyT59_2(.dout(w_dff_A_VWpPITbl1_2),.din(w_dff_A_VriCAyT59_2),.clk(gclk));
	jdff dff_A_9veWSEuW6_2(.dout(w_dff_A_VriCAyT59_2),.din(w_dff_A_9veWSEuW6_2),.clk(gclk));
	jdff dff_A_ESY4zw8P7_2(.dout(w_dff_A_9veWSEuW6_2),.din(w_dff_A_ESY4zw8P7_2),.clk(gclk));
	jdff dff_A_WrvQyqRj9_2(.dout(w_dff_A_ESY4zw8P7_2),.din(w_dff_A_WrvQyqRj9_2),.clk(gclk));
	jdff dff_A_34mx983w1_2(.dout(w_dff_A_WrvQyqRj9_2),.din(w_dff_A_34mx983w1_2),.clk(gclk));
	jdff dff_A_sj5abWxI0_2(.dout(w_dff_A_34mx983w1_2),.din(w_dff_A_sj5abWxI0_2),.clk(gclk));
	jdff dff_A_3ZL6epNk0_2(.dout(w_dff_A_sj5abWxI0_2),.din(w_dff_A_3ZL6epNk0_2),.clk(gclk));
	jdff dff_A_ETkTuboE4_2(.dout(w_dff_A_3ZL6epNk0_2),.din(w_dff_A_ETkTuboE4_2),.clk(gclk));
	jdff dff_A_8wZX448Z7_2(.dout(w_dff_A_ETkTuboE4_2),.din(w_dff_A_8wZX448Z7_2),.clk(gclk));
	jdff dff_A_xWdDvhNX3_1(.dout(w_n840_0[1]),.din(w_dff_A_xWdDvhNX3_1),.clk(gclk));
	jdff dff_A_sgeRwZNV6_1(.dout(w_dff_A_xWdDvhNX3_1),.din(w_dff_A_sgeRwZNV6_1),.clk(gclk));
	jdff dff_A_yd8p5ipB7_1(.dout(w_dff_A_sgeRwZNV6_1),.din(w_dff_A_yd8p5ipB7_1),.clk(gclk));
	jdff dff_A_TXkCGyfc9_1(.dout(w_dff_A_yd8p5ipB7_1),.din(w_dff_A_TXkCGyfc9_1),.clk(gclk));
	jdff dff_A_fbiWGzUq3_1(.dout(w_dff_A_TXkCGyfc9_1),.din(w_dff_A_fbiWGzUq3_1),.clk(gclk));
	jdff dff_A_1ysmOmuF8_1(.dout(w_dff_A_fbiWGzUq3_1),.din(w_dff_A_1ysmOmuF8_1),.clk(gclk));
	jdff dff_A_MNw5UL0q4_1(.dout(w_dff_A_1ysmOmuF8_1),.din(w_dff_A_MNw5UL0q4_1),.clk(gclk));
	jdff dff_A_XN9drVBE1_1(.dout(w_dff_A_MNw5UL0q4_1),.din(w_dff_A_XN9drVBE1_1),.clk(gclk));
	jdff dff_A_FOjqyKUo7_1(.dout(w_dff_A_XN9drVBE1_1),.din(w_dff_A_FOjqyKUo7_1),.clk(gclk));
	jdff dff_A_2QcyE6Bd0_1(.dout(w_dff_A_FOjqyKUo7_1),.din(w_dff_A_2QcyE6Bd0_1),.clk(gclk));
	jdff dff_A_Yw8dhu3K1_1(.dout(w_dff_A_2QcyE6Bd0_1),.din(w_dff_A_Yw8dhu3K1_1),.clk(gclk));
	jdff dff_A_MPqETHIJ7_2(.dout(w_n840_0[2]),.din(w_dff_A_MPqETHIJ7_2),.clk(gclk));
	jdff dff_A_MgUL0Bl02_2(.dout(w_dff_A_MPqETHIJ7_2),.din(w_dff_A_MgUL0Bl02_2),.clk(gclk));
	jdff dff_A_2s3zZm4n4_2(.dout(w_dff_A_MgUL0Bl02_2),.din(w_dff_A_2s3zZm4n4_2),.clk(gclk));
	jdff dff_A_1eiEKxGE0_2(.dout(w_dff_A_2s3zZm4n4_2),.din(w_dff_A_1eiEKxGE0_2),.clk(gclk));
	jdff dff_B_d13xtpX31_3(.din(n840),.dout(w_dff_B_d13xtpX31_3),.clk(gclk));
	jdff dff_B_46qk7RXw5_3(.din(w_dff_B_d13xtpX31_3),.dout(w_dff_B_46qk7RXw5_3),.clk(gclk));
	jdff dff_B_wGWUR7wr4_3(.din(w_dff_B_46qk7RXw5_3),.dout(w_dff_B_wGWUR7wr4_3),.clk(gclk));
	jdff dff_B_bByIaimR9_3(.din(w_dff_B_wGWUR7wr4_3),.dout(w_dff_B_bByIaimR9_3),.clk(gclk));
	jdff dff_B_7dhOLKPu5_3(.din(w_dff_B_bByIaimR9_3),.dout(w_dff_B_7dhOLKPu5_3),.clk(gclk));
	jdff dff_B_rXjKCc991_3(.din(w_dff_B_7dhOLKPu5_3),.dout(w_dff_B_rXjKCc991_3),.clk(gclk));
	jdff dff_B_ybEFOdHf6_3(.din(w_dff_B_rXjKCc991_3),.dout(w_dff_B_ybEFOdHf6_3),.clk(gclk));
	jdff dff_A_4CRskux41_1(.dout(w_G4090_0[1]),.din(w_dff_A_4CRskux41_1),.clk(gclk));
	jdff dff_A_SGVINllK6_2(.dout(w_G4089_0[2]),.din(w_dff_A_SGVINllK6_2),.clk(gclk));
	jdff dff_B_WDSJg6To0_1(.din(n1626),.dout(w_dff_B_WDSJg6To0_1),.clk(gclk));
	jdff dff_B_W0VuoQNR9_0(.din(n1637),.dout(w_dff_B_W0VuoQNR9_0),.clk(gclk));
	jdff dff_B_SJ2s7CJX8_0(.din(w_dff_B_W0VuoQNR9_0),.dout(w_dff_B_SJ2s7CJX8_0),.clk(gclk));
	jdff dff_B_H8iMtuMh1_0(.din(w_dff_B_SJ2s7CJX8_0),.dout(w_dff_B_H8iMtuMh1_0),.clk(gclk));
	jdff dff_B_0PYhF4O05_0(.din(w_dff_B_H8iMtuMh1_0),.dout(w_dff_B_0PYhF4O05_0),.clk(gclk));
	jdff dff_B_iEFiicFC9_0(.din(w_dff_B_0PYhF4O05_0),.dout(w_dff_B_iEFiicFC9_0),.clk(gclk));
	jdff dff_B_0qwySIf04_0(.din(w_dff_B_iEFiicFC9_0),.dout(w_dff_B_0qwySIf04_0),.clk(gclk));
	jdff dff_B_nODTLu8j8_0(.din(w_dff_B_0qwySIf04_0),.dout(w_dff_B_nODTLu8j8_0),.clk(gclk));
	jdff dff_B_hwZ2QBFM2_0(.din(w_dff_B_nODTLu8j8_0),.dout(w_dff_B_hwZ2QBFM2_0),.clk(gclk));
	jdff dff_B_cq9WxawO3_0(.din(w_dff_B_hwZ2QBFM2_0),.dout(w_dff_B_cq9WxawO3_0),.clk(gclk));
	jdff dff_B_guJLuw7V8_0(.din(w_dff_B_cq9WxawO3_0),.dout(w_dff_B_guJLuw7V8_0),.clk(gclk));
	jdff dff_B_ap0gar116_0(.din(w_dff_B_guJLuw7V8_0),.dout(w_dff_B_ap0gar116_0),.clk(gclk));
	jdff dff_B_ze3dQJQJ8_0(.din(w_dff_B_ap0gar116_0),.dout(w_dff_B_ze3dQJQJ8_0),.clk(gclk));
	jdff dff_B_N72LmPrQ6_0(.din(w_dff_B_ze3dQJQJ8_0),.dout(w_dff_B_N72LmPrQ6_0),.clk(gclk));
	jdff dff_B_MivFnubg2_0(.din(w_dff_B_N72LmPrQ6_0),.dout(w_dff_B_MivFnubg2_0),.clk(gclk));
	jdff dff_B_eEimXZ8n5_0(.din(w_dff_B_MivFnubg2_0),.dout(w_dff_B_eEimXZ8n5_0),.clk(gclk));
	jdff dff_B_8hT4PvgW8_0(.din(w_dff_B_eEimXZ8n5_0),.dout(w_dff_B_8hT4PvgW8_0),.clk(gclk));
	jdff dff_B_vLSC3Jhc8_0(.din(w_dff_B_8hT4PvgW8_0),.dout(w_dff_B_vLSC3Jhc8_0),.clk(gclk));
	jdff dff_B_0HFVwDKA1_0(.din(w_dff_B_vLSC3Jhc8_0),.dout(w_dff_B_0HFVwDKA1_0),.clk(gclk));
	jdff dff_B_fNWvu0Ba5_1(.din(n1633),.dout(w_dff_B_fNWvu0Ba5_1),.clk(gclk));
	jdff dff_B_Y8Kz8GFj8_1(.din(n1627),.dout(w_dff_B_Y8Kz8GFj8_1),.clk(gclk));
	jdff dff_B_SycmWz7h0_1(.din(w_dff_B_Y8Kz8GFj8_1),.dout(w_dff_B_SycmWz7h0_1),.clk(gclk));
	jdff dff_B_77Z1O1pc6_1(.din(w_dff_B_SycmWz7h0_1),.dout(w_dff_B_77Z1O1pc6_1),.clk(gclk));
	jdff dff_B_SLkzalUW6_1(.din(w_dff_B_77Z1O1pc6_1),.dout(w_dff_B_SLkzalUW6_1),.clk(gclk));
	jdff dff_B_WmxQRnwC7_1(.din(w_dff_B_SLkzalUW6_1),.dout(w_dff_B_WmxQRnwC7_1),.clk(gclk));
	jdff dff_B_Mq51PVmM5_1(.din(w_dff_B_WmxQRnwC7_1),.dout(w_dff_B_Mq51PVmM5_1),.clk(gclk));
	jdff dff_B_SHf0hWt57_1(.din(w_dff_B_Mq51PVmM5_1),.dout(w_dff_B_SHf0hWt57_1),.clk(gclk));
	jdff dff_B_4eLVmgno8_1(.din(w_dff_B_SHf0hWt57_1),.dout(w_dff_B_4eLVmgno8_1),.clk(gclk));
	jdff dff_B_ZJJK44hD6_1(.din(w_dff_B_4eLVmgno8_1),.dout(w_dff_B_ZJJK44hD6_1),.clk(gclk));
	jdff dff_B_OZcxFgxD3_1(.din(w_dff_B_ZJJK44hD6_1),.dout(w_dff_B_OZcxFgxD3_1),.clk(gclk));
	jdff dff_B_S8tdATFH8_1(.din(w_dff_B_OZcxFgxD3_1),.dout(w_dff_B_S8tdATFH8_1),.clk(gclk));
	jdff dff_B_RE3od9HI0_1(.din(w_dff_B_S8tdATFH8_1),.dout(w_dff_B_RE3od9HI0_1),.clk(gclk));
	jdff dff_B_ipm9Ljwo2_1(.din(w_dff_B_RE3od9HI0_1),.dout(w_dff_B_ipm9Ljwo2_1),.clk(gclk));
	jdff dff_B_pq6E21WS5_1(.din(w_dff_B_ipm9Ljwo2_1),.dout(w_dff_B_pq6E21WS5_1),.clk(gclk));
	jdff dff_B_SZKGjNZO4_1(.din(w_dff_B_pq6E21WS5_1),.dout(w_dff_B_SZKGjNZO4_1),.clk(gclk));
	jdff dff_B_f9O6MNGd0_1(.din(w_dff_B_SZKGjNZO4_1),.dout(w_dff_B_f9O6MNGd0_1),.clk(gclk));
	jdff dff_B_Y58RtSJ29_1(.din(w_dff_B_f9O6MNGd0_1),.dout(w_dff_B_Y58RtSJ29_1),.clk(gclk));
	jdff dff_B_wotfyTJE5_1(.din(w_dff_B_Y58RtSJ29_1),.dout(w_dff_B_wotfyTJE5_1),.clk(gclk));
	jdff dff_B_lU0gpBps2_1(.din(w_dff_B_wotfyTJE5_1),.dout(w_dff_B_lU0gpBps2_1),.clk(gclk));
	jdff dff_A_iHELKUG08_0(.dout(w_n988_1[0]),.din(w_dff_A_iHELKUG08_0),.clk(gclk));
	jdff dff_A_JLMDq7te7_0(.dout(w_dff_A_iHELKUG08_0),.din(w_dff_A_JLMDq7te7_0),.clk(gclk));
	jdff dff_A_XlXlueqR2_0(.dout(w_dff_A_JLMDq7te7_0),.din(w_dff_A_XlXlueqR2_0),.clk(gclk));
	jdff dff_A_C65bxzey1_0(.dout(w_dff_A_XlXlueqR2_0),.din(w_dff_A_C65bxzey1_0),.clk(gclk));
	jdff dff_A_jwdxQDeC6_0(.dout(w_dff_A_C65bxzey1_0),.din(w_dff_A_jwdxQDeC6_0),.clk(gclk));
	jdff dff_A_RS3E63ZZ8_0(.dout(w_dff_A_jwdxQDeC6_0),.din(w_dff_A_RS3E63ZZ8_0),.clk(gclk));
	jdff dff_A_zaEMJS5y1_2(.dout(w_n988_1[2]),.din(w_dff_A_zaEMJS5y1_2),.clk(gclk));
	jdff dff_A_f1Ac9L4z1_2(.dout(w_dff_A_zaEMJS5y1_2),.din(w_dff_A_f1Ac9L4z1_2),.clk(gclk));
	jdff dff_A_4Q7Rqo8r2_2(.dout(w_dff_A_f1Ac9L4z1_2),.din(w_dff_A_4Q7Rqo8r2_2),.clk(gclk));
	jdff dff_A_5S8BuSF53_2(.dout(w_dff_A_4Q7Rqo8r2_2),.din(w_dff_A_5S8BuSF53_2),.clk(gclk));
	jdff dff_A_n2SQzVNL3_2(.dout(w_dff_A_5S8BuSF53_2),.din(w_dff_A_n2SQzVNL3_2),.clk(gclk));
	jdff dff_A_KeYBZipT4_2(.dout(w_dff_A_n2SQzVNL3_2),.din(w_dff_A_KeYBZipT4_2),.clk(gclk));
	jdff dff_A_RMdziKXA7_2(.dout(w_dff_A_KeYBZipT4_2),.din(w_dff_A_RMdziKXA7_2),.clk(gclk));
	jdff dff_A_xs8At4Ad5_2(.dout(w_dff_A_RMdziKXA7_2),.din(w_dff_A_xs8At4Ad5_2),.clk(gclk));
	jdff dff_A_ssuHvV1x9_2(.dout(w_dff_A_xs8At4Ad5_2),.din(w_dff_A_ssuHvV1x9_2),.clk(gclk));
	jdff dff_A_YEuyJf9P2_2(.dout(w_dff_A_ssuHvV1x9_2),.din(w_dff_A_YEuyJf9P2_2),.clk(gclk));
	jdff dff_A_eZyDpLQi3_2(.dout(w_dff_A_YEuyJf9P2_2),.din(w_dff_A_eZyDpLQi3_2),.clk(gclk));
	jdff dff_A_3d2wZlUO0_2(.dout(w_dff_A_eZyDpLQi3_2),.din(w_dff_A_3d2wZlUO0_2),.clk(gclk));
	jdff dff_A_XBNuIOju5_2(.dout(w_dff_A_3d2wZlUO0_2),.din(w_dff_A_XBNuIOju5_2),.clk(gclk));
	jdff dff_A_wXEszY9E9_2(.dout(w_dff_A_XBNuIOju5_2),.din(w_dff_A_wXEszY9E9_2),.clk(gclk));
	jdff dff_A_Y4SC1a0I0_2(.dout(w_dff_A_wXEszY9E9_2),.din(w_dff_A_Y4SC1a0I0_2),.clk(gclk));
	jdff dff_A_QLIc4odz2_2(.dout(w_dff_A_Y4SC1a0I0_2),.din(w_dff_A_QLIc4odz2_2),.clk(gclk));
	jdff dff_A_IkYQX1ya8_2(.dout(w_dff_A_QLIc4odz2_2),.din(w_dff_A_IkYQX1ya8_2),.clk(gclk));
	jdff dff_A_WcX8CP5O4_2(.dout(w_dff_A_IkYQX1ya8_2),.din(w_dff_A_WcX8CP5O4_2),.clk(gclk));
	jdff dff_A_eXFg4IlW1_1(.dout(w_n988_0[1]),.din(w_dff_A_eXFg4IlW1_1),.clk(gclk));
	jdff dff_A_ScsDh4u38_1(.dout(w_dff_A_eXFg4IlW1_1),.din(w_dff_A_ScsDh4u38_1),.clk(gclk));
	jdff dff_A_xhc8N4CO3_1(.dout(w_dff_A_ScsDh4u38_1),.din(w_dff_A_xhc8N4CO3_1),.clk(gclk));
	jdff dff_A_V8lgoi8O3_1(.dout(w_dff_A_xhc8N4CO3_1),.din(w_dff_A_V8lgoi8O3_1),.clk(gclk));
	jdff dff_A_rqzMa1as8_1(.dout(w_dff_A_V8lgoi8O3_1),.din(w_dff_A_rqzMa1as8_1),.clk(gclk));
	jdff dff_A_vKmt0qfj2_1(.dout(w_dff_A_rqzMa1as8_1),.din(w_dff_A_vKmt0qfj2_1),.clk(gclk));
	jdff dff_A_SBDi12mP8_1(.dout(w_dff_A_vKmt0qfj2_1),.din(w_dff_A_SBDi12mP8_1),.clk(gclk));
	jdff dff_A_0n4bZYXa1_1(.dout(w_dff_A_SBDi12mP8_1),.din(w_dff_A_0n4bZYXa1_1),.clk(gclk));
	jdff dff_A_wQW1a9xD2_1(.dout(w_dff_A_0n4bZYXa1_1),.din(w_dff_A_wQW1a9xD2_1),.clk(gclk));
	jdff dff_A_gu81xreD1_1(.dout(w_dff_A_wQW1a9xD2_1),.din(w_dff_A_gu81xreD1_1),.clk(gclk));
	jdff dff_A_OxxtIKWa9_1(.dout(w_dff_A_gu81xreD1_1),.din(w_dff_A_OxxtIKWa9_1),.clk(gclk));
	jdff dff_A_3Vgv66q52_1(.dout(w_dff_A_OxxtIKWa9_1),.din(w_dff_A_3Vgv66q52_1),.clk(gclk));
	jdff dff_A_qB07bLz41_1(.dout(w_dff_A_3Vgv66q52_1),.din(w_dff_A_qB07bLz41_1),.clk(gclk));
	jdff dff_A_JNnxzt9i4_1(.dout(w_dff_A_qB07bLz41_1),.din(w_dff_A_JNnxzt9i4_1),.clk(gclk));
	jdff dff_A_SnYGJwgI1_1(.dout(w_dff_A_JNnxzt9i4_1),.din(w_dff_A_SnYGJwgI1_1),.clk(gclk));
	jdff dff_A_q74Muz0Z9_1(.dout(w_dff_A_SnYGJwgI1_1),.din(w_dff_A_q74Muz0Z9_1),.clk(gclk));
	jdff dff_A_FmQcAuyX1_2(.dout(w_n988_0[2]),.din(w_dff_A_FmQcAuyX1_2),.clk(gclk));
	jdff dff_A_bVDZBFzy6_2(.dout(w_dff_A_FmQcAuyX1_2),.din(w_dff_A_bVDZBFzy6_2),.clk(gclk));
	jdff dff_A_BJg2IT4b6_2(.dout(w_dff_A_bVDZBFzy6_2),.din(w_dff_A_BJg2IT4b6_2),.clk(gclk));
	jdff dff_A_PMsPWmz07_2(.dout(w_dff_A_BJg2IT4b6_2),.din(w_dff_A_PMsPWmz07_2),.clk(gclk));
	jdff dff_A_JVDka3Zi9_2(.dout(w_dff_A_PMsPWmz07_2),.din(w_dff_A_JVDka3Zi9_2),.clk(gclk));
	jdff dff_A_pmBhRDCS4_2(.dout(w_dff_A_JVDka3Zi9_2),.din(w_dff_A_pmBhRDCS4_2),.clk(gclk));
	jdff dff_A_srwLQ5c40_2(.dout(w_dff_A_pmBhRDCS4_2),.din(w_dff_A_srwLQ5c40_2),.clk(gclk));
	jdff dff_B_ADl4x1I67_1(.din(n1625),.dout(w_dff_B_ADl4x1I67_1),.clk(gclk));
	jdff dff_B_YIkN63ix3_1(.din(w_dff_B_ADl4x1I67_1),.dout(w_dff_B_YIkN63ix3_1),.clk(gclk));
	jdff dff_B_02i94erj1_1(.din(w_dff_B_YIkN63ix3_1),.dout(w_dff_B_02i94erj1_1),.clk(gclk));
	jdff dff_B_1RqGvp9P5_1(.din(w_dff_B_02i94erj1_1),.dout(w_dff_B_1RqGvp9P5_1),.clk(gclk));
	jdff dff_B_0ZkJsJOg0_1(.din(w_dff_B_1RqGvp9P5_1),.dout(w_dff_B_0ZkJsJOg0_1),.clk(gclk));
	jdff dff_B_xbZwIeDv3_1(.din(w_dff_B_0ZkJsJOg0_1),.dout(w_dff_B_xbZwIeDv3_1),.clk(gclk));
	jdff dff_B_CCf1sQqX0_1(.din(w_dff_B_xbZwIeDv3_1),.dout(w_dff_B_CCf1sQqX0_1),.clk(gclk));
	jdff dff_B_7i3JhJil5_1(.din(w_dff_B_CCf1sQqX0_1),.dout(w_dff_B_7i3JhJil5_1),.clk(gclk));
	jdff dff_B_WdTnOeSQ7_1(.din(w_dff_B_7i3JhJil5_1),.dout(w_dff_B_WdTnOeSQ7_1),.clk(gclk));
	jdff dff_B_ZILFCqnK7_1(.din(w_dff_B_WdTnOeSQ7_1),.dout(w_dff_B_ZILFCqnK7_1),.clk(gclk));
	jdff dff_B_s0jOnRZr4_1(.din(w_dff_B_ZILFCqnK7_1),.dout(w_dff_B_s0jOnRZr4_1),.clk(gclk));
	jdff dff_B_T0AZJEkz9_1(.din(w_dff_B_s0jOnRZr4_1),.dout(w_dff_B_T0AZJEkz9_1),.clk(gclk));
	jdff dff_B_H9PfolCh3_1(.din(w_dff_B_T0AZJEkz9_1),.dout(w_dff_B_H9PfolCh3_1),.clk(gclk));
	jdff dff_B_IFzlGp5n3_1(.din(w_dff_B_H9PfolCh3_1),.dout(w_dff_B_IFzlGp5n3_1),.clk(gclk));
	jdff dff_B_4dMFw2le9_1(.din(w_dff_B_IFzlGp5n3_1),.dout(w_dff_B_4dMFw2le9_1),.clk(gclk));
	jdff dff_B_N973HRmS5_1(.din(w_dff_B_4dMFw2le9_1),.dout(w_dff_B_N973HRmS5_1),.clk(gclk));
	jdff dff_B_gag6sJdH4_1(.din(w_dff_B_N973HRmS5_1),.dout(w_dff_B_gag6sJdH4_1),.clk(gclk));
	jdff dff_B_ZhBvSANF8_1(.din(w_dff_B_gag6sJdH4_1),.dout(w_dff_B_ZhBvSANF8_1),.clk(gclk));
	jdff dff_B_2TT89mhw0_1(.din(w_dff_B_ZhBvSANF8_1),.dout(w_dff_B_2TT89mhw0_1),.clk(gclk));
	jdff dff_A_KaS8Gjmp7_0(.dout(w_n985_1[0]),.din(w_dff_A_KaS8Gjmp7_0),.clk(gclk));
	jdff dff_A_YDSjYdWi1_0(.dout(w_dff_A_KaS8Gjmp7_0),.din(w_dff_A_YDSjYdWi1_0),.clk(gclk));
	jdff dff_A_6sNleYyk2_0(.dout(w_dff_A_YDSjYdWi1_0),.din(w_dff_A_6sNleYyk2_0),.clk(gclk));
	jdff dff_A_QeuITl8g9_0(.dout(w_dff_A_6sNleYyk2_0),.din(w_dff_A_QeuITl8g9_0),.clk(gclk));
	jdff dff_A_uopNGU9Q9_0(.dout(w_dff_A_QeuITl8g9_0),.din(w_dff_A_uopNGU9Q9_0),.clk(gclk));
	jdff dff_A_A64mu9WC9_0(.dout(w_dff_A_uopNGU9Q9_0),.din(w_dff_A_A64mu9WC9_0),.clk(gclk));
	jdff dff_A_Nky4KSlY5_0(.dout(w_dff_A_A64mu9WC9_0),.din(w_dff_A_Nky4KSlY5_0),.clk(gclk));
	jdff dff_A_YXbuRvEe6_2(.dout(w_n985_1[2]),.din(w_dff_A_YXbuRvEe6_2),.clk(gclk));
	jdff dff_A_E8b3whZb0_2(.dout(w_dff_A_YXbuRvEe6_2),.din(w_dff_A_E8b3whZb0_2),.clk(gclk));
	jdff dff_A_Z6sV74iU8_2(.dout(w_dff_A_E8b3whZb0_2),.din(w_dff_A_Z6sV74iU8_2),.clk(gclk));
	jdff dff_A_ygwnds2u5_2(.dout(w_dff_A_Z6sV74iU8_2),.din(w_dff_A_ygwnds2u5_2),.clk(gclk));
	jdff dff_A_BkgepQIr4_2(.dout(w_dff_A_ygwnds2u5_2),.din(w_dff_A_BkgepQIr4_2),.clk(gclk));
	jdff dff_A_EDUFbXmI6_2(.dout(w_dff_A_BkgepQIr4_2),.din(w_dff_A_EDUFbXmI6_2),.clk(gclk));
	jdff dff_A_Fqya9Ppc7_2(.dout(w_dff_A_EDUFbXmI6_2),.din(w_dff_A_Fqya9Ppc7_2),.clk(gclk));
	jdff dff_A_bvgAqDQA7_2(.dout(w_dff_A_Fqya9Ppc7_2),.din(w_dff_A_bvgAqDQA7_2),.clk(gclk));
	jdff dff_A_yYPMmlIl2_2(.dout(w_dff_A_bvgAqDQA7_2),.din(w_dff_A_yYPMmlIl2_2),.clk(gclk));
	jdff dff_A_Yp2IxehB0_2(.dout(w_dff_A_yYPMmlIl2_2),.din(w_dff_A_Yp2IxehB0_2),.clk(gclk));
	jdff dff_A_Gi0yjUwF7_2(.dout(w_dff_A_Yp2IxehB0_2),.din(w_dff_A_Gi0yjUwF7_2),.clk(gclk));
	jdff dff_A_7LVqeWkA3_2(.dout(w_dff_A_Gi0yjUwF7_2),.din(w_dff_A_7LVqeWkA3_2),.clk(gclk));
	jdff dff_A_OsZUJQAV4_2(.dout(w_dff_A_7LVqeWkA3_2),.din(w_dff_A_OsZUJQAV4_2),.clk(gclk));
	jdff dff_A_Vf9Gdczv3_2(.dout(w_dff_A_OsZUJQAV4_2),.din(w_dff_A_Vf9Gdczv3_2),.clk(gclk));
	jdff dff_A_LHry1Kob6_2(.dout(w_dff_A_Vf9Gdczv3_2),.din(w_dff_A_LHry1Kob6_2),.clk(gclk));
	jdff dff_A_yj4xZaDO9_2(.dout(w_dff_A_LHry1Kob6_2),.din(w_dff_A_yj4xZaDO9_2),.clk(gclk));
	jdff dff_A_qDdl9PUa3_2(.dout(w_dff_A_yj4xZaDO9_2),.din(w_dff_A_qDdl9PUa3_2),.clk(gclk));
	jdff dff_A_Gx3srTJB5_2(.dout(w_dff_A_qDdl9PUa3_2),.din(w_dff_A_Gx3srTJB5_2),.clk(gclk));
	jdff dff_A_9vZJQ24L1_2(.dout(w_dff_A_Gx3srTJB5_2),.din(w_dff_A_9vZJQ24L1_2),.clk(gclk));
	jdff dff_A_SzmOzkWV1_1(.dout(w_n985_0[1]),.din(w_dff_A_SzmOzkWV1_1),.clk(gclk));
	jdff dff_A_EawolTbo1_1(.dout(w_dff_A_SzmOzkWV1_1),.din(w_dff_A_EawolTbo1_1),.clk(gclk));
	jdff dff_A_c5kw5qj53_1(.dout(w_dff_A_EawolTbo1_1),.din(w_dff_A_c5kw5qj53_1),.clk(gclk));
	jdff dff_A_CySUXMTS8_1(.dout(w_dff_A_c5kw5qj53_1),.din(w_dff_A_CySUXMTS8_1),.clk(gclk));
	jdff dff_A_0FhMjHqI6_1(.dout(w_dff_A_CySUXMTS8_1),.din(w_dff_A_0FhMjHqI6_1),.clk(gclk));
	jdff dff_A_VUbQvf5T2_1(.dout(w_dff_A_0FhMjHqI6_1),.din(w_dff_A_VUbQvf5T2_1),.clk(gclk));
	jdff dff_A_KRZJpQur7_1(.dout(w_dff_A_VUbQvf5T2_1),.din(w_dff_A_KRZJpQur7_1),.clk(gclk));
	jdff dff_A_VewggG2H4_1(.dout(w_dff_A_KRZJpQur7_1),.din(w_dff_A_VewggG2H4_1),.clk(gclk));
	jdff dff_A_6QfcUjhk5_1(.dout(w_dff_A_VewggG2H4_1),.din(w_dff_A_6QfcUjhk5_1),.clk(gclk));
	jdff dff_A_qno6efzJ4_1(.dout(w_dff_A_6QfcUjhk5_1),.din(w_dff_A_qno6efzJ4_1),.clk(gclk));
	jdff dff_A_foLlheHq1_1(.dout(w_dff_A_qno6efzJ4_1),.din(w_dff_A_foLlheHq1_1),.clk(gclk));
	jdff dff_A_QOzIT3WG2_1(.dout(w_dff_A_foLlheHq1_1),.din(w_dff_A_QOzIT3WG2_1),.clk(gclk));
	jdff dff_A_DSCTJOUl1_1(.dout(w_dff_A_QOzIT3WG2_1),.din(w_dff_A_DSCTJOUl1_1),.clk(gclk));
	jdff dff_A_uKVMB4oG5_1(.dout(w_dff_A_DSCTJOUl1_1),.din(w_dff_A_uKVMB4oG5_1),.clk(gclk));
	jdff dff_A_4G2HRrGl2_1(.dout(w_dff_A_uKVMB4oG5_1),.din(w_dff_A_4G2HRrGl2_1),.clk(gclk));
	jdff dff_A_EoNtu0H00_1(.dout(w_dff_A_4G2HRrGl2_1),.din(w_dff_A_EoNtu0H00_1),.clk(gclk));
	jdff dff_A_RFQeJ0rj8_1(.dout(w_dff_A_EoNtu0H00_1),.din(w_dff_A_RFQeJ0rj8_1),.clk(gclk));
	jdff dff_A_MN9hvVqO9_2(.dout(w_n985_0[2]),.din(w_dff_A_MN9hvVqO9_2),.clk(gclk));
	jdff dff_A_zY7AvL4P7_2(.dout(w_dff_A_MN9hvVqO9_2),.din(w_dff_A_zY7AvL4P7_2),.clk(gclk));
	jdff dff_A_5tARJulS1_2(.dout(w_dff_A_zY7AvL4P7_2),.din(w_dff_A_5tARJulS1_2),.clk(gclk));
	jdff dff_A_iqPyKJ4v2_2(.dout(w_dff_A_5tARJulS1_2),.din(w_dff_A_iqPyKJ4v2_2),.clk(gclk));
	jdff dff_A_HPm1gUJ59_2(.dout(w_dff_A_iqPyKJ4v2_2),.din(w_dff_A_HPm1gUJ59_2),.clk(gclk));
	jdff dff_A_DF7xBQUR0_2(.dout(w_dff_A_HPm1gUJ59_2),.din(w_dff_A_DF7xBQUR0_2),.clk(gclk));
	jdff dff_A_KtPzDrIM2_2(.dout(w_dff_A_DF7xBQUR0_2),.din(w_dff_A_KtPzDrIM2_2),.clk(gclk));
	jdff dff_A_dwSHW1VY7_2(.dout(w_dff_A_KtPzDrIM2_2),.din(w_dff_A_dwSHW1VY7_2),.clk(gclk));
	jdff dff_A_TZqrMTYV7_2(.dout(w_dff_A_dwSHW1VY7_2),.din(w_dff_A_TZqrMTYV7_2),.clk(gclk));
	jdff dff_A_nShUj1GO1_2(.dout(w_dff_A_TZqrMTYV7_2),.din(w_dff_A_nShUj1GO1_2),.clk(gclk));
	jdff dff_A_XlHVV9RA6_2(.dout(w_dff_A_nShUj1GO1_2),.din(w_dff_A_XlHVV9RA6_2),.clk(gclk));
	jdff dff_A_kWN7fJzX1_1(.dout(w_G1690_0[1]),.din(w_dff_A_kWN7fJzX1_1),.clk(gclk));
	jdff dff_A_shACUS9a7_2(.dout(w_G1689_0[2]),.din(w_dff_A_shACUS9a7_2),.clk(gclk));
	jdff dff_B_kO1xlF5h5_1(.din(n1642),.dout(w_dff_B_kO1xlF5h5_1),.clk(gclk));
	jdff dff_B_LfIV5xTx3_0(.din(n1649),.dout(w_dff_B_LfIV5xTx3_0),.clk(gclk));
	jdff dff_B_UiMih9lw6_0(.din(w_dff_B_LfIV5xTx3_0),.dout(w_dff_B_UiMih9lw6_0),.clk(gclk));
	jdff dff_B_bmXPNjKx8_0(.din(w_dff_B_UiMih9lw6_0),.dout(w_dff_B_bmXPNjKx8_0),.clk(gclk));
	jdff dff_B_0XCAjgoC6_0(.din(w_dff_B_bmXPNjKx8_0),.dout(w_dff_B_0XCAjgoC6_0),.clk(gclk));
	jdff dff_B_7mLXmI0j0_0(.din(w_dff_B_0XCAjgoC6_0),.dout(w_dff_B_7mLXmI0j0_0),.clk(gclk));
	jdff dff_B_zibivfLm9_0(.din(w_dff_B_7mLXmI0j0_0),.dout(w_dff_B_zibivfLm9_0),.clk(gclk));
	jdff dff_B_rDNdzLCw9_0(.din(w_dff_B_zibivfLm9_0),.dout(w_dff_B_rDNdzLCw9_0),.clk(gclk));
	jdff dff_B_aCpFc6yW1_0(.din(w_dff_B_rDNdzLCw9_0),.dout(w_dff_B_aCpFc6yW1_0),.clk(gclk));
	jdff dff_B_xG6T76pF6_0(.din(w_dff_B_aCpFc6yW1_0),.dout(w_dff_B_xG6T76pF6_0),.clk(gclk));
	jdff dff_B_6ARhtCrO9_0(.din(w_dff_B_xG6T76pF6_0),.dout(w_dff_B_6ARhtCrO9_0),.clk(gclk));
	jdff dff_B_nLYEia8J2_0(.din(w_dff_B_6ARhtCrO9_0),.dout(w_dff_B_nLYEia8J2_0),.clk(gclk));
	jdff dff_B_sMYYjckc0_0(.din(w_dff_B_nLYEia8J2_0),.dout(w_dff_B_sMYYjckc0_0),.clk(gclk));
	jdff dff_B_lpK4u32E2_0(.din(w_dff_B_sMYYjckc0_0),.dout(w_dff_B_lpK4u32E2_0),.clk(gclk));
	jdff dff_B_Q6TBJCfg7_0(.din(w_dff_B_lpK4u32E2_0),.dout(w_dff_B_Q6TBJCfg7_0),.clk(gclk));
	jdff dff_B_DenSSNA57_0(.din(w_dff_B_Q6TBJCfg7_0),.dout(w_dff_B_DenSSNA57_0),.clk(gclk));
	jdff dff_B_i1VLYggP1_0(.din(w_dff_B_DenSSNA57_0),.dout(w_dff_B_i1VLYggP1_0),.clk(gclk));
	jdff dff_B_7zETgrhx6_0(.din(w_dff_B_i1VLYggP1_0),.dout(w_dff_B_7zETgrhx6_0),.clk(gclk));
	jdff dff_B_sUjayH6W6_0(.din(w_dff_B_7zETgrhx6_0),.dout(w_dff_B_sUjayH6W6_0),.clk(gclk));
	jdff dff_B_pjxcf6tk2_1(.din(n1646),.dout(w_dff_B_pjxcf6tk2_1),.clk(gclk));
	jdff dff_B_fnBqcRVL1_2(.din(n1634),.dout(w_dff_B_fnBqcRVL1_2),.clk(gclk));
	jdff dff_B_9ka1Ae2n2_2(.din(w_dff_B_fnBqcRVL1_2),.dout(w_dff_B_9ka1Ae2n2_2),.clk(gclk));
	jdff dff_B_uXGqDPoi2_2(.din(n1631),.dout(w_dff_B_uXGqDPoi2_2),.clk(gclk));
	jdff dff_B_5nRWFFqr8_1(.din(n1643),.dout(w_dff_B_5nRWFFqr8_1),.clk(gclk));
	jdff dff_B_BSIomkER9_1(.din(w_dff_B_5nRWFFqr8_1),.dout(w_dff_B_BSIomkER9_1),.clk(gclk));
	jdff dff_B_mRgcY9Nb7_1(.din(w_dff_B_BSIomkER9_1),.dout(w_dff_B_mRgcY9Nb7_1),.clk(gclk));
	jdff dff_B_nCoNP1I53_1(.din(w_dff_B_mRgcY9Nb7_1),.dout(w_dff_B_nCoNP1I53_1),.clk(gclk));
	jdff dff_B_jSEeUeMY0_1(.din(w_dff_B_nCoNP1I53_1),.dout(w_dff_B_jSEeUeMY0_1),.clk(gclk));
	jdff dff_B_DNB5IOhH3_1(.din(w_dff_B_jSEeUeMY0_1),.dout(w_dff_B_DNB5IOhH3_1),.clk(gclk));
	jdff dff_B_jcYqNVaM4_1(.din(w_dff_B_DNB5IOhH3_1),.dout(w_dff_B_jcYqNVaM4_1),.clk(gclk));
	jdff dff_B_bsWaEmUV7_1(.din(w_dff_B_jcYqNVaM4_1),.dout(w_dff_B_bsWaEmUV7_1),.clk(gclk));
	jdff dff_B_nvfFrwUp2_1(.din(w_dff_B_bsWaEmUV7_1),.dout(w_dff_B_nvfFrwUp2_1),.clk(gclk));
	jdff dff_B_oQwCSowM1_1(.din(w_dff_B_nvfFrwUp2_1),.dout(w_dff_B_oQwCSowM1_1),.clk(gclk));
	jdff dff_B_H4yjJnyj3_1(.din(w_dff_B_oQwCSowM1_1),.dout(w_dff_B_H4yjJnyj3_1),.clk(gclk));
	jdff dff_B_q7zrlhNy5_1(.din(w_dff_B_H4yjJnyj3_1),.dout(w_dff_B_q7zrlhNy5_1),.clk(gclk));
	jdff dff_B_IYsRfYYL9_1(.din(w_dff_B_q7zrlhNy5_1),.dout(w_dff_B_IYsRfYYL9_1),.clk(gclk));
	jdff dff_B_GTWJnPbN0_1(.din(w_dff_B_IYsRfYYL9_1),.dout(w_dff_B_GTWJnPbN0_1),.clk(gclk));
	jdff dff_B_3YKgXkRR4_1(.din(w_dff_B_GTWJnPbN0_1),.dout(w_dff_B_3YKgXkRR4_1),.clk(gclk));
	jdff dff_B_whtlgsNr0_1(.din(w_dff_B_3YKgXkRR4_1),.dout(w_dff_B_whtlgsNr0_1),.clk(gclk));
	jdff dff_B_iOwKKTv57_1(.din(w_dff_B_whtlgsNr0_1),.dout(w_dff_B_iOwKKTv57_1),.clk(gclk));
	jdff dff_B_Gt6abUR49_1(.din(w_dff_B_iOwKKTv57_1),.dout(w_dff_B_Gt6abUR49_1),.clk(gclk));
	jdff dff_B_QQQYwGwz9_1(.din(w_dff_B_Gt6abUR49_1),.dout(w_dff_B_QQQYwGwz9_1),.clk(gclk));
	jdff dff_B_nSyVskDI9_0(.din(n1628),.dout(w_dff_B_nSyVskDI9_0),.clk(gclk));
	jdff dff_B_8wF03YzM8_0(.din(w_dff_B_nSyVskDI9_0),.dout(w_dff_B_8wF03YzM8_0),.clk(gclk));
	jdff dff_B_aPuqufsa5_0(.din(w_dff_B_8wF03YzM8_0),.dout(w_dff_B_aPuqufsa5_0),.clk(gclk));
	jdff dff_B_8VUeNZon6_0(.din(w_dff_B_aPuqufsa5_0),.dout(w_dff_B_8VUeNZon6_0),.clk(gclk));
	jdff dff_B_yHoVVJiQ8_0(.din(w_dff_B_8VUeNZon6_0),.dout(w_dff_B_yHoVVJiQ8_0),.clk(gclk));
	jdff dff_B_WfVGL2fU4_0(.din(w_dff_B_yHoVVJiQ8_0),.dout(w_dff_B_WfVGL2fU4_0),.clk(gclk));
	jdff dff_B_GY4ZbLlM0_0(.din(w_dff_B_WfVGL2fU4_0),.dout(w_dff_B_GY4ZbLlM0_0),.clk(gclk));
	jdff dff_B_ITN3cMfV3_0(.din(w_dff_B_GY4ZbLlM0_0),.dout(w_dff_B_ITN3cMfV3_0),.clk(gclk));
	jdff dff_B_HrHYRHr98_0(.din(w_dff_B_ITN3cMfV3_0),.dout(w_dff_B_HrHYRHr98_0),.clk(gclk));
	jdff dff_B_cBe28yCV4_0(.din(w_dff_B_HrHYRHr98_0),.dout(w_dff_B_cBe28yCV4_0),.clk(gclk));
	jdff dff_B_XUgYyT8M9_0(.din(w_dff_B_cBe28yCV4_0),.dout(w_dff_B_XUgYyT8M9_0),.clk(gclk));
	jdff dff_B_R9gTmzsv8_0(.din(w_dff_B_XUgYyT8M9_0),.dout(w_dff_B_R9gTmzsv8_0),.clk(gclk));
	jdff dff_B_AWCXUrGL8_0(.din(w_dff_B_R9gTmzsv8_0),.dout(w_dff_B_AWCXUrGL8_0),.clk(gclk));
	jdff dff_B_zvaA5D1N9_0(.din(w_dff_B_AWCXUrGL8_0),.dout(w_dff_B_zvaA5D1N9_0),.clk(gclk));
	jdff dff_B_g8Zkx60P2_0(.din(w_dff_B_zvaA5D1N9_0),.dout(w_dff_B_g8Zkx60P2_0),.clk(gclk));
	jdff dff_B_5MZ4CJjg4_0(.din(w_dff_B_g8Zkx60P2_0),.dout(w_dff_B_5MZ4CJjg4_0),.clk(gclk));
	jdff dff_B_6rYAchRu8_0(.din(w_dff_B_5MZ4CJjg4_0),.dout(w_dff_B_6rYAchRu8_0),.clk(gclk));
	jdff dff_B_U9I6NSKP4_0(.din(w_dff_B_6rYAchRu8_0),.dout(w_dff_B_U9I6NSKP4_0),.clk(gclk));
	jdff dff_B_VkqJ4JdF2_0(.din(w_dff_B_U9I6NSKP4_0),.dout(w_dff_B_VkqJ4JdF2_0),.clk(gclk));
	jdff dff_A_2qNBQAAz1_1(.dout(w_n1609_0[1]),.din(w_dff_A_2qNBQAAz1_1),.clk(gclk));
	jdff dff_A_KXq6F43g4_1(.dout(w_dff_A_2qNBQAAz1_1),.din(w_dff_A_KXq6F43g4_1),.clk(gclk));
	jdff dff_A_M7eigc2J0_1(.dout(w_dff_A_KXq6F43g4_1),.din(w_dff_A_M7eigc2J0_1),.clk(gclk));
	jdff dff_A_mE0bREcL4_1(.dout(w_dff_A_M7eigc2J0_1),.din(w_dff_A_mE0bREcL4_1),.clk(gclk));
	jdff dff_A_e3XV9LNK4_1(.dout(w_dff_A_mE0bREcL4_1),.din(w_dff_A_e3XV9LNK4_1),.clk(gclk));
	jdff dff_A_vxnwc74m0_1(.dout(w_dff_A_e3XV9LNK4_1),.din(w_dff_A_vxnwc74m0_1),.clk(gclk));
	jdff dff_A_WlQMOzsc4_1(.dout(w_dff_A_vxnwc74m0_1),.din(w_dff_A_WlQMOzsc4_1),.clk(gclk));
	jdff dff_A_q6RkgbSP8_1(.dout(w_dff_A_WlQMOzsc4_1),.din(w_dff_A_q6RkgbSP8_1),.clk(gclk));
	jdff dff_A_XhfRU2u52_1(.dout(w_dff_A_q6RkgbSP8_1),.din(w_dff_A_XhfRU2u52_1),.clk(gclk));
	jdff dff_A_0V4Iu1L22_1(.dout(w_dff_A_XhfRU2u52_1),.din(w_dff_A_0V4Iu1L22_1),.clk(gclk));
	jdff dff_A_Y90mAvUv5_1(.dout(w_dff_A_0V4Iu1L22_1),.din(w_dff_A_Y90mAvUv5_1),.clk(gclk));
	jdff dff_A_1iWUyKb64_1(.dout(w_dff_A_Y90mAvUv5_1),.din(w_dff_A_1iWUyKb64_1),.clk(gclk));
	jdff dff_A_stdcJoPf5_1(.dout(w_dff_A_1iWUyKb64_1),.din(w_dff_A_stdcJoPf5_1),.clk(gclk));
	jdff dff_A_4erDwzrp7_1(.dout(w_dff_A_stdcJoPf5_1),.din(w_dff_A_4erDwzrp7_1),.clk(gclk));
	jdff dff_A_H93Uu6Zn8_1(.dout(w_dff_A_4erDwzrp7_1),.din(w_dff_A_H93Uu6Zn8_1),.clk(gclk));
	jdff dff_A_pR8iYj328_1(.dout(w_dff_A_H93Uu6Zn8_1),.din(w_dff_A_pR8iYj328_1),.clk(gclk));
	jdff dff_A_EAQwzC245_1(.dout(w_dff_A_pR8iYj328_1),.din(w_dff_A_EAQwzC245_1),.clk(gclk));
	jdff dff_A_cKvkMZMF8_1(.dout(w_dff_A_EAQwzC245_1),.din(w_dff_A_cKvkMZMF8_1),.clk(gclk));
	jdff dff_A_a0wee1C72_1(.dout(w_dff_A_cKvkMZMF8_1),.din(w_dff_A_a0wee1C72_1),.clk(gclk));
	jdff dff_A_lOfGrWq38_1(.dout(w_dff_A_a0wee1C72_1),.din(w_dff_A_lOfGrWq38_1),.clk(gclk));
	jdff dff_B_EiferPjr7_1(.din(n1392),.dout(w_dff_B_EiferPjr7_1),.clk(gclk));
	jdff dff_B_LEYSzV9g6_1(.din(w_dff_B_EiferPjr7_1),.dout(w_dff_B_LEYSzV9g6_1),.clk(gclk));
	jdff dff_B_WDjFJlta3_1(.din(w_dff_B_LEYSzV9g6_1),.dout(w_dff_B_WDjFJlta3_1),.clk(gclk));
	jdff dff_B_A5UV8FbO1_1(.din(w_dff_B_WDjFJlta3_1),.dout(w_dff_B_A5UV8FbO1_1),.clk(gclk));
	jdff dff_B_vPNP0QHB0_1(.din(w_dff_B_A5UV8FbO1_1),.dout(w_dff_B_vPNP0QHB0_1),.clk(gclk));
	jdff dff_B_srRKSC302_1(.din(w_dff_B_vPNP0QHB0_1),.dout(w_dff_B_srRKSC302_1),.clk(gclk));
	jdff dff_A_uP4cssC57_1(.dout(w_n1447_0[1]),.din(w_dff_A_uP4cssC57_1),.clk(gclk));
	jdff dff_B_zLvkXYvw7_1(.din(n1412),.dout(w_dff_B_zLvkXYvw7_1),.clk(gclk));
	jdff dff_B_Ctzvl1pv9_1(.din(w_dff_B_zLvkXYvw7_1),.dout(w_dff_B_Ctzvl1pv9_1),.clk(gclk));
	jdff dff_B_ccoYs86D7_1(.din(w_dff_B_Ctzvl1pv9_1),.dout(w_dff_B_ccoYs86D7_1),.clk(gclk));
	jdff dff_B_fAtLgESn2_1(.din(w_dff_B_ccoYs86D7_1),.dout(w_dff_B_fAtLgESn2_1),.clk(gclk));
	jdff dff_B_h2h6XhD24_1(.din(w_dff_B_fAtLgESn2_1),.dout(w_dff_B_h2h6XhD24_1),.clk(gclk));
	jdff dff_B_78h5uKli9_1(.din(w_dff_B_h2h6XhD24_1),.dout(w_dff_B_78h5uKli9_1),.clk(gclk));
	jdff dff_B_y4lPWIZM9_1(.din(w_dff_B_78h5uKli9_1),.dout(w_dff_B_y4lPWIZM9_1),.clk(gclk));
	jdff dff_B_Ycw62p2G9_1(.din(w_dff_B_y4lPWIZM9_1),.dout(w_dff_B_Ycw62p2G9_1),.clk(gclk));
	jdff dff_B_OKGcimLH4_1(.din(w_dff_B_Ycw62p2G9_1),.dout(w_dff_B_OKGcimLH4_1),.clk(gclk));
	jdff dff_B_T5OrYCv76_1(.din(w_dff_B_OKGcimLH4_1),.dout(w_dff_B_T5OrYCv76_1),.clk(gclk));
	jdff dff_B_B8p0AihC4_0(.din(n1443),.dout(w_dff_B_B8p0AihC4_0),.clk(gclk));
	jdff dff_B_rYpnkdck4_0(.din(n1440),.dout(w_dff_B_rYpnkdck4_0),.clk(gclk));
	jdff dff_A_DAnZjvDa5_1(.dout(w_n1438_0[1]),.din(w_dff_A_DAnZjvDa5_1),.clk(gclk));
	jdff dff_A_RU3PesLf9_1(.dout(w_dff_A_DAnZjvDa5_1),.din(w_dff_A_RU3PesLf9_1),.clk(gclk));
	jdff dff_A_i4tnNOao0_1(.dout(w_dff_A_RU3PesLf9_1),.din(w_dff_A_i4tnNOao0_1),.clk(gclk));
	jdff dff_B_JlEetKWX5_0(.din(n1437),.dout(w_dff_B_JlEetKWX5_0),.clk(gclk));
	jdff dff_B_93VvCCoL9_1(.din(n1427),.dout(w_dff_B_93VvCCoL9_1),.clk(gclk));
	jdff dff_B_fBAZfIPF1_1(.din(n1428),.dout(w_dff_B_fBAZfIPF1_1),.clk(gclk));
	jdff dff_B_CmMYRjGy6_1(.din(w_dff_B_fBAZfIPF1_1),.dout(w_dff_B_CmMYRjGy6_1),.clk(gclk));
	jdff dff_B_k8wkP7V45_1(.din(w_dff_B_CmMYRjGy6_1),.dout(w_dff_B_k8wkP7V45_1),.clk(gclk));
	jdff dff_B_l5805JJW3_1(.din(w_dff_B_k8wkP7V45_1),.dout(w_dff_B_l5805JJW3_1),.clk(gclk));
	jdff dff_B_qtoGbi9Q3_1(.din(w_dff_B_l5805JJW3_1),.dout(w_dff_B_qtoGbi9Q3_1),.clk(gclk));
	jdff dff_B_DvW9Xmlr0_1(.din(w_dff_B_qtoGbi9Q3_1),.dout(w_dff_B_DvW9Xmlr0_1),.clk(gclk));
	jdff dff_B_mn2IDOe53_1(.din(w_dff_B_DvW9Xmlr0_1),.dout(w_dff_B_mn2IDOe53_1),.clk(gclk));
	jdff dff_B_ImFpiWwF0_1(.din(w_dff_B_mn2IDOe53_1),.dout(w_dff_B_ImFpiWwF0_1),.clk(gclk));
	jdff dff_B_6ADLqYUy0_1(.din(w_dff_B_ImFpiWwF0_1),.dout(w_dff_B_6ADLqYUy0_1),.clk(gclk));
	jdff dff_B_8lN77ZZV8_1(.din(w_dff_B_6ADLqYUy0_1),.dout(w_dff_B_8lN77ZZV8_1),.clk(gclk));
	jdff dff_B_E8bw2Xc02_1(.din(w_dff_B_8lN77ZZV8_1),.dout(w_dff_B_E8bw2Xc02_1),.clk(gclk));
	jdff dff_B_5hVWzVVv8_1(.din(n1414),.dout(w_dff_B_5hVWzVVv8_1),.clk(gclk));
	jdff dff_B_xPpdEmg91_1(.din(w_dff_B_5hVWzVVv8_1),.dout(w_dff_B_xPpdEmg91_1),.clk(gclk));
	jdff dff_B_hahaZNaU7_1(.din(w_dff_B_xPpdEmg91_1),.dout(w_dff_B_hahaZNaU7_1),.clk(gclk));
	jdff dff_B_m1reyT1g6_1(.din(w_dff_B_hahaZNaU7_1),.dout(w_dff_B_m1reyT1g6_1),.clk(gclk));
	jdff dff_B_DZsrSaJC9_1(.din(n1423),.dout(w_dff_B_DZsrSaJC9_1),.clk(gclk));
	jdff dff_B_5XddWEBp3_0(.din(n1422),.dout(w_dff_B_5XddWEBp3_0),.clk(gclk));
	jdff dff_A_HcOHyT6M2_0(.dout(w_n1421_0[0]),.din(w_dff_A_HcOHyT6M2_0),.clk(gclk));
	jdff dff_A_X51ckPEc8_0(.dout(w_dff_A_HcOHyT6M2_0),.din(w_dff_A_X51ckPEc8_0),.clk(gclk));
	jdff dff_A_dwyuefgZ4_0(.dout(w_dff_A_X51ckPEc8_0),.din(w_dff_A_dwyuefgZ4_0),.clk(gclk));
	jdff dff_B_41D4gjXK6_1(.din(n1415),.dout(w_dff_B_41D4gjXK6_1),.clk(gclk));
	jdff dff_A_q39Y62Qo9_1(.dout(w_n829_0[1]),.din(w_dff_A_q39Y62Qo9_1),.clk(gclk));
	jdff dff_A_7U8dAIfM4_0(.dout(w_n614_1[0]),.din(w_dff_A_7U8dAIfM4_0),.clk(gclk));
	jdff dff_A_Dj08AoB85_0(.dout(w_dff_A_7U8dAIfM4_0),.din(w_dff_A_Dj08AoB85_0),.clk(gclk));
	jdff dff_A_3BqQ1vZL7_0(.dout(w_dff_A_Dj08AoB85_0),.din(w_dff_A_3BqQ1vZL7_0),.clk(gclk));
	jdff dff_A_GRkkIbkc5_0(.dout(w_dff_A_3BqQ1vZL7_0),.din(w_dff_A_GRkkIbkc5_0),.clk(gclk));
	jdff dff_A_yFlhvwaL7_0(.dout(w_dff_A_GRkkIbkc5_0),.din(w_dff_A_yFlhvwaL7_0),.clk(gclk));
	jdff dff_A_vMZcvEne7_2(.dout(w_n614_1[2]),.din(w_dff_A_vMZcvEne7_2),.clk(gclk));
	jdff dff_A_v8ccX43L2_2(.dout(w_dff_A_vMZcvEne7_2),.din(w_dff_A_v8ccX43L2_2),.clk(gclk));
	jdff dff_A_6R0eBoST5_2(.dout(w_dff_A_v8ccX43L2_2),.din(w_dff_A_6R0eBoST5_2),.clk(gclk));
	jdff dff_A_43kEHPEg7_2(.dout(w_dff_A_6R0eBoST5_2),.din(w_dff_A_43kEHPEg7_2),.clk(gclk));
	jdff dff_A_7VdfCcrB8_2(.dout(w_dff_A_43kEHPEg7_2),.din(w_dff_A_7VdfCcrB8_2),.clk(gclk));
	jdff dff_A_SfMgCxe87_2(.dout(w_dff_A_7VdfCcrB8_2),.din(w_dff_A_SfMgCxe87_2),.clk(gclk));
	jdff dff_A_J6xtzue03_1(.dout(w_n828_0[1]),.din(w_dff_A_J6xtzue03_1),.clk(gclk));
	jdff dff_A_exhrGTRb2_1(.dout(w_dff_A_J6xtzue03_1),.din(w_dff_A_exhrGTRb2_1),.clk(gclk));
	jdff dff_A_U8cEK5rx7_1(.dout(w_dff_A_exhrGTRb2_1),.din(w_dff_A_U8cEK5rx7_1),.clk(gclk));
	jdff dff_A_bsDESXrn1_1(.dout(w_dff_A_U8cEK5rx7_1),.din(w_dff_A_bsDESXrn1_1),.clk(gclk));
	jdff dff_A_Llzfcz2D6_1(.dout(w_dff_A_bsDESXrn1_1),.din(w_dff_A_Llzfcz2D6_1),.clk(gclk));
	jdff dff_A_9p8FwHgm0_1(.dout(w_dff_A_Llzfcz2D6_1),.din(w_dff_A_9p8FwHgm0_1),.clk(gclk));
	jdff dff_A_oFlFmqrn6_2(.dout(w_n828_0[2]),.din(w_dff_A_oFlFmqrn6_2),.clk(gclk));
	jdff dff_A_VZ74eUt02_2(.dout(w_dff_A_oFlFmqrn6_2),.din(w_dff_A_VZ74eUt02_2),.clk(gclk));
	jdff dff_B_3haLFshg7_2(.din(n787),.dout(w_dff_B_3haLFshg7_2),.clk(gclk));
	jdff dff_B_YNCr1ghA7_2(.din(w_dff_B_3haLFshg7_2),.dout(w_dff_B_YNCr1ghA7_2),.clk(gclk));
	jdff dff_B_H8r2rb7a7_2(.din(w_dff_B_YNCr1ghA7_2),.dout(w_dff_B_H8r2rb7a7_2),.clk(gclk));
	jdff dff_B_qSk3uBpR2_2(.din(w_dff_B_H8r2rb7a7_2),.dout(w_dff_B_qSk3uBpR2_2),.clk(gclk));
	jdff dff_B_kx3bsKHd9_2(.din(w_dff_B_qSk3uBpR2_2),.dout(w_dff_B_kx3bsKHd9_2),.clk(gclk));
	jdff dff_B_5c34sflw2_2(.din(w_dff_B_kx3bsKHd9_2),.dout(w_dff_B_5c34sflw2_2),.clk(gclk));
	jdff dff_B_YU7MduXM0_2(.din(w_dff_B_5c34sflw2_2),.dout(w_dff_B_YU7MduXM0_2),.clk(gclk));
	jdff dff_B_PlWYkjCq5_2(.din(w_dff_B_YU7MduXM0_2),.dout(w_dff_B_PlWYkjCq5_2),.clk(gclk));
	jdff dff_B_G0r8g5BP1_2(.din(w_dff_B_PlWYkjCq5_2),.dout(w_dff_B_G0r8g5BP1_2),.clk(gclk));
	jdff dff_A_p02ZZeyY1_1(.dout(w_n779_0[1]),.din(w_dff_A_p02ZZeyY1_1),.clk(gclk));
	jdff dff_A_PiutBOKW9_1(.dout(w_dff_A_p02ZZeyY1_1),.din(w_dff_A_PiutBOKW9_1),.clk(gclk));
	jdff dff_A_fo7ty2Ig3_1(.dout(w_dff_A_PiutBOKW9_1),.din(w_dff_A_fo7ty2Ig3_1),.clk(gclk));
	jdff dff_A_vi7fcVaA1_1(.dout(w_dff_A_fo7ty2Ig3_1),.din(w_dff_A_vi7fcVaA1_1),.clk(gclk));
	jdff dff_A_qyJST7g97_1(.dout(w_dff_A_vi7fcVaA1_1),.din(w_dff_A_qyJST7g97_1),.clk(gclk));
	jdff dff_A_T9XOHi6A6_1(.dout(w_dff_A_qyJST7g97_1),.din(w_dff_A_T9XOHi6A6_1),.clk(gclk));
	jdff dff_A_FmJG8Dnv8_1(.dout(w_dff_A_T9XOHi6A6_1),.din(w_dff_A_FmJG8Dnv8_1),.clk(gclk));
	jdff dff_A_19NKEVfM8_1(.dout(w_dff_A_FmJG8Dnv8_1),.din(w_dff_A_19NKEVfM8_1),.clk(gclk));
	jdff dff_A_zsOTnmHl7_1(.dout(w_dff_A_19NKEVfM8_1),.din(w_dff_A_zsOTnmHl7_1),.clk(gclk));
	jdff dff_A_8mvt0AeL9_1(.dout(w_dff_A_zsOTnmHl7_1),.din(w_dff_A_8mvt0AeL9_1),.clk(gclk));
	jdff dff_A_ZHVBNmEb4_1(.dout(w_dff_A_8mvt0AeL9_1),.din(w_dff_A_ZHVBNmEb4_1),.clk(gclk));
	jdff dff_A_oxz4LApm0_1(.dout(w_dff_A_ZHVBNmEb4_1),.din(w_dff_A_oxz4LApm0_1),.clk(gclk));
	jdff dff_A_2vLDGwbn1_1(.dout(w_n636_1[1]),.din(w_dff_A_2vLDGwbn1_1),.clk(gclk));
	jdff dff_A_YybsqF5R9_1(.dout(w_dff_A_2vLDGwbn1_1),.din(w_dff_A_YybsqF5R9_1),.clk(gclk));
	jdff dff_A_lDwR0oxZ1_2(.dout(w_n636_0[2]),.din(w_dff_A_lDwR0oxZ1_2),.clk(gclk));
	jdff dff_A_83I4TDbd0_0(.dout(w_n1411_0[0]),.din(w_dff_A_83I4TDbd0_0),.clk(gclk));
	jdff dff_A_VhoHiYwh2_0(.dout(w_dff_A_83I4TDbd0_0),.din(w_dff_A_VhoHiYwh2_0),.clk(gclk));
	jdff dff_A_XEg2A39h3_0(.dout(w_dff_A_VhoHiYwh2_0),.din(w_dff_A_XEg2A39h3_0),.clk(gclk));
	jdff dff_A_1MjHR3At8_0(.dout(w_dff_A_XEg2A39h3_0),.din(w_dff_A_1MjHR3At8_0),.clk(gclk));
	jdff dff_A_FKyPYXmF7_0(.dout(w_dff_A_1MjHR3At8_0),.din(w_dff_A_FKyPYXmF7_0),.clk(gclk));
	jdff dff_A_CRdPderv7_0(.dout(w_dff_A_FKyPYXmF7_0),.din(w_dff_A_CRdPderv7_0),.clk(gclk));
	jdff dff_A_nQxZ6Apw4_0(.dout(w_dff_A_CRdPderv7_0),.din(w_dff_A_nQxZ6Apw4_0),.clk(gclk));
	jdff dff_A_bInQ2ewd0_0(.dout(w_dff_A_nQxZ6Apw4_0),.din(w_dff_A_bInQ2ewd0_0),.clk(gclk));
	jdff dff_A_8aOzhEPB5_0(.dout(w_dff_A_bInQ2ewd0_0),.din(w_dff_A_8aOzhEPB5_0),.clk(gclk));
	jdff dff_A_9i10deTR1_0(.dout(w_dff_A_8aOzhEPB5_0),.din(w_dff_A_9i10deTR1_0),.clk(gclk));
	jdff dff_A_yQLIJlPF6_0(.dout(w_dff_A_9i10deTR1_0),.din(w_dff_A_yQLIJlPF6_0),.clk(gclk));
	jdff dff_A_07bBmpDT9_0(.dout(w_n1409_0[0]),.din(w_dff_A_07bBmpDT9_0),.clk(gclk));
	jdff dff_B_jKVjrq5X9_1(.din(n1405),.dout(w_dff_B_jKVjrq5X9_1),.clk(gclk));
	jdff dff_B_fhLSiVLT7_0(.din(n1407),.dout(w_dff_B_fhLSiVLT7_0),.clk(gclk));
	jdff dff_B_E6HVoo1T4_0(.din(w_dff_B_fhLSiVLT7_0),.dout(w_dff_B_E6HVoo1T4_0),.clk(gclk));
	jdff dff_B_TQRLK7av2_0(.din(w_dff_B_E6HVoo1T4_0),.dout(w_dff_B_TQRLK7av2_0),.clk(gclk));
	jdff dff_B_0jfqp2Sr6_0(.din(w_dff_B_TQRLK7av2_0),.dout(w_dff_B_0jfqp2Sr6_0),.clk(gclk));
	jdff dff_A_A7pyJF0q2_1(.dout(w_n968_0[1]),.din(w_dff_A_A7pyJF0q2_1),.clk(gclk));
	jdff dff_A_GIQAnLri7_1(.dout(w_dff_A_A7pyJF0q2_1),.din(w_dff_A_GIQAnLri7_1),.clk(gclk));
	jdff dff_A_c2uT18W97_1(.dout(w_dff_A_GIQAnLri7_1),.din(w_dff_A_c2uT18W97_1),.clk(gclk));
	jdff dff_A_h1JDWaJA3_1(.dout(w_dff_A_c2uT18W97_1),.din(w_dff_A_h1JDWaJA3_1),.clk(gclk));
	jdff dff_A_qkS26nqD6_1(.dout(w_dff_A_h1JDWaJA3_1),.din(w_dff_A_qkS26nqD6_1),.clk(gclk));
	jdff dff_B_M8L1t6OB9_2(.din(n968),.dout(w_dff_B_M8L1t6OB9_2),.clk(gclk));
	jdff dff_B_sCZfvn0t7_2(.din(w_dff_B_M8L1t6OB9_2),.dout(w_dff_B_sCZfvn0t7_2),.clk(gclk));
	jdff dff_B_Ki3Mc9955_2(.din(w_dff_B_sCZfvn0t7_2),.dout(w_dff_B_Ki3Mc9955_2),.clk(gclk));
	jdff dff_B_p2gEwM9Z5_2(.din(w_dff_B_Ki3Mc9955_2),.dout(w_dff_B_p2gEwM9Z5_2),.clk(gclk));
	jdff dff_B_qYv6NP3V6_2(.din(w_dff_B_p2gEwM9Z5_2),.dout(w_dff_B_qYv6NP3V6_2),.clk(gclk));
	jdff dff_B_246mbD024_0(.din(n1404),.dout(w_dff_B_246mbD024_0),.clk(gclk));
	jdff dff_B_IKKyRrnr9_0(.din(w_dff_B_246mbD024_0),.dout(w_dff_B_IKKyRrnr9_0),.clk(gclk));
	jdff dff_B_S1s3UIPE3_1(.din(n1401),.dout(w_dff_B_S1s3UIPE3_1),.clk(gclk));
	jdff dff_B_dh32HErn3_1(.din(w_dff_B_S1s3UIPE3_1),.dout(w_dff_B_dh32HErn3_1),.clk(gclk));
	jdff dff_B_Q5aEoJqx2_1(.din(w_dff_B_dh32HErn3_1),.dout(w_dff_B_Q5aEoJqx2_1),.clk(gclk));
	jdff dff_A_qLi9mKAP9_1(.dout(w_n651_0[1]),.din(w_dff_A_qLi9mKAP9_1),.clk(gclk));
	jdff dff_A_i29xRiPG6_1(.dout(w_dff_A_qLi9mKAP9_1),.din(w_dff_A_i29xRiPG6_1),.clk(gclk));
	jdff dff_A_MmFNpZCS8_1(.dout(w_dff_A_i29xRiPG6_1),.din(w_dff_A_MmFNpZCS8_1),.clk(gclk));
	jdff dff_A_HmG6Z6ho0_2(.dout(w_n651_0[2]),.din(w_dff_A_HmG6Z6ho0_2),.clk(gclk));
	jdff dff_A_2gdmoAsn9_2(.dout(w_dff_A_HmG6Z6ho0_2),.din(w_dff_A_2gdmoAsn9_2),.clk(gclk));
	jdff dff_A_6tH0pIWo0_2(.dout(w_dff_A_2gdmoAsn9_2),.din(w_dff_A_6tH0pIWo0_2),.clk(gclk));
	jdff dff_A_RMtnfA0Q2_2(.dout(w_dff_A_6tH0pIWo0_2),.din(w_dff_A_RMtnfA0Q2_2),.clk(gclk));
	jdff dff_A_Cx4XFVwu0_2(.dout(w_dff_A_RMtnfA0Q2_2),.din(w_dff_A_Cx4XFVwu0_2),.clk(gclk));
	jdff dff_A_ppNgcQAy5_2(.dout(w_dff_A_Cx4XFVwu0_2),.din(w_dff_A_ppNgcQAy5_2),.clk(gclk));
	jdff dff_A_uonOlQ6T0_2(.dout(w_dff_A_ppNgcQAy5_2),.din(w_dff_A_uonOlQ6T0_2),.clk(gclk));
	jdff dff_B_5M9btRQs8_3(.din(n651),.dout(w_dff_B_5M9btRQs8_3),.clk(gclk));
	jdff dff_A_l8vT5vQK1_0(.dout(w_n650_0[0]),.din(w_dff_A_l8vT5vQK1_0),.clk(gclk));
	jdff dff_A_VNLyh4yD4_0(.dout(w_dff_A_l8vT5vQK1_0),.din(w_dff_A_VNLyh4yD4_0),.clk(gclk));
	jdff dff_A_t9r41Nco3_0(.dout(w_dff_A_VNLyh4yD4_0),.din(w_dff_A_t9r41Nco3_0),.clk(gclk));
	jdff dff_A_vw1ZzAog0_0(.dout(w_dff_A_t9r41Nco3_0),.din(w_dff_A_vw1ZzAog0_0),.clk(gclk));
	jdff dff_A_kLsYy4kh4_0(.dout(w_dff_A_vw1ZzAog0_0),.din(w_dff_A_kLsYy4kh4_0),.clk(gclk));
	jdff dff_A_rhwnmWmK9_0(.dout(w_dff_A_kLsYy4kh4_0),.din(w_dff_A_rhwnmWmK9_0),.clk(gclk));
	jdff dff_A_ohl3pi0p0_0(.dout(w_dff_A_rhwnmWmK9_0),.din(w_dff_A_ohl3pi0p0_0),.clk(gclk));
	jdff dff_A_nXyAlhw77_0(.dout(w_dff_A_ohl3pi0p0_0),.din(w_dff_A_nXyAlhw77_0),.clk(gclk));
	jdff dff_A_KnkyxPvf7_0(.dout(w_dff_A_nXyAlhw77_0),.din(w_dff_A_KnkyxPvf7_0),.clk(gclk));
	jdff dff_B_1KEajjX92_1(.din(n1395),.dout(w_dff_B_1KEajjX92_1),.clk(gclk));
	jdff dff_A_kUQDiRdJ1_1(.dout(w_n740_0[1]),.din(w_dff_A_kUQDiRdJ1_1),.clk(gclk));
	jdff dff_A_JlBhJpDg0_0(.dout(w_n739_1[0]),.din(w_dff_A_JlBhJpDg0_0),.clk(gclk));
	jdff dff_A_d4qRLEDP4_0(.dout(w_dff_A_JlBhJpDg0_0),.din(w_dff_A_d4qRLEDP4_0),.clk(gclk));
	jdff dff_A_a3SyjLHw4_0(.dout(w_dff_A_d4qRLEDP4_0),.din(w_dff_A_a3SyjLHw4_0),.clk(gclk));
	jdff dff_A_sutFpcGy7_0(.dout(w_dff_A_a3SyjLHw4_0),.din(w_dff_A_sutFpcGy7_0),.clk(gclk));
	jdff dff_A_uCbpn1v40_0(.dout(w_dff_A_sutFpcGy7_0),.din(w_dff_A_uCbpn1v40_0),.clk(gclk));
	jdff dff_A_D8G3IhyY8_0(.dout(w_dff_A_uCbpn1v40_0),.din(w_dff_A_D8G3IhyY8_0),.clk(gclk));
	jdff dff_A_ye3YonQl8_0(.dout(w_dff_A_D8G3IhyY8_0),.din(w_dff_A_ye3YonQl8_0),.clk(gclk));
	jdff dff_A_wNlLgMxG5_0(.dout(w_dff_A_ye3YonQl8_0),.din(w_dff_A_wNlLgMxG5_0),.clk(gclk));
	jdff dff_A_yKP8tZG88_0(.dout(w_dff_A_wNlLgMxG5_0),.din(w_dff_A_yKP8tZG88_0),.clk(gclk));
	jdff dff_A_OuggQ7wO4_2(.dout(w_n739_0[2]),.din(w_dff_A_OuggQ7wO4_2),.clk(gclk));
	jdff dff_A_xoIC4ohq8_2(.dout(w_dff_A_OuggQ7wO4_2),.din(w_dff_A_xoIC4ohq8_2),.clk(gclk));
	jdff dff_A_cPVSayx24_2(.dout(w_dff_A_xoIC4ohq8_2),.din(w_dff_A_cPVSayx24_2),.clk(gclk));
	jdff dff_A_LSHlXkhS6_2(.dout(w_dff_A_cPVSayx24_2),.din(w_dff_A_LSHlXkhS6_2),.clk(gclk));
	jdff dff_A_FIgmJxWn2_2(.dout(w_dff_A_LSHlXkhS6_2),.din(w_dff_A_FIgmJxWn2_2),.clk(gclk));
	jdff dff_A_MlFFv0D18_2(.dout(w_n649_0[2]),.din(w_dff_A_MlFFv0D18_2),.clk(gclk));
	jdff dff_B_5BaMNZE13_0(.din(n648),.dout(w_dff_B_5BaMNZE13_0),.clk(gclk));
	jdff dff_B_d9S4yyXW1_1(.din(G323),.dout(w_dff_B_d9S4yyXW1_1),.clk(gclk));
	jdff dff_A_Ah5jx5xq6_0(.dout(w_n640_1[0]),.din(w_dff_A_Ah5jx5xq6_0),.clk(gclk));
	jdff dff_A_5FaKLTAu6_0(.dout(w_dff_A_Ah5jx5xq6_0),.din(w_dff_A_5FaKLTAu6_0),.clk(gclk));
	jdff dff_A_hdHaghVi9_0(.dout(w_dff_A_5FaKLTAu6_0),.din(w_dff_A_hdHaghVi9_0),.clk(gclk));
	jdff dff_A_7y3fmF6K9_0(.dout(w_dff_A_hdHaghVi9_0),.din(w_dff_A_7y3fmF6K9_0),.clk(gclk));
	jdff dff_A_KMCz86P61_0(.dout(w_dff_A_7y3fmF6K9_0),.din(w_dff_A_KMCz86P61_0),.clk(gclk));
	jdff dff_A_ZHwX3Y8X3_0(.dout(w_dff_A_KMCz86P61_0),.din(w_dff_A_ZHwX3Y8X3_0),.clk(gclk));
	jdff dff_A_T63qrX6K1_0(.dout(w_dff_A_ZHwX3Y8X3_0),.din(w_dff_A_T63qrX6K1_0),.clk(gclk));
	jdff dff_A_EgHcgpFC8_0(.dout(w_dff_A_T63qrX6K1_0),.din(w_dff_A_EgHcgpFC8_0),.clk(gclk));
	jdff dff_A_mB80jkcS5_0(.dout(w_dff_A_EgHcgpFC8_0),.din(w_dff_A_mB80jkcS5_0),.clk(gclk));
	jdff dff_A_zpxvzAgL6_0(.dout(w_dff_A_mB80jkcS5_0),.din(w_dff_A_zpxvzAgL6_0),.clk(gclk));
	jdff dff_A_OwxKxIKB0_0(.dout(w_dff_A_zpxvzAgL6_0),.din(w_dff_A_OwxKxIKB0_0),.clk(gclk));
	jdff dff_A_RZPL5dbr7_0(.dout(w_n646_0[0]),.din(w_dff_A_RZPL5dbr7_0),.clk(gclk));
	jdff dff_A_mdWYaNkU6_0(.dout(w_dff_A_RZPL5dbr7_0),.din(w_dff_A_mdWYaNkU6_0),.clk(gclk));
	jdff dff_B_kjeHPyV10_0(.din(n644),.dout(w_dff_B_kjeHPyV10_0),.clk(gclk));
	jdff dff_B_Ku26dCwl2_1(.din(G315),.dout(w_dff_B_Ku26dCwl2_1),.clk(gclk));
	jdff dff_A_7qnZTphL5_1(.dout(w_n640_0[1]),.din(w_dff_A_7qnZTphL5_1),.clk(gclk));
	jdff dff_A_BkVAH2ZV8_2(.dout(w_n640_0[2]),.din(w_dff_A_BkVAH2ZV8_2),.clk(gclk));
	jdff dff_A_vwcKKIkE5_2(.dout(w_dff_A_BkVAH2ZV8_2),.din(w_dff_A_vwcKKIkE5_2),.clk(gclk));
	jdff dff_A_VRwsdY0y4_2(.dout(w_dff_A_vwcKKIkE5_2),.din(w_dff_A_VRwsdY0y4_2),.clk(gclk));
	jdff dff_A_A3OPp8uX3_2(.dout(w_dff_A_VRwsdY0y4_2),.din(w_dff_A_A3OPp8uX3_2),.clk(gclk));
	jdff dff_A_azJ1Cwza1_2(.dout(w_dff_A_A3OPp8uX3_2),.din(w_dff_A_azJ1Cwza1_2),.clk(gclk));
	jdff dff_A_6qlwNx9c4_2(.dout(w_dff_A_azJ1Cwza1_2),.din(w_dff_A_6qlwNx9c4_2),.clk(gclk));
	jdff dff_A_BeDjNIWs3_2(.dout(w_dff_A_6qlwNx9c4_2),.din(w_dff_A_BeDjNIWs3_2),.clk(gclk));
	jdff dff_A_sp6qozvR2_2(.dout(w_dff_A_BeDjNIWs3_2),.din(w_dff_A_sp6qozvR2_2),.clk(gclk));
	jdff dff_A_tAJIxZZM3_2(.dout(w_dff_A_sp6qozvR2_2),.din(w_dff_A_tAJIxZZM3_2),.clk(gclk));
	jdff dff_A_zHqaBtl11_2(.dout(w_dff_A_tAJIxZZM3_2),.din(w_dff_A_zHqaBtl11_2),.clk(gclk));
	jdff dff_A_m2MJmds47_2(.dout(w_dff_A_zHqaBtl11_2),.din(w_dff_A_m2MJmds47_2),.clk(gclk));
	jdff dff_B_y2tM4x287_1(.din(n637),.dout(w_dff_B_y2tM4x287_1),.clk(gclk));
	jdff dff_B_9MSpMEdm3_1(.din(G307),.dout(w_dff_B_9MSpMEdm3_1),.clk(gclk));
	jdff dff_B_l1rPpzD15_0(.din(n1393),.dout(w_dff_B_l1rPpzD15_0),.clk(gclk));
	jdff dff_B_QJtKWBiP2_0(.din(w_dff_B_l1rPpzD15_0),.dout(w_dff_B_QJtKWBiP2_0),.clk(gclk));
	jdff dff_B_bavSCnqv8_0(.din(w_dff_B_QJtKWBiP2_0),.dout(w_dff_B_bavSCnqv8_0),.clk(gclk));
	jdff dff_A_607vqbmS9_0(.dout(w_n631_0[0]),.din(w_dff_A_607vqbmS9_0),.clk(gclk));
	jdff dff_A_0bob9csf8_0(.dout(w_dff_A_607vqbmS9_0),.din(w_dff_A_0bob9csf8_0),.clk(gclk));
	jdff dff_A_HIdUAKGh5_0(.dout(w_dff_A_0bob9csf8_0),.din(w_dff_A_HIdUAKGh5_0),.clk(gclk));
	jdff dff_A_nmDxEz0M2_1(.dout(w_n629_0[1]),.din(w_dff_A_nmDxEz0M2_1),.clk(gclk));
	jdff dff_A_YPqa7FE77_1(.dout(w_dff_A_nmDxEz0M2_1),.din(w_dff_A_YPqa7FE77_1),.clk(gclk));
	jdff dff_A_ArazxxYs6_1(.dout(w_dff_A_YPqa7FE77_1),.din(w_dff_A_ArazxxYs6_1),.clk(gclk));
	jdff dff_A_y078HFsd3_1(.dout(w_n628_0[1]),.din(w_dff_A_y078HFsd3_1),.clk(gclk));
	jdff dff_B_VrYukKn71_0(.din(n627),.dout(w_dff_B_VrYukKn71_0),.clk(gclk));
	jdff dff_A_PGqWpFTY3_0(.dout(w_n625_0[0]),.din(w_dff_A_PGqWpFTY3_0),.clk(gclk));
	jdff dff_A_ye7KwXvM9_2(.dout(w_n625_0[2]),.din(w_dff_A_ye7KwXvM9_2),.clk(gclk));
	jdff dff_A_rPjvbile5_0(.dout(w_n623_0[0]),.din(w_dff_A_rPjvbile5_0),.clk(gclk));
	jdff dff_B_rkiHOKfh7_0(.din(n616),.dout(w_dff_B_rkiHOKfh7_0),.clk(gclk));
	jdff dff_A_7yrUm62o8_0(.dout(w_G2174_0[0]),.din(w_dff_A_7yrUm62o8_0),.clk(gclk));
	jdff dff_A_zm4lqhY66_0(.dout(w_dff_A_7yrUm62o8_0),.din(w_dff_A_zm4lqhY66_0),.clk(gclk));
	jdff dff_A_5Xz5M9m92_0(.dout(w_dff_A_zm4lqhY66_0),.din(w_dff_A_5Xz5M9m92_0),.clk(gclk));
	jdff dff_A_ekf3WwRm4_0(.dout(w_dff_A_5Xz5M9m92_0),.din(w_dff_A_ekf3WwRm4_0),.clk(gclk));
	jdff dff_A_pqviEFAC5_0(.dout(w_dff_A_ekf3WwRm4_0),.din(w_dff_A_pqviEFAC5_0),.clk(gclk));
	jdff dff_A_rjfCWH7v3_0(.dout(w_dff_A_pqviEFAC5_0),.din(w_dff_A_rjfCWH7v3_0),.clk(gclk));
	jdff dff_A_JZRfTq6S6_0(.dout(w_dff_A_rjfCWH7v3_0),.din(w_dff_A_JZRfTq6S6_0),.clk(gclk));
	jdff dff_A_IBfCtatM8_0(.dout(w_dff_A_JZRfTq6S6_0),.din(w_dff_A_IBfCtatM8_0),.clk(gclk));
	jdff dff_A_tO8jjP8l6_0(.dout(w_dff_A_IBfCtatM8_0),.din(w_dff_A_tO8jjP8l6_0),.clk(gclk));
	jdff dff_A_5bV9BeUp6_0(.dout(w_dff_A_tO8jjP8l6_0),.din(w_dff_A_5bV9BeUp6_0),.clk(gclk));
	jdff dff_A_2PvgxPFn8_0(.dout(w_dff_A_5bV9BeUp6_0),.din(w_dff_A_2PvgxPFn8_0),.clk(gclk));
	jdff dff_A_J7IMqfUf0_2(.dout(w_G2174_0[2]),.din(w_dff_A_J7IMqfUf0_2),.clk(gclk));
	jdff dff_A_eqOLkfew4_2(.dout(w_dff_A_J7IMqfUf0_2),.din(w_dff_A_eqOLkfew4_2),.clk(gclk));
	jdff dff_A_bYIpvWPS6_2(.dout(w_dff_A_eqOLkfew4_2),.din(w_dff_A_bYIpvWPS6_2),.clk(gclk));
	jdff dff_A_G1x36azM6_2(.dout(w_dff_A_bYIpvWPS6_2),.din(w_dff_A_G1x36azM6_2),.clk(gclk));
	jdff dff_A_CNIbL2NR6_2(.dout(w_dff_A_G1x36azM6_2),.din(w_dff_A_CNIbL2NR6_2),.clk(gclk));
	jdff dff_A_wKjQFHTu1_2(.dout(w_dff_A_CNIbL2NR6_2),.din(w_dff_A_wKjQFHTu1_2),.clk(gclk));
	jdff dff_A_ESHT4cdV3_2(.dout(w_dff_A_wKjQFHTu1_2),.din(w_dff_A_ESHT4cdV3_2),.clk(gclk));
	jdff dff_A_yp2Uiusj4_2(.dout(w_dff_A_ESHT4cdV3_2),.din(w_dff_A_yp2Uiusj4_2),.clk(gclk));
	jdff dff_B_JGqAcsRr8_1(.din(n711),.dout(w_dff_B_JGqAcsRr8_1),.clk(gclk));
	jdff dff_B_GHUFqe1f3_1(.din(w_dff_B_JGqAcsRr8_1),.dout(w_dff_B_GHUFqe1f3_1),.clk(gclk));
	jdff dff_B_fulIQZQl7_1(.din(w_dff_B_GHUFqe1f3_1),.dout(w_dff_B_fulIQZQl7_1),.clk(gclk));
	jdff dff_B_9sooi4Uc8_1(.din(w_dff_B_fulIQZQl7_1),.dout(w_dff_B_9sooi4Uc8_1),.clk(gclk));
	jdff dff_B_8kjyRUHx5_1(.din(w_dff_B_9sooi4Uc8_1),.dout(w_dff_B_8kjyRUHx5_1),.clk(gclk));
	jdff dff_B_UwWcPl1b7_1(.din(w_dff_B_8kjyRUHx5_1),.dout(w_dff_B_UwWcPl1b7_1),.clk(gclk));
	jdff dff_B_SLHDcqRL3_1(.din(n712),.dout(w_dff_B_SLHDcqRL3_1),.clk(gclk));
	jdff dff_B_t1eZh6es9_1(.din(w_dff_B_SLHDcqRL3_1),.dout(w_dff_B_t1eZh6es9_1),.clk(gclk));
	jdff dff_B_b1MTaIZk2_1(.din(w_dff_B_t1eZh6es9_1),.dout(w_dff_B_b1MTaIZk2_1),.clk(gclk));
	jdff dff_B_LeAwGtZq7_1(.din(w_dff_B_b1MTaIZk2_1),.dout(w_dff_B_LeAwGtZq7_1),.clk(gclk));
	jdff dff_B_boRSAyMn0_1(.din(w_dff_B_LeAwGtZq7_1),.dout(w_dff_B_boRSAyMn0_1),.clk(gclk));
	jdff dff_B_WFuUAlZN4_1(.din(n713),.dout(w_dff_B_WFuUAlZN4_1),.clk(gclk));
	jdff dff_B_znUCkEJB4_1(.din(w_dff_B_WFuUAlZN4_1),.dout(w_dff_B_znUCkEJB4_1),.clk(gclk));
	jdff dff_B_W4dZU0oB8_1(.din(w_dff_B_znUCkEJB4_1),.dout(w_dff_B_W4dZU0oB8_1),.clk(gclk));
	jdff dff_B_J8ZZvl7V7_1(.din(w_dff_B_W4dZU0oB8_1),.dout(w_dff_B_J8ZZvl7V7_1),.clk(gclk));
	jdff dff_A_jDdGjmD57_0(.dout(w_n723_0[0]),.din(w_dff_A_jDdGjmD57_0),.clk(gclk));
	jdff dff_A_IFsxbyU17_0(.dout(w_n621_2[0]),.din(w_dff_A_IFsxbyU17_0),.clk(gclk));
	jdff dff_A_9v7IrxGW5_1(.dout(w_n721_0[1]),.din(w_dff_A_9v7IrxGW5_1),.clk(gclk));
	jdff dff_A_xwNgPe5F2_1(.dout(w_dff_A_9v7IrxGW5_1),.din(w_dff_A_xwNgPe5F2_1),.clk(gclk));
	jdff dff_A_QfJbN9cG1_1(.dout(w_dff_A_xwNgPe5F2_1),.din(w_dff_A_QfJbN9cG1_1),.clk(gclk));
	jdff dff_A_fZ1P4Zf60_1(.dout(w_dff_A_QfJbN9cG1_1),.din(w_dff_A_fZ1P4Zf60_1),.clk(gclk));
	jdff dff_A_c6KmzTiU9_1(.dout(w_dff_A_fZ1P4Zf60_1),.din(w_dff_A_c6KmzTiU9_1),.clk(gclk));
	jdff dff_A_BlrkuVzQ3_1(.dout(w_dff_A_c6KmzTiU9_1),.din(w_dff_A_BlrkuVzQ3_1),.clk(gclk));
	jdff dff_A_JD0BOWzY6_0(.dout(w_G358_0[0]),.din(w_dff_A_JD0BOWzY6_0),.clk(gclk));
	jdff dff_A_tNKKSYbO1_0(.dout(w_n388_1[0]),.din(w_dff_A_tNKKSYbO1_0),.clk(gclk));
	jdff dff_A_UvZHh7uC5_1(.dout(w_n388_1[1]),.din(w_dff_A_UvZHh7uC5_1),.clk(gclk));
	jdff dff_A_6QtFNhGn3_1(.dout(w_n717_0[1]),.din(w_dff_A_6QtFNhGn3_1),.clk(gclk));
	jdff dff_A_bRFzw5NC2_1(.dout(w_dff_A_6QtFNhGn3_1),.din(w_dff_A_bRFzw5NC2_1),.clk(gclk));
	jdff dff_A_HKufdfLD0_1(.dout(w_dff_A_bRFzw5NC2_1),.din(w_dff_A_HKufdfLD0_1),.clk(gclk));
	jdff dff_A_tGhsZud05_2(.dout(w_n717_0[2]),.din(w_dff_A_tGhsZud05_2),.clk(gclk));
	jdff dff_A_CKr4KLtG9_2(.dout(w_dff_A_tGhsZud05_2),.din(w_dff_A_CKr4KLtG9_2),.clk(gclk));
	jdff dff_A_IcUKXp9b7_0(.dout(w_G348_0[0]),.din(w_dff_A_IcUKXp9b7_0),.clk(gclk));
	jdff dff_A_IDL7tBGd6_0(.dout(w_G332_2[0]),.din(w_dff_A_IDL7tBGd6_0),.clk(gclk));
	jdff dff_A_n0fgwF552_0(.dout(w_n437_1[0]),.din(w_dff_A_n0fgwF552_0),.clk(gclk));
	jdff dff_A_S9nwTBvd1_1(.dout(w_n437_1[1]),.din(w_dff_A_S9nwTBvd1_1),.clk(gclk));
	jdff dff_A_289YKKsd7_0(.dout(w_G332_3[0]),.din(w_dff_A_289YKKsd7_0),.clk(gclk));
	jdff dff_A_5nV0ELg97_2(.dout(w_G332_3[2]),.din(w_dff_A_5nV0ELg97_2),.clk(gclk));
	jdff dff_A_gHKJPNrq2_0(.dout(w_n410_1[0]),.din(w_dff_A_gHKJPNrq2_0),.clk(gclk));
	jdff dff_A_tX71DhYN1_0(.dout(w_n614_2[0]),.din(w_dff_A_tX71DhYN1_0),.clk(gclk));
	jdff dff_A_vjaJejNG5_0(.dout(w_dff_A_tX71DhYN1_0),.din(w_dff_A_vjaJejNG5_0),.clk(gclk));
	jdff dff_A_JWom5X3a3_0(.dout(w_dff_A_vjaJejNG5_0),.din(w_dff_A_JWom5X3a3_0),.clk(gclk));
	jdff dff_A_2HCW811z8_1(.dout(w_n614_0[1]),.din(w_dff_A_2HCW811z8_1),.clk(gclk));
	jdff dff_A_MGTmNajW1_1(.dout(w_dff_A_2HCW811z8_1),.din(w_dff_A_MGTmNajW1_1),.clk(gclk));
	jdff dff_A_O8HdHmMk5_2(.dout(w_n614_0[2]),.din(w_dff_A_O8HdHmMk5_2),.clk(gclk));
	jdff dff_A_e2wFTsdm5_2(.dout(w_dff_A_O8HdHmMk5_2),.din(w_dff_A_e2wFTsdm5_2),.clk(gclk));
	jdff dff_A_sDamZIWu9_2(.dout(w_dff_A_e2wFTsdm5_2),.din(w_dff_A_sDamZIWu9_2),.clk(gclk));
	jdff dff_A_HBGiEuX35_2(.dout(w_dff_A_sDamZIWu9_2),.din(w_dff_A_HBGiEuX35_2),.clk(gclk));
	jdff dff_B_rYGqbmNG0_1(.din(n610),.dout(w_dff_B_rYGqbmNG0_1),.clk(gclk));
	jdff dff_A_LT5SgMpK3_0(.dout(w_G332_4[0]),.din(w_dff_A_LT5SgMpK3_0),.clk(gclk));
	jdff dff_A_TWNRPvyV2_2(.dout(w_G332_1[2]),.din(w_dff_A_TWNRPvyV2_2),.clk(gclk));
	jdff dff_A_7Eb9Jmja7_1(.dout(w_G331_0[1]),.din(w_dff_A_7Eb9Jmja7_1),.clk(gclk));
	jdff dff_A_dWzcPerA0_0(.dout(w_n1391_0[0]),.din(w_dff_A_dWzcPerA0_0),.clk(gclk));
	jdff dff_A_CaI8okV65_0(.dout(w_dff_A_dWzcPerA0_0),.din(w_dff_A_CaI8okV65_0),.clk(gclk));
	jdff dff_A_3PmkaxBr7_0(.dout(w_dff_A_CaI8okV65_0),.din(w_dff_A_3PmkaxBr7_0),.clk(gclk));
	jdff dff_A_Sg7RcbN19_0(.dout(w_dff_A_3PmkaxBr7_0),.din(w_dff_A_Sg7RcbN19_0),.clk(gclk));
	jdff dff_A_rjwvY9S35_0(.dout(w_dff_A_Sg7RcbN19_0),.din(w_dff_A_rjwvY9S35_0),.clk(gclk));
	jdff dff_A_ydPM95mj5_0(.dout(w_dff_A_rjwvY9S35_0),.din(w_dff_A_ydPM95mj5_0),.clk(gclk));
	jdff dff_A_2zAA9Umb0_0(.dout(w_dff_A_ydPM95mj5_0),.din(w_dff_A_2zAA9Umb0_0),.clk(gclk));
	jdff dff_B_SQxsLgcW7_1(.din(n1389),.dout(w_dff_B_SQxsLgcW7_1),.clk(gclk));
	jdff dff_B_fwDQ9fKU8_1(.din(w_dff_B_SQxsLgcW7_1),.dout(w_dff_B_fwDQ9fKU8_1),.clk(gclk));
	jdff dff_A_u6mEIkBT1_1(.dout(w_G4091_1[1]),.din(w_dff_A_u6mEIkBT1_1),.clk(gclk));
	jdff dff_A_YprWSQXl2_1(.dout(w_dff_A_u6mEIkBT1_1),.din(w_dff_A_YprWSQXl2_1),.clk(gclk));
	jdff dff_A_UQf0Whvu4_1(.dout(w_dff_A_YprWSQXl2_1),.din(w_dff_A_UQf0Whvu4_1),.clk(gclk));
	jdff dff_A_8JQLu9eK9_1(.dout(w_dff_A_UQf0Whvu4_1),.din(w_dff_A_8JQLu9eK9_1),.clk(gclk));
	jdff dff_A_MkKKhlk65_1(.dout(w_dff_A_8JQLu9eK9_1),.din(w_dff_A_MkKKhlk65_1),.clk(gclk));
	jdff dff_A_u5EHQxMO5_1(.dout(w_dff_A_MkKKhlk65_1),.din(w_dff_A_u5EHQxMO5_1),.clk(gclk));
	jdff dff_A_LNrO9Vr24_1(.dout(w_dff_A_u5EHQxMO5_1),.din(w_dff_A_LNrO9Vr24_1),.clk(gclk));
	jdff dff_A_dRdZwZm91_1(.dout(w_dff_A_LNrO9Vr24_1),.din(w_dff_A_dRdZwZm91_1),.clk(gclk));
	jdff dff_A_sUXL1Gpm1_1(.dout(w_dff_A_dRdZwZm91_1),.din(w_dff_A_sUXL1Gpm1_1),.clk(gclk));
	jdff dff_A_PSud7I7X4_1(.dout(w_dff_A_sUXL1Gpm1_1),.din(w_dff_A_PSud7I7X4_1),.clk(gclk));
	jdff dff_A_2nGnnnYf9_1(.dout(w_dff_A_PSud7I7X4_1),.din(w_dff_A_2nGnnnYf9_1),.clk(gclk));
	jdff dff_A_nArJsp985_1(.dout(w_dff_A_2nGnnnYf9_1),.din(w_dff_A_nArJsp985_1),.clk(gclk));
	jdff dff_A_h6TM1nLb0_1(.dout(w_dff_A_nArJsp985_1),.din(w_dff_A_h6TM1nLb0_1),.clk(gclk));
	jdff dff_A_jl11dvRb3_1(.dout(w_dff_A_h6TM1nLb0_1),.din(w_dff_A_jl11dvRb3_1),.clk(gclk));
	jdff dff_A_BuIuQJ7E7_1(.dout(w_dff_A_jl11dvRb3_1),.din(w_dff_A_BuIuQJ7E7_1),.clk(gclk));
	jdff dff_A_mlFn4RIz5_1(.dout(w_dff_A_BuIuQJ7E7_1),.din(w_dff_A_mlFn4RIz5_1),.clk(gclk));
	jdff dff_A_mJUPKJal7_1(.dout(w_dff_A_mlFn4RIz5_1),.din(w_dff_A_mJUPKJal7_1),.clk(gclk));
	jdff dff_A_kLbvHeRq5_1(.dout(w_dff_A_mJUPKJal7_1),.din(w_dff_A_kLbvHeRq5_1),.clk(gclk));
	jdff dff_A_WWz6kItk5_2(.dout(w_G4091_1[2]),.din(w_dff_A_WWz6kItk5_2),.clk(gclk));
	jdff dff_A_yoTy8XiB6_2(.dout(w_dff_A_WWz6kItk5_2),.din(w_dff_A_yoTy8XiB6_2),.clk(gclk));
	jdff dff_A_FO2LjoWX8_2(.dout(w_dff_A_yoTy8XiB6_2),.din(w_dff_A_FO2LjoWX8_2),.clk(gclk));
	jdff dff_A_jRCz178b5_2(.dout(w_dff_A_FO2LjoWX8_2),.din(w_dff_A_jRCz178b5_2),.clk(gclk));
	jdff dff_A_H3iU3qlg3_2(.dout(w_dff_A_jRCz178b5_2),.din(w_dff_A_H3iU3qlg3_2),.clk(gclk));
	jdff dff_A_iDrou3bl9_2(.dout(w_dff_A_H3iU3qlg3_2),.din(w_dff_A_iDrou3bl9_2),.clk(gclk));
	jdff dff_A_DVM9SFrA2_2(.dout(w_dff_A_iDrou3bl9_2),.din(w_dff_A_DVM9SFrA2_2),.clk(gclk));
	jdff dff_A_bD7SVp1N3_2(.dout(w_dff_A_DVM9SFrA2_2),.din(w_dff_A_bD7SVp1N3_2),.clk(gclk));
	jdff dff_A_fxY25Nyx7_2(.dout(w_dff_A_bD7SVp1N3_2),.din(w_dff_A_fxY25Nyx7_2),.clk(gclk));
	jdff dff_A_m8eHBqdZ6_2(.dout(w_dff_A_fxY25Nyx7_2),.din(w_dff_A_m8eHBqdZ6_2),.clk(gclk));
	jdff dff_A_vJ2Onia90_0(.dout(w_n1383_0[0]),.din(w_dff_A_vJ2Onia90_0),.clk(gclk));
	jdff dff_A_fOBNq5Es2_0(.dout(w_dff_A_vJ2Onia90_0),.din(w_dff_A_fOBNq5Es2_0),.clk(gclk));
	jdff dff_B_khmYPcgz9_1(.din(n1363),.dout(w_dff_B_khmYPcgz9_1),.clk(gclk));
	jdff dff_B_Cn27TpIJ0_1(.din(w_dff_B_khmYPcgz9_1),.dout(w_dff_B_Cn27TpIJ0_1),.clk(gclk));
	jdff dff_B_rhIZik0W9_1(.din(n1376),.dout(w_dff_B_rhIZik0W9_1),.clk(gclk));
	jdff dff_B_kRJT3wse7_1(.din(n1377),.dout(w_dff_B_kRJT3wse7_1),.clk(gclk));
	jdff dff_A_7Lv7AdWl5_1(.dout(w_n426_0[1]),.din(w_dff_A_7Lv7AdWl5_1),.clk(gclk));
	jdff dff_A_ddU9OMzw0_0(.dout(w_G503_1[0]),.din(w_dff_A_ddU9OMzw0_0),.clk(gclk));
	jdff dff_A_VW1wU9Xh5_0(.dout(w_dff_A_ddU9OMzw0_0),.din(w_dff_A_VW1wU9Xh5_0),.clk(gclk));
	jdff dff_A_wK71iNMU8_0(.dout(w_dff_A_VW1wU9Xh5_0),.din(w_dff_A_wK71iNMU8_0),.clk(gclk));
	jdff dff_A_t8pGFjp86_0(.dout(w_dff_A_wK71iNMU8_0),.din(w_dff_A_t8pGFjp86_0),.clk(gclk));
	jdff dff_A_MIQ1Y4FX5_1(.dout(w_G503_1[1]),.din(w_dff_A_MIQ1Y4FX5_1),.clk(gclk));
	jdff dff_A_THHCLd8W5_1(.dout(w_G503_0[1]),.din(w_dff_A_THHCLd8W5_1),.clk(gclk));
	jdff dff_A_uvjxOwaX1_1(.dout(w_dff_A_THHCLd8W5_1),.din(w_dff_A_uvjxOwaX1_1),.clk(gclk));
	jdff dff_A_C7If0JOz7_2(.dout(w_G503_0[2]),.din(w_dff_A_C7If0JOz7_2),.clk(gclk));
	jdff dff_A_y0LvTvBl1_2(.dout(w_dff_A_C7If0JOz7_2),.din(w_dff_A_y0LvTvBl1_2),.clk(gclk));
	jdff dff_A_TIFXSPOy5_2(.dout(w_dff_A_y0LvTvBl1_2),.din(w_dff_A_TIFXSPOy5_2),.clk(gclk));
	jdff dff_A_Pru7XwWy6_2(.dout(w_dff_A_TIFXSPOy5_2),.din(w_dff_A_Pru7XwWy6_2),.clk(gclk));
	jdff dff_A_2TCoX7101_1(.dout(w_G324_1[1]),.din(w_dff_A_2TCoX7101_1),.clk(gclk));
	jdff dff_A_o35FUYa91_1(.dout(w_G324_0[1]),.din(w_dff_A_o35FUYa91_1),.clk(gclk));
	jdff dff_B_j3XPcoFH2_1(.din(n1368),.dout(w_dff_B_j3XPcoFH2_1),.clk(gclk));
	jdff dff_B_5XAEIhWx1_1(.din(w_dff_B_j3XPcoFH2_1),.dout(w_dff_B_5XAEIhWx1_1),.clk(gclk));
	jdff dff_A_x1spk4jM5_2(.dout(w_n388_0[2]),.din(w_dff_A_x1spk4jM5_2),.clk(gclk));
	jdff dff_B_Q4dSipxa8_3(.din(n388),.dout(w_dff_B_Q4dSipxa8_3),.clk(gclk));
	jdff dff_A_5nmcFANn6_0(.dout(w_G534_1[0]),.din(w_dff_A_5nmcFANn6_0),.clk(gclk));
	jdff dff_A_gEgy98RR2_0(.dout(w_dff_A_5nmcFANn6_0),.din(w_dff_A_gEgy98RR2_0),.clk(gclk));
	jdff dff_A_hFq9wJpJ8_0(.dout(w_dff_A_gEgy98RR2_0),.din(w_dff_A_hFq9wJpJ8_0),.clk(gclk));
	jdff dff_A_5qhikpfe9_1(.dout(w_G534_1[1]),.din(w_dff_A_5qhikpfe9_1),.clk(gclk));
	jdff dff_B_aWUAzN4U2_1(.din(n1364),.dout(w_dff_B_aWUAzN4U2_1),.clk(gclk));
	jdff dff_A_kJ1VNvQG9_1(.dout(w_G351_2[1]),.din(w_dff_A_kJ1VNvQG9_1),.clk(gclk));
	jdff dff_A_cvrUomGe6_1(.dout(w_G534_0[1]),.din(w_dff_A_cvrUomGe6_1),.clk(gclk));
	jdff dff_A_1OY5sP727_1(.dout(w_dff_A_cvrUomGe6_1),.din(w_dff_A_1OY5sP727_1),.clk(gclk));
	jdff dff_A_VidaYrBB3_2(.dout(w_G534_0[2]),.din(w_dff_A_VidaYrBB3_2),.clk(gclk));
	jdff dff_A_xiyzJKe73_2(.dout(w_dff_A_VidaYrBB3_2),.din(w_dff_A_xiyzJKe73_2),.clk(gclk));
	jdff dff_A_0pFK2Ner1_2(.dout(w_dff_A_xiyzJKe73_2),.din(w_dff_A_0pFK2Ner1_2),.clk(gclk));
	jdff dff_A_OglsVBYO9_0(.dout(w_G351_1[0]),.din(w_dff_A_OglsVBYO9_0),.clk(gclk));
	jdff dff_A_Rtj5CWw78_2(.dout(w_n410_0[2]),.din(w_dff_A_Rtj5CWw78_2),.clk(gclk));
	jdff dff_A_6st0OpoW4_1(.dout(w_G514_0[1]),.din(w_dff_A_6st0OpoW4_1),.clk(gclk));
	jdff dff_A_FlZ0ONBZ3_2(.dout(w_G514_0[2]),.din(w_dff_A_FlZ0ONBZ3_2),.clk(gclk));
	jdff dff_A_rhNxgrBE4_2(.dout(w_dff_A_FlZ0ONBZ3_2),.din(w_dff_A_rhNxgrBE4_2),.clk(gclk));
	jdff dff_A_iMsQLFAt3_1(.dout(w_G361_0[1]),.din(w_dff_A_iMsQLFAt3_1),.clk(gclk));
	jdff dff_B_TBo6RMLm5_1(.din(n1354),.dout(w_dff_B_TBo6RMLm5_1),.clk(gclk));
	jdff dff_B_Ywm0ecfJ3_1(.din(w_dff_B_TBo6RMLm5_1),.dout(w_dff_B_Ywm0ecfJ3_1),.clk(gclk));
	jdff dff_B_lAeKIlEP8_1(.din(n1355),.dout(w_dff_B_lAeKIlEP8_1),.clk(gclk));
	jdff dff_B_Nsmg6kdC0_1(.din(n378),.dout(w_dff_B_Nsmg6kdC0_1),.clk(gclk));
	jdff dff_B_HrGeroVV9_1(.din(n379),.dout(w_dff_B_HrGeroVV9_1),.clk(gclk));
	jdff dff_A_T7u7M1HZ3_0(.dout(w_G490_1[0]),.din(w_dff_A_T7u7M1HZ3_0),.clk(gclk));
	jdff dff_A_TiknX4FY5_0(.dout(w_dff_A_T7u7M1HZ3_0),.din(w_dff_A_TiknX4FY5_0),.clk(gclk));
	jdff dff_A_4rgexoVy5_0(.dout(w_dff_A_TiknX4FY5_0),.din(w_dff_A_4rgexoVy5_0),.clk(gclk));
	jdff dff_A_FWhTANMH7_1(.dout(w_G490_1[1]),.din(w_dff_A_FWhTANMH7_1),.clk(gclk));
	jdff dff_A_sGs16ISw7_1(.dout(w_dff_A_FWhTANMH7_1),.din(w_dff_A_sGs16ISw7_1),.clk(gclk));
	jdff dff_A_yhl7EdmH5_1(.dout(w_G490_0[1]),.din(w_dff_A_yhl7EdmH5_1),.clk(gclk));
	jdff dff_A_gzcDVFSt0_1(.dout(w_dff_A_yhl7EdmH5_1),.din(w_dff_A_gzcDVFSt0_1),.clk(gclk));
	jdff dff_A_eREKj2st1_1(.dout(w_dff_A_gzcDVFSt0_1),.din(w_dff_A_eREKj2st1_1),.clk(gclk));
	jdff dff_A_LAxhXHmZ7_2(.dout(w_G490_0[2]),.din(w_dff_A_LAxhXHmZ7_2),.clk(gclk));
	jdff dff_A_fTEYH5MJ3_2(.dout(w_dff_A_LAxhXHmZ7_2),.din(w_dff_A_fTEYH5MJ3_2),.clk(gclk));
	jdff dff_A_4J7QjujL1_2(.dout(w_dff_A_fTEYH5MJ3_2),.din(w_dff_A_4J7QjujL1_2),.clk(gclk));
	jdff dff_A_msxUPXKl5_0(.dout(w_G316_1[0]),.din(w_dff_A_msxUPXKl5_0),.clk(gclk));
	jdff dff_B_DYaX8Hgu3_1(.din(n365),.dout(w_dff_B_DYaX8Hgu3_1),.clk(gclk));
	jdff dff_B_Ad7FIs4t6_1(.din(n367),.dout(w_dff_B_Ad7FIs4t6_1),.clk(gclk));
	jdff dff_A_HqRQQ5Dw3_0(.dout(w_n362_0[0]),.din(w_dff_A_HqRQQ5Dw3_0),.clk(gclk));
	jdff dff_A_v2PmSzza2_0(.dout(w_dff_A_HqRQQ5Dw3_0),.din(w_dff_A_v2PmSzza2_0),.clk(gclk));
	jdff dff_A_RvHiWXFc7_0(.dout(w_dff_A_v2PmSzza2_0),.din(w_dff_A_RvHiWXFc7_0),.clk(gclk));
	jdff dff_A_V2gQG1eZ7_0(.dout(w_G479_1[0]),.din(w_dff_A_V2gQG1eZ7_0),.clk(gclk));
	jdff dff_A_MvzDF7Oj4_0(.dout(w_dff_A_V2gQG1eZ7_0),.din(w_dff_A_MvzDF7Oj4_0),.clk(gclk));
	jdff dff_A_C5PijlUF7_1(.dout(w_G479_0[1]),.din(w_dff_A_C5PijlUF7_1),.clk(gclk));
	jdff dff_A_GTBQ4FCe4_1(.dout(w_dff_A_C5PijlUF7_1),.din(w_dff_A_GTBQ4FCe4_1),.clk(gclk));
	jdff dff_A_1kxmuCHH2_1(.dout(w_dff_A_GTBQ4FCe4_1),.din(w_dff_A_1kxmuCHH2_1),.clk(gclk));
	jdff dff_A_DtmHDySL8_2(.dout(w_G479_0[2]),.din(w_dff_A_DtmHDySL8_2),.clk(gclk));
	jdff dff_A_swKeyPw01_2(.dout(w_dff_A_DtmHDySL8_2),.din(w_dff_A_swKeyPw01_2),.clk(gclk));
	jdff dff_A_5hM7wWQg4_2(.dout(w_dff_A_swKeyPw01_2),.din(w_dff_A_5hM7wWQg4_2),.clk(gclk));
	jdff dff_A_77KRC1lc4_0(.dout(w_G308_1[0]),.din(w_dff_A_77KRC1lc4_0),.clk(gclk));
	jdff dff_A_4NWISi2H3_0(.dout(w_G302_0[0]),.din(w_dff_A_4NWISi2H3_0),.clk(gclk));
	jdff dff_A_j41D3iUL7_1(.dout(w_G302_0[1]),.din(w_dff_A_j41D3iUL7_1),.clk(gclk));
	jdff dff_A_9RxrP5xD1_0(.dout(w_n401_0[0]),.din(w_dff_A_9RxrP5xD1_0),.clk(gclk));
	jdff dff_A_USqn9juS4_2(.dout(w_n401_0[2]),.din(w_dff_A_USqn9juS4_2),.clk(gclk));
	jdff dff_A_rU5hIRg20_1(.dout(w_G293_0[1]),.din(w_dff_A_rU5hIRg20_1),.clk(gclk));
	jdff dff_B_a2v8VoHg4_1(.din(n1349),.dout(w_dff_B_a2v8VoHg4_1),.clk(gclk));
	jdff dff_B_nc06qPDF0_1(.din(n1350),.dout(w_dff_B_nc06qPDF0_1),.clk(gclk));
	jdff dff_A_X8JEPTvo8_0(.dout(w_n437_0[0]),.din(w_dff_A_X8JEPTvo8_0),.clk(gclk));
	jdff dff_A_SLhPDG6J2_2(.dout(w_n437_0[2]),.din(w_dff_A_SLhPDG6J2_2),.clk(gclk));
	jdff dff_A_rVsBUueX2_2(.dout(w_dff_A_SLhPDG6J2_2),.din(w_dff_A_rVsBUueX2_2),.clk(gclk));
	jdff dff_A_QGecVUIb6_0(.dout(w_G523_1[0]),.din(w_dff_A_QGecVUIb6_0),.clk(gclk));
	jdff dff_A_92YtTzxb0_1(.dout(w_G523_0[1]),.din(w_dff_A_92YtTzxb0_1),.clk(gclk));
	jdff dff_A_6KjX17et2_1(.dout(w_dff_A_92YtTzxb0_1),.din(w_dff_A_6KjX17et2_1),.clk(gclk));
	jdff dff_A_6PiK53K50_1(.dout(w_dff_A_6KjX17et2_1),.din(w_dff_A_6PiK53K50_1),.clk(gclk));
	jdff dff_A_RDUmUsws8_2(.dout(w_G523_0[2]),.din(w_dff_A_RDUmUsws8_2),.clk(gclk));
	jdff dff_A_zDMoByYg7_2(.dout(w_dff_A_RDUmUsws8_2),.din(w_dff_A_zDMoByYg7_2),.clk(gclk));
	jdff dff_A_bcnZ5QXg4_1(.dout(w_G341_2[1]),.din(w_dff_A_bcnZ5QXg4_1),.clk(gclk));
	jdff dff_A_8Kvxk1sW7_2(.dout(w_G341_0[2]),.din(w_dff_A_8Kvxk1sW7_2),.clk(gclk));
	jdff dff_A_aze7x1926_2(.dout(w_n746_0[2]),.din(w_dff_A_aze7x1926_2),.clk(gclk));
	jdff dff_A_pFPTIqm75_2(.dout(w_dff_A_aze7x1926_2),.din(w_dff_A_pFPTIqm75_2),.clk(gclk));
	jdff dff_A_uZpT0iYG7_2(.dout(w_dff_A_pFPTIqm75_2),.din(w_dff_A_uZpT0iYG7_2),.clk(gclk));
	jdff dff_A_hvkmYb9T5_2(.dout(w_dff_A_uZpT0iYG7_2),.din(w_dff_A_hvkmYb9T5_2),.clk(gclk));
	jdff dff_A_W4QeQyRj1_2(.dout(w_dff_A_hvkmYb9T5_2),.din(w_dff_A_W4QeQyRj1_2),.clk(gclk));
	jdff dff_A_yBmEkHR52_2(.dout(w_dff_A_W4QeQyRj1_2),.din(w_dff_A_yBmEkHR52_2),.clk(gclk));
	jdff dff_A_ph5qFrFO9_2(.dout(w_dff_A_yBmEkHR52_2),.din(w_dff_A_ph5qFrFO9_2),.clk(gclk));
	jdff dff_A_q9xs8aBf7_2(.dout(w_dff_A_ph5qFrFO9_2),.din(w_dff_A_q9xs8aBf7_2),.clk(gclk));
	jdff dff_A_IW8s2snX7_2(.dout(w_dff_A_q9xs8aBf7_2),.din(w_dff_A_IW8s2snX7_2),.clk(gclk));
	jdff dff_A_rxs8mDsb4_2(.dout(w_dff_A_IW8s2snX7_2),.din(w_dff_A_rxs8mDsb4_2),.clk(gclk));
	jdff dff_A_xCoe0Yxo1_2(.dout(w_dff_A_rxs8mDsb4_2),.din(w_dff_A_xCoe0Yxo1_2),.clk(gclk));
	jdff dff_A_NLKlnGtd4_0(.dout(w_n1002_1[0]),.din(w_dff_A_NLKlnGtd4_0),.clk(gclk));
	jdff dff_A_HYLUqFkp4_0(.dout(w_dff_A_NLKlnGtd4_0),.din(w_dff_A_HYLUqFkp4_0),.clk(gclk));
	jdff dff_A_GYLgjmw42_0(.dout(w_dff_A_HYLUqFkp4_0),.din(w_dff_A_GYLgjmw42_0),.clk(gclk));
	jdff dff_A_nm9NQ2Pf3_0(.dout(w_dff_A_GYLgjmw42_0),.din(w_dff_A_nm9NQ2Pf3_0),.clk(gclk));
	jdff dff_A_EfLg9am28_0(.dout(w_dff_A_nm9NQ2Pf3_0),.din(w_dff_A_EfLg9am28_0),.clk(gclk));
	jdff dff_A_LW7Mt9wV8_0(.dout(w_dff_A_EfLg9am28_0),.din(w_dff_A_LW7Mt9wV8_0),.clk(gclk));
	jdff dff_A_7eioFKEk0_2(.dout(w_n1002_1[2]),.din(w_dff_A_7eioFKEk0_2),.clk(gclk));
	jdff dff_A_ZuuYbSaV3_2(.dout(w_dff_A_7eioFKEk0_2),.din(w_dff_A_ZuuYbSaV3_2),.clk(gclk));
	jdff dff_A_h1nyXclN6_2(.dout(w_dff_A_ZuuYbSaV3_2),.din(w_dff_A_h1nyXclN6_2),.clk(gclk));
	jdff dff_A_fdlHF7ir3_2(.dout(w_dff_A_h1nyXclN6_2),.din(w_dff_A_fdlHF7ir3_2),.clk(gclk));
	jdff dff_A_HZ5IFSO28_2(.dout(w_dff_A_fdlHF7ir3_2),.din(w_dff_A_HZ5IFSO28_2),.clk(gclk));
	jdff dff_A_KF45V0xS4_2(.dout(w_dff_A_HZ5IFSO28_2),.din(w_dff_A_KF45V0xS4_2),.clk(gclk));
	jdff dff_A_bISymSaK6_2(.dout(w_dff_A_KF45V0xS4_2),.din(w_dff_A_bISymSaK6_2),.clk(gclk));
	jdff dff_A_taQFjGuE7_2(.dout(w_dff_A_bISymSaK6_2),.din(w_dff_A_taQFjGuE7_2),.clk(gclk));
	jdff dff_A_Voo3CxCM6_2(.dout(w_dff_A_taQFjGuE7_2),.din(w_dff_A_Voo3CxCM6_2),.clk(gclk));
	jdff dff_A_ND6PrY139_2(.dout(w_dff_A_Voo3CxCM6_2),.din(w_dff_A_ND6PrY139_2),.clk(gclk));
	jdff dff_A_Z9p8ucLv1_2(.dout(w_dff_A_ND6PrY139_2),.din(w_dff_A_Z9p8ucLv1_2),.clk(gclk));
	jdff dff_A_AIgbrBNr3_2(.dout(w_dff_A_Z9p8ucLv1_2),.din(w_dff_A_AIgbrBNr3_2),.clk(gclk));
	jdff dff_A_xLgZBadQ1_2(.dout(w_dff_A_AIgbrBNr3_2),.din(w_dff_A_xLgZBadQ1_2),.clk(gclk));
	jdff dff_A_RW3szw4Z4_2(.dout(w_dff_A_xLgZBadQ1_2),.din(w_dff_A_RW3szw4Z4_2),.clk(gclk));
	jdff dff_A_IjIs24Tj0_2(.dout(w_dff_A_RW3szw4Z4_2),.din(w_dff_A_IjIs24Tj0_2),.clk(gclk));
	jdff dff_A_kW6BxD995_2(.dout(w_dff_A_IjIs24Tj0_2),.din(w_dff_A_kW6BxD995_2),.clk(gclk));
	jdff dff_A_Ytz3WvXx7_2(.dout(w_dff_A_kW6BxD995_2),.din(w_dff_A_Ytz3WvXx7_2),.clk(gclk));
	jdff dff_A_IDxTqGVC1_2(.dout(w_dff_A_Ytz3WvXx7_2),.din(w_dff_A_IDxTqGVC1_2),.clk(gclk));
	jdff dff_A_Deyg2NPH8_1(.dout(w_n1002_0[1]),.din(w_dff_A_Deyg2NPH8_1),.clk(gclk));
	jdff dff_A_RMquG1VH5_1(.dout(w_dff_A_Deyg2NPH8_1),.din(w_dff_A_RMquG1VH5_1),.clk(gclk));
	jdff dff_A_qAkVl2KR2_1(.dout(w_dff_A_RMquG1VH5_1),.din(w_dff_A_qAkVl2KR2_1),.clk(gclk));
	jdff dff_A_S8Q5VEb37_1(.dout(w_dff_A_qAkVl2KR2_1),.din(w_dff_A_S8Q5VEb37_1),.clk(gclk));
	jdff dff_A_iGo2aX4h1_1(.dout(w_dff_A_S8Q5VEb37_1),.din(w_dff_A_iGo2aX4h1_1),.clk(gclk));
	jdff dff_A_QldryrM18_1(.dout(w_dff_A_iGo2aX4h1_1),.din(w_dff_A_QldryrM18_1),.clk(gclk));
	jdff dff_A_OmHXET6u8_1(.dout(w_dff_A_QldryrM18_1),.din(w_dff_A_OmHXET6u8_1),.clk(gclk));
	jdff dff_A_afAF2FrS8_1(.dout(w_dff_A_OmHXET6u8_1),.din(w_dff_A_afAF2FrS8_1),.clk(gclk));
	jdff dff_A_zWIkN5RY2_1(.dout(w_dff_A_afAF2FrS8_1),.din(w_dff_A_zWIkN5RY2_1),.clk(gclk));
	jdff dff_A_2CqVssKs0_1(.dout(w_dff_A_zWIkN5RY2_1),.din(w_dff_A_2CqVssKs0_1),.clk(gclk));
	jdff dff_A_JreCyYxF9_1(.dout(w_dff_A_2CqVssKs0_1),.din(w_dff_A_JreCyYxF9_1),.clk(gclk));
	jdff dff_A_wYxPPXOo4_1(.dout(w_dff_A_JreCyYxF9_1),.din(w_dff_A_wYxPPXOo4_1),.clk(gclk));
	jdff dff_A_7aE8ig800_1(.dout(w_dff_A_wYxPPXOo4_1),.din(w_dff_A_7aE8ig800_1),.clk(gclk));
	jdff dff_A_TH0PPm387_1(.dout(w_dff_A_7aE8ig800_1),.din(w_dff_A_TH0PPm387_1),.clk(gclk));
	jdff dff_A_zOfvnnl55_1(.dout(w_dff_A_TH0PPm387_1),.din(w_dff_A_zOfvnnl55_1),.clk(gclk));
	jdff dff_A_32D0wbyv8_1(.dout(w_dff_A_zOfvnnl55_1),.din(w_dff_A_32D0wbyv8_1),.clk(gclk));
	jdff dff_A_wsDP1bJN1_2(.dout(w_n1002_0[2]),.din(w_dff_A_wsDP1bJN1_2),.clk(gclk));
	jdff dff_A_QRo3H8Pp1_2(.dout(w_dff_A_wsDP1bJN1_2),.din(w_dff_A_QRo3H8Pp1_2),.clk(gclk));
	jdff dff_A_jk0adFD75_2(.dout(w_dff_A_QRo3H8Pp1_2),.din(w_dff_A_jk0adFD75_2),.clk(gclk));
	jdff dff_A_FaY6W2PO3_2(.dout(w_dff_A_jk0adFD75_2),.din(w_dff_A_FaY6W2PO3_2),.clk(gclk));
	jdff dff_A_xchrOceB9_2(.dout(w_dff_A_FaY6W2PO3_2),.din(w_dff_A_xchrOceB9_2),.clk(gclk));
	jdff dff_A_SA6K04Ui8_2(.dout(w_dff_A_xchrOceB9_2),.din(w_dff_A_SA6K04Ui8_2),.clk(gclk));
	jdff dff_A_wXW4sHwz1_2(.dout(w_dff_A_SA6K04Ui8_2),.din(w_dff_A_wXW4sHwz1_2),.clk(gclk));
	jdff dff_B_D0CWybsJ3_1(.din(n1641),.dout(w_dff_B_D0CWybsJ3_1),.clk(gclk));
	jdff dff_B_E9pVTg2h6_1(.din(w_dff_B_D0CWybsJ3_1),.dout(w_dff_B_E9pVTg2h6_1),.clk(gclk));
	jdff dff_B_gYfskHur3_1(.din(w_dff_B_E9pVTg2h6_1),.dout(w_dff_B_gYfskHur3_1),.clk(gclk));
	jdff dff_B_iYhTyRRk3_1(.din(w_dff_B_gYfskHur3_1),.dout(w_dff_B_iYhTyRRk3_1),.clk(gclk));
	jdff dff_B_Wik5T94l9_1(.din(w_dff_B_iYhTyRRk3_1),.dout(w_dff_B_Wik5T94l9_1),.clk(gclk));
	jdff dff_B_f7yEEDOe6_1(.din(w_dff_B_Wik5T94l9_1),.dout(w_dff_B_f7yEEDOe6_1),.clk(gclk));
	jdff dff_B_YNReeq394_1(.din(w_dff_B_f7yEEDOe6_1),.dout(w_dff_B_YNReeq394_1),.clk(gclk));
	jdff dff_B_266Bsybs0_1(.din(w_dff_B_YNReeq394_1),.dout(w_dff_B_266Bsybs0_1),.clk(gclk));
	jdff dff_B_U7qNGUDw4_1(.din(w_dff_B_266Bsybs0_1),.dout(w_dff_B_U7qNGUDw4_1),.clk(gclk));
	jdff dff_B_w8H034wv6_1(.din(w_dff_B_U7qNGUDw4_1),.dout(w_dff_B_w8H034wv6_1),.clk(gclk));
	jdff dff_B_obFN7baq1_1(.din(w_dff_B_w8H034wv6_1),.dout(w_dff_B_obFN7baq1_1),.clk(gclk));
	jdff dff_B_KqzyrakD9_1(.din(w_dff_B_obFN7baq1_1),.dout(w_dff_B_KqzyrakD9_1),.clk(gclk));
	jdff dff_B_qhIFKDUt1_1(.din(w_dff_B_KqzyrakD9_1),.dout(w_dff_B_qhIFKDUt1_1),.clk(gclk));
	jdff dff_B_403AIYZk7_1(.din(w_dff_B_qhIFKDUt1_1),.dout(w_dff_B_403AIYZk7_1),.clk(gclk));
	jdff dff_B_on9cbfOZ0_1(.din(w_dff_B_403AIYZk7_1),.dout(w_dff_B_on9cbfOZ0_1),.clk(gclk));
	jdff dff_B_AvbfHbsE0_1(.din(w_dff_B_on9cbfOZ0_1),.dout(w_dff_B_AvbfHbsE0_1),.clk(gclk));
	jdff dff_B_3cmqoIzR5_1(.din(w_dff_B_AvbfHbsE0_1),.dout(w_dff_B_3cmqoIzR5_1),.clk(gclk));
	jdff dff_B_BhU5I1SB5_1(.din(w_dff_B_3cmqoIzR5_1),.dout(w_dff_B_BhU5I1SB5_1),.clk(gclk));
	jdff dff_B_y6t5PHBq2_1(.din(w_dff_B_BhU5I1SB5_1),.dout(w_dff_B_y6t5PHBq2_1),.clk(gclk));
	jdff dff_B_m9RvD3KT2_0(.din(n1600),.dout(w_dff_B_m9RvD3KT2_0),.clk(gclk));
	jdff dff_B_bAjPbLHg5_0(.din(w_dff_B_m9RvD3KT2_0),.dout(w_dff_B_bAjPbLHg5_0),.clk(gclk));
	jdff dff_B_t283aIEp3_0(.din(w_dff_B_bAjPbLHg5_0),.dout(w_dff_B_t283aIEp3_0),.clk(gclk));
	jdff dff_B_07k7FyeT2_0(.din(w_dff_B_t283aIEp3_0),.dout(w_dff_B_07k7FyeT2_0),.clk(gclk));
	jdff dff_B_K80B8jMO0_0(.din(w_dff_B_07k7FyeT2_0),.dout(w_dff_B_K80B8jMO0_0),.clk(gclk));
	jdff dff_B_rThIxeqp0_0(.din(w_dff_B_K80B8jMO0_0),.dout(w_dff_B_rThIxeqp0_0),.clk(gclk));
	jdff dff_B_kbljello1_0(.din(w_dff_B_rThIxeqp0_0),.dout(w_dff_B_kbljello1_0),.clk(gclk));
	jdff dff_B_sqNmiUWR4_0(.din(w_dff_B_kbljello1_0),.dout(w_dff_B_sqNmiUWR4_0),.clk(gclk));
	jdff dff_B_oeJrBfkf2_0(.din(w_dff_B_sqNmiUWR4_0),.dout(w_dff_B_oeJrBfkf2_0),.clk(gclk));
	jdff dff_B_dj564phh1_0(.din(w_dff_B_oeJrBfkf2_0),.dout(w_dff_B_dj564phh1_0),.clk(gclk));
	jdff dff_B_eg3XnDXj7_0(.din(w_dff_B_dj564phh1_0),.dout(w_dff_B_eg3XnDXj7_0),.clk(gclk));
	jdff dff_B_ruonKnZQ4_0(.din(w_dff_B_eg3XnDXj7_0),.dout(w_dff_B_ruonKnZQ4_0),.clk(gclk));
	jdff dff_B_jZD2Stwo6_0(.din(w_dff_B_ruonKnZQ4_0),.dout(w_dff_B_jZD2Stwo6_0),.clk(gclk));
	jdff dff_B_sb0Pk6hN5_0(.din(w_dff_B_jZD2Stwo6_0),.dout(w_dff_B_sb0Pk6hN5_0),.clk(gclk));
	jdff dff_B_55jthq2E1_0(.din(w_dff_B_sb0Pk6hN5_0),.dout(w_dff_B_55jthq2E1_0),.clk(gclk));
	jdff dff_B_qSjIQnq75_0(.din(w_dff_B_55jthq2E1_0),.dout(w_dff_B_qSjIQnq75_0),.clk(gclk));
	jdff dff_B_ZCNmBO4p3_0(.din(w_dff_B_qSjIQnq75_0),.dout(w_dff_B_ZCNmBO4p3_0),.clk(gclk));
	jdff dff_B_bcAW2MU46_0(.din(w_dff_B_ZCNmBO4p3_0),.dout(w_dff_B_bcAW2MU46_0),.clk(gclk));
	jdff dff_B_CczamCeA6_0(.din(w_dff_B_bcAW2MU46_0),.dout(w_dff_B_CczamCeA6_0),.clk(gclk));
	jdff dff_B_y6eSBI4b3_1(.din(n1540),.dout(w_dff_B_y6eSBI4b3_1),.clk(gclk));
	jdff dff_B_cybQlxok1_1(.din(w_dff_B_y6eSBI4b3_1),.dout(w_dff_B_cybQlxok1_1),.clk(gclk));
	jdff dff_B_71f4yUDK4_1(.din(w_dff_B_cybQlxok1_1),.dout(w_dff_B_71f4yUDK4_1),.clk(gclk));
	jdff dff_B_cMGm7CZg8_1(.din(w_dff_B_71f4yUDK4_1),.dout(w_dff_B_cMGm7CZg8_1),.clk(gclk));
	jdff dff_B_5OhrnJ7w7_1(.din(w_dff_B_cMGm7CZg8_1),.dout(w_dff_B_5OhrnJ7w7_1),.clk(gclk));
	jdff dff_B_cEHmt6JV6_1(.din(w_dff_B_5OhrnJ7w7_1),.dout(w_dff_B_cEHmt6JV6_1),.clk(gclk));
	jdff dff_B_SSdPyBsD3_1(.din(w_dff_B_cEHmt6JV6_1),.dout(w_dff_B_SSdPyBsD3_1),.clk(gclk));
	jdff dff_B_JxnJFHBJ9_1(.din(w_dff_B_SSdPyBsD3_1),.dout(w_dff_B_JxnJFHBJ9_1),.clk(gclk));
	jdff dff_B_voDq9m3C7_0(.din(n1589),.dout(w_dff_B_voDq9m3C7_0),.clk(gclk));
	jdff dff_B_OBkh3hor7_0(.din(w_dff_B_voDq9m3C7_0),.dout(w_dff_B_OBkh3hor7_0),.clk(gclk));
	jdff dff_B_Y0KUzQp49_1(.din(n1579),.dout(w_dff_B_Y0KUzQp49_1),.clk(gclk));
	jdff dff_B_fDgFNn5p1_0(.din(n1586),.dout(w_dff_B_fDgFNn5p1_0),.clk(gclk));
	jdff dff_B_HmHRIsmj7_0(.din(w_dff_B_fDgFNn5p1_0),.dout(w_dff_B_HmHRIsmj7_0),.clk(gclk));
	jdff dff_B_13uFmaH52_0(.din(w_dff_B_HmHRIsmj7_0),.dout(w_dff_B_13uFmaH52_0),.clk(gclk));
	jdff dff_B_8LDZHcFf0_0(.din(n1584),.dout(w_dff_B_8LDZHcFf0_0),.clk(gclk));
	jdff dff_B_oHymJl9Z4_1(.din(n1567),.dout(w_dff_B_oHymJl9Z4_1),.clk(gclk));
	jdff dff_B_p0OjHqQ14_1(.din(w_dff_B_oHymJl9Z4_1),.dout(w_dff_B_p0OjHqQ14_1),.clk(gclk));
	jdff dff_B_Oo98Fwqg2_1(.din(w_dff_B_p0OjHqQ14_1),.dout(w_dff_B_Oo98Fwqg2_1),.clk(gclk));
	jdff dff_B_hvQyuDWe6_1(.din(w_dff_B_Oo98Fwqg2_1),.dout(w_dff_B_hvQyuDWe6_1),.clk(gclk));
	jdff dff_B_kfga65Hg1_1(.din(w_dff_B_hvQyuDWe6_1),.dout(w_dff_B_kfga65Hg1_1),.clk(gclk));
	jdff dff_B_oKx2tdWk3_1(.din(w_dff_B_kfga65Hg1_1),.dout(w_dff_B_oKx2tdWk3_1),.clk(gclk));
	jdff dff_B_s6FttiPF9_1(.din(w_dff_B_oKx2tdWk3_1),.dout(w_dff_B_s6FttiPF9_1),.clk(gclk));
	jdff dff_B_BK8bDYqc8_1(.din(w_dff_B_s6FttiPF9_1),.dout(w_dff_B_BK8bDYqc8_1),.clk(gclk));
	jdff dff_B_NRoWvbCT3_1(.din(w_dff_B_BK8bDYqc8_1),.dout(w_dff_B_NRoWvbCT3_1),.clk(gclk));
	jdff dff_B_zJkuUrqE1_1(.din(w_dff_B_NRoWvbCT3_1),.dout(w_dff_B_zJkuUrqE1_1),.clk(gclk));
	jdff dff_B_CPYGXWMg6_1(.din(w_dff_B_zJkuUrqE1_1),.dout(w_dff_B_CPYGXWMg6_1),.clk(gclk));
	jdff dff_B_gm7OfTpl8_1(.din(w_dff_B_CPYGXWMg6_1),.dout(w_dff_B_gm7OfTpl8_1),.clk(gclk));
	jdff dff_B_KRgvwtkw4_1(.din(w_dff_B_gm7OfTpl8_1),.dout(w_dff_B_KRgvwtkw4_1),.clk(gclk));
	jdff dff_B_TWtG4G4Q2_1(.din(n1570),.dout(w_dff_B_TWtG4G4Q2_1),.clk(gclk));
	jdff dff_B_m5YzHZ2X8_1(.din(w_dff_B_TWtG4G4Q2_1),.dout(w_dff_B_m5YzHZ2X8_1),.clk(gclk));
	jdff dff_B_WWxDy1XO9_1(.din(w_dff_B_m5YzHZ2X8_1),.dout(w_dff_B_WWxDy1XO9_1),.clk(gclk));
	jdff dff_B_ZEHe0Y898_1(.din(w_dff_B_WWxDy1XO9_1),.dout(w_dff_B_ZEHe0Y898_1),.clk(gclk));
	jdff dff_B_NyEhML011_1(.din(n1571),.dout(w_dff_B_NyEhML011_1),.clk(gclk));
	jdff dff_B_8v8wTRNY5_1(.din(w_dff_B_NyEhML011_1),.dout(w_dff_B_8v8wTRNY5_1),.clk(gclk));
	jdff dff_B_PtQ18N2B6_1(.din(w_dff_B_8v8wTRNY5_1),.dout(w_dff_B_PtQ18N2B6_1),.clk(gclk));
	jdff dff_B_XIfNXhkf4_1(.din(w_dff_B_PtQ18N2B6_1),.dout(w_dff_B_XIfNXhkf4_1),.clk(gclk));
	jdff dff_B_GIHZRyBw4_1(.din(w_dff_B_XIfNXhkf4_1),.dout(w_dff_B_GIHZRyBw4_1),.clk(gclk));
	jdff dff_B_LvevyD0u7_1(.din(w_dff_B_GIHZRyBw4_1),.dout(w_dff_B_LvevyD0u7_1),.clk(gclk));
	jdff dff_A_hEsPBp8w3_0(.dout(w_n855_0[0]),.din(w_dff_A_hEsPBp8w3_0),.clk(gclk));
	jdff dff_A_1lupsNG66_1(.dout(w_n853_0[1]),.din(w_dff_A_1lupsNG66_1),.clk(gclk));
	jdff dff_B_MtLqDPHt3_2(.din(n853),.dout(w_dff_B_MtLqDPHt3_2),.clk(gclk));
	jdff dff_B_Br1j1YCb7_2(.din(w_dff_B_MtLqDPHt3_2),.dout(w_dff_B_Br1j1YCb7_2),.clk(gclk));
	jdff dff_B_jurjrizg7_2(.din(w_dff_B_Br1j1YCb7_2),.dout(w_dff_B_jurjrizg7_2),.clk(gclk));
	jdff dff_B_kllcc4En5_2(.din(w_dff_B_jurjrizg7_2),.dout(w_dff_B_kllcc4En5_2),.clk(gclk));
	jdff dff_A_QxLJaRx41_0(.dout(w_n681_1[0]),.din(w_dff_A_QxLJaRx41_0),.clk(gclk));
	jdff dff_A_9O4EolNm4_0(.dout(w_dff_A_QxLJaRx41_0),.din(w_dff_A_9O4EolNm4_0),.clk(gclk));
	jdff dff_A_srsVW9Af9_0(.dout(w_dff_A_9O4EolNm4_0),.din(w_dff_A_srsVW9Af9_0),.clk(gclk));
	jdff dff_A_j8tzyT2m1_0(.dout(w_dff_A_srsVW9Af9_0),.din(w_dff_A_j8tzyT2m1_0),.clk(gclk));
	jdff dff_A_jHm2wTS61_1(.dout(w_n681_1[1]),.din(w_dff_A_jHm2wTS61_1),.clk(gclk));
	jdff dff_A_zKmaTsBv8_1(.dout(w_n1568_0[1]),.din(w_dff_A_zKmaTsBv8_1),.clk(gclk));
	jdff dff_B_fiDJVqRi0_1(.din(n1562),.dout(w_dff_B_fiDJVqRi0_1),.clk(gclk));
	jdff dff_B_9mibG71Y7_0(.din(n1563),.dout(w_dff_B_9mibG71Y7_0),.clk(gclk));
	jdff dff_B_IJNya5Rl8_1(.din(n1557),.dout(w_dff_B_IJNya5Rl8_1),.clk(gclk));
	jdff dff_A_ikduT0UA6_0(.dout(w_n1555_0[0]),.din(w_dff_A_ikduT0UA6_0),.clk(gclk));
	jdff dff_A_i0edykUa5_0(.dout(w_dff_A_ikduT0UA6_0),.din(w_dff_A_i0edykUa5_0),.clk(gclk));
	jdff dff_B_LOnslHMK5_2(.din(n1553),.dout(w_dff_B_LOnslHMK5_2),.clk(gclk));
	jdff dff_B_KrP6ACxw1_2(.din(w_dff_B_LOnslHMK5_2),.dout(w_dff_B_KrP6ACxw1_2),.clk(gclk));
	jdff dff_B_tMwK3bNH7_2(.din(w_dff_B_KrP6ACxw1_2),.dout(w_dff_B_tMwK3bNH7_2),.clk(gclk));
	jdff dff_B_JjpdH9y39_2(.din(w_dff_B_tMwK3bNH7_2),.dout(w_dff_B_JjpdH9y39_2),.clk(gclk));
	jdff dff_B_bsSRZaF56_2(.din(w_dff_B_JjpdH9y39_2),.dout(w_dff_B_bsSRZaF56_2),.clk(gclk));
	jdff dff_B_bK8R2NEB5_2(.din(w_dff_B_bsSRZaF56_2),.dout(w_dff_B_bK8R2NEB5_2),.clk(gclk));
	jdff dff_B_3kGxsvzi2_0(.din(n1551),.dout(w_dff_B_3kGxsvzi2_0),.clk(gclk));
	jdff dff_B_IknBggBW4_0(.din(w_dff_B_3kGxsvzi2_0),.dout(w_dff_B_IknBggBW4_0),.clk(gclk));
	jdff dff_B_wrBjtwS76_0(.din(w_dff_B_IknBggBW4_0),.dout(w_dff_B_wrBjtwS76_0),.clk(gclk));
	jdff dff_B_CCqndtHG8_0(.din(n1550),.dout(w_dff_B_CCqndtHG8_0),.clk(gclk));
	jdff dff_B_7ohlDYPp9_0(.din(w_dff_B_CCqndtHG8_0),.dout(w_dff_B_7ohlDYPp9_0),.clk(gclk));
	jdff dff_B_e0AiH9RI4_0(.din(w_dff_B_7ohlDYPp9_0),.dout(w_dff_B_e0AiH9RI4_0),.clk(gclk));
	jdff dff_B_SCPpuGLX7_0(.din(w_dff_B_e0AiH9RI4_0),.dout(w_dff_B_SCPpuGLX7_0),.clk(gclk));
	jdff dff_B_3TEKFXjF7_0(.din(w_dff_B_SCPpuGLX7_0),.dout(w_dff_B_3TEKFXjF7_0),.clk(gclk));
	jdff dff_A_BSIOabYs3_2(.dout(w_n605_1[2]),.din(w_dff_A_BSIOabYs3_2),.clk(gclk));
	jdff dff_A_y1EzK1zt2_2(.dout(w_dff_A_BSIOabYs3_2),.din(w_dff_A_y1EzK1zt2_2),.clk(gclk));
	jdff dff_A_wJ97G8MC0_2(.dout(w_dff_A_y1EzK1zt2_2),.din(w_dff_A_wJ97G8MC0_2),.clk(gclk));
	jdff dff_A_aKdImrnP2_2(.dout(w_dff_A_wJ97G8MC0_2),.din(w_dff_A_aKdImrnP2_2),.clk(gclk));
	jdff dff_A_SsmDP4dU2_2(.dout(w_dff_A_aKdImrnP2_2),.din(w_dff_A_SsmDP4dU2_2),.clk(gclk));
	jdff dff_A_l3KMi0Lf5_2(.dout(w_dff_A_SsmDP4dU2_2),.din(w_dff_A_l3KMi0Lf5_2),.clk(gclk));
	jdff dff_A_YPhObIO37_2(.dout(w_dff_A_l3KMi0Lf5_2),.din(w_dff_A_YPhObIO37_2),.clk(gclk));
	jdff dff_A_jWiQ0e9t3_2(.dout(w_dff_A_YPhObIO37_2),.din(w_dff_A_jWiQ0e9t3_2),.clk(gclk));
	jdff dff_A_YYDdGiXM6_2(.dout(w_dff_A_jWiQ0e9t3_2),.din(w_dff_A_YYDdGiXM6_2),.clk(gclk));
	jdff dff_A_aTQiV29g7_2(.dout(w_dff_A_YYDdGiXM6_2),.din(w_dff_A_aTQiV29g7_2),.clk(gclk));
	jdff dff_A_jLfgwm3B2_2(.dout(w_dff_A_aTQiV29g7_2),.din(w_dff_A_jLfgwm3B2_2),.clk(gclk));
	jdff dff_A_vtSVt5Ke4_2(.dout(w_dff_A_jLfgwm3B2_2),.din(w_dff_A_vtSVt5Ke4_2),.clk(gclk));
	jdff dff_A_oxQIZz4S9_1(.dout(w_n944_0[1]),.din(w_dff_A_oxQIZz4S9_1),.clk(gclk));
	jdff dff_A_GKLhhMUB8_1(.dout(w_dff_A_oxQIZz4S9_1),.din(w_dff_A_GKLhhMUB8_1),.clk(gclk));
	jdff dff_A_rrWg23Ee9_1(.dout(w_dff_A_GKLhhMUB8_1),.din(w_dff_A_rrWg23Ee9_1),.clk(gclk));
	jdff dff_A_ogIfQWlc6_1(.dout(w_dff_A_rrWg23Ee9_1),.din(w_dff_A_ogIfQWlc6_1),.clk(gclk));
	jdff dff_A_1syFJ1BI3_1(.dout(w_dff_A_ogIfQWlc6_1),.din(w_dff_A_1syFJ1BI3_1),.clk(gclk));
	jdff dff_A_wopdOaqf6_1(.dout(w_dff_A_1syFJ1BI3_1),.din(w_dff_A_wopdOaqf6_1),.clk(gclk));
	jdff dff_A_Zw8N9znH7_1(.dout(w_dff_A_wopdOaqf6_1),.din(w_dff_A_Zw8N9znH7_1),.clk(gclk));
	jdff dff_A_vvnwE0dB6_1(.dout(w_dff_A_Zw8N9znH7_1),.din(w_dff_A_vvnwE0dB6_1),.clk(gclk));
	jdff dff_A_JiOFjd856_1(.dout(w_dff_A_vvnwE0dB6_1),.din(w_dff_A_JiOFjd856_1),.clk(gclk));
	jdff dff_A_YA3kvibd3_2(.dout(w_n930_0[2]),.din(w_dff_A_YA3kvibd3_2),.clk(gclk));
	jdff dff_A_lcrB65fP0_2(.dout(w_dff_A_YA3kvibd3_2),.din(w_dff_A_lcrB65fP0_2),.clk(gclk));
	jdff dff_A_Dnw3qxl19_2(.dout(w_dff_A_lcrB65fP0_2),.din(w_dff_A_Dnw3qxl19_2),.clk(gclk));
	jdff dff_A_HhCA1haI8_2(.dout(w_dff_A_Dnw3qxl19_2),.din(w_dff_A_HhCA1haI8_2),.clk(gclk));
	jdff dff_A_myzx6miw8_2(.dout(w_dff_A_HhCA1haI8_2),.din(w_dff_A_myzx6miw8_2),.clk(gclk));
	jdff dff_A_SuTsqUUz7_2(.dout(w_dff_A_myzx6miw8_2),.din(w_dff_A_SuTsqUUz7_2),.clk(gclk));
	jdff dff_A_lTS9xalW3_2(.dout(w_dff_A_SuTsqUUz7_2),.din(w_dff_A_lTS9xalW3_2),.clk(gclk));
	jdff dff_A_xzbAIfva8_2(.dout(w_dff_A_lTS9xalW3_2),.din(w_dff_A_xzbAIfva8_2),.clk(gclk));
	jdff dff_A_DcNViKZO3_2(.dout(w_dff_A_xzbAIfva8_2),.din(w_dff_A_DcNViKZO3_2),.clk(gclk));
	jdff dff_B_8w9SjXgu8_3(.din(n930),.dout(w_dff_B_8w9SjXgu8_3),.clk(gclk));
	jdff dff_B_cNCEHzcg0_3(.din(w_dff_B_8w9SjXgu8_3),.dout(w_dff_B_cNCEHzcg0_3),.clk(gclk));
	jdff dff_A_QPJrCzQ94_1(.dout(w_n700_0[1]),.din(w_dff_A_QPJrCzQ94_1),.clk(gclk));
	jdff dff_A_uQWcp82E3_1(.dout(w_dff_A_QPJrCzQ94_1),.din(w_dff_A_uQWcp82E3_1),.clk(gclk));
	jdff dff_A_HcWZaaDr7_1(.dout(w_dff_A_uQWcp82E3_1),.din(w_dff_A_HcWZaaDr7_1),.clk(gclk));
	jdff dff_A_RabxUM5u6_0(.dout(w_n706_0[0]),.din(w_dff_A_RabxUM5u6_0),.clk(gclk));
	jdff dff_B_LWfr27by0_1(.din(n701),.dout(w_dff_B_LWfr27by0_1),.clk(gclk));
	jdff dff_B_zHdUCnVa4_1(.din(w_dff_B_LWfr27by0_1),.dout(w_dff_B_zHdUCnVa4_1),.clk(gclk));
	jdff dff_B_0rl6XDgm3_0(.din(n599),.dout(w_dff_B_0rl6XDgm3_0),.clk(gclk));
	jdff dff_B_PV5733b09_1(.din(G233),.dout(w_dff_B_PV5733b09_1),.clk(gclk));
	jdff dff_B_yJUIuqCl3_2(.din(n702),.dout(w_dff_B_yJUIuqCl3_2),.clk(gclk));
	jdff dff_A_d2qPCzLc6_0(.dout(w_n604_0[0]),.din(w_dff_A_d2qPCzLc6_0),.clk(gclk));
	jdff dff_B_IrYITDwn2_0(.din(n603),.dout(w_dff_B_IrYITDwn2_0),.clk(gclk));
	jdff dff_B_I4f65N7O1_1(.din(G225),.dout(w_dff_B_I4f65N7O1_1),.clk(gclk));
	jdff dff_A_BSGd3JMX3_1(.dout(w_n928_0[1]),.din(w_dff_A_BSGd3JMX3_1),.clk(gclk));
	jdff dff_A_3ESHHXks4_1(.dout(w_dff_A_BSGd3JMX3_1),.din(w_dff_A_3ESHHXks4_1),.clk(gclk));
	jdff dff_A_cwv6t5gy6_1(.dout(w_dff_A_3ESHHXks4_1),.din(w_dff_A_cwv6t5gy6_1),.clk(gclk));
	jdff dff_A_m14ZmyXb3_1(.dout(w_dff_A_cwv6t5gy6_1),.din(w_dff_A_m14ZmyXb3_1),.clk(gclk));
	jdff dff_A_SkQ9pSQd8_1(.dout(w_dff_A_m14ZmyXb3_1),.din(w_dff_A_SkQ9pSQd8_1),.clk(gclk));
	jdff dff_A_jEfh31XR7_1(.dout(w_dff_A_SkQ9pSQd8_1),.din(w_dff_A_jEfh31XR7_1),.clk(gclk));
	jdff dff_A_mLPZdrPX1_1(.dout(w_dff_A_jEfh31XR7_1),.din(w_dff_A_mLPZdrPX1_1),.clk(gclk));
	jdff dff_A_ifObSwrm4_1(.dout(w_dff_A_mLPZdrPX1_1),.din(w_dff_A_ifObSwrm4_1),.clk(gclk));
	jdff dff_A_pCOCpnTh6_1(.dout(w_dff_A_ifObSwrm4_1),.din(w_dff_A_pCOCpnTh6_1),.clk(gclk));
	jdff dff_B_jqKCjf4A8_2(.din(n928),.dout(w_dff_B_jqKCjf4A8_2),.clk(gclk));
	jdff dff_B_JLAvMhPP4_2(.din(w_dff_B_jqKCjf4A8_2),.dout(w_dff_B_JLAvMhPP4_2),.clk(gclk));
	jdff dff_B_tHW24P2b1_2(.din(w_dff_B_JLAvMhPP4_2),.dout(w_dff_B_tHW24P2b1_2),.clk(gclk));
	jdff dff_A_0flIumw26_0(.dout(w_n596_0[0]),.din(w_dff_A_0flIumw26_0),.clk(gclk));
	jdff dff_A_NFa9gf9t3_0(.dout(w_dff_A_0flIumw26_0),.din(w_dff_A_NFa9gf9t3_0),.clk(gclk));
	jdff dff_A_PfRuB1eH7_0(.dout(w_dff_A_NFa9gf9t3_0),.din(w_dff_A_PfRuB1eH7_0),.clk(gclk));
	jdff dff_A_S5K49NIm7_0(.dout(w_dff_A_PfRuB1eH7_0),.din(w_dff_A_S5K49NIm7_0),.clk(gclk));
	jdff dff_A_09eiEXdN9_0(.dout(w_dff_A_S5K49NIm7_0),.din(w_dff_A_09eiEXdN9_0),.clk(gclk));
	jdff dff_B_p3feOSO34_1(.din(n592),.dout(w_dff_B_p3feOSO34_1),.clk(gclk));
	jdff dff_B_WCFRpAvJ0_1(.din(G209),.dout(w_dff_B_WCFRpAvJ0_1),.clk(gclk));
	jdff dff_B_6kfQng679_0(.din(n1544),.dout(w_dff_B_6kfQng679_0),.clk(gclk));
	jdff dff_A_ZUHGbJNA8_0(.dout(w_n585_0[0]),.din(w_dff_A_ZUHGbJNA8_0),.clk(gclk));
	jdff dff_B_CbaEUmP63_0(.din(n584),.dout(w_dff_B_CbaEUmP63_0),.clk(gclk));
	jdff dff_B_SDAncjIu4_0(.din(w_dff_B_CbaEUmP63_0),.dout(w_dff_B_SDAncjIu4_0),.clk(gclk));
	jdff dff_A_7dpqGCjC5_0(.dout(w_n583_1[0]),.din(w_dff_A_7dpqGCjC5_0),.clk(gclk));
	jdff dff_A_x5NtLHI71_0(.dout(w_dff_A_7dpqGCjC5_0),.din(w_dff_A_x5NtLHI71_0),.clk(gclk));
	jdff dff_A_bnNVtO9w5_0(.dout(w_dff_A_x5NtLHI71_0),.din(w_dff_A_bnNVtO9w5_0),.clk(gclk));
	jdff dff_A_63KvYAOB7_0(.dout(w_n572_0[0]),.din(w_dff_A_63KvYAOB7_0),.clk(gclk));
	jdff dff_A_BPpn6oSc2_0(.dout(w_dff_A_63KvYAOB7_0),.din(w_dff_A_BPpn6oSc2_0),.clk(gclk));
	jdff dff_A_JRHCN90s7_0(.dout(w_dff_A_BPpn6oSc2_0),.din(w_dff_A_JRHCN90s7_0),.clk(gclk));
	jdff dff_A_EXbfzPrL4_0(.dout(w_dff_A_JRHCN90s7_0),.din(w_dff_A_EXbfzPrL4_0),.clk(gclk));
	jdff dff_A_P8xOK5uz1_1(.dout(w_n567_1[1]),.din(w_dff_A_P8xOK5uz1_1),.clk(gclk));
	jdff dff_A_uK6OIkPM0_1(.dout(w_n567_0[1]),.din(w_dff_A_uK6OIkPM0_1),.clk(gclk));
	jdff dff_A_wIlEuhuF7_1(.dout(w_dff_A_uK6OIkPM0_1),.din(w_dff_A_wIlEuhuF7_1),.clk(gclk));
	jdff dff_A_9WJodyuM8_1(.dout(w_dff_A_wIlEuhuF7_1),.din(w_dff_A_9WJodyuM8_1),.clk(gclk));
	jdff dff_A_IwN1l2Xb1_0(.dout(w_n497_1[0]),.din(w_dff_A_IwN1l2Xb1_0),.clk(gclk));
	jdff dff_A_fMctWRTU0_0(.dout(w_n562_0[0]),.din(w_dff_A_fMctWRTU0_0),.clk(gclk));
	jdff dff_A_92dWOa9m5_0(.dout(w_dff_A_fMctWRTU0_0),.din(w_dff_A_92dWOa9m5_0),.clk(gclk));
	jdff dff_A_zTGz7cTw7_0(.dout(w_dff_A_92dWOa9m5_0),.din(w_dff_A_zTGz7cTw7_0),.clk(gclk));
	jdff dff_A_mMMU0x3m6_0(.dout(w_dff_A_zTGz7cTw7_0),.din(w_dff_A_mMMU0x3m6_0),.clk(gclk));
	jdff dff_A_YLbN2nBA3_0(.dout(w_dff_A_mMMU0x3m6_0),.din(w_dff_A_YLbN2nBA3_0),.clk(gclk));
	jdff dff_B_Q17ELFLL2_2(.din(n562),.dout(w_dff_B_Q17ELFLL2_2),.clk(gclk));
	jdff dff_B_f1SPZpZX8_2(.din(w_dff_B_Q17ELFLL2_2),.dout(w_dff_B_f1SPZpZX8_2),.clk(gclk));
	jdff dff_A_LT7SfRtI1_0(.dout(w_n561_0[0]),.din(w_dff_A_LT7SfRtI1_0),.clk(gclk));
	jdff dff_A_QeGAPcQN6_1(.dout(w_n561_0[1]),.din(w_dff_A_QeGAPcQN6_1),.clk(gclk));
	jdff dff_A_TYKPX5VY6_1(.dout(w_dff_A_QeGAPcQN6_1),.din(w_dff_A_TYKPX5VY6_1),.clk(gclk));
	jdff dff_A_Q094VyXA8_1(.dout(w_dff_A_TYKPX5VY6_1),.din(w_dff_A_Q094VyXA8_1),.clk(gclk));
	jdff dff_A_ZrUszQjG6_0(.dout(w_G1497_0[0]),.din(w_dff_A_ZrUszQjG6_0),.clk(gclk));
	jdff dff_A_5X3yEdkl6_0(.dout(w_dff_A_ZrUszQjG6_0),.din(w_dff_A_5X3yEdkl6_0),.clk(gclk));
	jdff dff_A_GrRXcfIM7_0(.dout(w_dff_A_5X3yEdkl6_0),.din(w_dff_A_GrRXcfIM7_0),.clk(gclk));
	jdff dff_A_Bb9lsqzh5_0(.dout(w_dff_A_GrRXcfIM7_0),.din(w_dff_A_Bb9lsqzh5_0),.clk(gclk));
	jdff dff_A_kEMwIXIn5_0(.dout(w_dff_A_Bb9lsqzh5_0),.din(w_dff_A_kEMwIXIn5_0),.clk(gclk));
	jdff dff_A_0Fa8os3z7_0(.dout(w_dff_A_kEMwIXIn5_0),.din(w_dff_A_0Fa8os3z7_0),.clk(gclk));
	jdff dff_A_FS4Kxid42_0(.dout(w_dff_A_0Fa8os3z7_0),.din(w_dff_A_FS4Kxid42_0),.clk(gclk));
	jdff dff_A_oWUaqytK7_0(.dout(w_dff_A_FS4Kxid42_0),.din(w_dff_A_oWUaqytK7_0),.clk(gclk));
	jdff dff_A_dG2Mjsc11_0(.dout(w_dff_A_oWUaqytK7_0),.din(w_dff_A_dG2Mjsc11_0),.clk(gclk));
	jdff dff_A_eSrgxN3W7_0(.dout(w_dff_A_dG2Mjsc11_0),.din(w_dff_A_eSrgxN3W7_0),.clk(gclk));
	jdff dff_A_OYUQNdxS0_0(.dout(w_dff_A_eSrgxN3W7_0),.din(w_dff_A_OYUQNdxS0_0),.clk(gclk));
	jdff dff_A_JqaM0uqn6_0(.dout(w_dff_A_OYUQNdxS0_0),.din(w_dff_A_JqaM0uqn6_0),.clk(gclk));
	jdff dff_A_JIsGZ0Ow2_2(.dout(w_G1497_0[2]),.din(w_dff_A_JIsGZ0Ow2_2),.clk(gclk));
	jdff dff_A_UsYkc8JY3_2(.dout(w_dff_A_JIsGZ0Ow2_2),.din(w_dff_A_UsYkc8JY3_2),.clk(gclk));
	jdff dff_A_bFLN5keE7_2(.dout(w_dff_A_UsYkc8JY3_2),.din(w_dff_A_bFLN5keE7_2),.clk(gclk));
	jdff dff_A_2PVSg64j2_2(.dout(w_dff_A_bFLN5keE7_2),.din(w_dff_A_2PVSg64j2_2),.clk(gclk));
	jdff dff_A_kdVLLeTI5_2(.dout(w_dff_A_2PVSg64j2_2),.din(w_dff_A_kdVLLeTI5_2),.clk(gclk));
	jdff dff_A_t9pvmhFv2_2(.dout(w_dff_A_kdVLLeTI5_2),.din(w_dff_A_t9pvmhFv2_2),.clk(gclk));
	jdff dff_A_PU2cSZfk8_2(.dout(w_dff_A_t9pvmhFv2_2),.din(w_dff_A_PU2cSZfk8_2),.clk(gclk));
	jdff dff_A_pMmppbiq0_2(.dout(w_dff_A_PU2cSZfk8_2),.din(w_dff_A_pMmppbiq0_2),.clk(gclk));
	jdff dff_A_er9MN6VG4_2(.dout(w_dff_A_pMmppbiq0_2),.din(w_dff_A_er9MN6VG4_2),.clk(gclk));
	jdff dff_A_EWHZ9Osq4_2(.dout(w_dff_A_er9MN6VG4_2),.din(w_dff_A_EWHZ9Osq4_2),.clk(gclk));
	jdff dff_B_oq0Ywofd2_1(.din(n675),.dout(w_dff_B_oq0Ywofd2_1),.clk(gclk));
	jdff dff_B_gZDI64Ns3_1(.din(w_dff_B_oq0Ywofd2_1),.dout(w_dff_B_gZDI64Ns3_1),.clk(gclk));
	jdff dff_B_7T1LkwOg9_1(.din(w_dff_B_gZDI64Ns3_1),.dout(w_dff_B_7T1LkwOg9_1),.clk(gclk));
	jdff dff_B_ahsHh9Ol7_1(.din(w_dff_B_7T1LkwOg9_1),.dout(w_dff_B_ahsHh9Ol7_1),.clk(gclk));
	jdff dff_B_CbbG04359_1(.din(n676),.dout(w_dff_B_CbbG04359_1),.clk(gclk));
	jdff dff_B_bOYmoYFs5_1(.din(w_dff_B_CbbG04359_1),.dout(w_dff_B_bOYmoYFs5_1),.clk(gclk));
	jdff dff_B_Xz7zCVNm5_1(.din(w_dff_B_bOYmoYFs5_1),.dout(w_dff_B_Xz7zCVNm5_1),.clk(gclk));
	jdff dff_B_9hso8GXL7_1(.din(w_dff_B_Xz7zCVNm5_1),.dout(w_dff_B_9hso8GXL7_1),.clk(gclk));
	jdff dff_B_1PaqHFXG2_1(.din(w_dff_B_9hso8GXL7_1),.dout(w_dff_B_1PaqHFXG2_1),.clk(gclk));
	jdff dff_A_8v12xvBk6_1(.dout(w_n691_0[1]),.din(w_dff_A_8v12xvBk6_1),.clk(gclk));
	jdff dff_A_JOLCGD738_0(.dout(w_n689_0[0]),.din(w_dff_A_JOLCGD738_0),.clk(gclk));
	jdff dff_A_NiKCeGge1_0(.dout(w_n687_0[0]),.din(w_dff_A_NiKCeGge1_0),.clk(gclk));
	jdff dff_A_hVs7x4Xo4_1(.dout(w_n687_0[1]),.din(w_dff_A_hVs7x4Xo4_1),.clk(gclk));
	jdff dff_A_qTLdxIJi4_1(.dout(w_dff_A_hVs7x4Xo4_1),.din(w_dff_A_qTLdxIJi4_1),.clk(gclk));
	jdff dff_A_ssmlvYDc9_1(.dout(w_dff_A_qTLdxIJi4_1),.din(w_dff_A_ssmlvYDc9_1),.clk(gclk));
	jdff dff_A_EvD6p0zS9_1(.dout(w_dff_A_ssmlvYDc9_1),.din(w_dff_A_EvD6p0zS9_1),.clk(gclk));
	jdff dff_A_VD5hiWkc2_2(.dout(w_n571_0[2]),.din(w_dff_A_VD5hiWkc2_2),.clk(gclk));
	jdff dff_A_4yccVk0V6_2(.dout(w_dff_A_VD5hiWkc2_2),.din(w_dff_A_4yccVk0V6_2),.clk(gclk));
	jdff dff_A_9prX5OOG0_2(.dout(w_dff_A_4yccVk0V6_2),.din(w_dff_A_9prX5OOG0_2),.clk(gclk));
	jdff dff_A_SU22FOku6_1(.dout(w_n569_0[1]),.din(w_dff_A_SU22FOku6_1),.clk(gclk));
	jdff dff_A_dIXvuexv7_1(.dout(w_G280_0[1]),.din(w_dff_A_dIXvuexv7_1),.clk(gclk));
	jdff dff_A_iqc2tmVP1_0(.dout(w_n486_1[0]),.din(w_dff_A_iqc2tmVP1_0),.clk(gclk));
	jdff dff_A_pe5x4dCf1_0(.dout(w_n681_2[0]),.din(w_dff_A_pe5x4dCf1_0),.clk(gclk));
	jdff dff_A_CZu92rYw1_0(.dout(w_dff_A_pe5x4dCf1_0),.din(w_dff_A_CZu92rYw1_0),.clk(gclk));
	jdff dff_A_Vpom8c187_1(.dout(w_n680_0[1]),.din(w_dff_A_Vpom8c187_1),.clk(gclk));
	jdff dff_B_97Od1iLj9_2(.din(n680),.dout(w_dff_B_97Od1iLj9_2),.clk(gclk));
	jdff dff_A_rdwYEB797_0(.dout(w_n451_1[0]),.din(w_dff_A_rdwYEB797_0),.clk(gclk));
	jdff dff_A_BUnEjW585_1(.dout(w_n679_0[1]),.din(w_dff_A_BUnEjW585_1),.clk(gclk));
	jdff dff_A_EeOODEu20_1(.dout(w_dff_A_BUnEjW585_1),.din(w_dff_A_EeOODEu20_1),.clk(gclk));
	jdff dff_A_LoROC9dG1_1(.dout(w_n678_0[1]),.din(w_dff_A_LoROC9dG1_1),.clk(gclk));
	jdff dff_A_6jdQc28D4_1(.dout(w_dff_A_LoROC9dG1_1),.din(w_dff_A_6jdQc28D4_1),.clk(gclk));
	jdff dff_A_cdBdRrEJ6_1(.dout(w_dff_A_6jdQc28D4_1),.din(w_dff_A_cdBdRrEJ6_1),.clk(gclk));
	jdff dff_B_c5b0SisU2_1(.din(n557),.dout(w_dff_B_c5b0SisU2_1),.clk(gclk));
	jdff dff_B_OdDnxJVz1_1(.din(G241),.dout(w_dff_B_OdDnxJVz1_1),.clk(gclk));
	jdff dff_B_nYHrPa6X7_2(.din(n1543),.dout(w_dff_B_nYHrPa6X7_2),.clk(gclk));
	jdff dff_B_NCF2avyc2_2(.din(w_dff_B_nYHrPa6X7_2),.dout(w_dff_B_NCF2avyc2_2),.clk(gclk));
	jdff dff_B_70esU5vR8_2(.din(w_dff_B_NCF2avyc2_2),.dout(w_dff_B_70esU5vR8_2),.clk(gclk));
	jdff dff_B_8sWR1LZ04_2(.din(w_dff_B_70esU5vR8_2),.dout(w_dff_B_8sWR1LZ04_2),.clk(gclk));
	jdff dff_B_MNvJXFBW1_2(.din(w_dff_B_8sWR1LZ04_2),.dout(w_dff_B_MNvJXFBW1_2),.clk(gclk));
	jdff dff_B_rABvzCqa6_2(.din(w_dff_B_MNvJXFBW1_2),.dout(w_dff_B_rABvzCqa6_2),.clk(gclk));
	jdff dff_B_piFvOyF13_2(.din(w_dff_B_rABvzCqa6_2),.dout(w_dff_B_piFvOyF13_2),.clk(gclk));
	jdff dff_B_FvrOhXZl9_2(.din(w_dff_B_piFvOyF13_2),.dout(w_dff_B_FvrOhXZl9_2),.clk(gclk));
	jdff dff_B_BIDd6ZH78_2(.din(w_dff_B_FvrOhXZl9_2),.dout(w_dff_B_BIDd6ZH78_2),.clk(gclk));
	jdff dff_B_4ofr7wj29_2(.din(w_dff_B_BIDd6ZH78_2),.dout(w_dff_B_4ofr7wj29_2),.clk(gclk));
	jdff dff_A_fAbKqvX35_2(.dout(w_n583_0[2]),.din(w_dff_A_fAbKqvX35_2),.clk(gclk));
	jdff dff_A_OQaTlxtk6_2(.dout(w_dff_A_fAbKqvX35_2),.din(w_dff_A_OQaTlxtk6_2),.clk(gclk));
	jdff dff_A_uMBcqh5w8_2(.dout(w_dff_A_OQaTlxtk6_2),.din(w_dff_A_uMBcqh5w8_2),.clk(gclk));
	jdff dff_A_96EIOfti0_2(.dout(w_dff_A_uMBcqh5w8_2),.din(w_dff_A_96EIOfti0_2),.clk(gclk));
	jdff dff_A_OVx7vuIf6_2(.dout(w_dff_A_96EIOfti0_2),.din(w_dff_A_OVx7vuIf6_2),.clk(gclk));
	jdff dff_A_3W9nTXQe8_1(.dout(w_n578_0[1]),.din(w_dff_A_3W9nTXQe8_1),.clk(gclk));
	jdff dff_A_CZc7oxpZ0_1(.dout(w_dff_A_3W9nTXQe8_1),.din(w_dff_A_CZc7oxpZ0_1),.clk(gclk));
	jdff dff_A_p16N9eAf4_1(.dout(w_dff_A_CZc7oxpZ0_1),.din(w_dff_A_p16N9eAf4_1),.clk(gclk));
	jdff dff_A_IRvJ5n7H9_1(.dout(w_dff_A_p16N9eAf4_1),.din(w_dff_A_IRvJ5n7H9_1),.clk(gclk));
	jdff dff_A_mRHePuIw5_1(.dout(w_dff_A_IRvJ5n7H9_1),.din(w_dff_A_mRHePuIw5_1),.clk(gclk));
	jdff dff_A_ZM6t2rqF7_1(.dout(w_dff_A_mRHePuIw5_1),.din(w_dff_A_ZM6t2rqF7_1),.clk(gclk));
	jdff dff_A_nLtBEqxt1_1(.dout(w_dff_A_ZM6t2rqF7_1),.din(w_dff_A_nLtBEqxt1_1),.clk(gclk));
	jdff dff_B_y2DrAnYB0_0(.din(n576),.dout(w_dff_B_y2DrAnYB0_0),.clk(gclk));
	jdff dff_A_X5VE5Rn87_0(.dout(w_G335_3[0]),.din(w_dff_A_X5VE5Rn87_0),.clk(gclk));
	jdff dff_B_ex8iQiFj3_1(.din(G264),.dout(w_dff_B_ex8iQiFj3_1),.clk(gclk));
	jdff dff_A_I48WH7cW8_0(.dout(w_n473_1[0]),.din(w_dff_A_I48WH7cW8_0),.clk(gclk));
	jdff dff_A_xwueaaXp8_0(.dout(w_dff_A_I48WH7cW8_0),.din(w_dff_A_xwueaaXp8_0),.clk(gclk));
	jdff dff_A_3XYAaoiY3_1(.dout(w_n473_1[1]),.din(w_dff_A_3XYAaoiY3_1),.clk(gclk));
	jdff dff_A_BBMmeLKm0_1(.dout(w_n943_0[1]),.din(w_dff_A_BBMmeLKm0_1),.clk(gclk));
	jdff dff_A_rEbBXL8M5_1(.dout(w_dff_A_BBMmeLKm0_1),.din(w_dff_A_rEbBXL8M5_1),.clk(gclk));
	jdff dff_A_gq866Uyx9_1(.dout(w_dff_A_rEbBXL8M5_1),.din(w_dff_A_gq866Uyx9_1),.clk(gclk));
	jdff dff_A_iFiqIPSR9_1(.dout(w_dff_A_gq866Uyx9_1),.din(w_dff_A_iFiqIPSR9_1),.clk(gclk));
	jdff dff_A_pTzrZNO72_1(.dout(w_dff_A_iFiqIPSR9_1),.din(w_dff_A_pTzrZNO72_1),.clk(gclk));
	jdff dff_A_habZwT1r8_1(.dout(w_dff_A_pTzrZNO72_1),.din(w_dff_A_habZwT1r8_1),.clk(gclk));
	jdff dff_A_hLTnTAOU5_1(.dout(w_dff_A_habZwT1r8_1),.din(w_dff_A_hLTnTAOU5_1),.clk(gclk));
	jdff dff_A_huzUM75a1_1(.dout(w_dff_A_hLTnTAOU5_1),.din(w_dff_A_huzUM75a1_1),.clk(gclk));
	jdff dff_A_wi0ZbLkl6_1(.dout(w_dff_A_huzUM75a1_1),.din(w_dff_A_wi0ZbLkl6_1),.clk(gclk));
	jdff dff_A_n8KaUCZM2_1(.dout(w_dff_A_wi0ZbLkl6_1),.din(w_dff_A_n8KaUCZM2_1),.clk(gclk));
	jdff dff_A_3kVqWks17_1(.dout(w_dff_A_n8KaUCZM2_1),.din(w_dff_A_3kVqWks17_1),.clk(gclk));
	jdff dff_A_rc6cyPT01_1(.dout(w_dff_A_3kVqWks17_1),.din(w_dff_A_rc6cyPT01_1),.clk(gclk));
	jdff dff_A_nJ2td3iY0_1(.dout(w_n591_0[1]),.din(w_dff_A_nJ2td3iY0_1),.clk(gclk));
	jdff dff_A_Gt3ZoqjV6_1(.dout(w_n590_0[1]),.din(w_dff_A_Gt3ZoqjV6_1),.clk(gclk));
	jdff dff_A_K7sE6wq35_1(.dout(w_dff_A_Gt3ZoqjV6_1),.din(w_dff_A_K7sE6wq35_1),.clk(gclk));
	jdff dff_B_7O06H6yB2_0(.din(n589),.dout(w_dff_B_7O06H6yB2_0),.clk(gclk));
	jdff dff_B_oSc3NJlp1_1(.din(G217),.dout(w_dff_B_oSc3NJlp1_1),.clk(gclk));
	jdff dff_A_Y0C5iHwL0_0(.dout(w_G335_4[0]),.din(w_dff_A_Y0C5iHwL0_0),.clk(gclk));
	jdff dff_A_6CHDTV882_2(.dout(w_G335_1[2]),.din(w_dff_A_6CHDTV882_2),.clk(gclk));
	jdff dff_A_SJM3llbf3_1(.dout(w_n750_0[1]),.din(w_dff_A_SJM3llbf3_1),.clk(gclk));
	jdff dff_A_u8JSnDQi1_1(.dout(w_dff_A_SJM3llbf3_1),.din(w_dff_A_u8JSnDQi1_1),.clk(gclk));
	jdff dff_A_il7T7hol3_1(.dout(w_dff_A_u8JSnDQi1_1),.din(w_dff_A_il7T7hol3_1),.clk(gclk));
	jdff dff_A_IV7T04QO9_1(.dout(w_dff_A_il7T7hol3_1),.din(w_dff_A_IV7T04QO9_1),.clk(gclk));
	jdff dff_A_NgP28wni9_1(.dout(w_dff_A_IV7T04QO9_1),.din(w_dff_A_NgP28wni9_1),.clk(gclk));
	jdff dff_A_cuQLzaUW8_1(.dout(w_dff_A_NgP28wni9_1),.din(w_dff_A_cuQLzaUW8_1),.clk(gclk));
	jdff dff_A_bmyElyw24_1(.dout(w_dff_A_cuQLzaUW8_1),.din(w_dff_A_bmyElyw24_1),.clk(gclk));
	jdff dff_A_2ljb2NLh7_1(.dout(w_dff_A_bmyElyw24_1),.din(w_dff_A_2ljb2NLh7_1),.clk(gclk));
	jdff dff_A_1pPdm0Gj8_1(.dout(w_dff_A_2ljb2NLh7_1),.din(w_dff_A_1pPdm0Gj8_1),.clk(gclk));
	jdff dff_A_830R7nnO7_1(.dout(w_dff_A_1pPdm0Gj8_1),.din(w_dff_A_830R7nnO7_1),.clk(gclk));
	jdff dff_A_HWW4jZFn9_1(.dout(w_dff_A_830R7nnO7_1),.din(w_dff_A_HWW4jZFn9_1),.clk(gclk));
	jdff dff_A_nFQtPAcr9_1(.dout(w_dff_A_HWW4jZFn9_1),.din(w_dff_A_nFQtPAcr9_1),.clk(gclk));
	jdff dff_A_8s4z32cf7_1(.dout(w_dff_A_nFQtPAcr9_1),.din(w_dff_A_8s4z32cf7_1),.clk(gclk));
	jdff dff_A_zfGaarHY9_1(.dout(w_dff_A_8s4z32cf7_1),.din(w_dff_A_zfGaarHY9_1),.clk(gclk));
	jdff dff_A_EdWZtHnH2_1(.dout(w_dff_A_zfGaarHY9_1),.din(w_dff_A_EdWZtHnH2_1),.clk(gclk));
	jdff dff_A_zQQQTv6k9_1(.dout(w_dff_A_EdWZtHnH2_1),.din(w_dff_A_zQQQTv6k9_1),.clk(gclk));
	jdff dff_A_vGWoQ90w7_1(.dout(w_dff_A_zQQQTv6k9_1),.din(w_dff_A_vGWoQ90w7_1),.clk(gclk));
	jdff dff_A_HAUkrzKr3_2(.dout(w_n750_0[2]),.din(w_dff_A_HAUkrzKr3_2),.clk(gclk));
	jdff dff_A_U6v1aeNf5_2(.dout(w_dff_A_HAUkrzKr3_2),.din(w_dff_A_U6v1aeNf5_2),.clk(gclk));
	jdff dff_A_G3jFXJA17_2(.dout(w_dff_A_U6v1aeNf5_2),.din(w_dff_A_G3jFXJA17_2),.clk(gclk));
	jdff dff_A_n6Sv8eHr5_2(.dout(w_dff_A_G3jFXJA17_2),.din(w_dff_A_n6Sv8eHr5_2),.clk(gclk));
	jdff dff_A_uuHG5Q250_2(.dout(w_dff_A_n6Sv8eHr5_2),.din(w_dff_A_uuHG5Q250_2),.clk(gclk));
	jdff dff_A_Ru9HNxHt3_2(.dout(w_dff_A_uuHG5Q250_2),.din(w_dff_A_Ru9HNxHt3_2),.clk(gclk));
	jdff dff_A_uAOJH08I9_2(.dout(w_dff_A_Ru9HNxHt3_2),.din(w_dff_A_uAOJH08I9_2),.clk(gclk));
	jdff dff_A_NYquPSHS8_2(.dout(w_dff_A_uAOJH08I9_2),.din(w_dff_A_NYquPSHS8_2),.clk(gclk));
	jdff dff_A_5GaXf1406_2(.dout(w_G4091_2[2]),.din(w_dff_A_5GaXf1406_2),.clk(gclk));
	jdff dff_A_pMnAPbPy2_2(.dout(w_G4091_0[2]),.din(w_dff_A_pMnAPbPy2_2),.clk(gclk));
	jdff dff_A_fUn5nLBT4_2(.dout(w_dff_A_pMnAPbPy2_2),.din(w_dff_A_fUn5nLBT4_2),.clk(gclk));
	jdff dff_A_s5nuRzJv2_2(.dout(w_dff_A_fUn5nLBT4_2),.din(w_dff_A_s5nuRzJv2_2),.clk(gclk));
	jdff dff_A_VThthqik6_2(.dout(w_dff_A_s5nuRzJv2_2),.din(w_dff_A_VThthqik6_2),.clk(gclk));
	jdff dff_A_zxu4Y6xJ2_2(.dout(w_dff_A_VThthqik6_2),.din(w_dff_A_zxu4Y6xJ2_2),.clk(gclk));
	jdff dff_A_2vUuaBgp4_2(.dout(w_dff_A_zxu4Y6xJ2_2),.din(w_dff_A_2vUuaBgp4_2),.clk(gclk));
	jdff dff_A_wnUidp9P8_2(.dout(w_dff_A_2vUuaBgp4_2),.din(w_dff_A_wnUidp9P8_2),.clk(gclk));
	jdff dff_A_GkHTtTX37_2(.dout(w_dff_A_wnUidp9P8_2),.din(w_dff_A_GkHTtTX37_2),.clk(gclk));
	jdff dff_A_9KWaRm4D7_2(.dout(w_dff_A_GkHTtTX37_2),.din(w_dff_A_9KWaRm4D7_2),.clk(gclk));
	jdff dff_A_gV6NFZlV5_2(.dout(w_dff_A_9KWaRm4D7_2),.din(w_dff_A_gV6NFZlV5_2),.clk(gclk));
	jdff dff_A_vaajNmmr9_2(.dout(w_dff_A_gV6NFZlV5_2),.din(w_dff_A_vaajNmmr9_2),.clk(gclk));
	jdff dff_A_xCnhGROG9_2(.dout(w_dff_A_vaajNmmr9_2),.din(w_dff_A_xCnhGROG9_2),.clk(gclk));
	jdff dff_A_ydaMKyjA1_2(.dout(w_dff_A_xCnhGROG9_2),.din(w_dff_A_ydaMKyjA1_2),.clk(gclk));
	jdff dff_A_COWnrVOF2_2(.dout(w_dff_A_ydaMKyjA1_2),.din(w_dff_A_COWnrVOF2_2),.clk(gclk));
	jdff dff_A_0n8QOOed6_2(.dout(w_dff_A_COWnrVOF2_2),.din(w_dff_A_0n8QOOed6_2),.clk(gclk));
	jdff dff_A_QMHeXJpH0_2(.dout(w_dff_A_0n8QOOed6_2),.din(w_dff_A_QMHeXJpH0_2),.clk(gclk));
	jdff dff_A_2K3aXCom4_2(.dout(w_dff_A_QMHeXJpH0_2),.din(w_dff_A_2K3aXCom4_2),.clk(gclk));
	jdff dff_A_mDT9zZ7v2_2(.dout(w_dff_A_2K3aXCom4_2),.din(w_dff_A_mDT9zZ7v2_2),.clk(gclk));
	jdff dff_B_otbjf07u4_2(.din(n1533),.dout(w_dff_B_otbjf07u4_2),.clk(gclk));
	jdff dff_B_m1R52wP16_1(.din(n1526),.dout(w_dff_B_m1R52wP16_1),.clk(gclk));
	jdff dff_B_AJTqV7fd2_1(.din(n1527),.dout(w_dff_B_AJTqV7fd2_1),.clk(gclk));
	jdff dff_A_1YbHecmV2_0(.dout(w_n486_0[0]),.din(w_dff_A_1YbHecmV2_0),.clk(gclk));
	jdff dff_A_posRy3dw0_2(.dout(w_n486_0[2]),.din(w_dff_A_posRy3dw0_2),.clk(gclk));
	jdff dff_A_8RSXgteW1_2(.dout(w_dff_A_posRy3dw0_2),.din(w_dff_A_8RSXgteW1_2),.clk(gclk));
	jdff dff_A_d064H4t07_0(.dout(w_G411_0[0]),.din(w_dff_A_d064H4t07_0),.clk(gclk));
	jdff dff_A_Zw8gwf5R7_0(.dout(w_dff_A_d064H4t07_0),.din(w_dff_A_Zw8gwf5R7_0),.clk(gclk));
	jdff dff_A_6BR4DVNt6_1(.dout(w_G411_0[1]),.din(w_dff_A_6BR4DVNt6_1),.clk(gclk));
	jdff dff_A_HlJL891t2_1(.dout(w_G273_2[1]),.din(w_dff_A_HlJL891t2_1),.clk(gclk));
	jdff dff_A_rbLJ0fbJ2_2(.dout(w_G273_0[2]),.din(w_dff_A_rbLJ0fbJ2_2),.clk(gclk));
	jdff dff_B_YIiBl1PT1_1(.din(n1518),.dout(w_dff_B_YIiBl1PT1_1),.clk(gclk));
	jdff dff_B_pwRFMlrp9_1(.din(w_dff_B_YIiBl1PT1_1),.dout(w_dff_B_pwRFMlrp9_1),.clk(gclk));
	jdff dff_A_VieoZLRK7_2(.dout(w_n473_0[2]),.din(w_dff_A_VieoZLRK7_2),.clk(gclk));
	jdff dff_A_yQsZz6LY3_2(.dout(w_dff_A_VieoZLRK7_2),.din(w_dff_A_yQsZz6LY3_2),.clk(gclk));
	jdff dff_B_c5M0faWB5_3(.din(n473),.dout(w_dff_B_c5M0faWB5_3),.clk(gclk));
	jdff dff_B_s5CmWdDh1_1(.din(n1514),.dout(w_dff_B_s5CmWdDh1_1),.clk(gclk));
	jdff dff_A_KFQivGam9_1(.dout(w_G257_2[1]),.din(w_dff_A_KFQivGam9_1),.clk(gclk));
	jdff dff_A_PP7ffUZ67_0(.dout(w_G389_0[0]),.din(w_dff_A_PP7ffUZ67_0),.clk(gclk));
	jdff dff_A_ntbxNQMz8_0(.dout(w_dff_A_PP7ffUZ67_0),.din(w_dff_A_ntbxNQMz8_0),.clk(gclk));
	jdff dff_A_G0yvkdsE8_1(.dout(w_G389_0[1]),.din(w_dff_A_G0yvkdsE8_1),.clk(gclk));
	jdff dff_A_0vmrnqG67_0(.dout(w_G257_1[0]),.din(w_dff_A_0vmrnqG67_0),.clk(gclk));
	jdff dff_B_8WJiVgDg4_1(.din(n1507),.dout(w_dff_B_8WJiVgDg4_1),.clk(gclk));
	jdff dff_B_dA7S9O0q4_1(.din(n1508),.dout(w_dff_B_dA7S9O0q4_1),.clk(gclk));
	jdff dff_A_yzVfqSoE5_0(.dout(w_n451_0[0]),.din(w_dff_A_yzVfqSoE5_0),.clk(gclk));
	jdff dff_A_XPcdGorN6_2(.dout(w_n451_0[2]),.din(w_dff_A_XPcdGorN6_2),.clk(gclk));
	jdff dff_A_C9wiUB3i5_2(.dout(w_dff_A_XPcdGorN6_2),.din(w_dff_A_C9wiUB3i5_2),.clk(gclk));
	jdff dff_A_SQiowSOU1_0(.dout(w_G400_1[0]),.din(w_dff_A_SQiowSOU1_0),.clk(gclk));
	jdff dff_A_KwfjedKL4_1(.dout(w_G400_0[1]),.din(w_dff_A_KwfjedKL4_1),.clk(gclk));
	jdff dff_A_LR4UwY9l0_1(.dout(w_dff_A_KwfjedKL4_1),.din(w_dff_A_LR4UwY9l0_1),.clk(gclk));
	jdff dff_A_ttdzmNqI7_2(.dout(w_G400_0[2]),.din(w_dff_A_ttdzmNqI7_2),.clk(gclk));
	jdff dff_A_rSBlSYSC0_2(.dout(w_dff_A_ttdzmNqI7_2),.din(w_dff_A_rSBlSYSC0_2),.clk(gclk));
	jdff dff_A_bodr78eO0_2(.dout(w_dff_A_rSBlSYSC0_2),.din(w_dff_A_bodr78eO0_2),.clk(gclk));
	jdff dff_A_GHf1WuLw3_0(.dout(w_G265_2[0]),.din(w_dff_A_GHf1WuLw3_0),.clk(gclk));
	jdff dff_A_e3JIbNxC8_2(.dout(w_G265_0[2]),.din(w_dff_A_e3JIbNxC8_2),.clk(gclk));
	jdff dff_B_F7dSwWAA2_1(.din(n1498),.dout(w_dff_B_F7dSwWAA2_1),.clk(gclk));
	jdff dff_B_t4xIJt4T5_1(.din(n1499),.dout(w_dff_B_t4xIJt4T5_1),.clk(gclk));
	jdff dff_A_CQDvDQIN0_0(.dout(w_n497_0[0]),.din(w_dff_A_CQDvDQIN0_0),.clk(gclk));
	jdff dff_A_KbGIdVt48_2(.dout(w_n497_0[2]),.din(w_dff_A_KbGIdVt48_2),.clk(gclk));
	jdff dff_A_53wdL9Ic4_2(.dout(w_dff_A_KbGIdVt48_2),.din(w_dff_A_53wdL9Ic4_2),.clk(gclk));
	jdff dff_A_ZMRooXgA5_0(.dout(w_G374_0[0]),.din(w_dff_A_ZMRooXgA5_0),.clk(gclk));
	jdff dff_A_jk4Zfurw9_0(.dout(w_dff_A_ZMRooXgA5_0),.din(w_dff_A_jk4Zfurw9_0),.clk(gclk));
	jdff dff_A_rrQKLtgY1_1(.dout(w_G374_0[1]),.din(w_dff_A_rrQKLtgY1_1),.clk(gclk));
	jdff dff_A_zwQWhkLL1_0(.dout(w_G281_2[0]),.din(w_dff_A_zwQWhkLL1_0),.clk(gclk));
	jdff dff_A_Z2ld8Ms42_2(.dout(w_G281_0[2]),.din(w_dff_A_Z2ld8Ms42_2),.clk(gclk));
	jdff dff_B_CggUUJyJ9_1(.din(n1463),.dout(w_dff_B_CggUUJyJ9_1),.clk(gclk));
	jdff dff_B_McPhVsr13_1(.din(w_dff_B_CggUUJyJ9_1),.dout(w_dff_B_McPhVsr13_1),.clk(gclk));
	jdff dff_B_M2BfNANf4_1(.din(n1486),.dout(w_dff_B_M2BfNANf4_1),.clk(gclk));
	jdff dff_B_xqQZZMkN9_1(.din(n1487),.dout(w_dff_B_xqQZZMkN9_1),.clk(gclk));
	jdff dff_A_2Fos1n793_1(.dout(w_G210_1[1]),.din(w_dff_A_2Fos1n793_1),.clk(gclk));
	jdff dff_A_K1sSTTDM4_1(.dout(w_n543_0[1]),.din(w_dff_A_K1sSTTDM4_1),.clk(gclk));
	jdff dff_A_PpQBE0k26_0(.dout(w_G457_2[0]),.din(w_dff_A_PpQBE0k26_0),.clk(gclk));
	jdff dff_A_ikHJwaSR6_0(.dout(w_G457_0[0]),.din(w_dff_A_ikHJwaSR6_0),.clk(gclk));
	jdff dff_A_5utZaRT63_0(.dout(w_dff_A_ikHJwaSR6_0),.din(w_dff_A_5utZaRT63_0),.clk(gclk));
	jdff dff_A_kIlLJhno4_0(.dout(w_dff_A_5utZaRT63_0),.din(w_dff_A_kIlLJhno4_0),.clk(gclk));
	jdff dff_A_uzNAGVgL4_2(.dout(w_G457_0[2]),.din(w_dff_A_uzNAGVgL4_2),.clk(gclk));
	jdff dff_A_NIHaGDVF2_2(.dout(w_dff_A_uzNAGVgL4_2),.din(w_dff_A_NIHaGDVF2_2),.clk(gclk));
	jdff dff_A_Wvhep0ki2_1(.dout(w_G210_2[1]),.din(w_dff_A_Wvhep0ki2_1),.clk(gclk));
	jdff dff_A_W0Bp2O9F7_2(.dout(w_G210_0[2]),.din(w_dff_A_W0Bp2O9F7_2),.clk(gclk));
	jdff dff_B_drKLrYsS4_1(.din(n1478),.dout(w_dff_B_drKLrYsS4_1),.clk(gclk));
	jdff dff_B_p5kmLarl3_1(.din(w_dff_B_drKLrYsS4_1),.dout(w_dff_B_p5kmLarl3_1),.clk(gclk));
	jdff dff_B_juMTaES87_2(.din(n509),.dout(w_dff_B_juMTaES87_2),.clk(gclk));
	jdff dff_A_FCoTUeF00_0(.dout(w_G468_1[0]),.din(w_dff_A_FCoTUeF00_0),.clk(gclk));
	jdff dff_A_X5buWeyf0_0(.dout(w_dff_A_FCoTUeF00_0),.din(w_dff_A_X5buWeyf0_0),.clk(gclk));
	jdff dff_A_P62yhVsH3_0(.dout(w_dff_A_X5buWeyf0_0),.din(w_dff_A_P62yhVsH3_0),.clk(gclk));
	jdff dff_A_6D3Di4A10_1(.dout(w_G468_1[1]),.din(w_dff_A_6D3Di4A10_1),.clk(gclk));
	jdff dff_B_rzADqUVV1_1(.din(n1474),.dout(w_dff_B_rzADqUVV1_1),.clk(gclk));
	jdff dff_A_sblDCa1a4_1(.dout(w_G218_2[1]),.din(w_dff_A_sblDCa1a4_1),.clk(gclk));
	jdff dff_A_8XrAwFnq4_1(.dout(w_G468_0[1]),.din(w_dff_A_8XrAwFnq4_1),.clk(gclk));
	jdff dff_A_IcWadWZz6_1(.dout(w_dff_A_8XrAwFnq4_1),.din(w_dff_A_IcWadWZz6_1),.clk(gclk));
	jdff dff_A_u3XK0Zs11_2(.dout(w_G468_0[2]),.din(w_dff_A_u3XK0Zs11_2),.clk(gclk));
	jdff dff_A_KoCm3FHP7_2(.dout(w_dff_A_u3XK0Zs11_2),.din(w_dff_A_KoCm3FHP7_2),.clk(gclk));
	jdff dff_A_KNLrAf8K1_2(.dout(w_dff_A_KoCm3FHP7_2),.din(w_dff_A_KNLrAf8K1_2),.clk(gclk));
	jdff dff_A_9a9Fd7d06_0(.dout(w_G218_1[0]),.din(w_dff_A_9a9Fd7d06_0),.clk(gclk));
	jdff dff_B_vP9uQ1Iv3_1(.din(n1468),.dout(w_dff_B_vP9uQ1Iv3_1),.clk(gclk));
	jdff dff_B_Z0Onc9aE6_1(.din(w_dff_B_vP9uQ1Iv3_1),.dout(w_dff_B_Z0Onc9aE6_1),.clk(gclk));
	jdff dff_B_E0EfueVk5_2(.din(n532),.dout(w_dff_B_E0EfueVk5_2),.clk(gclk));
	jdff dff_A_dTobYgT19_0(.dout(w_G422_2[0]),.din(w_dff_A_dTobYgT19_0),.clk(gclk));
	jdff dff_B_PS8UhcAt3_1(.din(n1464),.dout(w_dff_B_PS8UhcAt3_1),.clk(gclk));
	jdff dff_A_8jIdLr0h7_1(.dout(w_G226_2[1]),.din(w_dff_A_8jIdLr0h7_1),.clk(gclk));
	jdff dff_A_Hs8KFHmw9_0(.dout(w_G422_0[0]),.din(w_dff_A_Hs8KFHmw9_0),.clk(gclk));
	jdff dff_A_bi0OmC4g3_0(.dout(w_dff_A_Hs8KFHmw9_0),.din(w_dff_A_bi0OmC4g3_0),.clk(gclk));
	jdff dff_A_dQHbuo6n9_0(.dout(w_dff_A_bi0OmC4g3_0),.din(w_dff_A_dQHbuo6n9_0),.clk(gclk));
	jdff dff_A_1yF74THA3_2(.dout(w_G422_0[2]),.din(w_dff_A_1yF74THA3_2),.clk(gclk));
	jdff dff_A_TPUCpvG71_2(.dout(w_dff_A_1yF74THA3_2),.din(w_dff_A_TPUCpvG71_2),.clk(gclk));
	jdff dff_A_g05iV4qr9_1(.dout(w_G251_4[1]),.din(w_dff_A_g05iV4qr9_1),.clk(gclk));
	jdff dff_A_umsvQfiS2_2(.dout(w_G251_4[2]),.din(w_dff_A_umsvQfiS2_2),.clk(gclk));
	jdff dff_A_K6d3lJfk5_1(.dout(w_G251_1[1]),.din(w_dff_A_K6d3lJfk5_1),.clk(gclk));
	jdff dff_A_CwMNRSJ39_2(.dout(w_G251_1[2]),.din(w_dff_A_CwMNRSJ39_2),.clk(gclk));
	jdff dff_A_6CZxVukQ2_0(.dout(w_G226_1[0]),.din(w_dff_A_6CZxVukQ2_0),.clk(gclk));
	jdff dff_B_J4fIGD0M8_1(.din(n523),.dout(w_dff_B_J4fIGD0M8_1),.clk(gclk));
	jdff dff_B_jPvxMSUl7_1(.din(n524),.dout(w_dff_B_jPvxMSUl7_1),.clk(gclk));
	jdff dff_A_a3DYy5kJ1_0(.dout(w_G446_1[0]),.din(w_dff_A_a3DYy5kJ1_0),.clk(gclk));
	jdff dff_A_WDwUZNW40_0(.dout(w_dff_A_a3DYy5kJ1_0),.din(w_dff_A_WDwUZNW40_0),.clk(gclk));
	jdff dff_A_JOkU9xyp2_0(.dout(w_dff_A_WDwUZNW40_0),.din(w_dff_A_JOkU9xyp2_0),.clk(gclk));
	jdff dff_A_5RAOQJeX5_0(.dout(w_dff_A_JOkU9xyp2_0),.din(w_dff_A_5RAOQJeX5_0),.clk(gclk));
	jdff dff_A_RDfsVM6X2_1(.dout(w_G446_1[1]),.din(w_dff_A_RDfsVM6X2_1),.clk(gclk));
	jdff dff_A_PjIXy07J6_1(.dout(w_dff_A_RDfsVM6X2_1),.din(w_dff_A_PjIXy07J6_1),.clk(gclk));
	jdff dff_A_L84Mh0M65_1(.dout(w_G446_0[1]),.din(w_dff_A_L84Mh0M65_1),.clk(gclk));
	jdff dff_A_1SfBBiXl2_1(.dout(w_dff_A_L84Mh0M65_1),.din(w_dff_A_1SfBBiXl2_1),.clk(gclk));
	jdff dff_A_WTBqrzoc1_1(.dout(w_dff_A_1SfBBiXl2_1),.din(w_dff_A_WTBqrzoc1_1),.clk(gclk));
	jdff dff_A_G6lbEGdA0_1(.dout(w_dff_A_WTBqrzoc1_1),.din(w_dff_A_G6lbEGdA0_1),.clk(gclk));
	jdff dff_A_pJCGRX3l2_2(.dout(w_G446_0[2]),.din(w_dff_A_pJCGRX3l2_2),.clk(gclk));
	jdff dff_A_WL2r15fE7_2(.dout(w_dff_A_pJCGRX3l2_2),.din(w_dff_A_WL2r15fE7_2),.clk(gclk));
	jdff dff_A_yGjiDEl32_2(.dout(w_dff_A_WL2r15fE7_2),.din(w_dff_A_yGjiDEl32_2),.clk(gclk));
	jdff dff_A_jWocplEn0_2(.dout(w_dff_A_yGjiDEl32_2),.din(w_dff_A_jWocplEn0_2),.clk(gclk));
	jdff dff_A_4WsIfzAC9_0(.dout(w_G206_0[0]),.din(w_dff_A_4WsIfzAC9_0),.clk(gclk));
	jdff dff_B_PzdBPeFS4_1(.din(n1458),.dout(w_dff_B_PzdBPeFS4_1),.clk(gclk));
	jdff dff_B_ESW2Jyin8_1(.din(n1459),.dout(w_dff_B_ESW2Jyin8_1),.clk(gclk));
	jdff dff_A_cQwm38V27_0(.dout(w_G242_1[0]),.din(w_dff_A_cQwm38V27_0),.clk(gclk));
	jdff dff_A_Q5zt9qC28_1(.dout(w_G242_1[1]),.din(w_dff_A_Q5zt9qC28_1),.clk(gclk));
	jdff dff_A_HpUvt8bN7_1(.dout(w_G242_0[1]),.din(w_dff_A_HpUvt8bN7_1),.clk(gclk));
	jdff dff_A_L1bi1yru6_2(.dout(w_G242_0[2]),.din(w_dff_A_L1bi1yru6_2),.clk(gclk));
	jdff dff_A_iVswdcIQ0_2(.dout(w_G248_3[2]),.din(w_dff_A_iVswdcIQ0_2),.clk(gclk));
	jdff dff_A_zsQn6rAz9_1(.dout(w_n462_0[1]),.din(w_dff_A_zsQn6rAz9_1),.clk(gclk));
	jdff dff_A_6xE1kp3C5_1(.dout(w_dff_A_zsQn6rAz9_1),.din(w_dff_A_6xE1kp3C5_1),.clk(gclk));
	jdff dff_A_yPEI7Z7s6_1(.dout(w_dff_A_6xE1kp3C5_1),.din(w_dff_A_yPEI7Z7s6_1),.clk(gclk));
	jdff dff_A_IxdqBATw2_1(.dout(w_dff_A_yPEI7Z7s6_1),.din(w_dff_A_IxdqBATw2_1),.clk(gclk));
	jdff dff_A_CvTLzAgQ6_2(.dout(w_n462_0[2]),.din(w_dff_A_CvTLzAgQ6_2),.clk(gclk));
	jdff dff_A_145FCC1R1_0(.dout(w_G435_1[0]),.din(w_dff_A_145FCC1R1_0),.clk(gclk));
	jdff dff_A_E0jDH5bB5_0(.dout(w_dff_A_145FCC1R1_0),.din(w_dff_A_E0jDH5bB5_0),.clk(gclk));
	jdff dff_A_9326LpdF4_0(.dout(w_dff_A_E0jDH5bB5_0),.din(w_dff_A_9326LpdF4_0),.clk(gclk));
	jdff dff_A_BKERlw5H5_0(.dout(w_dff_A_9326LpdF4_0),.din(w_dff_A_BKERlw5H5_0),.clk(gclk));
	jdff dff_A_93DnRBLx5_1(.dout(w_G435_1[1]),.din(w_dff_A_93DnRBLx5_1),.clk(gclk));
	jdff dff_A_6JXrWEu75_1(.dout(w_G435_0[1]),.din(w_dff_A_6JXrWEu75_1),.clk(gclk));
	jdff dff_A_fxjrjCh67_1(.dout(w_dff_A_6JXrWEu75_1),.din(w_dff_A_fxjrjCh67_1),.clk(gclk));
	jdff dff_A_jKyhf4HO5_2(.dout(w_G435_0[2]),.din(w_dff_A_jKyhf4HO5_2),.clk(gclk));
	jdff dff_A_3rQhbg9g1_2(.dout(w_dff_A_jKyhf4HO5_2),.din(w_dff_A_3rQhbg9g1_2),.clk(gclk));
	jdff dff_A_1AEaBP9I6_2(.dout(w_dff_A_3rQhbg9g1_2),.din(w_dff_A_1AEaBP9I6_2),.clk(gclk));
	jdff dff_A_93tWPI9q8_2(.dout(w_dff_A_1AEaBP9I6_2),.din(w_dff_A_93tWPI9q8_2),.clk(gclk));
	jdff dff_A_xBie47Qk2_1(.dout(w_G251_0[1]),.din(w_dff_A_xBie47Qk2_1),.clk(gclk));
	jdff dff_A_EmzcZY9t8_2(.dout(w_G251_0[2]),.din(w_dff_A_EmzcZY9t8_2),.clk(gclk));
	jdff dff_A_y5HQIe6X9_0(.dout(w_G234_2[0]),.din(w_dff_A_y5HQIe6X9_0),.clk(gclk));
	jdff dff_A_5gdKQzfI4_2(.dout(w_G234_0[2]),.din(w_dff_A_5gdKQzfI4_2),.clk(gclk));
	jdff dff_A_MYR8O7PY4_0(.dout(w_G4092_1[0]),.din(w_dff_A_MYR8O7PY4_0),.clk(gclk));
	jdff dff_A_tBnMUCjT0_0(.dout(w_dff_A_MYR8O7PY4_0),.din(w_dff_A_tBnMUCjT0_0),.clk(gclk));
	jdff dff_A_ca1oavqp1_0(.dout(w_dff_A_tBnMUCjT0_0),.din(w_dff_A_ca1oavqp1_0),.clk(gclk));
	jdff dff_A_gnnwhmDU5_0(.dout(w_dff_A_ca1oavqp1_0),.din(w_dff_A_gnnwhmDU5_0),.clk(gclk));
	jdff dff_A_mzXovG4n0_0(.dout(w_dff_A_gnnwhmDU5_0),.din(w_dff_A_mzXovG4n0_0),.clk(gclk));
	jdff dff_A_0hup6JtJ1_0(.dout(w_dff_A_mzXovG4n0_0),.din(w_dff_A_0hup6JtJ1_0),.clk(gclk));
	jdff dff_A_s8Cwsbp59_0(.dout(w_dff_A_0hup6JtJ1_0),.din(w_dff_A_s8Cwsbp59_0),.clk(gclk));
	jdff dff_A_9J9gV7LA9_0(.dout(w_dff_A_s8Cwsbp59_0),.din(w_dff_A_9J9gV7LA9_0),.clk(gclk));
	jdff dff_A_UMSDBrGl4_0(.dout(w_dff_A_9J9gV7LA9_0),.din(w_dff_A_UMSDBrGl4_0),.clk(gclk));
	jdff dff_A_vPrnZUAq7_0(.dout(w_dff_A_UMSDBrGl4_0),.din(w_dff_A_vPrnZUAq7_0),.clk(gclk));
	jdff dff_A_c9obuGxY8_0(.dout(w_dff_A_vPrnZUAq7_0),.din(w_dff_A_c9obuGxY8_0),.clk(gclk));
	jdff dff_A_zdrI3PDS9_1(.dout(w_G4092_1[1]),.din(w_dff_A_zdrI3PDS9_1),.clk(gclk));
	jdff dff_A_BoMi0olI2_0(.dout(w_n999_1[0]),.din(w_dff_A_BoMi0olI2_0),.clk(gclk));
	jdff dff_A_nvTaLphW4_0(.dout(w_dff_A_BoMi0olI2_0),.din(w_dff_A_nvTaLphW4_0),.clk(gclk));
	jdff dff_A_QsJjPFXN5_0(.dout(w_dff_A_nvTaLphW4_0),.din(w_dff_A_QsJjPFXN5_0),.clk(gclk));
	jdff dff_A_j3O89ShG0_0(.dout(w_dff_A_QsJjPFXN5_0),.din(w_dff_A_j3O89ShG0_0),.clk(gclk));
	jdff dff_A_S0vDBA0J9_0(.dout(w_dff_A_j3O89ShG0_0),.din(w_dff_A_S0vDBA0J9_0),.clk(gclk));
	jdff dff_A_iW9HFaD08_0(.dout(w_dff_A_S0vDBA0J9_0),.din(w_dff_A_iW9HFaD08_0),.clk(gclk));
	jdff dff_A_rrccWHtp0_0(.dout(w_dff_A_iW9HFaD08_0),.din(w_dff_A_rrccWHtp0_0),.clk(gclk));
	jdff dff_A_Ikjyje7n8_2(.dout(w_n999_1[2]),.din(w_dff_A_Ikjyje7n8_2),.clk(gclk));
	jdff dff_A_TOXxie9F4_2(.dout(w_dff_A_Ikjyje7n8_2),.din(w_dff_A_TOXxie9F4_2),.clk(gclk));
	jdff dff_A_apl4wpDY6_2(.dout(w_dff_A_TOXxie9F4_2),.din(w_dff_A_apl4wpDY6_2),.clk(gclk));
	jdff dff_A_WaRh8NRP3_2(.dout(w_dff_A_apl4wpDY6_2),.din(w_dff_A_WaRh8NRP3_2),.clk(gclk));
	jdff dff_A_fYJv7fYP2_2(.dout(w_dff_A_WaRh8NRP3_2),.din(w_dff_A_fYJv7fYP2_2),.clk(gclk));
	jdff dff_A_lIlX7Wn50_2(.dout(w_dff_A_fYJv7fYP2_2),.din(w_dff_A_lIlX7Wn50_2),.clk(gclk));
	jdff dff_A_LJliNtAy7_2(.dout(w_dff_A_lIlX7Wn50_2),.din(w_dff_A_LJliNtAy7_2),.clk(gclk));
	jdff dff_A_1bp8sStG3_2(.dout(w_dff_A_LJliNtAy7_2),.din(w_dff_A_1bp8sStG3_2),.clk(gclk));
	jdff dff_A_3DLSZKbP5_2(.dout(w_dff_A_1bp8sStG3_2),.din(w_dff_A_3DLSZKbP5_2),.clk(gclk));
	jdff dff_A_mYHbTfFD9_2(.dout(w_dff_A_3DLSZKbP5_2),.din(w_dff_A_mYHbTfFD9_2),.clk(gclk));
	jdff dff_A_szsVc30w8_2(.dout(w_dff_A_mYHbTfFD9_2),.din(w_dff_A_szsVc30w8_2),.clk(gclk));
	jdff dff_A_F3pXSx5e6_2(.dout(w_dff_A_szsVc30w8_2),.din(w_dff_A_F3pXSx5e6_2),.clk(gclk));
	jdff dff_A_MUqtxYMl0_2(.dout(w_dff_A_F3pXSx5e6_2),.din(w_dff_A_MUqtxYMl0_2),.clk(gclk));
	jdff dff_A_WcsDrtic9_2(.dout(w_dff_A_MUqtxYMl0_2),.din(w_dff_A_WcsDrtic9_2),.clk(gclk));
	jdff dff_A_IvX1SISW3_2(.dout(w_dff_A_WcsDrtic9_2),.din(w_dff_A_IvX1SISW3_2),.clk(gclk));
	jdff dff_A_lAQC2soE4_2(.dout(w_dff_A_IvX1SISW3_2),.din(w_dff_A_lAQC2soE4_2),.clk(gclk));
	jdff dff_A_tRXZgcD47_2(.dout(w_dff_A_lAQC2soE4_2),.din(w_dff_A_tRXZgcD47_2),.clk(gclk));
	jdff dff_A_ZKRb0Opf1_2(.dout(w_dff_A_tRXZgcD47_2),.din(w_dff_A_ZKRb0Opf1_2),.clk(gclk));
	jdff dff_A_A9I8q0GE3_2(.dout(w_dff_A_ZKRb0Opf1_2),.din(w_dff_A_A9I8q0GE3_2),.clk(gclk));
	jdff dff_A_ppyogrIt4_1(.dout(w_n999_0[1]),.din(w_dff_A_ppyogrIt4_1),.clk(gclk));
	jdff dff_A_8b3QS6fT7_1(.dout(w_dff_A_ppyogrIt4_1),.din(w_dff_A_8b3QS6fT7_1),.clk(gclk));
	jdff dff_A_uJdOCJWZ0_1(.dout(w_dff_A_8b3QS6fT7_1),.din(w_dff_A_uJdOCJWZ0_1),.clk(gclk));
	jdff dff_A_Ie5jSKVK5_1(.dout(w_dff_A_uJdOCJWZ0_1),.din(w_dff_A_Ie5jSKVK5_1),.clk(gclk));
	jdff dff_A_b6C8S39j3_1(.dout(w_dff_A_Ie5jSKVK5_1),.din(w_dff_A_b6C8S39j3_1),.clk(gclk));
	jdff dff_A_ciBTzmfd6_1(.dout(w_dff_A_b6C8S39j3_1),.din(w_dff_A_ciBTzmfd6_1),.clk(gclk));
	jdff dff_A_7wqJ9Bsa1_1(.dout(w_dff_A_ciBTzmfd6_1),.din(w_dff_A_7wqJ9Bsa1_1),.clk(gclk));
	jdff dff_A_VVDAx3uY1_1(.dout(w_dff_A_7wqJ9Bsa1_1),.din(w_dff_A_VVDAx3uY1_1),.clk(gclk));
	jdff dff_A_AD2tdsOF8_1(.dout(w_dff_A_VVDAx3uY1_1),.din(w_dff_A_AD2tdsOF8_1),.clk(gclk));
	jdff dff_A_4Xvbbywf5_1(.dout(w_dff_A_AD2tdsOF8_1),.din(w_dff_A_4Xvbbywf5_1),.clk(gclk));
	jdff dff_A_quyEqx870_1(.dout(w_dff_A_4Xvbbywf5_1),.din(w_dff_A_quyEqx870_1),.clk(gclk));
	jdff dff_A_SJc8o4by1_1(.dout(w_dff_A_quyEqx870_1),.din(w_dff_A_SJc8o4by1_1),.clk(gclk));
	jdff dff_A_M7vcgRzt2_1(.dout(w_dff_A_SJc8o4by1_1),.din(w_dff_A_M7vcgRzt2_1),.clk(gclk));
	jdff dff_A_oqBQk2bZ4_1(.dout(w_dff_A_M7vcgRzt2_1),.din(w_dff_A_oqBQk2bZ4_1),.clk(gclk));
	jdff dff_A_jXWACblp2_1(.dout(w_dff_A_oqBQk2bZ4_1),.din(w_dff_A_jXWACblp2_1),.clk(gclk));
	jdff dff_A_I0qaYEYe2_1(.dout(w_dff_A_jXWACblp2_1),.din(w_dff_A_I0qaYEYe2_1),.clk(gclk));
	jdff dff_A_YkaaOJ3u5_1(.dout(w_dff_A_I0qaYEYe2_1),.din(w_dff_A_YkaaOJ3u5_1),.clk(gclk));
	jdff dff_A_kmY6zEzX4_2(.dout(w_n999_0[2]),.din(w_dff_A_kmY6zEzX4_2),.clk(gclk));
	jdff dff_A_YSXjvyKU1_2(.dout(w_dff_A_kmY6zEzX4_2),.din(w_dff_A_YSXjvyKU1_2),.clk(gclk));
	jdff dff_A_WtJarjZg2_2(.dout(w_dff_A_YSXjvyKU1_2),.din(w_dff_A_WtJarjZg2_2),.clk(gclk));
	jdff dff_A_puxkd1286_2(.dout(w_dff_A_WtJarjZg2_2),.din(w_dff_A_puxkd1286_2),.clk(gclk));
	jdff dff_A_LBmRRY814_2(.dout(w_dff_A_puxkd1286_2),.din(w_dff_A_LBmRRY814_2),.clk(gclk));
	jdff dff_A_VQwgBGOY4_2(.dout(w_dff_A_LBmRRY814_2),.din(w_dff_A_VQwgBGOY4_2),.clk(gclk));
	jdff dff_A_Dhp9Osxv4_2(.dout(w_dff_A_VQwgBGOY4_2),.din(w_dff_A_Dhp9Osxv4_2),.clk(gclk));
	jdff dff_A_i7mXiXBc4_2(.dout(w_dff_A_Dhp9Osxv4_2),.din(w_dff_A_i7mXiXBc4_2),.clk(gclk));
	jdff dff_A_pal6TTlv8_2(.dout(w_dff_A_i7mXiXBc4_2),.din(w_dff_A_pal6TTlv8_2),.clk(gclk));
	jdff dff_A_c6gSTUhR6_2(.dout(w_dff_A_pal6TTlv8_2),.din(w_dff_A_c6gSTUhR6_2),.clk(gclk));
	jdff dff_A_KgaFGU7S5_2(.dout(w_dff_A_c6gSTUhR6_2),.din(w_dff_A_KgaFGU7S5_2),.clk(gclk));
	jdff dff_A_UygF6HbI1_1(.dout(w_G1694_0[1]),.din(w_dff_A_UygF6HbI1_1),.clk(gclk));
	jdff dff_A_T9Chpajb1_2(.dout(w_G1691_0[2]),.din(w_dff_A_T9Chpajb1_2),.clk(gclk));
	jdff dff_B_7NAwkOja3_2(.din(n1624),.dout(w_dff_B_7NAwkOja3_2),.clk(gclk));
	jdff dff_B_RNOSPl9T2_2(.din(w_dff_B_7NAwkOja3_2),.dout(w_dff_B_RNOSPl9T2_2),.clk(gclk));
	jdff dff_B_E8goaBHO6_2(.din(w_dff_B_RNOSPl9T2_2),.dout(w_dff_B_E8goaBHO6_2),.clk(gclk));
	jdff dff_B_kD7A8Gu39_2(.din(w_dff_B_E8goaBHO6_2),.dout(w_dff_B_kD7A8Gu39_2),.clk(gclk));
	jdff dff_B_5VSnKx8E3_2(.din(w_dff_B_kD7A8Gu39_2),.dout(w_dff_B_5VSnKx8E3_2),.clk(gclk));
	jdff dff_B_4MJXGFq35_2(.din(w_dff_B_5VSnKx8E3_2),.dout(w_dff_B_4MJXGFq35_2),.clk(gclk));
	jdff dff_B_IgrxV5K80_2(.din(w_dff_B_4MJXGFq35_2),.dout(w_dff_B_IgrxV5K80_2),.clk(gclk));
	jdff dff_B_SQ4edi7L6_2(.din(w_dff_B_IgrxV5K80_2),.dout(w_dff_B_SQ4edi7L6_2),.clk(gclk));
	jdff dff_B_XO2G3nyv7_2(.din(w_dff_B_SQ4edi7L6_2),.dout(w_dff_B_XO2G3nyv7_2),.clk(gclk));
	jdff dff_B_qrXm9Kl65_2(.din(w_dff_B_XO2G3nyv7_2),.dout(w_dff_B_qrXm9Kl65_2),.clk(gclk));
	jdff dff_B_0BJ2ic2B4_2(.din(w_dff_B_qrXm9Kl65_2),.dout(w_dff_B_0BJ2ic2B4_2),.clk(gclk));
	jdff dff_B_W6OUSo1Y4_2(.din(w_dff_B_0BJ2ic2B4_2),.dout(w_dff_B_W6OUSo1Y4_2),.clk(gclk));
	jdff dff_B_ZCsYp7Y29_2(.din(w_dff_B_W6OUSo1Y4_2),.dout(w_dff_B_ZCsYp7Y29_2),.clk(gclk));
	jdff dff_B_myZIM1NK6_2(.din(w_dff_B_ZCsYp7Y29_2),.dout(w_dff_B_myZIM1NK6_2),.clk(gclk));
	jdff dff_B_vet7eIdY0_2(.din(w_dff_B_myZIM1NK6_2),.dout(w_dff_B_vet7eIdY0_2),.clk(gclk));
	jdff dff_B_xwoFjAZC4_2(.din(w_dff_B_vet7eIdY0_2),.dout(w_dff_B_xwoFjAZC4_2),.clk(gclk));
	jdff dff_B_265D6Uep9_2(.din(w_dff_B_xwoFjAZC4_2),.dout(w_dff_B_265D6Uep9_2),.clk(gclk));
	jdff dff_B_ZbQa7PCp5_2(.din(w_dff_B_265D6Uep9_2),.dout(w_dff_B_ZbQa7PCp5_2),.clk(gclk));
	jdff dff_B_tzjSzFk76_2(.din(w_dff_B_ZbQa7PCp5_2),.dout(w_dff_B_tzjSzFk76_2),.clk(gclk));
	jdff dff_B_J7FJ6BEE5_2(.din(w_dff_B_tzjSzFk76_2),.dout(w_dff_B_J7FJ6BEE5_2),.clk(gclk));
	jdff dff_B_FNrz4wUl8_2(.din(w_dff_B_J7FJ6BEE5_2),.dout(w_dff_B_FNrz4wUl8_2),.clk(gclk));
	jdff dff_B_6IqE0GFm7_2(.din(w_dff_B_FNrz4wUl8_2),.dout(w_dff_B_6IqE0GFm7_2),.clk(gclk));
	jdff dff_B_jW1C4NRR4_2(.din(w_dff_B_6IqE0GFm7_2),.dout(w_dff_B_jW1C4NRR4_2),.clk(gclk));
	jdff dff_B_XDizpPKl7_2(.din(w_dff_B_jW1C4NRR4_2),.dout(w_dff_B_XDizpPKl7_2),.clk(gclk));
	jdff dff_A_PxRY2uzP1_2(.dout(w_G137_3[2]),.din(w_dff_A_PxRY2uzP1_2),.clk(gclk));
	jdff dff_A_RDqLBym93_2(.dout(w_dff_A_PxRY2uzP1_2),.din(w_dff_A_RDqLBym93_2),.clk(gclk));
	jdff dff_A_SsyNtHW39_2(.dout(w_dff_A_RDqLBym93_2),.din(w_dff_A_SsyNtHW39_2),.clk(gclk));
	jdff dff_A_5fuBd4Rc0_2(.dout(w_dff_A_SsyNtHW39_2),.din(w_dff_A_5fuBd4Rc0_2),.clk(gclk));
	jdff dff_A_2a4lBvd87_2(.dout(w_dff_A_5fuBd4Rc0_2),.din(w_dff_A_2a4lBvd87_2),.clk(gclk));
	jdff dff_A_lj9TLTIy0_2(.dout(w_dff_A_2a4lBvd87_2),.din(w_dff_A_lj9TLTIy0_2),.clk(gclk));
	jdff dff_A_0VuRgy847_2(.dout(w_dff_A_lj9TLTIy0_2),.din(w_dff_A_0VuRgy847_2),.clk(gclk));
	jdff dff_A_YrtCm23Q6_2(.dout(w_dff_A_0VuRgy847_2),.din(w_dff_A_YrtCm23Q6_2),.clk(gclk));
	jdff dff_A_WAFqwUEP9_2(.dout(w_dff_A_YrtCm23Q6_2),.din(w_dff_A_WAFqwUEP9_2),.clk(gclk));
	jdff dff_A_LD2TpBWz4_2(.dout(w_dff_A_WAFqwUEP9_2),.din(w_dff_A_LD2TpBWz4_2),.clk(gclk));
	jdff dff_A_k2vTd8Xu7_2(.dout(w_dff_A_LD2TpBWz4_2),.din(w_dff_A_k2vTd8Xu7_2),.clk(gclk));
	jdff dff_A_KA52KHCR6_2(.dout(w_dff_A_k2vTd8Xu7_2),.din(w_dff_A_KA52KHCR6_2),.clk(gclk));
	jdff dff_A_NGxsdPAI3_2(.dout(w_dff_A_KA52KHCR6_2),.din(w_dff_A_NGxsdPAI3_2),.clk(gclk));
	jdff dff_A_UaBDrsHk9_2(.dout(w_dff_A_NGxsdPAI3_2),.din(w_dff_A_UaBDrsHk9_2),.clk(gclk));
	jdff dff_A_Sz8mgOhv0_2(.dout(w_dff_A_UaBDrsHk9_2),.din(w_dff_A_Sz8mgOhv0_2),.clk(gclk));
	jdff dff_A_dUYkmnTs3_2(.dout(w_dff_A_Sz8mgOhv0_2),.din(w_dff_A_dUYkmnTs3_2),.clk(gclk));
	jdff dff_A_FGNPx9p15_2(.dout(w_dff_A_dUYkmnTs3_2),.din(w_dff_A_FGNPx9p15_2),.clk(gclk));
	jdff dff_A_i4GR8iVn4_2(.dout(w_dff_A_FGNPx9p15_2),.din(w_dff_A_i4GR8iVn4_2),.clk(gclk));
	jdff dff_A_DUw5Epjj0_2(.dout(w_dff_A_i4GR8iVn4_2),.din(w_dff_A_DUw5Epjj0_2),.clk(gclk));
	jdff dff_A_hhI9bfnN0_2(.dout(w_dff_A_DUw5Epjj0_2),.din(w_dff_A_hhI9bfnN0_2),.clk(gclk));
	jdff dff_A_zy1gQ3ov1_2(.dout(w_dff_A_hhI9bfnN0_2),.din(w_dff_A_zy1gQ3ov1_2),.clk(gclk));
	jdff dff_A_Uyj3YvV44_2(.dout(w_dff_A_zy1gQ3ov1_2),.din(w_dff_A_Uyj3YvV44_2),.clk(gclk));
	jdff dff_A_LoVGMRWh5_2(.dout(w_dff_A_Uyj3YvV44_2),.din(w_dff_A_LoVGMRWh5_2),.clk(gclk));
	jdff dff_A_fuRUgZwW6_0(.dout(w_G137_0[0]),.din(w_dff_A_fuRUgZwW6_0),.clk(gclk));
	jdff dff_A_pHqyWyMF6_0(.dout(w_dff_A_fuRUgZwW6_0),.din(w_dff_A_pHqyWyMF6_0),.clk(gclk));
	jdff dff_A_BA92vPRz0_0(.dout(w_dff_A_pHqyWyMF6_0),.din(w_dff_A_BA92vPRz0_0),.clk(gclk));
	jdff dff_A_bhah2Hxn6_0(.dout(w_dff_A_BA92vPRz0_0),.din(w_dff_A_bhah2Hxn6_0),.clk(gclk));
	jdff dff_A_sKt9M6kK5_0(.dout(w_dff_A_bhah2Hxn6_0),.din(w_dff_A_sKt9M6kK5_0),.clk(gclk));
	jdff dff_A_q9h7freb6_0(.dout(w_dff_A_sKt9M6kK5_0),.din(w_dff_A_q9h7freb6_0),.clk(gclk));
	jdff dff_A_e9Y3whVb1_0(.dout(w_dff_A_q9h7freb6_0),.din(w_dff_A_e9Y3whVb1_0),.clk(gclk));
	jdff dff_A_SscALKln3_0(.dout(w_dff_A_e9Y3whVb1_0),.din(w_dff_A_SscALKln3_0),.clk(gclk));
	jdff dff_A_mv9Qe9hZ8_0(.dout(w_dff_A_SscALKln3_0),.din(w_dff_A_mv9Qe9hZ8_0),.clk(gclk));
	jdff dff_A_5RacaMh79_0(.dout(w_dff_A_mv9Qe9hZ8_0),.din(w_dff_A_5RacaMh79_0),.clk(gclk));
	jdff dff_A_OhqbPePe9_0(.dout(w_dff_A_5RacaMh79_0),.din(w_dff_A_OhqbPePe9_0),.clk(gclk));
	jdff dff_A_yfeF5XSX1_0(.dout(w_dff_A_OhqbPePe9_0),.din(w_dff_A_yfeF5XSX1_0),.clk(gclk));
	jdff dff_A_hhoDlKC51_0(.dout(w_dff_A_yfeF5XSX1_0),.din(w_dff_A_hhoDlKC51_0),.clk(gclk));
	jdff dff_A_cag0b5qf4_0(.dout(w_dff_A_hhoDlKC51_0),.din(w_dff_A_cag0b5qf4_0),.clk(gclk));
	jdff dff_A_PasI4ITh8_0(.dout(w_dff_A_cag0b5qf4_0),.din(w_dff_A_PasI4ITh8_0),.clk(gclk));
	jdff dff_A_Y7lYWyOM7_0(.dout(w_dff_A_PasI4ITh8_0),.din(w_dff_A_Y7lYWyOM7_0),.clk(gclk));
	jdff dff_A_hyar6FWU7_1(.dout(w_G137_0[1]),.din(w_dff_A_hyar6FWU7_1),.clk(gclk));
	jdff dff_A_L5vcJehQ6_1(.dout(w_dff_A_hyar6FWU7_1),.din(w_dff_A_L5vcJehQ6_1),.clk(gclk));
	jdff dff_A_OCY1RXdO1_1(.dout(w_dff_A_L5vcJehQ6_1),.din(w_dff_A_OCY1RXdO1_1),.clk(gclk));
	jdff dff_A_jRZYI5ML9_1(.dout(w_dff_A_OCY1RXdO1_1),.din(w_dff_A_jRZYI5ML9_1),.clk(gclk));
	jdff dff_A_fN4BFm7N2_1(.dout(w_dff_A_jRZYI5ML9_1),.din(w_dff_A_fN4BFm7N2_1),.clk(gclk));
	jdff dff_A_KRs8Gbmq9_1(.dout(w_dff_A_fN4BFm7N2_1),.din(w_dff_A_KRs8Gbmq9_1),.clk(gclk));
	jdff dff_A_tgGPUvU04_1(.dout(w_dff_A_KRs8Gbmq9_1),.din(w_dff_A_tgGPUvU04_1),.clk(gclk));
	jdff dff_A_4elJ960V5_1(.dout(w_dff_A_tgGPUvU04_1),.din(w_dff_A_4elJ960V5_1),.clk(gclk));
	jdff dff_A_SxVrNxLb4_1(.dout(w_dff_A_4elJ960V5_1),.din(w_dff_A_SxVrNxLb4_1),.clk(gclk));
	jdff dff_A_QQuo31aY2_1(.dout(w_dff_A_SxVrNxLb4_1),.din(w_dff_A_QQuo31aY2_1),.clk(gclk));
	jdff dff_A_qfPzuRhQ3_1(.dout(w_dff_A_QQuo31aY2_1),.din(w_dff_A_qfPzuRhQ3_1),.clk(gclk));
	jdff dff_A_cb5G565l2_1(.dout(w_dff_A_3RHCVIMc4_0),.din(w_dff_A_cb5G565l2_1),.clk(gclk));
	jdff dff_A_3RHCVIMc4_0(.dout(w_dff_A_ISAWvOxo3_0),.din(w_dff_A_3RHCVIMc4_0),.clk(gclk));
	jdff dff_A_ISAWvOxo3_0(.dout(w_dff_A_9Y9yy8zR4_0),.din(w_dff_A_ISAWvOxo3_0),.clk(gclk));
	jdff dff_A_9Y9yy8zR4_0(.dout(w_dff_A_3irR0KP65_0),.din(w_dff_A_9Y9yy8zR4_0),.clk(gclk));
	jdff dff_A_3irR0KP65_0(.dout(w_dff_A_JhPOMwGL6_0),.din(w_dff_A_3irR0KP65_0),.clk(gclk));
	jdff dff_A_JhPOMwGL6_0(.dout(w_dff_A_hYbRxPIL1_0),.din(w_dff_A_JhPOMwGL6_0),.clk(gclk));
	jdff dff_A_hYbRxPIL1_0(.dout(w_dff_A_mSDgAZtS5_0),.din(w_dff_A_hYbRxPIL1_0),.clk(gclk));
	jdff dff_A_mSDgAZtS5_0(.dout(w_dff_A_1nelbSrb4_0),.din(w_dff_A_mSDgAZtS5_0),.clk(gclk));
	jdff dff_A_1nelbSrb4_0(.dout(w_dff_A_y309zFKo4_0),.din(w_dff_A_1nelbSrb4_0),.clk(gclk));
	jdff dff_A_y309zFKo4_0(.dout(w_dff_A_B5kI9FwV9_0),.din(w_dff_A_y309zFKo4_0),.clk(gclk));
	jdff dff_A_B5kI9FwV9_0(.dout(w_dff_A_ny7ajQjk6_0),.din(w_dff_A_B5kI9FwV9_0),.clk(gclk));
	jdff dff_A_ny7ajQjk6_0(.dout(w_dff_A_AJE5QduK8_0),.din(w_dff_A_ny7ajQjk6_0),.clk(gclk));
	jdff dff_A_AJE5QduK8_0(.dout(w_dff_A_t07HMYYV8_0),.din(w_dff_A_AJE5QduK8_0),.clk(gclk));
	jdff dff_A_t07HMYYV8_0(.dout(w_dff_A_Vn6bD5F74_0),.din(w_dff_A_t07HMYYV8_0),.clk(gclk));
	jdff dff_A_Vn6bD5F74_0(.dout(w_dff_A_sQKv8hqb0_0),.din(w_dff_A_Vn6bD5F74_0),.clk(gclk));
	jdff dff_A_sQKv8hqb0_0(.dout(w_dff_A_XFJScwnh8_0),.din(w_dff_A_sQKv8hqb0_0),.clk(gclk));
	jdff dff_A_XFJScwnh8_0(.dout(w_dff_A_PLWBdEet3_0),.din(w_dff_A_XFJScwnh8_0),.clk(gclk));
	jdff dff_A_PLWBdEet3_0(.dout(w_dff_A_xeKRPcYs3_0),.din(w_dff_A_PLWBdEet3_0),.clk(gclk));
	jdff dff_A_xeKRPcYs3_0(.dout(w_dff_A_p16RC3072_0),.din(w_dff_A_xeKRPcYs3_0),.clk(gclk));
	jdff dff_A_p16RC3072_0(.dout(w_dff_A_oizumvxp6_0),.din(w_dff_A_p16RC3072_0),.clk(gclk));
	jdff dff_A_oizumvxp6_0(.dout(w_dff_A_0HHe19PL3_0),.din(w_dff_A_oizumvxp6_0),.clk(gclk));
	jdff dff_A_0HHe19PL3_0(.dout(w_dff_A_AstgGGaD1_0),.din(w_dff_A_0HHe19PL3_0),.clk(gclk));
	jdff dff_A_AstgGGaD1_0(.dout(w_dff_A_pCLflLim8_0),.din(w_dff_A_AstgGGaD1_0),.clk(gclk));
	jdff dff_A_pCLflLim8_0(.dout(w_dff_A_4HYNfnur1_0),.din(w_dff_A_pCLflLim8_0),.clk(gclk));
	jdff dff_A_4HYNfnur1_0(.dout(G144),.din(w_dff_A_4HYNfnur1_0),.clk(gclk));
	jdff dff_A_HUppY1yx4_1(.dout(w_dff_A_JkxxEBys7_0),.din(w_dff_A_HUppY1yx4_1),.clk(gclk));
	jdff dff_A_JkxxEBys7_0(.dout(w_dff_A_q0n3POXW3_0),.din(w_dff_A_JkxxEBys7_0),.clk(gclk));
	jdff dff_A_q0n3POXW3_0(.dout(w_dff_A_cehktUxD0_0),.din(w_dff_A_q0n3POXW3_0),.clk(gclk));
	jdff dff_A_cehktUxD0_0(.dout(w_dff_A_M44KfxPO4_0),.din(w_dff_A_cehktUxD0_0),.clk(gclk));
	jdff dff_A_M44KfxPO4_0(.dout(w_dff_A_5bBBem6b8_0),.din(w_dff_A_M44KfxPO4_0),.clk(gclk));
	jdff dff_A_5bBBem6b8_0(.dout(w_dff_A_GPrB7LAM2_0),.din(w_dff_A_5bBBem6b8_0),.clk(gclk));
	jdff dff_A_GPrB7LAM2_0(.dout(w_dff_A_TGBFibZw6_0),.din(w_dff_A_GPrB7LAM2_0),.clk(gclk));
	jdff dff_A_TGBFibZw6_0(.dout(w_dff_A_apRmpxY45_0),.din(w_dff_A_TGBFibZw6_0),.clk(gclk));
	jdff dff_A_apRmpxY45_0(.dout(w_dff_A_T89OFW921_0),.din(w_dff_A_apRmpxY45_0),.clk(gclk));
	jdff dff_A_T89OFW921_0(.dout(w_dff_A_8yYH2IQ27_0),.din(w_dff_A_T89OFW921_0),.clk(gclk));
	jdff dff_A_8yYH2IQ27_0(.dout(w_dff_A_R4kJCjqO1_0),.din(w_dff_A_8yYH2IQ27_0),.clk(gclk));
	jdff dff_A_R4kJCjqO1_0(.dout(w_dff_A_q9P3EMcU5_0),.din(w_dff_A_R4kJCjqO1_0),.clk(gclk));
	jdff dff_A_q9P3EMcU5_0(.dout(w_dff_A_PCp7I8GM7_0),.din(w_dff_A_q9P3EMcU5_0),.clk(gclk));
	jdff dff_A_PCp7I8GM7_0(.dout(w_dff_A_VsAtRIEU7_0),.din(w_dff_A_PCp7I8GM7_0),.clk(gclk));
	jdff dff_A_VsAtRIEU7_0(.dout(w_dff_A_hIBPr7HU2_0),.din(w_dff_A_VsAtRIEU7_0),.clk(gclk));
	jdff dff_A_hIBPr7HU2_0(.dout(w_dff_A_0c2WevMi6_0),.din(w_dff_A_hIBPr7HU2_0),.clk(gclk));
	jdff dff_A_0c2WevMi6_0(.dout(w_dff_A_x2swy0xC4_0),.din(w_dff_A_0c2WevMi6_0),.clk(gclk));
	jdff dff_A_x2swy0xC4_0(.dout(w_dff_A_Q5s0T84Y1_0),.din(w_dff_A_x2swy0xC4_0),.clk(gclk));
	jdff dff_A_Q5s0T84Y1_0(.dout(w_dff_A_SZdqoSlS9_0),.din(w_dff_A_Q5s0T84Y1_0),.clk(gclk));
	jdff dff_A_SZdqoSlS9_0(.dout(w_dff_A_Ih4eRD3R7_0),.din(w_dff_A_SZdqoSlS9_0),.clk(gclk));
	jdff dff_A_Ih4eRD3R7_0(.dout(w_dff_A_ViwAE7JN3_0),.din(w_dff_A_Ih4eRD3R7_0),.clk(gclk));
	jdff dff_A_ViwAE7JN3_0(.dout(w_dff_A_wIcM7nXD6_0),.din(w_dff_A_ViwAE7JN3_0),.clk(gclk));
	jdff dff_A_wIcM7nXD6_0(.dout(w_dff_A_gR3xRhPa6_0),.din(w_dff_A_wIcM7nXD6_0),.clk(gclk));
	jdff dff_A_gR3xRhPa6_0(.dout(w_dff_A_s7fIBDsj0_0),.din(w_dff_A_gR3xRhPa6_0),.clk(gclk));
	jdff dff_A_s7fIBDsj0_0(.dout(G298),.din(w_dff_A_s7fIBDsj0_0),.clk(gclk));
	jdff dff_A_bgbfZxUg8_1(.dout(w_dff_A_3iukpOH64_0),.din(w_dff_A_bgbfZxUg8_1),.clk(gclk));
	jdff dff_A_3iukpOH64_0(.dout(w_dff_A_N2tLGc6e0_0),.din(w_dff_A_3iukpOH64_0),.clk(gclk));
	jdff dff_A_N2tLGc6e0_0(.dout(w_dff_A_382wXYrB6_0),.din(w_dff_A_N2tLGc6e0_0),.clk(gclk));
	jdff dff_A_382wXYrB6_0(.dout(w_dff_A_wognC2Q89_0),.din(w_dff_A_382wXYrB6_0),.clk(gclk));
	jdff dff_A_wognC2Q89_0(.dout(w_dff_A_DmT4I2r63_0),.din(w_dff_A_wognC2Q89_0),.clk(gclk));
	jdff dff_A_DmT4I2r63_0(.dout(w_dff_A_AQZkrOwm2_0),.din(w_dff_A_DmT4I2r63_0),.clk(gclk));
	jdff dff_A_AQZkrOwm2_0(.dout(w_dff_A_UTpaR8fz6_0),.din(w_dff_A_AQZkrOwm2_0),.clk(gclk));
	jdff dff_A_UTpaR8fz6_0(.dout(w_dff_A_wrgdHrHz8_0),.din(w_dff_A_UTpaR8fz6_0),.clk(gclk));
	jdff dff_A_wrgdHrHz8_0(.dout(w_dff_A_HdUoc6hb0_0),.din(w_dff_A_wrgdHrHz8_0),.clk(gclk));
	jdff dff_A_HdUoc6hb0_0(.dout(w_dff_A_Zwd2PX9a0_0),.din(w_dff_A_HdUoc6hb0_0),.clk(gclk));
	jdff dff_A_Zwd2PX9a0_0(.dout(w_dff_A_2BwNehvp7_0),.din(w_dff_A_Zwd2PX9a0_0),.clk(gclk));
	jdff dff_A_2BwNehvp7_0(.dout(w_dff_A_0h2tkLmC1_0),.din(w_dff_A_2BwNehvp7_0),.clk(gclk));
	jdff dff_A_0h2tkLmC1_0(.dout(w_dff_A_iXK43Zs41_0),.din(w_dff_A_0h2tkLmC1_0),.clk(gclk));
	jdff dff_A_iXK43Zs41_0(.dout(w_dff_A_OmLbW4Iy4_0),.din(w_dff_A_iXK43Zs41_0),.clk(gclk));
	jdff dff_A_OmLbW4Iy4_0(.dout(w_dff_A_HubVTvWd0_0),.din(w_dff_A_OmLbW4Iy4_0),.clk(gclk));
	jdff dff_A_HubVTvWd0_0(.dout(w_dff_A_KxWanDai5_0),.din(w_dff_A_HubVTvWd0_0),.clk(gclk));
	jdff dff_A_KxWanDai5_0(.dout(w_dff_A_hIH32iKu8_0),.din(w_dff_A_KxWanDai5_0),.clk(gclk));
	jdff dff_A_hIH32iKu8_0(.dout(w_dff_A_4PpY3odB6_0),.din(w_dff_A_hIH32iKu8_0),.clk(gclk));
	jdff dff_A_4PpY3odB6_0(.dout(w_dff_A_qb9watoE0_0),.din(w_dff_A_4PpY3odB6_0),.clk(gclk));
	jdff dff_A_qb9watoE0_0(.dout(w_dff_A_DDikxFB50_0),.din(w_dff_A_qb9watoE0_0),.clk(gclk));
	jdff dff_A_DDikxFB50_0(.dout(w_dff_A_0HXgrLo47_0),.din(w_dff_A_DDikxFB50_0),.clk(gclk));
	jdff dff_A_0HXgrLo47_0(.dout(w_dff_A_ioyeN63Z6_0),.din(w_dff_A_0HXgrLo47_0),.clk(gclk));
	jdff dff_A_ioyeN63Z6_0(.dout(w_dff_A_JN965QCk0_0),.din(w_dff_A_ioyeN63Z6_0),.clk(gclk));
	jdff dff_A_JN965QCk0_0(.dout(w_dff_A_a7Abiasf0_0),.din(w_dff_A_JN965QCk0_0),.clk(gclk));
	jdff dff_A_a7Abiasf0_0(.dout(G973),.din(w_dff_A_a7Abiasf0_0),.clk(gclk));
	jdff dff_A_xnuHcXtR9_1(.dout(w_dff_A_Spw7PSBT8_0),.din(w_dff_A_xnuHcXtR9_1),.clk(gclk));
	jdff dff_A_Spw7PSBT8_0(.dout(w_dff_A_Xd0gO3jg3_0),.din(w_dff_A_Spw7PSBT8_0),.clk(gclk));
	jdff dff_A_Xd0gO3jg3_0(.dout(w_dff_A_dYJW6aHA3_0),.din(w_dff_A_Xd0gO3jg3_0),.clk(gclk));
	jdff dff_A_dYJW6aHA3_0(.dout(w_dff_A_wyOinnPZ9_0),.din(w_dff_A_dYJW6aHA3_0),.clk(gclk));
	jdff dff_A_wyOinnPZ9_0(.dout(w_dff_A_FAJL4wXN9_0),.din(w_dff_A_wyOinnPZ9_0),.clk(gclk));
	jdff dff_A_FAJL4wXN9_0(.dout(w_dff_A_UqfFpiUn5_0),.din(w_dff_A_FAJL4wXN9_0),.clk(gclk));
	jdff dff_A_UqfFpiUn5_0(.dout(w_dff_A_waGytCvG3_0),.din(w_dff_A_UqfFpiUn5_0),.clk(gclk));
	jdff dff_A_waGytCvG3_0(.dout(w_dff_A_d59ubn9F1_0),.din(w_dff_A_waGytCvG3_0),.clk(gclk));
	jdff dff_A_d59ubn9F1_0(.dout(w_dff_A_NaNrlEHF1_0),.din(w_dff_A_d59ubn9F1_0),.clk(gclk));
	jdff dff_A_NaNrlEHF1_0(.dout(w_dff_A_seAYEsp76_0),.din(w_dff_A_NaNrlEHF1_0),.clk(gclk));
	jdff dff_A_seAYEsp76_0(.dout(w_dff_A_T1823c4M5_0),.din(w_dff_A_seAYEsp76_0),.clk(gclk));
	jdff dff_A_T1823c4M5_0(.dout(w_dff_A_PHux2mT88_0),.din(w_dff_A_T1823c4M5_0),.clk(gclk));
	jdff dff_A_PHux2mT88_0(.dout(w_dff_A_GkeuVsPt3_0),.din(w_dff_A_PHux2mT88_0),.clk(gclk));
	jdff dff_A_GkeuVsPt3_0(.dout(w_dff_A_LXypeAx94_0),.din(w_dff_A_GkeuVsPt3_0),.clk(gclk));
	jdff dff_A_LXypeAx94_0(.dout(w_dff_A_He3iXIhu0_0),.din(w_dff_A_LXypeAx94_0),.clk(gclk));
	jdff dff_A_He3iXIhu0_0(.dout(w_dff_A_dhrAaJGI9_0),.din(w_dff_A_He3iXIhu0_0),.clk(gclk));
	jdff dff_A_dhrAaJGI9_0(.dout(w_dff_A_5jo1I6l73_0),.din(w_dff_A_dhrAaJGI9_0),.clk(gclk));
	jdff dff_A_5jo1I6l73_0(.dout(w_dff_A_iVV58X7c6_0),.din(w_dff_A_5jo1I6l73_0),.clk(gclk));
	jdff dff_A_iVV58X7c6_0(.dout(w_dff_A_WSa20qeo2_0),.din(w_dff_A_iVV58X7c6_0),.clk(gclk));
	jdff dff_A_WSa20qeo2_0(.dout(w_dff_A_xkFAl7Fg1_0),.din(w_dff_A_WSa20qeo2_0),.clk(gclk));
	jdff dff_A_xkFAl7Fg1_0(.dout(w_dff_A_9CD5bB7k9_0),.din(w_dff_A_xkFAl7Fg1_0),.clk(gclk));
	jdff dff_A_9CD5bB7k9_0(.dout(w_dff_A_JVyna9ul2_0),.din(w_dff_A_9CD5bB7k9_0),.clk(gclk));
	jdff dff_A_JVyna9ul2_0(.dout(w_dff_A_RPmdp4rG3_0),.din(w_dff_A_JVyna9ul2_0),.clk(gclk));
	jdff dff_A_RPmdp4rG3_0(.dout(w_dff_A_S8O1fbJY7_0),.din(w_dff_A_RPmdp4rG3_0),.clk(gclk));
	jdff dff_A_S8O1fbJY7_0(.dout(G594),.din(w_dff_A_S8O1fbJY7_0),.clk(gclk));
	jdff dff_A_ywNt4EiO1_1(.dout(w_dff_A_VVNM3nxk7_0),.din(w_dff_A_ywNt4EiO1_1),.clk(gclk));
	jdff dff_A_VVNM3nxk7_0(.dout(w_dff_A_mmjtDoSM2_0),.din(w_dff_A_VVNM3nxk7_0),.clk(gclk));
	jdff dff_A_mmjtDoSM2_0(.dout(w_dff_A_b2Sh4jsb2_0),.din(w_dff_A_mmjtDoSM2_0),.clk(gclk));
	jdff dff_A_b2Sh4jsb2_0(.dout(w_dff_A_6hYJGPOL7_0),.din(w_dff_A_b2Sh4jsb2_0),.clk(gclk));
	jdff dff_A_6hYJGPOL7_0(.dout(w_dff_A_5umprcy05_0),.din(w_dff_A_6hYJGPOL7_0),.clk(gclk));
	jdff dff_A_5umprcy05_0(.dout(w_dff_A_D5UXYMnK7_0),.din(w_dff_A_5umprcy05_0),.clk(gclk));
	jdff dff_A_D5UXYMnK7_0(.dout(w_dff_A_bMwFVns33_0),.din(w_dff_A_D5UXYMnK7_0),.clk(gclk));
	jdff dff_A_bMwFVns33_0(.dout(w_dff_A_40wmxGgT3_0),.din(w_dff_A_bMwFVns33_0),.clk(gclk));
	jdff dff_A_40wmxGgT3_0(.dout(w_dff_A_fgKMQkj48_0),.din(w_dff_A_40wmxGgT3_0),.clk(gclk));
	jdff dff_A_fgKMQkj48_0(.dout(w_dff_A_0ZQxhR5e9_0),.din(w_dff_A_fgKMQkj48_0),.clk(gclk));
	jdff dff_A_0ZQxhR5e9_0(.dout(w_dff_A_8dPtbYpI0_0),.din(w_dff_A_0ZQxhR5e9_0),.clk(gclk));
	jdff dff_A_8dPtbYpI0_0(.dout(w_dff_A_Fq3HN0CL1_0),.din(w_dff_A_8dPtbYpI0_0),.clk(gclk));
	jdff dff_A_Fq3HN0CL1_0(.dout(w_dff_A_Bd05Wsy23_0),.din(w_dff_A_Fq3HN0CL1_0),.clk(gclk));
	jdff dff_A_Bd05Wsy23_0(.dout(w_dff_A_ALM58iN24_0),.din(w_dff_A_Bd05Wsy23_0),.clk(gclk));
	jdff dff_A_ALM58iN24_0(.dout(w_dff_A_6t3ZeJx36_0),.din(w_dff_A_ALM58iN24_0),.clk(gclk));
	jdff dff_A_6t3ZeJx36_0(.dout(w_dff_A_g3hPaqWW1_0),.din(w_dff_A_6t3ZeJx36_0),.clk(gclk));
	jdff dff_A_g3hPaqWW1_0(.dout(w_dff_A_vz1QgAqq4_0),.din(w_dff_A_g3hPaqWW1_0),.clk(gclk));
	jdff dff_A_vz1QgAqq4_0(.dout(w_dff_A_klPbOt779_0),.din(w_dff_A_vz1QgAqq4_0),.clk(gclk));
	jdff dff_A_klPbOt779_0(.dout(w_dff_A_XQsxFS3V8_0),.din(w_dff_A_klPbOt779_0),.clk(gclk));
	jdff dff_A_XQsxFS3V8_0(.dout(w_dff_A_iP1vrYH23_0),.din(w_dff_A_XQsxFS3V8_0),.clk(gclk));
	jdff dff_A_iP1vrYH23_0(.dout(w_dff_A_koqwoAFO7_0),.din(w_dff_A_iP1vrYH23_0),.clk(gclk));
	jdff dff_A_koqwoAFO7_0(.dout(w_dff_A_LkXpchdi4_0),.din(w_dff_A_koqwoAFO7_0),.clk(gclk));
	jdff dff_A_LkXpchdi4_0(.dout(w_dff_A_IOYig3dL4_0),.din(w_dff_A_LkXpchdi4_0),.clk(gclk));
	jdff dff_A_IOYig3dL4_0(.dout(w_dff_A_RiPmO5jO7_0),.din(w_dff_A_IOYig3dL4_0),.clk(gclk));
	jdff dff_A_RiPmO5jO7_0(.dout(G599),.din(w_dff_A_RiPmO5jO7_0),.clk(gclk));
	jdff dff_A_wEbXZwDn0_1(.dout(w_dff_A_HSvLcFhP5_0),.din(w_dff_A_wEbXZwDn0_1),.clk(gclk));
	jdff dff_A_HSvLcFhP5_0(.dout(w_dff_A_BCZSTrqm4_0),.din(w_dff_A_HSvLcFhP5_0),.clk(gclk));
	jdff dff_A_BCZSTrqm4_0(.dout(w_dff_A_311DW8Cb4_0),.din(w_dff_A_BCZSTrqm4_0),.clk(gclk));
	jdff dff_A_311DW8Cb4_0(.dout(w_dff_A_EM8T03Ww0_0),.din(w_dff_A_311DW8Cb4_0),.clk(gclk));
	jdff dff_A_EM8T03Ww0_0(.dout(w_dff_A_7mfxGjPM5_0),.din(w_dff_A_EM8T03Ww0_0),.clk(gclk));
	jdff dff_A_7mfxGjPM5_0(.dout(w_dff_A_yGoa4VFG3_0),.din(w_dff_A_7mfxGjPM5_0),.clk(gclk));
	jdff dff_A_yGoa4VFG3_0(.dout(w_dff_A_BCLyTzPz5_0),.din(w_dff_A_yGoa4VFG3_0),.clk(gclk));
	jdff dff_A_BCLyTzPz5_0(.dout(w_dff_A_dSxoOqCP5_0),.din(w_dff_A_BCLyTzPz5_0),.clk(gclk));
	jdff dff_A_dSxoOqCP5_0(.dout(w_dff_A_AaFa3NAg8_0),.din(w_dff_A_dSxoOqCP5_0),.clk(gclk));
	jdff dff_A_AaFa3NAg8_0(.dout(w_dff_A_onjYlMBl9_0),.din(w_dff_A_AaFa3NAg8_0),.clk(gclk));
	jdff dff_A_onjYlMBl9_0(.dout(w_dff_A_XfTgz1Vg6_0),.din(w_dff_A_onjYlMBl9_0),.clk(gclk));
	jdff dff_A_XfTgz1Vg6_0(.dout(w_dff_A_JncHxJWa5_0),.din(w_dff_A_XfTgz1Vg6_0),.clk(gclk));
	jdff dff_A_JncHxJWa5_0(.dout(w_dff_A_1g6dkrv70_0),.din(w_dff_A_JncHxJWa5_0),.clk(gclk));
	jdff dff_A_1g6dkrv70_0(.dout(w_dff_A_Yvh6AOlh0_0),.din(w_dff_A_1g6dkrv70_0),.clk(gclk));
	jdff dff_A_Yvh6AOlh0_0(.dout(w_dff_A_aSNyovvN8_0),.din(w_dff_A_Yvh6AOlh0_0),.clk(gclk));
	jdff dff_A_aSNyovvN8_0(.dout(w_dff_A_Ev5iRoSw1_0),.din(w_dff_A_aSNyovvN8_0),.clk(gclk));
	jdff dff_A_Ev5iRoSw1_0(.dout(w_dff_A_ENUbs8W56_0),.din(w_dff_A_Ev5iRoSw1_0),.clk(gclk));
	jdff dff_A_ENUbs8W56_0(.dout(w_dff_A_Wuoudu227_0),.din(w_dff_A_ENUbs8W56_0),.clk(gclk));
	jdff dff_A_Wuoudu227_0(.dout(w_dff_A_rJulTKrw4_0),.din(w_dff_A_Wuoudu227_0),.clk(gclk));
	jdff dff_A_rJulTKrw4_0(.dout(w_dff_A_gOIlfFh00_0),.din(w_dff_A_rJulTKrw4_0),.clk(gclk));
	jdff dff_A_gOIlfFh00_0(.dout(w_dff_A_NwZT58qA1_0),.din(w_dff_A_gOIlfFh00_0),.clk(gclk));
	jdff dff_A_NwZT58qA1_0(.dout(w_dff_A_shR6BZ6X7_0),.din(w_dff_A_NwZT58qA1_0),.clk(gclk));
	jdff dff_A_shR6BZ6X7_0(.dout(w_dff_A_YY9zUnjr2_0),.din(w_dff_A_shR6BZ6X7_0),.clk(gclk));
	jdff dff_A_YY9zUnjr2_0(.dout(w_dff_A_jrqvbr3c8_0),.din(w_dff_A_YY9zUnjr2_0),.clk(gclk));
	jdff dff_A_jrqvbr3c8_0(.dout(G600),.din(w_dff_A_jrqvbr3c8_0),.clk(gclk));
	jdff dff_A_XBKdFEY12_1(.dout(w_dff_A_W3blJKaT6_0),.din(w_dff_A_XBKdFEY12_1),.clk(gclk));
	jdff dff_A_W3blJKaT6_0(.dout(w_dff_A_m5lxHlBy9_0),.din(w_dff_A_W3blJKaT6_0),.clk(gclk));
	jdff dff_A_m5lxHlBy9_0(.dout(w_dff_A_hDxQ0zxn9_0),.din(w_dff_A_m5lxHlBy9_0),.clk(gclk));
	jdff dff_A_hDxQ0zxn9_0(.dout(w_dff_A_Hlx88qOv2_0),.din(w_dff_A_hDxQ0zxn9_0),.clk(gclk));
	jdff dff_A_Hlx88qOv2_0(.dout(w_dff_A_SRZmYHN44_0),.din(w_dff_A_Hlx88qOv2_0),.clk(gclk));
	jdff dff_A_SRZmYHN44_0(.dout(w_dff_A_j8WvfXCf3_0),.din(w_dff_A_SRZmYHN44_0),.clk(gclk));
	jdff dff_A_j8WvfXCf3_0(.dout(w_dff_A_hGPvJOyA4_0),.din(w_dff_A_j8WvfXCf3_0),.clk(gclk));
	jdff dff_A_hGPvJOyA4_0(.dout(w_dff_A_1CGvhTYl6_0),.din(w_dff_A_hGPvJOyA4_0),.clk(gclk));
	jdff dff_A_1CGvhTYl6_0(.dout(w_dff_A_y4T2JSsi1_0),.din(w_dff_A_1CGvhTYl6_0),.clk(gclk));
	jdff dff_A_y4T2JSsi1_0(.dout(w_dff_A_ghNw8vfW5_0),.din(w_dff_A_y4T2JSsi1_0),.clk(gclk));
	jdff dff_A_ghNw8vfW5_0(.dout(w_dff_A_lQLqOei06_0),.din(w_dff_A_ghNw8vfW5_0),.clk(gclk));
	jdff dff_A_lQLqOei06_0(.dout(w_dff_A_3un9PmG75_0),.din(w_dff_A_lQLqOei06_0),.clk(gclk));
	jdff dff_A_3un9PmG75_0(.dout(w_dff_A_U8ZpNnbz5_0),.din(w_dff_A_3un9PmG75_0),.clk(gclk));
	jdff dff_A_U8ZpNnbz5_0(.dout(w_dff_A_CQI7aj3O9_0),.din(w_dff_A_U8ZpNnbz5_0),.clk(gclk));
	jdff dff_A_CQI7aj3O9_0(.dout(w_dff_A_PymAOf9O4_0),.din(w_dff_A_CQI7aj3O9_0),.clk(gclk));
	jdff dff_A_PymAOf9O4_0(.dout(w_dff_A_WFBKwnf95_0),.din(w_dff_A_PymAOf9O4_0),.clk(gclk));
	jdff dff_A_WFBKwnf95_0(.dout(w_dff_A_bUgXr9FK0_0),.din(w_dff_A_WFBKwnf95_0),.clk(gclk));
	jdff dff_A_bUgXr9FK0_0(.dout(w_dff_A_5ga8yakY1_0),.din(w_dff_A_bUgXr9FK0_0),.clk(gclk));
	jdff dff_A_5ga8yakY1_0(.dout(w_dff_A_jyezGBJM0_0),.din(w_dff_A_5ga8yakY1_0),.clk(gclk));
	jdff dff_A_jyezGBJM0_0(.dout(w_dff_A_ADE6YPIK2_0),.din(w_dff_A_jyezGBJM0_0),.clk(gclk));
	jdff dff_A_ADE6YPIK2_0(.dout(w_dff_A_ZMSHaKc78_0),.din(w_dff_A_ADE6YPIK2_0),.clk(gclk));
	jdff dff_A_ZMSHaKc78_0(.dout(w_dff_A_StMOIgqG7_0),.din(w_dff_A_ZMSHaKc78_0),.clk(gclk));
	jdff dff_A_StMOIgqG7_0(.dout(w_dff_A_VVPO2BMh9_0),.din(w_dff_A_StMOIgqG7_0),.clk(gclk));
	jdff dff_A_VVPO2BMh9_0(.dout(w_dff_A_oe8Go6Nb7_0),.din(w_dff_A_VVPO2BMh9_0),.clk(gclk));
	jdff dff_A_oe8Go6Nb7_0(.dout(G601),.din(w_dff_A_oe8Go6Nb7_0),.clk(gclk));
	jdff dff_A_5UiApBuf0_1(.dout(w_dff_A_ZOfNn9lZ0_0),.din(w_dff_A_5UiApBuf0_1),.clk(gclk));
	jdff dff_A_ZOfNn9lZ0_0(.dout(w_dff_A_pCIAjKVy3_0),.din(w_dff_A_ZOfNn9lZ0_0),.clk(gclk));
	jdff dff_A_pCIAjKVy3_0(.dout(w_dff_A_lfRHEVvT8_0),.din(w_dff_A_pCIAjKVy3_0),.clk(gclk));
	jdff dff_A_lfRHEVvT8_0(.dout(w_dff_A_CCsFULqC1_0),.din(w_dff_A_lfRHEVvT8_0),.clk(gclk));
	jdff dff_A_CCsFULqC1_0(.dout(w_dff_A_q26Ia2Vz8_0),.din(w_dff_A_CCsFULqC1_0),.clk(gclk));
	jdff dff_A_q26Ia2Vz8_0(.dout(w_dff_A_txdgd2aV0_0),.din(w_dff_A_q26Ia2Vz8_0),.clk(gclk));
	jdff dff_A_txdgd2aV0_0(.dout(w_dff_A_Tqyn0PGs2_0),.din(w_dff_A_txdgd2aV0_0),.clk(gclk));
	jdff dff_A_Tqyn0PGs2_0(.dout(w_dff_A_PupEY9tU4_0),.din(w_dff_A_Tqyn0PGs2_0),.clk(gclk));
	jdff dff_A_PupEY9tU4_0(.dout(w_dff_A_GulXQyOr1_0),.din(w_dff_A_PupEY9tU4_0),.clk(gclk));
	jdff dff_A_GulXQyOr1_0(.dout(w_dff_A_VwJ7xpip8_0),.din(w_dff_A_GulXQyOr1_0),.clk(gclk));
	jdff dff_A_VwJ7xpip8_0(.dout(w_dff_A_JiNepxSR2_0),.din(w_dff_A_VwJ7xpip8_0),.clk(gclk));
	jdff dff_A_JiNepxSR2_0(.dout(w_dff_A_fdfoUjCQ8_0),.din(w_dff_A_JiNepxSR2_0),.clk(gclk));
	jdff dff_A_fdfoUjCQ8_0(.dout(w_dff_A_evjQ1GOQ6_0),.din(w_dff_A_fdfoUjCQ8_0),.clk(gclk));
	jdff dff_A_evjQ1GOQ6_0(.dout(w_dff_A_Ai2LZgHB2_0),.din(w_dff_A_evjQ1GOQ6_0),.clk(gclk));
	jdff dff_A_Ai2LZgHB2_0(.dout(w_dff_A_qkThCd3n6_0),.din(w_dff_A_Ai2LZgHB2_0),.clk(gclk));
	jdff dff_A_qkThCd3n6_0(.dout(w_dff_A_wP7OkQIs7_0),.din(w_dff_A_qkThCd3n6_0),.clk(gclk));
	jdff dff_A_wP7OkQIs7_0(.dout(w_dff_A_0gh7OFPG4_0),.din(w_dff_A_wP7OkQIs7_0),.clk(gclk));
	jdff dff_A_0gh7OFPG4_0(.dout(w_dff_A_Bc87HXuD6_0),.din(w_dff_A_0gh7OFPG4_0),.clk(gclk));
	jdff dff_A_Bc87HXuD6_0(.dout(w_dff_A_IXJSGref9_0),.din(w_dff_A_Bc87HXuD6_0),.clk(gclk));
	jdff dff_A_IXJSGref9_0(.dout(w_dff_A_3RJ4Z2zp8_0),.din(w_dff_A_IXJSGref9_0),.clk(gclk));
	jdff dff_A_3RJ4Z2zp8_0(.dout(w_dff_A_nZsYqJsJ8_0),.din(w_dff_A_3RJ4Z2zp8_0),.clk(gclk));
	jdff dff_A_nZsYqJsJ8_0(.dout(w_dff_A_jmvhyzkZ3_0),.din(w_dff_A_nZsYqJsJ8_0),.clk(gclk));
	jdff dff_A_jmvhyzkZ3_0(.dout(w_dff_A_TZvXZ9uQ0_0),.din(w_dff_A_jmvhyzkZ3_0),.clk(gclk));
	jdff dff_A_TZvXZ9uQ0_0(.dout(w_dff_A_uHLArAq26_0),.din(w_dff_A_TZvXZ9uQ0_0),.clk(gclk));
	jdff dff_A_uHLArAq26_0(.dout(G602),.din(w_dff_A_uHLArAq26_0),.clk(gclk));
	jdff dff_A_lAjJ6ntN2_1(.dout(w_dff_A_gX4l8LdO0_0),.din(w_dff_A_lAjJ6ntN2_1),.clk(gclk));
	jdff dff_A_gX4l8LdO0_0(.dout(w_dff_A_Ez6ANdeV7_0),.din(w_dff_A_gX4l8LdO0_0),.clk(gclk));
	jdff dff_A_Ez6ANdeV7_0(.dout(w_dff_A_0KZsZlnI4_0),.din(w_dff_A_Ez6ANdeV7_0),.clk(gclk));
	jdff dff_A_0KZsZlnI4_0(.dout(w_dff_A_dLJb00FY5_0),.din(w_dff_A_0KZsZlnI4_0),.clk(gclk));
	jdff dff_A_dLJb00FY5_0(.dout(w_dff_A_UJcq1LMn1_0),.din(w_dff_A_dLJb00FY5_0),.clk(gclk));
	jdff dff_A_UJcq1LMn1_0(.dout(w_dff_A_lD83Iwof9_0),.din(w_dff_A_UJcq1LMn1_0),.clk(gclk));
	jdff dff_A_lD83Iwof9_0(.dout(w_dff_A_Nx1kym4p3_0),.din(w_dff_A_lD83Iwof9_0),.clk(gclk));
	jdff dff_A_Nx1kym4p3_0(.dout(w_dff_A_QavivzIi6_0),.din(w_dff_A_Nx1kym4p3_0),.clk(gclk));
	jdff dff_A_QavivzIi6_0(.dout(w_dff_A_2t2VTaDi9_0),.din(w_dff_A_QavivzIi6_0),.clk(gclk));
	jdff dff_A_2t2VTaDi9_0(.dout(w_dff_A_CDtK9NDC3_0),.din(w_dff_A_2t2VTaDi9_0),.clk(gclk));
	jdff dff_A_CDtK9NDC3_0(.dout(w_dff_A_MJ9UoudK5_0),.din(w_dff_A_CDtK9NDC3_0),.clk(gclk));
	jdff dff_A_MJ9UoudK5_0(.dout(w_dff_A_btQjM91A6_0),.din(w_dff_A_MJ9UoudK5_0),.clk(gclk));
	jdff dff_A_btQjM91A6_0(.dout(w_dff_A_ncjZG1842_0),.din(w_dff_A_btQjM91A6_0),.clk(gclk));
	jdff dff_A_ncjZG1842_0(.dout(w_dff_A_BTtIqM3W0_0),.din(w_dff_A_ncjZG1842_0),.clk(gclk));
	jdff dff_A_BTtIqM3W0_0(.dout(w_dff_A_YPsrmVI95_0),.din(w_dff_A_BTtIqM3W0_0),.clk(gclk));
	jdff dff_A_YPsrmVI95_0(.dout(w_dff_A_efGUEy068_0),.din(w_dff_A_YPsrmVI95_0),.clk(gclk));
	jdff dff_A_efGUEy068_0(.dout(w_dff_A_XMI3Hs1t2_0),.din(w_dff_A_efGUEy068_0),.clk(gclk));
	jdff dff_A_XMI3Hs1t2_0(.dout(w_dff_A_43dXQUqv6_0),.din(w_dff_A_XMI3Hs1t2_0),.clk(gclk));
	jdff dff_A_43dXQUqv6_0(.dout(w_dff_A_c6UIM3pj6_0),.din(w_dff_A_43dXQUqv6_0),.clk(gclk));
	jdff dff_A_c6UIM3pj6_0(.dout(w_dff_A_t6VnbjB46_0),.din(w_dff_A_c6UIM3pj6_0),.clk(gclk));
	jdff dff_A_t6VnbjB46_0(.dout(w_dff_A_saPPbtAo1_0),.din(w_dff_A_t6VnbjB46_0),.clk(gclk));
	jdff dff_A_saPPbtAo1_0(.dout(w_dff_A_woxLorAt1_0),.din(w_dff_A_saPPbtAo1_0),.clk(gclk));
	jdff dff_A_woxLorAt1_0(.dout(w_dff_A_xC83BlN51_0),.din(w_dff_A_woxLorAt1_0),.clk(gclk));
	jdff dff_A_xC83BlN51_0(.dout(w_dff_A_yFnvOrBl4_0),.din(w_dff_A_xC83BlN51_0),.clk(gclk));
	jdff dff_A_yFnvOrBl4_0(.dout(G603),.din(w_dff_A_yFnvOrBl4_0),.clk(gclk));
	jdff dff_A_0HHr3PS48_1(.dout(w_dff_A_Qmt1iINc8_0),.din(w_dff_A_0HHr3PS48_1),.clk(gclk));
	jdff dff_A_Qmt1iINc8_0(.dout(w_dff_A_aEUtmnu55_0),.din(w_dff_A_Qmt1iINc8_0),.clk(gclk));
	jdff dff_A_aEUtmnu55_0(.dout(w_dff_A_68hFG8kh9_0),.din(w_dff_A_aEUtmnu55_0),.clk(gclk));
	jdff dff_A_68hFG8kh9_0(.dout(w_dff_A_i1ZtKfQ55_0),.din(w_dff_A_68hFG8kh9_0),.clk(gclk));
	jdff dff_A_i1ZtKfQ55_0(.dout(w_dff_A_02bHml4r6_0),.din(w_dff_A_i1ZtKfQ55_0),.clk(gclk));
	jdff dff_A_02bHml4r6_0(.dout(w_dff_A_1D89T5S51_0),.din(w_dff_A_02bHml4r6_0),.clk(gclk));
	jdff dff_A_1D89T5S51_0(.dout(w_dff_A_1eccpagy6_0),.din(w_dff_A_1D89T5S51_0),.clk(gclk));
	jdff dff_A_1eccpagy6_0(.dout(w_dff_A_69nOebat5_0),.din(w_dff_A_1eccpagy6_0),.clk(gclk));
	jdff dff_A_69nOebat5_0(.dout(w_dff_A_NrxZeAKF7_0),.din(w_dff_A_69nOebat5_0),.clk(gclk));
	jdff dff_A_NrxZeAKF7_0(.dout(w_dff_A_DhUKxEso9_0),.din(w_dff_A_NrxZeAKF7_0),.clk(gclk));
	jdff dff_A_DhUKxEso9_0(.dout(w_dff_A_IhPRGPGP1_0),.din(w_dff_A_DhUKxEso9_0),.clk(gclk));
	jdff dff_A_IhPRGPGP1_0(.dout(w_dff_A_RqErZqyq3_0),.din(w_dff_A_IhPRGPGP1_0),.clk(gclk));
	jdff dff_A_RqErZqyq3_0(.dout(w_dff_A_mvELn8jo3_0),.din(w_dff_A_RqErZqyq3_0),.clk(gclk));
	jdff dff_A_mvELn8jo3_0(.dout(w_dff_A_XLzwTO640_0),.din(w_dff_A_mvELn8jo3_0),.clk(gclk));
	jdff dff_A_XLzwTO640_0(.dout(w_dff_A_WbG5VX9j6_0),.din(w_dff_A_XLzwTO640_0),.clk(gclk));
	jdff dff_A_WbG5VX9j6_0(.dout(w_dff_A_PcQC7G1V9_0),.din(w_dff_A_WbG5VX9j6_0),.clk(gclk));
	jdff dff_A_PcQC7G1V9_0(.dout(w_dff_A_yXkrA4Gj0_0),.din(w_dff_A_PcQC7G1V9_0),.clk(gclk));
	jdff dff_A_yXkrA4Gj0_0(.dout(w_dff_A_lg24CHzt4_0),.din(w_dff_A_yXkrA4Gj0_0),.clk(gclk));
	jdff dff_A_lg24CHzt4_0(.dout(w_dff_A_U4yiVyUN6_0),.din(w_dff_A_lg24CHzt4_0),.clk(gclk));
	jdff dff_A_U4yiVyUN6_0(.dout(w_dff_A_IuxKDhvs7_0),.din(w_dff_A_U4yiVyUN6_0),.clk(gclk));
	jdff dff_A_IuxKDhvs7_0(.dout(w_dff_A_uJSbDNmw2_0),.din(w_dff_A_IuxKDhvs7_0),.clk(gclk));
	jdff dff_A_uJSbDNmw2_0(.dout(w_dff_A_9D16R5mB7_0),.din(w_dff_A_uJSbDNmw2_0),.clk(gclk));
	jdff dff_A_9D16R5mB7_0(.dout(w_dff_A_nqZkEy4U6_0),.din(w_dff_A_9D16R5mB7_0),.clk(gclk));
	jdff dff_A_nqZkEy4U6_0(.dout(w_dff_A_ALW4vH0j8_0),.din(w_dff_A_nqZkEy4U6_0),.clk(gclk));
	jdff dff_A_ALW4vH0j8_0(.dout(G604),.din(w_dff_A_ALW4vH0j8_0),.clk(gclk));
	jdff dff_A_pVw4klAf8_1(.dout(w_dff_A_QLZW3LF36_0),.din(w_dff_A_pVw4klAf8_1),.clk(gclk));
	jdff dff_A_QLZW3LF36_0(.dout(w_dff_A_U6fvBceE8_0),.din(w_dff_A_QLZW3LF36_0),.clk(gclk));
	jdff dff_A_U6fvBceE8_0(.dout(w_dff_A_j2UNdXJB2_0),.din(w_dff_A_U6fvBceE8_0),.clk(gclk));
	jdff dff_A_j2UNdXJB2_0(.dout(w_dff_A_mhqfB2Nq4_0),.din(w_dff_A_j2UNdXJB2_0),.clk(gclk));
	jdff dff_A_mhqfB2Nq4_0(.dout(w_dff_A_lvme9Jct0_0),.din(w_dff_A_mhqfB2Nq4_0),.clk(gclk));
	jdff dff_A_lvme9Jct0_0(.dout(w_dff_A_jJFicvkV8_0),.din(w_dff_A_lvme9Jct0_0),.clk(gclk));
	jdff dff_A_jJFicvkV8_0(.dout(w_dff_A_6YMLwFrZ2_0),.din(w_dff_A_jJFicvkV8_0),.clk(gclk));
	jdff dff_A_6YMLwFrZ2_0(.dout(w_dff_A_ja7oAzQ41_0),.din(w_dff_A_6YMLwFrZ2_0),.clk(gclk));
	jdff dff_A_ja7oAzQ41_0(.dout(w_dff_A_nGvgUjE06_0),.din(w_dff_A_ja7oAzQ41_0),.clk(gclk));
	jdff dff_A_nGvgUjE06_0(.dout(w_dff_A_24EAdmNA6_0),.din(w_dff_A_nGvgUjE06_0),.clk(gclk));
	jdff dff_A_24EAdmNA6_0(.dout(w_dff_A_GZdqD08q0_0),.din(w_dff_A_24EAdmNA6_0),.clk(gclk));
	jdff dff_A_GZdqD08q0_0(.dout(w_dff_A_4VY4z9Pt4_0),.din(w_dff_A_GZdqD08q0_0),.clk(gclk));
	jdff dff_A_4VY4z9Pt4_0(.dout(w_dff_A_il4hTyVm3_0),.din(w_dff_A_4VY4z9Pt4_0),.clk(gclk));
	jdff dff_A_il4hTyVm3_0(.dout(w_dff_A_ZEhDEe0d7_0),.din(w_dff_A_il4hTyVm3_0),.clk(gclk));
	jdff dff_A_ZEhDEe0d7_0(.dout(w_dff_A_RST6M91K4_0),.din(w_dff_A_ZEhDEe0d7_0),.clk(gclk));
	jdff dff_A_RST6M91K4_0(.dout(w_dff_A_NxDDcVaf2_0),.din(w_dff_A_RST6M91K4_0),.clk(gclk));
	jdff dff_A_NxDDcVaf2_0(.dout(w_dff_A_dvmq6JXW8_0),.din(w_dff_A_NxDDcVaf2_0),.clk(gclk));
	jdff dff_A_dvmq6JXW8_0(.dout(w_dff_A_NQkEYQCw9_0),.din(w_dff_A_dvmq6JXW8_0),.clk(gclk));
	jdff dff_A_NQkEYQCw9_0(.dout(w_dff_A_BKhPLSCs0_0),.din(w_dff_A_NQkEYQCw9_0),.clk(gclk));
	jdff dff_A_BKhPLSCs0_0(.dout(w_dff_A_JPzGiUwV2_0),.din(w_dff_A_BKhPLSCs0_0),.clk(gclk));
	jdff dff_A_JPzGiUwV2_0(.dout(w_dff_A_l2wvO4NR9_0),.din(w_dff_A_JPzGiUwV2_0),.clk(gclk));
	jdff dff_A_l2wvO4NR9_0(.dout(w_dff_A_W2E9JpJS4_0),.din(w_dff_A_l2wvO4NR9_0),.clk(gclk));
	jdff dff_A_W2E9JpJS4_0(.dout(w_dff_A_YI2X50pv5_0),.din(w_dff_A_W2E9JpJS4_0),.clk(gclk));
	jdff dff_A_YI2X50pv5_0(.dout(w_dff_A_XqTn1v4h0_0),.din(w_dff_A_YI2X50pv5_0),.clk(gclk));
	jdff dff_A_XqTn1v4h0_0(.dout(G611),.din(w_dff_A_XqTn1v4h0_0),.clk(gclk));
	jdff dff_A_Kl1VYOge1_1(.dout(w_dff_A_B3EwKRTa9_0),.din(w_dff_A_Kl1VYOge1_1),.clk(gclk));
	jdff dff_A_B3EwKRTa9_0(.dout(w_dff_A_rbVVryLn6_0),.din(w_dff_A_B3EwKRTa9_0),.clk(gclk));
	jdff dff_A_rbVVryLn6_0(.dout(w_dff_A_c6k24Z1B1_0),.din(w_dff_A_rbVVryLn6_0),.clk(gclk));
	jdff dff_A_c6k24Z1B1_0(.dout(w_dff_A_2SynLc0q1_0),.din(w_dff_A_c6k24Z1B1_0),.clk(gclk));
	jdff dff_A_2SynLc0q1_0(.dout(w_dff_A_O3rLhcNa3_0),.din(w_dff_A_2SynLc0q1_0),.clk(gclk));
	jdff dff_A_O3rLhcNa3_0(.dout(w_dff_A_YFCZmZn02_0),.din(w_dff_A_O3rLhcNa3_0),.clk(gclk));
	jdff dff_A_YFCZmZn02_0(.dout(w_dff_A_DE6c4i8X6_0),.din(w_dff_A_YFCZmZn02_0),.clk(gclk));
	jdff dff_A_DE6c4i8X6_0(.dout(w_dff_A_NeIydeCE1_0),.din(w_dff_A_DE6c4i8X6_0),.clk(gclk));
	jdff dff_A_NeIydeCE1_0(.dout(w_dff_A_2Gutarxx1_0),.din(w_dff_A_NeIydeCE1_0),.clk(gclk));
	jdff dff_A_2Gutarxx1_0(.dout(w_dff_A_NuPQ2fAM5_0),.din(w_dff_A_2Gutarxx1_0),.clk(gclk));
	jdff dff_A_NuPQ2fAM5_0(.dout(w_dff_A_GwN5urio6_0),.din(w_dff_A_NuPQ2fAM5_0),.clk(gclk));
	jdff dff_A_GwN5urio6_0(.dout(w_dff_A_k0m57NFn4_0),.din(w_dff_A_GwN5urio6_0),.clk(gclk));
	jdff dff_A_k0m57NFn4_0(.dout(w_dff_A_MRZmuARF4_0),.din(w_dff_A_k0m57NFn4_0),.clk(gclk));
	jdff dff_A_MRZmuARF4_0(.dout(w_dff_A_veRZFaGf5_0),.din(w_dff_A_MRZmuARF4_0),.clk(gclk));
	jdff dff_A_veRZFaGf5_0(.dout(w_dff_A_EXIBH7FF2_0),.din(w_dff_A_veRZFaGf5_0),.clk(gclk));
	jdff dff_A_EXIBH7FF2_0(.dout(w_dff_A_AtIWkV7A8_0),.din(w_dff_A_EXIBH7FF2_0),.clk(gclk));
	jdff dff_A_AtIWkV7A8_0(.dout(w_dff_A_TFfMWMZO1_0),.din(w_dff_A_AtIWkV7A8_0),.clk(gclk));
	jdff dff_A_TFfMWMZO1_0(.dout(w_dff_A_iLXbjr3R9_0),.din(w_dff_A_TFfMWMZO1_0),.clk(gclk));
	jdff dff_A_iLXbjr3R9_0(.dout(w_dff_A_d4aptmOa9_0),.din(w_dff_A_iLXbjr3R9_0),.clk(gclk));
	jdff dff_A_d4aptmOa9_0(.dout(w_dff_A_q2MZOYAs3_0),.din(w_dff_A_d4aptmOa9_0),.clk(gclk));
	jdff dff_A_q2MZOYAs3_0(.dout(w_dff_A_KMZPdXSE5_0),.din(w_dff_A_q2MZOYAs3_0),.clk(gclk));
	jdff dff_A_KMZPdXSE5_0(.dout(w_dff_A_BbSM9Wij0_0),.din(w_dff_A_KMZPdXSE5_0),.clk(gclk));
	jdff dff_A_BbSM9Wij0_0(.dout(w_dff_A_hlhQvUvX2_0),.din(w_dff_A_BbSM9Wij0_0),.clk(gclk));
	jdff dff_A_hlhQvUvX2_0(.dout(w_dff_A_6NRR88zZ4_0),.din(w_dff_A_hlhQvUvX2_0),.clk(gclk));
	jdff dff_A_6NRR88zZ4_0(.dout(G612),.din(w_dff_A_6NRR88zZ4_0),.clk(gclk));
	jdff dff_A_xWfJIjhY9_2(.dout(w_dff_A_W4QEECt23_0),.din(w_dff_A_xWfJIjhY9_2),.clk(gclk));
	jdff dff_A_W4QEECt23_0(.dout(w_dff_A_MXJCNFNP1_0),.din(w_dff_A_W4QEECt23_0),.clk(gclk));
	jdff dff_A_MXJCNFNP1_0(.dout(w_dff_A_cSP4Twnl9_0),.din(w_dff_A_MXJCNFNP1_0),.clk(gclk));
	jdff dff_A_cSP4Twnl9_0(.dout(w_dff_A_iXMe5Czr1_0),.din(w_dff_A_cSP4Twnl9_0),.clk(gclk));
	jdff dff_A_iXMe5Czr1_0(.dout(w_dff_A_xFIVFouJ1_0),.din(w_dff_A_iXMe5Czr1_0),.clk(gclk));
	jdff dff_A_xFIVFouJ1_0(.dout(w_dff_A_0gMiaVB54_0),.din(w_dff_A_xFIVFouJ1_0),.clk(gclk));
	jdff dff_A_0gMiaVB54_0(.dout(w_dff_A_9jo7rlqd1_0),.din(w_dff_A_0gMiaVB54_0),.clk(gclk));
	jdff dff_A_9jo7rlqd1_0(.dout(w_dff_A_3JCQ8Gq22_0),.din(w_dff_A_9jo7rlqd1_0),.clk(gclk));
	jdff dff_A_3JCQ8Gq22_0(.dout(w_dff_A_Ax7jbXJF4_0),.din(w_dff_A_3JCQ8Gq22_0),.clk(gclk));
	jdff dff_A_Ax7jbXJF4_0(.dout(w_dff_A_nFmYb7tG1_0),.din(w_dff_A_Ax7jbXJF4_0),.clk(gclk));
	jdff dff_A_nFmYb7tG1_0(.dout(w_dff_A_6VGXosrO9_0),.din(w_dff_A_nFmYb7tG1_0),.clk(gclk));
	jdff dff_A_6VGXosrO9_0(.dout(w_dff_A_R0wUTnBv8_0),.din(w_dff_A_6VGXosrO9_0),.clk(gclk));
	jdff dff_A_R0wUTnBv8_0(.dout(w_dff_A_qw6D6rlu2_0),.din(w_dff_A_R0wUTnBv8_0),.clk(gclk));
	jdff dff_A_qw6D6rlu2_0(.dout(w_dff_A_OioMYsVH6_0),.din(w_dff_A_qw6D6rlu2_0),.clk(gclk));
	jdff dff_A_OioMYsVH6_0(.dout(w_dff_A_Pfcmgsu95_0),.din(w_dff_A_OioMYsVH6_0),.clk(gclk));
	jdff dff_A_Pfcmgsu95_0(.dout(w_dff_A_i8mtKWq51_0),.din(w_dff_A_Pfcmgsu95_0),.clk(gclk));
	jdff dff_A_i8mtKWq51_0(.dout(w_dff_A_IsSgKvSD1_0),.din(w_dff_A_i8mtKWq51_0),.clk(gclk));
	jdff dff_A_IsSgKvSD1_0(.dout(w_dff_A_uzhGcz4w8_0),.din(w_dff_A_IsSgKvSD1_0),.clk(gclk));
	jdff dff_A_uzhGcz4w8_0(.dout(w_dff_A_HsMeHz2e6_0),.din(w_dff_A_uzhGcz4w8_0),.clk(gclk));
	jdff dff_A_HsMeHz2e6_0(.dout(w_dff_A_n5iaUi1I4_0),.din(w_dff_A_HsMeHz2e6_0),.clk(gclk));
	jdff dff_A_n5iaUi1I4_0(.dout(w_dff_A_TXXm7fNr1_0),.din(w_dff_A_n5iaUi1I4_0),.clk(gclk));
	jdff dff_A_TXXm7fNr1_0(.dout(w_dff_A_r6nBd33b4_0),.din(w_dff_A_TXXm7fNr1_0),.clk(gclk));
	jdff dff_A_r6nBd33b4_0(.dout(w_dff_A_7eHj7Vmb0_0),.din(w_dff_A_r6nBd33b4_0),.clk(gclk));
	jdff dff_A_7eHj7Vmb0_0(.dout(w_dff_A_aMOluZcQ8_0),.din(w_dff_A_7eHj7Vmb0_0),.clk(gclk));
	jdff dff_A_aMOluZcQ8_0(.dout(G810),.din(w_dff_A_aMOluZcQ8_0),.clk(gclk));
	jdff dff_A_DKH03zRr9_1(.dout(w_dff_A_V9Dl4hlm9_0),.din(w_dff_A_DKH03zRr9_1),.clk(gclk));
	jdff dff_A_V9Dl4hlm9_0(.dout(w_dff_A_ZevjiADK7_0),.din(w_dff_A_V9Dl4hlm9_0),.clk(gclk));
	jdff dff_A_ZevjiADK7_0(.dout(w_dff_A_YH5oIzoM3_0),.din(w_dff_A_ZevjiADK7_0),.clk(gclk));
	jdff dff_A_YH5oIzoM3_0(.dout(w_dff_A_TYuXSnAM2_0),.din(w_dff_A_YH5oIzoM3_0),.clk(gclk));
	jdff dff_A_TYuXSnAM2_0(.dout(w_dff_A_ubolZQDz4_0),.din(w_dff_A_TYuXSnAM2_0),.clk(gclk));
	jdff dff_A_ubolZQDz4_0(.dout(w_dff_A_J1c3ZeLx1_0),.din(w_dff_A_ubolZQDz4_0),.clk(gclk));
	jdff dff_A_J1c3ZeLx1_0(.dout(w_dff_A_OCHDOgu56_0),.din(w_dff_A_J1c3ZeLx1_0),.clk(gclk));
	jdff dff_A_OCHDOgu56_0(.dout(w_dff_A_wU3Gi6uw6_0),.din(w_dff_A_OCHDOgu56_0),.clk(gclk));
	jdff dff_A_wU3Gi6uw6_0(.dout(w_dff_A_5z0GlFRk3_0),.din(w_dff_A_wU3Gi6uw6_0),.clk(gclk));
	jdff dff_A_5z0GlFRk3_0(.dout(w_dff_A_ISNGNLqq6_0),.din(w_dff_A_5z0GlFRk3_0),.clk(gclk));
	jdff dff_A_ISNGNLqq6_0(.dout(w_dff_A_itNXrn802_0),.din(w_dff_A_ISNGNLqq6_0),.clk(gclk));
	jdff dff_A_itNXrn802_0(.dout(w_dff_A_Cjtrg6io1_0),.din(w_dff_A_itNXrn802_0),.clk(gclk));
	jdff dff_A_Cjtrg6io1_0(.dout(w_dff_A_xtaWXGfw8_0),.din(w_dff_A_Cjtrg6io1_0),.clk(gclk));
	jdff dff_A_xtaWXGfw8_0(.dout(w_dff_A_SugRY9d51_0),.din(w_dff_A_xtaWXGfw8_0),.clk(gclk));
	jdff dff_A_SugRY9d51_0(.dout(w_dff_A_fXetze8D1_0),.din(w_dff_A_SugRY9d51_0),.clk(gclk));
	jdff dff_A_fXetze8D1_0(.dout(w_dff_A_PoTC19mg5_0),.din(w_dff_A_fXetze8D1_0),.clk(gclk));
	jdff dff_A_PoTC19mg5_0(.dout(w_dff_A_dOIkIvFI4_0),.din(w_dff_A_PoTC19mg5_0),.clk(gclk));
	jdff dff_A_dOIkIvFI4_0(.dout(w_dff_A_qYYjo8Di4_0),.din(w_dff_A_dOIkIvFI4_0),.clk(gclk));
	jdff dff_A_qYYjo8Di4_0(.dout(w_dff_A_50UqEfcW1_0),.din(w_dff_A_qYYjo8Di4_0),.clk(gclk));
	jdff dff_A_50UqEfcW1_0(.dout(w_dff_A_enR1XClG3_0),.din(w_dff_A_50UqEfcW1_0),.clk(gclk));
	jdff dff_A_enR1XClG3_0(.dout(w_dff_A_9S2mwn7J5_0),.din(w_dff_A_enR1XClG3_0),.clk(gclk));
	jdff dff_A_9S2mwn7J5_0(.dout(w_dff_A_RpaTGwKC1_0),.din(w_dff_A_9S2mwn7J5_0),.clk(gclk));
	jdff dff_A_RpaTGwKC1_0(.dout(w_dff_A_lo72eVtF8_0),.din(w_dff_A_RpaTGwKC1_0),.clk(gclk));
	jdff dff_A_lo72eVtF8_0(.dout(w_dff_A_0TcMbMkW1_0),.din(w_dff_A_lo72eVtF8_0),.clk(gclk));
	jdff dff_A_0TcMbMkW1_0(.dout(G848),.din(w_dff_A_0TcMbMkW1_0),.clk(gclk));
	jdff dff_A_C4E6I9xm8_1(.dout(w_dff_A_J3wecKfl8_0),.din(w_dff_A_C4E6I9xm8_1),.clk(gclk));
	jdff dff_A_J3wecKfl8_0(.dout(w_dff_A_PVdshIEX2_0),.din(w_dff_A_J3wecKfl8_0),.clk(gclk));
	jdff dff_A_PVdshIEX2_0(.dout(w_dff_A_9tqw22TR0_0),.din(w_dff_A_PVdshIEX2_0),.clk(gclk));
	jdff dff_A_9tqw22TR0_0(.dout(w_dff_A_o3O10GqH6_0),.din(w_dff_A_9tqw22TR0_0),.clk(gclk));
	jdff dff_A_o3O10GqH6_0(.dout(w_dff_A_VKsIspZl5_0),.din(w_dff_A_o3O10GqH6_0),.clk(gclk));
	jdff dff_A_VKsIspZl5_0(.dout(w_dff_A_w7nMf7iq6_0),.din(w_dff_A_VKsIspZl5_0),.clk(gclk));
	jdff dff_A_w7nMf7iq6_0(.dout(w_dff_A_gD03OdNp1_0),.din(w_dff_A_w7nMf7iq6_0),.clk(gclk));
	jdff dff_A_gD03OdNp1_0(.dout(w_dff_A_pWObaypn4_0),.din(w_dff_A_gD03OdNp1_0),.clk(gclk));
	jdff dff_A_pWObaypn4_0(.dout(w_dff_A_JhTP2HUO8_0),.din(w_dff_A_pWObaypn4_0),.clk(gclk));
	jdff dff_A_JhTP2HUO8_0(.dout(w_dff_A_vNHZzIe48_0),.din(w_dff_A_JhTP2HUO8_0),.clk(gclk));
	jdff dff_A_vNHZzIe48_0(.dout(w_dff_A_LcUEyZrV4_0),.din(w_dff_A_vNHZzIe48_0),.clk(gclk));
	jdff dff_A_LcUEyZrV4_0(.dout(w_dff_A_tb1jacsR7_0),.din(w_dff_A_LcUEyZrV4_0),.clk(gclk));
	jdff dff_A_tb1jacsR7_0(.dout(w_dff_A_KIy3WwXd8_0),.din(w_dff_A_tb1jacsR7_0),.clk(gclk));
	jdff dff_A_KIy3WwXd8_0(.dout(w_dff_A_K1ZQVDtw3_0),.din(w_dff_A_KIy3WwXd8_0),.clk(gclk));
	jdff dff_A_K1ZQVDtw3_0(.dout(w_dff_A_JprNTZPk2_0),.din(w_dff_A_K1ZQVDtw3_0),.clk(gclk));
	jdff dff_A_JprNTZPk2_0(.dout(w_dff_A_QObp4Vzv6_0),.din(w_dff_A_JprNTZPk2_0),.clk(gclk));
	jdff dff_A_QObp4Vzv6_0(.dout(w_dff_A_uFxb5Z0a8_0),.din(w_dff_A_QObp4Vzv6_0),.clk(gclk));
	jdff dff_A_uFxb5Z0a8_0(.dout(w_dff_A_mfr59jnh5_0),.din(w_dff_A_uFxb5Z0a8_0),.clk(gclk));
	jdff dff_A_mfr59jnh5_0(.dout(w_dff_A_hmAAue0G0_0),.din(w_dff_A_mfr59jnh5_0),.clk(gclk));
	jdff dff_A_hmAAue0G0_0(.dout(w_dff_A_KhmX7SqM9_0),.din(w_dff_A_hmAAue0G0_0),.clk(gclk));
	jdff dff_A_KhmX7SqM9_0(.dout(w_dff_A_82TbgnjM3_0),.din(w_dff_A_KhmX7SqM9_0),.clk(gclk));
	jdff dff_A_82TbgnjM3_0(.dout(w_dff_A_qur3YhbT2_0),.din(w_dff_A_82TbgnjM3_0),.clk(gclk));
	jdff dff_A_qur3YhbT2_0(.dout(w_dff_A_PgAh9jYo8_0),.din(w_dff_A_qur3YhbT2_0),.clk(gclk));
	jdff dff_A_PgAh9jYo8_0(.dout(w_dff_A_vJqoAf853_0),.din(w_dff_A_PgAh9jYo8_0),.clk(gclk));
	jdff dff_A_vJqoAf853_0(.dout(G849),.din(w_dff_A_vJqoAf853_0),.clk(gclk));
	jdff dff_A_IneqafsU3_1(.dout(w_dff_A_bdp2HV5j4_0),.din(w_dff_A_IneqafsU3_1),.clk(gclk));
	jdff dff_A_bdp2HV5j4_0(.dout(w_dff_A_ZMxhpMte3_0),.din(w_dff_A_bdp2HV5j4_0),.clk(gclk));
	jdff dff_A_ZMxhpMte3_0(.dout(w_dff_A_T24lEb8t1_0),.din(w_dff_A_ZMxhpMte3_0),.clk(gclk));
	jdff dff_A_T24lEb8t1_0(.dout(w_dff_A_zDmCoZu30_0),.din(w_dff_A_T24lEb8t1_0),.clk(gclk));
	jdff dff_A_zDmCoZu30_0(.dout(w_dff_A_woHPVkCV7_0),.din(w_dff_A_zDmCoZu30_0),.clk(gclk));
	jdff dff_A_woHPVkCV7_0(.dout(w_dff_A_s6T66enI5_0),.din(w_dff_A_woHPVkCV7_0),.clk(gclk));
	jdff dff_A_s6T66enI5_0(.dout(w_dff_A_60S9acg72_0),.din(w_dff_A_s6T66enI5_0),.clk(gclk));
	jdff dff_A_60S9acg72_0(.dout(w_dff_A_IsYTu06N0_0),.din(w_dff_A_60S9acg72_0),.clk(gclk));
	jdff dff_A_IsYTu06N0_0(.dout(w_dff_A_CDoPbfqB5_0),.din(w_dff_A_IsYTu06N0_0),.clk(gclk));
	jdff dff_A_CDoPbfqB5_0(.dout(w_dff_A_wB8aa1u45_0),.din(w_dff_A_CDoPbfqB5_0),.clk(gclk));
	jdff dff_A_wB8aa1u45_0(.dout(w_dff_A_SpKjj8Rh2_0),.din(w_dff_A_wB8aa1u45_0),.clk(gclk));
	jdff dff_A_SpKjj8Rh2_0(.dout(w_dff_A_FiJF7Unv8_0),.din(w_dff_A_SpKjj8Rh2_0),.clk(gclk));
	jdff dff_A_FiJF7Unv8_0(.dout(w_dff_A_PUkP4kX68_0),.din(w_dff_A_FiJF7Unv8_0),.clk(gclk));
	jdff dff_A_PUkP4kX68_0(.dout(w_dff_A_HpCYed7l8_0),.din(w_dff_A_PUkP4kX68_0),.clk(gclk));
	jdff dff_A_HpCYed7l8_0(.dout(w_dff_A_HP3KpLfy3_0),.din(w_dff_A_HpCYed7l8_0),.clk(gclk));
	jdff dff_A_HP3KpLfy3_0(.dout(w_dff_A_utArNpwp5_0),.din(w_dff_A_HP3KpLfy3_0),.clk(gclk));
	jdff dff_A_utArNpwp5_0(.dout(w_dff_A_nn2F6oWB8_0),.din(w_dff_A_utArNpwp5_0),.clk(gclk));
	jdff dff_A_nn2F6oWB8_0(.dout(w_dff_A_wFixckNx2_0),.din(w_dff_A_nn2F6oWB8_0),.clk(gclk));
	jdff dff_A_wFixckNx2_0(.dout(w_dff_A_DcnDZqoU9_0),.din(w_dff_A_wFixckNx2_0),.clk(gclk));
	jdff dff_A_DcnDZqoU9_0(.dout(w_dff_A_fnWcAW433_0),.din(w_dff_A_DcnDZqoU9_0),.clk(gclk));
	jdff dff_A_fnWcAW433_0(.dout(w_dff_A_j6BIrdjI5_0),.din(w_dff_A_fnWcAW433_0),.clk(gclk));
	jdff dff_A_j6BIrdjI5_0(.dout(w_dff_A_zF1ysYqI0_0),.din(w_dff_A_j6BIrdjI5_0),.clk(gclk));
	jdff dff_A_zF1ysYqI0_0(.dout(w_dff_A_JSZIW3jV1_0),.din(w_dff_A_zF1ysYqI0_0),.clk(gclk));
	jdff dff_A_JSZIW3jV1_0(.dout(w_dff_A_kfRy5ahu9_0),.din(w_dff_A_JSZIW3jV1_0),.clk(gclk));
	jdff dff_A_kfRy5ahu9_0(.dout(G850),.din(w_dff_A_kfRy5ahu9_0),.clk(gclk));
	jdff dff_A_1xSfMYMt0_1(.dout(w_dff_A_9LKRB3f68_0),.din(w_dff_A_1xSfMYMt0_1),.clk(gclk));
	jdff dff_A_9LKRB3f68_0(.dout(w_dff_A_gc0i5aTx3_0),.din(w_dff_A_9LKRB3f68_0),.clk(gclk));
	jdff dff_A_gc0i5aTx3_0(.dout(w_dff_A_ZnFsmU7S4_0),.din(w_dff_A_gc0i5aTx3_0),.clk(gclk));
	jdff dff_A_ZnFsmU7S4_0(.dout(w_dff_A_LXhdFnde2_0),.din(w_dff_A_ZnFsmU7S4_0),.clk(gclk));
	jdff dff_A_LXhdFnde2_0(.dout(w_dff_A_OK9feKSz0_0),.din(w_dff_A_LXhdFnde2_0),.clk(gclk));
	jdff dff_A_OK9feKSz0_0(.dout(w_dff_A_teOyDpbz2_0),.din(w_dff_A_OK9feKSz0_0),.clk(gclk));
	jdff dff_A_teOyDpbz2_0(.dout(w_dff_A_P1SAHPB60_0),.din(w_dff_A_teOyDpbz2_0),.clk(gclk));
	jdff dff_A_P1SAHPB60_0(.dout(w_dff_A_agHq9Vxe8_0),.din(w_dff_A_P1SAHPB60_0),.clk(gclk));
	jdff dff_A_agHq9Vxe8_0(.dout(w_dff_A_W6mCaI3z2_0),.din(w_dff_A_agHq9Vxe8_0),.clk(gclk));
	jdff dff_A_W6mCaI3z2_0(.dout(w_dff_A_8vAThO435_0),.din(w_dff_A_W6mCaI3z2_0),.clk(gclk));
	jdff dff_A_8vAThO435_0(.dout(w_dff_A_eP8CBvWY0_0),.din(w_dff_A_8vAThO435_0),.clk(gclk));
	jdff dff_A_eP8CBvWY0_0(.dout(w_dff_A_lJPviwf89_0),.din(w_dff_A_eP8CBvWY0_0),.clk(gclk));
	jdff dff_A_lJPviwf89_0(.dout(w_dff_A_KQClxOC20_0),.din(w_dff_A_lJPviwf89_0),.clk(gclk));
	jdff dff_A_KQClxOC20_0(.dout(w_dff_A_xYtiwiq53_0),.din(w_dff_A_KQClxOC20_0),.clk(gclk));
	jdff dff_A_xYtiwiq53_0(.dout(w_dff_A_jROIc4bY6_0),.din(w_dff_A_xYtiwiq53_0),.clk(gclk));
	jdff dff_A_jROIc4bY6_0(.dout(w_dff_A_V1qaUMme6_0),.din(w_dff_A_jROIc4bY6_0),.clk(gclk));
	jdff dff_A_V1qaUMme6_0(.dout(w_dff_A_jAtJSnBV4_0),.din(w_dff_A_V1qaUMme6_0),.clk(gclk));
	jdff dff_A_jAtJSnBV4_0(.dout(w_dff_A_Q4j7EZNm1_0),.din(w_dff_A_jAtJSnBV4_0),.clk(gclk));
	jdff dff_A_Q4j7EZNm1_0(.dout(w_dff_A_dGN7hzBT7_0),.din(w_dff_A_Q4j7EZNm1_0),.clk(gclk));
	jdff dff_A_dGN7hzBT7_0(.dout(w_dff_A_hR5xHatP1_0),.din(w_dff_A_dGN7hzBT7_0),.clk(gclk));
	jdff dff_A_hR5xHatP1_0(.dout(w_dff_A_FszJodIF2_0),.din(w_dff_A_hR5xHatP1_0),.clk(gclk));
	jdff dff_A_FszJodIF2_0(.dout(w_dff_A_mAvnTKmL2_0),.din(w_dff_A_FszJodIF2_0),.clk(gclk));
	jdff dff_A_mAvnTKmL2_0(.dout(w_dff_A_S6IQxkHY2_0),.din(w_dff_A_mAvnTKmL2_0),.clk(gclk));
	jdff dff_A_S6IQxkHY2_0(.dout(w_dff_A_aqqtuCRt9_0),.din(w_dff_A_S6IQxkHY2_0),.clk(gclk));
	jdff dff_A_aqqtuCRt9_0(.dout(G851),.din(w_dff_A_aqqtuCRt9_0),.clk(gclk));
	jdff dff_A_ZCfZqptZ2_2(.dout(w_dff_A_AkxK3PXr7_0),.din(w_dff_A_ZCfZqptZ2_2),.clk(gclk));
	jdff dff_A_AkxK3PXr7_0(.dout(w_dff_A_j94OQCS04_0),.din(w_dff_A_AkxK3PXr7_0),.clk(gclk));
	jdff dff_A_j94OQCS04_0(.dout(w_dff_A_cQBw3GLb0_0),.din(w_dff_A_j94OQCS04_0),.clk(gclk));
	jdff dff_A_cQBw3GLb0_0(.dout(w_dff_A_ysenTGml1_0),.din(w_dff_A_cQBw3GLb0_0),.clk(gclk));
	jdff dff_A_ysenTGml1_0(.dout(w_dff_A_AxYT9JZM0_0),.din(w_dff_A_ysenTGml1_0),.clk(gclk));
	jdff dff_A_AxYT9JZM0_0(.dout(w_dff_A_hKYqQDsu7_0),.din(w_dff_A_AxYT9JZM0_0),.clk(gclk));
	jdff dff_A_hKYqQDsu7_0(.dout(w_dff_A_1r1Xn5aR6_0),.din(w_dff_A_hKYqQDsu7_0),.clk(gclk));
	jdff dff_A_1r1Xn5aR6_0(.dout(w_dff_A_q78m1Ni15_0),.din(w_dff_A_1r1Xn5aR6_0),.clk(gclk));
	jdff dff_A_q78m1Ni15_0(.dout(w_dff_A_FOJ9xqi72_0),.din(w_dff_A_q78m1Ni15_0),.clk(gclk));
	jdff dff_A_FOJ9xqi72_0(.dout(w_dff_A_oWZFgUY55_0),.din(w_dff_A_FOJ9xqi72_0),.clk(gclk));
	jdff dff_A_oWZFgUY55_0(.dout(w_dff_A_Zct95VyD4_0),.din(w_dff_A_oWZFgUY55_0),.clk(gclk));
	jdff dff_A_Zct95VyD4_0(.dout(w_dff_A_Yl725GGn9_0),.din(w_dff_A_Zct95VyD4_0),.clk(gclk));
	jdff dff_A_Yl725GGn9_0(.dout(w_dff_A_4vRX5qte9_0),.din(w_dff_A_Yl725GGn9_0),.clk(gclk));
	jdff dff_A_4vRX5qte9_0(.dout(w_dff_A_TzdtOuMs7_0),.din(w_dff_A_4vRX5qte9_0),.clk(gclk));
	jdff dff_A_TzdtOuMs7_0(.dout(w_dff_A_ZsjCNNIt6_0),.din(w_dff_A_TzdtOuMs7_0),.clk(gclk));
	jdff dff_A_ZsjCNNIt6_0(.dout(w_dff_A_sNtzgHPm3_0),.din(w_dff_A_ZsjCNNIt6_0),.clk(gclk));
	jdff dff_A_sNtzgHPm3_0(.dout(w_dff_A_W3L6Sddn7_0),.din(w_dff_A_sNtzgHPm3_0),.clk(gclk));
	jdff dff_A_W3L6Sddn7_0(.dout(w_dff_A_UAHvOLWt6_0),.din(w_dff_A_W3L6Sddn7_0),.clk(gclk));
	jdff dff_A_UAHvOLWt6_0(.dout(w_dff_A_J7uiRwTk6_0),.din(w_dff_A_UAHvOLWt6_0),.clk(gclk));
	jdff dff_A_J7uiRwTk6_0(.dout(w_dff_A_l6pT0S5f5_0),.din(w_dff_A_J7uiRwTk6_0),.clk(gclk));
	jdff dff_A_l6pT0S5f5_0(.dout(w_dff_A_yXpblTTG0_0),.din(w_dff_A_l6pT0S5f5_0),.clk(gclk));
	jdff dff_A_yXpblTTG0_0(.dout(w_dff_A_uS9K5RRB1_0),.din(w_dff_A_yXpblTTG0_0),.clk(gclk));
	jdff dff_A_uS9K5RRB1_0(.dout(w_dff_A_Xtw3kVUu5_0),.din(w_dff_A_uS9K5RRB1_0),.clk(gclk));
	jdff dff_A_Xtw3kVUu5_0(.dout(w_dff_A_dlMMGcj04_0),.din(w_dff_A_Xtw3kVUu5_0),.clk(gclk));
	jdff dff_A_dlMMGcj04_0(.dout(G634),.din(w_dff_A_dlMMGcj04_0),.clk(gclk));
	jdff dff_A_85EWI87F1_2(.dout(w_dff_A_wUlp3ZHb7_0),.din(w_dff_A_85EWI87F1_2),.clk(gclk));
	jdff dff_A_wUlp3ZHb7_0(.dout(w_dff_A_CtFMHTU65_0),.din(w_dff_A_wUlp3ZHb7_0),.clk(gclk));
	jdff dff_A_CtFMHTU65_0(.dout(w_dff_A_VRHQM1D97_0),.din(w_dff_A_CtFMHTU65_0),.clk(gclk));
	jdff dff_A_VRHQM1D97_0(.dout(w_dff_A_vuJDotK36_0),.din(w_dff_A_VRHQM1D97_0),.clk(gclk));
	jdff dff_A_vuJDotK36_0(.dout(w_dff_A_smtJ0N6p1_0),.din(w_dff_A_vuJDotK36_0),.clk(gclk));
	jdff dff_A_smtJ0N6p1_0(.dout(w_dff_A_nVzTU1wv0_0),.din(w_dff_A_smtJ0N6p1_0),.clk(gclk));
	jdff dff_A_nVzTU1wv0_0(.dout(w_dff_A_vgYyKTxe5_0),.din(w_dff_A_nVzTU1wv0_0),.clk(gclk));
	jdff dff_A_vgYyKTxe5_0(.dout(w_dff_A_CbaKDPNt4_0),.din(w_dff_A_vgYyKTxe5_0),.clk(gclk));
	jdff dff_A_CbaKDPNt4_0(.dout(w_dff_A_NJXZjmGw5_0),.din(w_dff_A_CbaKDPNt4_0),.clk(gclk));
	jdff dff_A_NJXZjmGw5_0(.dout(w_dff_A_U8hkgIES8_0),.din(w_dff_A_NJXZjmGw5_0),.clk(gclk));
	jdff dff_A_U8hkgIES8_0(.dout(w_dff_A_aCh7I36M3_0),.din(w_dff_A_U8hkgIES8_0),.clk(gclk));
	jdff dff_A_aCh7I36M3_0(.dout(w_dff_A_gVs8XcDN0_0),.din(w_dff_A_aCh7I36M3_0),.clk(gclk));
	jdff dff_A_gVs8XcDN0_0(.dout(w_dff_A_zkZJzAKK1_0),.din(w_dff_A_gVs8XcDN0_0),.clk(gclk));
	jdff dff_A_zkZJzAKK1_0(.dout(w_dff_A_2EEfBfON7_0),.din(w_dff_A_zkZJzAKK1_0),.clk(gclk));
	jdff dff_A_2EEfBfON7_0(.dout(w_dff_A_m8vJpnEV2_0),.din(w_dff_A_2EEfBfON7_0),.clk(gclk));
	jdff dff_A_m8vJpnEV2_0(.dout(w_dff_A_uUKXjEl93_0),.din(w_dff_A_m8vJpnEV2_0),.clk(gclk));
	jdff dff_A_uUKXjEl93_0(.dout(w_dff_A_RAsSNRWz7_0),.din(w_dff_A_uUKXjEl93_0),.clk(gclk));
	jdff dff_A_RAsSNRWz7_0(.dout(w_dff_A_NTzsG20u9_0),.din(w_dff_A_RAsSNRWz7_0),.clk(gclk));
	jdff dff_A_NTzsG20u9_0(.dout(w_dff_A_H8wcQRyh4_0),.din(w_dff_A_NTzsG20u9_0),.clk(gclk));
	jdff dff_A_H8wcQRyh4_0(.dout(w_dff_A_L6kVtjQ69_0),.din(w_dff_A_H8wcQRyh4_0),.clk(gclk));
	jdff dff_A_L6kVtjQ69_0(.dout(w_dff_A_RRt0yPzE5_0),.din(w_dff_A_L6kVtjQ69_0),.clk(gclk));
	jdff dff_A_RRt0yPzE5_0(.dout(w_dff_A_7o8UcTC54_0),.din(w_dff_A_RRt0yPzE5_0),.clk(gclk));
	jdff dff_A_7o8UcTC54_0(.dout(w_dff_A_0ncU4kYV4_0),.din(w_dff_A_7o8UcTC54_0),.clk(gclk));
	jdff dff_A_0ncU4kYV4_0(.dout(G815),.din(w_dff_A_0ncU4kYV4_0),.clk(gclk));
	jdff dff_A_wbIT1XPG9_2(.dout(w_dff_A_vgwIbBju5_0),.din(w_dff_A_wbIT1XPG9_2),.clk(gclk));
	jdff dff_A_vgwIbBju5_0(.dout(w_dff_A_bkFvrZ5J3_0),.din(w_dff_A_vgwIbBju5_0),.clk(gclk));
	jdff dff_A_bkFvrZ5J3_0(.dout(w_dff_A_xRcw8JG86_0),.din(w_dff_A_bkFvrZ5J3_0),.clk(gclk));
	jdff dff_A_xRcw8JG86_0(.dout(w_dff_A_kbBSzTe02_0),.din(w_dff_A_xRcw8JG86_0),.clk(gclk));
	jdff dff_A_kbBSzTe02_0(.dout(w_dff_A_7bH0luB35_0),.din(w_dff_A_kbBSzTe02_0),.clk(gclk));
	jdff dff_A_7bH0luB35_0(.dout(w_dff_A_zHxniMfJ0_0),.din(w_dff_A_7bH0luB35_0),.clk(gclk));
	jdff dff_A_zHxniMfJ0_0(.dout(w_dff_A_GXJk6YgY3_0),.din(w_dff_A_zHxniMfJ0_0),.clk(gclk));
	jdff dff_A_GXJk6YgY3_0(.dout(w_dff_A_DklyxYxz6_0),.din(w_dff_A_GXJk6YgY3_0),.clk(gclk));
	jdff dff_A_DklyxYxz6_0(.dout(w_dff_A_5J3lHr7j0_0),.din(w_dff_A_DklyxYxz6_0),.clk(gclk));
	jdff dff_A_5J3lHr7j0_0(.dout(w_dff_A_gkAYmFWb4_0),.din(w_dff_A_5J3lHr7j0_0),.clk(gclk));
	jdff dff_A_gkAYmFWb4_0(.dout(w_dff_A_Z9izDOnl8_0),.din(w_dff_A_gkAYmFWb4_0),.clk(gclk));
	jdff dff_A_Z9izDOnl8_0(.dout(w_dff_A_2UoyOGkc1_0),.din(w_dff_A_Z9izDOnl8_0),.clk(gclk));
	jdff dff_A_2UoyOGkc1_0(.dout(w_dff_A_besySP5H1_0),.din(w_dff_A_2UoyOGkc1_0),.clk(gclk));
	jdff dff_A_besySP5H1_0(.dout(w_dff_A_T1cYBKAv7_0),.din(w_dff_A_besySP5H1_0),.clk(gclk));
	jdff dff_A_T1cYBKAv7_0(.dout(w_dff_A_DWjNw2ar2_0),.din(w_dff_A_T1cYBKAv7_0),.clk(gclk));
	jdff dff_A_DWjNw2ar2_0(.dout(w_dff_A_yiRhqAu64_0),.din(w_dff_A_DWjNw2ar2_0),.clk(gclk));
	jdff dff_A_yiRhqAu64_0(.dout(w_dff_A_3s9vnMc08_0),.din(w_dff_A_yiRhqAu64_0),.clk(gclk));
	jdff dff_A_3s9vnMc08_0(.dout(w_dff_A_1XzhlFWJ2_0),.din(w_dff_A_3s9vnMc08_0),.clk(gclk));
	jdff dff_A_1XzhlFWJ2_0(.dout(w_dff_A_wSKLq0gu0_0),.din(w_dff_A_1XzhlFWJ2_0),.clk(gclk));
	jdff dff_A_wSKLq0gu0_0(.dout(w_dff_A_BCZp0mBa3_0),.din(w_dff_A_wSKLq0gu0_0),.clk(gclk));
	jdff dff_A_BCZp0mBa3_0(.dout(w_dff_A_uApHQBbg7_0),.din(w_dff_A_BCZp0mBa3_0),.clk(gclk));
	jdff dff_A_uApHQBbg7_0(.dout(w_dff_A_es2KX2yR9_0),.din(w_dff_A_uApHQBbg7_0),.clk(gclk));
	jdff dff_A_es2KX2yR9_0(.dout(w_dff_A_frJMrqSo1_0),.din(w_dff_A_es2KX2yR9_0),.clk(gclk));
	jdff dff_A_frJMrqSo1_0(.dout(G845),.din(w_dff_A_frJMrqSo1_0),.clk(gclk));
	jdff dff_A_baaaIop22_1(.dout(w_dff_A_qHT3LPmz5_0),.din(w_dff_A_baaaIop22_1),.clk(gclk));
	jdff dff_A_qHT3LPmz5_0(.dout(w_dff_A_zMglTbSo5_0),.din(w_dff_A_qHT3LPmz5_0),.clk(gclk));
	jdff dff_A_zMglTbSo5_0(.dout(w_dff_A_h9dnR1xR0_0),.din(w_dff_A_zMglTbSo5_0),.clk(gclk));
	jdff dff_A_h9dnR1xR0_0(.dout(w_dff_A_Wb0DyuPT7_0),.din(w_dff_A_h9dnR1xR0_0),.clk(gclk));
	jdff dff_A_Wb0DyuPT7_0(.dout(w_dff_A_rn7xnLiI9_0),.din(w_dff_A_Wb0DyuPT7_0),.clk(gclk));
	jdff dff_A_rn7xnLiI9_0(.dout(w_dff_A_gpoeS98b4_0),.din(w_dff_A_rn7xnLiI9_0),.clk(gclk));
	jdff dff_A_gpoeS98b4_0(.dout(w_dff_A_cJHceGsL9_0),.din(w_dff_A_gpoeS98b4_0),.clk(gclk));
	jdff dff_A_cJHceGsL9_0(.dout(w_dff_A_u3soHglQ8_0),.din(w_dff_A_cJHceGsL9_0),.clk(gclk));
	jdff dff_A_u3soHglQ8_0(.dout(w_dff_A_XrlUDqrv8_0),.din(w_dff_A_u3soHglQ8_0),.clk(gclk));
	jdff dff_A_XrlUDqrv8_0(.dout(w_dff_A_3yjouAZG0_0),.din(w_dff_A_XrlUDqrv8_0),.clk(gclk));
	jdff dff_A_3yjouAZG0_0(.dout(w_dff_A_jwnGBlz66_0),.din(w_dff_A_3yjouAZG0_0),.clk(gclk));
	jdff dff_A_jwnGBlz66_0(.dout(w_dff_A_NqnhHSnG4_0),.din(w_dff_A_jwnGBlz66_0),.clk(gclk));
	jdff dff_A_NqnhHSnG4_0(.dout(w_dff_A_ZzH1PtJZ5_0),.din(w_dff_A_NqnhHSnG4_0),.clk(gclk));
	jdff dff_A_ZzH1PtJZ5_0(.dout(w_dff_A_x7LHgaJv8_0),.din(w_dff_A_ZzH1PtJZ5_0),.clk(gclk));
	jdff dff_A_x7LHgaJv8_0(.dout(w_dff_A_VZvGSK4Y3_0),.din(w_dff_A_x7LHgaJv8_0),.clk(gclk));
	jdff dff_A_VZvGSK4Y3_0(.dout(w_dff_A_TYHC74x96_0),.din(w_dff_A_VZvGSK4Y3_0),.clk(gclk));
	jdff dff_A_TYHC74x96_0(.dout(w_dff_A_23nFjEDI6_0),.din(w_dff_A_TYHC74x96_0),.clk(gclk));
	jdff dff_A_23nFjEDI6_0(.dout(w_dff_A_ET4TfNhs6_0),.din(w_dff_A_23nFjEDI6_0),.clk(gclk));
	jdff dff_A_ET4TfNhs6_0(.dout(w_dff_A_yMhm8xQV2_0),.din(w_dff_A_ET4TfNhs6_0),.clk(gclk));
	jdff dff_A_yMhm8xQV2_0(.dout(w_dff_A_Pco2ROqo6_0),.din(w_dff_A_yMhm8xQV2_0),.clk(gclk));
	jdff dff_A_Pco2ROqo6_0(.dout(w_dff_A_pv6D1KCd8_0),.din(w_dff_A_Pco2ROqo6_0),.clk(gclk));
	jdff dff_A_pv6D1KCd8_0(.dout(w_dff_A_WHxedDe84_0),.din(w_dff_A_pv6D1KCd8_0),.clk(gclk));
	jdff dff_A_WHxedDe84_0(.dout(w_dff_A_Q52y1VST8_0),.din(w_dff_A_WHxedDe84_0),.clk(gclk));
	jdff dff_A_Q52y1VST8_0(.dout(G847),.din(w_dff_A_Q52y1VST8_0),.clk(gclk));
	jdff dff_A_0NtsHe4k0_1(.dout(w_dff_A_z8SEhmuw8_0),.din(w_dff_A_0NtsHe4k0_1),.clk(gclk));
	jdff dff_A_z8SEhmuw8_0(.dout(w_dff_A_0JW3qpPK1_0),.din(w_dff_A_z8SEhmuw8_0),.clk(gclk));
	jdff dff_A_0JW3qpPK1_0(.dout(w_dff_A_uZQRpj9u4_0),.din(w_dff_A_0JW3qpPK1_0),.clk(gclk));
	jdff dff_A_uZQRpj9u4_0(.dout(w_dff_A_UOWIhbIO6_0),.din(w_dff_A_uZQRpj9u4_0),.clk(gclk));
	jdff dff_A_UOWIhbIO6_0(.dout(w_dff_A_fcI1VUiZ9_0),.din(w_dff_A_UOWIhbIO6_0),.clk(gclk));
	jdff dff_A_fcI1VUiZ9_0(.dout(w_dff_A_BWbThhkX9_0),.din(w_dff_A_fcI1VUiZ9_0),.clk(gclk));
	jdff dff_A_BWbThhkX9_0(.dout(w_dff_A_4qtfWl6m2_0),.din(w_dff_A_BWbThhkX9_0),.clk(gclk));
	jdff dff_A_4qtfWl6m2_0(.dout(w_dff_A_UIUiWn8S4_0),.din(w_dff_A_4qtfWl6m2_0),.clk(gclk));
	jdff dff_A_UIUiWn8S4_0(.dout(w_dff_A_fvWGtN4H3_0),.din(w_dff_A_UIUiWn8S4_0),.clk(gclk));
	jdff dff_A_fvWGtN4H3_0(.dout(w_dff_A_VgWcOzhL8_0),.din(w_dff_A_fvWGtN4H3_0),.clk(gclk));
	jdff dff_A_VgWcOzhL8_0(.dout(w_dff_A_8VCmIRiZ1_0),.din(w_dff_A_VgWcOzhL8_0),.clk(gclk));
	jdff dff_A_8VCmIRiZ1_0(.dout(w_dff_A_aiG5mRhr7_0),.din(w_dff_A_8VCmIRiZ1_0),.clk(gclk));
	jdff dff_A_aiG5mRhr7_0(.dout(w_dff_A_rnff7rdv9_0),.din(w_dff_A_aiG5mRhr7_0),.clk(gclk));
	jdff dff_A_rnff7rdv9_0(.dout(w_dff_A_C5fA222u1_0),.din(w_dff_A_rnff7rdv9_0),.clk(gclk));
	jdff dff_A_C5fA222u1_0(.dout(w_dff_A_in6rFIyp5_0),.din(w_dff_A_C5fA222u1_0),.clk(gclk));
	jdff dff_A_in6rFIyp5_0(.dout(w_dff_A_xHmOpUZn8_0),.din(w_dff_A_in6rFIyp5_0),.clk(gclk));
	jdff dff_A_xHmOpUZn8_0(.dout(w_dff_A_ZO8cscaM6_0),.din(w_dff_A_xHmOpUZn8_0),.clk(gclk));
	jdff dff_A_ZO8cscaM6_0(.dout(w_dff_A_N8nSplsF6_0),.din(w_dff_A_ZO8cscaM6_0),.clk(gclk));
	jdff dff_A_N8nSplsF6_0(.dout(w_dff_A_22FwJYlc0_0),.din(w_dff_A_N8nSplsF6_0),.clk(gclk));
	jdff dff_A_22FwJYlc0_0(.dout(w_dff_A_xbtWDrRh7_0),.din(w_dff_A_22FwJYlc0_0),.clk(gclk));
	jdff dff_A_xbtWDrRh7_0(.dout(w_dff_A_JzC9FgC18_0),.din(w_dff_A_xbtWDrRh7_0),.clk(gclk));
	jdff dff_A_JzC9FgC18_0(.dout(w_dff_A_DhTOD46w3_0),.din(w_dff_A_JzC9FgC18_0),.clk(gclk));
	jdff dff_A_DhTOD46w3_0(.dout(w_dff_A_0lLBpF6k3_0),.din(w_dff_A_DhTOD46w3_0),.clk(gclk));
	jdff dff_A_0lLBpF6k3_0(.dout(w_dff_A_910Pao2f1_0),.din(w_dff_A_0lLBpF6k3_0),.clk(gclk));
	jdff dff_A_910Pao2f1_0(.dout(G926),.din(w_dff_A_910Pao2f1_0),.clk(gclk));
	jdff dff_A_U6IqrDOA3_1(.dout(w_dff_A_JFuCtzja3_0),.din(w_dff_A_U6IqrDOA3_1),.clk(gclk));
	jdff dff_A_JFuCtzja3_0(.dout(w_dff_A_gBl0FTYb2_0),.din(w_dff_A_JFuCtzja3_0),.clk(gclk));
	jdff dff_A_gBl0FTYb2_0(.dout(w_dff_A_1U6gpGID3_0),.din(w_dff_A_gBl0FTYb2_0),.clk(gclk));
	jdff dff_A_1U6gpGID3_0(.dout(w_dff_A_tzfrMzca0_0),.din(w_dff_A_1U6gpGID3_0),.clk(gclk));
	jdff dff_A_tzfrMzca0_0(.dout(w_dff_A_7nS1bCmI1_0),.din(w_dff_A_tzfrMzca0_0),.clk(gclk));
	jdff dff_A_7nS1bCmI1_0(.dout(w_dff_A_TxHYNhcK3_0),.din(w_dff_A_7nS1bCmI1_0),.clk(gclk));
	jdff dff_A_TxHYNhcK3_0(.dout(w_dff_A_6joH87FZ8_0),.din(w_dff_A_TxHYNhcK3_0),.clk(gclk));
	jdff dff_A_6joH87FZ8_0(.dout(w_dff_A_Q1vsS2BU7_0),.din(w_dff_A_6joH87FZ8_0),.clk(gclk));
	jdff dff_A_Q1vsS2BU7_0(.dout(w_dff_A_1lOXF1qY7_0),.din(w_dff_A_Q1vsS2BU7_0),.clk(gclk));
	jdff dff_A_1lOXF1qY7_0(.dout(w_dff_A_QxvhYoBx7_0),.din(w_dff_A_1lOXF1qY7_0),.clk(gclk));
	jdff dff_A_QxvhYoBx7_0(.dout(w_dff_A_SLCOGf525_0),.din(w_dff_A_QxvhYoBx7_0),.clk(gclk));
	jdff dff_A_SLCOGf525_0(.dout(w_dff_A_4roXJf559_0),.din(w_dff_A_SLCOGf525_0),.clk(gclk));
	jdff dff_A_4roXJf559_0(.dout(w_dff_A_r1zjsBTd8_0),.din(w_dff_A_4roXJf559_0),.clk(gclk));
	jdff dff_A_r1zjsBTd8_0(.dout(w_dff_A_CLtav2Qi1_0),.din(w_dff_A_r1zjsBTd8_0),.clk(gclk));
	jdff dff_A_CLtav2Qi1_0(.dout(w_dff_A_WF6cgsK41_0),.din(w_dff_A_CLtav2Qi1_0),.clk(gclk));
	jdff dff_A_WF6cgsK41_0(.dout(w_dff_A_dJChjvxg0_0),.din(w_dff_A_WF6cgsK41_0),.clk(gclk));
	jdff dff_A_dJChjvxg0_0(.dout(w_dff_A_8ofXVN961_0),.din(w_dff_A_dJChjvxg0_0),.clk(gclk));
	jdff dff_A_8ofXVN961_0(.dout(w_dff_A_2WY6iaes8_0),.din(w_dff_A_8ofXVN961_0),.clk(gclk));
	jdff dff_A_2WY6iaes8_0(.dout(w_dff_A_PhvR06020_0),.din(w_dff_A_2WY6iaes8_0),.clk(gclk));
	jdff dff_A_PhvR06020_0(.dout(w_dff_A_gZnyTgn10_0),.din(w_dff_A_PhvR06020_0),.clk(gclk));
	jdff dff_A_gZnyTgn10_0(.dout(w_dff_A_OovXxVAL4_0),.din(w_dff_A_gZnyTgn10_0),.clk(gclk));
	jdff dff_A_OovXxVAL4_0(.dout(w_dff_A_XeYo21uv6_0),.din(w_dff_A_OovXxVAL4_0),.clk(gclk));
	jdff dff_A_XeYo21uv6_0(.dout(w_dff_A_EoG4hnUo0_0),.din(w_dff_A_XeYo21uv6_0),.clk(gclk));
	jdff dff_A_EoG4hnUo0_0(.dout(w_dff_A_Xe6emeEV6_0),.din(w_dff_A_EoG4hnUo0_0),.clk(gclk));
	jdff dff_A_Xe6emeEV6_0(.dout(G923),.din(w_dff_A_Xe6emeEV6_0),.clk(gclk));
	jdff dff_A_NmT0XjCB0_1(.dout(w_dff_A_RZMcr9ml7_0),.din(w_dff_A_NmT0XjCB0_1),.clk(gclk));
	jdff dff_A_RZMcr9ml7_0(.dout(w_dff_A_n5rXPReW6_0),.din(w_dff_A_RZMcr9ml7_0),.clk(gclk));
	jdff dff_A_n5rXPReW6_0(.dout(w_dff_A_ixu9Ajnm3_0),.din(w_dff_A_n5rXPReW6_0),.clk(gclk));
	jdff dff_A_ixu9Ajnm3_0(.dout(w_dff_A_uawdFRIq5_0),.din(w_dff_A_ixu9Ajnm3_0),.clk(gclk));
	jdff dff_A_uawdFRIq5_0(.dout(w_dff_A_97KL3mNg1_0),.din(w_dff_A_uawdFRIq5_0),.clk(gclk));
	jdff dff_A_97KL3mNg1_0(.dout(w_dff_A_pms3kupZ5_0),.din(w_dff_A_97KL3mNg1_0),.clk(gclk));
	jdff dff_A_pms3kupZ5_0(.dout(w_dff_A_TRzUWzqA9_0),.din(w_dff_A_pms3kupZ5_0),.clk(gclk));
	jdff dff_A_TRzUWzqA9_0(.dout(w_dff_A_4GOOIoBm5_0),.din(w_dff_A_TRzUWzqA9_0),.clk(gclk));
	jdff dff_A_4GOOIoBm5_0(.dout(w_dff_A_ILzC5j1Y5_0),.din(w_dff_A_4GOOIoBm5_0),.clk(gclk));
	jdff dff_A_ILzC5j1Y5_0(.dout(w_dff_A_2KgoG5uF9_0),.din(w_dff_A_ILzC5j1Y5_0),.clk(gclk));
	jdff dff_A_2KgoG5uF9_0(.dout(w_dff_A_rCHZvA3y5_0),.din(w_dff_A_2KgoG5uF9_0),.clk(gclk));
	jdff dff_A_rCHZvA3y5_0(.dout(w_dff_A_Q8wagKWl2_0),.din(w_dff_A_rCHZvA3y5_0),.clk(gclk));
	jdff dff_A_Q8wagKWl2_0(.dout(w_dff_A_vlO09x095_0),.din(w_dff_A_Q8wagKWl2_0),.clk(gclk));
	jdff dff_A_vlO09x095_0(.dout(w_dff_A_hHuvKOIz6_0),.din(w_dff_A_vlO09x095_0),.clk(gclk));
	jdff dff_A_hHuvKOIz6_0(.dout(w_dff_A_3HceagY58_0),.din(w_dff_A_hHuvKOIz6_0),.clk(gclk));
	jdff dff_A_3HceagY58_0(.dout(w_dff_A_SlaJdS6O3_0),.din(w_dff_A_3HceagY58_0),.clk(gclk));
	jdff dff_A_SlaJdS6O3_0(.dout(w_dff_A_Z0wJn0BU4_0),.din(w_dff_A_SlaJdS6O3_0),.clk(gclk));
	jdff dff_A_Z0wJn0BU4_0(.dout(w_dff_A_PMJ4zAW60_0),.din(w_dff_A_Z0wJn0BU4_0),.clk(gclk));
	jdff dff_A_PMJ4zAW60_0(.dout(w_dff_A_0ZzEXFnr9_0),.din(w_dff_A_PMJ4zAW60_0),.clk(gclk));
	jdff dff_A_0ZzEXFnr9_0(.dout(w_dff_A_MVqRmjUv6_0),.din(w_dff_A_0ZzEXFnr9_0),.clk(gclk));
	jdff dff_A_MVqRmjUv6_0(.dout(w_dff_A_iNYzOTkj1_0),.din(w_dff_A_MVqRmjUv6_0),.clk(gclk));
	jdff dff_A_iNYzOTkj1_0(.dout(w_dff_A_zC9HvHJF1_0),.din(w_dff_A_iNYzOTkj1_0),.clk(gclk));
	jdff dff_A_zC9HvHJF1_0(.dout(w_dff_A_yEObtYBs5_0),.din(w_dff_A_zC9HvHJF1_0),.clk(gclk));
	jdff dff_A_yEObtYBs5_0(.dout(w_dff_A_2jxIV3B49_0),.din(w_dff_A_yEObtYBs5_0),.clk(gclk));
	jdff dff_A_2jxIV3B49_0(.dout(G921),.din(w_dff_A_2jxIV3B49_0),.clk(gclk));
	jdff dff_A_FwI0aGbj2_1(.dout(w_dff_A_XHPaJRCE4_0),.din(w_dff_A_FwI0aGbj2_1),.clk(gclk));
	jdff dff_A_XHPaJRCE4_0(.dout(w_dff_A_Mhc8ZdV60_0),.din(w_dff_A_XHPaJRCE4_0),.clk(gclk));
	jdff dff_A_Mhc8ZdV60_0(.dout(w_dff_A_InkJaXhL9_0),.din(w_dff_A_Mhc8ZdV60_0),.clk(gclk));
	jdff dff_A_InkJaXhL9_0(.dout(w_dff_A_3k09P2nw0_0),.din(w_dff_A_InkJaXhL9_0),.clk(gclk));
	jdff dff_A_3k09P2nw0_0(.dout(w_dff_A_ndQSjTAy5_0),.din(w_dff_A_3k09P2nw0_0),.clk(gclk));
	jdff dff_A_ndQSjTAy5_0(.dout(w_dff_A_z4Vz3Q9U8_0),.din(w_dff_A_ndQSjTAy5_0),.clk(gclk));
	jdff dff_A_z4Vz3Q9U8_0(.dout(w_dff_A_MolwkUZP4_0),.din(w_dff_A_z4Vz3Q9U8_0),.clk(gclk));
	jdff dff_A_MolwkUZP4_0(.dout(w_dff_A_lMu4vz877_0),.din(w_dff_A_MolwkUZP4_0),.clk(gclk));
	jdff dff_A_lMu4vz877_0(.dout(w_dff_A_1xNYFVuB7_0),.din(w_dff_A_lMu4vz877_0),.clk(gclk));
	jdff dff_A_1xNYFVuB7_0(.dout(w_dff_A_92MBFYl93_0),.din(w_dff_A_1xNYFVuB7_0),.clk(gclk));
	jdff dff_A_92MBFYl93_0(.dout(w_dff_A_A1R43ry02_0),.din(w_dff_A_92MBFYl93_0),.clk(gclk));
	jdff dff_A_A1R43ry02_0(.dout(w_dff_A_mi3U7mX09_0),.din(w_dff_A_A1R43ry02_0),.clk(gclk));
	jdff dff_A_mi3U7mX09_0(.dout(w_dff_A_J4z8VsmN4_0),.din(w_dff_A_mi3U7mX09_0),.clk(gclk));
	jdff dff_A_J4z8VsmN4_0(.dout(w_dff_A_cALNuMci9_0),.din(w_dff_A_J4z8VsmN4_0),.clk(gclk));
	jdff dff_A_cALNuMci9_0(.dout(w_dff_A_tHyB8OW05_0),.din(w_dff_A_cALNuMci9_0),.clk(gclk));
	jdff dff_A_tHyB8OW05_0(.dout(w_dff_A_cjPvDO8B7_0),.din(w_dff_A_tHyB8OW05_0),.clk(gclk));
	jdff dff_A_cjPvDO8B7_0(.dout(w_dff_A_1vUF3bQz3_0),.din(w_dff_A_cjPvDO8B7_0),.clk(gclk));
	jdff dff_A_1vUF3bQz3_0(.dout(w_dff_A_OwwzloIQ9_0),.din(w_dff_A_1vUF3bQz3_0),.clk(gclk));
	jdff dff_A_OwwzloIQ9_0(.dout(w_dff_A_YYP46nOo1_0),.din(w_dff_A_OwwzloIQ9_0),.clk(gclk));
	jdff dff_A_YYP46nOo1_0(.dout(w_dff_A_SuKMQElZ8_0),.din(w_dff_A_YYP46nOo1_0),.clk(gclk));
	jdff dff_A_SuKMQElZ8_0(.dout(w_dff_A_SeUcB0pi6_0),.din(w_dff_A_SuKMQElZ8_0),.clk(gclk));
	jdff dff_A_SeUcB0pi6_0(.dout(w_dff_A_TSnMP6gk0_0),.din(w_dff_A_SeUcB0pi6_0),.clk(gclk));
	jdff dff_A_TSnMP6gk0_0(.dout(w_dff_A_mIPC2zON9_0),.din(w_dff_A_TSnMP6gk0_0),.clk(gclk));
	jdff dff_A_mIPC2zON9_0(.dout(w_dff_A_9Ueuxn9R0_0),.din(w_dff_A_mIPC2zON9_0),.clk(gclk));
	jdff dff_A_9Ueuxn9R0_0(.dout(G892),.din(w_dff_A_9Ueuxn9R0_0),.clk(gclk));
	jdff dff_A_IM6ysSsv4_1(.dout(w_dff_A_zY63OBZr1_0),.din(w_dff_A_IM6ysSsv4_1),.clk(gclk));
	jdff dff_A_zY63OBZr1_0(.dout(w_dff_A_ktX1edDQ1_0),.din(w_dff_A_zY63OBZr1_0),.clk(gclk));
	jdff dff_A_ktX1edDQ1_0(.dout(w_dff_A_QJZkZGhW5_0),.din(w_dff_A_ktX1edDQ1_0),.clk(gclk));
	jdff dff_A_QJZkZGhW5_0(.dout(w_dff_A_WAeZpLlO6_0),.din(w_dff_A_QJZkZGhW5_0),.clk(gclk));
	jdff dff_A_WAeZpLlO6_0(.dout(w_dff_A_A7bdGS0l1_0),.din(w_dff_A_WAeZpLlO6_0),.clk(gclk));
	jdff dff_A_A7bdGS0l1_0(.dout(w_dff_A_XlA4f5kQ4_0),.din(w_dff_A_A7bdGS0l1_0),.clk(gclk));
	jdff dff_A_XlA4f5kQ4_0(.dout(w_dff_A_e4AlmKNp9_0),.din(w_dff_A_XlA4f5kQ4_0),.clk(gclk));
	jdff dff_A_e4AlmKNp9_0(.dout(w_dff_A_aKQt76y24_0),.din(w_dff_A_e4AlmKNp9_0),.clk(gclk));
	jdff dff_A_aKQt76y24_0(.dout(w_dff_A_a3EsAeRB6_0),.din(w_dff_A_aKQt76y24_0),.clk(gclk));
	jdff dff_A_a3EsAeRB6_0(.dout(w_dff_A_PoGMbfkG8_0),.din(w_dff_A_a3EsAeRB6_0),.clk(gclk));
	jdff dff_A_PoGMbfkG8_0(.dout(w_dff_A_QJOSBcQ79_0),.din(w_dff_A_PoGMbfkG8_0),.clk(gclk));
	jdff dff_A_QJOSBcQ79_0(.dout(w_dff_A_qh2QGmt83_0),.din(w_dff_A_QJOSBcQ79_0),.clk(gclk));
	jdff dff_A_qh2QGmt83_0(.dout(w_dff_A_tPJmWqXF3_0),.din(w_dff_A_qh2QGmt83_0),.clk(gclk));
	jdff dff_A_tPJmWqXF3_0(.dout(w_dff_A_6j2Kddnx8_0),.din(w_dff_A_tPJmWqXF3_0),.clk(gclk));
	jdff dff_A_6j2Kddnx8_0(.dout(w_dff_A_VJkgFuuW7_0),.din(w_dff_A_6j2Kddnx8_0),.clk(gclk));
	jdff dff_A_VJkgFuuW7_0(.dout(w_dff_A_NmESWnZK6_0),.din(w_dff_A_VJkgFuuW7_0),.clk(gclk));
	jdff dff_A_NmESWnZK6_0(.dout(w_dff_A_SHBUuRdc2_0),.din(w_dff_A_NmESWnZK6_0),.clk(gclk));
	jdff dff_A_SHBUuRdc2_0(.dout(w_dff_A_JV1R3ej42_0),.din(w_dff_A_SHBUuRdc2_0),.clk(gclk));
	jdff dff_A_JV1R3ej42_0(.dout(w_dff_A_7uLaISER7_0),.din(w_dff_A_JV1R3ej42_0),.clk(gclk));
	jdff dff_A_7uLaISER7_0(.dout(w_dff_A_Gl01ovTA0_0),.din(w_dff_A_7uLaISER7_0),.clk(gclk));
	jdff dff_A_Gl01ovTA0_0(.dout(w_dff_A_c9eWRvHJ3_0),.din(w_dff_A_Gl01ovTA0_0),.clk(gclk));
	jdff dff_A_c9eWRvHJ3_0(.dout(w_dff_A_2zS9LLHd5_0),.din(w_dff_A_c9eWRvHJ3_0),.clk(gclk));
	jdff dff_A_2zS9LLHd5_0(.dout(w_dff_A_q7TqjPED9_0),.din(w_dff_A_2zS9LLHd5_0),.clk(gclk));
	jdff dff_A_q7TqjPED9_0(.dout(w_dff_A_r9Ba313H0_0),.din(w_dff_A_q7TqjPED9_0),.clk(gclk));
	jdff dff_A_r9Ba313H0_0(.dout(G887),.din(w_dff_A_r9Ba313H0_0),.clk(gclk));
	jdff dff_A_ELUGCjOB6_1(.dout(w_dff_A_nCOVKXJW4_0),.din(w_dff_A_ELUGCjOB6_1),.clk(gclk));
	jdff dff_A_nCOVKXJW4_0(.dout(w_dff_A_gDFQfVk81_0),.din(w_dff_A_nCOVKXJW4_0),.clk(gclk));
	jdff dff_A_gDFQfVk81_0(.dout(w_dff_A_x1x58NKi6_0),.din(w_dff_A_gDFQfVk81_0),.clk(gclk));
	jdff dff_A_x1x58NKi6_0(.dout(w_dff_A_DADGKog67_0),.din(w_dff_A_x1x58NKi6_0),.clk(gclk));
	jdff dff_A_DADGKog67_0(.dout(w_dff_A_s3y8BDx91_0),.din(w_dff_A_DADGKog67_0),.clk(gclk));
	jdff dff_A_s3y8BDx91_0(.dout(w_dff_A_adgIwvf93_0),.din(w_dff_A_s3y8BDx91_0),.clk(gclk));
	jdff dff_A_adgIwvf93_0(.dout(w_dff_A_uQ4JskQk3_0),.din(w_dff_A_adgIwvf93_0),.clk(gclk));
	jdff dff_A_uQ4JskQk3_0(.dout(w_dff_A_DdINJAaW6_0),.din(w_dff_A_uQ4JskQk3_0),.clk(gclk));
	jdff dff_A_DdINJAaW6_0(.dout(w_dff_A_3n3LtgKK4_0),.din(w_dff_A_DdINJAaW6_0),.clk(gclk));
	jdff dff_A_3n3LtgKK4_0(.dout(w_dff_A_6ZgYHm3y4_0),.din(w_dff_A_3n3LtgKK4_0),.clk(gclk));
	jdff dff_A_6ZgYHm3y4_0(.dout(w_dff_A_mBmZXUZ80_0),.din(w_dff_A_6ZgYHm3y4_0),.clk(gclk));
	jdff dff_A_mBmZXUZ80_0(.dout(w_dff_A_rsAcAc5H9_0),.din(w_dff_A_mBmZXUZ80_0),.clk(gclk));
	jdff dff_A_rsAcAc5H9_0(.dout(w_dff_A_XtXrAGbu0_0),.din(w_dff_A_rsAcAc5H9_0),.clk(gclk));
	jdff dff_A_XtXrAGbu0_0(.dout(w_dff_A_tyukI0qE2_0),.din(w_dff_A_XtXrAGbu0_0),.clk(gclk));
	jdff dff_A_tyukI0qE2_0(.dout(w_dff_A_DsSsIf3L7_0),.din(w_dff_A_tyukI0qE2_0),.clk(gclk));
	jdff dff_A_DsSsIf3L7_0(.dout(w_dff_A_qHLc86ct6_0),.din(w_dff_A_DsSsIf3L7_0),.clk(gclk));
	jdff dff_A_qHLc86ct6_0(.dout(w_dff_A_shdq50ZH0_0),.din(w_dff_A_qHLc86ct6_0),.clk(gclk));
	jdff dff_A_shdq50ZH0_0(.dout(w_dff_A_j5IFX4Zg0_0),.din(w_dff_A_shdq50ZH0_0),.clk(gclk));
	jdff dff_A_j5IFX4Zg0_0(.dout(w_dff_A_vCy38a642_0),.din(w_dff_A_j5IFX4Zg0_0),.clk(gclk));
	jdff dff_A_vCy38a642_0(.dout(w_dff_A_VD7wn6bm6_0),.din(w_dff_A_vCy38a642_0),.clk(gclk));
	jdff dff_A_VD7wn6bm6_0(.dout(w_dff_A_TJXtEoKU1_0),.din(w_dff_A_VD7wn6bm6_0),.clk(gclk));
	jdff dff_A_TJXtEoKU1_0(.dout(w_dff_A_JO5766qF6_0),.din(w_dff_A_TJXtEoKU1_0),.clk(gclk));
	jdff dff_A_JO5766qF6_0(.dout(w_dff_A_4rNpAa2X8_0),.din(w_dff_A_JO5766qF6_0),.clk(gclk));
	jdff dff_A_4rNpAa2X8_0(.dout(w_dff_A_Z42TPgXx5_0),.din(w_dff_A_4rNpAa2X8_0),.clk(gclk));
	jdff dff_A_Z42TPgXx5_0(.dout(G606),.din(w_dff_A_Z42TPgXx5_0),.clk(gclk));
	jdff dff_A_keD9V7g93_2(.dout(w_dff_A_6No7jZ3l5_0),.din(w_dff_A_keD9V7g93_2),.clk(gclk));
	jdff dff_A_6No7jZ3l5_0(.dout(w_dff_A_YwCOvnJB1_0),.din(w_dff_A_6No7jZ3l5_0),.clk(gclk));
	jdff dff_A_YwCOvnJB1_0(.dout(w_dff_A_e2Zwj5m62_0),.din(w_dff_A_YwCOvnJB1_0),.clk(gclk));
	jdff dff_A_e2Zwj5m62_0(.dout(w_dff_A_jj23SIgP4_0),.din(w_dff_A_e2Zwj5m62_0),.clk(gclk));
	jdff dff_A_jj23SIgP4_0(.dout(w_dff_A_IpvWiYMh2_0),.din(w_dff_A_jj23SIgP4_0),.clk(gclk));
	jdff dff_A_IpvWiYMh2_0(.dout(w_dff_A_RRAU7Feh9_0),.din(w_dff_A_IpvWiYMh2_0),.clk(gclk));
	jdff dff_A_RRAU7Feh9_0(.dout(w_dff_A_Rs4lQiv80_0),.din(w_dff_A_RRAU7Feh9_0),.clk(gclk));
	jdff dff_A_Rs4lQiv80_0(.dout(w_dff_A_TaIA0Syt7_0),.din(w_dff_A_Rs4lQiv80_0),.clk(gclk));
	jdff dff_A_TaIA0Syt7_0(.dout(w_dff_A_Xl2iu4F66_0),.din(w_dff_A_TaIA0Syt7_0),.clk(gclk));
	jdff dff_A_Xl2iu4F66_0(.dout(w_dff_A_vTMnpaNz6_0),.din(w_dff_A_Xl2iu4F66_0),.clk(gclk));
	jdff dff_A_vTMnpaNz6_0(.dout(w_dff_A_D9yertSl6_0),.din(w_dff_A_vTMnpaNz6_0),.clk(gclk));
	jdff dff_A_D9yertSl6_0(.dout(w_dff_A_Yb8R0NBp9_0),.din(w_dff_A_D9yertSl6_0),.clk(gclk));
	jdff dff_A_Yb8R0NBp9_0(.dout(w_dff_A_zoiV8HqI0_0),.din(w_dff_A_Yb8R0NBp9_0),.clk(gclk));
	jdff dff_A_zoiV8HqI0_0(.dout(w_dff_A_frH1zcVH3_0),.din(w_dff_A_zoiV8HqI0_0),.clk(gclk));
	jdff dff_A_frH1zcVH3_0(.dout(w_dff_A_jlSvN7Gi6_0),.din(w_dff_A_frH1zcVH3_0),.clk(gclk));
	jdff dff_A_jlSvN7Gi6_0(.dout(w_dff_A_l2yUoy9h5_0),.din(w_dff_A_jlSvN7Gi6_0),.clk(gclk));
	jdff dff_A_l2yUoy9h5_0(.dout(w_dff_A_zoYPNHe88_0),.din(w_dff_A_l2yUoy9h5_0),.clk(gclk));
	jdff dff_A_zoYPNHe88_0(.dout(w_dff_A_bwEjAIaO7_0),.din(w_dff_A_zoYPNHe88_0),.clk(gclk));
	jdff dff_A_bwEjAIaO7_0(.dout(w_dff_A_w7sR6eES9_0),.din(w_dff_A_bwEjAIaO7_0),.clk(gclk));
	jdff dff_A_w7sR6eES9_0(.dout(w_dff_A_AsVarqsG3_0),.din(w_dff_A_w7sR6eES9_0),.clk(gclk));
	jdff dff_A_AsVarqsG3_0(.dout(w_dff_A_uJzgPcEF4_0),.din(w_dff_A_AsVarqsG3_0),.clk(gclk));
	jdff dff_A_uJzgPcEF4_0(.dout(w_dff_A_PeVg3iqd4_0),.din(w_dff_A_uJzgPcEF4_0),.clk(gclk));
	jdff dff_A_PeVg3iqd4_0(.dout(G656),.din(w_dff_A_PeVg3iqd4_0),.clk(gclk));
	jdff dff_A_x86FEGCI7_2(.dout(w_dff_A_QZa27yH73_0),.din(w_dff_A_x86FEGCI7_2),.clk(gclk));
	jdff dff_A_QZa27yH73_0(.dout(w_dff_A_b9fGvEec6_0),.din(w_dff_A_QZa27yH73_0),.clk(gclk));
	jdff dff_A_b9fGvEec6_0(.dout(w_dff_A_iGk5muXF6_0),.din(w_dff_A_b9fGvEec6_0),.clk(gclk));
	jdff dff_A_iGk5muXF6_0(.dout(w_dff_A_Gh3424E94_0),.din(w_dff_A_iGk5muXF6_0),.clk(gclk));
	jdff dff_A_Gh3424E94_0(.dout(w_dff_A_LCebUzlT4_0),.din(w_dff_A_Gh3424E94_0),.clk(gclk));
	jdff dff_A_LCebUzlT4_0(.dout(w_dff_A_PxdHmspX4_0),.din(w_dff_A_LCebUzlT4_0),.clk(gclk));
	jdff dff_A_PxdHmspX4_0(.dout(w_dff_A_TivC2nGk7_0),.din(w_dff_A_PxdHmspX4_0),.clk(gclk));
	jdff dff_A_TivC2nGk7_0(.dout(w_dff_A_u9Lazg1R2_0),.din(w_dff_A_TivC2nGk7_0),.clk(gclk));
	jdff dff_A_u9Lazg1R2_0(.dout(w_dff_A_Vsi66rb35_0),.din(w_dff_A_u9Lazg1R2_0),.clk(gclk));
	jdff dff_A_Vsi66rb35_0(.dout(w_dff_A_Z1fiM0vR6_0),.din(w_dff_A_Vsi66rb35_0),.clk(gclk));
	jdff dff_A_Z1fiM0vR6_0(.dout(w_dff_A_3NZ0yDjb3_0),.din(w_dff_A_Z1fiM0vR6_0),.clk(gclk));
	jdff dff_A_3NZ0yDjb3_0(.dout(w_dff_A_6SUEWyFS5_0),.din(w_dff_A_3NZ0yDjb3_0),.clk(gclk));
	jdff dff_A_6SUEWyFS5_0(.dout(w_dff_A_YSCxAza49_0),.din(w_dff_A_6SUEWyFS5_0),.clk(gclk));
	jdff dff_A_YSCxAza49_0(.dout(w_dff_A_BlGFREtI4_0),.din(w_dff_A_YSCxAza49_0),.clk(gclk));
	jdff dff_A_BlGFREtI4_0(.dout(w_dff_A_s5FtIMzv5_0),.din(w_dff_A_BlGFREtI4_0),.clk(gclk));
	jdff dff_A_s5FtIMzv5_0(.dout(w_dff_A_00AvwFTZ2_0),.din(w_dff_A_s5FtIMzv5_0),.clk(gclk));
	jdff dff_A_00AvwFTZ2_0(.dout(w_dff_A_hhMxq2Tc8_0),.din(w_dff_A_00AvwFTZ2_0),.clk(gclk));
	jdff dff_A_hhMxq2Tc8_0(.dout(w_dff_A_fMEkWrrV5_0),.din(w_dff_A_hhMxq2Tc8_0),.clk(gclk));
	jdff dff_A_fMEkWrrV5_0(.dout(w_dff_A_rkNNEXs64_0),.din(w_dff_A_fMEkWrrV5_0),.clk(gclk));
	jdff dff_A_rkNNEXs64_0(.dout(w_dff_A_aOJlDXK89_0),.din(w_dff_A_rkNNEXs64_0),.clk(gclk));
	jdff dff_A_aOJlDXK89_0(.dout(w_dff_A_vS5vbLYA1_0),.din(w_dff_A_aOJlDXK89_0),.clk(gclk));
	jdff dff_A_vS5vbLYA1_0(.dout(w_dff_A_KofkMd3a9_0),.din(w_dff_A_vS5vbLYA1_0),.clk(gclk));
	jdff dff_A_KofkMd3a9_0(.dout(w_dff_A_0g7TGgoS7_0),.din(w_dff_A_KofkMd3a9_0),.clk(gclk));
	jdff dff_A_0g7TGgoS7_0(.dout(G809),.din(w_dff_A_0g7TGgoS7_0),.clk(gclk));
	jdff dff_A_YeaIpaov7_1(.dout(w_dff_A_jiXK9IhC9_0),.din(w_dff_A_YeaIpaov7_1),.clk(gclk));
	jdff dff_A_jiXK9IhC9_0(.dout(w_dff_A_0iaZKLE90_0),.din(w_dff_A_jiXK9IhC9_0),.clk(gclk));
	jdff dff_A_0iaZKLE90_0(.dout(w_dff_A_o39kVAQT8_0),.din(w_dff_A_0iaZKLE90_0),.clk(gclk));
	jdff dff_A_o39kVAQT8_0(.dout(w_dff_A_BtRLGDEP0_0),.din(w_dff_A_o39kVAQT8_0),.clk(gclk));
	jdff dff_A_BtRLGDEP0_0(.dout(w_dff_A_99i7LAPF7_0),.din(w_dff_A_BtRLGDEP0_0),.clk(gclk));
	jdff dff_A_99i7LAPF7_0(.dout(w_dff_A_57O3sZWL4_0),.din(w_dff_A_99i7LAPF7_0),.clk(gclk));
	jdff dff_A_57O3sZWL4_0(.dout(w_dff_A_xlNFVysj3_0),.din(w_dff_A_57O3sZWL4_0),.clk(gclk));
	jdff dff_A_xlNFVysj3_0(.dout(w_dff_A_XrLXivbj2_0),.din(w_dff_A_xlNFVysj3_0),.clk(gclk));
	jdff dff_A_XrLXivbj2_0(.dout(w_dff_A_L6iGirEZ7_0),.din(w_dff_A_XrLXivbj2_0),.clk(gclk));
	jdff dff_A_L6iGirEZ7_0(.dout(w_dff_A_2JxubHvP6_0),.din(w_dff_A_L6iGirEZ7_0),.clk(gclk));
	jdff dff_A_2JxubHvP6_0(.dout(w_dff_A_BZKSH1bR1_0),.din(w_dff_A_2JxubHvP6_0),.clk(gclk));
	jdff dff_A_BZKSH1bR1_0(.dout(w_dff_A_o1MoDGsA2_0),.din(w_dff_A_BZKSH1bR1_0),.clk(gclk));
	jdff dff_A_o1MoDGsA2_0(.dout(w_dff_A_MkJoJj2e9_0),.din(w_dff_A_o1MoDGsA2_0),.clk(gclk));
	jdff dff_A_MkJoJj2e9_0(.dout(w_dff_A_948uc08y8_0),.din(w_dff_A_MkJoJj2e9_0),.clk(gclk));
	jdff dff_A_948uc08y8_0(.dout(w_dff_A_zRXXoYv12_0),.din(w_dff_A_948uc08y8_0),.clk(gclk));
	jdff dff_A_zRXXoYv12_0(.dout(w_dff_A_Z9DbpMDw3_0),.din(w_dff_A_zRXXoYv12_0),.clk(gclk));
	jdff dff_A_Z9DbpMDw3_0(.dout(w_dff_A_wFCG80GU4_0),.din(w_dff_A_Z9DbpMDw3_0),.clk(gclk));
	jdff dff_A_wFCG80GU4_0(.dout(w_dff_A_aygIYzC69_0),.din(w_dff_A_wFCG80GU4_0),.clk(gclk));
	jdff dff_A_aygIYzC69_0(.dout(w_dff_A_xwJ2ZW0q4_0),.din(w_dff_A_aygIYzC69_0),.clk(gclk));
	jdff dff_A_xwJ2ZW0q4_0(.dout(w_dff_A_KwXllmL38_0),.din(w_dff_A_xwJ2ZW0q4_0),.clk(gclk));
	jdff dff_A_KwXllmL38_0(.dout(w_dff_A_Ebnw4n3T0_0),.din(w_dff_A_KwXllmL38_0),.clk(gclk));
	jdff dff_A_Ebnw4n3T0_0(.dout(w_dff_A_GLVGhJ037_0),.din(w_dff_A_Ebnw4n3T0_0),.clk(gclk));
	jdff dff_A_GLVGhJ037_0(.dout(w_dff_A_jcMUFEnB7_0),.din(w_dff_A_GLVGhJ037_0),.clk(gclk));
	jdff dff_A_jcMUFEnB7_0(.dout(w_dff_A_TvHVLmIo4_0),.din(w_dff_A_jcMUFEnB7_0),.clk(gclk));
	jdff dff_A_TvHVLmIo4_0(.dout(G993),.din(w_dff_A_TvHVLmIo4_0),.clk(gclk));
	jdff dff_A_SpO2BMhM3_1(.dout(w_dff_A_jCo04NMI5_0),.din(w_dff_A_SpO2BMhM3_1),.clk(gclk));
	jdff dff_A_jCo04NMI5_0(.dout(w_dff_A_47nucgNw2_0),.din(w_dff_A_jCo04NMI5_0),.clk(gclk));
	jdff dff_A_47nucgNw2_0(.dout(w_dff_A_kWzdgH5L4_0),.din(w_dff_A_47nucgNw2_0),.clk(gclk));
	jdff dff_A_kWzdgH5L4_0(.dout(w_dff_A_UqajSPWh9_0),.din(w_dff_A_kWzdgH5L4_0),.clk(gclk));
	jdff dff_A_UqajSPWh9_0(.dout(w_dff_A_JKzZdKFE9_0),.din(w_dff_A_UqajSPWh9_0),.clk(gclk));
	jdff dff_A_JKzZdKFE9_0(.dout(w_dff_A_jJba68X70_0),.din(w_dff_A_JKzZdKFE9_0),.clk(gclk));
	jdff dff_A_jJba68X70_0(.dout(w_dff_A_4GlW8KNG1_0),.din(w_dff_A_jJba68X70_0),.clk(gclk));
	jdff dff_A_4GlW8KNG1_0(.dout(w_dff_A_uFgZRCcw0_0),.din(w_dff_A_4GlW8KNG1_0),.clk(gclk));
	jdff dff_A_uFgZRCcw0_0(.dout(w_dff_A_X5fIxnN13_0),.din(w_dff_A_uFgZRCcw0_0),.clk(gclk));
	jdff dff_A_X5fIxnN13_0(.dout(w_dff_A_UXfhf2CA5_0),.din(w_dff_A_X5fIxnN13_0),.clk(gclk));
	jdff dff_A_UXfhf2CA5_0(.dout(w_dff_A_nRP8m8mD1_0),.din(w_dff_A_UXfhf2CA5_0),.clk(gclk));
	jdff dff_A_nRP8m8mD1_0(.dout(w_dff_A_aiFZ5ciw2_0),.din(w_dff_A_nRP8m8mD1_0),.clk(gclk));
	jdff dff_A_aiFZ5ciw2_0(.dout(w_dff_A_qHkjQACn7_0),.din(w_dff_A_aiFZ5ciw2_0),.clk(gclk));
	jdff dff_A_qHkjQACn7_0(.dout(w_dff_A_qjEkwSO13_0),.din(w_dff_A_qHkjQACn7_0),.clk(gclk));
	jdff dff_A_qjEkwSO13_0(.dout(w_dff_A_s81eWuvH7_0),.din(w_dff_A_qjEkwSO13_0),.clk(gclk));
	jdff dff_A_s81eWuvH7_0(.dout(w_dff_A_Mw9uFUtC9_0),.din(w_dff_A_s81eWuvH7_0),.clk(gclk));
	jdff dff_A_Mw9uFUtC9_0(.dout(w_dff_A_8PszQ2VZ8_0),.din(w_dff_A_Mw9uFUtC9_0),.clk(gclk));
	jdff dff_A_8PszQ2VZ8_0(.dout(w_dff_A_kQXK6ufu9_0),.din(w_dff_A_8PszQ2VZ8_0),.clk(gclk));
	jdff dff_A_kQXK6ufu9_0(.dout(w_dff_A_03d5zdZt4_0),.din(w_dff_A_kQXK6ufu9_0),.clk(gclk));
	jdff dff_A_03d5zdZt4_0(.dout(w_dff_A_meMuVMTn9_0),.din(w_dff_A_03d5zdZt4_0),.clk(gclk));
	jdff dff_A_meMuVMTn9_0(.dout(w_dff_A_4VSEAS7z3_0),.din(w_dff_A_meMuVMTn9_0),.clk(gclk));
	jdff dff_A_4VSEAS7z3_0(.dout(w_dff_A_OhWZ7Kp21_0),.din(w_dff_A_4VSEAS7z3_0),.clk(gclk));
	jdff dff_A_OhWZ7Kp21_0(.dout(w_dff_A_L5bNWsc53_0),.din(w_dff_A_OhWZ7Kp21_0),.clk(gclk));
	jdff dff_A_L5bNWsc53_0(.dout(w_dff_A_OtBO3pev2_0),.din(w_dff_A_L5bNWsc53_0),.clk(gclk));
	jdff dff_A_OtBO3pev2_0(.dout(G978),.din(w_dff_A_OtBO3pev2_0),.clk(gclk));
	jdff dff_A_abVhkHvY7_1(.dout(w_dff_A_V85JZFxw4_0),.din(w_dff_A_abVhkHvY7_1),.clk(gclk));
	jdff dff_A_V85JZFxw4_0(.dout(w_dff_A_d3Gpi8Jc0_0),.din(w_dff_A_V85JZFxw4_0),.clk(gclk));
	jdff dff_A_d3Gpi8Jc0_0(.dout(w_dff_A_jcmEfclu4_0),.din(w_dff_A_d3Gpi8Jc0_0),.clk(gclk));
	jdff dff_A_jcmEfclu4_0(.dout(w_dff_A_Yb6Nbclj0_0),.din(w_dff_A_jcmEfclu4_0),.clk(gclk));
	jdff dff_A_Yb6Nbclj0_0(.dout(w_dff_A_R1AK6bSL6_0),.din(w_dff_A_Yb6Nbclj0_0),.clk(gclk));
	jdff dff_A_R1AK6bSL6_0(.dout(w_dff_A_R8FvGvkB6_0),.din(w_dff_A_R1AK6bSL6_0),.clk(gclk));
	jdff dff_A_R8FvGvkB6_0(.dout(w_dff_A_kcFAIxA96_0),.din(w_dff_A_R8FvGvkB6_0),.clk(gclk));
	jdff dff_A_kcFAIxA96_0(.dout(w_dff_A_qZIX0z0i8_0),.din(w_dff_A_kcFAIxA96_0),.clk(gclk));
	jdff dff_A_qZIX0z0i8_0(.dout(w_dff_A_famX9DUw0_0),.din(w_dff_A_qZIX0z0i8_0),.clk(gclk));
	jdff dff_A_famX9DUw0_0(.dout(w_dff_A_gNC84Z308_0),.din(w_dff_A_famX9DUw0_0),.clk(gclk));
	jdff dff_A_gNC84Z308_0(.dout(w_dff_A_ofIv66Zj4_0),.din(w_dff_A_gNC84Z308_0),.clk(gclk));
	jdff dff_A_ofIv66Zj4_0(.dout(w_dff_A_w6uY1qWn7_0),.din(w_dff_A_ofIv66Zj4_0),.clk(gclk));
	jdff dff_A_w6uY1qWn7_0(.dout(w_dff_A_6LpPMPaN4_0),.din(w_dff_A_w6uY1qWn7_0),.clk(gclk));
	jdff dff_A_6LpPMPaN4_0(.dout(w_dff_A_xEfkJmnA8_0),.din(w_dff_A_6LpPMPaN4_0),.clk(gclk));
	jdff dff_A_xEfkJmnA8_0(.dout(w_dff_A_8G9h2CEO0_0),.din(w_dff_A_xEfkJmnA8_0),.clk(gclk));
	jdff dff_A_8G9h2CEO0_0(.dout(w_dff_A_XKpVDc3B3_0),.din(w_dff_A_8G9h2CEO0_0),.clk(gclk));
	jdff dff_A_XKpVDc3B3_0(.dout(w_dff_A_ebKE19mp1_0),.din(w_dff_A_XKpVDc3B3_0),.clk(gclk));
	jdff dff_A_ebKE19mp1_0(.dout(w_dff_A_lBxUdizI1_0),.din(w_dff_A_ebKE19mp1_0),.clk(gclk));
	jdff dff_A_lBxUdizI1_0(.dout(w_dff_A_XRZtbF221_0),.din(w_dff_A_lBxUdizI1_0),.clk(gclk));
	jdff dff_A_XRZtbF221_0(.dout(w_dff_A_FUWpOhri7_0),.din(w_dff_A_XRZtbF221_0),.clk(gclk));
	jdff dff_A_FUWpOhri7_0(.dout(w_dff_A_eOzo2qa53_0),.din(w_dff_A_FUWpOhri7_0),.clk(gclk));
	jdff dff_A_eOzo2qa53_0(.dout(w_dff_A_jznu23Zk0_0),.din(w_dff_A_eOzo2qa53_0),.clk(gclk));
	jdff dff_A_jznu23Zk0_0(.dout(w_dff_A_9YXdI7EP2_0),.din(w_dff_A_jznu23Zk0_0),.clk(gclk));
	jdff dff_A_9YXdI7EP2_0(.dout(w_dff_A_ML9mQqH98_0),.din(w_dff_A_9YXdI7EP2_0),.clk(gclk));
	jdff dff_A_ML9mQqH98_0(.dout(G949),.din(w_dff_A_ML9mQqH98_0),.clk(gclk));
	jdff dff_A_qpWbjoOy4_1(.dout(w_dff_A_oaFPvoaF5_0),.din(w_dff_A_qpWbjoOy4_1),.clk(gclk));
	jdff dff_A_oaFPvoaF5_0(.dout(w_dff_A_TrKS8yWm2_0),.din(w_dff_A_oaFPvoaF5_0),.clk(gclk));
	jdff dff_A_TrKS8yWm2_0(.dout(w_dff_A_E4VJRHTl3_0),.din(w_dff_A_TrKS8yWm2_0),.clk(gclk));
	jdff dff_A_E4VJRHTl3_0(.dout(w_dff_A_mXSY4zYP5_0),.din(w_dff_A_E4VJRHTl3_0),.clk(gclk));
	jdff dff_A_mXSY4zYP5_0(.dout(w_dff_A_w9A5TP2H2_0),.din(w_dff_A_mXSY4zYP5_0),.clk(gclk));
	jdff dff_A_w9A5TP2H2_0(.dout(w_dff_A_VlZUHRa21_0),.din(w_dff_A_w9A5TP2H2_0),.clk(gclk));
	jdff dff_A_VlZUHRa21_0(.dout(w_dff_A_IvtZ7P7g1_0),.din(w_dff_A_VlZUHRa21_0),.clk(gclk));
	jdff dff_A_IvtZ7P7g1_0(.dout(w_dff_A_BfS3k26j9_0),.din(w_dff_A_IvtZ7P7g1_0),.clk(gclk));
	jdff dff_A_BfS3k26j9_0(.dout(w_dff_A_JOfFvtra7_0),.din(w_dff_A_BfS3k26j9_0),.clk(gclk));
	jdff dff_A_JOfFvtra7_0(.dout(w_dff_A_KvfZLhqi5_0),.din(w_dff_A_JOfFvtra7_0),.clk(gclk));
	jdff dff_A_KvfZLhqi5_0(.dout(w_dff_A_9y1c4S6c9_0),.din(w_dff_A_KvfZLhqi5_0),.clk(gclk));
	jdff dff_A_9y1c4S6c9_0(.dout(w_dff_A_ZojNuHXZ5_0),.din(w_dff_A_9y1c4S6c9_0),.clk(gclk));
	jdff dff_A_ZojNuHXZ5_0(.dout(w_dff_A_xpH9CXJM5_0),.din(w_dff_A_ZojNuHXZ5_0),.clk(gclk));
	jdff dff_A_xpH9CXJM5_0(.dout(w_dff_A_fKaLlKz50_0),.din(w_dff_A_xpH9CXJM5_0),.clk(gclk));
	jdff dff_A_fKaLlKz50_0(.dout(w_dff_A_6MgvSZpQ6_0),.din(w_dff_A_fKaLlKz50_0),.clk(gclk));
	jdff dff_A_6MgvSZpQ6_0(.dout(w_dff_A_AqsUbGqI2_0),.din(w_dff_A_6MgvSZpQ6_0),.clk(gclk));
	jdff dff_A_AqsUbGqI2_0(.dout(w_dff_A_sHrKWhtn6_0),.din(w_dff_A_AqsUbGqI2_0),.clk(gclk));
	jdff dff_A_sHrKWhtn6_0(.dout(w_dff_A_k4QmlshR7_0),.din(w_dff_A_sHrKWhtn6_0),.clk(gclk));
	jdff dff_A_k4QmlshR7_0(.dout(w_dff_A_ptLqqP2h2_0),.din(w_dff_A_k4QmlshR7_0),.clk(gclk));
	jdff dff_A_ptLqqP2h2_0(.dout(w_dff_A_TiUNK2D95_0),.din(w_dff_A_ptLqqP2h2_0),.clk(gclk));
	jdff dff_A_TiUNK2D95_0(.dout(w_dff_A_uKi4mG2o3_0),.din(w_dff_A_TiUNK2D95_0),.clk(gclk));
	jdff dff_A_uKi4mG2o3_0(.dout(w_dff_A_EstgPHQC2_0),.din(w_dff_A_uKi4mG2o3_0),.clk(gclk));
	jdff dff_A_EstgPHQC2_0(.dout(w_dff_A_TkpcScS52_0),.din(w_dff_A_EstgPHQC2_0),.clk(gclk));
	jdff dff_A_TkpcScS52_0(.dout(w_dff_A_wsNhdpVO8_0),.din(w_dff_A_TkpcScS52_0),.clk(gclk));
	jdff dff_A_wsNhdpVO8_0(.dout(G939),.din(w_dff_A_wsNhdpVO8_0),.clk(gclk));
	jdff dff_A_lD6XExhc7_1(.dout(w_dff_A_Jl4ZNpnA1_0),.din(w_dff_A_lD6XExhc7_1),.clk(gclk));
	jdff dff_A_Jl4ZNpnA1_0(.dout(w_dff_A_YRcS2ikS6_0),.din(w_dff_A_Jl4ZNpnA1_0),.clk(gclk));
	jdff dff_A_YRcS2ikS6_0(.dout(w_dff_A_c9n10fjS4_0),.din(w_dff_A_YRcS2ikS6_0),.clk(gclk));
	jdff dff_A_c9n10fjS4_0(.dout(w_dff_A_QTjUCbq50_0),.din(w_dff_A_c9n10fjS4_0),.clk(gclk));
	jdff dff_A_QTjUCbq50_0(.dout(w_dff_A_XMibHe3f4_0),.din(w_dff_A_QTjUCbq50_0),.clk(gclk));
	jdff dff_A_XMibHe3f4_0(.dout(w_dff_A_Hgy08DiC8_0),.din(w_dff_A_XMibHe3f4_0),.clk(gclk));
	jdff dff_A_Hgy08DiC8_0(.dout(w_dff_A_ty6mWJ6Y6_0),.din(w_dff_A_Hgy08DiC8_0),.clk(gclk));
	jdff dff_A_ty6mWJ6Y6_0(.dout(w_dff_A_NcpEUnwM2_0),.din(w_dff_A_ty6mWJ6Y6_0),.clk(gclk));
	jdff dff_A_NcpEUnwM2_0(.dout(w_dff_A_zHy5uA2U5_0),.din(w_dff_A_NcpEUnwM2_0),.clk(gclk));
	jdff dff_A_zHy5uA2U5_0(.dout(w_dff_A_k6LFJOLP7_0),.din(w_dff_A_zHy5uA2U5_0),.clk(gclk));
	jdff dff_A_k6LFJOLP7_0(.dout(w_dff_A_GQGhDm5G4_0),.din(w_dff_A_k6LFJOLP7_0),.clk(gclk));
	jdff dff_A_GQGhDm5G4_0(.dout(w_dff_A_iiw7dC0S9_0),.din(w_dff_A_GQGhDm5G4_0),.clk(gclk));
	jdff dff_A_iiw7dC0S9_0(.dout(w_dff_A_pGv4YvHQ3_0),.din(w_dff_A_iiw7dC0S9_0),.clk(gclk));
	jdff dff_A_pGv4YvHQ3_0(.dout(w_dff_A_ReWdVeme4_0),.din(w_dff_A_pGv4YvHQ3_0),.clk(gclk));
	jdff dff_A_ReWdVeme4_0(.dout(w_dff_A_IDiLCvME8_0),.din(w_dff_A_ReWdVeme4_0),.clk(gclk));
	jdff dff_A_IDiLCvME8_0(.dout(w_dff_A_ATyGnFjX3_0),.din(w_dff_A_IDiLCvME8_0),.clk(gclk));
	jdff dff_A_ATyGnFjX3_0(.dout(w_dff_A_FsvZQZ7i2_0),.din(w_dff_A_ATyGnFjX3_0),.clk(gclk));
	jdff dff_A_FsvZQZ7i2_0(.dout(w_dff_A_RsX6UkSY0_0),.din(w_dff_A_FsvZQZ7i2_0),.clk(gclk));
	jdff dff_A_RsX6UkSY0_0(.dout(w_dff_A_EsQzUZc85_0),.din(w_dff_A_RsX6UkSY0_0),.clk(gclk));
	jdff dff_A_EsQzUZc85_0(.dout(w_dff_A_brVQAggx3_0),.din(w_dff_A_EsQzUZc85_0),.clk(gclk));
	jdff dff_A_brVQAggx3_0(.dout(w_dff_A_cwqWPGr07_0),.din(w_dff_A_brVQAggx3_0),.clk(gclk));
	jdff dff_A_cwqWPGr07_0(.dout(w_dff_A_dVrG7hGV7_0),.din(w_dff_A_cwqWPGr07_0),.clk(gclk));
	jdff dff_A_dVrG7hGV7_0(.dout(w_dff_A_FrYoED5t0_0),.din(w_dff_A_dVrG7hGV7_0),.clk(gclk));
	jdff dff_A_FrYoED5t0_0(.dout(w_dff_A_TpleHrMc4_0),.din(w_dff_A_FrYoED5t0_0),.clk(gclk));
	jdff dff_A_TpleHrMc4_0(.dout(G889),.din(w_dff_A_TpleHrMc4_0),.clk(gclk));
	jdff dff_A_4e4EIA5N1_1(.dout(w_dff_A_NNj3eLVc1_0),.din(w_dff_A_4e4EIA5N1_1),.clk(gclk));
	jdff dff_A_NNj3eLVc1_0(.dout(w_dff_A_3HlQ2bnD6_0),.din(w_dff_A_NNj3eLVc1_0),.clk(gclk));
	jdff dff_A_3HlQ2bnD6_0(.dout(w_dff_A_K0APsira4_0),.din(w_dff_A_3HlQ2bnD6_0),.clk(gclk));
	jdff dff_A_K0APsira4_0(.dout(w_dff_A_5mirhI067_0),.din(w_dff_A_K0APsira4_0),.clk(gclk));
	jdff dff_A_5mirhI067_0(.dout(w_dff_A_SgChimeS9_0),.din(w_dff_A_5mirhI067_0),.clk(gclk));
	jdff dff_A_SgChimeS9_0(.dout(w_dff_A_I7tJAHJo4_0),.din(w_dff_A_SgChimeS9_0),.clk(gclk));
	jdff dff_A_I7tJAHJo4_0(.dout(w_dff_A_jEORaBQ79_0),.din(w_dff_A_I7tJAHJo4_0),.clk(gclk));
	jdff dff_A_jEORaBQ79_0(.dout(w_dff_A_981HW88k6_0),.din(w_dff_A_jEORaBQ79_0),.clk(gclk));
	jdff dff_A_981HW88k6_0(.dout(w_dff_A_rAG8wnC35_0),.din(w_dff_A_981HW88k6_0),.clk(gclk));
	jdff dff_A_rAG8wnC35_0(.dout(w_dff_A_yEMSOdVg2_0),.din(w_dff_A_rAG8wnC35_0),.clk(gclk));
	jdff dff_A_yEMSOdVg2_0(.dout(w_dff_A_7H2nFOht3_0),.din(w_dff_A_yEMSOdVg2_0),.clk(gclk));
	jdff dff_A_7H2nFOht3_0(.dout(w_dff_A_0fRBeq0C1_0),.din(w_dff_A_7H2nFOht3_0),.clk(gclk));
	jdff dff_A_0fRBeq0C1_0(.dout(w_dff_A_8X4qeEpt1_0),.din(w_dff_A_0fRBeq0C1_0),.clk(gclk));
	jdff dff_A_8X4qeEpt1_0(.dout(w_dff_A_ja6OvJz09_0),.din(w_dff_A_8X4qeEpt1_0),.clk(gclk));
	jdff dff_A_ja6OvJz09_0(.dout(w_dff_A_FpJLk7TL0_0),.din(w_dff_A_ja6OvJz09_0),.clk(gclk));
	jdff dff_A_FpJLk7TL0_0(.dout(w_dff_A_LzWbjckA9_0),.din(w_dff_A_FpJLk7TL0_0),.clk(gclk));
	jdff dff_A_LzWbjckA9_0(.dout(w_dff_A_s9R8RfWi8_0),.din(w_dff_A_LzWbjckA9_0),.clk(gclk));
	jdff dff_A_s9R8RfWi8_0(.dout(w_dff_A_pqgIY3NN1_0),.din(w_dff_A_s9R8RfWi8_0),.clk(gclk));
	jdff dff_A_pqgIY3NN1_0(.dout(w_dff_A_26dtetRk3_0),.din(w_dff_A_pqgIY3NN1_0),.clk(gclk));
	jdff dff_A_26dtetRk3_0(.dout(w_dff_A_h3Zg1kjR9_0),.din(w_dff_A_26dtetRk3_0),.clk(gclk));
	jdff dff_A_h3Zg1kjR9_0(.dout(w_dff_A_EtvJhjP99_0),.din(w_dff_A_h3Zg1kjR9_0),.clk(gclk));
	jdff dff_A_EtvJhjP99_0(.dout(w_dff_A_yiqcB09d7_0),.din(w_dff_A_EtvJhjP99_0),.clk(gclk));
	jdff dff_A_yiqcB09d7_0(.dout(w_dff_A_iCRYLmRz2_0),.din(w_dff_A_yiqcB09d7_0),.clk(gclk));
	jdff dff_A_iCRYLmRz2_0(.dout(w_dff_A_Uhx4mFUf4_0),.din(w_dff_A_iCRYLmRz2_0),.clk(gclk));
	jdff dff_A_Uhx4mFUf4_0(.dout(G593),.din(w_dff_A_Uhx4mFUf4_0),.clk(gclk));
	jdff dff_A_5DKWnxSc5_2(.dout(w_dff_A_xVQWH6Tr1_0),.din(w_dff_A_5DKWnxSc5_2),.clk(gclk));
	jdff dff_A_xVQWH6Tr1_0(.dout(w_dff_A_uI2A11gr1_0),.din(w_dff_A_xVQWH6Tr1_0),.clk(gclk));
	jdff dff_A_uI2A11gr1_0(.dout(w_dff_A_xr7y9Smy1_0),.din(w_dff_A_uI2A11gr1_0),.clk(gclk));
	jdff dff_A_xr7y9Smy1_0(.dout(w_dff_A_E4DmUa6Y8_0),.din(w_dff_A_xr7y9Smy1_0),.clk(gclk));
	jdff dff_A_E4DmUa6Y8_0(.dout(w_dff_A_KCPLWmcP4_0),.din(w_dff_A_E4DmUa6Y8_0),.clk(gclk));
	jdff dff_A_KCPLWmcP4_0(.dout(w_dff_A_6WVWdltR0_0),.din(w_dff_A_KCPLWmcP4_0),.clk(gclk));
	jdff dff_A_6WVWdltR0_0(.dout(w_dff_A_ahA86vOb6_0),.din(w_dff_A_6WVWdltR0_0),.clk(gclk));
	jdff dff_A_ahA86vOb6_0(.dout(w_dff_A_6KcVJOQL8_0),.din(w_dff_A_ahA86vOb6_0),.clk(gclk));
	jdff dff_A_6KcVJOQL8_0(.dout(w_dff_A_oIjlbJoV5_0),.din(w_dff_A_6KcVJOQL8_0),.clk(gclk));
	jdff dff_A_oIjlbJoV5_0(.dout(w_dff_A_x57fBEvW9_0),.din(w_dff_A_oIjlbJoV5_0),.clk(gclk));
	jdff dff_A_x57fBEvW9_0(.dout(w_dff_A_YwmGE3Am3_0),.din(w_dff_A_x57fBEvW9_0),.clk(gclk));
	jdff dff_A_YwmGE3Am3_0(.dout(w_dff_A_pd1p2vGz2_0),.din(w_dff_A_YwmGE3Am3_0),.clk(gclk));
	jdff dff_A_pd1p2vGz2_0(.dout(w_dff_A_nKTgTCH18_0),.din(w_dff_A_pd1p2vGz2_0),.clk(gclk));
	jdff dff_A_nKTgTCH18_0(.dout(w_dff_A_QP5hFykY0_0),.din(w_dff_A_nKTgTCH18_0),.clk(gclk));
	jdff dff_A_QP5hFykY0_0(.dout(w_dff_A_WeoXHbwr4_0),.din(w_dff_A_QP5hFykY0_0),.clk(gclk));
	jdff dff_A_WeoXHbwr4_0(.dout(w_dff_A_Ydk4Ner15_0),.din(w_dff_A_WeoXHbwr4_0),.clk(gclk));
	jdff dff_A_Ydk4Ner15_0(.dout(w_dff_A_uI1fL5E10_0),.din(w_dff_A_Ydk4Ner15_0),.clk(gclk));
	jdff dff_A_uI1fL5E10_0(.dout(w_dff_A_NhiN46YI3_0),.din(w_dff_A_uI1fL5E10_0),.clk(gclk));
	jdff dff_A_NhiN46YI3_0(.dout(w_dff_A_BvVZYSyB5_0),.din(w_dff_A_NhiN46YI3_0),.clk(gclk));
	jdff dff_A_BvVZYSyB5_0(.dout(w_dff_A_CPpuDR8l0_0),.din(w_dff_A_BvVZYSyB5_0),.clk(gclk));
	jdff dff_A_CPpuDR8l0_0(.dout(w_dff_A_2AJPeBJv2_0),.din(w_dff_A_CPpuDR8l0_0),.clk(gclk));
	jdff dff_A_2AJPeBJv2_0(.dout(G636),.din(w_dff_A_2AJPeBJv2_0),.clk(gclk));
	jdff dff_A_CXKw5YL30_2(.dout(w_dff_A_sN8DakQO6_0),.din(w_dff_A_CXKw5YL30_2),.clk(gclk));
	jdff dff_A_sN8DakQO6_0(.dout(w_dff_A_JcOoUIoU0_0),.din(w_dff_A_sN8DakQO6_0),.clk(gclk));
	jdff dff_A_JcOoUIoU0_0(.dout(w_dff_A_AMQ9nWoi5_0),.din(w_dff_A_JcOoUIoU0_0),.clk(gclk));
	jdff dff_A_AMQ9nWoi5_0(.dout(w_dff_A_ffv8D3iP0_0),.din(w_dff_A_AMQ9nWoi5_0),.clk(gclk));
	jdff dff_A_ffv8D3iP0_0(.dout(w_dff_A_NLkBdWcm3_0),.din(w_dff_A_ffv8D3iP0_0),.clk(gclk));
	jdff dff_A_NLkBdWcm3_0(.dout(w_dff_A_rkUBQDy35_0),.din(w_dff_A_NLkBdWcm3_0),.clk(gclk));
	jdff dff_A_rkUBQDy35_0(.dout(w_dff_A_gYFtotOP3_0),.din(w_dff_A_rkUBQDy35_0),.clk(gclk));
	jdff dff_A_gYFtotOP3_0(.dout(w_dff_A_WHcSynkR0_0),.din(w_dff_A_gYFtotOP3_0),.clk(gclk));
	jdff dff_A_WHcSynkR0_0(.dout(w_dff_A_lBDItlpU6_0),.din(w_dff_A_WHcSynkR0_0),.clk(gclk));
	jdff dff_A_lBDItlpU6_0(.dout(w_dff_A_07oRUG598_0),.din(w_dff_A_lBDItlpU6_0),.clk(gclk));
	jdff dff_A_07oRUG598_0(.dout(w_dff_A_luXZfeUs5_0),.din(w_dff_A_07oRUG598_0),.clk(gclk));
	jdff dff_A_luXZfeUs5_0(.dout(w_dff_A_zVtXFOHs9_0),.din(w_dff_A_luXZfeUs5_0),.clk(gclk));
	jdff dff_A_zVtXFOHs9_0(.dout(w_dff_A_WGsCsiRH9_0),.din(w_dff_A_zVtXFOHs9_0),.clk(gclk));
	jdff dff_A_WGsCsiRH9_0(.dout(w_dff_A_NweTt4l64_0),.din(w_dff_A_WGsCsiRH9_0),.clk(gclk));
	jdff dff_A_NweTt4l64_0(.dout(w_dff_A_if2qgv0H6_0),.din(w_dff_A_NweTt4l64_0),.clk(gclk));
	jdff dff_A_if2qgv0H6_0(.dout(w_dff_A_wAsJxjbj2_0),.din(w_dff_A_if2qgv0H6_0),.clk(gclk));
	jdff dff_A_wAsJxjbj2_0(.dout(w_dff_A_9xIy5x3z4_0),.din(w_dff_A_wAsJxjbj2_0),.clk(gclk));
	jdff dff_A_9xIy5x3z4_0(.dout(w_dff_A_6JOjYtxb7_0),.din(w_dff_A_9xIy5x3z4_0),.clk(gclk));
	jdff dff_A_6JOjYtxb7_0(.dout(w_dff_A_cRKkT0PC0_0),.din(w_dff_A_6JOjYtxb7_0),.clk(gclk));
	jdff dff_A_cRKkT0PC0_0(.dout(w_dff_A_aItKAicj2_0),.din(w_dff_A_cRKkT0PC0_0),.clk(gclk));
	jdff dff_A_aItKAicj2_0(.dout(w_dff_A_wTQCLBXD0_0),.din(w_dff_A_aItKAicj2_0),.clk(gclk));
	jdff dff_A_wTQCLBXD0_0(.dout(G704),.din(w_dff_A_wTQCLBXD0_0),.clk(gclk));
	jdff dff_A_TR3QSKJ91_2(.dout(w_dff_A_RkLtvXpE6_0),.din(w_dff_A_TR3QSKJ91_2),.clk(gclk));
	jdff dff_A_RkLtvXpE6_0(.dout(w_dff_A_z0TMj8TG3_0),.din(w_dff_A_RkLtvXpE6_0),.clk(gclk));
	jdff dff_A_z0TMj8TG3_0(.dout(w_dff_A_64wFIkQ95_0),.din(w_dff_A_z0TMj8TG3_0),.clk(gclk));
	jdff dff_A_64wFIkQ95_0(.dout(w_dff_A_puWSMKTF7_0),.din(w_dff_A_64wFIkQ95_0),.clk(gclk));
	jdff dff_A_puWSMKTF7_0(.dout(w_dff_A_dk9tfpKv2_0),.din(w_dff_A_puWSMKTF7_0),.clk(gclk));
	jdff dff_A_dk9tfpKv2_0(.dout(w_dff_A_8tTZc8Kw2_0),.din(w_dff_A_dk9tfpKv2_0),.clk(gclk));
	jdff dff_A_8tTZc8Kw2_0(.dout(w_dff_A_Xevm6M2H3_0),.din(w_dff_A_8tTZc8Kw2_0),.clk(gclk));
	jdff dff_A_Xevm6M2H3_0(.dout(w_dff_A_FyPeZUxw6_0),.din(w_dff_A_Xevm6M2H3_0),.clk(gclk));
	jdff dff_A_FyPeZUxw6_0(.dout(w_dff_A_9aTbQNIu4_0),.din(w_dff_A_FyPeZUxw6_0),.clk(gclk));
	jdff dff_A_9aTbQNIu4_0(.dout(w_dff_A_nzxuVn7x7_0),.din(w_dff_A_9aTbQNIu4_0),.clk(gclk));
	jdff dff_A_nzxuVn7x7_0(.dout(w_dff_A_gLUPRY4w4_0),.din(w_dff_A_nzxuVn7x7_0),.clk(gclk));
	jdff dff_A_gLUPRY4w4_0(.dout(w_dff_A_PBKA6CSE2_0),.din(w_dff_A_gLUPRY4w4_0),.clk(gclk));
	jdff dff_A_PBKA6CSE2_0(.dout(w_dff_A_40L5QOHL3_0),.din(w_dff_A_PBKA6CSE2_0),.clk(gclk));
	jdff dff_A_40L5QOHL3_0(.dout(w_dff_A_VDZx6CGd6_0),.din(w_dff_A_40L5QOHL3_0),.clk(gclk));
	jdff dff_A_VDZx6CGd6_0(.dout(w_dff_A_wr4CqXl23_0),.din(w_dff_A_VDZx6CGd6_0),.clk(gclk));
	jdff dff_A_wr4CqXl23_0(.dout(w_dff_A_TjeCiBd20_0),.din(w_dff_A_wr4CqXl23_0),.clk(gclk));
	jdff dff_A_TjeCiBd20_0(.dout(w_dff_A_jh06xNKB8_0),.din(w_dff_A_TjeCiBd20_0),.clk(gclk));
	jdff dff_A_jh06xNKB8_0(.dout(w_dff_A_xpbmMFm96_0),.din(w_dff_A_jh06xNKB8_0),.clk(gclk));
	jdff dff_A_xpbmMFm96_0(.dout(w_dff_A_3X92xAxM1_0),.din(w_dff_A_xpbmMFm96_0),.clk(gclk));
	jdff dff_A_3X92xAxM1_0(.dout(w_dff_A_3aVTff5Z7_0),.din(w_dff_A_3X92xAxM1_0),.clk(gclk));
	jdff dff_A_3aVTff5Z7_0(.dout(w_dff_A_wISkywuW2_0),.din(w_dff_A_3aVTff5Z7_0),.clk(gclk));
	jdff dff_A_wISkywuW2_0(.dout(G717),.din(w_dff_A_wISkywuW2_0),.clk(gclk));
	jdff dff_A_9yC0VVfO7_2(.dout(w_dff_A_jFXPlW4o6_0),.din(w_dff_A_9yC0VVfO7_2),.clk(gclk));
	jdff dff_A_jFXPlW4o6_0(.dout(w_dff_A_xJpXaXBX8_0),.din(w_dff_A_jFXPlW4o6_0),.clk(gclk));
	jdff dff_A_xJpXaXBX8_0(.dout(w_dff_A_5kSP9aBD0_0),.din(w_dff_A_xJpXaXBX8_0),.clk(gclk));
	jdff dff_A_5kSP9aBD0_0(.dout(w_dff_A_zNTpmbIP0_0),.din(w_dff_A_5kSP9aBD0_0),.clk(gclk));
	jdff dff_A_zNTpmbIP0_0(.dout(w_dff_A_a2AJYJZY2_0),.din(w_dff_A_zNTpmbIP0_0),.clk(gclk));
	jdff dff_A_a2AJYJZY2_0(.dout(w_dff_A_S7QEW4ah1_0),.din(w_dff_A_a2AJYJZY2_0),.clk(gclk));
	jdff dff_A_S7QEW4ah1_0(.dout(w_dff_A_9NJzThi50_0),.din(w_dff_A_S7QEW4ah1_0),.clk(gclk));
	jdff dff_A_9NJzThi50_0(.dout(w_dff_A_ilQaAq009_0),.din(w_dff_A_9NJzThi50_0),.clk(gclk));
	jdff dff_A_ilQaAq009_0(.dout(w_dff_A_I6OnOS4L9_0),.din(w_dff_A_ilQaAq009_0),.clk(gclk));
	jdff dff_A_I6OnOS4L9_0(.dout(w_dff_A_Kqfm5GjQ8_0),.din(w_dff_A_I6OnOS4L9_0),.clk(gclk));
	jdff dff_A_Kqfm5GjQ8_0(.dout(w_dff_A_DQQxTDK83_0),.din(w_dff_A_Kqfm5GjQ8_0),.clk(gclk));
	jdff dff_A_DQQxTDK83_0(.dout(w_dff_A_2z7dsrkQ1_0),.din(w_dff_A_DQQxTDK83_0),.clk(gclk));
	jdff dff_A_2z7dsrkQ1_0(.dout(w_dff_A_7xiub2BF7_0),.din(w_dff_A_2z7dsrkQ1_0),.clk(gclk));
	jdff dff_A_7xiub2BF7_0(.dout(w_dff_A_pj51po7o9_0),.din(w_dff_A_7xiub2BF7_0),.clk(gclk));
	jdff dff_A_pj51po7o9_0(.dout(w_dff_A_jekEyZBi1_0),.din(w_dff_A_pj51po7o9_0),.clk(gclk));
	jdff dff_A_jekEyZBi1_0(.dout(w_dff_A_1mn3SqOD2_0),.din(w_dff_A_jekEyZBi1_0),.clk(gclk));
	jdff dff_A_1mn3SqOD2_0(.dout(w_dff_A_A90jU8Hx4_0),.din(w_dff_A_1mn3SqOD2_0),.clk(gclk));
	jdff dff_A_A90jU8Hx4_0(.dout(w_dff_A_NS9tbqK98_0),.din(w_dff_A_A90jU8Hx4_0),.clk(gclk));
	jdff dff_A_NS9tbqK98_0(.dout(w_dff_A_TGZ9z4nW7_0),.din(w_dff_A_NS9tbqK98_0),.clk(gclk));
	jdff dff_A_TGZ9z4nW7_0(.dout(w_dff_A_ymbLtiM65_0),.din(w_dff_A_TGZ9z4nW7_0),.clk(gclk));
	jdff dff_A_ymbLtiM65_0(.dout(w_dff_A_D3s1irdO4_0),.din(w_dff_A_ymbLtiM65_0),.clk(gclk));
	jdff dff_A_D3s1irdO4_0(.dout(w_dff_A_lQWDjGuG1_0),.din(w_dff_A_D3s1irdO4_0),.clk(gclk));
	jdff dff_A_lQWDjGuG1_0(.dout(G820),.din(w_dff_A_lQWDjGuG1_0),.clk(gclk));
	jdff dff_A_rizW0C430_2(.dout(w_dff_A_KgAAbwuH8_0),.din(w_dff_A_rizW0C430_2),.clk(gclk));
	jdff dff_A_KgAAbwuH8_0(.dout(w_dff_A_7nnuyk1Q2_0),.din(w_dff_A_KgAAbwuH8_0),.clk(gclk));
	jdff dff_A_7nnuyk1Q2_0(.dout(w_dff_A_vYgPw98P2_0),.din(w_dff_A_7nnuyk1Q2_0),.clk(gclk));
	jdff dff_A_vYgPw98P2_0(.dout(w_dff_A_GiHiMhTQ7_0),.din(w_dff_A_vYgPw98P2_0),.clk(gclk));
	jdff dff_A_GiHiMhTQ7_0(.dout(w_dff_A_AUqkSgAN4_0),.din(w_dff_A_GiHiMhTQ7_0),.clk(gclk));
	jdff dff_A_AUqkSgAN4_0(.dout(w_dff_A_aDDEqaYT7_0),.din(w_dff_A_AUqkSgAN4_0),.clk(gclk));
	jdff dff_A_aDDEqaYT7_0(.dout(w_dff_A_wChBvq3p6_0),.din(w_dff_A_aDDEqaYT7_0),.clk(gclk));
	jdff dff_A_wChBvq3p6_0(.dout(w_dff_A_vJm1Pm654_0),.din(w_dff_A_wChBvq3p6_0),.clk(gclk));
	jdff dff_A_vJm1Pm654_0(.dout(w_dff_A_MQroQ7IC1_0),.din(w_dff_A_vJm1Pm654_0),.clk(gclk));
	jdff dff_A_MQroQ7IC1_0(.dout(w_dff_A_GiyvZx260_0),.din(w_dff_A_MQroQ7IC1_0),.clk(gclk));
	jdff dff_A_GiyvZx260_0(.dout(w_dff_A_jcrhMJgS8_0),.din(w_dff_A_GiyvZx260_0),.clk(gclk));
	jdff dff_A_jcrhMJgS8_0(.dout(w_dff_A_gs4gCJG75_0),.din(w_dff_A_jcrhMJgS8_0),.clk(gclk));
	jdff dff_A_gs4gCJG75_0(.dout(w_dff_A_43PrkEhK8_0),.din(w_dff_A_gs4gCJG75_0),.clk(gclk));
	jdff dff_A_43PrkEhK8_0(.dout(w_dff_A_blgBBLO64_0),.din(w_dff_A_43PrkEhK8_0),.clk(gclk));
	jdff dff_A_blgBBLO64_0(.dout(w_dff_A_Mn3y9pAO6_0),.din(w_dff_A_blgBBLO64_0),.clk(gclk));
	jdff dff_A_Mn3y9pAO6_0(.dout(w_dff_A_OmwUq7pT7_0),.din(w_dff_A_Mn3y9pAO6_0),.clk(gclk));
	jdff dff_A_OmwUq7pT7_0(.dout(w_dff_A_wTIzYJdY3_0),.din(w_dff_A_OmwUq7pT7_0),.clk(gclk));
	jdff dff_A_wTIzYJdY3_0(.dout(w_dff_A_X6fMt0Zj0_0),.din(w_dff_A_wTIzYJdY3_0),.clk(gclk));
	jdff dff_A_X6fMt0Zj0_0(.dout(w_dff_A_kU02qcPQ1_0),.din(w_dff_A_X6fMt0Zj0_0),.clk(gclk));
	jdff dff_A_kU02qcPQ1_0(.dout(w_dff_A_adtuXUxE0_0),.din(w_dff_A_kU02qcPQ1_0),.clk(gclk));
	jdff dff_A_adtuXUxE0_0(.dout(G639),.din(w_dff_A_adtuXUxE0_0),.clk(gclk));
	jdff dff_A_elugQIR87_2(.dout(w_dff_A_vjOvb3W06_0),.din(w_dff_A_elugQIR87_2),.clk(gclk));
	jdff dff_A_vjOvb3W06_0(.dout(w_dff_A_f7oJb32k4_0),.din(w_dff_A_vjOvb3W06_0),.clk(gclk));
	jdff dff_A_f7oJb32k4_0(.dout(w_dff_A_cGLVsDBl2_0),.din(w_dff_A_f7oJb32k4_0),.clk(gclk));
	jdff dff_A_cGLVsDBl2_0(.dout(w_dff_A_LAicCfTh9_0),.din(w_dff_A_cGLVsDBl2_0),.clk(gclk));
	jdff dff_A_LAicCfTh9_0(.dout(w_dff_A_zPpsueOZ2_0),.din(w_dff_A_LAicCfTh9_0),.clk(gclk));
	jdff dff_A_zPpsueOZ2_0(.dout(w_dff_A_ncAURSH36_0),.din(w_dff_A_zPpsueOZ2_0),.clk(gclk));
	jdff dff_A_ncAURSH36_0(.dout(w_dff_A_kCSS4AZq0_0),.din(w_dff_A_ncAURSH36_0),.clk(gclk));
	jdff dff_A_kCSS4AZq0_0(.dout(w_dff_A_NYHD2jE67_0),.din(w_dff_A_kCSS4AZq0_0),.clk(gclk));
	jdff dff_A_NYHD2jE67_0(.dout(w_dff_A_oYi4of0D3_0),.din(w_dff_A_NYHD2jE67_0),.clk(gclk));
	jdff dff_A_oYi4of0D3_0(.dout(w_dff_A_Hb4ytExg0_0),.din(w_dff_A_oYi4of0D3_0),.clk(gclk));
	jdff dff_A_Hb4ytExg0_0(.dout(w_dff_A_mhiIvyDJ5_0),.din(w_dff_A_Hb4ytExg0_0),.clk(gclk));
	jdff dff_A_mhiIvyDJ5_0(.dout(w_dff_A_GMirbeNl4_0),.din(w_dff_A_mhiIvyDJ5_0),.clk(gclk));
	jdff dff_A_GMirbeNl4_0(.dout(w_dff_A_6PHqUvff5_0),.din(w_dff_A_GMirbeNl4_0),.clk(gclk));
	jdff dff_A_6PHqUvff5_0(.dout(w_dff_A_NhBUSYdt2_0),.din(w_dff_A_6PHqUvff5_0),.clk(gclk));
	jdff dff_A_NhBUSYdt2_0(.dout(w_dff_A_njyrBR860_0),.din(w_dff_A_NhBUSYdt2_0),.clk(gclk));
	jdff dff_A_njyrBR860_0(.dout(w_dff_A_0fI8E1tn5_0),.din(w_dff_A_njyrBR860_0),.clk(gclk));
	jdff dff_A_0fI8E1tn5_0(.dout(w_dff_A_LjAQVpdm0_0),.din(w_dff_A_0fI8E1tn5_0),.clk(gclk));
	jdff dff_A_LjAQVpdm0_0(.dout(w_dff_A_hOjv7GI27_0),.din(w_dff_A_LjAQVpdm0_0),.clk(gclk));
	jdff dff_A_hOjv7GI27_0(.dout(w_dff_A_fvRySZuu8_0),.din(w_dff_A_hOjv7GI27_0),.clk(gclk));
	jdff dff_A_fvRySZuu8_0(.dout(w_dff_A_FrydKVP70_0),.din(w_dff_A_fvRySZuu8_0),.clk(gclk));
	jdff dff_A_FrydKVP70_0(.dout(G673),.din(w_dff_A_FrydKVP70_0),.clk(gclk));
	jdff dff_A_FaokHENP3_2(.dout(w_dff_A_0QcR0jCY9_0),.din(w_dff_A_FaokHENP3_2),.clk(gclk));
	jdff dff_A_0QcR0jCY9_0(.dout(w_dff_A_fkXPbOey1_0),.din(w_dff_A_0QcR0jCY9_0),.clk(gclk));
	jdff dff_A_fkXPbOey1_0(.dout(w_dff_A_FBlijyyz1_0),.din(w_dff_A_fkXPbOey1_0),.clk(gclk));
	jdff dff_A_FBlijyyz1_0(.dout(w_dff_A_oaAOkGXK3_0),.din(w_dff_A_FBlijyyz1_0),.clk(gclk));
	jdff dff_A_oaAOkGXK3_0(.dout(w_dff_A_K7S56rVT4_0),.din(w_dff_A_oaAOkGXK3_0),.clk(gclk));
	jdff dff_A_K7S56rVT4_0(.dout(w_dff_A_KCQuRw3E0_0),.din(w_dff_A_K7S56rVT4_0),.clk(gclk));
	jdff dff_A_KCQuRw3E0_0(.dout(w_dff_A_fgZNn9MB6_0),.din(w_dff_A_KCQuRw3E0_0),.clk(gclk));
	jdff dff_A_fgZNn9MB6_0(.dout(w_dff_A_TbSvztVd9_0),.din(w_dff_A_fgZNn9MB6_0),.clk(gclk));
	jdff dff_A_TbSvztVd9_0(.dout(w_dff_A_S7lPsxhh1_0),.din(w_dff_A_TbSvztVd9_0),.clk(gclk));
	jdff dff_A_S7lPsxhh1_0(.dout(w_dff_A_xOKC3ko35_0),.din(w_dff_A_S7lPsxhh1_0),.clk(gclk));
	jdff dff_A_xOKC3ko35_0(.dout(w_dff_A_d3Ip3zeE9_0),.din(w_dff_A_xOKC3ko35_0),.clk(gclk));
	jdff dff_A_d3Ip3zeE9_0(.dout(w_dff_A_64YrB5C19_0),.din(w_dff_A_d3Ip3zeE9_0),.clk(gclk));
	jdff dff_A_64YrB5C19_0(.dout(w_dff_A_iSOwSdHN7_0),.din(w_dff_A_64YrB5C19_0),.clk(gclk));
	jdff dff_A_iSOwSdHN7_0(.dout(w_dff_A_n29ScSW67_0),.din(w_dff_A_iSOwSdHN7_0),.clk(gclk));
	jdff dff_A_n29ScSW67_0(.dout(w_dff_A_xQwsdKbI5_0),.din(w_dff_A_n29ScSW67_0),.clk(gclk));
	jdff dff_A_xQwsdKbI5_0(.dout(w_dff_A_XqEADTOL7_0),.din(w_dff_A_xQwsdKbI5_0),.clk(gclk));
	jdff dff_A_XqEADTOL7_0(.dout(w_dff_A_QXQ2Bv1S2_0),.din(w_dff_A_XqEADTOL7_0),.clk(gclk));
	jdff dff_A_QXQ2Bv1S2_0(.dout(w_dff_A_ao6Jk5qP6_0),.din(w_dff_A_QXQ2Bv1S2_0),.clk(gclk));
	jdff dff_A_ao6Jk5qP6_0(.dout(w_dff_A_xTYZkzUF4_0),.din(w_dff_A_ao6Jk5qP6_0),.clk(gclk));
	jdff dff_A_xTYZkzUF4_0(.dout(w_dff_A_K4tG1aVx5_0),.din(w_dff_A_xTYZkzUF4_0),.clk(gclk));
	jdff dff_A_K4tG1aVx5_0(.dout(G707),.din(w_dff_A_K4tG1aVx5_0),.clk(gclk));
	jdff dff_A_xsbWQ4I27_2(.dout(w_dff_A_ZmxnlbO75_0),.din(w_dff_A_xsbWQ4I27_2),.clk(gclk));
	jdff dff_A_ZmxnlbO75_0(.dout(w_dff_A_pGGRNlkO6_0),.din(w_dff_A_ZmxnlbO75_0),.clk(gclk));
	jdff dff_A_pGGRNlkO6_0(.dout(w_dff_A_vT2fL17A8_0),.din(w_dff_A_pGGRNlkO6_0),.clk(gclk));
	jdff dff_A_vT2fL17A8_0(.dout(w_dff_A_HyQ7vQWy2_0),.din(w_dff_A_vT2fL17A8_0),.clk(gclk));
	jdff dff_A_HyQ7vQWy2_0(.dout(w_dff_A_gUlXqVgu7_0),.din(w_dff_A_HyQ7vQWy2_0),.clk(gclk));
	jdff dff_A_gUlXqVgu7_0(.dout(w_dff_A_mFipyJM54_0),.din(w_dff_A_gUlXqVgu7_0),.clk(gclk));
	jdff dff_A_mFipyJM54_0(.dout(w_dff_A_vnhY7zrE0_0),.din(w_dff_A_mFipyJM54_0),.clk(gclk));
	jdff dff_A_vnhY7zrE0_0(.dout(w_dff_A_zvh8j5m56_0),.din(w_dff_A_vnhY7zrE0_0),.clk(gclk));
	jdff dff_A_zvh8j5m56_0(.dout(w_dff_A_NX87CFfs2_0),.din(w_dff_A_zvh8j5m56_0),.clk(gclk));
	jdff dff_A_NX87CFfs2_0(.dout(w_dff_A_bMeo0Xii2_0),.din(w_dff_A_NX87CFfs2_0),.clk(gclk));
	jdff dff_A_bMeo0Xii2_0(.dout(w_dff_A_0gDixBLJ5_0),.din(w_dff_A_bMeo0Xii2_0),.clk(gclk));
	jdff dff_A_0gDixBLJ5_0(.dout(w_dff_A_ShcqrH7E4_0),.din(w_dff_A_0gDixBLJ5_0),.clk(gclk));
	jdff dff_A_ShcqrH7E4_0(.dout(w_dff_A_uXKUj2lM3_0),.din(w_dff_A_ShcqrH7E4_0),.clk(gclk));
	jdff dff_A_uXKUj2lM3_0(.dout(w_dff_A_ayzisLxe1_0),.din(w_dff_A_uXKUj2lM3_0),.clk(gclk));
	jdff dff_A_ayzisLxe1_0(.dout(w_dff_A_B7C4cCNj4_0),.din(w_dff_A_ayzisLxe1_0),.clk(gclk));
	jdff dff_A_B7C4cCNj4_0(.dout(w_dff_A_VyHL6giX3_0),.din(w_dff_A_B7C4cCNj4_0),.clk(gclk));
	jdff dff_A_VyHL6giX3_0(.dout(w_dff_A_p7En6qza1_0),.din(w_dff_A_VyHL6giX3_0),.clk(gclk));
	jdff dff_A_p7En6qza1_0(.dout(w_dff_A_wlaTIjaE6_0),.din(w_dff_A_p7En6qza1_0),.clk(gclk));
	jdff dff_A_wlaTIjaE6_0(.dout(w_dff_A_ASPWIk2T1_0),.din(w_dff_A_wlaTIjaE6_0),.clk(gclk));
	jdff dff_A_ASPWIk2T1_0(.dout(w_dff_A_6SUGHeB62_0),.din(w_dff_A_ASPWIk2T1_0),.clk(gclk));
	jdff dff_A_6SUGHeB62_0(.dout(G715),.din(w_dff_A_6SUGHeB62_0),.clk(gclk));
	jdff dff_A_BEb53Iaq1_2(.dout(w_dff_A_oloWKfMa0_0),.din(w_dff_A_BEb53Iaq1_2),.clk(gclk));
	jdff dff_A_oloWKfMa0_0(.dout(w_dff_A_pqD3GZ3g8_0),.din(w_dff_A_oloWKfMa0_0),.clk(gclk));
	jdff dff_A_pqD3GZ3g8_0(.dout(w_dff_A_EYGuIKep0_0),.din(w_dff_A_pqD3GZ3g8_0),.clk(gclk));
	jdff dff_A_EYGuIKep0_0(.dout(w_dff_A_9LMeRw9x6_0),.din(w_dff_A_EYGuIKep0_0),.clk(gclk));
	jdff dff_A_9LMeRw9x6_0(.dout(w_dff_A_deNX8pML9_0),.din(w_dff_A_9LMeRw9x6_0),.clk(gclk));
	jdff dff_A_deNX8pML9_0(.dout(w_dff_A_MxDtdVQe0_0),.din(w_dff_A_deNX8pML9_0),.clk(gclk));
	jdff dff_A_MxDtdVQe0_0(.dout(w_dff_A_nl4mcWAu4_0),.din(w_dff_A_MxDtdVQe0_0),.clk(gclk));
	jdff dff_A_nl4mcWAu4_0(.dout(w_dff_A_ewEv8Ybp9_0),.din(w_dff_A_nl4mcWAu4_0),.clk(gclk));
	jdff dff_A_ewEv8Ybp9_0(.dout(w_dff_A_U6aBBlE37_0),.din(w_dff_A_ewEv8Ybp9_0),.clk(gclk));
	jdff dff_A_U6aBBlE37_0(.dout(w_dff_A_sgeIN7sc3_0),.din(w_dff_A_U6aBBlE37_0),.clk(gclk));
	jdff dff_A_sgeIN7sc3_0(.dout(w_dff_A_P1ICeaaJ8_0),.din(w_dff_A_sgeIN7sc3_0),.clk(gclk));
	jdff dff_A_P1ICeaaJ8_0(.dout(w_dff_A_QA7VTbku3_0),.din(w_dff_A_P1ICeaaJ8_0),.clk(gclk));
	jdff dff_A_QA7VTbku3_0(.dout(w_dff_A_sgG74Gx40_0),.din(w_dff_A_QA7VTbku3_0),.clk(gclk));
	jdff dff_A_sgG74Gx40_0(.dout(w_dff_A_CUgQ3iz31_0),.din(w_dff_A_sgG74Gx40_0),.clk(gclk));
	jdff dff_A_CUgQ3iz31_0(.dout(w_dff_A_aJMDk6zR2_0),.din(w_dff_A_CUgQ3iz31_0),.clk(gclk));
	jdff dff_A_aJMDk6zR2_0(.dout(w_dff_A_SUtsIFMm6_0),.din(w_dff_A_aJMDk6zR2_0),.clk(gclk));
	jdff dff_A_SUtsIFMm6_0(.dout(G598),.din(w_dff_A_SUtsIFMm6_0),.clk(gclk));
	jdff dff_A_j4efVi3O6_2(.dout(w_dff_A_Yq0pu1wW0_0),.din(w_dff_A_j4efVi3O6_2),.clk(gclk));
	jdff dff_A_Yq0pu1wW0_0(.dout(w_dff_A_GOBiuBFn1_0),.din(w_dff_A_Yq0pu1wW0_0),.clk(gclk));
	jdff dff_A_GOBiuBFn1_0(.dout(w_dff_A_WbbPGbyL9_0),.din(w_dff_A_GOBiuBFn1_0),.clk(gclk));
	jdff dff_A_WbbPGbyL9_0(.dout(w_dff_A_QUDDyT3N6_0),.din(w_dff_A_WbbPGbyL9_0),.clk(gclk));
	jdff dff_A_QUDDyT3N6_0(.dout(w_dff_A_SRlVGceg3_0),.din(w_dff_A_QUDDyT3N6_0),.clk(gclk));
	jdff dff_A_SRlVGceg3_0(.dout(w_dff_A_uALdLlXS3_0),.din(w_dff_A_SRlVGceg3_0),.clk(gclk));
	jdff dff_A_uALdLlXS3_0(.dout(w_dff_A_5DWrPsbL7_0),.din(w_dff_A_uALdLlXS3_0),.clk(gclk));
	jdff dff_A_5DWrPsbL7_0(.dout(w_dff_A_TJ8wjj571_0),.din(w_dff_A_5DWrPsbL7_0),.clk(gclk));
	jdff dff_A_TJ8wjj571_0(.dout(w_dff_A_g4gbUWNR7_0),.din(w_dff_A_TJ8wjj571_0),.clk(gclk));
	jdff dff_A_g4gbUWNR7_0(.dout(w_dff_A_awoE7okF8_0),.din(w_dff_A_g4gbUWNR7_0),.clk(gclk));
	jdff dff_A_awoE7okF8_0(.dout(w_dff_A_lUxuw5nY6_0),.din(w_dff_A_awoE7okF8_0),.clk(gclk));
	jdff dff_A_lUxuw5nY6_0(.dout(w_dff_A_HON1Q2SL5_0),.din(w_dff_A_lUxuw5nY6_0),.clk(gclk));
	jdff dff_A_HON1Q2SL5_0(.dout(w_dff_A_VA68RU7z1_0),.din(w_dff_A_HON1Q2SL5_0),.clk(gclk));
	jdff dff_A_VA68RU7z1_0(.dout(w_dff_A_iT40JmC66_0),.din(w_dff_A_VA68RU7z1_0),.clk(gclk));
	jdff dff_A_iT40JmC66_0(.dout(w_dff_A_U5oLsT2f1_0),.din(w_dff_A_iT40JmC66_0),.clk(gclk));
	jdff dff_A_U5oLsT2f1_0(.dout(w_dff_A_I4bktKWu6_0),.din(w_dff_A_U5oLsT2f1_0),.clk(gclk));
	jdff dff_A_I4bktKWu6_0(.dout(G610),.din(w_dff_A_I4bktKWu6_0),.clk(gclk));
	jdff dff_A_4Xgg3Wdu6_2(.dout(w_dff_A_1M4z8uvC6_0),.din(w_dff_A_4Xgg3Wdu6_2),.clk(gclk));
	jdff dff_A_1M4z8uvC6_0(.dout(w_dff_A_5FiHU8d02_0),.din(w_dff_A_1M4z8uvC6_0),.clk(gclk));
	jdff dff_A_5FiHU8d02_0(.dout(w_dff_A_tjm3Ww215_0),.din(w_dff_A_5FiHU8d02_0),.clk(gclk));
	jdff dff_A_tjm3Ww215_0(.dout(w_dff_A_71ej5SFX2_0),.din(w_dff_A_tjm3Ww215_0),.clk(gclk));
	jdff dff_A_71ej5SFX2_0(.dout(w_dff_A_TkQReInG0_0),.din(w_dff_A_71ej5SFX2_0),.clk(gclk));
	jdff dff_A_TkQReInG0_0(.dout(w_dff_A_3Nz5jTUP4_0),.din(w_dff_A_TkQReInG0_0),.clk(gclk));
	jdff dff_A_3Nz5jTUP4_0(.dout(w_dff_A_GuaHMZHy1_0),.din(w_dff_A_3Nz5jTUP4_0),.clk(gclk));
	jdff dff_A_GuaHMZHy1_0(.dout(w_dff_A_G3Nt3byh6_0),.din(w_dff_A_GuaHMZHy1_0),.clk(gclk));
	jdff dff_A_G3Nt3byh6_0(.dout(w_dff_A_CJkqSmBs2_0),.din(w_dff_A_G3Nt3byh6_0),.clk(gclk));
	jdff dff_A_CJkqSmBs2_0(.dout(w_dff_A_MN2Ias6m6_0),.din(w_dff_A_CJkqSmBs2_0),.clk(gclk));
	jdff dff_A_MN2Ias6m6_0(.dout(w_dff_A_aWeCwI952_0),.din(w_dff_A_MN2Ias6m6_0),.clk(gclk));
	jdff dff_A_aWeCwI952_0(.dout(w_dff_A_KD0XfKV14_0),.din(w_dff_A_aWeCwI952_0),.clk(gclk));
	jdff dff_A_KD0XfKV14_0(.dout(w_dff_A_IiaX7pO55_0),.din(w_dff_A_KD0XfKV14_0),.clk(gclk));
	jdff dff_A_IiaX7pO55_0(.dout(w_dff_A_LnHzd7tf5_0),.din(w_dff_A_IiaX7pO55_0),.clk(gclk));
	jdff dff_A_LnHzd7tf5_0(.dout(G588),.din(w_dff_A_LnHzd7tf5_0),.clk(gclk));
	jdff dff_A_n3GGxwow0_2(.dout(w_dff_A_BC4hp5hS2_0),.din(w_dff_A_n3GGxwow0_2),.clk(gclk));
	jdff dff_A_BC4hp5hS2_0(.dout(w_dff_A_8Tk9dvqi4_0),.din(w_dff_A_BC4hp5hS2_0),.clk(gclk));
	jdff dff_A_8Tk9dvqi4_0(.dout(w_dff_A_35g2JW3m8_0),.din(w_dff_A_8Tk9dvqi4_0),.clk(gclk));
	jdff dff_A_35g2JW3m8_0(.dout(w_dff_A_HCgQiUjK2_0),.din(w_dff_A_35g2JW3m8_0),.clk(gclk));
	jdff dff_A_HCgQiUjK2_0(.dout(w_dff_A_wzBljx7g8_0),.din(w_dff_A_HCgQiUjK2_0),.clk(gclk));
	jdff dff_A_wzBljx7g8_0(.dout(w_dff_A_t0eXidmG0_0),.din(w_dff_A_wzBljx7g8_0),.clk(gclk));
	jdff dff_A_t0eXidmG0_0(.dout(w_dff_A_Vz2gVHAS2_0),.din(w_dff_A_t0eXidmG0_0),.clk(gclk));
	jdff dff_A_Vz2gVHAS2_0(.dout(w_dff_A_igQvbAAg2_0),.din(w_dff_A_Vz2gVHAS2_0),.clk(gclk));
	jdff dff_A_igQvbAAg2_0(.dout(w_dff_A_dNQgYKEB7_0),.din(w_dff_A_igQvbAAg2_0),.clk(gclk));
	jdff dff_A_dNQgYKEB7_0(.dout(w_dff_A_HZi5PSZl0_0),.din(w_dff_A_dNQgYKEB7_0),.clk(gclk));
	jdff dff_A_HZi5PSZl0_0(.dout(w_dff_A_Y3j9diA04_0),.din(w_dff_A_HZi5PSZl0_0),.clk(gclk));
	jdff dff_A_Y3j9diA04_0(.dout(w_dff_A_tSL6M70X7_0),.din(w_dff_A_Y3j9diA04_0),.clk(gclk));
	jdff dff_A_tSL6M70X7_0(.dout(w_dff_A_KL55QyXJ1_0),.din(w_dff_A_tSL6M70X7_0),.clk(gclk));
	jdff dff_A_KL55QyXJ1_0(.dout(w_dff_A_Svx5lZzP2_0),.din(w_dff_A_KL55QyXJ1_0),.clk(gclk));
	jdff dff_A_Svx5lZzP2_0(.dout(w_dff_A_58pnp1Fr3_0),.din(w_dff_A_Svx5lZzP2_0),.clk(gclk));
	jdff dff_A_58pnp1Fr3_0(.dout(w_dff_A_Qysn4twB7_0),.din(w_dff_A_58pnp1Fr3_0),.clk(gclk));
	jdff dff_A_Qysn4twB7_0(.dout(G615),.din(w_dff_A_Qysn4twB7_0),.clk(gclk));
	jdff dff_A_QmKqJRIv2_2(.dout(w_dff_A_qkdo91Fi2_0),.din(w_dff_A_QmKqJRIv2_2),.clk(gclk));
	jdff dff_A_qkdo91Fi2_0(.dout(w_dff_A_OGCZ5huo7_0),.din(w_dff_A_qkdo91Fi2_0),.clk(gclk));
	jdff dff_A_OGCZ5huo7_0(.dout(w_dff_A_5UvpBk0r5_0),.din(w_dff_A_OGCZ5huo7_0),.clk(gclk));
	jdff dff_A_5UvpBk0r5_0(.dout(w_dff_A_x0JF5A1q7_0),.din(w_dff_A_5UvpBk0r5_0),.clk(gclk));
	jdff dff_A_x0JF5A1q7_0(.dout(w_dff_A_QL1opl1b8_0),.din(w_dff_A_x0JF5A1q7_0),.clk(gclk));
	jdff dff_A_QL1opl1b8_0(.dout(w_dff_A_3OlaC27m3_0),.din(w_dff_A_QL1opl1b8_0),.clk(gclk));
	jdff dff_A_3OlaC27m3_0(.dout(w_dff_A_vVvcsjH78_0),.din(w_dff_A_3OlaC27m3_0),.clk(gclk));
	jdff dff_A_vVvcsjH78_0(.dout(w_dff_A_6eBH2sMQ8_0),.din(w_dff_A_vVvcsjH78_0),.clk(gclk));
	jdff dff_A_6eBH2sMQ8_0(.dout(w_dff_A_0fdM7YKm5_0),.din(w_dff_A_6eBH2sMQ8_0),.clk(gclk));
	jdff dff_A_0fdM7YKm5_0(.dout(w_dff_A_iDGcRBmp4_0),.din(w_dff_A_0fdM7YKm5_0),.clk(gclk));
	jdff dff_A_iDGcRBmp4_0(.dout(w_dff_A_jEyBLj9Q6_0),.din(w_dff_A_iDGcRBmp4_0),.clk(gclk));
	jdff dff_A_jEyBLj9Q6_0(.dout(w_dff_A_pU8QpZRt2_0),.din(w_dff_A_jEyBLj9Q6_0),.clk(gclk));
	jdff dff_A_pU8QpZRt2_0(.dout(w_dff_A_yW1sngvI9_0),.din(w_dff_A_pU8QpZRt2_0),.clk(gclk));
	jdff dff_A_yW1sngvI9_0(.dout(w_dff_A_j1vu3Yto4_0),.din(w_dff_A_yW1sngvI9_0),.clk(gclk));
	jdff dff_A_j1vu3Yto4_0(.dout(w_dff_A_zMkrSvUF8_0),.din(w_dff_A_j1vu3Yto4_0),.clk(gclk));
	jdff dff_A_zMkrSvUF8_0(.dout(w_dff_A_silvTFXx7_0),.din(w_dff_A_zMkrSvUF8_0),.clk(gclk));
	jdff dff_A_silvTFXx7_0(.dout(G626),.din(w_dff_A_silvTFXx7_0),.clk(gclk));
	jdff dff_A_t4OEWpbI4_2(.dout(w_dff_A_XSGwYZJ66_0),.din(w_dff_A_t4OEWpbI4_2),.clk(gclk));
	jdff dff_A_XSGwYZJ66_0(.dout(w_dff_A_qKUKWfzu2_0),.din(w_dff_A_XSGwYZJ66_0),.clk(gclk));
	jdff dff_A_qKUKWfzu2_0(.dout(w_dff_A_qxukhu7v4_0),.din(w_dff_A_qKUKWfzu2_0),.clk(gclk));
	jdff dff_A_qxukhu7v4_0(.dout(w_dff_A_qBLwA6M94_0),.din(w_dff_A_qxukhu7v4_0),.clk(gclk));
	jdff dff_A_qBLwA6M94_0(.dout(w_dff_A_JG0L87Ww6_0),.din(w_dff_A_qBLwA6M94_0),.clk(gclk));
	jdff dff_A_JG0L87Ww6_0(.dout(w_dff_A_2E0x3VZI3_0),.din(w_dff_A_JG0L87Ww6_0),.clk(gclk));
	jdff dff_A_2E0x3VZI3_0(.dout(w_dff_A_fuXWis3a2_0),.din(w_dff_A_2E0x3VZI3_0),.clk(gclk));
	jdff dff_A_fuXWis3a2_0(.dout(w_dff_A_0ReWyaKS8_0),.din(w_dff_A_fuXWis3a2_0),.clk(gclk));
	jdff dff_A_0ReWyaKS8_0(.dout(w_dff_A_fKGZCOfD7_0),.din(w_dff_A_0ReWyaKS8_0),.clk(gclk));
	jdff dff_A_fKGZCOfD7_0(.dout(w_dff_A_PF4yy7YQ5_0),.din(w_dff_A_fKGZCOfD7_0),.clk(gclk));
	jdff dff_A_PF4yy7YQ5_0(.dout(w_dff_A_EPhcu3l71_0),.din(w_dff_A_PF4yy7YQ5_0),.clk(gclk));
	jdff dff_A_EPhcu3l71_0(.dout(w_dff_A_84XnLP5F1_0),.din(w_dff_A_EPhcu3l71_0),.clk(gclk));
	jdff dff_A_84XnLP5F1_0(.dout(w_dff_A_DW0i6k8X9_0),.din(w_dff_A_84XnLP5F1_0),.clk(gclk));
	jdff dff_A_DW0i6k8X9_0(.dout(w_dff_A_Vto4TfUX5_0),.din(w_dff_A_DW0i6k8X9_0),.clk(gclk));
	jdff dff_A_Vto4TfUX5_0(.dout(G632),.din(w_dff_A_Vto4TfUX5_0),.clk(gclk));
	jdff dff_A_8MThqmXy2_1(.dout(w_dff_A_DifVr3Om1_0),.din(w_dff_A_8MThqmXy2_1),.clk(gclk));
	jdff dff_A_DifVr3Om1_0(.dout(w_dff_A_Ng0oECXB3_0),.din(w_dff_A_DifVr3Om1_0),.clk(gclk));
	jdff dff_A_Ng0oECXB3_0(.dout(w_dff_A_l0AW4AGy0_0),.din(w_dff_A_Ng0oECXB3_0),.clk(gclk));
	jdff dff_A_l0AW4AGy0_0(.dout(w_dff_A_mmWYF7Z63_0),.din(w_dff_A_l0AW4AGy0_0),.clk(gclk));
	jdff dff_A_mmWYF7Z63_0(.dout(w_dff_A_G1z6TzYy4_0),.din(w_dff_A_mmWYF7Z63_0),.clk(gclk));
	jdff dff_A_G1z6TzYy4_0(.dout(w_dff_A_z7M6r6dH6_0),.din(w_dff_A_G1z6TzYy4_0),.clk(gclk));
	jdff dff_A_z7M6r6dH6_0(.dout(w_dff_A_ttc7DjDN3_0),.din(w_dff_A_z7M6r6dH6_0),.clk(gclk));
	jdff dff_A_ttc7DjDN3_0(.dout(w_dff_A_njPV4DTd3_0),.din(w_dff_A_ttc7DjDN3_0),.clk(gclk));
	jdff dff_A_njPV4DTd3_0(.dout(w_dff_A_JqmkJdmq5_0),.din(w_dff_A_njPV4DTd3_0),.clk(gclk));
	jdff dff_A_JqmkJdmq5_0(.dout(w_dff_A_2tof4Dml2_0),.din(w_dff_A_JqmkJdmq5_0),.clk(gclk));
	jdff dff_A_2tof4Dml2_0(.dout(w_dff_A_QK0QUSLo3_0),.din(w_dff_A_2tof4Dml2_0),.clk(gclk));
	jdff dff_A_QK0QUSLo3_0(.dout(w_dff_A_W8pZpPQW0_0),.din(w_dff_A_QK0QUSLo3_0),.clk(gclk));
	jdff dff_A_W8pZpPQW0_0(.dout(w_dff_A_hwvb23Lb6_0),.din(w_dff_A_W8pZpPQW0_0),.clk(gclk));
	jdff dff_A_hwvb23Lb6_0(.dout(w_dff_A_7ZzzLzVy7_0),.din(w_dff_A_hwvb23Lb6_0),.clk(gclk));
	jdff dff_A_7ZzzLzVy7_0(.dout(w_dff_A_Y9LsZRIZ3_0),.din(w_dff_A_7ZzzLzVy7_0),.clk(gclk));
	jdff dff_A_Y9LsZRIZ3_0(.dout(w_dff_A_R3Bi5i7L2_0),.din(w_dff_A_Y9LsZRIZ3_0),.clk(gclk));
	jdff dff_A_R3Bi5i7L2_0(.dout(w_dff_A_dJA0b8xC9_0),.din(w_dff_A_R3Bi5i7L2_0),.clk(gclk));
	jdff dff_A_dJA0b8xC9_0(.dout(w_dff_A_Ez533ZU05_0),.din(w_dff_A_dJA0b8xC9_0),.clk(gclk));
	jdff dff_A_Ez533ZU05_0(.dout(w_dff_A_yP86I3PT5_0),.din(w_dff_A_Ez533ZU05_0),.clk(gclk));
	jdff dff_A_yP86I3PT5_0(.dout(w_dff_A_pheM8mO71_0),.din(w_dff_A_yP86I3PT5_0),.clk(gclk));
	jdff dff_A_pheM8mO71_0(.dout(G1002),.din(w_dff_A_pheM8mO71_0),.clk(gclk));
	jdff dff_A_FM7ga7ou8_1(.dout(w_dff_A_liYurLTQ9_0),.din(w_dff_A_FM7ga7ou8_1),.clk(gclk));
	jdff dff_A_liYurLTQ9_0(.dout(w_dff_A_n80DzAQ95_0),.din(w_dff_A_liYurLTQ9_0),.clk(gclk));
	jdff dff_A_n80DzAQ95_0(.dout(w_dff_A_TkSX4e669_0),.din(w_dff_A_n80DzAQ95_0),.clk(gclk));
	jdff dff_A_TkSX4e669_0(.dout(w_dff_A_V1PAS0K72_0),.din(w_dff_A_TkSX4e669_0),.clk(gclk));
	jdff dff_A_V1PAS0K72_0(.dout(w_dff_A_86hg12ZQ9_0),.din(w_dff_A_V1PAS0K72_0),.clk(gclk));
	jdff dff_A_86hg12ZQ9_0(.dout(w_dff_A_zseMmEC93_0),.din(w_dff_A_86hg12ZQ9_0),.clk(gclk));
	jdff dff_A_zseMmEC93_0(.dout(w_dff_A_bYF9qzDW2_0),.din(w_dff_A_zseMmEC93_0),.clk(gclk));
	jdff dff_A_bYF9qzDW2_0(.dout(w_dff_A_ZRANlNYg9_0),.din(w_dff_A_bYF9qzDW2_0),.clk(gclk));
	jdff dff_A_ZRANlNYg9_0(.dout(w_dff_A_IK7n4Vwj6_0),.din(w_dff_A_ZRANlNYg9_0),.clk(gclk));
	jdff dff_A_IK7n4Vwj6_0(.dout(w_dff_A_ttrUmXIN0_0),.din(w_dff_A_IK7n4Vwj6_0),.clk(gclk));
	jdff dff_A_ttrUmXIN0_0(.dout(w_dff_A_UkrFsFir7_0),.din(w_dff_A_ttrUmXIN0_0),.clk(gclk));
	jdff dff_A_UkrFsFir7_0(.dout(w_dff_A_NHS2pa075_0),.din(w_dff_A_UkrFsFir7_0),.clk(gclk));
	jdff dff_A_NHS2pa075_0(.dout(w_dff_A_dxCAVoLL3_0),.din(w_dff_A_NHS2pa075_0),.clk(gclk));
	jdff dff_A_dxCAVoLL3_0(.dout(w_dff_A_Q1qsc3s55_0),.din(w_dff_A_dxCAVoLL3_0),.clk(gclk));
	jdff dff_A_Q1qsc3s55_0(.dout(w_dff_A_4e1Us7Ku2_0),.din(w_dff_A_Q1qsc3s55_0),.clk(gclk));
	jdff dff_A_4e1Us7Ku2_0(.dout(w_dff_A_hfWDkREK5_0),.din(w_dff_A_4e1Us7Ku2_0),.clk(gclk));
	jdff dff_A_hfWDkREK5_0(.dout(w_dff_A_iqOjJnuo3_0),.din(w_dff_A_hfWDkREK5_0),.clk(gclk));
	jdff dff_A_iqOjJnuo3_0(.dout(w_dff_A_ntWxwqQK1_0),.din(w_dff_A_iqOjJnuo3_0),.clk(gclk));
	jdff dff_A_ntWxwqQK1_0(.dout(w_dff_A_2xFGmuuI8_0),.din(w_dff_A_ntWxwqQK1_0),.clk(gclk));
	jdff dff_A_2xFGmuuI8_0(.dout(w_dff_A_JRAIqznC6_0),.din(w_dff_A_2xFGmuuI8_0),.clk(gclk));
	jdff dff_A_JRAIqznC6_0(.dout(G1004),.din(w_dff_A_JRAIqznC6_0),.clk(gclk));
	jdff dff_A_x5Bdeqtt8_2(.dout(w_dff_A_hPhp5Y865_0),.din(w_dff_A_x5Bdeqtt8_2),.clk(gclk));
	jdff dff_A_hPhp5Y865_0(.dout(w_dff_A_b14ek91s8_0),.din(w_dff_A_hPhp5Y865_0),.clk(gclk));
	jdff dff_A_b14ek91s8_0(.dout(w_dff_A_ZfCVIXFP5_0),.din(w_dff_A_b14ek91s8_0),.clk(gclk));
	jdff dff_A_ZfCVIXFP5_0(.dout(w_dff_A_zGLOD5nD8_0),.din(w_dff_A_ZfCVIXFP5_0),.clk(gclk));
	jdff dff_A_zGLOD5nD8_0(.dout(w_dff_A_ANbg6Wwm2_0),.din(w_dff_A_zGLOD5nD8_0),.clk(gclk));
	jdff dff_A_ANbg6Wwm2_0(.dout(w_dff_A_rG5dGwXV3_0),.din(w_dff_A_ANbg6Wwm2_0),.clk(gclk));
	jdff dff_A_rG5dGwXV3_0(.dout(w_dff_A_yI5iJGLK9_0),.din(w_dff_A_rG5dGwXV3_0),.clk(gclk));
	jdff dff_A_yI5iJGLK9_0(.dout(w_dff_A_g6nfOlMj9_0),.din(w_dff_A_yI5iJGLK9_0),.clk(gclk));
	jdff dff_A_g6nfOlMj9_0(.dout(w_dff_A_DemqSCnw7_0),.din(w_dff_A_g6nfOlMj9_0),.clk(gclk));
	jdff dff_A_DemqSCnw7_0(.dout(w_dff_A_VCVhWC6d6_0),.din(w_dff_A_DemqSCnw7_0),.clk(gclk));
	jdff dff_A_VCVhWC6d6_0(.dout(w_dff_A_7iGFQniU7_0),.din(w_dff_A_VCVhWC6d6_0),.clk(gclk));
	jdff dff_A_7iGFQniU7_0(.dout(G591),.din(w_dff_A_7iGFQniU7_0),.clk(gclk));
	jdff dff_A_dUvFZuI17_2(.dout(w_dff_A_XDTo9of91_0),.din(w_dff_A_dUvFZuI17_2),.clk(gclk));
	jdff dff_A_XDTo9of91_0(.dout(w_dff_A_k3CyBxZC2_0),.din(w_dff_A_XDTo9of91_0),.clk(gclk));
	jdff dff_A_k3CyBxZC2_0(.dout(w_dff_A_n1DUMr9q9_0),.din(w_dff_A_k3CyBxZC2_0),.clk(gclk));
	jdff dff_A_n1DUMr9q9_0(.dout(w_dff_A_1TzUogFk7_0),.din(w_dff_A_n1DUMr9q9_0),.clk(gclk));
	jdff dff_A_1TzUogFk7_0(.dout(w_dff_A_1lDnUSeg9_0),.din(w_dff_A_1TzUogFk7_0),.clk(gclk));
	jdff dff_A_1lDnUSeg9_0(.dout(w_dff_A_mGNG4H3s8_0),.din(w_dff_A_1lDnUSeg9_0),.clk(gclk));
	jdff dff_A_mGNG4H3s8_0(.dout(w_dff_A_Y6F9dhiL1_0),.din(w_dff_A_mGNG4H3s8_0),.clk(gclk));
	jdff dff_A_Y6F9dhiL1_0(.dout(w_dff_A_3Br8LzRX7_0),.din(w_dff_A_Y6F9dhiL1_0),.clk(gclk));
	jdff dff_A_3Br8LzRX7_0(.dout(w_dff_A_g7JJJbif9_0),.din(w_dff_A_3Br8LzRX7_0),.clk(gclk));
	jdff dff_A_g7JJJbif9_0(.dout(w_dff_A_9YmxPRjd2_0),.din(w_dff_A_g7JJJbif9_0),.clk(gclk));
	jdff dff_A_9YmxPRjd2_0(.dout(w_dff_A_dVFojz512_0),.din(w_dff_A_9YmxPRjd2_0),.clk(gclk));
	jdff dff_A_dVFojz512_0(.dout(G618),.din(w_dff_A_dVFojz512_0),.clk(gclk));
	jdff dff_A_KD56kTfy9_2(.dout(w_dff_A_d4narGFS4_0),.din(w_dff_A_KD56kTfy9_2),.clk(gclk));
	jdff dff_A_d4narGFS4_0(.dout(w_dff_A_R5rS28be5_0),.din(w_dff_A_d4narGFS4_0),.clk(gclk));
	jdff dff_A_R5rS28be5_0(.dout(w_dff_A_a4yXc90U1_0),.din(w_dff_A_R5rS28be5_0),.clk(gclk));
	jdff dff_A_a4yXc90U1_0(.dout(w_dff_A_x4bT6BTj0_0),.din(w_dff_A_a4yXc90U1_0),.clk(gclk));
	jdff dff_A_x4bT6BTj0_0(.dout(w_dff_A_XVnWRPNy5_0),.din(w_dff_A_x4bT6BTj0_0),.clk(gclk));
	jdff dff_A_XVnWRPNy5_0(.dout(w_dff_A_8vHnto142_0),.din(w_dff_A_XVnWRPNy5_0),.clk(gclk));
	jdff dff_A_8vHnto142_0(.dout(w_dff_A_NkyevxkC1_0),.din(w_dff_A_8vHnto142_0),.clk(gclk));
	jdff dff_A_NkyevxkC1_0(.dout(w_dff_A_i7NRLqUr7_0),.din(w_dff_A_NkyevxkC1_0),.clk(gclk));
	jdff dff_A_i7NRLqUr7_0(.dout(w_dff_A_PkvviMUt2_0),.din(w_dff_A_i7NRLqUr7_0),.clk(gclk));
	jdff dff_A_PkvviMUt2_0(.dout(w_dff_A_YmyiEMt48_0),.din(w_dff_A_PkvviMUt2_0),.clk(gclk));
	jdff dff_A_YmyiEMt48_0(.dout(w_dff_A_YsqjyaXh4_0),.din(w_dff_A_YmyiEMt48_0),.clk(gclk));
	jdff dff_A_YsqjyaXh4_0(.dout(G621),.din(w_dff_A_YsqjyaXh4_0),.clk(gclk));
	jdff dff_A_Cy9lkNbV7_2(.dout(w_dff_A_NhrnOveV2_0),.din(w_dff_A_Cy9lkNbV7_2),.clk(gclk));
	jdff dff_A_NhrnOveV2_0(.dout(w_dff_A_7Yvj5zxD4_0),.din(w_dff_A_NhrnOveV2_0),.clk(gclk));
	jdff dff_A_7Yvj5zxD4_0(.dout(w_dff_A_X3xuNiyw9_0),.din(w_dff_A_7Yvj5zxD4_0),.clk(gclk));
	jdff dff_A_X3xuNiyw9_0(.dout(w_dff_A_Qvyp2K459_0),.din(w_dff_A_X3xuNiyw9_0),.clk(gclk));
	jdff dff_A_Qvyp2K459_0(.dout(w_dff_A_c7vrLhPU0_0),.din(w_dff_A_Qvyp2K459_0),.clk(gclk));
	jdff dff_A_c7vrLhPU0_0(.dout(w_dff_A_sUSzQodi5_0),.din(w_dff_A_c7vrLhPU0_0),.clk(gclk));
	jdff dff_A_sUSzQodi5_0(.dout(w_dff_A_uPhWfkZE8_0),.din(w_dff_A_sUSzQodi5_0),.clk(gclk));
	jdff dff_A_uPhWfkZE8_0(.dout(w_dff_A_2NiPPrNn4_0),.din(w_dff_A_uPhWfkZE8_0),.clk(gclk));
	jdff dff_A_2NiPPrNn4_0(.dout(w_dff_A_XryDxHHc7_0),.din(w_dff_A_2NiPPrNn4_0),.clk(gclk));
	jdff dff_A_XryDxHHc7_0(.dout(w_dff_A_b0E8rjz12_0),.din(w_dff_A_XryDxHHc7_0),.clk(gclk));
	jdff dff_A_b0E8rjz12_0(.dout(w_dff_A_cZ9PTVaY6_0),.din(w_dff_A_b0E8rjz12_0),.clk(gclk));
	jdff dff_A_cZ9PTVaY6_0(.dout(G629),.din(w_dff_A_cZ9PTVaY6_0),.clk(gclk));
	jdff dff_A_snZJi9ST6_1(.dout(w_dff_A_aq8I2DKO3_0),.din(w_dff_A_snZJi9ST6_1),.clk(gclk));
	jdff dff_A_aq8I2DKO3_0(.dout(w_dff_A_7cy1O96o3_0),.din(w_dff_A_aq8I2DKO3_0),.clk(gclk));
	jdff dff_A_7cy1O96o3_0(.dout(w_dff_A_IOaltbKl6_0),.din(w_dff_A_7cy1O96o3_0),.clk(gclk));
	jdff dff_A_IOaltbKl6_0(.dout(w_dff_A_EMmGKFik4_0),.din(w_dff_A_IOaltbKl6_0),.clk(gclk));
	jdff dff_A_EMmGKFik4_0(.dout(w_dff_A_nz9wzjG16_0),.din(w_dff_A_EMmGKFik4_0),.clk(gclk));
	jdff dff_A_nz9wzjG16_0(.dout(w_dff_A_X8V0nYfi7_0),.din(w_dff_A_nz9wzjG16_0),.clk(gclk));
	jdff dff_A_X8V0nYfi7_0(.dout(w_dff_A_TajhmYGg3_0),.din(w_dff_A_X8V0nYfi7_0),.clk(gclk));
	jdff dff_A_TajhmYGg3_0(.dout(w_dff_A_Y0a6UnnT6_0),.din(w_dff_A_TajhmYGg3_0),.clk(gclk));
	jdff dff_A_Y0a6UnnT6_0(.dout(w_dff_A_ao25x0TM2_0),.din(w_dff_A_Y0a6UnnT6_0),.clk(gclk));
	jdff dff_A_ao25x0TM2_0(.dout(w_dff_A_yASrjxQ85_0),.din(w_dff_A_ao25x0TM2_0),.clk(gclk));
	jdff dff_A_yASrjxQ85_0(.dout(w_dff_A_7qI3Ea5C9_0),.din(w_dff_A_yASrjxQ85_0),.clk(gclk));
	jdff dff_A_7qI3Ea5C9_0(.dout(w_dff_A_9tdBiNxn1_0),.din(w_dff_A_7qI3Ea5C9_0),.clk(gclk));
	jdff dff_A_9tdBiNxn1_0(.dout(w_dff_A_4pz3WHHu2_0),.din(w_dff_A_9tdBiNxn1_0),.clk(gclk));
	jdff dff_A_4pz3WHHu2_0(.dout(w_dff_A_q7fYNNpk5_0),.din(w_dff_A_4pz3WHHu2_0),.clk(gclk));
	jdff dff_A_q7fYNNpk5_0(.dout(w_dff_A_VFHKjjf15_0),.din(w_dff_A_q7fYNNpk5_0),.clk(gclk));
	jdff dff_A_VFHKjjf15_0(.dout(w_dff_A_iRbCYIBv5_0),.din(w_dff_A_VFHKjjf15_0),.clk(gclk));
	jdff dff_A_iRbCYIBv5_0(.dout(w_dff_A_NoqhdNf00_0),.din(w_dff_A_iRbCYIBv5_0),.clk(gclk));
	jdff dff_A_NoqhdNf00_0(.dout(w_dff_A_DEjCMjYR1_0),.din(w_dff_A_NoqhdNf00_0),.clk(gclk));
	jdff dff_A_DEjCMjYR1_0(.dout(G822),.din(w_dff_A_DEjCMjYR1_0),.clk(gclk));
	jdff dff_A_NU9RSijT7_1(.dout(w_dff_A_Ep3zLD1i4_0),.din(w_dff_A_NU9RSijT7_1),.clk(gclk));
	jdff dff_A_Ep3zLD1i4_0(.dout(w_dff_A_Ybo5zWwy2_0),.din(w_dff_A_Ep3zLD1i4_0),.clk(gclk));
	jdff dff_A_Ybo5zWwy2_0(.dout(w_dff_A_isKRucTK0_0),.din(w_dff_A_Ybo5zWwy2_0),.clk(gclk));
	jdff dff_A_isKRucTK0_0(.dout(w_dff_A_QAWQtNTc2_0),.din(w_dff_A_isKRucTK0_0),.clk(gclk));
	jdff dff_A_QAWQtNTc2_0(.dout(w_dff_A_Uw61XWbZ4_0),.din(w_dff_A_QAWQtNTc2_0),.clk(gclk));
	jdff dff_A_Uw61XWbZ4_0(.dout(w_dff_A_2OaVpKAG8_0),.din(w_dff_A_Uw61XWbZ4_0),.clk(gclk));
	jdff dff_A_2OaVpKAG8_0(.dout(w_dff_A_E8YSR3hE2_0),.din(w_dff_A_2OaVpKAG8_0),.clk(gclk));
	jdff dff_A_E8YSR3hE2_0(.dout(w_dff_A_1vQVqcdV0_0),.din(w_dff_A_E8YSR3hE2_0),.clk(gclk));
	jdff dff_A_1vQVqcdV0_0(.dout(w_dff_A_E420atvZ0_0),.din(w_dff_A_1vQVqcdV0_0),.clk(gclk));
	jdff dff_A_E420atvZ0_0(.dout(w_dff_A_lO8HBcVh6_0),.din(w_dff_A_E420atvZ0_0),.clk(gclk));
	jdff dff_A_lO8HBcVh6_0(.dout(w_dff_A_CC1DrSrT2_0),.din(w_dff_A_lO8HBcVh6_0),.clk(gclk));
	jdff dff_A_CC1DrSrT2_0(.dout(w_dff_A_kkH6UtBj1_0),.din(w_dff_A_CC1DrSrT2_0),.clk(gclk));
	jdff dff_A_kkH6UtBj1_0(.dout(w_dff_A_vOZGE8vc3_0),.din(w_dff_A_kkH6UtBj1_0),.clk(gclk));
	jdff dff_A_vOZGE8vc3_0(.dout(w_dff_A_lqf1ogiV1_0),.din(w_dff_A_vOZGE8vc3_0),.clk(gclk));
	jdff dff_A_lqf1ogiV1_0(.dout(w_dff_A_k1dgeqFz8_0),.din(w_dff_A_lqf1ogiV1_0),.clk(gclk));
	jdff dff_A_k1dgeqFz8_0(.dout(w_dff_A_0NMOQF9m1_0),.din(w_dff_A_k1dgeqFz8_0),.clk(gclk));
	jdff dff_A_0NMOQF9m1_0(.dout(w_dff_A_wVNaNbx41_0),.din(w_dff_A_0NMOQF9m1_0),.clk(gclk));
	jdff dff_A_wVNaNbx41_0(.dout(G838),.din(w_dff_A_wVNaNbx41_0),.clk(gclk));
	jdff dff_A_ZXolT0V26_1(.dout(w_dff_A_ZZq4kYo64_0),.din(w_dff_A_ZXolT0V26_1),.clk(gclk));
	jdff dff_A_ZZq4kYo64_0(.dout(w_dff_A_kldSVPQ84_0),.din(w_dff_A_ZZq4kYo64_0),.clk(gclk));
	jdff dff_A_kldSVPQ84_0(.dout(w_dff_A_kqFFAjy18_0),.din(w_dff_A_kldSVPQ84_0),.clk(gclk));
	jdff dff_A_kqFFAjy18_0(.dout(w_dff_A_df8MVVbc5_0),.din(w_dff_A_kqFFAjy18_0),.clk(gclk));
	jdff dff_A_df8MVVbc5_0(.dout(w_dff_A_gjHY7BFg2_0),.din(w_dff_A_df8MVVbc5_0),.clk(gclk));
	jdff dff_A_gjHY7BFg2_0(.dout(w_dff_A_N1YpechW1_0),.din(w_dff_A_gjHY7BFg2_0),.clk(gclk));
	jdff dff_A_N1YpechW1_0(.dout(w_dff_A_Xs2t9kTr4_0),.din(w_dff_A_N1YpechW1_0),.clk(gclk));
	jdff dff_A_Xs2t9kTr4_0(.dout(w_dff_A_JN19R1lq1_0),.din(w_dff_A_Xs2t9kTr4_0),.clk(gclk));
	jdff dff_A_JN19R1lq1_0(.dout(w_dff_A_v9VaeYR98_0),.din(w_dff_A_JN19R1lq1_0),.clk(gclk));
	jdff dff_A_v9VaeYR98_0(.dout(w_dff_A_2WGcBnbR7_0),.din(w_dff_A_v9VaeYR98_0),.clk(gclk));
	jdff dff_A_2WGcBnbR7_0(.dout(w_dff_A_ipFZ34Lt1_0),.din(w_dff_A_2WGcBnbR7_0),.clk(gclk));
	jdff dff_A_ipFZ34Lt1_0(.dout(w_dff_A_iTZPwjIH7_0),.din(w_dff_A_ipFZ34Lt1_0),.clk(gclk));
	jdff dff_A_iTZPwjIH7_0(.dout(w_dff_A_kXYckNTh4_0),.din(w_dff_A_iTZPwjIH7_0),.clk(gclk));
	jdff dff_A_kXYckNTh4_0(.dout(w_dff_A_gww8E7655_0),.din(w_dff_A_kXYckNTh4_0),.clk(gclk));
	jdff dff_A_gww8E7655_0(.dout(w_dff_A_oOE0Yfsj3_0),.din(w_dff_A_gww8E7655_0),.clk(gclk));
	jdff dff_A_oOE0Yfsj3_0(.dout(w_dff_A_ya5AUVCw8_0),.din(w_dff_A_oOE0Yfsj3_0),.clk(gclk));
	jdff dff_A_ya5AUVCw8_0(.dout(w_dff_A_hTLAoxsz8_0),.din(w_dff_A_ya5AUVCw8_0),.clk(gclk));
	jdff dff_A_hTLAoxsz8_0(.dout(G861),.din(w_dff_A_hTLAoxsz8_0),.clk(gclk));
	jdff dff_A_ThmdqykU8_1(.dout(w_dff_A_dh5p1ikk2_0),.din(w_dff_A_ThmdqykU8_1),.clk(gclk));
	jdff dff_A_dh5p1ikk2_0(.dout(w_dff_A_pEqBSy1B5_0),.din(w_dff_A_dh5p1ikk2_0),.clk(gclk));
	jdff dff_A_pEqBSy1B5_0(.dout(w_dff_A_vGTJbVse1_0),.din(w_dff_A_pEqBSy1B5_0),.clk(gclk));
	jdff dff_A_vGTJbVse1_0(.dout(w_dff_A_MhaL0zvK2_0),.din(w_dff_A_vGTJbVse1_0),.clk(gclk));
	jdff dff_A_MhaL0zvK2_0(.dout(w_dff_A_3tpwft3G5_0),.din(w_dff_A_MhaL0zvK2_0),.clk(gclk));
	jdff dff_A_3tpwft3G5_0(.dout(w_dff_A_VkYGSsx51_0),.din(w_dff_A_3tpwft3G5_0),.clk(gclk));
	jdff dff_A_VkYGSsx51_0(.dout(G623),.din(w_dff_A_VkYGSsx51_0),.clk(gclk));
	jdff dff_A_ZHMTSP3i6_2(.dout(w_dff_A_V4EC7Dd53_0),.din(w_dff_A_ZHMTSP3i6_2),.clk(gclk));
	jdff dff_A_V4EC7Dd53_0(.dout(w_dff_A_aYgdNbkN9_0),.din(w_dff_A_V4EC7Dd53_0),.clk(gclk));
	jdff dff_A_aYgdNbkN9_0(.dout(w_dff_A_UNBiD9eu9_0),.din(w_dff_A_aYgdNbkN9_0),.clk(gclk));
	jdff dff_A_UNBiD9eu9_0(.dout(w_dff_A_9oNu4w210_0),.din(w_dff_A_UNBiD9eu9_0),.clk(gclk));
	jdff dff_A_9oNu4w210_0(.dout(w_dff_A_h3ZyZ3hk0_0),.din(w_dff_A_9oNu4w210_0),.clk(gclk));
	jdff dff_A_h3ZyZ3hk0_0(.dout(w_dff_A_umIRhdYr8_0),.din(w_dff_A_h3ZyZ3hk0_0),.clk(gclk));
	jdff dff_A_umIRhdYr8_0(.dout(w_dff_A_cKv4AR9w0_0),.din(w_dff_A_umIRhdYr8_0),.clk(gclk));
	jdff dff_A_cKv4AR9w0_0(.dout(w_dff_A_jMxXD8LX8_0),.din(w_dff_A_cKv4AR9w0_0),.clk(gclk));
	jdff dff_A_jMxXD8LX8_0(.dout(w_dff_A_7d04FC6Z1_0),.din(w_dff_A_jMxXD8LX8_0),.clk(gclk));
	jdff dff_A_7d04FC6Z1_0(.dout(w_dff_A_CQB6sj5B2_0),.din(w_dff_A_7d04FC6Z1_0),.clk(gclk));
	jdff dff_A_CQB6sj5B2_0(.dout(w_dff_A_VvWL19su1_0),.din(w_dff_A_CQB6sj5B2_0),.clk(gclk));
	jdff dff_A_VvWL19su1_0(.dout(w_dff_A_UOiucRSY6_0),.din(w_dff_A_VvWL19su1_0),.clk(gclk));
	jdff dff_A_UOiucRSY6_0(.dout(w_dff_A_br8hVELs5_0),.din(w_dff_A_UOiucRSY6_0),.clk(gclk));
	jdff dff_A_br8hVELs5_0(.dout(w_dff_A_IbBxoM2o5_0),.din(w_dff_A_br8hVELs5_0),.clk(gclk));
	jdff dff_A_IbBxoM2o5_0(.dout(G722),.din(w_dff_A_IbBxoM2o5_0),.clk(gclk));
	jdff dff_A_wR17c80c2_1(.dout(w_dff_A_XfJEjMF64_0),.din(w_dff_A_wR17c80c2_1),.clk(gclk));
	jdff dff_A_XfJEjMF64_0(.dout(w_dff_A_og1H0ZN97_0),.din(w_dff_A_XfJEjMF64_0),.clk(gclk));
	jdff dff_A_og1H0ZN97_0(.dout(w_dff_A_SM2wA2Wy3_0),.din(w_dff_A_og1H0ZN97_0),.clk(gclk));
	jdff dff_A_SM2wA2Wy3_0(.dout(w_dff_A_MUGDUylO6_0),.din(w_dff_A_SM2wA2Wy3_0),.clk(gclk));
	jdff dff_A_MUGDUylO6_0(.dout(w_dff_A_bBuWOqqy7_0),.din(w_dff_A_MUGDUylO6_0),.clk(gclk));
	jdff dff_A_bBuWOqqy7_0(.dout(w_dff_A_c2vFd4CO8_0),.din(w_dff_A_bBuWOqqy7_0),.clk(gclk));
	jdff dff_A_c2vFd4CO8_0(.dout(w_dff_A_PSykAM4I7_0),.din(w_dff_A_c2vFd4CO8_0),.clk(gclk));
	jdff dff_A_PSykAM4I7_0(.dout(w_dff_A_bkq4kN653_0),.din(w_dff_A_PSykAM4I7_0),.clk(gclk));
	jdff dff_A_bkq4kN653_0(.dout(w_dff_A_rB5l1Dxt4_0),.din(w_dff_A_bkq4kN653_0),.clk(gclk));
	jdff dff_A_rB5l1Dxt4_0(.dout(w_dff_A_7WDLAm422_0),.din(w_dff_A_rB5l1Dxt4_0),.clk(gclk));
	jdff dff_A_7WDLAm422_0(.dout(w_dff_A_FdOzntpk3_0),.din(w_dff_A_7WDLAm422_0),.clk(gclk));
	jdff dff_A_FdOzntpk3_0(.dout(G832),.din(w_dff_A_FdOzntpk3_0),.clk(gclk));
	jdff dff_A_5Xx6TgKH7_1(.dout(w_dff_A_lMOqQ0rS8_0),.din(w_dff_A_5Xx6TgKH7_1),.clk(gclk));
	jdff dff_A_lMOqQ0rS8_0(.dout(w_dff_A_t7z3xsnm6_0),.din(w_dff_A_lMOqQ0rS8_0),.clk(gclk));
	jdff dff_A_t7z3xsnm6_0(.dout(w_dff_A_OetBEDxM9_0),.din(w_dff_A_t7z3xsnm6_0),.clk(gclk));
	jdff dff_A_OetBEDxM9_0(.dout(w_dff_A_icOXVjl64_0),.din(w_dff_A_OetBEDxM9_0),.clk(gclk));
	jdff dff_A_icOXVjl64_0(.dout(w_dff_A_shiYJbDp9_0),.din(w_dff_A_icOXVjl64_0),.clk(gclk));
	jdff dff_A_shiYJbDp9_0(.dout(w_dff_A_rAXf54PX9_0),.din(w_dff_A_shiYJbDp9_0),.clk(gclk));
	jdff dff_A_rAXf54PX9_0(.dout(w_dff_A_Jg4vQ9HV2_0),.din(w_dff_A_rAXf54PX9_0),.clk(gclk));
	jdff dff_A_Jg4vQ9HV2_0(.dout(w_dff_A_WcamD9mg6_0),.din(w_dff_A_Jg4vQ9HV2_0),.clk(gclk));
	jdff dff_A_WcamD9mg6_0(.dout(w_dff_A_JuZhTEyw5_0),.din(w_dff_A_WcamD9mg6_0),.clk(gclk));
	jdff dff_A_JuZhTEyw5_0(.dout(w_dff_A_goRRc3wp5_0),.din(w_dff_A_JuZhTEyw5_0),.clk(gclk));
	jdff dff_A_goRRc3wp5_0(.dout(w_dff_A_DDmMEMTW2_0),.din(w_dff_A_goRRc3wp5_0),.clk(gclk));
	jdff dff_A_DDmMEMTW2_0(.dout(w_dff_A_8MZY8CUr4_0),.din(w_dff_A_DDmMEMTW2_0),.clk(gclk));
	jdff dff_A_8MZY8CUr4_0(.dout(w_dff_A_AA3ph8CU2_0),.din(w_dff_A_8MZY8CUr4_0),.clk(gclk));
	jdff dff_A_AA3ph8CU2_0(.dout(G834),.din(w_dff_A_AA3ph8CU2_0),.clk(gclk));
	jdff dff_A_qqGvtkqc6_1(.dout(w_dff_A_qGoG3T8h0_0),.din(w_dff_A_qqGvtkqc6_1),.clk(gclk));
	jdff dff_A_qGoG3T8h0_0(.dout(w_dff_A_Ii5ZwzAM5_0),.din(w_dff_A_qGoG3T8h0_0),.clk(gclk));
	jdff dff_A_Ii5ZwzAM5_0(.dout(w_dff_A_ybg4YFsM6_0),.din(w_dff_A_Ii5ZwzAM5_0),.clk(gclk));
	jdff dff_A_ybg4YFsM6_0(.dout(w_dff_A_PWBe3cmi9_0),.din(w_dff_A_ybg4YFsM6_0),.clk(gclk));
	jdff dff_A_PWBe3cmi9_0(.dout(w_dff_A_9jv2sYF36_0),.din(w_dff_A_PWBe3cmi9_0),.clk(gclk));
	jdff dff_A_9jv2sYF36_0(.dout(w_dff_A_18j6Fyyx0_0),.din(w_dff_A_9jv2sYF36_0),.clk(gclk));
	jdff dff_A_18j6Fyyx0_0(.dout(w_dff_A_389TtBxd9_0),.din(w_dff_A_18j6Fyyx0_0),.clk(gclk));
	jdff dff_A_389TtBxd9_0(.dout(w_dff_A_2IXg8DsH0_0),.din(w_dff_A_389TtBxd9_0),.clk(gclk));
	jdff dff_A_2IXg8DsH0_0(.dout(w_dff_A_oXW4n89S0_0),.din(w_dff_A_2IXg8DsH0_0),.clk(gclk));
	jdff dff_A_oXW4n89S0_0(.dout(w_dff_A_LqJlf77v3_0),.din(w_dff_A_oXW4n89S0_0),.clk(gclk));
	jdff dff_A_LqJlf77v3_0(.dout(w_dff_A_SBVJSIm32_0),.din(w_dff_A_LqJlf77v3_0),.clk(gclk));
	jdff dff_A_SBVJSIm32_0(.dout(w_dff_A_0ulM0GLY8_0),.din(w_dff_A_SBVJSIm32_0),.clk(gclk));
	jdff dff_A_0ulM0GLY8_0(.dout(w_dff_A_jPf8QPi70_0),.din(w_dff_A_0ulM0GLY8_0),.clk(gclk));
	jdff dff_A_jPf8QPi70_0(.dout(w_dff_A_NzPM8eWl4_0),.din(w_dff_A_jPf8QPi70_0),.clk(gclk));
	jdff dff_A_NzPM8eWl4_0(.dout(w_dff_A_r7DH87ma9_0),.din(w_dff_A_NzPM8eWl4_0),.clk(gclk));
	jdff dff_A_r7DH87ma9_0(.dout(G836),.din(w_dff_A_r7DH87ma9_0),.clk(gclk));
	jdff dff_A_7O2wzkaw1_2(.dout(w_dff_A_ilQmmqJD0_0),.din(w_dff_A_7O2wzkaw1_2),.clk(gclk));
	jdff dff_A_ilQmmqJD0_0(.dout(w_dff_A_IYtFxu9W0_0),.din(w_dff_A_ilQmmqJD0_0),.clk(gclk));
	jdff dff_A_IYtFxu9W0_0(.dout(w_dff_A_e2k2DRdl7_0),.din(w_dff_A_IYtFxu9W0_0),.clk(gclk));
	jdff dff_A_e2k2DRdl7_0(.dout(w_dff_A_WeGYUlUa8_0),.din(w_dff_A_e2k2DRdl7_0),.clk(gclk));
	jdff dff_A_WeGYUlUa8_0(.dout(w_dff_A_cr3jm7j96_0),.din(w_dff_A_WeGYUlUa8_0),.clk(gclk));
	jdff dff_A_cr3jm7j96_0(.dout(w_dff_A_WFMfEKIz5_0),.din(w_dff_A_cr3jm7j96_0),.clk(gclk));
	jdff dff_A_WFMfEKIz5_0(.dout(w_dff_A_6Etd3qUY3_0),.din(w_dff_A_WFMfEKIz5_0),.clk(gclk));
	jdff dff_A_6Etd3qUY3_0(.dout(w_dff_A_BHu1VUKb9_0),.din(w_dff_A_6Etd3qUY3_0),.clk(gclk));
	jdff dff_A_BHu1VUKb9_0(.dout(w_dff_A_yykVMFx44_0),.din(w_dff_A_BHu1VUKb9_0),.clk(gclk));
	jdff dff_A_yykVMFx44_0(.dout(w_dff_A_rarOqqIw2_0),.din(w_dff_A_yykVMFx44_0),.clk(gclk));
	jdff dff_A_rarOqqIw2_0(.dout(w_dff_A_h2U5pKVg1_0),.din(w_dff_A_rarOqqIw2_0),.clk(gclk));
	jdff dff_A_h2U5pKVg1_0(.dout(w_dff_A_pbVMcsM92_0),.din(w_dff_A_h2U5pKVg1_0),.clk(gclk));
	jdff dff_A_pbVMcsM92_0(.dout(w_dff_A_MuzgbhDl3_0),.din(w_dff_A_pbVMcsM92_0),.clk(gclk));
	jdff dff_A_MuzgbhDl3_0(.dout(w_dff_A_1jIKfZT23_0),.din(w_dff_A_MuzgbhDl3_0),.clk(gclk));
	jdff dff_A_1jIKfZT23_0(.dout(G859),.din(w_dff_A_1jIKfZT23_0),.clk(gclk));
	jdff dff_A_N7LHGUu06_1(.dout(w_dff_A_Uqa9WElK9_0),.din(w_dff_A_N7LHGUu06_1),.clk(gclk));
	jdff dff_A_Uqa9WElK9_0(.dout(w_dff_A_drEy0vdf7_0),.din(w_dff_A_Uqa9WElK9_0),.clk(gclk));
	jdff dff_A_drEy0vdf7_0(.dout(w_dff_A_vCOILdJZ5_0),.din(w_dff_A_drEy0vdf7_0),.clk(gclk));
	jdff dff_A_vCOILdJZ5_0(.dout(w_dff_A_RV1WwCaw6_0),.din(w_dff_A_vCOILdJZ5_0),.clk(gclk));
	jdff dff_A_RV1WwCaw6_0(.dout(w_dff_A_ISZ4NYmR7_0),.din(w_dff_A_RV1WwCaw6_0),.clk(gclk));
	jdff dff_A_ISZ4NYmR7_0(.dout(w_dff_A_Hpj30Ax63_0),.din(w_dff_A_ISZ4NYmR7_0),.clk(gclk));
	jdff dff_A_Hpj30Ax63_0(.dout(w_dff_A_mFOiPj4c2_0),.din(w_dff_A_Hpj30Ax63_0),.clk(gclk));
	jdff dff_A_mFOiPj4c2_0(.dout(w_dff_A_ppkBLltQ7_0),.din(w_dff_A_mFOiPj4c2_0),.clk(gclk));
	jdff dff_A_ppkBLltQ7_0(.dout(w_dff_A_dPMgjU3R7_0),.din(w_dff_A_ppkBLltQ7_0),.clk(gclk));
	jdff dff_A_dPMgjU3R7_0(.dout(G871),.din(w_dff_A_dPMgjU3R7_0),.clk(gclk));
	jdff dff_A_Z21vggDg8_1(.dout(w_dff_A_c64wwYKJ4_0),.din(w_dff_A_Z21vggDg8_1),.clk(gclk));
	jdff dff_A_c64wwYKJ4_0(.dout(w_dff_A_ypNE6hvh7_0),.din(w_dff_A_c64wwYKJ4_0),.clk(gclk));
	jdff dff_A_ypNE6hvh7_0(.dout(w_dff_A_CvZYO3aI0_0),.din(w_dff_A_ypNE6hvh7_0),.clk(gclk));
	jdff dff_A_CvZYO3aI0_0(.dout(w_dff_A_g94nGanx7_0),.din(w_dff_A_CvZYO3aI0_0),.clk(gclk));
	jdff dff_A_g94nGanx7_0(.dout(w_dff_A_p1vJkx1M8_0),.din(w_dff_A_g94nGanx7_0),.clk(gclk));
	jdff dff_A_p1vJkx1M8_0(.dout(w_dff_A_A7pY0dpX1_0),.din(w_dff_A_p1vJkx1M8_0),.clk(gclk));
	jdff dff_A_A7pY0dpX1_0(.dout(w_dff_A_hYyeh1fV6_0),.din(w_dff_A_A7pY0dpX1_0),.clk(gclk));
	jdff dff_A_hYyeh1fV6_0(.dout(w_dff_A_ZAVSQPGH8_0),.din(w_dff_A_hYyeh1fV6_0),.clk(gclk));
	jdff dff_A_ZAVSQPGH8_0(.dout(w_dff_A_p11MuTuQ9_0),.din(w_dff_A_ZAVSQPGH8_0),.clk(gclk));
	jdff dff_A_p11MuTuQ9_0(.dout(w_dff_A_PZOjwCQ04_0),.din(w_dff_A_p11MuTuQ9_0),.clk(gclk));
	jdff dff_A_PZOjwCQ04_0(.dout(w_dff_A_hq6ePeyd7_0),.din(w_dff_A_PZOjwCQ04_0),.clk(gclk));
	jdff dff_A_hq6ePeyd7_0(.dout(G873),.din(w_dff_A_hq6ePeyd7_0),.clk(gclk));
	jdff dff_A_5zsUPBA47_1(.dout(w_dff_A_VYoBtlWz3_0),.din(w_dff_A_5zsUPBA47_1),.clk(gclk));
	jdff dff_A_VYoBtlWz3_0(.dout(w_dff_A_RkhlHoH04_0),.din(w_dff_A_VYoBtlWz3_0),.clk(gclk));
	jdff dff_A_RkhlHoH04_0(.dout(w_dff_A_m9DOy8Tk0_0),.din(w_dff_A_RkhlHoH04_0),.clk(gclk));
	jdff dff_A_m9DOy8Tk0_0(.dout(w_dff_A_U50f7xEO2_0),.din(w_dff_A_m9DOy8Tk0_0),.clk(gclk));
	jdff dff_A_U50f7xEO2_0(.dout(w_dff_A_pgJa7A665_0),.din(w_dff_A_U50f7xEO2_0),.clk(gclk));
	jdff dff_A_pgJa7A665_0(.dout(w_dff_A_93DO8Yf21_0),.din(w_dff_A_pgJa7A665_0),.clk(gclk));
	jdff dff_A_93DO8Yf21_0(.dout(w_dff_A_jwa96Fl75_0),.din(w_dff_A_93DO8Yf21_0),.clk(gclk));
	jdff dff_A_jwa96Fl75_0(.dout(w_dff_A_HnAfBtkG4_0),.din(w_dff_A_jwa96Fl75_0),.clk(gclk));
	jdff dff_A_HnAfBtkG4_0(.dout(w_dff_A_Fulb2dLV5_0),.din(w_dff_A_HnAfBtkG4_0),.clk(gclk));
	jdff dff_A_Fulb2dLV5_0(.dout(w_dff_A_Zp2sodSg8_0),.din(w_dff_A_Fulb2dLV5_0),.clk(gclk));
	jdff dff_A_Zp2sodSg8_0(.dout(w_dff_A_6hDRUkCX4_0),.din(w_dff_A_Zp2sodSg8_0),.clk(gclk));
	jdff dff_A_6hDRUkCX4_0(.dout(w_dff_A_Q01r9AYR6_0),.din(w_dff_A_6hDRUkCX4_0),.clk(gclk));
	jdff dff_A_Q01r9AYR6_0(.dout(G875),.din(w_dff_A_Q01r9AYR6_0),.clk(gclk));
	jdff dff_A_M2r8JevI0_1(.dout(w_dff_A_4NKiSx5A2_0),.din(w_dff_A_M2r8JevI0_1),.clk(gclk));
	jdff dff_A_4NKiSx5A2_0(.dout(w_dff_A_VWi6s1Jw2_0),.din(w_dff_A_4NKiSx5A2_0),.clk(gclk));
	jdff dff_A_VWi6s1Jw2_0(.dout(w_dff_A_podGFzGD8_0),.din(w_dff_A_VWi6s1Jw2_0),.clk(gclk));
	jdff dff_A_podGFzGD8_0(.dout(w_dff_A_dBpxepUG6_0),.din(w_dff_A_podGFzGD8_0),.clk(gclk));
	jdff dff_A_dBpxepUG6_0(.dout(w_dff_A_k5ZtWuAc5_0),.din(w_dff_A_dBpxepUG6_0),.clk(gclk));
	jdff dff_A_k5ZtWuAc5_0(.dout(w_dff_A_ODIXZ89F6_0),.din(w_dff_A_k5ZtWuAc5_0),.clk(gclk));
	jdff dff_A_ODIXZ89F6_0(.dout(w_dff_A_JAenVpx02_0),.din(w_dff_A_ODIXZ89F6_0),.clk(gclk));
	jdff dff_A_JAenVpx02_0(.dout(w_dff_A_IHvtxObP5_0),.din(w_dff_A_JAenVpx02_0),.clk(gclk));
	jdff dff_A_IHvtxObP5_0(.dout(w_dff_A_bMf3h5LL5_0),.din(w_dff_A_IHvtxObP5_0),.clk(gclk));
	jdff dff_A_bMf3h5LL5_0(.dout(w_dff_A_b4ooQjrS2_0),.din(w_dff_A_bMf3h5LL5_0),.clk(gclk));
	jdff dff_A_b4ooQjrS2_0(.dout(w_dff_A_gUT7qUu26_0),.din(w_dff_A_b4ooQjrS2_0),.clk(gclk));
	jdff dff_A_gUT7qUu26_0(.dout(w_dff_A_ufoCXX3U0_0),.din(w_dff_A_gUT7qUu26_0),.clk(gclk));
	jdff dff_A_ufoCXX3U0_0(.dout(w_dff_A_3QUBX8Qt3_0),.din(w_dff_A_ufoCXX3U0_0),.clk(gclk));
	jdff dff_A_3QUBX8Qt3_0(.dout(G877),.din(w_dff_A_3QUBX8Qt3_0),.clk(gclk));
	jdff dff_A_rsHUFwPC0_1(.dout(w_dff_A_T9asdqcq4_0),.din(w_dff_A_rsHUFwPC0_1),.clk(gclk));
	jdff dff_A_T9asdqcq4_0(.dout(w_dff_A_ixcoWCSO2_0),.din(w_dff_A_T9asdqcq4_0),.clk(gclk));
	jdff dff_A_ixcoWCSO2_0(.dout(w_dff_A_PtOWfpMy2_0),.din(w_dff_A_ixcoWCSO2_0),.clk(gclk));
	jdff dff_A_PtOWfpMy2_0(.dout(w_dff_A_DBRdP60S9_0),.din(w_dff_A_PtOWfpMy2_0),.clk(gclk));
	jdff dff_A_DBRdP60S9_0(.dout(w_dff_A_Yc6tf6mU9_0),.din(w_dff_A_DBRdP60S9_0),.clk(gclk));
	jdff dff_A_Yc6tf6mU9_0(.dout(w_dff_A_tMCRbGHo2_0),.din(w_dff_A_Yc6tf6mU9_0),.clk(gclk));
	jdff dff_A_tMCRbGHo2_0(.dout(w_dff_A_rz5qe9ya3_0),.din(w_dff_A_tMCRbGHo2_0),.clk(gclk));
	jdff dff_A_rz5qe9ya3_0(.dout(w_dff_A_x6hpU3qV9_0),.din(w_dff_A_rz5qe9ya3_0),.clk(gclk));
	jdff dff_A_x6hpU3qV9_0(.dout(w_dff_A_CAcrCyCy6_0),.din(w_dff_A_x6hpU3qV9_0),.clk(gclk));
	jdff dff_A_CAcrCyCy6_0(.dout(w_dff_A_UlofxvGN3_0),.din(w_dff_A_CAcrCyCy6_0),.clk(gclk));
	jdff dff_A_UlofxvGN3_0(.dout(w_dff_A_MB8Gfrb67_0),.din(w_dff_A_UlofxvGN3_0),.clk(gclk));
	jdff dff_A_MB8Gfrb67_0(.dout(w_dff_A_TmORDFHX5_0),.din(w_dff_A_MB8Gfrb67_0),.clk(gclk));
	jdff dff_A_TmORDFHX5_0(.dout(w_dff_A_3d3sMt6m5_0),.din(w_dff_A_TmORDFHX5_0),.clk(gclk));
	jdff dff_A_3d3sMt6m5_0(.dout(w_dff_A_PUJJon1W6_0),.din(w_dff_A_3d3sMt6m5_0),.clk(gclk));
	jdff dff_A_PUJJon1W6_0(.dout(w_dff_A_Gz5Kq3nn1_0),.din(w_dff_A_PUJJon1W6_0),.clk(gclk));
	jdff dff_A_Gz5Kq3nn1_0(.dout(w_dff_A_xJCTIBfG9_0),.din(w_dff_A_Gz5Kq3nn1_0),.clk(gclk));
	jdff dff_A_xJCTIBfG9_0(.dout(G998),.din(w_dff_A_xJCTIBfG9_0),.clk(gclk));
	jdff dff_A_vxWk0kuz4_1(.dout(w_dff_A_lol7tGyc9_0),.din(w_dff_A_vxWk0kuz4_1),.clk(gclk));
	jdff dff_A_lol7tGyc9_0(.dout(w_dff_A_iKEkTV5t6_0),.din(w_dff_A_lol7tGyc9_0),.clk(gclk));
	jdff dff_A_iKEkTV5t6_0(.dout(w_dff_A_o0iOlF0S9_0),.din(w_dff_A_iKEkTV5t6_0),.clk(gclk));
	jdff dff_A_o0iOlF0S9_0(.dout(w_dff_A_txTUDvuk0_0),.din(w_dff_A_o0iOlF0S9_0),.clk(gclk));
	jdff dff_A_txTUDvuk0_0(.dout(w_dff_A_gpSSDnqP8_0),.din(w_dff_A_txTUDvuk0_0),.clk(gclk));
	jdff dff_A_gpSSDnqP8_0(.dout(w_dff_A_gKKBMyGH2_0),.din(w_dff_A_gpSSDnqP8_0),.clk(gclk));
	jdff dff_A_gKKBMyGH2_0(.dout(w_dff_A_ujXf7ey06_0),.din(w_dff_A_gKKBMyGH2_0),.clk(gclk));
	jdff dff_A_ujXf7ey06_0(.dout(w_dff_A_qdLImWtr9_0),.din(w_dff_A_ujXf7ey06_0),.clk(gclk));
	jdff dff_A_qdLImWtr9_0(.dout(w_dff_A_a52EhNS14_0),.din(w_dff_A_qdLImWtr9_0),.clk(gclk));
	jdff dff_A_a52EhNS14_0(.dout(w_dff_A_C11h4Fyo7_0),.din(w_dff_A_a52EhNS14_0),.clk(gclk));
	jdff dff_A_C11h4Fyo7_0(.dout(w_dff_A_z4QWg72y8_0),.din(w_dff_A_C11h4Fyo7_0),.clk(gclk));
	jdff dff_A_z4QWg72y8_0(.dout(w_dff_A_18nj1Z018_0),.din(w_dff_A_z4QWg72y8_0),.clk(gclk));
	jdff dff_A_18nj1Z018_0(.dout(w_dff_A_P057rDQ20_0),.din(w_dff_A_18nj1Z018_0),.clk(gclk));
	jdff dff_A_P057rDQ20_0(.dout(w_dff_A_lqnMz7y54_0),.din(w_dff_A_P057rDQ20_0),.clk(gclk));
	jdff dff_A_lqnMz7y54_0(.dout(w_dff_A_TscTtr5T5_0),.din(w_dff_A_lqnMz7y54_0),.clk(gclk));
	jdff dff_A_TscTtr5T5_0(.dout(w_dff_A_WFluOpEp0_0),.din(w_dff_A_TscTtr5T5_0),.clk(gclk));
	jdff dff_A_WFluOpEp0_0(.dout(w_dff_A_v6IyGWyY9_0),.din(w_dff_A_WFluOpEp0_0),.clk(gclk));
	jdff dff_A_v6IyGWyY9_0(.dout(w_dff_A_UkYV04p32_0),.din(w_dff_A_v6IyGWyY9_0),.clk(gclk));
	jdff dff_A_UkYV04p32_0(.dout(G1000),.din(w_dff_A_UkYV04p32_0),.clk(gclk));
	jdff dff_A_ZwVSUgu01_2(.dout(w_dff_A_cx4CKnL32_0),.din(w_dff_A_ZwVSUgu01_2),.clk(gclk));
	jdff dff_A_cx4CKnL32_0(.dout(w_dff_A_PlH2NXOH3_0),.din(w_dff_A_cx4CKnL32_0),.clk(gclk));
	jdff dff_A_PlH2NXOH3_0(.dout(w_dff_A_XoYOnOg67_0),.din(w_dff_A_PlH2NXOH3_0),.clk(gclk));
	jdff dff_A_XoYOnOg67_0(.dout(w_dff_A_51s5SvMF4_0),.din(w_dff_A_XoYOnOg67_0),.clk(gclk));
	jdff dff_A_51s5SvMF4_0(.dout(G575),.din(w_dff_A_51s5SvMF4_0),.clk(gclk));
	jdff dff_A_aPAHZ5LL4_2(.dout(w_dff_A_1nQkdxS48_0),.din(w_dff_A_aPAHZ5LL4_2),.clk(gclk));
	jdff dff_A_1nQkdxS48_0(.dout(w_dff_A_SYXW0W7J6_0),.din(w_dff_A_1nQkdxS48_0),.clk(gclk));
	jdff dff_A_SYXW0W7J6_0(.dout(w_dff_A_JNkxd2Je5_0),.din(w_dff_A_SYXW0W7J6_0),.clk(gclk));
	jdff dff_A_JNkxd2Je5_0(.dout(w_dff_A_1sFFBQuW9_0),.din(w_dff_A_JNkxd2Je5_0),.clk(gclk));
	jdff dff_A_1sFFBQuW9_0(.dout(w_dff_A_UbtI2DGo5_0),.din(w_dff_A_1sFFBQuW9_0),.clk(gclk));
	jdff dff_A_UbtI2DGo5_0(.dout(w_dff_A_G63HbYJb4_0),.din(w_dff_A_UbtI2DGo5_0),.clk(gclk));
	jdff dff_A_G63HbYJb4_0(.dout(w_dff_A_FqGrfaly0_0),.din(w_dff_A_G63HbYJb4_0),.clk(gclk));
	jdff dff_A_FqGrfaly0_0(.dout(G585),.din(w_dff_A_FqGrfaly0_0),.clk(gclk));
	jdff dff_A_BjvcmaIf8_2(.dout(w_dff_A_O1uS5i5W7_0),.din(w_dff_A_BjvcmaIf8_2),.clk(gclk));
	jdff dff_A_O1uS5i5W7_0(.dout(w_dff_A_Iyon78Eh2_0),.din(w_dff_A_O1uS5i5W7_0),.clk(gclk));
	jdff dff_A_Iyon78Eh2_0(.dout(w_dff_A_PSu94Fp34_0),.din(w_dff_A_Iyon78Eh2_0),.clk(gclk));
	jdff dff_A_PSu94Fp34_0(.dout(w_dff_A_FJ6BLk6H5_0),.din(w_dff_A_PSu94Fp34_0),.clk(gclk));
	jdff dff_A_FJ6BLk6H5_0(.dout(w_dff_A_t8fnELcm5_0),.din(w_dff_A_FJ6BLk6H5_0),.clk(gclk));
	jdff dff_A_t8fnELcm5_0(.dout(w_dff_A_Qy9pUNkj4_0),.din(w_dff_A_t8fnELcm5_0),.clk(gclk));
	jdff dff_A_Qy9pUNkj4_0(.dout(w_dff_A_yw6LOFQ46_0),.din(w_dff_A_Qy9pUNkj4_0),.clk(gclk));
	jdff dff_A_yw6LOFQ46_0(.dout(w_dff_A_wvNU9kS00_0),.din(w_dff_A_yw6LOFQ46_0),.clk(gclk));
	jdff dff_A_wvNU9kS00_0(.dout(w_dff_A_1sDO05d45_0),.din(w_dff_A_wvNU9kS00_0),.clk(gclk));
	jdff dff_A_1sDO05d45_0(.dout(w_dff_A_gF1yE8Rg5_0),.din(w_dff_A_1sDO05d45_0),.clk(gclk));
	jdff dff_A_gF1yE8Rg5_0(.dout(w_dff_A_Y8i03vy06_0),.din(w_dff_A_gF1yE8Rg5_0),.clk(gclk));
	jdff dff_A_Y8i03vy06_0(.dout(w_dff_A_ONibe0tZ3_0),.din(w_dff_A_Y8i03vy06_0),.clk(gclk));
	jdff dff_A_ONibe0tZ3_0(.dout(w_dff_A_jjXailx57_0),.din(w_dff_A_ONibe0tZ3_0),.clk(gclk));
	jdff dff_A_jjXailx57_0(.dout(G661),.din(w_dff_A_jjXailx57_0),.clk(gclk));
	jdff dff_A_T2PMMgd24_2(.dout(w_dff_A_mZ8pUlFz5_0),.din(w_dff_A_T2PMMgd24_2),.clk(gclk));
	jdff dff_A_mZ8pUlFz5_0(.dout(w_dff_A_TNXH6GIs1_0),.din(w_dff_A_mZ8pUlFz5_0),.clk(gclk));
	jdff dff_A_TNXH6GIs1_0(.dout(w_dff_A_1ej4X1Vz2_0),.din(w_dff_A_TNXH6GIs1_0),.clk(gclk));
	jdff dff_A_1ej4X1Vz2_0(.dout(w_dff_A_KkGM2XdS9_0),.din(w_dff_A_1ej4X1Vz2_0),.clk(gclk));
	jdff dff_A_KkGM2XdS9_0(.dout(w_dff_A_I4WTF1c89_0),.din(w_dff_A_KkGM2XdS9_0),.clk(gclk));
	jdff dff_A_I4WTF1c89_0(.dout(w_dff_A_8IpmZLyl1_0),.din(w_dff_A_I4WTF1c89_0),.clk(gclk));
	jdff dff_A_8IpmZLyl1_0(.dout(w_dff_A_ncsfzng79_0),.din(w_dff_A_8IpmZLyl1_0),.clk(gclk));
	jdff dff_A_ncsfzng79_0(.dout(w_dff_A_I7zMWBsM7_0),.din(w_dff_A_ncsfzng79_0),.clk(gclk));
	jdff dff_A_I7zMWBsM7_0(.dout(w_dff_A_dHBnbEgv2_0),.din(w_dff_A_I7zMWBsM7_0),.clk(gclk));
	jdff dff_A_dHBnbEgv2_0(.dout(w_dff_A_7dbf1h419_0),.din(w_dff_A_dHBnbEgv2_0),.clk(gclk));
	jdff dff_A_7dbf1h419_0(.dout(w_dff_A_fTI4crZ25_0),.din(w_dff_A_7dbf1h419_0),.clk(gclk));
	jdff dff_A_fTI4crZ25_0(.dout(w_dff_A_3h2XP5c53_0),.din(w_dff_A_fTI4crZ25_0),.clk(gclk));
	jdff dff_A_3h2XP5c53_0(.dout(w_dff_A_MjH02BQJ1_0),.din(w_dff_A_3h2XP5c53_0),.clk(gclk));
	jdff dff_A_MjH02BQJ1_0(.dout(G693),.din(w_dff_A_MjH02BQJ1_0),.clk(gclk));
	jdff dff_A_xNgk3bJf2_2(.dout(w_dff_A_W2BFYOlt5_0),.din(w_dff_A_xNgk3bJf2_2),.clk(gclk));
	jdff dff_A_W2BFYOlt5_0(.dout(w_dff_A_s48iNXK05_0),.din(w_dff_A_W2BFYOlt5_0),.clk(gclk));
	jdff dff_A_s48iNXK05_0(.dout(w_dff_A_bKoO846w1_0),.din(w_dff_A_s48iNXK05_0),.clk(gclk));
	jdff dff_A_bKoO846w1_0(.dout(w_dff_A_VhQuBeBX9_0),.din(w_dff_A_bKoO846w1_0),.clk(gclk));
	jdff dff_A_VhQuBeBX9_0(.dout(w_dff_A_pP2OPXy75_0),.din(w_dff_A_VhQuBeBX9_0),.clk(gclk));
	jdff dff_A_pP2OPXy75_0(.dout(w_dff_A_UcorWion6_0),.din(w_dff_A_pP2OPXy75_0),.clk(gclk));
	jdff dff_A_UcorWion6_0(.dout(G747),.din(w_dff_A_UcorWion6_0),.clk(gclk));
	jdff dff_A_g0IwlMxo1_2(.dout(w_dff_A_lwtRUbdz2_0),.din(w_dff_A_g0IwlMxo1_2),.clk(gclk));
	jdff dff_A_lwtRUbdz2_0(.dout(w_dff_A_M8Yz6tkD9_0),.din(w_dff_A_lwtRUbdz2_0),.clk(gclk));
	jdff dff_A_M8Yz6tkD9_0(.dout(w_dff_A_jeVaUGCm4_0),.din(w_dff_A_M8Yz6tkD9_0),.clk(gclk));
	jdff dff_A_jeVaUGCm4_0(.dout(w_dff_A_ADLXexMg5_0),.din(w_dff_A_jeVaUGCm4_0),.clk(gclk));
	jdff dff_A_ADLXexMg5_0(.dout(w_dff_A_Ec8wgNHe0_0),.din(w_dff_A_ADLXexMg5_0),.clk(gclk));
	jdff dff_A_Ec8wgNHe0_0(.dout(w_dff_A_q1ZP4Ju71_0),.din(w_dff_A_Ec8wgNHe0_0),.clk(gclk));
	jdff dff_A_q1ZP4Ju71_0(.dout(w_dff_A_CWPC1Hao1_0),.din(w_dff_A_q1ZP4Ju71_0),.clk(gclk));
	jdff dff_A_CWPC1Hao1_0(.dout(w_dff_A_E9glpBty5_0),.din(w_dff_A_CWPC1Hao1_0),.clk(gclk));
	jdff dff_A_E9glpBty5_0(.dout(G752),.din(w_dff_A_E9glpBty5_0),.clk(gclk));
	jdff dff_A_m9mvQOBB9_2(.dout(w_dff_A_ksAJL9kY7_0),.din(w_dff_A_m9mvQOBB9_2),.clk(gclk));
	jdff dff_A_ksAJL9kY7_0(.dout(w_dff_A_1Y3wWmRJ0_0),.din(w_dff_A_ksAJL9kY7_0),.clk(gclk));
	jdff dff_A_1Y3wWmRJ0_0(.dout(w_dff_A_aPagkDPs1_0),.din(w_dff_A_1Y3wWmRJ0_0),.clk(gclk));
	jdff dff_A_aPagkDPs1_0(.dout(w_dff_A_QWdDj9Qn7_0),.din(w_dff_A_aPagkDPs1_0),.clk(gclk));
	jdff dff_A_QWdDj9Qn7_0(.dout(w_dff_A_njL2hrF09_0),.din(w_dff_A_QWdDj9Qn7_0),.clk(gclk));
	jdff dff_A_njL2hrF09_0(.dout(w_dff_A_xDSaxUyy4_0),.din(w_dff_A_njL2hrF09_0),.clk(gclk));
	jdff dff_A_xDSaxUyy4_0(.dout(w_dff_A_ltxeGomy7_0),.din(w_dff_A_xDSaxUyy4_0),.clk(gclk));
	jdff dff_A_ltxeGomy7_0(.dout(w_dff_A_2YYotMmc5_0),.din(w_dff_A_ltxeGomy7_0),.clk(gclk));
	jdff dff_A_2YYotMmc5_0(.dout(w_dff_A_yHFZUxf10_0),.din(w_dff_A_2YYotMmc5_0),.clk(gclk));
	jdff dff_A_yHFZUxf10_0(.dout(G757),.din(w_dff_A_yHFZUxf10_0),.clk(gclk));
	jdff dff_A_V5IgNeJF5_2(.dout(w_dff_A_WpKOQMgU6_0),.din(w_dff_A_V5IgNeJF5_2),.clk(gclk));
	jdff dff_A_WpKOQMgU6_0(.dout(w_dff_A_Q4LeZp0o5_0),.din(w_dff_A_WpKOQMgU6_0),.clk(gclk));
	jdff dff_A_Q4LeZp0o5_0(.dout(w_dff_A_FvOsX6rh2_0),.din(w_dff_A_Q4LeZp0o5_0),.clk(gclk));
	jdff dff_A_FvOsX6rh2_0(.dout(w_dff_A_7BkNzJCb6_0),.din(w_dff_A_FvOsX6rh2_0),.clk(gclk));
	jdff dff_A_7BkNzJCb6_0(.dout(w_dff_A_BJ3sBhf47_0),.din(w_dff_A_7BkNzJCb6_0),.clk(gclk));
	jdff dff_A_BJ3sBhf47_0(.dout(w_dff_A_eEZWHRGO0_0),.din(w_dff_A_BJ3sBhf47_0),.clk(gclk));
	jdff dff_A_eEZWHRGO0_0(.dout(w_dff_A_bC9aoJ696_0),.din(w_dff_A_eEZWHRGO0_0),.clk(gclk));
	jdff dff_A_bC9aoJ696_0(.dout(w_dff_A_XblsMeDR1_0),.din(w_dff_A_bC9aoJ696_0),.clk(gclk));
	jdff dff_A_XblsMeDR1_0(.dout(w_dff_A_EuGEL2YL8_0),.din(w_dff_A_XblsMeDR1_0),.clk(gclk));
	jdff dff_A_EuGEL2YL8_0(.dout(w_dff_A_psBQKyDZ2_0),.din(w_dff_A_EuGEL2YL8_0),.clk(gclk));
	jdff dff_A_psBQKyDZ2_0(.dout(G762),.din(w_dff_A_psBQKyDZ2_0),.clk(gclk));
	jdff dff_A_cPQHNv5B9_2(.dout(w_dff_A_Ex4eapIB2_0),.din(w_dff_A_cPQHNv5B9_2),.clk(gclk));
	jdff dff_A_Ex4eapIB2_0(.dout(w_dff_A_CDNEXem76_0),.din(w_dff_A_Ex4eapIB2_0),.clk(gclk));
	jdff dff_A_CDNEXem76_0(.dout(w_dff_A_j2MpnEKC7_0),.din(w_dff_A_CDNEXem76_0),.clk(gclk));
	jdff dff_A_j2MpnEKC7_0(.dout(w_dff_A_ccbMY84v3_0),.din(w_dff_A_j2MpnEKC7_0),.clk(gclk));
	jdff dff_A_ccbMY84v3_0(.dout(w_dff_A_jIVTXgdV8_0),.din(w_dff_A_ccbMY84v3_0),.clk(gclk));
	jdff dff_A_jIVTXgdV8_0(.dout(w_dff_A_HNL4anZJ1_0),.din(w_dff_A_jIVTXgdV8_0),.clk(gclk));
	jdff dff_A_HNL4anZJ1_0(.dout(G787),.din(w_dff_A_HNL4anZJ1_0),.clk(gclk));
	jdff dff_A_oRgwlr2S2_2(.dout(w_dff_A_uz6TL8Fv8_0),.din(w_dff_A_oRgwlr2S2_2),.clk(gclk));
	jdff dff_A_uz6TL8Fv8_0(.dout(w_dff_A_SU6dX10N2_0),.din(w_dff_A_uz6TL8Fv8_0),.clk(gclk));
	jdff dff_A_SU6dX10N2_0(.dout(w_dff_A_e658WdM31_0),.din(w_dff_A_SU6dX10N2_0),.clk(gclk));
	jdff dff_A_e658WdM31_0(.dout(w_dff_A_pGhyNCH50_0),.din(w_dff_A_e658WdM31_0),.clk(gclk));
	jdff dff_A_pGhyNCH50_0(.dout(w_dff_A_WJQibS2G0_0),.din(w_dff_A_pGhyNCH50_0),.clk(gclk));
	jdff dff_A_WJQibS2G0_0(.dout(w_dff_A_HUolGx9D6_0),.din(w_dff_A_WJQibS2G0_0),.clk(gclk));
	jdff dff_A_HUolGx9D6_0(.dout(w_dff_A_ICfuHqFr6_0),.din(w_dff_A_HUolGx9D6_0),.clk(gclk));
	jdff dff_A_ICfuHqFr6_0(.dout(w_dff_A_P7pf4Vfe9_0),.din(w_dff_A_ICfuHqFr6_0),.clk(gclk));
	jdff dff_A_P7pf4Vfe9_0(.dout(G792),.din(w_dff_A_P7pf4Vfe9_0),.clk(gclk));
	jdff dff_A_7sYsf6TN1_2(.dout(w_dff_A_vNqj2az50_0),.din(w_dff_A_7sYsf6TN1_2),.clk(gclk));
	jdff dff_A_vNqj2az50_0(.dout(w_dff_A_WyJvKw7E0_0),.din(w_dff_A_vNqj2az50_0),.clk(gclk));
	jdff dff_A_WyJvKw7E0_0(.dout(w_dff_A_7onYI73d0_0),.din(w_dff_A_WyJvKw7E0_0),.clk(gclk));
	jdff dff_A_7onYI73d0_0(.dout(w_dff_A_IqxEx9ys7_0),.din(w_dff_A_7onYI73d0_0),.clk(gclk));
	jdff dff_A_IqxEx9ys7_0(.dout(w_dff_A_XDTDN5YN7_0),.din(w_dff_A_IqxEx9ys7_0),.clk(gclk));
	jdff dff_A_XDTDN5YN7_0(.dout(w_dff_A_8xqp0GbX0_0),.din(w_dff_A_XDTDN5YN7_0),.clk(gclk));
	jdff dff_A_8xqp0GbX0_0(.dout(w_dff_A_7cTf1T4i3_0),.din(w_dff_A_8xqp0GbX0_0),.clk(gclk));
	jdff dff_A_7cTf1T4i3_0(.dout(w_dff_A_AGcDh32s5_0),.din(w_dff_A_7cTf1T4i3_0),.clk(gclk));
	jdff dff_A_AGcDh32s5_0(.dout(w_dff_A_NQrAO3Rv3_0),.din(w_dff_A_AGcDh32s5_0),.clk(gclk));
	jdff dff_A_NQrAO3Rv3_0(.dout(G797),.din(w_dff_A_NQrAO3Rv3_0),.clk(gclk));
	jdff dff_A_axuI5cBD5_2(.dout(w_dff_A_6qTWw12u7_0),.din(w_dff_A_axuI5cBD5_2),.clk(gclk));
	jdff dff_A_6qTWw12u7_0(.dout(w_dff_A_nlQVr92Q0_0),.din(w_dff_A_6qTWw12u7_0),.clk(gclk));
	jdff dff_A_nlQVr92Q0_0(.dout(w_dff_A_r8CcTp2v1_0),.din(w_dff_A_nlQVr92Q0_0),.clk(gclk));
	jdff dff_A_r8CcTp2v1_0(.dout(w_dff_A_FiW4QVMn3_0),.din(w_dff_A_r8CcTp2v1_0),.clk(gclk));
	jdff dff_A_FiW4QVMn3_0(.dout(w_dff_A_1Zb7RLc86_0),.din(w_dff_A_FiW4QVMn3_0),.clk(gclk));
	jdff dff_A_1Zb7RLc86_0(.dout(w_dff_A_OUTDsZUk6_0),.din(w_dff_A_1Zb7RLc86_0),.clk(gclk));
	jdff dff_A_OUTDsZUk6_0(.dout(w_dff_A_89UOq2Qy0_0),.din(w_dff_A_OUTDsZUk6_0),.clk(gclk));
	jdff dff_A_89UOq2Qy0_0(.dout(w_dff_A_l9nTWXBB3_0),.din(w_dff_A_89UOq2Qy0_0),.clk(gclk));
	jdff dff_A_l9nTWXBB3_0(.dout(w_dff_A_CYnA1xGP9_0),.din(w_dff_A_l9nTWXBB3_0),.clk(gclk));
	jdff dff_A_CYnA1xGP9_0(.dout(w_dff_A_aQZEqZ2H8_0),.din(w_dff_A_CYnA1xGP9_0),.clk(gclk));
	jdff dff_A_aQZEqZ2H8_0(.dout(G802),.din(w_dff_A_aQZEqZ2H8_0),.clk(gclk));
	jdff dff_A_6rpt8BSf5_2(.dout(w_dff_A_z17Rcdpv0_0),.din(w_dff_A_6rpt8BSf5_2),.clk(gclk));
	jdff dff_A_z17Rcdpv0_0(.dout(w_dff_A_KyNOtPHU3_0),.din(w_dff_A_z17Rcdpv0_0),.clk(gclk));
	jdff dff_A_KyNOtPHU3_0(.dout(w_dff_A_yawDQFw12_0),.din(w_dff_A_KyNOtPHU3_0),.clk(gclk));
	jdff dff_A_yawDQFw12_0(.dout(w_dff_A_cSrNiilW2_0),.din(w_dff_A_yawDQFw12_0),.clk(gclk));
	jdff dff_A_cSrNiilW2_0(.dout(w_dff_A_utYL87sS2_0),.din(w_dff_A_cSrNiilW2_0),.clk(gclk));
	jdff dff_A_utYL87sS2_0(.dout(G642),.din(w_dff_A_utYL87sS2_0),.clk(gclk));
	jdff dff_A_8re8Z0rV0_2(.dout(w_dff_A_GRR10IgP0_0),.din(w_dff_A_8re8Z0rV0_2),.clk(gclk));
	jdff dff_A_GRR10IgP0_0(.dout(w_dff_A_cJNFi75R8_0),.din(w_dff_A_GRR10IgP0_0),.clk(gclk));
	jdff dff_A_cJNFi75R8_0(.dout(w_dff_A_ndU0ew5q3_0),.din(w_dff_A_cJNFi75R8_0),.clk(gclk));
	jdff dff_A_ndU0ew5q3_0(.dout(w_dff_A_5tssc9dj5_0),.din(w_dff_A_ndU0ew5q3_0),.clk(gclk));
	jdff dff_A_5tssc9dj5_0(.dout(w_dff_A_6Ux2QBei0_0),.din(w_dff_A_5tssc9dj5_0),.clk(gclk));
	jdff dff_A_6Ux2QBei0_0(.dout(w_dff_A_cW0sIP7H9_0),.din(w_dff_A_6Ux2QBei0_0),.clk(gclk));
	jdff dff_A_cW0sIP7H9_0(.dout(w_dff_A_yZQ2yunU8_0),.din(w_dff_A_cW0sIP7H9_0),.clk(gclk));
	jdff dff_A_yZQ2yunU8_0(.dout(w_dff_A_inf7Of335_0),.din(w_dff_A_yZQ2yunU8_0),.clk(gclk));
	jdff dff_A_inf7Of335_0(.dout(w_dff_A_pTC26Tiz3_0),.din(w_dff_A_inf7Of335_0),.clk(gclk));
	jdff dff_A_pTC26Tiz3_0(.dout(G664),.din(w_dff_A_pTC26Tiz3_0),.clk(gclk));
	jdff dff_A_3hWNAct47_2(.dout(w_dff_A_vRwhH48E3_0),.din(w_dff_A_3hWNAct47_2),.clk(gclk));
	jdff dff_A_vRwhH48E3_0(.dout(w_dff_A_Cy3dTs2N4_0),.din(w_dff_A_vRwhH48E3_0),.clk(gclk));
	jdff dff_A_Cy3dTs2N4_0(.dout(w_dff_A_CdPWBX9T4_0),.din(w_dff_A_Cy3dTs2N4_0),.clk(gclk));
	jdff dff_A_CdPWBX9T4_0(.dout(w_dff_A_pNUKCvzA0_0),.din(w_dff_A_CdPWBX9T4_0),.clk(gclk));
	jdff dff_A_pNUKCvzA0_0(.dout(w_dff_A_yJUKYI1N5_0),.din(w_dff_A_pNUKCvzA0_0),.clk(gclk));
	jdff dff_A_yJUKYI1N5_0(.dout(w_dff_A_T2bI25Oj5_0),.din(w_dff_A_yJUKYI1N5_0),.clk(gclk));
	jdff dff_A_T2bI25Oj5_0(.dout(w_dff_A_zsBSBdfK1_0),.din(w_dff_A_T2bI25Oj5_0),.clk(gclk));
	jdff dff_A_zsBSBdfK1_0(.dout(w_dff_A_NK31XUtu1_0),.din(w_dff_A_zsBSBdfK1_0),.clk(gclk));
	jdff dff_A_NK31XUtu1_0(.dout(G667),.din(w_dff_A_NK31XUtu1_0),.clk(gclk));
	jdff dff_A_BCHA1aqF8_2(.dout(w_dff_A_4tbiLbgq2_0),.din(w_dff_A_BCHA1aqF8_2),.clk(gclk));
	jdff dff_A_4tbiLbgq2_0(.dout(w_dff_A_0rAlDyUm2_0),.din(w_dff_A_4tbiLbgq2_0),.clk(gclk));
	jdff dff_A_0rAlDyUm2_0(.dout(w_dff_A_ZpX5zIOT4_0),.din(w_dff_A_0rAlDyUm2_0),.clk(gclk));
	jdff dff_A_ZpX5zIOT4_0(.dout(w_dff_A_EAuFQQyb3_0),.din(w_dff_A_ZpX5zIOT4_0),.clk(gclk));
	jdff dff_A_EAuFQQyb3_0(.dout(w_dff_A_F4PkPkyH6_0),.din(w_dff_A_EAuFQQyb3_0),.clk(gclk));
	jdff dff_A_F4PkPkyH6_0(.dout(w_dff_A_c9VTKL0p0_0),.din(w_dff_A_F4PkPkyH6_0),.clk(gclk));
	jdff dff_A_c9VTKL0p0_0(.dout(w_dff_A_4ZYvl2q66_0),.din(w_dff_A_c9VTKL0p0_0),.clk(gclk));
	jdff dff_A_4ZYvl2q66_0(.dout(G670),.din(w_dff_A_4ZYvl2q66_0),.clk(gclk));
	jdff dff_A_Dt6jwWtM8_2(.dout(w_dff_A_X8y2MPUc5_0),.din(w_dff_A_Dt6jwWtM8_2),.clk(gclk));
	jdff dff_A_X8y2MPUc5_0(.dout(w_dff_A_01xYAUnS3_0),.din(w_dff_A_X8y2MPUc5_0),.clk(gclk));
	jdff dff_A_01xYAUnS3_0(.dout(w_dff_A_HRPcuduB5_0),.din(w_dff_A_01xYAUnS3_0),.clk(gclk));
	jdff dff_A_HRPcuduB5_0(.dout(w_dff_A_Wbt5YpQd5_0),.din(w_dff_A_HRPcuduB5_0),.clk(gclk));
	jdff dff_A_Wbt5YpQd5_0(.dout(w_dff_A_t38XyCSz3_0),.din(w_dff_A_Wbt5YpQd5_0),.clk(gclk));
	jdff dff_A_t38XyCSz3_0(.dout(G676),.din(w_dff_A_t38XyCSz3_0),.clk(gclk));
	jdff dff_A_MqQBwMxU9_2(.dout(w_dff_A_8PyI6sKE1_0),.din(w_dff_A_MqQBwMxU9_2),.clk(gclk));
	jdff dff_A_8PyI6sKE1_0(.dout(w_dff_A_KosG7yld5_0),.din(w_dff_A_8PyI6sKE1_0),.clk(gclk));
	jdff dff_A_KosG7yld5_0(.dout(w_dff_A_Ei7LzMha6_0),.din(w_dff_A_KosG7yld5_0),.clk(gclk));
	jdff dff_A_Ei7LzMha6_0(.dout(w_dff_A_I4j4iM1L0_0),.din(w_dff_A_Ei7LzMha6_0),.clk(gclk));
	jdff dff_A_I4j4iM1L0_0(.dout(w_dff_A_LhURLAYy2_0),.din(w_dff_A_I4j4iM1L0_0),.clk(gclk));
	jdff dff_A_LhURLAYy2_0(.dout(w_dff_A_H303VnPt9_0),.din(w_dff_A_LhURLAYy2_0),.clk(gclk));
	jdff dff_A_H303VnPt9_0(.dout(w_dff_A_Pgb2sB8L8_0),.din(w_dff_A_H303VnPt9_0),.clk(gclk));
	jdff dff_A_Pgb2sB8L8_0(.dout(w_dff_A_jOZEJrWW1_0),.din(w_dff_A_Pgb2sB8L8_0),.clk(gclk));
	jdff dff_A_jOZEJrWW1_0(.dout(w_dff_A_RYqammxv7_0),.din(w_dff_A_jOZEJrWW1_0),.clk(gclk));
	jdff dff_A_RYqammxv7_0(.dout(G696),.din(w_dff_A_RYqammxv7_0),.clk(gclk));
	jdff dff_A_AX6UZEQe8_2(.dout(w_dff_A_JGwoNHNd1_0),.din(w_dff_A_AX6UZEQe8_2),.clk(gclk));
	jdff dff_A_JGwoNHNd1_0(.dout(w_dff_A_DLSBcTjB7_0),.din(w_dff_A_JGwoNHNd1_0),.clk(gclk));
	jdff dff_A_DLSBcTjB7_0(.dout(w_dff_A_60WASzlJ6_0),.din(w_dff_A_DLSBcTjB7_0),.clk(gclk));
	jdff dff_A_60WASzlJ6_0(.dout(w_dff_A_5DR4MYjN6_0),.din(w_dff_A_60WASzlJ6_0),.clk(gclk));
	jdff dff_A_5DR4MYjN6_0(.dout(w_dff_A_1fEYA2CO0_0),.din(w_dff_A_5DR4MYjN6_0),.clk(gclk));
	jdff dff_A_1fEYA2CO0_0(.dout(w_dff_A_VEesDnjg3_0),.din(w_dff_A_1fEYA2CO0_0),.clk(gclk));
	jdff dff_A_VEesDnjg3_0(.dout(w_dff_A_w0wt9ylw3_0),.din(w_dff_A_VEesDnjg3_0),.clk(gclk));
	jdff dff_A_w0wt9ylw3_0(.dout(w_dff_A_74UZtK6D7_0),.din(w_dff_A_w0wt9ylw3_0),.clk(gclk));
	jdff dff_A_74UZtK6D7_0(.dout(G699),.din(w_dff_A_74UZtK6D7_0),.clk(gclk));
	jdff dff_A_pI4UzbjX7_2(.dout(w_dff_A_PD7GVt7w3_0),.din(w_dff_A_pI4UzbjX7_2),.clk(gclk));
	jdff dff_A_PD7GVt7w3_0(.dout(w_dff_A_VIbBDNCn6_0),.din(w_dff_A_PD7GVt7w3_0),.clk(gclk));
	jdff dff_A_VIbBDNCn6_0(.dout(w_dff_A_W0P9SmEA4_0),.din(w_dff_A_VIbBDNCn6_0),.clk(gclk));
	jdff dff_A_W0P9SmEA4_0(.dout(w_dff_A_Ny37ee9D9_0),.din(w_dff_A_W0P9SmEA4_0),.clk(gclk));
	jdff dff_A_Ny37ee9D9_0(.dout(w_dff_A_q0FWV8NW2_0),.din(w_dff_A_Ny37ee9D9_0),.clk(gclk));
	jdff dff_A_q0FWV8NW2_0(.dout(w_dff_A_ShpImyfo3_0),.din(w_dff_A_q0FWV8NW2_0),.clk(gclk));
	jdff dff_A_ShpImyfo3_0(.dout(w_dff_A_NbP1wXAe0_0),.din(w_dff_A_ShpImyfo3_0),.clk(gclk));
	jdff dff_A_NbP1wXAe0_0(.dout(G702),.din(w_dff_A_NbP1wXAe0_0),.clk(gclk));
	jdff dff_A_PL0nReCd3_2(.dout(w_dff_A_u6EqJ3Cf5_0),.din(w_dff_A_PL0nReCd3_2),.clk(gclk));
	jdff dff_A_u6EqJ3Cf5_0(.dout(w_dff_A_irnvtUxB4_0),.din(w_dff_A_u6EqJ3Cf5_0),.clk(gclk));
	jdff dff_A_irnvtUxB4_0(.dout(w_dff_A_Nmyz9r8A8_0),.din(w_dff_A_irnvtUxB4_0),.clk(gclk));
	jdff dff_A_Nmyz9r8A8_0(.dout(w_dff_A_0pY5zyR49_0),.din(w_dff_A_Nmyz9r8A8_0),.clk(gclk));
	jdff dff_A_0pY5zyR49_0(.dout(G818),.din(w_dff_A_0pY5zyR49_0),.clk(gclk));
	jdff dff_A_wjwk8NfH6_2(.dout(w_dff_A_xgw7p0Rd0_0),.din(w_dff_A_wjwk8NfH6_2),.clk(gclk));
	jdff dff_A_xgw7p0Rd0_0(.dout(w_dff_A_2MfCMQnB8_0),.din(w_dff_A_xgw7p0Rd0_0),.clk(gclk));
	jdff dff_A_2MfCMQnB8_0(.dout(w_dff_A_osVvMOyj5_0),.din(w_dff_A_2MfCMQnB8_0),.clk(gclk));
	jdff dff_A_osVvMOyj5_0(.dout(w_dff_A_pWQMjWgi5_0),.din(w_dff_A_osVvMOyj5_0),.clk(gclk));
	jdff dff_A_pWQMjWgi5_0(.dout(w_dff_A_MgBElAsh9_0),.din(w_dff_A_pWQMjWgi5_0),.clk(gclk));
	jdff dff_A_MgBElAsh9_0(.dout(w_dff_A_Fc2CDHyE3_0),.din(w_dff_A_MgBElAsh9_0),.clk(gclk));
	jdff dff_A_Fc2CDHyE3_0(.dout(w_dff_A_KEmcbVxm3_0),.din(w_dff_A_Fc2CDHyE3_0),.clk(gclk));
	jdff dff_A_KEmcbVxm3_0(.dout(w_dff_A_r5dLtpmm2_0),.din(w_dff_A_KEmcbVxm3_0),.clk(gclk));
	jdff dff_A_r5dLtpmm2_0(.dout(G813),.din(w_dff_A_r5dLtpmm2_0),.clk(gclk));
	jdff dff_A_H9l19U0M7_1(.dout(w_dff_A_sXU9p2Em6_0),.din(w_dff_A_H9l19U0M7_1),.clk(gclk));
	jdff dff_A_sXU9p2Em6_0(.dout(w_dff_A_s63tS9o31_0),.din(w_dff_A_sXU9p2Em6_0),.clk(gclk));
	jdff dff_A_s63tS9o31_0(.dout(w_dff_A_ll0iwTxF4_0),.din(w_dff_A_s63tS9o31_0),.clk(gclk));
	jdff dff_A_ll0iwTxF4_0(.dout(w_dff_A_BS2SFMqn9_0),.din(w_dff_A_ll0iwTxF4_0),.clk(gclk));
	jdff dff_A_BS2SFMqn9_0(.dout(G824),.din(w_dff_A_BS2SFMqn9_0),.clk(gclk));
	jdff dff_A_G7R4DQMb4_1(.dout(w_dff_A_YL4vOG652_0),.din(w_dff_A_G7R4DQMb4_1),.clk(gclk));
	jdff dff_A_YL4vOG652_0(.dout(w_dff_A_bDH0qyyM4_0),.din(w_dff_A_YL4vOG652_0),.clk(gclk));
	jdff dff_A_bDH0qyyM4_0(.dout(w_dff_A_wEHEWSJm2_0),.din(w_dff_A_bDH0qyyM4_0),.clk(gclk));
	jdff dff_A_wEHEWSJm2_0(.dout(w_dff_A_SjK7TBBe2_0),.din(w_dff_A_wEHEWSJm2_0),.clk(gclk));
	jdff dff_A_SjK7TBBe2_0(.dout(w_dff_A_AR8ckWXU8_0),.din(w_dff_A_SjK7TBBe2_0),.clk(gclk));
	jdff dff_A_AR8ckWXU8_0(.dout(w_dff_A_ju0hEPEo9_0),.din(w_dff_A_AR8ckWXU8_0),.clk(gclk));
	jdff dff_A_ju0hEPEo9_0(.dout(w_dff_A_5aEQ9g5v0_0),.din(w_dff_A_ju0hEPEo9_0),.clk(gclk));
	jdff dff_A_5aEQ9g5v0_0(.dout(G826),.din(w_dff_A_5aEQ9g5v0_0),.clk(gclk));
	jdff dff_A_Bmlo6mAl5_1(.dout(w_dff_A_U8enSGN17_0),.din(w_dff_A_Bmlo6mAl5_1),.clk(gclk));
	jdff dff_A_U8enSGN17_0(.dout(w_dff_A_AZMS5jDx8_0),.din(w_dff_A_U8enSGN17_0),.clk(gclk));
	jdff dff_A_AZMS5jDx8_0(.dout(w_dff_A_XlDDOS1I0_0),.din(w_dff_A_AZMS5jDx8_0),.clk(gclk));
	jdff dff_A_XlDDOS1I0_0(.dout(w_dff_A_EC7USFKY8_0),.din(w_dff_A_XlDDOS1I0_0),.clk(gclk));
	jdff dff_A_EC7USFKY8_0(.dout(w_dff_A_QdSxRkTV5_0),.din(w_dff_A_EC7USFKY8_0),.clk(gclk));
	jdff dff_A_QdSxRkTV5_0(.dout(w_dff_A_IPO3asO77_0),.din(w_dff_A_QdSxRkTV5_0),.clk(gclk));
	jdff dff_A_IPO3asO77_0(.dout(w_dff_A_IEdhuDou6_0),.din(w_dff_A_IPO3asO77_0),.clk(gclk));
	jdff dff_A_IEdhuDou6_0(.dout(G828),.din(w_dff_A_IEdhuDou6_0),.clk(gclk));
	jdff dff_A_FIVSn6jT5_1(.dout(w_dff_A_Qi12p23v0_0),.din(w_dff_A_FIVSn6jT5_1),.clk(gclk));
	jdff dff_A_Qi12p23v0_0(.dout(w_dff_A_nTf3kGoq3_0),.din(w_dff_A_Qi12p23v0_0),.clk(gclk));
	jdff dff_A_nTf3kGoq3_0(.dout(w_dff_A_aqjkUbL88_0),.din(w_dff_A_nTf3kGoq3_0),.clk(gclk));
	jdff dff_A_aqjkUbL88_0(.dout(w_dff_A_eJEjRJto9_0),.din(w_dff_A_aqjkUbL88_0),.clk(gclk));
	jdff dff_A_eJEjRJto9_0(.dout(w_dff_A_hqvWELcf9_0),.din(w_dff_A_eJEjRJto9_0),.clk(gclk));
	jdff dff_A_hqvWELcf9_0(.dout(w_dff_A_oW4Mql2N5_0),.din(w_dff_A_hqvWELcf9_0),.clk(gclk));
	jdff dff_A_oW4Mql2N5_0(.dout(w_dff_A_CGCd2iDo0_0),.din(w_dff_A_oW4Mql2N5_0),.clk(gclk));
	jdff dff_A_CGCd2iDo0_0(.dout(w_dff_A_vkIbfGlh2_0),.din(w_dff_A_CGCd2iDo0_0),.clk(gclk));
	jdff dff_A_vkIbfGlh2_0(.dout(G830),.din(w_dff_A_vkIbfGlh2_0),.clk(gclk));
	jdff dff_A_kppvDxAs8_2(.dout(w_dff_A_CJc1MQX59_0),.din(w_dff_A_kppvDxAs8_2),.clk(gclk));
	jdff dff_A_CJc1MQX59_0(.dout(w_dff_A_NHzDBLZ10_0),.din(w_dff_A_CJc1MQX59_0),.clk(gclk));
	jdff dff_A_NHzDBLZ10_0(.dout(w_dff_A_0kZnrD8X5_0),.din(w_dff_A_NHzDBLZ10_0),.clk(gclk));
	jdff dff_A_0kZnrD8X5_0(.dout(w_dff_A_FQcx36GC3_0),.din(w_dff_A_0kZnrD8X5_0),.clk(gclk));
	jdff dff_A_FQcx36GC3_0(.dout(w_dff_A_7HfiSwIN0_0),.din(w_dff_A_FQcx36GC3_0),.clk(gclk));
	jdff dff_A_7HfiSwIN0_0(.dout(w_dff_A_K4h0biQT9_0),.din(w_dff_A_7HfiSwIN0_0),.clk(gclk));
	jdff dff_A_K4h0biQT9_0(.dout(w_dff_A_OIHn8raU3_0),.din(w_dff_A_K4h0biQT9_0),.clk(gclk));
	jdff dff_A_OIHn8raU3_0(.dout(w_dff_A_zwbI27Zl7_0),.din(w_dff_A_OIHn8raU3_0),.clk(gclk));
	jdff dff_A_zwbI27Zl7_0(.dout(w_dff_A_qiqBJ46L3_0),.din(w_dff_A_zwbI27Zl7_0),.clk(gclk));
	jdff dff_A_qiqBJ46L3_0(.dout(w_dff_A_JuBUJKWv1_0),.din(w_dff_A_qiqBJ46L3_0),.clk(gclk));
	jdff dff_A_JuBUJKWv1_0(.dout(w_dff_A_a2gz8XBV4_0),.din(w_dff_A_JuBUJKWv1_0),.clk(gclk));
	jdff dff_A_a2gz8XBV4_0(.dout(w_dff_A_fBGxTbSY1_0),.din(w_dff_A_a2gz8XBV4_0),.clk(gclk));
	jdff dff_A_fBGxTbSY1_0(.dout(w_dff_A_vLnah9Nh3_0),.din(w_dff_A_fBGxTbSY1_0),.clk(gclk));
	jdff dff_A_vLnah9Nh3_0(.dout(w_dff_A_zEGDd7WI3_0),.din(w_dff_A_vLnah9Nh3_0),.clk(gclk));
	jdff dff_A_zEGDd7WI3_0(.dout(w_dff_A_G2xREmvo6_0),.din(w_dff_A_zEGDd7WI3_0),.clk(gclk));
	jdff dff_A_G2xREmvo6_0(.dout(G854),.din(w_dff_A_G2xREmvo6_0),.clk(gclk));
	jdff dff_A_Db0Se1s10_1(.dout(w_dff_A_0yPptQX48_0),.din(w_dff_A_Db0Se1s10_1),.clk(gclk));
	jdff dff_A_0yPptQX48_0(.dout(w_dff_A_ve4s6jcr8_0),.din(w_dff_A_0yPptQX48_0),.clk(gclk));
	jdff dff_A_ve4s6jcr8_0(.dout(w_dff_A_ybX7Iq9q0_0),.din(w_dff_A_ve4s6jcr8_0),.clk(gclk));
	jdff dff_A_ybX7Iq9q0_0(.dout(G863),.din(w_dff_A_ybX7Iq9q0_0),.clk(gclk));
	jdff dff_A_Xvirj3x92_1(.dout(w_dff_A_9HLefwsM7_0),.din(w_dff_A_Xvirj3x92_1),.clk(gclk));
	jdff dff_A_9HLefwsM7_0(.dout(w_dff_A_ZKR4KOu15_0),.din(w_dff_A_9HLefwsM7_0),.clk(gclk));
	jdff dff_A_ZKR4KOu15_0(.dout(w_dff_A_1vfEAqKj1_0),.din(w_dff_A_ZKR4KOu15_0),.clk(gclk));
	jdff dff_A_1vfEAqKj1_0(.dout(w_dff_A_UTqRB3JZ8_0),.din(w_dff_A_1vfEAqKj1_0),.clk(gclk));
	jdff dff_A_UTqRB3JZ8_0(.dout(G865),.din(w_dff_A_UTqRB3JZ8_0),.clk(gclk));
	jdff dff_A_0gsqbsOX9_1(.dout(w_dff_A_2MU3zQs79_0),.din(w_dff_A_0gsqbsOX9_1),.clk(gclk));
	jdff dff_A_2MU3zQs79_0(.dout(w_dff_A_8YV8pcFe0_0),.din(w_dff_A_2MU3zQs79_0),.clk(gclk));
	jdff dff_A_8YV8pcFe0_0(.dout(w_dff_A_clG1kHoL9_0),.din(w_dff_A_8YV8pcFe0_0),.clk(gclk));
	jdff dff_A_clG1kHoL9_0(.dout(w_dff_A_DN5dca3V1_0),.din(w_dff_A_clG1kHoL9_0),.clk(gclk));
	jdff dff_A_DN5dca3V1_0(.dout(w_dff_A_0s4VnOCC6_0),.din(w_dff_A_DN5dca3V1_0),.clk(gclk));
	jdff dff_A_0s4VnOCC6_0(.dout(w_dff_A_2JE9l8j69_0),.din(w_dff_A_0s4VnOCC6_0),.clk(gclk));
	jdff dff_A_2JE9l8j69_0(.dout(G867),.din(w_dff_A_2JE9l8j69_0),.clk(gclk));
	jdff dff_A_Y9DXbQ481_1(.dout(w_dff_A_kyD7zK7U1_0),.din(w_dff_A_Y9DXbQ481_1),.clk(gclk));
	jdff dff_A_kyD7zK7U1_0(.dout(w_dff_A_1rSdnZCe4_0),.din(w_dff_A_kyD7zK7U1_0),.clk(gclk));
	jdff dff_A_1rSdnZCe4_0(.dout(w_dff_A_xdEoz0CS8_0),.din(w_dff_A_1rSdnZCe4_0),.clk(gclk));
	jdff dff_A_xdEoz0CS8_0(.dout(w_dff_A_3jeAbU1w5_0),.din(w_dff_A_xdEoz0CS8_0),.clk(gclk));
	jdff dff_A_3jeAbU1w5_0(.dout(w_dff_A_NjzqUsoA9_0),.din(w_dff_A_3jeAbU1w5_0),.clk(gclk));
	jdff dff_A_NjzqUsoA9_0(.dout(w_dff_A_6yUTm2Ws8_0),.din(w_dff_A_NjzqUsoA9_0),.clk(gclk));
	jdff dff_A_6yUTm2Ws8_0(.dout(w_dff_A_rCo1GP2Y6_0),.din(w_dff_A_6yUTm2Ws8_0),.clk(gclk));
	jdff dff_A_rCo1GP2Y6_0(.dout(G869),.din(w_dff_A_rCo1GP2Y6_0),.clk(gclk));
	jdff dff_A_UTwmXiJV5_2(.dout(w_dff_A_TXy3L1NG6_0),.din(w_dff_A_UTwmXiJV5_2),.clk(gclk));
	jdff dff_A_TXy3L1NG6_0(.dout(w_dff_A_fWRL19Y44_0),.din(w_dff_A_TXy3L1NG6_0),.clk(gclk));
	jdff dff_A_fWRL19Y44_0(.dout(G712),.din(w_dff_A_fWRL19Y44_0),.clk(gclk));
	jdff dff_A_cpxnTtkT7_2(.dout(w_dff_A_DkB9eyZc1_0),.din(w_dff_A_cpxnTtkT7_2),.clk(gclk));
	jdff dff_A_DkB9eyZc1_0(.dout(w_dff_A_vkSUaR3g5_0),.din(w_dff_A_DkB9eyZc1_0),.clk(gclk));
	jdff dff_A_vkSUaR3g5_0(.dout(G727),.din(w_dff_A_vkSUaR3g5_0),.clk(gclk));
	jdff dff_A_zT3XBVAo1_2(.dout(w_dff_A_DUQ5RHt73_0),.din(w_dff_A_zT3XBVAo1_2),.clk(gclk));
	jdff dff_A_DUQ5RHt73_0(.dout(w_dff_A_3mGJs6Ph6_0),.din(w_dff_A_DUQ5RHt73_0),.clk(gclk));
	jdff dff_A_3mGJs6Ph6_0(.dout(w_dff_A_Wh7K7oZ84_0),.din(w_dff_A_3mGJs6Ph6_0),.clk(gclk));
	jdff dff_A_Wh7K7oZ84_0(.dout(G732),.din(w_dff_A_Wh7K7oZ84_0),.clk(gclk));
	jdff dff_A_8UD0c5Ru2_2(.dout(w_dff_A_tWlDItD29_0),.din(w_dff_A_8UD0c5Ru2_2),.clk(gclk));
	jdff dff_A_tWlDItD29_0(.dout(w_dff_A_AqPdayHI6_0),.din(w_dff_A_tWlDItD29_0),.clk(gclk));
	jdff dff_A_AqPdayHI6_0(.dout(w_dff_A_nF3iWpjD1_0),.din(w_dff_A_AqPdayHI6_0),.clk(gclk));
	jdff dff_A_nF3iWpjD1_0(.dout(G737),.din(w_dff_A_nF3iWpjD1_0),.clk(gclk));
	jdff dff_A_PIldz9RX9_2(.dout(w_dff_A_sD9RiPX72_0),.din(w_dff_A_PIldz9RX9_2),.clk(gclk));
	jdff dff_A_sD9RiPX72_0(.dout(w_dff_A_WO8lGLWg1_0),.din(w_dff_A_sD9RiPX72_0),.clk(gclk));
	jdff dff_A_WO8lGLWg1_0(.dout(w_dff_A_u65Zf4pJ9_0),.din(w_dff_A_WO8lGLWg1_0),.clk(gclk));
	jdff dff_A_u65Zf4pJ9_0(.dout(w_dff_A_EWnvNPoH7_0),.din(w_dff_A_u65Zf4pJ9_0),.clk(gclk));
	jdff dff_A_EWnvNPoH7_0(.dout(G742),.din(w_dff_A_EWnvNPoH7_0),.clk(gclk));
	jdff dff_A_zLFP5pWE0_2(.dout(w_dff_A_ngOjbvSY8_0),.din(w_dff_A_zLFP5pWE0_2),.clk(gclk));
	jdff dff_A_ngOjbvSY8_0(.dout(w_dff_A_YB3NsWiX5_0),.din(w_dff_A_ngOjbvSY8_0),.clk(gclk));
	jdff dff_A_YB3NsWiX5_0(.dout(w_dff_A_4jrRbgWU5_0),.din(w_dff_A_YB3NsWiX5_0),.clk(gclk));
	jdff dff_A_4jrRbgWU5_0(.dout(G772),.din(w_dff_A_4jrRbgWU5_0),.clk(gclk));
	jdff dff_A_Jc6Rpzbn3_2(.dout(w_dff_A_USWGTGjs0_0),.din(w_dff_A_Jc6Rpzbn3_2),.clk(gclk));
	jdff dff_A_USWGTGjs0_0(.dout(w_dff_A_AYIiujB36_0),.din(w_dff_A_USWGTGjs0_0),.clk(gclk));
	jdff dff_A_AYIiujB36_0(.dout(w_dff_A_2oSbqiNS6_0),.din(w_dff_A_AYIiujB36_0),.clk(gclk));
	jdff dff_A_2oSbqiNS6_0(.dout(G777),.din(w_dff_A_2oSbqiNS6_0),.clk(gclk));
	jdff dff_A_W3LY4oTh8_2(.dout(w_dff_A_p4Z6OHCa9_0),.din(w_dff_A_W3LY4oTh8_2),.clk(gclk));
	jdff dff_A_p4Z6OHCa9_0(.dout(w_dff_A_Uh9DHK8c5_0),.din(w_dff_A_p4Z6OHCa9_0),.clk(gclk));
	jdff dff_A_Uh9DHK8c5_0(.dout(w_dff_A_mtX3FGsz2_0),.din(w_dff_A_Uh9DHK8c5_0),.clk(gclk));
	jdff dff_A_mtX3FGsz2_0(.dout(w_dff_A_TCsuykfJ9_0),.din(w_dff_A_mtX3FGsz2_0),.clk(gclk));
	jdff dff_A_TCsuykfJ9_0(.dout(G782),.din(w_dff_A_TCsuykfJ9_0),.clk(gclk));
	jdff dff_A_FMg1FwX22_2(.dout(w_dff_A_oMhcGBxd0_0),.din(w_dff_A_FMg1FwX22_2),.clk(gclk));
	jdff dff_A_oMhcGBxd0_0(.dout(w_dff_A_DlsGPHEV0_0),.din(w_dff_A_oMhcGBxd0_0),.clk(gclk));
	jdff dff_A_DlsGPHEV0_0(.dout(w_dff_A_R2caKM6X3_0),.din(w_dff_A_DlsGPHEV0_0),.clk(gclk));
	jdff dff_A_R2caKM6X3_0(.dout(G645),.din(w_dff_A_R2caKM6X3_0),.clk(gclk));
	jdff dff_A_1QlhlnXk4_2(.dout(w_dff_A_0phmmXY59_0),.din(w_dff_A_1QlhlnXk4_2),.clk(gclk));
	jdff dff_A_0phmmXY59_0(.dout(w_dff_A_9HeNAnN46_0),.din(w_dff_A_0phmmXY59_0),.clk(gclk));
	jdff dff_A_9HeNAnN46_0(.dout(G648),.din(w_dff_A_9HeNAnN46_0),.clk(gclk));
	jdff dff_A_yqoRBsWS7_2(.dout(w_dff_A_HJOc8wDx5_0),.din(w_dff_A_yqoRBsWS7_2),.clk(gclk));
	jdff dff_A_HJOc8wDx5_0(.dout(w_dff_A_wNH9s7Zb0_0),.din(w_dff_A_HJOc8wDx5_0),.clk(gclk));
	jdff dff_A_wNH9s7Zb0_0(.dout(G651),.din(w_dff_A_wNH9s7Zb0_0),.clk(gclk));
	jdff dff_A_GDUy23aV8_2(.dout(w_dff_A_3cv1kEqb2_0),.din(w_dff_A_GDUy23aV8_2),.clk(gclk));
	jdff dff_A_3cv1kEqb2_0(.dout(G654),.din(w_dff_A_3cv1kEqb2_0),.clk(gclk));
	jdff dff_A_Koy1Jatt2_2(.dout(w_dff_A_2UHCS21P1_0),.din(w_dff_A_Koy1Jatt2_2),.clk(gclk));
	jdff dff_A_2UHCS21P1_0(.dout(w_dff_A_gmRVeP8O9_0),.din(w_dff_A_2UHCS21P1_0),.clk(gclk));
	jdff dff_A_gmRVeP8O9_0(.dout(w_dff_A_TAD277UN8_0),.din(w_dff_A_gmRVeP8O9_0),.clk(gclk));
	jdff dff_A_TAD277UN8_0(.dout(G679),.din(w_dff_A_TAD277UN8_0),.clk(gclk));
	jdff dff_A_pBwC6pVv9_2(.dout(w_dff_A_uRcD19pB1_0),.din(w_dff_A_pBwC6pVv9_2),.clk(gclk));
	jdff dff_A_uRcD19pB1_0(.dout(w_dff_A_gRXC4Tr85_0),.din(w_dff_A_uRcD19pB1_0),.clk(gclk));
	jdff dff_A_gRXC4Tr85_0(.dout(G682),.din(w_dff_A_gRXC4Tr85_0),.clk(gclk));
	jdff dff_A_R1XS5Ihe0_2(.dout(w_dff_A_gk80YyZu3_0),.din(w_dff_A_R1XS5Ihe0_2),.clk(gclk));
	jdff dff_A_gk80YyZu3_0(.dout(w_dff_A_tBzr0fGn3_0),.din(w_dff_A_gk80YyZu3_0),.clk(gclk));
	jdff dff_A_tBzr0fGn3_0(.dout(G685),.din(w_dff_A_tBzr0fGn3_0),.clk(gclk));
	jdff dff_A_8T6yUygj4_2(.dout(w_dff_A_83ihCwOD9_0),.din(w_dff_A_8T6yUygj4_2),.clk(gclk));
	jdff dff_A_83ihCwOD9_0(.dout(G688),.din(w_dff_A_83ihCwOD9_0),.clk(gclk));
	jdff dff_A_SURhQcVE9_2(.dout(w_dff_A_5JQSpGdh3_0),.din(w_dff_A_SURhQcVE9_2),.clk(gclk));
	jdff dff_A_5JQSpGdh3_0(.dout(w_dff_A_IphPcu077_0),.din(w_dff_A_5JQSpGdh3_0),.clk(gclk));
	jdff dff_A_IphPcu077_0(.dout(w_dff_A_pNCoGSMR1_0),.din(w_dff_A_IphPcu077_0),.clk(gclk));
	jdff dff_A_pNCoGSMR1_0(.dout(G843),.din(w_dff_A_pNCoGSMR1_0),.clk(gclk));
	jdff dff_A_uG8smKgl3_2(.dout(w_dff_A_YDRa4Cqv9_0),.din(w_dff_A_uG8smKgl3_2),.clk(gclk));
	jdff dff_A_YDRa4Cqv9_0(.dout(w_dff_A_Gb01iVMQ7_0),.din(w_dff_A_YDRa4Cqv9_0),.clk(gclk));
	jdff dff_A_Gb01iVMQ7_0(.dout(w_dff_A_B66RrRug7_0),.din(w_dff_A_Gb01iVMQ7_0),.clk(gclk));
	jdff dff_A_B66RrRug7_0(.dout(G882),.din(w_dff_A_B66RrRug7_0),.clk(gclk));
	jdff dff_A_jKaG1UkO8_2(.dout(G767),.din(w_dff_A_jKaG1UkO8_2),.clk(gclk));
	jdff dff_A_1hgo6KA25_2(.dout(G807),.din(w_dff_A_1hgo6KA25_2),.clk(gclk));
endmodule

