/*
gf_c880:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1588
	jand: 151
	jor: 122

Summary:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1588
	jand: 151
	jor: 122

The maximum logic level gap of any gate:
	gf_c880: 5
*/

module gf_c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n103;
	wire n104;
	wire n105;
	wire n107;
	wire n108;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n119;
	wire n120;
	wire n122;
	wire n123;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [2:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [1:0] w_G201gat_1;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [2:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [1:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [2:0] w_n95_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n113_0;
	wire [2:0] w_n119_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n144_0;
	wire [1:0] w_n146_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [1:0] w_n149_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n164_0;
	wire [2:0] w_n164_1;
	wire [2:0] w_n164_2;
	wire [1:0] w_n164_3;
	wire [1:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [2:0] w_n170_0;
	wire [1:0] w_n170_1;
	wire [1:0] w_n173_0;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n178_2;
	wire [1:0] w_n178_3;
	wire [2:0] w_n181_0;
	wire [1:0] w_n185_0;
	wire [2:0] w_n197_0;
	wire [2:0] w_n198_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [2:0] w_n219_0;
	wire [2:0] w_n222_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n234_0;
	wire [1:0] w_n235_0;
	wire [2:0] w_n239_0;
	wire [1:0] w_n239_1;
	wire [1:0] w_n240_0;
	wire [1:0] w_n241_0;
	wire [1:0] w_n242_0;
	wire [1:0] w_n245_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n258_0;
	wire [1:0] w_n260_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n267_0;
	wire [2:0] w_n285_0;
	wire [2:0] w_n303_0;
	wire [1:0] w_n303_1;
	wire [2:0] w_n306_0;
	wire [1:0] w_n306_1;
	wire [2:0] w_n311_0;
	wire [2:0] w_n311_1;
	wire [2:0] w_n319_0;
	wire [2:0] w_n319_1;
	wire [1:0] w_n320_0;
	wire [1:0] w_n321_0;
	wire [2:0] w_n327_0;
	wire [2:0] w_n327_1;
	wire [1:0] w_n328_0;
	wire [1:0] w_n329_0;
	wire [2:0] w_n335_0;
	wire [1:0] w_n335_1;
	wire [2:0] w_n336_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n346_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n352_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n361_0;
	wire [2:0] w_n377_0;
	wire [1:0] w_n391_0;
	wire [1:0] w_n393_0;
	wire [2:0] w_n404_0;
	wire [2:0] w_n420_0;
	wire w_dff_B_GSIaywte5_2;
	wire w_dff_B_tAReGijg0_1;
	wire w_dff_B_zHSEY54C2_1;
	wire w_dff_B_kiZvJ92o9_1;
	wire w_dff_A_xHbkrqDb3_1;
	wire w_dff_A_6u0KVS2n6_1;
	wire w_dff_B_p7UUrr9R3_1;
	wire w_dff_B_N3gDhnya0_1;
	wire w_dff_B_kggM7kW44_1;
	wire w_dff_B_qVLElNTY8_1;
	wire w_dff_B_rs6GoOFe1_1;
	wire w_dff_B_IYnRNLZA4_1;
	wire w_dff_B_CaTEttEE8_1;
	wire w_dff_A_VbHs2Mun8_1;
	wire w_dff_B_xZ4cSpAA9_1;
	wire w_dff_B_MsViwyTq7_1;
	wire w_dff_B_KBWPjDHB7_1;
	wire w_dff_B_lBXbOrwb0_1;
	wire w_dff_B_ZpbdFtNi8_1;
	wire w_dff_B_EPAe0jse5_1;
	wire w_dff_B_yeiXuvcf0_0;
	wire w_dff_B_UGuoYXmm1_0;
	wire w_dff_B_NiLdjS6E0_0;
	wire w_dff_B_iODpJsBp4_0;
	wire w_dff_B_CqEcUHpB6_0;
	wire w_dff_B_13NRcRbk2_0;
	wire w_dff_B_PRsgJq3f1_0;
	wire w_dff_B_ldYpc67U9_0;
	wire w_dff_B_qzjTKzz27_0;
	wire w_dff_B_4Awn7C4E9_0;
	wire w_dff_B_7yALASj83_0;
	wire w_dff_B_RU1Eypu97_0;
	wire w_dff_B_aDLR7Kvq2_0;
	wire w_dff_B_glchsX2h6_0;
	wire w_dff_A_lbbwU5MU8_0;
	wire w_dff_A_ovymAdQG1_0;
	wire w_dff_A_SmruBy2C7_0;
	wire w_dff_A_jJiEuFvK4_0;
	wire w_dff_B_KRXK0BIK7_1;
	wire w_dff_B_JS8AxjnQ2_1;
	wire w_dff_B_CcigUWsG8_1;
	wire w_dff_B_Y30hR4Xq7_1;
	wire w_dff_B_cmC4qDUJ6_1;
	wire w_dff_B_4rqCsIZw9_1;
	wire w_dff_B_fDhPSzWG5_1;
	wire w_dff_B_5tPrt5TS0_1;
	wire w_dff_B_DMUQEEkT6_1;
	wire w_dff_B_5RxU2FrA5_1;
	wire w_dff_B_dQ96iAXH6_1;
	wire w_dff_B_8yNUeOwK7_1;
	wire w_dff_B_7UJ5sV2m1_1;
	wire w_dff_B_6pSDPMc78_1;
	wire w_dff_B_7gnwILmQ9_1;
	wire w_dff_B_9AMMAbma1_1;
	wire w_dff_B_RMJa3JFY2_1;
	wire w_dff_B_V2HBIQJY9_1;
	wire w_dff_B_7TXgyzlL9_1;
	wire w_dff_B_jQkrUx4e0_1;
	wire w_dff_B_84n8DlGf3_1;
	wire w_dff_B_uIXJncuN6_0;
	wire w_dff_B_oVL95WD29_0;
	wire w_dff_B_BEQmc9da3_0;
	wire w_dff_B_mzBl8A180_0;
	wire w_dff_B_ff64FpwW7_0;
	wire w_dff_B_YFBtf0H28_0;
	wire w_dff_B_nqqmaY0D9_0;
	wire w_dff_B_7PLyaIN99_0;
	wire w_dff_A_EAMIyyQt3_1;
	wire w_dff_A_CXvq3uDD5_1;
	wire w_dff_A_RKnVw1t78_1;
	wire w_dff_A_LS30gOEK1_1;
	wire w_dff_A_XCbuhe4z0_1;
	wire w_dff_A_JtT7Xivj8_1;
	wire w_dff_A_YIUMp9I11_1;
	wire w_dff_A_qgTNje5x7_1;
	wire w_dff_A_HzVUopj19_1;
	wire w_dff_A_IaniZYls9_0;
	wire w_dff_A_o46JxSdL2_0;
	wire w_dff_A_8hignWYJ0_0;
	wire w_dff_A_SYl1ZTaK7_0;
	wire w_dff_A_foXrpMJg4_1;
	wire w_dff_A_QQFj4ndL4_1;
	wire w_dff_A_0uaWIG1l7_1;
	wire w_dff_A_NLAVdITU2_1;
	wire w_dff_A_ODHcvoO50_1;
	wire w_dff_A_dGtI2dac5_1;
	wire w_dff_A_84Y2JVtx4_1;
	wire w_dff_A_0099FcX74_1;
	wire w_dff_A_j14IaQH59_1;
	wire w_dff_B_tPIYVKvH9_1;
	wire w_dff_B_F0f1ClMC4_1;
	wire w_dff_B_A932LBmu1_1;
	wire w_dff_B_ijtp4fIJ1_1;
	wire w_dff_B_lTkxRn4p5_1;
	wire w_dff_B_FU6iXRqU8_1;
	wire w_dff_B_Hu5j9bju6_0;
	wire w_dff_B_TLrXwqyY7_0;
	wire w_dff_B_P7XkTJJ67_0;
	wire w_dff_B_JIUTpmJ50_0;
	wire w_dff_A_jO3Qq5u22_0;
	wire w_dff_A_I47TRL0K7_0;
	wire w_dff_A_cswhGIzL9_0;
	wire w_dff_A_aF2RwkzK0_1;
	wire w_dff_A_PVgGCB742_1;
	wire w_dff_A_HcTM1GVX3_1;
	wire w_dff_A_kEdOAhc04_1;
	wire w_dff_A_jC3o60vi7_1;
	wire w_dff_B_s73pqaah1_1;
	wire w_dff_B_nn6wMOGk0_0;
	wire w_dff_B_7cjJs6LO5_0;
	wire w_dff_B_20CebZ979_0;
	wire w_dff_B_6E7KgVIu3_0;
	wire w_dff_B_9r22lERW4_1;
	wire w_dff_B_OmeFB6pZ1_1;
	wire w_dff_B_H0zx1ZtW2_1;
	wire w_dff_B_3ZMkq8Hj4_1;
	wire w_dff_B_x3DtjL5f7_1;
	wire w_dff_B_1a2TZAgG4_1;
	wire w_dff_B_Y1cVy0MP9_1;
	wire w_dff_B_D8OM8Dun0_1;
	wire w_dff_B_nomCx90E8_1;
	wire w_dff_B_rBgMgBtT9_1;
	wire w_dff_B_WCr7dEsS6_1;
	wire w_dff_B_eALMfTKs8_1;
	wire w_dff_B_WS4odQnb5_0;
	wire w_dff_B_iQF6CmOP3_0;
	wire w_dff_B_eNyofXta8_0;
	wire w_dff_B_5LYf5VqB1_0;
	wire w_dff_B_mXgbvMDp2_0;
	wire w_dff_B_XpaDHBzu2_0;
	wire w_dff_A_ma28hyni2_1;
	wire w_dff_A_ryLF9ho38_1;
	wire w_dff_A_MICi2kaS5_1;
	wire w_dff_A_oPYePDtu1_1;
	wire w_dff_A_Ld9vuEK63_1;
	wire w_dff_B_sv0h8F5G0_1;
	wire w_dff_B_doZbIsdq4_1;
	wire w_dff_B_quorBJTR4_1;
	wire w_dff_B_FdyFEEuq6_1;
	wire w_dff_B_yFZnzdM23_0;
	wire w_dff_B_uQCll2v58_0;
	wire w_dff_B_uYfs2cxK6_1;
	wire w_dff_B_hQhrmT7l8_0;
	wire w_dff_B_vqXqbZSx8_0;
	wire w_dff_B_zCUSekvJ1_0;
	wire w_dff_B_9QPYehDS4_0;
	wire w_dff_B_pfDKVsB08_0;
	wire w_dff_B_N6L8NkBI2_0;
	wire w_dff_B_itdv4hEJ5_0;
	wire w_dff_B_pg4cL8EJ9_0;
	wire w_dff_B_A16QuiJk1_1;
	wire w_dff_B_D1GtwHkq2_1;
	wire w_dff_B_lbCEY3NP1_1;
	wire w_dff_B_TY17PhMk2_1;
	wire w_dff_B_BJwEZ6133_1;
	wire w_dff_B_dDcipXBN9_1;
	wire w_dff_B_6OVoBhBC5_1;
	wire w_dff_B_Cx9viwQK4_1;
	wire w_dff_B_KKr6Xmht4_0;
	wire w_dff_B_oFbHHbPU4_0;
	wire w_dff_B_IJ1xQlMV2_0;
	wire w_dff_B_XSdgvg7a2_0;
	wire w_dff_B_WGeQ4lVH4_0;
	wire w_dff_B_Cy6GudwD7_0;
	wire w_dff_A_A6pBvmPj2_1;
	wire w_dff_A_uSC7OrEy1_1;
	wire w_dff_A_KWSQz0Ql4_1;
	wire w_dff_B_Rbgx2vm75_1;
	wire w_dff_B_3eNKzKk52_1;
	wire w_dff_B_AzUGH2hI5_1;
	wire w_dff_B_ml8j43294_1;
	wire w_dff_B_VakEVg175_1;
	wire w_dff_B_20wcC6Ne3_1;
	wire w_dff_B_g8o3Zviv8_1;
	wire w_dff_B_5cFhrUcq6_1;
	wire w_dff_B_QKePrQ611_1;
	wire w_dff_B_ghwV2H0S0_1;
	wire w_dff_B_eJ50nooN0_1;
	wire w_dff_B_HEUlk5BE9_1;
	wire w_dff_B_voHXs2Qa4_1;
	wire w_dff_B_8r6bEAey5_1;
	wire w_dff_B_vSOUwK2N3_1;
	wire w_dff_B_efrgUlBb8_1;
	wire w_dff_B_fFyNbHDS8_1;
	wire w_dff_B_LbgnQHev8_1;
	wire w_dff_B_P8gRLnd94_1;
	wire w_dff_B_JeXEp6s22_1;
	wire w_dff_B_cK3e9Z3T8_1;
	wire w_dff_B_BUnj0QyW7_1;
	wire w_dff_B_0f3GhMrc8_1;
	wire w_dff_B_agPU4M1E7_1;
	wire w_dff_B_yxqbIcDq2_1;
	wire w_dff_B_RmIz27ih2_1;
	wire w_dff_B_TCubaHiW8_1;
	wire w_dff_B_Crsi5cq54_1;
	wire w_dff_B_G5W7pFqL9_1;
	wire w_dff_A_xVCbd2lf1_0;
	wire w_dff_A_HC0x09Pj9_0;
	wire w_dff_A_kR5YIjbe0_0;
	wire w_dff_A_ATAq18RA7_0;
	wire w_dff_A_568KjyB94_0;
	wire w_dff_A_DqioWgSz5_0;
	wire w_dff_A_es7kT23C2_0;
	wire w_dff_A_1BKxyyK10_0;
	wire w_dff_A_O8Vklup97_0;
	wire w_dff_A_DFUfRgTK0_1;
	wire w_dff_A_t2TQ3gLM1_1;
	wire w_dff_A_ULzcb9f16_1;
	wire w_dff_A_Exgb0kkr0_1;
	wire w_dff_A_LLlRukt87_1;
	wire w_dff_A_gnkWmC5J5_1;
	wire w_dff_A_Cz0Cu0aV2_1;
	wire w_dff_A_jFhtMyKy5_1;
	wire w_dff_A_5rMxZFOJ6_1;
	wire w_dff_B_GPhE9peD1_1;
	wire w_dff_B_dDZMWDgu2_1;
	wire w_dff_B_FN5MSQz78_0;
	wire w_dff_B_JOYH0Xz12_0;
	wire w_dff_B_FuOOvbjw1_0;
	wire w_dff_B_nhK3TEkx1_0;
	wire w_dff_B_YJfwExrU1_0;
	wire w_dff_B_1pV9Y5bC2_0;
	wire w_dff_B_oM4e1fGD4_0;
	wire w_dff_B_oYpqn9Si8_0;
	wire w_dff_B_KIQzMffs8_0;
	wire w_dff_B_45YLzm8C4_0;
	wire w_dff_B_t1lwdvkp9_0;
	wire w_dff_B_mCEZtpVI8_0;
	wire w_dff_B_3ejL3m9E0_0;
	wire w_dff_B_gpVBdfsV2_1;
	wire w_dff_B_3nLihxdL9_1;
	wire w_dff_B_1r9sycvd2_1;
	wire w_dff_B_C2QS22wE8_1;
	wire w_dff_A_59789IK71_0;
	wire w_dff_A_vxoLuX1Q7_0;
	wire w_dff_A_JhfWkjJ38_0;
	wire w_dff_A_7VJLBtPY3_0;
	wire w_dff_A_sGzLHVee3_0;
	wire w_dff_A_g8THXuPB6_0;
	wire w_dff_A_tNk60cMu8_0;
	wire w_dff_A_h4gHO2iu9_0;
	wire w_dff_A_eThL9HM11_0;
	wire w_dff_A_gDlbk4Ia6_0;
	wire w_dff_A_ch7dmcIp8_0;
	wire w_dff_A_2UGetOFz2_0;
	wire w_dff_A_u2asBRF63_0;
	wire w_dff_A_MSP3JsP91_0;
	wire w_dff_A_Fb5zEkqL0_0;
	wire w_dff_A_zu6g0c7R2_0;
	wire w_dff_A_1LorvZwg6_0;
	wire w_dff_A_Gs7sp7nX6_0;
	wire w_dff_A_lBzLUwpW9_0;
	wire w_dff_A_G51sbAmz5_0;
	wire w_dff_A_nDEMpseI7_0;
	wire w_dff_A_BUhkNS0b3_0;
	wire w_dff_A_tIFLXirb2_0;
	wire w_dff_A_Oe9a0CGt2_0;
	wire w_dff_A_REtwFYfb2_0;
	wire w_dff_A_XYTdUqX19_0;
	wire w_dff_A_W48Xm7nX1_0;
	wire w_dff_A_XHTaupih4_0;
	wire w_dff_B_n2gwc0Wj5_1;
	wire w_dff_B_b8rYDj6P0_1;
	wire w_dff_B_3TSyV1bV3_1;
	wire w_dff_B_GuAntEwq1_1;
	wire w_dff_B_j7SlwgB99_1;
	wire w_dff_B_kh9VxO0k5_1;
	wire w_dff_B_ndfcPuaT1_1;
	wire w_dff_B_bYpKujEX4_1;
	wire w_dff_A_bJ3daH7s7_0;
	wire w_dff_A_FFFIshbQ3_0;
	wire w_dff_A_qtemNoQF6_0;
	wire w_dff_A_GArnw1Hh2_0;
	wire w_dff_A_veE51J5r6_0;
	wire w_dff_A_sidqFTyr6_1;
	wire w_dff_A_q8r5PICu7_1;
	wire w_dff_A_MoxOgXXi2_1;
	wire w_dff_A_5ThYq8HY6_1;
	wire w_dff_A_HdP8i38R0_1;
	wire w_dff_A_tSxS8ex92_0;
	wire w_dff_A_9HdxmpXx7_0;
	wire w_dff_A_k2Q75X6R6_0;
	wire w_dff_A_7iYUx3bS4_0;
	wire w_dff_A_c2ulKy9Q7_0;
	wire w_dff_A_zxLR4eFD5_0;
	wire w_dff_A_MuNfmDZT5_0;
	wire w_dff_A_LCf2uBmQ9_0;
	wire w_dff_A_9Z1wnDuS3_0;
	wire w_dff_A_WTmwzHhH3_0;
	wire w_dff_B_70CWGrjI8_1;
	wire w_dff_B_K4KwPQzj4_1;
	wire w_dff_B_elh2Lk664_1;
	wire w_dff_B_QJXJPvJC7_1;
	wire w_dff_B_JcgMogmf8_1;
	wire w_dff_B_TAxAW1TE0_1;
	wire w_dff_B_p6qSeAFm5_1;
	wire w_dff_B_UBdkgCNo1_1;
	wire w_dff_B_3TIzWT7q7_1;
	wire w_dff_B_jllHzEmu8_1;
	wire w_dff_B_dZ8btkFc7_1;
	wire w_dff_B_ZJiliUBo6_1;
	wire w_dff_B_ijMSrt5x0_1;
	wire w_dff_B_mfXSlU7j1_1;
	wire w_dff_B_gjEntSGG0_0;
	wire w_dff_B_TtY3cPI91_0;
	wire w_dff_B_eeKoyiNY8_0;
	wire w_dff_B_0UUyqVNO3_0;
	wire w_dff_B_nS0kYOT68_0;
	wire w_dff_B_LavBUcDn8_0;
	wire w_dff_B_x7scORUO7_0;
	wire w_dff_B_bnIP7UBA7_0;
	wire w_dff_B_dEFVNWWr4_0;
	wire w_dff_B_E5dNJnVk6_0;
	wire w_dff_B_ekhsX9qf0_0;
	wire w_dff_B_zyDzmDZh4_0;
	wire w_dff_B_1H8axePV9_0;
	wire w_dff_B_fp7LMI6Y1_1;
	wire w_dff_B_2NjnirCd9_1;
	wire w_dff_B_ecR09ZOB4_1;
	wire w_dff_B_bRMTJVsK4_1;
	wire w_dff_B_y3lGjh756_1;
	wire w_dff_B_jU7pNuAJ5_1;
	wire w_dff_B_WFd4YglH5_1;
	wire w_dff_B_Di7pQTo20_1;
	wire w_dff_B_OBxQareG3_1;
	wire w_dff_B_dcIdBJQX2_1;
	wire w_dff_B_yueMlWGZ3_1;
	wire w_dff_B_YkK2LiLL9_1;
	wire w_dff_B_aHvNFreD1_1;
	wire w_dff_B_CSXGgycY4_1;
	wire w_dff_B_Up8wcUm81_1;
	wire w_dff_B_xRKcFhbq1_1;
	wire w_dff_B_jubtWu7l6_1;
	wire w_dff_B_kSzUQxZW4_1;
	wire w_dff_B_O0Co4cgu7_1;
	wire w_dff_B_N6UCPSSF5_1;
	wire w_dff_B_aKNoyOfg5_1;
	wire w_dff_B_eDgVJC478_1;
	wire w_dff_B_ORnpkLBA5_1;
	wire w_dff_A_SPd4hQoH9_1;
	wire w_dff_A_alXJXg7B6_1;
	wire w_dff_A_dHrcjvzZ0_1;
	wire w_dff_A_5zOnVWgp5_1;
	wire w_dff_A_WtDQ0C6I6_1;
	wire w_dff_A_MN2wCX0R6_1;
	wire w_dff_A_kiWtPUaK0_1;
	wire w_dff_A_kDsYcmTD4_1;
	wire w_dff_A_S0lkKPoz1_1;
	wire w_dff_A_k27b6J7i0_1;
	wire w_dff_A_xpGovbfh8_1;
	wire w_dff_A_uy3vY4jq6_1;
	wire w_dff_A_i3iRedDT1_1;
	wire w_dff_A_Vtb3yNv80_1;
	wire w_dff_A_NB21JOM31_1;
	wire w_dff_A_8FnFl0Ka1_1;
	wire w_dff_A_Bfh220527_1;
	wire w_dff_A_Bd3YpNBu6_1;
	wire w_dff_A_L2jm9TSj8_1;
	wire w_dff_A_RzrELDkc0_1;
	wire w_dff_A_5DNRdYme2_1;
	wire w_dff_A_rwqahejY1_1;
	wire w_dff_A_Wm0Jxyom7_1;
	wire w_dff_A_P7w0ZNjN8_1;
	wire w_dff_A_pcKRiF3c5_1;
	wire w_dff_A_f0Tnz2Rf4_0;
	wire w_dff_A_hYU0cSRm4_0;
	wire w_dff_A_IKgKATdn5_0;
	wire w_dff_A_0392metA6_0;
	wire w_dff_A_hfHBCBrd4_0;
	wire w_dff_A_mwI5hC6T4_0;
	wire w_dff_A_BjfqaBXx3_0;
	wire w_dff_A_e8Ofl2I68_0;
	wire w_dff_A_C391u25s3_1;
	wire w_dff_A_zPqbXuor2_1;
	wire w_dff_A_cx3u6k8U7_1;
	wire w_dff_A_EZKn2qb88_1;
	wire w_dff_A_Rm1vi7Dm2_1;
	wire w_dff_A_T6MFeb4P1_1;
	wire w_dff_A_Ubtbp1NT0_1;
	wire w_dff_A_gCsMnsrE5_1;
	wire w_dff_B_TnSxArNL8_1;
	wire w_dff_B_KipvtkXk5_0;
	wire w_dff_B_dhwGUi4C4_0;
	wire w_dff_B_MHrCsJvJ9_0;
	wire w_dff_B_CpbJkFt88_0;
	wire w_dff_B_HtzshIPQ6_0;
	wire w_dff_B_Its1ghR50_0;
	wire w_dff_B_qBnUhGcF5_0;
	wire w_dff_B_7sJIehnG8_0;
	wire w_dff_B_3ohoTttX1_0;
	wire w_dff_B_BYWnBMy53_0;
	wire w_dff_B_VrBGeUMi8_0;
	wire w_dff_B_bwf0huTv8_0;
	wire w_dff_A_7ATrk8lA0_1;
	wire w_dff_A_fI0k704R3_1;
	wire w_dff_A_FTX2Vn1G9_1;
	wire w_dff_A_oTX2lA851_1;
	wire w_dff_A_6elblald0_1;
	wire w_dff_A_wOf0Vs3J2_1;
	wire w_dff_A_rEdaWlZD6_1;
	wire w_dff_A_wpFhUrYf7_1;
	wire w_dff_A_1zoxcUQz6_1;
	wire w_dff_A_5uR6ew4C1_1;
	wire w_dff_A_PzTRTfC43_1;
	wire w_dff_A_QWIExkVG9_1;
	wire w_dff_A_xHEuLEKk9_1;
	wire w_dff_A_L9BAJdW84_1;
	wire w_dff_B_CLxBbHRk0_1;
	wire w_dff_B_mE57rEnW3_0;
	wire w_dff_B_JyLV2Q8U5_0;
	wire w_dff_B_iqj695lP5_0;
	wire w_dff_B_I7u5Bzyw3_0;
	wire w_dff_B_hAr2lqVH2_0;
	wire w_dff_B_gNuOt0Qh5_0;
	wire w_dff_B_mf2zHNDT5_1;
	wire w_dff_A_RPvBiwtN1_1;
	wire w_dff_A_AhNfZjqw4_1;
	wire w_dff_A_ii5jO80d8_1;
	wire w_dff_A_FRKPHSb78_1;
	wire w_dff_A_xfzsnMIv6_1;
	wire w_dff_A_BAHIDpAU2_1;
	wire w_dff_A_KrKVBosd4_1;
	wire w_dff_A_mztmAX8J0_1;
	wire w_dff_A_Cdh1RHdS9_1;
	wire w_dff_A_Lq5lGMV70_2;
	wire w_dff_A_mS6P4vMk2_2;
	wire w_dff_A_zjTxZgD94_2;
	wire w_dff_A_D4q2zQEj8_2;
	wire w_dff_A_OiQ2ftAf5_2;
	wire w_dff_A_LA9QaM5A7_2;
	wire w_dff_A_U6k3qrq82_2;
	wire w_dff_A_l6nWrpZy7_2;
	wire w_dff_A_WIZqdezD2_2;
	wire w_dff_A_Gj1DOGlz4_2;
	wire w_dff_A_ooxJvQMe3_2;
	wire w_dff_B_IxmWWaaA2_1;
	wire w_dff_B_6niYvNzb6_1;
	wire w_dff_B_Kpy8p9277_1;
	wire w_dff_B_Fr1O2fo07_1;
	wire w_dff_B_o3W47Yud8_1;
	wire w_dff_B_ZQQbyMHB4_1;
	wire w_dff_B_SpTcmguP0_1;
	wire w_dff_B_ThYCInlC6_1;
	wire w_dff_B_TgmfaMBk4_1;
	wire w_dff_B_8fNxos089_1;
	wire w_dff_B_b77xlsdY5_1;
	wire w_dff_B_mebxrYF86_1;
	wire w_dff_B_5sJrgmDu4_0;
	wire w_dff_B_1pydwt8Y6_0;
	wire w_dff_B_BzkI7QOS5_0;
	wire w_dff_B_ObuiwlhG6_0;
	wire w_dff_B_uQgBBIEg4_0;
	wire w_dff_B_mi3XB9ba4_0;
	wire w_dff_B_P6C7vMeD7_0;
	wire w_dff_B_VKR7baJS2_0;
	wire w_dff_B_D9jll0ar0_0;
	wire w_dff_B_6pyf0hvZ3_0;
	wire w_dff_B_2CBrTZA57_0;
	wire w_dff_B_UZNijE2z1_1;
	wire w_dff_B_3LU1e96R4_1;
	wire w_dff_B_XRT4DgV51_1;
	wire w_dff_B_YLPxsV2m2_1;
	wire w_dff_B_eF1gTHkW1_1;
	wire w_dff_B_E0dRo7Ap4_1;
	wire w_dff_B_pwYc6g3t5_1;
	wire w_dff_B_1LJfeufW8_1;
	wire w_dff_B_0NfAE29N8_1;
	wire w_dff_B_BPEUKfMy0_1;
	wire w_dff_B_oEAOUbTH8_1;
	wire w_dff_B_gJRVFlMj1_1;
	wire w_dff_B_E5vJf1TA7_1;
	wire w_dff_B_PQc7fllE3_1;
	wire w_dff_B_9ixuTAQ49_1;
	wire w_dff_B_UtgkDoeP8_1;
	wire w_dff_B_qejEdbeU3_1;
	wire w_dff_B_rmn6hfnz2_1;
	wire w_dff_B_A3NTip0I7_1;
	wire w_dff_A_d2q87DtS4_1;
	wire w_dff_A_XFTT5lTa1_1;
	wire w_dff_A_DAZQY4LC8_1;
	wire w_dff_A_rxU9HR7l9_1;
	wire w_dff_A_NFzSnkBu4_1;
	wire w_dff_A_hzmtlQNW0_1;
	wire w_dff_A_XLbgnOm52_1;
	wire w_dff_A_TBEbmUIM3_1;
	wire w_dff_A_92L2Is1y1_1;
	wire w_dff_A_g1NKNY736_1;
	wire w_dff_A_9ojVpIRN3_1;
	wire w_dff_A_08R7Lev64_1;
	wire w_dff_A_WdjsqJVn3_1;
	wire w_dff_A_n8CJ7ICn0_1;
	wire w_dff_A_R8Vs0EG03_1;
	wire w_dff_A_mV0FOiNZ9_1;
	wire w_dff_A_CMxlevNE6_1;
	wire w_dff_A_RUTyJ0s48_1;
	wire w_dff_A_MM3tbpEL4_1;
	wire w_dff_A_l4Ds0gqY9_1;
	wire w_dff_A_GAhtxgvl0_1;
	wire w_dff_A_yf3Es2g00_0;
	wire w_dff_A_USrduznW5_0;
	wire w_dff_A_RyCpXcoG7_0;
	wire w_dff_A_RlEP8WcD4_0;
	wire w_dff_A_19Wqj0xR3_0;
	wire w_dff_A_LfoXiNxK0_0;
	wire w_dff_A_5l1pAPm48_0;
	wire w_dff_A_XRapL5ry9_0;
	wire w_dff_A_5UnxKDUu8_0;
	wire w_dff_A_ppOcJGmE8_1;
	wire w_dff_A_pioUJZBQ7_1;
	wire w_dff_A_JYwpyw1R4_1;
	wire w_dff_A_Xyx0mOje4_1;
	wire w_dff_A_OzXuUR4n4_1;
	wire w_dff_A_4Fo6cjNh2_1;
	wire w_dff_A_TS9LzjdN2_1;
	wire w_dff_A_yrGGfm964_1;
	wire w_dff_A_SDHk0Ayh3_1;
	wire w_dff_B_em656vaO0_1;
	wire w_dff_B_LNaa5wLb6_0;
	wire w_dff_B_6GQCrwjA3_0;
	wire w_dff_B_0VR8D4NB0_0;
	wire w_dff_B_LH3CBpk42_0;
	wire w_dff_B_Qr1Exhr47_0;
	wire w_dff_B_vXtvioYj5_0;
	wire w_dff_B_WNAWS9qW8_0;
	wire w_dff_B_BWDOHGqr9_0;
	wire w_dff_B_LAuNqCAH6_0;
	wire w_dff_B_ZlYS1TIf0_0;
	wire w_dff_B_8yfsx2nm3_0;
	wire w_dff_B_wTQ1267p5_0;
	wire w_dff_A_YiYdZcsI5_1;
	wire w_dff_A_lIdggpTg7_1;
	wire w_dff_A_Bx15hbLn1_1;
	wire w_dff_A_z2n6usdp9_1;
	wire w_dff_A_hHT4DfCN8_1;
	wire w_dff_A_pSUFoYvh7_1;
	wire w_dff_A_BcMDqKgm5_1;
	wire w_dff_A_SCgwyVPp8_1;
	wire w_dff_A_86jZxEJm1_1;
	wire w_dff_A_iFAjw0GP6_1;
	wire w_dff_A_BvksVKM82_1;
	wire w_dff_A_zHL6klVf2_1;
	wire w_dff_A_ogtdX02Z2_1;
	wire w_dff_A_f7gAH5oF8_1;
	wire w_dff_A_lcXQg14O7_1;
	wire w_dff_A_FodcDkDs4_1;
	wire w_dff_A_JJoZkWO27_1;
	wire w_dff_A_Xa5F2hGi1_1;
	wire w_dff_B_py9DwAIB7_0;
	wire w_dff_B_ME3aqBur3_0;
	wire w_dff_B_FGhC9g0D4_0;
	wire w_dff_B_8IAzCC8t9_0;
	wire w_dff_B_sDlKO3YR9_0;
	wire w_dff_A_aNQIUORM4_0;
	wire w_dff_A_6ZGK6Eos5_0;
	wire w_dff_A_f16D6L1E6_1;
	wire w_dff_A_VMDtzSMh3_1;
	wire w_dff_A_2H6Iw6yB7_1;
	wire w_dff_A_di2SfrFP5_1;
	wire w_dff_A_ugTcDXZo3_1;
	wire w_dff_A_ZzoTFIye8_1;
	wire w_dff_A_pfeKiM682_1;
	wire w_dff_A_D05oNxKZ1_1;
	wire w_dff_A_gV8tk6AY7_2;
	wire w_dff_A_FCaw76er3_2;
	wire w_dff_A_ZTSQR2WJ0_2;
	wire w_dff_A_6KPCu3Km9_2;
	wire w_dff_A_ItNotLYK3_2;
	wire w_dff_A_wwwFtVNb1_2;
	wire w_dff_A_38dpMtXr9_2;
	wire w_dff_A_md0ncrWr1_2;
	wire w_dff_A_BTy1ECCB1_2;
	wire w_dff_A_ZuaxcF6B6_2;
	wire w_dff_B_epr6vjWz6_3;
	wire w_dff_B_TjZuYqWm5_1;
	wire w_dff_B_RQ8n5l5u4_1;
	wire w_dff_B_8YmqLXfr9_1;
	wire w_dff_B_SsrziKMG3_1;
	wire w_dff_B_9DIcCkY60_1;
	wire w_dff_B_nUPNL3Do2_1;
	wire w_dff_B_7T0nKnwn6_1;
	wire w_dff_B_Ypdj6s0X1_1;
	wire w_dff_B_lvNTZ2L67_1;
	wire w_dff_B_EwFU9vN70_1;
	wire w_dff_B_W3z3T0lt7_1;
	wire w_dff_B_YvFDfzdB1_1;
	wire w_dff_B_OXuQGpJw2_1;
	wire w_dff_B_6DpSRe6W7_1;
	wire w_dff_B_pcnzQFld0_1;
	wire w_dff_B_8Q9L2Ugr5_1;
	wire w_dff_B_GmmfPo5h3_1;
	wire w_dff_B_EY4aSTkf0_1;
	wire w_dff_B_yoby2iPW5_1;
	wire w_dff_B_id5kLjQl1_1;
	wire w_dff_B_vbu4v1jM8_1;
	wire w_dff_B_rl9Vq7JE8_0;
	wire w_dff_A_rWOHNZkG3_1;
	wire w_dff_A_sqprAlgC0_1;
	wire w_dff_A_lslrCMJR3_2;
	wire w_dff_A_UUauDlHl2_2;
	wire w_dff_A_QObBHfh02_2;
	wire w_dff_A_4Sd4npID9_2;
	wire w_dff_A_O1Lucx3I5_0;
	wire w_dff_A_uzqWPfXI1_0;
	wire w_dff_A_a1FPNMpL1_0;
	wire w_dff_A_asF04T9x1_0;
	wire w_dff_A_edw16gTV5_0;
	wire w_dff_A_kOUkT3XB5_0;
	wire w_dff_A_jtlU4Qz41_0;
	wire w_dff_A_yV2b8S5z8_0;
	wire w_dff_A_SfnO8thz7_0;
	wire w_dff_A_sMiNjPDH1_1;
	wire w_dff_B_PLaI4vFA4_3;
	wire w_dff_B_UIDBElnm6_3;
	wire w_dff_B_wqnAYARH5_3;
	wire w_dff_B_BfeD4erD1_3;
	wire w_dff_B_R9hstALJ1_3;
	wire w_dff_B_o3Pi5RmB4_3;
	wire w_dff_B_ptPcvAMe1_3;
	wire w_dff_B_q7NuIUaE4_3;
	wire w_dff_B_2xljmZZE0_3;
	wire w_dff_B_R3Xi5MM07_3;
	wire w_dff_B_cexpfoTi9_3;
	wire w_dff_B_kEi3TNjC8_3;
	wire w_dff_B_9wLbiQPo5_0;
	wire w_dff_B_KjaHok4l3_0;
	wire w_dff_B_CgkK8ZDX5_0;
	wire w_dff_B_cvEIrjfx2_0;
	wire w_dff_B_onPodhm80_0;
	wire w_dff_B_csD3o8sT0_0;
	wire w_dff_B_TnQ6bYOD9_0;
	wire w_dff_B_WB2r8z254_0;
	wire w_dff_B_bOfGwb3m3_0;
	wire w_dff_B_WSMxIz7D4_1;
	wire w_dff_B_xeCAAGe97_1;
	wire w_dff_B_wPr6t00I9_1;
	wire w_dff_B_oQvKxCeK5_1;
	wire w_dff_B_rBwTdNrd7_1;
	wire w_dff_B_MIa4ORsT9_1;
	wire w_dff_B_eALyMLm19_1;
	wire w_dff_B_9YbA9GZ99_1;
	wire w_dff_B_2niJCX933_1;
	wire w_dff_B_2tdBkyD23_1;
	wire w_dff_B_L7mGhCgb8_1;
	wire w_dff_B_YBwhKsRa3_1;
	wire w_dff_B_NjjmpL1C0_1;
	wire w_dff_B_axRcZCmb1_1;
	wire w_dff_B_Y9ex9KpT5_1;
	wire w_dff_B_qKC3uJD64_1;
	wire w_dff_B_VXLgkgsg4_1;
	wire w_dff_B_IGXkI59T7_1;
	wire w_dff_B_ZEdnkMpZ5_1;
	wire w_dff_B_XRitnMuY1_1;
	wire w_dff_B_BjzQLaOI5_1;
	wire w_dff_B_YfHJEGy66_1;
	wire w_dff_B_EXS4HU1R9_1;
	wire w_dff_B_a0X6tw2p1_1;
	wire w_dff_B_LVXLDEJp9_1;
	wire w_dff_B_5z8THAnV5_1;
	wire w_dff_B_E84IDsFC6_1;
	wire w_dff_B_a8bqaFgB0_1;
	wire w_dff_B_E40CS4Av2_1;
	wire w_dff_A_r3WANGgp2_1;
	wire w_dff_B_TcBGh5e38_2;
	wire w_dff_B_GZI1XtSJ9_2;
	wire w_dff_B_qJeypqZ09_2;
	wire w_dff_B_GdrfCwyA0_2;
	wire w_dff_B_gjPcV6FL6_2;
	wire w_dff_B_Od2j9ylF8_2;
	wire w_dff_B_hmAaJchv4_2;
	wire w_dff_B_yM4KmRWJ9_2;
	wire w_dff_B_OnztqHNG8_2;
	wire w_dff_A_3MnImfhx0_0;
	wire w_dff_A_hbDEDvy40_0;
	wire w_dff_A_96Mgs9Aq8_0;
	wire w_dff_A_URHxRA7b2_0;
	wire w_dff_A_5gUO1yCr0_0;
	wire w_dff_A_LAyl2Q3X3_0;
	wire w_dff_A_AhYmlxv09_0;
	wire w_dff_A_dGt58nX79_0;
	wire w_dff_A_GVhlbfMO6_0;
	wire w_dff_A_ccCzQTdh6_0;
	wire w_dff_A_xhCMx9Wp1_2;
	wire w_dff_A_gQCTnKEc5_2;
	wire w_dff_A_Oo3s6GkZ7_2;
	wire w_dff_A_Utk7lrqA7_2;
	wire w_dff_A_HNm7eEoG8_2;
	wire w_dff_A_zV5pQmm24_2;
	wire w_dff_A_mPWFUcQR4_2;
	wire w_dff_A_QeE2dAfw5_2;
	wire w_dff_A_GcNMlFBW8_2;
	wire w_dff_A_TBAA5QPO6_2;
	wire w_dff_A_DB211iR03_0;
	wire w_dff_B_f9PFycb75_1;
	wire w_dff_B_02REkNbb6_1;
	wire w_dff_B_y2AXDNAR1_1;
	wire w_dff_B_7CUkmzZD5_1;
	wire w_dff_B_ObvjXfyc0_1;
	wire w_dff_B_kvx6MqsJ7_1;
	wire w_dff_B_HnluH0Uh6_1;
	wire w_dff_B_901NAY6l2_1;
	wire w_dff_B_XmavlbES5_1;
	wire w_dff_B_hKw61krO9_1;
	wire w_dff_B_jn0YtmUD9_1;
	wire w_dff_B_BJriCuaR1_1;
	wire w_dff_A_dU3YKqVA4_1;
	wire w_dff_A_7iacd3fw9_1;
	wire w_dff_A_HyAzXTRm3_1;
	wire w_dff_A_7HQPvZec9_1;
	wire w_dff_A_RGLzaIRm5_1;
	wire w_dff_A_IxPp00Gn2_1;
	wire w_dff_B_0z4F70Dg9_3;
	wire w_dff_B_Ythl7dYS6_3;
	wire w_dff_B_WZmIcOnv1_3;
	wire w_dff_B_xcZpoV7G9_3;
	wire w_dff_B_Mh9Rh9t26_3;
	wire w_dff_B_AyRVInel9_3;
	wire w_dff_B_zrgDDyU05_3;
	wire w_dff_B_juyi9VzG8_3;
	wire w_dff_A_WAOntSsh3_1;
	wire w_dff_A_PKGxXbie3_1;
	wire w_dff_A_SnGcm0yV3_1;
	wire w_dff_A_eT09wCdN9_1;
	wire w_dff_A_lyUuIx8R6_1;
	wire w_dff_A_9ZGB39M65_1;
	wire w_dff_A_VkU8dekx9_1;
	wire w_dff_A_25R4wEmD7_1;
	wire w_dff_A_DVUZWOLC3_1;
	wire w_dff_A_ZsvT9tFg9_1;
	wire w_dff_A_vnB3XQGd9_1;
	wire w_dff_A_HtD9ivyS4_1;
	wire w_dff_A_X388gADN1_1;
	wire w_dff_A_nFZrfz888_1;
	wire w_dff_A_75Z0Ttk17_1;
	wire w_dff_A_JkpUGZBf2_1;
	wire w_dff_A_Piy7sRBc7_1;
	wire w_dff_A_bI3C978E9_1;
	wire w_dff_A_DZOh1sNt7_1;
	wire w_dff_A_TKBNZ3Sl1_1;
	wire w_dff_A_oB8wX8y63_2;
	wire w_dff_A_KD6KpCBg7_2;
	wire w_dff_A_TyLearqF5_2;
	wire w_dff_A_dHwoZXZW7_2;
	wire w_dff_A_GldfbQnw1_2;
	wire w_dff_A_YhlLimJq7_2;
	wire w_dff_A_0L2Xkrqe9_2;
	wire w_dff_A_FKwPJQjV2_2;
	wire w_dff_A_RcHTt1r62_1;
	wire w_dff_A_Q4NqfTz41_1;
	wire w_dff_A_LfhSIsyo9_1;
	wire w_dff_A_P4zV80J80_1;
	wire w_dff_A_zB6Gv0j14_0;
	wire w_dff_A_4TbRHPQ64_0;
	wire w_dff_A_K2ZbbhQx8_0;
	wire w_dff_A_DGPwAcHs4_0;
	wire w_dff_A_PdUsLsWK7_0;
	wire w_dff_A_2O2Q4pOl4_0;
	wire w_dff_A_4e58sPPQ2_0;
	wire w_dff_A_vAJMRL0o8_0;
	wire w_dff_A_e8keUhLf1_0;
	wire w_dff_A_yBKCEkH24_0;
	wire w_dff_A_XjCVYkKl7_0;
	wire w_dff_A_SKoyFyBL6_0;
	wire w_dff_A_a1EvICEe9_0;
	wire w_dff_A_gzSCnwQh6_0;
	wire w_dff_A_58KEmVE42_2;
	wire w_dff_A_Gz0ZKhMP3_2;
	wire w_dff_A_hsRqyjQF2_2;
	wire w_dff_A_7I1OU8ZZ1_2;
	wire w_dff_A_HQIrl6Va9_1;
	wire w_dff_A_T7BVjZmB1_1;
	wire w_dff_A_KorqsZZp3_1;
	wire w_dff_A_KtvHNEcG6_1;
	wire w_dff_A_CB2CKF6I5_1;
	wire w_dff_A_H6T3bKCf7_1;
	wire w_dff_A_68Es0FZV4_1;
	wire w_dff_A_iIdqfS259_1;
	wire w_dff_A_mW1Fgj0O8_1;
	wire w_dff_A_panc784W4_1;
	wire w_dff_A_mkV3RWMw8_1;
	wire w_dff_A_0RWsyMFv1_1;
	wire w_dff_A_JQ4JKKZN3_1;
	wire w_dff_A_3kGgvMV84_2;
	wire w_dff_A_gFPaDQdq1_2;
	wire w_dff_A_zjrh4Zhi9_2;
	wire w_dff_A_N1dGASNL1_2;
	wire w_dff_A_Qeh2TP0d5_2;
	wire w_dff_A_TiRiaqpM7_2;
	wire w_dff_A_fJHNsO0G1_2;
	wire w_dff_A_BONYvIGV9_2;
	wire w_dff_A_biPzaajY5_1;
	wire w_dff_A_CdGEj5VR7_1;
	wire w_dff_A_xeuZn17I5_1;
	wire w_dff_A_UucWkXq47_1;
	wire w_dff_A_3lnmUeB01_1;
	wire w_dff_A_k3roUDba9_1;
	wire w_dff_A_RgrZBGyU8_1;
	wire w_dff_B_43DQC57i3_2;
	wire w_dff_B_XqQFUiyg4_2;
	wire w_dff_B_dQhxHCWz2_2;
	wire w_dff_B_ELVxRGg83_2;
	wire w_dff_A_6nBN1ogq9_1;
	wire w_dff_A_ROKh5EhK0_1;
	wire w_dff_A_1kIFFkiw8_1;
	wire w_dff_A_gw22SdBI6_1;
	wire w_dff_A_cYPOGd2v4_1;
	wire w_dff_A_d6biRXab9_1;
	wire w_dff_A_CRKecSso3_0;
	wire w_dff_A_T6ccq5hL7_0;
	wire w_dff_A_p5d4la7a7_0;
	wire w_dff_A_J9Wi2rGg5_0;
	wire w_dff_A_Yf6uo45Z9_0;
	wire w_dff_A_xCZKXQlo2_0;
	wire w_dff_A_6wM7kc4N2_0;
	wire w_dff_A_15PxcqHD1_0;
	wire w_dff_A_zOXzmiA46_2;
	wire w_dff_A_ptCLX6vO7_2;
	wire w_dff_A_IKVk7OZN7_2;
	wire w_dff_A_OWu9GO5M9_2;
	wire w_dff_A_EGJT6SzF8_0;
	wire w_dff_A_vpcGVEZ13_0;
	wire w_dff_A_zljUsMXi2_0;
	wire w_dff_A_DdnYctoD0_0;
	wire w_dff_A_wAhB5Dpr9_0;
	wire w_dff_A_SfACn2Ng8_0;
	wire w_dff_B_17GVwLMI4_1;
	wire w_dff_B_NXo4Vcax5_1;
	wire w_dff_B_pklLYb6D2_1;
	wire w_dff_B_zMH2pYu61_1;
	wire w_dff_B_Xnfmz8m85_1;
	wire w_dff_B_IsHlgTDw1_1;
	wire w_dff_B_rYhg64yR0_1;
	wire w_dff_B_THrVAbF30_1;
	wire w_dff_A_7s7pj6yq6_1;
	wire w_dff_A_4CdHw3xI2_1;
	wire w_dff_A_IKaGLcQx4_1;
	wire w_dff_A_yX7WiixN2_1;
	wire w_dff_A_w0TsZFF95_1;
	wire w_dff_A_hFE75WfB3_1;
	wire w_dff_A_QCIoRFPs4_1;
	wire w_dff_A_uyfWmlS52_1;
	wire w_dff_A_nQJVdCYi2_0;
	wire w_dff_A_QqjlHKmk1_0;
	wire w_dff_A_6GAsQtzw5_0;
	wire w_dff_A_PH8TGeuR4_1;
	wire w_dff_B_ckQ37O4F2_2;
	wire w_dff_B_tJWrjoTV0_2;
	wire w_dff_B_pvufKJtW7_2;
	wire w_dff_B_65QB3twe0_2;
	wire w_dff_A_x0AiMJPD2_2;
	wire w_dff_A_yVEYHzL20_2;
	wire w_dff_A_zd94hS645_1;
	wire w_dff_A_XFB29Rx80_1;
	wire w_dff_A_0ss6Ng1O9_1;
	wire w_dff_A_z2blFpm61_1;
	wire w_dff_A_bjp8xU1K8_1;
	wire w_dff_A_cThWVYcY6_1;
	wire w_dff_A_QqaogmRE3_2;
	wire w_dff_A_gRlOYoRF9_2;
	wire w_dff_A_0EMUVmRj6_2;
	wire w_dff_A_soEfiLC39_2;
	wire w_dff_A_RJlScyza6_2;
	wire w_dff_A_pOLLdz346_2;
	wire w_dff_A_3Cz6OzwJ3_2;
	wire w_dff_A_54e5qKsY5_2;
	wire w_dff_A_w73sto869_0;
	wire w_dff_A_pwpjSjNC8_0;
	wire w_dff_A_paMU3kcr5_0;
	wire w_dff_A_DhIYGIoK8_0;
	wire w_dff_A_zFIWgomP6_0;
	wire w_dff_A_p742Ppg74_0;
	wire w_dff_A_lyr1kNRw7_0;
	wire w_dff_B_BHrdnGlM6_1;
	wire w_dff_B_GWM0xa6L8_1;
	wire w_dff_B_T713Ti4e7_1;
	wire w_dff_B_2JnXiDwJ0_1;
	wire w_dff_B_j8ejU5395_1;
	wire w_dff_B_1BnI7T5Q0_1;
	wire w_dff_B_TBWOYx9H7_1;
	wire w_dff_B_GQdyiRzL9_1;
	wire w_dff_B_zRWcyhoV2_1;
	wire w_dff_A_iaarpLbz1_2;
	wire w_dff_A_aeWtvHSd9_2;
	wire w_dff_A_siMNGYZJ1_2;
	wire w_dff_A_szMHMi966_2;
	wire w_dff_A_j8R3cMdQ2_2;
	wire w_dff_A_DPPJxwXO3_2;
	wire w_dff_A_qyfsu4mV1_2;
	wire w_dff_A_wzlfTpSR4_2;
	wire w_dff_A_SexcC3WA1_2;
	wire w_dff_B_6GSYaz0e9_0;
	wire w_dff_B_XR90HrZC3_0;
	wire w_dff_B_eOwpGUK18_0;
	wire w_dff_B_4eSsaiJV7_0;
	wire w_dff_B_Kn1FYWoV5_0;
	wire w_dff_A_X3qLaOM47_0;
	wire w_dff_A_2meL8y736_0;
	wire w_dff_A_64HgHN3Q9_0;
	wire w_dff_A_fWbf8oFC2_0;
	wire w_dff_A_1tJh7omA6_2;
	wire w_dff_A_wqRgMnMr2_2;
	wire w_dff_A_cKVQ8j5j7_2;
	wire w_dff_A_1Sr3NbGH3_2;
	wire w_dff_A_kiWkekqw1_2;
	wire w_dff_A_CUbpgPGn2_0;
	wire w_dff_A_s3zAHzsd5_0;
	wire w_dff_A_eB2W1GEJ3_0;
	wire w_dff_A_c2a3JZsZ6_0;
	wire w_dff_A_6EYbj9qD5_0;
	wire w_dff_A_URmQRko84_0;
	wire w_dff_A_jwCTRDKo0_1;
	wire w_dff_A_KHqIG8Ny1_1;
	wire w_dff_A_l7HuiG969_1;
	wire w_dff_A_1Tv02Wh29_1;
	wire w_dff_A_HJjv8p6k1_1;
	wire w_dff_A_5rAKIP7Z4_1;
	wire w_dff_A_eAq0ZszF3_1;
	wire w_dff_A_Tfb3Se8u8_1;
	wire w_dff_A_NT7xUXH68_1;
	wire w_dff_A_ST8w2acz9_1;
	wire w_dff_A_Zlcc1WBo6_1;
	wire w_dff_A_R26fKNaK3_1;
	wire w_dff_A_VewlEDL70_1;
	wire w_dff_A_yyUdDatr8_2;
	wire w_dff_A_KgHjpYpx2_2;
	wire w_dff_A_WLRj8K4X0_2;
	wire w_dff_A_h308vyhu8_2;
	wire w_dff_A_j7fqDAxq3_2;
	wire w_dff_A_C8L4BNUS5_2;
	wire w_dff_A_nYV1IXK00_2;
	wire w_dff_A_sX7oZQmF4_2;
	wire w_dff_A_eyk3KoDE9_2;
	wire w_dff_B_9BWndEVS6_1;
	wire w_dff_B_JDVZwhDt8_0;
	wire w_dff_B_guRjmfLS2_0;
	wire w_dff_A_YoFWnBwt3_0;
	wire w_dff_A_d1HhWs9R1_0;
	wire w_dff_A_jYjxtVsY3_0;
	wire w_dff_A_fIGaozpt2_0;
	wire w_dff_A_sv7ef6nn8_0;
	wire w_dff_A_uvliav676_0;
	wire w_dff_A_Bm7VBKl85_0;
	wire w_dff_A_pRmQpTHG9_0;
	wire w_dff_A_v2wpW7I60_2;
	wire w_dff_A_HYAAvPMU0_2;
	wire w_dff_A_q812jhGF1_2;
	wire w_dff_A_wYIuQO3E2_2;
	wire w_dff_A_6yWhX6pT4_2;
	wire w_dff_A_8823zXGq1_2;
	wire w_dff_A_zoxLnd2T6_2;
	wire w_dff_B_FbsYManE5_3;
	wire w_dff_B_tPbzwCid2_0;
	wire w_dff_B_DkZqUcE39_0;
	wire w_dff_B_iyOm5jen4_0;
	wire w_dff_B_fJz966m29_0;
	wire w_dff_B_0xpvP6Sy8_0;
	wire w_dff_B_yzzNuLNe8_0;
	wire w_dff_B_auaD2fl65_0;
	wire w_dff_B_HS5mRapg2_0;
	wire w_dff_B_spCLzmLV8_0;
	wire w_dff_B_q5Ktwy8s3_0;
	wire w_dff_A_SqO57Zob2_1;
	wire w_dff_A_sCOXXYkL6_1;
	wire w_dff_A_JhEi1HTD5_1;
	wire w_dff_A_ENmqCqTt3_1;
	wire w_dff_A_6TrxxOM32_1;
	wire w_dff_A_i58d2qx50_1;
	wire w_dff_A_WBLbT3Mu9_0;
	wire w_dff_A_3b3TYrUP1_0;
	wire w_dff_A_jiIgGLHY5_0;
	wire w_dff_A_CjbDfE3e9_0;
	wire w_dff_A_cODPshmq1_0;
	wire w_dff_A_JDBYFYWt7_0;
	wire w_dff_A_e6nOEHk31_0;
	wire w_dff_A_HOXSNJxj9_0;
	wire w_dff_A_oeP4XS5h4_0;
	wire w_dff_A_H1gPzLXb4_0;
	wire w_dff_A_HlfwhfIe3_0;
	wire w_dff_B_WkQ1Z08U2_3;
	wire w_dff_B_yj19BfzW4_3;
	wire w_dff_B_jcyjnR323_3;
	wire w_dff_B_9P6gXs5P0_3;
	wire w_dff_B_Jlkm723F3_3;
	wire w_dff_B_vFDnUJ2v2_3;
	wire w_dff_B_aw3uN2ng6_3;
	wire w_dff_B_MkHlyEnr7_3;
	wire w_dff_B_QR0EmBkX8_3;
	wire w_dff_B_s45QQpiD1_0;
	wire w_dff_B_Uv6o4uxD1_0;
	wire w_dff_B_ZJXg71DB7_0;
	wire w_dff_B_nqHDBrNL8_0;
	wire w_dff_B_QzdtIJtd4_0;
	wire w_dff_A_VIBDWbqU0_1;
	wire w_dff_B_jGyfQp2c6_2;
	wire w_dff_B_aJ6kLBXZ2_2;
	wire w_dff_B_ZvYqvzJP6_2;
	wire w_dff_B_rozhVQNP3_2;
	wire w_dff_A_3dL30TBv8_0;
	wire w_dff_B_XXbV3zQw3_1;
	wire w_dff_B_hMdlKyK58_1;
	wire w_dff_A_cSLTPijy3_0;
	wire w_dff_A_srPCK7nJ5_0;
	wire w_dff_B_Yh1MOgGx9_2;
	wire w_dff_A_O39kA17A9_0;
	wire w_dff_A_H2GZtF6F1_0;
	wire w_dff_A_FcRWR8m76_1;
	wire w_dff_A_7Xsqoc8r5_0;
	wire w_dff_A_vFzjVfJl1_0;
	wire w_dff_A_CJ6pJ0Sd6_0;
	wire w_dff_A_883qTqWJ8_0;
	wire w_dff_A_RYpoHz774_2;
	wire w_dff_A_SWS8zYQ67_2;
	wire w_dff_A_BJqiOklz3_2;
	wire w_dff_A_uzkzW8UG4_2;
	wire w_dff_A_QNvHU31e7_1;
	wire w_dff_A_Q8n0dWw79_1;
	wire w_dff_A_7H4wQV9e9_1;
	wire w_dff_A_T9ZOG8LW8_1;
	wire w_dff_A_AsnBQUSc1_1;
	wire w_dff_A_Kq8CvxTw7_1;
	wire w_dff_A_tmgnPL9s8_1;
	wire w_dff_A_WZEDCsWq4_1;
	wire w_dff_A_bYVKdZ3g4_2;
	wire w_dff_A_vg7FDJnQ3_2;
	wire w_dff_A_QRFb94mw6_2;
	wire w_dff_A_udxixTEL4_1;
	wire w_dff_A_qjh96vI27_0;
	wire w_dff_A_fzqXj6HD0_0;
	wire w_dff_A_gsqSXBtL6_2;
	wire w_dff_A_inIXd7Eh8_0;
	wire w_dff_A_ChJmihjf4_0;
	wire w_dff_A_eFGwfiAL1_0;
	wire w_dff_A_WzQeFSph6_0;
	wire w_dff_A_6lqp49I31_0;
	wire w_dff_A_d0pgtZvo9_0;
	wire w_dff_A_6a7MvcJ44_0;
	wire w_dff_A_47CLtQ8n0_0;
	wire w_dff_A_pLKY32TV0_0;
	wire w_dff_A_9QSAiuJY3_1;
	wire w_dff_A_hAcwclaT7_1;
	wire w_dff_A_tABhtonR0_1;
	wire w_dff_B_bGky21ci8_2;
	wire w_dff_B_ZRqV7zKa0_2;
	wire w_dff_B_hXi4GvvB5_2;
	wire w_dff_B_kzHPPf338_2;
	wire w_dff_A_ur5K87AI0_0;
	wire w_dff_A_oFPbvM8S9_0;
	wire w_dff_A_6s5JWaOQ9_0;
	wire w_dff_A_FQ3gAwJT5_0;
	wire w_dff_A_1lCmjEwm4_0;
	wire w_dff_A_KpHEoisX1_0;
	wire w_dff_A_2PZPIQRa0_0;
	wire w_dff_A_H81VmuLa9_0;
	wire w_dff_A_JCmb31hf1_0;
	wire w_dff_A_4fkzmxwA3_2;
	wire w_dff_A_0cSXR2PC0_2;
	wire w_dff_A_UmHC5iqM7_2;
	wire w_dff_A_epP6TRl44_2;
	wire w_dff_A_yZveYZra3_2;
	wire w_dff_A_KkiWDRZQ4_2;
	wire w_dff_A_xjav24r93_2;
	wire w_dff_A_xjJ1q6HZ2_2;
	wire w_dff_A_5Xt0KupC1_2;
	wire w_dff_A_BANckRck8_0;
	wire w_dff_A_kXUfKTBt6_0;
	wire w_dff_A_hZhmGr6N0_0;
	wire w_dff_A_yKn7Acjc5_0;
	wire w_dff_A_QnxKz3Rl1_0;
	wire w_dff_A_nABzgguu0_0;
	wire w_dff_B_neQ6GObu2_0;
	wire w_dff_A_qGEjEI2b9_1;
	wire w_dff_A_bQ1HpIsw9_1;
	wire w_dff_A_QqoOc1Jz9_1;
	wire w_dff_A_1bJBU0Ea0_1;
	wire w_dff_A_CJN7BoNr6_1;
	wire w_dff_A_fOOkhVnI6_1;
	wire w_dff_A_dADlnIYC6_1;
	wire w_dff_A_fVb50uyJ6_1;
	wire w_dff_A_FaerhiMT4_2;
	wire w_dff_A_T7TLZoUt2_1;
	wire w_dff_A_qO7i5XFD5_1;
	wire w_dff_A_y1OnYwrt7_1;
	wire w_dff_A_Xok89pFc6_1;
	wire w_dff_A_Lst0McxJ1_1;
	wire w_dff_A_QxIfccYM2_1;
	wire w_dff_A_egK1zrPp8_0;
	wire w_dff_A_rW7uXXy70_1;
	wire w_dff_A_5WA9MwRB4_1;
	wire w_dff_B_244tRTRv6_3;
	wire w_dff_B_lEMQTvZA9_3;
	wire w_dff_A_OrDC34Ke6_1;
	wire w_dff_A_sh3SKIBB9_1;
	wire w_dff_A_K3NLT9Ak4_1;
	wire w_dff_A_k3sAJFMy3_1;
	wire w_dff_A_V3aHJn8o0_1;
	wire w_dff_A_2f98JMSZ7_1;
	wire w_dff_A_foFC6nAh4_1;
	wire w_dff_A_6PmdFaOp5_1;
	wire w_dff_A_aWmdXhqw4_1;
	wire w_dff_A_vx1IlplW0_2;
	wire w_dff_A_UCXNWv1U7_2;
	wire w_dff_A_0qBQ3hYR1_2;
	wire w_dff_A_2crjAIGA0_2;
	wire w_dff_A_IqrXtOF58_2;
	wire w_dff_A_IMua5r6F0_2;
	wire w_dff_A_M6cJgRvz3_2;
	wire w_dff_A_bnf6zr3H2_2;
	wire w_dff_A_cyJN6K3q5_2;
	wire w_dff_A_MchCa0XT1_2;
	wire w_dff_A_YEa8x4XB1_2;
	wire w_dff_A_wF8Cl85X4_2;
	wire w_dff_A_ClLJEkci1_0;
	wire w_dff_A_f6kzESnr4_0;
	wire w_dff_A_tKHLe5Cw2_0;
	wire w_dff_A_JWwv185I6_0;
	wire w_dff_A_FC34CPBS3_0;
	wire w_dff_A_QqRuJ6Mz7_0;
	wire w_dff_A_hPp50bWJ9_0;
	wire w_dff_A_ClnPAPNM7_0;
	wire w_dff_A_mFisWiIl3_0;
	wire w_dff_A_LQZ9fwxO8_0;
	wire w_dff_A_sZJoyY4C3_0;
	wire w_dff_A_IK1gHZ8x6_0;
	wire w_dff_A_joFkzNBo9_0;
	wire w_dff_A_EME01GPk3_0;
	wire w_dff_A_2KG3pNHw2_0;
	wire w_dff_A_evZ0erhW1_0;
	wire w_dff_A_6lm5GJZU3_0;
	wire w_dff_A_4RpFJ8NO5_0;
	wire w_dff_A_Db8WX77x7_0;
	wire w_dff_A_oUv0FQ8Q0_0;
	wire w_dff_A_1vk4U44o1_0;
	wire w_dff_A_TlymtKvy7_0;
	wire w_dff_A_bZ5MyR6O9_0;
	wire w_dff_A_6rixA4pP6_0;
	wire w_dff_A_HsDIHK2K7_0;
	wire w_dff_A_URn4EI0h7_2;
	wire w_dff_A_XU4X6X4G4_0;
	wire w_dff_A_eN3cOpU68_0;
	wire w_dff_A_Phqa3cVI6_0;
	wire w_dff_A_WMxX7sO32_0;
	wire w_dff_A_VsfHtiiX0_0;
	wire w_dff_A_YygaCAQN5_0;
	wire w_dff_A_6gY5i48W2_0;
	wire w_dff_A_Gfwt14mj8_0;
	wire w_dff_A_k34j0FCu9_0;
	wire w_dff_A_v20MPbiG9_0;
	wire w_dff_A_gjGv3n1a4_0;
	wire w_dff_A_g5vGD8Aq1_0;
	wire w_dff_A_4ZouqCnj2_0;
	wire w_dff_A_1DA1D5Mc6_0;
	wire w_dff_A_drPR7nGB2_0;
	wire w_dff_A_UKTifiP88_0;
	wire w_dff_A_gycEUIEt7_0;
	wire w_dff_A_qbSLaw9U7_0;
	wire w_dff_A_sRsqK2Np6_0;
	wire w_dff_A_2h9Grpbb5_0;
	wire w_dff_A_kjPyLyTg1_0;
	wire w_dff_A_hqqkMEyB7_0;
	wire w_dff_A_j95b8i4I1_0;
	wire w_dff_A_MpPJ47RF0_0;
	wire w_dff_A_CkOdEVXw9_0;
	wire w_dff_A_DCUnLUjN5_2;
	wire w_dff_A_LK3B1J3Q0_0;
	wire w_dff_A_4UCHGtCy9_0;
	wire w_dff_A_L5lWpIQT0_0;
	wire w_dff_A_YpNPzlTs9_0;
	wire w_dff_A_vvj60zCk8_0;
	wire w_dff_A_J9zBqNvc1_0;
	wire w_dff_A_VuZSqEM76_0;
	wire w_dff_A_ySaquppi4_0;
	wire w_dff_A_QOoTBZhk3_0;
	wire w_dff_A_4pUseqsY3_0;
	wire w_dff_A_vuKy39YH7_0;
	wire w_dff_A_O6bLVEVt0_0;
	wire w_dff_A_ORTJY1pH6_0;
	wire w_dff_A_lQDhlEbv0_0;
	wire w_dff_A_Pyv83LjJ3_0;
	wire w_dff_A_sQ48iNgC9_0;
	wire w_dff_A_6XZ86Acu6_0;
	wire w_dff_A_35EwFhGE1_0;
	wire w_dff_A_6Yz27eOL3_0;
	wire w_dff_A_T5XnaazA0_0;
	wire w_dff_A_EPCzY0nk0_0;
	wire w_dff_A_ySH44Wtm2_0;
	wire w_dff_A_HVtHdww27_0;
	wire w_dff_A_XoQZlwbF4_0;
	wire w_dff_A_f97qhAPz3_0;
	wire w_dff_A_8pBCiBMs8_2;
	wire w_dff_A_clRKRtNn5_0;
	wire w_dff_A_F1xYbvEk6_0;
	wire w_dff_A_mwbhn23q5_0;
	wire w_dff_A_F4CG209h0_0;
	wire w_dff_A_6SrCwavk3_0;
	wire w_dff_A_erjEthf31_0;
	wire w_dff_A_a68gOB9j7_0;
	wire w_dff_A_WB4HwnZq6_0;
	wire w_dff_A_Zxswmoi59_0;
	wire w_dff_A_rHv7T4Nd0_0;
	wire w_dff_A_2ZAVattz3_0;
	wire w_dff_A_p3eZOdir1_0;
	wire w_dff_A_o6NAy5RB9_0;
	wire w_dff_A_hBWVZAPV9_0;
	wire w_dff_A_K71kYyS69_0;
	wire w_dff_A_ssp9WvJv0_0;
	wire w_dff_A_ZwAROs2J7_0;
	wire w_dff_A_Ebv1GTbQ8_0;
	wire w_dff_A_S0BYbNXc0_0;
	wire w_dff_A_tgchaNDi7_0;
	wire w_dff_A_1V4BEQ3z7_0;
	wire w_dff_A_8u12CGUO6_0;
	wire w_dff_A_KD0GetWJ0_0;
	wire w_dff_A_LhUQn7548_0;
	wire w_dff_A_04EcVYd20_0;
	wire w_dff_A_te6HLR6I3_0;
	wire w_dff_A_h8jo52As9_2;
	wire w_dff_A_R75aPu7G3_0;
	wire w_dff_A_EwHYCa2j3_0;
	wire w_dff_A_3hOOZs231_0;
	wire w_dff_A_UNaLyMaH6_0;
	wire w_dff_A_tNThjERl2_0;
	wire w_dff_A_uHLHGbMT5_0;
	wire w_dff_A_HTYfIR785_0;
	wire w_dff_A_M9YJ3cWh0_0;
	wire w_dff_A_8SPFwIRK5_0;
	wire w_dff_A_XoWZiUEt3_0;
	wire w_dff_A_2uGbiMSz7_0;
	wire w_dff_A_XJMQcD9b0_0;
	wire w_dff_A_tCtRc8VJ8_0;
	wire w_dff_A_UNHayenH9_0;
	wire w_dff_A_YRDJ7zfO1_0;
	wire w_dff_A_RE4s87sI8_0;
	wire w_dff_A_H1e0lKX53_0;
	wire w_dff_A_9sVH2EWT8_0;
	wire w_dff_A_UJ29qjt87_0;
	wire w_dff_A_j6E1AQjs1_0;
	wire w_dff_A_ywOoEXd11_0;
	wire w_dff_A_rEkvsX6m7_0;
	wire w_dff_A_xTDZk3NR1_0;
	wire w_dff_A_gyR8xsKb6_0;
	wire w_dff_A_laVyLnLT1_2;
	wire w_dff_A_DIISTH446_0;
	wire w_dff_A_z5pexYFN7_0;
	wire w_dff_A_C7NokHXA2_0;
	wire w_dff_A_cDGkuiuT6_0;
	wire w_dff_A_lopyjr0n8_0;
	wire w_dff_A_dHbgcKoN5_0;
	wire w_dff_A_YrhhiGQw7_0;
	wire w_dff_A_RtdbOFHE2_0;
	wire w_dff_A_C6d8BV7I8_0;
	wire w_dff_A_qopnCWSg8_0;
	wire w_dff_A_C3l1wK7Q2_0;
	wire w_dff_A_NPaJ6teP8_0;
	wire w_dff_A_lMVnUSQa9_0;
	wire w_dff_A_VwATLboz1_0;
	wire w_dff_A_Ov7GXoYI1_0;
	wire w_dff_A_w1fPEtm99_0;
	wire w_dff_A_mMXNLHmQ0_0;
	wire w_dff_A_WHGfAUfB5_0;
	wire w_dff_A_bePrq1Ae9_0;
	wire w_dff_A_gJZmO8AF9_0;
	wire w_dff_A_fFKp0A8X8_0;
	wire w_dff_A_nBLlvPvN3_0;
	wire w_dff_A_deOSyrnr7_2;
	wire w_dff_A_a4fwSDdu0_0;
	wire w_dff_A_Bjl15bpH7_0;
	wire w_dff_A_b8SdHcNp8_0;
	wire w_dff_A_Ovob1aRK7_0;
	wire w_dff_A_SQXgrj802_0;
	wire w_dff_A_gfpiyVsr9_0;
	wire w_dff_A_q9RiCr198_0;
	wire w_dff_A_6cGXUVLp6_0;
	wire w_dff_A_NBR5S5FV9_0;
	wire w_dff_A_tgussN988_0;
	wire w_dff_A_kLK4FU254_0;
	wire w_dff_A_S0tChvUW8_0;
	wire w_dff_A_vNXHHIjf9_0;
	wire w_dff_A_H937d63b3_0;
	wire w_dff_A_EUn111oZ0_0;
	wire w_dff_A_ioefZaX57_0;
	wire w_dff_A_9H0l3MS87_0;
	wire w_dff_A_xBDueBwD2_0;
	wire w_dff_A_CuuDcqMy7_0;
	wire w_dff_A_b0mAXX6M5_0;
	wire w_dff_A_akTJ28XZ2_0;
	wire w_dff_A_fVpoRMzG0_0;
	wire w_dff_A_QEwcGjuL7_0;
	wire w_dff_A_K9G3agmX4_0;
	wire w_dff_A_lrqAObpH1_2;
	wire w_dff_A_GcKxzyGJ6_0;
	wire w_dff_A_GmhPtNCE3_0;
	wire w_dff_A_nwps0OYt5_0;
	wire w_dff_A_PiJuzgoU7_0;
	wire w_dff_A_nLm44Rnf1_0;
	wire w_dff_A_IZBxedDW6_0;
	wire w_dff_A_yXKPRIBm4_0;
	wire w_dff_A_UanwxyNM5_0;
	wire w_dff_A_hnWstzmq3_0;
	wire w_dff_A_rEqdIL1A6_0;
	wire w_dff_A_aDdIWWAw5_0;
	wire w_dff_A_nC26oicF6_0;
	wire w_dff_A_6uET4wis0_0;
	wire w_dff_A_AEDBBR8K6_0;
	wire w_dff_A_5eQrw2qB3_0;
	wire w_dff_A_i8KaPZQ84_0;
	wire w_dff_A_9BbMzB5n3_0;
	wire w_dff_A_nTfYHYpn1_0;
	wire w_dff_A_glGd2eIY0_0;
	wire w_dff_A_kFXj5wby9_0;
	wire w_dff_A_FR4YFsJa2_0;
	wire w_dff_A_bZpnLv9f9_0;
	wire w_dff_A_o90m62D30_0;
	wire w_dff_A_vUia2Ft49_0;
	wire w_dff_A_wFW2ch691_2;
	wire w_dff_A_nUq230zl4_0;
	wire w_dff_A_qSwWXXuX5_0;
	wire w_dff_A_JYnFWZ4p0_0;
	wire w_dff_A_6Tbd5IY18_0;
	wire w_dff_A_dFpr3Elq1_0;
	wire w_dff_A_RyCOhIiE7_0;
	wire w_dff_A_oimxdRd20_0;
	wire w_dff_A_eBcUOe005_0;
	wire w_dff_A_x3WlSW253_0;
	wire w_dff_A_heONL2uT7_0;
	wire w_dff_A_EV4S88b56_0;
	wire w_dff_A_rgZALcik5_0;
	wire w_dff_A_4eWjyWWv5_0;
	wire w_dff_A_VNptx7qK4_0;
	wire w_dff_A_iUn7dDuR6_0;
	wire w_dff_A_Ut4nLxxv1_0;
	wire w_dff_A_BJQ5DKvF3_0;
	wire w_dff_A_lTPtvgTj5_0;
	wire w_dff_A_l0yD8ZRM2_0;
	wire w_dff_A_y02V02D96_0;
	wire w_dff_A_ycCJAbyC0_0;
	wire w_dff_A_8ejQo4jA0_0;
	wire w_dff_A_ljXSKrKm8_0;
	wire w_dff_A_yAVcfKPP6_0;
	wire w_dff_A_EI1AbcoC2_2;
	wire w_dff_A_8JD0Pdk98_0;
	wire w_dff_A_osCCU1Yc0_0;
	wire w_dff_A_QiF03HjA7_0;
	wire w_dff_A_Cl8U4e6d0_0;
	wire w_dff_A_X0ZFpbfj8_0;
	wire w_dff_A_QCHUAAkh1_0;
	wire w_dff_A_tNR47FzG2_0;
	wire w_dff_A_SEEB3kFx5_0;
	wire w_dff_A_Wj5wxuFc3_0;
	wire w_dff_A_7dVf7Ssj6_0;
	wire w_dff_A_wy33EccP1_0;
	wire w_dff_A_vShCL3cO4_0;
	wire w_dff_A_oj45jCHk3_0;
	wire w_dff_A_GM5B2vaZ3_0;
	wire w_dff_A_eonXjgxS2_0;
	wire w_dff_A_MxmfaX7b7_0;
	wire w_dff_A_PGsUldvm8_0;
	wire w_dff_A_iXOBFjoF4_0;
	wire w_dff_A_Et2Sl7yz8_0;
	wire w_dff_A_gXPrIarz7_0;
	wire w_dff_A_yJanGnWa1_0;
	wire w_dff_A_JU2DrTmE6_0;
	wire w_dff_A_niZrNab53_0;
	wire w_dff_A_yjBKcbmZ0_0;
	wire w_dff_A_V3bxT7gL2_0;
	wire w_dff_A_O6jn1Gue3_2;
	wire w_dff_A_kgsD6hKS3_0;
	wire w_dff_A_5IvpyKGc3_0;
	wire w_dff_A_fu73RqIQ8_0;
	wire w_dff_A_X9OVA8s22_0;
	wire w_dff_A_EZqJvrRG6_0;
	wire w_dff_A_Rps1wixn1_0;
	wire w_dff_A_r5whXDcm0_0;
	wire w_dff_A_oGwqlfyY7_0;
	wire w_dff_A_f0kZlnSr0_0;
	wire w_dff_A_lUJL6bqw8_0;
	wire w_dff_A_lW3LOW715_0;
	wire w_dff_A_cIiEsxtk6_0;
	wire w_dff_A_5uFhLSaM2_0;
	wire w_dff_A_uqrlZ0w69_0;
	wire w_dff_A_aUBDG2uL6_0;
	wire w_dff_A_ovWTiWeL1_0;
	wire w_dff_A_uDPFbiSV5_0;
	wire w_dff_A_PFnYDDsh9_0;
	wire w_dff_A_LyxSbZFw9_0;
	wire w_dff_A_6auhD7d33_0;
	wire w_dff_A_gK4yLJSg5_0;
	wire w_dff_A_NFlCp7eI0_0;
	wire w_dff_A_bDsVM3Cz7_1;
	wire w_dff_A_BEa6ECR94_0;
	wire w_dff_A_j8BSzuoO5_0;
	wire w_dff_A_wqewGXlq4_0;
	wire w_dff_A_Xrjtlo7x2_0;
	wire w_dff_A_JygVPBNZ0_0;
	wire w_dff_A_4gQ4kPKd2_0;
	wire w_dff_A_UjBAK97Z1_0;
	wire w_dff_A_v6i9W8d93_0;
	wire w_dff_A_dReMKxeq8_0;
	wire w_dff_A_hBzNvfgR7_0;
	wire w_dff_A_9IfKUUth2_0;
	wire w_dff_A_ecr7qeEJ3_0;
	wire w_dff_A_vfAaOUuf3_0;
	wire w_dff_A_r5YP6lXY8_0;
	wire w_dff_A_83NxtOxK1_0;
	wire w_dff_A_ee9mZmBx6_0;
	wire w_dff_A_QXu8jWsX3_0;
	wire w_dff_A_AKZURNN02_0;
	wire w_dff_A_WvwA8LiT6_0;
	wire w_dff_A_Krl3ZUX24_0;
	wire w_dff_A_bPIcYI5T0_0;
	wire w_dff_A_6iYzJI2M5_0;
	wire w_dff_A_YCHX3iBi0_0;
	wire w_dff_A_Ptv9l8jB6_0;
	wire w_dff_A_JveD93U55_0;
	wire w_dff_A_d7DwcygA1_2;
	wire w_dff_A_MhstYeIf3_0;
	wire w_dff_A_Yl5exmZf3_0;
	wire w_dff_A_72IKoJsn0_0;
	wire w_dff_A_6PQ7w8RY1_0;
	wire w_dff_A_8RtDEWQX2_0;
	wire w_dff_A_LcxT1DII1_0;
	wire w_dff_A_zM3QRekq3_0;
	wire w_dff_A_Md0LfRkU8_0;
	wire w_dff_A_yII40mDR7_0;
	wire w_dff_A_3wsZMJIN8_0;
	wire w_dff_A_mdki67i10_0;
	wire w_dff_A_K6ykE9Es0_0;
	wire w_dff_A_S4xidspa6_0;
	wire w_dff_A_KSV1Dyqt8_0;
	wire w_dff_A_8dZ3D4dc2_0;
	wire w_dff_A_U2k9AOlS6_0;
	wire w_dff_A_um8nsU6v7_0;
	wire w_dff_A_VdSaoWRT1_0;
	wire w_dff_A_Q3xRzlFV7_0;
	wire w_dff_A_EJJpLg9J1_0;
	wire w_dff_A_07fLWie52_0;
	wire w_dff_A_eu2X2mip2_0;
	wire w_dff_A_VbVzM2jM1_2;
	wire w_dff_A_CgoddBim3_0;
	wire w_dff_A_Jgo03Sv45_0;
	wire w_dff_A_wFDivU5a4_0;
	wire w_dff_A_ZwYGWjRz5_0;
	wire w_dff_A_50WfZlRv9_0;
	wire w_dff_A_HtYxp3CU8_0;
	wire w_dff_A_GvkBVEZY7_0;
	wire w_dff_A_B5NMwLW42_0;
	wire w_dff_A_ZEsUSQyw7_0;
	wire w_dff_A_xuXfIYyy9_0;
	wire w_dff_A_3qJoRJzD0_0;
	wire w_dff_A_HFBl8UVZ8_0;
	wire w_dff_A_AggPnzlb1_0;
	wire w_dff_A_z9iQBznL7_0;
	wire w_dff_A_rqYgT0Dl0_0;
	wire w_dff_A_Vnn3D59h3_0;
	wire w_dff_A_fVFkq9qw8_0;
	wire w_dff_A_gvAHydQ76_0;
	wire w_dff_A_4N8IUoXA7_0;
	wire w_dff_A_AqquzEvy1_0;
	wire w_dff_A_Retbe4sH3_0;
	wire w_dff_A_4P6xKnKW5_0;
	wire w_dff_A_46oFJh5I3_2;
	wire w_dff_A_C0PghwRv6_0;
	wire w_dff_A_wgptwsmK8_0;
	wire w_dff_A_9jwx3rml7_0;
	wire w_dff_A_JdOCm0dx1_0;
	wire w_dff_A_MLGMIGu43_0;
	wire w_dff_A_8B4y4y9K3_0;
	wire w_dff_A_pkjTEZjv2_0;
	wire w_dff_A_Ml5hqJBm4_0;
	wire w_dff_A_q6NT3oCv1_0;
	wire w_dff_A_pgP4yugU0_0;
	wire w_dff_A_qd0YjtjN5_0;
	wire w_dff_A_hQgmV7lM8_0;
	wire w_dff_A_COVMCks73_0;
	wire w_dff_A_uISI1WsD5_0;
	wire w_dff_A_QikJSJ3d1_0;
	wire w_dff_A_4c9L0DV80_0;
	wire w_dff_A_0RQkebOo9_0;
	wire w_dff_A_2vQiqEB96_0;
	wire w_dff_A_YaBG4oSU9_0;
	wire w_dff_A_MdzUCVzI6_0;
	wire w_dff_A_lQ1dH66v6_0;
	wire w_dff_A_QMKe07Im0_0;
	wire w_dff_A_McwYecOY1_0;
	wire w_dff_A_D604cKvP7_0;
	wire w_dff_A_vyrLqLGJ4_0;
	wire w_dff_A_U7erAsDQ5_2;
	wire w_dff_A_TM5MgPuX3_0;
	wire w_dff_A_Mz9qLphq2_0;
	wire w_dff_A_2As3Gp9u4_0;
	wire w_dff_A_vXcrQt8P2_0;
	wire w_dff_A_yrZBHJd72_0;
	wire w_dff_A_HDSOKIyw3_0;
	wire w_dff_A_dA3HrudG7_0;
	wire w_dff_A_oSp4Wycw9_0;
	wire w_dff_A_l10DnAiv7_0;
	wire w_dff_A_zCXOxBdL0_0;
	wire w_dff_A_mgNFwFQI6_0;
	wire w_dff_A_KL22KnRp0_0;
	wire w_dff_A_M4wox5Ln1_0;
	wire w_dff_A_lKvVqxvf2_0;
	wire w_dff_A_VtjWYBoD7_0;
	wire w_dff_A_nRN3mXyO0_0;
	wire w_dff_A_f4YfKqPQ5_0;
	wire w_dff_A_lJZCFmRb2_0;
	wire w_dff_A_4cghf02G5_0;
	wire w_dff_A_zayDYMAC9_0;
	wire w_dff_A_MhpwNvY03_0;
	wire w_dff_A_pRnNxhi55_0;
	wire w_dff_A_GaIMETuo0_0;
	wire w_dff_A_kFURueqb2_2;
	wire w_dff_A_tfJCnvsX0_0;
	wire w_dff_A_4MHuud4Z4_0;
	wire w_dff_A_rFqSc2Fp3_0;
	wire w_dff_A_0sGc09mi4_0;
	wire w_dff_A_COMTXygF4_0;
	wire w_dff_A_pHqeztw50_0;
	wire w_dff_A_R7Y3MG942_0;
	wire w_dff_A_xRYGPthN0_0;
	wire w_dff_A_M4Z4rDQt2_0;
	wire w_dff_A_kFyR0jOj6_0;
	wire w_dff_A_DyDUDH0p4_0;
	wire w_dff_A_xqnlnMaR6_0;
	wire w_dff_A_rJVwUmKk0_0;
	wire w_dff_A_qRogF6Ix9_0;
	wire w_dff_A_IJZegaBq5_0;
	wire w_dff_A_uq1pQA367_0;
	wire w_dff_A_2vWaFgIl2_0;
	wire w_dff_A_1TKF6j2i2_0;
	wire w_dff_A_Kankvch38_0;
	wire w_dff_A_f6YJmiCl1_0;
	wire w_dff_A_ikFvfpAo1_0;
	wire w_dff_A_MyBrPLSD4_0;
	wire w_dff_A_154bAPmV3_0;
	wire w_dff_A_0bei3kWP7_2;
	wire w_dff_A_FW3tNPOQ3_0;
	wire w_dff_A_p3rjj3bx0_0;
	wire w_dff_A_DDv9Ri6O3_0;
	wire w_dff_A_7AnUinVD1_0;
	wire w_dff_A_BjlvJ0cv9_0;
	wire w_dff_A_RDyqs1ny6_0;
	wire w_dff_A_0sjJb1qh1_0;
	wire w_dff_A_SC86Nwwo5_0;
	wire w_dff_A_2TSW3xlc0_0;
	wire w_dff_A_Q8RntV027_0;
	wire w_dff_A_zisxz3fN4_0;
	wire w_dff_A_z2UgFbIY1_0;
	wire w_dff_A_kOlKxf7O4_2;
	wire w_dff_A_WifP3QV35_0;
	wire w_dff_A_rCvrwCWK4_0;
	wire w_dff_A_tWQhGJB15_0;
	wire w_dff_A_iJBFqXoD7_0;
	wire w_dff_A_FIPprnkS9_0;
	wire w_dff_A_o0Ti0cIn1_0;
	wire w_dff_A_bfi6CDsu0_0;
	wire w_dff_A_EaLwtXtj9_2;
	wire w_dff_A_Yw8WOXeD3_0;
	wire w_dff_A_rihFLxqu4_0;
	wire w_dff_A_Kl7a5jAB0_0;
	wire w_dff_A_pCjPIYbn1_0;
	wire w_dff_A_gWtLxFGp7_0;
	wire w_dff_A_8iMkopc76_0;
	wire w_dff_A_luZJ4B4N8_0;
	wire w_dff_A_CZ2WFe3r6_0;
	wire w_dff_A_a8gxr0EZ7_0;
	wire w_dff_A_i7fpZ1qg5_2;
	wire w_dff_A_rvjWJORW9_0;
	wire w_dff_A_T2UfIs6M5_0;
	wire w_dff_A_nAlhdSUP5_0;
	wire w_dff_A_xvs9Erk25_0;
	wire w_dff_A_UxxXG8wq0_0;
	wire w_dff_A_IulKnn1f1_0;
	wire w_dff_A_1sEohxXZ4_0;
	wire w_dff_A_OKY0dIbs7_0;
	wire w_dff_A_VdkCCeHd8_0;
	wire w_dff_A_vdT0ciDk9_0;
	wire w_dff_A_OWy0ZP7R1_0;
	wire w_dff_A_uu90gjxu6_2;
	wire w_dff_A_TgbimvxW0_0;
	wire w_dff_A_59cdx3DS7_2;
	wire w_dff_A_HlFeHme37_0;
	wire w_dff_A_Qci0cMBR4_0;
	wire w_dff_A_t0q54zPC0_0;
	wire w_dff_A_k6q6b7sE7_0;
	wire w_dff_A_j2wVWtWp7_2;
	wire w_dff_A_peHDjjEc4_0;
	wire w_dff_A_yvuvlarN9_2;
	wire w_dff_A_hKsJVxjJ0_0;
	wire w_dff_A_ToHw2GrJ1_0;
	wire w_dff_A_RrvOc9bb9_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_wF8Cl85X4_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_URn4EI0h7_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_8pBCiBMs8_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_n92_0[1]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_G17gat_2[2]),.dout(w_dff_A_h8jo52As9_2),.clk(gclk));
	jnot g009(.din(w_G17gat_2[1]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G13gat_0[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G1gat_1[0]),.dout(n97),.clk(gclk));
	jnot g012(.din(w_G26gat_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(n98),.dinb(w_n97_0[1]),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_dff_B_kiZvJ92o9_1),.dout(n100),.clk(gclk));
	jor g015(.dina(n100),.dinb(w_n95_0[2]),.dout(n101),.clk(gclk));
	jor g016(.dina(w_n101_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_laVyLnLT1_2),.clk(gclk));
	jnot g017(.din(w_G80gat_0[1]),.dout(n103),.clk(gclk));
	jand g018(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n104),.clk(gclk));
	jnot g019(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jor g020(.dina(n105),.dinb(w_n103_0[1]),.dout(w_dff_A_deOSyrnr7_2),.clk(gclk));
	jnot g021(.din(w_G36gat_0[0]),.dout(n107),.clk(gclk));
	jnot g022(.din(w_G59gat_1[0]),.dout(n108),.clk(gclk));
	jor g023(.dina(w_n108_0[1]),.dinb(n107),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n109_0[1]),.dinb(w_n103_0[0]),.dout(w_dff_A_lrqAObpH1_2),.clk(gclk));
	jnot g025(.din(w_G42gat_1[2]),.dout(n111),.clk(gclk));
	jor g026(.dina(w_n109_0[0]),.dinb(w_n111_0[1]),.dout(w_dff_A_wFW2ch691_2),.clk(gclk));
	jor g027(.dina(G88gat),.dinb(G87gat),.dout(n113),.clk(gclk));
	jand g028(.dina(w_n113_0[1]),.dinb(w_dff_B_tAReGijg0_1),.dout(w_dff_A_EI1AbcoC2_2),.clk(gclk));
	jnot g029(.din(w_G390gat_0[0]),.dout(n115),.clk(gclk));
	jor g030(.dina(w_n101_0[0]),.dinb(w_dff_B_zHSEY54C2_1),.dout(w_dff_A_O6jn1Gue3_2),.clk(gclk));
	jand g031(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g033(.dina(w_n93_0[0]),.dinb(w_G55gat_0[2]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_n119_0[2]),.dinb(w_G29gat_0[0]),.dout(n120),.clk(gclk));
	jand g035(.dina(n120),.dinb(w_G68gat_0[1]),.dout(w_dff_A_d7DwcygA1_2),.clk(gclk));
	jand g036(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n122),.clk(gclk));
	jand g037(.dina(w_n119_0[1]),.dinb(w_dff_B_kggM7kW44_1),.dout(n123),.clk(gclk));
	jand g038(.dina(n123),.dinb(w_n122_0[1]),.dout(w_dff_A_VbVzM2jM1_2),.clk(gclk));
	jand g039(.dina(w_n113_0[0]),.dinb(w_dff_B_qVLElNTY8_1),.dout(w_dff_A_46oFJh5I3_2),.clk(gclk));
	jxor g040(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n126),.clk(gclk));
	jxor g041(.dina(n126),.dinb(w_dff_B_IYnRNLZA4_1),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n128),.clk(gclk));
	jxor g043(.dina(n128),.dinb(w_G130gat_0[1]),.dout(n129),.clk(gclk));
	jxor g044(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G126gat_0[2]),.dinb(w_G121gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(n131),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n129),.dout(n133),.clk(gclk));
	jxor g048(.dina(n133),.dinb(w_dff_B_rs6GoOFe1_1),.dout(w_dff_A_U7erAsDQ5_2),.clk(gclk));
	jxor g049(.dina(w_G189gat_2[1]),.dinb(w_G183gat_1[2]),.dout(n135),.clk(gclk));
	jxor g050(.dina(n135),.dinb(w_dff_B_xZ4cSpAA9_1),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_G159gat_1[2]),.dinb(w_G130gat_0[0]),.dout(n137),.clk(gclk));
	jxor g052(.dina(n137),.dinb(w_G165gat_1[2]),.dout(n138),.clk(gclk));
	jxor g053(.dina(w_G177gat_1[2]),.dinb(w_G171gat_1[2]),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G201gat_1[1]),.dinb(w_G195gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g057(.dina(n142),.dinb(w_dff_B_CaTEttEE8_1),.dout(w_dff_A_kFURueqb2_2),.clk(gclk));
	jnot g058(.din(w_G268gat_0[1]),.dout(n144),.clk(gclk));
	jand g059(.dina(w_G447gat_1),.dinb(w_G80gat_0[0]),.dout(n145),.clk(gclk));
	jand g060(.dina(n145),.dinb(w_n86_0[0]),.dout(n146),.clk(gclk));
	jand g061(.dina(w_n146_0[1]),.dinb(w_G55gat_0[1]),.dout(n147),.clk(gclk));
	jand g062(.dina(n147),.dinb(w_n144_0[1]),.dout(n148),.clk(gclk));
	jand g063(.dina(w_n111_0[0]),.dinb(w_n95_0[1]),.dout(n149),.clk(gclk));
	jnot g064(.din(w_n149_0[1]),.dout(n150),.clk(gclk));
	jand g065(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(w_G42gat_1[1]),.dinb(w_G17gat_2[0]),.dout(n152),.clk(gclk));
	jnot g067(.din(w_n152_0[1]),.dout(n153),.clk(gclk));
	jand g068(.dina(n153),.dinb(w_n151_0[1]),.dout(n154),.clk(gclk));
	jand g069(.dina(n154),.dinb(w_G447gat_0[2]),.dout(n155),.clk(gclk));
	jand g070(.dina(n155),.dinb(w_dff_B_hMdlKyK58_1),.dout(n156),.clk(gclk));
	jnot g071(.din(w_n92_0[0]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n104_0[0]),.dinb(w_G42gat_1[0]),.dout(n158),.clk(gclk));
	jand g073(.dina(w_G51gat_1[0]),.dinb(w_G17gat_1[2]),.dout(n159),.clk(gclk));
	jnot g074(.din(n159),.dout(n160),.clk(gclk));
	jor g075(.dina(n160),.dinb(n158),.dout(n161),.clk(gclk));
	jor g076(.dina(n161),.dinb(w_dff_B_XXbV3zQw3_1),.dout(n162),.clk(gclk));
	jnot g077(.din(w_n162_0[1]),.dout(n163),.clk(gclk));
	jor g078(.dina(n163),.dinb(n156),.dout(n164),.clk(gclk));
	jand g079(.dina(w_n164_3[1]),.dinb(w_G126gat_0[1]),.dout(n165),.clk(gclk));
	jnot g080(.din(w_G156gat_0[0]),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n108_0[0]),.dout(n167),.clk(gclk));
	jand g082(.dina(w_n167_0[1]),.dinb(w_G447gat_0[1]),.dout(n168),.clk(gclk));
	jand g083(.dina(w_n168_0[1]),.dinb(w_G17gat_1[1]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n97_0[0]),.dout(n170),.clk(gclk));
	jand g085(.dina(w_n170_1[1]),.dinb(w_G153gat_0[2]),.dout(n171),.clk(gclk));
	jor g086(.dina(w_dff_B_rl9Vq7JE8_0),.dinb(n165),.dout(n172),.clk(gclk));
	jor g087(.dina(n172),.dinb(w_n148_1[2]),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n173_0[1]),.dinb(w_G246gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_n122_0[0]),.dinb(w_G42gat_0[2]),.dout(n175),.clk(gclk));
	jand g090(.dina(G73gat),.dinb(G72gat),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_neQ6GObu2_0),.dinb(n175),.dout(n177),.clk(gclk));
	jand g092(.dina(n177),.dinb(w_n119_0[0]),.dout(n178),.clk(gclk));
	jand g093(.dina(w_n178_3[1]),.dinb(w_G201gat_1[0]),.dout(n179),.clk(gclk));
	jor g094(.dina(w_dff_B_glchsX2h6_0),.dinb(n174),.dout(n180),.clk(gclk));
	jnot g095(.din(w_G201gat_0[2]),.dout(n181),.clk(gclk));
	jnot g096(.din(w_n148_1[1]),.dout(n182),.clk(gclk));
	jnot g097(.din(w_G126gat_0[0]),.dout(n183),.clk(gclk));
	jnot g098(.din(w_G51gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(w_n99_0[0]),.dinb(w_dff_B_BJriCuaR1_1),.dout(n185),.clk(gclk));
	jor g100(.dina(w_n152_0[0]),.dinb(w_n167_0[0]),.dout(n186),.clk(gclk));
	jor g101(.dina(n186),.dinb(w_n185_0[1]),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(w_n149_0[0]),.dout(n188),.clk(gclk));
	jand g103(.dina(w_n162_0[0]),.dinb(n188),.dout(n189),.clk(gclk));
	jor g104(.dina(n189),.dinb(w_dff_B_jn0YtmUD9_1),.dout(n190),.clk(gclk));
	jnot g105(.din(w_G153gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(w_n151_0[0]),.dinb(w_n185_0[0]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_n95_0[0]),.dout(n193),.clk(gclk));
	jand g108(.dina(n193),.dinb(w_G1gat_0[1]),.dout(n194),.clk(gclk));
	jor g109(.dina(n194),.dinb(w_dff_B_kvx6MqsJ7_1),.dout(n195),.clk(gclk));
	jand g110(.dina(n195),.dinb(n190),.dout(n196),.clk(gclk));
	jand g111(.dina(n196),.dinb(w_dff_B_f9PFycb75_1),.dout(n197),.clk(gclk));
	jxor g112(.dina(w_n197_0[2]),.dinb(w_n181_0[2]),.dout(n198),.clk(gclk));
	jand g113(.dina(w_n198_0[2]),.dinb(w_G228gat_3[1]),.dout(n199),.clk(gclk));
	jand g114(.dina(w_n173_0[0]),.dinb(w_G201gat_0[1]),.dout(n200),.clk(gclk));
	jand g115(.dina(w_n200_0[1]),.dinb(w_G237gat_3[1]),.dout(n201),.clk(gclk));
	jand g116(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n202),.clk(gclk));
	jand g117(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n203),.clk(gclk));
	jor g118(.dina(n203),.dinb(n202),.dout(n204),.clk(gclk));
	jor g119(.dina(w_dff_B_qzjTKzz27_0),.dinb(n201),.dout(n205),.clk(gclk));
	jor g120(.dina(n205),.dinb(w_dff_B_EPAe0jse5_1),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_ZpbdFtNi8_1),.dout(n207),.clk(gclk));
	jor g122(.dina(w_n198_0[1]),.dinb(w_G261gat_0[2]),.dout(n208),.clk(gclk));
	jnot g123(.din(w_G261gat_0[1]),.dout(n209),.clk(gclk));
	jnot g124(.din(w_n198_0[0]),.dout(n210),.clk(gclk));
	jor g125(.dina(n210),.dinb(w_n209_0[1]),.dout(n211),.clk(gclk));
	jand g126(.dina(n211),.dinb(w_G219gat_3[2]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_KBWPjDHB7_1),.dout(n213),.clk(gclk));
	jor g128(.dina(n213),.dinb(n207),.dout(w_dff_A_0bei3kWP7_2),.clk(gclk));
	jand g129(.dina(w_n164_3[0]),.dinb(w_G111gat_0[1]),.dout(n215),.clk(gclk));
	jand g130(.dina(w_n170_1[0]),.dinb(w_G143gat_0[1]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_n148_1[0]),.dout(n217),.clk(gclk));
	jor g132(.dina(n217),.dinb(n215),.dout(n218),.clk(gclk));
	jxor g133(.dina(w_n218_1[1]),.dinb(w_G183gat_1[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n219_0[2]),.dinb(w_G228gat_3[0]),.dout(n220),.clk(gclk));
	jand g135(.dina(w_n178_3[0]),.dinb(w_G183gat_1[0]),.dout(n221),.clk(gclk));
	jand g136(.dina(w_n218_1[0]),.dinb(w_G183gat_0[2]),.dout(n222),.clk(gclk));
	jand g137(.dina(w_n222_0[2]),.dinb(w_G237gat_3[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n218_0[2]),.dinb(w_G246gat_3[0]),.dout(n224),.clk(gclk));
	jand g139(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_7PLyaIN99_0),.dinb(n224),.dout(n226),.clk(gclk));
	jor g141(.dina(n226),.dinb(n223),.dout(n227),.clk(gclk));
	jor g142(.dina(n227),.dinb(w_dff_B_84n8DlGf3_1),.dout(n228),.clk(gclk));
	jor g143(.dina(n228),.dinb(w_dff_B_7gnwILmQ9_1),.dout(n229),.clk(gclk));
	jand g144(.dina(w_n164_2[2]),.dinb(w_G116gat_0[1]),.dout(n230),.clk(gclk));
	jand g145(.dina(w_n170_0[2]),.dinb(w_G146gat_0[1]),.dout(n231),.clk(gclk));
	jor g146(.dina(n231),.dinb(w_n148_0[2]),.dout(n232),.clk(gclk));
	jor g147(.dina(n232),.dinb(n230),.dout(n233),.clk(gclk));
	jand g148(.dina(w_n233_1[1]),.dinb(w_G189gat_2[0]),.dout(n234),.clk(gclk));
	jor g149(.dina(w_n233_1[0]),.dinb(w_G189gat_1[2]),.dout(n235),.clk(gclk));
	jand g150(.dina(w_n164_2[1]),.dinb(w_G121gat_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n170_0[1]),.dinb(w_G149gat_0[1]),.dout(n237),.clk(gclk));
	jor g152(.dina(n237),.dinb(w_n148_0[1]),.dout(n238),.clk(gclk));
	jor g153(.dina(n238),.dinb(n236),.dout(n239),.clk(gclk));
	jand g154(.dina(w_n239_1[1]),.dinb(w_G195gat_2[0]),.dout(n240),.clk(gclk));
	jor g155(.dina(w_n239_1[0]),.dinb(w_G195gat_1[2]),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n197_0[1]),.dinb(w_n181_0[1]),.dout(n242),.clk(gclk));
	jnot g157(.din(w_n242_0[1]),.dout(n243),.clk(gclk));
	jor g158(.dina(w_n200_0[0]),.dinb(w_G261gat_0[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(n244),.dinb(n243),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n245_0[1]),.dinb(w_n241_0[1]),.dout(n246),.clk(gclk));
	jor g161(.dina(n246),.dinb(w_n240_0[1]),.dout(n247),.clk(gclk));
	jand g162(.dina(w_n247_0[1]),.dinb(w_n235_0[1]),.dout(n248),.clk(gclk));
	jor g163(.dina(n248),.dinb(w_n234_0[1]),.dout(n249),.clk(gclk));
	jor g164(.dina(w_n249_0[1]),.dinb(w_n219_0[1]),.dout(n250),.clk(gclk));
	jnot g165(.din(w_n219_0[0]),.dout(n251),.clk(gclk));
	jnot g166(.din(w_n234_0[0]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n235_0[0]),.dout(n253),.clk(gclk));
	jnot g168(.din(w_n240_0[0]),.dout(n254),.clk(gclk));
	jnot g169(.din(w_n241_0[0]),.dout(n255),.clk(gclk));
	jor g170(.dina(w_n197_0[0]),.dinb(w_n181_0[0]),.dout(n256),.clk(gclk));
	jand g171(.dina(n256),.dinb(w_n209_0[0]),.dout(n257),.clk(gclk));
	jor g172(.dina(n257),.dinb(w_n242_0[0]),.dout(n258),.clk(gclk));
	jor g173(.dina(w_n258_0[1]),.dinb(w_dff_B_E40CS4Av2_1),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(w_dff_B_E84IDsFC6_1),.dout(n260),.clk(gclk));
	jor g175(.dina(w_n260_0[1]),.dinb(w_dff_B_a0X6tw2p1_1),.dout(n261),.clk(gclk));
	jand g176(.dina(n261),.dinb(w_dff_B_XRitnMuY1_1),.dout(n262),.clk(gclk));
	jor g177(.dina(w_n262_0[1]),.dinb(w_dff_B_7UJ5sV2m1_1),.dout(n263),.clk(gclk));
	jand g178(.dina(n263),.dinb(w_G219gat_3[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(n264),.dinb(w_dff_B_fDhPSzWG5_1),.dout(n265),.clk(gclk));
	jor g180(.dina(n265),.dinb(w_dff_B_4rqCsIZw9_1),.dout(w_dff_A_kOlKxf7O4_2),.clk(gclk));
	jxor g181(.dina(w_n233_0[2]),.dinb(w_G189gat_1[1]),.dout(n267),.clk(gclk));
	jand g182(.dina(w_n267_0[2]),.dinb(w_G228gat_2[2]),.dout(n268),.clk(gclk));
	jand g183(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n269),.clk(gclk));
	jand g184(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(w_G246gat_2[2]),.dout(n271),.clk(gclk));
	jand g186(.dina(w_dff_B_XpaDHBzu2_0),.dinb(w_n233_0[1]),.dout(n272),.clk(gclk));
	jor g187(.dina(n272),.dinb(w_dff_B_eALMfTKs8_1),.dout(n273),.clk(gclk));
	jand g188(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n274),.clk(gclk));
	jand g189(.dina(w_n178_2[2]),.dinb(w_G189gat_0[2]),.dout(n275),.clk(gclk));
	jor g190(.dina(n275),.dinb(w_dff_B_3ZMkq8Hj4_1),.dout(n276),.clk(gclk));
	jor g191(.dina(w_dff_B_6E7KgVIu3_0),.dinb(n273),.dout(n277),.clk(gclk));
	jor g192(.dina(n277),.dinb(w_dff_B_s73pqaah1_1),.dout(n278),.clk(gclk));
	jor g193(.dina(w_n267_0[1]),.dinb(w_n247_0[0]),.dout(n279),.clk(gclk));
	jnot g194(.din(w_n267_0[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(w_dff_B_JIUTpmJ50_0),.dinb(w_n260_0[0]),.dout(n281),.clk(gclk));
	jand g196(.dina(n281),.dinb(w_G219gat_3[0]),.dout(n282),.clk(gclk));
	jand g197(.dina(n282),.dinb(w_dff_B_FU6iXRqU8_1),.dout(n283),.clk(gclk));
	jor g198(.dina(n283),.dinb(w_dff_B_lTkxRn4p5_1),.dout(w_dff_A_EaLwtXtj9_2),.clk(gclk));
	jxor g199(.dina(w_n239_0[2]),.dinb(w_G195gat_1[1]),.dout(n285),.clk(gclk));
	jand g200(.dina(w_n285_0[2]),.dinb(w_G228gat_2[1]),.dout(n286),.clk(gclk));
	jand g201(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n287),.clk(gclk));
	jand g202(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(w_G246gat_2[1]),.dout(n289),.clk(gclk));
	jand g204(.dina(w_dff_B_Cy6GudwD7_0),.dinb(w_n239_0[1]),.dout(n290),.clk(gclk));
	jor g205(.dina(n290),.dinb(w_dff_B_Cx9viwQK4_1),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n178_2[1]),.dinb(w_G195gat_0[2]),.dout(n292),.clk(gclk));
	jand g207(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n293),.clk(gclk));
	jor g208(.dina(w_dff_B_pg4cL8EJ9_0),.dinb(n292),.dout(n294),.clk(gclk));
	jor g209(.dina(w_dff_B_9QPYehDS4_0),.dinb(n291),.dout(n295),.clk(gclk));
	jor g210(.dina(n295),.dinb(w_dff_B_uYfs2cxK6_1),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n285_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g212(.din(w_n285_0[0]),.dout(n298),.clk(gclk));
	jor g213(.dina(w_dff_B_uQCll2v58_0),.dinb(w_n258_0[0]),.dout(n299),.clk(gclk));
	jand g214(.dina(n299),.dinb(w_G219gat_2[2]),.dout(n300),.clk(gclk));
	jand g215(.dina(n300),.dinb(w_dff_B_FdyFEEuq6_1),.dout(n301),.clk(gclk));
	jor g216(.dina(n301),.dinb(w_dff_B_quorBJTR4_1),.dout(w_dff_A_i7fpZ1qg5_2),.clk(gclk));
	jand g217(.dina(w_n168_0[0]),.dinb(w_G55gat_0[0]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n303_1[1]),.dinb(w_G143gat_0[0]),.dout(n304),.clk(gclk));
	jand g219(.dina(w_n146_0[0]),.dinb(w_G17gat_1[0]),.dout(n305),.clk(gclk));
	jand g220(.dina(n305),.dinb(w_n144_0[0]),.dout(n306),.clk(gclk));
	jor g221(.dina(w_n306_1[1]),.dinb(w_dff_B_mf2zHNDT5_1),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n164_2[0]),.dinb(w_G91gat_0[1]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_gNuOt0Qh5_0),.dinb(n308),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(w_dff_B_CLxBbHRk0_1),.dout(n311),.clk(gclk));
	jand g226(.dina(w_n311_1[2]),.dinb(w_G159gat_1[1]),.dout(n312),.clk(gclk));
	jor g227(.dina(w_n311_1[1]),.dinb(w_G159gat_1[0]),.dout(n313),.clk(gclk));
	jand g228(.dina(w_n164_1[2]),.dinb(w_G96gat_0[1]),.dout(n314),.clk(gclk));
	jand g229(.dina(w_n303_1[0]),.dinb(w_G146gat_0[0]),.dout(n315),.clk(gclk));
	jand g230(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n316),.clk(gclk));
	jor g231(.dina(w_dff_B_sDlKO3YR9_0),.dinb(n315),.dout(n317),.clk(gclk));
	jor g232(.dina(w_dff_B_py9DwAIB7_0),.dinb(n314),.dout(n318),.clk(gclk));
	jor g233(.dina(n318),.dinb(w_n306_1[0]),.dout(n319),.clk(gclk));
	jand g234(.dina(w_n319_1[2]),.dinb(w_G165gat_1[1]),.dout(n320),.clk(gclk));
	jor g235(.dina(w_n319_1[1]),.dinb(w_G165gat_1[0]),.dout(n321),.clk(gclk));
	jand g236(.dina(w_n164_1[1]),.dinb(w_G101gat_0[1]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n303_0[2]),.dinb(w_G149gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n324),.clk(gclk));
	jor g239(.dina(w_dff_B_QzdtIJtd4_0),.dinb(n323),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_s45QQpiD1_0),.dinb(n322),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(w_n306_0[2]),.dout(n327),.clk(gclk));
	jand g242(.dina(w_n327_1[2]),.dinb(w_G171gat_1[1]),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n327_1[1]),.dinb(w_G171gat_1[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n164_1[0]),.dinb(w_G106gat_0[0]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n303_0[1]),.dinb(w_G153gat_0[0]),.dout(n331),.clk(gclk));
	jand g246(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n332),.clk(gclk));
	jor g247(.dina(w_dff_B_Kn1FYWoV5_0),.dinb(n331),.dout(n333),.clk(gclk));
	jor g248(.dina(w_dff_B_6GSYaz0e9_0),.dinb(n330),.dout(n334),.clk(gclk));
	jor g249(.dina(n334),.dinb(w_n306_0[1]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_1[1]),.dinb(w_G177gat_1[1]),.dout(n336),.clk(gclk));
	jnot g251(.din(w_G177gat_1[0]),.dout(n337),.clk(gclk));
	jnot g252(.din(w_n335_1[0]),.dout(n338),.clk(gclk));
	jand g253(.dina(n338),.dinb(w_dff_B_zRWcyhoV2_1),.dout(n339),.clk(gclk));
	jnot g254(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jnot g255(.din(w_G183gat_0[1]),.dout(n341),.clk(gclk));
	jnot g256(.din(w_n218_0[1]),.dout(n342),.clk(gclk));
	jand g257(.dina(n342),.dinb(w_dff_B_THrVAbF30_1),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n343_0[1]),.dout(n344),.clk(gclk));
	jand g259(.dina(w_n249_0[0]),.dinb(w_dff_B_vbu4v1jM8_1),.dout(n345),.clk(gclk));
	jor g260(.dina(n345),.dinb(w_n222_0[1]),.dout(n346),.clk(gclk));
	jand g261(.dina(w_n346_0[1]),.dinb(w_dff_B_8Q9L2Ugr5_1),.dout(n347),.clk(gclk));
	jor g262(.dina(n347),.dinb(w_n336_0[2]),.dout(n348),.clk(gclk));
	jand g263(.dina(w_n348_0[1]),.dinb(w_n329_0[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(n349),.dinb(w_n328_0[1]),.dout(n350),.clk(gclk));
	jand g265(.dina(w_n350_0[1]),.dinb(w_n321_0[1]),.dout(n351),.clk(gclk));
	jor g266(.dina(n351),.dinb(w_n320_0[1]),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n352_0[1]),.dinb(w_dff_B_G5W7pFqL9_1),.dout(n353),.clk(gclk));
	jor g268(.dina(n353),.dinb(w_dff_B_vSOUwK2N3_1),.dout(w_dff_A_uu90gjxu6_2),.clk(gclk));
	jxor g269(.dina(w_n335_0[2]),.dinb(w_G177gat_0[2]),.dout(n355),.clk(gclk));
	jnot g270(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n346_0[0]),.dinb(w_G219gat_2[1]),.dout(n357),.clk(gclk));
	jand g272(.dina(n357),.dinb(w_dff_B_bYpKujEX4_1),.dout(n358),.clk(gclk));
	jnot g273(.din(w_n222_0[0]),.dout(n359),.clk(gclk));
	jor g274(.dina(w_n262_0[0]),.dinb(w_n343_0[0]),.dout(n360),.clk(gclk));
	jand g275(.dina(n360),.dinb(w_dff_B_Y9ex9KpT5_1),.dout(n361),.clk(gclk));
	jand g276(.dina(w_n361_0[1]),.dinb(w_G219gat_2[0]),.dout(n362),.clk(gclk));
	jor g277(.dina(n362),.dinb(w_G228gat_2[0]),.dout(n363),.clk(gclk));
	jand g278(.dina(n363),.dinb(w_n355_0[0]),.dout(n364),.clk(gclk));
	jand g279(.dina(w_n336_0[1]),.dinb(w_G237gat_2[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_n335_0[1]),.dinb(w_G246gat_2[0]),.dout(n366),.clk(gclk));
	jand g281(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n367),.clk(gclk));
	jand g282(.dina(w_n178_2[0]),.dinb(w_G177gat_0[1]),.dout(n368),.clk(gclk));
	jor g283(.dina(n368),.dinb(w_dff_B_C2QS22wE8_1),.dout(n369),.clk(gclk));
	jor g284(.dina(w_dff_B_3ejL3m9E0_0),.dinb(n366),.dout(n370),.clk(gclk));
	jor g285(.dina(n370),.dinb(n365),.dout(n371),.clk(gclk));
	jor g286(.dina(w_dff_B_KIQzMffs8_0),.dinb(n364),.dout(n372),.clk(gclk));
	jor g287(.dina(n372),.dinb(w_dff_B_dDZMWDgu2_1),.dout(w_dff_A_59cdx3DS7_2),.clk(gclk));
	jand g288(.dina(w_n311_1[0]),.dinb(w_G237gat_1[2]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_n178_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(n375),.dinb(w_G159gat_0[2]),.dout(n376),.clk(gclk));
	jxor g291(.dina(w_n311_0[2]),.dinb(w_G159gat_0[1]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_n377_0[2]),.dinb(w_G228gat_1[2]),.dout(n378),.clk(gclk));
	jand g293(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_bwf0huTv8_0),.dinb(n378),.dout(n380),.clk(gclk));
	jand g295(.dina(w_n311_0[1]),.dinb(w_G246gat_1[2]),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_dhwGUi4C4_0),.dinb(n380),.dout(n382),.clk(gclk));
	jor g297(.dina(n382),.dinb(w_dff_B_TnSxArNL8_1),.dout(n383),.clk(gclk));
	jor g298(.dina(w_n377_0[1]),.dinb(w_n352_0[0]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n320_0[0]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n321_0[0]),.dout(n386),.clk(gclk));
	jnot g301(.din(w_n328_0[0]),.dout(n387),.clk(gclk));
	jnot g302(.din(w_n329_0[0]),.dout(n388),.clk(gclk));
	jnot g303(.din(w_n336_0[0]),.dout(n389),.clk(gclk));
	jor g304(.dina(w_n361_0[0]),.dinb(w_n339_0[0]),.dout(n390),.clk(gclk));
	jand g305(.dina(n390),.dinb(w_dff_B_9YbA9GZ99_1),.dout(n391),.clk(gclk));
	jor g306(.dina(w_n391_0[1]),.dinb(w_dff_B_A3NTip0I7_1),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_dff_B_BPEUKfMy0_1),.dout(n393),.clk(gclk));
	jor g308(.dina(w_n393_0[1]),.dinb(w_dff_B_ORnpkLBA5_1),.dout(n394),.clk(gclk));
	jand g309(.dina(n394),.dinb(w_dff_B_YkK2LiLL9_1),.dout(n395),.clk(gclk));
	jnot g310(.din(w_n377_0[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(w_dff_B_1H8axePV9_0),.dinb(n395),.dout(n397),.clk(gclk));
	jand g312(.dina(n397),.dinb(w_G219gat_1[2]),.dout(n398),.clk(gclk));
	jand g313(.dina(n398),.dinb(w_dff_B_mfXSlU7j1_1),.dout(n399),.clk(gclk));
	jor g314(.dina(n399),.dinb(w_dff_B_ijMSrt5x0_1),.dout(G878gat),.clk(gclk));
	jand g315(.dina(w_n319_1[0]),.dinb(w_G237gat_1[1]),.dout(n401),.clk(gclk));
	jor g316(.dina(n401),.dinb(w_n178_1[1]),.dout(n402),.clk(gclk));
	jand g317(.dina(n402),.dinb(w_G165gat_0[2]),.dout(n403),.clk(gclk));
	jxor g318(.dina(w_n319_0[2]),.dinb(w_G165gat_0[1]),.dout(n404),.clk(gclk));
	jand g319(.dina(w_n404_0[2]),.dinb(w_G228gat_1[1]),.dout(n405),.clk(gclk));
	jand g320(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n406),.clk(gclk));
	jor g321(.dina(w_dff_B_wTQ1267p5_0),.dinb(n405),.dout(n407),.clk(gclk));
	jand g322(.dina(w_n319_0[1]),.dinb(w_G246gat_1[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_6GQCrwjA3_0),.dinb(n407),.dout(n409),.clk(gclk));
	jor g324(.dina(n409),.dinb(w_dff_B_em656vaO0_1),.dout(n410),.clk(gclk));
	jor g325(.dina(w_n404_0[1]),.dinb(w_n350_0[0]),.dout(n411),.clk(gclk));
	jnot g326(.din(w_n404_0[0]),.dout(n412),.clk(gclk));
	jor g327(.dina(w_dff_B_2CBrTZA57_0),.dinb(w_n393_0[0]),.dout(n413),.clk(gclk));
	jand g328(.dina(n413),.dinb(w_G219gat_1[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_dff_B_mebxrYF86_1),.dout(n415),.clk(gclk));
	jor g330(.dina(n415),.dinb(w_dff_B_b77xlsdY5_1),.dout(w_dff_A_j2wVWtWp7_2),.clk(gclk));
	jand g331(.dina(w_n327_1[0]),.dinb(w_G237gat_1[0]),.dout(n417),.clk(gclk));
	jor g332(.dina(n417),.dinb(w_n178_1[0]),.dout(n418),.clk(gclk));
	jand g333(.dina(n418),.dinb(w_G171gat_0[2]),.dout(n419),.clk(gclk));
	jxor g334(.dina(w_n327_0[2]),.dinb(w_G171gat_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n420_0[2]),.dinb(w_G228gat_1[0]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_q5Ktwy8s3_0),.dinb(n421),.dout(n423),.clk(gclk));
	jand g338(.dina(w_n327_0[1]),.dinb(w_G246gat_1[0]),.dout(n424),.clk(gclk));
	jor g339(.dina(w_dff_B_guRjmfLS2_0),.dinb(n423),.dout(n425),.clk(gclk));
	jor g340(.dina(n425),.dinb(w_dff_B_9BWndEVS6_1),.dout(n426),.clk(gclk));
	jnot g341(.din(w_n420_0[1]),.dout(n427),.clk(gclk));
	jor g342(.dina(w_dff_B_bOfGwb3m3_0),.dinb(w_n391_0[0]),.dout(n428),.clk(gclk));
	jor g343(.dina(w_n420_0[0]),.dinb(w_n348_0[0]),.dout(n429),.clk(gclk));
	jand g344(.dina(n429),.dinb(w_G219gat_1[0]),.dout(n430),.clk(gclk));
	jand g345(.dina(n430),.dinb(w_dff_B_EwFU9vN70_1),.dout(n431),.clk(gclk));
	jor g346(.dina(n431),.dinb(w_dff_B_lvNTZ2L67_1),.dout(w_dff_A_yvuvlarN9_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_Lst0McxJ1_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_dff_A_QxIfccYM2_1),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_pLKY32TV0_0),.doutb(w_dff_A_tABhtonR0_1),.doutc(w_G17gat_1[2]),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_dff_A_uzkzW8UG4_2),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_6lqp49I31_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_fVb50uyJ6_1),.doutc(w_dff_A_FaerhiMT4_2),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_dff_A_7Xsqoc8r5_0),.doutb(w_G42gat_1[1]),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_udxixTEL4_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_egK1zrPp8_0),.doutb(w_dff_A_5WA9MwRB4_1),.doutc(w_G55gat_0[2]),.din(w_dff_B_lEMQTvZA9_3));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_dff_A_dADlnIYC6_1),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_fzqXj6HD0_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_gsqSXBtL6_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_pSUFoYvh7_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_i58d2qx50_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_Kq8CvxTw7_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_URmQRko84_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_cThWVYcY6_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_d6biRXab9_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_2O2Q4pOl4_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl3 jspl3_w_G126gat_0(.douta(w_G126gat_0[0]),.doutb(w_dff_A_IxPp00Gn2_1),.doutc(w_G126gat_0[2]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_dff_A_VbHs2Mun8_1),.din(G130gat));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_PH8TGeuR4_1),.din(w_dff_B_65QB3twe0_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_RgrZBGyU8_1),.din(w_dff_B_ELVxRGg83_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_VIBDWbqU0_1),.din(w_dff_B_rozhVQNP3_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_fWbf8oFC2_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_kiWkekqw1_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_dff_A_Cdh1RHdS9_1),.doutc(w_dff_A_ooxJvQMe3_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_dff_A_O8Vklup97_0),.doutb(w_dff_A_5rMxZFOJ6_1),.doutc(w_G159gat_1[2]),.din(w_G159gat_0[0]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_dff_A_D05oNxKZ1_1),.doutc(w_dff_A_ZuaxcF6B6_2),.din(w_dff_B_epr6vjWz6_3));
	jspl3 jspl3_w_G165gat_1(.douta(w_dff_A_e8Ofl2I68_0),.doutb(w_dff_A_gCsMnsrE5_1),.doutc(w_G165gat_1[2]),.din(w_G165gat_0[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_dff_A_aWmdXhqw4_1),.doutc(w_dff_A_YEa8x4XB1_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_dff_A_5UnxKDUu8_0),.doutb(w_dff_A_SDHk0Ayh3_1),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_dff_A_VewlEDL70_1),.doutc(w_dff_A_eyk3KoDE9_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_NT7xUXH68_1),.doutc(w_G177gat_1[2]),.din(w_G177gat_0[0]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_54e5qKsY5_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_SYl1ZTaK7_0),.doutb(w_dff_A_0099FcX74_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_OWu9GO5M9_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_JQ4JKKZN3_1),.doutc(w_dff_A_BONYvIGV9_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_15PxcqHD1_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_7I1OU8ZZ1_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_TKBNZ3Sl1_1),.doutc(w_dff_A_FKwPJQjV2_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_gzSCnwQh6_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_dff_A_DVUZWOLC3_1),.doutc(w_G201gat_0[2]),.din(G201gat));
	jspl jspl_w_G201gat_1(.douta(w_dff_A_jJiEuFvK4_0),.doutb(w_G201gat_1[1]),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_SfnO8thz7_0),.doutb(w_dff_A_sMiNjPDH1_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_kEi3TNjC8_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_dff_A_sqprAlgC0_1),.doutc(w_dff_A_4Sd4npID9_2),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_veE51J5r6_0),.doutb(w_dff_A_HdP8i38R0_1),.doutc(w_G219gat_2[2]),.din(w_G219gat_0[1]));
	jspl3 jspl3_w_G219gat_3(.douta(w_dff_A_cswhGIzL9_0),.doutb(w_dff_A_jC3o60vi7_1),.doutc(w_G219gat_3[2]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_dff_A_HlfwhfIe3_0),.doutb(w_G228gat_0[1]),.doutc(w_G228gat_0[2]),.din(w_dff_B_QR0EmBkX8_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_dff_A_XHTaupih4_0),.doutb(w_G228gat_2[1]),.doutc(w_G228gat_2[2]),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_dff_A_j14IaQH59_1),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_dff_A_JCmb31hf1_0),.doutb(w_G237gat_0[1]),.doutc(w_dff_A_5Xt0KupC1_2),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_dff_A_Gs7sp7nX6_0),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_dff_A_CXvq3uDD5_1),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_dff_A_pRmQpTHG9_0),.doutb(w_G246gat_0[1]),.doutc(w_dff_A_zoxLnd2T6_2),.din(w_dff_B_FbsYManE5_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_dff_A_h4gHO2iu9_0),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_dff_A_EAMIyyQt3_1),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_ccCzQTdh6_0),.doutb(w_G261gat_0[1]),.doutc(w_dff_A_TBAA5QPO6_2),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_6u0KVS2n6_1),.doutc(w_dff_A_DCUnLUjN5_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_dff_A_QRFb94mw6_2),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_bDsVM3Cz7_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_dff_A_ChJmihjf4_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_883qTqWJ8_0),.doutb(w_n95_0[1]),.doutc(w_dff_A_SWS8zYQ67_2),.din(n95));
	jspl jspl_w_n97_0(.douta(w_dff_A_6GAsQtzw5_0),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(w_dff_B_GSIaywte5_2));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_dff_A_FcRWR8m76_1),.din(n111));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.din(n113));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_QqoOc1Jz9_1),.din(n122));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_kzHPPf338_2));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.doutc(w_dff_A_yVEYHzL20_2),.din(w_n148_0[0]));
	jspl jspl_w_n149_0(.douta(w_dff_A_H2GZtF6F1_0),.doutb(w_n149_0[1]),.din(n149));
	jspl jspl_w_n151_0(.douta(w_dff_A_srPCK7nJ5_0),.doutb(w_n151_0[1]),.din(w_dff_B_Yh1MOgGx9_2));
	jspl jspl_w_n152_0(.douta(w_dff_A_cSLTPijy3_0),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n162_0(.douta(w_dff_A_3dL30TBv8_0),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_n164_1[0]),.doutb(w_n164_1[1]),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n164_2(.douta(w_n164_2[0]),.doutb(w_n164_2[1]),.doutc(w_n164_2[2]),.din(w_n164_0[1]));
	jspl jspl_w_n164_3(.douta(w_n164_3[0]),.doutb(w_n164_3[1]),.din(w_n164_0[2]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n170_1(.douta(w_n170_1[0]),.doutb(w_n170_1[1]),.din(w_n170_0[0]));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_nABzgguu0_0),.doutb(w_n178_0[1]),.doutc(w_n178_0[2]),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n178_2(.douta(w_n178_2[0]),.doutb(w_n178_2[1]),.doutc(w_n178_2[2]),.din(w_n178_0[1]));
	jspl jspl_w_n178_3(.douta(w_n178_3[0]),.doutb(w_n178_3[1]),.din(w_n178_0[2]));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(w_dff_B_juyi9VzG8_3));
	jspl jspl_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.din(n185));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_r3WANGgp2_1),.din(w_dff_B_OnztqHNG8_2));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_HzVUopj19_1),.doutc(w_n219_0[2]),.din(n219));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_dff_A_uyfWmlS52_1),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_k3roUDba9_1),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_dff_A_CB2CKF6I5_1),.din(n235));
	jspl3 jspl3_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.doutc(w_n239_0[2]),.din(n239));
	jspl jspl_w_n239_1(.douta(w_n239_1[0]),.doutb(w_n239_1[1]),.din(w_n239_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_dff_A_P4zV80J80_1),.din(n240));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_dff_A_HtD9ivyS4_1),.din(n241));
	jspl jspl_w_n242_0(.douta(w_dff_A_DB211iR03_0),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_dff_A_Ld9vuEK63_1),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_dff_A_KWSQz0Ql4_1),.doutc(w_n285_0[2]),.din(n285));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl jspl_w_n303_1(.douta(w_n303_1[0]),.doutb(w_n303_1[1]),.din(w_n303_0[0]));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_dff_A_WZEDCsWq4_1),.doutc(w_dff_A_vg7FDJnQ3_2),.din(n306));
	jspl jspl_w_n306_1(.douta(w_dff_A_6ZGK6Eos5_0),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n311_1(.douta(w_n311_1[0]),.doutb(w_n311_1[1]),.doutc(w_n311_1[2]),.din(w_n311_0[0]));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(n319));
	jspl3 jspl3_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.doutc(w_n319_1[2]),.din(w_n319_0[0]));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_dff_A_pcKRiF3c5_1),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_uy3vY4jq6_1),.din(n321));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_dff_A_GAhtxgvl0_1),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_dff_A_g1NKNY736_1),.din(n329));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl jspl_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.din(w_n335_0[0]));
	jspl3 jspl3_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.doutc(w_dff_A_SexcC3WA1_2),.din(n336));
	jspl jspl_w_n339_0(.douta(w_dff_A_lyr1kNRw7_0),.doutb(w_n339_0[1]),.din(n339));
	jspl jspl_w_n343_0(.douta(w_dff_A_SfACn2Ng8_0),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.din(n352));
	jspl jspl_w_n355_0(.douta(w_dff_A_WTmwzHhH3_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_L9BAJdW84_1),.doutc(w_n377_0[2]),.din(n377));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_dff_A_Xa5F2hGi1_1),.doutc(w_n404_0[2]),.din(n404));
	jspl3 jspl3_w_n420_0(.douta(w_dff_A_H1gPzLXb4_0),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jdff dff_B_GSIaywte5_2(.din(n103),.dout(w_dff_B_GSIaywte5_2),.clk(gclk));
	jdff dff_B_tAReGijg0_1(.din(G90gat),.dout(w_dff_B_tAReGijg0_1),.clk(gclk));
	jdff dff_B_zHSEY54C2_1(.din(n115),.dout(w_dff_B_zHSEY54C2_1),.clk(gclk));
	jdff dff_B_kiZvJ92o9_1(.din(n96),.dout(w_dff_B_kiZvJ92o9_1),.clk(gclk));
	jdff dff_A_xHbkrqDb3_1(.dout(w_G390gat_0[1]),.din(w_dff_A_xHbkrqDb3_1),.clk(gclk));
	jdff dff_A_6u0KVS2n6_1(.dout(w_dff_A_xHbkrqDb3_1),.din(w_dff_A_6u0KVS2n6_1),.clk(gclk));
	jdff dff_B_p7UUrr9R3_1(.din(G74gat),.dout(w_dff_B_p7UUrr9R3_1),.clk(gclk));
	jdff dff_B_N3gDhnya0_1(.din(w_dff_B_p7UUrr9R3_1),.dout(w_dff_B_N3gDhnya0_1),.clk(gclk));
	jdff dff_B_kggM7kW44_1(.din(w_dff_B_N3gDhnya0_1),.dout(w_dff_B_kggM7kW44_1),.clk(gclk));
	jdff dff_B_qVLElNTY8_1(.din(G89gat),.dout(w_dff_B_qVLElNTY8_1),.clk(gclk));
	jdff dff_B_rs6GoOFe1_1(.din(n127),.dout(w_dff_B_rs6GoOFe1_1),.clk(gclk));
	jdff dff_B_IYnRNLZA4_1(.din(G135gat),.dout(w_dff_B_IYnRNLZA4_1),.clk(gclk));
	jdff dff_B_CaTEttEE8_1(.din(n136),.dout(w_dff_B_CaTEttEE8_1),.clk(gclk));
	jdff dff_A_VbHs2Mun8_1(.dout(w_G130gat_0[1]),.din(w_dff_A_VbHs2Mun8_1),.clk(gclk));
	jdff dff_B_xZ4cSpAA9_1(.din(G207gat),.dout(w_dff_B_xZ4cSpAA9_1),.clk(gclk));
	jdff dff_B_MsViwyTq7_1(.din(n208),.dout(w_dff_B_MsViwyTq7_1),.clk(gclk));
	jdff dff_B_KBWPjDHB7_1(.din(w_dff_B_MsViwyTq7_1),.dout(w_dff_B_KBWPjDHB7_1),.clk(gclk));
	jdff dff_B_lBXbOrwb0_1(.din(n180),.dout(w_dff_B_lBXbOrwb0_1),.clk(gclk));
	jdff dff_B_ZpbdFtNi8_1(.din(w_dff_B_lBXbOrwb0_1),.dout(w_dff_B_ZpbdFtNi8_1),.clk(gclk));
	jdff dff_B_EPAe0jse5_1(.din(n199),.dout(w_dff_B_EPAe0jse5_1),.clk(gclk));
	jdff dff_B_yeiXuvcf0_0(.din(n204),.dout(w_dff_B_yeiXuvcf0_0),.clk(gclk));
	jdff dff_B_UGuoYXmm1_0(.din(w_dff_B_yeiXuvcf0_0),.dout(w_dff_B_UGuoYXmm1_0),.clk(gclk));
	jdff dff_B_NiLdjS6E0_0(.din(w_dff_B_UGuoYXmm1_0),.dout(w_dff_B_NiLdjS6E0_0),.clk(gclk));
	jdff dff_B_iODpJsBp4_0(.din(w_dff_B_NiLdjS6E0_0),.dout(w_dff_B_iODpJsBp4_0),.clk(gclk));
	jdff dff_B_CqEcUHpB6_0(.din(w_dff_B_iODpJsBp4_0),.dout(w_dff_B_CqEcUHpB6_0),.clk(gclk));
	jdff dff_B_13NRcRbk2_0(.din(w_dff_B_CqEcUHpB6_0),.dout(w_dff_B_13NRcRbk2_0),.clk(gclk));
	jdff dff_B_PRsgJq3f1_0(.din(w_dff_B_13NRcRbk2_0),.dout(w_dff_B_PRsgJq3f1_0),.clk(gclk));
	jdff dff_B_ldYpc67U9_0(.din(w_dff_B_PRsgJq3f1_0),.dout(w_dff_B_ldYpc67U9_0),.clk(gclk));
	jdff dff_B_qzjTKzz27_0(.din(w_dff_B_ldYpc67U9_0),.dout(w_dff_B_qzjTKzz27_0),.clk(gclk));
	jdff dff_B_4Awn7C4E9_0(.din(n179),.dout(w_dff_B_4Awn7C4E9_0),.clk(gclk));
	jdff dff_B_7yALASj83_0(.din(w_dff_B_4Awn7C4E9_0),.dout(w_dff_B_7yALASj83_0),.clk(gclk));
	jdff dff_B_RU1Eypu97_0(.din(w_dff_B_7yALASj83_0),.dout(w_dff_B_RU1Eypu97_0),.clk(gclk));
	jdff dff_B_aDLR7Kvq2_0(.din(w_dff_B_RU1Eypu97_0),.dout(w_dff_B_aDLR7Kvq2_0),.clk(gclk));
	jdff dff_B_glchsX2h6_0(.din(w_dff_B_aDLR7Kvq2_0),.dout(w_dff_B_glchsX2h6_0),.clk(gclk));
	jdff dff_A_lbbwU5MU8_0(.dout(w_G201gat_1[0]),.din(w_dff_A_lbbwU5MU8_0),.clk(gclk));
	jdff dff_A_ovymAdQG1_0(.dout(w_dff_A_lbbwU5MU8_0),.din(w_dff_A_ovymAdQG1_0),.clk(gclk));
	jdff dff_A_SmruBy2C7_0(.dout(w_dff_A_ovymAdQG1_0),.din(w_dff_A_SmruBy2C7_0),.clk(gclk));
	jdff dff_A_jJiEuFvK4_0(.dout(w_dff_A_SmruBy2C7_0),.din(w_dff_A_jJiEuFvK4_0),.clk(gclk));
	jdff dff_B_KRXK0BIK7_1(.din(n229),.dout(w_dff_B_KRXK0BIK7_1),.clk(gclk));
	jdff dff_B_JS8AxjnQ2_1(.din(w_dff_B_KRXK0BIK7_1),.dout(w_dff_B_JS8AxjnQ2_1),.clk(gclk));
	jdff dff_B_CcigUWsG8_1(.din(w_dff_B_JS8AxjnQ2_1),.dout(w_dff_B_CcigUWsG8_1),.clk(gclk));
	jdff dff_B_Y30hR4Xq7_1(.din(w_dff_B_CcigUWsG8_1),.dout(w_dff_B_Y30hR4Xq7_1),.clk(gclk));
	jdff dff_B_cmC4qDUJ6_1(.din(w_dff_B_Y30hR4Xq7_1),.dout(w_dff_B_cmC4qDUJ6_1),.clk(gclk));
	jdff dff_B_4rqCsIZw9_1(.din(w_dff_B_cmC4qDUJ6_1),.dout(w_dff_B_4rqCsIZw9_1),.clk(gclk));
	jdff dff_B_fDhPSzWG5_1(.din(n250),.dout(w_dff_B_fDhPSzWG5_1),.clk(gclk));
	jdff dff_B_5tPrt5TS0_1(.din(n251),.dout(w_dff_B_5tPrt5TS0_1),.clk(gclk));
	jdff dff_B_DMUQEEkT6_1(.din(w_dff_B_5tPrt5TS0_1),.dout(w_dff_B_DMUQEEkT6_1),.clk(gclk));
	jdff dff_B_5RxU2FrA5_1(.din(w_dff_B_DMUQEEkT6_1),.dout(w_dff_B_5RxU2FrA5_1),.clk(gclk));
	jdff dff_B_dQ96iAXH6_1(.din(w_dff_B_5RxU2FrA5_1),.dout(w_dff_B_dQ96iAXH6_1),.clk(gclk));
	jdff dff_B_8yNUeOwK7_1(.din(w_dff_B_dQ96iAXH6_1),.dout(w_dff_B_8yNUeOwK7_1),.clk(gclk));
	jdff dff_B_7UJ5sV2m1_1(.din(w_dff_B_8yNUeOwK7_1),.dout(w_dff_B_7UJ5sV2m1_1),.clk(gclk));
	jdff dff_B_6pSDPMc78_1(.din(n220),.dout(w_dff_B_6pSDPMc78_1),.clk(gclk));
	jdff dff_B_7gnwILmQ9_1(.din(w_dff_B_6pSDPMc78_1),.dout(w_dff_B_7gnwILmQ9_1),.clk(gclk));
	jdff dff_B_9AMMAbma1_1(.din(n221),.dout(w_dff_B_9AMMAbma1_1),.clk(gclk));
	jdff dff_B_RMJa3JFY2_1(.din(w_dff_B_9AMMAbma1_1),.dout(w_dff_B_RMJa3JFY2_1),.clk(gclk));
	jdff dff_B_V2HBIQJY9_1(.din(w_dff_B_RMJa3JFY2_1),.dout(w_dff_B_V2HBIQJY9_1),.clk(gclk));
	jdff dff_B_7TXgyzlL9_1(.din(w_dff_B_V2HBIQJY9_1),.dout(w_dff_B_7TXgyzlL9_1),.clk(gclk));
	jdff dff_B_jQkrUx4e0_1(.din(w_dff_B_7TXgyzlL9_1),.dout(w_dff_B_jQkrUx4e0_1),.clk(gclk));
	jdff dff_B_84n8DlGf3_1(.din(w_dff_B_jQkrUx4e0_1),.dout(w_dff_B_84n8DlGf3_1),.clk(gclk));
	jdff dff_B_uIXJncuN6_0(.din(n225),.dout(w_dff_B_uIXJncuN6_0),.clk(gclk));
	jdff dff_B_oVL95WD29_0(.din(w_dff_B_uIXJncuN6_0),.dout(w_dff_B_oVL95WD29_0),.clk(gclk));
	jdff dff_B_BEQmc9da3_0(.din(w_dff_B_oVL95WD29_0),.dout(w_dff_B_BEQmc9da3_0),.clk(gclk));
	jdff dff_B_mzBl8A180_0(.din(w_dff_B_BEQmc9da3_0),.dout(w_dff_B_mzBl8A180_0),.clk(gclk));
	jdff dff_B_ff64FpwW7_0(.din(w_dff_B_mzBl8A180_0),.dout(w_dff_B_ff64FpwW7_0),.clk(gclk));
	jdff dff_B_YFBtf0H28_0(.din(w_dff_B_ff64FpwW7_0),.dout(w_dff_B_YFBtf0H28_0),.clk(gclk));
	jdff dff_B_nqqmaY0D9_0(.din(w_dff_B_YFBtf0H28_0),.dout(w_dff_B_nqqmaY0D9_0),.clk(gclk));
	jdff dff_B_7PLyaIN99_0(.din(w_dff_B_nqqmaY0D9_0),.dout(w_dff_B_7PLyaIN99_0),.clk(gclk));
	jdff dff_A_EAMIyyQt3_1(.dout(w_G246gat_3[1]),.din(w_dff_A_EAMIyyQt3_1),.clk(gclk));
	jdff dff_A_CXvq3uDD5_1(.dout(w_G237gat_3[1]),.din(w_dff_A_CXvq3uDD5_1),.clk(gclk));
	jdff dff_A_RKnVw1t78_1(.dout(w_n219_0[1]),.din(w_dff_A_RKnVw1t78_1),.clk(gclk));
	jdff dff_A_LS30gOEK1_1(.dout(w_dff_A_RKnVw1t78_1),.din(w_dff_A_LS30gOEK1_1),.clk(gclk));
	jdff dff_A_XCbuhe4z0_1(.dout(w_dff_A_LS30gOEK1_1),.din(w_dff_A_XCbuhe4z0_1),.clk(gclk));
	jdff dff_A_JtT7Xivj8_1(.dout(w_dff_A_XCbuhe4z0_1),.din(w_dff_A_JtT7Xivj8_1),.clk(gclk));
	jdff dff_A_YIUMp9I11_1(.dout(w_dff_A_JtT7Xivj8_1),.din(w_dff_A_YIUMp9I11_1),.clk(gclk));
	jdff dff_A_qgTNje5x7_1(.dout(w_dff_A_YIUMp9I11_1),.din(w_dff_A_qgTNje5x7_1),.clk(gclk));
	jdff dff_A_HzVUopj19_1(.dout(w_dff_A_qgTNje5x7_1),.din(w_dff_A_HzVUopj19_1),.clk(gclk));
	jdff dff_A_IaniZYls9_0(.dout(w_G183gat_1[0]),.din(w_dff_A_IaniZYls9_0),.clk(gclk));
	jdff dff_A_o46JxSdL2_0(.dout(w_dff_A_IaniZYls9_0),.din(w_dff_A_o46JxSdL2_0),.clk(gclk));
	jdff dff_A_8hignWYJ0_0(.dout(w_dff_A_o46JxSdL2_0),.din(w_dff_A_8hignWYJ0_0),.clk(gclk));
	jdff dff_A_SYl1ZTaK7_0(.dout(w_dff_A_8hignWYJ0_0),.din(w_dff_A_SYl1ZTaK7_0),.clk(gclk));
	jdff dff_A_foXrpMJg4_1(.dout(w_G183gat_1[1]),.din(w_dff_A_foXrpMJg4_1),.clk(gclk));
	jdff dff_A_QQFj4ndL4_1(.dout(w_dff_A_foXrpMJg4_1),.din(w_dff_A_QQFj4ndL4_1),.clk(gclk));
	jdff dff_A_0uaWIG1l7_1(.dout(w_dff_A_QQFj4ndL4_1),.din(w_dff_A_0uaWIG1l7_1),.clk(gclk));
	jdff dff_A_NLAVdITU2_1(.dout(w_dff_A_0uaWIG1l7_1),.din(w_dff_A_NLAVdITU2_1),.clk(gclk));
	jdff dff_A_ODHcvoO50_1(.dout(w_dff_A_NLAVdITU2_1),.din(w_dff_A_ODHcvoO50_1),.clk(gclk));
	jdff dff_A_dGtI2dac5_1(.dout(w_dff_A_ODHcvoO50_1),.din(w_dff_A_dGtI2dac5_1),.clk(gclk));
	jdff dff_A_84Y2JVtx4_1(.dout(w_dff_A_dGtI2dac5_1),.din(w_dff_A_84Y2JVtx4_1),.clk(gclk));
	jdff dff_A_0099FcX74_1(.dout(w_dff_A_84Y2JVtx4_1),.din(w_dff_A_0099FcX74_1),.clk(gclk));
	jdff dff_A_j14IaQH59_1(.dout(w_G228gat_3[1]),.din(w_dff_A_j14IaQH59_1),.clk(gclk));
	jdff dff_B_tPIYVKvH9_1(.din(n278),.dout(w_dff_B_tPIYVKvH9_1),.clk(gclk));
	jdff dff_B_F0f1ClMC4_1(.din(w_dff_B_tPIYVKvH9_1),.dout(w_dff_B_F0f1ClMC4_1),.clk(gclk));
	jdff dff_B_A932LBmu1_1(.din(w_dff_B_F0f1ClMC4_1),.dout(w_dff_B_A932LBmu1_1),.clk(gclk));
	jdff dff_B_ijtp4fIJ1_1(.din(w_dff_B_A932LBmu1_1),.dout(w_dff_B_ijtp4fIJ1_1),.clk(gclk));
	jdff dff_B_lTkxRn4p5_1(.din(w_dff_B_ijtp4fIJ1_1),.dout(w_dff_B_lTkxRn4p5_1),.clk(gclk));
	jdff dff_B_FU6iXRqU8_1(.din(n279),.dout(w_dff_B_FU6iXRqU8_1),.clk(gclk));
	jdff dff_B_Hu5j9bju6_0(.din(n280),.dout(w_dff_B_Hu5j9bju6_0),.clk(gclk));
	jdff dff_B_TLrXwqyY7_0(.din(w_dff_B_Hu5j9bju6_0),.dout(w_dff_B_TLrXwqyY7_0),.clk(gclk));
	jdff dff_B_P7XkTJJ67_0(.din(w_dff_B_TLrXwqyY7_0),.dout(w_dff_B_P7XkTJJ67_0),.clk(gclk));
	jdff dff_B_JIUTpmJ50_0(.din(w_dff_B_P7XkTJJ67_0),.dout(w_dff_B_JIUTpmJ50_0),.clk(gclk));
	jdff dff_A_jO3Qq5u22_0(.dout(w_G219gat_3[0]),.din(w_dff_A_jO3Qq5u22_0),.clk(gclk));
	jdff dff_A_I47TRL0K7_0(.dout(w_dff_A_jO3Qq5u22_0),.din(w_dff_A_I47TRL0K7_0),.clk(gclk));
	jdff dff_A_cswhGIzL9_0(.dout(w_dff_A_I47TRL0K7_0),.din(w_dff_A_cswhGIzL9_0),.clk(gclk));
	jdff dff_A_aF2RwkzK0_1(.dout(w_G219gat_3[1]),.din(w_dff_A_aF2RwkzK0_1),.clk(gclk));
	jdff dff_A_PVgGCB742_1(.dout(w_dff_A_aF2RwkzK0_1),.din(w_dff_A_PVgGCB742_1),.clk(gclk));
	jdff dff_A_HcTM1GVX3_1(.dout(w_dff_A_PVgGCB742_1),.din(w_dff_A_HcTM1GVX3_1),.clk(gclk));
	jdff dff_A_kEdOAhc04_1(.dout(w_dff_A_HcTM1GVX3_1),.din(w_dff_A_kEdOAhc04_1),.clk(gclk));
	jdff dff_A_jC3o60vi7_1(.dout(w_dff_A_kEdOAhc04_1),.din(w_dff_A_jC3o60vi7_1),.clk(gclk));
	jdff dff_B_s73pqaah1_1(.din(n268),.dout(w_dff_B_s73pqaah1_1),.clk(gclk));
	jdff dff_B_nn6wMOGk0_0(.din(n276),.dout(w_dff_B_nn6wMOGk0_0),.clk(gclk));
	jdff dff_B_7cjJs6LO5_0(.din(w_dff_B_nn6wMOGk0_0),.dout(w_dff_B_7cjJs6LO5_0),.clk(gclk));
	jdff dff_B_20CebZ979_0(.din(w_dff_B_7cjJs6LO5_0),.dout(w_dff_B_20CebZ979_0),.clk(gclk));
	jdff dff_B_6E7KgVIu3_0(.din(w_dff_B_20CebZ979_0),.dout(w_dff_B_6E7KgVIu3_0),.clk(gclk));
	jdff dff_B_9r22lERW4_1(.din(n274),.dout(w_dff_B_9r22lERW4_1),.clk(gclk));
	jdff dff_B_OmeFB6pZ1_1(.din(w_dff_B_9r22lERW4_1),.dout(w_dff_B_OmeFB6pZ1_1),.clk(gclk));
	jdff dff_B_H0zx1ZtW2_1(.din(w_dff_B_OmeFB6pZ1_1),.dout(w_dff_B_H0zx1ZtW2_1),.clk(gclk));
	jdff dff_B_3ZMkq8Hj4_1(.din(w_dff_B_H0zx1ZtW2_1),.dout(w_dff_B_3ZMkq8Hj4_1),.clk(gclk));
	jdff dff_B_x3DtjL5f7_1(.din(n269),.dout(w_dff_B_x3DtjL5f7_1),.clk(gclk));
	jdff dff_B_1a2TZAgG4_1(.din(w_dff_B_x3DtjL5f7_1),.dout(w_dff_B_1a2TZAgG4_1),.clk(gclk));
	jdff dff_B_Y1cVy0MP9_1(.din(w_dff_B_1a2TZAgG4_1),.dout(w_dff_B_Y1cVy0MP9_1),.clk(gclk));
	jdff dff_B_D8OM8Dun0_1(.din(w_dff_B_Y1cVy0MP9_1),.dout(w_dff_B_D8OM8Dun0_1),.clk(gclk));
	jdff dff_B_nomCx90E8_1(.din(w_dff_B_D8OM8Dun0_1),.dout(w_dff_B_nomCx90E8_1),.clk(gclk));
	jdff dff_B_rBgMgBtT9_1(.din(w_dff_B_nomCx90E8_1),.dout(w_dff_B_rBgMgBtT9_1),.clk(gclk));
	jdff dff_B_WCr7dEsS6_1(.din(w_dff_B_rBgMgBtT9_1),.dout(w_dff_B_WCr7dEsS6_1),.clk(gclk));
	jdff dff_B_eALMfTKs8_1(.din(w_dff_B_WCr7dEsS6_1),.dout(w_dff_B_eALMfTKs8_1),.clk(gclk));
	jdff dff_B_WS4odQnb5_0(.din(n271),.dout(w_dff_B_WS4odQnb5_0),.clk(gclk));
	jdff dff_B_iQF6CmOP3_0(.din(w_dff_B_WS4odQnb5_0),.dout(w_dff_B_iQF6CmOP3_0),.clk(gclk));
	jdff dff_B_eNyofXta8_0(.din(w_dff_B_iQF6CmOP3_0),.dout(w_dff_B_eNyofXta8_0),.clk(gclk));
	jdff dff_B_5LYf5VqB1_0(.din(w_dff_B_eNyofXta8_0),.dout(w_dff_B_5LYf5VqB1_0),.clk(gclk));
	jdff dff_B_mXgbvMDp2_0(.din(w_dff_B_5LYf5VqB1_0),.dout(w_dff_B_mXgbvMDp2_0),.clk(gclk));
	jdff dff_B_XpaDHBzu2_0(.din(w_dff_B_mXgbvMDp2_0),.dout(w_dff_B_XpaDHBzu2_0),.clk(gclk));
	jdff dff_A_ma28hyni2_1(.dout(w_n267_0[1]),.din(w_dff_A_ma28hyni2_1),.clk(gclk));
	jdff dff_A_ryLF9ho38_1(.dout(w_dff_A_ma28hyni2_1),.din(w_dff_A_ryLF9ho38_1),.clk(gclk));
	jdff dff_A_MICi2kaS5_1(.dout(w_dff_A_ryLF9ho38_1),.din(w_dff_A_MICi2kaS5_1),.clk(gclk));
	jdff dff_A_oPYePDtu1_1(.dout(w_dff_A_MICi2kaS5_1),.din(w_dff_A_oPYePDtu1_1),.clk(gclk));
	jdff dff_A_Ld9vuEK63_1(.dout(w_dff_A_oPYePDtu1_1),.din(w_dff_A_Ld9vuEK63_1),.clk(gclk));
	jdff dff_B_sv0h8F5G0_1(.din(n296),.dout(w_dff_B_sv0h8F5G0_1),.clk(gclk));
	jdff dff_B_doZbIsdq4_1(.din(w_dff_B_sv0h8F5G0_1),.dout(w_dff_B_doZbIsdq4_1),.clk(gclk));
	jdff dff_B_quorBJTR4_1(.din(w_dff_B_doZbIsdq4_1),.dout(w_dff_B_quorBJTR4_1),.clk(gclk));
	jdff dff_B_FdyFEEuq6_1(.din(n297),.dout(w_dff_B_FdyFEEuq6_1),.clk(gclk));
	jdff dff_B_yFZnzdM23_0(.din(n298),.dout(w_dff_B_yFZnzdM23_0),.clk(gclk));
	jdff dff_B_uQCll2v58_0(.din(w_dff_B_yFZnzdM23_0),.dout(w_dff_B_uQCll2v58_0),.clk(gclk));
	jdff dff_B_uYfs2cxK6_1(.din(n286),.dout(w_dff_B_uYfs2cxK6_1),.clk(gclk));
	jdff dff_B_hQhrmT7l8_0(.din(n294),.dout(w_dff_B_hQhrmT7l8_0),.clk(gclk));
	jdff dff_B_vqXqbZSx8_0(.din(w_dff_B_hQhrmT7l8_0),.dout(w_dff_B_vqXqbZSx8_0),.clk(gclk));
	jdff dff_B_zCUSekvJ1_0(.din(w_dff_B_vqXqbZSx8_0),.dout(w_dff_B_zCUSekvJ1_0),.clk(gclk));
	jdff dff_B_9QPYehDS4_0(.din(w_dff_B_zCUSekvJ1_0),.dout(w_dff_B_9QPYehDS4_0),.clk(gclk));
	jdff dff_B_pfDKVsB08_0(.din(n293),.dout(w_dff_B_pfDKVsB08_0),.clk(gclk));
	jdff dff_B_N6L8NkBI2_0(.din(w_dff_B_pfDKVsB08_0),.dout(w_dff_B_N6L8NkBI2_0),.clk(gclk));
	jdff dff_B_itdv4hEJ5_0(.din(w_dff_B_N6L8NkBI2_0),.dout(w_dff_B_itdv4hEJ5_0),.clk(gclk));
	jdff dff_B_pg4cL8EJ9_0(.din(w_dff_B_itdv4hEJ5_0),.dout(w_dff_B_pg4cL8EJ9_0),.clk(gclk));
	jdff dff_B_A16QuiJk1_1(.din(n287),.dout(w_dff_B_A16QuiJk1_1),.clk(gclk));
	jdff dff_B_D1GtwHkq2_1(.din(w_dff_B_A16QuiJk1_1),.dout(w_dff_B_D1GtwHkq2_1),.clk(gclk));
	jdff dff_B_lbCEY3NP1_1(.din(w_dff_B_D1GtwHkq2_1),.dout(w_dff_B_lbCEY3NP1_1),.clk(gclk));
	jdff dff_B_TY17PhMk2_1(.din(w_dff_B_lbCEY3NP1_1),.dout(w_dff_B_TY17PhMk2_1),.clk(gclk));
	jdff dff_B_BJwEZ6133_1(.din(w_dff_B_TY17PhMk2_1),.dout(w_dff_B_BJwEZ6133_1),.clk(gclk));
	jdff dff_B_dDcipXBN9_1(.din(w_dff_B_BJwEZ6133_1),.dout(w_dff_B_dDcipXBN9_1),.clk(gclk));
	jdff dff_B_6OVoBhBC5_1(.din(w_dff_B_dDcipXBN9_1),.dout(w_dff_B_6OVoBhBC5_1),.clk(gclk));
	jdff dff_B_Cx9viwQK4_1(.din(w_dff_B_6OVoBhBC5_1),.dout(w_dff_B_Cx9viwQK4_1),.clk(gclk));
	jdff dff_B_KKr6Xmht4_0(.din(n289),.dout(w_dff_B_KKr6Xmht4_0),.clk(gclk));
	jdff dff_B_oFbHHbPU4_0(.din(w_dff_B_KKr6Xmht4_0),.dout(w_dff_B_oFbHHbPU4_0),.clk(gclk));
	jdff dff_B_IJ1xQlMV2_0(.din(w_dff_B_oFbHHbPU4_0),.dout(w_dff_B_IJ1xQlMV2_0),.clk(gclk));
	jdff dff_B_XSdgvg7a2_0(.din(w_dff_B_IJ1xQlMV2_0),.dout(w_dff_B_XSdgvg7a2_0),.clk(gclk));
	jdff dff_B_WGeQ4lVH4_0(.din(w_dff_B_XSdgvg7a2_0),.dout(w_dff_B_WGeQ4lVH4_0),.clk(gclk));
	jdff dff_B_Cy6GudwD7_0(.din(w_dff_B_WGeQ4lVH4_0),.dout(w_dff_B_Cy6GudwD7_0),.clk(gclk));
	jdff dff_A_A6pBvmPj2_1(.dout(w_n285_0[1]),.din(w_dff_A_A6pBvmPj2_1),.clk(gclk));
	jdff dff_A_uSC7OrEy1_1(.dout(w_dff_A_A6pBvmPj2_1),.din(w_dff_A_uSC7OrEy1_1),.clk(gclk));
	jdff dff_A_KWSQz0Ql4_1(.dout(w_dff_A_uSC7OrEy1_1),.din(w_dff_A_KWSQz0Ql4_1),.clk(gclk));
	jdff dff_B_Rbgx2vm75_1(.din(n312),.dout(w_dff_B_Rbgx2vm75_1),.clk(gclk));
	jdff dff_B_3eNKzKk52_1(.din(w_dff_B_Rbgx2vm75_1),.dout(w_dff_B_3eNKzKk52_1),.clk(gclk));
	jdff dff_B_AzUGH2hI5_1(.din(w_dff_B_3eNKzKk52_1),.dout(w_dff_B_AzUGH2hI5_1),.clk(gclk));
	jdff dff_B_ml8j43294_1(.din(w_dff_B_AzUGH2hI5_1),.dout(w_dff_B_ml8j43294_1),.clk(gclk));
	jdff dff_B_VakEVg175_1(.din(w_dff_B_ml8j43294_1),.dout(w_dff_B_VakEVg175_1),.clk(gclk));
	jdff dff_B_20wcC6Ne3_1(.din(w_dff_B_VakEVg175_1),.dout(w_dff_B_20wcC6Ne3_1),.clk(gclk));
	jdff dff_B_g8o3Zviv8_1(.din(w_dff_B_20wcC6Ne3_1),.dout(w_dff_B_g8o3Zviv8_1),.clk(gclk));
	jdff dff_B_5cFhrUcq6_1(.din(w_dff_B_g8o3Zviv8_1),.dout(w_dff_B_5cFhrUcq6_1),.clk(gclk));
	jdff dff_B_QKePrQ611_1(.din(w_dff_B_5cFhrUcq6_1),.dout(w_dff_B_QKePrQ611_1),.clk(gclk));
	jdff dff_B_ghwV2H0S0_1(.din(w_dff_B_QKePrQ611_1),.dout(w_dff_B_ghwV2H0S0_1),.clk(gclk));
	jdff dff_B_eJ50nooN0_1(.din(w_dff_B_ghwV2H0S0_1),.dout(w_dff_B_eJ50nooN0_1),.clk(gclk));
	jdff dff_B_HEUlk5BE9_1(.din(w_dff_B_eJ50nooN0_1),.dout(w_dff_B_HEUlk5BE9_1),.clk(gclk));
	jdff dff_B_voHXs2Qa4_1(.din(w_dff_B_HEUlk5BE9_1),.dout(w_dff_B_voHXs2Qa4_1),.clk(gclk));
	jdff dff_B_8r6bEAey5_1(.din(w_dff_B_voHXs2Qa4_1),.dout(w_dff_B_8r6bEAey5_1),.clk(gclk));
	jdff dff_B_vSOUwK2N3_1(.din(w_dff_B_8r6bEAey5_1),.dout(w_dff_B_vSOUwK2N3_1),.clk(gclk));
	jdff dff_B_efrgUlBb8_1(.din(n313),.dout(w_dff_B_efrgUlBb8_1),.clk(gclk));
	jdff dff_B_fFyNbHDS8_1(.din(w_dff_B_efrgUlBb8_1),.dout(w_dff_B_fFyNbHDS8_1),.clk(gclk));
	jdff dff_B_LbgnQHev8_1(.din(w_dff_B_fFyNbHDS8_1),.dout(w_dff_B_LbgnQHev8_1),.clk(gclk));
	jdff dff_B_P8gRLnd94_1(.din(w_dff_B_LbgnQHev8_1),.dout(w_dff_B_P8gRLnd94_1),.clk(gclk));
	jdff dff_B_JeXEp6s22_1(.din(w_dff_B_P8gRLnd94_1),.dout(w_dff_B_JeXEp6s22_1),.clk(gclk));
	jdff dff_B_cK3e9Z3T8_1(.din(w_dff_B_JeXEp6s22_1),.dout(w_dff_B_cK3e9Z3T8_1),.clk(gclk));
	jdff dff_B_BUnj0QyW7_1(.din(w_dff_B_cK3e9Z3T8_1),.dout(w_dff_B_BUnj0QyW7_1),.clk(gclk));
	jdff dff_B_0f3GhMrc8_1(.din(w_dff_B_BUnj0QyW7_1),.dout(w_dff_B_0f3GhMrc8_1),.clk(gclk));
	jdff dff_B_agPU4M1E7_1(.din(w_dff_B_0f3GhMrc8_1),.dout(w_dff_B_agPU4M1E7_1),.clk(gclk));
	jdff dff_B_yxqbIcDq2_1(.din(w_dff_B_agPU4M1E7_1),.dout(w_dff_B_yxqbIcDq2_1),.clk(gclk));
	jdff dff_B_RmIz27ih2_1(.din(w_dff_B_yxqbIcDq2_1),.dout(w_dff_B_RmIz27ih2_1),.clk(gclk));
	jdff dff_B_TCubaHiW8_1(.din(w_dff_B_RmIz27ih2_1),.dout(w_dff_B_TCubaHiW8_1),.clk(gclk));
	jdff dff_B_Crsi5cq54_1(.din(w_dff_B_TCubaHiW8_1),.dout(w_dff_B_Crsi5cq54_1),.clk(gclk));
	jdff dff_B_G5W7pFqL9_1(.din(w_dff_B_Crsi5cq54_1),.dout(w_dff_B_G5W7pFqL9_1),.clk(gclk));
	jdff dff_A_xVCbd2lf1_0(.dout(w_G159gat_1[0]),.din(w_dff_A_xVCbd2lf1_0),.clk(gclk));
	jdff dff_A_HC0x09Pj9_0(.dout(w_dff_A_xVCbd2lf1_0),.din(w_dff_A_HC0x09Pj9_0),.clk(gclk));
	jdff dff_A_kR5YIjbe0_0(.dout(w_dff_A_HC0x09Pj9_0),.din(w_dff_A_kR5YIjbe0_0),.clk(gclk));
	jdff dff_A_ATAq18RA7_0(.dout(w_dff_A_kR5YIjbe0_0),.din(w_dff_A_ATAq18RA7_0),.clk(gclk));
	jdff dff_A_568KjyB94_0(.dout(w_dff_A_ATAq18RA7_0),.din(w_dff_A_568KjyB94_0),.clk(gclk));
	jdff dff_A_DqioWgSz5_0(.dout(w_dff_A_568KjyB94_0),.din(w_dff_A_DqioWgSz5_0),.clk(gclk));
	jdff dff_A_es7kT23C2_0(.dout(w_dff_A_DqioWgSz5_0),.din(w_dff_A_es7kT23C2_0),.clk(gclk));
	jdff dff_A_1BKxyyK10_0(.dout(w_dff_A_es7kT23C2_0),.din(w_dff_A_1BKxyyK10_0),.clk(gclk));
	jdff dff_A_O8Vklup97_0(.dout(w_dff_A_1BKxyyK10_0),.din(w_dff_A_O8Vklup97_0),.clk(gclk));
	jdff dff_A_DFUfRgTK0_1(.dout(w_G159gat_1[1]),.din(w_dff_A_DFUfRgTK0_1),.clk(gclk));
	jdff dff_A_t2TQ3gLM1_1(.dout(w_dff_A_DFUfRgTK0_1),.din(w_dff_A_t2TQ3gLM1_1),.clk(gclk));
	jdff dff_A_ULzcb9f16_1(.dout(w_dff_A_t2TQ3gLM1_1),.din(w_dff_A_ULzcb9f16_1),.clk(gclk));
	jdff dff_A_Exgb0kkr0_1(.dout(w_dff_A_ULzcb9f16_1),.din(w_dff_A_Exgb0kkr0_1),.clk(gclk));
	jdff dff_A_LLlRukt87_1(.dout(w_dff_A_Exgb0kkr0_1),.din(w_dff_A_LLlRukt87_1),.clk(gclk));
	jdff dff_A_gnkWmC5J5_1(.dout(w_dff_A_LLlRukt87_1),.din(w_dff_A_gnkWmC5J5_1),.clk(gclk));
	jdff dff_A_Cz0Cu0aV2_1(.dout(w_dff_A_gnkWmC5J5_1),.din(w_dff_A_Cz0Cu0aV2_1),.clk(gclk));
	jdff dff_A_jFhtMyKy5_1(.dout(w_dff_A_Cz0Cu0aV2_1),.din(w_dff_A_jFhtMyKy5_1),.clk(gclk));
	jdff dff_A_5rMxZFOJ6_1(.dout(w_dff_A_jFhtMyKy5_1),.din(w_dff_A_5rMxZFOJ6_1),.clk(gclk));
	jdff dff_B_GPhE9peD1_1(.din(n358),.dout(w_dff_B_GPhE9peD1_1),.clk(gclk));
	jdff dff_B_dDZMWDgu2_1(.din(w_dff_B_GPhE9peD1_1),.dout(w_dff_B_dDZMWDgu2_1),.clk(gclk));
	jdff dff_B_FN5MSQz78_0(.din(n371),.dout(w_dff_B_FN5MSQz78_0),.clk(gclk));
	jdff dff_B_JOYH0Xz12_0(.din(w_dff_B_FN5MSQz78_0),.dout(w_dff_B_JOYH0Xz12_0),.clk(gclk));
	jdff dff_B_FuOOvbjw1_0(.din(w_dff_B_JOYH0Xz12_0),.dout(w_dff_B_FuOOvbjw1_0),.clk(gclk));
	jdff dff_B_nhK3TEkx1_0(.din(w_dff_B_FuOOvbjw1_0),.dout(w_dff_B_nhK3TEkx1_0),.clk(gclk));
	jdff dff_B_YJfwExrU1_0(.din(w_dff_B_nhK3TEkx1_0),.dout(w_dff_B_YJfwExrU1_0),.clk(gclk));
	jdff dff_B_1pV9Y5bC2_0(.din(w_dff_B_YJfwExrU1_0),.dout(w_dff_B_1pV9Y5bC2_0),.clk(gclk));
	jdff dff_B_oM4e1fGD4_0(.din(w_dff_B_1pV9Y5bC2_0),.dout(w_dff_B_oM4e1fGD4_0),.clk(gclk));
	jdff dff_B_oYpqn9Si8_0(.din(w_dff_B_oM4e1fGD4_0),.dout(w_dff_B_oYpqn9Si8_0),.clk(gclk));
	jdff dff_B_KIQzMffs8_0(.din(w_dff_B_oYpqn9Si8_0),.dout(w_dff_B_KIQzMffs8_0),.clk(gclk));
	jdff dff_B_45YLzm8C4_0(.din(n369),.dout(w_dff_B_45YLzm8C4_0),.clk(gclk));
	jdff dff_B_t1lwdvkp9_0(.din(w_dff_B_45YLzm8C4_0),.dout(w_dff_B_t1lwdvkp9_0),.clk(gclk));
	jdff dff_B_mCEZtpVI8_0(.din(w_dff_B_t1lwdvkp9_0),.dout(w_dff_B_mCEZtpVI8_0),.clk(gclk));
	jdff dff_B_3ejL3m9E0_0(.din(w_dff_B_mCEZtpVI8_0),.dout(w_dff_B_3ejL3m9E0_0),.clk(gclk));
	jdff dff_B_gpVBdfsV2_1(.din(n367),.dout(w_dff_B_gpVBdfsV2_1),.clk(gclk));
	jdff dff_B_3nLihxdL9_1(.din(w_dff_B_gpVBdfsV2_1),.dout(w_dff_B_3nLihxdL9_1),.clk(gclk));
	jdff dff_B_1r9sycvd2_1(.din(w_dff_B_3nLihxdL9_1),.dout(w_dff_B_1r9sycvd2_1),.clk(gclk));
	jdff dff_B_C2QS22wE8_1(.din(w_dff_B_1r9sycvd2_1),.dout(w_dff_B_C2QS22wE8_1),.clk(gclk));
	jdff dff_A_59789IK71_0(.dout(w_G246gat_2[0]),.din(w_dff_A_59789IK71_0),.clk(gclk));
	jdff dff_A_vxoLuX1Q7_0(.dout(w_dff_A_59789IK71_0),.din(w_dff_A_vxoLuX1Q7_0),.clk(gclk));
	jdff dff_A_JhfWkjJ38_0(.dout(w_dff_A_vxoLuX1Q7_0),.din(w_dff_A_JhfWkjJ38_0),.clk(gclk));
	jdff dff_A_7VJLBtPY3_0(.dout(w_dff_A_JhfWkjJ38_0),.din(w_dff_A_7VJLBtPY3_0),.clk(gclk));
	jdff dff_A_sGzLHVee3_0(.dout(w_dff_A_7VJLBtPY3_0),.din(w_dff_A_sGzLHVee3_0),.clk(gclk));
	jdff dff_A_g8THXuPB6_0(.dout(w_dff_A_sGzLHVee3_0),.din(w_dff_A_g8THXuPB6_0),.clk(gclk));
	jdff dff_A_tNk60cMu8_0(.dout(w_dff_A_g8THXuPB6_0),.din(w_dff_A_tNk60cMu8_0),.clk(gclk));
	jdff dff_A_h4gHO2iu9_0(.dout(w_dff_A_tNk60cMu8_0),.din(w_dff_A_h4gHO2iu9_0),.clk(gclk));
	jdff dff_A_eThL9HM11_0(.dout(w_G237gat_2[0]),.din(w_dff_A_eThL9HM11_0),.clk(gclk));
	jdff dff_A_gDlbk4Ia6_0(.dout(w_dff_A_eThL9HM11_0),.din(w_dff_A_gDlbk4Ia6_0),.clk(gclk));
	jdff dff_A_ch7dmcIp8_0(.dout(w_dff_A_gDlbk4Ia6_0),.din(w_dff_A_ch7dmcIp8_0),.clk(gclk));
	jdff dff_A_2UGetOFz2_0(.dout(w_dff_A_ch7dmcIp8_0),.din(w_dff_A_2UGetOFz2_0),.clk(gclk));
	jdff dff_A_u2asBRF63_0(.dout(w_dff_A_2UGetOFz2_0),.din(w_dff_A_u2asBRF63_0),.clk(gclk));
	jdff dff_A_MSP3JsP91_0(.dout(w_dff_A_u2asBRF63_0),.din(w_dff_A_MSP3JsP91_0),.clk(gclk));
	jdff dff_A_Fb5zEkqL0_0(.dout(w_dff_A_MSP3JsP91_0),.din(w_dff_A_Fb5zEkqL0_0),.clk(gclk));
	jdff dff_A_zu6g0c7R2_0(.dout(w_dff_A_Fb5zEkqL0_0),.din(w_dff_A_zu6g0c7R2_0),.clk(gclk));
	jdff dff_A_1LorvZwg6_0(.dout(w_dff_A_zu6g0c7R2_0),.din(w_dff_A_1LorvZwg6_0),.clk(gclk));
	jdff dff_A_Gs7sp7nX6_0(.dout(w_dff_A_1LorvZwg6_0),.din(w_dff_A_Gs7sp7nX6_0),.clk(gclk));
	jdff dff_A_lBzLUwpW9_0(.dout(w_G228gat_2[0]),.din(w_dff_A_lBzLUwpW9_0),.clk(gclk));
	jdff dff_A_G51sbAmz5_0(.dout(w_dff_A_lBzLUwpW9_0),.din(w_dff_A_G51sbAmz5_0),.clk(gclk));
	jdff dff_A_nDEMpseI7_0(.dout(w_dff_A_G51sbAmz5_0),.din(w_dff_A_nDEMpseI7_0),.clk(gclk));
	jdff dff_A_BUhkNS0b3_0(.dout(w_dff_A_nDEMpseI7_0),.din(w_dff_A_BUhkNS0b3_0),.clk(gclk));
	jdff dff_A_tIFLXirb2_0(.dout(w_dff_A_BUhkNS0b3_0),.din(w_dff_A_tIFLXirb2_0),.clk(gclk));
	jdff dff_A_Oe9a0CGt2_0(.dout(w_dff_A_tIFLXirb2_0),.din(w_dff_A_Oe9a0CGt2_0),.clk(gclk));
	jdff dff_A_REtwFYfb2_0(.dout(w_dff_A_Oe9a0CGt2_0),.din(w_dff_A_REtwFYfb2_0),.clk(gclk));
	jdff dff_A_XYTdUqX19_0(.dout(w_dff_A_REtwFYfb2_0),.din(w_dff_A_XYTdUqX19_0),.clk(gclk));
	jdff dff_A_W48Xm7nX1_0(.dout(w_dff_A_XYTdUqX19_0),.din(w_dff_A_W48Xm7nX1_0),.clk(gclk));
	jdff dff_A_XHTaupih4_0(.dout(w_dff_A_W48Xm7nX1_0),.din(w_dff_A_XHTaupih4_0),.clk(gclk));
	jdff dff_B_n2gwc0Wj5_1(.din(n356),.dout(w_dff_B_n2gwc0Wj5_1),.clk(gclk));
	jdff dff_B_b8rYDj6P0_1(.din(w_dff_B_n2gwc0Wj5_1),.dout(w_dff_B_b8rYDj6P0_1),.clk(gclk));
	jdff dff_B_3TSyV1bV3_1(.din(w_dff_B_b8rYDj6P0_1),.dout(w_dff_B_3TSyV1bV3_1),.clk(gclk));
	jdff dff_B_GuAntEwq1_1(.din(w_dff_B_3TSyV1bV3_1),.dout(w_dff_B_GuAntEwq1_1),.clk(gclk));
	jdff dff_B_j7SlwgB99_1(.din(w_dff_B_GuAntEwq1_1),.dout(w_dff_B_j7SlwgB99_1),.clk(gclk));
	jdff dff_B_kh9VxO0k5_1(.din(w_dff_B_j7SlwgB99_1),.dout(w_dff_B_kh9VxO0k5_1),.clk(gclk));
	jdff dff_B_ndfcPuaT1_1(.din(w_dff_B_kh9VxO0k5_1),.dout(w_dff_B_ndfcPuaT1_1),.clk(gclk));
	jdff dff_B_bYpKujEX4_1(.din(w_dff_B_ndfcPuaT1_1),.dout(w_dff_B_bYpKujEX4_1),.clk(gclk));
	jdff dff_A_bJ3daH7s7_0(.dout(w_G219gat_2[0]),.din(w_dff_A_bJ3daH7s7_0),.clk(gclk));
	jdff dff_A_FFFIshbQ3_0(.dout(w_dff_A_bJ3daH7s7_0),.din(w_dff_A_FFFIshbQ3_0),.clk(gclk));
	jdff dff_A_qtemNoQF6_0(.dout(w_dff_A_FFFIshbQ3_0),.din(w_dff_A_qtemNoQF6_0),.clk(gclk));
	jdff dff_A_GArnw1Hh2_0(.dout(w_dff_A_qtemNoQF6_0),.din(w_dff_A_GArnw1Hh2_0),.clk(gclk));
	jdff dff_A_veE51J5r6_0(.dout(w_dff_A_GArnw1Hh2_0),.din(w_dff_A_veE51J5r6_0),.clk(gclk));
	jdff dff_A_sidqFTyr6_1(.dout(w_G219gat_2[1]),.din(w_dff_A_sidqFTyr6_1),.clk(gclk));
	jdff dff_A_q8r5PICu7_1(.dout(w_dff_A_sidqFTyr6_1),.din(w_dff_A_q8r5PICu7_1),.clk(gclk));
	jdff dff_A_MoxOgXXi2_1(.dout(w_dff_A_q8r5PICu7_1),.din(w_dff_A_MoxOgXXi2_1),.clk(gclk));
	jdff dff_A_5ThYq8HY6_1(.dout(w_dff_A_MoxOgXXi2_1),.din(w_dff_A_5ThYq8HY6_1),.clk(gclk));
	jdff dff_A_HdP8i38R0_1(.dout(w_dff_A_5ThYq8HY6_1),.din(w_dff_A_HdP8i38R0_1),.clk(gclk));
	jdff dff_A_tSxS8ex92_0(.dout(w_n355_0[0]),.din(w_dff_A_tSxS8ex92_0),.clk(gclk));
	jdff dff_A_9HdxmpXx7_0(.dout(w_dff_A_tSxS8ex92_0),.din(w_dff_A_9HdxmpXx7_0),.clk(gclk));
	jdff dff_A_k2Q75X6R6_0(.dout(w_dff_A_9HdxmpXx7_0),.din(w_dff_A_k2Q75X6R6_0),.clk(gclk));
	jdff dff_A_7iYUx3bS4_0(.dout(w_dff_A_k2Q75X6R6_0),.din(w_dff_A_7iYUx3bS4_0),.clk(gclk));
	jdff dff_A_c2ulKy9Q7_0(.dout(w_dff_A_7iYUx3bS4_0),.din(w_dff_A_c2ulKy9Q7_0),.clk(gclk));
	jdff dff_A_zxLR4eFD5_0(.dout(w_dff_A_c2ulKy9Q7_0),.din(w_dff_A_zxLR4eFD5_0),.clk(gclk));
	jdff dff_A_MuNfmDZT5_0(.dout(w_dff_A_zxLR4eFD5_0),.din(w_dff_A_MuNfmDZT5_0),.clk(gclk));
	jdff dff_A_LCf2uBmQ9_0(.dout(w_dff_A_MuNfmDZT5_0),.din(w_dff_A_LCf2uBmQ9_0),.clk(gclk));
	jdff dff_A_9Z1wnDuS3_0(.dout(w_dff_A_LCf2uBmQ9_0),.din(w_dff_A_9Z1wnDuS3_0),.clk(gclk));
	jdff dff_A_WTmwzHhH3_0(.dout(w_dff_A_9Z1wnDuS3_0),.din(w_dff_A_WTmwzHhH3_0),.clk(gclk));
	jdff dff_B_70CWGrjI8_1(.din(n383),.dout(w_dff_B_70CWGrjI8_1),.clk(gclk));
	jdff dff_B_K4KwPQzj4_1(.din(w_dff_B_70CWGrjI8_1),.dout(w_dff_B_K4KwPQzj4_1),.clk(gclk));
	jdff dff_B_elh2Lk664_1(.din(w_dff_B_K4KwPQzj4_1),.dout(w_dff_B_elh2Lk664_1),.clk(gclk));
	jdff dff_B_QJXJPvJC7_1(.din(w_dff_B_elh2Lk664_1),.dout(w_dff_B_QJXJPvJC7_1),.clk(gclk));
	jdff dff_B_JcgMogmf8_1(.din(w_dff_B_QJXJPvJC7_1),.dout(w_dff_B_JcgMogmf8_1),.clk(gclk));
	jdff dff_B_TAxAW1TE0_1(.din(w_dff_B_JcgMogmf8_1),.dout(w_dff_B_TAxAW1TE0_1),.clk(gclk));
	jdff dff_B_p6qSeAFm5_1(.din(w_dff_B_TAxAW1TE0_1),.dout(w_dff_B_p6qSeAFm5_1),.clk(gclk));
	jdff dff_B_UBdkgCNo1_1(.din(w_dff_B_p6qSeAFm5_1),.dout(w_dff_B_UBdkgCNo1_1),.clk(gclk));
	jdff dff_B_3TIzWT7q7_1(.din(w_dff_B_UBdkgCNo1_1),.dout(w_dff_B_3TIzWT7q7_1),.clk(gclk));
	jdff dff_B_jllHzEmu8_1(.din(w_dff_B_3TIzWT7q7_1),.dout(w_dff_B_jllHzEmu8_1),.clk(gclk));
	jdff dff_B_dZ8btkFc7_1(.din(w_dff_B_jllHzEmu8_1),.dout(w_dff_B_dZ8btkFc7_1),.clk(gclk));
	jdff dff_B_ZJiliUBo6_1(.din(w_dff_B_dZ8btkFc7_1),.dout(w_dff_B_ZJiliUBo6_1),.clk(gclk));
	jdff dff_B_ijMSrt5x0_1(.din(w_dff_B_ZJiliUBo6_1),.dout(w_dff_B_ijMSrt5x0_1),.clk(gclk));
	jdff dff_B_mfXSlU7j1_1(.din(n384),.dout(w_dff_B_mfXSlU7j1_1),.clk(gclk));
	jdff dff_B_gjEntSGG0_0(.din(n396),.dout(w_dff_B_gjEntSGG0_0),.clk(gclk));
	jdff dff_B_TtY3cPI91_0(.din(w_dff_B_gjEntSGG0_0),.dout(w_dff_B_TtY3cPI91_0),.clk(gclk));
	jdff dff_B_eeKoyiNY8_0(.din(w_dff_B_TtY3cPI91_0),.dout(w_dff_B_eeKoyiNY8_0),.clk(gclk));
	jdff dff_B_0UUyqVNO3_0(.din(w_dff_B_eeKoyiNY8_0),.dout(w_dff_B_0UUyqVNO3_0),.clk(gclk));
	jdff dff_B_nS0kYOT68_0(.din(w_dff_B_0UUyqVNO3_0),.dout(w_dff_B_nS0kYOT68_0),.clk(gclk));
	jdff dff_B_LavBUcDn8_0(.din(w_dff_B_nS0kYOT68_0),.dout(w_dff_B_LavBUcDn8_0),.clk(gclk));
	jdff dff_B_x7scORUO7_0(.din(w_dff_B_LavBUcDn8_0),.dout(w_dff_B_x7scORUO7_0),.clk(gclk));
	jdff dff_B_bnIP7UBA7_0(.din(w_dff_B_x7scORUO7_0),.dout(w_dff_B_bnIP7UBA7_0),.clk(gclk));
	jdff dff_B_dEFVNWWr4_0(.din(w_dff_B_bnIP7UBA7_0),.dout(w_dff_B_dEFVNWWr4_0),.clk(gclk));
	jdff dff_B_E5dNJnVk6_0(.din(w_dff_B_dEFVNWWr4_0),.dout(w_dff_B_E5dNJnVk6_0),.clk(gclk));
	jdff dff_B_ekhsX9qf0_0(.din(w_dff_B_E5dNJnVk6_0),.dout(w_dff_B_ekhsX9qf0_0),.clk(gclk));
	jdff dff_B_zyDzmDZh4_0(.din(w_dff_B_ekhsX9qf0_0),.dout(w_dff_B_zyDzmDZh4_0),.clk(gclk));
	jdff dff_B_1H8axePV9_0(.din(w_dff_B_zyDzmDZh4_0),.dout(w_dff_B_1H8axePV9_0),.clk(gclk));
	jdff dff_B_fp7LMI6Y1_1(.din(n385),.dout(w_dff_B_fp7LMI6Y1_1),.clk(gclk));
	jdff dff_B_2NjnirCd9_1(.din(w_dff_B_fp7LMI6Y1_1),.dout(w_dff_B_2NjnirCd9_1),.clk(gclk));
	jdff dff_B_ecR09ZOB4_1(.din(w_dff_B_2NjnirCd9_1),.dout(w_dff_B_ecR09ZOB4_1),.clk(gclk));
	jdff dff_B_bRMTJVsK4_1(.din(w_dff_B_ecR09ZOB4_1),.dout(w_dff_B_bRMTJVsK4_1),.clk(gclk));
	jdff dff_B_y3lGjh756_1(.din(w_dff_B_bRMTJVsK4_1),.dout(w_dff_B_y3lGjh756_1),.clk(gclk));
	jdff dff_B_jU7pNuAJ5_1(.din(w_dff_B_y3lGjh756_1),.dout(w_dff_B_jU7pNuAJ5_1),.clk(gclk));
	jdff dff_B_WFd4YglH5_1(.din(w_dff_B_jU7pNuAJ5_1),.dout(w_dff_B_WFd4YglH5_1),.clk(gclk));
	jdff dff_B_Di7pQTo20_1(.din(w_dff_B_WFd4YglH5_1),.dout(w_dff_B_Di7pQTo20_1),.clk(gclk));
	jdff dff_B_OBxQareG3_1(.din(w_dff_B_Di7pQTo20_1),.dout(w_dff_B_OBxQareG3_1),.clk(gclk));
	jdff dff_B_dcIdBJQX2_1(.din(w_dff_B_OBxQareG3_1),.dout(w_dff_B_dcIdBJQX2_1),.clk(gclk));
	jdff dff_B_yueMlWGZ3_1(.din(w_dff_B_dcIdBJQX2_1),.dout(w_dff_B_yueMlWGZ3_1),.clk(gclk));
	jdff dff_B_YkK2LiLL9_1(.din(w_dff_B_yueMlWGZ3_1),.dout(w_dff_B_YkK2LiLL9_1),.clk(gclk));
	jdff dff_B_aHvNFreD1_1(.din(n386),.dout(w_dff_B_aHvNFreD1_1),.clk(gclk));
	jdff dff_B_CSXGgycY4_1(.din(w_dff_B_aHvNFreD1_1),.dout(w_dff_B_CSXGgycY4_1),.clk(gclk));
	jdff dff_B_Up8wcUm81_1(.din(w_dff_B_CSXGgycY4_1),.dout(w_dff_B_Up8wcUm81_1),.clk(gclk));
	jdff dff_B_xRKcFhbq1_1(.din(w_dff_B_Up8wcUm81_1),.dout(w_dff_B_xRKcFhbq1_1),.clk(gclk));
	jdff dff_B_jubtWu7l6_1(.din(w_dff_B_xRKcFhbq1_1),.dout(w_dff_B_jubtWu7l6_1),.clk(gclk));
	jdff dff_B_kSzUQxZW4_1(.din(w_dff_B_jubtWu7l6_1),.dout(w_dff_B_kSzUQxZW4_1),.clk(gclk));
	jdff dff_B_O0Co4cgu7_1(.din(w_dff_B_kSzUQxZW4_1),.dout(w_dff_B_O0Co4cgu7_1),.clk(gclk));
	jdff dff_B_N6UCPSSF5_1(.din(w_dff_B_O0Co4cgu7_1),.dout(w_dff_B_N6UCPSSF5_1),.clk(gclk));
	jdff dff_B_aKNoyOfg5_1(.din(w_dff_B_N6UCPSSF5_1),.dout(w_dff_B_aKNoyOfg5_1),.clk(gclk));
	jdff dff_B_eDgVJC478_1(.din(w_dff_B_aKNoyOfg5_1),.dout(w_dff_B_eDgVJC478_1),.clk(gclk));
	jdff dff_B_ORnpkLBA5_1(.din(w_dff_B_eDgVJC478_1),.dout(w_dff_B_ORnpkLBA5_1),.clk(gclk));
	jdff dff_A_SPd4hQoH9_1(.dout(w_n321_0[1]),.din(w_dff_A_SPd4hQoH9_1),.clk(gclk));
	jdff dff_A_alXJXg7B6_1(.dout(w_dff_A_SPd4hQoH9_1),.din(w_dff_A_alXJXg7B6_1),.clk(gclk));
	jdff dff_A_dHrcjvzZ0_1(.dout(w_dff_A_alXJXg7B6_1),.din(w_dff_A_dHrcjvzZ0_1),.clk(gclk));
	jdff dff_A_5zOnVWgp5_1(.dout(w_dff_A_dHrcjvzZ0_1),.din(w_dff_A_5zOnVWgp5_1),.clk(gclk));
	jdff dff_A_WtDQ0C6I6_1(.dout(w_dff_A_5zOnVWgp5_1),.din(w_dff_A_WtDQ0C6I6_1),.clk(gclk));
	jdff dff_A_MN2wCX0R6_1(.dout(w_dff_A_WtDQ0C6I6_1),.din(w_dff_A_MN2wCX0R6_1),.clk(gclk));
	jdff dff_A_kiWtPUaK0_1(.dout(w_dff_A_MN2wCX0R6_1),.din(w_dff_A_kiWtPUaK0_1),.clk(gclk));
	jdff dff_A_kDsYcmTD4_1(.dout(w_dff_A_kiWtPUaK0_1),.din(w_dff_A_kDsYcmTD4_1),.clk(gclk));
	jdff dff_A_S0lkKPoz1_1(.dout(w_dff_A_kDsYcmTD4_1),.din(w_dff_A_S0lkKPoz1_1),.clk(gclk));
	jdff dff_A_k27b6J7i0_1(.dout(w_dff_A_S0lkKPoz1_1),.din(w_dff_A_k27b6J7i0_1),.clk(gclk));
	jdff dff_A_xpGovbfh8_1(.dout(w_dff_A_k27b6J7i0_1),.din(w_dff_A_xpGovbfh8_1),.clk(gclk));
	jdff dff_A_uy3vY4jq6_1(.dout(w_dff_A_xpGovbfh8_1),.din(w_dff_A_uy3vY4jq6_1),.clk(gclk));
	jdff dff_A_i3iRedDT1_1(.dout(w_n320_0[1]),.din(w_dff_A_i3iRedDT1_1),.clk(gclk));
	jdff dff_A_Vtb3yNv80_1(.dout(w_dff_A_i3iRedDT1_1),.din(w_dff_A_Vtb3yNv80_1),.clk(gclk));
	jdff dff_A_NB21JOM31_1(.dout(w_dff_A_Vtb3yNv80_1),.din(w_dff_A_NB21JOM31_1),.clk(gclk));
	jdff dff_A_8FnFl0Ka1_1(.dout(w_dff_A_NB21JOM31_1),.din(w_dff_A_8FnFl0Ka1_1),.clk(gclk));
	jdff dff_A_Bfh220527_1(.dout(w_dff_A_8FnFl0Ka1_1),.din(w_dff_A_Bfh220527_1),.clk(gclk));
	jdff dff_A_Bd3YpNBu6_1(.dout(w_dff_A_Bfh220527_1),.din(w_dff_A_Bd3YpNBu6_1),.clk(gclk));
	jdff dff_A_L2jm9TSj8_1(.dout(w_dff_A_Bd3YpNBu6_1),.din(w_dff_A_L2jm9TSj8_1),.clk(gclk));
	jdff dff_A_RzrELDkc0_1(.dout(w_dff_A_L2jm9TSj8_1),.din(w_dff_A_RzrELDkc0_1),.clk(gclk));
	jdff dff_A_5DNRdYme2_1(.dout(w_dff_A_RzrELDkc0_1),.din(w_dff_A_5DNRdYme2_1),.clk(gclk));
	jdff dff_A_rwqahejY1_1(.dout(w_dff_A_5DNRdYme2_1),.din(w_dff_A_rwqahejY1_1),.clk(gclk));
	jdff dff_A_Wm0Jxyom7_1(.dout(w_dff_A_rwqahejY1_1),.din(w_dff_A_Wm0Jxyom7_1),.clk(gclk));
	jdff dff_A_P7w0ZNjN8_1(.dout(w_dff_A_Wm0Jxyom7_1),.din(w_dff_A_P7w0ZNjN8_1),.clk(gclk));
	jdff dff_A_pcKRiF3c5_1(.dout(w_dff_A_P7w0ZNjN8_1),.din(w_dff_A_pcKRiF3c5_1),.clk(gclk));
	jdff dff_A_f0Tnz2Rf4_0(.dout(w_G165gat_1[0]),.din(w_dff_A_f0Tnz2Rf4_0),.clk(gclk));
	jdff dff_A_hYU0cSRm4_0(.dout(w_dff_A_f0Tnz2Rf4_0),.din(w_dff_A_hYU0cSRm4_0),.clk(gclk));
	jdff dff_A_IKgKATdn5_0(.dout(w_dff_A_hYU0cSRm4_0),.din(w_dff_A_IKgKATdn5_0),.clk(gclk));
	jdff dff_A_0392metA6_0(.dout(w_dff_A_IKgKATdn5_0),.din(w_dff_A_0392metA6_0),.clk(gclk));
	jdff dff_A_hfHBCBrd4_0(.dout(w_dff_A_0392metA6_0),.din(w_dff_A_hfHBCBrd4_0),.clk(gclk));
	jdff dff_A_mwI5hC6T4_0(.dout(w_dff_A_hfHBCBrd4_0),.din(w_dff_A_mwI5hC6T4_0),.clk(gclk));
	jdff dff_A_BjfqaBXx3_0(.dout(w_dff_A_mwI5hC6T4_0),.din(w_dff_A_BjfqaBXx3_0),.clk(gclk));
	jdff dff_A_e8Ofl2I68_0(.dout(w_dff_A_BjfqaBXx3_0),.din(w_dff_A_e8Ofl2I68_0),.clk(gclk));
	jdff dff_A_C391u25s3_1(.dout(w_G165gat_1[1]),.din(w_dff_A_C391u25s3_1),.clk(gclk));
	jdff dff_A_zPqbXuor2_1(.dout(w_dff_A_C391u25s3_1),.din(w_dff_A_zPqbXuor2_1),.clk(gclk));
	jdff dff_A_cx3u6k8U7_1(.dout(w_dff_A_zPqbXuor2_1),.din(w_dff_A_cx3u6k8U7_1),.clk(gclk));
	jdff dff_A_EZKn2qb88_1(.dout(w_dff_A_cx3u6k8U7_1),.din(w_dff_A_EZKn2qb88_1),.clk(gclk));
	jdff dff_A_Rm1vi7Dm2_1(.dout(w_dff_A_EZKn2qb88_1),.din(w_dff_A_Rm1vi7Dm2_1),.clk(gclk));
	jdff dff_A_T6MFeb4P1_1(.dout(w_dff_A_Rm1vi7Dm2_1),.din(w_dff_A_T6MFeb4P1_1),.clk(gclk));
	jdff dff_A_Ubtbp1NT0_1(.dout(w_dff_A_T6MFeb4P1_1),.din(w_dff_A_Ubtbp1NT0_1),.clk(gclk));
	jdff dff_A_gCsMnsrE5_1(.dout(w_dff_A_Ubtbp1NT0_1),.din(w_dff_A_gCsMnsrE5_1),.clk(gclk));
	jdff dff_B_TnSxArNL8_1(.din(n376),.dout(w_dff_B_TnSxArNL8_1),.clk(gclk));
	jdff dff_B_KipvtkXk5_0(.din(n381),.dout(w_dff_B_KipvtkXk5_0),.clk(gclk));
	jdff dff_B_dhwGUi4C4_0(.din(w_dff_B_KipvtkXk5_0),.dout(w_dff_B_dhwGUi4C4_0),.clk(gclk));
	jdff dff_B_MHrCsJvJ9_0(.din(n379),.dout(w_dff_B_MHrCsJvJ9_0),.clk(gclk));
	jdff dff_B_CpbJkFt88_0(.din(w_dff_B_MHrCsJvJ9_0),.dout(w_dff_B_CpbJkFt88_0),.clk(gclk));
	jdff dff_B_HtzshIPQ6_0(.din(w_dff_B_CpbJkFt88_0),.dout(w_dff_B_HtzshIPQ6_0),.clk(gclk));
	jdff dff_B_Its1ghR50_0(.din(w_dff_B_HtzshIPQ6_0),.dout(w_dff_B_Its1ghR50_0),.clk(gclk));
	jdff dff_B_qBnUhGcF5_0(.din(w_dff_B_Its1ghR50_0),.dout(w_dff_B_qBnUhGcF5_0),.clk(gclk));
	jdff dff_B_7sJIehnG8_0(.din(w_dff_B_qBnUhGcF5_0),.dout(w_dff_B_7sJIehnG8_0),.clk(gclk));
	jdff dff_B_3ohoTttX1_0(.din(w_dff_B_7sJIehnG8_0),.dout(w_dff_B_3ohoTttX1_0),.clk(gclk));
	jdff dff_B_BYWnBMy53_0(.din(w_dff_B_3ohoTttX1_0),.dout(w_dff_B_BYWnBMy53_0),.clk(gclk));
	jdff dff_B_VrBGeUMi8_0(.din(w_dff_B_BYWnBMy53_0),.dout(w_dff_B_VrBGeUMi8_0),.clk(gclk));
	jdff dff_B_bwf0huTv8_0(.din(w_dff_B_VrBGeUMi8_0),.dout(w_dff_B_bwf0huTv8_0),.clk(gclk));
	jdff dff_A_7ATrk8lA0_1(.dout(w_n377_0[1]),.din(w_dff_A_7ATrk8lA0_1),.clk(gclk));
	jdff dff_A_fI0k704R3_1(.dout(w_dff_A_7ATrk8lA0_1),.din(w_dff_A_fI0k704R3_1),.clk(gclk));
	jdff dff_A_FTX2Vn1G9_1(.dout(w_dff_A_fI0k704R3_1),.din(w_dff_A_FTX2Vn1G9_1),.clk(gclk));
	jdff dff_A_oTX2lA851_1(.dout(w_dff_A_FTX2Vn1G9_1),.din(w_dff_A_oTX2lA851_1),.clk(gclk));
	jdff dff_A_6elblald0_1(.dout(w_dff_A_oTX2lA851_1),.din(w_dff_A_6elblald0_1),.clk(gclk));
	jdff dff_A_wOf0Vs3J2_1(.dout(w_dff_A_6elblald0_1),.din(w_dff_A_wOf0Vs3J2_1),.clk(gclk));
	jdff dff_A_rEdaWlZD6_1(.dout(w_dff_A_wOf0Vs3J2_1),.din(w_dff_A_rEdaWlZD6_1),.clk(gclk));
	jdff dff_A_wpFhUrYf7_1(.dout(w_dff_A_rEdaWlZD6_1),.din(w_dff_A_wpFhUrYf7_1),.clk(gclk));
	jdff dff_A_1zoxcUQz6_1(.dout(w_dff_A_wpFhUrYf7_1),.din(w_dff_A_1zoxcUQz6_1),.clk(gclk));
	jdff dff_A_5uR6ew4C1_1(.dout(w_dff_A_1zoxcUQz6_1),.din(w_dff_A_5uR6ew4C1_1),.clk(gclk));
	jdff dff_A_PzTRTfC43_1(.dout(w_dff_A_5uR6ew4C1_1),.din(w_dff_A_PzTRTfC43_1),.clk(gclk));
	jdff dff_A_QWIExkVG9_1(.dout(w_dff_A_PzTRTfC43_1),.din(w_dff_A_QWIExkVG9_1),.clk(gclk));
	jdff dff_A_xHEuLEKk9_1(.dout(w_dff_A_QWIExkVG9_1),.din(w_dff_A_xHEuLEKk9_1),.clk(gclk));
	jdff dff_A_L9BAJdW84_1(.dout(w_dff_A_xHEuLEKk9_1),.din(w_dff_A_L9BAJdW84_1),.clk(gclk));
	jdff dff_B_CLxBbHRk0_1(.din(n307),.dout(w_dff_B_CLxBbHRk0_1),.clk(gclk));
	jdff dff_B_mE57rEnW3_0(.din(n309),.dout(w_dff_B_mE57rEnW3_0),.clk(gclk));
	jdff dff_B_JyLV2Q8U5_0(.din(w_dff_B_mE57rEnW3_0),.dout(w_dff_B_JyLV2Q8U5_0),.clk(gclk));
	jdff dff_B_iqj695lP5_0(.din(w_dff_B_JyLV2Q8U5_0),.dout(w_dff_B_iqj695lP5_0),.clk(gclk));
	jdff dff_B_I7u5Bzyw3_0(.din(w_dff_B_iqj695lP5_0),.dout(w_dff_B_I7u5Bzyw3_0),.clk(gclk));
	jdff dff_B_hAr2lqVH2_0(.din(w_dff_B_I7u5Bzyw3_0),.dout(w_dff_B_hAr2lqVH2_0),.clk(gclk));
	jdff dff_B_gNuOt0Qh5_0(.din(w_dff_B_hAr2lqVH2_0),.dout(w_dff_B_gNuOt0Qh5_0),.clk(gclk));
	jdff dff_B_mf2zHNDT5_1(.din(n304),.dout(w_dff_B_mf2zHNDT5_1),.clk(gclk));
	jdff dff_A_RPvBiwtN1_1(.dout(w_G159gat_0[1]),.din(w_dff_A_RPvBiwtN1_1),.clk(gclk));
	jdff dff_A_AhNfZjqw4_1(.dout(w_dff_A_RPvBiwtN1_1),.din(w_dff_A_AhNfZjqw4_1),.clk(gclk));
	jdff dff_A_ii5jO80d8_1(.dout(w_dff_A_AhNfZjqw4_1),.din(w_dff_A_ii5jO80d8_1),.clk(gclk));
	jdff dff_A_FRKPHSb78_1(.dout(w_dff_A_ii5jO80d8_1),.din(w_dff_A_FRKPHSb78_1),.clk(gclk));
	jdff dff_A_xfzsnMIv6_1(.dout(w_dff_A_FRKPHSb78_1),.din(w_dff_A_xfzsnMIv6_1),.clk(gclk));
	jdff dff_A_BAHIDpAU2_1(.dout(w_dff_A_xfzsnMIv6_1),.din(w_dff_A_BAHIDpAU2_1),.clk(gclk));
	jdff dff_A_KrKVBosd4_1(.dout(w_dff_A_BAHIDpAU2_1),.din(w_dff_A_KrKVBosd4_1),.clk(gclk));
	jdff dff_A_mztmAX8J0_1(.dout(w_dff_A_KrKVBosd4_1),.din(w_dff_A_mztmAX8J0_1),.clk(gclk));
	jdff dff_A_Cdh1RHdS9_1(.dout(w_dff_A_mztmAX8J0_1),.din(w_dff_A_Cdh1RHdS9_1),.clk(gclk));
	jdff dff_A_Lq5lGMV70_2(.dout(w_G159gat_0[2]),.din(w_dff_A_Lq5lGMV70_2),.clk(gclk));
	jdff dff_A_mS6P4vMk2_2(.dout(w_dff_A_Lq5lGMV70_2),.din(w_dff_A_mS6P4vMk2_2),.clk(gclk));
	jdff dff_A_zjTxZgD94_2(.dout(w_dff_A_mS6P4vMk2_2),.din(w_dff_A_zjTxZgD94_2),.clk(gclk));
	jdff dff_A_D4q2zQEj8_2(.dout(w_dff_A_zjTxZgD94_2),.din(w_dff_A_D4q2zQEj8_2),.clk(gclk));
	jdff dff_A_OiQ2ftAf5_2(.dout(w_dff_A_D4q2zQEj8_2),.din(w_dff_A_OiQ2ftAf5_2),.clk(gclk));
	jdff dff_A_LA9QaM5A7_2(.dout(w_dff_A_OiQ2ftAf5_2),.din(w_dff_A_LA9QaM5A7_2),.clk(gclk));
	jdff dff_A_U6k3qrq82_2(.dout(w_dff_A_LA9QaM5A7_2),.din(w_dff_A_U6k3qrq82_2),.clk(gclk));
	jdff dff_A_l6nWrpZy7_2(.dout(w_dff_A_U6k3qrq82_2),.din(w_dff_A_l6nWrpZy7_2),.clk(gclk));
	jdff dff_A_WIZqdezD2_2(.dout(w_dff_A_l6nWrpZy7_2),.din(w_dff_A_WIZqdezD2_2),.clk(gclk));
	jdff dff_A_Gj1DOGlz4_2(.dout(w_dff_A_WIZqdezD2_2),.din(w_dff_A_Gj1DOGlz4_2),.clk(gclk));
	jdff dff_A_ooxJvQMe3_2(.dout(w_dff_A_Gj1DOGlz4_2),.din(w_dff_A_ooxJvQMe3_2),.clk(gclk));
	jdff dff_B_IxmWWaaA2_1(.din(n410),.dout(w_dff_B_IxmWWaaA2_1),.clk(gclk));
	jdff dff_B_6niYvNzb6_1(.din(w_dff_B_IxmWWaaA2_1),.dout(w_dff_B_6niYvNzb6_1),.clk(gclk));
	jdff dff_B_Kpy8p9277_1(.din(w_dff_B_6niYvNzb6_1),.dout(w_dff_B_Kpy8p9277_1),.clk(gclk));
	jdff dff_B_Fr1O2fo07_1(.din(w_dff_B_Kpy8p9277_1),.dout(w_dff_B_Fr1O2fo07_1),.clk(gclk));
	jdff dff_B_o3W47Yud8_1(.din(w_dff_B_Fr1O2fo07_1),.dout(w_dff_B_o3W47Yud8_1),.clk(gclk));
	jdff dff_B_ZQQbyMHB4_1(.din(w_dff_B_o3W47Yud8_1),.dout(w_dff_B_ZQQbyMHB4_1),.clk(gclk));
	jdff dff_B_SpTcmguP0_1(.din(w_dff_B_ZQQbyMHB4_1),.dout(w_dff_B_SpTcmguP0_1),.clk(gclk));
	jdff dff_B_ThYCInlC6_1(.din(w_dff_B_SpTcmguP0_1),.dout(w_dff_B_ThYCInlC6_1),.clk(gclk));
	jdff dff_B_TgmfaMBk4_1(.din(w_dff_B_ThYCInlC6_1),.dout(w_dff_B_TgmfaMBk4_1),.clk(gclk));
	jdff dff_B_8fNxos089_1(.din(w_dff_B_TgmfaMBk4_1),.dout(w_dff_B_8fNxos089_1),.clk(gclk));
	jdff dff_B_b77xlsdY5_1(.din(w_dff_B_8fNxos089_1),.dout(w_dff_B_b77xlsdY5_1),.clk(gclk));
	jdff dff_B_mebxrYF86_1(.din(n411),.dout(w_dff_B_mebxrYF86_1),.clk(gclk));
	jdff dff_B_5sJrgmDu4_0(.din(n412),.dout(w_dff_B_5sJrgmDu4_0),.clk(gclk));
	jdff dff_B_1pydwt8Y6_0(.din(w_dff_B_5sJrgmDu4_0),.dout(w_dff_B_1pydwt8Y6_0),.clk(gclk));
	jdff dff_B_BzkI7QOS5_0(.din(w_dff_B_1pydwt8Y6_0),.dout(w_dff_B_BzkI7QOS5_0),.clk(gclk));
	jdff dff_B_ObuiwlhG6_0(.din(w_dff_B_BzkI7QOS5_0),.dout(w_dff_B_ObuiwlhG6_0),.clk(gclk));
	jdff dff_B_uQgBBIEg4_0(.din(w_dff_B_ObuiwlhG6_0),.dout(w_dff_B_uQgBBIEg4_0),.clk(gclk));
	jdff dff_B_mi3XB9ba4_0(.din(w_dff_B_uQgBBIEg4_0),.dout(w_dff_B_mi3XB9ba4_0),.clk(gclk));
	jdff dff_B_P6C7vMeD7_0(.din(w_dff_B_mi3XB9ba4_0),.dout(w_dff_B_P6C7vMeD7_0),.clk(gclk));
	jdff dff_B_VKR7baJS2_0(.din(w_dff_B_P6C7vMeD7_0),.dout(w_dff_B_VKR7baJS2_0),.clk(gclk));
	jdff dff_B_D9jll0ar0_0(.din(w_dff_B_VKR7baJS2_0),.dout(w_dff_B_D9jll0ar0_0),.clk(gclk));
	jdff dff_B_6pyf0hvZ3_0(.din(w_dff_B_D9jll0ar0_0),.dout(w_dff_B_6pyf0hvZ3_0),.clk(gclk));
	jdff dff_B_2CBrTZA57_0(.din(w_dff_B_6pyf0hvZ3_0),.dout(w_dff_B_2CBrTZA57_0),.clk(gclk));
	jdff dff_B_UZNijE2z1_1(.din(n387),.dout(w_dff_B_UZNijE2z1_1),.clk(gclk));
	jdff dff_B_3LU1e96R4_1(.din(w_dff_B_UZNijE2z1_1),.dout(w_dff_B_3LU1e96R4_1),.clk(gclk));
	jdff dff_B_XRT4DgV51_1(.din(w_dff_B_3LU1e96R4_1),.dout(w_dff_B_XRT4DgV51_1),.clk(gclk));
	jdff dff_B_YLPxsV2m2_1(.din(w_dff_B_XRT4DgV51_1),.dout(w_dff_B_YLPxsV2m2_1),.clk(gclk));
	jdff dff_B_eF1gTHkW1_1(.din(w_dff_B_YLPxsV2m2_1),.dout(w_dff_B_eF1gTHkW1_1),.clk(gclk));
	jdff dff_B_E0dRo7Ap4_1(.din(w_dff_B_eF1gTHkW1_1),.dout(w_dff_B_E0dRo7Ap4_1),.clk(gclk));
	jdff dff_B_pwYc6g3t5_1(.din(w_dff_B_E0dRo7Ap4_1),.dout(w_dff_B_pwYc6g3t5_1),.clk(gclk));
	jdff dff_B_1LJfeufW8_1(.din(w_dff_B_pwYc6g3t5_1),.dout(w_dff_B_1LJfeufW8_1),.clk(gclk));
	jdff dff_B_0NfAE29N8_1(.din(w_dff_B_1LJfeufW8_1),.dout(w_dff_B_0NfAE29N8_1),.clk(gclk));
	jdff dff_B_BPEUKfMy0_1(.din(w_dff_B_0NfAE29N8_1),.dout(w_dff_B_BPEUKfMy0_1),.clk(gclk));
	jdff dff_B_oEAOUbTH8_1(.din(n388),.dout(w_dff_B_oEAOUbTH8_1),.clk(gclk));
	jdff dff_B_gJRVFlMj1_1(.din(w_dff_B_oEAOUbTH8_1),.dout(w_dff_B_gJRVFlMj1_1),.clk(gclk));
	jdff dff_B_E5vJf1TA7_1(.din(w_dff_B_gJRVFlMj1_1),.dout(w_dff_B_E5vJf1TA7_1),.clk(gclk));
	jdff dff_B_PQc7fllE3_1(.din(w_dff_B_E5vJf1TA7_1),.dout(w_dff_B_PQc7fllE3_1),.clk(gclk));
	jdff dff_B_9ixuTAQ49_1(.din(w_dff_B_PQc7fllE3_1),.dout(w_dff_B_9ixuTAQ49_1),.clk(gclk));
	jdff dff_B_UtgkDoeP8_1(.din(w_dff_B_9ixuTAQ49_1),.dout(w_dff_B_UtgkDoeP8_1),.clk(gclk));
	jdff dff_B_qejEdbeU3_1(.din(w_dff_B_UtgkDoeP8_1),.dout(w_dff_B_qejEdbeU3_1),.clk(gclk));
	jdff dff_B_rmn6hfnz2_1(.din(w_dff_B_qejEdbeU3_1),.dout(w_dff_B_rmn6hfnz2_1),.clk(gclk));
	jdff dff_B_A3NTip0I7_1(.din(w_dff_B_rmn6hfnz2_1),.dout(w_dff_B_A3NTip0I7_1),.clk(gclk));
	jdff dff_A_d2q87DtS4_1(.dout(w_n329_0[1]),.din(w_dff_A_d2q87DtS4_1),.clk(gclk));
	jdff dff_A_XFTT5lTa1_1(.dout(w_dff_A_d2q87DtS4_1),.din(w_dff_A_XFTT5lTa1_1),.clk(gclk));
	jdff dff_A_DAZQY4LC8_1(.dout(w_dff_A_XFTT5lTa1_1),.din(w_dff_A_DAZQY4LC8_1),.clk(gclk));
	jdff dff_A_rxU9HR7l9_1(.dout(w_dff_A_DAZQY4LC8_1),.din(w_dff_A_rxU9HR7l9_1),.clk(gclk));
	jdff dff_A_NFzSnkBu4_1(.dout(w_dff_A_rxU9HR7l9_1),.din(w_dff_A_NFzSnkBu4_1),.clk(gclk));
	jdff dff_A_hzmtlQNW0_1(.dout(w_dff_A_NFzSnkBu4_1),.din(w_dff_A_hzmtlQNW0_1),.clk(gclk));
	jdff dff_A_XLbgnOm52_1(.dout(w_dff_A_hzmtlQNW0_1),.din(w_dff_A_XLbgnOm52_1),.clk(gclk));
	jdff dff_A_TBEbmUIM3_1(.dout(w_dff_A_XLbgnOm52_1),.din(w_dff_A_TBEbmUIM3_1),.clk(gclk));
	jdff dff_A_92L2Is1y1_1(.dout(w_dff_A_TBEbmUIM3_1),.din(w_dff_A_92L2Is1y1_1),.clk(gclk));
	jdff dff_A_g1NKNY736_1(.dout(w_dff_A_92L2Is1y1_1),.din(w_dff_A_g1NKNY736_1),.clk(gclk));
	jdff dff_A_9ojVpIRN3_1(.dout(w_n328_0[1]),.din(w_dff_A_9ojVpIRN3_1),.clk(gclk));
	jdff dff_A_08R7Lev64_1(.dout(w_dff_A_9ojVpIRN3_1),.din(w_dff_A_08R7Lev64_1),.clk(gclk));
	jdff dff_A_WdjsqJVn3_1(.dout(w_dff_A_08R7Lev64_1),.din(w_dff_A_WdjsqJVn3_1),.clk(gclk));
	jdff dff_A_n8CJ7ICn0_1(.dout(w_dff_A_WdjsqJVn3_1),.din(w_dff_A_n8CJ7ICn0_1),.clk(gclk));
	jdff dff_A_R8Vs0EG03_1(.dout(w_dff_A_n8CJ7ICn0_1),.din(w_dff_A_R8Vs0EG03_1),.clk(gclk));
	jdff dff_A_mV0FOiNZ9_1(.dout(w_dff_A_R8Vs0EG03_1),.din(w_dff_A_mV0FOiNZ9_1),.clk(gclk));
	jdff dff_A_CMxlevNE6_1(.dout(w_dff_A_mV0FOiNZ9_1),.din(w_dff_A_CMxlevNE6_1),.clk(gclk));
	jdff dff_A_RUTyJ0s48_1(.dout(w_dff_A_CMxlevNE6_1),.din(w_dff_A_RUTyJ0s48_1),.clk(gclk));
	jdff dff_A_MM3tbpEL4_1(.dout(w_dff_A_RUTyJ0s48_1),.din(w_dff_A_MM3tbpEL4_1),.clk(gclk));
	jdff dff_A_l4Ds0gqY9_1(.dout(w_dff_A_MM3tbpEL4_1),.din(w_dff_A_l4Ds0gqY9_1),.clk(gclk));
	jdff dff_A_GAhtxgvl0_1(.dout(w_dff_A_l4Ds0gqY9_1),.din(w_dff_A_GAhtxgvl0_1),.clk(gclk));
	jdff dff_A_yf3Es2g00_0(.dout(w_G171gat_1[0]),.din(w_dff_A_yf3Es2g00_0),.clk(gclk));
	jdff dff_A_USrduznW5_0(.dout(w_dff_A_yf3Es2g00_0),.din(w_dff_A_USrduznW5_0),.clk(gclk));
	jdff dff_A_RyCpXcoG7_0(.dout(w_dff_A_USrduznW5_0),.din(w_dff_A_RyCpXcoG7_0),.clk(gclk));
	jdff dff_A_RlEP8WcD4_0(.dout(w_dff_A_RyCpXcoG7_0),.din(w_dff_A_RlEP8WcD4_0),.clk(gclk));
	jdff dff_A_19Wqj0xR3_0(.dout(w_dff_A_RlEP8WcD4_0),.din(w_dff_A_19Wqj0xR3_0),.clk(gclk));
	jdff dff_A_LfoXiNxK0_0(.dout(w_dff_A_19Wqj0xR3_0),.din(w_dff_A_LfoXiNxK0_0),.clk(gclk));
	jdff dff_A_5l1pAPm48_0(.dout(w_dff_A_LfoXiNxK0_0),.din(w_dff_A_5l1pAPm48_0),.clk(gclk));
	jdff dff_A_XRapL5ry9_0(.dout(w_dff_A_5l1pAPm48_0),.din(w_dff_A_XRapL5ry9_0),.clk(gclk));
	jdff dff_A_5UnxKDUu8_0(.dout(w_dff_A_XRapL5ry9_0),.din(w_dff_A_5UnxKDUu8_0),.clk(gclk));
	jdff dff_A_ppOcJGmE8_1(.dout(w_G171gat_1[1]),.din(w_dff_A_ppOcJGmE8_1),.clk(gclk));
	jdff dff_A_pioUJZBQ7_1(.dout(w_dff_A_ppOcJGmE8_1),.din(w_dff_A_pioUJZBQ7_1),.clk(gclk));
	jdff dff_A_JYwpyw1R4_1(.dout(w_dff_A_pioUJZBQ7_1),.din(w_dff_A_JYwpyw1R4_1),.clk(gclk));
	jdff dff_A_Xyx0mOje4_1(.dout(w_dff_A_JYwpyw1R4_1),.din(w_dff_A_Xyx0mOje4_1),.clk(gclk));
	jdff dff_A_OzXuUR4n4_1(.dout(w_dff_A_Xyx0mOje4_1),.din(w_dff_A_OzXuUR4n4_1),.clk(gclk));
	jdff dff_A_4Fo6cjNh2_1(.dout(w_dff_A_OzXuUR4n4_1),.din(w_dff_A_4Fo6cjNh2_1),.clk(gclk));
	jdff dff_A_TS9LzjdN2_1(.dout(w_dff_A_4Fo6cjNh2_1),.din(w_dff_A_TS9LzjdN2_1),.clk(gclk));
	jdff dff_A_yrGGfm964_1(.dout(w_dff_A_TS9LzjdN2_1),.din(w_dff_A_yrGGfm964_1),.clk(gclk));
	jdff dff_A_SDHk0Ayh3_1(.dout(w_dff_A_yrGGfm964_1),.din(w_dff_A_SDHk0Ayh3_1),.clk(gclk));
	jdff dff_B_em656vaO0_1(.din(n403),.dout(w_dff_B_em656vaO0_1),.clk(gclk));
	jdff dff_B_LNaa5wLb6_0(.din(n408),.dout(w_dff_B_LNaa5wLb6_0),.clk(gclk));
	jdff dff_B_6GQCrwjA3_0(.din(w_dff_B_LNaa5wLb6_0),.dout(w_dff_B_6GQCrwjA3_0),.clk(gclk));
	jdff dff_B_0VR8D4NB0_0(.din(n406),.dout(w_dff_B_0VR8D4NB0_0),.clk(gclk));
	jdff dff_B_LH3CBpk42_0(.din(w_dff_B_0VR8D4NB0_0),.dout(w_dff_B_LH3CBpk42_0),.clk(gclk));
	jdff dff_B_Qr1Exhr47_0(.din(w_dff_B_LH3CBpk42_0),.dout(w_dff_B_Qr1Exhr47_0),.clk(gclk));
	jdff dff_B_vXtvioYj5_0(.din(w_dff_B_Qr1Exhr47_0),.dout(w_dff_B_vXtvioYj5_0),.clk(gclk));
	jdff dff_B_WNAWS9qW8_0(.din(w_dff_B_vXtvioYj5_0),.dout(w_dff_B_WNAWS9qW8_0),.clk(gclk));
	jdff dff_B_BWDOHGqr9_0(.din(w_dff_B_WNAWS9qW8_0),.dout(w_dff_B_BWDOHGqr9_0),.clk(gclk));
	jdff dff_B_LAuNqCAH6_0(.din(w_dff_B_BWDOHGqr9_0),.dout(w_dff_B_LAuNqCAH6_0),.clk(gclk));
	jdff dff_B_ZlYS1TIf0_0(.din(w_dff_B_LAuNqCAH6_0),.dout(w_dff_B_ZlYS1TIf0_0),.clk(gclk));
	jdff dff_B_8yfsx2nm3_0(.din(w_dff_B_ZlYS1TIf0_0),.dout(w_dff_B_8yfsx2nm3_0),.clk(gclk));
	jdff dff_B_wTQ1267p5_0(.din(w_dff_B_8yfsx2nm3_0),.dout(w_dff_B_wTQ1267p5_0),.clk(gclk));
	jdff dff_A_YiYdZcsI5_1(.dout(w_G91gat_0[1]),.din(w_dff_A_YiYdZcsI5_1),.clk(gclk));
	jdff dff_A_lIdggpTg7_1(.dout(w_dff_A_YiYdZcsI5_1),.din(w_dff_A_lIdggpTg7_1),.clk(gclk));
	jdff dff_A_Bx15hbLn1_1(.dout(w_dff_A_lIdggpTg7_1),.din(w_dff_A_Bx15hbLn1_1),.clk(gclk));
	jdff dff_A_z2n6usdp9_1(.dout(w_dff_A_Bx15hbLn1_1),.din(w_dff_A_z2n6usdp9_1),.clk(gclk));
	jdff dff_A_hHT4DfCN8_1(.dout(w_dff_A_z2n6usdp9_1),.din(w_dff_A_hHT4DfCN8_1),.clk(gclk));
	jdff dff_A_pSUFoYvh7_1(.dout(w_dff_A_hHT4DfCN8_1),.din(w_dff_A_pSUFoYvh7_1),.clk(gclk));
	jdff dff_A_BcMDqKgm5_1(.dout(w_n404_0[1]),.din(w_dff_A_BcMDqKgm5_1),.clk(gclk));
	jdff dff_A_SCgwyVPp8_1(.dout(w_dff_A_BcMDqKgm5_1),.din(w_dff_A_SCgwyVPp8_1),.clk(gclk));
	jdff dff_A_86jZxEJm1_1(.dout(w_dff_A_SCgwyVPp8_1),.din(w_dff_A_86jZxEJm1_1),.clk(gclk));
	jdff dff_A_iFAjw0GP6_1(.dout(w_dff_A_86jZxEJm1_1),.din(w_dff_A_iFAjw0GP6_1),.clk(gclk));
	jdff dff_A_BvksVKM82_1(.dout(w_dff_A_iFAjw0GP6_1),.din(w_dff_A_BvksVKM82_1),.clk(gclk));
	jdff dff_A_zHL6klVf2_1(.dout(w_dff_A_BvksVKM82_1),.din(w_dff_A_zHL6klVf2_1),.clk(gclk));
	jdff dff_A_ogtdX02Z2_1(.dout(w_dff_A_zHL6klVf2_1),.din(w_dff_A_ogtdX02Z2_1),.clk(gclk));
	jdff dff_A_f7gAH5oF8_1(.dout(w_dff_A_ogtdX02Z2_1),.din(w_dff_A_f7gAH5oF8_1),.clk(gclk));
	jdff dff_A_lcXQg14O7_1(.dout(w_dff_A_f7gAH5oF8_1),.din(w_dff_A_lcXQg14O7_1),.clk(gclk));
	jdff dff_A_FodcDkDs4_1(.dout(w_dff_A_lcXQg14O7_1),.din(w_dff_A_FodcDkDs4_1),.clk(gclk));
	jdff dff_A_JJoZkWO27_1(.dout(w_dff_A_FodcDkDs4_1),.din(w_dff_A_JJoZkWO27_1),.clk(gclk));
	jdff dff_A_Xa5F2hGi1_1(.dout(w_dff_A_JJoZkWO27_1),.din(w_dff_A_Xa5F2hGi1_1),.clk(gclk));
	jdff dff_B_py9DwAIB7_0(.din(n317),.dout(w_dff_B_py9DwAIB7_0),.clk(gclk));
	jdff dff_B_ME3aqBur3_0(.din(n316),.dout(w_dff_B_ME3aqBur3_0),.clk(gclk));
	jdff dff_B_FGhC9g0D4_0(.din(w_dff_B_ME3aqBur3_0),.dout(w_dff_B_FGhC9g0D4_0),.clk(gclk));
	jdff dff_B_8IAzCC8t9_0(.din(w_dff_B_FGhC9g0D4_0),.dout(w_dff_B_8IAzCC8t9_0),.clk(gclk));
	jdff dff_B_sDlKO3YR9_0(.din(w_dff_B_8IAzCC8t9_0),.dout(w_dff_B_sDlKO3YR9_0),.clk(gclk));
	jdff dff_A_aNQIUORM4_0(.dout(w_n306_1[0]),.din(w_dff_A_aNQIUORM4_0),.clk(gclk));
	jdff dff_A_6ZGK6Eos5_0(.dout(w_dff_A_aNQIUORM4_0),.din(w_dff_A_6ZGK6Eos5_0),.clk(gclk));
	jdff dff_A_f16D6L1E6_1(.dout(w_G165gat_0[1]),.din(w_dff_A_f16D6L1E6_1),.clk(gclk));
	jdff dff_A_VMDtzSMh3_1(.dout(w_dff_A_f16D6L1E6_1),.din(w_dff_A_VMDtzSMh3_1),.clk(gclk));
	jdff dff_A_2H6Iw6yB7_1(.dout(w_dff_A_VMDtzSMh3_1),.din(w_dff_A_2H6Iw6yB7_1),.clk(gclk));
	jdff dff_A_di2SfrFP5_1(.dout(w_dff_A_2H6Iw6yB7_1),.din(w_dff_A_di2SfrFP5_1),.clk(gclk));
	jdff dff_A_ugTcDXZo3_1(.dout(w_dff_A_di2SfrFP5_1),.din(w_dff_A_ugTcDXZo3_1),.clk(gclk));
	jdff dff_A_ZzoTFIye8_1(.dout(w_dff_A_ugTcDXZo3_1),.din(w_dff_A_ZzoTFIye8_1),.clk(gclk));
	jdff dff_A_pfeKiM682_1(.dout(w_dff_A_ZzoTFIye8_1),.din(w_dff_A_pfeKiM682_1),.clk(gclk));
	jdff dff_A_D05oNxKZ1_1(.dout(w_dff_A_pfeKiM682_1),.din(w_dff_A_D05oNxKZ1_1),.clk(gclk));
	jdff dff_A_gV8tk6AY7_2(.dout(w_G165gat_0[2]),.din(w_dff_A_gV8tk6AY7_2),.clk(gclk));
	jdff dff_A_FCaw76er3_2(.dout(w_dff_A_gV8tk6AY7_2),.din(w_dff_A_FCaw76er3_2),.clk(gclk));
	jdff dff_A_ZTSQR2WJ0_2(.dout(w_dff_A_FCaw76er3_2),.din(w_dff_A_ZTSQR2WJ0_2),.clk(gclk));
	jdff dff_A_6KPCu3Km9_2(.dout(w_dff_A_ZTSQR2WJ0_2),.din(w_dff_A_6KPCu3Km9_2),.clk(gclk));
	jdff dff_A_ItNotLYK3_2(.dout(w_dff_A_6KPCu3Km9_2),.din(w_dff_A_ItNotLYK3_2),.clk(gclk));
	jdff dff_A_wwwFtVNb1_2(.dout(w_dff_A_ItNotLYK3_2),.din(w_dff_A_wwwFtVNb1_2),.clk(gclk));
	jdff dff_A_38dpMtXr9_2(.dout(w_dff_A_wwwFtVNb1_2),.din(w_dff_A_38dpMtXr9_2),.clk(gclk));
	jdff dff_A_md0ncrWr1_2(.dout(w_dff_A_38dpMtXr9_2),.din(w_dff_A_md0ncrWr1_2),.clk(gclk));
	jdff dff_A_BTy1ECCB1_2(.dout(w_dff_A_md0ncrWr1_2),.din(w_dff_A_BTy1ECCB1_2),.clk(gclk));
	jdff dff_A_ZuaxcF6B6_2(.dout(w_dff_A_BTy1ECCB1_2),.din(w_dff_A_ZuaxcF6B6_2),.clk(gclk));
	jdff dff_B_epr6vjWz6_3(.din(G165gat),.dout(w_dff_B_epr6vjWz6_3),.clk(gclk));
	jdff dff_B_TjZuYqWm5_1(.din(n426),.dout(w_dff_B_TjZuYqWm5_1),.clk(gclk));
	jdff dff_B_RQ8n5l5u4_1(.din(w_dff_B_TjZuYqWm5_1),.dout(w_dff_B_RQ8n5l5u4_1),.clk(gclk));
	jdff dff_B_8YmqLXfr9_1(.din(w_dff_B_RQ8n5l5u4_1),.dout(w_dff_B_8YmqLXfr9_1),.clk(gclk));
	jdff dff_B_SsrziKMG3_1(.din(w_dff_B_8YmqLXfr9_1),.dout(w_dff_B_SsrziKMG3_1),.clk(gclk));
	jdff dff_B_9DIcCkY60_1(.din(w_dff_B_SsrziKMG3_1),.dout(w_dff_B_9DIcCkY60_1),.clk(gclk));
	jdff dff_B_nUPNL3Do2_1(.din(w_dff_B_9DIcCkY60_1),.dout(w_dff_B_nUPNL3Do2_1),.clk(gclk));
	jdff dff_B_7T0nKnwn6_1(.din(w_dff_B_nUPNL3Do2_1),.dout(w_dff_B_7T0nKnwn6_1),.clk(gclk));
	jdff dff_B_Ypdj6s0X1_1(.din(w_dff_B_7T0nKnwn6_1),.dout(w_dff_B_Ypdj6s0X1_1),.clk(gclk));
	jdff dff_B_lvNTZ2L67_1(.din(w_dff_B_Ypdj6s0X1_1),.dout(w_dff_B_lvNTZ2L67_1),.clk(gclk));
	jdff dff_B_EwFU9vN70_1(.din(n428),.dout(w_dff_B_EwFU9vN70_1),.clk(gclk));
	jdff dff_B_W3z3T0lt7_1(.din(n340),.dout(w_dff_B_W3z3T0lt7_1),.clk(gclk));
	jdff dff_B_YvFDfzdB1_1(.din(w_dff_B_W3z3T0lt7_1),.dout(w_dff_B_YvFDfzdB1_1),.clk(gclk));
	jdff dff_B_OXuQGpJw2_1(.din(w_dff_B_YvFDfzdB1_1),.dout(w_dff_B_OXuQGpJw2_1),.clk(gclk));
	jdff dff_B_6DpSRe6W7_1(.din(w_dff_B_OXuQGpJw2_1),.dout(w_dff_B_6DpSRe6W7_1),.clk(gclk));
	jdff dff_B_pcnzQFld0_1(.din(w_dff_B_6DpSRe6W7_1),.dout(w_dff_B_pcnzQFld0_1),.clk(gclk));
	jdff dff_B_8Q9L2Ugr5_1(.din(w_dff_B_pcnzQFld0_1),.dout(w_dff_B_8Q9L2Ugr5_1),.clk(gclk));
	jdff dff_B_GmmfPo5h3_1(.din(n344),.dout(w_dff_B_GmmfPo5h3_1),.clk(gclk));
	jdff dff_B_EY4aSTkf0_1(.din(w_dff_B_GmmfPo5h3_1),.dout(w_dff_B_EY4aSTkf0_1),.clk(gclk));
	jdff dff_B_yoby2iPW5_1(.din(w_dff_B_EY4aSTkf0_1),.dout(w_dff_B_yoby2iPW5_1),.clk(gclk));
	jdff dff_B_id5kLjQl1_1(.din(w_dff_B_yoby2iPW5_1),.dout(w_dff_B_id5kLjQl1_1),.clk(gclk));
	jdff dff_B_vbu4v1jM8_1(.din(w_dff_B_id5kLjQl1_1),.dout(w_dff_B_vbu4v1jM8_1),.clk(gclk));
	jdff dff_B_rl9Vq7JE8_0(.din(n171),.dout(w_dff_B_rl9Vq7JE8_0),.clk(gclk));
	jdff dff_A_rWOHNZkG3_1(.dout(w_G219gat_1[1]),.din(w_dff_A_rWOHNZkG3_1),.clk(gclk));
	jdff dff_A_sqprAlgC0_1(.dout(w_dff_A_rWOHNZkG3_1),.din(w_dff_A_sqprAlgC0_1),.clk(gclk));
	jdff dff_A_lslrCMJR3_2(.dout(w_G219gat_1[2]),.din(w_dff_A_lslrCMJR3_2),.clk(gclk));
	jdff dff_A_UUauDlHl2_2(.dout(w_dff_A_lslrCMJR3_2),.din(w_dff_A_UUauDlHl2_2),.clk(gclk));
	jdff dff_A_QObBHfh02_2(.dout(w_dff_A_UUauDlHl2_2),.din(w_dff_A_QObBHfh02_2),.clk(gclk));
	jdff dff_A_4Sd4npID9_2(.dout(w_dff_A_QObBHfh02_2),.din(w_dff_A_4Sd4npID9_2),.clk(gclk));
	jdff dff_A_O1Lucx3I5_0(.dout(w_G219gat_0[0]),.din(w_dff_A_O1Lucx3I5_0),.clk(gclk));
	jdff dff_A_uzqWPfXI1_0(.dout(w_dff_A_O1Lucx3I5_0),.din(w_dff_A_uzqWPfXI1_0),.clk(gclk));
	jdff dff_A_a1FPNMpL1_0(.dout(w_dff_A_uzqWPfXI1_0),.din(w_dff_A_a1FPNMpL1_0),.clk(gclk));
	jdff dff_A_asF04T9x1_0(.dout(w_dff_A_a1FPNMpL1_0),.din(w_dff_A_asF04T9x1_0),.clk(gclk));
	jdff dff_A_edw16gTV5_0(.dout(w_dff_A_asF04T9x1_0),.din(w_dff_A_edw16gTV5_0),.clk(gclk));
	jdff dff_A_kOUkT3XB5_0(.dout(w_dff_A_edw16gTV5_0),.din(w_dff_A_kOUkT3XB5_0),.clk(gclk));
	jdff dff_A_jtlU4Qz41_0(.dout(w_dff_A_kOUkT3XB5_0),.din(w_dff_A_jtlU4Qz41_0),.clk(gclk));
	jdff dff_A_yV2b8S5z8_0(.dout(w_dff_A_jtlU4Qz41_0),.din(w_dff_A_yV2b8S5z8_0),.clk(gclk));
	jdff dff_A_SfnO8thz7_0(.dout(w_dff_A_yV2b8S5z8_0),.din(w_dff_A_SfnO8thz7_0),.clk(gclk));
	jdff dff_A_sMiNjPDH1_1(.dout(w_G219gat_0[1]),.din(w_dff_A_sMiNjPDH1_1),.clk(gclk));
	jdff dff_B_PLaI4vFA4_3(.din(G219gat),.dout(w_dff_B_PLaI4vFA4_3),.clk(gclk));
	jdff dff_B_UIDBElnm6_3(.din(w_dff_B_PLaI4vFA4_3),.dout(w_dff_B_UIDBElnm6_3),.clk(gclk));
	jdff dff_B_wqnAYARH5_3(.din(w_dff_B_UIDBElnm6_3),.dout(w_dff_B_wqnAYARH5_3),.clk(gclk));
	jdff dff_B_BfeD4erD1_3(.din(w_dff_B_wqnAYARH5_3),.dout(w_dff_B_BfeD4erD1_3),.clk(gclk));
	jdff dff_B_R9hstALJ1_3(.din(w_dff_B_BfeD4erD1_3),.dout(w_dff_B_R9hstALJ1_3),.clk(gclk));
	jdff dff_B_o3Pi5RmB4_3(.din(w_dff_B_R9hstALJ1_3),.dout(w_dff_B_o3Pi5RmB4_3),.clk(gclk));
	jdff dff_B_ptPcvAMe1_3(.din(w_dff_B_o3Pi5RmB4_3),.dout(w_dff_B_ptPcvAMe1_3),.clk(gclk));
	jdff dff_B_q7NuIUaE4_3(.din(w_dff_B_ptPcvAMe1_3),.dout(w_dff_B_q7NuIUaE4_3),.clk(gclk));
	jdff dff_B_2xljmZZE0_3(.din(w_dff_B_q7NuIUaE4_3),.dout(w_dff_B_2xljmZZE0_3),.clk(gclk));
	jdff dff_B_R3Xi5MM07_3(.din(w_dff_B_2xljmZZE0_3),.dout(w_dff_B_R3Xi5MM07_3),.clk(gclk));
	jdff dff_B_cexpfoTi9_3(.din(w_dff_B_R3Xi5MM07_3),.dout(w_dff_B_cexpfoTi9_3),.clk(gclk));
	jdff dff_B_kEi3TNjC8_3(.din(w_dff_B_cexpfoTi9_3),.dout(w_dff_B_kEi3TNjC8_3),.clk(gclk));
	jdff dff_B_9wLbiQPo5_0(.din(n427),.dout(w_dff_B_9wLbiQPo5_0),.clk(gclk));
	jdff dff_B_KjaHok4l3_0(.din(w_dff_B_9wLbiQPo5_0),.dout(w_dff_B_KjaHok4l3_0),.clk(gclk));
	jdff dff_B_CgkK8ZDX5_0(.din(w_dff_B_KjaHok4l3_0),.dout(w_dff_B_CgkK8ZDX5_0),.clk(gclk));
	jdff dff_B_cvEIrjfx2_0(.din(w_dff_B_CgkK8ZDX5_0),.dout(w_dff_B_cvEIrjfx2_0),.clk(gclk));
	jdff dff_B_onPodhm80_0(.din(w_dff_B_cvEIrjfx2_0),.dout(w_dff_B_onPodhm80_0),.clk(gclk));
	jdff dff_B_csD3o8sT0_0(.din(w_dff_B_onPodhm80_0),.dout(w_dff_B_csD3o8sT0_0),.clk(gclk));
	jdff dff_B_TnQ6bYOD9_0(.din(w_dff_B_csD3o8sT0_0),.dout(w_dff_B_TnQ6bYOD9_0),.clk(gclk));
	jdff dff_B_WB2r8z254_0(.din(w_dff_B_TnQ6bYOD9_0),.dout(w_dff_B_WB2r8z254_0),.clk(gclk));
	jdff dff_B_bOfGwb3m3_0(.din(w_dff_B_WB2r8z254_0),.dout(w_dff_B_bOfGwb3m3_0),.clk(gclk));
	jdff dff_B_WSMxIz7D4_1(.din(n389),.dout(w_dff_B_WSMxIz7D4_1),.clk(gclk));
	jdff dff_B_xeCAAGe97_1(.din(w_dff_B_WSMxIz7D4_1),.dout(w_dff_B_xeCAAGe97_1),.clk(gclk));
	jdff dff_B_wPr6t00I9_1(.din(w_dff_B_xeCAAGe97_1),.dout(w_dff_B_wPr6t00I9_1),.clk(gclk));
	jdff dff_B_oQvKxCeK5_1(.din(w_dff_B_wPr6t00I9_1),.dout(w_dff_B_oQvKxCeK5_1),.clk(gclk));
	jdff dff_B_rBwTdNrd7_1(.din(w_dff_B_oQvKxCeK5_1),.dout(w_dff_B_rBwTdNrd7_1),.clk(gclk));
	jdff dff_B_MIa4ORsT9_1(.din(w_dff_B_rBwTdNrd7_1),.dout(w_dff_B_MIa4ORsT9_1),.clk(gclk));
	jdff dff_B_eALyMLm19_1(.din(w_dff_B_MIa4ORsT9_1),.dout(w_dff_B_eALyMLm19_1),.clk(gclk));
	jdff dff_B_9YbA9GZ99_1(.din(w_dff_B_eALyMLm19_1),.dout(w_dff_B_9YbA9GZ99_1),.clk(gclk));
	jdff dff_B_2niJCX933_1(.din(n359),.dout(w_dff_B_2niJCX933_1),.clk(gclk));
	jdff dff_B_2tdBkyD23_1(.din(w_dff_B_2niJCX933_1),.dout(w_dff_B_2tdBkyD23_1),.clk(gclk));
	jdff dff_B_L7mGhCgb8_1(.din(w_dff_B_2tdBkyD23_1),.dout(w_dff_B_L7mGhCgb8_1),.clk(gclk));
	jdff dff_B_YBwhKsRa3_1(.din(w_dff_B_L7mGhCgb8_1),.dout(w_dff_B_YBwhKsRa3_1),.clk(gclk));
	jdff dff_B_NjjmpL1C0_1(.din(w_dff_B_YBwhKsRa3_1),.dout(w_dff_B_NjjmpL1C0_1),.clk(gclk));
	jdff dff_B_axRcZCmb1_1(.din(w_dff_B_NjjmpL1C0_1),.dout(w_dff_B_axRcZCmb1_1),.clk(gclk));
	jdff dff_B_Y9ex9KpT5_1(.din(w_dff_B_axRcZCmb1_1),.dout(w_dff_B_Y9ex9KpT5_1),.clk(gclk));
	jdff dff_B_qKC3uJD64_1(.din(n252),.dout(w_dff_B_qKC3uJD64_1),.clk(gclk));
	jdff dff_B_VXLgkgsg4_1(.din(w_dff_B_qKC3uJD64_1),.dout(w_dff_B_VXLgkgsg4_1),.clk(gclk));
	jdff dff_B_IGXkI59T7_1(.din(w_dff_B_VXLgkgsg4_1),.dout(w_dff_B_IGXkI59T7_1),.clk(gclk));
	jdff dff_B_ZEdnkMpZ5_1(.din(w_dff_B_IGXkI59T7_1),.dout(w_dff_B_ZEdnkMpZ5_1),.clk(gclk));
	jdff dff_B_XRitnMuY1_1(.din(w_dff_B_ZEdnkMpZ5_1),.dout(w_dff_B_XRitnMuY1_1),.clk(gclk));
	jdff dff_B_BjzQLaOI5_1(.din(n253),.dout(w_dff_B_BjzQLaOI5_1),.clk(gclk));
	jdff dff_B_YfHJEGy66_1(.din(w_dff_B_BjzQLaOI5_1),.dout(w_dff_B_YfHJEGy66_1),.clk(gclk));
	jdff dff_B_EXS4HU1R9_1(.din(w_dff_B_YfHJEGy66_1),.dout(w_dff_B_EXS4HU1R9_1),.clk(gclk));
	jdff dff_B_a0X6tw2p1_1(.din(w_dff_B_EXS4HU1R9_1),.dout(w_dff_B_a0X6tw2p1_1),.clk(gclk));
	jdff dff_B_LVXLDEJp9_1(.din(n254),.dout(w_dff_B_LVXLDEJp9_1),.clk(gclk));
	jdff dff_B_5z8THAnV5_1(.din(w_dff_B_LVXLDEJp9_1),.dout(w_dff_B_5z8THAnV5_1),.clk(gclk));
	jdff dff_B_E84IDsFC6_1(.din(w_dff_B_5z8THAnV5_1),.dout(w_dff_B_E84IDsFC6_1),.clk(gclk));
	jdff dff_B_a8bqaFgB0_1(.din(n255),.dout(w_dff_B_a8bqaFgB0_1),.clk(gclk));
	jdff dff_B_E40CS4Av2_1(.din(w_dff_B_a8bqaFgB0_1),.dout(w_dff_B_E40CS4Av2_1),.clk(gclk));
	jdff dff_A_r3WANGgp2_1(.dout(w_n209_0[1]),.din(w_dff_A_r3WANGgp2_1),.clk(gclk));
	jdff dff_B_TcBGh5e38_2(.din(n209),.dout(w_dff_B_TcBGh5e38_2),.clk(gclk));
	jdff dff_B_GZI1XtSJ9_2(.din(w_dff_B_TcBGh5e38_2),.dout(w_dff_B_GZI1XtSJ9_2),.clk(gclk));
	jdff dff_B_qJeypqZ09_2(.din(w_dff_B_GZI1XtSJ9_2),.dout(w_dff_B_qJeypqZ09_2),.clk(gclk));
	jdff dff_B_GdrfCwyA0_2(.din(w_dff_B_qJeypqZ09_2),.dout(w_dff_B_GdrfCwyA0_2),.clk(gclk));
	jdff dff_B_gjPcV6FL6_2(.din(w_dff_B_GdrfCwyA0_2),.dout(w_dff_B_gjPcV6FL6_2),.clk(gclk));
	jdff dff_B_Od2j9ylF8_2(.din(w_dff_B_gjPcV6FL6_2),.dout(w_dff_B_Od2j9ylF8_2),.clk(gclk));
	jdff dff_B_hmAaJchv4_2(.din(w_dff_B_Od2j9ylF8_2),.dout(w_dff_B_hmAaJchv4_2),.clk(gclk));
	jdff dff_B_yM4KmRWJ9_2(.din(w_dff_B_hmAaJchv4_2),.dout(w_dff_B_yM4KmRWJ9_2),.clk(gclk));
	jdff dff_B_OnztqHNG8_2(.din(w_dff_B_yM4KmRWJ9_2),.dout(w_dff_B_OnztqHNG8_2),.clk(gclk));
	jdff dff_A_3MnImfhx0_0(.dout(w_G261gat_0[0]),.din(w_dff_A_3MnImfhx0_0),.clk(gclk));
	jdff dff_A_hbDEDvy40_0(.dout(w_dff_A_3MnImfhx0_0),.din(w_dff_A_hbDEDvy40_0),.clk(gclk));
	jdff dff_A_96Mgs9Aq8_0(.dout(w_dff_A_hbDEDvy40_0),.din(w_dff_A_96Mgs9Aq8_0),.clk(gclk));
	jdff dff_A_URHxRA7b2_0(.dout(w_dff_A_96Mgs9Aq8_0),.din(w_dff_A_URHxRA7b2_0),.clk(gclk));
	jdff dff_A_5gUO1yCr0_0(.dout(w_dff_A_URHxRA7b2_0),.din(w_dff_A_5gUO1yCr0_0),.clk(gclk));
	jdff dff_A_LAyl2Q3X3_0(.dout(w_dff_A_5gUO1yCr0_0),.din(w_dff_A_LAyl2Q3X3_0),.clk(gclk));
	jdff dff_A_AhYmlxv09_0(.dout(w_dff_A_LAyl2Q3X3_0),.din(w_dff_A_AhYmlxv09_0),.clk(gclk));
	jdff dff_A_dGt58nX79_0(.dout(w_dff_A_AhYmlxv09_0),.din(w_dff_A_dGt58nX79_0),.clk(gclk));
	jdff dff_A_GVhlbfMO6_0(.dout(w_dff_A_dGt58nX79_0),.din(w_dff_A_GVhlbfMO6_0),.clk(gclk));
	jdff dff_A_ccCzQTdh6_0(.dout(w_dff_A_GVhlbfMO6_0),.din(w_dff_A_ccCzQTdh6_0),.clk(gclk));
	jdff dff_A_xhCMx9Wp1_2(.dout(w_G261gat_0[2]),.din(w_dff_A_xhCMx9Wp1_2),.clk(gclk));
	jdff dff_A_gQCTnKEc5_2(.dout(w_dff_A_xhCMx9Wp1_2),.din(w_dff_A_gQCTnKEc5_2),.clk(gclk));
	jdff dff_A_Oo3s6GkZ7_2(.dout(w_dff_A_gQCTnKEc5_2),.din(w_dff_A_Oo3s6GkZ7_2),.clk(gclk));
	jdff dff_A_Utk7lrqA7_2(.dout(w_dff_A_Oo3s6GkZ7_2),.din(w_dff_A_Utk7lrqA7_2),.clk(gclk));
	jdff dff_A_HNm7eEoG8_2(.dout(w_dff_A_Utk7lrqA7_2),.din(w_dff_A_HNm7eEoG8_2),.clk(gclk));
	jdff dff_A_zV5pQmm24_2(.dout(w_dff_A_HNm7eEoG8_2),.din(w_dff_A_zV5pQmm24_2),.clk(gclk));
	jdff dff_A_mPWFUcQR4_2(.dout(w_dff_A_zV5pQmm24_2),.din(w_dff_A_mPWFUcQR4_2),.clk(gclk));
	jdff dff_A_QeE2dAfw5_2(.dout(w_dff_A_mPWFUcQR4_2),.din(w_dff_A_QeE2dAfw5_2),.clk(gclk));
	jdff dff_A_GcNMlFBW8_2(.dout(w_dff_A_QeE2dAfw5_2),.din(w_dff_A_GcNMlFBW8_2),.clk(gclk));
	jdff dff_A_TBAA5QPO6_2(.dout(w_dff_A_GcNMlFBW8_2),.din(w_dff_A_TBAA5QPO6_2),.clk(gclk));
	jdff dff_A_DB211iR03_0(.dout(w_n242_0[0]),.din(w_dff_A_DB211iR03_0),.clk(gclk));
	jdff dff_B_f9PFycb75_1(.din(n182),.dout(w_dff_B_f9PFycb75_1),.clk(gclk));
	jdff dff_B_02REkNbb6_1(.din(n191),.dout(w_dff_B_02REkNbb6_1),.clk(gclk));
	jdff dff_B_y2AXDNAR1_1(.din(w_dff_B_02REkNbb6_1),.dout(w_dff_B_y2AXDNAR1_1),.clk(gclk));
	jdff dff_B_7CUkmzZD5_1(.din(w_dff_B_y2AXDNAR1_1),.dout(w_dff_B_7CUkmzZD5_1),.clk(gclk));
	jdff dff_B_ObvjXfyc0_1(.din(w_dff_B_7CUkmzZD5_1),.dout(w_dff_B_ObvjXfyc0_1),.clk(gclk));
	jdff dff_B_kvx6MqsJ7_1(.din(w_dff_B_ObvjXfyc0_1),.dout(w_dff_B_kvx6MqsJ7_1),.clk(gclk));
	jdff dff_B_HnluH0Uh6_1(.din(n183),.dout(w_dff_B_HnluH0Uh6_1),.clk(gclk));
	jdff dff_B_901NAY6l2_1(.din(w_dff_B_HnluH0Uh6_1),.dout(w_dff_B_901NAY6l2_1),.clk(gclk));
	jdff dff_B_XmavlbES5_1(.din(w_dff_B_901NAY6l2_1),.dout(w_dff_B_XmavlbES5_1),.clk(gclk));
	jdff dff_B_hKw61krO9_1(.din(w_dff_B_XmavlbES5_1),.dout(w_dff_B_hKw61krO9_1),.clk(gclk));
	jdff dff_B_jn0YtmUD9_1(.din(w_dff_B_hKw61krO9_1),.dout(w_dff_B_jn0YtmUD9_1),.clk(gclk));
	jdff dff_B_BJriCuaR1_1(.din(n184),.dout(w_dff_B_BJriCuaR1_1),.clk(gclk));
	jdff dff_A_dU3YKqVA4_1(.dout(w_G126gat_0[1]),.din(w_dff_A_dU3YKqVA4_1),.clk(gclk));
	jdff dff_A_7iacd3fw9_1(.dout(w_dff_A_dU3YKqVA4_1),.din(w_dff_A_7iacd3fw9_1),.clk(gclk));
	jdff dff_A_HyAzXTRm3_1(.dout(w_dff_A_7iacd3fw9_1),.din(w_dff_A_HyAzXTRm3_1),.clk(gclk));
	jdff dff_A_7HQPvZec9_1(.dout(w_dff_A_HyAzXTRm3_1),.din(w_dff_A_7HQPvZec9_1),.clk(gclk));
	jdff dff_A_RGLzaIRm5_1(.dout(w_dff_A_7HQPvZec9_1),.din(w_dff_A_RGLzaIRm5_1),.clk(gclk));
	jdff dff_A_IxPp00Gn2_1(.dout(w_dff_A_RGLzaIRm5_1),.din(w_dff_A_IxPp00Gn2_1),.clk(gclk));
	jdff dff_B_0z4F70Dg9_3(.din(n181),.dout(w_dff_B_0z4F70Dg9_3),.clk(gclk));
	jdff dff_B_Ythl7dYS6_3(.din(w_dff_B_0z4F70Dg9_3),.dout(w_dff_B_Ythl7dYS6_3),.clk(gclk));
	jdff dff_B_WZmIcOnv1_3(.din(w_dff_B_Ythl7dYS6_3),.dout(w_dff_B_WZmIcOnv1_3),.clk(gclk));
	jdff dff_B_xcZpoV7G9_3(.din(w_dff_B_WZmIcOnv1_3),.dout(w_dff_B_xcZpoV7G9_3),.clk(gclk));
	jdff dff_B_Mh9Rh9t26_3(.din(w_dff_B_xcZpoV7G9_3),.dout(w_dff_B_Mh9Rh9t26_3),.clk(gclk));
	jdff dff_B_AyRVInel9_3(.din(w_dff_B_Mh9Rh9t26_3),.dout(w_dff_B_AyRVInel9_3),.clk(gclk));
	jdff dff_B_zrgDDyU05_3(.din(w_dff_B_AyRVInel9_3),.dout(w_dff_B_zrgDDyU05_3),.clk(gclk));
	jdff dff_B_juyi9VzG8_3(.din(w_dff_B_zrgDDyU05_3),.dout(w_dff_B_juyi9VzG8_3),.clk(gclk));
	jdff dff_A_WAOntSsh3_1(.dout(w_G201gat_0[1]),.din(w_dff_A_WAOntSsh3_1),.clk(gclk));
	jdff dff_A_PKGxXbie3_1(.dout(w_dff_A_WAOntSsh3_1),.din(w_dff_A_PKGxXbie3_1),.clk(gclk));
	jdff dff_A_SnGcm0yV3_1(.dout(w_dff_A_PKGxXbie3_1),.din(w_dff_A_SnGcm0yV3_1),.clk(gclk));
	jdff dff_A_eT09wCdN9_1(.dout(w_dff_A_SnGcm0yV3_1),.din(w_dff_A_eT09wCdN9_1),.clk(gclk));
	jdff dff_A_lyUuIx8R6_1(.dout(w_dff_A_eT09wCdN9_1),.din(w_dff_A_lyUuIx8R6_1),.clk(gclk));
	jdff dff_A_9ZGB39M65_1(.dout(w_dff_A_lyUuIx8R6_1),.din(w_dff_A_9ZGB39M65_1),.clk(gclk));
	jdff dff_A_VkU8dekx9_1(.dout(w_dff_A_9ZGB39M65_1),.din(w_dff_A_VkU8dekx9_1),.clk(gclk));
	jdff dff_A_25R4wEmD7_1(.dout(w_dff_A_VkU8dekx9_1),.din(w_dff_A_25R4wEmD7_1),.clk(gclk));
	jdff dff_A_DVUZWOLC3_1(.dout(w_dff_A_25R4wEmD7_1),.din(w_dff_A_DVUZWOLC3_1),.clk(gclk));
	jdff dff_A_ZsvT9tFg9_1(.dout(w_n241_0[1]),.din(w_dff_A_ZsvT9tFg9_1),.clk(gclk));
	jdff dff_A_vnB3XQGd9_1(.dout(w_dff_A_ZsvT9tFg9_1),.din(w_dff_A_vnB3XQGd9_1),.clk(gclk));
	jdff dff_A_HtD9ivyS4_1(.dout(w_dff_A_vnB3XQGd9_1),.din(w_dff_A_HtD9ivyS4_1),.clk(gclk));
	jdff dff_A_X388gADN1_1(.dout(w_G195gat_1[1]),.din(w_dff_A_X388gADN1_1),.clk(gclk));
	jdff dff_A_nFZrfz888_1(.dout(w_dff_A_X388gADN1_1),.din(w_dff_A_nFZrfz888_1),.clk(gclk));
	jdff dff_A_75Z0Ttk17_1(.dout(w_dff_A_nFZrfz888_1),.din(w_dff_A_75Z0Ttk17_1),.clk(gclk));
	jdff dff_A_JkpUGZBf2_1(.dout(w_dff_A_75Z0Ttk17_1),.din(w_dff_A_JkpUGZBf2_1),.clk(gclk));
	jdff dff_A_Piy7sRBc7_1(.dout(w_dff_A_JkpUGZBf2_1),.din(w_dff_A_Piy7sRBc7_1),.clk(gclk));
	jdff dff_A_bI3C978E9_1(.dout(w_dff_A_Piy7sRBc7_1),.din(w_dff_A_bI3C978E9_1),.clk(gclk));
	jdff dff_A_DZOh1sNt7_1(.dout(w_dff_A_bI3C978E9_1),.din(w_dff_A_DZOh1sNt7_1),.clk(gclk));
	jdff dff_A_TKBNZ3Sl1_1(.dout(w_dff_A_DZOh1sNt7_1),.din(w_dff_A_TKBNZ3Sl1_1),.clk(gclk));
	jdff dff_A_oB8wX8y63_2(.dout(w_G195gat_1[2]),.din(w_dff_A_oB8wX8y63_2),.clk(gclk));
	jdff dff_A_KD6KpCBg7_2(.dout(w_dff_A_oB8wX8y63_2),.din(w_dff_A_KD6KpCBg7_2),.clk(gclk));
	jdff dff_A_TyLearqF5_2(.dout(w_dff_A_KD6KpCBg7_2),.din(w_dff_A_TyLearqF5_2),.clk(gclk));
	jdff dff_A_dHwoZXZW7_2(.dout(w_dff_A_TyLearqF5_2),.din(w_dff_A_dHwoZXZW7_2),.clk(gclk));
	jdff dff_A_GldfbQnw1_2(.dout(w_dff_A_dHwoZXZW7_2),.din(w_dff_A_GldfbQnw1_2),.clk(gclk));
	jdff dff_A_YhlLimJq7_2(.dout(w_dff_A_GldfbQnw1_2),.din(w_dff_A_YhlLimJq7_2),.clk(gclk));
	jdff dff_A_0L2Xkrqe9_2(.dout(w_dff_A_YhlLimJq7_2),.din(w_dff_A_0L2Xkrqe9_2),.clk(gclk));
	jdff dff_A_FKwPJQjV2_2(.dout(w_dff_A_0L2Xkrqe9_2),.din(w_dff_A_FKwPJQjV2_2),.clk(gclk));
	jdff dff_A_RcHTt1r62_1(.dout(w_n240_0[1]),.din(w_dff_A_RcHTt1r62_1),.clk(gclk));
	jdff dff_A_Q4NqfTz41_1(.dout(w_dff_A_RcHTt1r62_1),.din(w_dff_A_Q4NqfTz41_1),.clk(gclk));
	jdff dff_A_LfhSIsyo9_1(.dout(w_dff_A_Q4NqfTz41_1),.din(w_dff_A_LfhSIsyo9_1),.clk(gclk));
	jdff dff_A_P4zV80J80_1(.dout(w_dff_A_LfhSIsyo9_1),.din(w_dff_A_P4zV80J80_1),.clk(gclk));
	jdff dff_A_zB6Gv0j14_0(.dout(w_G121gat_0[0]),.din(w_dff_A_zB6Gv0j14_0),.clk(gclk));
	jdff dff_A_4TbRHPQ64_0(.dout(w_dff_A_zB6Gv0j14_0),.din(w_dff_A_4TbRHPQ64_0),.clk(gclk));
	jdff dff_A_K2ZbbhQx8_0(.dout(w_dff_A_4TbRHPQ64_0),.din(w_dff_A_K2ZbbhQx8_0),.clk(gclk));
	jdff dff_A_DGPwAcHs4_0(.dout(w_dff_A_K2ZbbhQx8_0),.din(w_dff_A_DGPwAcHs4_0),.clk(gclk));
	jdff dff_A_PdUsLsWK7_0(.dout(w_dff_A_DGPwAcHs4_0),.din(w_dff_A_PdUsLsWK7_0),.clk(gclk));
	jdff dff_A_2O2Q4pOl4_0(.dout(w_dff_A_PdUsLsWK7_0),.din(w_dff_A_2O2Q4pOl4_0),.clk(gclk));
	jdff dff_A_4e58sPPQ2_0(.dout(w_G195gat_2[0]),.din(w_dff_A_4e58sPPQ2_0),.clk(gclk));
	jdff dff_A_vAJMRL0o8_0(.dout(w_dff_A_4e58sPPQ2_0),.din(w_dff_A_vAJMRL0o8_0),.clk(gclk));
	jdff dff_A_e8keUhLf1_0(.dout(w_dff_A_vAJMRL0o8_0),.din(w_dff_A_e8keUhLf1_0),.clk(gclk));
	jdff dff_A_yBKCEkH24_0(.dout(w_dff_A_e8keUhLf1_0),.din(w_dff_A_yBKCEkH24_0),.clk(gclk));
	jdff dff_A_XjCVYkKl7_0(.dout(w_dff_A_yBKCEkH24_0),.din(w_dff_A_XjCVYkKl7_0),.clk(gclk));
	jdff dff_A_SKoyFyBL6_0(.dout(w_dff_A_XjCVYkKl7_0),.din(w_dff_A_SKoyFyBL6_0),.clk(gclk));
	jdff dff_A_a1EvICEe9_0(.dout(w_dff_A_SKoyFyBL6_0),.din(w_dff_A_a1EvICEe9_0),.clk(gclk));
	jdff dff_A_gzSCnwQh6_0(.dout(w_dff_A_a1EvICEe9_0),.din(w_dff_A_gzSCnwQh6_0),.clk(gclk));
	jdff dff_A_58KEmVE42_2(.dout(w_G195gat_0[2]),.din(w_dff_A_58KEmVE42_2),.clk(gclk));
	jdff dff_A_Gz0ZKhMP3_2(.dout(w_dff_A_58KEmVE42_2),.din(w_dff_A_Gz0ZKhMP3_2),.clk(gclk));
	jdff dff_A_hsRqyjQF2_2(.dout(w_dff_A_Gz0ZKhMP3_2),.din(w_dff_A_hsRqyjQF2_2),.clk(gclk));
	jdff dff_A_7I1OU8ZZ1_2(.dout(w_dff_A_hsRqyjQF2_2),.din(w_dff_A_7I1OU8ZZ1_2),.clk(gclk));
	jdff dff_A_HQIrl6Va9_1(.dout(w_n235_0[1]),.din(w_dff_A_HQIrl6Va9_1),.clk(gclk));
	jdff dff_A_T7BVjZmB1_1(.dout(w_dff_A_HQIrl6Va9_1),.din(w_dff_A_T7BVjZmB1_1),.clk(gclk));
	jdff dff_A_KorqsZZp3_1(.dout(w_dff_A_T7BVjZmB1_1),.din(w_dff_A_KorqsZZp3_1),.clk(gclk));
	jdff dff_A_KtvHNEcG6_1(.dout(w_dff_A_KorqsZZp3_1),.din(w_dff_A_KtvHNEcG6_1),.clk(gclk));
	jdff dff_A_CB2CKF6I5_1(.dout(w_dff_A_KtvHNEcG6_1),.din(w_dff_A_CB2CKF6I5_1),.clk(gclk));
	jdff dff_A_H6T3bKCf7_1(.dout(w_G189gat_1[1]),.din(w_dff_A_H6T3bKCf7_1),.clk(gclk));
	jdff dff_A_68Es0FZV4_1(.dout(w_dff_A_H6T3bKCf7_1),.din(w_dff_A_68Es0FZV4_1),.clk(gclk));
	jdff dff_A_iIdqfS259_1(.dout(w_dff_A_68Es0FZV4_1),.din(w_dff_A_iIdqfS259_1),.clk(gclk));
	jdff dff_A_mW1Fgj0O8_1(.dout(w_dff_A_iIdqfS259_1),.din(w_dff_A_mW1Fgj0O8_1),.clk(gclk));
	jdff dff_A_panc784W4_1(.dout(w_dff_A_mW1Fgj0O8_1),.din(w_dff_A_panc784W4_1),.clk(gclk));
	jdff dff_A_mkV3RWMw8_1(.dout(w_dff_A_panc784W4_1),.din(w_dff_A_mkV3RWMw8_1),.clk(gclk));
	jdff dff_A_0RWsyMFv1_1(.dout(w_dff_A_mkV3RWMw8_1),.din(w_dff_A_0RWsyMFv1_1),.clk(gclk));
	jdff dff_A_JQ4JKKZN3_1(.dout(w_dff_A_0RWsyMFv1_1),.din(w_dff_A_JQ4JKKZN3_1),.clk(gclk));
	jdff dff_A_3kGgvMV84_2(.dout(w_G189gat_1[2]),.din(w_dff_A_3kGgvMV84_2),.clk(gclk));
	jdff dff_A_gFPaDQdq1_2(.dout(w_dff_A_3kGgvMV84_2),.din(w_dff_A_gFPaDQdq1_2),.clk(gclk));
	jdff dff_A_zjrh4Zhi9_2(.dout(w_dff_A_gFPaDQdq1_2),.din(w_dff_A_zjrh4Zhi9_2),.clk(gclk));
	jdff dff_A_N1dGASNL1_2(.dout(w_dff_A_zjrh4Zhi9_2),.din(w_dff_A_N1dGASNL1_2),.clk(gclk));
	jdff dff_A_Qeh2TP0d5_2(.dout(w_dff_A_N1dGASNL1_2),.din(w_dff_A_Qeh2TP0d5_2),.clk(gclk));
	jdff dff_A_TiRiaqpM7_2(.dout(w_dff_A_Qeh2TP0d5_2),.din(w_dff_A_TiRiaqpM7_2),.clk(gclk));
	jdff dff_A_fJHNsO0G1_2(.dout(w_dff_A_TiRiaqpM7_2),.din(w_dff_A_fJHNsO0G1_2),.clk(gclk));
	jdff dff_A_BONYvIGV9_2(.dout(w_dff_A_fJHNsO0G1_2),.din(w_dff_A_BONYvIGV9_2),.clk(gclk));
	jdff dff_A_biPzaajY5_1(.dout(w_n234_0[1]),.din(w_dff_A_biPzaajY5_1),.clk(gclk));
	jdff dff_A_CdGEj5VR7_1(.dout(w_dff_A_biPzaajY5_1),.din(w_dff_A_CdGEj5VR7_1),.clk(gclk));
	jdff dff_A_xeuZn17I5_1(.dout(w_dff_A_CdGEj5VR7_1),.din(w_dff_A_xeuZn17I5_1),.clk(gclk));
	jdff dff_A_UucWkXq47_1(.dout(w_dff_A_xeuZn17I5_1),.din(w_dff_A_UucWkXq47_1),.clk(gclk));
	jdff dff_A_3lnmUeB01_1(.dout(w_dff_A_UucWkXq47_1),.din(w_dff_A_3lnmUeB01_1),.clk(gclk));
	jdff dff_A_k3roUDba9_1(.dout(w_dff_A_3lnmUeB01_1),.din(w_dff_A_k3roUDba9_1),.clk(gclk));
	jdff dff_A_RgrZBGyU8_1(.dout(w_G146gat_0[1]),.din(w_dff_A_RgrZBGyU8_1),.clk(gclk));
	jdff dff_B_43DQC57i3_2(.din(G146gat),.dout(w_dff_B_43DQC57i3_2),.clk(gclk));
	jdff dff_B_XqQFUiyg4_2(.din(w_dff_B_43DQC57i3_2),.dout(w_dff_B_XqQFUiyg4_2),.clk(gclk));
	jdff dff_B_dQhxHCWz2_2(.din(w_dff_B_XqQFUiyg4_2),.dout(w_dff_B_dQhxHCWz2_2),.clk(gclk));
	jdff dff_B_ELVxRGg83_2(.din(w_dff_B_dQhxHCWz2_2),.dout(w_dff_B_ELVxRGg83_2),.clk(gclk));
	jdff dff_A_6nBN1ogq9_1(.dout(w_G116gat_0[1]),.din(w_dff_A_6nBN1ogq9_1),.clk(gclk));
	jdff dff_A_ROKh5EhK0_1(.dout(w_dff_A_6nBN1ogq9_1),.din(w_dff_A_ROKh5EhK0_1),.clk(gclk));
	jdff dff_A_1kIFFkiw8_1(.dout(w_dff_A_ROKh5EhK0_1),.din(w_dff_A_1kIFFkiw8_1),.clk(gclk));
	jdff dff_A_gw22SdBI6_1(.dout(w_dff_A_1kIFFkiw8_1),.din(w_dff_A_gw22SdBI6_1),.clk(gclk));
	jdff dff_A_cYPOGd2v4_1(.dout(w_dff_A_gw22SdBI6_1),.din(w_dff_A_cYPOGd2v4_1),.clk(gclk));
	jdff dff_A_d6biRXab9_1(.dout(w_dff_A_cYPOGd2v4_1),.din(w_dff_A_d6biRXab9_1),.clk(gclk));
	jdff dff_A_CRKecSso3_0(.dout(w_G189gat_2[0]),.din(w_dff_A_CRKecSso3_0),.clk(gclk));
	jdff dff_A_T6ccq5hL7_0(.dout(w_dff_A_CRKecSso3_0),.din(w_dff_A_T6ccq5hL7_0),.clk(gclk));
	jdff dff_A_p5d4la7a7_0(.dout(w_dff_A_T6ccq5hL7_0),.din(w_dff_A_p5d4la7a7_0),.clk(gclk));
	jdff dff_A_J9Wi2rGg5_0(.dout(w_dff_A_p5d4la7a7_0),.din(w_dff_A_J9Wi2rGg5_0),.clk(gclk));
	jdff dff_A_Yf6uo45Z9_0(.dout(w_dff_A_J9Wi2rGg5_0),.din(w_dff_A_Yf6uo45Z9_0),.clk(gclk));
	jdff dff_A_xCZKXQlo2_0(.dout(w_dff_A_Yf6uo45Z9_0),.din(w_dff_A_xCZKXQlo2_0),.clk(gclk));
	jdff dff_A_6wM7kc4N2_0(.dout(w_dff_A_xCZKXQlo2_0),.din(w_dff_A_6wM7kc4N2_0),.clk(gclk));
	jdff dff_A_15PxcqHD1_0(.dout(w_dff_A_6wM7kc4N2_0),.din(w_dff_A_15PxcqHD1_0),.clk(gclk));
	jdff dff_A_zOXzmiA46_2(.dout(w_G189gat_0[2]),.din(w_dff_A_zOXzmiA46_2),.clk(gclk));
	jdff dff_A_ptCLX6vO7_2(.dout(w_dff_A_zOXzmiA46_2),.din(w_dff_A_ptCLX6vO7_2),.clk(gclk));
	jdff dff_A_IKVk7OZN7_2(.dout(w_dff_A_ptCLX6vO7_2),.din(w_dff_A_IKVk7OZN7_2),.clk(gclk));
	jdff dff_A_OWu9GO5M9_2(.dout(w_dff_A_IKVk7OZN7_2),.din(w_dff_A_OWu9GO5M9_2),.clk(gclk));
	jdff dff_A_EGJT6SzF8_0(.dout(w_n343_0[0]),.din(w_dff_A_EGJT6SzF8_0),.clk(gclk));
	jdff dff_A_vpcGVEZ13_0(.dout(w_dff_A_EGJT6SzF8_0),.din(w_dff_A_vpcGVEZ13_0),.clk(gclk));
	jdff dff_A_zljUsMXi2_0(.dout(w_dff_A_vpcGVEZ13_0),.din(w_dff_A_zljUsMXi2_0),.clk(gclk));
	jdff dff_A_DdnYctoD0_0(.dout(w_dff_A_zljUsMXi2_0),.din(w_dff_A_DdnYctoD0_0),.clk(gclk));
	jdff dff_A_wAhB5Dpr9_0(.dout(w_dff_A_DdnYctoD0_0),.din(w_dff_A_wAhB5Dpr9_0),.clk(gclk));
	jdff dff_A_SfACn2Ng8_0(.dout(w_dff_A_wAhB5Dpr9_0),.din(w_dff_A_SfACn2Ng8_0),.clk(gclk));
	jdff dff_B_17GVwLMI4_1(.din(n341),.dout(w_dff_B_17GVwLMI4_1),.clk(gclk));
	jdff dff_B_NXo4Vcax5_1(.din(w_dff_B_17GVwLMI4_1),.dout(w_dff_B_NXo4Vcax5_1),.clk(gclk));
	jdff dff_B_pklLYb6D2_1(.din(w_dff_B_NXo4Vcax5_1),.dout(w_dff_B_pklLYb6D2_1),.clk(gclk));
	jdff dff_B_zMH2pYu61_1(.din(w_dff_B_pklLYb6D2_1),.dout(w_dff_B_zMH2pYu61_1),.clk(gclk));
	jdff dff_B_Xnfmz8m85_1(.din(w_dff_B_zMH2pYu61_1),.dout(w_dff_B_Xnfmz8m85_1),.clk(gclk));
	jdff dff_B_IsHlgTDw1_1(.din(w_dff_B_Xnfmz8m85_1),.dout(w_dff_B_IsHlgTDw1_1),.clk(gclk));
	jdff dff_B_rYhg64yR0_1(.din(w_dff_B_IsHlgTDw1_1),.dout(w_dff_B_rYhg64yR0_1),.clk(gclk));
	jdff dff_B_THrVAbF30_1(.din(w_dff_B_rYhg64yR0_1),.dout(w_dff_B_THrVAbF30_1),.clk(gclk));
	jdff dff_A_7s7pj6yq6_1(.dout(w_n222_0[1]),.din(w_dff_A_7s7pj6yq6_1),.clk(gclk));
	jdff dff_A_4CdHw3xI2_1(.dout(w_dff_A_7s7pj6yq6_1),.din(w_dff_A_4CdHw3xI2_1),.clk(gclk));
	jdff dff_A_IKaGLcQx4_1(.dout(w_dff_A_4CdHw3xI2_1),.din(w_dff_A_IKaGLcQx4_1),.clk(gclk));
	jdff dff_A_yX7WiixN2_1(.dout(w_dff_A_IKaGLcQx4_1),.din(w_dff_A_yX7WiixN2_1),.clk(gclk));
	jdff dff_A_w0TsZFF95_1(.dout(w_dff_A_yX7WiixN2_1),.din(w_dff_A_w0TsZFF95_1),.clk(gclk));
	jdff dff_A_hFE75WfB3_1(.dout(w_dff_A_w0TsZFF95_1),.din(w_dff_A_hFE75WfB3_1),.clk(gclk));
	jdff dff_A_QCIoRFPs4_1(.dout(w_dff_A_hFE75WfB3_1),.din(w_dff_A_QCIoRFPs4_1),.clk(gclk));
	jdff dff_A_uyfWmlS52_1(.dout(w_dff_A_QCIoRFPs4_1),.din(w_dff_A_uyfWmlS52_1),.clk(gclk));
	jdff dff_A_nQJVdCYi2_0(.dout(w_n97_0[0]),.din(w_dff_A_nQJVdCYi2_0),.clk(gclk));
	jdff dff_A_QqjlHKmk1_0(.dout(w_dff_A_nQJVdCYi2_0),.din(w_dff_A_QqjlHKmk1_0),.clk(gclk));
	jdff dff_A_6GAsQtzw5_0(.dout(w_dff_A_QqjlHKmk1_0),.din(w_dff_A_6GAsQtzw5_0),.clk(gclk));
	jdff dff_A_PH8TGeuR4_1(.dout(w_G143gat_0[1]),.din(w_dff_A_PH8TGeuR4_1),.clk(gclk));
	jdff dff_B_ckQ37O4F2_2(.din(G143gat),.dout(w_dff_B_ckQ37O4F2_2),.clk(gclk));
	jdff dff_B_tJWrjoTV0_2(.din(w_dff_B_ckQ37O4F2_2),.dout(w_dff_B_tJWrjoTV0_2),.clk(gclk));
	jdff dff_B_pvufKJtW7_2(.din(w_dff_B_tJWrjoTV0_2),.dout(w_dff_B_pvufKJtW7_2),.clk(gclk));
	jdff dff_B_65QB3twe0_2(.din(w_dff_B_pvufKJtW7_2),.dout(w_dff_B_65QB3twe0_2),.clk(gclk));
	jdff dff_A_x0AiMJPD2_2(.dout(w_n148_1[2]),.din(w_dff_A_x0AiMJPD2_2),.clk(gclk));
	jdff dff_A_yVEYHzL20_2(.dout(w_dff_A_x0AiMJPD2_2),.din(w_dff_A_yVEYHzL20_2),.clk(gclk));
	jdff dff_A_zd94hS645_1(.dout(w_G111gat_0[1]),.din(w_dff_A_zd94hS645_1),.clk(gclk));
	jdff dff_A_XFB29Rx80_1(.dout(w_dff_A_zd94hS645_1),.din(w_dff_A_XFB29Rx80_1),.clk(gclk));
	jdff dff_A_0ss6Ng1O9_1(.dout(w_dff_A_XFB29Rx80_1),.din(w_dff_A_0ss6Ng1O9_1),.clk(gclk));
	jdff dff_A_z2blFpm61_1(.dout(w_dff_A_0ss6Ng1O9_1),.din(w_dff_A_z2blFpm61_1),.clk(gclk));
	jdff dff_A_bjp8xU1K8_1(.dout(w_dff_A_z2blFpm61_1),.din(w_dff_A_bjp8xU1K8_1),.clk(gclk));
	jdff dff_A_cThWVYcY6_1(.dout(w_dff_A_bjp8xU1K8_1),.din(w_dff_A_cThWVYcY6_1),.clk(gclk));
	jdff dff_A_QqaogmRE3_2(.dout(w_G183gat_0[2]),.din(w_dff_A_QqaogmRE3_2),.clk(gclk));
	jdff dff_A_gRlOYoRF9_2(.dout(w_dff_A_QqaogmRE3_2),.din(w_dff_A_gRlOYoRF9_2),.clk(gclk));
	jdff dff_A_0EMUVmRj6_2(.dout(w_dff_A_gRlOYoRF9_2),.din(w_dff_A_0EMUVmRj6_2),.clk(gclk));
	jdff dff_A_soEfiLC39_2(.dout(w_dff_A_0EMUVmRj6_2),.din(w_dff_A_soEfiLC39_2),.clk(gclk));
	jdff dff_A_RJlScyza6_2(.dout(w_dff_A_soEfiLC39_2),.din(w_dff_A_RJlScyza6_2),.clk(gclk));
	jdff dff_A_pOLLdz346_2(.dout(w_dff_A_RJlScyza6_2),.din(w_dff_A_pOLLdz346_2),.clk(gclk));
	jdff dff_A_3Cz6OzwJ3_2(.dout(w_dff_A_pOLLdz346_2),.din(w_dff_A_3Cz6OzwJ3_2),.clk(gclk));
	jdff dff_A_54e5qKsY5_2(.dout(w_dff_A_3Cz6OzwJ3_2),.din(w_dff_A_54e5qKsY5_2),.clk(gclk));
	jdff dff_A_w73sto869_0(.dout(w_n339_0[0]),.din(w_dff_A_w73sto869_0),.clk(gclk));
	jdff dff_A_pwpjSjNC8_0(.dout(w_dff_A_w73sto869_0),.din(w_dff_A_pwpjSjNC8_0),.clk(gclk));
	jdff dff_A_paMU3kcr5_0(.dout(w_dff_A_pwpjSjNC8_0),.din(w_dff_A_paMU3kcr5_0),.clk(gclk));
	jdff dff_A_DhIYGIoK8_0(.dout(w_dff_A_paMU3kcr5_0),.din(w_dff_A_DhIYGIoK8_0),.clk(gclk));
	jdff dff_A_zFIWgomP6_0(.dout(w_dff_A_DhIYGIoK8_0),.din(w_dff_A_zFIWgomP6_0),.clk(gclk));
	jdff dff_A_p742Ppg74_0(.dout(w_dff_A_zFIWgomP6_0),.din(w_dff_A_p742Ppg74_0),.clk(gclk));
	jdff dff_A_lyr1kNRw7_0(.dout(w_dff_A_p742Ppg74_0),.din(w_dff_A_lyr1kNRw7_0),.clk(gclk));
	jdff dff_B_BHrdnGlM6_1(.din(n337),.dout(w_dff_B_BHrdnGlM6_1),.clk(gclk));
	jdff dff_B_GWM0xa6L8_1(.din(w_dff_B_BHrdnGlM6_1),.dout(w_dff_B_GWM0xa6L8_1),.clk(gclk));
	jdff dff_B_T713Ti4e7_1(.din(w_dff_B_GWM0xa6L8_1),.dout(w_dff_B_T713Ti4e7_1),.clk(gclk));
	jdff dff_B_2JnXiDwJ0_1(.din(w_dff_B_T713Ti4e7_1),.dout(w_dff_B_2JnXiDwJ0_1),.clk(gclk));
	jdff dff_B_j8ejU5395_1(.din(w_dff_B_2JnXiDwJ0_1),.dout(w_dff_B_j8ejU5395_1),.clk(gclk));
	jdff dff_B_1BnI7T5Q0_1(.din(w_dff_B_j8ejU5395_1),.dout(w_dff_B_1BnI7T5Q0_1),.clk(gclk));
	jdff dff_B_TBWOYx9H7_1(.din(w_dff_B_1BnI7T5Q0_1),.dout(w_dff_B_TBWOYx9H7_1),.clk(gclk));
	jdff dff_B_GQdyiRzL9_1(.din(w_dff_B_TBWOYx9H7_1),.dout(w_dff_B_GQdyiRzL9_1),.clk(gclk));
	jdff dff_B_zRWcyhoV2_1(.din(w_dff_B_GQdyiRzL9_1),.dout(w_dff_B_zRWcyhoV2_1),.clk(gclk));
	jdff dff_A_iaarpLbz1_2(.dout(w_n336_0[2]),.din(w_dff_A_iaarpLbz1_2),.clk(gclk));
	jdff dff_A_aeWtvHSd9_2(.dout(w_dff_A_iaarpLbz1_2),.din(w_dff_A_aeWtvHSd9_2),.clk(gclk));
	jdff dff_A_siMNGYZJ1_2(.dout(w_dff_A_aeWtvHSd9_2),.din(w_dff_A_siMNGYZJ1_2),.clk(gclk));
	jdff dff_A_szMHMi966_2(.dout(w_dff_A_siMNGYZJ1_2),.din(w_dff_A_szMHMi966_2),.clk(gclk));
	jdff dff_A_j8R3cMdQ2_2(.dout(w_dff_A_szMHMi966_2),.din(w_dff_A_j8R3cMdQ2_2),.clk(gclk));
	jdff dff_A_DPPJxwXO3_2(.dout(w_dff_A_j8R3cMdQ2_2),.din(w_dff_A_DPPJxwXO3_2),.clk(gclk));
	jdff dff_A_qyfsu4mV1_2(.dout(w_dff_A_DPPJxwXO3_2),.din(w_dff_A_qyfsu4mV1_2),.clk(gclk));
	jdff dff_A_wzlfTpSR4_2(.dout(w_dff_A_qyfsu4mV1_2),.din(w_dff_A_wzlfTpSR4_2),.clk(gclk));
	jdff dff_A_SexcC3WA1_2(.dout(w_dff_A_wzlfTpSR4_2),.din(w_dff_A_SexcC3WA1_2),.clk(gclk));
	jdff dff_B_6GSYaz0e9_0(.din(n333),.dout(w_dff_B_6GSYaz0e9_0),.clk(gclk));
	jdff dff_B_XR90HrZC3_0(.din(n332),.dout(w_dff_B_XR90HrZC3_0),.clk(gclk));
	jdff dff_B_eOwpGUK18_0(.din(w_dff_B_XR90HrZC3_0),.dout(w_dff_B_eOwpGUK18_0),.clk(gclk));
	jdff dff_B_4eSsaiJV7_0(.din(w_dff_B_eOwpGUK18_0),.dout(w_dff_B_4eSsaiJV7_0),.clk(gclk));
	jdff dff_B_Kn1FYWoV5_0(.din(w_dff_B_4eSsaiJV7_0),.dout(w_dff_B_Kn1FYWoV5_0),.clk(gclk));
	jdff dff_A_X3qLaOM47_0(.dout(w_G153gat_0[0]),.din(w_dff_A_X3qLaOM47_0),.clk(gclk));
	jdff dff_A_2meL8y736_0(.dout(w_dff_A_X3qLaOM47_0),.din(w_dff_A_2meL8y736_0),.clk(gclk));
	jdff dff_A_64HgHN3Q9_0(.dout(w_dff_A_2meL8y736_0),.din(w_dff_A_64HgHN3Q9_0),.clk(gclk));
	jdff dff_A_fWbf8oFC2_0(.dout(w_dff_A_64HgHN3Q9_0),.din(w_dff_A_fWbf8oFC2_0),.clk(gclk));
	jdff dff_A_1tJh7omA6_2(.dout(w_G153gat_0[2]),.din(w_dff_A_1tJh7omA6_2),.clk(gclk));
	jdff dff_A_wqRgMnMr2_2(.dout(w_dff_A_1tJh7omA6_2),.din(w_dff_A_wqRgMnMr2_2),.clk(gclk));
	jdff dff_A_cKVQ8j5j7_2(.dout(w_dff_A_wqRgMnMr2_2),.din(w_dff_A_cKVQ8j5j7_2),.clk(gclk));
	jdff dff_A_1Sr3NbGH3_2(.dout(w_dff_A_cKVQ8j5j7_2),.din(w_dff_A_1Sr3NbGH3_2),.clk(gclk));
	jdff dff_A_kiWkekqw1_2(.dout(w_dff_A_1Sr3NbGH3_2),.din(w_dff_A_kiWkekqw1_2),.clk(gclk));
	jdff dff_A_CUbpgPGn2_0(.dout(w_G106gat_0[0]),.din(w_dff_A_CUbpgPGn2_0),.clk(gclk));
	jdff dff_A_s3zAHzsd5_0(.dout(w_dff_A_CUbpgPGn2_0),.din(w_dff_A_s3zAHzsd5_0),.clk(gclk));
	jdff dff_A_eB2W1GEJ3_0(.dout(w_dff_A_s3zAHzsd5_0),.din(w_dff_A_eB2W1GEJ3_0),.clk(gclk));
	jdff dff_A_c2a3JZsZ6_0(.dout(w_dff_A_eB2W1GEJ3_0),.din(w_dff_A_c2a3JZsZ6_0),.clk(gclk));
	jdff dff_A_6EYbj9qD5_0(.dout(w_dff_A_c2a3JZsZ6_0),.din(w_dff_A_6EYbj9qD5_0),.clk(gclk));
	jdff dff_A_URmQRko84_0(.dout(w_dff_A_6EYbj9qD5_0),.din(w_dff_A_URmQRko84_0),.clk(gclk));
	jdff dff_A_jwCTRDKo0_1(.dout(w_G177gat_1[1]),.din(w_dff_A_jwCTRDKo0_1),.clk(gclk));
	jdff dff_A_KHqIG8Ny1_1(.dout(w_dff_A_jwCTRDKo0_1),.din(w_dff_A_KHqIG8Ny1_1),.clk(gclk));
	jdff dff_A_l7HuiG969_1(.dout(w_dff_A_KHqIG8Ny1_1),.din(w_dff_A_l7HuiG969_1),.clk(gclk));
	jdff dff_A_1Tv02Wh29_1(.dout(w_dff_A_l7HuiG969_1),.din(w_dff_A_1Tv02Wh29_1),.clk(gclk));
	jdff dff_A_HJjv8p6k1_1(.dout(w_dff_A_1Tv02Wh29_1),.din(w_dff_A_HJjv8p6k1_1),.clk(gclk));
	jdff dff_A_5rAKIP7Z4_1(.dout(w_dff_A_HJjv8p6k1_1),.din(w_dff_A_5rAKIP7Z4_1),.clk(gclk));
	jdff dff_A_eAq0ZszF3_1(.dout(w_dff_A_5rAKIP7Z4_1),.din(w_dff_A_eAq0ZszF3_1),.clk(gclk));
	jdff dff_A_Tfb3Se8u8_1(.dout(w_dff_A_eAq0ZszF3_1),.din(w_dff_A_Tfb3Se8u8_1),.clk(gclk));
	jdff dff_A_NT7xUXH68_1(.dout(w_dff_A_Tfb3Se8u8_1),.din(w_dff_A_NT7xUXH68_1),.clk(gclk));
	jdff dff_A_ST8w2acz9_1(.dout(w_G177gat_0[1]),.din(w_dff_A_ST8w2acz9_1),.clk(gclk));
	jdff dff_A_Zlcc1WBo6_1(.dout(w_dff_A_ST8w2acz9_1),.din(w_dff_A_Zlcc1WBo6_1),.clk(gclk));
	jdff dff_A_R26fKNaK3_1(.dout(w_dff_A_Zlcc1WBo6_1),.din(w_dff_A_R26fKNaK3_1),.clk(gclk));
	jdff dff_A_VewlEDL70_1(.dout(w_dff_A_R26fKNaK3_1),.din(w_dff_A_VewlEDL70_1),.clk(gclk));
	jdff dff_A_yyUdDatr8_2(.dout(w_G177gat_0[2]),.din(w_dff_A_yyUdDatr8_2),.clk(gclk));
	jdff dff_A_KgHjpYpx2_2(.dout(w_dff_A_yyUdDatr8_2),.din(w_dff_A_KgHjpYpx2_2),.clk(gclk));
	jdff dff_A_WLRj8K4X0_2(.dout(w_dff_A_KgHjpYpx2_2),.din(w_dff_A_WLRj8K4X0_2),.clk(gclk));
	jdff dff_A_h308vyhu8_2(.dout(w_dff_A_WLRj8K4X0_2),.din(w_dff_A_h308vyhu8_2),.clk(gclk));
	jdff dff_A_j7fqDAxq3_2(.dout(w_dff_A_h308vyhu8_2),.din(w_dff_A_j7fqDAxq3_2),.clk(gclk));
	jdff dff_A_C8L4BNUS5_2(.dout(w_dff_A_j7fqDAxq3_2),.din(w_dff_A_C8L4BNUS5_2),.clk(gclk));
	jdff dff_A_nYV1IXK00_2(.dout(w_dff_A_C8L4BNUS5_2),.din(w_dff_A_nYV1IXK00_2),.clk(gclk));
	jdff dff_A_sX7oZQmF4_2(.dout(w_dff_A_nYV1IXK00_2),.din(w_dff_A_sX7oZQmF4_2),.clk(gclk));
	jdff dff_A_eyk3KoDE9_2(.dout(w_dff_A_sX7oZQmF4_2),.din(w_dff_A_eyk3KoDE9_2),.clk(gclk));
	jdff dff_B_9BWndEVS6_1(.din(n419),.dout(w_dff_B_9BWndEVS6_1),.clk(gclk));
	jdff dff_B_JDVZwhDt8_0(.din(n424),.dout(w_dff_B_JDVZwhDt8_0),.clk(gclk));
	jdff dff_B_guRjmfLS2_0(.din(w_dff_B_JDVZwhDt8_0),.dout(w_dff_B_guRjmfLS2_0),.clk(gclk));
	jdff dff_A_YoFWnBwt3_0(.dout(w_G246gat_0[0]),.din(w_dff_A_YoFWnBwt3_0),.clk(gclk));
	jdff dff_A_d1HhWs9R1_0(.dout(w_dff_A_YoFWnBwt3_0),.din(w_dff_A_d1HhWs9R1_0),.clk(gclk));
	jdff dff_A_jYjxtVsY3_0(.dout(w_dff_A_d1HhWs9R1_0),.din(w_dff_A_jYjxtVsY3_0),.clk(gclk));
	jdff dff_A_fIGaozpt2_0(.dout(w_dff_A_jYjxtVsY3_0),.din(w_dff_A_fIGaozpt2_0),.clk(gclk));
	jdff dff_A_sv7ef6nn8_0(.dout(w_dff_A_fIGaozpt2_0),.din(w_dff_A_sv7ef6nn8_0),.clk(gclk));
	jdff dff_A_uvliav676_0(.dout(w_dff_A_sv7ef6nn8_0),.din(w_dff_A_uvliav676_0),.clk(gclk));
	jdff dff_A_Bm7VBKl85_0(.dout(w_dff_A_uvliav676_0),.din(w_dff_A_Bm7VBKl85_0),.clk(gclk));
	jdff dff_A_pRmQpTHG9_0(.dout(w_dff_A_Bm7VBKl85_0),.din(w_dff_A_pRmQpTHG9_0),.clk(gclk));
	jdff dff_A_v2wpW7I60_2(.dout(w_G246gat_0[2]),.din(w_dff_A_v2wpW7I60_2),.clk(gclk));
	jdff dff_A_HYAAvPMU0_2(.dout(w_dff_A_v2wpW7I60_2),.din(w_dff_A_HYAAvPMU0_2),.clk(gclk));
	jdff dff_A_q812jhGF1_2(.dout(w_dff_A_HYAAvPMU0_2),.din(w_dff_A_q812jhGF1_2),.clk(gclk));
	jdff dff_A_wYIuQO3E2_2(.dout(w_dff_A_q812jhGF1_2),.din(w_dff_A_wYIuQO3E2_2),.clk(gclk));
	jdff dff_A_6yWhX6pT4_2(.dout(w_dff_A_wYIuQO3E2_2),.din(w_dff_A_6yWhX6pT4_2),.clk(gclk));
	jdff dff_A_8823zXGq1_2(.dout(w_dff_A_6yWhX6pT4_2),.din(w_dff_A_8823zXGq1_2),.clk(gclk));
	jdff dff_A_zoxLnd2T6_2(.dout(w_dff_A_8823zXGq1_2),.din(w_dff_A_zoxLnd2T6_2),.clk(gclk));
	jdff dff_B_FbsYManE5_3(.din(G246gat),.dout(w_dff_B_FbsYManE5_3),.clk(gclk));
	jdff dff_B_tPbzwCid2_0(.din(n422),.dout(w_dff_B_tPbzwCid2_0),.clk(gclk));
	jdff dff_B_DkZqUcE39_0(.din(w_dff_B_tPbzwCid2_0),.dout(w_dff_B_DkZqUcE39_0),.clk(gclk));
	jdff dff_B_iyOm5jen4_0(.din(w_dff_B_DkZqUcE39_0),.dout(w_dff_B_iyOm5jen4_0),.clk(gclk));
	jdff dff_B_fJz966m29_0(.din(w_dff_B_iyOm5jen4_0),.dout(w_dff_B_fJz966m29_0),.clk(gclk));
	jdff dff_B_0xpvP6Sy8_0(.din(w_dff_B_fJz966m29_0),.dout(w_dff_B_0xpvP6Sy8_0),.clk(gclk));
	jdff dff_B_yzzNuLNe8_0(.din(w_dff_B_0xpvP6Sy8_0),.dout(w_dff_B_yzzNuLNe8_0),.clk(gclk));
	jdff dff_B_auaD2fl65_0(.din(w_dff_B_yzzNuLNe8_0),.dout(w_dff_B_auaD2fl65_0),.clk(gclk));
	jdff dff_B_HS5mRapg2_0(.din(w_dff_B_auaD2fl65_0),.dout(w_dff_B_HS5mRapg2_0),.clk(gclk));
	jdff dff_B_spCLzmLV8_0(.din(w_dff_B_HS5mRapg2_0),.dout(w_dff_B_spCLzmLV8_0),.clk(gclk));
	jdff dff_B_q5Ktwy8s3_0(.din(w_dff_B_spCLzmLV8_0),.dout(w_dff_B_q5Ktwy8s3_0),.clk(gclk));
	jdff dff_A_SqO57Zob2_1(.dout(w_G96gat_0[1]),.din(w_dff_A_SqO57Zob2_1),.clk(gclk));
	jdff dff_A_sCOXXYkL6_1(.dout(w_dff_A_SqO57Zob2_1),.din(w_dff_A_sCOXXYkL6_1),.clk(gclk));
	jdff dff_A_JhEi1HTD5_1(.dout(w_dff_A_sCOXXYkL6_1),.din(w_dff_A_JhEi1HTD5_1),.clk(gclk));
	jdff dff_A_ENmqCqTt3_1(.dout(w_dff_A_JhEi1HTD5_1),.din(w_dff_A_ENmqCqTt3_1),.clk(gclk));
	jdff dff_A_6TrxxOM32_1(.dout(w_dff_A_ENmqCqTt3_1),.din(w_dff_A_6TrxxOM32_1),.clk(gclk));
	jdff dff_A_i58d2qx50_1(.dout(w_dff_A_6TrxxOM32_1),.din(w_dff_A_i58d2qx50_1),.clk(gclk));
	jdff dff_A_WBLbT3Mu9_0(.dout(w_n420_0[0]),.din(w_dff_A_WBLbT3Mu9_0),.clk(gclk));
	jdff dff_A_3b3TYrUP1_0(.dout(w_dff_A_WBLbT3Mu9_0),.din(w_dff_A_3b3TYrUP1_0),.clk(gclk));
	jdff dff_A_jiIgGLHY5_0(.dout(w_dff_A_3b3TYrUP1_0),.din(w_dff_A_jiIgGLHY5_0),.clk(gclk));
	jdff dff_A_CjbDfE3e9_0(.dout(w_dff_A_jiIgGLHY5_0),.din(w_dff_A_CjbDfE3e9_0),.clk(gclk));
	jdff dff_A_cODPshmq1_0(.dout(w_dff_A_CjbDfE3e9_0),.din(w_dff_A_cODPshmq1_0),.clk(gclk));
	jdff dff_A_JDBYFYWt7_0(.dout(w_dff_A_cODPshmq1_0),.din(w_dff_A_JDBYFYWt7_0),.clk(gclk));
	jdff dff_A_e6nOEHk31_0(.dout(w_dff_A_JDBYFYWt7_0),.din(w_dff_A_e6nOEHk31_0),.clk(gclk));
	jdff dff_A_HOXSNJxj9_0(.dout(w_dff_A_e6nOEHk31_0),.din(w_dff_A_HOXSNJxj9_0),.clk(gclk));
	jdff dff_A_oeP4XS5h4_0(.dout(w_dff_A_HOXSNJxj9_0),.din(w_dff_A_oeP4XS5h4_0),.clk(gclk));
	jdff dff_A_H1gPzLXb4_0(.dout(w_dff_A_oeP4XS5h4_0),.din(w_dff_A_H1gPzLXb4_0),.clk(gclk));
	jdff dff_A_HlfwhfIe3_0(.dout(w_G228gat_0[0]),.din(w_dff_A_HlfwhfIe3_0),.clk(gclk));
	jdff dff_B_WkQ1Z08U2_3(.din(G228gat),.dout(w_dff_B_WkQ1Z08U2_3),.clk(gclk));
	jdff dff_B_yj19BfzW4_3(.din(w_dff_B_WkQ1Z08U2_3),.dout(w_dff_B_yj19BfzW4_3),.clk(gclk));
	jdff dff_B_jcyjnR323_3(.din(w_dff_B_yj19BfzW4_3),.dout(w_dff_B_jcyjnR323_3),.clk(gclk));
	jdff dff_B_9P6gXs5P0_3(.din(w_dff_B_jcyjnR323_3),.dout(w_dff_B_9P6gXs5P0_3),.clk(gclk));
	jdff dff_B_Jlkm723F3_3(.din(w_dff_B_9P6gXs5P0_3),.dout(w_dff_B_Jlkm723F3_3),.clk(gclk));
	jdff dff_B_vFDnUJ2v2_3(.din(w_dff_B_Jlkm723F3_3),.dout(w_dff_B_vFDnUJ2v2_3),.clk(gclk));
	jdff dff_B_aw3uN2ng6_3(.din(w_dff_B_vFDnUJ2v2_3),.dout(w_dff_B_aw3uN2ng6_3),.clk(gclk));
	jdff dff_B_MkHlyEnr7_3(.din(w_dff_B_aw3uN2ng6_3),.dout(w_dff_B_MkHlyEnr7_3),.clk(gclk));
	jdff dff_B_QR0EmBkX8_3(.din(w_dff_B_MkHlyEnr7_3),.dout(w_dff_B_QR0EmBkX8_3),.clk(gclk));
	jdff dff_B_s45QQpiD1_0(.din(n325),.dout(w_dff_B_s45QQpiD1_0),.clk(gclk));
	jdff dff_B_Uv6o4uxD1_0(.din(n324),.dout(w_dff_B_Uv6o4uxD1_0),.clk(gclk));
	jdff dff_B_ZJXg71DB7_0(.din(w_dff_B_Uv6o4uxD1_0),.dout(w_dff_B_ZJXg71DB7_0),.clk(gclk));
	jdff dff_B_nqHDBrNL8_0(.din(w_dff_B_ZJXg71DB7_0),.dout(w_dff_B_nqHDBrNL8_0),.clk(gclk));
	jdff dff_B_QzdtIJtd4_0(.din(w_dff_B_nqHDBrNL8_0),.dout(w_dff_B_QzdtIJtd4_0),.clk(gclk));
	jdff dff_A_VIBDWbqU0_1(.dout(w_G149gat_0[1]),.din(w_dff_A_VIBDWbqU0_1),.clk(gclk));
	jdff dff_B_jGyfQp2c6_2(.din(G149gat),.dout(w_dff_B_jGyfQp2c6_2),.clk(gclk));
	jdff dff_B_aJ6kLBXZ2_2(.din(w_dff_B_jGyfQp2c6_2),.dout(w_dff_B_aJ6kLBXZ2_2),.clk(gclk));
	jdff dff_B_ZvYqvzJP6_2(.din(w_dff_B_aJ6kLBXZ2_2),.dout(w_dff_B_ZvYqvzJP6_2),.clk(gclk));
	jdff dff_B_rozhVQNP3_2(.din(w_dff_B_ZvYqvzJP6_2),.dout(w_dff_B_rozhVQNP3_2),.clk(gclk));
	jdff dff_A_3dL30TBv8_0(.dout(w_n162_0[0]),.din(w_dff_A_3dL30TBv8_0),.clk(gclk));
	jdff dff_B_XXbV3zQw3_1(.din(n157),.dout(w_dff_B_XXbV3zQw3_1),.clk(gclk));
	jdff dff_B_hMdlKyK58_1(.din(n150),.dout(w_dff_B_hMdlKyK58_1),.clk(gclk));
	jdff dff_A_cSLTPijy3_0(.dout(w_n152_0[0]),.din(w_dff_A_cSLTPijy3_0),.clk(gclk));
	jdff dff_A_srPCK7nJ5_0(.dout(w_n151_0[0]),.din(w_dff_A_srPCK7nJ5_0),.clk(gclk));
	jdff dff_B_Yh1MOgGx9_2(.din(n151),.dout(w_dff_B_Yh1MOgGx9_2),.clk(gclk));
	jdff dff_A_O39kA17A9_0(.dout(w_n149_0[0]),.din(w_dff_A_O39kA17A9_0),.clk(gclk));
	jdff dff_A_H2GZtF6F1_0(.dout(w_dff_A_O39kA17A9_0),.din(w_dff_A_H2GZtF6F1_0),.clk(gclk));
	jdff dff_A_FcRWR8m76_1(.dout(w_n111_0[1]),.din(w_dff_A_FcRWR8m76_1),.clk(gclk));
	jdff dff_A_7Xsqoc8r5_0(.dout(w_G42gat_1[0]),.din(w_dff_A_7Xsqoc8r5_0),.clk(gclk));
	jdff dff_A_vFzjVfJl1_0(.dout(w_n95_0[0]),.din(w_dff_A_vFzjVfJl1_0),.clk(gclk));
	jdff dff_A_CJ6pJ0Sd6_0(.dout(w_dff_A_vFzjVfJl1_0),.din(w_dff_A_CJ6pJ0Sd6_0),.clk(gclk));
	jdff dff_A_883qTqWJ8_0(.dout(w_dff_A_CJ6pJ0Sd6_0),.din(w_dff_A_883qTqWJ8_0),.clk(gclk));
	jdff dff_A_RYpoHz774_2(.dout(w_n95_0[2]),.din(w_dff_A_RYpoHz774_2),.clk(gclk));
	jdff dff_A_SWS8zYQ67_2(.dout(w_dff_A_RYpoHz774_2),.din(w_dff_A_SWS8zYQ67_2),.clk(gclk));
	jdff dff_A_BJqiOklz3_2(.dout(w_G17gat_2[2]),.din(w_dff_A_BJqiOklz3_2),.clk(gclk));
	jdff dff_A_uzkzW8UG4_2(.dout(w_dff_A_BJqiOklz3_2),.din(w_dff_A_uzkzW8UG4_2),.clk(gclk));
	jdff dff_A_QNvHU31e7_1(.dout(w_G101gat_0[1]),.din(w_dff_A_QNvHU31e7_1),.clk(gclk));
	jdff dff_A_Q8n0dWw79_1(.dout(w_dff_A_QNvHU31e7_1),.din(w_dff_A_Q8n0dWw79_1),.clk(gclk));
	jdff dff_A_7H4wQV9e9_1(.dout(w_dff_A_Q8n0dWw79_1),.din(w_dff_A_7H4wQV9e9_1),.clk(gclk));
	jdff dff_A_T9ZOG8LW8_1(.dout(w_dff_A_7H4wQV9e9_1),.din(w_dff_A_T9ZOG8LW8_1),.clk(gclk));
	jdff dff_A_AsnBQUSc1_1(.dout(w_dff_A_T9ZOG8LW8_1),.din(w_dff_A_AsnBQUSc1_1),.clk(gclk));
	jdff dff_A_Kq8CvxTw7_1(.dout(w_dff_A_AsnBQUSc1_1),.din(w_dff_A_Kq8CvxTw7_1),.clk(gclk));
	jdff dff_A_tmgnPL9s8_1(.dout(w_n306_0[1]),.din(w_dff_A_tmgnPL9s8_1),.clk(gclk));
	jdff dff_A_WZEDCsWq4_1(.dout(w_dff_A_tmgnPL9s8_1),.din(w_dff_A_WZEDCsWq4_1),.clk(gclk));
	jdff dff_A_bYVKdZ3g4_2(.dout(w_n306_0[2]),.din(w_dff_A_bYVKdZ3g4_2),.clk(gclk));
	jdff dff_A_vg7FDJnQ3_2(.dout(w_dff_A_bYVKdZ3g4_2),.din(w_dff_A_vg7FDJnQ3_2),.clk(gclk));
	jdff dff_A_QRFb94mw6_2(.dout(w_G447gat_0[2]),.din(w_dff_A_QRFb94mw6_2),.clk(gclk));
	jdff dff_A_udxixTEL4_1(.dout(w_G51gat_1[1]),.din(w_dff_A_udxixTEL4_1),.clk(gclk));
	jdff dff_A_qjh96vI27_0(.dout(w_G80gat_0[0]),.din(w_dff_A_qjh96vI27_0),.clk(gclk));
	jdff dff_A_fzqXj6HD0_0(.dout(w_dff_A_qjh96vI27_0),.din(w_dff_A_fzqXj6HD0_0),.clk(gclk));
	jdff dff_A_gsqSXBtL6_2(.dout(w_G80gat_0[2]),.din(w_dff_A_gsqSXBtL6_2),.clk(gclk));
	jdff dff_A_inIXd7Eh8_0(.dout(w_n86_0[0]),.din(w_dff_A_inIXd7Eh8_0),.clk(gclk));
	jdff dff_A_ChJmihjf4_0(.dout(w_dff_A_inIXd7Eh8_0),.din(w_dff_A_ChJmihjf4_0),.clk(gclk));
	jdff dff_A_eFGwfiAL1_0(.dout(w_G29gat_0[0]),.din(w_dff_A_eFGwfiAL1_0),.clk(gclk));
	jdff dff_A_WzQeFSph6_0(.dout(w_dff_A_eFGwfiAL1_0),.din(w_dff_A_WzQeFSph6_0),.clk(gclk));
	jdff dff_A_6lqp49I31_0(.dout(w_dff_A_WzQeFSph6_0),.din(w_dff_A_6lqp49I31_0),.clk(gclk));
	jdff dff_A_d0pgtZvo9_0(.dout(w_G17gat_1[0]),.din(w_dff_A_d0pgtZvo9_0),.clk(gclk));
	jdff dff_A_6a7MvcJ44_0(.dout(w_dff_A_d0pgtZvo9_0),.din(w_dff_A_6a7MvcJ44_0),.clk(gclk));
	jdff dff_A_47CLtQ8n0_0(.dout(w_dff_A_6a7MvcJ44_0),.din(w_dff_A_47CLtQ8n0_0),.clk(gclk));
	jdff dff_A_pLKY32TV0_0(.dout(w_dff_A_47CLtQ8n0_0),.din(w_dff_A_pLKY32TV0_0),.clk(gclk));
	jdff dff_A_9QSAiuJY3_1(.dout(w_G17gat_1[1]),.din(w_dff_A_9QSAiuJY3_1),.clk(gclk));
	jdff dff_A_hAcwclaT7_1(.dout(w_dff_A_9QSAiuJY3_1),.din(w_dff_A_hAcwclaT7_1),.clk(gclk));
	jdff dff_A_tABhtonR0_1(.dout(w_dff_A_hAcwclaT7_1),.din(w_dff_A_tABhtonR0_1),.clk(gclk));
	jdff dff_B_bGky21ci8_2(.din(n144),.dout(w_dff_B_bGky21ci8_2),.clk(gclk));
	jdff dff_B_ZRqV7zKa0_2(.din(w_dff_B_bGky21ci8_2),.dout(w_dff_B_ZRqV7zKa0_2),.clk(gclk));
	jdff dff_B_hXi4GvvB5_2(.din(w_dff_B_ZRqV7zKa0_2),.dout(w_dff_B_hXi4GvvB5_2),.clk(gclk));
	jdff dff_B_kzHPPf338_2(.din(w_dff_B_hXi4GvvB5_2),.dout(w_dff_B_kzHPPf338_2),.clk(gclk));
	jdff dff_A_ur5K87AI0_0(.dout(w_G237gat_0[0]),.din(w_dff_A_ur5K87AI0_0),.clk(gclk));
	jdff dff_A_oFPbvM8S9_0(.dout(w_dff_A_ur5K87AI0_0),.din(w_dff_A_oFPbvM8S9_0),.clk(gclk));
	jdff dff_A_6s5JWaOQ9_0(.dout(w_dff_A_oFPbvM8S9_0),.din(w_dff_A_6s5JWaOQ9_0),.clk(gclk));
	jdff dff_A_FQ3gAwJT5_0(.dout(w_dff_A_6s5JWaOQ9_0),.din(w_dff_A_FQ3gAwJT5_0),.clk(gclk));
	jdff dff_A_1lCmjEwm4_0(.dout(w_dff_A_FQ3gAwJT5_0),.din(w_dff_A_1lCmjEwm4_0),.clk(gclk));
	jdff dff_A_KpHEoisX1_0(.dout(w_dff_A_1lCmjEwm4_0),.din(w_dff_A_KpHEoisX1_0),.clk(gclk));
	jdff dff_A_2PZPIQRa0_0(.dout(w_dff_A_KpHEoisX1_0),.din(w_dff_A_2PZPIQRa0_0),.clk(gclk));
	jdff dff_A_H81VmuLa9_0(.dout(w_dff_A_2PZPIQRa0_0),.din(w_dff_A_H81VmuLa9_0),.clk(gclk));
	jdff dff_A_JCmb31hf1_0(.dout(w_dff_A_H81VmuLa9_0),.din(w_dff_A_JCmb31hf1_0),.clk(gclk));
	jdff dff_A_4fkzmxwA3_2(.dout(w_G237gat_0[2]),.din(w_dff_A_4fkzmxwA3_2),.clk(gclk));
	jdff dff_A_0cSXR2PC0_2(.dout(w_dff_A_4fkzmxwA3_2),.din(w_dff_A_0cSXR2PC0_2),.clk(gclk));
	jdff dff_A_UmHC5iqM7_2(.dout(w_dff_A_0cSXR2PC0_2),.din(w_dff_A_UmHC5iqM7_2),.clk(gclk));
	jdff dff_A_epP6TRl44_2(.dout(w_dff_A_UmHC5iqM7_2),.din(w_dff_A_epP6TRl44_2),.clk(gclk));
	jdff dff_A_yZveYZra3_2(.dout(w_dff_A_epP6TRl44_2),.din(w_dff_A_yZveYZra3_2),.clk(gclk));
	jdff dff_A_KkiWDRZQ4_2(.dout(w_dff_A_yZveYZra3_2),.din(w_dff_A_KkiWDRZQ4_2),.clk(gclk));
	jdff dff_A_xjav24r93_2(.dout(w_dff_A_KkiWDRZQ4_2),.din(w_dff_A_xjav24r93_2),.clk(gclk));
	jdff dff_A_xjJ1q6HZ2_2(.dout(w_dff_A_xjav24r93_2),.din(w_dff_A_xjJ1q6HZ2_2),.clk(gclk));
	jdff dff_A_5Xt0KupC1_2(.dout(w_dff_A_xjJ1q6HZ2_2),.din(w_dff_A_5Xt0KupC1_2),.clk(gclk));
	jdff dff_A_BANckRck8_0(.dout(w_n178_0[0]),.din(w_dff_A_BANckRck8_0),.clk(gclk));
	jdff dff_A_kXUfKTBt6_0(.dout(w_dff_A_BANckRck8_0),.din(w_dff_A_kXUfKTBt6_0),.clk(gclk));
	jdff dff_A_hZhmGr6N0_0(.dout(w_dff_A_kXUfKTBt6_0),.din(w_dff_A_hZhmGr6N0_0),.clk(gclk));
	jdff dff_A_yKn7Acjc5_0(.dout(w_dff_A_hZhmGr6N0_0),.din(w_dff_A_yKn7Acjc5_0),.clk(gclk));
	jdff dff_A_QnxKz3Rl1_0(.dout(w_dff_A_yKn7Acjc5_0),.din(w_dff_A_QnxKz3Rl1_0),.clk(gclk));
	jdff dff_A_nABzgguu0_0(.dout(w_dff_A_QnxKz3Rl1_0),.din(w_dff_A_nABzgguu0_0),.clk(gclk));
	jdff dff_B_neQ6GObu2_0(.din(n176),.dout(w_dff_B_neQ6GObu2_0),.clk(gclk));
	jdff dff_A_qGEjEI2b9_1(.dout(w_n122_0[1]),.din(w_dff_A_qGEjEI2b9_1),.clk(gclk));
	jdff dff_A_bQ1HpIsw9_1(.dout(w_dff_A_qGEjEI2b9_1),.din(w_dff_A_bQ1HpIsw9_1),.clk(gclk));
	jdff dff_A_QqoOc1Jz9_1(.dout(w_dff_A_bQ1HpIsw9_1),.din(w_dff_A_QqoOc1Jz9_1),.clk(gclk));
	jdff dff_A_1bJBU0Ea0_1(.dout(w_G68gat_0[1]),.din(w_dff_A_1bJBU0Ea0_1),.clk(gclk));
	jdff dff_A_CJN7BoNr6_1(.dout(w_dff_A_1bJBU0Ea0_1),.din(w_dff_A_CJN7BoNr6_1),.clk(gclk));
	jdff dff_A_fOOkhVnI6_1(.dout(w_dff_A_CJN7BoNr6_1),.din(w_dff_A_fOOkhVnI6_1),.clk(gclk));
	jdff dff_A_dADlnIYC6_1(.dout(w_dff_A_fOOkhVnI6_1),.din(w_dff_A_dADlnIYC6_1),.clk(gclk));
	jdff dff_A_fVb50uyJ6_1(.dout(w_G42gat_0[1]),.din(w_dff_A_fVb50uyJ6_1),.clk(gclk));
	jdff dff_A_FaerhiMT4_2(.dout(w_G42gat_0[2]),.din(w_dff_A_FaerhiMT4_2),.clk(gclk));
	jdff dff_A_T7TLZoUt2_1(.dout(w_G1gat_0[1]),.din(w_dff_A_T7TLZoUt2_1),.clk(gclk));
	jdff dff_A_qO7i5XFD5_1(.dout(w_dff_A_T7TLZoUt2_1),.din(w_dff_A_qO7i5XFD5_1),.clk(gclk));
	jdff dff_A_y1OnYwrt7_1(.dout(w_dff_A_qO7i5XFD5_1),.din(w_dff_A_y1OnYwrt7_1),.clk(gclk));
	jdff dff_A_Xok89pFc6_1(.dout(w_dff_A_y1OnYwrt7_1),.din(w_dff_A_Xok89pFc6_1),.clk(gclk));
	jdff dff_A_Lst0McxJ1_1(.dout(w_dff_A_Xok89pFc6_1),.din(w_dff_A_Lst0McxJ1_1),.clk(gclk));
	jdff dff_A_QxIfccYM2_1(.dout(w_G13gat_0[1]),.din(w_dff_A_QxIfccYM2_1),.clk(gclk));
	jdff dff_A_egK1zrPp8_0(.dout(w_G55gat_0[0]),.din(w_dff_A_egK1zrPp8_0),.clk(gclk));
	jdff dff_A_rW7uXXy70_1(.dout(w_G55gat_0[1]),.din(w_dff_A_rW7uXXy70_1),.clk(gclk));
	jdff dff_A_5WA9MwRB4_1(.dout(w_dff_A_rW7uXXy70_1),.din(w_dff_A_5WA9MwRB4_1),.clk(gclk));
	jdff dff_B_244tRTRv6_3(.din(G55gat),.dout(w_dff_B_244tRTRv6_3),.clk(gclk));
	jdff dff_B_lEMQTvZA9_3(.din(w_dff_B_244tRTRv6_3),.dout(w_dff_B_lEMQTvZA9_3),.clk(gclk));
	jdff dff_A_OrDC34Ke6_1(.dout(w_G171gat_0[1]),.din(w_dff_A_OrDC34Ke6_1),.clk(gclk));
	jdff dff_A_sh3SKIBB9_1(.dout(w_dff_A_OrDC34Ke6_1),.din(w_dff_A_sh3SKIBB9_1),.clk(gclk));
	jdff dff_A_K3NLT9Ak4_1(.dout(w_dff_A_sh3SKIBB9_1),.din(w_dff_A_K3NLT9Ak4_1),.clk(gclk));
	jdff dff_A_k3sAJFMy3_1(.dout(w_dff_A_K3NLT9Ak4_1),.din(w_dff_A_k3sAJFMy3_1),.clk(gclk));
	jdff dff_A_V3aHJn8o0_1(.dout(w_dff_A_k3sAJFMy3_1),.din(w_dff_A_V3aHJn8o0_1),.clk(gclk));
	jdff dff_A_2f98JMSZ7_1(.dout(w_dff_A_V3aHJn8o0_1),.din(w_dff_A_2f98JMSZ7_1),.clk(gclk));
	jdff dff_A_foFC6nAh4_1(.dout(w_dff_A_2f98JMSZ7_1),.din(w_dff_A_foFC6nAh4_1),.clk(gclk));
	jdff dff_A_6PmdFaOp5_1(.dout(w_dff_A_foFC6nAh4_1),.din(w_dff_A_6PmdFaOp5_1),.clk(gclk));
	jdff dff_A_aWmdXhqw4_1(.dout(w_dff_A_6PmdFaOp5_1),.din(w_dff_A_aWmdXhqw4_1),.clk(gclk));
	jdff dff_A_vx1IlplW0_2(.dout(w_G171gat_0[2]),.din(w_dff_A_vx1IlplW0_2),.clk(gclk));
	jdff dff_A_UCXNWv1U7_2(.dout(w_dff_A_vx1IlplW0_2),.din(w_dff_A_UCXNWv1U7_2),.clk(gclk));
	jdff dff_A_0qBQ3hYR1_2(.dout(w_dff_A_UCXNWv1U7_2),.din(w_dff_A_0qBQ3hYR1_2),.clk(gclk));
	jdff dff_A_2crjAIGA0_2(.dout(w_dff_A_0qBQ3hYR1_2),.din(w_dff_A_2crjAIGA0_2),.clk(gclk));
	jdff dff_A_IqrXtOF58_2(.dout(w_dff_A_2crjAIGA0_2),.din(w_dff_A_IqrXtOF58_2),.clk(gclk));
	jdff dff_A_IMua5r6F0_2(.dout(w_dff_A_IqrXtOF58_2),.din(w_dff_A_IMua5r6F0_2),.clk(gclk));
	jdff dff_A_M6cJgRvz3_2(.dout(w_dff_A_IMua5r6F0_2),.din(w_dff_A_M6cJgRvz3_2),.clk(gclk));
	jdff dff_A_bnf6zr3H2_2(.dout(w_dff_A_M6cJgRvz3_2),.din(w_dff_A_bnf6zr3H2_2),.clk(gclk));
	jdff dff_A_cyJN6K3q5_2(.dout(w_dff_A_bnf6zr3H2_2),.din(w_dff_A_cyJN6K3q5_2),.clk(gclk));
	jdff dff_A_MchCa0XT1_2(.dout(w_dff_A_cyJN6K3q5_2),.din(w_dff_A_MchCa0XT1_2),.clk(gclk));
	jdff dff_A_YEa8x4XB1_2(.dout(w_dff_A_MchCa0XT1_2),.din(w_dff_A_YEa8x4XB1_2),.clk(gclk));
	jdff dff_A_wF8Cl85X4_2(.dout(w_dff_A_ClLJEkci1_0),.din(w_dff_A_wF8Cl85X4_2),.clk(gclk));
	jdff dff_A_ClLJEkci1_0(.dout(w_dff_A_f6kzESnr4_0),.din(w_dff_A_ClLJEkci1_0),.clk(gclk));
	jdff dff_A_f6kzESnr4_0(.dout(w_dff_A_tKHLe5Cw2_0),.din(w_dff_A_f6kzESnr4_0),.clk(gclk));
	jdff dff_A_tKHLe5Cw2_0(.dout(w_dff_A_JWwv185I6_0),.din(w_dff_A_tKHLe5Cw2_0),.clk(gclk));
	jdff dff_A_JWwv185I6_0(.dout(w_dff_A_FC34CPBS3_0),.din(w_dff_A_JWwv185I6_0),.clk(gclk));
	jdff dff_A_FC34CPBS3_0(.dout(w_dff_A_QqRuJ6Mz7_0),.din(w_dff_A_FC34CPBS3_0),.clk(gclk));
	jdff dff_A_QqRuJ6Mz7_0(.dout(w_dff_A_hPp50bWJ9_0),.din(w_dff_A_QqRuJ6Mz7_0),.clk(gclk));
	jdff dff_A_hPp50bWJ9_0(.dout(w_dff_A_ClnPAPNM7_0),.din(w_dff_A_hPp50bWJ9_0),.clk(gclk));
	jdff dff_A_ClnPAPNM7_0(.dout(w_dff_A_mFisWiIl3_0),.din(w_dff_A_ClnPAPNM7_0),.clk(gclk));
	jdff dff_A_mFisWiIl3_0(.dout(w_dff_A_LQZ9fwxO8_0),.din(w_dff_A_mFisWiIl3_0),.clk(gclk));
	jdff dff_A_LQZ9fwxO8_0(.dout(w_dff_A_sZJoyY4C3_0),.din(w_dff_A_LQZ9fwxO8_0),.clk(gclk));
	jdff dff_A_sZJoyY4C3_0(.dout(w_dff_A_IK1gHZ8x6_0),.din(w_dff_A_sZJoyY4C3_0),.clk(gclk));
	jdff dff_A_IK1gHZ8x6_0(.dout(w_dff_A_joFkzNBo9_0),.din(w_dff_A_IK1gHZ8x6_0),.clk(gclk));
	jdff dff_A_joFkzNBo9_0(.dout(w_dff_A_EME01GPk3_0),.din(w_dff_A_joFkzNBo9_0),.clk(gclk));
	jdff dff_A_EME01GPk3_0(.dout(w_dff_A_2KG3pNHw2_0),.din(w_dff_A_EME01GPk3_0),.clk(gclk));
	jdff dff_A_2KG3pNHw2_0(.dout(w_dff_A_evZ0erhW1_0),.din(w_dff_A_2KG3pNHw2_0),.clk(gclk));
	jdff dff_A_evZ0erhW1_0(.dout(w_dff_A_6lm5GJZU3_0),.din(w_dff_A_evZ0erhW1_0),.clk(gclk));
	jdff dff_A_6lm5GJZU3_0(.dout(w_dff_A_4RpFJ8NO5_0),.din(w_dff_A_6lm5GJZU3_0),.clk(gclk));
	jdff dff_A_4RpFJ8NO5_0(.dout(w_dff_A_Db8WX77x7_0),.din(w_dff_A_4RpFJ8NO5_0),.clk(gclk));
	jdff dff_A_Db8WX77x7_0(.dout(w_dff_A_oUv0FQ8Q0_0),.din(w_dff_A_Db8WX77x7_0),.clk(gclk));
	jdff dff_A_oUv0FQ8Q0_0(.dout(w_dff_A_1vk4U44o1_0),.din(w_dff_A_oUv0FQ8Q0_0),.clk(gclk));
	jdff dff_A_1vk4U44o1_0(.dout(w_dff_A_TlymtKvy7_0),.din(w_dff_A_1vk4U44o1_0),.clk(gclk));
	jdff dff_A_TlymtKvy7_0(.dout(w_dff_A_bZ5MyR6O9_0),.din(w_dff_A_TlymtKvy7_0),.clk(gclk));
	jdff dff_A_bZ5MyR6O9_0(.dout(w_dff_A_6rixA4pP6_0),.din(w_dff_A_bZ5MyR6O9_0),.clk(gclk));
	jdff dff_A_6rixA4pP6_0(.dout(w_dff_A_HsDIHK2K7_0),.din(w_dff_A_6rixA4pP6_0),.clk(gclk));
	jdff dff_A_HsDIHK2K7_0(.dout(G388gat),.din(w_dff_A_HsDIHK2K7_0),.clk(gclk));
	jdff dff_A_URn4EI0h7_2(.dout(w_dff_A_XU4X6X4G4_0),.din(w_dff_A_URn4EI0h7_2),.clk(gclk));
	jdff dff_A_XU4X6X4G4_0(.dout(w_dff_A_eN3cOpU68_0),.din(w_dff_A_XU4X6X4G4_0),.clk(gclk));
	jdff dff_A_eN3cOpU68_0(.dout(w_dff_A_Phqa3cVI6_0),.din(w_dff_A_eN3cOpU68_0),.clk(gclk));
	jdff dff_A_Phqa3cVI6_0(.dout(w_dff_A_WMxX7sO32_0),.din(w_dff_A_Phqa3cVI6_0),.clk(gclk));
	jdff dff_A_WMxX7sO32_0(.dout(w_dff_A_VsfHtiiX0_0),.din(w_dff_A_WMxX7sO32_0),.clk(gclk));
	jdff dff_A_VsfHtiiX0_0(.dout(w_dff_A_YygaCAQN5_0),.din(w_dff_A_VsfHtiiX0_0),.clk(gclk));
	jdff dff_A_YygaCAQN5_0(.dout(w_dff_A_6gY5i48W2_0),.din(w_dff_A_YygaCAQN5_0),.clk(gclk));
	jdff dff_A_6gY5i48W2_0(.dout(w_dff_A_Gfwt14mj8_0),.din(w_dff_A_6gY5i48W2_0),.clk(gclk));
	jdff dff_A_Gfwt14mj8_0(.dout(w_dff_A_k34j0FCu9_0),.din(w_dff_A_Gfwt14mj8_0),.clk(gclk));
	jdff dff_A_k34j0FCu9_0(.dout(w_dff_A_v20MPbiG9_0),.din(w_dff_A_k34j0FCu9_0),.clk(gclk));
	jdff dff_A_v20MPbiG9_0(.dout(w_dff_A_gjGv3n1a4_0),.din(w_dff_A_v20MPbiG9_0),.clk(gclk));
	jdff dff_A_gjGv3n1a4_0(.dout(w_dff_A_g5vGD8Aq1_0),.din(w_dff_A_gjGv3n1a4_0),.clk(gclk));
	jdff dff_A_g5vGD8Aq1_0(.dout(w_dff_A_4ZouqCnj2_0),.din(w_dff_A_g5vGD8Aq1_0),.clk(gclk));
	jdff dff_A_4ZouqCnj2_0(.dout(w_dff_A_1DA1D5Mc6_0),.din(w_dff_A_4ZouqCnj2_0),.clk(gclk));
	jdff dff_A_1DA1D5Mc6_0(.dout(w_dff_A_drPR7nGB2_0),.din(w_dff_A_1DA1D5Mc6_0),.clk(gclk));
	jdff dff_A_drPR7nGB2_0(.dout(w_dff_A_UKTifiP88_0),.din(w_dff_A_drPR7nGB2_0),.clk(gclk));
	jdff dff_A_UKTifiP88_0(.dout(w_dff_A_gycEUIEt7_0),.din(w_dff_A_UKTifiP88_0),.clk(gclk));
	jdff dff_A_gycEUIEt7_0(.dout(w_dff_A_qbSLaw9U7_0),.din(w_dff_A_gycEUIEt7_0),.clk(gclk));
	jdff dff_A_qbSLaw9U7_0(.dout(w_dff_A_sRsqK2Np6_0),.din(w_dff_A_qbSLaw9U7_0),.clk(gclk));
	jdff dff_A_sRsqK2Np6_0(.dout(w_dff_A_2h9Grpbb5_0),.din(w_dff_A_sRsqK2Np6_0),.clk(gclk));
	jdff dff_A_2h9Grpbb5_0(.dout(w_dff_A_kjPyLyTg1_0),.din(w_dff_A_2h9Grpbb5_0),.clk(gclk));
	jdff dff_A_kjPyLyTg1_0(.dout(w_dff_A_hqqkMEyB7_0),.din(w_dff_A_kjPyLyTg1_0),.clk(gclk));
	jdff dff_A_hqqkMEyB7_0(.dout(w_dff_A_j95b8i4I1_0),.din(w_dff_A_hqqkMEyB7_0),.clk(gclk));
	jdff dff_A_j95b8i4I1_0(.dout(w_dff_A_MpPJ47RF0_0),.din(w_dff_A_j95b8i4I1_0),.clk(gclk));
	jdff dff_A_MpPJ47RF0_0(.dout(w_dff_A_CkOdEVXw9_0),.din(w_dff_A_MpPJ47RF0_0),.clk(gclk));
	jdff dff_A_CkOdEVXw9_0(.dout(G389gat),.din(w_dff_A_CkOdEVXw9_0),.clk(gclk));
	jdff dff_A_DCUnLUjN5_2(.dout(w_dff_A_LK3B1J3Q0_0),.din(w_dff_A_DCUnLUjN5_2),.clk(gclk));
	jdff dff_A_LK3B1J3Q0_0(.dout(w_dff_A_4UCHGtCy9_0),.din(w_dff_A_LK3B1J3Q0_0),.clk(gclk));
	jdff dff_A_4UCHGtCy9_0(.dout(w_dff_A_L5lWpIQT0_0),.din(w_dff_A_4UCHGtCy9_0),.clk(gclk));
	jdff dff_A_L5lWpIQT0_0(.dout(w_dff_A_YpNPzlTs9_0),.din(w_dff_A_L5lWpIQT0_0),.clk(gclk));
	jdff dff_A_YpNPzlTs9_0(.dout(w_dff_A_vvj60zCk8_0),.din(w_dff_A_YpNPzlTs9_0),.clk(gclk));
	jdff dff_A_vvj60zCk8_0(.dout(w_dff_A_J9zBqNvc1_0),.din(w_dff_A_vvj60zCk8_0),.clk(gclk));
	jdff dff_A_J9zBqNvc1_0(.dout(w_dff_A_VuZSqEM76_0),.din(w_dff_A_J9zBqNvc1_0),.clk(gclk));
	jdff dff_A_VuZSqEM76_0(.dout(w_dff_A_ySaquppi4_0),.din(w_dff_A_VuZSqEM76_0),.clk(gclk));
	jdff dff_A_ySaquppi4_0(.dout(w_dff_A_QOoTBZhk3_0),.din(w_dff_A_ySaquppi4_0),.clk(gclk));
	jdff dff_A_QOoTBZhk3_0(.dout(w_dff_A_4pUseqsY3_0),.din(w_dff_A_QOoTBZhk3_0),.clk(gclk));
	jdff dff_A_4pUseqsY3_0(.dout(w_dff_A_vuKy39YH7_0),.din(w_dff_A_4pUseqsY3_0),.clk(gclk));
	jdff dff_A_vuKy39YH7_0(.dout(w_dff_A_O6bLVEVt0_0),.din(w_dff_A_vuKy39YH7_0),.clk(gclk));
	jdff dff_A_O6bLVEVt0_0(.dout(w_dff_A_ORTJY1pH6_0),.din(w_dff_A_O6bLVEVt0_0),.clk(gclk));
	jdff dff_A_ORTJY1pH6_0(.dout(w_dff_A_lQDhlEbv0_0),.din(w_dff_A_ORTJY1pH6_0),.clk(gclk));
	jdff dff_A_lQDhlEbv0_0(.dout(w_dff_A_Pyv83LjJ3_0),.din(w_dff_A_lQDhlEbv0_0),.clk(gclk));
	jdff dff_A_Pyv83LjJ3_0(.dout(w_dff_A_sQ48iNgC9_0),.din(w_dff_A_Pyv83LjJ3_0),.clk(gclk));
	jdff dff_A_sQ48iNgC9_0(.dout(w_dff_A_6XZ86Acu6_0),.din(w_dff_A_sQ48iNgC9_0),.clk(gclk));
	jdff dff_A_6XZ86Acu6_0(.dout(w_dff_A_35EwFhGE1_0),.din(w_dff_A_6XZ86Acu6_0),.clk(gclk));
	jdff dff_A_35EwFhGE1_0(.dout(w_dff_A_6Yz27eOL3_0),.din(w_dff_A_35EwFhGE1_0),.clk(gclk));
	jdff dff_A_6Yz27eOL3_0(.dout(w_dff_A_T5XnaazA0_0),.din(w_dff_A_6Yz27eOL3_0),.clk(gclk));
	jdff dff_A_T5XnaazA0_0(.dout(w_dff_A_EPCzY0nk0_0),.din(w_dff_A_T5XnaazA0_0),.clk(gclk));
	jdff dff_A_EPCzY0nk0_0(.dout(w_dff_A_ySH44Wtm2_0),.din(w_dff_A_EPCzY0nk0_0),.clk(gclk));
	jdff dff_A_ySH44Wtm2_0(.dout(w_dff_A_HVtHdww27_0),.din(w_dff_A_ySH44Wtm2_0),.clk(gclk));
	jdff dff_A_HVtHdww27_0(.dout(w_dff_A_XoQZlwbF4_0),.din(w_dff_A_HVtHdww27_0),.clk(gclk));
	jdff dff_A_XoQZlwbF4_0(.dout(w_dff_A_f97qhAPz3_0),.din(w_dff_A_XoQZlwbF4_0),.clk(gclk));
	jdff dff_A_f97qhAPz3_0(.dout(G390gat),.din(w_dff_A_f97qhAPz3_0),.clk(gclk));
	jdff dff_A_8pBCiBMs8_2(.dout(w_dff_A_clRKRtNn5_0),.din(w_dff_A_8pBCiBMs8_2),.clk(gclk));
	jdff dff_A_clRKRtNn5_0(.dout(w_dff_A_F1xYbvEk6_0),.din(w_dff_A_clRKRtNn5_0),.clk(gclk));
	jdff dff_A_F1xYbvEk6_0(.dout(w_dff_A_mwbhn23q5_0),.din(w_dff_A_F1xYbvEk6_0),.clk(gclk));
	jdff dff_A_mwbhn23q5_0(.dout(w_dff_A_F4CG209h0_0),.din(w_dff_A_mwbhn23q5_0),.clk(gclk));
	jdff dff_A_F4CG209h0_0(.dout(w_dff_A_6SrCwavk3_0),.din(w_dff_A_F4CG209h0_0),.clk(gclk));
	jdff dff_A_6SrCwavk3_0(.dout(w_dff_A_erjEthf31_0),.din(w_dff_A_6SrCwavk3_0),.clk(gclk));
	jdff dff_A_erjEthf31_0(.dout(w_dff_A_a68gOB9j7_0),.din(w_dff_A_erjEthf31_0),.clk(gclk));
	jdff dff_A_a68gOB9j7_0(.dout(w_dff_A_WB4HwnZq6_0),.din(w_dff_A_a68gOB9j7_0),.clk(gclk));
	jdff dff_A_WB4HwnZq6_0(.dout(w_dff_A_Zxswmoi59_0),.din(w_dff_A_WB4HwnZq6_0),.clk(gclk));
	jdff dff_A_Zxswmoi59_0(.dout(w_dff_A_rHv7T4Nd0_0),.din(w_dff_A_Zxswmoi59_0),.clk(gclk));
	jdff dff_A_rHv7T4Nd0_0(.dout(w_dff_A_2ZAVattz3_0),.din(w_dff_A_rHv7T4Nd0_0),.clk(gclk));
	jdff dff_A_2ZAVattz3_0(.dout(w_dff_A_p3eZOdir1_0),.din(w_dff_A_2ZAVattz3_0),.clk(gclk));
	jdff dff_A_p3eZOdir1_0(.dout(w_dff_A_o6NAy5RB9_0),.din(w_dff_A_p3eZOdir1_0),.clk(gclk));
	jdff dff_A_o6NAy5RB9_0(.dout(w_dff_A_hBWVZAPV9_0),.din(w_dff_A_o6NAy5RB9_0),.clk(gclk));
	jdff dff_A_hBWVZAPV9_0(.dout(w_dff_A_K71kYyS69_0),.din(w_dff_A_hBWVZAPV9_0),.clk(gclk));
	jdff dff_A_K71kYyS69_0(.dout(w_dff_A_ssp9WvJv0_0),.din(w_dff_A_K71kYyS69_0),.clk(gclk));
	jdff dff_A_ssp9WvJv0_0(.dout(w_dff_A_ZwAROs2J7_0),.din(w_dff_A_ssp9WvJv0_0),.clk(gclk));
	jdff dff_A_ZwAROs2J7_0(.dout(w_dff_A_Ebv1GTbQ8_0),.din(w_dff_A_ZwAROs2J7_0),.clk(gclk));
	jdff dff_A_Ebv1GTbQ8_0(.dout(w_dff_A_S0BYbNXc0_0),.din(w_dff_A_Ebv1GTbQ8_0),.clk(gclk));
	jdff dff_A_S0BYbNXc0_0(.dout(w_dff_A_tgchaNDi7_0),.din(w_dff_A_S0BYbNXc0_0),.clk(gclk));
	jdff dff_A_tgchaNDi7_0(.dout(w_dff_A_1V4BEQ3z7_0),.din(w_dff_A_tgchaNDi7_0),.clk(gclk));
	jdff dff_A_1V4BEQ3z7_0(.dout(w_dff_A_8u12CGUO6_0),.din(w_dff_A_1V4BEQ3z7_0),.clk(gclk));
	jdff dff_A_8u12CGUO6_0(.dout(w_dff_A_KD0GetWJ0_0),.din(w_dff_A_8u12CGUO6_0),.clk(gclk));
	jdff dff_A_KD0GetWJ0_0(.dout(w_dff_A_LhUQn7548_0),.din(w_dff_A_KD0GetWJ0_0),.clk(gclk));
	jdff dff_A_LhUQn7548_0(.dout(w_dff_A_04EcVYd20_0),.din(w_dff_A_LhUQn7548_0),.clk(gclk));
	jdff dff_A_04EcVYd20_0(.dout(w_dff_A_te6HLR6I3_0),.din(w_dff_A_04EcVYd20_0),.clk(gclk));
	jdff dff_A_te6HLR6I3_0(.dout(G391gat),.din(w_dff_A_te6HLR6I3_0),.clk(gclk));
	jdff dff_A_h8jo52As9_2(.dout(w_dff_A_R75aPu7G3_0),.din(w_dff_A_h8jo52As9_2),.clk(gclk));
	jdff dff_A_R75aPu7G3_0(.dout(w_dff_A_EwHYCa2j3_0),.din(w_dff_A_R75aPu7G3_0),.clk(gclk));
	jdff dff_A_EwHYCa2j3_0(.dout(w_dff_A_3hOOZs231_0),.din(w_dff_A_EwHYCa2j3_0),.clk(gclk));
	jdff dff_A_3hOOZs231_0(.dout(w_dff_A_UNaLyMaH6_0),.din(w_dff_A_3hOOZs231_0),.clk(gclk));
	jdff dff_A_UNaLyMaH6_0(.dout(w_dff_A_tNThjERl2_0),.din(w_dff_A_UNaLyMaH6_0),.clk(gclk));
	jdff dff_A_tNThjERl2_0(.dout(w_dff_A_uHLHGbMT5_0),.din(w_dff_A_tNThjERl2_0),.clk(gclk));
	jdff dff_A_uHLHGbMT5_0(.dout(w_dff_A_HTYfIR785_0),.din(w_dff_A_uHLHGbMT5_0),.clk(gclk));
	jdff dff_A_HTYfIR785_0(.dout(w_dff_A_M9YJ3cWh0_0),.din(w_dff_A_HTYfIR785_0),.clk(gclk));
	jdff dff_A_M9YJ3cWh0_0(.dout(w_dff_A_8SPFwIRK5_0),.din(w_dff_A_M9YJ3cWh0_0),.clk(gclk));
	jdff dff_A_8SPFwIRK5_0(.dout(w_dff_A_XoWZiUEt3_0),.din(w_dff_A_8SPFwIRK5_0),.clk(gclk));
	jdff dff_A_XoWZiUEt3_0(.dout(w_dff_A_2uGbiMSz7_0),.din(w_dff_A_XoWZiUEt3_0),.clk(gclk));
	jdff dff_A_2uGbiMSz7_0(.dout(w_dff_A_XJMQcD9b0_0),.din(w_dff_A_2uGbiMSz7_0),.clk(gclk));
	jdff dff_A_XJMQcD9b0_0(.dout(w_dff_A_tCtRc8VJ8_0),.din(w_dff_A_XJMQcD9b0_0),.clk(gclk));
	jdff dff_A_tCtRc8VJ8_0(.dout(w_dff_A_UNHayenH9_0),.din(w_dff_A_tCtRc8VJ8_0),.clk(gclk));
	jdff dff_A_UNHayenH9_0(.dout(w_dff_A_YRDJ7zfO1_0),.din(w_dff_A_UNHayenH9_0),.clk(gclk));
	jdff dff_A_YRDJ7zfO1_0(.dout(w_dff_A_RE4s87sI8_0),.din(w_dff_A_YRDJ7zfO1_0),.clk(gclk));
	jdff dff_A_RE4s87sI8_0(.dout(w_dff_A_H1e0lKX53_0),.din(w_dff_A_RE4s87sI8_0),.clk(gclk));
	jdff dff_A_H1e0lKX53_0(.dout(w_dff_A_9sVH2EWT8_0),.din(w_dff_A_H1e0lKX53_0),.clk(gclk));
	jdff dff_A_9sVH2EWT8_0(.dout(w_dff_A_UJ29qjt87_0),.din(w_dff_A_9sVH2EWT8_0),.clk(gclk));
	jdff dff_A_UJ29qjt87_0(.dout(w_dff_A_j6E1AQjs1_0),.din(w_dff_A_UJ29qjt87_0),.clk(gclk));
	jdff dff_A_j6E1AQjs1_0(.dout(w_dff_A_ywOoEXd11_0),.din(w_dff_A_j6E1AQjs1_0),.clk(gclk));
	jdff dff_A_ywOoEXd11_0(.dout(w_dff_A_rEkvsX6m7_0),.din(w_dff_A_ywOoEXd11_0),.clk(gclk));
	jdff dff_A_rEkvsX6m7_0(.dout(w_dff_A_xTDZk3NR1_0),.din(w_dff_A_rEkvsX6m7_0),.clk(gclk));
	jdff dff_A_xTDZk3NR1_0(.dout(w_dff_A_gyR8xsKb6_0),.din(w_dff_A_xTDZk3NR1_0),.clk(gclk));
	jdff dff_A_gyR8xsKb6_0(.dout(G418gat),.din(w_dff_A_gyR8xsKb6_0),.clk(gclk));
	jdff dff_A_laVyLnLT1_2(.dout(w_dff_A_DIISTH446_0),.din(w_dff_A_laVyLnLT1_2),.clk(gclk));
	jdff dff_A_DIISTH446_0(.dout(w_dff_A_z5pexYFN7_0),.din(w_dff_A_DIISTH446_0),.clk(gclk));
	jdff dff_A_z5pexYFN7_0(.dout(w_dff_A_C7NokHXA2_0),.din(w_dff_A_z5pexYFN7_0),.clk(gclk));
	jdff dff_A_C7NokHXA2_0(.dout(w_dff_A_cDGkuiuT6_0),.din(w_dff_A_C7NokHXA2_0),.clk(gclk));
	jdff dff_A_cDGkuiuT6_0(.dout(w_dff_A_lopyjr0n8_0),.din(w_dff_A_cDGkuiuT6_0),.clk(gclk));
	jdff dff_A_lopyjr0n8_0(.dout(w_dff_A_dHbgcKoN5_0),.din(w_dff_A_lopyjr0n8_0),.clk(gclk));
	jdff dff_A_dHbgcKoN5_0(.dout(w_dff_A_YrhhiGQw7_0),.din(w_dff_A_dHbgcKoN5_0),.clk(gclk));
	jdff dff_A_YrhhiGQw7_0(.dout(w_dff_A_RtdbOFHE2_0),.din(w_dff_A_YrhhiGQw7_0),.clk(gclk));
	jdff dff_A_RtdbOFHE2_0(.dout(w_dff_A_C6d8BV7I8_0),.din(w_dff_A_RtdbOFHE2_0),.clk(gclk));
	jdff dff_A_C6d8BV7I8_0(.dout(w_dff_A_qopnCWSg8_0),.din(w_dff_A_C6d8BV7I8_0),.clk(gclk));
	jdff dff_A_qopnCWSg8_0(.dout(w_dff_A_C3l1wK7Q2_0),.din(w_dff_A_qopnCWSg8_0),.clk(gclk));
	jdff dff_A_C3l1wK7Q2_0(.dout(w_dff_A_NPaJ6teP8_0),.din(w_dff_A_C3l1wK7Q2_0),.clk(gclk));
	jdff dff_A_NPaJ6teP8_0(.dout(w_dff_A_lMVnUSQa9_0),.din(w_dff_A_NPaJ6teP8_0),.clk(gclk));
	jdff dff_A_lMVnUSQa9_0(.dout(w_dff_A_VwATLboz1_0),.din(w_dff_A_lMVnUSQa9_0),.clk(gclk));
	jdff dff_A_VwATLboz1_0(.dout(w_dff_A_Ov7GXoYI1_0),.din(w_dff_A_VwATLboz1_0),.clk(gclk));
	jdff dff_A_Ov7GXoYI1_0(.dout(w_dff_A_w1fPEtm99_0),.din(w_dff_A_Ov7GXoYI1_0),.clk(gclk));
	jdff dff_A_w1fPEtm99_0(.dout(w_dff_A_mMXNLHmQ0_0),.din(w_dff_A_w1fPEtm99_0),.clk(gclk));
	jdff dff_A_mMXNLHmQ0_0(.dout(w_dff_A_WHGfAUfB5_0),.din(w_dff_A_mMXNLHmQ0_0),.clk(gclk));
	jdff dff_A_WHGfAUfB5_0(.dout(w_dff_A_bePrq1Ae9_0),.din(w_dff_A_WHGfAUfB5_0),.clk(gclk));
	jdff dff_A_bePrq1Ae9_0(.dout(w_dff_A_gJZmO8AF9_0),.din(w_dff_A_bePrq1Ae9_0),.clk(gclk));
	jdff dff_A_gJZmO8AF9_0(.dout(w_dff_A_fFKp0A8X8_0),.din(w_dff_A_gJZmO8AF9_0),.clk(gclk));
	jdff dff_A_fFKp0A8X8_0(.dout(w_dff_A_nBLlvPvN3_0),.din(w_dff_A_fFKp0A8X8_0),.clk(gclk));
	jdff dff_A_nBLlvPvN3_0(.dout(G419gat),.din(w_dff_A_nBLlvPvN3_0),.clk(gclk));
	jdff dff_A_deOSyrnr7_2(.dout(w_dff_A_a4fwSDdu0_0),.din(w_dff_A_deOSyrnr7_2),.clk(gclk));
	jdff dff_A_a4fwSDdu0_0(.dout(w_dff_A_Bjl15bpH7_0),.din(w_dff_A_a4fwSDdu0_0),.clk(gclk));
	jdff dff_A_Bjl15bpH7_0(.dout(w_dff_A_b8SdHcNp8_0),.din(w_dff_A_Bjl15bpH7_0),.clk(gclk));
	jdff dff_A_b8SdHcNp8_0(.dout(w_dff_A_Ovob1aRK7_0),.din(w_dff_A_b8SdHcNp8_0),.clk(gclk));
	jdff dff_A_Ovob1aRK7_0(.dout(w_dff_A_SQXgrj802_0),.din(w_dff_A_Ovob1aRK7_0),.clk(gclk));
	jdff dff_A_SQXgrj802_0(.dout(w_dff_A_gfpiyVsr9_0),.din(w_dff_A_SQXgrj802_0),.clk(gclk));
	jdff dff_A_gfpiyVsr9_0(.dout(w_dff_A_q9RiCr198_0),.din(w_dff_A_gfpiyVsr9_0),.clk(gclk));
	jdff dff_A_q9RiCr198_0(.dout(w_dff_A_6cGXUVLp6_0),.din(w_dff_A_q9RiCr198_0),.clk(gclk));
	jdff dff_A_6cGXUVLp6_0(.dout(w_dff_A_NBR5S5FV9_0),.din(w_dff_A_6cGXUVLp6_0),.clk(gclk));
	jdff dff_A_NBR5S5FV9_0(.dout(w_dff_A_tgussN988_0),.din(w_dff_A_NBR5S5FV9_0),.clk(gclk));
	jdff dff_A_tgussN988_0(.dout(w_dff_A_kLK4FU254_0),.din(w_dff_A_tgussN988_0),.clk(gclk));
	jdff dff_A_kLK4FU254_0(.dout(w_dff_A_S0tChvUW8_0),.din(w_dff_A_kLK4FU254_0),.clk(gclk));
	jdff dff_A_S0tChvUW8_0(.dout(w_dff_A_vNXHHIjf9_0),.din(w_dff_A_S0tChvUW8_0),.clk(gclk));
	jdff dff_A_vNXHHIjf9_0(.dout(w_dff_A_H937d63b3_0),.din(w_dff_A_vNXHHIjf9_0),.clk(gclk));
	jdff dff_A_H937d63b3_0(.dout(w_dff_A_EUn111oZ0_0),.din(w_dff_A_H937d63b3_0),.clk(gclk));
	jdff dff_A_EUn111oZ0_0(.dout(w_dff_A_ioefZaX57_0),.din(w_dff_A_EUn111oZ0_0),.clk(gclk));
	jdff dff_A_ioefZaX57_0(.dout(w_dff_A_9H0l3MS87_0),.din(w_dff_A_ioefZaX57_0),.clk(gclk));
	jdff dff_A_9H0l3MS87_0(.dout(w_dff_A_xBDueBwD2_0),.din(w_dff_A_9H0l3MS87_0),.clk(gclk));
	jdff dff_A_xBDueBwD2_0(.dout(w_dff_A_CuuDcqMy7_0),.din(w_dff_A_xBDueBwD2_0),.clk(gclk));
	jdff dff_A_CuuDcqMy7_0(.dout(w_dff_A_b0mAXX6M5_0),.din(w_dff_A_CuuDcqMy7_0),.clk(gclk));
	jdff dff_A_b0mAXX6M5_0(.dout(w_dff_A_akTJ28XZ2_0),.din(w_dff_A_b0mAXX6M5_0),.clk(gclk));
	jdff dff_A_akTJ28XZ2_0(.dout(w_dff_A_fVpoRMzG0_0),.din(w_dff_A_akTJ28XZ2_0),.clk(gclk));
	jdff dff_A_fVpoRMzG0_0(.dout(w_dff_A_QEwcGjuL7_0),.din(w_dff_A_fVpoRMzG0_0),.clk(gclk));
	jdff dff_A_QEwcGjuL7_0(.dout(w_dff_A_K9G3agmX4_0),.din(w_dff_A_QEwcGjuL7_0),.clk(gclk));
	jdff dff_A_K9G3agmX4_0(.dout(G420gat),.din(w_dff_A_K9G3agmX4_0),.clk(gclk));
	jdff dff_A_lrqAObpH1_2(.dout(w_dff_A_GcKxzyGJ6_0),.din(w_dff_A_lrqAObpH1_2),.clk(gclk));
	jdff dff_A_GcKxzyGJ6_0(.dout(w_dff_A_GmhPtNCE3_0),.din(w_dff_A_GcKxzyGJ6_0),.clk(gclk));
	jdff dff_A_GmhPtNCE3_0(.dout(w_dff_A_nwps0OYt5_0),.din(w_dff_A_GmhPtNCE3_0),.clk(gclk));
	jdff dff_A_nwps0OYt5_0(.dout(w_dff_A_PiJuzgoU7_0),.din(w_dff_A_nwps0OYt5_0),.clk(gclk));
	jdff dff_A_PiJuzgoU7_0(.dout(w_dff_A_nLm44Rnf1_0),.din(w_dff_A_PiJuzgoU7_0),.clk(gclk));
	jdff dff_A_nLm44Rnf1_0(.dout(w_dff_A_IZBxedDW6_0),.din(w_dff_A_nLm44Rnf1_0),.clk(gclk));
	jdff dff_A_IZBxedDW6_0(.dout(w_dff_A_yXKPRIBm4_0),.din(w_dff_A_IZBxedDW6_0),.clk(gclk));
	jdff dff_A_yXKPRIBm4_0(.dout(w_dff_A_UanwxyNM5_0),.din(w_dff_A_yXKPRIBm4_0),.clk(gclk));
	jdff dff_A_UanwxyNM5_0(.dout(w_dff_A_hnWstzmq3_0),.din(w_dff_A_UanwxyNM5_0),.clk(gclk));
	jdff dff_A_hnWstzmq3_0(.dout(w_dff_A_rEqdIL1A6_0),.din(w_dff_A_hnWstzmq3_0),.clk(gclk));
	jdff dff_A_rEqdIL1A6_0(.dout(w_dff_A_aDdIWWAw5_0),.din(w_dff_A_rEqdIL1A6_0),.clk(gclk));
	jdff dff_A_aDdIWWAw5_0(.dout(w_dff_A_nC26oicF6_0),.din(w_dff_A_aDdIWWAw5_0),.clk(gclk));
	jdff dff_A_nC26oicF6_0(.dout(w_dff_A_6uET4wis0_0),.din(w_dff_A_nC26oicF6_0),.clk(gclk));
	jdff dff_A_6uET4wis0_0(.dout(w_dff_A_AEDBBR8K6_0),.din(w_dff_A_6uET4wis0_0),.clk(gclk));
	jdff dff_A_AEDBBR8K6_0(.dout(w_dff_A_5eQrw2qB3_0),.din(w_dff_A_AEDBBR8K6_0),.clk(gclk));
	jdff dff_A_5eQrw2qB3_0(.dout(w_dff_A_i8KaPZQ84_0),.din(w_dff_A_5eQrw2qB3_0),.clk(gclk));
	jdff dff_A_i8KaPZQ84_0(.dout(w_dff_A_9BbMzB5n3_0),.din(w_dff_A_i8KaPZQ84_0),.clk(gclk));
	jdff dff_A_9BbMzB5n3_0(.dout(w_dff_A_nTfYHYpn1_0),.din(w_dff_A_9BbMzB5n3_0),.clk(gclk));
	jdff dff_A_nTfYHYpn1_0(.dout(w_dff_A_glGd2eIY0_0),.din(w_dff_A_nTfYHYpn1_0),.clk(gclk));
	jdff dff_A_glGd2eIY0_0(.dout(w_dff_A_kFXj5wby9_0),.din(w_dff_A_glGd2eIY0_0),.clk(gclk));
	jdff dff_A_kFXj5wby9_0(.dout(w_dff_A_FR4YFsJa2_0),.din(w_dff_A_kFXj5wby9_0),.clk(gclk));
	jdff dff_A_FR4YFsJa2_0(.dout(w_dff_A_bZpnLv9f9_0),.din(w_dff_A_FR4YFsJa2_0),.clk(gclk));
	jdff dff_A_bZpnLv9f9_0(.dout(w_dff_A_o90m62D30_0),.din(w_dff_A_bZpnLv9f9_0),.clk(gclk));
	jdff dff_A_o90m62D30_0(.dout(w_dff_A_vUia2Ft49_0),.din(w_dff_A_o90m62D30_0),.clk(gclk));
	jdff dff_A_vUia2Ft49_0(.dout(G421gat),.din(w_dff_A_vUia2Ft49_0),.clk(gclk));
	jdff dff_A_wFW2ch691_2(.dout(w_dff_A_nUq230zl4_0),.din(w_dff_A_wFW2ch691_2),.clk(gclk));
	jdff dff_A_nUq230zl4_0(.dout(w_dff_A_qSwWXXuX5_0),.din(w_dff_A_nUq230zl4_0),.clk(gclk));
	jdff dff_A_qSwWXXuX5_0(.dout(w_dff_A_JYnFWZ4p0_0),.din(w_dff_A_qSwWXXuX5_0),.clk(gclk));
	jdff dff_A_JYnFWZ4p0_0(.dout(w_dff_A_6Tbd5IY18_0),.din(w_dff_A_JYnFWZ4p0_0),.clk(gclk));
	jdff dff_A_6Tbd5IY18_0(.dout(w_dff_A_dFpr3Elq1_0),.din(w_dff_A_6Tbd5IY18_0),.clk(gclk));
	jdff dff_A_dFpr3Elq1_0(.dout(w_dff_A_RyCOhIiE7_0),.din(w_dff_A_dFpr3Elq1_0),.clk(gclk));
	jdff dff_A_RyCOhIiE7_0(.dout(w_dff_A_oimxdRd20_0),.din(w_dff_A_RyCOhIiE7_0),.clk(gclk));
	jdff dff_A_oimxdRd20_0(.dout(w_dff_A_eBcUOe005_0),.din(w_dff_A_oimxdRd20_0),.clk(gclk));
	jdff dff_A_eBcUOe005_0(.dout(w_dff_A_x3WlSW253_0),.din(w_dff_A_eBcUOe005_0),.clk(gclk));
	jdff dff_A_x3WlSW253_0(.dout(w_dff_A_heONL2uT7_0),.din(w_dff_A_x3WlSW253_0),.clk(gclk));
	jdff dff_A_heONL2uT7_0(.dout(w_dff_A_EV4S88b56_0),.din(w_dff_A_heONL2uT7_0),.clk(gclk));
	jdff dff_A_EV4S88b56_0(.dout(w_dff_A_rgZALcik5_0),.din(w_dff_A_EV4S88b56_0),.clk(gclk));
	jdff dff_A_rgZALcik5_0(.dout(w_dff_A_4eWjyWWv5_0),.din(w_dff_A_rgZALcik5_0),.clk(gclk));
	jdff dff_A_4eWjyWWv5_0(.dout(w_dff_A_VNptx7qK4_0),.din(w_dff_A_4eWjyWWv5_0),.clk(gclk));
	jdff dff_A_VNptx7qK4_0(.dout(w_dff_A_iUn7dDuR6_0),.din(w_dff_A_VNptx7qK4_0),.clk(gclk));
	jdff dff_A_iUn7dDuR6_0(.dout(w_dff_A_Ut4nLxxv1_0),.din(w_dff_A_iUn7dDuR6_0),.clk(gclk));
	jdff dff_A_Ut4nLxxv1_0(.dout(w_dff_A_BJQ5DKvF3_0),.din(w_dff_A_Ut4nLxxv1_0),.clk(gclk));
	jdff dff_A_BJQ5DKvF3_0(.dout(w_dff_A_lTPtvgTj5_0),.din(w_dff_A_BJQ5DKvF3_0),.clk(gclk));
	jdff dff_A_lTPtvgTj5_0(.dout(w_dff_A_l0yD8ZRM2_0),.din(w_dff_A_lTPtvgTj5_0),.clk(gclk));
	jdff dff_A_l0yD8ZRM2_0(.dout(w_dff_A_y02V02D96_0),.din(w_dff_A_l0yD8ZRM2_0),.clk(gclk));
	jdff dff_A_y02V02D96_0(.dout(w_dff_A_ycCJAbyC0_0),.din(w_dff_A_y02V02D96_0),.clk(gclk));
	jdff dff_A_ycCJAbyC0_0(.dout(w_dff_A_8ejQo4jA0_0),.din(w_dff_A_ycCJAbyC0_0),.clk(gclk));
	jdff dff_A_8ejQo4jA0_0(.dout(w_dff_A_ljXSKrKm8_0),.din(w_dff_A_8ejQo4jA0_0),.clk(gclk));
	jdff dff_A_ljXSKrKm8_0(.dout(w_dff_A_yAVcfKPP6_0),.din(w_dff_A_ljXSKrKm8_0),.clk(gclk));
	jdff dff_A_yAVcfKPP6_0(.dout(G422gat),.din(w_dff_A_yAVcfKPP6_0),.clk(gclk));
	jdff dff_A_EI1AbcoC2_2(.dout(w_dff_A_8JD0Pdk98_0),.din(w_dff_A_EI1AbcoC2_2),.clk(gclk));
	jdff dff_A_8JD0Pdk98_0(.dout(w_dff_A_osCCU1Yc0_0),.din(w_dff_A_8JD0Pdk98_0),.clk(gclk));
	jdff dff_A_osCCU1Yc0_0(.dout(w_dff_A_QiF03HjA7_0),.din(w_dff_A_osCCU1Yc0_0),.clk(gclk));
	jdff dff_A_QiF03HjA7_0(.dout(w_dff_A_Cl8U4e6d0_0),.din(w_dff_A_QiF03HjA7_0),.clk(gclk));
	jdff dff_A_Cl8U4e6d0_0(.dout(w_dff_A_X0ZFpbfj8_0),.din(w_dff_A_Cl8U4e6d0_0),.clk(gclk));
	jdff dff_A_X0ZFpbfj8_0(.dout(w_dff_A_QCHUAAkh1_0),.din(w_dff_A_X0ZFpbfj8_0),.clk(gclk));
	jdff dff_A_QCHUAAkh1_0(.dout(w_dff_A_tNR47FzG2_0),.din(w_dff_A_QCHUAAkh1_0),.clk(gclk));
	jdff dff_A_tNR47FzG2_0(.dout(w_dff_A_SEEB3kFx5_0),.din(w_dff_A_tNR47FzG2_0),.clk(gclk));
	jdff dff_A_SEEB3kFx5_0(.dout(w_dff_A_Wj5wxuFc3_0),.din(w_dff_A_SEEB3kFx5_0),.clk(gclk));
	jdff dff_A_Wj5wxuFc3_0(.dout(w_dff_A_7dVf7Ssj6_0),.din(w_dff_A_Wj5wxuFc3_0),.clk(gclk));
	jdff dff_A_7dVf7Ssj6_0(.dout(w_dff_A_wy33EccP1_0),.din(w_dff_A_7dVf7Ssj6_0),.clk(gclk));
	jdff dff_A_wy33EccP1_0(.dout(w_dff_A_vShCL3cO4_0),.din(w_dff_A_wy33EccP1_0),.clk(gclk));
	jdff dff_A_vShCL3cO4_0(.dout(w_dff_A_oj45jCHk3_0),.din(w_dff_A_vShCL3cO4_0),.clk(gclk));
	jdff dff_A_oj45jCHk3_0(.dout(w_dff_A_GM5B2vaZ3_0),.din(w_dff_A_oj45jCHk3_0),.clk(gclk));
	jdff dff_A_GM5B2vaZ3_0(.dout(w_dff_A_eonXjgxS2_0),.din(w_dff_A_GM5B2vaZ3_0),.clk(gclk));
	jdff dff_A_eonXjgxS2_0(.dout(w_dff_A_MxmfaX7b7_0),.din(w_dff_A_eonXjgxS2_0),.clk(gclk));
	jdff dff_A_MxmfaX7b7_0(.dout(w_dff_A_PGsUldvm8_0),.din(w_dff_A_MxmfaX7b7_0),.clk(gclk));
	jdff dff_A_PGsUldvm8_0(.dout(w_dff_A_iXOBFjoF4_0),.din(w_dff_A_PGsUldvm8_0),.clk(gclk));
	jdff dff_A_iXOBFjoF4_0(.dout(w_dff_A_Et2Sl7yz8_0),.din(w_dff_A_iXOBFjoF4_0),.clk(gclk));
	jdff dff_A_Et2Sl7yz8_0(.dout(w_dff_A_gXPrIarz7_0),.din(w_dff_A_Et2Sl7yz8_0),.clk(gclk));
	jdff dff_A_gXPrIarz7_0(.dout(w_dff_A_yJanGnWa1_0),.din(w_dff_A_gXPrIarz7_0),.clk(gclk));
	jdff dff_A_yJanGnWa1_0(.dout(w_dff_A_JU2DrTmE6_0),.din(w_dff_A_yJanGnWa1_0),.clk(gclk));
	jdff dff_A_JU2DrTmE6_0(.dout(w_dff_A_niZrNab53_0),.din(w_dff_A_JU2DrTmE6_0),.clk(gclk));
	jdff dff_A_niZrNab53_0(.dout(w_dff_A_yjBKcbmZ0_0),.din(w_dff_A_niZrNab53_0),.clk(gclk));
	jdff dff_A_yjBKcbmZ0_0(.dout(w_dff_A_V3bxT7gL2_0),.din(w_dff_A_yjBKcbmZ0_0),.clk(gclk));
	jdff dff_A_V3bxT7gL2_0(.dout(G423gat),.din(w_dff_A_V3bxT7gL2_0),.clk(gclk));
	jdff dff_A_O6jn1Gue3_2(.dout(w_dff_A_kgsD6hKS3_0),.din(w_dff_A_O6jn1Gue3_2),.clk(gclk));
	jdff dff_A_kgsD6hKS3_0(.dout(w_dff_A_5IvpyKGc3_0),.din(w_dff_A_kgsD6hKS3_0),.clk(gclk));
	jdff dff_A_5IvpyKGc3_0(.dout(w_dff_A_fu73RqIQ8_0),.din(w_dff_A_5IvpyKGc3_0),.clk(gclk));
	jdff dff_A_fu73RqIQ8_0(.dout(w_dff_A_X9OVA8s22_0),.din(w_dff_A_fu73RqIQ8_0),.clk(gclk));
	jdff dff_A_X9OVA8s22_0(.dout(w_dff_A_EZqJvrRG6_0),.din(w_dff_A_X9OVA8s22_0),.clk(gclk));
	jdff dff_A_EZqJvrRG6_0(.dout(w_dff_A_Rps1wixn1_0),.din(w_dff_A_EZqJvrRG6_0),.clk(gclk));
	jdff dff_A_Rps1wixn1_0(.dout(w_dff_A_r5whXDcm0_0),.din(w_dff_A_Rps1wixn1_0),.clk(gclk));
	jdff dff_A_r5whXDcm0_0(.dout(w_dff_A_oGwqlfyY7_0),.din(w_dff_A_r5whXDcm0_0),.clk(gclk));
	jdff dff_A_oGwqlfyY7_0(.dout(w_dff_A_f0kZlnSr0_0),.din(w_dff_A_oGwqlfyY7_0),.clk(gclk));
	jdff dff_A_f0kZlnSr0_0(.dout(w_dff_A_lUJL6bqw8_0),.din(w_dff_A_f0kZlnSr0_0),.clk(gclk));
	jdff dff_A_lUJL6bqw8_0(.dout(w_dff_A_lW3LOW715_0),.din(w_dff_A_lUJL6bqw8_0),.clk(gclk));
	jdff dff_A_lW3LOW715_0(.dout(w_dff_A_cIiEsxtk6_0),.din(w_dff_A_lW3LOW715_0),.clk(gclk));
	jdff dff_A_cIiEsxtk6_0(.dout(w_dff_A_5uFhLSaM2_0),.din(w_dff_A_cIiEsxtk6_0),.clk(gclk));
	jdff dff_A_5uFhLSaM2_0(.dout(w_dff_A_uqrlZ0w69_0),.din(w_dff_A_5uFhLSaM2_0),.clk(gclk));
	jdff dff_A_uqrlZ0w69_0(.dout(w_dff_A_aUBDG2uL6_0),.din(w_dff_A_uqrlZ0w69_0),.clk(gclk));
	jdff dff_A_aUBDG2uL6_0(.dout(w_dff_A_ovWTiWeL1_0),.din(w_dff_A_aUBDG2uL6_0),.clk(gclk));
	jdff dff_A_ovWTiWeL1_0(.dout(w_dff_A_uDPFbiSV5_0),.din(w_dff_A_ovWTiWeL1_0),.clk(gclk));
	jdff dff_A_uDPFbiSV5_0(.dout(w_dff_A_PFnYDDsh9_0),.din(w_dff_A_uDPFbiSV5_0),.clk(gclk));
	jdff dff_A_PFnYDDsh9_0(.dout(w_dff_A_LyxSbZFw9_0),.din(w_dff_A_PFnYDDsh9_0),.clk(gclk));
	jdff dff_A_LyxSbZFw9_0(.dout(w_dff_A_6auhD7d33_0),.din(w_dff_A_LyxSbZFw9_0),.clk(gclk));
	jdff dff_A_6auhD7d33_0(.dout(w_dff_A_gK4yLJSg5_0),.din(w_dff_A_6auhD7d33_0),.clk(gclk));
	jdff dff_A_gK4yLJSg5_0(.dout(w_dff_A_NFlCp7eI0_0),.din(w_dff_A_gK4yLJSg5_0),.clk(gclk));
	jdff dff_A_NFlCp7eI0_0(.dout(G446gat),.din(w_dff_A_NFlCp7eI0_0),.clk(gclk));
	jdff dff_A_bDsVM3Cz7_1(.dout(w_dff_A_BEa6ECR94_0),.din(w_dff_A_bDsVM3Cz7_1),.clk(gclk));
	jdff dff_A_BEa6ECR94_0(.dout(w_dff_A_j8BSzuoO5_0),.din(w_dff_A_BEa6ECR94_0),.clk(gclk));
	jdff dff_A_j8BSzuoO5_0(.dout(w_dff_A_wqewGXlq4_0),.din(w_dff_A_j8BSzuoO5_0),.clk(gclk));
	jdff dff_A_wqewGXlq4_0(.dout(w_dff_A_Xrjtlo7x2_0),.din(w_dff_A_wqewGXlq4_0),.clk(gclk));
	jdff dff_A_Xrjtlo7x2_0(.dout(w_dff_A_JygVPBNZ0_0),.din(w_dff_A_Xrjtlo7x2_0),.clk(gclk));
	jdff dff_A_JygVPBNZ0_0(.dout(w_dff_A_4gQ4kPKd2_0),.din(w_dff_A_JygVPBNZ0_0),.clk(gclk));
	jdff dff_A_4gQ4kPKd2_0(.dout(w_dff_A_UjBAK97Z1_0),.din(w_dff_A_4gQ4kPKd2_0),.clk(gclk));
	jdff dff_A_UjBAK97Z1_0(.dout(w_dff_A_v6i9W8d93_0),.din(w_dff_A_UjBAK97Z1_0),.clk(gclk));
	jdff dff_A_v6i9W8d93_0(.dout(w_dff_A_dReMKxeq8_0),.din(w_dff_A_v6i9W8d93_0),.clk(gclk));
	jdff dff_A_dReMKxeq8_0(.dout(w_dff_A_hBzNvfgR7_0),.din(w_dff_A_dReMKxeq8_0),.clk(gclk));
	jdff dff_A_hBzNvfgR7_0(.dout(w_dff_A_9IfKUUth2_0),.din(w_dff_A_hBzNvfgR7_0),.clk(gclk));
	jdff dff_A_9IfKUUth2_0(.dout(w_dff_A_ecr7qeEJ3_0),.din(w_dff_A_9IfKUUth2_0),.clk(gclk));
	jdff dff_A_ecr7qeEJ3_0(.dout(w_dff_A_vfAaOUuf3_0),.din(w_dff_A_ecr7qeEJ3_0),.clk(gclk));
	jdff dff_A_vfAaOUuf3_0(.dout(w_dff_A_r5YP6lXY8_0),.din(w_dff_A_vfAaOUuf3_0),.clk(gclk));
	jdff dff_A_r5YP6lXY8_0(.dout(w_dff_A_83NxtOxK1_0),.din(w_dff_A_r5YP6lXY8_0),.clk(gclk));
	jdff dff_A_83NxtOxK1_0(.dout(w_dff_A_ee9mZmBx6_0),.din(w_dff_A_83NxtOxK1_0),.clk(gclk));
	jdff dff_A_ee9mZmBx6_0(.dout(w_dff_A_QXu8jWsX3_0),.din(w_dff_A_ee9mZmBx6_0),.clk(gclk));
	jdff dff_A_QXu8jWsX3_0(.dout(w_dff_A_AKZURNN02_0),.din(w_dff_A_QXu8jWsX3_0),.clk(gclk));
	jdff dff_A_AKZURNN02_0(.dout(w_dff_A_WvwA8LiT6_0),.din(w_dff_A_AKZURNN02_0),.clk(gclk));
	jdff dff_A_WvwA8LiT6_0(.dout(w_dff_A_Krl3ZUX24_0),.din(w_dff_A_WvwA8LiT6_0),.clk(gclk));
	jdff dff_A_Krl3ZUX24_0(.dout(w_dff_A_bPIcYI5T0_0),.din(w_dff_A_Krl3ZUX24_0),.clk(gclk));
	jdff dff_A_bPIcYI5T0_0(.dout(w_dff_A_6iYzJI2M5_0),.din(w_dff_A_bPIcYI5T0_0),.clk(gclk));
	jdff dff_A_6iYzJI2M5_0(.dout(w_dff_A_YCHX3iBi0_0),.din(w_dff_A_6iYzJI2M5_0),.clk(gclk));
	jdff dff_A_YCHX3iBi0_0(.dout(w_dff_A_Ptv9l8jB6_0),.din(w_dff_A_YCHX3iBi0_0),.clk(gclk));
	jdff dff_A_Ptv9l8jB6_0(.dout(w_dff_A_JveD93U55_0),.din(w_dff_A_Ptv9l8jB6_0),.clk(gclk));
	jdff dff_A_JveD93U55_0(.dout(G447gat),.din(w_dff_A_JveD93U55_0),.clk(gclk));
	jdff dff_A_d7DwcygA1_2(.dout(w_dff_A_MhstYeIf3_0),.din(w_dff_A_d7DwcygA1_2),.clk(gclk));
	jdff dff_A_MhstYeIf3_0(.dout(w_dff_A_Yl5exmZf3_0),.din(w_dff_A_MhstYeIf3_0),.clk(gclk));
	jdff dff_A_Yl5exmZf3_0(.dout(w_dff_A_72IKoJsn0_0),.din(w_dff_A_Yl5exmZf3_0),.clk(gclk));
	jdff dff_A_72IKoJsn0_0(.dout(w_dff_A_6PQ7w8RY1_0),.din(w_dff_A_72IKoJsn0_0),.clk(gclk));
	jdff dff_A_6PQ7w8RY1_0(.dout(w_dff_A_8RtDEWQX2_0),.din(w_dff_A_6PQ7w8RY1_0),.clk(gclk));
	jdff dff_A_8RtDEWQX2_0(.dout(w_dff_A_LcxT1DII1_0),.din(w_dff_A_8RtDEWQX2_0),.clk(gclk));
	jdff dff_A_LcxT1DII1_0(.dout(w_dff_A_zM3QRekq3_0),.din(w_dff_A_LcxT1DII1_0),.clk(gclk));
	jdff dff_A_zM3QRekq3_0(.dout(w_dff_A_Md0LfRkU8_0),.din(w_dff_A_zM3QRekq3_0),.clk(gclk));
	jdff dff_A_Md0LfRkU8_0(.dout(w_dff_A_yII40mDR7_0),.din(w_dff_A_Md0LfRkU8_0),.clk(gclk));
	jdff dff_A_yII40mDR7_0(.dout(w_dff_A_3wsZMJIN8_0),.din(w_dff_A_yII40mDR7_0),.clk(gclk));
	jdff dff_A_3wsZMJIN8_0(.dout(w_dff_A_mdki67i10_0),.din(w_dff_A_3wsZMJIN8_0),.clk(gclk));
	jdff dff_A_mdki67i10_0(.dout(w_dff_A_K6ykE9Es0_0),.din(w_dff_A_mdki67i10_0),.clk(gclk));
	jdff dff_A_K6ykE9Es0_0(.dout(w_dff_A_S4xidspa6_0),.din(w_dff_A_K6ykE9Es0_0),.clk(gclk));
	jdff dff_A_S4xidspa6_0(.dout(w_dff_A_KSV1Dyqt8_0),.din(w_dff_A_S4xidspa6_0),.clk(gclk));
	jdff dff_A_KSV1Dyqt8_0(.dout(w_dff_A_8dZ3D4dc2_0),.din(w_dff_A_KSV1Dyqt8_0),.clk(gclk));
	jdff dff_A_8dZ3D4dc2_0(.dout(w_dff_A_U2k9AOlS6_0),.din(w_dff_A_8dZ3D4dc2_0),.clk(gclk));
	jdff dff_A_U2k9AOlS6_0(.dout(w_dff_A_um8nsU6v7_0),.din(w_dff_A_U2k9AOlS6_0),.clk(gclk));
	jdff dff_A_um8nsU6v7_0(.dout(w_dff_A_VdSaoWRT1_0),.din(w_dff_A_um8nsU6v7_0),.clk(gclk));
	jdff dff_A_VdSaoWRT1_0(.dout(w_dff_A_Q3xRzlFV7_0),.din(w_dff_A_VdSaoWRT1_0),.clk(gclk));
	jdff dff_A_Q3xRzlFV7_0(.dout(w_dff_A_EJJpLg9J1_0),.din(w_dff_A_Q3xRzlFV7_0),.clk(gclk));
	jdff dff_A_EJJpLg9J1_0(.dout(w_dff_A_07fLWie52_0),.din(w_dff_A_EJJpLg9J1_0),.clk(gclk));
	jdff dff_A_07fLWie52_0(.dout(w_dff_A_eu2X2mip2_0),.din(w_dff_A_07fLWie52_0),.clk(gclk));
	jdff dff_A_eu2X2mip2_0(.dout(G448gat),.din(w_dff_A_eu2X2mip2_0),.clk(gclk));
	jdff dff_A_VbVzM2jM1_2(.dout(w_dff_A_CgoddBim3_0),.din(w_dff_A_VbVzM2jM1_2),.clk(gclk));
	jdff dff_A_CgoddBim3_0(.dout(w_dff_A_Jgo03Sv45_0),.din(w_dff_A_CgoddBim3_0),.clk(gclk));
	jdff dff_A_Jgo03Sv45_0(.dout(w_dff_A_wFDivU5a4_0),.din(w_dff_A_Jgo03Sv45_0),.clk(gclk));
	jdff dff_A_wFDivU5a4_0(.dout(w_dff_A_ZwYGWjRz5_0),.din(w_dff_A_wFDivU5a4_0),.clk(gclk));
	jdff dff_A_ZwYGWjRz5_0(.dout(w_dff_A_50WfZlRv9_0),.din(w_dff_A_ZwYGWjRz5_0),.clk(gclk));
	jdff dff_A_50WfZlRv9_0(.dout(w_dff_A_HtYxp3CU8_0),.din(w_dff_A_50WfZlRv9_0),.clk(gclk));
	jdff dff_A_HtYxp3CU8_0(.dout(w_dff_A_GvkBVEZY7_0),.din(w_dff_A_HtYxp3CU8_0),.clk(gclk));
	jdff dff_A_GvkBVEZY7_0(.dout(w_dff_A_B5NMwLW42_0),.din(w_dff_A_GvkBVEZY7_0),.clk(gclk));
	jdff dff_A_B5NMwLW42_0(.dout(w_dff_A_ZEsUSQyw7_0),.din(w_dff_A_B5NMwLW42_0),.clk(gclk));
	jdff dff_A_ZEsUSQyw7_0(.dout(w_dff_A_xuXfIYyy9_0),.din(w_dff_A_ZEsUSQyw7_0),.clk(gclk));
	jdff dff_A_xuXfIYyy9_0(.dout(w_dff_A_3qJoRJzD0_0),.din(w_dff_A_xuXfIYyy9_0),.clk(gclk));
	jdff dff_A_3qJoRJzD0_0(.dout(w_dff_A_HFBl8UVZ8_0),.din(w_dff_A_3qJoRJzD0_0),.clk(gclk));
	jdff dff_A_HFBl8UVZ8_0(.dout(w_dff_A_AggPnzlb1_0),.din(w_dff_A_HFBl8UVZ8_0),.clk(gclk));
	jdff dff_A_AggPnzlb1_0(.dout(w_dff_A_z9iQBznL7_0),.din(w_dff_A_AggPnzlb1_0),.clk(gclk));
	jdff dff_A_z9iQBznL7_0(.dout(w_dff_A_rqYgT0Dl0_0),.din(w_dff_A_z9iQBznL7_0),.clk(gclk));
	jdff dff_A_rqYgT0Dl0_0(.dout(w_dff_A_Vnn3D59h3_0),.din(w_dff_A_rqYgT0Dl0_0),.clk(gclk));
	jdff dff_A_Vnn3D59h3_0(.dout(w_dff_A_fVFkq9qw8_0),.din(w_dff_A_Vnn3D59h3_0),.clk(gclk));
	jdff dff_A_fVFkq9qw8_0(.dout(w_dff_A_gvAHydQ76_0),.din(w_dff_A_fVFkq9qw8_0),.clk(gclk));
	jdff dff_A_gvAHydQ76_0(.dout(w_dff_A_4N8IUoXA7_0),.din(w_dff_A_gvAHydQ76_0),.clk(gclk));
	jdff dff_A_4N8IUoXA7_0(.dout(w_dff_A_AqquzEvy1_0),.din(w_dff_A_4N8IUoXA7_0),.clk(gclk));
	jdff dff_A_AqquzEvy1_0(.dout(w_dff_A_Retbe4sH3_0),.din(w_dff_A_AqquzEvy1_0),.clk(gclk));
	jdff dff_A_Retbe4sH3_0(.dout(w_dff_A_4P6xKnKW5_0),.din(w_dff_A_Retbe4sH3_0),.clk(gclk));
	jdff dff_A_4P6xKnKW5_0(.dout(G449gat),.din(w_dff_A_4P6xKnKW5_0),.clk(gclk));
	jdff dff_A_46oFJh5I3_2(.dout(w_dff_A_C0PghwRv6_0),.din(w_dff_A_46oFJh5I3_2),.clk(gclk));
	jdff dff_A_C0PghwRv6_0(.dout(w_dff_A_wgptwsmK8_0),.din(w_dff_A_C0PghwRv6_0),.clk(gclk));
	jdff dff_A_wgptwsmK8_0(.dout(w_dff_A_9jwx3rml7_0),.din(w_dff_A_wgptwsmK8_0),.clk(gclk));
	jdff dff_A_9jwx3rml7_0(.dout(w_dff_A_JdOCm0dx1_0),.din(w_dff_A_9jwx3rml7_0),.clk(gclk));
	jdff dff_A_JdOCm0dx1_0(.dout(w_dff_A_MLGMIGu43_0),.din(w_dff_A_JdOCm0dx1_0),.clk(gclk));
	jdff dff_A_MLGMIGu43_0(.dout(w_dff_A_8B4y4y9K3_0),.din(w_dff_A_MLGMIGu43_0),.clk(gclk));
	jdff dff_A_8B4y4y9K3_0(.dout(w_dff_A_pkjTEZjv2_0),.din(w_dff_A_8B4y4y9K3_0),.clk(gclk));
	jdff dff_A_pkjTEZjv2_0(.dout(w_dff_A_Ml5hqJBm4_0),.din(w_dff_A_pkjTEZjv2_0),.clk(gclk));
	jdff dff_A_Ml5hqJBm4_0(.dout(w_dff_A_q6NT3oCv1_0),.din(w_dff_A_Ml5hqJBm4_0),.clk(gclk));
	jdff dff_A_q6NT3oCv1_0(.dout(w_dff_A_pgP4yugU0_0),.din(w_dff_A_q6NT3oCv1_0),.clk(gclk));
	jdff dff_A_pgP4yugU0_0(.dout(w_dff_A_qd0YjtjN5_0),.din(w_dff_A_pgP4yugU0_0),.clk(gclk));
	jdff dff_A_qd0YjtjN5_0(.dout(w_dff_A_hQgmV7lM8_0),.din(w_dff_A_qd0YjtjN5_0),.clk(gclk));
	jdff dff_A_hQgmV7lM8_0(.dout(w_dff_A_COVMCks73_0),.din(w_dff_A_hQgmV7lM8_0),.clk(gclk));
	jdff dff_A_COVMCks73_0(.dout(w_dff_A_uISI1WsD5_0),.din(w_dff_A_COVMCks73_0),.clk(gclk));
	jdff dff_A_uISI1WsD5_0(.dout(w_dff_A_QikJSJ3d1_0),.din(w_dff_A_uISI1WsD5_0),.clk(gclk));
	jdff dff_A_QikJSJ3d1_0(.dout(w_dff_A_4c9L0DV80_0),.din(w_dff_A_QikJSJ3d1_0),.clk(gclk));
	jdff dff_A_4c9L0DV80_0(.dout(w_dff_A_0RQkebOo9_0),.din(w_dff_A_4c9L0DV80_0),.clk(gclk));
	jdff dff_A_0RQkebOo9_0(.dout(w_dff_A_2vQiqEB96_0),.din(w_dff_A_0RQkebOo9_0),.clk(gclk));
	jdff dff_A_2vQiqEB96_0(.dout(w_dff_A_YaBG4oSU9_0),.din(w_dff_A_2vQiqEB96_0),.clk(gclk));
	jdff dff_A_YaBG4oSU9_0(.dout(w_dff_A_MdzUCVzI6_0),.din(w_dff_A_YaBG4oSU9_0),.clk(gclk));
	jdff dff_A_MdzUCVzI6_0(.dout(w_dff_A_lQ1dH66v6_0),.din(w_dff_A_MdzUCVzI6_0),.clk(gclk));
	jdff dff_A_lQ1dH66v6_0(.dout(w_dff_A_QMKe07Im0_0),.din(w_dff_A_lQ1dH66v6_0),.clk(gclk));
	jdff dff_A_QMKe07Im0_0(.dout(w_dff_A_McwYecOY1_0),.din(w_dff_A_QMKe07Im0_0),.clk(gclk));
	jdff dff_A_McwYecOY1_0(.dout(w_dff_A_D604cKvP7_0),.din(w_dff_A_McwYecOY1_0),.clk(gclk));
	jdff dff_A_D604cKvP7_0(.dout(w_dff_A_vyrLqLGJ4_0),.din(w_dff_A_D604cKvP7_0),.clk(gclk));
	jdff dff_A_vyrLqLGJ4_0(.dout(G450gat),.din(w_dff_A_vyrLqLGJ4_0),.clk(gclk));
	jdff dff_A_U7erAsDQ5_2(.dout(w_dff_A_TM5MgPuX3_0),.din(w_dff_A_U7erAsDQ5_2),.clk(gclk));
	jdff dff_A_TM5MgPuX3_0(.dout(w_dff_A_Mz9qLphq2_0),.din(w_dff_A_TM5MgPuX3_0),.clk(gclk));
	jdff dff_A_Mz9qLphq2_0(.dout(w_dff_A_2As3Gp9u4_0),.din(w_dff_A_Mz9qLphq2_0),.clk(gclk));
	jdff dff_A_2As3Gp9u4_0(.dout(w_dff_A_vXcrQt8P2_0),.din(w_dff_A_2As3Gp9u4_0),.clk(gclk));
	jdff dff_A_vXcrQt8P2_0(.dout(w_dff_A_yrZBHJd72_0),.din(w_dff_A_vXcrQt8P2_0),.clk(gclk));
	jdff dff_A_yrZBHJd72_0(.dout(w_dff_A_HDSOKIyw3_0),.din(w_dff_A_yrZBHJd72_0),.clk(gclk));
	jdff dff_A_HDSOKIyw3_0(.dout(w_dff_A_dA3HrudG7_0),.din(w_dff_A_HDSOKIyw3_0),.clk(gclk));
	jdff dff_A_dA3HrudG7_0(.dout(w_dff_A_oSp4Wycw9_0),.din(w_dff_A_dA3HrudG7_0),.clk(gclk));
	jdff dff_A_oSp4Wycw9_0(.dout(w_dff_A_l10DnAiv7_0),.din(w_dff_A_oSp4Wycw9_0),.clk(gclk));
	jdff dff_A_l10DnAiv7_0(.dout(w_dff_A_zCXOxBdL0_0),.din(w_dff_A_l10DnAiv7_0),.clk(gclk));
	jdff dff_A_zCXOxBdL0_0(.dout(w_dff_A_mgNFwFQI6_0),.din(w_dff_A_zCXOxBdL0_0),.clk(gclk));
	jdff dff_A_mgNFwFQI6_0(.dout(w_dff_A_KL22KnRp0_0),.din(w_dff_A_mgNFwFQI6_0),.clk(gclk));
	jdff dff_A_KL22KnRp0_0(.dout(w_dff_A_M4wox5Ln1_0),.din(w_dff_A_KL22KnRp0_0),.clk(gclk));
	jdff dff_A_M4wox5Ln1_0(.dout(w_dff_A_lKvVqxvf2_0),.din(w_dff_A_M4wox5Ln1_0),.clk(gclk));
	jdff dff_A_lKvVqxvf2_0(.dout(w_dff_A_VtjWYBoD7_0),.din(w_dff_A_lKvVqxvf2_0),.clk(gclk));
	jdff dff_A_VtjWYBoD7_0(.dout(w_dff_A_nRN3mXyO0_0),.din(w_dff_A_VtjWYBoD7_0),.clk(gclk));
	jdff dff_A_nRN3mXyO0_0(.dout(w_dff_A_f4YfKqPQ5_0),.din(w_dff_A_nRN3mXyO0_0),.clk(gclk));
	jdff dff_A_f4YfKqPQ5_0(.dout(w_dff_A_lJZCFmRb2_0),.din(w_dff_A_f4YfKqPQ5_0),.clk(gclk));
	jdff dff_A_lJZCFmRb2_0(.dout(w_dff_A_4cghf02G5_0),.din(w_dff_A_lJZCFmRb2_0),.clk(gclk));
	jdff dff_A_4cghf02G5_0(.dout(w_dff_A_zayDYMAC9_0),.din(w_dff_A_4cghf02G5_0),.clk(gclk));
	jdff dff_A_zayDYMAC9_0(.dout(w_dff_A_MhpwNvY03_0),.din(w_dff_A_zayDYMAC9_0),.clk(gclk));
	jdff dff_A_MhpwNvY03_0(.dout(w_dff_A_pRnNxhi55_0),.din(w_dff_A_MhpwNvY03_0),.clk(gclk));
	jdff dff_A_pRnNxhi55_0(.dout(w_dff_A_GaIMETuo0_0),.din(w_dff_A_pRnNxhi55_0),.clk(gclk));
	jdff dff_A_GaIMETuo0_0(.dout(G767gat),.din(w_dff_A_GaIMETuo0_0),.clk(gclk));
	jdff dff_A_kFURueqb2_2(.dout(w_dff_A_tfJCnvsX0_0),.din(w_dff_A_kFURueqb2_2),.clk(gclk));
	jdff dff_A_tfJCnvsX0_0(.dout(w_dff_A_4MHuud4Z4_0),.din(w_dff_A_tfJCnvsX0_0),.clk(gclk));
	jdff dff_A_4MHuud4Z4_0(.dout(w_dff_A_rFqSc2Fp3_0),.din(w_dff_A_4MHuud4Z4_0),.clk(gclk));
	jdff dff_A_rFqSc2Fp3_0(.dout(w_dff_A_0sGc09mi4_0),.din(w_dff_A_rFqSc2Fp3_0),.clk(gclk));
	jdff dff_A_0sGc09mi4_0(.dout(w_dff_A_COMTXygF4_0),.din(w_dff_A_0sGc09mi4_0),.clk(gclk));
	jdff dff_A_COMTXygF4_0(.dout(w_dff_A_pHqeztw50_0),.din(w_dff_A_COMTXygF4_0),.clk(gclk));
	jdff dff_A_pHqeztw50_0(.dout(w_dff_A_R7Y3MG942_0),.din(w_dff_A_pHqeztw50_0),.clk(gclk));
	jdff dff_A_R7Y3MG942_0(.dout(w_dff_A_xRYGPthN0_0),.din(w_dff_A_R7Y3MG942_0),.clk(gclk));
	jdff dff_A_xRYGPthN0_0(.dout(w_dff_A_M4Z4rDQt2_0),.din(w_dff_A_xRYGPthN0_0),.clk(gclk));
	jdff dff_A_M4Z4rDQt2_0(.dout(w_dff_A_kFyR0jOj6_0),.din(w_dff_A_M4Z4rDQt2_0),.clk(gclk));
	jdff dff_A_kFyR0jOj6_0(.dout(w_dff_A_DyDUDH0p4_0),.din(w_dff_A_kFyR0jOj6_0),.clk(gclk));
	jdff dff_A_DyDUDH0p4_0(.dout(w_dff_A_xqnlnMaR6_0),.din(w_dff_A_DyDUDH0p4_0),.clk(gclk));
	jdff dff_A_xqnlnMaR6_0(.dout(w_dff_A_rJVwUmKk0_0),.din(w_dff_A_xqnlnMaR6_0),.clk(gclk));
	jdff dff_A_rJVwUmKk0_0(.dout(w_dff_A_qRogF6Ix9_0),.din(w_dff_A_rJVwUmKk0_0),.clk(gclk));
	jdff dff_A_qRogF6Ix9_0(.dout(w_dff_A_IJZegaBq5_0),.din(w_dff_A_qRogF6Ix9_0),.clk(gclk));
	jdff dff_A_IJZegaBq5_0(.dout(w_dff_A_uq1pQA367_0),.din(w_dff_A_IJZegaBq5_0),.clk(gclk));
	jdff dff_A_uq1pQA367_0(.dout(w_dff_A_2vWaFgIl2_0),.din(w_dff_A_uq1pQA367_0),.clk(gclk));
	jdff dff_A_2vWaFgIl2_0(.dout(w_dff_A_1TKF6j2i2_0),.din(w_dff_A_2vWaFgIl2_0),.clk(gclk));
	jdff dff_A_1TKF6j2i2_0(.dout(w_dff_A_Kankvch38_0),.din(w_dff_A_1TKF6j2i2_0),.clk(gclk));
	jdff dff_A_Kankvch38_0(.dout(w_dff_A_f6YJmiCl1_0),.din(w_dff_A_Kankvch38_0),.clk(gclk));
	jdff dff_A_f6YJmiCl1_0(.dout(w_dff_A_ikFvfpAo1_0),.din(w_dff_A_f6YJmiCl1_0),.clk(gclk));
	jdff dff_A_ikFvfpAo1_0(.dout(w_dff_A_MyBrPLSD4_0),.din(w_dff_A_ikFvfpAo1_0),.clk(gclk));
	jdff dff_A_MyBrPLSD4_0(.dout(w_dff_A_154bAPmV3_0),.din(w_dff_A_MyBrPLSD4_0),.clk(gclk));
	jdff dff_A_154bAPmV3_0(.dout(G768gat),.din(w_dff_A_154bAPmV3_0),.clk(gclk));
	jdff dff_A_0bei3kWP7_2(.dout(w_dff_A_FW3tNPOQ3_0),.din(w_dff_A_0bei3kWP7_2),.clk(gclk));
	jdff dff_A_FW3tNPOQ3_0(.dout(w_dff_A_p3rjj3bx0_0),.din(w_dff_A_FW3tNPOQ3_0),.clk(gclk));
	jdff dff_A_p3rjj3bx0_0(.dout(w_dff_A_DDv9Ri6O3_0),.din(w_dff_A_p3rjj3bx0_0),.clk(gclk));
	jdff dff_A_DDv9Ri6O3_0(.dout(w_dff_A_7AnUinVD1_0),.din(w_dff_A_DDv9Ri6O3_0),.clk(gclk));
	jdff dff_A_7AnUinVD1_0(.dout(w_dff_A_BjlvJ0cv9_0),.din(w_dff_A_7AnUinVD1_0),.clk(gclk));
	jdff dff_A_BjlvJ0cv9_0(.dout(w_dff_A_RDyqs1ny6_0),.din(w_dff_A_BjlvJ0cv9_0),.clk(gclk));
	jdff dff_A_RDyqs1ny6_0(.dout(w_dff_A_0sjJb1qh1_0),.din(w_dff_A_RDyqs1ny6_0),.clk(gclk));
	jdff dff_A_0sjJb1qh1_0(.dout(w_dff_A_SC86Nwwo5_0),.din(w_dff_A_0sjJb1qh1_0),.clk(gclk));
	jdff dff_A_SC86Nwwo5_0(.dout(w_dff_A_2TSW3xlc0_0),.din(w_dff_A_SC86Nwwo5_0),.clk(gclk));
	jdff dff_A_2TSW3xlc0_0(.dout(w_dff_A_Q8RntV027_0),.din(w_dff_A_2TSW3xlc0_0),.clk(gclk));
	jdff dff_A_Q8RntV027_0(.dout(w_dff_A_zisxz3fN4_0),.din(w_dff_A_Q8RntV027_0),.clk(gclk));
	jdff dff_A_zisxz3fN4_0(.dout(w_dff_A_z2UgFbIY1_0),.din(w_dff_A_zisxz3fN4_0),.clk(gclk));
	jdff dff_A_z2UgFbIY1_0(.dout(G850gat),.din(w_dff_A_z2UgFbIY1_0),.clk(gclk));
	jdff dff_A_kOlKxf7O4_2(.dout(w_dff_A_WifP3QV35_0),.din(w_dff_A_kOlKxf7O4_2),.clk(gclk));
	jdff dff_A_WifP3QV35_0(.dout(w_dff_A_rCvrwCWK4_0),.din(w_dff_A_WifP3QV35_0),.clk(gclk));
	jdff dff_A_rCvrwCWK4_0(.dout(w_dff_A_tWQhGJB15_0),.din(w_dff_A_rCvrwCWK4_0),.clk(gclk));
	jdff dff_A_tWQhGJB15_0(.dout(w_dff_A_iJBFqXoD7_0),.din(w_dff_A_tWQhGJB15_0),.clk(gclk));
	jdff dff_A_iJBFqXoD7_0(.dout(w_dff_A_FIPprnkS9_0),.din(w_dff_A_iJBFqXoD7_0),.clk(gclk));
	jdff dff_A_FIPprnkS9_0(.dout(w_dff_A_o0Ti0cIn1_0),.din(w_dff_A_FIPprnkS9_0),.clk(gclk));
	jdff dff_A_o0Ti0cIn1_0(.dout(w_dff_A_bfi6CDsu0_0),.din(w_dff_A_o0Ti0cIn1_0),.clk(gclk));
	jdff dff_A_bfi6CDsu0_0(.dout(G863gat),.din(w_dff_A_bfi6CDsu0_0),.clk(gclk));
	jdff dff_A_EaLwtXtj9_2(.dout(w_dff_A_Yw8WOXeD3_0),.din(w_dff_A_EaLwtXtj9_2),.clk(gclk));
	jdff dff_A_Yw8WOXeD3_0(.dout(w_dff_A_rihFLxqu4_0),.din(w_dff_A_Yw8WOXeD3_0),.clk(gclk));
	jdff dff_A_rihFLxqu4_0(.dout(w_dff_A_Kl7a5jAB0_0),.din(w_dff_A_rihFLxqu4_0),.clk(gclk));
	jdff dff_A_Kl7a5jAB0_0(.dout(w_dff_A_pCjPIYbn1_0),.din(w_dff_A_Kl7a5jAB0_0),.clk(gclk));
	jdff dff_A_pCjPIYbn1_0(.dout(w_dff_A_gWtLxFGp7_0),.din(w_dff_A_pCjPIYbn1_0),.clk(gclk));
	jdff dff_A_gWtLxFGp7_0(.dout(w_dff_A_8iMkopc76_0),.din(w_dff_A_gWtLxFGp7_0),.clk(gclk));
	jdff dff_A_8iMkopc76_0(.dout(w_dff_A_luZJ4B4N8_0),.din(w_dff_A_8iMkopc76_0),.clk(gclk));
	jdff dff_A_luZJ4B4N8_0(.dout(w_dff_A_CZ2WFe3r6_0),.din(w_dff_A_luZJ4B4N8_0),.clk(gclk));
	jdff dff_A_CZ2WFe3r6_0(.dout(w_dff_A_a8gxr0EZ7_0),.din(w_dff_A_CZ2WFe3r6_0),.clk(gclk));
	jdff dff_A_a8gxr0EZ7_0(.dout(G864gat),.din(w_dff_A_a8gxr0EZ7_0),.clk(gclk));
	jdff dff_A_i7fpZ1qg5_2(.dout(w_dff_A_rvjWJORW9_0),.din(w_dff_A_i7fpZ1qg5_2),.clk(gclk));
	jdff dff_A_rvjWJORW9_0(.dout(w_dff_A_T2UfIs6M5_0),.din(w_dff_A_rvjWJORW9_0),.clk(gclk));
	jdff dff_A_T2UfIs6M5_0(.dout(w_dff_A_nAlhdSUP5_0),.din(w_dff_A_T2UfIs6M5_0),.clk(gclk));
	jdff dff_A_nAlhdSUP5_0(.dout(w_dff_A_xvs9Erk25_0),.din(w_dff_A_nAlhdSUP5_0),.clk(gclk));
	jdff dff_A_xvs9Erk25_0(.dout(w_dff_A_UxxXG8wq0_0),.din(w_dff_A_xvs9Erk25_0),.clk(gclk));
	jdff dff_A_UxxXG8wq0_0(.dout(w_dff_A_IulKnn1f1_0),.din(w_dff_A_UxxXG8wq0_0),.clk(gclk));
	jdff dff_A_IulKnn1f1_0(.dout(w_dff_A_1sEohxXZ4_0),.din(w_dff_A_IulKnn1f1_0),.clk(gclk));
	jdff dff_A_1sEohxXZ4_0(.dout(w_dff_A_OKY0dIbs7_0),.din(w_dff_A_1sEohxXZ4_0),.clk(gclk));
	jdff dff_A_OKY0dIbs7_0(.dout(w_dff_A_VdkCCeHd8_0),.din(w_dff_A_OKY0dIbs7_0),.clk(gclk));
	jdff dff_A_VdkCCeHd8_0(.dout(w_dff_A_vdT0ciDk9_0),.din(w_dff_A_VdkCCeHd8_0),.clk(gclk));
	jdff dff_A_vdT0ciDk9_0(.dout(w_dff_A_OWy0ZP7R1_0),.din(w_dff_A_vdT0ciDk9_0),.clk(gclk));
	jdff dff_A_OWy0ZP7R1_0(.dout(G865gat),.din(w_dff_A_OWy0ZP7R1_0),.clk(gclk));
	jdff dff_A_uu90gjxu6_2(.dout(w_dff_A_TgbimvxW0_0),.din(w_dff_A_uu90gjxu6_2),.clk(gclk));
	jdff dff_A_TgbimvxW0_0(.dout(G866gat),.din(w_dff_A_TgbimvxW0_0),.clk(gclk));
	jdff dff_A_59cdx3DS7_2(.dout(w_dff_A_HlFeHme37_0),.din(w_dff_A_59cdx3DS7_2),.clk(gclk));
	jdff dff_A_HlFeHme37_0(.dout(w_dff_A_Qci0cMBR4_0),.din(w_dff_A_HlFeHme37_0),.clk(gclk));
	jdff dff_A_Qci0cMBR4_0(.dout(w_dff_A_t0q54zPC0_0),.din(w_dff_A_Qci0cMBR4_0),.clk(gclk));
	jdff dff_A_t0q54zPC0_0(.dout(w_dff_A_k6q6b7sE7_0),.din(w_dff_A_t0q54zPC0_0),.clk(gclk));
	jdff dff_A_k6q6b7sE7_0(.dout(G874gat),.din(w_dff_A_k6q6b7sE7_0),.clk(gclk));
	jdff dff_A_j2wVWtWp7_2(.dout(w_dff_A_peHDjjEc4_0),.din(w_dff_A_j2wVWtWp7_2),.clk(gclk));
	jdff dff_A_peHDjjEc4_0(.dout(G879gat),.din(w_dff_A_peHDjjEc4_0),.clk(gclk));
	jdff dff_A_yvuvlarN9_2(.dout(w_dff_A_hKsJVxjJ0_0),.din(w_dff_A_yvuvlarN9_2),.clk(gclk));
	jdff dff_A_hKsJVxjJ0_0(.dout(w_dff_A_ToHw2GrJ1_0),.din(w_dff_A_hKsJVxjJ0_0),.clk(gclk));
	jdff dff_A_ToHw2GrJ1_0(.dout(w_dff_A_RrvOc9bb9_0),.din(w_dff_A_ToHw2GrJ1_0),.clk(gclk));
	jdff dff_A_RrvOc9bb9_0(.dout(G880gat),.din(w_dff_A_RrvOc9bb9_0),.clk(gclk));
endmodule

