/*

c1355:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 509
	jand: 65
	jor: 6

Summary:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 509
	jand: 65
	jor: 6
*/

module c1355(gclk, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat, G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat, G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat, G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat, G1352gat, G1353gat, G1354gat, G1355gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G15gat;
	input G22gat;
	input G29gat;
	input G36gat;
	input G43gat;
	input G50gat;
	input G57gat;
	input G64gat;
	input G71gat;
	input G78gat;
	input G85gat;
	input G92gat;
	input G99gat;
	input G106gat;
	input G113gat;
	input G120gat;
	input G127gat;
	input G134gat;
	input G141gat;
	input G148gat;
	input G155gat;
	input G162gat;
	input G169gat;
	input G176gat;
	input G183gat;
	input G190gat;
	input G197gat;
	input G204gat;
	input G211gat;
	input G218gat;
	input G225gat;
	input G226gat;
	input G227gat;
	input G228gat;
	input G229gat;
	input G230gat;
	input G231gat;
	input G232gat;
	input G233gat;
	output G1324gat;
	output G1325gat;
	output G1326gat;
	output G1327gat;
	output G1328gat;
	output G1329gat;
	output G1330gat;
	output G1331gat;
	output G1332gat;
	output G1333gat;
	output G1334gat;
	output G1335gat;
	output G1336gat;
	output G1337gat;
	output G1338gat;
	output G1339gat;
	output G1340gat;
	output G1341gat;
	output G1342gat;
	output G1343gat;
	output G1344gat;
	output G1345gat;
	output G1346gat;
	output G1347gat;
	output G1348gat;
	output G1349gat;
	output G1350gat;
	output G1351gat;
	output G1352gat;
	output G1353gat;
	output G1354gat;
	output G1355gat;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n178;
	wire n179;
	wire n181;
	wire n182;
	wire n184;
	wire n185;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n193;
	wire n195;
	wire n197;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n205;
	wire n207;
	wire n209;
	wire n211;
	wire n212;
	wire n214;
	wire n216;
	wire n218;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n233;
	wire n235;
	wire n237;
	wire n239;
	wire n240;
	wire n241;
	wire n243;
	wire n245;
	wire n247;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n254;
	wire n256;
	wire n258;
	wire n260;
	wire n261;
	wire n263;
	wire n265;
	wire n267;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G15gat_0;
	wire [2:0] w_G22gat_0;
	wire [2:0] w_G29gat_0;
	wire [2:0] w_G36gat_0;
	wire [2:0] w_G43gat_0;
	wire [2:0] w_G50gat_0;
	wire [2:0] w_G57gat_0;
	wire [2:0] w_G64gat_0;
	wire [2:0] w_G71gat_0;
	wire [2:0] w_G78gat_0;
	wire [2:0] w_G85gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G113gat_0;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G127gat_0;
	wire [2:0] w_G134gat_0;
	wire [2:0] w_G141gat_0;
	wire [2:0] w_G148gat_0;
	wire [2:0] w_G155gat_0;
	wire [2:0] w_G162gat_0;
	wire [2:0] w_G169gat_0;
	wire [2:0] w_G176gat_0;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G190gat_0;
	wire [2:0] w_G197gat_0;
	wire [2:0] w_G204gat_0;
	wire [2:0] w_G211gat_0;
	wire [2:0] w_G218gat_0;
	wire [2:0] w_G233gat_0;
	wire [2:0] w_G233gat_1;
	wire [1:0] w_n78_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n86_0;
	wire [1:0] w_n86_1;
	wire [2:0] w_n87_0;
	wire [2:0] w_n87_1;
	wire [1:0] w_n93_0;
	wire [2:0] w_n96_0;
	wire [1:0] w_n96_1;
	wire [1:0] w_n100_0;
	wire [2:0] w_n102_0;
	wire [1:0] w_n102_1;
	wire [1:0] w_n108_0;
	wire [1:0] w_n114_0;
	wire [2:0] w_n116_0;
	wire [1:0] w_n116_1;
	wire [2:0] w_n117_0;
	wire [2:0] w_n117_1;
	wire [1:0] w_n118_0;
	wire [1:0] w_n124_0;
	wire [1:0] w_n130_0;
	wire [2:0] w_n132_0;
	wire [1:0] w_n132_1;
	wire [2:0] w_n141_0;
	wire [1:0] w_n141_1;
	wire [2:0] w_n149_0;
	wire [1:0] w_n149_1;
	wire [2:0] w_n155_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [2:0] w_n164_0;
	wire [2:0] w_n164_1;
	wire [2:0] w_n172_0;
	wire [1:0] w_n172_1;
	wire [1:0] w_n173_0;
	wire [2:0] w_n175_0;
	wire [1:0] w_n175_1;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n184_0;
	wire [2:0] w_n184_1;
	wire [2:0] w_n187_0;
	wire [2:0] w_n187_1;
	wire [1:0] w_n189_0;
	wire [2:0] w_n190_0;
	wire [1:0] w_n190_1;
	wire [2:0] w_n199_0;
	wire [2:0] w_n199_1;
	wire [1:0] w_n200_0;
	wire [2:0] w_n202_0;
	wire [1:0] w_n202_1;
	wire [2:0] w_n211_0;
	wire [1:0] w_n211_1;
	wire [1:0] w_n220_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n229_0;
	wire [2:0] w_n230_0;
	wire [1:0] w_n230_1;
	wire [1:0] w_n239_0;
	wire [2:0] w_n240_0;
	wire [1:0] w_n240_1;
	wire [1:0] w_n250_0;
	wire [2:0] w_n251_0;
	wire [1:0] w_n251_1;
	wire [2:0] w_n260_0;
	wire [1:0] w_n260_1;
	wire w_dff_A_8JuFjjCQ2_0;
	wire w_dff_B_8NUdgw8m9_2;
	wire w_dff_B_am6g3HwZ6_2;
	wire w_dff_A_AS5DiFPi6_1;
	wire w_dff_B_icqtxdVr5_2;
	wire w_dff_B_zvAI8Bn44_2;
	wire w_dff_B_HX8pgkMt4_2;
	wire w_dff_B_Ao3mF6jD5_2;
	wire w_dff_B_xvKMKOjR6_2;
	wire w_dff_B_5mJw1h9l2_0;
	wire w_dff_B_HukrD1ZN6_0;
	wire w_dff_B_L8hwV9M20_1;
	wire w_dff_A_CuTx14e61_0;
	wire w_dff_A_Sdvdv2ww4_0;
	wire w_dff_A_q9i9M5zw9_0;
	wire w_dff_A_bBfmBw576_0;
	wire w_dff_A_CYjvTZXb0_0;
	wire w_dff_A_qrJVjDxM4_0;
	wire w_dff_A_FyMtaAU47_0;
	wire w_dff_A_fT9dh2oP6_1;
	wire w_dff_A_a7y40y1C5_1;
	wire w_dff_A_mYLiq6mY2_1;
	wire w_dff_A_6X2jNa6m2_1;
	wire w_dff_A_vgv1IbVN6_1;
	wire w_dff_A_L20QRunt7_0;
	wire w_dff_A_zaRGelBp6_0;
	wire w_dff_A_9Y8Y2EZM4_0;
	wire w_dff_A_pHHr8qCy1_0;
	wire w_dff_A_SWUusfbe4_0;
	wire w_dff_A_O57MIXbh7_1;
	wire w_dff_A_bz85RdKA4_1;
	wire w_dff_A_STu1RUb93_1;
	wire w_dff_A_LXuHtb6K8_1;
	wire w_dff_A_9dMBYRhg5_1;
	wire w_dff_A_sEZ1BWzB8_0;
	wire w_dff_A_Fh30niyP0_0;
	wire w_dff_A_2lnlPTc33_0;
	wire w_dff_A_NTJGSX5p8_0;
	wire w_dff_A_fozk3laX3_0;
	wire w_dff_A_GTG0p0QH6_1;
	wire w_dff_A_KWRa1ulO8_1;
	wire w_dff_A_vy53priu5_1;
	wire w_dff_A_A6Z2XqIo9_1;
	wire w_dff_A_Xb55nq249_1;
	wire w_dff_B_yIG8Xxhd6_1;
	wire w_dff_B_e4ssjTZ55_1;
	wire w_dff_A_9TBx4ji69_0;
	wire w_dff_A_noTTOzMr3_0;
	wire w_dff_A_oX3TABZB0_0;
	wire w_dff_A_Wn2kC3ox6_0;
	wire w_dff_A_9LSOWbPS8_0;
	wire w_dff_A_VhTbhjy14_2;
	wire w_dff_A_EeJvPDNh1_2;
	wire w_dff_A_Q9hIvtog2_2;
	wire w_dff_A_CrbgB4IN2_2;
	wire w_dff_A_bfNkBzqG1_2;
	wire w_dff_A_WIcU59q00_0;
	wire w_dff_A_vNqZzioz3_0;
	wire w_dff_A_3fjB3M6l9_0;
	wire w_dff_A_YvSJDBRq8_0;
	wire w_dff_A_1EwuVeVU7_0;
	wire w_dff_A_Y5gXd9006_1;
	wire w_dff_A_XRZTSRNe1_1;
	wire w_dff_A_0HTn2Dt71_1;
	wire w_dff_A_72m1i4TZ8_1;
	wire w_dff_A_QQ4lHGA13_1;
	wire w_dff_B_nemRtXzG4_2;
	wire w_dff_B_cNMapHAP6_2;
	wire w_dff_B_YnP07Vuw0_2;
	wire w_dff_A_5OuMraU69_0;
	wire w_dff_A_TLbyTtBw5_0;
	wire w_dff_A_4klv3bXp6_0;
	wire w_dff_A_9FEDRJlK1_0;
	wire w_dff_A_eb0E6ue46_0;
	wire w_dff_A_0Joc3Vii4_2;
	wire w_dff_A_qng5xjpf1_2;
	wire w_dff_A_K1OUCfD43_2;
	wire w_dff_A_9HRfUdej9_2;
	wire w_dff_A_JsXhfJE76_2;
	wire w_dff_A_EWZzrm5V2_1;
	wire w_dff_A_w8oUgXdQ0_1;
	wire w_dff_A_lJoPA1BP5_1;
	wire w_dff_A_JG5HPrIz9_1;
	wire w_dff_A_I29TAoUH3_1;
	wire w_dff_A_qM65IoOa8_2;
	wire w_dff_A_ZI4Jn9Nr1_2;
	wire w_dff_A_KBequAQw6_2;
	wire w_dff_A_wOdA5qfh8_2;
	wire w_dff_A_aKl7Y1CB7_2;
	wire w_dff_A_nApm0Jzs2_0;
	wire w_dff_A_nDFyIYZ49_1;
	wire w_dff_A_esT7zxR70_1;
	wire w_dff_A_k2S79Kwl5_1;
	wire w_dff_A_ED9ixB6q2_1;
	wire w_dff_A_RKWXYvMO3_1;
	wire w_dff_A_YtOrFiTv2_2;
	wire w_dff_A_hZgvwz5H1_2;
	wire w_dff_A_olcDohVr6_2;
	wire w_dff_A_0pmU4C2a3_2;
	wire w_dff_A_nCJDKVfu2_2;
	wire w_dff_A_1KuXAB0J0_1;
	wire w_dff_A_xTJyjQSd0_1;
	wire w_dff_A_sFsaMdu40_1;
	wire w_dff_A_8fbEma5R7_1;
	wire w_dff_A_0owp1E3X3_1;
	wire w_dff_A_3Rfm1gUM6_1;
	wire w_dff_A_dNaCs9U53_2;
	wire w_dff_A_DJ03KHzt2_2;
	wire w_dff_A_7KyCDYpz0_2;
	wire w_dff_A_ggwqiEHo5_2;
	wire w_dff_A_TTNNcIoX3_2;
	wire w_dff_A_lQZyNmHG3_0;
	wire w_dff_B_cpb3gZPs5_1;
	wire w_dff_B_C9BeA8KM7_1;
	wire w_dff_B_xzTrjmVV4_0;
	wire w_dff_A_BgzgqeGf9_2;
	wire w_dff_A_oF1y5N940_2;
	wire w_dff_A_EyhmX1MY6_2;
	wire w_dff_A_28Nizbl97_0;
	wire w_dff_A_q8tswYZT7_0;
	wire w_dff_A_1BnerfKd7_0;
	wire w_dff_A_8VSuDl4t1_0;
	wire w_dff_A_oS4wZYHo2_0;
	wire w_dff_A_Gc94o9pn1_2;
	wire w_dff_A_rUMWj6Xa2_2;
	wire w_dff_A_ta2rhT3d4_2;
	wire w_dff_A_1EWKPCFS3_2;
	wire w_dff_A_ZWHn74Gi5_2;
	wire w_dff_A_bMqIfJaP7_1;
	wire w_dff_A_Gy2CJJnj2_0;
	wire w_dff_A_Waq2GnRU5_0;
	wire w_dff_A_rIbPlINT4_0;
	wire w_dff_A_mYQpjEIT1_0;
	wire w_dff_A_MUecw0188_0;
	wire w_dff_A_rp1YaFq33_0;
	wire w_dff_A_9ql2u9ZS2_0;
	wire w_dff_A_VEU5HbcK8_0;
	wire w_dff_A_2OfhNg3O0_0;
	wire w_dff_A_GuJuuoNy3_0;
	wire w_dff_A_mMj5LMFW2_0;
	wire w_dff_A_RTpFpdC09_0;
	wire w_dff_A_6vFxHHfd4_0;
	wire w_dff_A_oZG3wzxO0_0;
	wire w_dff_A_Ag32BBoU1_0;
	wire w_dff_A_VQr5k33k2_0;
	wire w_dff_A_iu6nTUdv9_0;
	wire w_dff_A_MxUjFTQs7_0;
	wire w_dff_A_9clkR7LB8_0;
	wire w_dff_A_Y4yvmXJ00_0;
	wire w_dff_A_kUkOPeyL7_0;
	wire w_dff_A_zxy5Nh8h9_0;
	wire w_dff_A_JeFRJKoD5_1;
	wire w_dff_A_YsSOuQPd4_2;
	wire w_dff_A_fjyD841N9_0;
	wire w_dff_A_avJj2ftp0_0;
	wire w_dff_A_tuYWeo190_0;
	wire w_dff_A_bYbJAC8d0_0;
	wire w_dff_A_UhrEUqlX9_0;
	wire w_dff_A_ipxFgEKq0_0;
	wire w_dff_A_bayfh9BD1_0;
	wire w_dff_A_kXsHjL2F7_0;
	wire w_dff_A_gZJUWUz46_0;
	wire w_dff_A_C7ey6viR4_0;
	wire w_dff_A_q3IXA9W52_0;
	wire w_dff_A_c8M1Daca4_0;
	wire w_dff_A_DeYvB5iv4_0;
	wire w_dff_A_8x6vm9N22_0;
	wire w_dff_A_a8nYAgs06_0;
	wire w_dff_A_RVttjQKE7_0;
	wire w_dff_A_9mHACmty0_0;
	wire w_dff_A_lrmPbqPV3_0;
	wire w_dff_A_9Zndlanj0_0;
	wire w_dff_A_ojE9KtrR0_0;
	wire w_dff_A_HIeUN9hn4_0;
	wire w_dff_A_9XxXW3xX6_0;
	wire w_dff_B_FN6x3i5p4_2;
	wire w_dff_B_DZK3WZP06_2;
	wire w_dff_B_mgU9srBl5_2;
	wire w_dff_A_5rpBHZ9Y5_0;
	wire w_dff_A_wS3rMX7Z2_0;
	wire w_dff_A_obZl66Kp2_0;
	wire w_dff_A_b3ZU5CRD9_0;
	wire w_dff_A_A5YsYjkw6_0;
	wire w_dff_A_6ksQyobo0_2;
	wire w_dff_A_FW6K1mqG8_2;
	wire w_dff_A_fFLvYv756_2;
	wire w_dff_A_hNg3QhNa1_2;
	wire w_dff_A_GTn9ZlPg9_2;
	wire w_dff_A_mOfIDB2G0_1;
	wire w_dff_A_IBrKcLNG2_0;
	wire w_dff_A_9kJParzG4_0;
	wire w_dff_A_v5B8dYbp6_0;
	wire w_dff_A_3JJvdBJw4_0;
	wire w_dff_A_mGkbc5EB5_0;
	wire w_dff_A_cS1pVD993_0;
	wire w_dff_A_a1uA0RCw3_0;
	wire w_dff_A_hoHB0SEm3_0;
	wire w_dff_A_CscjWyJh9_0;
	wire w_dff_A_298x2fhx8_0;
	wire w_dff_A_QUevK6dp3_0;
	wire w_dff_A_GrMeMyZF1_0;
	wire w_dff_A_3uUohaPd7_0;
	wire w_dff_A_vPVttXBf1_0;
	wire w_dff_A_ZenmOmLK7_0;
	wire w_dff_A_VCQ27pGC2_0;
	wire w_dff_A_WcmBgBec0_0;
	wire w_dff_A_rxSUfTEa1_0;
	wire w_dff_A_jrftIraZ8_0;
	wire w_dff_A_5zQR7pOJ1_0;
	wire w_dff_A_IyqTxqZr5_0;
	wire w_dff_A_jysE7TwX7_0;
	wire w_dff_A_Wjup1IRw4_0;
	wire w_dff_A_LXkA0udj3_0;
	wire w_dff_A_sNOjqHPW9_0;
	wire w_dff_A_HH4SlpT82_0;
	wire w_dff_A_2TxDSsYj0_0;
	wire w_dff_A_AoQqhtKp4_0;
	wire w_dff_A_hvEi9KZs8_0;
	wire w_dff_A_Ws3QqX2U4_0;
	wire w_dff_A_CSyVbtZr0_0;
	wire w_dff_A_60vNMrCt1_0;
	wire w_dff_A_ngdY3SaI8_0;
	wire w_dff_A_dUlmOZCS9_0;
	wire w_dff_A_t88rpmNf5_0;
	wire w_dff_A_05NRixIk1_0;
	wire w_dff_A_qFwhbF090_0;
	wire w_dff_A_62pxMxPT3_0;
	wire w_dff_A_gIvEyhlY3_0;
	wire w_dff_A_IrNsnhhT7_0;
	wire w_dff_A_BsFFiPo78_0;
	wire w_dff_A_VtflH0ef6_0;
	wire w_dff_A_kLAoUdji0_0;
	wire w_dff_A_9QQ3fZkz9_0;
	wire w_dff_A_F1ag4jyI7_0;
	wire w_dff_A_7Ad9wT1O1_0;
	wire w_dff_A_6zZSLCky6_0;
	wire w_dff_A_WS9y7ycB1_0;
	wire w_dff_A_dTzzst487_0;
	wire w_dff_A_w5eDU67r2_0;
	wire w_dff_A_7gg6dw5F5_0;
	wire w_dff_A_TTbcbWoG6_0;
	wire w_dff_A_6dhh8FJW0_0;
	wire w_dff_A_v4rVVFR89_0;
	wire w_dff_A_BwzKoTGC1_0;
	wire w_dff_A_ltmQRJef6_0;
	wire w_dff_A_2wmY0NjK8_0;
	wire w_dff_A_jWcYPu8D1_0;
	wire w_dff_A_WbFxjA5x8_0;
	wire w_dff_A_aOxQvsnk3_0;
	wire w_dff_A_VnaQW3wC7_0;
	wire w_dff_A_msJfL2z22_0;
	wire w_dff_A_syAWKpDS8_0;
	wire w_dff_A_F9ivLoom3_0;
	wire w_dff_A_AYXiWdPm5_0;
	wire w_dff_A_KrOmtTGV2_0;
	wire w_dff_A_b39vc3QZ9_0;
	wire w_dff_A_J9bzhHzr3_0;
	wire w_dff_A_mBQ4E0OV7_0;
	wire w_dff_A_BhhvN9zP2_0;
	wire w_dff_A_zNvTAT2H4_0;
	wire w_dff_A_XYOFRBsW9_0;
	wire w_dff_A_u0Vo8dHc9_0;
	wire w_dff_A_8sJHAHMa8_0;
	wire w_dff_A_YvDo8HyO0_0;
	wire w_dff_A_fOyPEcy97_0;
	wire w_dff_A_Gwy7oFm21_0;
	wire w_dff_A_9hFN8fiq0_0;
	wire w_dff_A_29a9GGBp5_0;
	wire w_dff_A_sLB8Djhu8_0;
	wire w_dff_A_b0BNUmcL6_0;
	wire w_dff_A_ZBxHxwk98_0;
	wire w_dff_A_SOqBOHeV2_0;
	wire w_dff_A_9peYCn8v9_0;
	wire w_dff_A_eUmG3bzi4_0;
	wire w_dff_A_nDGzSmq67_0;
	wire w_dff_A_Z2bMR47X9_0;
	wire w_dff_A_lMiBnJV77_0;
	wire w_dff_A_ijYXtsu43_1;
	wire w_dff_A_Lb6kz2pA7_0;
	wire w_dff_A_sbVzrm911_0;
	wire w_dff_A_NEf6hx670_0;
	wire w_dff_A_zN7s2WAX1_0;
	wire w_dff_A_EcDuipzG7_0;
	wire w_dff_A_BIttUVuv5_0;
	wire w_dff_A_HE2q2hQk9_0;
	wire w_dff_A_l4ZNmGCZ2_0;
	wire w_dff_A_pBytW4Ve6_0;
	wire w_dff_A_EIa4wKO89_0;
	wire w_dff_A_ZuYfv5UA5_0;
	wire w_dff_A_isSYifqF7_0;
	wire w_dff_A_RUmCfxN44_0;
	wire w_dff_A_wWNqEg6X7_0;
	wire w_dff_A_Pp61Fpnw7_0;
	wire w_dff_A_pTWFA8Of1_0;
	wire w_dff_A_FzCodUre2_0;
	wire w_dff_A_ooi2NbM65_0;
	wire w_dff_A_CjkmQe6O8_0;
	wire w_dff_A_pNXEIKWR9_0;
	wire w_dff_A_aR24SEHt8_0;
	wire w_dff_A_uiifWNTX9_0;
	wire w_dff_A_IlsdWfLE1_0;
	wire w_dff_A_WLrUWIod0_0;
	wire w_dff_A_F99SQd835_0;
	wire w_dff_A_b3MpnxRj6_0;
	wire w_dff_A_AzpbqCB43_0;
	wire w_dff_A_9XpmKFk98_0;
	wire w_dff_A_FASDJSlH3_0;
	wire w_dff_A_jgB2nQ7x2_0;
	wire w_dff_A_4Wki2hco9_0;
	wire w_dff_A_ZXMVv5bR9_0;
	wire w_dff_A_k98m0A6N9_0;
	wire w_dff_A_ZNghoZoP8_0;
	wire w_dff_A_bDis0Ej32_0;
	wire w_dff_A_nfbbIKTc1_0;
	wire w_dff_A_hC9ErcYS1_0;
	wire w_dff_A_hcP8IOIL7_0;
	wire w_dff_A_N4nYGrpn9_0;
	wire w_dff_A_iWCToGTf4_0;
	wire w_dff_A_OKp1P4BM3_0;
	wire w_dff_A_44dvDDGH3_0;
	wire w_dff_A_1A3pKgdw0_0;
	wire w_dff_A_9Zmys9zm8_0;
	wire w_dff_A_F5f0KTTL2_0;
	wire w_dff_A_1zeN642C6_0;
	wire w_dff_A_tVwf1G7g4_0;
	wire w_dff_A_amEVcshH5_0;
	wire w_dff_A_6q4EgFg07_0;
	wire w_dff_A_P024Q8QK2_0;
	wire w_dff_A_jWQzdFGG2_0;
	wire w_dff_A_iIdzb1Zl8_0;
	wire w_dff_A_GBzglkQJ2_0;
	wire w_dff_A_bFixfnyz9_0;
	wire w_dff_A_wNbvbPej9_0;
	wire w_dff_A_FkeL3ixr3_0;
	wire w_dff_A_md2Y4LjD5_0;
	wire w_dff_A_YRE9P2K52_0;
	wire w_dff_A_dLDKf2tP4_0;
	wire w_dff_A_btBz3Pw79_0;
	wire w_dff_A_L7Opz9Ul2_0;
	wire w_dff_A_rQeAf3kD2_0;
	wire w_dff_A_D6sWsJ3m5_0;
	wire w_dff_A_OpM7NSH44_0;
	wire w_dff_A_b7D4FyFS5_0;
	wire w_dff_A_DXT6JGjF6_0;
	wire w_dff_A_TZkhoD105_0;
	wire w_dff_A_nnUOQRxn3_0;
	wire w_dff_A_uEx2BNFk1_0;
	wire w_dff_A_ojGlo7Fo9_0;
	wire w_dff_A_fMUtyY8P0_0;
	wire w_dff_A_DF38NtLE4_0;
	wire w_dff_A_Fycx3Eoy4_0;
	wire w_dff_A_cMorxdi31_0;
	wire w_dff_A_HMzP6F4k3_0;
	wire w_dff_A_eCzi1cYe3_0;
	wire w_dff_A_FKRrwreq2_0;
	wire w_dff_A_XLv82hXB4_0;
	wire w_dff_A_tfMOTZAD1_0;
	wire w_dff_A_L4eZFemM2_0;
	wire w_dff_A_mzaJ5xL68_0;
	wire w_dff_A_rLx6zcib2_0;
	wire w_dff_A_bS4eyqfj1_0;
	wire w_dff_A_6htZAKQQ3_0;
	wire w_dff_A_jzfnpbd26_0;
	wire w_dff_A_rLBsRemY7_0;
	wire w_dff_A_adApjwo32_0;
	wire w_dff_A_l7QUQJ4y2_0;
	wire w_dff_A_wu2Fi6xf5_1;
	wire w_dff_A_QHtTSUqp2_1;
	wire w_dff_A_UhfF8zm33_1;
	wire w_dff_A_vlAdmt1s4_1;
	wire w_dff_A_4G4z2rLk7_1;
	wire w_dff_A_3fJI5Gln5_2;
	wire w_dff_A_P3ilw5YH3_2;
	wire w_dff_A_JpauP8u43_2;
	wire w_dff_A_MO0shkh64_2;
	wire w_dff_A_TWxn2FOh5_2;
	wire w_dff_A_ObRYbEa95_1;
	wire w_dff_A_eeBMqcSL9_0;
	wire w_dff_A_81y54dIb4_0;
	wire w_dff_A_99p2sCA35_0;
	wire w_dff_A_vuXmwXtk2_0;
	wire w_dff_A_zU1yKGA75_0;
	wire w_dff_A_nN6CIYEv6_0;
	wire w_dff_A_zupqc8xA8_0;
	wire w_dff_A_R6QXTkRz7_0;
	wire w_dff_A_AcC6QKlA7_0;
	wire w_dff_A_Aw6xG1tM9_0;
	wire w_dff_A_M9pBSjVC9_0;
	wire w_dff_A_NEQrfpyP2_0;
	wire w_dff_A_dNzug4h47_0;
	wire w_dff_A_JbObE0ED8_0;
	wire w_dff_A_4ePAcUgm1_0;
	wire w_dff_A_Z2FUtYC02_0;
	wire w_dff_A_k1syVgTO2_0;
	wire w_dff_A_gxRxyFBv0_0;
	wire w_dff_A_XtD5lwcV3_0;
	wire w_dff_A_UBMdbGhA9_0;
	wire w_dff_A_zPTZq0wv6_0;
	wire w_dff_A_i5GnN5Yd6_0;
	wire w_dff_A_ZHwhbieb2_0;
	wire w_dff_A_mBUG7djK3_0;
	wire w_dff_A_a8TreNbt2_0;
	wire w_dff_A_cNds3O5H4_0;
	wire w_dff_A_WSi4d5NM0_0;
	wire w_dff_A_FMY34EcV9_0;
	wire w_dff_A_UOYNfn8m1_0;
	wire w_dff_A_da63xLHh9_0;
	wire w_dff_A_IMc9dQrW2_0;
	wire w_dff_A_5WiMBiUZ1_0;
	wire w_dff_A_horf3TtB3_0;
	wire w_dff_A_O07U9qP48_0;
	wire w_dff_A_dDPdfrUH9_0;
	wire w_dff_A_SxLffwx60_0;
	wire w_dff_A_7AGBAL0J9_0;
	wire w_dff_A_gZc4VdEM7_0;
	wire w_dff_A_28NRwmeY6_0;
	wire w_dff_A_9kuC86Nm8_0;
	wire w_dff_A_ER1xiWRB0_0;
	wire w_dff_A_j0gRPcQX1_0;
	wire w_dff_A_OomMhRsY9_0;
	wire w_dff_A_iqz6IBc73_0;
	wire w_dff_A_fKZ0sX0M6_0;
	wire w_dff_A_l9dYyST45_0;
	wire w_dff_A_zjdxJQMp2_0;
	wire w_dff_A_1PUk7Ety7_0;
	wire w_dff_A_LgyQ6g5M7_0;
	wire w_dff_A_vEnIl3od7_0;
	wire w_dff_A_M6rDpDZN8_0;
	wire w_dff_A_vFOH2N399_0;
	wire w_dff_A_mbP7sAWu4_0;
	wire w_dff_A_6l3GUOco6_0;
	wire w_dff_A_J8e7MW7e3_0;
	wire w_dff_A_9TFueqTW3_0;
	wire w_dff_A_UTDp6bgi1_0;
	wire w_dff_A_WI44idSQ7_0;
	wire w_dff_A_duHRM7dn9_0;
	wire w_dff_A_wdC1AY5R5_0;
	wire w_dff_A_ThnwJJzD5_0;
	wire w_dff_A_Lih1vTLs0_0;
	wire w_dff_A_t73Q1kH36_0;
	wire w_dff_A_G7YnaCet8_0;
	wire w_dff_A_539bRIsv3_0;
	wire w_dff_A_ogvUz4vm1_0;
	wire w_dff_A_WGUmRrbA4_0;
	wire w_dff_A_4XW7jGFD4_0;
	wire w_dff_A_V1JfakCo9_0;
	wire w_dff_A_pLFom1cO5_0;
	wire w_dff_A_a7OoHm4U7_0;
	wire w_dff_A_v4vRyEaP1_0;
	wire w_dff_A_EL1XSLtn3_0;
	wire w_dff_A_pvUwuCBL8_0;
	wire w_dff_A_FKu71oGJ6_0;
	wire w_dff_A_abmM5fXE4_0;
	wire w_dff_A_zEYHoXXM2_0;
	wire w_dff_A_jxH1okq01_0;
	wire w_dff_A_KACfGxsG0_0;
	wire w_dff_A_MKCBvkUz4_0;
	wire w_dff_A_MzSnlUK85_0;
	wire w_dff_A_XvIpWAEw2_0;
	wire w_dff_A_KyC6agDj9_0;
	wire w_dff_A_bekBbxnn6_0;
	wire w_dff_A_4aA0BhyM5_0;
	wire w_dff_A_G4XyztvT0_0;
	wire w_dff_A_Mw7a1sut3_0;
	wire w_dff_A_p1F05AkQ9_0;
	wire w_dff_A_60qy12T34_0;
	wire w_dff_A_RgSEkwA58_0;
	wire w_dff_A_PoS3Xb0E1_0;
	wire w_dff_A_oLIAvyFR7_0;
	wire w_dff_A_QW4mBDm74_0;
	wire w_dff_A_y4Sd6yUH4_0;
	wire w_dff_A_3CTHyfGu1_0;
	wire w_dff_A_eXDMBhMJ3_0;
	wire w_dff_A_jgWMoFNs0_0;
	wire w_dff_A_p16PEy079_0;
	wire w_dff_A_XAMCx2EQ4_0;
	wire w_dff_A_drjs0qgZ6_0;
	wire w_dff_A_w4W9N0gC2_0;
	wire w_dff_A_s5uTdpFC1_0;
	wire w_dff_A_zn0AjZ8j1_0;
	wire w_dff_A_HjSzdfsR2_0;
	wire w_dff_A_8EvGxAog9_0;
	wire w_dff_A_ndqVGKcx9_0;
	wire w_dff_A_TN4iO5KY6_0;
	wire w_dff_A_THdEW0hn9_0;
	wire w_dff_A_UF18l7zG8_0;
	wire w_dff_A_veYjb4335_0;
	wire w_dff_A_k9ckY6gO7_0;
	wire w_dff_A_HSPjeVkt8_0;
	wire w_dff_A_676eCCUB0_0;
	wire w_dff_A_lh4CpKCC9_0;
	wire w_dff_A_kbc9h4uc7_0;
	wire w_dff_A_3Mkj6noc0_0;
	wire w_dff_A_1Tym3ah83_0;
	wire w_dff_A_Fk7Z8YEN9_0;
	wire w_dff_A_62MbArOl0_0;
	wire w_dff_A_MiIvMP0N9_0;
	wire w_dff_A_odWp6WvU9_0;
	wire w_dff_A_SU5SE6Es6_0;
	wire w_dff_A_UvXJo7II8_0;
	wire w_dff_A_SVfkbTlp9_0;
	wire w_dff_A_yByDrXlw0_0;
	wire w_dff_A_lNUBuyqd2_0;
	wire w_dff_A_Sqv5eqQ09_0;
	wire w_dff_A_XVXoWrNB6_0;
	wire w_dff_A_YDslV3Dm6_0;
	wire w_dff_A_u5d3WRZt3_0;
	wire w_dff_A_Tt4PlzHN7_0;
	wire w_dff_A_9BZA5ENF8_0;
	jxor g000(.dina(w_G85gat_0[2]),.dinb(w_G57gat_0[2]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_G29gat_0[2]),.dinb(w_G1gat_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(n74),.dinb(n73),.dout(n75),.clk(gclk));
	jxor g003(.dina(w_G162gat_0[2]),.dinb(w_G155gat_0[2]),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_G148gat_0[2]),.dinb(w_G141gat_0[2]),.dout(n77),.clk(gclk));
	jxor g005(.dina(n77),.dinb(n76),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_n78_0[1]),.dinb(n75),.dout(n79),.clk(gclk));
	jand g007(.dina(w_G233gat_1[2]),.dinb(G225gat),.dout(n80),.clk(gclk));
	jnot g008(.din(n80),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_G134gat_0[2]),.dinb(w_G127gat_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(w_G120gat_0[2]),.dinb(w_G113gat_0[2]),.dout(n83),.clk(gclk));
	jxor g011(.dina(n83),.dinb(n82),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n81),.dout(n85),.clk(gclk));
	jxor g013(.dina(n85),.dinb(n79),.dout(n86),.clk(gclk));
	jnot g014(.din(w_n86_1[1]),.dout(n87),.clk(gclk));
	jxor g015(.dina(w_G218gat_0[2]),.dinb(w_G190gat_0[2]),.dout(n88),.clk(gclk));
	jxor g016(.dina(w_G162gat_0[1]),.dinb(w_G134gat_0[1]),.dout(n89),.clk(gclk));
	jxor g017(.dina(n89),.dinb(n88),.dout(n90),.clk(gclk));
	jxor g018(.dina(w_G106gat_0[2]),.dinb(w_G99gat_0[2]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_G92gat_0[2]),.dinb(w_G85gat_0[1]),.dout(n92),.clk(gclk));
	jxor g020(.dina(n92),.dinb(n91),.dout(n93),.clk(gclk));
	jxor g021(.dina(w_n93_0[1]),.dinb(n90),.dout(n94),.clk(gclk));
	jnot g022(.din(G232gat),.dout(n95),.clk(gclk));
	jnot g023(.din(w_G233gat_1[1]),.dout(n96),.clk(gclk));
	jor g024(.dina(w_n96_1[1]),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_G50gat_0[2]),.dinb(w_G43gat_0[2]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_G36gat_0[2]),.dinb(w_G29gat_0[1]),.dout(n99),.clk(gclk));
	jxor g027(.dina(n99),.dinb(n98),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_n100_0[1]),.dinb(n97),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n94),.dout(n102),.clk(gclk));
	jxor g030(.dina(w_G211gat_0[2]),.dinb(w_G183gat_0[2]),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_G155gat_0[1]),.dinb(w_G127gat_0[1]),.dout(n104),.clk(gclk));
	jxor g032(.dina(n104),.dinb(n103),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_G78gat_0[2]),.dinb(w_G71gat_0[2]),.dout(n106),.clk(gclk));
	jxor g034(.dina(w_G64gat_0[2]),.dinb(w_G57gat_0[1]),.dout(n107),.clk(gclk));
	jxor g035(.dina(n107),.dinb(n106),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_n108_0[1]),.dinb(n105),.dout(n109),.clk(gclk));
	jnot g037(.din(G231gat),.dout(n110),.clk(gclk));
	jor g038(.dina(w_n96_1[0]),.dinb(n110),.dout(n111),.clk(gclk));
	jxor g039(.dina(w_G22gat_0[2]),.dinb(w_G15gat_0[2]),.dout(n112),.clk(gclk));
	jxor g040(.dina(w_G8gat_0[2]),.dinb(w_G1gat_0[1]),.dout(n113),.clk(gclk));
	jxor g041(.dina(n113),.dinb(n112),.dout(n114),.clk(gclk));
	jxor g042(.dina(w_n114_0[1]),.dinb(n111),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n109),.dout(n116),.clk(gclk));
	jnot g044(.din(w_n116_1[1]),.dout(n117),.clk(gclk));
	jand g045(.dina(w_n117_1[2]),.dinb(w_n102_1[1]),.dout(n118),.clk(gclk));
	jxor g046(.dina(w_G92gat_0[1]),.dinb(w_G64gat_0[1]),.dout(n119),.clk(gclk));
	jxor g047(.dina(w_G36gat_0[1]),.dinb(w_G8gat_0[1]),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(n119),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_G190gat_0[1]),.dinb(w_G183gat_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_G176gat_0[2]),.dinb(w_G169gat_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(w_n124_0[1]),.dinb(n121),.dout(n125),.clk(gclk));
	jand g053(.dina(w_G233gat_1[0]),.dinb(G226gat),.dout(n126),.clk(gclk));
	jnot g054(.din(n126),.dout(n127),.clk(gclk));
	jxor g055(.dina(w_G218gat_0[1]),.dinb(w_G211gat_0[1]),.dout(n128),.clk(gclk));
	jxor g056(.dina(w_G204gat_0[2]),.dinb(w_G197gat_0[2]),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(n128),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_n130_0[1]),.dinb(n127),.dout(n131),.clk(gclk));
	jxor g059(.dina(n131),.dinb(n125),.dout(n132),.clk(gclk));
	jxor g060(.dina(w_n132_1[1]),.dinb(w_n86_1[0]),.dout(n133),.clk(gclk));
	jxor g061(.dina(w_G99gat_0[1]),.dinb(w_G71gat_0[1]),.dout(n134),.clk(gclk));
	jxor g062(.dina(w_G43gat_0[1]),.dinb(w_G15gat_0[1]),.dout(n135),.clk(gclk));
	jxor g063(.dina(n135),.dinb(n134),.dout(n136),.clk(gclk));
	jxor g064(.dina(n136),.dinb(w_n124_0[0]),.dout(n137),.clk(gclk));
	jnot g065(.din(G227gat),.dout(n138),.clk(gclk));
	jor g066(.dina(w_n96_0[2]),.dinb(n138),.dout(n139),.clk(gclk));
	jxor g067(.dina(n139),.dinb(w_n84_0[0]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n137),.dout(n141),.clk(gclk));
	jxor g069(.dina(w_G106gat_0[1]),.dinb(w_G78gat_0[1]),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_G50gat_0[1]),.dinb(w_G22gat_0[1]),.dout(n143),.clk(gclk));
	jxor g071(.dina(n143),.dinb(n142),.dout(n144),.clk(gclk));
	jxor g072(.dina(n144),.dinb(w_n130_0[0]),.dout(n145),.clk(gclk));
	jnot g073(.din(G228gat),.dout(n146),.clk(gclk));
	jor g074(.dina(w_n96_0[1]),.dinb(n146),.dout(n147),.clk(gclk));
	jxor g075(.dina(n147),.dinb(w_n78_0[0]),.dout(n148),.clk(gclk));
	jxor g076(.dina(n148),.dinb(n145),.dout(n149),.clk(gclk));
	jand g077(.dina(w_n149_1[1]),.dinb(w_n141_1[1]),.dout(n150),.clk(gclk));
	jand g078(.dina(n150),.dinb(n133),.dout(n151),.clk(gclk));
	jxor g079(.dina(w_n149_1[0]),.dinb(w_n141_1[0]),.dout(n152),.clk(gclk));
	jand g080(.dina(n152),.dinb(w_n86_0[2]),.dout(n153),.clk(gclk));
	jand g081(.dina(n153),.dinb(w_n132_1[0]),.dout(n154),.clk(gclk));
	jor g082(.dina(n154),.dinb(w_dff_B_L8hwV9M20_1),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_G197gat_0[1]),.dinb(w_G169gat_0[1]),.dout(n156),.clk(gclk));
	jxor g084(.dina(w_G141gat_0[1]),.dinb(w_G113gat_0[1]),.dout(n157),.clk(gclk));
	jxor g085(.dina(n157),.dinb(n156),.dout(n158),.clk(gclk));
	jxor g086(.dina(n158),.dinb(w_n114_0[0]),.dout(n159),.clk(gclk));
	jand g087(.dina(w_G233gat_0[2]),.dinb(G229gat),.dout(n160),.clk(gclk));
	jnot g088(.din(n160),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(w_n100_0[0]),.dout(n162),.clk(gclk));
	jxor g090(.dina(n162),.dinb(n159),.dout(n163),.clk(gclk));
	jnot g091(.din(w_n163_1[1]),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_G204gat_0[1]),.dinb(w_G176gat_0[1]),.dout(n165),.clk(gclk));
	jxor g093(.dina(w_G148gat_0[1]),.dinb(w_G120gat_0[1]),.dout(n166),.clk(gclk));
	jxor g094(.dina(n166),.dinb(n165),.dout(n167),.clk(gclk));
	jxor g095(.dina(n167),.dinb(w_n108_0[0]),.dout(n168),.clk(gclk));
	jand g096(.dina(w_G233gat_0[1]),.dinb(G230gat),.dout(n169),.clk(gclk));
	jnot g097(.din(n169),.dout(n170),.clk(gclk));
	jxor g098(.dina(n170),.dinb(w_n93_0[0]),.dout(n171),.clk(gclk));
	jxor g099(.dina(n171),.dinb(n168),.dout(n172),.clk(gclk));
	jand g100(.dina(w_n172_1[1]),.dinb(w_n164_1[2]),.dout(n173),.clk(gclk));
	jand g101(.dina(w_n173_0[1]),.dinb(w_n155_0[2]),.dout(n174),.clk(gclk));
	jand g102(.dina(n174),.dinb(w_n118_0[1]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_1[1]),.dinb(w_n87_1[2]),.dout(n176),.clk(gclk));
	jxor g104(.dina(n176),.dinb(w_G1gat_0[0]),.dout(G1324gat),.clk(gclk));
	jnot g105(.din(w_n132_0[2]),.dout(n178),.clk(gclk));
	jand g106(.dina(w_n175_1[0]),.dinb(w_n178_1[2]),.dout(n179),.clk(gclk));
	jxor g107(.dina(n179),.dinb(w_G8gat_0[0]),.dout(G1325gat),.clk(gclk));
	jnot g108(.din(w_n141_0[2]),.dout(n181),.clk(gclk));
	jand g109(.dina(w_n175_0[2]),.dinb(w_n181_1[2]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_G15gat_0[0]),.dout(G1326gat),.clk(gclk));
	jnot g111(.din(w_n149_0[2]),.dout(n184),.clk(gclk));
	jand g112(.dina(w_n175_0[1]),.dinb(w_n184_1[2]),.dout(n185),.clk(gclk));
	jxor g113(.dina(n185),.dinb(w_G22gat_0[0]),.dout(G1327gat),.clk(gclk));
	jnot g114(.din(w_n102_1[0]),.dout(n187),.clk(gclk));
	jand g115(.dina(w_n116_1[0]),.dinb(w_n187_1[2]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_dff_B_HukrD1ZN6_0),.dinb(w_n155_0[1]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_n189_0[1]),.dinb(w_n173_0[0]),.dout(n190),.clk(gclk));
	jand g118(.dina(w_n190_1[1]),.dinb(w_n87_1[1]),.dout(n191),.clk(gclk));
	jxor g119(.dina(n191),.dinb(w_G29gat_0[0]),.dout(G1328gat),.clk(gclk));
	jand g120(.dina(w_n190_1[0]),.dinb(w_n178_1[1]),.dout(n193),.clk(gclk));
	jxor g121(.dina(n193),.dinb(w_G36gat_0[0]),.dout(G1329gat),.clk(gclk));
	jand g122(.dina(w_n190_0[2]),.dinb(w_n181_1[1]),.dout(n195),.clk(gclk));
	jxor g123(.dina(n195),.dinb(w_G43gat_0[0]),.dout(G1330gat),.clk(gclk));
	jand g124(.dina(w_n190_0[1]),.dinb(w_n184_1[1]),.dout(n197),.clk(gclk));
	jxor g125(.dina(n197),.dinb(w_G50gat_0[0]),.dout(G1331gat),.clk(gclk));
	jnot g126(.din(w_n172_1[0]),.dout(n199),.clk(gclk));
	jand g127(.dina(w_n199_1[2]),.dinb(w_n163_1[0]),.dout(n200),.clk(gclk));
	jand g128(.dina(w_n155_0[0]),.dinb(w_n118_0[0]),.dout(n201),.clk(gclk));
	jand g129(.dina(n201),.dinb(w_n200_0[1]),.dout(n202),.clk(gclk));
	jand g130(.dina(w_n202_1[1]),.dinb(w_n87_1[0]),.dout(n203),.clk(gclk));
	jxor g131(.dina(n203),.dinb(w_G57gat_0[0]),.dout(G1332gat),.clk(gclk));
	jand g132(.dina(w_n202_1[0]),.dinb(w_n178_1[0]),.dout(n205),.clk(gclk));
	jxor g133(.dina(n205),.dinb(w_G64gat_0[0]),.dout(G1333gat),.clk(gclk));
	jand g134(.dina(w_n202_0[2]),.dinb(w_n181_1[0]),.dout(n207),.clk(gclk));
	jxor g135(.dina(n207),.dinb(w_G71gat_0[0]),.dout(G1334gat),.clk(gclk));
	jand g136(.dina(w_n202_0[1]),.dinb(w_n184_1[0]),.dout(n209),.clk(gclk));
	jxor g137(.dina(n209),.dinb(w_G78gat_0[0]),.dout(G1335gat),.clk(gclk));
	jand g138(.dina(w_n200_0[0]),.dinb(w_n189_0[0]),.dout(n211),.clk(gclk));
	jand g139(.dina(w_n211_1[1]),.dinb(w_n87_0[2]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_G85gat_0[0]),.dout(G1336gat),.clk(gclk));
	jand g141(.dina(w_n211_1[0]),.dinb(w_n178_0[2]),.dout(n214),.clk(gclk));
	jxor g142(.dina(n214),.dinb(w_G92gat_0[0]),.dout(G1337gat),.clk(gclk));
	jand g143(.dina(w_n211_0[2]),.dinb(w_n181_0[2]),.dout(n216),.clk(gclk));
	jxor g144(.dina(n216),.dinb(w_G99gat_0[0]),.dout(G1338gat),.clk(gclk));
	jand g145(.dina(w_n211_0[1]),.dinb(w_n184_0[2]),.dout(n218),.clk(gclk));
	jxor g146(.dina(n218),.dinb(w_G106gat_0[0]),.dout(G1339gat),.clk(gclk));
	jand g147(.dina(w_n149_0[1]),.dinb(w_n181_0[1]),.dout(n220),.clk(gclk));
	jand g148(.dina(w_n132_0[1]),.dinb(w_n87_0[1]),.dout(n221),.clk(gclk));
	jxor g149(.dina(w_n116_0[2]),.dinb(w_n102_0[2]),.dout(n222),.clk(gclk));
	jand g150(.dina(n222),.dinb(w_n163_0[2]),.dout(n223),.clk(gclk));
	jand g151(.dina(n223),.dinb(w_n172_0[2]),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n172_0[1]),.dinb(w_n163_0[1]),.dout(n225),.clk(gclk));
	jand g153(.dina(w_n116_0[1]),.dinb(w_n102_0[1]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(n225),.dout(n227),.clk(gclk));
	jor g155(.dina(w_dff_B_xzTrjmVV4_0),.dinb(n224),.dout(n228),.clk(gclk));
	jand g156(.dina(w_n228_0[1]),.dinb(w_dff_B_e4ssjTZ55_1),.dout(n229),.clk(gclk));
	jand g157(.dina(w_n229_0[1]),.dinb(w_n220_0[1]),.dout(n230),.clk(gclk));
	jand g158(.dina(w_n230_1[1]),.dinb(w_n164_1[1]),.dout(n231),.clk(gclk));
	jxor g159(.dina(n231),.dinb(w_G113gat_0[0]),.dout(G1340gat),.clk(gclk));
	jand g160(.dina(w_n230_1[0]),.dinb(w_n199_1[1]),.dout(n233),.clk(gclk));
	jxor g161(.dina(n233),.dinb(w_G120gat_0[0]),.dout(G1341gat),.clk(gclk));
	jand g162(.dina(w_n230_0[2]),.dinb(w_n117_1[1]),.dout(n235),.clk(gclk));
	jxor g163(.dina(n235),.dinb(w_G127gat_0[0]),.dout(G1342gat),.clk(gclk));
	jand g164(.dina(w_n230_0[1]),.dinb(w_n187_1[1]),.dout(n237),.clk(gclk));
	jxor g165(.dina(n237),.dinb(w_G134gat_0[0]),.dout(G1343gat),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n141_0[1]),.dout(n239),.clk(gclk));
	jand g167(.dina(w_n229_0[0]),.dinb(w_n239_0[1]),.dout(n240),.clk(gclk));
	jand g168(.dina(w_n240_1[1]),.dinb(w_n164_1[0]),.dout(n241),.clk(gclk));
	jxor g169(.dina(n241),.dinb(w_G141gat_0[0]),.dout(G1344gat),.clk(gclk));
	jand g170(.dina(w_n240_1[0]),.dinb(w_n199_1[0]),.dout(n243),.clk(gclk));
	jxor g171(.dina(n243),.dinb(w_G148gat_0[0]),.dout(G1345gat),.clk(gclk));
	jand g172(.dina(w_n240_0[2]),.dinb(w_n117_1[0]),.dout(n245),.clk(gclk));
	jxor g173(.dina(n245),.dinb(w_G155gat_0[0]),.dout(G1346gat),.clk(gclk));
	jand g174(.dina(w_n240_0[1]),.dinb(w_n187_1[0]),.dout(n247),.clk(gclk));
	jxor g175(.dina(n247),.dinb(w_G162gat_0[0]),.dout(G1347gat),.clk(gclk));
	jand g176(.dina(w_n178_0[1]),.dinb(w_n86_0[1]),.dout(n249),.clk(gclk));
	jand g177(.dina(w_n228_0[0]),.dinb(w_dff_B_C9BeA8KM7_1),.dout(n250),.clk(gclk));
	jand g178(.dina(w_n250_0[1]),.dinb(w_n220_0[0]),.dout(n251),.clk(gclk));
	jand g179(.dina(w_n251_1[1]),.dinb(w_n164_0[2]),.dout(n252),.clk(gclk));
	jxor g180(.dina(n252),.dinb(w_G169gat_0[0]),.dout(G1348gat),.clk(gclk));
	jand g181(.dina(w_n251_1[0]),.dinb(w_n199_0[2]),.dout(n254),.clk(gclk));
	jxor g182(.dina(n254),.dinb(w_G176gat_0[0]),.dout(G1349gat),.clk(gclk));
	jand g183(.dina(w_n251_0[2]),.dinb(w_n117_0[2]),.dout(n256),.clk(gclk));
	jxor g184(.dina(n256),.dinb(w_G183gat_0[0]),.dout(G1350gat),.clk(gclk));
	jand g185(.dina(w_n251_0[1]),.dinb(w_n187_0[2]),.dout(n258),.clk(gclk));
	jxor g186(.dina(n258),.dinb(w_G190gat_0[0]),.dout(G1351gat),.clk(gclk));
	jand g187(.dina(w_n250_0[0]),.dinb(w_n239_0[0]),.dout(n260),.clk(gclk));
	jand g188(.dina(w_n260_1[1]),.dinb(w_n164_0[1]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_G197gat_0[0]),.dout(G1352gat),.clk(gclk));
	jand g190(.dina(w_n260_1[0]),.dinb(w_n199_0[1]),.dout(n263),.clk(gclk));
	jxor g191(.dina(n263),.dinb(w_G204gat_0[0]),.dout(G1353gat),.clk(gclk));
	jand g192(.dina(w_n260_0[2]),.dinb(w_n117_0[1]),.dout(n265),.clk(gclk));
	jxor g193(.dina(n265),.dinb(w_G211gat_0[0]),.dout(G1354gat),.clk(gclk));
	jand g194(.dina(w_n260_0[1]),.dinb(w_n187_0[1]),.dout(n267),.clk(gclk));
	jxor g195(.dina(n267),.dinb(w_G218gat_0[0]),.dout(G1355gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_q3IXA9W52_0),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_mMj5LMFW2_0),.doutb(w_G8gat_0[1]),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G15gat_0(.douta(w_dff_A_9Zmys9zm8_0),.doutb(w_G15gat_0[1]),.doutc(w_G15gat_0[2]),.din(G15gat));
	jspl3 jspl3_w_G22gat_0(.douta(w_dff_A_9QQ3fZkz9_0),.doutb(w_G22gat_0[1]),.doutc(w_G22gat_0[2]),.din(G22gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_i5GnN5Yd6_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl3 jspl3_w_G36gat_0(.douta(w_dff_A_M9pBSjVC9_0),.doutb(w_G36gat_0[1]),.doutc(w_G36gat_0[2]),.din(G36gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_dff_A_iqz6IBc73_0),.doutb(w_G43gat_0[1]),.doutc(w_G43gat_0[2]),.din(G43gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_horf3TtB3_0),.doutb(w_G50gat_0[1]),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl3 jspl3_w_G57gat_0(.douta(w_dff_A_9XxXW3xX6_0),.doutb(w_G57gat_0[1]),.doutc(w_G57gat_0[2]),.din(G57gat));
	jspl3 jspl3_w_G64gat_0(.douta(w_dff_A_zxy5Nh8h9_0),.doutb(w_G64gat_0[1]),.doutc(w_G64gat_0[2]),.din(G64gat));
	jspl3 jspl3_w_G71gat_0(.douta(w_dff_A_wNbvbPej9_0),.doutb(w_G71gat_0[1]),.doutc(w_G71gat_0[2]),.din(G71gat));
	jspl3 jspl3_w_G78gat_0(.douta(w_dff_A_BwzKoTGC1_0),.doutb(w_G78gat_0[1]),.doutc(w_G78gat_0[2]),.din(G78gat));
	jspl3 jspl3_w_G85gat_0(.douta(w_dff_A_ogvUz4vm1_0),.doutb(w_G85gat_0[1]),.doutc(w_G85gat_0[2]),.din(G85gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_J8e7MW7e3_0),.doutb(w_G92gat_0[1]),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_p1F05AkQ9_0),.doutb(w_G99gat_0[1]),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_zEYHoXXM2_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G113gat_0(.douta(w_dff_A_uiifWNTX9_0),.doutb(w_G113gat_0[1]),.doutc(w_G113gat_0[2]),.din(G113gat));
	jspl3 jspl3_w_G120gat_0(.douta(w_dff_A_ZuYfv5UA5_0),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G127gat_0(.douta(w_dff_A_k98m0A6N9_0),.doutb(w_G127gat_0[1]),.doutc(w_G127gat_0[2]),.din(G127gat));
	jspl3 jspl3_w_G134gat_0(.douta(w_dff_A_veYjb4335_0),.doutb(w_G134gat_0[1]),.doutc(w_G134gat_0[2]),.din(G134gat));
	jspl3 jspl3_w_G141gat_0(.douta(w_dff_A_jysE7TwX7_0),.doutb(w_G141gat_0[1]),.doutc(w_G141gat_0[2]),.din(G141gat));
	jspl3 jspl3_w_G148gat_0(.douta(w_dff_A_QUevK6dp3_0),.doutb(w_G148gat_0[1]),.doutc(w_G148gat_0[2]),.din(G148gat));
	jspl3 jspl3_w_G155gat_0(.douta(w_dff_A_ngdY3SaI8_0),.doutb(w_G155gat_0[1]),.doutc(w_G155gat_0[2]),.din(G155gat));
	jspl3 jspl3_w_G162gat_0(.douta(w_dff_A_XAMCx2EQ4_0),.doutb(w_G162gat_0[1]),.doutc(w_G162gat_0[2]),.din(G162gat));
	jspl3 jspl3_w_G169gat_0(.douta(w_dff_A_FKRrwreq2_0),.doutb(w_G169gat_0[1]),.doutc(w_G169gat_0[2]),.din(G169gat));
	jspl3 jspl3_w_G176gat_0(.douta(w_dff_A_DXT6JGjF6_0),.doutb(w_G176gat_0[1]),.doutc(w_G176gat_0[2]),.din(G176gat));
	jspl3 jspl3_w_G183gat_0(.douta(w_dff_A_l7QUQJ4y2_0),.doutb(w_G183gat_0[1]),.doutc(w_G183gat_0[2]),.din(G183gat));
	jspl3 jspl3_w_G190gat_0(.douta(w_dff_A_9BZA5ENF8_0),.doutb(w_G190gat_0[1]),.doutc(w_G190gat_0[2]),.din(G190gat));
	jspl3 jspl3_w_G197gat_0(.douta(w_dff_A_Gwy7oFm21_0),.doutb(w_G197gat_0[1]),.doutc(w_G197gat_0[2]),.din(G197gat));
	jspl3 jspl3_w_G204gat_0(.douta(w_dff_A_KrOmtTGV2_0),.doutb(w_G204gat_0[1]),.doutc(w_G204gat_0[2]),.din(G204gat));
	jspl3 jspl3_w_G211gat_0(.douta(w_dff_A_lMiBnJV77_0),.doutb(w_G211gat_0[1]),.doutc(w_G211gat_0[2]),.din(G211gat));
	jspl3 jspl3_w_G218gat_0(.douta(w_dff_A_odWp6WvU9_0),.doutb(w_G218gat_0[1]),.doutc(w_G218gat_0[2]),.din(G218gat));
	jspl3 jspl3_w_G233gat_0(.douta(w_G233gat_0[0]),.doutb(w_G233gat_0[1]),.doutc(w_G233gat_0[2]),.din(G233gat));
	jspl3 jspl3_w_G233gat_1(.douta(w_G233gat_1[0]),.doutb(w_G233gat_1[1]),.doutc(w_G233gat_1[2]),.din(w_G233gat_0[0]));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n86_0(.douta(w_n86_0[0]),.doutb(w_dff_A_JeFRJKoD5_1),.doutc(w_dff_A_YsSOuQPd4_2),.din(n86));
	jspl jspl_w_n86_1(.douta(w_n86_1[0]),.doutb(w_n86_1[1]),.din(w_n86_0[0]));
	jspl3 jspl3_w_n87_0(.douta(w_dff_A_9LSOWbPS8_0),.doutb(w_n87_0[1]),.doutc(w_dff_A_bfNkBzqG1_2),.din(n87));
	jspl3 jspl3_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.doutc(w_n87_1[2]),.din(w_n87_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl jspl_w_n96_1(.douta(w_n96_1[0]),.doutb(w_n96_1[1]),.din(w_n96_0[0]));
	jspl jspl_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.din(n100));
	jspl3 jspl3_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.doutc(w_n102_0[2]),.din(n102));
	jspl jspl_w_n102_1(.douta(w_n102_1[0]),.doutb(w_dff_A_ObRYbEa95_1),.din(w_n102_0[0]));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n114_0(.douta(w_n114_0[0]),.doutb(w_n114_0[1]),.din(n114));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl jspl_w_n116_1(.douta(w_dff_A_lQZyNmHG3_0),.doutb(w_n116_1[1]),.din(w_n116_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_3Rfm1gUM6_1),.doutc(w_dff_A_TTNNcIoX3_2),.din(n117));
	jspl3 jspl3_w_n117_1(.douta(w_dff_A_fozk3laX3_0),.doutb(w_dff_A_Xb55nq249_1),.doutc(w_n117_1[2]),.din(w_n117_0[0]));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_dff_A_AS5DiFPi6_1),.din(w_dff_B_zvAI8Bn44_2));
	jspl jspl_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.din(n124));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_dff_A_bMqIfJaP7_1),.doutc(w_n132_0[2]),.din(n132));
	jspl jspl_w_n132_1(.douta(w_dff_A_Sdvdv2ww4_0),.doutb(w_n132_1[1]),.din(w_n132_0[0]));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_dff_A_ijYXtsu43_1),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_dff_A_mOfIDB2G0_1),.doutc(w_n149_0[2]),.din(n149));
	jspl jspl_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.din(w_n149_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_dff_A_BgzgqeGf9_2),.din(n163));
	jspl jspl_w_n163_1(.douta(w_dff_A_nApm0Jzs2_0),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_dff_A_I29TAoUH3_1),.doutc(w_dff_A_aKl7Y1CB7_2),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_dff_A_FyMtaAU47_0),.doutb(w_dff_A_vgv1IbVN6_1),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.doutc(w_dff_A_EyhmX1MY6_2),.din(n172));
	jspl jspl_w_n172_1(.douta(w_n172_1[0]),.doutb(w_dff_A_1KuXAB0J0_1),.din(w_n172_0[0]));
	jspl jspl_w_n173_0(.douta(w_dff_A_8JuFjjCQ2_0),.doutb(w_n173_0[1]),.din(w_dff_B_am6g3HwZ6_2));
	jspl3 jspl3_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.doutc(w_n175_0[2]),.din(n175));
	jspl jspl_w_n175_1(.douta(w_n175_1[0]),.doutb(w_n175_1[1]),.din(w_n175_0[0]));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_oS4wZYHo2_0),.doutb(w_n178_0[1]),.doutc(w_dff_A_ZWHn74Gi5_2),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n181_0(.douta(w_dff_A_eb0E6ue46_0),.doutb(w_n181_0[1]),.doutc(w_dff_A_JsXhfJE76_2),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n184_0(.douta(w_dff_A_A5YsYjkw6_0),.doutb(w_n184_0[1]),.doutc(w_dff_A_GTn9ZlPg9_2),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.doutc(w_n184_1[2]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_n187_0[0]),.doutb(w_dff_A_4G4z2rLk7_1),.doutc(w_dff_A_TWxn2FOh5_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_dff_A_1EwuVeVU7_0),.doutb(w_dff_A_QQ4lHGA13_1),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl jspl_w_n190_1(.douta(w_n190_1[0]),.doutb(w_n190_1[1]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_dff_A_RKWXYvMO3_1),.doutc(w_dff_A_nCJDKVfu2_2),.din(n199));
	jspl3 jspl3_w_n199_1(.douta(w_dff_A_SWUusfbe4_0),.doutb(w_dff_A_9dMBYRhg5_1),.doutc(w_n199_1[2]),.din(w_n199_0[0]));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(w_dff_B_xvKMKOjR6_2));
	jspl3 jspl3_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.doutc(w_n202_0[2]),.din(n202));
	jspl jspl_w_n202_1(.douta(w_n202_1[0]),.doutb(w_n202_1[1]),.din(w_n202_0[0]));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(w_dff_B_YnP07Vuw0_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl jspl_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.din(w_n230_0[0]));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(w_dff_B_mgU9srBl5_2));
	jspl3 jspl3_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.doutc(w_n240_0[2]),.din(n240));
	jspl jspl_w_n240_1(.douta(w_n240_1[0]),.doutb(w_n240_1[1]),.din(w_n240_0[0]));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl jspl_w_n251_1(.douta(w_n251_1[0]),.doutb(w_n251_1[1]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.doutc(w_n260_0[2]),.din(n260));
	jspl jspl_w_n260_1(.douta(w_n260_1[0]),.doutb(w_n260_1[1]),.din(w_n260_0[0]));
	jdff dff_A_8JuFjjCQ2_0(.dout(w_n173_0[0]),.din(w_dff_A_8JuFjjCQ2_0),.clk(gclk));
	jdff dff_B_8NUdgw8m9_2(.din(n173),.dout(w_dff_B_8NUdgw8m9_2),.clk(gclk));
	jdff dff_B_am6g3HwZ6_2(.din(w_dff_B_8NUdgw8m9_2),.dout(w_dff_B_am6g3HwZ6_2),.clk(gclk));
	jdff dff_A_AS5DiFPi6_1(.dout(w_n118_0[1]),.din(w_dff_A_AS5DiFPi6_1),.clk(gclk));
	jdff dff_B_icqtxdVr5_2(.din(n118),.dout(w_dff_B_icqtxdVr5_2),.clk(gclk));
	jdff dff_B_zvAI8Bn44_2(.din(w_dff_B_icqtxdVr5_2),.dout(w_dff_B_zvAI8Bn44_2),.clk(gclk));
	jdff dff_B_HX8pgkMt4_2(.din(n200),.dout(w_dff_B_HX8pgkMt4_2),.clk(gclk));
	jdff dff_B_Ao3mF6jD5_2(.din(w_dff_B_HX8pgkMt4_2),.dout(w_dff_B_Ao3mF6jD5_2),.clk(gclk));
	jdff dff_B_xvKMKOjR6_2(.din(w_dff_B_Ao3mF6jD5_2),.dout(w_dff_B_xvKMKOjR6_2),.clk(gclk));
	jdff dff_B_5mJw1h9l2_0(.din(n188),.dout(w_dff_B_5mJw1h9l2_0),.clk(gclk));
	jdff dff_B_HukrD1ZN6_0(.din(w_dff_B_5mJw1h9l2_0),.dout(w_dff_B_HukrD1ZN6_0),.clk(gclk));
	jdff dff_B_L8hwV9M20_1(.din(n151),.dout(w_dff_B_L8hwV9M20_1),.clk(gclk));
	jdff dff_A_CuTx14e61_0(.dout(w_n132_1[0]),.din(w_dff_A_CuTx14e61_0),.clk(gclk));
	jdff dff_A_Sdvdv2ww4_0(.dout(w_dff_A_CuTx14e61_0),.din(w_dff_A_Sdvdv2ww4_0),.clk(gclk));
	jdff dff_A_q9i9M5zw9_0(.dout(w_n164_1[0]),.din(w_dff_A_q9i9M5zw9_0),.clk(gclk));
	jdff dff_A_bBfmBw576_0(.dout(w_dff_A_q9i9M5zw9_0),.din(w_dff_A_bBfmBw576_0),.clk(gclk));
	jdff dff_A_CYjvTZXb0_0(.dout(w_dff_A_bBfmBw576_0),.din(w_dff_A_CYjvTZXb0_0),.clk(gclk));
	jdff dff_A_qrJVjDxM4_0(.dout(w_dff_A_CYjvTZXb0_0),.din(w_dff_A_qrJVjDxM4_0),.clk(gclk));
	jdff dff_A_FyMtaAU47_0(.dout(w_dff_A_qrJVjDxM4_0),.din(w_dff_A_FyMtaAU47_0),.clk(gclk));
	jdff dff_A_fT9dh2oP6_1(.dout(w_n164_1[1]),.din(w_dff_A_fT9dh2oP6_1),.clk(gclk));
	jdff dff_A_a7y40y1C5_1(.dout(w_dff_A_fT9dh2oP6_1),.din(w_dff_A_a7y40y1C5_1),.clk(gclk));
	jdff dff_A_mYLiq6mY2_1(.dout(w_dff_A_a7y40y1C5_1),.din(w_dff_A_mYLiq6mY2_1),.clk(gclk));
	jdff dff_A_6X2jNa6m2_1(.dout(w_dff_A_mYLiq6mY2_1),.din(w_dff_A_6X2jNa6m2_1),.clk(gclk));
	jdff dff_A_vgv1IbVN6_1(.dout(w_dff_A_6X2jNa6m2_1),.din(w_dff_A_vgv1IbVN6_1),.clk(gclk));
	jdff dff_A_L20QRunt7_0(.dout(w_n199_1[0]),.din(w_dff_A_L20QRunt7_0),.clk(gclk));
	jdff dff_A_zaRGelBp6_0(.dout(w_dff_A_L20QRunt7_0),.din(w_dff_A_zaRGelBp6_0),.clk(gclk));
	jdff dff_A_9Y8Y2EZM4_0(.dout(w_dff_A_zaRGelBp6_0),.din(w_dff_A_9Y8Y2EZM4_0),.clk(gclk));
	jdff dff_A_pHHr8qCy1_0(.dout(w_dff_A_9Y8Y2EZM4_0),.din(w_dff_A_pHHr8qCy1_0),.clk(gclk));
	jdff dff_A_SWUusfbe4_0(.dout(w_dff_A_pHHr8qCy1_0),.din(w_dff_A_SWUusfbe4_0),.clk(gclk));
	jdff dff_A_O57MIXbh7_1(.dout(w_n199_1[1]),.din(w_dff_A_O57MIXbh7_1),.clk(gclk));
	jdff dff_A_bz85RdKA4_1(.dout(w_dff_A_O57MIXbh7_1),.din(w_dff_A_bz85RdKA4_1),.clk(gclk));
	jdff dff_A_STu1RUb93_1(.dout(w_dff_A_bz85RdKA4_1),.din(w_dff_A_STu1RUb93_1),.clk(gclk));
	jdff dff_A_LXuHtb6K8_1(.dout(w_dff_A_STu1RUb93_1),.din(w_dff_A_LXuHtb6K8_1),.clk(gclk));
	jdff dff_A_9dMBYRhg5_1(.dout(w_dff_A_LXuHtb6K8_1),.din(w_dff_A_9dMBYRhg5_1),.clk(gclk));
	jdff dff_A_sEZ1BWzB8_0(.dout(w_n117_1[0]),.din(w_dff_A_sEZ1BWzB8_0),.clk(gclk));
	jdff dff_A_Fh30niyP0_0(.dout(w_dff_A_sEZ1BWzB8_0),.din(w_dff_A_Fh30niyP0_0),.clk(gclk));
	jdff dff_A_2lnlPTc33_0(.dout(w_dff_A_Fh30niyP0_0),.din(w_dff_A_2lnlPTc33_0),.clk(gclk));
	jdff dff_A_NTJGSX5p8_0(.dout(w_dff_A_2lnlPTc33_0),.din(w_dff_A_NTJGSX5p8_0),.clk(gclk));
	jdff dff_A_fozk3laX3_0(.dout(w_dff_A_NTJGSX5p8_0),.din(w_dff_A_fozk3laX3_0),.clk(gclk));
	jdff dff_A_GTG0p0QH6_1(.dout(w_n117_1[1]),.din(w_dff_A_GTG0p0QH6_1),.clk(gclk));
	jdff dff_A_KWRa1ulO8_1(.dout(w_dff_A_GTG0p0QH6_1),.din(w_dff_A_KWRa1ulO8_1),.clk(gclk));
	jdff dff_A_vy53priu5_1(.dout(w_dff_A_KWRa1ulO8_1),.din(w_dff_A_vy53priu5_1),.clk(gclk));
	jdff dff_A_A6Z2XqIo9_1(.dout(w_dff_A_vy53priu5_1),.din(w_dff_A_A6Z2XqIo9_1),.clk(gclk));
	jdff dff_A_Xb55nq249_1(.dout(w_dff_A_A6Z2XqIo9_1),.din(w_dff_A_Xb55nq249_1),.clk(gclk));
	jdff dff_B_yIG8Xxhd6_1(.din(n221),.dout(w_dff_B_yIG8Xxhd6_1),.clk(gclk));
	jdff dff_B_e4ssjTZ55_1(.din(w_dff_B_yIG8Xxhd6_1),.dout(w_dff_B_e4ssjTZ55_1),.clk(gclk));
	jdff dff_A_9TBx4ji69_0(.dout(w_n87_0[0]),.din(w_dff_A_9TBx4ji69_0),.clk(gclk));
	jdff dff_A_noTTOzMr3_0(.dout(w_dff_A_9TBx4ji69_0),.din(w_dff_A_noTTOzMr3_0),.clk(gclk));
	jdff dff_A_oX3TABZB0_0(.dout(w_dff_A_noTTOzMr3_0),.din(w_dff_A_oX3TABZB0_0),.clk(gclk));
	jdff dff_A_Wn2kC3ox6_0(.dout(w_dff_A_oX3TABZB0_0),.din(w_dff_A_Wn2kC3ox6_0),.clk(gclk));
	jdff dff_A_9LSOWbPS8_0(.dout(w_dff_A_Wn2kC3ox6_0),.din(w_dff_A_9LSOWbPS8_0),.clk(gclk));
	jdff dff_A_VhTbhjy14_2(.dout(w_n87_0[2]),.din(w_dff_A_VhTbhjy14_2),.clk(gclk));
	jdff dff_A_EeJvPDNh1_2(.dout(w_dff_A_VhTbhjy14_2),.din(w_dff_A_EeJvPDNh1_2),.clk(gclk));
	jdff dff_A_Q9hIvtog2_2(.dout(w_dff_A_EeJvPDNh1_2),.din(w_dff_A_Q9hIvtog2_2),.clk(gclk));
	jdff dff_A_CrbgB4IN2_2(.dout(w_dff_A_Q9hIvtog2_2),.din(w_dff_A_CrbgB4IN2_2),.clk(gclk));
	jdff dff_A_bfNkBzqG1_2(.dout(w_dff_A_CrbgB4IN2_2),.din(w_dff_A_bfNkBzqG1_2),.clk(gclk));
	jdff dff_A_WIcU59q00_0(.dout(w_n187_1[0]),.din(w_dff_A_WIcU59q00_0),.clk(gclk));
	jdff dff_A_vNqZzioz3_0(.dout(w_dff_A_WIcU59q00_0),.din(w_dff_A_vNqZzioz3_0),.clk(gclk));
	jdff dff_A_3fjB3M6l9_0(.dout(w_dff_A_vNqZzioz3_0),.din(w_dff_A_3fjB3M6l9_0),.clk(gclk));
	jdff dff_A_YvSJDBRq8_0(.dout(w_dff_A_3fjB3M6l9_0),.din(w_dff_A_YvSJDBRq8_0),.clk(gclk));
	jdff dff_A_1EwuVeVU7_0(.dout(w_dff_A_YvSJDBRq8_0),.din(w_dff_A_1EwuVeVU7_0),.clk(gclk));
	jdff dff_A_Y5gXd9006_1(.dout(w_n187_1[1]),.din(w_dff_A_Y5gXd9006_1),.clk(gclk));
	jdff dff_A_XRZTSRNe1_1(.dout(w_dff_A_Y5gXd9006_1),.din(w_dff_A_XRZTSRNe1_1),.clk(gclk));
	jdff dff_A_0HTn2Dt71_1(.dout(w_dff_A_XRZTSRNe1_1),.din(w_dff_A_0HTn2Dt71_1),.clk(gclk));
	jdff dff_A_72m1i4TZ8_1(.dout(w_dff_A_0HTn2Dt71_1),.din(w_dff_A_72m1i4TZ8_1),.clk(gclk));
	jdff dff_A_QQ4lHGA13_1(.dout(w_dff_A_72m1i4TZ8_1),.din(w_dff_A_QQ4lHGA13_1),.clk(gclk));
	jdff dff_B_nemRtXzG4_2(.din(n220),.dout(w_dff_B_nemRtXzG4_2),.clk(gclk));
	jdff dff_B_cNMapHAP6_2(.din(w_dff_B_nemRtXzG4_2),.dout(w_dff_B_cNMapHAP6_2),.clk(gclk));
	jdff dff_B_YnP07Vuw0_2(.din(w_dff_B_cNMapHAP6_2),.dout(w_dff_B_YnP07Vuw0_2),.clk(gclk));
	jdff dff_A_5OuMraU69_0(.dout(w_n181_0[0]),.din(w_dff_A_5OuMraU69_0),.clk(gclk));
	jdff dff_A_TLbyTtBw5_0(.dout(w_dff_A_5OuMraU69_0),.din(w_dff_A_TLbyTtBw5_0),.clk(gclk));
	jdff dff_A_4klv3bXp6_0(.dout(w_dff_A_TLbyTtBw5_0),.din(w_dff_A_4klv3bXp6_0),.clk(gclk));
	jdff dff_A_9FEDRJlK1_0(.dout(w_dff_A_4klv3bXp6_0),.din(w_dff_A_9FEDRJlK1_0),.clk(gclk));
	jdff dff_A_eb0E6ue46_0(.dout(w_dff_A_9FEDRJlK1_0),.din(w_dff_A_eb0E6ue46_0),.clk(gclk));
	jdff dff_A_0Joc3Vii4_2(.dout(w_n181_0[2]),.din(w_dff_A_0Joc3Vii4_2),.clk(gclk));
	jdff dff_A_qng5xjpf1_2(.dout(w_dff_A_0Joc3Vii4_2),.din(w_dff_A_qng5xjpf1_2),.clk(gclk));
	jdff dff_A_K1OUCfD43_2(.dout(w_dff_A_qng5xjpf1_2),.din(w_dff_A_K1OUCfD43_2),.clk(gclk));
	jdff dff_A_9HRfUdej9_2(.dout(w_dff_A_K1OUCfD43_2),.din(w_dff_A_9HRfUdej9_2),.clk(gclk));
	jdff dff_A_JsXhfJE76_2(.dout(w_dff_A_9HRfUdej9_2),.din(w_dff_A_JsXhfJE76_2),.clk(gclk));
	jdff dff_A_EWZzrm5V2_1(.dout(w_n164_0[1]),.din(w_dff_A_EWZzrm5V2_1),.clk(gclk));
	jdff dff_A_w8oUgXdQ0_1(.dout(w_dff_A_EWZzrm5V2_1),.din(w_dff_A_w8oUgXdQ0_1),.clk(gclk));
	jdff dff_A_lJoPA1BP5_1(.dout(w_dff_A_w8oUgXdQ0_1),.din(w_dff_A_lJoPA1BP5_1),.clk(gclk));
	jdff dff_A_JG5HPrIz9_1(.dout(w_dff_A_lJoPA1BP5_1),.din(w_dff_A_JG5HPrIz9_1),.clk(gclk));
	jdff dff_A_I29TAoUH3_1(.dout(w_dff_A_JG5HPrIz9_1),.din(w_dff_A_I29TAoUH3_1),.clk(gclk));
	jdff dff_A_qM65IoOa8_2(.dout(w_n164_0[2]),.din(w_dff_A_qM65IoOa8_2),.clk(gclk));
	jdff dff_A_ZI4Jn9Nr1_2(.dout(w_dff_A_qM65IoOa8_2),.din(w_dff_A_ZI4Jn9Nr1_2),.clk(gclk));
	jdff dff_A_KBequAQw6_2(.dout(w_dff_A_ZI4Jn9Nr1_2),.din(w_dff_A_KBequAQw6_2),.clk(gclk));
	jdff dff_A_wOdA5qfh8_2(.dout(w_dff_A_KBequAQw6_2),.din(w_dff_A_wOdA5qfh8_2),.clk(gclk));
	jdff dff_A_aKl7Y1CB7_2(.dout(w_dff_A_wOdA5qfh8_2),.din(w_dff_A_aKl7Y1CB7_2),.clk(gclk));
	jdff dff_A_nApm0Jzs2_0(.dout(w_n163_1[0]),.din(w_dff_A_nApm0Jzs2_0),.clk(gclk));
	jdff dff_A_nDFyIYZ49_1(.dout(w_n199_0[1]),.din(w_dff_A_nDFyIYZ49_1),.clk(gclk));
	jdff dff_A_esT7zxR70_1(.dout(w_dff_A_nDFyIYZ49_1),.din(w_dff_A_esT7zxR70_1),.clk(gclk));
	jdff dff_A_k2S79Kwl5_1(.dout(w_dff_A_esT7zxR70_1),.din(w_dff_A_k2S79Kwl5_1),.clk(gclk));
	jdff dff_A_ED9ixB6q2_1(.dout(w_dff_A_k2S79Kwl5_1),.din(w_dff_A_ED9ixB6q2_1),.clk(gclk));
	jdff dff_A_RKWXYvMO3_1(.dout(w_dff_A_ED9ixB6q2_1),.din(w_dff_A_RKWXYvMO3_1),.clk(gclk));
	jdff dff_A_YtOrFiTv2_2(.dout(w_n199_0[2]),.din(w_dff_A_YtOrFiTv2_2),.clk(gclk));
	jdff dff_A_hZgvwz5H1_2(.dout(w_dff_A_YtOrFiTv2_2),.din(w_dff_A_hZgvwz5H1_2),.clk(gclk));
	jdff dff_A_olcDohVr6_2(.dout(w_dff_A_hZgvwz5H1_2),.din(w_dff_A_olcDohVr6_2),.clk(gclk));
	jdff dff_A_0pmU4C2a3_2(.dout(w_dff_A_olcDohVr6_2),.din(w_dff_A_0pmU4C2a3_2),.clk(gclk));
	jdff dff_A_nCJDKVfu2_2(.dout(w_dff_A_0pmU4C2a3_2),.din(w_dff_A_nCJDKVfu2_2),.clk(gclk));
	jdff dff_A_1KuXAB0J0_1(.dout(w_n172_1[1]),.din(w_dff_A_1KuXAB0J0_1),.clk(gclk));
	jdff dff_A_xTJyjQSd0_1(.dout(w_n117_0[1]),.din(w_dff_A_xTJyjQSd0_1),.clk(gclk));
	jdff dff_A_sFsaMdu40_1(.dout(w_dff_A_xTJyjQSd0_1),.din(w_dff_A_sFsaMdu40_1),.clk(gclk));
	jdff dff_A_8fbEma5R7_1(.dout(w_dff_A_sFsaMdu40_1),.din(w_dff_A_8fbEma5R7_1),.clk(gclk));
	jdff dff_A_0owp1E3X3_1(.dout(w_dff_A_8fbEma5R7_1),.din(w_dff_A_0owp1E3X3_1),.clk(gclk));
	jdff dff_A_3Rfm1gUM6_1(.dout(w_dff_A_0owp1E3X3_1),.din(w_dff_A_3Rfm1gUM6_1),.clk(gclk));
	jdff dff_A_dNaCs9U53_2(.dout(w_n117_0[2]),.din(w_dff_A_dNaCs9U53_2),.clk(gclk));
	jdff dff_A_DJ03KHzt2_2(.dout(w_dff_A_dNaCs9U53_2),.din(w_dff_A_DJ03KHzt2_2),.clk(gclk));
	jdff dff_A_7KyCDYpz0_2(.dout(w_dff_A_DJ03KHzt2_2),.din(w_dff_A_7KyCDYpz0_2),.clk(gclk));
	jdff dff_A_ggwqiEHo5_2(.dout(w_dff_A_7KyCDYpz0_2),.din(w_dff_A_ggwqiEHo5_2),.clk(gclk));
	jdff dff_A_TTNNcIoX3_2(.dout(w_dff_A_ggwqiEHo5_2),.din(w_dff_A_TTNNcIoX3_2),.clk(gclk));
	jdff dff_A_lQZyNmHG3_0(.dout(w_n116_1[0]),.din(w_dff_A_lQZyNmHG3_0),.clk(gclk));
	jdff dff_B_cpb3gZPs5_1(.din(n249),.dout(w_dff_B_cpb3gZPs5_1),.clk(gclk));
	jdff dff_B_C9BeA8KM7_1(.din(w_dff_B_cpb3gZPs5_1),.dout(w_dff_B_C9BeA8KM7_1),.clk(gclk));
	jdff dff_B_xzTrjmVV4_0(.din(n227),.dout(w_dff_B_xzTrjmVV4_0),.clk(gclk));
	jdff dff_A_BgzgqeGf9_2(.dout(w_n163_0[2]),.din(w_dff_A_BgzgqeGf9_2),.clk(gclk));
	jdff dff_A_oF1y5N940_2(.dout(w_n172_0[2]),.din(w_dff_A_oF1y5N940_2),.clk(gclk));
	jdff dff_A_EyhmX1MY6_2(.dout(w_dff_A_oF1y5N940_2),.din(w_dff_A_EyhmX1MY6_2),.clk(gclk));
	jdff dff_A_28Nizbl97_0(.dout(w_n178_0[0]),.din(w_dff_A_28Nizbl97_0),.clk(gclk));
	jdff dff_A_q8tswYZT7_0(.dout(w_dff_A_28Nizbl97_0),.din(w_dff_A_q8tswYZT7_0),.clk(gclk));
	jdff dff_A_1BnerfKd7_0(.dout(w_dff_A_q8tswYZT7_0),.din(w_dff_A_1BnerfKd7_0),.clk(gclk));
	jdff dff_A_8VSuDl4t1_0(.dout(w_dff_A_1BnerfKd7_0),.din(w_dff_A_8VSuDl4t1_0),.clk(gclk));
	jdff dff_A_oS4wZYHo2_0(.dout(w_dff_A_8VSuDl4t1_0),.din(w_dff_A_oS4wZYHo2_0),.clk(gclk));
	jdff dff_A_Gc94o9pn1_2(.dout(w_n178_0[2]),.din(w_dff_A_Gc94o9pn1_2),.clk(gclk));
	jdff dff_A_rUMWj6Xa2_2(.dout(w_dff_A_Gc94o9pn1_2),.din(w_dff_A_rUMWj6Xa2_2),.clk(gclk));
	jdff dff_A_ta2rhT3d4_2(.dout(w_dff_A_rUMWj6Xa2_2),.din(w_dff_A_ta2rhT3d4_2),.clk(gclk));
	jdff dff_A_1EWKPCFS3_2(.dout(w_dff_A_ta2rhT3d4_2),.din(w_dff_A_1EWKPCFS3_2),.clk(gclk));
	jdff dff_A_ZWHn74Gi5_2(.dout(w_dff_A_1EWKPCFS3_2),.din(w_dff_A_ZWHn74Gi5_2),.clk(gclk));
	jdff dff_A_bMqIfJaP7_1(.dout(w_n132_0[1]),.din(w_dff_A_bMqIfJaP7_1),.clk(gclk));
	jdff dff_A_Gy2CJJnj2_0(.dout(w_G8gat_0[0]),.din(w_dff_A_Gy2CJJnj2_0),.clk(gclk));
	jdff dff_A_Waq2GnRU5_0(.dout(w_dff_A_Gy2CJJnj2_0),.din(w_dff_A_Waq2GnRU5_0),.clk(gclk));
	jdff dff_A_rIbPlINT4_0(.dout(w_dff_A_Waq2GnRU5_0),.din(w_dff_A_rIbPlINT4_0),.clk(gclk));
	jdff dff_A_mYQpjEIT1_0(.dout(w_dff_A_rIbPlINT4_0),.din(w_dff_A_mYQpjEIT1_0),.clk(gclk));
	jdff dff_A_MUecw0188_0(.dout(w_dff_A_mYQpjEIT1_0),.din(w_dff_A_MUecw0188_0),.clk(gclk));
	jdff dff_A_rp1YaFq33_0(.dout(w_dff_A_MUecw0188_0),.din(w_dff_A_rp1YaFq33_0),.clk(gclk));
	jdff dff_A_9ql2u9ZS2_0(.dout(w_dff_A_rp1YaFq33_0),.din(w_dff_A_9ql2u9ZS2_0),.clk(gclk));
	jdff dff_A_VEU5HbcK8_0(.dout(w_dff_A_9ql2u9ZS2_0),.din(w_dff_A_VEU5HbcK8_0),.clk(gclk));
	jdff dff_A_2OfhNg3O0_0(.dout(w_dff_A_VEU5HbcK8_0),.din(w_dff_A_2OfhNg3O0_0),.clk(gclk));
	jdff dff_A_GuJuuoNy3_0(.dout(w_dff_A_2OfhNg3O0_0),.din(w_dff_A_GuJuuoNy3_0),.clk(gclk));
	jdff dff_A_mMj5LMFW2_0(.dout(w_dff_A_GuJuuoNy3_0),.din(w_dff_A_mMj5LMFW2_0),.clk(gclk));
	jdff dff_A_RTpFpdC09_0(.dout(w_G64gat_0[0]),.din(w_dff_A_RTpFpdC09_0),.clk(gclk));
	jdff dff_A_6vFxHHfd4_0(.dout(w_dff_A_RTpFpdC09_0),.din(w_dff_A_6vFxHHfd4_0),.clk(gclk));
	jdff dff_A_oZG3wzxO0_0(.dout(w_dff_A_6vFxHHfd4_0),.din(w_dff_A_oZG3wzxO0_0),.clk(gclk));
	jdff dff_A_Ag32BBoU1_0(.dout(w_dff_A_oZG3wzxO0_0),.din(w_dff_A_Ag32BBoU1_0),.clk(gclk));
	jdff dff_A_VQr5k33k2_0(.dout(w_dff_A_Ag32BBoU1_0),.din(w_dff_A_VQr5k33k2_0),.clk(gclk));
	jdff dff_A_iu6nTUdv9_0(.dout(w_dff_A_VQr5k33k2_0),.din(w_dff_A_iu6nTUdv9_0),.clk(gclk));
	jdff dff_A_MxUjFTQs7_0(.dout(w_dff_A_iu6nTUdv9_0),.din(w_dff_A_MxUjFTQs7_0),.clk(gclk));
	jdff dff_A_9clkR7LB8_0(.dout(w_dff_A_MxUjFTQs7_0),.din(w_dff_A_9clkR7LB8_0),.clk(gclk));
	jdff dff_A_Y4yvmXJ00_0(.dout(w_dff_A_9clkR7LB8_0),.din(w_dff_A_Y4yvmXJ00_0),.clk(gclk));
	jdff dff_A_kUkOPeyL7_0(.dout(w_dff_A_Y4yvmXJ00_0),.din(w_dff_A_kUkOPeyL7_0),.clk(gclk));
	jdff dff_A_zxy5Nh8h9_0(.dout(w_dff_A_kUkOPeyL7_0),.din(w_dff_A_zxy5Nh8h9_0),.clk(gclk));
	jdff dff_A_JeFRJKoD5_1(.dout(w_n86_0[1]),.din(w_dff_A_JeFRJKoD5_1),.clk(gclk));
	jdff dff_A_YsSOuQPd4_2(.dout(w_n86_0[2]),.din(w_dff_A_YsSOuQPd4_2),.clk(gclk));
	jdff dff_A_fjyD841N9_0(.dout(w_G1gat_0[0]),.din(w_dff_A_fjyD841N9_0),.clk(gclk));
	jdff dff_A_avJj2ftp0_0(.dout(w_dff_A_fjyD841N9_0),.din(w_dff_A_avJj2ftp0_0),.clk(gclk));
	jdff dff_A_tuYWeo190_0(.dout(w_dff_A_avJj2ftp0_0),.din(w_dff_A_tuYWeo190_0),.clk(gclk));
	jdff dff_A_bYbJAC8d0_0(.dout(w_dff_A_tuYWeo190_0),.din(w_dff_A_bYbJAC8d0_0),.clk(gclk));
	jdff dff_A_UhrEUqlX9_0(.dout(w_dff_A_bYbJAC8d0_0),.din(w_dff_A_UhrEUqlX9_0),.clk(gclk));
	jdff dff_A_ipxFgEKq0_0(.dout(w_dff_A_UhrEUqlX9_0),.din(w_dff_A_ipxFgEKq0_0),.clk(gclk));
	jdff dff_A_bayfh9BD1_0(.dout(w_dff_A_ipxFgEKq0_0),.din(w_dff_A_bayfh9BD1_0),.clk(gclk));
	jdff dff_A_kXsHjL2F7_0(.dout(w_dff_A_bayfh9BD1_0),.din(w_dff_A_kXsHjL2F7_0),.clk(gclk));
	jdff dff_A_gZJUWUz46_0(.dout(w_dff_A_kXsHjL2F7_0),.din(w_dff_A_gZJUWUz46_0),.clk(gclk));
	jdff dff_A_C7ey6viR4_0(.dout(w_dff_A_gZJUWUz46_0),.din(w_dff_A_C7ey6viR4_0),.clk(gclk));
	jdff dff_A_q3IXA9W52_0(.dout(w_dff_A_C7ey6viR4_0),.din(w_dff_A_q3IXA9W52_0),.clk(gclk));
	jdff dff_A_c8M1Daca4_0(.dout(w_G57gat_0[0]),.din(w_dff_A_c8M1Daca4_0),.clk(gclk));
	jdff dff_A_DeYvB5iv4_0(.dout(w_dff_A_c8M1Daca4_0),.din(w_dff_A_DeYvB5iv4_0),.clk(gclk));
	jdff dff_A_8x6vm9N22_0(.dout(w_dff_A_DeYvB5iv4_0),.din(w_dff_A_8x6vm9N22_0),.clk(gclk));
	jdff dff_A_a8nYAgs06_0(.dout(w_dff_A_8x6vm9N22_0),.din(w_dff_A_a8nYAgs06_0),.clk(gclk));
	jdff dff_A_RVttjQKE7_0(.dout(w_dff_A_a8nYAgs06_0),.din(w_dff_A_RVttjQKE7_0),.clk(gclk));
	jdff dff_A_9mHACmty0_0(.dout(w_dff_A_RVttjQKE7_0),.din(w_dff_A_9mHACmty0_0),.clk(gclk));
	jdff dff_A_lrmPbqPV3_0(.dout(w_dff_A_9mHACmty0_0),.din(w_dff_A_lrmPbqPV3_0),.clk(gclk));
	jdff dff_A_9Zndlanj0_0(.dout(w_dff_A_lrmPbqPV3_0),.din(w_dff_A_9Zndlanj0_0),.clk(gclk));
	jdff dff_A_ojE9KtrR0_0(.dout(w_dff_A_9Zndlanj0_0),.din(w_dff_A_ojE9KtrR0_0),.clk(gclk));
	jdff dff_A_HIeUN9hn4_0(.dout(w_dff_A_ojE9KtrR0_0),.din(w_dff_A_HIeUN9hn4_0),.clk(gclk));
	jdff dff_A_9XxXW3xX6_0(.dout(w_dff_A_HIeUN9hn4_0),.din(w_dff_A_9XxXW3xX6_0),.clk(gclk));
	jdff dff_B_FN6x3i5p4_2(.din(n239),.dout(w_dff_B_FN6x3i5p4_2),.clk(gclk));
	jdff dff_B_DZK3WZP06_2(.din(w_dff_B_FN6x3i5p4_2),.dout(w_dff_B_DZK3WZP06_2),.clk(gclk));
	jdff dff_B_mgU9srBl5_2(.din(w_dff_B_DZK3WZP06_2),.dout(w_dff_B_mgU9srBl5_2),.clk(gclk));
	jdff dff_A_5rpBHZ9Y5_0(.dout(w_n184_0[0]),.din(w_dff_A_5rpBHZ9Y5_0),.clk(gclk));
	jdff dff_A_wS3rMX7Z2_0(.dout(w_dff_A_5rpBHZ9Y5_0),.din(w_dff_A_wS3rMX7Z2_0),.clk(gclk));
	jdff dff_A_obZl66Kp2_0(.dout(w_dff_A_wS3rMX7Z2_0),.din(w_dff_A_obZl66Kp2_0),.clk(gclk));
	jdff dff_A_b3ZU5CRD9_0(.dout(w_dff_A_obZl66Kp2_0),.din(w_dff_A_b3ZU5CRD9_0),.clk(gclk));
	jdff dff_A_A5YsYjkw6_0(.dout(w_dff_A_b3ZU5CRD9_0),.din(w_dff_A_A5YsYjkw6_0),.clk(gclk));
	jdff dff_A_6ksQyobo0_2(.dout(w_n184_0[2]),.din(w_dff_A_6ksQyobo0_2),.clk(gclk));
	jdff dff_A_FW6K1mqG8_2(.dout(w_dff_A_6ksQyobo0_2),.din(w_dff_A_FW6K1mqG8_2),.clk(gclk));
	jdff dff_A_fFLvYv756_2(.dout(w_dff_A_FW6K1mqG8_2),.din(w_dff_A_fFLvYv756_2),.clk(gclk));
	jdff dff_A_hNg3QhNa1_2(.dout(w_dff_A_fFLvYv756_2),.din(w_dff_A_hNg3QhNa1_2),.clk(gclk));
	jdff dff_A_GTn9ZlPg9_2(.dout(w_dff_A_hNg3QhNa1_2),.din(w_dff_A_GTn9ZlPg9_2),.clk(gclk));
	jdff dff_A_mOfIDB2G0_1(.dout(w_n149_0[1]),.din(w_dff_A_mOfIDB2G0_1),.clk(gclk));
	jdff dff_A_IBrKcLNG2_0(.dout(w_G148gat_0[0]),.din(w_dff_A_IBrKcLNG2_0),.clk(gclk));
	jdff dff_A_9kJParzG4_0(.dout(w_dff_A_IBrKcLNG2_0),.din(w_dff_A_9kJParzG4_0),.clk(gclk));
	jdff dff_A_v5B8dYbp6_0(.dout(w_dff_A_9kJParzG4_0),.din(w_dff_A_v5B8dYbp6_0),.clk(gclk));
	jdff dff_A_3JJvdBJw4_0(.dout(w_dff_A_v5B8dYbp6_0),.din(w_dff_A_3JJvdBJw4_0),.clk(gclk));
	jdff dff_A_mGkbc5EB5_0(.dout(w_dff_A_3JJvdBJw4_0),.din(w_dff_A_mGkbc5EB5_0),.clk(gclk));
	jdff dff_A_cS1pVD993_0(.dout(w_dff_A_mGkbc5EB5_0),.din(w_dff_A_cS1pVD993_0),.clk(gclk));
	jdff dff_A_a1uA0RCw3_0(.dout(w_dff_A_cS1pVD993_0),.din(w_dff_A_a1uA0RCw3_0),.clk(gclk));
	jdff dff_A_hoHB0SEm3_0(.dout(w_dff_A_a1uA0RCw3_0),.din(w_dff_A_hoHB0SEm3_0),.clk(gclk));
	jdff dff_A_CscjWyJh9_0(.dout(w_dff_A_hoHB0SEm3_0),.din(w_dff_A_CscjWyJh9_0),.clk(gclk));
	jdff dff_A_298x2fhx8_0(.dout(w_dff_A_CscjWyJh9_0),.din(w_dff_A_298x2fhx8_0),.clk(gclk));
	jdff dff_A_QUevK6dp3_0(.dout(w_dff_A_298x2fhx8_0),.din(w_dff_A_QUevK6dp3_0),.clk(gclk));
	jdff dff_A_GrMeMyZF1_0(.dout(w_G141gat_0[0]),.din(w_dff_A_GrMeMyZF1_0),.clk(gclk));
	jdff dff_A_3uUohaPd7_0(.dout(w_dff_A_GrMeMyZF1_0),.din(w_dff_A_3uUohaPd7_0),.clk(gclk));
	jdff dff_A_vPVttXBf1_0(.dout(w_dff_A_3uUohaPd7_0),.din(w_dff_A_vPVttXBf1_0),.clk(gclk));
	jdff dff_A_ZenmOmLK7_0(.dout(w_dff_A_vPVttXBf1_0),.din(w_dff_A_ZenmOmLK7_0),.clk(gclk));
	jdff dff_A_VCQ27pGC2_0(.dout(w_dff_A_ZenmOmLK7_0),.din(w_dff_A_VCQ27pGC2_0),.clk(gclk));
	jdff dff_A_WcmBgBec0_0(.dout(w_dff_A_VCQ27pGC2_0),.din(w_dff_A_WcmBgBec0_0),.clk(gclk));
	jdff dff_A_rxSUfTEa1_0(.dout(w_dff_A_WcmBgBec0_0),.din(w_dff_A_rxSUfTEa1_0),.clk(gclk));
	jdff dff_A_jrftIraZ8_0(.dout(w_dff_A_rxSUfTEa1_0),.din(w_dff_A_jrftIraZ8_0),.clk(gclk));
	jdff dff_A_5zQR7pOJ1_0(.dout(w_dff_A_jrftIraZ8_0),.din(w_dff_A_5zQR7pOJ1_0),.clk(gclk));
	jdff dff_A_IyqTxqZr5_0(.dout(w_dff_A_5zQR7pOJ1_0),.din(w_dff_A_IyqTxqZr5_0),.clk(gclk));
	jdff dff_A_jysE7TwX7_0(.dout(w_dff_A_IyqTxqZr5_0),.din(w_dff_A_jysE7TwX7_0),.clk(gclk));
	jdff dff_A_Wjup1IRw4_0(.dout(w_G155gat_0[0]),.din(w_dff_A_Wjup1IRw4_0),.clk(gclk));
	jdff dff_A_LXkA0udj3_0(.dout(w_dff_A_Wjup1IRw4_0),.din(w_dff_A_LXkA0udj3_0),.clk(gclk));
	jdff dff_A_sNOjqHPW9_0(.dout(w_dff_A_LXkA0udj3_0),.din(w_dff_A_sNOjqHPW9_0),.clk(gclk));
	jdff dff_A_HH4SlpT82_0(.dout(w_dff_A_sNOjqHPW9_0),.din(w_dff_A_HH4SlpT82_0),.clk(gclk));
	jdff dff_A_2TxDSsYj0_0(.dout(w_dff_A_HH4SlpT82_0),.din(w_dff_A_2TxDSsYj0_0),.clk(gclk));
	jdff dff_A_AoQqhtKp4_0(.dout(w_dff_A_2TxDSsYj0_0),.din(w_dff_A_AoQqhtKp4_0),.clk(gclk));
	jdff dff_A_hvEi9KZs8_0(.dout(w_dff_A_AoQqhtKp4_0),.din(w_dff_A_hvEi9KZs8_0),.clk(gclk));
	jdff dff_A_Ws3QqX2U4_0(.dout(w_dff_A_hvEi9KZs8_0),.din(w_dff_A_Ws3QqX2U4_0),.clk(gclk));
	jdff dff_A_CSyVbtZr0_0(.dout(w_dff_A_Ws3QqX2U4_0),.din(w_dff_A_CSyVbtZr0_0),.clk(gclk));
	jdff dff_A_60vNMrCt1_0(.dout(w_dff_A_CSyVbtZr0_0),.din(w_dff_A_60vNMrCt1_0),.clk(gclk));
	jdff dff_A_ngdY3SaI8_0(.dout(w_dff_A_60vNMrCt1_0),.din(w_dff_A_ngdY3SaI8_0),.clk(gclk));
	jdff dff_A_dUlmOZCS9_0(.dout(w_G22gat_0[0]),.din(w_dff_A_dUlmOZCS9_0),.clk(gclk));
	jdff dff_A_t88rpmNf5_0(.dout(w_dff_A_dUlmOZCS9_0),.din(w_dff_A_t88rpmNf5_0),.clk(gclk));
	jdff dff_A_05NRixIk1_0(.dout(w_dff_A_t88rpmNf5_0),.din(w_dff_A_05NRixIk1_0),.clk(gclk));
	jdff dff_A_qFwhbF090_0(.dout(w_dff_A_05NRixIk1_0),.din(w_dff_A_qFwhbF090_0),.clk(gclk));
	jdff dff_A_62pxMxPT3_0(.dout(w_dff_A_qFwhbF090_0),.din(w_dff_A_62pxMxPT3_0),.clk(gclk));
	jdff dff_A_gIvEyhlY3_0(.dout(w_dff_A_62pxMxPT3_0),.din(w_dff_A_gIvEyhlY3_0),.clk(gclk));
	jdff dff_A_IrNsnhhT7_0(.dout(w_dff_A_gIvEyhlY3_0),.din(w_dff_A_IrNsnhhT7_0),.clk(gclk));
	jdff dff_A_BsFFiPo78_0(.dout(w_dff_A_IrNsnhhT7_0),.din(w_dff_A_BsFFiPo78_0),.clk(gclk));
	jdff dff_A_VtflH0ef6_0(.dout(w_dff_A_BsFFiPo78_0),.din(w_dff_A_VtflH0ef6_0),.clk(gclk));
	jdff dff_A_kLAoUdji0_0(.dout(w_dff_A_VtflH0ef6_0),.din(w_dff_A_kLAoUdji0_0),.clk(gclk));
	jdff dff_A_9QQ3fZkz9_0(.dout(w_dff_A_kLAoUdji0_0),.din(w_dff_A_9QQ3fZkz9_0),.clk(gclk));
	jdff dff_A_F1ag4jyI7_0(.dout(w_G78gat_0[0]),.din(w_dff_A_F1ag4jyI7_0),.clk(gclk));
	jdff dff_A_7Ad9wT1O1_0(.dout(w_dff_A_F1ag4jyI7_0),.din(w_dff_A_7Ad9wT1O1_0),.clk(gclk));
	jdff dff_A_6zZSLCky6_0(.dout(w_dff_A_7Ad9wT1O1_0),.din(w_dff_A_6zZSLCky6_0),.clk(gclk));
	jdff dff_A_WS9y7ycB1_0(.dout(w_dff_A_6zZSLCky6_0),.din(w_dff_A_WS9y7ycB1_0),.clk(gclk));
	jdff dff_A_dTzzst487_0(.dout(w_dff_A_WS9y7ycB1_0),.din(w_dff_A_dTzzst487_0),.clk(gclk));
	jdff dff_A_w5eDU67r2_0(.dout(w_dff_A_dTzzst487_0),.din(w_dff_A_w5eDU67r2_0),.clk(gclk));
	jdff dff_A_7gg6dw5F5_0(.dout(w_dff_A_w5eDU67r2_0),.din(w_dff_A_7gg6dw5F5_0),.clk(gclk));
	jdff dff_A_TTbcbWoG6_0(.dout(w_dff_A_7gg6dw5F5_0),.din(w_dff_A_TTbcbWoG6_0),.clk(gclk));
	jdff dff_A_6dhh8FJW0_0(.dout(w_dff_A_TTbcbWoG6_0),.din(w_dff_A_6dhh8FJW0_0),.clk(gclk));
	jdff dff_A_v4rVVFR89_0(.dout(w_dff_A_6dhh8FJW0_0),.din(w_dff_A_v4rVVFR89_0),.clk(gclk));
	jdff dff_A_BwzKoTGC1_0(.dout(w_dff_A_v4rVVFR89_0),.din(w_dff_A_BwzKoTGC1_0),.clk(gclk));
	jdff dff_A_ltmQRJef6_0(.dout(w_G204gat_0[0]),.din(w_dff_A_ltmQRJef6_0),.clk(gclk));
	jdff dff_A_2wmY0NjK8_0(.dout(w_dff_A_ltmQRJef6_0),.din(w_dff_A_2wmY0NjK8_0),.clk(gclk));
	jdff dff_A_jWcYPu8D1_0(.dout(w_dff_A_2wmY0NjK8_0),.din(w_dff_A_jWcYPu8D1_0),.clk(gclk));
	jdff dff_A_WbFxjA5x8_0(.dout(w_dff_A_jWcYPu8D1_0),.din(w_dff_A_WbFxjA5x8_0),.clk(gclk));
	jdff dff_A_aOxQvsnk3_0(.dout(w_dff_A_WbFxjA5x8_0),.din(w_dff_A_aOxQvsnk3_0),.clk(gclk));
	jdff dff_A_VnaQW3wC7_0(.dout(w_dff_A_aOxQvsnk3_0),.din(w_dff_A_VnaQW3wC7_0),.clk(gclk));
	jdff dff_A_msJfL2z22_0(.dout(w_dff_A_VnaQW3wC7_0),.din(w_dff_A_msJfL2z22_0),.clk(gclk));
	jdff dff_A_syAWKpDS8_0(.dout(w_dff_A_msJfL2z22_0),.din(w_dff_A_syAWKpDS8_0),.clk(gclk));
	jdff dff_A_F9ivLoom3_0(.dout(w_dff_A_syAWKpDS8_0),.din(w_dff_A_F9ivLoom3_0),.clk(gclk));
	jdff dff_A_AYXiWdPm5_0(.dout(w_dff_A_F9ivLoom3_0),.din(w_dff_A_AYXiWdPm5_0),.clk(gclk));
	jdff dff_A_KrOmtTGV2_0(.dout(w_dff_A_AYXiWdPm5_0),.din(w_dff_A_KrOmtTGV2_0),.clk(gclk));
	jdff dff_A_b39vc3QZ9_0(.dout(w_G197gat_0[0]),.din(w_dff_A_b39vc3QZ9_0),.clk(gclk));
	jdff dff_A_J9bzhHzr3_0(.dout(w_dff_A_b39vc3QZ9_0),.din(w_dff_A_J9bzhHzr3_0),.clk(gclk));
	jdff dff_A_mBQ4E0OV7_0(.dout(w_dff_A_J9bzhHzr3_0),.din(w_dff_A_mBQ4E0OV7_0),.clk(gclk));
	jdff dff_A_BhhvN9zP2_0(.dout(w_dff_A_mBQ4E0OV7_0),.din(w_dff_A_BhhvN9zP2_0),.clk(gclk));
	jdff dff_A_zNvTAT2H4_0(.dout(w_dff_A_BhhvN9zP2_0),.din(w_dff_A_zNvTAT2H4_0),.clk(gclk));
	jdff dff_A_XYOFRBsW9_0(.dout(w_dff_A_zNvTAT2H4_0),.din(w_dff_A_XYOFRBsW9_0),.clk(gclk));
	jdff dff_A_u0Vo8dHc9_0(.dout(w_dff_A_XYOFRBsW9_0),.din(w_dff_A_u0Vo8dHc9_0),.clk(gclk));
	jdff dff_A_8sJHAHMa8_0(.dout(w_dff_A_u0Vo8dHc9_0),.din(w_dff_A_8sJHAHMa8_0),.clk(gclk));
	jdff dff_A_YvDo8HyO0_0(.dout(w_dff_A_8sJHAHMa8_0),.din(w_dff_A_YvDo8HyO0_0),.clk(gclk));
	jdff dff_A_fOyPEcy97_0(.dout(w_dff_A_YvDo8HyO0_0),.din(w_dff_A_fOyPEcy97_0),.clk(gclk));
	jdff dff_A_Gwy7oFm21_0(.dout(w_dff_A_fOyPEcy97_0),.din(w_dff_A_Gwy7oFm21_0),.clk(gclk));
	jdff dff_A_9hFN8fiq0_0(.dout(w_G211gat_0[0]),.din(w_dff_A_9hFN8fiq0_0),.clk(gclk));
	jdff dff_A_29a9GGBp5_0(.dout(w_dff_A_9hFN8fiq0_0),.din(w_dff_A_29a9GGBp5_0),.clk(gclk));
	jdff dff_A_sLB8Djhu8_0(.dout(w_dff_A_29a9GGBp5_0),.din(w_dff_A_sLB8Djhu8_0),.clk(gclk));
	jdff dff_A_b0BNUmcL6_0(.dout(w_dff_A_sLB8Djhu8_0),.din(w_dff_A_b0BNUmcL6_0),.clk(gclk));
	jdff dff_A_ZBxHxwk98_0(.dout(w_dff_A_b0BNUmcL6_0),.din(w_dff_A_ZBxHxwk98_0),.clk(gclk));
	jdff dff_A_SOqBOHeV2_0(.dout(w_dff_A_ZBxHxwk98_0),.din(w_dff_A_SOqBOHeV2_0),.clk(gclk));
	jdff dff_A_9peYCn8v9_0(.dout(w_dff_A_SOqBOHeV2_0),.din(w_dff_A_9peYCn8v9_0),.clk(gclk));
	jdff dff_A_eUmG3bzi4_0(.dout(w_dff_A_9peYCn8v9_0),.din(w_dff_A_eUmG3bzi4_0),.clk(gclk));
	jdff dff_A_nDGzSmq67_0(.dout(w_dff_A_eUmG3bzi4_0),.din(w_dff_A_nDGzSmq67_0),.clk(gclk));
	jdff dff_A_Z2bMR47X9_0(.dout(w_dff_A_nDGzSmq67_0),.din(w_dff_A_Z2bMR47X9_0),.clk(gclk));
	jdff dff_A_lMiBnJV77_0(.dout(w_dff_A_Z2bMR47X9_0),.din(w_dff_A_lMiBnJV77_0),.clk(gclk));
	jdff dff_A_ijYXtsu43_1(.dout(w_n141_0[1]),.din(w_dff_A_ijYXtsu43_1),.clk(gclk));
	jdff dff_A_Lb6kz2pA7_0(.dout(w_G120gat_0[0]),.din(w_dff_A_Lb6kz2pA7_0),.clk(gclk));
	jdff dff_A_sbVzrm911_0(.dout(w_dff_A_Lb6kz2pA7_0),.din(w_dff_A_sbVzrm911_0),.clk(gclk));
	jdff dff_A_NEf6hx670_0(.dout(w_dff_A_sbVzrm911_0),.din(w_dff_A_NEf6hx670_0),.clk(gclk));
	jdff dff_A_zN7s2WAX1_0(.dout(w_dff_A_NEf6hx670_0),.din(w_dff_A_zN7s2WAX1_0),.clk(gclk));
	jdff dff_A_EcDuipzG7_0(.dout(w_dff_A_zN7s2WAX1_0),.din(w_dff_A_EcDuipzG7_0),.clk(gclk));
	jdff dff_A_BIttUVuv5_0(.dout(w_dff_A_EcDuipzG7_0),.din(w_dff_A_BIttUVuv5_0),.clk(gclk));
	jdff dff_A_HE2q2hQk9_0(.dout(w_dff_A_BIttUVuv5_0),.din(w_dff_A_HE2q2hQk9_0),.clk(gclk));
	jdff dff_A_l4ZNmGCZ2_0(.dout(w_dff_A_HE2q2hQk9_0),.din(w_dff_A_l4ZNmGCZ2_0),.clk(gclk));
	jdff dff_A_pBytW4Ve6_0(.dout(w_dff_A_l4ZNmGCZ2_0),.din(w_dff_A_pBytW4Ve6_0),.clk(gclk));
	jdff dff_A_EIa4wKO89_0(.dout(w_dff_A_pBytW4Ve6_0),.din(w_dff_A_EIa4wKO89_0),.clk(gclk));
	jdff dff_A_ZuYfv5UA5_0(.dout(w_dff_A_EIa4wKO89_0),.din(w_dff_A_ZuYfv5UA5_0),.clk(gclk));
	jdff dff_A_isSYifqF7_0(.dout(w_G113gat_0[0]),.din(w_dff_A_isSYifqF7_0),.clk(gclk));
	jdff dff_A_RUmCfxN44_0(.dout(w_dff_A_isSYifqF7_0),.din(w_dff_A_RUmCfxN44_0),.clk(gclk));
	jdff dff_A_wWNqEg6X7_0(.dout(w_dff_A_RUmCfxN44_0),.din(w_dff_A_wWNqEg6X7_0),.clk(gclk));
	jdff dff_A_Pp61Fpnw7_0(.dout(w_dff_A_wWNqEg6X7_0),.din(w_dff_A_Pp61Fpnw7_0),.clk(gclk));
	jdff dff_A_pTWFA8Of1_0(.dout(w_dff_A_Pp61Fpnw7_0),.din(w_dff_A_pTWFA8Of1_0),.clk(gclk));
	jdff dff_A_FzCodUre2_0(.dout(w_dff_A_pTWFA8Of1_0),.din(w_dff_A_FzCodUre2_0),.clk(gclk));
	jdff dff_A_ooi2NbM65_0(.dout(w_dff_A_FzCodUre2_0),.din(w_dff_A_ooi2NbM65_0),.clk(gclk));
	jdff dff_A_CjkmQe6O8_0(.dout(w_dff_A_ooi2NbM65_0),.din(w_dff_A_CjkmQe6O8_0),.clk(gclk));
	jdff dff_A_pNXEIKWR9_0(.dout(w_dff_A_CjkmQe6O8_0),.din(w_dff_A_pNXEIKWR9_0),.clk(gclk));
	jdff dff_A_aR24SEHt8_0(.dout(w_dff_A_pNXEIKWR9_0),.din(w_dff_A_aR24SEHt8_0),.clk(gclk));
	jdff dff_A_uiifWNTX9_0(.dout(w_dff_A_aR24SEHt8_0),.din(w_dff_A_uiifWNTX9_0),.clk(gclk));
	jdff dff_A_IlsdWfLE1_0(.dout(w_G127gat_0[0]),.din(w_dff_A_IlsdWfLE1_0),.clk(gclk));
	jdff dff_A_WLrUWIod0_0(.dout(w_dff_A_IlsdWfLE1_0),.din(w_dff_A_WLrUWIod0_0),.clk(gclk));
	jdff dff_A_F99SQd835_0(.dout(w_dff_A_WLrUWIod0_0),.din(w_dff_A_F99SQd835_0),.clk(gclk));
	jdff dff_A_b3MpnxRj6_0(.dout(w_dff_A_F99SQd835_0),.din(w_dff_A_b3MpnxRj6_0),.clk(gclk));
	jdff dff_A_AzpbqCB43_0(.dout(w_dff_A_b3MpnxRj6_0),.din(w_dff_A_AzpbqCB43_0),.clk(gclk));
	jdff dff_A_9XpmKFk98_0(.dout(w_dff_A_AzpbqCB43_0),.din(w_dff_A_9XpmKFk98_0),.clk(gclk));
	jdff dff_A_FASDJSlH3_0(.dout(w_dff_A_9XpmKFk98_0),.din(w_dff_A_FASDJSlH3_0),.clk(gclk));
	jdff dff_A_jgB2nQ7x2_0(.dout(w_dff_A_FASDJSlH3_0),.din(w_dff_A_jgB2nQ7x2_0),.clk(gclk));
	jdff dff_A_4Wki2hco9_0(.dout(w_dff_A_jgB2nQ7x2_0),.din(w_dff_A_4Wki2hco9_0),.clk(gclk));
	jdff dff_A_ZXMVv5bR9_0(.dout(w_dff_A_4Wki2hco9_0),.din(w_dff_A_ZXMVv5bR9_0),.clk(gclk));
	jdff dff_A_k98m0A6N9_0(.dout(w_dff_A_ZXMVv5bR9_0),.din(w_dff_A_k98m0A6N9_0),.clk(gclk));
	jdff dff_A_ZNghoZoP8_0(.dout(w_G15gat_0[0]),.din(w_dff_A_ZNghoZoP8_0),.clk(gclk));
	jdff dff_A_bDis0Ej32_0(.dout(w_dff_A_ZNghoZoP8_0),.din(w_dff_A_bDis0Ej32_0),.clk(gclk));
	jdff dff_A_nfbbIKTc1_0(.dout(w_dff_A_bDis0Ej32_0),.din(w_dff_A_nfbbIKTc1_0),.clk(gclk));
	jdff dff_A_hC9ErcYS1_0(.dout(w_dff_A_nfbbIKTc1_0),.din(w_dff_A_hC9ErcYS1_0),.clk(gclk));
	jdff dff_A_hcP8IOIL7_0(.dout(w_dff_A_hC9ErcYS1_0),.din(w_dff_A_hcP8IOIL7_0),.clk(gclk));
	jdff dff_A_N4nYGrpn9_0(.dout(w_dff_A_hcP8IOIL7_0),.din(w_dff_A_N4nYGrpn9_0),.clk(gclk));
	jdff dff_A_iWCToGTf4_0(.dout(w_dff_A_N4nYGrpn9_0),.din(w_dff_A_iWCToGTf4_0),.clk(gclk));
	jdff dff_A_OKp1P4BM3_0(.dout(w_dff_A_iWCToGTf4_0),.din(w_dff_A_OKp1P4BM3_0),.clk(gclk));
	jdff dff_A_44dvDDGH3_0(.dout(w_dff_A_OKp1P4BM3_0),.din(w_dff_A_44dvDDGH3_0),.clk(gclk));
	jdff dff_A_1A3pKgdw0_0(.dout(w_dff_A_44dvDDGH3_0),.din(w_dff_A_1A3pKgdw0_0),.clk(gclk));
	jdff dff_A_9Zmys9zm8_0(.dout(w_dff_A_1A3pKgdw0_0),.din(w_dff_A_9Zmys9zm8_0),.clk(gclk));
	jdff dff_A_F5f0KTTL2_0(.dout(w_G71gat_0[0]),.din(w_dff_A_F5f0KTTL2_0),.clk(gclk));
	jdff dff_A_1zeN642C6_0(.dout(w_dff_A_F5f0KTTL2_0),.din(w_dff_A_1zeN642C6_0),.clk(gclk));
	jdff dff_A_tVwf1G7g4_0(.dout(w_dff_A_1zeN642C6_0),.din(w_dff_A_tVwf1G7g4_0),.clk(gclk));
	jdff dff_A_amEVcshH5_0(.dout(w_dff_A_tVwf1G7g4_0),.din(w_dff_A_amEVcshH5_0),.clk(gclk));
	jdff dff_A_6q4EgFg07_0(.dout(w_dff_A_amEVcshH5_0),.din(w_dff_A_6q4EgFg07_0),.clk(gclk));
	jdff dff_A_P024Q8QK2_0(.dout(w_dff_A_6q4EgFg07_0),.din(w_dff_A_P024Q8QK2_0),.clk(gclk));
	jdff dff_A_jWQzdFGG2_0(.dout(w_dff_A_P024Q8QK2_0),.din(w_dff_A_jWQzdFGG2_0),.clk(gclk));
	jdff dff_A_iIdzb1Zl8_0(.dout(w_dff_A_jWQzdFGG2_0),.din(w_dff_A_iIdzb1Zl8_0),.clk(gclk));
	jdff dff_A_GBzglkQJ2_0(.dout(w_dff_A_iIdzb1Zl8_0),.din(w_dff_A_GBzglkQJ2_0),.clk(gclk));
	jdff dff_A_bFixfnyz9_0(.dout(w_dff_A_GBzglkQJ2_0),.din(w_dff_A_bFixfnyz9_0),.clk(gclk));
	jdff dff_A_wNbvbPej9_0(.dout(w_dff_A_bFixfnyz9_0),.din(w_dff_A_wNbvbPej9_0),.clk(gclk));
	jdff dff_A_FkeL3ixr3_0(.dout(w_G176gat_0[0]),.din(w_dff_A_FkeL3ixr3_0),.clk(gclk));
	jdff dff_A_md2Y4LjD5_0(.dout(w_dff_A_FkeL3ixr3_0),.din(w_dff_A_md2Y4LjD5_0),.clk(gclk));
	jdff dff_A_YRE9P2K52_0(.dout(w_dff_A_md2Y4LjD5_0),.din(w_dff_A_YRE9P2K52_0),.clk(gclk));
	jdff dff_A_dLDKf2tP4_0(.dout(w_dff_A_YRE9P2K52_0),.din(w_dff_A_dLDKf2tP4_0),.clk(gclk));
	jdff dff_A_btBz3Pw79_0(.dout(w_dff_A_dLDKf2tP4_0),.din(w_dff_A_btBz3Pw79_0),.clk(gclk));
	jdff dff_A_L7Opz9Ul2_0(.dout(w_dff_A_btBz3Pw79_0),.din(w_dff_A_L7Opz9Ul2_0),.clk(gclk));
	jdff dff_A_rQeAf3kD2_0(.dout(w_dff_A_L7Opz9Ul2_0),.din(w_dff_A_rQeAf3kD2_0),.clk(gclk));
	jdff dff_A_D6sWsJ3m5_0(.dout(w_dff_A_rQeAf3kD2_0),.din(w_dff_A_D6sWsJ3m5_0),.clk(gclk));
	jdff dff_A_OpM7NSH44_0(.dout(w_dff_A_D6sWsJ3m5_0),.din(w_dff_A_OpM7NSH44_0),.clk(gclk));
	jdff dff_A_b7D4FyFS5_0(.dout(w_dff_A_OpM7NSH44_0),.din(w_dff_A_b7D4FyFS5_0),.clk(gclk));
	jdff dff_A_DXT6JGjF6_0(.dout(w_dff_A_b7D4FyFS5_0),.din(w_dff_A_DXT6JGjF6_0),.clk(gclk));
	jdff dff_A_TZkhoD105_0(.dout(w_G169gat_0[0]),.din(w_dff_A_TZkhoD105_0),.clk(gclk));
	jdff dff_A_nnUOQRxn3_0(.dout(w_dff_A_TZkhoD105_0),.din(w_dff_A_nnUOQRxn3_0),.clk(gclk));
	jdff dff_A_uEx2BNFk1_0(.dout(w_dff_A_nnUOQRxn3_0),.din(w_dff_A_uEx2BNFk1_0),.clk(gclk));
	jdff dff_A_ojGlo7Fo9_0(.dout(w_dff_A_uEx2BNFk1_0),.din(w_dff_A_ojGlo7Fo9_0),.clk(gclk));
	jdff dff_A_fMUtyY8P0_0(.dout(w_dff_A_ojGlo7Fo9_0),.din(w_dff_A_fMUtyY8P0_0),.clk(gclk));
	jdff dff_A_DF38NtLE4_0(.dout(w_dff_A_fMUtyY8P0_0),.din(w_dff_A_DF38NtLE4_0),.clk(gclk));
	jdff dff_A_Fycx3Eoy4_0(.dout(w_dff_A_DF38NtLE4_0),.din(w_dff_A_Fycx3Eoy4_0),.clk(gclk));
	jdff dff_A_cMorxdi31_0(.dout(w_dff_A_Fycx3Eoy4_0),.din(w_dff_A_cMorxdi31_0),.clk(gclk));
	jdff dff_A_HMzP6F4k3_0(.dout(w_dff_A_cMorxdi31_0),.din(w_dff_A_HMzP6F4k3_0),.clk(gclk));
	jdff dff_A_eCzi1cYe3_0(.dout(w_dff_A_HMzP6F4k3_0),.din(w_dff_A_eCzi1cYe3_0),.clk(gclk));
	jdff dff_A_FKRrwreq2_0(.dout(w_dff_A_eCzi1cYe3_0),.din(w_dff_A_FKRrwreq2_0),.clk(gclk));
	jdff dff_A_XLv82hXB4_0(.dout(w_G183gat_0[0]),.din(w_dff_A_XLv82hXB4_0),.clk(gclk));
	jdff dff_A_tfMOTZAD1_0(.dout(w_dff_A_XLv82hXB4_0),.din(w_dff_A_tfMOTZAD1_0),.clk(gclk));
	jdff dff_A_L4eZFemM2_0(.dout(w_dff_A_tfMOTZAD1_0),.din(w_dff_A_L4eZFemM2_0),.clk(gclk));
	jdff dff_A_mzaJ5xL68_0(.dout(w_dff_A_L4eZFemM2_0),.din(w_dff_A_mzaJ5xL68_0),.clk(gclk));
	jdff dff_A_rLx6zcib2_0(.dout(w_dff_A_mzaJ5xL68_0),.din(w_dff_A_rLx6zcib2_0),.clk(gclk));
	jdff dff_A_bS4eyqfj1_0(.dout(w_dff_A_rLx6zcib2_0),.din(w_dff_A_bS4eyqfj1_0),.clk(gclk));
	jdff dff_A_6htZAKQQ3_0(.dout(w_dff_A_bS4eyqfj1_0),.din(w_dff_A_6htZAKQQ3_0),.clk(gclk));
	jdff dff_A_jzfnpbd26_0(.dout(w_dff_A_6htZAKQQ3_0),.din(w_dff_A_jzfnpbd26_0),.clk(gclk));
	jdff dff_A_rLBsRemY7_0(.dout(w_dff_A_jzfnpbd26_0),.din(w_dff_A_rLBsRemY7_0),.clk(gclk));
	jdff dff_A_adApjwo32_0(.dout(w_dff_A_rLBsRemY7_0),.din(w_dff_A_adApjwo32_0),.clk(gclk));
	jdff dff_A_l7QUQJ4y2_0(.dout(w_dff_A_adApjwo32_0),.din(w_dff_A_l7QUQJ4y2_0),.clk(gclk));
	jdff dff_A_wu2Fi6xf5_1(.dout(w_n187_0[1]),.din(w_dff_A_wu2Fi6xf5_1),.clk(gclk));
	jdff dff_A_QHtTSUqp2_1(.dout(w_dff_A_wu2Fi6xf5_1),.din(w_dff_A_QHtTSUqp2_1),.clk(gclk));
	jdff dff_A_UhfF8zm33_1(.dout(w_dff_A_QHtTSUqp2_1),.din(w_dff_A_UhfF8zm33_1),.clk(gclk));
	jdff dff_A_vlAdmt1s4_1(.dout(w_dff_A_UhfF8zm33_1),.din(w_dff_A_vlAdmt1s4_1),.clk(gclk));
	jdff dff_A_4G4z2rLk7_1(.dout(w_dff_A_vlAdmt1s4_1),.din(w_dff_A_4G4z2rLk7_1),.clk(gclk));
	jdff dff_A_3fJI5Gln5_2(.dout(w_n187_0[2]),.din(w_dff_A_3fJI5Gln5_2),.clk(gclk));
	jdff dff_A_P3ilw5YH3_2(.dout(w_dff_A_3fJI5Gln5_2),.din(w_dff_A_P3ilw5YH3_2),.clk(gclk));
	jdff dff_A_JpauP8u43_2(.dout(w_dff_A_P3ilw5YH3_2),.din(w_dff_A_JpauP8u43_2),.clk(gclk));
	jdff dff_A_MO0shkh64_2(.dout(w_dff_A_JpauP8u43_2),.din(w_dff_A_MO0shkh64_2),.clk(gclk));
	jdff dff_A_TWxn2FOh5_2(.dout(w_dff_A_MO0shkh64_2),.din(w_dff_A_TWxn2FOh5_2),.clk(gclk));
	jdff dff_A_ObRYbEa95_1(.dout(w_n102_1[1]),.din(w_dff_A_ObRYbEa95_1),.clk(gclk));
	jdff dff_A_eeBMqcSL9_0(.dout(w_G36gat_0[0]),.din(w_dff_A_eeBMqcSL9_0),.clk(gclk));
	jdff dff_A_81y54dIb4_0(.dout(w_dff_A_eeBMqcSL9_0),.din(w_dff_A_81y54dIb4_0),.clk(gclk));
	jdff dff_A_99p2sCA35_0(.dout(w_dff_A_81y54dIb4_0),.din(w_dff_A_99p2sCA35_0),.clk(gclk));
	jdff dff_A_vuXmwXtk2_0(.dout(w_dff_A_99p2sCA35_0),.din(w_dff_A_vuXmwXtk2_0),.clk(gclk));
	jdff dff_A_zU1yKGA75_0(.dout(w_dff_A_vuXmwXtk2_0),.din(w_dff_A_zU1yKGA75_0),.clk(gclk));
	jdff dff_A_nN6CIYEv6_0(.dout(w_dff_A_zU1yKGA75_0),.din(w_dff_A_nN6CIYEv6_0),.clk(gclk));
	jdff dff_A_zupqc8xA8_0(.dout(w_dff_A_nN6CIYEv6_0),.din(w_dff_A_zupqc8xA8_0),.clk(gclk));
	jdff dff_A_R6QXTkRz7_0(.dout(w_dff_A_zupqc8xA8_0),.din(w_dff_A_R6QXTkRz7_0),.clk(gclk));
	jdff dff_A_AcC6QKlA7_0(.dout(w_dff_A_R6QXTkRz7_0),.din(w_dff_A_AcC6QKlA7_0),.clk(gclk));
	jdff dff_A_Aw6xG1tM9_0(.dout(w_dff_A_AcC6QKlA7_0),.din(w_dff_A_Aw6xG1tM9_0),.clk(gclk));
	jdff dff_A_M9pBSjVC9_0(.dout(w_dff_A_Aw6xG1tM9_0),.din(w_dff_A_M9pBSjVC9_0),.clk(gclk));
	jdff dff_A_NEQrfpyP2_0(.dout(w_G29gat_0[0]),.din(w_dff_A_NEQrfpyP2_0),.clk(gclk));
	jdff dff_A_dNzug4h47_0(.dout(w_dff_A_NEQrfpyP2_0),.din(w_dff_A_dNzug4h47_0),.clk(gclk));
	jdff dff_A_JbObE0ED8_0(.dout(w_dff_A_dNzug4h47_0),.din(w_dff_A_JbObE0ED8_0),.clk(gclk));
	jdff dff_A_4ePAcUgm1_0(.dout(w_dff_A_JbObE0ED8_0),.din(w_dff_A_4ePAcUgm1_0),.clk(gclk));
	jdff dff_A_Z2FUtYC02_0(.dout(w_dff_A_4ePAcUgm1_0),.din(w_dff_A_Z2FUtYC02_0),.clk(gclk));
	jdff dff_A_k1syVgTO2_0(.dout(w_dff_A_Z2FUtYC02_0),.din(w_dff_A_k1syVgTO2_0),.clk(gclk));
	jdff dff_A_gxRxyFBv0_0(.dout(w_dff_A_k1syVgTO2_0),.din(w_dff_A_gxRxyFBv0_0),.clk(gclk));
	jdff dff_A_XtD5lwcV3_0(.dout(w_dff_A_gxRxyFBv0_0),.din(w_dff_A_XtD5lwcV3_0),.clk(gclk));
	jdff dff_A_UBMdbGhA9_0(.dout(w_dff_A_XtD5lwcV3_0),.din(w_dff_A_UBMdbGhA9_0),.clk(gclk));
	jdff dff_A_zPTZq0wv6_0(.dout(w_dff_A_UBMdbGhA9_0),.din(w_dff_A_zPTZq0wv6_0),.clk(gclk));
	jdff dff_A_i5GnN5Yd6_0(.dout(w_dff_A_zPTZq0wv6_0),.din(w_dff_A_i5GnN5Yd6_0),.clk(gclk));
	jdff dff_A_ZHwhbieb2_0(.dout(w_G50gat_0[0]),.din(w_dff_A_ZHwhbieb2_0),.clk(gclk));
	jdff dff_A_mBUG7djK3_0(.dout(w_dff_A_ZHwhbieb2_0),.din(w_dff_A_mBUG7djK3_0),.clk(gclk));
	jdff dff_A_a8TreNbt2_0(.dout(w_dff_A_mBUG7djK3_0),.din(w_dff_A_a8TreNbt2_0),.clk(gclk));
	jdff dff_A_cNds3O5H4_0(.dout(w_dff_A_a8TreNbt2_0),.din(w_dff_A_cNds3O5H4_0),.clk(gclk));
	jdff dff_A_WSi4d5NM0_0(.dout(w_dff_A_cNds3O5H4_0),.din(w_dff_A_WSi4d5NM0_0),.clk(gclk));
	jdff dff_A_FMY34EcV9_0(.dout(w_dff_A_WSi4d5NM0_0),.din(w_dff_A_FMY34EcV9_0),.clk(gclk));
	jdff dff_A_UOYNfn8m1_0(.dout(w_dff_A_FMY34EcV9_0),.din(w_dff_A_UOYNfn8m1_0),.clk(gclk));
	jdff dff_A_da63xLHh9_0(.dout(w_dff_A_UOYNfn8m1_0),.din(w_dff_A_da63xLHh9_0),.clk(gclk));
	jdff dff_A_IMc9dQrW2_0(.dout(w_dff_A_da63xLHh9_0),.din(w_dff_A_IMc9dQrW2_0),.clk(gclk));
	jdff dff_A_5WiMBiUZ1_0(.dout(w_dff_A_IMc9dQrW2_0),.din(w_dff_A_5WiMBiUZ1_0),.clk(gclk));
	jdff dff_A_horf3TtB3_0(.dout(w_dff_A_5WiMBiUZ1_0),.din(w_dff_A_horf3TtB3_0),.clk(gclk));
	jdff dff_A_O07U9qP48_0(.dout(w_G43gat_0[0]),.din(w_dff_A_O07U9qP48_0),.clk(gclk));
	jdff dff_A_dDPdfrUH9_0(.dout(w_dff_A_O07U9qP48_0),.din(w_dff_A_dDPdfrUH9_0),.clk(gclk));
	jdff dff_A_SxLffwx60_0(.dout(w_dff_A_dDPdfrUH9_0),.din(w_dff_A_SxLffwx60_0),.clk(gclk));
	jdff dff_A_7AGBAL0J9_0(.dout(w_dff_A_SxLffwx60_0),.din(w_dff_A_7AGBAL0J9_0),.clk(gclk));
	jdff dff_A_gZc4VdEM7_0(.dout(w_dff_A_7AGBAL0J9_0),.din(w_dff_A_gZc4VdEM7_0),.clk(gclk));
	jdff dff_A_28NRwmeY6_0(.dout(w_dff_A_gZc4VdEM7_0),.din(w_dff_A_28NRwmeY6_0),.clk(gclk));
	jdff dff_A_9kuC86Nm8_0(.dout(w_dff_A_28NRwmeY6_0),.din(w_dff_A_9kuC86Nm8_0),.clk(gclk));
	jdff dff_A_ER1xiWRB0_0(.dout(w_dff_A_9kuC86Nm8_0),.din(w_dff_A_ER1xiWRB0_0),.clk(gclk));
	jdff dff_A_j0gRPcQX1_0(.dout(w_dff_A_ER1xiWRB0_0),.din(w_dff_A_j0gRPcQX1_0),.clk(gclk));
	jdff dff_A_OomMhRsY9_0(.dout(w_dff_A_j0gRPcQX1_0),.din(w_dff_A_OomMhRsY9_0),.clk(gclk));
	jdff dff_A_iqz6IBc73_0(.dout(w_dff_A_OomMhRsY9_0),.din(w_dff_A_iqz6IBc73_0),.clk(gclk));
	jdff dff_A_fKZ0sX0M6_0(.dout(w_G92gat_0[0]),.din(w_dff_A_fKZ0sX0M6_0),.clk(gclk));
	jdff dff_A_l9dYyST45_0(.dout(w_dff_A_fKZ0sX0M6_0),.din(w_dff_A_l9dYyST45_0),.clk(gclk));
	jdff dff_A_zjdxJQMp2_0(.dout(w_dff_A_l9dYyST45_0),.din(w_dff_A_zjdxJQMp2_0),.clk(gclk));
	jdff dff_A_1PUk7Ety7_0(.dout(w_dff_A_zjdxJQMp2_0),.din(w_dff_A_1PUk7Ety7_0),.clk(gclk));
	jdff dff_A_LgyQ6g5M7_0(.dout(w_dff_A_1PUk7Ety7_0),.din(w_dff_A_LgyQ6g5M7_0),.clk(gclk));
	jdff dff_A_vEnIl3od7_0(.dout(w_dff_A_LgyQ6g5M7_0),.din(w_dff_A_vEnIl3od7_0),.clk(gclk));
	jdff dff_A_M6rDpDZN8_0(.dout(w_dff_A_vEnIl3od7_0),.din(w_dff_A_M6rDpDZN8_0),.clk(gclk));
	jdff dff_A_vFOH2N399_0(.dout(w_dff_A_M6rDpDZN8_0),.din(w_dff_A_vFOH2N399_0),.clk(gclk));
	jdff dff_A_mbP7sAWu4_0(.dout(w_dff_A_vFOH2N399_0),.din(w_dff_A_mbP7sAWu4_0),.clk(gclk));
	jdff dff_A_6l3GUOco6_0(.dout(w_dff_A_mbP7sAWu4_0),.din(w_dff_A_6l3GUOco6_0),.clk(gclk));
	jdff dff_A_J8e7MW7e3_0(.dout(w_dff_A_6l3GUOco6_0),.din(w_dff_A_J8e7MW7e3_0),.clk(gclk));
	jdff dff_A_9TFueqTW3_0(.dout(w_G85gat_0[0]),.din(w_dff_A_9TFueqTW3_0),.clk(gclk));
	jdff dff_A_UTDp6bgi1_0(.dout(w_dff_A_9TFueqTW3_0),.din(w_dff_A_UTDp6bgi1_0),.clk(gclk));
	jdff dff_A_WI44idSQ7_0(.dout(w_dff_A_UTDp6bgi1_0),.din(w_dff_A_WI44idSQ7_0),.clk(gclk));
	jdff dff_A_duHRM7dn9_0(.dout(w_dff_A_WI44idSQ7_0),.din(w_dff_A_duHRM7dn9_0),.clk(gclk));
	jdff dff_A_wdC1AY5R5_0(.dout(w_dff_A_duHRM7dn9_0),.din(w_dff_A_wdC1AY5R5_0),.clk(gclk));
	jdff dff_A_ThnwJJzD5_0(.dout(w_dff_A_wdC1AY5R5_0),.din(w_dff_A_ThnwJJzD5_0),.clk(gclk));
	jdff dff_A_Lih1vTLs0_0(.dout(w_dff_A_ThnwJJzD5_0),.din(w_dff_A_Lih1vTLs0_0),.clk(gclk));
	jdff dff_A_t73Q1kH36_0(.dout(w_dff_A_Lih1vTLs0_0),.din(w_dff_A_t73Q1kH36_0),.clk(gclk));
	jdff dff_A_G7YnaCet8_0(.dout(w_dff_A_t73Q1kH36_0),.din(w_dff_A_G7YnaCet8_0),.clk(gclk));
	jdff dff_A_539bRIsv3_0(.dout(w_dff_A_G7YnaCet8_0),.din(w_dff_A_539bRIsv3_0),.clk(gclk));
	jdff dff_A_ogvUz4vm1_0(.dout(w_dff_A_539bRIsv3_0),.din(w_dff_A_ogvUz4vm1_0),.clk(gclk));
	jdff dff_A_WGUmRrbA4_0(.dout(w_G106gat_0[0]),.din(w_dff_A_WGUmRrbA4_0),.clk(gclk));
	jdff dff_A_4XW7jGFD4_0(.dout(w_dff_A_WGUmRrbA4_0),.din(w_dff_A_4XW7jGFD4_0),.clk(gclk));
	jdff dff_A_V1JfakCo9_0(.dout(w_dff_A_4XW7jGFD4_0),.din(w_dff_A_V1JfakCo9_0),.clk(gclk));
	jdff dff_A_pLFom1cO5_0(.dout(w_dff_A_V1JfakCo9_0),.din(w_dff_A_pLFom1cO5_0),.clk(gclk));
	jdff dff_A_a7OoHm4U7_0(.dout(w_dff_A_pLFom1cO5_0),.din(w_dff_A_a7OoHm4U7_0),.clk(gclk));
	jdff dff_A_v4vRyEaP1_0(.dout(w_dff_A_a7OoHm4U7_0),.din(w_dff_A_v4vRyEaP1_0),.clk(gclk));
	jdff dff_A_EL1XSLtn3_0(.dout(w_dff_A_v4vRyEaP1_0),.din(w_dff_A_EL1XSLtn3_0),.clk(gclk));
	jdff dff_A_pvUwuCBL8_0(.dout(w_dff_A_EL1XSLtn3_0),.din(w_dff_A_pvUwuCBL8_0),.clk(gclk));
	jdff dff_A_FKu71oGJ6_0(.dout(w_dff_A_pvUwuCBL8_0),.din(w_dff_A_FKu71oGJ6_0),.clk(gclk));
	jdff dff_A_abmM5fXE4_0(.dout(w_dff_A_FKu71oGJ6_0),.din(w_dff_A_abmM5fXE4_0),.clk(gclk));
	jdff dff_A_zEYHoXXM2_0(.dout(w_dff_A_abmM5fXE4_0),.din(w_dff_A_zEYHoXXM2_0),.clk(gclk));
	jdff dff_A_jxH1okq01_0(.dout(w_G99gat_0[0]),.din(w_dff_A_jxH1okq01_0),.clk(gclk));
	jdff dff_A_KACfGxsG0_0(.dout(w_dff_A_jxH1okq01_0),.din(w_dff_A_KACfGxsG0_0),.clk(gclk));
	jdff dff_A_MKCBvkUz4_0(.dout(w_dff_A_KACfGxsG0_0),.din(w_dff_A_MKCBvkUz4_0),.clk(gclk));
	jdff dff_A_MzSnlUK85_0(.dout(w_dff_A_MKCBvkUz4_0),.din(w_dff_A_MzSnlUK85_0),.clk(gclk));
	jdff dff_A_XvIpWAEw2_0(.dout(w_dff_A_MzSnlUK85_0),.din(w_dff_A_XvIpWAEw2_0),.clk(gclk));
	jdff dff_A_KyC6agDj9_0(.dout(w_dff_A_XvIpWAEw2_0),.din(w_dff_A_KyC6agDj9_0),.clk(gclk));
	jdff dff_A_bekBbxnn6_0(.dout(w_dff_A_KyC6agDj9_0),.din(w_dff_A_bekBbxnn6_0),.clk(gclk));
	jdff dff_A_4aA0BhyM5_0(.dout(w_dff_A_bekBbxnn6_0),.din(w_dff_A_4aA0BhyM5_0),.clk(gclk));
	jdff dff_A_G4XyztvT0_0(.dout(w_dff_A_4aA0BhyM5_0),.din(w_dff_A_G4XyztvT0_0),.clk(gclk));
	jdff dff_A_Mw7a1sut3_0(.dout(w_dff_A_G4XyztvT0_0),.din(w_dff_A_Mw7a1sut3_0),.clk(gclk));
	jdff dff_A_p1F05AkQ9_0(.dout(w_dff_A_Mw7a1sut3_0),.din(w_dff_A_p1F05AkQ9_0),.clk(gclk));
	jdff dff_A_60qy12T34_0(.dout(w_G162gat_0[0]),.din(w_dff_A_60qy12T34_0),.clk(gclk));
	jdff dff_A_RgSEkwA58_0(.dout(w_dff_A_60qy12T34_0),.din(w_dff_A_RgSEkwA58_0),.clk(gclk));
	jdff dff_A_PoS3Xb0E1_0(.dout(w_dff_A_RgSEkwA58_0),.din(w_dff_A_PoS3Xb0E1_0),.clk(gclk));
	jdff dff_A_oLIAvyFR7_0(.dout(w_dff_A_PoS3Xb0E1_0),.din(w_dff_A_oLIAvyFR7_0),.clk(gclk));
	jdff dff_A_QW4mBDm74_0(.dout(w_dff_A_oLIAvyFR7_0),.din(w_dff_A_QW4mBDm74_0),.clk(gclk));
	jdff dff_A_y4Sd6yUH4_0(.dout(w_dff_A_QW4mBDm74_0),.din(w_dff_A_y4Sd6yUH4_0),.clk(gclk));
	jdff dff_A_3CTHyfGu1_0(.dout(w_dff_A_y4Sd6yUH4_0),.din(w_dff_A_3CTHyfGu1_0),.clk(gclk));
	jdff dff_A_eXDMBhMJ3_0(.dout(w_dff_A_3CTHyfGu1_0),.din(w_dff_A_eXDMBhMJ3_0),.clk(gclk));
	jdff dff_A_jgWMoFNs0_0(.dout(w_dff_A_eXDMBhMJ3_0),.din(w_dff_A_jgWMoFNs0_0),.clk(gclk));
	jdff dff_A_p16PEy079_0(.dout(w_dff_A_jgWMoFNs0_0),.din(w_dff_A_p16PEy079_0),.clk(gclk));
	jdff dff_A_XAMCx2EQ4_0(.dout(w_dff_A_p16PEy079_0),.din(w_dff_A_XAMCx2EQ4_0),.clk(gclk));
	jdff dff_A_drjs0qgZ6_0(.dout(w_G134gat_0[0]),.din(w_dff_A_drjs0qgZ6_0),.clk(gclk));
	jdff dff_A_w4W9N0gC2_0(.dout(w_dff_A_drjs0qgZ6_0),.din(w_dff_A_w4W9N0gC2_0),.clk(gclk));
	jdff dff_A_s5uTdpFC1_0(.dout(w_dff_A_w4W9N0gC2_0),.din(w_dff_A_s5uTdpFC1_0),.clk(gclk));
	jdff dff_A_zn0AjZ8j1_0(.dout(w_dff_A_s5uTdpFC1_0),.din(w_dff_A_zn0AjZ8j1_0),.clk(gclk));
	jdff dff_A_HjSzdfsR2_0(.dout(w_dff_A_zn0AjZ8j1_0),.din(w_dff_A_HjSzdfsR2_0),.clk(gclk));
	jdff dff_A_8EvGxAog9_0(.dout(w_dff_A_HjSzdfsR2_0),.din(w_dff_A_8EvGxAog9_0),.clk(gclk));
	jdff dff_A_ndqVGKcx9_0(.dout(w_dff_A_8EvGxAog9_0),.din(w_dff_A_ndqVGKcx9_0),.clk(gclk));
	jdff dff_A_TN4iO5KY6_0(.dout(w_dff_A_ndqVGKcx9_0),.din(w_dff_A_TN4iO5KY6_0),.clk(gclk));
	jdff dff_A_THdEW0hn9_0(.dout(w_dff_A_TN4iO5KY6_0),.din(w_dff_A_THdEW0hn9_0),.clk(gclk));
	jdff dff_A_UF18l7zG8_0(.dout(w_dff_A_THdEW0hn9_0),.din(w_dff_A_UF18l7zG8_0),.clk(gclk));
	jdff dff_A_veYjb4335_0(.dout(w_dff_A_UF18l7zG8_0),.din(w_dff_A_veYjb4335_0),.clk(gclk));
	jdff dff_A_k9ckY6gO7_0(.dout(w_G218gat_0[0]),.din(w_dff_A_k9ckY6gO7_0),.clk(gclk));
	jdff dff_A_HSPjeVkt8_0(.dout(w_dff_A_k9ckY6gO7_0),.din(w_dff_A_HSPjeVkt8_0),.clk(gclk));
	jdff dff_A_676eCCUB0_0(.dout(w_dff_A_HSPjeVkt8_0),.din(w_dff_A_676eCCUB0_0),.clk(gclk));
	jdff dff_A_lh4CpKCC9_0(.dout(w_dff_A_676eCCUB0_0),.din(w_dff_A_lh4CpKCC9_0),.clk(gclk));
	jdff dff_A_kbc9h4uc7_0(.dout(w_dff_A_lh4CpKCC9_0),.din(w_dff_A_kbc9h4uc7_0),.clk(gclk));
	jdff dff_A_3Mkj6noc0_0(.dout(w_dff_A_kbc9h4uc7_0),.din(w_dff_A_3Mkj6noc0_0),.clk(gclk));
	jdff dff_A_1Tym3ah83_0(.dout(w_dff_A_3Mkj6noc0_0),.din(w_dff_A_1Tym3ah83_0),.clk(gclk));
	jdff dff_A_Fk7Z8YEN9_0(.dout(w_dff_A_1Tym3ah83_0),.din(w_dff_A_Fk7Z8YEN9_0),.clk(gclk));
	jdff dff_A_62MbArOl0_0(.dout(w_dff_A_Fk7Z8YEN9_0),.din(w_dff_A_62MbArOl0_0),.clk(gclk));
	jdff dff_A_MiIvMP0N9_0(.dout(w_dff_A_62MbArOl0_0),.din(w_dff_A_MiIvMP0N9_0),.clk(gclk));
	jdff dff_A_odWp6WvU9_0(.dout(w_dff_A_MiIvMP0N9_0),.din(w_dff_A_odWp6WvU9_0),.clk(gclk));
	jdff dff_A_SU5SE6Es6_0(.dout(w_G190gat_0[0]),.din(w_dff_A_SU5SE6Es6_0),.clk(gclk));
	jdff dff_A_UvXJo7II8_0(.dout(w_dff_A_SU5SE6Es6_0),.din(w_dff_A_UvXJo7II8_0),.clk(gclk));
	jdff dff_A_SVfkbTlp9_0(.dout(w_dff_A_UvXJo7II8_0),.din(w_dff_A_SVfkbTlp9_0),.clk(gclk));
	jdff dff_A_yByDrXlw0_0(.dout(w_dff_A_SVfkbTlp9_0),.din(w_dff_A_yByDrXlw0_0),.clk(gclk));
	jdff dff_A_lNUBuyqd2_0(.dout(w_dff_A_yByDrXlw0_0),.din(w_dff_A_lNUBuyqd2_0),.clk(gclk));
	jdff dff_A_Sqv5eqQ09_0(.dout(w_dff_A_lNUBuyqd2_0),.din(w_dff_A_Sqv5eqQ09_0),.clk(gclk));
	jdff dff_A_XVXoWrNB6_0(.dout(w_dff_A_Sqv5eqQ09_0),.din(w_dff_A_XVXoWrNB6_0),.clk(gclk));
	jdff dff_A_YDslV3Dm6_0(.dout(w_dff_A_XVXoWrNB6_0),.din(w_dff_A_YDslV3Dm6_0),.clk(gclk));
	jdff dff_A_u5d3WRZt3_0(.dout(w_dff_A_YDslV3Dm6_0),.din(w_dff_A_u5d3WRZt3_0),.clk(gclk));
	jdff dff_A_Tt4PlzHN7_0(.dout(w_dff_A_u5d3WRZt3_0),.din(w_dff_A_Tt4PlzHN7_0),.clk(gclk));
	jdff dff_A_9BZA5ENF8_0(.dout(w_dff_A_Tt4PlzHN7_0),.din(w_dff_A_9BZA5ENF8_0),.clk(gclk));
endmodule

