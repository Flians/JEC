module gf_c1355(G233gat, G228gat, G229gat, G227gat, G218gat, G211gat, G197gat, G50gat, G64gat, G43gat, G232gat, G22gat, G36gat, G127gat, G29gat, G78gat, G230gat, G15gat, G8gat, G71gat, G120gat, G226gat, G162gat, G85gat, G57gat, G92gat, G1gat, G190gat, G148gat, G99gat, G155gat, G106gat, G225gat, G113gat, G134gat, G141gat, G204gat, G169gat, G176gat, G231gat, G183gat, G1353gat, G1355gat, G1335gat, G1338gat, G1334gat, G1332gat, G1340gat, G1354gat, G1331gat, G1329gat, G1350gat, G1352gat, G1328gat, G1327gat, G1336gat, G1326gat, G1341gat, G1344gat, G1333gat, G1325gat, G1343gat, G1330gat, G1339gat, G1337gat, G1342gat, G1324gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1351gat);
    input G233gat, G228gat, G229gat, G227gat, G218gat, G211gat, G197gat, G50gat, G64gat, G43gat, G232gat, G22gat, G36gat, G127gat, G29gat, G78gat, G230gat, G15gat, G8gat, G71gat, G120gat, G226gat, G162gat, G85gat, G57gat, G92gat, G1gat, G190gat, G148gat, G99gat, G155gat, G106gat, G225gat, G113gat, G134gat, G141gat, G204gat, G169gat, G176gat, G231gat, G183gat;
    output G1353gat, G1355gat, G1335gat, G1338gat, G1334gat, G1332gat, G1340gat, G1354gat, G1331gat, G1329gat, G1350gat, G1352gat, G1328gat, G1327gat, G1336gat, G1326gat, G1341gat, G1344gat, G1333gat, G1325gat, G1343gat, G1330gat, G1339gat, G1337gat, G1342gat, G1324gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1351gat;
    wire n76;
    wire n80;
    wire n84;
    wire n88;
    wire n92;
    wire n96;
    wire n100;
    wire n104;
    wire n107;
    wire n111;
    wire n115;
    wire n119;
    wire n123;
    wire n127;
    wire n130;
    wire n134;
    wire n138;
    wire n142;
    wire n146;
    wire n150;
    wire n154;
    wire n158;
    wire n161;
    wire n164;
    wire n168;
    wire n172;
    wire n176;
    wire n180;
    wire n184;
    wire n188;
    wire n192;
    wire n196;
    wire n200;
    wire n204;
    wire n208;
    wire n212;
    wire n216;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n243;
    wire n246;
    wire n250;
    wire n254;
    wire n258;
    wire n262;
    wire n266;
    wire n270;
    wire n274;
    wire n278;
    wire n282;
    wire n285;
    wire n289;
    wire n293;
    wire n297;
    wire n301;
    wire n305;
    wire n309;
    wire n313;
    wire n317;
    wire n321;
    wire n325;
    wire n328;
    wire n332;
    wire n336;
    wire n340;
    wire n344;
    wire n348;
    wire n352;
    wire n356;
    wire n359;
    wire n363;
    wire n367;
    wire n371;
    wire n375;
    wire n379;
    wire n383;
    wire n387;
    wire n391;
    wire n395;
    wire n399;
    wire n403;
    wire n407;
    wire n411;
    wire n415;
    wire n418;
    wire n422;
    wire n426;
    wire n429;
    wire n433;
    wire n437;
    wire n441;
    wire n445;
    wire n449;
    wire n452;
    wire n456;
    wire n460;
    wire n464;
    wire n468;
    wire n472;
    wire n476;
    wire n483;
    wire n487;
    wire n494;
    wire n498;
    wire n505;
    wire n509;
    wire n516;
    wire n520;
    wire n524;
    wire n528;
    wire n532;
    wire n540;
    wire n548;
    wire n556;
    wire n563;
    wire n567;
    wire n571;
    wire n575;
    wire n579;
    wire n587;
    wire n595;
    wire n603;
    wire n611;
    wire n615;
    wire n623;
    wire n631;
    wire n639;
    wire n647;
    wire n651;
    wire n655;
    wire n659;
    wire n663;
    wire n667;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n699;
    wire n707;
    wire n715;
    wire n723;
    wire n727;
    wire n731;
    wire n739;
    wire n747;
    wire n755;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n783;
    wire n791;
    wire n799;
    wire n807;
    wire n811;
    wire n819;
    wire n827;
    wire n835;
    wire n1215;
    wire n1219;
    wire n1222;
    wire n1224;
    wire n1228;
    wire n1231;
    wire n1234;
    wire n1237;
    wire n1240;
    wire n1243;
    wire n1246;
    wire n1249;
    wire n1251;
    wire n1254;
    wire n1257;
    wire n1260;
    wire n1263;
    wire n1266;
    wire n1269;
    wire n1272;
    wire n1275;
    wire n1278;
    wire n1281;
    wire n1284;
    wire n1287;
    wire n1290;
    wire n1293;
    wire n1296;
    wire n1299;
    wire n1302;
    wire n1305;
    wire n1308;
    wire n1311;
    wire n1314;
    wire n1317;
    wire n1320;
    wire n1323;
    wire n1326;
    wire n1329;
    wire n1332;
    wire n1335;
    wire n1338;
    wire n1341;
    wire n1344;
    wire n1348;
    wire n1351;
    wire n1353;
    wire n1356;
    wire n1359;
    wire n1362;
    wire n1365;
    wire n1368;
    wire n1371;
    wire n1374;
    wire n1377;
    wire n1380;
    wire n1383;
    wire n1386;
    wire n1389;
    wire n1392;
    wire n1395;
    wire n1398;
    wire n1401;
    wire n1404;
    wire n1407;
    wire n1410;
    wire n1414;
    wire n1417;
    wire n1420;
    wire n1422;
    wire n1425;
    wire n1428;
    wire n1431;
    wire n1434;
    wire n1437;
    wire n1440;
    wire n1443;
    wire n1446;
    wire n1449;
    wire n1452;
    wire n1455;
    wire n1458;
    wire n1461;
    wire n1464;
    wire n1467;
    wire n1470;
    wire n1473;
    wire n1476;
    wire n1479;
    wire n1482;
    wire n1485;
    wire n1488;
    wire n1491;
    wire n1494;
    wire n1497;
    wire n1500;
    wire n1503;
    wire n1506;
    wire n1509;
    wire n1512;
    wire n1515;
    wire n1518;
    wire n1521;
    wire n1524;
    wire n1527;
    wire n1530;
    wire n1533;
    wire n1536;
    wire n1539;
    wire n1542;
    wire n1545;
    wire n1548;
    wire n1552;
    wire n1555;
    wire n1558;
    wire n1560;
    wire n1563;
    wire n1566;
    wire n1569;
    wire n1572;
    wire n1575;
    wire n1578;
    wire n1581;
    wire n1584;
    wire n1587;
    wire n1590;
    wire n1593;
    wire n1596;
    wire n1599;
    wire n1602;
    wire n1605;
    wire n1608;
    wire n1611;
    wire n1614;
    wire n1617;
    wire n1620;
    wire n1623;
    wire n1626;
    wire n1629;
    wire n1632;
    wire n1635;
    wire n1638;
    wire n1641;
    wire n1644;
    wire n1647;
    wire n1650;
    wire n1653;
    wire n1656;
    wire n1659;
    wire n1662;
    wire n1665;
    wire n1668;
    wire n1671;
    wire n1674;
    wire n1677;
    wire n1680;
    wire n1683;
    wire n1686;
    wire n1689;
    wire n1692;
    wire n1695;
    wire n1698;
    wire n1701;
    wire n1704;
    wire n1707;
    wire n1710;
    wire n1713;
    wire n1716;
    wire n1719;
    wire n1722;
    wire n1725;
    wire n1728;
    wire n1731;
    wire n1734;
    wire n1737;
    wire n1741;
    wire n1744;
    wire n1747;
    wire n1749;
    wire n1752;
    wire n1755;
    wire n1758;
    wire n1761;
    wire n1764;
    wire n1767;
    wire n1770;
    wire n1773;
    wire n1776;
    wire n1779;
    wire n1782;
    wire n1785;
    wire n1788;
    wire n1791;
    wire n1794;
    wire n1797;
    wire n1800;
    wire n1803;
    wire n1806;
    wire n1809;
    wire n1812;
    wire n1815;
    wire n1818;
    wire n1821;
    wire n1824;
    wire n1827;
    wire n1830;
    wire n1833;
    wire n1836;
    wire n1839;
    wire n1842;
    wire n1845;
    wire n1848;
    wire n1851;
    wire n1854;
    wire n1857;
    wire n1860;
    wire n1863;
    wire n1866;
    wire n1869;
    wire n1872;
    wire n1875;
    wire n1878;
    wire n1881;
    wire n1884;
    wire n1887;
    wire n1890;
    wire n1893;
    wire n1896;
    wire n1899;
    wire n1902;
    wire n1905;
    wire n1908;
    wire n1911;
    wire n1914;
    wire n1917;
    wire n1920;
    wire n1923;
    wire n1926;
    wire n1929;
    wire n1932;
    wire n1935;
    wire n1938;
    wire n1941;
    wire n1944;
    wire n1947;
    wire n1950;
    wire n1953;
    wire n1956;
    wire n1959;
    wire n1962;
    wire n1965;
    wire n1968;
    wire n1971;
    wire n1974;
    wire n1977;
    wire n1980;
    wire n1983;
    wire n1986;
    wire n1989;
    wire n1992;
    wire n1995;
    wire n1998;
    wire n2001;
    wire n2004;
    wire n2007;
    wire n2010;
    wire n2013;
    wire n2016;
    wire n2019;
    wire n2022;
    wire n2025;
    wire n2028;
    wire n2031;
    wire n2034;
    wire n2037;
    wire n2040;
    wire n2043;
    wire n2046;
    wire n2049;
    wire n2052;
    wire n2055;
    wire n2058;
    wire n2061;
    wire n2064;
    wire n2067;
    wire n2070;
    wire n2073;
    wire n2076;
    wire n2079;
    wire n2082;
    wire n2085;
    wire n2088;
    wire n2091;
    wire n2094;
    wire n2097;
    wire n2100;
    wire n2103;
    wire n2106;
    wire n2109;
    wire n2112;
    wire n2115;
    wire n2118;
    wire n2121;
    wire n2124;
    wire n2127;
    wire n2130;
    wire n2133;
    wire n2136;
    wire n2139;
    wire n2142;
    wire n2145;
    wire n2148;
    wire n2151;
    wire n2154;
    wire n2157;
    wire n2160;
    wire n2163;
    wire n2166;
    wire n2169;
    wire n2172;
    wire n2175;
    wire n2178;
    wire n2181;
    wire n2184;
    wire n2187;
    wire n2190;
    wire n2193;
    wire n2196;
    wire n2199;
    wire n2202;
    wire n2205;
    wire n2208;
    wire n2211;
    wire n2214;
    wire n2217;
    wire n2220;
    wire n2223;
    wire n2226;
    wire n2229;
    wire n2232;
    wire n2235;
    wire n2238;
    wire n2241;
    wire n2244;
    wire n2247;
    wire n2250;
    wire n2253;
    wire n2256;
    wire n2259;
    wire n2262;
    wire n2265;
    wire n2268;
    wire n2271;
    wire n2274;
    wire n2277;
    wire n2280;
    wire n2283;
    wire n2286;
    wire n2289;
    wire n2292;
    wire n2295;
    wire n2298;
    wire n2301;
    wire n2304;
    wire n2307;
    wire n2310;
    wire n2313;
    wire n2316;
    wire n2319;
    wire n2322;
    wire n2325;
    wire n2328;
    wire n2331;
    wire n2334;
    wire n2337;
    wire n2340;
    wire n2343;
    wire n2346;
    wire n2349;
    wire n2352;
    wire n2355;
    wire n2358;
    wire n2361;
    wire n2364;
    wire n2367;
    wire n2370;
    wire n2373;
    wire n2376;
    wire n2379;
    wire n2382;
    wire n2385;
    wire n2388;
    wire n2391;
    wire n2394;
    wire n2397;
    wire n2400;
    wire n2403;
    wire n2406;
    wire n2409;
    wire n2412;
    wire n2415;
    wire n2418;
    wire n2421;
    wire n2424;
    wire n2427;
    wire n2430;
    wire n2433;
    wire n2436;
    wire n2439;
    wire n2442;
    wire n2445;
    wire n2448;
    wire n2451;
    wire n2454;
    wire n2457;
    wire n2460;
    wire n2463;
    wire n2466;
    wire n2469;
    wire n2472;
    wire n2475;
    wire n2478;
    wire n2481;
    wire n2484;
    wire n2487;
    wire n2490;
    wire n2493;
    wire n2496;
    wire n2499;
    wire n2502;
    wire n2505;
    wire n2508;
    wire n2511;
    wire n2514;
    wire n2517;
    wire n2520;
    wire n2523;
    wire n2526;
    wire n2529;
    wire n2532;
    wire n2535;
    wire n2538;
    wire n2541;
    wire n2544;
    wire n2547;
    wire n2550;
    wire n2553;
    wire n2556;
    wire n2559;
    wire n2562;
    wire n2565;
    wire n2568;
    wire n2571;
    wire n2574;
    wire n2577;
    wire n2580;
    wire n2583;
    wire n2586;
    wire n2589;
    wire n2592;
    wire n2595;
    wire n2598;
    wire n2601;
    wire n2604;
    wire n2607;
    wire n2610;
    wire n2613;
    wire n2616;
    wire n2619;
    wire n2622;
    wire n2625;
    wire n2628;
    wire n2631;
    wire n2634;
    wire n2637;
    wire n2640;
    wire n2643;
    wire n2646;
    wire n2649;
    wire n2652;
    wire n2655;
    wire n2658;
    wire n2661;
    wire n2664;
    wire n2667;
    wire n2670;
    wire n2673;
    wire n2676;
    wire n2679;
    wire n2682;
    wire n2685;
    wire n2688;
    wire n2691;
    wire n2694;
    wire n2697;
    wire n2700;
    wire n2703;
    wire n2706;
    wire n2709;
    wire n2712;
    wire n2715;
    wire n2718;
    wire n2721;
    wire n2724;
    wire n2727;
    wire n2730;
    wire n2733;
    wire n2736;
    wire n2739;
    jxor g000(.dinb(G57gat), .dina(G85gat), .dout(n76));
    jxor g001(.dinb(G1gat), .dina(G29gat), .dout(n80));
    jxor g002(.dinb(n76), .dina(n80), .dout(n84));
    jxor g003(.dinb(G155gat), .dina(G162gat), .dout(n88));
    jxor g004(.dinb(G141gat), .dina(G148gat), .dout(n92));
    jxor g005(.dinb(n88), .dina(n92), .dout(n96));
    jxor g006(.dinb(n84), .dina(n96), .dout(n100));
    jand g007(.dinb(G225gat), .dina(G233gat), .dout(n104));
    jnot g008(.din(n104), .dout(n107));
    jxor g009(.dinb(G127gat), .dina(G134gat), .dout(n111));
    jxor g010(.dinb(G113gat), .dina(G120gat), .dout(n115));
    jxor g011(.dinb(n111), .dina(n115), .dout(n119));
    jxor g012(.dinb(n107), .dina(n119), .dout(n123));
    jxor g013(.dinb(n100), .dina(n123), .dout(n127));
    jnot g014(.din(n127), .dout(n130));
    jxor g015(.dinb(G190gat), .dina(G218gat), .dout(n134));
    jxor g016(.dinb(G134gat), .dina(G162gat), .dout(n138));
    jxor g017(.dinb(n134), .dina(n138), .dout(n142));
    jxor g018(.dinb(G99gat), .dina(G106gat), .dout(n146));
    jxor g019(.dinb(G85gat), .dina(G92gat), .dout(n150));
    jxor g020(.dinb(n146), .dina(n150), .dout(n154));
    jxor g021(.dinb(n142), .dina(n154), .dout(n158));
    jnot g022(.din(G232gat), .dout(n161));
    jnot g023(.din(G233gat), .dout(n164));
    jor g024(.dinb(n161), .dina(n164), .dout(n168));
    jxor g025(.dinb(G43gat), .dina(G50gat), .dout(n172));
    jxor g026(.dinb(G29gat), .dina(G36gat), .dout(n176));
    jxor g027(.dinb(n172), .dina(n176), .dout(n180));
    jxor g028(.dinb(n168), .dina(n180), .dout(n184));
    jxor g029(.dinb(n158), .dina(n184), .dout(n188));
    jxor g030(.dinb(G183gat), .dina(G211gat), .dout(n192));
    jxor g031(.dinb(G127gat), .dina(G155gat), .dout(n196));
    jxor g032(.dinb(n192), .dina(n196), .dout(n200));
    jxor g033(.dinb(G71gat), .dina(G78gat), .dout(n204));
    jxor g034(.dinb(G57gat), .dina(G64gat), .dout(n208));
    jxor g035(.dinb(n204), .dina(n208), .dout(n212));
    jxor g036(.dinb(n200), .dina(n212), .dout(n216));
    jnot g037(.din(G231gat), .dout(n219));
    jor g038(.dinb(n219), .dina(n164), .dout(n223));
    jxor g039(.dinb(G15gat), .dina(G22gat), .dout(n227));
    jxor g040(.dinb(G1gat), .dina(G8gat), .dout(n231));
    jxor g041(.dinb(n227), .dina(n231), .dout(n235));
    jxor g042(.dinb(n223), .dina(n235), .dout(n239));
    jxor g043(.dinb(n216), .dina(n239), .dout(n243));
    jnot g044(.din(n243), .dout(n246));
    jand g045(.dinb(n2343), .dina(n246), .dout(n250));
    jxor g046(.dinb(G64gat), .dina(G92gat), .dout(n254));
    jxor g047(.dinb(G8gat), .dina(G36gat), .dout(n258));
    jxor g048(.dinb(n254), .dina(n258), .dout(n262));
    jxor g049(.dinb(G183gat), .dina(G190gat), .dout(n266));
    jxor g050(.dinb(G169gat), .dina(G176gat), .dout(n270));
    jxor g051(.dinb(n266), .dina(n270), .dout(n274));
    jxor g052(.dinb(n262), .dina(n274), .dout(n278));
    jand g053(.dinb(G226gat), .dina(G233gat), .dout(n282));
    jnot g054(.din(n282), .dout(n285));
    jxor g055(.dinb(G211gat), .dina(G218gat), .dout(n289));
    jxor g056(.dinb(G197gat), .dina(G204gat), .dout(n293));
    jxor g057(.dinb(n289), .dina(n293), .dout(n297));
    jxor g058(.dinb(n285), .dina(n297), .dout(n301));
    jxor g059(.dinb(n278), .dina(n301), .dout(n305));
    jxor g060(.dinb(n127), .dina(n305), .dout(n309));
    jxor g061(.dinb(G71gat), .dina(G99gat), .dout(n313));
    jxor g062(.dinb(G15gat), .dina(G43gat), .dout(n317));
    jxor g063(.dinb(n313), .dina(n317), .dout(n321));
    jxor g064(.dinb(n274), .dina(n321), .dout(n325));
    jnot g065(.din(G227gat), .dout(n328));
    jor g066(.dinb(n328), .dina(n164), .dout(n332));
    jxor g067(.dinb(n119), .dina(n332), .dout(n336));
    jxor g068(.dinb(n325), .dina(n336), .dout(n340));
    jxor g069(.dinb(G78gat), .dina(G106gat), .dout(n344));
    jxor g070(.dinb(G22gat), .dina(G50gat), .dout(n348));
    jxor g071(.dinb(n344), .dina(n348), .dout(n352));
    jxor g072(.dinb(n297), .dina(n352), .dout(n356));
    jnot g073(.din(G228gat), .dout(n359));
    jor g074(.dinb(n359), .dina(n164), .dout(n363));
    jxor g075(.dinb(n96), .dina(n363), .dout(n367));
    jxor g076(.dinb(n356), .dina(n367), .dout(n371));
    jand g077(.dinb(n340), .dina(n371), .dout(n375));
    jand g078(.dinb(n309), .dina(n375), .dout(n379));
    jxor g079(.dinb(n340), .dina(n371), .dout(n383));
    jand g080(.dinb(n1671), .dina(n383), .dout(n387));
    jand g081(.dinb(n1251), .dina(n387), .dout(n391));
    jor g082(.dinb(n1249), .dina(n391), .dout(n395));
    jxor g083(.dinb(G169gat), .dina(G197gat), .dout(n399));
    jxor g084(.dinb(G113gat), .dina(G141gat), .dout(n403));
    jxor g085(.dinb(n399), .dina(n403), .dout(n407));
    jxor g086(.dinb(n235), .dina(n407), .dout(n411));
    jand g087(.dinb(G229gat), .dina(G233gat), .dout(n415));
    jnot g088(.din(n415), .dout(n418));
    jxor g089(.dinb(n180), .dina(n418), .dout(n422));
    jxor g090(.dinb(n411), .dina(n422), .dout(n426));
    jnot g091(.din(n426), .dout(n429));
    jxor g092(.dinb(G176gat), .dina(G204gat), .dout(n433));
    jxor g093(.dinb(G120gat), .dina(G148gat), .dout(n437));
    jxor g094(.dinb(n433), .dina(n437), .dout(n441));
    jxor g095(.dinb(n212), .dina(n441), .dout(n445));
    jand g096(.dinb(G230gat), .dina(G233gat), .dout(n449));
    jnot g097(.din(n449), .dout(n452));
    jxor g098(.dinb(n154), .dina(n452), .dout(n456));
    jxor g099(.dinb(n445), .dina(n456), .dout(n460));
    jand g100(.dinb(n429), .dina(n1515), .dout(n464));
    jand g101(.dinb(n395), .dina(n1222), .dout(n468));
    jand g102(.dinb(n1224), .dina(n468), .dout(n472));
    jand g103(.dinb(n1353), .dina(n472), .dout(n476));
    jxor g104(.dinb(n1674), .dina(n476), .dout(G1324gat));
    jnot g105(.din(n305), .dout(n483));
    jand g106(.dinb(n1569), .dina(n472), .dout(n487));
    jxor g107(.dinb(n1602), .dina(n487), .dout(G1325gat));
    jnot g108(.din(n340), .dout(n494));
    jand g109(.dinb(n1422), .dina(n472), .dout(n498));
    jxor g110(.dinb(n2148), .dina(n498), .dout(G1326gat));
    jnot g111(.din(n371), .dout(n505));
    jand g112(.dinb(n1749), .dina(n472), .dout(n509));
    jxor g113(.dinb(n1881), .dina(n509), .dout(G1327gat));
    jnot g114(.din(n188), .dout(n516));
    jand g115(.dinb(n516), .dina(n1548), .dout(n520));
    jand g116(.dinb(n395), .dina(n1246), .dout(n524));
    jand g117(.dinb(n1215), .dina(n524), .dout(n528));
    jand g118(.dinb(n1353), .dina(n528), .dout(n532));
    jxor g119(.dinb(n2379), .dina(n532), .dout(G1328gat));
    jand g120(.dinb(n1569), .dina(n528), .dout(n540));
    jxor g121(.dinb(n2346), .dina(n540), .dout(G1329gat));
    jand g122(.dinb(n1422), .dina(n528), .dout(n548));
    jxor g123(.dinb(n2445), .dina(n548), .dout(G1330gat));
    jand g124(.dinb(n1749), .dina(n528), .dout(n556));
    jxor g125(.dinb(n2412), .dina(n556), .dout(G1331gat));
    jnot g126(.din(n460), .dout(n563));
    jand g127(.dinb(n1482), .dina(n563), .dout(n567));
    jand g128(.dinb(n1231), .dina(n395), .dout(n571));
    jand g129(.dinb(n1240), .dina(n571), .dout(n575));
    jand g130(.dinb(n1353), .dina(n575), .dout(n579));
    jxor g131(.dinb(n1707), .dina(n579), .dout(G1332gat));
    jand g132(.dinb(n1569), .dina(n575), .dout(n587));
    jxor g133(.dinb(n1635), .dina(n587), .dout(G1333gat));
    jand g134(.dinb(n1422), .dina(n575), .dout(n595));
    jxor g135(.dinb(n2181), .dina(n595), .dout(G1334gat));
    jand g136(.dinb(n1749), .dina(n575), .dout(n603));
    jxor g137(.dinb(n1914), .dina(n603), .dout(G1335gat));
    jand g138(.dinb(n524), .dina(n1240), .dout(n611));
    jand g139(.dinb(n1368), .dina(n611), .dout(n615));
    jxor g140(.dinb(n2511), .dina(n615), .dout(G1336gat));
    jand g141(.dinb(n1584), .dina(n611), .dout(n623));
    jxor g142(.dinb(n2478), .dina(n623), .dout(G1337gat));
    jand g143(.dinb(n1437), .dina(n611), .dout(n631));
    jxor g144(.dinb(n2577), .dina(n631), .dout(G1338gat));
    jand g145(.dinb(n1764), .dina(n611), .dout(n639));
    jxor g146(.dinb(n2544), .dina(n639), .dout(G1339gat));
    jand g147(.dinb(n494), .dina(n1779), .dout(n647));
    jand g148(.dinb(n130), .dina(n1599), .dout(n651));
    jxor g149(.dinb(n188), .dina(n243), .dout(n655));
    jand g150(.dinb(n1560), .dina(n655), .dout(n659));
    jand g151(.dinb(n1563), .dina(n659), .dout(n663));
    jxor g152(.dinb(n426), .dina(n460), .dout(n667));
    jand g153(.dinb(n188), .dina(n243), .dout(n671));
    jand g154(.dinb(n667), .dina(n671), .dout(n675));
    jor g155(.dinb(n663), .dina(n1558), .dout(n679));
    jand g156(.dinb(n1351), .dina(n679), .dout(n683));
    jand g157(.dinb(n1420), .dina(n683), .dout(n687));
    jand g158(.dinb(n1272), .dina(n687), .dout(n691));
    jxor g159(.dinb(n2082), .dina(n691), .dout(G1340gat));
    jand g160(.dinb(n1302), .dina(n687), .dout(n699));
    jxor g161(.dinb(n2049), .dina(n699), .dout(G1341gat));
    jand g162(.dinb(n1332), .dina(n687), .dout(n707));
    jxor g163(.dinb(n2115), .dina(n707), .dout(G1342gat));
    jand g164(.dinb(n1398), .dina(n687), .dout(n715));
    jxor g165(.dinb(n2643), .dina(n715), .dout(G1343gat));
    jand g166(.dinb(n2046), .dina(n505), .dout(n723));
    jand g167(.dinb(n1747), .dina(n683), .dout(n727));
    jand g168(.dinb(n1257), .dina(n727), .dout(n731));
    jxor g169(.dinb(n1815), .dina(n731), .dout(G1344gat));
    jand g170(.dinb(n1287), .dina(n727), .dout(n739));
    jxor g171(.dinb(n1782), .dina(n739), .dout(G1345gat));
    jand g172(.dinb(n1317), .dina(n727), .dout(n747));
    jxor g173(.dinb(n1848), .dina(n747), .dout(G1346gat));
    jand g174(.dinb(n1383), .dina(n727), .dout(n755));
    jxor g175(.dinb(n2610), .dina(n755), .dout(G1347gat));
    jand g176(.dinb(n1668), .dina(n483), .dout(n763));
    jand g177(.dinb(n1555), .dina(n679), .dout(n767));
    jand g178(.dinb(n1420), .dina(n767), .dout(n771));
    jand g179(.dinb(n1467), .dina(n771), .dout(n775));
    jxor g180(.dinb(n2247), .dina(n775), .dout(G1348gat));
    jand g181(.dinb(n1500), .dina(n771), .dout(n783));
    jxor g182(.dinb(n2214), .dina(n783), .dout(G1349gat));
    jand g183(.dinb(n1533), .dina(n771), .dout(n791));
    jxor g184(.dinb(n2280), .dina(n791), .dout(G1350gat));
    jand g185(.dinb(n2328), .dina(n771), .dout(n799));
    jxor g186(.dinb(n2709), .dina(n799), .dout(G1351gat));
    jand g187(.dinb(n1747), .dina(n767), .dout(n807));
    jand g188(.dinb(n1452), .dina(n807), .dout(n811));
    jxor g189(.dinb(n1980), .dina(n811), .dout(G1352gat));
    jand g190(.dinb(n1485), .dina(n807), .dout(n819));
    jxor g191(.dinb(n1947), .dina(n819), .dout(G1353gat));
    jand g192(.dinb(n1518), .dina(n807), .dout(n827));
    jxor g193(.dinb(n2013), .dina(n827), .dout(G1354gat));
    jand g194(.dinb(n2313), .dina(n807), .dout(n835));
    jxor g195(.dinb(n2676), .dina(n835), .dout(G1355gat));
    jdff dff_A_KQTvHfr49_0(.din(G190gat), .dout(n2739));
    jdff dff_A_ioNA677y0_0(.din(n2739), .dout(n2736));
    jdff dff_A_zZHpXqXw9_0(.din(n2736), .dout(n2733));
    jdff dff_A_fMsTXQ4I3_0(.din(n2733), .dout(n2730));
    jdff dff_A_metjIlrp0_0(.din(n2730), .dout(n2727));
    jdff dff_A_HIZilLLr7_0(.din(n2727), .dout(n2724));
    jdff dff_A_PxWIvayd9_0(.din(n2724), .dout(n2721));
    jdff dff_A_WtTdz0lC0_0(.din(n2721), .dout(n2718));
    jdff dff_A_FqwzPC3E8_0(.din(n2718), .dout(n2715));
    jdff dff_A_uK1a1sii7_0(.din(n2715), .dout(n2712));
    jdff dff_A_FapeOVY95_0(.din(n2712), .dout(n2709));
    jdff dff_A_jkYTbfyn8_0(.din(G218gat), .dout(n2706));
    jdff dff_A_sRof27eR9_0(.din(n2706), .dout(n2703));
    jdff dff_A_F1eypsoi6_0(.din(n2703), .dout(n2700));
    jdff dff_A_iIiGKZl39_0(.din(n2700), .dout(n2697));
    jdff dff_A_pkKkitfx9_0(.din(n2697), .dout(n2694));
    jdff dff_A_YT6aLnYY2_0(.din(n2694), .dout(n2691));
    jdff dff_A_m43anPMI1_0(.din(n2691), .dout(n2688));
    jdff dff_A_3tq7bs351_0(.din(n2688), .dout(n2685));
    jdff dff_A_Ckrg3HfM2_0(.din(n2685), .dout(n2682));
    jdff dff_A_wxcsNfRJ6_0(.din(n2682), .dout(n2679));
    jdff dff_A_deLr8FPU4_0(.din(n2679), .dout(n2676));
    jdff dff_A_vKv8bSYv9_0(.din(G134gat), .dout(n2673));
    jdff dff_A_IjZ9WPvP0_0(.din(n2673), .dout(n2670));
    jdff dff_A_nQYkzxOf3_0(.din(n2670), .dout(n2667));
    jdff dff_A_XtmNMhD51_0(.din(n2667), .dout(n2664));
    jdff dff_A_o1QY7sx44_0(.din(n2664), .dout(n2661));
    jdff dff_A_6S06bhx94_0(.din(n2661), .dout(n2658));
    jdff dff_A_S6I0eFoT7_0(.din(n2658), .dout(n2655));
    jdff dff_A_d7lTRz1w1_0(.din(n2655), .dout(n2652));
    jdff dff_A_ydDsvXT58_0(.din(n2652), .dout(n2649));
    jdff dff_A_moTWRqlj4_0(.din(n2649), .dout(n2646));
    jdff dff_A_6FqbQmRT9_0(.din(n2646), .dout(n2643));
    jdff dff_A_M94Wx5ES3_0(.din(G162gat), .dout(n2640));
    jdff dff_A_9kXPIB2g0_0(.din(n2640), .dout(n2637));
    jdff dff_A_XylOKzOO5_0(.din(n2637), .dout(n2634));
    jdff dff_A_0Hk51g9W6_0(.din(n2634), .dout(n2631));
    jdff dff_A_6iyMxZ369_0(.din(n2631), .dout(n2628));
    jdff dff_A_7OnIDFpU2_0(.din(n2628), .dout(n2625));
    jdff dff_A_5PlTz9Gj5_0(.din(n2625), .dout(n2622));
    jdff dff_A_lH4RvTb54_0(.din(n2622), .dout(n2619));
    jdff dff_A_uYZ9ddvD0_0(.din(n2619), .dout(n2616));
    jdff dff_A_VWJb7aaj1_0(.din(n2616), .dout(n2613));
    jdff dff_A_8SAwAT9O2_0(.din(n2613), .dout(n2610));
    jdff dff_A_qsVz5g8R4_0(.din(G99gat), .dout(n2607));
    jdff dff_A_7rpyD8io6_0(.din(n2607), .dout(n2604));
    jdff dff_A_wxeVzPs08_0(.din(n2604), .dout(n2601));
    jdff dff_A_asTS1FeR3_0(.din(n2601), .dout(n2598));
    jdff dff_A_MWMyUdxS1_0(.din(n2598), .dout(n2595));
    jdff dff_A_aRgEUGVX7_0(.din(n2595), .dout(n2592));
    jdff dff_A_JAZzS8LO5_0(.din(n2592), .dout(n2589));
    jdff dff_A_zG7HLKGw9_0(.din(n2589), .dout(n2586));
    jdff dff_A_Qs8IxPQU4_0(.din(n2586), .dout(n2583));
    jdff dff_A_ekdPj6c14_0(.din(n2583), .dout(n2580));
    jdff dff_A_qbVd0D6m1_0(.din(n2580), .dout(n2577));
    jdff dff_A_1TLSdQqz3_0(.din(G106gat), .dout(n2574));
    jdff dff_A_iHtSzie08_0(.din(n2574), .dout(n2571));
    jdff dff_A_qcu5Rdl66_0(.din(n2571), .dout(n2568));
    jdff dff_A_AurYlREi0_0(.din(n2568), .dout(n2565));
    jdff dff_A_avvZpOWE5_0(.din(n2565), .dout(n2562));
    jdff dff_A_CqkDwW2h5_0(.din(n2562), .dout(n2559));
    jdff dff_A_0nrKv9xc9_0(.din(n2559), .dout(n2556));
    jdff dff_A_XMDCLix27_0(.din(n2556), .dout(n2553));
    jdff dff_A_3bjSki6M1_0(.din(n2553), .dout(n2550));
    jdff dff_A_LlqxGvMB3_0(.din(n2550), .dout(n2547));
    jdff dff_A_ptDHawF33_0(.din(n2547), .dout(n2544));
    jdff dff_A_ScOY6LQa6_0(.din(G85gat), .dout(n2541));
    jdff dff_A_9v7HP2XB4_0(.din(n2541), .dout(n2538));
    jdff dff_A_Z5xDBAup9_0(.din(n2538), .dout(n2535));
    jdff dff_A_yQ2U1kXz8_0(.din(n2535), .dout(n2532));
    jdff dff_A_7cCj6nXZ7_0(.din(n2532), .dout(n2529));
    jdff dff_A_v9i7mDaN7_0(.din(n2529), .dout(n2526));
    jdff dff_A_5cf0d9z87_0(.din(n2526), .dout(n2523));
    jdff dff_A_VJFhodmT2_0(.din(n2523), .dout(n2520));
    jdff dff_A_9WyYmbh25_0(.din(n2520), .dout(n2517));
    jdff dff_A_KIflMu126_0(.din(n2517), .dout(n2514));
    jdff dff_A_Pxm2Hynp3_0(.din(n2514), .dout(n2511));
    jdff dff_A_fOGk2Zs59_0(.din(G92gat), .dout(n2508));
    jdff dff_A_1WTtnRBD1_0(.din(n2508), .dout(n2505));
    jdff dff_A_8jt1bLpO0_0(.din(n2505), .dout(n2502));
    jdff dff_A_4iVMijiM8_0(.din(n2502), .dout(n2499));
    jdff dff_A_5qgA06l26_0(.din(n2499), .dout(n2496));
    jdff dff_A_e6HsgDU97_0(.din(n2496), .dout(n2493));
    jdff dff_A_33XygtPg9_0(.din(n2493), .dout(n2490));
    jdff dff_A_N5Ot1bJF0_0(.din(n2490), .dout(n2487));
    jdff dff_A_N5jH4jXA9_0(.din(n2487), .dout(n2484));
    jdff dff_A_4xUDPzTL8_0(.din(n2484), .dout(n2481));
    jdff dff_A_oghYpZ7M3_0(.din(n2481), .dout(n2478));
    jdff dff_A_EWk6wSym1_0(.din(G43gat), .dout(n2475));
    jdff dff_A_W5moqzen2_0(.din(n2475), .dout(n2472));
    jdff dff_A_rXxZgoZN9_0(.din(n2472), .dout(n2469));
    jdff dff_A_iVB6eI8q1_0(.din(n2469), .dout(n2466));
    jdff dff_A_vEymCU7L9_0(.din(n2466), .dout(n2463));
    jdff dff_A_mvr7PKmQ0_0(.din(n2463), .dout(n2460));
    jdff dff_A_dBIHdzLw4_0(.din(n2460), .dout(n2457));
    jdff dff_A_EagGbAgF2_0(.din(n2457), .dout(n2454));
    jdff dff_A_jkxtHo3y3_0(.din(n2454), .dout(n2451));
    jdff dff_A_Hr4RJzin2_0(.din(n2451), .dout(n2448));
    jdff dff_A_tKZgqRDz6_0(.din(n2448), .dout(n2445));
    jdff dff_A_6CKFAuNy6_0(.din(G50gat), .dout(n2442));
    jdff dff_A_Cry3SQuq9_0(.din(n2442), .dout(n2439));
    jdff dff_A_n8FL9cNI3_0(.din(n2439), .dout(n2436));
    jdff dff_A_g7fWtRC34_0(.din(n1222), .dout(n1215));
    jdff dff_B_UbdA9TpT0_2(.din(n464), .dout(n1219));
    jdff dff_B_XLzfbrYo1_2(.din(n1219), .dout(n1222));
    jdff dff_A_XFMs5PF89_1(.din(n1231), .dout(n1224));
    jdff dff_B_C82Ol07Z2_2(.din(n250), .dout(n1228));
    jdff dff_B_cMdmeUqR9_2(.din(n1228), .dout(n1231));
    jdff dff_B_oD2VeBYI1_2(.din(n567), .dout(n1234));
    jdff dff_B_uXMssaTF3_2(.din(n1234), .dout(n1237));
    jdff dff_B_ictF7VVB8_2(.din(n1237), .dout(n1240));
    jdff dff_B_fEXmCUEr6_0(.din(n520), .dout(n1243));
    jdff dff_B_qvVbhgQM2_0(.din(n1243), .dout(n1246));
    jdff dff_B_IfNW47ib0_1(.din(n379), .dout(n1249));
    jdff dff_A_4kRfFieY2_0(.din(n1254), .dout(n1251));
    jdff dff_A_qvU4pT7M9_0(.din(n305), .dout(n1254));
    jdff dff_A_w5BUOEI76_0(.din(n1260), .dout(n1257));
    jdff dff_A_WOeCCUnT6_0(.din(n1263), .dout(n1260));
    jdff dff_A_pjcl3KMO5_0(.din(n1266), .dout(n1263));
    jdff dff_A_bM5Ydb574_0(.din(n1269), .dout(n1266));
    jdff dff_A_FZGlmU2N4_0(.din(n429), .dout(n1269));
    jdff dff_A_GY3GUQUV5_1(.din(n1275), .dout(n1272));
    jdff dff_A_bbxDdLtV6_1(.din(n1278), .dout(n1275));
    jdff dff_A_a0vgmC6X2_1(.din(n1281), .dout(n1278));
    jdff dff_A_xdfdtWBd6_1(.din(n1284), .dout(n1281));
    jdff dff_A_sFVdG6WN0_1(.din(n429), .dout(n1284));
    jdff dff_A_qJ5zHxs81_0(.din(n1290), .dout(n1287));
    jdff dff_A_K1PQJV6P4_0(.din(n1293), .dout(n1290));
    jdff dff_A_Fo4NdyDl9_0(.din(n1296), .dout(n1293));
    jdff dff_A_cNwRv10B6_0(.din(n1299), .dout(n1296));
    jdff dff_A_iuTgCrL40_0(.din(n563), .dout(n1299));
    jdff dff_A_0mjTla9J4_1(.din(n1305), .dout(n1302));
    jdff dff_A_MkIJKXmu7_1(.din(n1308), .dout(n1305));
    jdff dff_A_Br5tP2ke6_1(.din(n1311), .dout(n1308));
    jdff dff_A_kJVItLlC5_1(.din(n1314), .dout(n1311));
    jdff dff_A_pFx1qlrF2_1(.din(n563), .dout(n1314));
    jdff dff_A_NyHcnITN2_0(.din(n1320), .dout(n1317));
    jdff dff_A_PjEsC2Nt6_0(.din(n1323), .dout(n1320));
    jdff dff_A_9hMNiwAr7_0(.din(n1326), .dout(n1323));
    jdff dff_A_3FNVJZ6b6_0(.din(n1329), .dout(n1326));
    jdff dff_A_BvcpixTz4_0(.din(n246), .dout(n1329));
    jdff dff_A_OhMm5bUl1_1(.din(n1335), .dout(n1332));
    jdff dff_A_FNmPuiPJ4_1(.din(n1338), .dout(n1335));
    jdff dff_A_wzYEryQA7_1(.din(n1341), .dout(n1338));
    jdff dff_A_NlQU0y8n4_1(.din(n1344), .dout(n1341));
    jdff dff_A_ANbbw8Pr3_1(.din(n246), .dout(n1344));
    jdff dff_B_I3NQ9kWv8_1(.din(n651), .dout(n1348));
    jdff dff_B_X2Im87NO5_1(.din(n1348), .dout(n1351));
    jdff dff_A_nkRXkBK28_0(.din(n1356), .dout(n1353));
    jdff dff_A_y2E5kge90_0(.din(n1359), .dout(n1356));
    jdff dff_A_N0Qm4qx03_0(.din(n1362), .dout(n1359));
    jdff dff_A_KE3xKRPJ8_0(.din(n1365), .dout(n1362));
    jdff dff_A_HDvR5fGe3_0(.din(n130), .dout(n1365));
    jdff dff_A_r5DYRlB56_2(.din(n1371), .dout(n1368));
    jdff dff_A_EXqygMbt8_2(.din(n1374), .dout(n1371));
    jdff dff_A_8TN8oAwb5_2(.din(n1377), .dout(n1374));
    jdff dff_A_kg3pIg939_2(.din(n1380), .dout(n1377));
    jdff dff_A_7DImgA5K9_2(.din(n130), .dout(n1380));
    jdff dff_A_oCgw7TMx6_0(.din(n1386), .dout(n1383));
    jdff dff_A_I1aMf9ZZ5_0(.din(n1389), .dout(n1386));
    jdff dff_A_YeY29Oym9_0(.din(n1392), .dout(n1389));
    jdff dff_A_zBAy3kXJ3_0(.din(n1395), .dout(n1392));
    jdff dff_A_pFG4FcaY0_0(.din(n516), .dout(n1395));
    jdff dff_A_OnF2YcdG6_1(.din(n1401), .dout(n1398));
    jdff dff_A_mPYlZrow8_1(.din(n1404), .dout(n1401));
    jdff dff_A_fx5E7a5D4_1(.din(n1407), .dout(n1404));
    jdff dff_A_CitHGTA41_1(.din(n1410), .dout(n1407));
    jdff dff_A_2DYJGpGs2_1(.din(n516), .dout(n1410));
    jdff dff_B_Bvp8kghG2_2(.din(n647), .dout(n1414));
    jdff dff_B_hw1dCfcE1_2(.din(n1414), .dout(n1417));
    jdff dff_B_ZnnCJ2u80_2(.din(n1417), .dout(n1420));
    jdff dff_A_tAxc8FNh3_0(.din(n1425), .dout(n1422));
    jdff dff_A_H9RAuYj59_0(.din(n1428), .dout(n1425));
    jdff dff_A_zhKE0ORh8_0(.din(n1431), .dout(n1428));
    jdff dff_A_978ixOg97_0(.din(n1434), .dout(n1431));
    jdff dff_A_Z09T7J496_0(.din(n494), .dout(n1434));
    jdff dff_A_9vEsrmUR1_2(.din(n1440), .dout(n1437));
    jdff dff_A_3GTNAkxF1_2(.din(n1443), .dout(n1440));
    jdff dff_A_S26JRI2o8_2(.din(n1446), .dout(n1443));
    jdff dff_A_hf96O2073_2(.din(n1449), .dout(n1446));
    jdff dff_A_KepHnE5C4_2(.din(n494), .dout(n1449));
    jdff dff_A_Pq1Q8flQ6_1(.din(n1455), .dout(n1452));
    jdff dff_A_tiXy71DX0_1(.din(n1458), .dout(n1455));
    jdff dff_A_J1RAxLIK9_1(.din(n1461), .dout(n1458));
    jdff dff_A_xA55UyWX5_1(.din(n1464), .dout(n1461));
    jdff dff_A_fiIPpVW66_1(.din(n429), .dout(n1464));
    jdff dff_A_IZxkOlFJ1_2(.din(n1470), .dout(n1467));
    jdff dff_A_PRQAdJrd6_2(.din(n1473), .dout(n1470));
    jdff dff_A_ruYlIlni4_2(.din(n1476), .dout(n1473));
    jdff dff_A_OatywFOG1_2(.din(n1479), .dout(n1476));
    jdff dff_A_neoNnWwU3_2(.din(n429), .dout(n1479));
    jdff dff_A_9woERz7Z9_0(.din(n426), .dout(n1482));
    jdff dff_A_cI7o6xKU6_1(.din(n1488), .dout(n1485));
    jdff dff_A_p6IPhVq52_1(.din(n1491), .dout(n1488));
    jdff dff_A_x5ATtBGA0_1(.din(n1494), .dout(n1491));
    jdff dff_A_s89WmVE65_1(.din(n1497), .dout(n1494));
    jdff dff_A_Pt4jPtr59_1(.din(n563), .dout(n1497));
    jdff dff_A_jw7x2tkw3_2(.din(n1503), .dout(n1500));
    jdff dff_A_6WsW1NfW8_2(.din(n1506), .dout(n1503));
    jdff dff_A_ShANqaSA1_2(.din(n1509), .dout(n1506));
    jdff dff_A_qOihlfpz6_2(.din(n1512), .dout(n1509));
    jdff dff_A_dDSIcMPD8_2(.din(n563), .dout(n1512));
    jdff dff_A_Y51j7kVV7_1(.din(n460), .dout(n1515));
    jdff dff_A_NqSOUP0c2_1(.din(n1521), .dout(n1518));
    jdff dff_A_G3ZB9A949_1(.din(n1524), .dout(n1521));
    jdff dff_A_chUHDdp50_1(.din(n1527), .dout(n1524));
    jdff dff_A_kjcJgFsq5_1(.din(n1530), .dout(n1527));
    jdff dff_A_C2tRsLlm2_1(.din(n246), .dout(n1530));
    jdff dff_A_7ayfKDEO3_2(.din(n1536), .dout(n1533));
    jdff dff_A_2uRtdZbc2_2(.din(n1539), .dout(n1536));
    jdff dff_A_4uP4cjSF1_2(.din(n1542), .dout(n1539));
    jdff dff_A_grZsy7Tu6_2(.din(n1545), .dout(n1542));
    jdff dff_A_6rL5Wax43_2(.din(n246), .dout(n1545));
    jdff dff_A_rIYE9OzL2_0(.din(n243), .dout(n1548));
    jdff dff_B_qyGoOx4d0_1(.din(n763), .dout(n1552));
    jdff dff_B_gMAT52TG0_1(.din(n1552), .dout(n1555));
    jdff dff_B_kBn5VUQX0_0(.din(n675), .dout(n1558));
    jdff dff_A_xsODTihY7_2(.din(n426), .dout(n1560));
    jdff dff_A_k2sYJBL53_2(.din(n1566), .dout(n1563));
    jdff dff_A_xz3I73mA6_2(.din(n460), .dout(n1566));
    jdff dff_A_g5l9RMl53_0(.din(n1572), .dout(n1569));
    jdff dff_A_y8KyCeV62_0(.din(n1575), .dout(n1572));
    jdff dff_A_ifxEZZu00_0(.din(n1578), .dout(n1575));
    jdff dff_A_SBY2aqI75_0(.din(n1581), .dout(n1578));
    jdff dff_A_awOn1qiS3_0(.din(n483), .dout(n1581));
    jdff dff_A_PzVgNCOy3_2(.din(n1587), .dout(n1584));
    jdff dff_A_kj68dVfq5_2(.din(n1590), .dout(n1587));
    jdff dff_A_BI0MT9n17_2(.din(n1593), .dout(n1590));
    jdff dff_A_45F2Wfbn4_2(.din(n1596), .dout(n1593));
    jdff dff_A_IBdGzWN69_2(.din(n483), .dout(n1596));
    jdff dff_A_bOqX34r50_1(.din(n305), .dout(n1599));
    jdff dff_A_nRDA2vYG6_0(.din(n1605), .dout(n1602));
    jdff dff_A_Mym3gcbE7_0(.din(n1608), .dout(n1605));
    jdff dff_A_gRCIq3DY7_0(.din(n1611), .dout(n1608));
    jdff dff_A_tfc7ibsH7_0(.din(n1614), .dout(n1611));
    jdff dff_A_pNPAEwfB1_0(.din(n1617), .dout(n1614));
    jdff dff_A_H3vghLHm2_0(.din(n1620), .dout(n1617));
    jdff dff_A_XkM3NqXz1_0(.din(n1623), .dout(n1620));
    jdff dff_A_UTLB9La62_0(.din(n1626), .dout(n1623));
    jdff dff_A_nvOZlLyp4_0(.din(n1629), .dout(n1626));
    jdff dff_A_eKpGKkJK3_0(.din(n1632), .dout(n1629));
    jdff dff_A_iq1FECP85_0(.din(G8gat), .dout(n1632));
    jdff dff_A_LLwYrFqp7_0(.din(n1638), .dout(n1635));
    jdff dff_A_VMHuDbXW2_0(.din(n1641), .dout(n1638));
    jdff dff_A_6k0ZNcJS5_0(.din(n1644), .dout(n1641));
    jdff dff_A_MY4xu2Sr4_0(.din(n1647), .dout(n1644));
    jdff dff_A_d58reL1z1_0(.din(n1650), .dout(n1647));
    jdff dff_A_57UHzbkQ8_0(.din(n1653), .dout(n1650));
    jdff dff_A_817YCMfQ3_0(.din(n1656), .dout(n1653));
    jdff dff_A_IG27HCOo2_0(.din(n1659), .dout(n1656));
    jdff dff_A_p8E3sw4r8_0(.din(n1662), .dout(n1659));
    jdff dff_A_tEUrMgvT0_0(.din(n1665), .dout(n1662));
    jdff dff_A_D3IYoDKs3_0(.din(G64gat), .dout(n1665));
    jdff dff_A_wHstNy2b2_1(.din(n127), .dout(n1668));
    jdff dff_A_5WUuWzmE9_2(.din(n127), .dout(n1671));
    jdff dff_A_aMsv7RJo4_0(.din(n1677), .dout(n1674));
    jdff dff_A_fqzMkq1x0_0(.din(n1680), .dout(n1677));
    jdff dff_A_mnjIAAwl1_0(.din(n1683), .dout(n1680));
    jdff dff_A_Q0rJsq7D2_0(.din(n1686), .dout(n1683));
    jdff dff_A_zwJqievP9_0(.din(n1689), .dout(n1686));
    jdff dff_A_8rcd7bQa7_0(.din(n1692), .dout(n1689));
    jdff dff_A_nXwlvstj8_0(.din(n1695), .dout(n1692));
    jdff dff_A_HLWbYNWE0_0(.din(n1698), .dout(n1695));
    jdff dff_A_FSgxPSWq7_0(.din(n1701), .dout(n1698));
    jdff dff_A_JCZNzEoJ9_0(.din(n1704), .dout(n1701));
    jdff dff_A_UcmzbQkh5_0(.din(G1gat), .dout(n1704));
    jdff dff_A_B88P9Sez4_0(.din(n1710), .dout(n1707));
    jdff dff_A_FnxcZ3DO9_0(.din(n1713), .dout(n1710));
    jdff dff_A_46g3VgXk0_0(.din(n1716), .dout(n1713));
    jdff dff_A_e3Uxfk0L0_0(.din(n1719), .dout(n1716));
    jdff dff_A_D6pRyXT40_0(.din(n1722), .dout(n1719));
    jdff dff_A_AiXwK1vd9_0(.din(n1725), .dout(n1722));
    jdff dff_A_z5VEzgME0_0(.din(n1728), .dout(n1725));
    jdff dff_A_5sV6vwcA1_0(.din(n1731), .dout(n1728));
    jdff dff_A_8Uo2JvBy7_0(.din(n1734), .dout(n1731));
    jdff dff_A_sADhmOWS6_0(.din(n1737), .dout(n1734));
    jdff dff_A_l9rnSSI04_0(.din(G57gat), .dout(n1737));
    jdff dff_B_HSHaE9Ih2_2(.din(n723), .dout(n1741));
    jdff dff_B_XNRly9na4_2(.din(n1741), .dout(n1744));
    jdff dff_B_nHxscb9U4_2(.din(n1744), .dout(n1747));
    jdff dff_A_y1RUfWp32_0(.din(n1752), .dout(n1749));
    jdff dff_A_j7cpPJAr6_0(.din(n1755), .dout(n1752));
    jdff dff_A_YIskqoSz7_0(.din(n1758), .dout(n1755));
    jdff dff_A_mmKCDQrv0_0(.din(n1761), .dout(n1758));
    jdff dff_A_QkSzTCdN3_0(.din(n505), .dout(n1761));
    jdff dff_A_M1aNCpEq0_2(.din(n1767), .dout(n1764));
    jdff dff_A_xxP5WCIH0_2(.din(n1770), .dout(n1767));
    jdff dff_A_5wqRAZPE4_2(.din(n1773), .dout(n1770));
    jdff dff_A_3ECLkrun6_2(.din(n1776), .dout(n1773));
    jdff dff_A_JKedJh0d4_2(.din(n505), .dout(n1776));
    jdff dff_A_GSwAHdKK6_1(.din(n371), .dout(n1779));
    jdff dff_A_ddD5a0Aw5_0(.din(n1785), .dout(n1782));
    jdff dff_A_hvyyoF785_0(.din(n1788), .dout(n1785));
    jdff dff_A_vOxg2hAo2_0(.din(n1791), .dout(n1788));
    jdff dff_A_ptyxYr8f2_0(.din(n1794), .dout(n1791));
    jdff dff_A_BSBT0qQK9_0(.din(n1797), .dout(n1794));
    jdff dff_A_7QY9nNvq6_0(.din(n1800), .dout(n1797));
    jdff dff_A_np3P7awH0_0(.din(n1803), .dout(n1800));
    jdff dff_A_gixtXHhu8_0(.din(n1806), .dout(n1803));
    jdff dff_A_16IA2rWe6_0(.din(n1809), .dout(n1806));
    jdff dff_A_XwxqnrD51_0(.din(n1812), .dout(n1809));
    jdff dff_A_rrqo86Nk9_0(.din(G148gat), .dout(n1812));
    jdff dff_A_5ZT7LSoQ0_0(.din(n1818), .dout(n1815));
    jdff dff_A_bTiiKfGM2_0(.din(n1821), .dout(n1818));
    jdff dff_A_fZCFhG694_0(.din(n1824), .dout(n1821));
    jdff dff_A_sNfeIk8T6_0(.din(n1827), .dout(n1824));
    jdff dff_A_d1EHCy0X4_0(.din(n1830), .dout(n1827));
    jdff dff_A_7ulYWxJU5_0(.din(n1833), .dout(n1830));
    jdff dff_A_sRQ6aVyO3_0(.din(n1836), .dout(n1833));
    jdff dff_A_fDNR9epd3_0(.din(n1839), .dout(n1836));
    jdff dff_A_wBEH4Wj33_0(.din(n1842), .dout(n1839));
    jdff dff_A_DeyXqbRp9_0(.din(n1845), .dout(n1842));
    jdff dff_A_4US1ySSH8_0(.din(G141gat), .dout(n1845));
    jdff dff_A_lnIce6xP3_0(.din(n1851), .dout(n1848));
    jdff dff_A_sic6zVz01_0(.din(n1854), .dout(n1851));
    jdff dff_A_rwoTpeUC7_0(.din(n1857), .dout(n1854));
    jdff dff_A_ZGUuCZRu1_0(.din(n1860), .dout(n1857));
    jdff dff_A_uamd48YW7_0(.din(n1863), .dout(n1860));
    jdff dff_A_8UeOxRJh2_0(.din(n1866), .dout(n1863));
    jdff dff_A_LNp6Muz40_0(.din(n1869), .dout(n1866));
    jdff dff_A_s02xCIfa1_0(.din(n1872), .dout(n1869));
    jdff dff_A_TKIVSopJ8_0(.din(n1875), .dout(n1872));
    jdff dff_A_U2BrVfOt1_0(.din(n1878), .dout(n1875));
    jdff dff_A_Q9CXhgde5_0(.din(G155gat), .dout(n1878));
    jdff dff_A_53kmCpTX7_0(.din(n1884), .dout(n1881));
    jdff dff_A_hyBkMIIC4_0(.din(n1887), .dout(n1884));
    jdff dff_A_wiS5E5NZ3_0(.din(n1890), .dout(n1887));
    jdff dff_A_85Ht0P2y9_0(.din(n1893), .dout(n1890));
    jdff dff_A_rdvvKlaS2_0(.din(n1896), .dout(n1893));
    jdff dff_A_EDDOjM8Z0_0(.din(n1899), .dout(n1896));
    jdff dff_A_vDLbXTvY4_0(.din(n1902), .dout(n1899));
    jdff dff_A_qmiZIMVd8_0(.din(n1905), .dout(n1902));
    jdff dff_A_nv0TeVXs4_0(.din(n1908), .dout(n1905));
    jdff dff_A_8e3J57y30_0(.din(n1911), .dout(n1908));
    jdff dff_A_axs5ry7q1_0(.din(G22gat), .dout(n1911));
    jdff dff_A_x43OYFnI8_0(.din(n1917), .dout(n1914));
    jdff dff_A_9WX8LZch9_0(.din(n1920), .dout(n1917));
    jdff dff_A_vkyOKHke5_0(.din(n1923), .dout(n1920));
    jdff dff_A_2NzI4PPC1_0(.din(n1926), .dout(n1923));
    jdff dff_A_W5cq667D0_0(.din(n1929), .dout(n1926));
    jdff dff_A_QDoA0WXj3_0(.din(n1932), .dout(n1929));
    jdff dff_A_bJzb9TiQ3_0(.din(n1935), .dout(n1932));
    jdff dff_A_KiDbmSMU7_0(.din(n1938), .dout(n1935));
    jdff dff_A_IRWXDphX8_0(.din(n1941), .dout(n1938));
    jdff dff_A_Rv7Ika1y6_0(.din(n1944), .dout(n1941));
    jdff dff_A_RaPgyqEB0_0(.din(G78gat), .dout(n1944));
    jdff dff_A_8UClQlks9_0(.din(n1950), .dout(n1947));
    jdff dff_A_aDxvsTPX7_0(.din(n1953), .dout(n1950));
    jdff dff_A_oFeujOQt1_0(.din(n1956), .dout(n1953));
    jdff dff_A_10V6IQla6_0(.din(n1959), .dout(n1956));
    jdff dff_A_76AAjDM61_0(.din(n1962), .dout(n1959));
    jdff dff_A_4OFky0sv7_0(.din(n1965), .dout(n1962));
    jdff dff_A_DrSqs3n32_0(.din(n1968), .dout(n1965));
    jdff dff_A_AjUdYfVM5_0(.din(n1971), .dout(n1968));
    jdff dff_A_4tQryBox6_0(.din(n1974), .dout(n1971));
    jdff dff_A_zRUc7yJH0_0(.din(n1977), .dout(n1974));
    jdff dff_A_NpQuwQpU9_0(.din(G204gat), .dout(n1977));
    jdff dff_A_0kag68kR1_0(.din(n1983), .dout(n1980));
    jdff dff_A_zjPOeu2C6_0(.din(n1986), .dout(n1983));
    jdff dff_A_Bc0fjxVV8_0(.din(n1989), .dout(n1986));
    jdff dff_A_VWomtTTY1_0(.din(n1992), .dout(n1989));
    jdff dff_A_RgvbKDty8_0(.din(n1995), .dout(n1992));
    jdff dff_A_EH6tmStE3_0(.din(n1998), .dout(n1995));
    jdff dff_A_2WpoxvPT7_0(.din(n2001), .dout(n1998));
    jdff dff_A_F3OywF0E2_0(.din(n2004), .dout(n2001));
    jdff dff_A_ZYFOHQcy8_0(.din(n2007), .dout(n2004));
    jdff dff_A_lVVieE0z3_0(.din(n2010), .dout(n2007));
    jdff dff_A_vfHsKIz05_0(.din(G197gat), .dout(n2010));
    jdff dff_A_tUPJ8xBQ2_0(.din(n2016), .dout(n2013));
    jdff dff_A_qJpb2hhC9_0(.din(n2019), .dout(n2016));
    jdff dff_A_mZlViL2C3_0(.din(n2022), .dout(n2019));
    jdff dff_A_dIzhVf4v7_0(.din(n2025), .dout(n2022));
    jdff dff_A_JhQ1WFom2_0(.din(n2028), .dout(n2025));
    jdff dff_A_HrFpJHTX4_0(.din(n2031), .dout(n2028));
    jdff dff_A_i1uTj3yO9_0(.din(n2034), .dout(n2031));
    jdff dff_A_Kdk8Zcjt9_0(.din(n2037), .dout(n2034));
    jdff dff_A_zsblTJ4d8_0(.din(n2040), .dout(n2037));
    jdff dff_A_dU3kP5r20_0(.din(n2043), .dout(n2040));
    jdff dff_A_yreAeIPE7_0(.din(G211gat), .dout(n2043));
    jdff dff_A_gx2kTY761_1(.din(n340), .dout(n2046));
    jdff dff_A_KvbXou8D0_0(.din(n2052), .dout(n2049));
    jdff dff_A_RvvEEplq5_0(.din(n2055), .dout(n2052));
    jdff dff_A_RSoabOWz8_0(.din(n2058), .dout(n2055));
    jdff dff_A_A6blB7S96_0(.din(n2061), .dout(n2058));
    jdff dff_A_zNJAKhRu8_0(.din(n2064), .dout(n2061));
    jdff dff_A_ef7t8ovF2_0(.din(n2067), .dout(n2064));
    jdff dff_A_6EwLDQLU9_0(.din(n2070), .dout(n2067));
    jdff dff_A_GOkfIyGo4_0(.din(n2073), .dout(n2070));
    jdff dff_A_Pu10F1fI7_0(.din(n2076), .dout(n2073));
    jdff dff_A_VpVb5lPW9_0(.din(n2079), .dout(n2076));
    jdff dff_A_RNbr4DrG7_0(.din(G120gat), .dout(n2079));
    jdff dff_A_Uvq2ISC13_0(.din(n2085), .dout(n2082));
    jdff dff_A_7NHM8MYj7_0(.din(n2088), .dout(n2085));
    jdff dff_A_2B33gQmD1_0(.din(n2091), .dout(n2088));
    jdff dff_A_VU7Wfq9c0_0(.din(n2094), .dout(n2091));
    jdff dff_A_E64gVZvF1_0(.din(n2097), .dout(n2094));
    jdff dff_A_oTj1Gib57_0(.din(n2100), .dout(n2097));
    jdff dff_A_3QTYpOlI5_0(.din(n2103), .dout(n2100));
    jdff dff_A_InFSudi49_0(.din(n2106), .dout(n2103));
    jdff dff_A_cckRExhv2_0(.din(n2109), .dout(n2106));
    jdff dff_A_FDtq2BbX6_0(.din(n2112), .dout(n2109));
    jdff dff_A_9ZJCqNHa9_0(.din(G113gat), .dout(n2112));
    jdff dff_A_xLHFZHh25_0(.din(n2118), .dout(n2115));
    jdff dff_A_jH5hUEm57_0(.din(n2121), .dout(n2118));
    jdff dff_A_k2y2WbVO4_0(.din(n2124), .dout(n2121));
    jdff dff_A_KPvoMPps7_0(.din(n2127), .dout(n2124));
    jdff dff_A_zoXmEvjH7_0(.din(n2130), .dout(n2127));
    jdff dff_A_I9ltBUix1_0(.din(n2133), .dout(n2130));
    jdff dff_A_8rerxCpB2_0(.din(n2136), .dout(n2133));
    jdff dff_A_zOoOuxQo5_0(.din(n2139), .dout(n2136));
    jdff dff_A_dyUIIFQ78_0(.din(n2142), .dout(n2139));
    jdff dff_A_NW3saaZP9_0(.din(n2145), .dout(n2142));
    jdff dff_A_WzdV4eai8_0(.din(G127gat), .dout(n2145));
    jdff dff_A_e4m04q3B9_0(.din(n2151), .dout(n2148));
    jdff dff_A_aJENA3Po1_0(.din(n2154), .dout(n2151));
    jdff dff_A_CnrwW58Q0_0(.din(n2157), .dout(n2154));
    jdff dff_A_aITPlvab5_0(.din(n2160), .dout(n2157));
    jdff dff_A_1UeYkWGW6_0(.din(n2163), .dout(n2160));
    jdff dff_A_mnYtbXEY3_0(.din(n2166), .dout(n2163));
    jdff dff_A_AfU7IXd18_0(.din(n2169), .dout(n2166));
    jdff dff_A_57nUM4lY3_0(.din(n2172), .dout(n2169));
    jdff dff_A_7qUonzYj2_0(.din(n2175), .dout(n2172));
    jdff dff_A_JAcdjA6v9_0(.din(n2178), .dout(n2175));
    jdff dff_A_DGF6gZJt9_0(.din(G15gat), .dout(n2178));
    jdff dff_A_iWPGaqeT9_0(.din(n2184), .dout(n2181));
    jdff dff_A_tHhgsdKJ8_0(.din(n2187), .dout(n2184));
    jdff dff_A_XLpT9dqa2_0(.din(n2190), .dout(n2187));
    jdff dff_A_j4B1sx2o1_0(.din(n2193), .dout(n2190));
    jdff dff_A_AbQnepcZ1_0(.din(n2196), .dout(n2193));
    jdff dff_A_k9osiVcG7_0(.din(n2199), .dout(n2196));
    jdff dff_A_VFCyZIEE9_0(.din(n2202), .dout(n2199));
    jdff dff_A_QFLZhNPM4_0(.din(n2205), .dout(n2202));
    jdff dff_A_h6RqiRQ63_0(.din(n2208), .dout(n2205));
    jdff dff_A_tPOqLmLd3_0(.din(n2211), .dout(n2208));
    jdff dff_A_tVGFvDGq0_0(.din(G71gat), .dout(n2211));
    jdff dff_A_V7659hYV8_0(.din(n2217), .dout(n2214));
    jdff dff_A_904aWuNT2_0(.din(n2220), .dout(n2217));
    jdff dff_A_dkWeLLyS6_0(.din(n2223), .dout(n2220));
    jdff dff_A_t7yj3dmV4_0(.din(n2226), .dout(n2223));
    jdff dff_A_tKFWOP2H5_0(.din(n2229), .dout(n2226));
    jdff dff_A_TcfeqVxa7_0(.din(n2232), .dout(n2229));
    jdff dff_A_0nMjYDmr2_0(.din(n2235), .dout(n2232));
    jdff dff_A_zret7jSo2_0(.din(n2238), .dout(n2235));
    jdff dff_A_YIBYXjAd8_0(.din(n2241), .dout(n2238));
    jdff dff_A_J88dYbRL2_0(.din(n2244), .dout(n2241));
    jdff dff_A_7v7dT4Ll9_0(.din(G176gat), .dout(n2244));
    jdff dff_A_KjBgybxO9_0(.din(n2250), .dout(n2247));
    jdff dff_A_luIVE5603_0(.din(n2253), .dout(n2250));
    jdff dff_A_rTeWKTuK5_0(.din(n2256), .dout(n2253));
    jdff dff_A_UqGw2XlN2_0(.din(n2259), .dout(n2256));
    jdff dff_A_CENrdQJ84_0(.din(n2262), .dout(n2259));
    jdff dff_A_PmM4NndX9_0(.din(n2265), .dout(n2262));
    jdff dff_A_RHrH6hO82_0(.din(n2268), .dout(n2265));
    jdff dff_A_fue47tCg2_0(.din(n2271), .dout(n2268));
    jdff dff_A_8NznfdDM5_0(.din(n2274), .dout(n2271));
    jdff dff_A_CuWHA5Yp4_0(.din(n2277), .dout(n2274));
    jdff dff_A_M6HBiUCH5_0(.din(G169gat), .dout(n2277));
    jdff dff_A_oJO62Rp16_0(.din(n2283), .dout(n2280));
    jdff dff_A_z7UbHL3d5_0(.din(n2286), .dout(n2283));
    jdff dff_A_1aYYLMj23_0(.din(n2289), .dout(n2286));
    jdff dff_A_ZyrqKgsj1_0(.din(n2292), .dout(n2289));
    jdff dff_A_Z1jwAMuK9_0(.din(n2295), .dout(n2292));
    jdff dff_A_tPPdVKKG0_0(.din(n2298), .dout(n2295));
    jdff dff_A_sfJWps624_0(.din(n2301), .dout(n2298));
    jdff dff_A_EJdh07eS4_0(.din(n2304), .dout(n2301));
    jdff dff_A_cJdhGI191_0(.din(n2307), .dout(n2304));
    jdff dff_A_ocWcBmRt3_0(.din(n2310), .dout(n2307));
    jdff dff_A_ZQIL4zOV3_0(.din(G183gat), .dout(n2310));
    jdff dff_A_TnMHhmql2_1(.din(n2316), .dout(n2313));
    jdff dff_A_CxeUrvIJ4_1(.din(n2319), .dout(n2316));
    jdff dff_A_JCTjOkmL1_1(.din(n2322), .dout(n2319));
    jdff dff_A_PrT1bVMz2_1(.din(n2325), .dout(n2322));
    jdff dff_A_oKvAYkiG8_1(.din(n516), .dout(n2325));
    jdff dff_A_DSe6qKbN2_2(.din(n2331), .dout(n2328));
    jdff dff_A_lkQsU6Fo1_2(.din(n2334), .dout(n2331));
    jdff dff_A_hFQ7RFzM3_2(.din(n2337), .dout(n2334));
    jdff dff_A_TYAYYZlu6_2(.din(n2340), .dout(n2337));
    jdff dff_A_oeYXzT0W7_2(.din(n516), .dout(n2340));
    jdff dff_A_XXy1jOTI2_1(.din(n188), .dout(n2343));
    jdff dff_A_JWYMyi2G2_0(.din(n2349), .dout(n2346));
    jdff dff_A_YhzLEPzi5_0(.din(n2352), .dout(n2349));
    jdff dff_A_laAcwvOq2_0(.din(n2355), .dout(n2352));
    jdff dff_A_HfW89dTG3_0(.din(n2358), .dout(n2355));
    jdff dff_A_uloYN7lo4_0(.din(n2361), .dout(n2358));
    jdff dff_A_Z1pFR60o7_0(.din(n2364), .dout(n2361));
    jdff dff_A_gOBFhiLk5_0(.din(n2367), .dout(n2364));
    jdff dff_A_Tih0hyYL3_0(.din(n2370), .dout(n2367));
    jdff dff_A_YgeUGz0u3_0(.din(n2373), .dout(n2370));
    jdff dff_A_952dId8H4_0(.din(n2376), .dout(n2373));
    jdff dff_A_drLvg0bw5_0(.din(G36gat), .dout(n2376));
    jdff dff_A_8NgL0byW5_0(.din(n2382), .dout(n2379));
    jdff dff_A_jhBVRKmS9_0(.din(n2385), .dout(n2382));
    jdff dff_A_ajgQ6ECf4_0(.din(n2388), .dout(n2385));
    jdff dff_A_M3mEFDcA5_0(.din(n2391), .dout(n2388));
    jdff dff_A_xjhhtLpD2_0(.din(n2394), .dout(n2391));
    jdff dff_A_lgbpSjju5_0(.din(n2397), .dout(n2394));
    jdff dff_A_Xf7ek1yO6_0(.din(n2400), .dout(n2397));
    jdff dff_A_ZBlzI3ey8_0(.din(n2403), .dout(n2400));
    jdff dff_A_8fY33f0s7_0(.din(n2406), .dout(n2403));
    jdff dff_A_eBECbbOr7_0(.din(n2409), .dout(n2406));
    jdff dff_A_OB7GilfJ9_0(.din(G29gat), .dout(n2409));
    jdff dff_A_PifLK1KF9_0(.din(n2415), .dout(n2412));
    jdff dff_A_lN9CVWBF2_0(.din(n2418), .dout(n2415));
    jdff dff_A_zcT3cTsb7_0(.din(n2421), .dout(n2418));
    jdff dff_A_E5vlx3Ay8_0(.din(n2424), .dout(n2421));
    jdff dff_A_c1PhGR751_0(.din(n2427), .dout(n2424));
    jdff dff_A_9QnLx7LZ2_0(.din(n2430), .dout(n2427));
    jdff dff_A_XFIyex0l2_0(.din(n2433), .dout(n2430));
    jdff dff_A_OGklGDSh0_0(.din(n2436), .dout(n2433));
endmodule

