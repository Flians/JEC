// Benchmark "top" written by ABC on Thu May 28 22:01:20 2020

module gf_square ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] ;
  wire n193, n195, n196, n197, n198, n200, n201, n202, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632, n633, n634, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
    n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
    n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
    n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
    n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
    n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
    n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
    n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
    n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
    n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
    n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
    n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
    n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
    n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
    n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
    n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3532, n3533,
    n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
    n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
    n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
    n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
    n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
    n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
    n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
    n4770, n4771, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
    n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
    n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
    n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
    n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
    n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
    n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
    n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
    n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
    n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
    n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
    n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5579, n5580, n5581, n5582, n5583, n5584,
    n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
    n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
    n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5794, n5795,
    n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
    n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
    n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
    n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
    n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
    n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
    n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
    n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
    n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011, n6013, n6014, n6015, n6016,
    n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
    n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
    n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
    n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
    n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
    n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
    n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
    n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
    n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
    n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
    n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
    n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
    n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
    n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
    n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
    n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
    n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
    n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
    n6438, n6439, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
    n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
    n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
    n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
    n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
    n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
    n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
    n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
    n6659, n6660, n6661, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
    n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
    n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
    n6870, n6871, n6872, n6873, n6874, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
    n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
    n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
    n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
    n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
    n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
    n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
    n7322, n7323, n7324, n7325, n7326, n7327, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
    n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
    n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
    n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
    n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
    n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
    n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
    n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
    n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
    n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
    n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
    n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
    n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
    n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
    n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
    n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
    n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582, n8584, n8585, n8586, n8587,
    n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
    n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
    n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
    n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
    n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
    n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
    n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
    n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
    n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
    n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
    n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
    n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
    n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
    n8808, n8809, n8810, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
    n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
    n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
    n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
    n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
    n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
    n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
    n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
    n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
    n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
    n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
    n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
    n9270, n9271, n9272, n9273, n9274, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
    n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
    n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9496, n9497, n9498, n9499, n9500, n9501,
    n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
    n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
    n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
    n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
    n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
    n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
    n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
    n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
    n9712, n9713, n9714, n9715, n9716, n9717, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
    n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
    n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
    n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
    n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
    n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
    n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
    n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9939, n9940, n9941, n9942, n9943,
    n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
    n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
    n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
    n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
    n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10143, n10144, n10145, n10146, n10147,
    n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
    n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
    n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
    n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
    n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
    n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
    n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
    n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
    n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
    n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
    n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
    n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
    n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
    n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
    n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
    n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
    n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
    n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
    n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
    n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
    n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
    n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
    n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
    n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
    n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
    n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
    n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
    n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
    n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
    n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
    n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
    n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
    n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
    n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
    n10744, n10745, n10746, n10747, n10748, n10749, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
    n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
    n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
    n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
    n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
    n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
    n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129, n11131, n11132, n11133,
    n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
    n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
    n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
    n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
    n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
    n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
    n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
    n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
    n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
    n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
    n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
    n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
    n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
    n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
    n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
    n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
    n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
    n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
    n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
    n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
    n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
    n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
    n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
    n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
    n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
    n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
    n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
    n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
    n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
    n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
    n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
    n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
    n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
    n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
    n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
    n11857, n11858, n11859, n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
    n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
    n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
    n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
    n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
    n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
    n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
    n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
    n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
    n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
    n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
    n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
    n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
    n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
    n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
    n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
    n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
    n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
    n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
    n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
    n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
    n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
    n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
    n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
    n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
    n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
    n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
    n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
    n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
    n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
    n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
    n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
    n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
    n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
    n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
    n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
    n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
    n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
    n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
    n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
    n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
    n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
    n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
    n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
    n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
    n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
    n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
    n13279, n13280, n13281, n13283, n13284, n13285, n13286, n13287, n13288,
    n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
    n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
    n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
    n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
    n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
    n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556, n13558, n13559, n13560,
    n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
    n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
    n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
    n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
    n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
    n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
    n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
    n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
    n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
    n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
    n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
    n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
    n13687, n13688, n13689, n13690, n13691, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
    n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
    n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
    n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
    n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13937, n13938, n13939, n13940, n13941,
    n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
    n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
    n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
    n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
    n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
    n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
    n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
    n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
    n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
    n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
    n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
    n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
    n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
    n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
    n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
    n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
    n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
    n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
    n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
    n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
    n14177, n14178, n14179, n14180, n14181, n14182, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
    n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
    n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
    n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
    n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
    n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
    n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
    n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
    n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
    n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
    n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
    n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
    n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
    n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
    n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14421, n14422,
    n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
    n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
    n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
    n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
    n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
    n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
    n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
    n14531, n14532, n14533, n14534, n14535, n14536, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
    n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
    n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
    n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
    n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
    n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
    n14640, n14641, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
    n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
    n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
    n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
    n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
    n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
    n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
    n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
    n14731, n14732, n14733, n14734, n14735, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
    n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
    n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
    n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
    n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
    n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
    n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
    n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
    n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
    n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
    n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
    n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
    n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
    n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
    n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
    n15095, n15096, n15097, n15098, n15099, n15100, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
    n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
    n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
    n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
    n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
    n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
    n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
    n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
    n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
    n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
    n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
    n15250, n15251, n15252, n15253, n15254, n15255, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
    n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
    n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
    n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
    n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
    n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
    n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
    n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
    n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
    n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
    n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
    n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
    n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
    n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
    n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
    n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
    n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
    n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
    n15524, n15525, n15526, n15527, n15528, n15530, n15531, n15532, n15533,
    n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
    n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
    n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
    n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
    n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
    n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
    n15625, n15626, n15627, n15628, n15629, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
    n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
    n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15723, n15724, n15725, n15726,
    n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
    n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
    n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
    n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15763,
    n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
    n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
    n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
    n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15808, n15809,
    n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
    n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15836, n15837,
    n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
    n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
    n15856, n15857, n15858, n15859, n15860, n15861, n15863, n15864, n15865,
    n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
    n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
    n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
    n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15908, n15909, n15910, n15911, n15912,
    n15913, n15914, n15915, n15916, n15917, n15918, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
    n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
    n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
    n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16241;
  zero g00000(.dout(\asquared[1] ));
  jnot g00001(.din(\a[0] ), .dout(n193));
  jand g00002(.dina(\a[1] ), .dinb(n193), .dout(\asquared[2] ));
  jand g00003(.dina(\a[2] ), .dinb(\a[1] ), .dout(n195));
  jnot g00004(.din(n195), .dout(n196));
  jor  g00005(.dina(\a[2] ), .dinb(\a[1] ), .dout(n197));
  jand g00006(.dina(n197), .dinb(\a[0] ), .dout(n198));
  jand g00007(.dina(n198), .dinb(n196), .dout(\asquared[3] ));
  jnot g00008(.din(\asquared[2] ), .dout(n200));
  jand g00009(.dina(\a[3] ), .dinb(\a[0] ), .dout(n201));
  jxor g00010(.dina(n201), .dinb(\a[2] ), .dout(n202));
  jand g00011(.dina(n202), .dinb(n200), .dout(\asquared[4] ));
  jand g00012(.dina(n201), .dinb(\a[2] ), .dout(n204));
  jnot g00013(.din(\a[3] ), .dout(n205));
  jor  g00014(.dina(n205), .dinb(n193), .dout(n206));
  jnot g00015(.din(\a[1] ), .dout(n207));
  jnot g00016(.din(\a[4] ), .dout(n208));
  jor  g00017(.dina(n208), .dinb(n207), .dout(n209));
  jor  g00018(.dina(n209), .dinb(n206), .dout(n210));
  jand g00019(.dina(\a[3] ), .dinb(\a[1] ), .dout(n211));
  jand g00020(.dina(\a[4] ), .dinb(\a[0] ), .dout(n212));
  jor  g00021(.dina(n212), .dinb(n211), .dout(n213));
  jand g00022(.dina(n213), .dinb(n210), .dout(n214));
  jxor g00023(.dina(n214), .dinb(n195), .dout(n215));
  jxor g00024(.dina(n215), .dinb(n204), .dout(\asquared[5] ));
  jnot g00025(.din(\a[2] ), .dout(n217));
  jand g00026(.dina(\a[3] ), .dinb(n217), .dout(n218));
  jnot g00027(.din(n218), .dout(n219));
  jand g00028(.dina(\a[4] ), .dinb(\a[1] ), .dout(n220));
  jand g00029(.dina(n220), .dinb(n201), .dout(n221));
  jand g00030(.dina(\a[5] ), .dinb(\a[0] ), .dout(n222));
  jor  g00031(.dina(n222), .dinb(n220), .dout(n223));
  jand g00032(.dina(\a[5] ), .dinb(\a[1] ), .dout(n224));
  jand g00033(.dina(n224), .dinb(n212), .dout(n225));
  jnot g00034(.din(n225), .dout(n226));
  jand g00035(.dina(n226), .dinb(n223), .dout(n227));
  jxor g00036(.dina(n227), .dinb(n221), .dout(n228));
  jxor g00037(.dina(n228), .dinb(n219), .dout(n229));
  jor  g00038(.dina(n205), .dinb(n207), .dout(n230));
  jor  g00039(.dina(n208), .dinb(n193), .dout(n231));
  jand g00040(.dina(n231), .dinb(n230), .dout(n232));
  jor  g00041(.dina(n232), .dinb(n221), .dout(n233));
  jor  g00042(.dina(n233), .dinb(n196), .dout(n234));
  jnot g00043(.din(n204), .dout(n235));
  jand g00044(.dina(n233), .dinb(n196), .dout(n236));
  jor  g00045(.dina(n236), .dinb(n235), .dout(n237));
  jand g00046(.dina(n237), .dinb(n234), .dout(n238));
  jxor g00047(.dina(n238), .dinb(n229), .dout(\asquared[6] ));
  jand g00048(.dina(n227), .dinb(n221), .dout(n240));
  jor  g00049(.dina(n240), .dinb(n225), .dout(n241));
  jand g00050(.dina(\a[5] ), .dinb(\a[4] ), .dout(n242));
  jand g00051(.dina(n242), .dinb(n195), .dout(n243));
  jnot g00052(.din(n243), .dout(n244));
  jand g00053(.dina(\a[4] ), .dinb(\a[2] ), .dout(n245));
  jor  g00054(.dina(n245), .dinb(n224), .dout(n246));
  jand g00055(.dina(n246), .dinb(n244), .dout(n247));
  jand g00056(.dina(\a[3] ), .dinb(\a[2] ), .dout(n248));
  jand g00057(.dina(\a[6] ), .dinb(\a[0] ), .dout(n249));
  jxor g00058(.dina(n249), .dinb(n248), .dout(n250));
  jxor g00059(.dina(n250), .dinb(n247), .dout(n251));
  jor  g00060(.dina(n251), .dinb(n241), .dout(n252));
  jnot g00061(.din(n252), .dout(n253));
  jand g00062(.dina(n251), .dinb(n241), .dout(n254));
  jor  g00063(.dina(n254), .dinb(n253), .dout(n255));
  jand g00064(.dina(n228), .dinb(n218), .dout(n256));
  jnot g00065(.din(n256), .dout(n257));
  jxor g00066(.dina(n227), .dinb(n210), .dout(n258));
  jand g00067(.dina(n258), .dinb(n219), .dout(n259));
  jor  g00068(.dina(n238), .dinb(n259), .dout(n260));
  jand g00069(.dina(n260), .dinb(n257), .dout(n261));
  jxor g00070(.dina(n261), .dinb(n255), .dout(\asquared[7] ));
  jand g00071(.dina(n242), .dinb(n248), .dout(n263));
  jnot g00072(.din(n263), .dout(n264));
  jand g00073(.dina(\a[4] ), .dinb(\a[3] ), .dout(n265));
  jand g00074(.dina(\a[7] ), .dinb(\a[0] ), .dout(n266));
  jand g00075(.dina(n266), .dinb(n265), .dout(n267));
  jand g00076(.dina(\a[7] ), .dinb(\a[2] ), .dout(n268));
  jand g00077(.dina(n268), .dinb(n222), .dout(n269));
  jor  g00078(.dina(n269), .dinb(n267), .dout(n270));
  jnot g00079(.din(n270), .dout(n271));
  jand g00080(.dina(n271), .dinb(n264), .dout(n272));
  jand g00081(.dina(\a[5] ), .dinb(\a[2] ), .dout(n273));
  jor  g00082(.dina(n273), .dinb(n265), .dout(n274));
  jand g00083(.dina(n274), .dinb(n272), .dout(n275));
  jand g00084(.dina(n270), .dinb(n264), .dout(n276));
  jnot g00085(.din(n276), .dout(n277));
  jand g00086(.dina(n277), .dinb(n266), .dout(n278));
  jor  g00087(.dina(n278), .dinb(n275), .dout(n279));
  jnot g00088(.din(n279), .dout(n280));
  jand g00089(.dina(n249), .dinb(n248), .dout(n281));
  jand g00090(.dina(n250), .dinb(n247), .dout(n282));
  jor  g00091(.dina(n282), .dinb(n281), .dout(n283));
  jnot g00092(.din(\a[6] ), .dout(n284));
  jand g00093(.dina(n243), .dinb(n284), .dout(n285));
  jnot g00094(.din(n285), .dout(n286));
  jand g00095(.dina(\a[6] ), .dinb(\a[1] ), .dout(n287));
  jxor g00096(.dina(n287), .dinb(\a[4] ), .dout(n288));
  jor  g00097(.dina(n288), .dinb(n243), .dout(n289));
  jand g00098(.dina(n289), .dinb(n286), .dout(n290));
  jxor g00099(.dina(n290), .dinb(n283), .dout(n291));
  jxor g00100(.dina(n291), .dinb(n280), .dout(n292));
  jnot g00101(.din(n254), .dout(n293));
  jor  g00102(.dina(n261), .dinb(n253), .dout(n294));
  jand g00103(.dina(n294), .dinb(n293), .dout(n295));
  jxor g00104(.dina(n295), .dinb(n292), .dout(\asquared[8] ));
  jand g00105(.dina(n290), .dinb(n283), .dout(n297));
  jor  g00106(.dina(n297), .dinb(n285), .dout(n298));
  jand g00107(.dina(n287), .dinb(\a[4] ), .dout(n299));
  jand g00108(.dina(\a[8] ), .dinb(\a[0] ), .dout(n300));
  jand g00109(.dina(\a[6] ), .dinb(\a[2] ), .dout(n301));
  jor  g00110(.dina(n301), .dinb(n300), .dout(n302));
  jand g00111(.dina(\a[8] ), .dinb(\a[2] ), .dout(n303));
  jand g00112(.dina(n303), .dinb(n249), .dout(n304));
  jnot g00113(.din(n304), .dout(n305));
  jand g00114(.dina(n305), .dinb(n302), .dout(n306));
  jxor g00115(.dina(n306), .dinb(n299), .dout(n307));
  jnot g00116(.din(n272), .dout(n308));
  jand g00117(.dina(\a[7] ), .dinb(\a[1] ), .dout(n309));
  jand g00118(.dina(\a[5] ), .dinb(\a[3] ), .dout(n310));
  jxor g00119(.dina(n310), .dinb(n309), .dout(n311));
  jxor g00120(.dina(n311), .dinb(n308), .dout(n312));
  jxor g00121(.dina(n312), .dinb(n307), .dout(n313));
  jor  g00122(.dina(n313), .dinb(n298), .dout(n314));
  jnot g00123(.din(n314), .dout(n315));
  jand g00124(.dina(n313), .dinb(n298), .dout(n316));
  jor  g00125(.dina(n316), .dinb(n315), .dout(n317));
  jand g00126(.dina(n291), .dinb(n279), .dout(n318));
  jnot g00127(.din(n318), .dout(n319));
  jnot g00128(.din(n291), .dout(n320));
  jand g00129(.dina(n320), .dinb(n280), .dout(n321));
  jor  g00130(.dina(n295), .dinb(n321), .dout(n322));
  jand g00131(.dina(n322), .dinb(n319), .dout(n323));
  jxor g00132(.dina(n323), .dinb(n317), .dout(\asquared[9] ));
  jand g00133(.dina(n311), .dinb(n308), .dout(n325));
  jand g00134(.dina(n312), .dinb(n307), .dout(n326));
  jor  g00135(.dina(n326), .dinb(n325), .dout(n327));
  jand g00136(.dina(n310), .dinb(n309), .dout(n328));
  jand g00137(.dina(\a[9] ), .dinb(\a[0] ), .dout(n329));
  jxor g00138(.dina(n329), .dinb(n328), .dout(n330));
  jand g00139(.dina(n224), .dinb(\a[8] ), .dout(n331));
  jnot g00140(.din(n331), .dout(n332));
  jand g00141(.dina(\a[8] ), .dinb(\a[1] ), .dout(n333));
  jor  g00142(.dina(n333), .dinb(\a[5] ), .dout(n334));
  jand g00143(.dina(n334), .dinb(n332), .dout(n335));
  jxor g00144(.dina(n335), .dinb(n330), .dout(n336));
  jand g00145(.dina(n306), .dinb(n299), .dout(n337));
  jor  g00146(.dina(n337), .dinb(n304), .dout(n338));
  jand g00147(.dina(\a[6] ), .dinb(\a[5] ), .dout(n339));
  jand g00148(.dina(n339), .dinb(n265), .dout(n340));
  jnot g00149(.din(n340), .dout(n341));
  jand g00150(.dina(\a[6] ), .dinb(\a[3] ), .dout(n342));
  jor  g00151(.dina(n342), .dinb(n242), .dout(n343));
  jand g00152(.dina(n343), .dinb(n341), .dout(n344));
  jxor g00153(.dina(n344), .dinb(n268), .dout(n345));
  jxor g00154(.dina(n345), .dinb(n338), .dout(n346));
  jxor g00155(.dina(n346), .dinb(n336), .dout(n347));
  jand g00156(.dina(n347), .dinb(n327), .dout(n348));
  jor  g00157(.dina(n347), .dinb(n327), .dout(n349));
  jnot g00158(.din(n349), .dout(n350));
  jor  g00159(.dina(n350), .dinb(n348), .dout(n351));
  jnot g00160(.din(n316), .dout(n352));
  jor  g00161(.dina(n323), .dinb(n315), .dout(n353));
  jand g00162(.dina(n353), .dinb(n352), .dout(n354));
  jxor g00163(.dina(n354), .dinb(n351), .dout(\asquared[10] ));
  jand g00164(.dina(n345), .dinb(n338), .dout(n356));
  jand g00165(.dina(n346), .dinb(n336), .dout(n357));
  jor  g00166(.dina(n357), .dinb(n356), .dout(n358));
  jand g00167(.dina(n344), .dinb(n268), .dout(n359));
  jor  g00168(.dina(n359), .dinb(n340), .dout(n360));
  jand g00169(.dina(\a[9] ), .dinb(\a[1] ), .dout(n361));
  jand g00170(.dina(\a[6] ), .dinb(\a[4] ), .dout(n362));
  jxor g00171(.dina(n362), .dinb(n361), .dout(n363));
  jxor g00172(.dina(n363), .dinb(n331), .dout(n364));
  jxor g00173(.dina(n364), .dinb(n360), .dout(n365));
  jand g00174(.dina(n329), .dinb(n328), .dout(n366));
  jand g00175(.dina(n335), .dinb(n330), .dout(n367));
  jor  g00176(.dina(n367), .dinb(n366), .dout(n368));
  jand g00177(.dina(\a[10] ), .dinb(\a[0] ), .dout(n369));
  jand g00178(.dina(\a[7] ), .dinb(\a[3] ), .dout(n370));
  jxor g00179(.dina(n370), .dinb(n369), .dout(n371));
  jxor g00180(.dina(n371), .dinb(n303), .dout(n372));
  jxor g00181(.dina(n372), .dinb(n368), .dout(n373));
  jxor g00182(.dina(n373), .dinb(n365), .dout(n374));
  jnot g00183(.din(n374), .dout(n375));
  jxor g00184(.dina(n375), .dinb(n358), .dout(n376));
  jnot g00185(.din(n348), .dout(n377));
  jor  g00186(.dina(n354), .dinb(n350), .dout(n378));
  jand g00187(.dina(n378), .dinb(n377), .dout(n379));
  jxor g00188(.dina(n379), .dinb(n376), .dout(\asquared[11] ));
  jand g00189(.dina(n372), .dinb(n368), .dout(n381));
  jand g00190(.dina(n373), .dinb(n365), .dout(n382));
  jor  g00191(.dina(n382), .dinb(n381), .dout(n383));
  jnot g00192(.din(n383), .dout(n384));
  jand g00193(.dina(n370), .dinb(n369), .dout(n385));
  jand g00194(.dina(n371), .dinb(n303), .dout(n386));
  jor  g00195(.dina(n386), .dinb(n385), .dout(n387));
  jand g00196(.dina(n287), .dinb(\a[10] ), .dout(n388));
  jnot g00197(.din(n388), .dout(n389));
  jand g00198(.dina(\a[10] ), .dinb(\a[1] ), .dout(n390));
  jor  g00199(.dina(n390), .dinb(\a[6] ), .dout(n391));
  jand g00200(.dina(n391), .dinb(n389), .dout(n392));
  jxor g00201(.dina(n392), .dinb(n387), .dout(n393));
  jand g00202(.dina(n362), .dinb(n361), .dout(n394));
  jand g00203(.dina(\a[9] ), .dinb(\a[8] ), .dout(n395));
  jand g00204(.dina(n395), .dinb(n248), .dout(n396));
  jnot g00205(.din(n396), .dout(n397));
  jand g00206(.dina(\a[9] ), .dinb(\a[2] ), .dout(n398));
  jand g00207(.dina(\a[8] ), .dinb(\a[3] ), .dout(n399));
  jor  g00208(.dina(n399), .dinb(n398), .dout(n400));
  jand g00209(.dina(n400), .dinb(n397), .dout(n401));
  jxor g00210(.dina(n401), .dinb(n394), .dout(n402));
  jxor g00211(.dina(n402), .dinb(n393), .dout(n403));
  jand g00212(.dina(n363), .dinb(n331), .dout(n404));
  jand g00213(.dina(n364), .dinb(n360), .dout(n405));
  jor  g00214(.dina(n405), .dinb(n404), .dout(n406));
  jand g00215(.dina(\a[11] ), .dinb(\a[0] ), .dout(n407));
  jand g00216(.dina(\a[7] ), .dinb(\a[4] ), .dout(n408));
  jor  g00217(.dina(n408), .dinb(n339), .dout(n409));
  jand g00218(.dina(\a[7] ), .dinb(\a[6] ), .dout(n410));
  jand g00219(.dina(n410), .dinb(n242), .dout(n411));
  jnot g00220(.din(n411), .dout(n412));
  jand g00221(.dina(n412), .dinb(n409), .dout(n413));
  jxor g00222(.dina(n413), .dinb(n407), .dout(n414));
  jxor g00223(.dina(n414), .dinb(n406), .dout(n415));
  jxor g00224(.dina(n415), .dinb(n403), .dout(n416));
  jxor g00225(.dina(n416), .dinb(n384), .dout(n417));
  jand g00226(.dina(n374), .dinb(n358), .dout(n418));
  jnot g00227(.din(n418), .dout(n419));
  jnot g00228(.din(n358), .dout(n420));
  jand g00229(.dina(n375), .dinb(n420), .dout(n421));
  jor  g00230(.dina(n379), .dinb(n421), .dout(n422));
  jand g00231(.dina(n422), .dinb(n419), .dout(n423));
  jxor g00232(.dina(n423), .dinb(n417), .dout(\asquared[12] ));
  jand g00233(.dina(n414), .dinb(n406), .dout(n425));
  jand g00234(.dina(n415), .dinb(n403), .dout(n426));
  jor  g00235(.dina(n426), .dinb(n425), .dout(n427));
  jand g00236(.dina(n392), .dinb(n387), .dout(n428));
  jand g00237(.dina(n402), .dinb(n393), .dout(n429));
  jor  g00238(.dina(n429), .dinb(n428), .dout(n430));
  jand g00239(.dina(\a[7] ), .dinb(\a[5] ), .dout(n431));
  jand g00240(.dina(\a[11] ), .dinb(\a[1] ), .dout(n432));
  jxor g00241(.dina(n432), .dinb(n431), .dout(n433));
  jand g00242(.dina(\a[8] ), .dinb(\a[4] ), .dout(n434));
  jor  g00243(.dina(n434), .dinb(n388), .dout(n435));
  jand g00244(.dina(\a[10] ), .dinb(\a[8] ), .dout(n436));
  jand g00245(.dina(n436), .dinb(n299), .dout(n437));
  jnot g00246(.din(n437), .dout(n438));
  jand g00247(.dina(n438), .dinb(n435), .dout(n439));
  jxor g00248(.dina(n439), .dinb(n433), .dout(n440));
  jxor g00249(.dina(n440), .dinb(n430), .dout(n441));
  jand g00250(.dina(n401), .dinb(n394), .dout(n442));
  jor  g00251(.dina(n442), .dinb(n396), .dout(n443));
  jand g00252(.dina(n413), .dinb(n407), .dout(n444));
  jor  g00253(.dina(n444), .dinb(n411), .dout(n445));
  jxor g00254(.dina(n445), .dinb(n443), .dout(n446));
  jand g00255(.dina(\a[9] ), .dinb(\a[3] ), .dout(n447));
  jand g00256(.dina(\a[12] ), .dinb(\a[2] ), .dout(n448));
  jand g00257(.dina(n448), .dinb(n369), .dout(n449));
  jnot g00258(.din(n449), .dout(n450));
  jand g00259(.dina(\a[12] ), .dinb(\a[0] ), .dout(n451));
  jand g00260(.dina(n451), .dinb(n447), .dout(n452));
  jand g00261(.dina(\a[10] ), .dinb(\a[9] ), .dout(n453));
  jand g00262(.dina(n453), .dinb(n248), .dout(n454));
  jor  g00263(.dina(n454), .dinb(n452), .dout(n455));
  jand g00264(.dina(n455), .dinb(n450), .dout(n456));
  jnot g00265(.din(n456), .dout(n457));
  jand g00266(.dina(n457), .dinb(n447), .dout(n458));
  jor  g00267(.dina(n455), .dinb(n449), .dout(n459));
  jnot g00268(.din(n459), .dout(n460));
  jand g00269(.dina(\a[10] ), .dinb(\a[2] ), .dout(n461));
  jor  g00270(.dina(n461), .dinb(n451), .dout(n462));
  jand g00271(.dina(n462), .dinb(n460), .dout(n463));
  jor  g00272(.dina(n463), .dinb(n458), .dout(n464));
  jxor g00273(.dina(n464), .dinb(n446), .dout(n465));
  jxor g00274(.dina(n465), .dinb(n441), .dout(n466));
  jnot g00275(.din(n466), .dout(n467));
  jxor g00276(.dina(n467), .dinb(n427), .dout(n468));
  jand g00277(.dina(n416), .dinb(n383), .dout(n469));
  jnot g00278(.din(n469), .dout(n470));
  jnot g00279(.din(n416), .dout(n471));
  jand g00280(.dina(n471), .dinb(n384), .dout(n472));
  jor  g00281(.dina(n423), .dinb(n472), .dout(n473));
  jand g00282(.dina(n473), .dinb(n470), .dout(n474));
  jxor g00283(.dina(n474), .dinb(n468), .dout(\asquared[13] ));
  jand g00284(.dina(n439), .dinb(n433), .dout(n476));
  jor  g00285(.dina(n476), .dinb(n437), .dout(n477));
  jand g00286(.dina(\a[10] ), .dinb(\a[3] ), .dout(n478));
  jand g00287(.dina(\a[13] ), .dinb(\a[9] ), .dout(n479));
  jand g00288(.dina(n479), .dinb(n212), .dout(n480));
  jnot g00289(.din(n480), .dout(n481));
  jand g00290(.dina(n453), .dinb(n265), .dout(n482));
  jand g00291(.dina(\a[13] ), .dinb(\a[0] ), .dout(n483));
  jand g00292(.dina(n483), .dinb(n478), .dout(n484));
  jor  g00293(.dina(n484), .dinb(n482), .dout(n485));
  jand g00294(.dina(n485), .dinb(n481), .dout(n486));
  jnot g00295(.din(n486), .dout(n487));
  jand g00296(.dina(n487), .dinb(n478), .dout(n488));
  jor  g00297(.dina(n485), .dinb(n480), .dout(n489));
  jnot g00298(.din(n489), .dout(n490));
  jand g00299(.dina(\a[9] ), .dinb(\a[4] ), .dout(n491));
  jor  g00300(.dina(n491), .dinb(n483), .dout(n492));
  jand g00301(.dina(n492), .dinb(n490), .dout(n493));
  jor  g00302(.dina(n493), .dinb(n488), .dout(n494));
  jxor g00303(.dina(n494), .dinb(n477), .dout(n495));
  jnot g00304(.din(n495), .dout(n496));
  jand g00305(.dina(\a[11] ), .dinb(\a[2] ), .dout(n497));
  jnot g00306(.din(n497), .dout(n498));
  jand g00307(.dina(\a[8] ), .dinb(\a[7] ), .dout(n499));
  jand g00308(.dina(n499), .dinb(n339), .dout(n500));
  jnot g00309(.din(n500), .dout(n501));
  jand g00310(.dina(\a[8] ), .dinb(\a[5] ), .dout(n502));
  jor  g00311(.dina(n502), .dinb(n410), .dout(n503));
  jand g00312(.dina(n503), .dinb(n501), .dout(n504));
  jxor g00313(.dina(n504), .dinb(n498), .dout(n505));
  jxor g00314(.dina(n505), .dinb(n496), .dout(n506));
  jnot g00315(.din(n506), .dout(n507));
  jand g00316(.dina(n445), .dinb(n443), .dout(n508));
  jand g00317(.dina(n464), .dinb(n446), .dout(n509));
  jor  g00318(.dina(n509), .dinb(n508), .dout(n510));
  jnot g00319(.din(\a[12] ), .dout(n511));
  jand g00320(.dina(n432), .dinb(n431), .dout(n512));
  jand g00321(.dina(n512), .dinb(n511), .dout(n513));
  jnot g00322(.din(n513), .dout(n514));
  jand g00323(.dina(n309), .dinb(\a[12] ), .dout(n515));
  jnot g00324(.din(n515), .dout(n516));
  jand g00325(.dina(\a[12] ), .dinb(\a[1] ), .dout(n517));
  jor  g00326(.dina(n517), .dinb(\a[7] ), .dout(n518));
  jand g00327(.dina(n518), .dinb(n516), .dout(n519));
  jor  g00328(.dina(n519), .dinb(n512), .dout(n520));
  jand g00329(.dina(n520), .dinb(n514), .dout(n521));
  jxor g00330(.dina(n521), .dinb(n459), .dout(n522));
  jxor g00331(.dina(n522), .dinb(n510), .dout(n523));
  jand g00332(.dina(n440), .dinb(n430), .dout(n524));
  jand g00333(.dina(n465), .dinb(n441), .dout(n525));
  jor  g00334(.dina(n525), .dinb(n524), .dout(n526));
  jxor g00335(.dina(n526), .dinb(n523), .dout(n527));
  jxor g00336(.dina(n527), .dinb(n507), .dout(n528));
  jand g00337(.dina(n466), .dinb(n427), .dout(n529));
  jnot g00338(.din(n529), .dout(n530));
  jnot g00339(.din(n427), .dout(n531));
  jand g00340(.dina(n467), .dinb(n531), .dout(n532));
  jor  g00341(.dina(n474), .dinb(n532), .dout(n533));
  jand g00342(.dina(n533), .dinb(n530), .dout(n534));
  jxor g00343(.dina(n534), .dinb(n528), .dout(\asquared[14] ));
  jand g00344(.dina(n522), .dinb(n510), .dout(n536));
  jand g00345(.dina(n526), .dinb(n523), .dout(n537));
  jor  g00346(.dina(n537), .dinb(n536), .dout(n538));
  jand g00347(.dina(n494), .dinb(n477), .dout(n539));
  jnot g00348(.din(n539), .dout(n540));
  jor  g00349(.dina(n505), .dinb(n496), .dout(n541));
  jand g00350(.dina(n541), .dinb(n540), .dout(n542));
  jnot g00351(.din(n542), .dout(n543));
  jand g00352(.dina(\a[8] ), .dinb(\a[6] ), .dout(n544));
  jand g00353(.dina(\a[13] ), .dinb(\a[1] ), .dout(n545));
  jxor g00354(.dina(n545), .dinb(n544), .dout(n546));
  jand g00355(.dina(n501), .dinb(n498), .dout(n547));
  jnot g00356(.din(n547), .dout(n548));
  jand g00357(.dina(n548), .dinb(n503), .dout(n549));
  jxor g00358(.dina(n549), .dinb(n546), .dout(n550));
  jxor g00359(.dina(n550), .dinb(n489), .dout(n551));
  jxor g00360(.dina(n551), .dinb(n543), .dout(n552));
  jand g00361(.dina(n521), .dinb(n459), .dout(n553));
  jor  g00362(.dina(n553), .dinb(n513), .dout(n554));
  jand g00363(.dina(\a[12] ), .dinb(\a[11] ), .dout(n555));
  jand g00364(.dina(n555), .dinb(n248), .dout(n556));
  jnot g00365(.din(n556), .dout(n557));
  jand g00366(.dina(\a[11] ), .dinb(\a[3] ), .dout(n558));
  jand g00367(.dina(\a[14] ), .dinb(\a[0] ), .dout(n559));
  jand g00368(.dina(n559), .dinb(n558), .dout(n560));
  jand g00369(.dina(\a[14] ), .dinb(\a[2] ), .dout(n561));
  jand g00370(.dina(n561), .dinb(n451), .dout(n562));
  jor  g00371(.dina(n562), .dinb(n560), .dout(n563));
  jnot g00372(.din(n563), .dout(n564));
  jand g00373(.dina(n564), .dinb(n557), .dout(n565));
  jor  g00374(.dina(n558), .dinb(n448), .dout(n566));
  jand g00375(.dina(n566), .dinb(n565), .dout(n567));
  jand g00376(.dina(n563), .dinb(n557), .dout(n568));
  jnot g00377(.din(n568), .dout(n569));
  jand g00378(.dina(n569), .dinb(n559), .dout(n570));
  jor  g00379(.dina(n570), .dinb(n567), .dout(n571));
  jand g00380(.dina(n453), .dinb(n242), .dout(n572));
  jnot g00381(.din(n572), .dout(n573));
  jand g00382(.dina(\a[10] ), .dinb(\a[4] ), .dout(n574));
  jand g00383(.dina(\a[9] ), .dinb(\a[5] ), .dout(n575));
  jor  g00384(.dina(n575), .dinb(n574), .dout(n576));
  jand g00385(.dina(n576), .dinb(n573), .dout(n577));
  jxor g00386(.dina(n577), .dinb(n515), .dout(n578));
  jxor g00387(.dina(n578), .dinb(n571), .dout(n579));
  jxor g00388(.dina(n579), .dinb(n554), .dout(n580));
  jxor g00389(.dina(n580), .dinb(n552), .dout(n581));
  jand g00390(.dina(n581), .dinb(n538), .dout(n582));
  jor  g00391(.dina(n581), .dinb(n538), .dout(n583));
  jnot g00392(.din(n583), .dout(n584));
  jor  g00393(.dina(n584), .dinb(n582), .dout(n585));
  jand g00394(.dina(n527), .dinb(n506), .dout(n586));
  jnot g00395(.din(n586), .dout(n587));
  jnot g00396(.din(n527), .dout(n588));
  jand g00397(.dina(n588), .dinb(n507), .dout(n589));
  jor  g00398(.dina(n534), .dinb(n589), .dout(n590));
  jand g00399(.dina(n590), .dinb(n587), .dout(n591));
  jxor g00400(.dina(n591), .dinb(n585), .dout(\asquared[15] ));
  jand g00401(.dina(n551), .dinb(n543), .dout(n593));
  jand g00402(.dina(n580), .dinb(n552), .dout(n594));
  jor  g00403(.dina(n594), .dinb(n593), .dout(n595));
  jand g00404(.dina(n549), .dinb(n546), .dout(n596));
  jand g00405(.dina(n550), .dinb(n489), .dout(n597));
  jor  g00406(.dina(n597), .dinb(n596), .dout(n598));
  jand g00407(.dina(\a[14] ), .dinb(\a[1] ), .dout(n599));
  jxor g00408(.dina(n599), .dinb(\a[8] ), .dout(n600));
  jand g00409(.dina(n545), .dinb(n544), .dout(n601));
  jand g00410(.dina(\a[11] ), .dinb(\a[4] ), .dout(n602));
  jxor g00411(.dina(n602), .dinb(n601), .dout(n603));
  jxor g00412(.dina(n603), .dinb(n600), .dout(n604));
  jand g00413(.dina(\a[13] ), .dinb(\a[2] ), .dout(n605));
  jand g00414(.dina(\a[9] ), .dinb(\a[6] ), .dout(n606));
  jxor g00415(.dina(n606), .dinb(n499), .dout(n607));
  jxor g00416(.dina(n607), .dinb(n605), .dout(n608));
  jxor g00417(.dina(n608), .dinb(n604), .dout(n609));
  jxor g00418(.dina(n609), .dinb(n598), .dout(n610));
  jand g00419(.dina(n578), .dinb(n571), .dout(n611));
  jand g00420(.dina(n579), .dinb(n554), .dout(n612));
  jor  g00421(.dina(n612), .dinb(n611), .dout(n613));
  jnot g00422(.din(n565), .dout(n614));
  jand g00423(.dina(n577), .dinb(n515), .dout(n615));
  jor  g00424(.dina(n615), .dinb(n572), .dout(n616));
  jxor g00425(.dina(n616), .dinb(n614), .dout(n617));
  jnot g00426(.din(n617), .dout(n618));
  jand g00427(.dina(\a[10] ), .dinb(\a[5] ), .dout(n619));
  jnot g00428(.din(n619), .dout(n620));
  jand g00429(.dina(\a[15] ), .dinb(\a[0] ), .dout(n621));
  jand g00430(.dina(\a[12] ), .dinb(\a[3] ), .dout(n622));
  jxor g00431(.dina(n622), .dinb(n621), .dout(n623));
  jxor g00432(.dina(n623), .dinb(n620), .dout(n624));
  jxor g00433(.dina(n624), .dinb(n618), .dout(n625));
  jxor g00434(.dina(n625), .dinb(n613), .dout(n626));
  jxor g00435(.dina(n626), .dinb(n610), .dout(n627));
  jand g00436(.dina(n627), .dinb(n595), .dout(n628));
  jor  g00437(.dina(n627), .dinb(n595), .dout(n629));
  jnot g00438(.din(n629), .dout(n630));
  jor  g00439(.dina(n630), .dinb(n628), .dout(n631));
  jnot g00440(.din(n582), .dout(n632));
  jor  g00441(.dina(n591), .dinb(n584), .dout(n633));
  jand g00442(.dina(n633), .dinb(n632), .dout(n634));
  jxor g00443(.dina(n634), .dinb(n631), .dout(\asquared[16] ));
  jand g00444(.dina(n625), .dinb(n613), .dout(n636));
  jand g00445(.dina(n626), .dinb(n610), .dout(n637));
  jor  g00446(.dina(n637), .dinb(n636), .dout(n638));
  jand g00447(.dina(n608), .dinb(n604), .dout(n639));
  jand g00448(.dina(n609), .dinb(n598), .dout(n640));
  jor  g00449(.dina(n640), .dinb(n639), .dout(n641));
  jand g00450(.dina(n602), .dinb(n601), .dout(n642));
  jand g00451(.dina(n603), .dinb(n600), .dout(n643));
  jor  g00452(.dina(n643), .dinb(n642), .dout(n644));
  jor  g00453(.dina(n622), .dinb(n621), .dout(n645));
  jand g00454(.dina(n622), .dinb(n621), .dout(n646));
  jor  g00455(.dina(n646), .dinb(n619), .dout(n647));
  jand g00456(.dina(n647), .dinb(n645), .dout(n648));
  jxor g00457(.dina(n648), .dinb(n644), .dout(n649));
  jand g00458(.dina(\a[11] ), .dinb(\a[5] ), .dout(n650));
  jand g00459(.dina(\a[10] ), .dinb(\a[6] ), .dout(n651));
  jand g00460(.dina(\a[16] ), .dinb(\a[0] ), .dout(n652));
  jand g00461(.dina(n652), .dinb(n651), .dout(n653));
  jnot g00462(.din(n653), .dout(n654));
  jand g00463(.dina(\a[11] ), .dinb(\a[10] ), .dout(n655));
  jand g00464(.dina(n655), .dinb(n339), .dout(n656));
  jand g00465(.dina(n652), .dinb(n650), .dout(n657));
  jor  g00466(.dina(n657), .dinb(n656), .dout(n658));
  jand g00467(.dina(n658), .dinb(n654), .dout(n659));
  jnot g00468(.din(n659), .dout(n660));
  jand g00469(.dina(n660), .dinb(n650), .dout(n661));
  jor  g00470(.dina(n658), .dinb(n653), .dout(n662));
  jnot g00471(.din(n662), .dout(n663));
  jor  g00472(.dina(n652), .dinb(n651), .dout(n664));
  jand g00473(.dina(n664), .dinb(n663), .dout(n665));
  jor  g00474(.dina(n665), .dinb(n661), .dout(n666));
  jxor g00475(.dina(n666), .dinb(n649), .dout(n667));
  jxor g00476(.dina(n667), .dinb(n641), .dout(n668));
  jand g00477(.dina(n616), .dinb(n614), .dout(n669));
  jnot g00478(.din(n669), .dout(n670));
  jor  g00479(.dina(n624), .dinb(n618), .dout(n671));
  jand g00480(.dina(n671), .dinb(n670), .dout(n672));
  jnot g00481(.din(n672), .dout(n673));
  jand g00482(.dina(\a[12] ), .dinb(\a[4] ), .dout(n674));
  jand g00483(.dina(\a[14] ), .dinb(\a[13] ), .dout(n675));
  jand g00484(.dina(n675), .dinb(n248), .dout(n676));
  jnot g00485(.din(n676), .dout(n677));
  jand g00486(.dina(\a[13] ), .dinb(\a[3] ), .dout(n678));
  jor  g00487(.dina(n678), .dinb(n561), .dout(n679));
  jand g00488(.dina(n679), .dinb(n677), .dout(n680));
  jxor g00489(.dina(n680), .dinb(n674), .dout(n681));
  jxor g00490(.dina(n681), .dinb(n673), .dout(n682));
  jand g00491(.dina(n599), .dinb(\a[8] ), .dout(n683));
  jand g00492(.dina(\a[9] ), .dinb(\a[7] ), .dout(n684));
  jand g00493(.dina(\a[15] ), .dinb(\a[1] ), .dout(n685));
  jxor g00494(.dina(n685), .dinb(n684), .dout(n686));
  jxor g00495(.dina(n686), .dinb(n683), .dout(n687));
  jor  g00496(.dina(n606), .dinb(n499), .dout(n688));
  jand g00497(.dina(n606), .dinb(n499), .dout(n689));
  jor  g00498(.dina(n689), .dinb(n605), .dout(n690));
  jand g00499(.dina(n690), .dinb(n688), .dout(n691));
  jxor g00500(.dina(n691), .dinb(n687), .dout(n692));
  jxor g00501(.dina(n692), .dinb(n682), .dout(n693));
  jxor g00502(.dina(n693), .dinb(n668), .dout(n694));
  jand g00503(.dina(n694), .dinb(n638), .dout(n695));
  jor  g00504(.dina(n694), .dinb(n638), .dout(n696));
  jnot g00505(.din(n696), .dout(n697));
  jor  g00506(.dina(n697), .dinb(n695), .dout(n698));
  jnot g00507(.din(n628), .dout(n699));
  jor  g00508(.dina(n634), .dinb(n630), .dout(n700));
  jand g00509(.dina(n700), .dinb(n699), .dout(n701));
  jxor g00510(.dina(n701), .dinb(n698), .dout(\asquared[17] ));
  jand g00511(.dina(n667), .dinb(n641), .dout(n703));
  jand g00512(.dina(n693), .dinb(n668), .dout(n704));
  jor  g00513(.dina(n704), .dinb(n703), .dout(n705));
  jand g00514(.dina(n681), .dinb(n673), .dout(n706));
  jand g00515(.dina(n692), .dinb(n682), .dout(n707));
  jor  g00516(.dina(n707), .dinb(n706), .dout(n708));
  jand g00517(.dina(n685), .dinb(n684), .dout(n709));
  jand g00518(.dina(\a[12] ), .dinb(\a[5] ), .dout(n710));
  jand g00519(.dina(\a[17] ), .dinb(\a[0] ), .dout(n711));
  jnot g00520(.din(n711), .dout(n712));
  jxor g00521(.dina(n712), .dinb(n710), .dout(n713));
  jxor g00522(.dina(n713), .dinb(n709), .dout(n714));
  jand g00523(.dina(\a[14] ), .dinb(\a[3] ), .dout(n715));
  jnot g00524(.din(n715), .dout(n716));
  jand g00525(.dina(n499), .dinb(n453), .dout(n717));
  jnot g00526(.din(n717), .dout(n718));
  jand g00527(.dina(\a[10] ), .dinb(\a[7] ), .dout(n719));
  jor  g00528(.dina(n719), .dinb(n395), .dout(n720));
  jand g00529(.dina(n720), .dinb(n718), .dout(n721));
  jxor g00530(.dina(n721), .dinb(n716), .dout(n722));
  jxor g00531(.dina(n722), .dinb(n714), .dout(n723));
  jnot g00532(.din(n723), .dout(n724));
  jand g00533(.dina(\a[11] ), .dinb(\a[6] ), .dout(n725));
  jnot g00534(.din(n725), .dout(n726));
  jand g00535(.dina(\a[15] ), .dinb(\a[13] ), .dout(n727));
  jand g00536(.dina(n727), .dinb(n245), .dout(n728));
  jnot g00537(.din(n728), .dout(n729));
  jand g00538(.dina(\a[15] ), .dinb(\a[2] ), .dout(n730));
  jand g00539(.dina(\a[13] ), .dinb(\a[4] ), .dout(n731));
  jor  g00540(.dina(n731), .dinb(n730), .dout(n732));
  jand g00541(.dina(n732), .dinb(n729), .dout(n733));
  jxor g00542(.dina(n733), .dinb(n726), .dout(n734));
  jxor g00543(.dina(n734), .dinb(n724), .dout(n735));
  jxor g00544(.dina(n735), .dinb(n708), .dout(n736));
  jand g00545(.dina(n686), .dinb(n683), .dout(n737));
  jand g00546(.dina(n691), .dinb(n687), .dout(n738));
  jor  g00547(.dina(n738), .dinb(n737), .dout(n739));
  jand g00548(.dina(n648), .dinb(n644), .dout(n740));
  jand g00549(.dina(n666), .dinb(n649), .dout(n741));
  jor  g00550(.dina(n741), .dinb(n740), .dout(n742));
  jxor g00551(.dina(n742), .dinb(n739), .dout(n743));
  jand g00552(.dina(\a[16] ), .dinb(\a[1] ), .dout(n744));
  jor  g00553(.dina(n744), .dinb(\a[9] ), .dout(n745));
  jand g00554(.dina(n361), .dinb(\a[16] ), .dout(n746));
  jnot g00555(.din(n746), .dout(n747));
  jand g00556(.dina(n747), .dinb(n745), .dout(n748));
  jnot g00557(.din(n674), .dout(n749));
  jand g00558(.dina(n677), .dinb(n749), .dout(n750));
  jnot g00559(.din(n750), .dout(n751));
  jand g00560(.dina(n751), .dinb(n679), .dout(n752));
  jxor g00561(.dina(n752), .dinb(n748), .dout(n753));
  jxor g00562(.dina(n753), .dinb(n662), .dout(n754));
  jxor g00563(.dina(n754), .dinb(n743), .dout(n755));
  jxor g00564(.dina(n755), .dinb(n736), .dout(n756));
  jand g00565(.dina(n756), .dinb(n705), .dout(n757));
  jor  g00566(.dina(n756), .dinb(n705), .dout(n758));
  jnot g00567(.din(n758), .dout(n759));
  jor  g00568(.dina(n759), .dinb(n757), .dout(n760));
  jnot g00569(.din(n695), .dout(n761));
  jor  g00570(.dina(n701), .dinb(n697), .dout(n762));
  jand g00571(.dina(n762), .dinb(n761), .dout(n763));
  jxor g00572(.dina(n763), .dinb(n760), .dout(\asquared[18] ));
  jand g00573(.dina(n735), .dinb(n708), .dout(n765));
  jand g00574(.dina(n755), .dinb(n736), .dout(n766));
  jor  g00575(.dina(n766), .dinb(n765), .dout(n767));
  jand g00576(.dina(n729), .dinb(n726), .dout(n768));
  jnot g00577(.din(n768), .dout(n769));
  jand g00578(.dina(n769), .dinb(n732), .dout(n770));
  jand g00579(.dina(n718), .dinb(n716), .dout(n771));
  jnot g00580(.din(n771), .dout(n772));
  jand g00581(.dina(n772), .dinb(n720), .dout(n773));
  jxor g00582(.dina(n773), .dinb(n770), .dout(n774));
  jnot g00583(.din(n710), .dout(n775));
  jand g00584(.dina(n712), .dinb(n775), .dout(n776));
  jnot g00585(.din(n776), .dout(n777));
  jand g00586(.dina(n711), .dinb(n710), .dout(n778));
  jor  g00587(.dina(n778), .dinb(n709), .dout(n779));
  jand g00588(.dina(n779), .dinb(n777), .dout(n780));
  jxor g00589(.dina(n780), .dinb(n774), .dout(n781));
  jand g00590(.dina(n752), .dinb(n748), .dout(n782));
  jand g00591(.dina(n753), .dinb(n662), .dout(n783));
  jor  g00592(.dina(n783), .dinb(n782), .dout(n784));
  jnot g00593(.din(n784), .dout(n785));
  jor  g00594(.dina(n722), .dinb(n714), .dout(n786));
  jor  g00595(.dina(n734), .dinb(n724), .dout(n787));
  jand g00596(.dina(n787), .dinb(n786), .dout(n788));
  jxor g00597(.dina(n788), .dinb(n785), .dout(n789));
  jxor g00598(.dina(n789), .dinb(n781), .dout(n790));
  jand g00599(.dina(n742), .dinb(n739), .dout(n791));
  jand g00600(.dina(n754), .dinb(n743), .dout(n792));
  jor  g00601(.dina(n792), .dinb(n791), .dout(n793));
  jand g00602(.dina(\a[17] ), .dinb(\a[1] ), .dout(n794));
  jxor g00603(.dina(n794), .dinb(n436), .dout(n795));
  jnot g00604(.din(n795), .dout(n796));
  jand g00605(.dina(\a[12] ), .dinb(\a[6] ), .dout(n797));
  jxor g00606(.dina(n797), .dinb(n746), .dout(n798));
  jor  g00607(.dina(n798), .dinb(n796), .dout(n799));
  jnot g00608(.din(n797), .dout(n800));
  jand g00609(.dina(n800), .dinb(n747), .dout(n801));
  jnot g00610(.din(n801), .dout(n802));
  jand g00611(.dina(n797), .dinb(n746), .dout(n803));
  jor  g00612(.dina(n803), .dinb(n795), .dout(n804));
  jnot g00613(.din(n804), .dout(n805));
  jand g00614(.dina(n805), .dinb(n802), .dout(n806));
  jnot g00615(.din(n806), .dout(n807));
  jand g00616(.dina(n807), .dinb(n799), .dout(n808));
  jnot g00617(.din(n808), .dout(n809));
  jand g00618(.dina(\a[13] ), .dinb(\a[5] ), .dout(n810));
  jand g00619(.dina(\a[18] ), .dinb(\a[0] ), .dout(n811));
  jand g00620(.dina(n811), .dinb(n810), .dout(n812));
  jnot g00621(.din(n812), .dout(n813));
  jand g00622(.dina(\a[11] ), .dinb(\a[7] ), .dout(n814));
  jand g00623(.dina(n814), .dinb(n811), .dout(n815));
  jand g00624(.dina(\a[13] ), .dinb(\a[11] ), .dout(n816));
  jand g00625(.dina(n816), .dinb(n431), .dout(n817));
  jor  g00626(.dina(n817), .dinb(n815), .dout(n818));
  jnot g00627(.din(n818), .dout(n819));
  jand g00628(.dina(n819), .dinb(n813), .dout(n820));
  jor  g00629(.dina(n811), .dinb(n810), .dout(n821));
  jand g00630(.dina(n821), .dinb(n820), .dout(n822));
  jand g00631(.dina(n818), .dinb(n813), .dout(n823));
  jnot g00632(.din(n823), .dout(n824));
  jand g00633(.dina(n824), .dinb(n814), .dout(n825));
  jor  g00634(.dina(n825), .dinb(n822), .dout(n826));
  jand g00635(.dina(\a[14] ), .dinb(\a[4] ), .dout(n827));
  jnot g00636(.din(n827), .dout(n828));
  jand g00637(.dina(\a[16] ), .dinb(\a[15] ), .dout(n829));
  jand g00638(.dina(n829), .dinb(n248), .dout(n830));
  jnot g00639(.din(n830), .dout(n831));
  jand g00640(.dina(\a[15] ), .dinb(\a[3] ), .dout(n832));
  jand g00641(.dina(\a[16] ), .dinb(\a[2] ), .dout(n833));
  jor  g00642(.dina(n833), .dinb(n832), .dout(n834));
  jand g00643(.dina(n834), .dinb(n831), .dout(n835));
  jxor g00644(.dina(n835), .dinb(n828), .dout(n836));
  jnot g00645(.din(n836), .dout(n837));
  jxor g00646(.dina(n837), .dinb(n826), .dout(n838));
  jxor g00647(.dina(n838), .dinb(n809), .dout(n839));
  jxor g00648(.dina(n839), .dinb(n793), .dout(n840));
  jxor g00649(.dina(n840), .dinb(n790), .dout(n841));
  jand g00650(.dina(n841), .dinb(n767), .dout(n842));
  jor  g00651(.dina(n841), .dinb(n767), .dout(n843));
  jnot g00652(.din(n843), .dout(n844));
  jor  g00653(.dina(n844), .dinb(n842), .dout(n845));
  jnot g00654(.din(n757), .dout(n846));
  jor  g00655(.dina(n763), .dinb(n759), .dout(n847));
  jand g00656(.dina(n847), .dinb(n846), .dout(n848));
  jxor g00657(.dina(n848), .dinb(n845), .dout(\asquared[19] ));
  jand g00658(.dina(n837), .dinb(n826), .dout(n850));
  jand g00659(.dina(n838), .dinb(n809), .dout(n851));
  jor  g00660(.dina(n851), .dinb(n850), .dout(n852));
  jnot g00661(.din(\a[18] ), .dout(n853));
  jand g00662(.dina(n794), .dinb(n436), .dout(n854));
  jand g00663(.dina(n854), .dinb(n853), .dout(n855));
  jnot g00664(.din(n855), .dout(n856));
  jand g00665(.dina(\a[18] ), .dinb(\a[1] ), .dout(n857));
  jxor g00666(.dina(n857), .dinb(\a[10] ), .dout(n858));
  jor  g00667(.dina(n858), .dinb(n854), .dout(n859));
  jand g00668(.dina(n859), .dinb(n856), .dout(n860));
  jand g00669(.dina(n831), .dinb(n828), .dout(n861));
  jnot g00670(.din(n861), .dout(n862));
  jand g00671(.dina(n862), .dinb(n834), .dout(n863));
  jxor g00672(.dina(n863), .dinb(n860), .dout(n864));
  jxor g00673(.dina(n864), .dinb(n852), .dout(n865));
  jnot g00674(.din(n820), .dout(n866));
  jand g00675(.dina(n804), .dinb(n802), .dout(n867));
  jxor g00676(.dina(n867), .dinb(n866), .dout(n868));
  jand g00677(.dina(\a[16] ), .dinb(\a[3] ), .dout(n869));
  jand g00678(.dina(\a[11] ), .dinb(\a[8] ), .dout(n870));
  jxor g00679(.dina(n870), .dinb(n453), .dout(n871));
  jxor g00680(.dina(n871), .dinb(n869), .dout(n872));
  jxor g00681(.dina(n872), .dinb(n868), .dout(n873));
  jxor g00682(.dina(n873), .dinb(n865), .dout(n874));
  jand g00683(.dina(n773), .dinb(n770), .dout(n875));
  jand g00684(.dina(n780), .dinb(n774), .dout(n876));
  jor  g00685(.dina(n876), .dinb(n875), .dout(n877));
  jand g00686(.dina(\a[17] ), .dinb(\a[15] ), .dout(n878));
  jand g00687(.dina(n878), .dinb(n245), .dout(n879));
  jand g00688(.dina(n212), .dinb(\a[15] ), .dout(n880));
  jand g00689(.dina(\a[17] ), .dinb(\a[2] ), .dout(n881));
  jand g00690(.dina(n881), .dinb(\a[0] ), .dout(n882));
  jor  g00691(.dina(n882), .dinb(n880), .dout(n883));
  jand g00692(.dina(n883), .dinb(\a[19] ), .dout(n884));
  jor  g00693(.dina(n884), .dinb(n879), .dout(n885));
  jnot g00694(.din(n885), .dout(n886));
  jand g00695(.dina(\a[15] ), .dinb(\a[4] ), .dout(n887));
  jor  g00696(.dina(n887), .dinb(n881), .dout(n888));
  jand g00697(.dina(n888), .dinb(n886), .dout(n889));
  jnot g00698(.din(n889), .dout(n890));
  jnot g00699(.din(\a[19] ), .dout(n891));
  jnot g00700(.din(n879), .dout(n892));
  jand g00701(.dina(n883), .dinb(n892), .dout(n893));
  jor  g00702(.dina(n893), .dinb(n891), .dout(n894));
  jor  g00703(.dina(n894), .dinb(n193), .dout(n895));
  jand g00704(.dina(n895), .dinb(n890), .dout(n896));
  jand g00705(.dina(\a[14] ), .dinb(\a[5] ), .dout(n897));
  jnot g00706(.din(n897), .dout(n898));
  jand g00707(.dina(\a[13] ), .dinb(\a[12] ), .dout(n899));
  jand g00708(.dina(n899), .dinb(n410), .dout(n900));
  jnot g00709(.din(n900), .dout(n901));
  jand g00710(.dina(\a[13] ), .dinb(\a[6] ), .dout(n902));
  jand g00711(.dina(\a[12] ), .dinb(\a[7] ), .dout(n903));
  jor  g00712(.dina(n903), .dinb(n902), .dout(n904));
  jand g00713(.dina(n904), .dinb(n901), .dout(n905));
  jxor g00714(.dina(n905), .dinb(n898), .dout(n906));
  jxor g00715(.dina(n906), .dinb(n896), .dout(n907));
  jxor g00716(.dina(n907), .dinb(n877), .dout(n908));
  jnot g00717(.din(n908), .dout(n909));
  jor  g00718(.dina(n788), .dinb(n785), .dout(n910));
  jand g00719(.dina(n789), .dinb(n781), .dout(n911));
  jnot g00720(.din(n911), .dout(n912));
  jand g00721(.dina(n912), .dinb(n910), .dout(n913));
  jxor g00722(.dina(n913), .dinb(n909), .dout(n914));
  jxor g00723(.dina(n914), .dinb(n874), .dout(n915));
  jand g00724(.dina(n839), .dinb(n793), .dout(n916));
  jand g00725(.dina(n840), .dinb(n790), .dout(n917));
  jor  g00726(.dina(n917), .dinb(n916), .dout(n918));
  jnot g00727(.din(n918), .dout(n919));
  jxor g00728(.dina(n919), .dinb(n915), .dout(n920));
  jnot g00729(.din(n842), .dout(n921));
  jor  g00730(.dina(n848), .dinb(n844), .dout(n922));
  jand g00731(.dina(n922), .dinb(n921), .dout(n923));
  jxor g00732(.dina(n923), .dinb(n920), .dout(\asquared[20] ));
  jor  g00733(.dina(n913), .dinb(n909), .dout(n925));
  jand g00734(.dina(n914), .dinb(n874), .dout(n926));
  jnot g00735(.din(n926), .dout(n927));
  jand g00736(.dina(n927), .dinb(n925), .dout(n928));
  jand g00737(.dina(n867), .dinb(n866), .dout(n929));
  jand g00738(.dina(n872), .dinb(n868), .dout(n930));
  jor  g00739(.dina(n930), .dinb(n929), .dout(n931));
  jand g00740(.dina(n863), .dinb(n860), .dout(n932));
  jor  g00741(.dina(n932), .dinb(n855), .dout(n933));
  jnot g00742(.din(n933), .dout(n934));
  jand g00743(.dina(\a[18] ), .dinb(\a[2] ), .dout(n935));
  jnot g00744(.din(n935), .dout(n936));
  jand g00745(.dina(\a[17] ), .dinb(\a[16] ), .dout(n937));
  jand g00746(.dina(n937), .dinb(n265), .dout(n938));
  jnot g00747(.din(n938), .dout(n939));
  jand g00748(.dina(\a[17] ), .dinb(\a[3] ), .dout(n940));
  jand g00749(.dina(\a[16] ), .dinb(\a[4] ), .dout(n941));
  jor  g00750(.dina(n941), .dinb(n940), .dout(n942));
  jand g00751(.dina(n942), .dinb(n939), .dout(n943));
  jxor g00752(.dina(n943), .dinb(n936), .dout(n944));
  jxor g00753(.dina(n944), .dinb(n934), .dout(n945));
  jxor g00754(.dina(n945), .dinb(n931), .dout(n946));
  jand g00755(.dina(n864), .dinb(n852), .dout(n947));
  jand g00756(.dina(n873), .dinb(n865), .dout(n948));
  jor  g00757(.dina(n948), .dinb(n947), .dout(n949));
  jxor g00758(.dina(n949), .dinb(n946), .dout(n950));
  jor  g00759(.dina(n906), .dinb(n896), .dout(n951));
  jand g00760(.dina(n907), .dinb(n877), .dout(n952));
  jnot g00761(.din(n952), .dout(n953));
  jand g00762(.dina(n953), .dinb(n951), .dout(n954));
  jnot g00763(.din(n954), .dout(n955));
  jand g00764(.dina(n870), .dinb(n453), .dout(n956));
  jand g00765(.dina(n871), .dinb(n869), .dout(n957));
  jor  g00766(.dina(n957), .dinb(n956), .dout(n958));
  jand g00767(.dina(\a[11] ), .dinb(\a[9] ), .dout(n959));
  jand g00768(.dina(\a[19] ), .dinb(\a[1] ), .dout(n960));
  jxor g00769(.dina(n960), .dinb(n959), .dout(n961));
  jxor g00770(.dina(n961), .dinb(n958), .dout(n962));
  jxor g00771(.dina(n962), .dinb(n885), .dout(n963));
  jxor g00772(.dina(n963), .dinb(n955), .dout(n964));
  jand g00773(.dina(n857), .dinb(\a[10] ), .dout(n965));
  jand g00774(.dina(\a[20] ), .dinb(\a[0] ), .dout(n966));
  jand g00775(.dina(\a[13] ), .dinb(\a[7] ), .dout(n967));
  jxor g00776(.dina(n967), .dinb(n966), .dout(n968));
  jxor g00777(.dina(n968), .dinb(n965), .dout(n969));
  jand g00778(.dina(n901), .dinb(n898), .dout(n970));
  jnot g00779(.din(n970), .dout(n971));
  jand g00780(.dina(n971), .dinb(n904), .dout(n972));
  jxor g00781(.dina(n972), .dinb(n969), .dout(n973));
  jnot g00782(.din(n973), .dout(n974));
  jand g00783(.dina(\a[12] ), .dinb(\a[8] ), .dout(n975));
  jand g00784(.dina(\a[15] ), .dinb(\a[14] ), .dout(n976));
  jand g00785(.dina(n976), .dinb(n339), .dout(n977));
  jnot g00786(.din(n977), .dout(n978));
  jand g00787(.dina(\a[14] ), .dinb(\a[12] ), .dout(n979));
  jand g00788(.dina(n979), .dinb(n544), .dout(n980));
  jand g00789(.dina(\a[15] ), .dinb(\a[5] ), .dout(n981));
  jand g00790(.dina(n981), .dinb(n975), .dout(n982));
  jor  g00791(.dina(n982), .dinb(n980), .dout(n983));
  jand g00792(.dina(n983), .dinb(n978), .dout(n984));
  jnot g00793(.din(n984), .dout(n985));
  jand g00794(.dina(n985), .dinb(n975), .dout(n986));
  jnot g00795(.din(n986), .dout(n987));
  jor  g00796(.dina(n983), .dinb(n977), .dout(n988));
  jnot g00797(.din(n981), .dout(n989));
  jand g00798(.dina(\a[14] ), .dinb(\a[6] ), .dout(n990));
  jnot g00799(.din(n990), .dout(n991));
  jand g00800(.dina(n991), .dinb(n989), .dout(n992));
  jor  g00801(.dina(n992), .dinb(n988), .dout(n993));
  jand g00802(.dina(n993), .dinb(n987), .dout(n994));
  jxor g00803(.dina(n994), .dinb(n974), .dout(n995));
  jxor g00804(.dina(n995), .dinb(n964), .dout(n996));
  jxor g00805(.dina(n996), .dinb(n950), .dout(n997));
  jxor g00806(.dina(n997), .dinb(n928), .dout(n998));
  jand g00807(.dina(n918), .dinb(n915), .dout(n999));
  jnot g00808(.din(n999), .dout(n1000));
  jnot g00809(.din(n915), .dout(n1001));
  jand g00810(.dina(n919), .dinb(n1001), .dout(n1002));
  jor  g00811(.dina(n923), .dinb(n1002), .dout(n1003));
  jand g00812(.dina(n1003), .dinb(n1000), .dout(n1004));
  jxor g00813(.dina(n1004), .dinb(n998), .dout(\asquared[21] ));
  jand g00814(.dina(n949), .dinb(n946), .dout(n1006));
  jand g00815(.dina(n996), .dinb(n950), .dout(n1007));
  jor  g00816(.dina(n1007), .dinb(n1006), .dout(n1008));
  jand g00817(.dina(n939), .dinb(n936), .dout(n1009));
  jnot g00818(.din(n1009), .dout(n1010));
  jand g00819(.dina(n1010), .dinb(n942), .dout(n1011));
  jxor g00820(.dina(n1011), .dinb(n988), .dout(n1012));
  jand g00821(.dina(n967), .dinb(n966), .dout(n1013));
  jand g00822(.dina(n968), .dinb(n965), .dout(n1014));
  jor  g00823(.dina(n1014), .dinb(n1013), .dout(n1015));
  jxor g00824(.dina(n1015), .dinb(n1012), .dout(n1016));
  jnot g00825(.din(n1016), .dout(n1017));
  jor  g00826(.dina(n944), .dinb(n934), .dout(n1018));
  jand g00827(.dina(n945), .dinb(n931), .dout(n1019));
  jnot g00828(.din(n1019), .dout(n1020));
  jand g00829(.dina(n1020), .dinb(n1018), .dout(n1021));
  jxor g00830(.dina(n1021), .dinb(n1017), .dout(n1022));
  jand g00831(.dina(\a[16] ), .dinb(\a[5] ), .dout(n1023));
  jand g00832(.dina(\a[19] ), .dinb(\a[18] ), .dout(n1024));
  jand g00833(.dina(n1024), .dinb(n248), .dout(n1025));
  jnot g00834(.din(n1025), .dout(n1026));
  jand g00835(.dina(\a[19] ), .dinb(\a[2] ), .dout(n1027));
  jand g00836(.dina(\a[18] ), .dinb(\a[3] ), .dout(n1028));
  jor  g00837(.dina(n1028), .dinb(n1027), .dout(n1029));
  jand g00838(.dina(n1029), .dinb(n1026), .dout(n1030));
  jxor g00839(.dina(n1030), .dinb(n1023), .dout(n1031));
  jnot g00840(.din(n1031), .dout(n1032));
  jand g00841(.dina(\a[15] ), .dinb(\a[6] ), .dout(n1033));
  jnot g00842(.din(n1033), .dout(n1034));
  jand g00843(.dina(n675), .dinb(n499), .dout(n1035));
  jnot g00844(.din(n1035), .dout(n1036));
  jand g00845(.dina(\a[13] ), .dinb(\a[8] ), .dout(n1037));
  jand g00846(.dina(\a[14] ), .dinb(\a[7] ), .dout(n1038));
  jor  g00847(.dina(n1038), .dinb(n1037), .dout(n1039));
  jand g00848(.dina(n1039), .dinb(n1036), .dout(n1040));
  jxor g00849(.dina(n1040), .dinb(n1034), .dout(n1041));
  jxor g00850(.dina(n1041), .dinb(n1032), .dout(n1042));
  jnot g00851(.din(n1042), .dout(n1043));
  jand g00852(.dina(\a[17] ), .dinb(\a[4] ), .dout(n1044));
  jnot g00853(.din(n1044), .dout(n1045));
  jand g00854(.dina(n555), .dinb(n453), .dout(n1046));
  jnot g00855(.din(n1046), .dout(n1047));
  jand g00856(.dina(\a[12] ), .dinb(\a[9] ), .dout(n1048));
  jor  g00857(.dina(n1048), .dinb(n655), .dout(n1049));
  jand g00858(.dina(n1049), .dinb(n1047), .dout(n1050));
  jxor g00859(.dina(n1050), .dinb(n1045), .dout(n1051));
  jxor g00860(.dina(n1051), .dinb(n1043), .dout(n1052));
  jxor g00861(.dina(n1052), .dinb(n1022), .dout(n1053));
  jand g00862(.dina(n961), .dinb(n958), .dout(n1054));
  jand g00863(.dina(n962), .dinb(n885), .dout(n1055));
  jor  g00864(.dina(n1055), .dinb(n1054), .dout(n1056));
  jand g00865(.dina(n960), .dinb(n959), .dout(n1057));
  jand g00866(.dina(\a[21] ), .dinb(\a[0] ), .dout(n1058));
  jxor g00867(.dina(n1058), .dinb(n1057), .dout(n1059));
  jand g00868(.dina(\a[20] ), .dinb(\a[1] ), .dout(n1060));
  jxor g00869(.dina(n1060), .dinb(\a[11] ), .dout(n1061));
  jxor g00870(.dina(n1061), .dinb(n1059), .dout(n1062));
  jxor g00871(.dina(n1062), .dinb(n1056), .dout(n1063));
  jnot g00872(.din(n1063), .dout(n1064));
  jand g00873(.dina(n972), .dinb(n969), .dout(n1065));
  jnot g00874(.din(n1065), .dout(n1066));
  jor  g00875(.dina(n994), .dinb(n974), .dout(n1067));
  jand g00876(.dina(n1067), .dinb(n1066), .dout(n1068));
  jxor g00877(.dina(n1068), .dinb(n1064), .dout(n1069));
  jand g00878(.dina(n963), .dinb(n955), .dout(n1070));
  jand g00879(.dina(n995), .dinb(n964), .dout(n1071));
  jor  g00880(.dina(n1071), .dinb(n1070), .dout(n1072));
  jxor g00881(.dina(n1072), .dinb(n1069), .dout(n1073));
  jxor g00882(.dina(n1073), .dinb(n1053), .dout(n1074));
  jand g00883(.dina(n1074), .dinb(n1008), .dout(n1075));
  jor  g00884(.dina(n1074), .dinb(n1008), .dout(n1076));
  jnot g00885(.din(n1076), .dout(n1077));
  jor  g00886(.dina(n1077), .dinb(n1075), .dout(n1078));
  jnot g00887(.din(n928), .dout(n1079));
  jand g00888(.dina(n997), .dinb(n1079), .dout(n1080));
  jnot g00889(.din(n1080), .dout(n1081));
  jor  g00890(.dina(n997), .dinb(n1079), .dout(n1082));
  jnot g00891(.din(n1082), .dout(n1083));
  jor  g00892(.dina(n1004), .dinb(n1083), .dout(n1084));
  jand g00893(.dina(n1084), .dinb(n1081), .dout(n1085));
  jxor g00894(.dina(n1085), .dinb(n1078), .dout(\asquared[22] ));
  jand g00895(.dina(n1072), .dinb(n1069), .dout(n1087));
  jand g00896(.dina(n1073), .dinb(n1053), .dout(n1088));
  jor  g00897(.dina(n1088), .dinb(n1087), .dout(n1089));
  jand g00898(.dina(n1030), .dinb(n1023), .dout(n1090));
  jor  g00899(.dina(n1090), .dinb(n1025), .dout(n1091));
  jand g00900(.dina(n1036), .dinb(n1034), .dout(n1092));
  jnot g00901(.din(n1092), .dout(n1093));
  jand g00902(.dina(n1093), .dinb(n1039), .dout(n1094));
  jxor g00903(.dina(n1094), .dinb(n1091), .dout(n1095));
  jand g00904(.dina(n1058), .dinb(n1057), .dout(n1096));
  jand g00905(.dina(n1061), .dinb(n1059), .dout(n1097));
  jor  g00906(.dina(n1097), .dinb(n1096), .dout(n1098));
  jxor g00907(.dina(n1098), .dinb(n1095), .dout(n1099));
  jnot g00908(.din(n1099), .dout(n1100));
  jand g00909(.dina(n1062), .dinb(n1056), .dout(n1101));
  jnot g00910(.din(n1101), .dout(n1102));
  jor  g00911(.dina(n1068), .dinb(n1064), .dout(n1103));
  jand g00912(.dina(n1103), .dinb(n1102), .dout(n1104));
  jxor g00913(.dina(n1104), .dinb(n1100), .dout(n1105));
  jand g00914(.dina(\a[19] ), .dinb(\a[3] ), .dout(n1106));
  jand g00915(.dina(\a[18] ), .dinb(\a[17] ), .dout(n1107));
  jand g00916(.dina(n1107), .dinb(n242), .dout(n1108));
  jnot g00917(.din(n1108), .dout(n1109));
  jand g00918(.dina(n1024), .dinb(n265), .dout(n1110));
  jand g00919(.dina(\a[17] ), .dinb(\a[5] ), .dout(n1111));
  jand g00920(.dina(n1111), .dinb(n1106), .dout(n1112));
  jor  g00921(.dina(n1112), .dinb(n1110), .dout(n1113));
  jand g00922(.dina(n1113), .dinb(n1109), .dout(n1114));
  jnot g00923(.din(n1114), .dout(n1115));
  jand g00924(.dina(n1115), .dinb(n1106), .dout(n1116));
  jor  g00925(.dina(n1113), .dinb(n1108), .dout(n1117));
  jnot g00926(.din(n1117), .dout(n1118));
  jand g00927(.dina(\a[18] ), .dinb(\a[4] ), .dout(n1119));
  jor  g00928(.dina(n1119), .dinb(n1111), .dout(n1120));
  jand g00929(.dina(n1120), .dinb(n1118), .dout(n1121));
  jor  g00930(.dina(n1121), .dinb(n1116), .dout(n1122));
  jand g00931(.dina(\a[22] ), .dinb(\a[0] ), .dout(n1123));
  jand g00932(.dina(\a[15] ), .dinb(\a[7] ), .dout(n1124));
  jand g00933(.dina(\a[14] ), .dinb(\a[8] ), .dout(n1125));
  jor  g00934(.dina(n1125), .dinb(n1124), .dout(n1126));
  jand g00935(.dina(n976), .dinb(n499), .dout(n1127));
  jnot g00936(.din(n1127), .dout(n1128));
  jand g00937(.dina(n1128), .dinb(n1126), .dout(n1129));
  jxor g00938(.dina(n1129), .dinb(n1123), .dout(n1130));
  jand g00939(.dina(\a[16] ), .dinb(\a[6] ), .dout(n1131));
  jand g00940(.dina(\a[20] ), .dinb(\a[2] ), .dout(n1132));
  jxor g00941(.dina(n1132), .dinb(n1131), .dout(n1133));
  jxor g00942(.dina(n1133), .dinb(n479), .dout(n1134));
  jxor g00943(.dina(n1134), .dinb(n1130), .dout(n1135));
  jxor g00944(.dina(n1135), .dinb(n1122), .dout(n1136));
  jxor g00945(.dina(n1136), .dinb(n1105), .dout(n1137));
  jor  g00946(.dina(n1021), .dinb(n1017), .dout(n1138));
  jand g00947(.dina(n1052), .dinb(n1022), .dout(n1139));
  jnot g00948(.din(n1139), .dout(n1140));
  jand g00949(.dina(n1140), .dinb(n1138), .dout(n1141));
  jnot g00950(.din(n1141), .dout(n1142));
  jor  g00951(.dina(n1041), .dinb(n1032), .dout(n1143));
  jor  g00952(.dina(n1051), .dinb(n1043), .dout(n1144));
  jand g00953(.dina(n1144), .dinb(n1143), .dout(n1145));
  jnot g00954(.din(n1145), .dout(n1146));
  jand g00955(.dina(n1011), .dinb(n988), .dout(n1147));
  jand g00956(.dina(n1015), .dinb(n1012), .dout(n1148));
  jor  g00957(.dina(n1148), .dinb(n1147), .dout(n1149));
  jand g00958(.dina(n1060), .dinb(\a[11] ), .dout(n1150));
  jand g00959(.dina(\a[12] ), .dinb(\a[10] ), .dout(n1151));
  jand g00960(.dina(\a[21] ), .dinb(\a[1] ), .dout(n1152));
  jxor g00961(.dina(n1152), .dinb(n1151), .dout(n1153));
  jxor g00962(.dina(n1153), .dinb(n1150), .dout(n1154));
  jand g00963(.dina(n1047), .dinb(n1045), .dout(n1155));
  jnot g00964(.din(n1155), .dout(n1156));
  jand g00965(.dina(n1156), .dinb(n1049), .dout(n1157));
  jxor g00966(.dina(n1157), .dinb(n1154), .dout(n1158));
  jxor g00967(.dina(n1158), .dinb(n1149), .dout(n1159));
  jxor g00968(.dina(n1159), .dinb(n1146), .dout(n1160));
  jxor g00969(.dina(n1160), .dinb(n1142), .dout(n1161));
  jxor g00970(.dina(n1161), .dinb(n1137), .dout(n1162));
  jand g00971(.dina(n1162), .dinb(n1089), .dout(n1163));
  jor  g00972(.dina(n1162), .dinb(n1089), .dout(n1164));
  jnot g00973(.din(n1164), .dout(n1165));
  jor  g00974(.dina(n1165), .dinb(n1163), .dout(n1166));
  jnot g00975(.din(n1075), .dout(n1167));
  jor  g00976(.dina(n1085), .dinb(n1077), .dout(n1168));
  jand g00977(.dina(n1168), .dinb(n1167), .dout(n1169));
  jxor g00978(.dina(n1169), .dinb(n1166), .dout(\asquared[23] ));
  jand g00979(.dina(n1160), .dinb(n1142), .dout(n1171));
  jand g00980(.dina(n1161), .dinb(n1137), .dout(n1172));
  jor  g00981(.dina(n1172), .dinb(n1171), .dout(n1173));
  jand g00982(.dina(n1158), .dinb(n1149), .dout(n1174));
  jand g00983(.dina(n1159), .dinb(n1146), .dout(n1175));
  jor  g00984(.dina(n1175), .dinb(n1174), .dout(n1176));
  jand g00985(.dina(n1153), .dinb(n1150), .dout(n1177));
  jand g00986(.dina(n1157), .dinb(n1154), .dout(n1178));
  jor  g00987(.dina(n1178), .dinb(n1177), .dout(n1179));
  jand g00988(.dina(\a[17] ), .dinb(\a[6] ), .dout(n1180));
  jand g00989(.dina(\a[20] ), .dinb(\a[18] ), .dout(n1181));
  jand g00990(.dina(n1181), .dinb(n310), .dout(n1182));
  jnot g00991(.din(n1182), .dout(n1183));
  jand g00992(.dina(\a[20] ), .dinb(\a[3] ), .dout(n1184));
  jand g00993(.dina(\a[18] ), .dinb(\a[5] ), .dout(n1185));
  jor  g00994(.dina(n1185), .dinb(n1184), .dout(n1186));
  jand g00995(.dina(n1186), .dinb(n1183), .dout(n1187));
  jxor g00996(.dina(n1187), .dinb(n1180), .dout(n1188));
  jnot g00997(.din(n1188), .dout(n1189));
  jand g00998(.dina(\a[19] ), .dinb(\a[4] ), .dout(n1190));
  jnot g00999(.din(n1190), .dout(n1191));
  jand g01000(.dina(n899), .dinb(n655), .dout(n1192));
  jnot g01001(.din(n1192), .dout(n1193));
  jand g01002(.dina(\a[13] ), .dinb(\a[10] ), .dout(n1194));
  jor  g01003(.dina(n1194), .dinb(n555), .dout(n1195));
  jand g01004(.dina(n1195), .dinb(n1193), .dout(n1196));
  jxor g01005(.dina(n1196), .dinb(n1191), .dout(n1197));
  jxor g01006(.dina(n1197), .dinb(n1189), .dout(n1198));
  jxor g01007(.dina(n1198), .dinb(n1179), .dout(n1199));
  jand g01008(.dina(n1129), .dinb(n1123), .dout(n1200));
  jor  g01009(.dina(n1200), .dinb(n1127), .dout(n1201));
  jand g01010(.dina(n1152), .dinb(n1151), .dout(n1202));
  jand g01011(.dina(\a[23] ), .dinb(\a[0] ), .dout(n1203));
  jand g01012(.dina(\a[21] ), .dinb(\a[2] ), .dout(n1204));
  jor  g01013(.dina(n1204), .dinb(n1203), .dout(n1205));
  jand g01014(.dina(\a[23] ), .dinb(\a[2] ), .dout(n1206));
  jand g01015(.dina(n1206), .dinb(n1058), .dout(n1207));
  jnot g01016(.din(n1207), .dout(n1208));
  jand g01017(.dina(n1208), .dinb(n1205), .dout(n1209));
  jxor g01018(.dina(n1209), .dinb(n1202), .dout(n1210));
  jxor g01019(.dina(n1210), .dinb(n1201), .dout(n1211));
  jand g01020(.dina(\a[16] ), .dinb(\a[7] ), .dout(n1212));
  jand g01021(.dina(n976), .dinb(n395), .dout(n1213));
  jnot g01022(.din(n1213), .dout(n1214));
  jand g01023(.dina(\a[15] ), .dinb(\a[8] ), .dout(n1215));
  jand g01024(.dina(\a[14] ), .dinb(\a[9] ), .dout(n1216));
  jor  g01025(.dina(n1216), .dinb(n1215), .dout(n1217));
  jand g01026(.dina(n1217), .dinb(n1214), .dout(n1218));
  jxor g01027(.dina(n1218), .dinb(n1212), .dout(n1219));
  jxor g01028(.dina(n1219), .dinb(n1211), .dout(n1220));
  jxor g01029(.dina(n1220), .dinb(n1199), .dout(n1221));
  jxor g01030(.dina(n1221), .dinb(n1176), .dout(n1222));
  jor  g01031(.dina(n1104), .dinb(n1100), .dout(n1223));
  jand g01032(.dina(n1136), .dinb(n1105), .dout(n1224));
  jnot g01033(.din(n1224), .dout(n1225));
  jand g01034(.dina(n1225), .dinb(n1223), .dout(n1226));
  jnot g01035(.din(n1226), .dout(n1227));
  jand g01036(.dina(n1094), .dinb(n1091), .dout(n1228));
  jand g01037(.dina(n1098), .dinb(n1095), .dout(n1229));
  jor  g01038(.dina(n1229), .dinb(n1228), .dout(n1230));
  jand g01039(.dina(n1134), .dinb(n1130), .dout(n1231));
  jand g01040(.dina(n1135), .dinb(n1122), .dout(n1232));
  jor  g01041(.dina(n1232), .dinb(n1231), .dout(n1233));
  jxor g01042(.dina(n1233), .dinb(n1230), .dout(n1234));
  jand g01043(.dina(n1132), .dinb(n1131), .dout(n1235));
  jand g01044(.dina(n1133), .dinb(n479), .dout(n1236));
  jor  g01045(.dina(n1236), .dinb(n1235), .dout(n1237));
  jand g01046(.dina(\a[22] ), .dinb(\a[1] ), .dout(n1238));
  jxor g01047(.dina(n1238), .dinb(\a[12] ), .dout(n1239));
  jxor g01048(.dina(n1239), .dinb(n1117), .dout(n1240));
  jxor g01049(.dina(n1240), .dinb(n1237), .dout(n1241));
  jxor g01050(.dina(n1241), .dinb(n1234), .dout(n1242));
  jxor g01051(.dina(n1242), .dinb(n1227), .dout(n1243));
  jxor g01052(.dina(n1243), .dinb(n1222), .dout(n1244));
  jnot g01053(.din(n1244), .dout(n1245));
  jxor g01054(.dina(n1245), .dinb(n1173), .dout(n1246));
  jnot g01055(.din(n1163), .dout(n1247));
  jor  g01056(.dina(n1169), .dinb(n1165), .dout(n1248));
  jand g01057(.dina(n1248), .dinb(n1247), .dout(n1249));
  jxor g01058(.dina(n1249), .dinb(n1246), .dout(\asquared[24] ));
  jand g01059(.dina(n1242), .dinb(n1227), .dout(n1251));
  jand g01060(.dina(n1243), .dinb(n1222), .dout(n1252));
  jor  g01061(.dina(n1252), .dinb(n1251), .dout(n1253));
  jand g01062(.dina(n1239), .dinb(n1117), .dout(n1254));
  jand g01063(.dina(n1240), .dinb(n1237), .dout(n1255));
  jor  g01064(.dina(n1255), .dinb(n1254), .dout(n1256));
  jand g01065(.dina(\a[17] ), .dinb(\a[7] ), .dout(n1257));
  jand g01066(.dina(\a[22] ), .dinb(\a[18] ), .dout(n1258));
  jand g01067(.dina(n1258), .dinb(n301), .dout(n1259));
  jnot g01068(.din(n1259), .dout(n1260));
  jand g01069(.dina(n1107), .dinb(n410), .dout(n1261));
  jand g01070(.dina(\a[22] ), .dinb(\a[2] ), .dout(n1262));
  jand g01071(.dina(n1262), .dinb(n1257), .dout(n1263));
  jor  g01072(.dina(n1263), .dinb(n1261), .dout(n1264));
  jand g01073(.dina(n1264), .dinb(n1260), .dout(n1265));
  jnot g01074(.din(n1265), .dout(n1266));
  jand g01075(.dina(n1266), .dinb(n1257), .dout(n1267));
  jor  g01076(.dina(n1264), .dinb(n1259), .dout(n1268));
  jnot g01077(.din(n1268), .dout(n1269));
  jand g01078(.dina(\a[18] ), .dinb(\a[6] ), .dout(n1270));
  jor  g01079(.dina(n1270), .dinb(n1262), .dout(n1271));
  jand g01080(.dina(n1271), .dinb(n1269), .dout(n1272));
  jor  g01081(.dina(n1272), .dinb(n1267), .dout(n1273));
  jand g01082(.dina(n1238), .dinb(\a[12] ), .dout(n1274));
  jand g01083(.dina(\a[24] ), .dinb(\a[0] ), .dout(n1275));
  jxor g01084(.dina(n1275), .dinb(n1274), .dout(n1276));
  jand g01085(.dina(\a[23] ), .dinb(\a[1] ), .dout(n1277));
  jxor g01086(.dina(n1277), .dinb(n816), .dout(n1278));
  jxor g01087(.dina(n1278), .dinb(n1276), .dout(n1279));
  jxor g01088(.dina(n1279), .dinb(n1273), .dout(n1280));
  jxor g01089(.dina(n1280), .dinb(n1256), .dout(n1281));
  jand g01090(.dina(n1209), .dinb(n1202), .dout(n1282));
  jor  g01091(.dina(n1282), .dinb(n1207), .dout(n1283));
  jnot g01092(.din(n1283), .dout(n1284));
  jand g01093(.dina(\a[21] ), .dinb(\a[3] ), .dout(n1285));
  jnot g01094(.din(n1285), .dout(n1286));
  jand g01095(.dina(\a[20] ), .dinb(\a[19] ), .dout(n1287));
  jand g01096(.dina(n1287), .dinb(n242), .dout(n1288));
  jnot g01097(.din(n1288), .dout(n1289));
  jand g01098(.dina(\a[20] ), .dinb(\a[4] ), .dout(n1290));
  jand g01099(.dina(\a[19] ), .dinb(\a[5] ), .dout(n1291));
  jor  g01100(.dina(n1291), .dinb(n1290), .dout(n1292));
  jand g01101(.dina(n1292), .dinb(n1289), .dout(n1293));
  jxor g01102(.dina(n1293), .dinb(n1286), .dout(n1294));
  jxor g01103(.dina(n1294), .dinb(n1284), .dout(n1295));
  jnot g01104(.din(n1295), .dout(n1296));
  jand g01105(.dina(\a[16] ), .dinb(\a[8] ), .dout(n1297));
  jnot g01106(.din(n1297), .dout(n1298));
  jand g01107(.dina(n976), .dinb(n453), .dout(n1299));
  jnot g01108(.din(n1299), .dout(n1300));
  jand g01109(.dina(\a[15] ), .dinb(\a[9] ), .dout(n1301));
  jand g01110(.dina(\a[14] ), .dinb(\a[10] ), .dout(n1302));
  jor  g01111(.dina(n1302), .dinb(n1301), .dout(n1303));
  jand g01112(.dina(n1303), .dinb(n1300), .dout(n1304));
  jxor g01113(.dina(n1304), .dinb(n1298), .dout(n1305));
  jxor g01114(.dina(n1305), .dinb(n1296), .dout(n1306));
  jxor g01115(.dina(n1306), .dinb(n1281), .dout(n1307));
  jand g01116(.dina(n1233), .dinb(n1230), .dout(n1308));
  jand g01117(.dina(n1241), .dinb(n1234), .dout(n1309));
  jor  g01118(.dina(n1309), .dinb(n1308), .dout(n1310));
  jxor g01119(.dina(n1310), .dinb(n1307), .dout(n1311));
  jand g01120(.dina(n1220), .dinb(n1199), .dout(n1312));
  jand g01121(.dina(n1221), .dinb(n1176), .dout(n1313));
  jor  g01122(.dina(n1313), .dinb(n1312), .dout(n1314));
  jand g01123(.dina(n1217), .dinb(n1212), .dout(n1315));
  jor  g01124(.dina(n1315), .dinb(n1213), .dout(n1316));
  jand g01125(.dina(n1187), .dinb(n1180), .dout(n1317));
  jor  g01126(.dina(n1317), .dinb(n1182), .dout(n1318));
  jand g01127(.dina(n1193), .dinb(n1191), .dout(n1319));
  jnot g01128(.din(n1319), .dout(n1320));
  jand g01129(.dina(n1320), .dinb(n1195), .dout(n1321));
  jxor g01130(.dina(n1321), .dinb(n1318), .dout(n1322));
  jxor g01131(.dina(n1322), .dinb(n1316), .dout(n1323));
  jor  g01132(.dina(n1197), .dinb(n1189), .dout(n1324));
  jand g01133(.dina(n1198), .dinb(n1179), .dout(n1325));
  jnot g01134(.din(n1325), .dout(n1326));
  jand g01135(.dina(n1326), .dinb(n1324), .dout(n1327));
  jnot g01136(.din(n1327), .dout(n1328));
  jand g01137(.dina(n1210), .dinb(n1201), .dout(n1329));
  jand g01138(.dina(n1219), .dinb(n1211), .dout(n1330));
  jor  g01139(.dina(n1330), .dinb(n1329), .dout(n1331));
  jxor g01140(.dina(n1331), .dinb(n1328), .dout(n1332));
  jxor g01141(.dina(n1332), .dinb(n1323), .dout(n1333));
  jxor g01142(.dina(n1333), .dinb(n1314), .dout(n1334));
  jxor g01143(.dina(n1334), .dinb(n1311), .dout(n1335));
  jand g01144(.dina(n1335), .dinb(n1253), .dout(n1336));
  jor  g01145(.dina(n1335), .dinb(n1253), .dout(n1337));
  jnot g01146(.din(n1337), .dout(n1338));
  jor  g01147(.dina(n1338), .dinb(n1336), .dout(n1339));
  jand g01148(.dina(n1244), .dinb(n1173), .dout(n1340));
  jnot g01149(.din(n1340), .dout(n1341));
  jnot g01150(.din(n1173), .dout(n1342));
  jand g01151(.dina(n1245), .dinb(n1342), .dout(n1343));
  jor  g01152(.dina(n1249), .dinb(n1343), .dout(n1344));
  jand g01153(.dina(n1344), .dinb(n1341), .dout(n1345));
  jxor g01154(.dina(n1345), .dinb(n1339), .dout(\asquared[25] ));
  jand g01155(.dina(n1333), .dinb(n1314), .dout(n1347));
  jand g01156(.dina(n1334), .dinb(n1311), .dout(n1348));
  jor  g01157(.dina(n1348), .dinb(n1347), .dout(n1349));
  jnot g01158(.din(n1349), .dout(n1350));
  jand g01159(.dina(n1331), .dinb(n1328), .dout(n1351));
  jand g01160(.dina(n1332), .dinb(n1323), .dout(n1352));
  jor  g01161(.dina(n1352), .dinb(n1351), .dout(n1353));
  jand g01162(.dina(\a[15] ), .dinb(\a[10] ), .dout(n1354));
  jand g01163(.dina(\a[25] ), .dinb(\a[0] ), .dout(n1355));
  jor  g01164(.dina(n1355), .dinb(n1206), .dout(n1356));
  jand g01165(.dina(\a[25] ), .dinb(\a[2] ), .dout(n1357));
  jand g01166(.dina(n1357), .dinb(n1203), .dout(n1358));
  jnot g01167(.din(n1358), .dout(n1359));
  jand g01168(.dina(n1359), .dinb(n1356), .dout(n1360));
  jxor g01169(.dina(n1360), .dinb(n1354), .dout(n1361));
  jnot g01170(.din(n1361), .dout(n1362));
  jand g01171(.dina(\a[18] ), .dinb(\a[7] ), .dout(n1363));
  jnot g01172(.din(n1363), .dout(n1364));
  jand g01173(.dina(n937), .dinb(n395), .dout(n1365));
  jnot g01174(.din(n1365), .dout(n1366));
  jand g01175(.dina(\a[16] ), .dinb(\a[9] ), .dout(n1367));
  jand g01176(.dina(\a[17] ), .dinb(\a[8] ), .dout(n1368));
  jor  g01177(.dina(n1368), .dinb(n1367), .dout(n1369));
  jand g01178(.dina(n1369), .dinb(n1366), .dout(n1370));
  jxor g01179(.dina(n1370), .dinb(n1364), .dout(n1371));
  jxor g01180(.dina(n1371), .dinb(n1362), .dout(n1372));
  jnot g01181(.din(n1372), .dout(n1373));
  jand g01182(.dina(\a[19] ), .dinb(\a[6] ), .dout(n1374));
  jnot g01183(.din(n1374), .dout(n1375));
  jand g01184(.dina(\a[22] ), .dinb(\a[21] ), .dout(n1376));
  jand g01185(.dina(n1376), .dinb(n265), .dout(n1377));
  jnot g01186(.din(n1377), .dout(n1378));
  jand g01187(.dina(\a[22] ), .dinb(\a[3] ), .dout(n1379));
  jand g01188(.dina(\a[21] ), .dinb(\a[4] ), .dout(n1380));
  jor  g01189(.dina(n1380), .dinb(n1379), .dout(n1381));
  jand g01190(.dina(n1381), .dinb(n1378), .dout(n1382));
  jxor g01191(.dina(n1382), .dinb(n1375), .dout(n1383));
  jxor g01192(.dina(n1383), .dinb(n1373), .dout(n1384));
  jxor g01193(.dina(n1384), .dinb(n1353), .dout(n1385));
  jand g01194(.dina(\a[24] ), .dinb(\a[1] ), .dout(n1386));
  jnot g01195(.din(n1386), .dout(n1387));
  jnot g01196(.din(\a[13] ), .dout(n1388));
  jand g01197(.dina(n1277), .dinb(n816), .dout(n1389));
  jor  g01198(.dina(n1389), .dinb(n1388), .dout(n1390));
  jxor g01199(.dina(n1390), .dinb(n1387), .dout(n1391));
  jand g01200(.dina(n1289), .dinb(n1286), .dout(n1392));
  jnot g01201(.din(n1392), .dout(n1393));
  jand g01202(.dina(n1393), .dinb(n1292), .dout(n1394));
  jxor g01203(.dina(n1394), .dinb(n1391), .dout(n1395));
  jand g01204(.dina(n1321), .dinb(n1318), .dout(n1396));
  jand g01205(.dina(n1322), .dinb(n1316), .dout(n1397));
  jor  g01206(.dina(n1397), .dinb(n1396), .dout(n1398));
  jand g01207(.dina(\a[20] ), .dinb(\a[5] ), .dout(n1399));
  jand g01208(.dina(\a[14] ), .dinb(\a[11] ), .dout(n1400));
  jxor g01209(.dina(n1400), .dinb(n899), .dout(n1401));
  jxor g01210(.dina(n1401), .dinb(n1399), .dout(n1402));
  jxor g01211(.dina(n1402), .dinb(n1398), .dout(n1403));
  jxor g01212(.dina(n1403), .dinb(n1395), .dout(n1404));
  jxor g01213(.dina(n1404), .dinb(n1385), .dout(n1405));
  jand g01214(.dina(n1300), .dinb(n1298), .dout(n1406));
  jnot g01215(.din(n1406), .dout(n1407));
  jand g01216(.dina(n1407), .dinb(n1303), .dout(n1408));
  jxor g01217(.dina(n1408), .dinb(n1268), .dout(n1409));
  jand g01218(.dina(n1275), .dinb(n1274), .dout(n1410));
  jand g01219(.dina(n1278), .dinb(n1276), .dout(n1411));
  jor  g01220(.dina(n1411), .dinb(n1410), .dout(n1412));
  jxor g01221(.dina(n1412), .dinb(n1409), .dout(n1413));
  jnot g01222(.din(n1413), .dout(n1414));
  jor  g01223(.dina(n1294), .dinb(n1284), .dout(n1415));
  jor  g01224(.dina(n1305), .dinb(n1296), .dout(n1416));
  jand g01225(.dina(n1416), .dinb(n1415), .dout(n1417));
  jxor g01226(.dina(n1417), .dinb(n1414), .dout(n1418));
  jand g01227(.dina(n1279), .dinb(n1273), .dout(n1419));
  jand g01228(.dina(n1280), .dinb(n1256), .dout(n1420));
  jor  g01229(.dina(n1420), .dinb(n1419), .dout(n1421));
  jxor g01230(.dina(n1421), .dinb(n1418), .dout(n1422));
  jand g01231(.dina(n1306), .dinb(n1281), .dout(n1423));
  jand g01232(.dina(n1310), .dinb(n1307), .dout(n1424));
  jor  g01233(.dina(n1424), .dinb(n1423), .dout(n1425));
  jxor g01234(.dina(n1425), .dinb(n1422), .dout(n1426));
  jxor g01235(.dina(n1426), .dinb(n1405), .dout(n1427));
  jxor g01236(.dina(n1427), .dinb(n1350), .dout(n1428));
  jnot g01237(.din(n1336), .dout(n1429));
  jor  g01238(.dina(n1345), .dinb(n1338), .dout(n1430));
  jand g01239(.dina(n1430), .dinb(n1429), .dout(n1431));
  jxor g01240(.dina(n1431), .dinb(n1428), .dout(\asquared[26] ));
  jand g01241(.dina(n1425), .dinb(n1422), .dout(n1433));
  jand g01242(.dina(n1426), .dinb(n1405), .dout(n1434));
  jor  g01243(.dina(n1434), .dinb(n1433), .dout(n1435));
  jand g01244(.dina(n1384), .dinb(n1353), .dout(n1436));
  jand g01245(.dina(n1404), .dinb(n1385), .dout(n1437));
  jor  g01246(.dina(n1437), .dinb(n1436), .dout(n1438));
  jand g01247(.dina(n1402), .dinb(n1398), .dout(n1439));
  jand g01248(.dina(n1403), .dinb(n1395), .dout(n1440));
  jor  g01249(.dina(n1440), .dinb(n1439), .dout(n1441));
  jor  g01250(.dina(n1371), .dinb(n1362), .dout(n1442));
  jor  g01251(.dina(n1383), .dinb(n1373), .dout(n1443));
  jand g01252(.dina(n1443), .dinb(n1442), .dout(n1444));
  jnot g01253(.din(n1444), .dout(n1445));
  jand g01254(.dina(\a[25] ), .dinb(\a[1] ), .dout(n1446));
  jxor g01255(.dina(n1446), .dinb(n979), .dout(n1447));
  jor  g01256(.dina(n1400), .dinb(n899), .dout(n1448));
  jand g01257(.dina(n1400), .dinb(n899), .dout(n1449));
  jor  g01258(.dina(n1449), .dinb(n1399), .dout(n1450));
  jand g01259(.dina(n1450), .dinb(n1448), .dout(n1451));
  jxor g01260(.dina(n1451), .dinb(n1447), .dout(n1452));
  jand g01261(.dina(n1378), .dinb(n1375), .dout(n1453));
  jnot g01262(.din(n1453), .dout(n1454));
  jand g01263(.dina(n1454), .dinb(n1381), .dout(n1455));
  jxor g01264(.dina(n1455), .dinb(n1452), .dout(n1456));
  jxor g01265(.dina(n1456), .dinb(n1445), .dout(n1457));
  jxor g01266(.dina(n1457), .dinb(n1441), .dout(n1458));
  jxor g01267(.dina(n1458), .dinb(n1438), .dout(n1459));
  jor  g01268(.dina(n1417), .dinb(n1414), .dout(n1460));
  jand g01269(.dina(n1421), .dinb(n1418), .dout(n1461));
  jnot g01270(.din(n1461), .dout(n1462));
  jand g01271(.dina(n1462), .dinb(n1460), .dout(n1463));
  jnot g01272(.din(n1463), .dout(n1464));
  jand g01273(.dina(\a[17] ), .dinb(\a[9] ), .dout(n1465));
  jnot g01274(.din(n1465), .dout(n1466));
  jand g01275(.dina(n829), .dinb(n655), .dout(n1467));
  jnot g01276(.din(n1467), .dout(n1468));
  jand g01277(.dina(\a[15] ), .dinb(\a[11] ), .dout(n1469));
  jand g01278(.dina(n1469), .dinb(n1465), .dout(n1470));
  jand g01279(.dina(n937), .dinb(n453), .dout(n1471));
  jor  g01280(.dina(n1471), .dinb(n1470), .dout(n1472));
  jand g01281(.dina(n1472), .dinb(n1468), .dout(n1473));
  jor  g01282(.dina(n1473), .dinb(n1466), .dout(n1474));
  jor  g01283(.dina(n1472), .dinb(n1467), .dout(n1475));
  jnot g01284(.din(n1475), .dout(n1476));
  jand g01285(.dina(\a[16] ), .dinb(\a[10] ), .dout(n1477));
  jor  g01286(.dina(n1477), .dinb(n1469), .dout(n1478));
  jand g01287(.dina(n1478), .dinb(n1476), .dout(n1479));
  jnot g01288(.din(n1479), .dout(n1480));
  jand g01289(.dina(n1480), .dinb(n1474), .dout(n1481));
  jand g01290(.dina(\a[24] ), .dinb(\a[2] ), .dout(n1482));
  jand g01291(.dina(\a[23] ), .dinb(\a[3] ), .dout(n1483));
  jand g01292(.dina(\a[19] ), .dinb(\a[7] ), .dout(n1484));
  jxor g01293(.dina(n1484), .dinb(n1483), .dout(n1485));
  jxor g01294(.dina(n1485), .dinb(n1482), .dout(n1486));
  jnot g01295(.din(n1486), .dout(n1487));
  jxor g01296(.dina(n1487), .dinb(n1481), .dout(n1488));
  jand g01297(.dina(\a[22] ), .dinb(\a[4] ), .dout(n1489));
  jand g01298(.dina(\a[21] ), .dinb(\a[20] ), .dout(n1490));
  jand g01299(.dina(n1490), .dinb(n339), .dout(n1491));
  jnot g01300(.din(n1491), .dout(n1492));
  jand g01301(.dina(\a[21] ), .dinb(\a[5] ), .dout(n1493));
  jand g01302(.dina(\a[20] ), .dinb(\a[6] ), .dout(n1494));
  jor  g01303(.dina(n1494), .dinb(n1493), .dout(n1495));
  jand g01304(.dina(n1495), .dinb(n1492), .dout(n1496));
  jxor g01305(.dina(n1496), .dinb(n1489), .dout(n1497));
  jxor g01306(.dina(n1497), .dinb(n1488), .dout(n1498));
  jxor g01307(.dina(n1498), .dinb(n1464), .dout(n1499));
  jand g01308(.dina(n1408), .dinb(n1268), .dout(n1500));
  jand g01309(.dina(n1412), .dinb(n1409), .dout(n1501));
  jor  g01310(.dina(n1501), .dinb(n1500), .dout(n1502));
  jand g01311(.dina(n1394), .dinb(n1391), .dout(n1503));
  jand g01312(.dina(n1387), .dinb(n1389), .dout(n1504));
  jor  g01313(.dina(n1504), .dinb(n1503), .dout(n1505));
  jxor g01314(.dina(n1505), .dinb(n1502), .dout(n1506));
  jand g01315(.dina(n1360), .dinb(n1354), .dout(n1507));
  jor  g01316(.dina(n1507), .dinb(n1358), .dout(n1508));
  jand g01317(.dina(n1366), .dinb(n1364), .dout(n1509));
  jnot g01318(.din(n1509), .dout(n1510));
  jand g01319(.dina(n1510), .dinb(n1369), .dout(n1511));
  jxor g01320(.dina(n1511), .dinb(n1508), .dout(n1512));
  jand g01321(.dina(n1386), .dinb(\a[13] ), .dout(n1513));
  jand g01322(.dina(\a[26] ), .dinb(\a[0] ), .dout(n1514));
  jand g01323(.dina(\a[18] ), .dinb(\a[8] ), .dout(n1515));
  jxor g01324(.dina(n1515), .dinb(n1514), .dout(n1516));
  jxor g01325(.dina(n1516), .dinb(n1513), .dout(n1517));
  jxor g01326(.dina(n1517), .dinb(n1512), .dout(n1518));
  jxor g01327(.dina(n1518), .dinb(n1506), .dout(n1519));
  jxor g01328(.dina(n1519), .dinb(n1499), .dout(n1520));
  jxor g01329(.dina(n1520), .dinb(n1459), .dout(n1521));
  jand g01330(.dina(n1521), .dinb(n1435), .dout(n1522));
  jor  g01331(.dina(n1521), .dinb(n1435), .dout(n1523));
  jnot g01332(.din(n1523), .dout(n1524));
  jor  g01333(.dina(n1524), .dinb(n1522), .dout(n1525));
  jand g01334(.dina(n1427), .dinb(n1349), .dout(n1526));
  jnot g01335(.din(n1526), .dout(n1527));
  jnot g01336(.din(n1427), .dout(n1528));
  jand g01337(.dina(n1528), .dinb(n1350), .dout(n1529));
  jor  g01338(.dina(n1431), .dinb(n1529), .dout(n1530));
  jand g01339(.dina(n1530), .dinb(n1527), .dout(n1531));
  jxor g01340(.dina(n1531), .dinb(n1525), .dout(\asquared[27] ));
  jand g01341(.dina(n1458), .dinb(n1438), .dout(n1533));
  jand g01342(.dina(n1520), .dinb(n1459), .dout(n1534));
  jor  g01343(.dina(n1534), .dinb(n1533), .dout(n1535));
  jand g01344(.dina(n1498), .dinb(n1464), .dout(n1536));
  jand g01345(.dina(n1519), .dinb(n1499), .dout(n1537));
  jor  g01346(.dina(n1537), .dinb(n1536), .dout(n1538));
  jand g01347(.dina(n1484), .dinb(n1483), .dout(n1539));
  jand g01348(.dina(n1485), .dinb(n1482), .dout(n1540));
  jor  g01349(.dina(n1540), .dinb(n1539), .dout(n1541));
  jor  g01350(.dina(n1491), .dinb(n1489), .dout(n1542));
  jand g01351(.dina(n1542), .dinb(n1495), .dout(n1543));
  jxor g01352(.dina(n1543), .dinb(n1475), .dout(n1544));
  jxor g01353(.dina(n1544), .dinb(n1541), .dout(n1545));
  jand g01354(.dina(n1505), .dinb(n1502), .dout(n1546));
  jand g01355(.dina(n1518), .dinb(n1506), .dout(n1547));
  jor  g01356(.dina(n1547), .dinb(n1546), .dout(n1548));
  jxor g01357(.dina(n1548), .dinb(n1545), .dout(n1549));
  jand g01358(.dina(n1446), .dinb(n979), .dout(n1550));
  jand g01359(.dina(\a[27] ), .dinb(\a[0] ), .dout(n1551));
  jxor g01360(.dina(n1551), .dinb(n1550), .dout(n1552));
  jand g01361(.dina(n599), .dinb(\a[26] ), .dout(n1553));
  jnot g01362(.din(n1553), .dout(n1554));
  jand g01363(.dina(\a[26] ), .dinb(\a[1] ), .dout(n1555));
  jor  g01364(.dina(n1555), .dinb(\a[14] ), .dout(n1556));
  jand g01365(.dina(n1556), .dinb(n1554), .dout(n1557));
  jxor g01366(.dina(n1557), .dinb(n1552), .dout(n1558));
  jand g01367(.dina(\a[24] ), .dinb(\a[3] ), .dout(n1559));
  jand g01368(.dina(\a[23] ), .dinb(\a[4] ), .dout(n1560));
  jand g01369(.dina(\a[21] ), .dinb(\a[6] ), .dout(n1561));
  jxor g01370(.dina(n1561), .dinb(n1560), .dout(n1562));
  jxor g01371(.dina(n1562), .dinb(n1559), .dout(n1563));
  jnot g01372(.din(n1563), .dout(n1564));
  jand g01373(.dina(\a[22] ), .dinb(\a[5] ), .dout(n1565));
  jnot g01374(.din(n1565), .dout(n1566));
  jand g01375(.dina(n976), .dinb(n899), .dout(n1567));
  jnot g01376(.din(n1567), .dout(n1568));
  jand g01377(.dina(\a[15] ), .dinb(\a[12] ), .dout(n1569));
  jor  g01378(.dina(n1569), .dinb(n675), .dout(n1570));
  jand g01379(.dina(n1570), .dinb(n1568), .dout(n1571));
  jxor g01380(.dina(n1571), .dinb(n1566), .dout(n1572));
  jxor g01381(.dina(n1572), .dinb(n1564), .dout(n1573));
  jxor g01382(.dina(n1573), .dinb(n1558), .dout(n1574));
  jxor g01383(.dina(n1574), .dinb(n1549), .dout(n1575));
  jxor g01384(.dina(n1575), .dinb(n1538), .dout(n1576));
  jand g01385(.dina(n1456), .dinb(n1445), .dout(n1577));
  jand g01386(.dina(n1457), .dinb(n1441), .dout(n1578));
  jor  g01387(.dina(n1578), .dinb(n1577), .dout(n1579));
  jand g01388(.dina(\a[16] ), .dinb(\a[11] ), .dout(n1580));
  jand g01389(.dina(\a[25] ), .dinb(\a[20] ), .dout(n1581));
  jand g01390(.dina(n1581), .dinb(n268), .dout(n1582));
  jnot g01391(.din(n1582), .dout(n1583));
  jand g01392(.dina(\a[20] ), .dinb(\a[7] ), .dout(n1584));
  jor  g01393(.dina(n1584), .dinb(n1357), .dout(n1585));
  jand g01394(.dina(n1585), .dinb(n1583), .dout(n1586));
  jxor g01395(.dina(n1586), .dinb(n1580), .dout(n1587));
  jnot g01396(.din(n1514), .dout(n1588));
  jnot g01397(.din(n1515), .dout(n1589));
  jand g01398(.dina(n1589), .dinb(n1588), .dout(n1590));
  jnot g01399(.din(n1590), .dout(n1591));
  jand g01400(.dina(n1515), .dinb(n1514), .dout(n1592));
  jor  g01401(.dina(n1592), .dinb(n1513), .dout(n1593));
  jand g01402(.dina(n1593), .dinb(n1591), .dout(n1594));
  jxor g01403(.dina(n1594), .dinb(n1587), .dout(n1595));
  jnot g01404(.din(n1595), .dout(n1596));
  jand g01405(.dina(\a[19] ), .dinb(\a[8] ), .dout(n1597));
  jnot g01406(.din(n1597), .dout(n1598));
  jand g01407(.dina(n1107), .dinb(n453), .dout(n1599));
  jnot g01408(.din(n1599), .dout(n1600));
  jand g01409(.dina(\a[17] ), .dinb(\a[10] ), .dout(n1601));
  jand g01410(.dina(n1601), .dinb(n1597), .dout(n1602));
  jand g01411(.dina(n1024), .dinb(n395), .dout(n1603));
  jor  g01412(.dina(n1603), .dinb(n1602), .dout(n1604));
  jand g01413(.dina(n1604), .dinb(n1600), .dout(n1605));
  jor  g01414(.dina(n1605), .dinb(n1598), .dout(n1606));
  jor  g01415(.dina(n1604), .dinb(n1599), .dout(n1607));
  jnot g01416(.din(n1607), .dout(n1608));
  jand g01417(.dina(\a[18] ), .dinb(\a[9] ), .dout(n1609));
  jor  g01418(.dina(n1609), .dinb(n1601), .dout(n1610));
  jand g01419(.dina(n1610), .dinb(n1608), .dout(n1611));
  jnot g01420(.din(n1611), .dout(n1612));
  jand g01421(.dina(n1612), .dinb(n1606), .dout(n1613));
  jxor g01422(.dina(n1613), .dinb(n1596), .dout(n1614));
  jxor g01423(.dina(n1614), .dinb(n1579), .dout(n1615));
  jand g01424(.dina(n1451), .dinb(n1447), .dout(n1616));
  jand g01425(.dina(n1455), .dinb(n1452), .dout(n1617));
  jor  g01426(.dina(n1617), .dinb(n1616), .dout(n1618));
  jand g01427(.dina(n1511), .dinb(n1508), .dout(n1619));
  jand g01428(.dina(n1517), .dinb(n1512), .dout(n1620));
  jor  g01429(.dina(n1620), .dinb(n1619), .dout(n1621));
  jxor g01430(.dina(n1621), .dinb(n1618), .dout(n1622));
  jnot g01431(.din(n1622), .dout(n1623));
  jor  g01432(.dina(n1487), .dinb(n1481), .dout(n1624));
  jand g01433(.dina(n1497), .dinb(n1488), .dout(n1625));
  jnot g01434(.din(n1625), .dout(n1626));
  jand g01435(.dina(n1626), .dinb(n1624), .dout(n1627));
  jxor g01436(.dina(n1627), .dinb(n1623), .dout(n1628));
  jxor g01437(.dina(n1628), .dinb(n1615), .dout(n1629));
  jxor g01438(.dina(n1629), .dinb(n1576), .dout(n1630));
  jand g01439(.dina(n1630), .dinb(n1535), .dout(n1631));
  jor  g01440(.dina(n1630), .dinb(n1535), .dout(n1632));
  jnot g01441(.din(n1632), .dout(n1633));
  jor  g01442(.dina(n1633), .dinb(n1631), .dout(n1634));
  jnot g01443(.din(n1522), .dout(n1635));
  jor  g01444(.dina(n1531), .dinb(n1524), .dout(n1636));
  jand g01445(.dina(n1636), .dinb(n1635), .dout(n1637));
  jxor g01446(.dina(n1637), .dinb(n1634), .dout(\asquared[28] ));
  jand g01447(.dina(n1548), .dinb(n1545), .dout(n1639));
  jand g01448(.dina(n1574), .dinb(n1549), .dout(n1640));
  jor  g01449(.dina(n1640), .dinb(n1639), .dout(n1641));
  jand g01450(.dina(n1551), .dinb(n1550), .dout(n1642));
  jand g01451(.dina(n1557), .dinb(n1552), .dout(n1643));
  jor  g01452(.dina(n1643), .dinb(n1642), .dout(n1644));
  jnot g01453(.din(n1644), .dout(n1645));
  jand g01454(.dina(\a[20] ), .dinb(\a[8] ), .dout(n1646));
  jnot g01455(.din(n1646), .dout(n1647));
  jand g01456(.dina(\a[25] ), .dinb(\a[24] ), .dout(n1648));
  jand g01457(.dina(n1648), .dinb(n265), .dout(n1649));
  jnot g01458(.din(n1649), .dout(n1650));
  jand g01459(.dina(\a[25] ), .dinb(\a[3] ), .dout(n1651));
  jand g01460(.dina(\a[24] ), .dinb(\a[4] ), .dout(n1652));
  jor  g01461(.dina(n1652), .dinb(n1651), .dout(n1653));
  jand g01462(.dina(n1653), .dinb(n1650), .dout(n1654));
  jxor g01463(.dina(n1654), .dinb(n1647), .dout(n1655));
  jxor g01464(.dina(n1655), .dinb(n1645), .dout(n1656));
  jand g01465(.dina(\a[21] ), .dinb(\a[7] ), .dout(n1657));
  jand g01466(.dina(\a[23] ), .dinb(\a[22] ), .dout(n1658));
  jand g01467(.dina(n1658), .dinb(n339), .dout(n1659));
  jnot g01468(.din(n1659), .dout(n1660));
  jand g01469(.dina(\a[23] ), .dinb(\a[5] ), .dout(n1661));
  jand g01470(.dina(\a[22] ), .dinb(\a[6] ), .dout(n1662));
  jor  g01471(.dina(n1662), .dinb(n1661), .dout(n1663));
  jand g01472(.dina(n1663), .dinb(n1660), .dout(n1664));
  jxor g01473(.dina(n1664), .dinb(n1657), .dout(n1665));
  jxor g01474(.dina(n1665), .dinb(n1656), .dout(n1666));
  jxor g01475(.dina(n1666), .dinb(n1641), .dout(n1667));
  jor  g01476(.dina(n1572), .dinb(n1564), .dout(n1668));
  jand g01477(.dina(n1573), .dinb(n1558), .dout(n1669));
  jnot g01478(.din(n1669), .dout(n1670));
  jand g01479(.dina(n1670), .dinb(n1668), .dout(n1671));
  jnot g01480(.din(n1671), .dout(n1672));
  jand g01481(.dina(n1594), .dinb(n1587), .dout(n1673));
  jnot g01482(.din(n1673), .dout(n1674));
  jor  g01483(.dina(n1613), .dinb(n1596), .dout(n1675));
  jand g01484(.dina(n1675), .dinb(n1674), .dout(n1676));
  jand g01485(.dina(\a[27] ), .dinb(\a[1] ), .dout(n1677));
  jxor g01486(.dina(n1677), .dinb(n727), .dout(n1678));
  jxor g01487(.dina(n1678), .dinb(n1553), .dout(n1679));
  jand g01488(.dina(n1568), .dinb(n1566), .dout(n1680));
  jnot g01489(.din(n1680), .dout(n1681));
  jand g01490(.dina(n1681), .dinb(n1570), .dout(n1682));
  jxor g01491(.dina(n1682), .dinb(n1679), .dout(n1683));
  jnot g01492(.din(n1683), .dout(n1684));
  jxor g01493(.dina(n1684), .dinb(n1676), .dout(n1685));
  jxor g01494(.dina(n1685), .dinb(n1672), .dout(n1686));
  jxor g01495(.dina(n1686), .dinb(n1667), .dout(n1687));
  jnot g01496(.din(n1687), .dout(n1688));
  jand g01497(.dina(n1575), .dinb(n1538), .dout(n1689));
  jand g01498(.dina(n1629), .dinb(n1576), .dout(n1690));
  jor  g01499(.dina(n1690), .dinb(n1689), .dout(n1691));
  jand g01500(.dina(n1614), .dinb(n1579), .dout(n1692));
  jand g01501(.dina(n1628), .dinb(n1615), .dout(n1693));
  jor  g01502(.dina(n1693), .dinb(n1692), .dout(n1694));
  jand g01503(.dina(n1561), .dinb(n1560), .dout(n1695));
  jand g01504(.dina(n1562), .dinb(n1559), .dout(n1696));
  jor  g01505(.dina(n1696), .dinb(n1695), .dout(n1697));
  jxor g01506(.dina(n1697), .dinb(n1607), .dout(n1698));
  jand g01507(.dina(n1586), .dinb(n1580), .dout(n1699));
  jor  g01508(.dina(n1699), .dinb(n1582), .dout(n1700));
  jxor g01509(.dina(n1700), .dinb(n1698), .dout(n1701));
  jnot g01510(.din(n1701), .dout(n1702));
  jand g01511(.dina(n1621), .dinb(n1618), .dout(n1703));
  jnot g01512(.din(n1703), .dout(n1704));
  jor  g01513(.dina(n1627), .dinb(n1623), .dout(n1705));
  jand g01514(.dina(n1705), .dinb(n1704), .dout(n1706));
  jxor g01515(.dina(n1706), .dinb(n1702), .dout(n1707));
  jand g01516(.dina(n1543), .dinb(n1475), .dout(n1708));
  jand g01517(.dina(n1544), .dinb(n1541), .dout(n1709));
  jor  g01518(.dina(n1709), .dinb(n1708), .dout(n1710));
  jand g01519(.dina(\a[16] ), .dinb(\a[12] ), .dout(n1711));
  jand g01520(.dina(\a[28] ), .dinb(\a[0] ), .dout(n1712));
  jand g01521(.dina(n1712), .dinb(n1711), .dout(n1713));
  jnot g01522(.din(n1713), .dout(n1714));
  jand g01523(.dina(\a[17] ), .dinb(\a[11] ), .dout(n1715));
  jand g01524(.dina(n1715), .dinb(n1712), .dout(n1716));
  jand g01525(.dina(n937), .dinb(n555), .dout(n1717));
  jor  g01526(.dina(n1717), .dinb(n1716), .dout(n1718));
  jnot g01527(.din(n1718), .dout(n1719));
  jand g01528(.dina(n1719), .dinb(n1714), .dout(n1720));
  jor  g01529(.dina(n1712), .dinb(n1711), .dout(n1721));
  jand g01530(.dina(n1721), .dinb(n1720), .dout(n1722));
  jand g01531(.dina(n1718), .dinb(n1714), .dout(n1723));
  jnot g01532(.din(n1723), .dout(n1724));
  jand g01533(.dina(n1724), .dinb(n1715), .dout(n1725));
  jor  g01534(.dina(n1725), .dinb(n1722), .dout(n1726));
  jand g01535(.dina(\a[26] ), .dinb(\a[2] ), .dout(n1727));
  jand g01536(.dina(n1024), .dinb(n453), .dout(n1728));
  jnot g01537(.din(n1728), .dout(n1729));
  jand g01538(.dina(\a[19] ), .dinb(\a[9] ), .dout(n1730));
  jand g01539(.dina(\a[18] ), .dinb(\a[10] ), .dout(n1731));
  jor  g01540(.dina(n1731), .dinb(n1730), .dout(n1732));
  jand g01541(.dina(n1732), .dinb(n1729), .dout(n1733));
  jxor g01542(.dina(n1733), .dinb(n1727), .dout(n1734));
  jxor g01543(.dina(n1734), .dinb(n1726), .dout(n1735));
  jxor g01544(.dina(n1735), .dinb(n1710), .dout(n1736));
  jxor g01545(.dina(n1736), .dinb(n1707), .dout(n1737));
  jxor g01546(.dina(n1737), .dinb(n1694), .dout(n1738));
  jxor g01547(.dina(n1738), .dinb(n1691), .dout(n1739));
  jxor g01548(.dina(n1739), .dinb(n1688), .dout(n1740));
  jnot g01549(.din(n1631), .dout(n1741));
  jor  g01550(.dina(n1637), .dinb(n1633), .dout(n1742));
  jand g01551(.dina(n1742), .dinb(n1741), .dout(n1743));
  jxor g01552(.dina(n1743), .dinb(n1740), .dout(\asquared[29] ));
  jand g01553(.dina(n1737), .dinb(n1694), .dout(n1745));
  jand g01554(.dina(n1738), .dinb(n1691), .dout(n1746));
  jor  g01555(.dina(n1746), .dinb(n1745), .dout(n1747));
  jor  g01556(.dina(n1706), .dinb(n1702), .dout(n1748));
  jand g01557(.dina(n1736), .dinb(n1707), .dout(n1749));
  jnot g01558(.din(n1749), .dout(n1750));
  jand g01559(.dina(n1750), .dinb(n1748), .dout(n1751));
  jor  g01560(.dina(n1684), .dinb(n1676), .dout(n1752));
  jand g01561(.dina(n1685), .dinb(n1672), .dout(n1753));
  jnot g01562(.din(n1753), .dout(n1754));
  jand g01563(.dina(n1754), .dinb(n1752), .dout(n1755));
  jxor g01564(.dina(n1755), .dinb(n1751), .dout(n1756));
  jand g01565(.dina(n1734), .dinb(n1726), .dout(n1757));
  jand g01566(.dina(n1735), .dinb(n1710), .dout(n1758));
  jor  g01567(.dina(n1758), .dinb(n1757), .dout(n1759));
  jor  g01568(.dina(n1655), .dinb(n1645), .dout(n1760));
  jand g01569(.dina(n1665), .dinb(n1656), .dout(n1761));
  jnot g01570(.din(n1761), .dout(n1762));
  jand g01571(.dina(n1762), .dinb(n1760), .dout(n1763));
  jnot g01572(.din(n1763), .dout(n1764));
  jxor g01573(.dina(n1764), .dinb(n1759), .dout(n1765));
  jnot g01574(.din(n1720), .dout(n1766));
  jor  g01575(.dina(n1728), .dinb(n1727), .dout(n1767));
  jand g01576(.dina(n1767), .dinb(n1732), .dout(n1768));
  jxor g01577(.dina(n1768), .dinb(n1766), .dout(n1769));
  jand g01578(.dina(n1677), .dinb(n727), .dout(n1770));
  jnot g01579(.din(n1770), .dout(n1771));
  jand g01580(.dina(\a[29] ), .dinb(\a[2] ), .dout(n1772));
  jand g01581(.dina(n1772), .dinb(n1551), .dout(n1773));
  jnot g01582(.din(n1773), .dout(n1774));
  jand g01583(.dina(\a[29] ), .dinb(\a[0] ), .dout(n1775));
  jand g01584(.dina(\a[27] ), .dinb(\a[2] ), .dout(n1776));
  jor  g01585(.dina(n1776), .dinb(n1775), .dout(n1777));
  jand g01586(.dina(n1777), .dinb(n1774), .dout(n1778));
  jxor g01587(.dina(n1778), .dinb(n1771), .dout(n1779));
  jnot g01588(.din(n1779), .dout(n1780));
  jxor g01589(.dina(n1780), .dinb(n1769), .dout(n1781));
  jxor g01590(.dina(n1781), .dinb(n1765), .dout(n1782));
  jxor g01591(.dina(n1782), .dinb(n1756), .dout(n1783));
  jand g01592(.dina(n1666), .dinb(n1641), .dout(n1784));
  jand g01593(.dina(n1686), .dinb(n1667), .dout(n1785));
  jor  g01594(.dina(n1785), .dinb(n1784), .dout(n1786));
  jand g01595(.dina(n1697), .dinb(n1607), .dout(n1787));
  jand g01596(.dina(n1700), .dinb(n1698), .dout(n1788));
  jor  g01597(.dina(n1788), .dinb(n1787), .dout(n1789));
  jand g01598(.dina(n1678), .dinb(n1553), .dout(n1790));
  jand g01599(.dina(n1682), .dinb(n1679), .dout(n1791));
  jor  g01600(.dina(n1791), .dinb(n1790), .dout(n1792));
  jand g01601(.dina(\a[23] ), .dinb(\a[6] ), .dout(n1793));
  jand g01602(.dina(\a[16] ), .dinb(\a[13] ), .dout(n1794));
  jxor g01603(.dina(n1794), .dinb(n976), .dout(n1795));
  jxor g01604(.dina(n1795), .dinb(n1793), .dout(n1796));
  jxor g01605(.dina(n1796), .dinb(n1792), .dout(n1797));
  jxor g01606(.dina(n1797), .dinb(n1789), .dout(n1798));
  jand g01607(.dina(n1663), .dinb(n1657), .dout(n1799));
  jor  g01608(.dina(n1799), .dinb(n1659), .dout(n1800));
  jand g01609(.dina(n685), .dinb(\a[28] ), .dout(n1801));
  jnot g01610(.din(\a[15] ), .dout(n1802));
  jand g01611(.dina(\a[28] ), .dinb(\a[1] ), .dout(n1803));
  jnot g01612(.din(n1803), .dout(n1804));
  jand g01613(.dina(n1804), .dinb(n1802), .dout(n1805));
  jor  g01614(.dina(n1805), .dinb(n1801), .dout(n1806));
  jnot g01615(.din(n1806), .dout(n1807));
  jxor g01616(.dina(n1807), .dinb(n1800), .dout(n1808));
  jand g01617(.dina(n1650), .dinb(n1647), .dout(n1809));
  jnot g01618(.din(n1809), .dout(n1810));
  jand g01619(.dina(n1810), .dinb(n1653), .dout(n1811));
  jxor g01620(.dina(n1811), .dinb(n1808), .dout(n1812));
  jand g01621(.dina(\a[25] ), .dinb(\a[4] ), .dout(n1813));
  jand g01622(.dina(\a[24] ), .dinb(\a[22] ), .dout(n1814));
  jand g01623(.dina(n1814), .dinb(n431), .dout(n1815));
  jnot g01624(.din(n1815), .dout(n1816));
  jand g01625(.dina(n1648), .dinb(n242), .dout(n1817));
  jand g01626(.dina(\a[22] ), .dinb(\a[7] ), .dout(n1818));
  jand g01627(.dina(n1818), .dinb(n1813), .dout(n1819));
  jor  g01628(.dina(n1819), .dinb(n1817), .dout(n1820));
  jand g01629(.dina(n1820), .dinb(n1816), .dout(n1821));
  jnot g01630(.din(n1821), .dout(n1822));
  jand g01631(.dina(n1822), .dinb(n1813), .dout(n1823));
  jor  g01632(.dina(n1820), .dinb(n1815), .dout(n1824));
  jnot g01633(.din(n1824), .dout(n1825));
  jand g01634(.dina(\a[24] ), .dinb(\a[5] ), .dout(n1826));
  jor  g01635(.dina(n1826), .dinb(n1818), .dout(n1827));
  jand g01636(.dina(n1827), .dinb(n1825), .dout(n1828));
  jor  g01637(.dina(n1828), .dinb(n1823), .dout(n1829));
  jand g01638(.dina(\a[17] ), .dinb(\a[12] ), .dout(n1830));
  jand g01639(.dina(\a[26] ), .dinb(\a[3] ), .dout(n1831));
  jand g01640(.dina(\a[21] ), .dinb(\a[8] ), .dout(n1832));
  jor  g01641(.dina(n1832), .dinb(n1831), .dout(n1833));
  jand g01642(.dina(\a[26] ), .dinb(\a[21] ), .dout(n1834));
  jand g01643(.dina(n1834), .dinb(n399), .dout(n1835));
  jnot g01644(.din(n1835), .dout(n1836));
  jand g01645(.dina(n1836), .dinb(n1833), .dout(n1837));
  jxor g01646(.dina(n1837), .dinb(n1830), .dout(n1838));
  jnot g01647(.din(n1838), .dout(n1839));
  jand g01648(.dina(\a[20] ), .dinb(\a[9] ), .dout(n1840));
  jnot g01649(.din(n1840), .dout(n1841));
  jand g01650(.dina(n1024), .dinb(n655), .dout(n1842));
  jnot g01651(.din(n1842), .dout(n1843));
  jand g01652(.dina(\a[18] ), .dinb(\a[11] ), .dout(n1844));
  jand g01653(.dina(\a[19] ), .dinb(\a[10] ), .dout(n1845));
  jor  g01654(.dina(n1845), .dinb(n1844), .dout(n1846));
  jand g01655(.dina(n1846), .dinb(n1843), .dout(n1847));
  jxor g01656(.dina(n1847), .dinb(n1841), .dout(n1848));
  jxor g01657(.dina(n1848), .dinb(n1839), .dout(n1849));
  jxor g01658(.dina(n1849), .dinb(n1829), .dout(n1850));
  jxor g01659(.dina(n1850), .dinb(n1812), .dout(n1851));
  jxor g01660(.dina(n1851), .dinb(n1798), .dout(n1852));
  jxor g01661(.dina(n1852), .dinb(n1786), .dout(n1853));
  jxor g01662(.dina(n1853), .dinb(n1783), .dout(n1854));
  jand g01663(.dina(n1854), .dinb(n1747), .dout(n1855));
  jor  g01664(.dina(n1854), .dinb(n1747), .dout(n1856));
  jnot g01665(.din(n1856), .dout(n1857));
  jor  g01666(.dina(n1857), .dinb(n1855), .dout(n1858));
  jand g01667(.dina(n1739), .dinb(n1687), .dout(n1859));
  jnot g01668(.din(n1859), .dout(n1860));
  jnot g01669(.din(n1739), .dout(n1861));
  jand g01670(.dina(n1861), .dinb(n1688), .dout(n1862));
  jor  g01671(.dina(n1743), .dinb(n1862), .dout(n1863));
  jand g01672(.dina(n1863), .dinb(n1860), .dout(n1864));
  jxor g01673(.dina(n1864), .dinb(n1858), .dout(\asquared[30] ));
  jand g01674(.dina(n1852), .dinb(n1786), .dout(n1866));
  jand g01675(.dina(n1853), .dinb(n1783), .dout(n1867));
  jor  g01676(.dina(n1867), .dinb(n1866), .dout(n1868));
  jand g01677(.dina(n1807), .dinb(n1800), .dout(n1869));
  jand g01678(.dina(n1811), .dinb(n1808), .dout(n1870));
  jor  g01679(.dina(n1870), .dinb(n1869), .dout(n1871));
  jand g01680(.dina(\a[30] ), .dinb(\a[0] ), .dout(n1872));
  jxor g01681(.dina(n1872), .dinb(n1801), .dout(n1873));
  jand g01682(.dina(\a[16] ), .dinb(\a[14] ), .dout(n1874));
  jand g01683(.dina(\a[29] ), .dinb(\a[1] ), .dout(n1875));
  jxor g01684(.dina(n1875), .dinb(n1874), .dout(n1876));
  jxor g01685(.dina(n1876), .dinb(n1873), .dout(n1877));
  jxor g01686(.dina(n1877), .dinb(n1871), .dout(n1878));
  jand g01687(.dina(n1768), .dinb(n1766), .dout(n1879));
  jand g01688(.dina(n1780), .dinb(n1769), .dout(n1880));
  jor  g01689(.dina(n1880), .dinb(n1879), .dout(n1881));
  jxor g01690(.dina(n1881), .dinb(n1878), .dout(n1882));
  jand g01691(.dina(n1850), .dinb(n1812), .dout(n1883));
  jand g01692(.dina(n1851), .dinb(n1798), .dout(n1884));
  jor  g01693(.dina(n1884), .dinb(n1883), .dout(n1885));
  jxor g01694(.dina(n1885), .dinb(n1882), .dout(n1886));
  jor  g01695(.dina(n1848), .dinb(n1839), .dout(n1887));
  jand g01696(.dina(n1849), .dinb(n1829), .dout(n1888));
  jnot g01697(.din(n1888), .dout(n1889));
  jand g01698(.dina(n1889), .dinb(n1887), .dout(n1890));
  jand g01699(.dina(n1794), .dinb(n976), .dout(n1891));
  jand g01700(.dina(n1795), .dinb(n1793), .dout(n1892));
  jor  g01701(.dina(n1892), .dinb(n1891), .dout(n1893));
  jxor g01702(.dina(n1893), .dinb(n1824), .dout(n1894));
  jand g01703(.dina(\a[17] ), .dinb(\a[13] ), .dout(n1895));
  jand g01704(.dina(\a[28] ), .dinb(\a[2] ), .dout(n1896));
  jand g01705(.dina(\a[21] ), .dinb(\a[9] ), .dout(n1897));
  jxor g01706(.dina(n1897), .dinb(n1896), .dout(n1898));
  jxor g01707(.dina(n1898), .dinb(n1895), .dout(n1899));
  jxor g01708(.dina(n1899), .dinb(n1894), .dout(n1900));
  jnot g01709(.din(n1900), .dout(n1901));
  jxor g01710(.dina(n1901), .dinb(n1890), .dout(n1902));
  jand g01711(.dina(n1837), .dinb(n1830), .dout(n1903));
  jor  g01712(.dina(n1903), .dinb(n1835), .dout(n1904));
  jand g01713(.dina(n1843), .dinb(n1841), .dout(n1905));
  jnot g01714(.din(n1905), .dout(n1906));
  jand g01715(.dina(n1906), .dinb(n1846), .dout(n1907));
  jxor g01716(.dina(n1907), .dinb(n1904), .dout(n1908));
  jand g01717(.dina(n1774), .dinb(n1771), .dout(n1909));
  jnot g01718(.din(n1909), .dout(n1910));
  jand g01719(.dina(n1910), .dinb(n1777), .dout(n1911));
  jxor g01720(.dina(n1911), .dinb(n1908), .dout(n1912));
  jxor g01721(.dina(n1912), .dinb(n1902), .dout(n1913));
  jxor g01722(.dina(n1913), .dinb(n1886), .dout(n1914));
  jor  g01723(.dina(n1755), .dinb(n1751), .dout(n1915));
  jand g01724(.dina(n1782), .dinb(n1756), .dout(n1916));
  jnot g01725(.din(n1916), .dout(n1917));
  jand g01726(.dina(n1917), .dinb(n1915), .dout(n1918));
  jnot g01727(.din(n1918), .dout(n1919));
  jand g01728(.dina(n1796), .dinb(n1792), .dout(n1920));
  jand g01729(.dina(n1797), .dinb(n1789), .dout(n1921));
  jor  g01730(.dina(n1921), .dinb(n1920), .dout(n1922));
  jand g01731(.dina(\a[26] ), .dinb(\a[4] ), .dout(n1923));
  jand g01732(.dina(\a[22] ), .dinb(\a[8] ), .dout(n1924));
  jand g01733(.dina(n1924), .dinb(n1923), .dout(n1925));
  jnot g01734(.din(n1925), .dout(n1926));
  jand g01735(.dina(\a[27] ), .dinb(\a[26] ), .dout(n1927));
  jand g01736(.dina(n1927), .dinb(n265), .dout(n1928));
  jand g01737(.dina(\a[27] ), .dinb(\a[3] ), .dout(n1929));
  jand g01738(.dina(n1929), .dinb(n1924), .dout(n1930));
  jor  g01739(.dina(n1930), .dinb(n1928), .dout(n1931));
  jnot g01740(.din(n1931), .dout(n1932));
  jand g01741(.dina(n1932), .dinb(n1926), .dout(n1933));
  jor  g01742(.dina(n1924), .dinb(n1923), .dout(n1934));
  jand g01743(.dina(n1934), .dinb(n1933), .dout(n1935));
  jand g01744(.dina(n1931), .dinb(n1926), .dout(n1936));
  jnot g01745(.din(n1936), .dout(n1937));
  jand g01746(.dina(n1937), .dinb(n1929), .dout(n1938));
  jor  g01747(.dina(n1938), .dinb(n1935), .dout(n1939));
  jand g01748(.dina(\a[25] ), .dinb(\a[5] ), .dout(n1940));
  jnot g01749(.din(n1940), .dout(n1941));
  jand g01750(.dina(\a[24] ), .dinb(\a[23] ), .dout(n1942));
  jand g01751(.dina(n1942), .dinb(n410), .dout(n1943));
  jnot g01752(.din(n1943), .dout(n1944));
  jand g01753(.dina(\a[24] ), .dinb(\a[6] ), .dout(n1945));
  jand g01754(.dina(\a[23] ), .dinb(\a[7] ), .dout(n1946));
  jor  g01755(.dina(n1946), .dinb(n1945), .dout(n1947));
  jand g01756(.dina(n1947), .dinb(n1944), .dout(n1948));
  jxor g01757(.dina(n1948), .dinb(n1941), .dout(n1949));
  jnot g01758(.din(n1949), .dout(n1950));
  jxor g01759(.dina(n1950), .dinb(n1939), .dout(n1951));
  jnot g01760(.din(n1951), .dout(n1952));
  jand g01761(.dina(\a[20] ), .dinb(\a[10] ), .dout(n1953));
  jnot g01762(.din(n1953), .dout(n1954));
  jand g01763(.dina(n1024), .dinb(n555), .dout(n1955));
  jnot g01764(.din(n1955), .dout(n1956));
  jand g01765(.dina(\a[19] ), .dinb(\a[11] ), .dout(n1957));
  jand g01766(.dina(\a[18] ), .dinb(\a[12] ), .dout(n1958));
  jor  g01767(.dina(n1958), .dinb(n1957), .dout(n1959));
  jand g01768(.dina(n1959), .dinb(n1956), .dout(n1960));
  jxor g01769(.dina(n1960), .dinb(n1954), .dout(n1961));
  jxor g01770(.dina(n1961), .dinb(n1952), .dout(n1962));
  jxor g01771(.dina(n1962), .dinb(n1922), .dout(n1963));
  jand g01772(.dina(n1764), .dinb(n1759), .dout(n1964));
  jand g01773(.dina(n1781), .dinb(n1765), .dout(n1965));
  jor  g01774(.dina(n1965), .dinb(n1964), .dout(n1966));
  jxor g01775(.dina(n1966), .dinb(n1963), .dout(n1967));
  jxor g01776(.dina(n1967), .dinb(n1919), .dout(n1968));
  jxor g01777(.dina(n1968), .dinb(n1914), .dout(n1969));
  jand g01778(.dina(n1969), .dinb(n1868), .dout(n1970));
  jor  g01779(.dina(n1969), .dinb(n1868), .dout(n1971));
  jnot g01780(.din(n1971), .dout(n1972));
  jor  g01781(.dina(n1972), .dinb(n1970), .dout(n1973));
  jnot g01782(.din(n1855), .dout(n1974));
  jor  g01783(.dina(n1864), .dinb(n1857), .dout(n1975));
  jand g01784(.dina(n1975), .dinb(n1974), .dout(n1976));
  jxor g01785(.dina(n1976), .dinb(n1973), .dout(\asquared[31] ));
  jand g01786(.dina(n1967), .dinb(n1919), .dout(n1978));
  jand g01787(.dina(n1968), .dinb(n1914), .dout(n1979));
  jor  g01788(.dina(n1979), .dinb(n1978), .dout(n1980));
  jand g01789(.dina(n1885), .dinb(n1882), .dout(n1981));
  jand g01790(.dina(n1913), .dinb(n1886), .dout(n1982));
  jor  g01791(.dina(n1982), .dinb(n1981), .dout(n1983));
  jor  g01792(.dina(n1901), .dinb(n1890), .dout(n1984));
  jand g01793(.dina(n1912), .dinb(n1902), .dout(n1985));
  jnot g01794(.din(n1985), .dout(n1986));
  jand g01795(.dina(n1986), .dinb(n1984), .dout(n1987));
  jnot g01796(.din(n1987), .dout(n1988));
  jand g01797(.dina(\a[31] ), .dinb(\a[22] ), .dout(n1989));
  jand g01798(.dina(n1989), .dinb(n329), .dout(n1990));
  jnot g01799(.din(n1990), .dout(n1991));
  jand g01800(.dina(\a[31] ), .dinb(\a[0] ), .dout(n1992));
  jand g01801(.dina(\a[21] ), .dinb(\a[10] ), .dout(n1993));
  jand g01802(.dina(n1993), .dinb(n1992), .dout(n1994));
  jand g01803(.dina(n1376), .dinb(n453), .dout(n1995));
  jor  g01804(.dina(n1995), .dinb(n1994), .dout(n1996));
  jnot g01805(.din(n1996), .dout(n1997));
  jand g01806(.dina(n1997), .dinb(n1991), .dout(n1998));
  jand g01807(.dina(\a[22] ), .dinb(\a[9] ), .dout(n1999));
  jor  g01808(.dina(n1999), .dinb(n1992), .dout(n2000));
  jand g01809(.dina(n2000), .dinb(n1998), .dout(n2001));
  jand g01810(.dina(n1996), .dinb(n1991), .dout(n2002));
  jnot g01811(.din(n2002), .dout(n2003));
  jand g01812(.dina(n2003), .dinb(n1993), .dout(n2004));
  jor  g01813(.dina(n2004), .dinb(n2001), .dout(n2005));
  jand g01814(.dina(n1872), .dinb(n1801), .dout(n2006));
  jand g01815(.dina(n1876), .dinb(n1873), .dout(n2007));
  jor  g01816(.dina(n2007), .dinb(n2006), .dout(n2008));
  jnot g01817(.din(n2008), .dout(n2009));
  jand g01818(.dina(\a[20] ), .dinb(\a[11] ), .dout(n2010));
  jnot g01819(.din(n2010), .dout(n2011));
  jand g01820(.dina(n1024), .dinb(n899), .dout(n2012));
  jnot g01821(.din(n2012), .dout(n2013));
  jand g01822(.dina(\a[18] ), .dinb(\a[13] ), .dout(n2014));
  jand g01823(.dina(\a[19] ), .dinb(\a[12] ), .dout(n2015));
  jor  g01824(.dina(n2015), .dinb(n2014), .dout(n2016));
  jand g01825(.dina(n2016), .dinb(n2013), .dout(n2017));
  jxor g01826(.dina(n2017), .dinb(n2011), .dout(n2018));
  jxor g01827(.dina(n2018), .dinb(n2009), .dout(n2019));
  jxor g01828(.dina(n2019), .dinb(n2005), .dout(n2020));
  jand g01829(.dina(\a[23] ), .dinb(\a[8] ), .dout(n2021));
  jand g01830(.dina(\a[26] ), .dinb(\a[24] ), .dout(n2022));
  jand g01831(.dina(n2022), .dinb(n431), .dout(n2023));
  jnot g01832(.din(n2023), .dout(n2024));
  jand g01833(.dina(\a[26] ), .dinb(\a[5] ), .dout(n2025));
  jand g01834(.dina(\a[24] ), .dinb(\a[7] ), .dout(n2026));
  jor  g01835(.dina(n2026), .dinb(n2025), .dout(n2027));
  jand g01836(.dina(n2027), .dinb(n2024), .dout(n2028));
  jxor g01837(.dina(n2028), .dinb(n2021), .dout(n2029));
  jnot g01838(.din(n2029), .dout(n2030));
  jand g01839(.dina(\a[25] ), .dinb(\a[6] ), .dout(n2031));
  jnot g01840(.din(n2031), .dout(n2032));
  jand g01841(.dina(n976), .dinb(n937), .dout(n2033));
  jnot g01842(.din(n2033), .dout(n2034));
  jand g01843(.dina(\a[17] ), .dinb(\a[14] ), .dout(n2035));
  jor  g01844(.dina(n2035), .dinb(n829), .dout(n2036));
  jand g01845(.dina(n2036), .dinb(n2034), .dout(n2037));
  jxor g01846(.dina(n2037), .dinb(n2032), .dout(n2038));
  jxor g01847(.dina(n2038), .dinb(n2030), .dout(n2039));
  jnot g01848(.din(n2039), .dout(n2040));
  jnot g01849(.din(n1772), .dout(n2041));
  jand g01850(.dina(\a[28] ), .dinb(\a[27] ), .dout(n2042));
  jand g01851(.dina(n2042), .dinb(n265), .dout(n2043));
  jnot g01852(.din(n2043), .dout(n2044));
  jand g01853(.dina(\a[28] ), .dinb(\a[3] ), .dout(n2045));
  jand g01854(.dina(\a[27] ), .dinb(\a[4] ), .dout(n2046));
  jor  g01855(.dina(n2046), .dinb(n2045), .dout(n2047));
  jand g01856(.dina(n2047), .dinb(n2044), .dout(n2048));
  jxor g01857(.dina(n2048), .dinb(n2041), .dout(n2049));
  jxor g01858(.dina(n2049), .dinb(n2040), .dout(n2050));
  jxor g01859(.dina(n2050), .dinb(n2020), .dout(n2051));
  jxor g01860(.dina(n2051), .dinb(n1988), .dout(n2052));
  jxor g01861(.dina(n2052), .dinb(n1983), .dout(n2053));
  jand g01862(.dina(n1962), .dinb(n1922), .dout(n2054));
  jand g01863(.dina(n1966), .dinb(n1963), .dout(n2055));
  jor  g01864(.dina(n2055), .dinb(n2054), .dout(n2056));
  jand g01865(.dina(n1893), .dinb(n1824), .dout(n2057));
  jand g01866(.dina(n1899), .dinb(n1894), .dout(n2058));
  jor  g01867(.dina(n2058), .dinb(n2057), .dout(n2059));
  jand g01868(.dina(n1907), .dinb(n1904), .dout(n2060));
  jand g01869(.dina(n1911), .dinb(n1908), .dout(n2061));
  jor  g01870(.dina(n2061), .dinb(n2060), .dout(n2062));
  jxor g01871(.dina(n2062), .dinb(n2059), .dout(n2063));
  jand g01872(.dina(\a[30] ), .dinb(\a[1] ), .dout(n2064));
  jnot g01873(.din(n2064), .dout(n2065));
  jnot g01874(.din(\a[16] ), .dout(n2066));
  jand g01875(.dina(n1875), .dinb(n1874), .dout(n2067));
  jor  g01876(.dina(n2067), .dinb(n2066), .dout(n2068));
  jxor g01877(.dina(n2068), .dinb(n2065), .dout(n2069));
  jand g01878(.dina(n1944), .dinb(n1941), .dout(n2070));
  jnot g01879(.din(n2070), .dout(n2071));
  jand g01880(.dina(n2071), .dinb(n1947), .dout(n2072));
  jxor g01881(.dina(n2072), .dinb(n2069), .dout(n2073));
  jxor g01882(.dina(n2073), .dinb(n2063), .dout(n2074));
  jxor g01883(.dina(n2074), .dinb(n2056), .dout(n2075));
  jnot g01884(.din(n1933), .dout(n2076));
  jand g01885(.dina(n1897), .dinb(n1896), .dout(n2077));
  jand g01886(.dina(n1898), .dinb(n1895), .dout(n2078));
  jor  g01887(.dina(n2078), .dinb(n2077), .dout(n2079));
  jxor g01888(.dina(n2079), .dinb(n2076), .dout(n2080));
  jand g01889(.dina(n1956), .dinb(n1954), .dout(n2081));
  jnot g01890(.din(n2081), .dout(n2082));
  jand g01891(.dina(n2082), .dinb(n1959), .dout(n2083));
  jxor g01892(.dina(n2083), .dinb(n2080), .dout(n2084));
  jnot g01893(.din(n2084), .dout(n2085));
  jand g01894(.dina(n1950), .dinb(n1939), .dout(n2086));
  jnot g01895(.din(n2086), .dout(n2087));
  jor  g01896(.dina(n1961), .dinb(n1952), .dout(n2088));
  jand g01897(.dina(n2088), .dinb(n2087), .dout(n2089));
  jxor g01898(.dina(n2089), .dinb(n2085), .dout(n2090));
  jand g01899(.dina(n1877), .dinb(n1871), .dout(n2091));
  jand g01900(.dina(n1881), .dinb(n1878), .dout(n2092));
  jor  g01901(.dina(n2092), .dinb(n2091), .dout(n2093));
  jxor g01902(.dina(n2093), .dinb(n2090), .dout(n2094));
  jxor g01903(.dina(n2094), .dinb(n2075), .dout(n2095));
  jxor g01904(.dina(n2095), .dinb(n2053), .dout(n2096));
  jand g01905(.dina(n2096), .dinb(n1980), .dout(n2097));
  jor  g01906(.dina(n2096), .dinb(n1980), .dout(n2098));
  jnot g01907(.din(n2098), .dout(n2099));
  jor  g01908(.dina(n2099), .dinb(n2097), .dout(n2100));
  jnot g01909(.din(n1970), .dout(n2101));
  jor  g01910(.dina(n1976), .dinb(n1972), .dout(n2102));
  jand g01911(.dina(n2102), .dinb(n2101), .dout(n2103));
  jxor g01912(.dina(n2103), .dinb(n2100), .dout(\asquared[32] ));
  jand g01913(.dina(n2052), .dinb(n1983), .dout(n2105));
  jand g01914(.dina(n2095), .dinb(n2053), .dout(n2106));
  jor  g01915(.dina(n2106), .dinb(n2105), .dout(n2107));
  jand g01916(.dina(n2074), .dinb(n2056), .dout(n2108));
  jand g01917(.dina(n2094), .dinb(n2075), .dout(n2109));
  jor  g01918(.dina(n2109), .dinb(n2108), .dout(n2110));
  jor  g01919(.dina(n2089), .dinb(n2085), .dout(n2111));
  jand g01920(.dina(n2093), .dinb(n2090), .dout(n2112));
  jnot g01921(.din(n2112), .dout(n2113));
  jand g01922(.dina(n2113), .dinb(n2111), .dout(n2114));
  jnot g01923(.din(n2114), .dout(n2115));
  jand g01924(.dina(n2072), .dinb(n2069), .dout(n2116));
  jand g01925(.dina(n2065), .dinb(n2067), .dout(n2117));
  jor  g01926(.dina(n2117), .dinb(n2116), .dout(n2118));
  jand g01927(.dina(\a[23] ), .dinb(\a[9] ), .dout(n2119));
  jand g01928(.dina(\a[27] ), .dinb(\a[5] ), .dout(n2120));
  jand g01929(.dina(\a[28] ), .dinb(\a[4] ), .dout(n2121));
  jor  g01930(.dina(n2121), .dinb(n2120), .dout(n2122));
  jand g01931(.dina(n2042), .dinb(n242), .dout(n2123));
  jnot g01932(.din(n2123), .dout(n2124));
  jand g01933(.dina(n2124), .dinb(n2122), .dout(n2125));
  jxor g01934(.dina(n2125), .dinb(n2119), .dout(n2126));
  jand g01935(.dina(\a[24] ), .dinb(\a[8] ), .dout(n2127));
  jand g01936(.dina(\a[26] ), .dinb(\a[25] ), .dout(n2128));
  jand g01937(.dina(n2128), .dinb(n410), .dout(n2129));
  jnot g01938(.din(n2129), .dout(n2130));
  jand g01939(.dina(\a[26] ), .dinb(\a[6] ), .dout(n2131));
  jand g01940(.dina(\a[25] ), .dinb(\a[7] ), .dout(n2132));
  jor  g01941(.dina(n2132), .dinb(n2131), .dout(n2133));
  jand g01942(.dina(n2133), .dinb(n2130), .dout(n2134));
  jxor g01943(.dina(n2134), .dinb(n2127), .dout(n2135));
  jxor g01944(.dina(n2135), .dinb(n2126), .dout(n2136));
  jxor g01945(.dina(n2136), .dinb(n2118), .dout(n2137));
  jand g01946(.dina(n2064), .dinb(\a[16] ), .dout(n2138));
  jand g01947(.dina(\a[32] ), .dinb(\a[0] ), .dout(n2139));
  jand g01948(.dina(\a[30] ), .dinb(\a[2] ), .dout(n2140));
  jor  g01949(.dina(n2140), .dinb(n2139), .dout(n2141));
  jand g01950(.dina(\a[32] ), .dinb(\a[2] ), .dout(n2142));
  jand g01951(.dina(n2142), .dinb(n1872), .dout(n2143));
  jnot g01952(.din(n2143), .dout(n2144));
  jand g01953(.dina(n2144), .dinb(n2141), .dout(n2145));
  jxor g01954(.dina(n2145), .dinb(n2138), .dout(n2146));
  jand g01955(.dina(\a[21] ), .dinb(\a[11] ), .dout(n2147));
  jand g01956(.dina(n1287), .dinb(n899), .dout(n2148));
  jnot g01957(.din(n2148), .dout(n2149));
  jand g01958(.dina(\a[20] ), .dinb(\a[12] ), .dout(n2150));
  jand g01959(.dina(\a[19] ), .dinb(\a[13] ), .dout(n2151));
  jor  g01960(.dina(n2151), .dinb(n2150), .dout(n2152));
  jand g01961(.dina(n2152), .dinb(n2149), .dout(n2153));
  jxor g01962(.dina(n2153), .dinb(n2147), .dout(n2154));
  jxor g01963(.dina(n2154), .dinb(n2146), .dout(n2155));
  jand g01964(.dina(\a[18] ), .dinb(\a[14] ), .dout(n2156));
  jand g01965(.dina(\a[29] ), .dinb(\a[3] ), .dout(n2157));
  jand g01966(.dina(\a[22] ), .dinb(\a[10] ), .dout(n2158));
  jxor g01967(.dina(n2158), .dinb(n2157), .dout(n2159));
  jxor g01968(.dina(n2159), .dinb(n2156), .dout(n2160));
  jxor g01969(.dina(n2160), .dinb(n2155), .dout(n2161));
  jxor g01970(.dina(n2161), .dinb(n2137), .dout(n2162));
  jxor g01971(.dina(n2162), .dinb(n2115), .dout(n2163));
  jxor g01972(.dina(n2163), .dinb(n2110), .dout(n2164));
  jand g01973(.dina(n2062), .dinb(n2059), .dout(n2165));
  jand g01974(.dina(n2073), .dinb(n2063), .dout(n2166));
  jor  g01975(.dina(n2166), .dinb(n2165), .dout(n2167));
  jnot g01976(.din(n1998), .dout(n2168));
  jand g01977(.dina(n2013), .dinb(n2011), .dout(n2169));
  jnot g01978(.din(n2169), .dout(n2170));
  jand g01979(.dina(n2170), .dinb(n2016), .dout(n2171));
  jxor g01980(.dina(n2171), .dinb(n2168), .dout(n2172));
  jand g01981(.dina(n2044), .dinb(n2041), .dout(n2173));
  jnot g01982(.din(n2173), .dout(n2174));
  jand g01983(.dina(n2174), .dinb(n2047), .dout(n2175));
  jxor g01984(.dina(n2175), .dinb(n2172), .dout(n2176));
  jand g01985(.dina(n2028), .dinb(n2021), .dout(n2177));
  jor  g01986(.dina(n2177), .dinb(n2023), .dout(n2178));
  jand g01987(.dina(\a[31] ), .dinb(\a[1] ), .dout(n2179));
  jxor g01988(.dina(n2179), .dinb(n878), .dout(n2180));
  jand g01989(.dina(n2034), .dinb(n2032), .dout(n2181));
  jnot g01990(.din(n2181), .dout(n2182));
  jand g01991(.dina(n2182), .dinb(n2036), .dout(n2183));
  jxor g01992(.dina(n2183), .dinb(n2180), .dout(n2184));
  jxor g01993(.dina(n2184), .dinb(n2178), .dout(n2185));
  jxor g01994(.dina(n2185), .dinb(n2176), .dout(n2186));
  jxor g01995(.dina(n2186), .dinb(n2167), .dout(n2187));
  jor  g01996(.dina(n2018), .dinb(n2009), .dout(n2188));
  jand g01997(.dina(n2019), .dinb(n2005), .dout(n2189));
  jnot g01998(.din(n2189), .dout(n2190));
  jand g01999(.dina(n2190), .dinb(n2188), .dout(n2191));
  jand g02000(.dina(n2079), .dinb(n2076), .dout(n2192));
  jand g02001(.dina(n2083), .dinb(n2080), .dout(n2193));
  jor  g02002(.dina(n2193), .dinb(n2192), .dout(n2194));
  jnot g02003(.din(n2194), .dout(n2195));
  jxor g02004(.dina(n2195), .dinb(n2191), .dout(n2196));
  jnot g02005(.din(n2196), .dout(n2197));
  jor  g02006(.dina(n2038), .dinb(n2030), .dout(n2198));
  jor  g02007(.dina(n2049), .dinb(n2040), .dout(n2199));
  jand g02008(.dina(n2199), .dinb(n2198), .dout(n2200));
  jxor g02009(.dina(n2200), .dinb(n2197), .dout(n2201));
  jand g02010(.dina(n2050), .dinb(n2020), .dout(n2202));
  jand g02011(.dina(n2051), .dinb(n1988), .dout(n2203));
  jor  g02012(.dina(n2203), .dinb(n2202), .dout(n2204));
  jxor g02013(.dina(n2204), .dinb(n2201), .dout(n2205));
  jxor g02014(.dina(n2205), .dinb(n2187), .dout(n2206));
  jxor g02015(.dina(n2206), .dinb(n2164), .dout(n2207));
  jand g02016(.dina(n2207), .dinb(n2107), .dout(n2208));
  jor  g02017(.dina(n2207), .dinb(n2107), .dout(n2209));
  jnot g02018(.din(n2209), .dout(n2210));
  jor  g02019(.dina(n2210), .dinb(n2208), .dout(n2211));
  jnot g02020(.din(n2097), .dout(n2212));
  jor  g02021(.dina(n2103), .dinb(n2099), .dout(n2213));
  jand g02022(.dina(n2213), .dinb(n2212), .dout(n2214));
  jxor g02023(.dina(n2214), .dinb(n2211), .dout(\asquared[33] ));
  jand g02024(.dina(n2171), .dinb(n2168), .dout(n2216));
  jand g02025(.dina(n2175), .dinb(n2172), .dout(n2217));
  jor  g02026(.dina(n2217), .dinb(n2216), .dout(n2218));
  jand g02027(.dina(n2154), .dinb(n2146), .dout(n2219));
  jand g02028(.dina(n2160), .dinb(n2155), .dout(n2220));
  jor  g02029(.dina(n2220), .dinb(n2219), .dout(n2221));
  jxor g02030(.dina(n2221), .dinb(n2218), .dout(n2222));
  jand g02031(.dina(n2135), .dinb(n2126), .dout(n2223));
  jand g02032(.dina(n2136), .dinb(n2118), .dout(n2224));
  jor  g02033(.dina(n2224), .dinb(n2223), .dout(n2225));
  jxor g02034(.dina(n2225), .dinb(n2222), .dout(n2226));
  jand g02035(.dina(n2161), .dinb(n2137), .dout(n2227));
  jand g02036(.dina(n2162), .dinb(n2115), .dout(n2228));
  jor  g02037(.dina(n2228), .dinb(n2227), .dout(n2229));
  jxor g02038(.dina(n2229), .dinb(n2226), .dout(n2230));
  jand g02039(.dina(n2158), .dinb(n2157), .dout(n2231));
  jand g02040(.dina(n2159), .dinb(n2156), .dout(n2232));
  jor  g02041(.dina(n2232), .dinb(n2231), .dout(n2233));
  jand g02042(.dina(n2145), .dinb(n2138), .dout(n2234));
  jor  g02043(.dina(n2234), .dinb(n2143), .dout(n2235));
  jor  g02044(.dina(n2148), .dinb(n2147), .dout(n2236));
  jand g02045(.dina(n2236), .dinb(n2152), .dout(n2237));
  jxor g02046(.dina(n2237), .dinb(n2235), .dout(n2238));
  jxor g02047(.dina(n2238), .dinb(n2233), .dout(n2239));
  jand g02048(.dina(n2125), .dinb(n2119), .dout(n2240));
  jor  g02049(.dina(n2240), .dinb(n2123), .dout(n2241));
  jor  g02050(.dina(n2129), .dinb(n2127), .dout(n2242));
  jand g02051(.dina(n2242), .dinb(n2133), .dout(n2243));
  jxor g02052(.dina(n2243), .dinb(n2241), .dout(n2244));
  jnot g02053(.din(n2244), .dout(n2245));
  jand g02054(.dina(\a[31] ), .dinb(\a[2] ), .dout(n2246));
  jnot g02055(.din(n2246), .dout(n2247));
  jand g02056(.dina(\a[33] ), .dinb(\a[22] ), .dout(n2248));
  jand g02057(.dina(n2248), .dinb(n407), .dout(n2249));
  jnot g02058(.din(n2249), .dout(n2250));
  jand g02059(.dina(\a[33] ), .dinb(\a[0] ), .dout(n2251));
  jand g02060(.dina(\a[22] ), .dinb(\a[11] ), .dout(n2252));
  jor  g02061(.dina(n2252), .dinb(n2251), .dout(n2253));
  jand g02062(.dina(n2253), .dinb(n2250), .dout(n2254));
  jxor g02063(.dina(n2254), .dinb(n2247), .dout(n2255));
  jxor g02064(.dina(n2255), .dinb(n2245), .dout(n2256));
  jxor g02065(.dina(n2256), .dinb(n2239), .dout(n2257));
  jand g02066(.dina(\a[28] ), .dinb(\a[5] ), .dout(n2258));
  jand g02067(.dina(\a[27] ), .dinb(\a[25] ), .dout(n2259));
  jand g02068(.dina(n2259), .dinb(n544), .dout(n2260));
  jnot g02069(.din(n2260), .dout(n2261));
  jand g02070(.dina(n2042), .dinb(n339), .dout(n2262));
  jand g02071(.dina(\a[25] ), .dinb(\a[8] ), .dout(n2263));
  jand g02072(.dina(n2263), .dinb(n2258), .dout(n2264));
  jor  g02073(.dina(n2264), .dinb(n2262), .dout(n2265));
  jand g02074(.dina(n2265), .dinb(n2261), .dout(n2266));
  jnot g02075(.din(n2266), .dout(n2267));
  jand g02076(.dina(n2267), .dinb(n2258), .dout(n2268));
  jand g02077(.dina(\a[27] ), .dinb(\a[6] ), .dout(n2269));
  jor  g02078(.dina(n2269), .dinb(n2263), .dout(n2270));
  jor  g02079(.dina(n2265), .dinb(n2260), .dout(n2271));
  jnot g02080(.din(n2271), .dout(n2272));
  jand g02081(.dina(n2272), .dinb(n2270), .dout(n2273));
  jor  g02082(.dina(n2273), .dinb(n2268), .dout(n2274));
  jand g02083(.dina(\a[30] ), .dinb(\a[3] ), .dout(n2275));
  jand g02084(.dina(\a[29] ), .dinb(\a[4] ), .dout(n2276));
  jand g02085(.dina(\a[24] ), .dinb(\a[9] ), .dout(n2277));
  jxor g02086(.dina(n2277), .dinb(n2276), .dout(n2278));
  jxor g02087(.dina(n2278), .dinb(n2275), .dout(n2279));
  jxor g02088(.dina(n2279), .dinb(n2274), .dout(n2280));
  jnot g02089(.din(n2280), .dout(n2281));
  jand g02090(.dina(\a[26] ), .dinb(\a[7] ), .dout(n2282));
  jnot g02091(.din(n2282), .dout(n2283));
  jand g02092(.dina(n1107), .dinb(n829), .dout(n2284));
  jnot g02093(.din(n2284), .dout(n2285));
  jand g02094(.dina(\a[18] ), .dinb(\a[15] ), .dout(n2286));
  jor  g02095(.dina(n2286), .dinb(n937), .dout(n2287));
  jand g02096(.dina(n2287), .dinb(n2285), .dout(n2288));
  jxor g02097(.dina(n2288), .dinb(n2283), .dout(n2289));
  jxor g02098(.dina(n2289), .dinb(n2281), .dout(n2290));
  jxor g02099(.dina(n2290), .dinb(n2257), .dout(n2291));
  jxor g02100(.dina(n2291), .dinb(n2230), .dout(n2292));
  jand g02101(.dina(n2183), .dinb(n2180), .dout(n2293));
  jand g02102(.dina(n2184), .dinb(n2178), .dout(n2294));
  jor  g02103(.dina(n2294), .dinb(n2293), .dout(n2295));
  jand g02104(.dina(\a[32] ), .dinb(\a[1] ), .dout(n2296));
  jxor g02105(.dina(n2296), .dinb(\a[17] ), .dout(n2297));
  jand g02106(.dina(n2179), .dinb(n878), .dout(n2298));
  jand g02107(.dina(\a[23] ), .dinb(\a[10] ), .dout(n2299));
  jxor g02108(.dina(n2299), .dinb(n2298), .dout(n2300));
  jxor g02109(.dina(n2300), .dinb(n2297), .dout(n2301));
  jnot g02110(.din(n2301), .dout(n2302));
  jand g02111(.dina(\a[21] ), .dinb(\a[12] ), .dout(n2303));
  jnot g02112(.din(n2303), .dout(n2304));
  jand g02113(.dina(n1287), .dinb(n675), .dout(n2305));
  jnot g02114(.din(n2305), .dout(n2306));
  jand g02115(.dina(\a[20] ), .dinb(\a[13] ), .dout(n2307));
  jand g02116(.dina(\a[19] ), .dinb(\a[14] ), .dout(n2308));
  jor  g02117(.dina(n2308), .dinb(n2307), .dout(n2309));
  jand g02118(.dina(n2309), .dinb(n2306), .dout(n2310));
  jxor g02119(.dina(n2310), .dinb(n2304), .dout(n2311));
  jxor g02120(.dina(n2311), .dinb(n2302), .dout(n2312));
  jxor g02121(.dina(n2312), .dinb(n2295), .dout(n2313));
  jnot g02122(.din(n2313), .dout(n2314));
  jor  g02123(.dina(n2195), .dinb(n2191), .dout(n2315));
  jor  g02124(.dina(n2200), .dinb(n2197), .dout(n2316));
  jand g02125(.dina(n2316), .dinb(n2315), .dout(n2317));
  jxor g02126(.dina(n2317), .dinb(n2314), .dout(n2318));
  jand g02127(.dina(n2185), .dinb(n2176), .dout(n2319));
  jand g02128(.dina(n2186), .dinb(n2167), .dout(n2320));
  jor  g02129(.dina(n2320), .dinb(n2319), .dout(n2321));
  jxor g02130(.dina(n2321), .dinb(n2318), .dout(n2322));
  jand g02131(.dina(n2204), .dinb(n2201), .dout(n2323));
  jand g02132(.dina(n2205), .dinb(n2187), .dout(n2324));
  jor  g02133(.dina(n2324), .dinb(n2323), .dout(n2325));
  jxor g02134(.dina(n2325), .dinb(n2322), .dout(n2326));
  jxor g02135(.dina(n2326), .dinb(n2292), .dout(n2327));
  jnot g02136(.din(n2327), .dout(n2328));
  jand g02137(.dina(n2163), .dinb(n2110), .dout(n2329));
  jand g02138(.dina(n2206), .dinb(n2164), .dout(n2330));
  jor  g02139(.dina(n2330), .dinb(n2329), .dout(n2331));
  jxor g02140(.dina(n2331), .dinb(n2328), .dout(n2332));
  jnot g02141(.din(n2208), .dout(n2333));
  jor  g02142(.dina(n2214), .dinb(n2210), .dout(n2334));
  jand g02143(.dina(n2334), .dinb(n2333), .dout(n2335));
  jxor g02144(.dina(n2335), .dinb(n2332), .dout(\asquared[34] ));
  jand g02145(.dina(n2325), .dinb(n2322), .dout(n2337));
  jand g02146(.dina(n2326), .dinb(n2292), .dout(n2338));
  jor  g02147(.dina(n2338), .dinb(n2337), .dout(n2339));
  jor  g02148(.dina(n2317), .dinb(n2314), .dout(n2340));
  jand g02149(.dina(n2321), .dinb(n2318), .dout(n2341));
  jnot g02150(.din(n2341), .dout(n2342));
  jand g02151(.dina(n2342), .dinb(n2340), .dout(n2343));
  jnot g02152(.din(n2343), .dout(n2344));
  jand g02153(.dina(n2277), .dinb(n2276), .dout(n2345));
  jand g02154(.dina(n2278), .dinb(n2275), .dout(n2346));
  jor  g02155(.dina(n2346), .dinb(n2345), .dout(n2347));
  jand g02156(.dina(n2250), .dinb(n2247), .dout(n2348));
  jnot g02157(.din(n2348), .dout(n2349));
  jand g02158(.dina(n2349), .dinb(n2253), .dout(n2350));
  jxor g02159(.dina(n2350), .dinb(n2347), .dout(n2351));
  jxor g02160(.dina(n2351), .dinb(n2271), .dout(n2352));
  jand g02161(.dina(n2279), .dinb(n2274), .dout(n2353));
  jnot g02162(.din(n2353), .dout(n2354));
  jor  g02163(.dina(n2289), .dinb(n2281), .dout(n2355));
  jand g02164(.dina(n2355), .dinb(n2354), .dout(n2356));
  jnot g02165(.din(n2356), .dout(n2357));
  jand g02166(.dina(n2296), .dinb(\a[17] ), .dout(n2358));
  jand g02167(.dina(\a[18] ), .dinb(\a[16] ), .dout(n2359));
  jand g02168(.dina(\a[33] ), .dinb(\a[1] ), .dout(n2360));
  jxor g02169(.dina(n2360), .dinb(n2359), .dout(n2361));
  jxor g02170(.dina(n2361), .dinb(n2358), .dout(n2362));
  jand g02171(.dina(n2285), .dinb(n2283), .dout(n2363));
  jnot g02172(.din(n2363), .dout(n2364));
  jand g02173(.dina(n2364), .dinb(n2287), .dout(n2365));
  jxor g02174(.dina(n2365), .dinb(n2362), .dout(n2366));
  jxor g02175(.dina(n2366), .dinb(n2357), .dout(n2367));
  jxor g02176(.dina(n2367), .dinb(n2352), .dout(n2368));
  jor  g02177(.dina(n2311), .dinb(n2302), .dout(n2369));
  jand g02178(.dina(n2312), .dinb(n2295), .dout(n2370));
  jnot g02179(.din(n2370), .dout(n2371));
  jand g02180(.dina(n2371), .dinb(n2369), .dout(n2372));
  jnot g02181(.din(n2372), .dout(n2373));
  jand g02182(.dina(n2299), .dinb(n2298), .dout(n2374));
  jand g02183(.dina(n2300), .dinb(n2297), .dout(n2375));
  jor  g02184(.dina(n2375), .dinb(n2374), .dout(n2376));
  jand g02185(.dina(n2306), .dinb(n2304), .dout(n2377));
  jnot g02186(.din(n2377), .dout(n2378));
  jand g02187(.dina(n2378), .dinb(n2309), .dout(n2379));
  jxor g02188(.dina(n2379), .dinb(n2376), .dout(n2380));
  jnot g02189(.din(n2380), .dout(n2381));
  jnot g02190(.din(n2142), .dout(n2382));
  jand g02191(.dina(n1658), .dinb(n555), .dout(n2383));
  jnot g02192(.din(n2383), .dout(n2384));
  jand g02193(.dina(\a[23] ), .dinb(\a[11] ), .dout(n2385));
  jand g02194(.dina(\a[22] ), .dinb(\a[12] ), .dout(n2386));
  jor  g02195(.dina(n2386), .dinb(n2385), .dout(n2387));
  jand g02196(.dina(n2387), .dinb(n2384), .dout(n2388));
  jxor g02197(.dina(n2388), .dinb(n2382), .dout(n2389));
  jxor g02198(.dina(n2389), .dinb(n2381), .dout(n2390));
  jxor g02199(.dina(n2390), .dinb(n2373), .dout(n2391));
  jand g02200(.dina(\a[24] ), .dinb(\a[10] ), .dout(n2392));
  jand g02201(.dina(\a[29] ), .dinb(\a[5] ), .dout(n2393));
  jand g02202(.dina(\a[25] ), .dinb(\a[9] ), .dout(n2394));
  jxor g02203(.dina(n2394), .dinb(n2393), .dout(n2395));
  jxor g02204(.dina(n2395), .dinb(n2392), .dout(n2396));
  jnot g02205(.din(n2396), .dout(n2397));
  jand g02206(.dina(\a[21] ), .dinb(\a[13] ), .dout(n2398));
  jnot g02207(.din(n2398), .dout(n2399));
  jand g02208(.dina(n1287), .dinb(n976), .dout(n2400));
  jnot g02209(.din(n2400), .dout(n2401));
  jand g02210(.dina(\a[20] ), .dinb(\a[14] ), .dout(n2402));
  jand g02211(.dina(\a[19] ), .dinb(\a[15] ), .dout(n2403));
  jor  g02212(.dina(n2403), .dinb(n2402), .dout(n2404));
  jand g02213(.dina(n2404), .dinb(n2401), .dout(n2405));
  jxor g02214(.dina(n2405), .dinb(n2399), .dout(n2406));
  jxor g02215(.dina(n2406), .dinb(n2397), .dout(n2407));
  jnot g02216(.din(n2407), .dout(n2408));
  jand g02217(.dina(\a[28] ), .dinb(\a[6] ), .dout(n2409));
  jnot g02218(.din(n2409), .dout(n2410));
  jand g02219(.dina(n1927), .dinb(n499), .dout(n2411));
  jnot g02220(.din(n2411), .dout(n2412));
  jand g02221(.dina(\a[27] ), .dinb(\a[7] ), .dout(n2413));
  jand g02222(.dina(\a[26] ), .dinb(\a[8] ), .dout(n2414));
  jor  g02223(.dina(n2414), .dinb(n2413), .dout(n2415));
  jand g02224(.dina(n2415), .dinb(n2412), .dout(n2416));
  jxor g02225(.dina(n2416), .dinb(n2410), .dout(n2417));
  jxor g02226(.dina(n2417), .dinb(n2408), .dout(n2418));
  jxor g02227(.dina(n2418), .dinb(n2391), .dout(n2419));
  jxor g02228(.dina(n2419), .dinb(n2368), .dout(n2420));
  jxor g02229(.dina(n2420), .dinb(n2344), .dout(n2421));
  jand g02230(.dina(n2229), .dinb(n2226), .dout(n2422));
  jand g02231(.dina(n2291), .dinb(n2230), .dout(n2423));
  jor  g02232(.dina(n2423), .dinb(n2422), .dout(n2424));
  jand g02233(.dina(n2256), .dinb(n2239), .dout(n2425));
  jand g02234(.dina(n2290), .dinb(n2257), .dout(n2426));
  jor  g02235(.dina(n2426), .dinb(n2425), .dout(n2427));
  jand g02236(.dina(n2221), .dinb(n2218), .dout(n2428));
  jand g02237(.dina(n2225), .dinb(n2222), .dout(n2429));
  jor  g02238(.dina(n2429), .dinb(n2428), .dout(n2430));
  jxor g02239(.dina(n2430), .dinb(n2427), .dout(n2431));
  jand g02240(.dina(n2243), .dinb(n2241), .dout(n2432));
  jnot g02241(.din(n2432), .dout(n2433));
  jor  g02242(.dina(n2255), .dinb(n2245), .dout(n2434));
  jand g02243(.dina(n2434), .dinb(n2433), .dout(n2435));
  jnot g02244(.din(n2435), .dout(n2436));
  jand g02245(.dina(n2237), .dinb(n2235), .dout(n2437));
  jand g02246(.dina(n2238), .dinb(n2233), .dout(n2438));
  jor  g02247(.dina(n2438), .dinb(n2437), .dout(n2439));
  jand g02248(.dina(\a[31] ), .dinb(\a[30] ), .dout(n2440));
  jand g02249(.dina(n2440), .dinb(n265), .dout(n2441));
  jnot g02250(.din(n2441), .dout(n2442));
  jand g02251(.dina(n201), .dinb(\a[31] ), .dout(n2443));
  jand g02252(.dina(n2443), .dinb(\a[34] ), .dout(n2444));
  jand g02253(.dina(\a[30] ), .dinb(\a[4] ), .dout(n2445));
  jand g02254(.dina(\a[34] ), .dinb(\a[0] ), .dout(n2446));
  jand g02255(.dina(n2446), .dinb(n2445), .dout(n2447));
  jor  g02256(.dina(n2447), .dinb(n2444), .dout(n2448));
  jand g02257(.dina(n2448), .dinb(n2442), .dout(n2449));
  jnot g02258(.din(n2449), .dout(n2450));
  jand g02259(.dina(\a[31] ), .dinb(\a[3] ), .dout(n2451));
  jor  g02260(.dina(n2451), .dinb(n2445), .dout(n2452));
  jand g02261(.dina(n2452), .dinb(n2442), .dout(n2453));
  jor  g02262(.dina(n2453), .dinb(n2446), .dout(n2454));
  jand g02263(.dina(n2454), .dinb(n2450), .dout(n2455));
  jxor g02264(.dina(n2455), .dinb(n2439), .dout(n2456));
  jxor g02265(.dina(n2456), .dinb(n2436), .dout(n2457));
  jxor g02266(.dina(n2457), .dinb(n2431), .dout(n2458));
  jxor g02267(.dina(n2458), .dinb(n2424), .dout(n2459));
  jxor g02268(.dina(n2459), .dinb(n2421), .dout(n2460));
  jand g02269(.dina(n2460), .dinb(n2339), .dout(n2461));
  jor  g02270(.dina(n2460), .dinb(n2339), .dout(n2462));
  jnot g02271(.din(n2462), .dout(n2463));
  jor  g02272(.dina(n2463), .dinb(n2461), .dout(n2464));
  jand g02273(.dina(n2331), .dinb(n2327), .dout(n2465));
  jnot g02274(.din(n2465), .dout(n2466));
  jnot g02275(.din(n2331), .dout(n2467));
  jand g02276(.dina(n2467), .dinb(n2328), .dout(n2468));
  jor  g02277(.dina(n2335), .dinb(n2468), .dout(n2469));
  jand g02278(.dina(n2469), .dinb(n2466), .dout(n2470));
  jxor g02279(.dina(n2470), .dinb(n2464), .dout(\asquared[35] ));
  jand g02280(.dina(n2458), .dinb(n2424), .dout(n2472));
  jand g02281(.dina(n2459), .dinb(n2421), .dout(n2473));
  jor  g02282(.dina(n2473), .dinb(n2472), .dout(n2474));
  jand g02283(.dina(n2419), .dinb(n2368), .dout(n2475));
  jand g02284(.dina(n2420), .dinb(n2344), .dout(n2476));
  jor  g02285(.dina(n2476), .dinb(n2475), .dout(n2477));
  jand g02286(.dina(n2350), .dinb(n2347), .dout(n2478));
  jand g02287(.dina(n2351), .dinb(n2271), .dout(n2479));
  jor  g02288(.dina(n2479), .dinb(n2478), .dout(n2480));
  jand g02289(.dina(n2361), .dinb(n2358), .dout(n2481));
  jand g02290(.dina(n2365), .dinb(n2362), .dout(n2482));
  jor  g02291(.dina(n2482), .dinb(n2481), .dout(n2483));
  jxor g02292(.dina(n2483), .dinb(n2480), .dout(n2484));
  jnot g02293(.din(n2484), .dout(n2485));
  jand g02294(.dina(n2379), .dinb(n2376), .dout(n2486));
  jnot g02295(.din(n2486), .dout(n2487));
  jor  g02296(.dina(n2389), .dinb(n2381), .dout(n2488));
  jand g02297(.dina(n2488), .dinb(n2487), .dout(n2489));
  jxor g02298(.dina(n2489), .dinb(n2485), .dout(n2490));
  jand g02299(.dina(n2366), .dinb(n2357), .dout(n2491));
  jand g02300(.dina(n2367), .dinb(n2352), .dout(n2492));
  jor  g02301(.dina(n2492), .dinb(n2491), .dout(n2493));
  jxor g02302(.dina(n2493), .dinb(n2490), .dout(n2494));
  jand g02303(.dina(n2390), .dinb(n2373), .dout(n2495));
  jand g02304(.dina(n2418), .dinb(n2391), .dout(n2496));
  jor  g02305(.dina(n2496), .dinb(n2495), .dout(n2497));
  jxor g02306(.dina(n2497), .dinb(n2494), .dout(n2498));
  jxor g02307(.dina(n2498), .dinb(n2477), .dout(n2499));
  jand g02308(.dina(n2430), .dinb(n2427), .dout(n2500));
  jand g02309(.dina(n2457), .dinb(n2431), .dout(n2501));
  jor  g02310(.dina(n2501), .dinb(n2500), .dout(n2502));
  jand g02311(.dina(n2384), .dinb(n2382), .dout(n2503));
  jnot g02312(.din(n2503), .dout(n2504));
  jand g02313(.dina(n2504), .dinb(n2387), .dout(n2505));
  jand g02314(.dina(n2401), .dinb(n2399), .dout(n2506));
  jnot g02315(.din(n2506), .dout(n2507));
  jand g02316(.dina(n2507), .dinb(n2404), .dout(n2508));
  jxor g02317(.dina(n2508), .dinb(n2505), .dout(n2509));
  jor  g02318(.dina(n2448), .dinb(n2441), .dout(n2510));
  jxor g02319(.dina(n2510), .dinb(n2509), .dout(n2511));
  jor  g02320(.dina(n2406), .dinb(n2397), .dout(n2512));
  jor  g02321(.dina(n2417), .dinb(n2408), .dout(n2513));
  jand g02322(.dina(n2513), .dinb(n2512), .dout(n2514));
  jnot g02323(.din(n2514), .dout(n2515));
  jand g02324(.dina(n2394), .dinb(n2393), .dout(n2516));
  jand g02325(.dina(n2395), .dinb(n2392), .dout(n2517));
  jor  g02326(.dina(n2517), .dinb(n2516), .dout(n2518));
  jand g02327(.dina(n857), .dinb(\a[34] ), .dout(n2519));
  jnot g02328(.din(n2519), .dout(n2520));
  jand g02329(.dina(\a[34] ), .dinb(\a[1] ), .dout(n2521));
  jor  g02330(.dina(n2521), .dinb(\a[18] ), .dout(n2522));
  jand g02331(.dina(n2522), .dinb(n2520), .dout(n2523));
  jand g02332(.dina(n2412), .dinb(n2410), .dout(n2524));
  jnot g02333(.din(n2524), .dout(n2525));
  jand g02334(.dina(n2525), .dinb(n2415), .dout(n2526));
  jxor g02335(.dina(n2526), .dinb(n2523), .dout(n2527));
  jxor g02336(.dina(n2527), .dinb(n2518), .dout(n2528));
  jxor g02337(.dina(n2528), .dinb(n2515), .dout(n2529));
  jxor g02338(.dina(n2529), .dinb(n2511), .dout(n2530));
  jxor g02339(.dina(n2530), .dinb(n2502), .dout(n2531));
  jand g02340(.dina(n2455), .dinb(n2439), .dout(n2532));
  jand g02341(.dina(n2456), .dinb(n2436), .dout(n2533));
  jor  g02342(.dina(n2533), .dinb(n2532), .dout(n2534));
  jand g02343(.dina(\a[30] ), .dinb(\a[5] ), .dout(n2535));
  jand g02344(.dina(\a[29] ), .dinb(\a[27] ), .dout(n2536));
  jand g02345(.dina(n2536), .dinb(n544), .dout(n2537));
  jnot g02346(.din(n2537), .dout(n2538));
  jand g02347(.dina(\a[27] ), .dinb(\a[8] ), .dout(n2539));
  jand g02348(.dina(\a[29] ), .dinb(\a[6] ), .dout(n2540));
  jor  g02349(.dina(n2540), .dinb(n2539), .dout(n2541));
  jand g02350(.dina(n2541), .dinb(n2538), .dout(n2542));
  jxor g02351(.dina(n2542), .dinb(n2535), .dout(n2543));
  jand g02352(.dina(\a[28] ), .dinb(\a[7] ), .dout(n2544));
  jand g02353(.dina(\a[19] ), .dinb(\a[16] ), .dout(n2545));
  jxor g02354(.dina(n2545), .dinb(n1107), .dout(n2546));
  jxor g02355(.dina(n2546), .dinb(n2544), .dout(n2547));
  jxor g02356(.dina(n2547), .dinb(n2543), .dout(n2548));
  jnot g02357(.din(n2548), .dout(n2549));
  jand g02358(.dina(\a[31] ), .dinb(\a[4] ), .dout(n2550));
  jnot g02359(.din(n2550), .dout(n2551));
  jand g02360(.dina(n2128), .dinb(n453), .dout(n2552));
  jnot g02361(.din(n2552), .dout(n2553));
  jand g02362(.dina(\a[26] ), .dinb(\a[9] ), .dout(n2554));
  jand g02363(.dina(\a[25] ), .dinb(\a[10] ), .dout(n2555));
  jor  g02364(.dina(n2555), .dinb(n2554), .dout(n2556));
  jand g02365(.dina(n2556), .dinb(n2553), .dout(n2557));
  jxor g02366(.dina(n2557), .dinb(n2551), .dout(n2558));
  jxor g02367(.dina(n2558), .dinb(n2549), .dout(n2559));
  jxor g02368(.dina(n2559), .dinb(n2534), .dout(n2560));
  jand g02369(.dina(n2360), .dinb(n2359), .dout(n2561));
  jand g02370(.dina(\a[35] ), .dinb(\a[0] ), .dout(n2562));
  jand g02371(.dina(\a[33] ), .dinb(\a[2] ), .dout(n2563));
  jor  g02372(.dina(n2563), .dinb(n2562), .dout(n2564));
  jand g02373(.dina(\a[35] ), .dinb(\a[2] ), .dout(n2565));
  jand g02374(.dina(n2565), .dinb(n2251), .dout(n2566));
  jnot g02375(.din(n2566), .dout(n2567));
  jand g02376(.dina(n2567), .dinb(n2564), .dout(n2568));
  jxor g02377(.dina(n2568), .dinb(n2561), .dout(n2569));
  jnot g02378(.din(n2569), .dout(n2570));
  jand g02379(.dina(\a[32] ), .dinb(\a[3] ), .dout(n2571));
  jnot g02380(.din(n2571), .dout(n2572));
  jand g02381(.dina(n1942), .dinb(n555), .dout(n2573));
  jnot g02382(.din(n2573), .dout(n2574));
  jand g02383(.dina(\a[24] ), .dinb(\a[11] ), .dout(n2575));
  jand g02384(.dina(\a[23] ), .dinb(\a[12] ), .dout(n2576));
  jor  g02385(.dina(n2576), .dinb(n2575), .dout(n2577));
  jand g02386(.dina(n2577), .dinb(n2574), .dout(n2578));
  jxor g02387(.dina(n2578), .dinb(n2572), .dout(n2579));
  jxor g02388(.dina(n2579), .dinb(n2570), .dout(n2580));
  jnot g02389(.din(n2580), .dout(n2581));
  jand g02390(.dina(\a[22] ), .dinb(\a[13] ), .dout(n2582));
  jnot g02391(.din(n2582), .dout(n2583));
  jand g02392(.dina(n1490), .dinb(n976), .dout(n2584));
  jnot g02393(.din(n2584), .dout(n2585));
  jand g02394(.dina(\a[21] ), .dinb(\a[14] ), .dout(n2586));
  jand g02395(.dina(\a[20] ), .dinb(\a[15] ), .dout(n2587));
  jor  g02396(.dina(n2587), .dinb(n2586), .dout(n2588));
  jand g02397(.dina(n2588), .dinb(n2585), .dout(n2589));
  jxor g02398(.dina(n2589), .dinb(n2583), .dout(n2590));
  jxor g02399(.dina(n2590), .dinb(n2581), .dout(n2591));
  jxor g02400(.dina(n2591), .dinb(n2560), .dout(n2592));
  jxor g02401(.dina(n2592), .dinb(n2531), .dout(n2593));
  jxor g02402(.dina(n2593), .dinb(n2499), .dout(n2594));
  jnot g02403(.din(n2594), .dout(n2595));
  jxor g02404(.dina(n2595), .dinb(n2474), .dout(n2596));
  jnot g02405(.din(n2461), .dout(n2597));
  jor  g02406(.dina(n2470), .dinb(n2463), .dout(n2598));
  jand g02407(.dina(n2598), .dinb(n2597), .dout(n2599));
  jxor g02408(.dina(n2599), .dinb(n2596), .dout(\asquared[36] ));
  jand g02409(.dina(n2498), .dinb(n2477), .dout(n2601));
  jand g02410(.dina(n2593), .dinb(n2499), .dout(n2602));
  jor  g02411(.dina(n2602), .dinb(n2601), .dout(n2603));
  jand g02412(.dina(n2530), .dinb(n2502), .dout(n2604));
  jand g02413(.dina(n2592), .dinb(n2531), .dout(n2605));
  jor  g02414(.dina(n2605), .dinb(n2604), .dout(n2606));
  jand g02415(.dina(n2508), .dinb(n2505), .dout(n2607));
  jand g02416(.dina(n2510), .dinb(n2509), .dout(n2608));
  jor  g02417(.dina(n2608), .dinb(n2607), .dout(n2609));
  jand g02418(.dina(n2526), .dinb(n2523), .dout(n2610));
  jand g02419(.dina(n2527), .dinb(n2518), .dout(n2611));
  jor  g02420(.dina(n2611), .dinb(n2610), .dout(n2612));
  jxor g02421(.dina(n2612), .dinb(n2609), .dout(n2613));
  jnot g02422(.din(n2613), .dout(n2614));
  jor  g02423(.dina(n2579), .dinb(n2570), .dout(n2615));
  jor  g02424(.dina(n2590), .dinb(n2581), .dout(n2616));
  jand g02425(.dina(n2616), .dinb(n2615), .dout(n2617));
  jxor g02426(.dina(n2617), .dinb(n2614), .dout(n2618));
  jand g02427(.dina(n2528), .dinb(n2515), .dout(n2619));
  jand g02428(.dina(n2529), .dinb(n2511), .dout(n2620));
  jor  g02429(.dina(n2620), .dinb(n2619), .dout(n2621));
  jxor g02430(.dina(n2621), .dinb(n2618), .dout(n2622));
  jand g02431(.dina(n2559), .dinb(n2534), .dout(n2623));
  jand g02432(.dina(n2591), .dinb(n2560), .dout(n2624));
  jor  g02433(.dina(n2624), .dinb(n2623), .dout(n2625));
  jxor g02434(.dina(n2625), .dinb(n2622), .dout(n2626));
  jxor g02435(.dina(n2626), .dinb(n2606), .dout(n2627));
  jand g02436(.dina(\a[34] ), .dinb(\a[2] ), .dout(n2628));
  jand g02437(.dina(\a[23] ), .dinb(\a[13] ), .dout(n2629));
  jand g02438(.dina(\a[24] ), .dinb(\a[12] ), .dout(n2630));
  jor  g02439(.dina(n2630), .dinb(n2629), .dout(n2631));
  jand g02440(.dina(n1942), .dinb(n899), .dout(n2632));
  jnot g02441(.din(n2632), .dout(n2633));
  jand g02442(.dina(n2633), .dinb(n2631), .dout(n2634));
  jxor g02443(.dina(n2634), .dinb(n2628), .dout(n2635));
  jand g02444(.dina(\a[27] ), .dinb(\a[9] ), .dout(n2636));
  jand g02445(.dina(\a[31] ), .dinb(\a[5] ), .dout(n2637));
  jand g02446(.dina(n2637), .dinb(n2636), .dout(n2638));
  jnot g02447(.din(n2638), .dout(n2639));
  jand g02448(.dina(n1927), .dinb(n453), .dout(n2640));
  jand g02449(.dina(\a[26] ), .dinb(\a[10] ), .dout(n2641));
  jand g02450(.dina(n2641), .dinb(n2637), .dout(n2642));
  jor  g02451(.dina(n2642), .dinb(n2640), .dout(n2643));
  jand g02452(.dina(n2643), .dinb(n2639), .dout(n2644));
  jnot g02453(.din(n2644), .dout(n2645));
  jxor g02454(.dina(n2637), .dinb(n2636), .dout(n2646));
  jor  g02455(.dina(n2646), .dinb(n2641), .dout(n2647));
  jand g02456(.dina(n2647), .dinb(n2645), .dout(n2648));
  jxor g02457(.dina(n2648), .dinb(n2635), .dout(n2649));
  jnot g02458(.din(n2649), .dout(n2650));
  jand g02459(.dina(\a[30] ), .dinb(\a[6] ), .dout(n2651));
  jnot g02460(.din(n2651), .dout(n2652));
  jand g02461(.dina(\a[29] ), .dinb(\a[28] ), .dout(n2653));
  jand g02462(.dina(n2653), .dinb(n499), .dout(n2654));
  jnot g02463(.din(n2654), .dout(n2655));
  jand g02464(.dina(\a[29] ), .dinb(\a[7] ), .dout(n2656));
  jand g02465(.dina(\a[28] ), .dinb(\a[8] ), .dout(n2657));
  jor  g02466(.dina(n2657), .dinb(n2656), .dout(n2658));
  jand g02467(.dina(n2658), .dinb(n2655), .dout(n2659));
  jxor g02468(.dina(n2659), .dinb(n2652), .dout(n2660));
  jxor g02469(.dina(n2660), .dinb(n2650), .dout(n2661));
  jand g02470(.dina(n2483), .dinb(n2480), .dout(n2662));
  jnot g02471(.din(n2662), .dout(n2663));
  jor  g02472(.dina(n2489), .dinb(n2485), .dout(n2664));
  jand g02473(.dina(n2664), .dinb(n2663), .dout(n2665));
  jnot g02474(.din(n2665), .dout(n2666));
  jand g02475(.dina(\a[32] ), .dinb(\a[4] ), .dout(n2667));
  jand g02476(.dina(\a[25] ), .dinb(\a[11] ), .dout(n2668));
  jand g02477(.dina(n2668), .dinb(n2667), .dout(n2669));
  jnot g02478(.din(n2669), .dout(n2670));
  jand g02479(.dina(\a[33] ), .dinb(\a[32] ), .dout(n2671));
  jand g02480(.dina(n2671), .dinb(n265), .dout(n2672));
  jand g02481(.dina(\a[33] ), .dinb(\a[3] ), .dout(n2673));
  jand g02482(.dina(n2673), .dinb(n2668), .dout(n2674));
  jor  g02483(.dina(n2674), .dinb(n2672), .dout(n2675));
  jnot g02484(.din(n2675), .dout(n2676));
  jand g02485(.dina(n2676), .dinb(n2670), .dout(n2677));
  jor  g02486(.dina(n2668), .dinb(n2667), .dout(n2678));
  jand g02487(.dina(n2678), .dinb(n2677), .dout(n2679));
  jand g02488(.dina(n2675), .dinb(n2670), .dout(n2680));
  jnot g02489(.din(n2680), .dout(n2681));
  jand g02490(.dina(n2681), .dinb(n2673), .dout(n2682));
  jor  g02491(.dina(n2682), .dinb(n2679), .dout(n2683));
  jand g02492(.dina(\a[22] ), .dinb(\a[14] ), .dout(n2684));
  jnot g02493(.din(n2684), .dout(n2685));
  jand g02494(.dina(n1490), .dinb(n829), .dout(n2686));
  jnot g02495(.din(n2686), .dout(n2687));
  jand g02496(.dina(\a[20] ), .dinb(\a[16] ), .dout(n2688));
  jand g02497(.dina(\a[21] ), .dinb(\a[15] ), .dout(n2689));
  jor  g02498(.dina(n2689), .dinb(n2688), .dout(n2690));
  jand g02499(.dina(n2690), .dinb(n2687), .dout(n2691));
  jxor g02500(.dina(n2691), .dinb(n2685), .dout(n2692));
  jnot g02501(.din(n2692), .dout(n2693));
  jxor g02502(.dina(n2693), .dinb(n2683), .dout(n2694));
  jand g02503(.dina(\a[36] ), .dinb(\a[0] ), .dout(n2695));
  jxor g02504(.dina(n2695), .dinb(n2519), .dout(n2696));
  jand g02505(.dina(\a[19] ), .dinb(\a[17] ), .dout(n2697));
  jand g02506(.dina(\a[35] ), .dinb(\a[1] ), .dout(n2698));
  jxor g02507(.dina(n2698), .dinb(n2697), .dout(n2699));
  jxor g02508(.dina(n2699), .dinb(n2696), .dout(n2700));
  jxor g02509(.dina(n2700), .dinb(n2694), .dout(n2701));
  jxor g02510(.dina(n2701), .dinb(n2666), .dout(n2702));
  jxor g02511(.dina(n2702), .dinb(n2661), .dout(n2703));
  jand g02512(.dina(n2493), .dinb(n2490), .dout(n2704));
  jand g02513(.dina(n2497), .dinb(n2494), .dout(n2705));
  jor  g02514(.dina(n2705), .dinb(n2704), .dout(n2706));
  jand g02515(.dina(n2545), .dinb(n1107), .dout(n2707));
  jand g02516(.dina(n2546), .dinb(n2544), .dout(n2708));
  jor  g02517(.dina(n2708), .dinb(n2707), .dout(n2709));
  jand g02518(.dina(n2542), .dinb(n2535), .dout(n2710));
  jor  g02519(.dina(n2710), .dinb(n2537), .dout(n2711));
  jand g02520(.dina(n2553), .dinb(n2551), .dout(n2712));
  jnot g02521(.din(n2712), .dout(n2713));
  jand g02522(.dina(n2713), .dinb(n2556), .dout(n2714));
  jxor g02523(.dina(n2714), .dinb(n2711), .dout(n2715));
  jxor g02524(.dina(n2715), .dinb(n2709), .dout(n2716));
  jand g02525(.dina(n2568), .dinb(n2561), .dout(n2717));
  jor  g02526(.dina(n2717), .dinb(n2566), .dout(n2718));
  jand g02527(.dina(n2585), .dinb(n2583), .dout(n2719));
  jnot g02528(.din(n2719), .dout(n2720));
  jand g02529(.dina(n2720), .dinb(n2588), .dout(n2721));
  jand g02530(.dina(n2574), .dinb(n2572), .dout(n2722));
  jnot g02531(.din(n2722), .dout(n2723));
  jand g02532(.dina(n2723), .dinb(n2577), .dout(n2724));
  jxor g02533(.dina(n2724), .dinb(n2721), .dout(n2725));
  jxor g02534(.dina(n2725), .dinb(n2718), .dout(n2726));
  jnot g02535(.din(n2726), .dout(n2727));
  jand g02536(.dina(n2547), .dinb(n2543), .dout(n2728));
  jnot g02537(.din(n2728), .dout(n2729));
  jor  g02538(.dina(n2558), .dinb(n2549), .dout(n2730));
  jand g02539(.dina(n2730), .dinb(n2729), .dout(n2731));
  jxor g02540(.dina(n2731), .dinb(n2727), .dout(n2732));
  jxor g02541(.dina(n2732), .dinb(n2716), .dout(n2733));
  jxor g02542(.dina(n2733), .dinb(n2706), .dout(n2734));
  jxor g02543(.dina(n2734), .dinb(n2703), .dout(n2735));
  jxor g02544(.dina(n2735), .dinb(n2627), .dout(n2736));
  jnot g02545(.din(n2736), .dout(n2737));
  jxor g02546(.dina(n2737), .dinb(n2603), .dout(n2738));
  jand g02547(.dina(n2594), .dinb(n2474), .dout(n2739));
  jnot g02548(.din(n2739), .dout(n2740));
  jnot g02549(.din(n2474), .dout(n2741));
  jand g02550(.dina(n2595), .dinb(n2741), .dout(n2742));
  jor  g02551(.dina(n2599), .dinb(n2742), .dout(n2743));
  jand g02552(.dina(n2743), .dinb(n2740), .dout(n2744));
  jxor g02553(.dina(n2744), .dinb(n2738), .dout(\asquared[37] ));
  jand g02554(.dina(n2626), .dinb(n2606), .dout(n2746));
  jand g02555(.dina(n2735), .dinb(n2627), .dout(n2747));
  jor  g02556(.dina(n2747), .dinb(n2746), .dout(n2748));
  jand g02557(.dina(n2621), .dinb(n2618), .dout(n2749));
  jand g02558(.dina(n2625), .dinb(n2622), .dout(n2750));
  jor  g02559(.dina(n2750), .dinb(n2749), .dout(n2751));
  jand g02560(.dina(n2634), .dinb(n2628), .dout(n2752));
  jor  g02561(.dina(n2752), .dinb(n2632), .dout(n2753));
  jnot g02562(.din(n2677), .dout(n2754));
  jand g02563(.dina(n2687), .dinb(n2685), .dout(n2755));
  jnot g02564(.din(n2755), .dout(n2756));
  jand g02565(.dina(n2756), .dinb(n2690), .dout(n2757));
  jxor g02566(.dina(n2757), .dinb(n2754), .dout(n2758));
  jxor g02567(.dina(n2758), .dinb(n2753), .dout(n2759));
  jand g02568(.dina(n2693), .dinb(n2683), .dout(n2760));
  jand g02569(.dina(n2700), .dinb(n2694), .dout(n2761));
  jor  g02570(.dina(n2761), .dinb(n2760), .dout(n2762));
  jxor g02571(.dina(n2762), .dinb(n2759), .dout(n2763));
  jor  g02572(.dina(n2643), .dinb(n2638), .dout(n2764));
  jand g02573(.dina(n2695), .dinb(n2519), .dout(n2765));
  jand g02574(.dina(n2699), .dinb(n2696), .dout(n2766));
  jor  g02575(.dina(n2766), .dinb(n2765), .dout(n2767));
  jxor g02576(.dina(n2767), .dinb(n2764), .dout(n2768));
  jnot g02577(.din(n2768), .dout(n2769));
  jand g02578(.dina(\a[24] ), .dinb(\a[13] ), .dout(n2770));
  jnot g02579(.din(n2770), .dout(n2771));
  jand g02580(.dina(n1658), .dinb(n976), .dout(n2772));
  jnot g02581(.din(n2772), .dout(n2773));
  jand g02582(.dina(\a[23] ), .dinb(\a[14] ), .dout(n2774));
  jand g02583(.dina(\a[22] ), .dinb(\a[15] ), .dout(n2775));
  jor  g02584(.dina(n2775), .dinb(n2774), .dout(n2776));
  jand g02585(.dina(n2776), .dinb(n2773), .dout(n2777));
  jxor g02586(.dina(n2777), .dinb(n2771), .dout(n2778));
  jxor g02587(.dina(n2778), .dinb(n2769), .dout(n2779));
  jxor g02588(.dina(n2779), .dinb(n2763), .dout(n2780));
  jxor g02589(.dina(n2780), .dinb(n2751), .dout(n2781));
  jand g02590(.dina(n2724), .dinb(n2721), .dout(n2782));
  jand g02591(.dina(n2725), .dinb(n2718), .dout(n2783));
  jor  g02592(.dina(n2783), .dinb(n2782), .dout(n2784));
  jand g02593(.dina(\a[26] ), .dinb(\a[11] ), .dout(n2785));
  jand g02594(.dina(\a[32] ), .dinb(\a[5] ), .dout(n2786));
  jand g02595(.dina(\a[27] ), .dinb(\a[10] ), .dout(n2787));
  jxor g02596(.dina(n2787), .dinb(n2786), .dout(n2788));
  jxor g02597(.dina(n2788), .dinb(n2785), .dout(n2789));
  jnot g02598(.din(n2789), .dout(n2790));
  jand g02599(.dina(\a[29] ), .dinb(\a[8] ), .dout(n2791));
  jnot g02600(.din(n2791), .dout(n2792));
  jand g02601(.dina(n1287), .dinb(n1107), .dout(n2793));
  jnot g02602(.din(n2793), .dout(n2794));
  jand g02603(.dina(\a[20] ), .dinb(\a[17] ), .dout(n2795));
  jor  g02604(.dina(n2795), .dinb(n1024), .dout(n2796));
  jand g02605(.dina(n2796), .dinb(n2794), .dout(n2797));
  jxor g02606(.dina(n2797), .dinb(n2792), .dout(n2798));
  jxor g02607(.dina(n2798), .dinb(n2790), .dout(n2799));
  jxor g02608(.dina(n2799), .dinb(n2784), .dout(n2800));
  jnot g02609(.din(n2800), .dout(n2801));
  jand g02610(.dina(n2612), .dinb(n2609), .dout(n2802));
  jnot g02611(.din(n2802), .dout(n2803));
  jor  g02612(.dina(n2617), .dinb(n2614), .dout(n2804));
  jand g02613(.dina(n2804), .dinb(n2803), .dout(n2805));
  jxor g02614(.dina(n2805), .dinb(n2801), .dout(n2806));
  jand g02615(.dina(\a[28] ), .dinb(\a[9] ), .dout(n2807));
  jand g02616(.dina(n2440), .dinb(n410), .dout(n2808));
  jnot g02617(.din(n2808), .dout(n2809));
  jand g02618(.dina(\a[30] ), .dinb(\a[28] ), .dout(n2810));
  jand g02619(.dina(n2810), .dinb(n684), .dout(n2811));
  jand g02620(.dina(\a[31] ), .dinb(\a[6] ), .dout(n2812));
  jand g02621(.dina(n2812), .dinb(n2807), .dout(n2813));
  jor  g02622(.dina(n2813), .dinb(n2811), .dout(n2814));
  jand g02623(.dina(n2814), .dinb(n2809), .dout(n2815));
  jnot g02624(.din(n2815), .dout(n2816));
  jand g02625(.dina(n2816), .dinb(n2807), .dout(n2817));
  jor  g02626(.dina(n2814), .dinb(n2808), .dout(n2818));
  jnot g02627(.din(n2818), .dout(n2819));
  jand g02628(.dina(\a[30] ), .dinb(\a[7] ), .dout(n2820));
  jor  g02629(.dina(n2820), .dinb(n2812), .dout(n2821));
  jand g02630(.dina(n2821), .dinb(n2819), .dout(n2822));
  jor  g02631(.dina(n2822), .dinb(n2817), .dout(n2823));
  jand g02632(.dina(\a[33] ), .dinb(\a[25] ), .dout(n2824));
  jand g02633(.dina(n2824), .dinb(n674), .dout(n2825));
  jand g02634(.dina(n451), .dinb(\a[25] ), .dout(n2826));
  jand g02635(.dina(\a[33] ), .dinb(\a[4] ), .dout(n2827));
  jand g02636(.dina(n2827), .dinb(\a[0] ), .dout(n2828));
  jor  g02637(.dina(n2828), .dinb(n2826), .dout(n2829));
  jand g02638(.dina(n2829), .dinb(\a[37] ), .dout(n2830));
  jor  g02639(.dina(n2830), .dinb(n2825), .dout(n2831));
  jnot g02640(.din(n2831), .dout(n2832));
  jand g02641(.dina(\a[25] ), .dinb(\a[12] ), .dout(n2833));
  jor  g02642(.dina(n2833), .dinb(n2827), .dout(n2834));
  jand g02643(.dina(n2834), .dinb(n2832), .dout(n2835));
  jnot g02644(.din(n2835), .dout(n2836));
  jnot g02645(.din(\a[37] ), .dout(n2837));
  jnot g02646(.din(n2825), .dout(n2838));
  jand g02647(.dina(n2829), .dinb(n2838), .dout(n2839));
  jor  g02648(.dina(n2839), .dinb(n2837), .dout(n2840));
  jor  g02649(.dina(n2840), .dinb(n193), .dout(n2841));
  jand g02650(.dina(n2841), .dinb(n2836), .dout(n2842));
  jand g02651(.dina(\a[21] ), .dinb(\a[16] ), .dout(n2843));
  jnot g02652(.din(n2843), .dout(n2844));
  jand g02653(.dina(\a[35] ), .dinb(\a[34] ), .dout(n2845));
  jand g02654(.dina(n2845), .dinb(n248), .dout(n2846));
  jnot g02655(.din(n2846), .dout(n2847));
  jand g02656(.dina(\a[34] ), .dinb(\a[3] ), .dout(n2848));
  jor  g02657(.dina(n2848), .dinb(n2565), .dout(n2849));
  jand g02658(.dina(n2849), .dinb(n2847), .dout(n2850));
  jxor g02659(.dina(n2850), .dinb(n2844), .dout(n2851));
  jxor g02660(.dina(n2851), .dinb(n2842), .dout(n2852));
  jxor g02661(.dina(n2852), .dinb(n2823), .dout(n2853));
  jxor g02662(.dina(n2853), .dinb(n2806), .dout(n2854));
  jxor g02663(.dina(n2854), .dinb(n2781), .dout(n2855));
  jand g02664(.dina(n2733), .dinb(n2706), .dout(n2856));
  jand g02665(.dina(n2734), .dinb(n2703), .dout(n2857));
  jor  g02666(.dina(n2857), .dinb(n2856), .dout(n2858));
  jand g02667(.dina(n2701), .dinb(n2666), .dout(n2859));
  jand g02668(.dina(n2702), .dinb(n2661), .dout(n2860));
  jor  g02669(.dina(n2860), .dinb(n2859), .dout(n2861));
  jor  g02670(.dina(n2731), .dinb(n2727), .dout(n2862));
  jand g02671(.dina(n2732), .dinb(n2716), .dout(n2863));
  jnot g02672(.din(n2863), .dout(n2864));
  jand g02673(.dina(n2864), .dinb(n2862), .dout(n2865));
  jnot g02674(.din(n2865), .dout(n2866));
  jand g02675(.dina(n2648), .dinb(n2635), .dout(n2867));
  jnot g02676(.din(n2867), .dout(n2868));
  jor  g02677(.dina(n2660), .dinb(n2650), .dout(n2869));
  jand g02678(.dina(n2869), .dinb(n2868), .dout(n2870));
  jnot g02679(.din(n2870), .dout(n2871));
  jand g02680(.dina(n2714), .dinb(n2711), .dout(n2872));
  jand g02681(.dina(n2715), .dinb(n2709), .dout(n2873));
  jor  g02682(.dina(n2873), .dinb(n2872), .dout(n2874));
  jand g02683(.dina(\a[36] ), .dinb(\a[1] ), .dout(n2875));
  jand g02684(.dina(n2698), .dinb(n2697), .dout(n2876));
  jor  g02685(.dina(n2876), .dinb(n891), .dout(n2877));
  jxor g02686(.dina(n2877), .dinb(n2875), .dout(n2878));
  jnot g02687(.din(n2878), .dout(n2879));
  jand g02688(.dina(n2655), .dinb(n2652), .dout(n2880));
  jnot g02689(.din(n2880), .dout(n2881));
  jand g02690(.dina(n2881), .dinb(n2658), .dout(n2882));
  jxor g02691(.dina(n2882), .dinb(n2879), .dout(n2883));
  jxor g02692(.dina(n2883), .dinb(n2874), .dout(n2884));
  jxor g02693(.dina(n2884), .dinb(n2871), .dout(n2885));
  jxor g02694(.dina(n2885), .dinb(n2866), .dout(n2886));
  jxor g02695(.dina(n2886), .dinb(n2861), .dout(n2887));
  jxor g02696(.dina(n2887), .dinb(n2858), .dout(n2888));
  jxor g02697(.dina(n2888), .dinb(n2855), .dout(n2889));
  jand g02698(.dina(n2889), .dinb(n2748), .dout(n2890));
  jor  g02699(.dina(n2889), .dinb(n2748), .dout(n2891));
  jnot g02700(.din(n2891), .dout(n2892));
  jor  g02701(.dina(n2892), .dinb(n2890), .dout(n2893));
  jand g02702(.dina(n2736), .dinb(n2603), .dout(n2894));
  jnot g02703(.din(n2894), .dout(n2895));
  jnot g02704(.din(n2603), .dout(n2896));
  jand g02705(.dina(n2737), .dinb(n2896), .dout(n2897));
  jor  g02706(.dina(n2744), .dinb(n2897), .dout(n2898));
  jand g02707(.dina(n2898), .dinb(n2895), .dout(n2899));
  jxor g02708(.dina(n2899), .dinb(n2893), .dout(\asquared[38] ));
  jand g02709(.dina(n2887), .dinb(n2858), .dout(n2901));
  jand g02710(.dina(n2888), .dinb(n2855), .dout(n2902));
  jor  g02711(.dina(n2902), .dinb(n2901), .dout(n2903));
  jand g02712(.dina(n2780), .dinb(n2751), .dout(n2904));
  jand g02713(.dina(n2854), .dinb(n2781), .dout(n2905));
  jor  g02714(.dina(n2905), .dinb(n2904), .dout(n2906));
  jor  g02715(.dina(n2805), .dinb(n2801), .dout(n2907));
  jand g02716(.dina(n2853), .dinb(n2806), .dout(n2908));
  jnot g02717(.din(n2908), .dout(n2909));
  jand g02718(.dina(n2909), .dinb(n2907), .dout(n2910));
  jnot g02719(.din(n2910), .dout(n2911));
  jand g02720(.dina(n2762), .dinb(n2759), .dout(n2912));
  jand g02721(.dina(n2779), .dinb(n2763), .dout(n2913));
  jor  g02722(.dina(n2913), .dinb(n2912), .dout(n2914));
  jxor g02723(.dina(n2914), .dinb(n2911), .dout(n2915));
  jand g02724(.dina(n2847), .dinb(n2844), .dout(n2916));
  jnot g02725(.din(n2916), .dout(n2917));
  jand g02726(.dina(n2917), .dinb(n2849), .dout(n2918));
  jxor g02727(.dina(n2918), .dinb(n2831), .dout(n2919));
  jand g02728(.dina(n2773), .dinb(n2771), .dout(n2920));
  jnot g02729(.din(n2920), .dout(n2921));
  jand g02730(.dina(n2921), .dinb(n2776), .dout(n2922));
  jxor g02731(.dina(n2922), .dinb(n2919), .dout(n2923));
  jnot g02732(.din(n2923), .dout(n2924));
  jor  g02733(.dina(n2798), .dinb(n2790), .dout(n2925));
  jand g02734(.dina(n2799), .dinb(n2784), .dout(n2926));
  jnot g02735(.din(n2926), .dout(n2927));
  jand g02736(.dina(n2927), .dinb(n2925), .dout(n2928));
  jxor g02737(.dina(n2928), .dinb(n2924), .dout(n2929));
  jand g02738(.dina(\a[32] ), .dinb(\a[6] ), .dout(n2930));
  jnot g02739(.din(n2930), .dout(n2931));
  jand g02740(.dina(\a[28] ), .dinb(\a[10] ), .dout(n2932));
  jnot g02741(.din(n2932), .dout(n2933));
  jand g02742(.dina(n2933), .dinb(n2931), .dout(n2934));
  jand g02743(.dina(n2932), .dinb(n2930), .dout(n2935));
  jnot g02744(.din(n2935), .dout(n2936));
  jand g02745(.dina(n2671), .dinb(n339), .dout(n2937));
  jand g02746(.dina(\a[33] ), .dinb(\a[5] ), .dout(n2938));
  jand g02747(.dina(n2938), .dinb(n2932), .dout(n2939));
  jor  g02748(.dina(n2939), .dinb(n2937), .dout(n2940));
  jnot g02749(.din(n2940), .dout(n2941));
  jand g02750(.dina(n2941), .dinb(n2936), .dout(n2942));
  jnot g02751(.din(n2942), .dout(n2943));
  jor  g02752(.dina(n2943), .dinb(n2934), .dout(n2944));
  jand g02753(.dina(n2940), .dinb(n2936), .dout(n2945));
  jnot g02754(.din(n2945), .dout(n2946));
  jand g02755(.dina(n2946), .dinb(n2938), .dout(n2947));
  jnot g02756(.din(n2947), .dout(n2948));
  jand g02757(.dina(n2948), .dinb(n2944), .dout(n2949));
  jand g02758(.dina(n1376), .dinb(n937), .dout(n2950));
  jnot g02759(.din(n2950), .dout(n2951));
  jand g02760(.dina(n1658), .dinb(n829), .dout(n2952));
  jand g02761(.dina(\a[23] ), .dinb(\a[15] ), .dout(n2953));
  jand g02762(.dina(\a[21] ), .dinb(\a[17] ), .dout(n2954));
  jand g02763(.dina(n2954), .dinb(n2953), .dout(n2955));
  jor  g02764(.dina(n2955), .dinb(n2952), .dout(n2956));
  jand g02765(.dina(n2956), .dinb(n2951), .dout(n2957));
  jnot g02766(.din(n2957), .dout(n2958));
  jand g02767(.dina(\a[22] ), .dinb(\a[16] ), .dout(n2959));
  jor  g02768(.dina(n2959), .dinb(n2954), .dout(n2960));
  jand g02769(.dina(n2960), .dinb(n2951), .dout(n2961));
  jor  g02770(.dina(n2961), .dinb(n2953), .dout(n2962));
  jand g02771(.dina(n2962), .dinb(n2958), .dout(n2963));
  jnot g02772(.din(n2963), .dout(n2964));
  jxor g02773(.dina(n2964), .dinb(n2949), .dout(n2965));
  jnot g02774(.din(n2965), .dout(n2966));
  jand g02775(.dina(\a[29] ), .dinb(\a[9] ), .dout(n2967));
  jnot g02776(.din(n2967), .dout(n2968));
  jand g02777(.dina(n2440), .dinb(n499), .dout(n2969));
  jnot g02778(.din(n2969), .dout(n2970));
  jand g02779(.dina(\a[31] ), .dinb(\a[7] ), .dout(n2971));
  jand g02780(.dina(\a[30] ), .dinb(\a[8] ), .dout(n2972));
  jor  g02781(.dina(n2972), .dinb(n2971), .dout(n2973));
  jand g02782(.dina(n2973), .dinb(n2970), .dout(n2974));
  jxor g02783(.dina(n2974), .dinb(n2968), .dout(n2975));
  jxor g02784(.dina(n2975), .dinb(n2966), .dout(n2976));
  jxor g02785(.dina(n2976), .dinb(n2929), .dout(n2977));
  jxor g02786(.dina(n2977), .dinb(n2915), .dout(n2978));
  jxor g02787(.dina(n2978), .dinb(n2906), .dout(n2979));
  jand g02788(.dina(n2885), .dinb(n2866), .dout(n2980));
  jand g02789(.dina(n2886), .dinb(n2861), .dout(n2981));
  jor  g02790(.dina(n2981), .dinb(n2980), .dout(n2982));
  jand g02791(.dina(n2767), .dinb(n2764), .dout(n2983));
  jnot g02792(.din(n2983), .dout(n2984));
  jor  g02793(.dina(n2778), .dinb(n2769), .dout(n2985));
  jand g02794(.dina(n2985), .dinb(n2984), .dout(n2986));
  jor  g02795(.dina(n2851), .dinb(n2842), .dout(n2987));
  jand g02796(.dina(n2852), .dinb(n2823), .dout(n2988));
  jnot g02797(.din(n2988), .dout(n2989));
  jand g02798(.dina(n2989), .dinb(n2987), .dout(n2990));
  jxor g02799(.dina(n2990), .dinb(n2986), .dout(n2991));
  jand g02800(.dina(\a[37] ), .dinb(\a[1] ), .dout(n2992));
  jxor g02801(.dina(n2992), .dinb(n1181), .dout(n2993));
  jand g02802(.dina(n2794), .dinb(n2792), .dout(n2994));
  jnot g02803(.din(n2994), .dout(n2995));
  jand g02804(.dina(n2995), .dinb(n2796), .dout(n2996));
  jxor g02805(.dina(n2996), .dinb(n2993), .dout(n2997));
  jxor g02806(.dina(n2997), .dinb(n2818), .dout(n2998));
  jxor g02807(.dina(n2998), .dinb(n2991), .dout(n2999));
  jxor g02808(.dina(n2999), .dinb(n2982), .dout(n3000));
  jand g02809(.dina(n2757), .dinb(n2754), .dout(n3001));
  jand g02810(.dina(n2758), .dinb(n2753), .dout(n3002));
  jor  g02811(.dina(n3002), .dinb(n3001), .dout(n3003));
  jand g02812(.dina(n2882), .dinb(n2879), .dout(n3004));
  jnot g02813(.din(\a[36] ), .dout(n3005));
  jand g02814(.dina(n2876), .dinb(n3005), .dout(n3006));
  jor  g02815(.dina(n3006), .dinb(n3004), .dout(n3007));
  jand g02816(.dina(\a[26] ), .dinb(\a[12] ), .dout(n3008));
  jand g02817(.dina(\a[34] ), .dinb(\a[27] ), .dout(n3009));
  jand g02818(.dina(n3009), .dinb(n602), .dout(n3010));
  jnot g02819(.din(n3010), .dout(n3011));
  jand g02820(.dina(n1927), .dinb(n555), .dout(n3012));
  jand g02821(.dina(\a[34] ), .dinb(\a[4] ), .dout(n3013));
  jand g02822(.dina(n3013), .dinb(n3008), .dout(n3014));
  jor  g02823(.dina(n3014), .dinb(n3012), .dout(n3015));
  jand g02824(.dina(n3015), .dinb(n3011), .dout(n3016));
  jnot g02825(.din(n3016), .dout(n3017));
  jand g02826(.dina(n3017), .dinb(n3008), .dout(n3018));
  jor  g02827(.dina(n3015), .dinb(n3010), .dout(n3019));
  jnot g02828(.din(n3019), .dout(n3020));
  jand g02829(.dina(\a[27] ), .dinb(\a[11] ), .dout(n3021));
  jor  g02830(.dina(n3021), .dinb(n3013), .dout(n3022));
  jand g02831(.dina(n3022), .dinb(n3020), .dout(n3023));
  jor  g02832(.dina(n3023), .dinb(n3018), .dout(n3024));
  jxor g02833(.dina(n3024), .dinb(n3007), .dout(n3025));
  jxor g02834(.dina(n3025), .dinb(n3003), .dout(n3026));
  jand g02835(.dina(n2883), .dinb(n2874), .dout(n3027));
  jand g02836(.dina(n2884), .dinb(n2871), .dout(n3028));
  jor  g02837(.dina(n3028), .dinb(n3027), .dout(n3029));
  jand g02838(.dina(n2787), .dinb(n2786), .dout(n3030));
  jand g02839(.dina(n2788), .dinb(n2785), .dout(n3031));
  jor  g02840(.dina(n3031), .dinb(n3030), .dout(n3032));
  jand g02841(.dina(n960), .dinb(\a[36] ), .dout(n3033));
  jand g02842(.dina(\a[38] ), .dinb(\a[0] ), .dout(n3034));
  jand g02843(.dina(\a[36] ), .dinb(\a[2] ), .dout(n3035));
  jor  g02844(.dina(n3035), .dinb(n3034), .dout(n3036));
  jand g02845(.dina(\a[38] ), .dinb(\a[2] ), .dout(n3037));
  jand g02846(.dina(n3037), .dinb(n2695), .dout(n3038));
  jnot g02847(.din(n3038), .dout(n3039));
  jand g02848(.dina(n3039), .dinb(n3036), .dout(n3040));
  jxor g02849(.dina(n3040), .dinb(n3033), .dout(n3041));
  jxor g02850(.dina(n3041), .dinb(n3032), .dout(n3042));
  jnot g02851(.din(n3042), .dout(n3043));
  jand g02852(.dina(\a[35] ), .dinb(\a[3] ), .dout(n3044));
  jnot g02853(.din(n3044), .dout(n3045));
  jand g02854(.dina(n1648), .dinb(n675), .dout(n3046));
  jnot g02855(.din(n3046), .dout(n3047));
  jand g02856(.dina(\a[25] ), .dinb(\a[13] ), .dout(n3048));
  jand g02857(.dina(\a[24] ), .dinb(\a[14] ), .dout(n3049));
  jor  g02858(.dina(n3049), .dinb(n3048), .dout(n3050));
  jand g02859(.dina(n3050), .dinb(n3047), .dout(n3051));
  jxor g02860(.dina(n3051), .dinb(n3045), .dout(n3052));
  jxor g02861(.dina(n3052), .dinb(n3043), .dout(n3053));
  jxor g02862(.dina(n3053), .dinb(n3029), .dout(n3054));
  jxor g02863(.dina(n3054), .dinb(n3026), .dout(n3055));
  jxor g02864(.dina(n3055), .dinb(n3000), .dout(n3056));
  jxor g02865(.dina(n3056), .dinb(n2979), .dout(n3057));
  jand g02866(.dina(n3057), .dinb(n2903), .dout(n3058));
  jor  g02867(.dina(n3057), .dinb(n2903), .dout(n3059));
  jnot g02868(.din(n3059), .dout(n3060));
  jor  g02869(.dina(n3060), .dinb(n3058), .dout(n3061));
  jnot g02870(.din(n2890), .dout(n3062));
  jor  g02871(.dina(n2899), .dinb(n2892), .dout(n3063));
  jand g02872(.dina(n3063), .dinb(n3062), .dout(n3064));
  jxor g02873(.dina(n3064), .dinb(n3061), .dout(\asquared[39] ));
  jand g02874(.dina(n2978), .dinb(n2906), .dout(n3066));
  jand g02875(.dina(n3056), .dinb(n2979), .dout(n3067));
  jor  g02876(.dina(n3067), .dinb(n3066), .dout(n3068));
  jand g02877(.dina(n2999), .dinb(n2982), .dout(n3069));
  jand g02878(.dina(n3055), .dinb(n3000), .dout(n3070));
  jor  g02879(.dina(n3070), .dinb(n3069), .dout(n3071));
  jand g02880(.dina(n3053), .dinb(n3029), .dout(n3072));
  jand g02881(.dina(n3054), .dinb(n3026), .dout(n3073));
  jor  g02882(.dina(n3073), .dinb(n3072), .dout(n3074));
  jand g02883(.dina(n2996), .dinb(n2993), .dout(n3075));
  jand g02884(.dina(n2997), .dinb(n2818), .dout(n3076));
  jor  g02885(.dina(n3076), .dinb(n3075), .dout(n3077));
  jand g02886(.dina(n2992), .dinb(n1181), .dout(n3078));
  jand g02887(.dina(\a[39] ), .dinb(\a[0] ), .dout(n3079));
  jxor g02888(.dina(n3079), .dinb(n3078), .dout(n3080));
  jand g02889(.dina(n1060), .dinb(\a[38] ), .dout(n3081));
  jnot g02890(.din(n3081), .dout(n3082));
  jand g02891(.dina(\a[38] ), .dinb(\a[1] ), .dout(n3083));
  jor  g02892(.dina(n3083), .dinb(\a[20] ), .dout(n3084));
  jand g02893(.dina(n3084), .dinb(n3082), .dout(n3085));
  jxor g02894(.dina(n3085), .dinb(n3080), .dout(n3086));
  jxor g02895(.dina(n3086), .dinb(n3077), .dout(n3087));
  jand g02896(.dina(n2918), .dinb(n2831), .dout(n3088));
  jand g02897(.dina(n2922), .dinb(n2919), .dout(n3089));
  jor  g02898(.dina(n3089), .dinb(n3088), .dout(n3090));
  jxor g02899(.dina(n3090), .dinb(n3087), .dout(n3091));
  jor  g02900(.dina(n2956), .dinb(n2950), .dout(n3092));
  jand g02901(.dina(n3040), .dinb(n3033), .dout(n3093));
  jor  g02902(.dina(n3093), .dinb(n3038), .dout(n3094));
  jand g02903(.dina(n3047), .dinb(n3045), .dout(n3095));
  jnot g02904(.din(n3095), .dout(n3096));
  jand g02905(.dina(n3096), .dinb(n3050), .dout(n3097));
  jxor g02906(.dina(n3097), .dinb(n3094), .dout(n3098));
  jxor g02907(.dina(n3098), .dinb(n3092), .dout(n3099));
  jor  g02908(.dina(n2964), .dinb(n2949), .dout(n3100));
  jor  g02909(.dina(n2975), .dinb(n2966), .dout(n3101));
  jand g02910(.dina(n3101), .dinb(n3100), .dout(n3102));
  jand g02911(.dina(n3041), .dinb(n3032), .dout(n3103));
  jnot g02912(.din(n3103), .dout(n3104));
  jor  g02913(.dina(n3052), .dinb(n3043), .dout(n3105));
  jand g02914(.dina(n3105), .dinb(n3104), .dout(n3106));
  jxor g02915(.dina(n3106), .dinb(n3102), .dout(n3107));
  jxor g02916(.dina(n3107), .dinb(n3099), .dout(n3108));
  jxor g02917(.dina(n3108), .dinb(n3091), .dout(n3109));
  jxor g02918(.dina(n3109), .dinb(n3074), .dout(n3110));
  jxor g02919(.dina(n3110), .dinb(n3071), .dout(n3111));
  jor  g02920(.dina(n2990), .dinb(n2986), .dout(n3112));
  jand g02921(.dina(n2998), .dinb(n2991), .dout(n3113));
  jnot g02922(.din(n3113), .dout(n3114));
  jand g02923(.dina(n3114), .dinb(n3112), .dout(n3115));
  jnot g02924(.din(n3115), .dout(n3116));
  jand g02925(.dina(\a[33] ), .dinb(\a[6] ), .dout(n3117));
  jand g02926(.dina(\a[32] ), .dinb(\a[30] ), .dout(n3118));
  jand g02927(.dina(n3118), .dinb(n684), .dout(n3119));
  jnot g02928(.din(n3119), .dout(n3120));
  jand g02929(.dina(n2671), .dinb(n410), .dout(n3121));
  jand g02930(.dina(\a[30] ), .dinb(\a[9] ), .dout(n3122));
  jand g02931(.dina(n3122), .dinb(n3117), .dout(n3123));
  jor  g02932(.dina(n3123), .dinb(n3121), .dout(n3124));
  jand g02933(.dina(n3124), .dinb(n3120), .dout(n3125));
  jnot g02934(.din(n3125), .dout(n3126));
  jand g02935(.dina(n3126), .dinb(n3117), .dout(n3127));
  jor  g02936(.dina(n3124), .dinb(n3119), .dout(n3128));
  jnot g02937(.din(n3128), .dout(n3129));
  jand g02938(.dina(\a[32] ), .dinb(\a[7] ), .dout(n3130));
  jor  g02939(.dina(n3130), .dinb(n3122), .dout(n3131));
  jand g02940(.dina(n3131), .dinb(n3129), .dout(n3132));
  jor  g02941(.dina(n3132), .dinb(n3127), .dout(n3133));
  jand g02942(.dina(\a[36] ), .dinb(\a[3] ), .dout(n3134));
  jand g02943(.dina(\a[26] ), .dinb(\a[13] ), .dout(n3135));
  jand g02944(.dina(n3135), .dinb(n3134), .dout(n3136));
  jnot g02945(.din(n3136), .dout(n3137));
  jand g02946(.dina(\a[37] ), .dinb(\a[36] ), .dout(n3138));
  jand g02947(.dina(n3138), .dinb(n248), .dout(n3139));
  jand g02948(.dina(\a[37] ), .dinb(\a[2] ), .dout(n3140));
  jand g02949(.dina(n3140), .dinb(n3135), .dout(n3141));
  jor  g02950(.dina(n3141), .dinb(n3139), .dout(n3142));
  jnot g02951(.din(n3142), .dout(n3143));
  jand g02952(.dina(n3143), .dinb(n3137), .dout(n3144));
  jor  g02953(.dina(n3135), .dinb(n3134), .dout(n3145));
  jand g02954(.dina(n3145), .dinb(n3144), .dout(n3146));
  jand g02955(.dina(n3142), .dinb(n3137), .dout(n3147));
  jnot g02956(.din(n3147), .dout(n3148));
  jand g02957(.dina(n3148), .dinb(n3140), .dout(n3149));
  jor  g02958(.dina(n3149), .dinb(n3146), .dout(n3150));
  jand g02959(.dina(\a[25] ), .dinb(\a[14] ), .dout(n3151));
  jnot g02960(.din(n3151), .dout(n3152));
  jand g02961(.dina(n1942), .dinb(n829), .dout(n3153));
  jnot g02962(.din(n3153), .dout(n3154));
  jand g02963(.dina(\a[24] ), .dinb(\a[15] ), .dout(n3155));
  jand g02964(.dina(\a[23] ), .dinb(\a[16] ), .dout(n3156));
  jor  g02965(.dina(n3156), .dinb(n3155), .dout(n3157));
  jand g02966(.dina(n3157), .dinb(n3154), .dout(n3158));
  jxor g02967(.dina(n3158), .dinb(n3152), .dout(n3159));
  jnot g02968(.din(n3159), .dout(n3160));
  jxor g02969(.dina(n3160), .dinb(n3150), .dout(n3161));
  jxor g02970(.dina(n3161), .dinb(n3133), .dout(n3162));
  jxor g02971(.dina(n3162), .dinb(n3116), .dout(n3163));
  jnot g02972(.din(n3163), .dout(n3164));
  jor  g02973(.dina(n2928), .dinb(n2924), .dout(n3165));
  jand g02974(.dina(n2976), .dinb(n2929), .dout(n3166));
  jnot g02975(.din(n3166), .dout(n3167));
  jand g02976(.dina(n3167), .dinb(n3165), .dout(n3168));
  jxor g02977(.dina(n3168), .dinb(n3164), .dout(n3169));
  jand g02978(.dina(n2914), .dinb(n2911), .dout(n3170));
  jand g02979(.dina(n2977), .dinb(n2915), .dout(n3171));
  jor  g02980(.dina(n3171), .dinb(n3170), .dout(n3172));
  jand g02981(.dina(n2970), .dinb(n2968), .dout(n3173));
  jnot g02982(.din(n3173), .dout(n3174));
  jand g02983(.dina(n3174), .dinb(n2973), .dout(n3175));
  jxor g02984(.dina(n3175), .dinb(n3019), .dout(n3176));
  jxor g02985(.dina(n3176), .dinb(n2943), .dout(n3177));
  jand g02986(.dina(n3024), .dinb(n3007), .dout(n3178));
  jand g02987(.dina(n3025), .dinb(n3003), .dout(n3179));
  jor  g02988(.dina(n3179), .dinb(n3178), .dout(n3180));
  jxor g02989(.dina(n3180), .dinb(n3177), .dout(n3181));
  jand g02990(.dina(\a[28] ), .dinb(\a[11] ), .dout(n3182));
  jand g02991(.dina(\a[34] ), .dinb(\a[29] ), .dout(n3183));
  jand g02992(.dina(n3183), .dinb(n619), .dout(n3184));
  jnot g02993(.din(n3184), .dout(n3185));
  jand g02994(.dina(\a[34] ), .dinb(\a[5] ), .dout(n3186));
  jand g02995(.dina(n3186), .dinb(n3182), .dout(n3187));
  jand g02996(.dina(n2653), .dinb(n655), .dout(n3188));
  jor  g02997(.dina(n3188), .dinb(n3187), .dout(n3189));
  jand g02998(.dina(n3189), .dinb(n3185), .dout(n3190));
  jnot g02999(.din(n3190), .dout(n3191));
  jand g03000(.dina(n3191), .dinb(n3182), .dout(n3192));
  jor  g03001(.dina(n3189), .dinb(n3184), .dout(n3193));
  jnot g03002(.din(n3193), .dout(n3194));
  jand g03003(.dina(\a[29] ), .dinb(\a[10] ), .dout(n3195));
  jor  g03004(.dina(n3195), .dinb(n3186), .dout(n3196));
  jand g03005(.dina(n3196), .dinb(n3194), .dout(n3197));
  jor  g03006(.dina(n3197), .dinb(n3192), .dout(n3198));
  jand g03007(.dina(\a[22] ), .dinb(\a[17] ), .dout(n3199));
  jand g03008(.dina(\a[35] ), .dinb(\a[4] ), .dout(n3200));
  jand g03009(.dina(\a[27] ), .dinb(\a[12] ), .dout(n3201));
  jxor g03010(.dina(n3201), .dinb(n3200), .dout(n3202));
  jxor g03011(.dina(n3202), .dinb(n3199), .dout(n3203));
  jnot g03012(.din(n3203), .dout(n3204));
  jand g03013(.dina(\a[31] ), .dinb(\a[8] ), .dout(n3205));
  jnot g03014(.din(n3205), .dout(n3206));
  jand g03015(.dina(n1490), .dinb(n1024), .dout(n3207));
  jnot g03016(.din(n3207), .dout(n3208));
  jand g03017(.dina(\a[21] ), .dinb(\a[18] ), .dout(n3209));
  jor  g03018(.dina(n3209), .dinb(n1287), .dout(n3210));
  jand g03019(.dina(n3210), .dinb(n3208), .dout(n3211));
  jxor g03020(.dina(n3211), .dinb(n3206), .dout(n3212));
  jxor g03021(.dina(n3212), .dinb(n3204), .dout(n3213));
  jxor g03022(.dina(n3213), .dinb(n3198), .dout(n3214));
  jxor g03023(.dina(n3214), .dinb(n3181), .dout(n3215));
  jxor g03024(.dina(n3215), .dinb(n3172), .dout(n3216));
  jxor g03025(.dina(n3216), .dinb(n3169), .dout(n3217));
  jxor g03026(.dina(n3217), .dinb(n3111), .dout(n3218));
  jand g03027(.dina(n3218), .dinb(n3068), .dout(n3219));
  jor  g03028(.dina(n3218), .dinb(n3068), .dout(n3220));
  jnot g03029(.din(n3220), .dout(n3221));
  jor  g03030(.dina(n3221), .dinb(n3219), .dout(n3222));
  jnot g03031(.din(n3058), .dout(n3223));
  jor  g03032(.dina(n3064), .dinb(n3060), .dout(n3224));
  jand g03033(.dina(n3224), .dinb(n3223), .dout(n3225));
  jxor g03034(.dina(n3225), .dinb(n3222), .dout(\asquared[40] ));
  jand g03035(.dina(n3110), .dinb(n3071), .dout(n3227));
  jand g03036(.dina(n3217), .dinb(n3111), .dout(n3228));
  jor  g03037(.dina(n3228), .dinb(n3227), .dout(n3229));
  jand g03038(.dina(n3154), .dinb(n3152), .dout(n3230));
  jnot g03039(.din(n3230), .dout(n3231));
  jand g03040(.dina(n3231), .dinb(n3157), .dout(n3232));
  jxor g03041(.dina(n3232), .dinb(n3128), .dout(n3233));
  jand g03042(.dina(n3079), .dinb(n3078), .dout(n3234));
  jand g03043(.dina(n3085), .dinb(n3080), .dout(n3235));
  jor  g03044(.dina(n3235), .dinb(n3234), .dout(n3236));
  jxor g03045(.dina(n3236), .dinb(n3233), .dout(n3237));
  jand g03046(.dina(n3086), .dinb(n3077), .dout(n3238));
  jand g03047(.dina(n3090), .dinb(n3087), .dout(n3239));
  jor  g03048(.dina(n3239), .dinb(n3238), .dout(n3240));
  jxor g03049(.dina(n3240), .dinb(n3237), .dout(n3241));
  jand g03050(.dina(\a[36] ), .dinb(\a[4] ), .dout(n3242));
  jand g03051(.dina(\a[36] ), .dinb(\a[35] ), .dout(n3243));
  jand g03052(.dina(n3243), .dinb(n242), .dout(n3244));
  jand g03053(.dina(\a[28] ), .dinb(\a[12] ), .dout(n3245));
  jand g03054(.dina(n3245), .dinb(n3242), .dout(n3246));
  jor  g03055(.dina(n3246), .dinb(n3244), .dout(n3247));
  jand g03056(.dina(\a[35] ), .dinb(\a[5] ), .dout(n3248));
  jand g03057(.dina(n3248), .dinb(n3245), .dout(n3249));
  jnot g03058(.din(n3249), .dout(n3250));
  jand g03059(.dina(n3250), .dinb(n3247), .dout(n3251));
  jnot g03060(.din(n3251), .dout(n3252));
  jand g03061(.dina(n3252), .dinb(n3242), .dout(n3253));
  jor  g03062(.dina(n3249), .dinb(n3247), .dout(n3254));
  jnot g03063(.din(n3254), .dout(n3255));
  jor  g03064(.dina(n3248), .dinb(n3245), .dout(n3256));
  jand g03065(.dina(n3256), .dinb(n3255), .dout(n3257));
  jor  g03066(.dina(n3257), .dinb(n3253), .dout(n3258));
  jand g03067(.dina(\a[40] ), .dinb(\a[0] ), .dout(n3259));
  jor  g03068(.dina(n3259), .dinb(n3037), .dout(n3260));
  jand g03069(.dina(\a[40] ), .dinb(\a[2] ), .dout(n3261));
  jand g03070(.dina(n3261), .dinb(n3034), .dout(n3262));
  jnot g03071(.din(n3262), .dout(n3263));
  jand g03072(.dina(n3263), .dinb(n3260), .dout(n3264));
  jxor g03073(.dina(n3264), .dinb(n1258), .dout(n3265));
  jnot g03074(.din(n3265), .dout(n3266));
  jand g03075(.dina(\a[33] ), .dinb(\a[7] ), .dout(n3267));
  jnot g03076(.din(n3267), .dout(n3268));
  jand g03077(.dina(\a[32] ), .dinb(\a[31] ), .dout(n3269));
  jand g03078(.dina(n3269), .dinb(n395), .dout(n3270));
  jnot g03079(.din(n3270), .dout(n3271));
  jand g03080(.dina(\a[31] ), .dinb(\a[9] ), .dout(n3272));
  jand g03081(.dina(\a[32] ), .dinb(\a[8] ), .dout(n3273));
  jor  g03082(.dina(n3273), .dinb(n3272), .dout(n3274));
  jand g03083(.dina(n3274), .dinb(n3271), .dout(n3275));
  jxor g03084(.dina(n3275), .dinb(n3268), .dout(n3276));
  jxor g03085(.dina(n3276), .dinb(n3266), .dout(n3277));
  jxor g03086(.dina(n3277), .dinb(n3258), .dout(n3278));
  jxor g03087(.dina(n3278), .dinb(n3241), .dout(n3279));
  jand g03088(.dina(n3108), .dinb(n3091), .dout(n3280));
  jand g03089(.dina(n3109), .dinb(n3074), .dout(n3281));
  jor  g03090(.dina(n3281), .dinb(n3280), .dout(n3282));
  jxor g03091(.dina(n3282), .dinb(n3279), .dout(n3283));
  jor  g03092(.dina(n3106), .dinb(n3102), .dout(n3284));
  jand g03093(.dina(n3107), .dinb(n3099), .dout(n3285));
  jnot g03094(.din(n3285), .dout(n3286));
  jand g03095(.dina(n3286), .dinb(n3284), .dout(n3287));
  jnot g03096(.din(n3287), .dout(n3288));
  jand g03097(.dina(\a[29] ), .dinb(\a[11] ), .dout(n3289));
  jand g03098(.dina(\a[30] ), .dinb(\a[10] ), .dout(n3290));
  jand g03099(.dina(\a[34] ), .dinb(\a[6] ), .dout(n3291));
  jand g03100(.dina(n3291), .dinb(n3290), .dout(n3292));
  jnot g03101(.din(n3292), .dout(n3293));
  jand g03102(.dina(\a[30] ), .dinb(\a[29] ), .dout(n3294));
  jand g03103(.dina(n3294), .dinb(n655), .dout(n3295));
  jand g03104(.dina(n3291), .dinb(n3289), .dout(n3296));
  jor  g03105(.dina(n3296), .dinb(n3295), .dout(n3297));
  jand g03106(.dina(n3297), .dinb(n3293), .dout(n3298));
  jnot g03107(.din(n3298), .dout(n3299));
  jand g03108(.dina(n3299), .dinb(n3289), .dout(n3300));
  jor  g03109(.dina(n3297), .dinb(n3292), .dout(n3301));
  jnot g03110(.din(n3301), .dout(n3302));
  jor  g03111(.dina(n3291), .dinb(n3290), .dout(n3303));
  jand g03112(.dina(n3303), .dinb(n3302), .dout(n3304));
  jor  g03113(.dina(n3304), .dinb(n3300), .dout(n3305));
  jand g03114(.dina(\a[37] ), .dinb(\a[3] ), .dout(n3306));
  jand g03115(.dina(\a[27] ), .dinb(\a[13] ), .dout(n3307));
  jand g03116(.dina(\a[26] ), .dinb(\a[14] ), .dout(n3308));
  jor  g03117(.dina(n3308), .dinb(n3307), .dout(n3309));
  jand g03118(.dina(n1927), .dinb(n675), .dout(n3310));
  jnot g03119(.din(n3310), .dout(n3311));
  jand g03120(.dina(n3311), .dinb(n3309), .dout(n3312));
  jxor g03121(.dina(n3312), .dinb(n3306), .dout(n3313));
  jnot g03122(.din(n3313), .dout(n3314));
  jand g03123(.dina(\a[25] ), .dinb(\a[15] ), .dout(n3315));
  jnot g03124(.din(n3315), .dout(n3316));
  jand g03125(.dina(n1942), .dinb(n937), .dout(n3317));
  jnot g03126(.din(n3317), .dout(n3318));
  jand g03127(.dina(\a[23] ), .dinb(\a[17] ), .dout(n3319));
  jand g03128(.dina(\a[24] ), .dinb(\a[16] ), .dout(n3320));
  jor  g03129(.dina(n3320), .dinb(n3319), .dout(n3321));
  jand g03130(.dina(n3321), .dinb(n3318), .dout(n3322));
  jxor g03131(.dina(n3322), .dinb(n3316), .dout(n3323));
  jxor g03132(.dina(n3323), .dinb(n3314), .dout(n3324));
  jxor g03133(.dina(n3324), .dinb(n3305), .dout(n3325));
  jxor g03134(.dina(n3325), .dinb(n3288), .dout(n3326));
  jand g03135(.dina(n3175), .dinb(n3019), .dout(n3327));
  jand g03136(.dina(n3176), .dinb(n2943), .dout(n3328));
  jor  g03137(.dina(n3328), .dinb(n3327), .dout(n3329));
  jand g03138(.dina(n3097), .dinb(n3094), .dout(n3330));
  jand g03139(.dina(n3098), .dinb(n3092), .dout(n3331));
  jor  g03140(.dina(n3331), .dinb(n3330), .dout(n3332));
  jxor g03141(.dina(n3332), .dinb(n3329), .dout(n3333));
  jand g03142(.dina(\a[21] ), .dinb(\a[19] ), .dout(n3334));
  jand g03143(.dina(\a[39] ), .dinb(\a[1] ), .dout(n3335));
  jxor g03144(.dina(n3335), .dinb(n3334), .dout(n3336));
  jxor g03145(.dina(n3336), .dinb(n3081), .dout(n3337));
  jand g03146(.dina(n3208), .dinb(n3206), .dout(n3338));
  jnot g03147(.din(n3338), .dout(n3339));
  jand g03148(.dina(n3339), .dinb(n3210), .dout(n3340));
  jxor g03149(.dina(n3340), .dinb(n3337), .dout(n3341));
  jxor g03150(.dina(n3341), .dinb(n3333), .dout(n3342));
  jxor g03151(.dina(n3342), .dinb(n3326), .dout(n3343));
  jxor g03152(.dina(n3343), .dinb(n3283), .dout(n3344));
  jand g03153(.dina(n3162), .dinb(n3116), .dout(n3345));
  jnot g03154(.din(n3345), .dout(n3346));
  jor  g03155(.dina(n3168), .dinb(n3164), .dout(n3347));
  jand g03156(.dina(n3347), .dinb(n3346), .dout(n3348));
  jnot g03157(.din(n3348), .dout(n3349));
  jand g03158(.dina(n3180), .dinb(n3177), .dout(n3350));
  jand g03159(.dina(n3214), .dinb(n3181), .dout(n3351));
  jor  g03160(.dina(n3351), .dinb(n3350), .dout(n3352));
  jand g03161(.dina(n3201), .dinb(n3200), .dout(n3353));
  jand g03162(.dina(n3202), .dinb(n3199), .dout(n3354));
  jor  g03163(.dina(n3354), .dinb(n3353), .dout(n3355));
  jxor g03164(.dina(n3194), .dinb(n3144), .dout(n3356));
  jxor g03165(.dina(n3356), .dinb(n3355), .dout(n3357));
  jor  g03166(.dina(n3212), .dinb(n3204), .dout(n3358));
  jand g03167(.dina(n3213), .dinb(n3198), .dout(n3359));
  jnot g03168(.din(n3359), .dout(n3360));
  jand g03169(.dina(n3360), .dinb(n3358), .dout(n3361));
  jnot g03170(.din(n3361), .dout(n3362));
  jand g03171(.dina(n3160), .dinb(n3150), .dout(n3363));
  jand g03172(.dina(n3161), .dinb(n3133), .dout(n3364));
  jor  g03173(.dina(n3364), .dinb(n3363), .dout(n3365));
  jxor g03174(.dina(n3365), .dinb(n3362), .dout(n3366));
  jxor g03175(.dina(n3366), .dinb(n3357), .dout(n3367));
  jxor g03176(.dina(n3367), .dinb(n3352), .dout(n3368));
  jxor g03177(.dina(n3368), .dinb(n3349), .dout(n3369));
  jand g03178(.dina(n3215), .dinb(n3172), .dout(n3370));
  jand g03179(.dina(n3216), .dinb(n3169), .dout(n3371));
  jor  g03180(.dina(n3371), .dinb(n3370), .dout(n3372));
  jxor g03181(.dina(n3372), .dinb(n3369), .dout(n3373));
  jxor g03182(.dina(n3373), .dinb(n3344), .dout(n3374));
  jand g03183(.dina(n3374), .dinb(n3229), .dout(n3375));
  jor  g03184(.dina(n3374), .dinb(n3229), .dout(n3376));
  jnot g03185(.din(n3376), .dout(n3377));
  jor  g03186(.dina(n3377), .dinb(n3375), .dout(n3378));
  jnot g03187(.din(n3219), .dout(n3379));
  jor  g03188(.dina(n3225), .dinb(n3221), .dout(n3380));
  jand g03189(.dina(n3380), .dinb(n3379), .dout(n3381));
  jxor g03190(.dina(n3381), .dinb(n3378), .dout(\asquared[41] ));
  jand g03191(.dina(n3372), .dinb(n3369), .dout(n3383));
  jand g03192(.dina(n3373), .dinb(n3344), .dout(n3384));
  jor  g03193(.dina(n3384), .dinb(n3383), .dout(n3385));
  jnot g03194(.din(n3385), .dout(n3386));
  jand g03195(.dina(n3325), .dinb(n3288), .dout(n3387));
  jand g03196(.dina(n3342), .dinb(n3326), .dout(n3388));
  jor  g03197(.dina(n3388), .dinb(n3387), .dout(n3389));
  jand g03198(.dina(n3240), .dinb(n3237), .dout(n3390));
  jand g03199(.dina(n3278), .dinb(n3241), .dout(n3391));
  jor  g03200(.dina(n3391), .dinb(n3390), .dout(n3392));
  jand g03201(.dina(n3312), .dinb(n3306), .dout(n3393));
  jor  g03202(.dina(n3393), .dinb(n3310), .dout(n3394));
  jand g03203(.dina(n3264), .dinb(n1258), .dout(n3395));
  jor  g03204(.dina(n3395), .dinb(n3262), .dout(n3396));
  jand g03205(.dina(n3318), .dinb(n3316), .dout(n3397));
  jnot g03206(.din(n3397), .dout(n3398));
  jand g03207(.dina(n3398), .dinb(n3321), .dout(n3399));
  jxor g03208(.dina(n3399), .dinb(n3396), .dout(n3400));
  jxor g03209(.dina(n3400), .dinb(n3394), .dout(n3401));
  jnot g03210(.din(n3401), .dout(n3402));
  jor  g03211(.dina(n3276), .dinb(n3266), .dout(n3403));
  jand g03212(.dina(n3277), .dinb(n3258), .dout(n3404));
  jnot g03213(.din(n3404), .dout(n3405));
  jand g03214(.dina(n3405), .dinb(n3403), .dout(n3406));
  jxor g03215(.dina(n3406), .dinb(n3402), .dout(n3407));
  jand g03216(.dina(n1152), .dinb(\a[40] ), .dout(n3408));
  jnot g03217(.din(n3408), .dout(n3409));
  jand g03218(.dina(\a[40] ), .dinb(\a[1] ), .dout(n3410));
  jor  g03219(.dina(n3410), .dinb(\a[21] ), .dout(n3411));
  jand g03220(.dina(n3411), .dinb(n3409), .dout(n3412));
  jand g03221(.dina(n3271), .dinb(n3268), .dout(n3413));
  jnot g03222(.din(n3413), .dout(n3414));
  jand g03223(.dina(n3414), .dinb(n3274), .dout(n3415));
  jxor g03224(.dina(n3415), .dinb(n3412), .dout(n3416));
  jxor g03225(.dina(n3416), .dinb(n3301), .dout(n3417));
  jxor g03226(.dina(n3417), .dinb(n3407), .dout(n3418));
  jxor g03227(.dina(n3418), .dinb(n3392), .dout(n3419));
  jxor g03228(.dina(n3419), .dinb(n3389), .dout(n3420));
  jand g03229(.dina(n3282), .dinb(n3279), .dout(n3421));
  jand g03230(.dina(n3343), .dinb(n3283), .dout(n3422));
  jor  g03231(.dina(n3422), .dinb(n3421), .dout(n3423));
  jxor g03232(.dina(n3423), .dinb(n3420), .dout(n3424));
  jand g03233(.dina(n3232), .dinb(n3128), .dout(n3425));
  jand g03234(.dina(n3236), .dinb(n3233), .dout(n3426));
  jor  g03235(.dina(n3426), .dinb(n3425), .dout(n3427));
  jnot g03236(.din(n3144), .dout(n3428));
  jand g03237(.dina(n3193), .dinb(n3428), .dout(n3429));
  jand g03238(.dina(n3356), .dinb(n3355), .dout(n3430));
  jor  g03239(.dina(n3430), .dinb(n3429), .dout(n3431));
  jxor g03240(.dina(n3431), .dinb(n3427), .dout(n3432));
  jnot g03241(.din(n3432), .dout(n3433));
  jor  g03242(.dina(n3323), .dinb(n3314), .dout(n3434));
  jand g03243(.dina(n3324), .dinb(n3305), .dout(n3435));
  jnot g03244(.din(n3435), .dout(n3436));
  jand g03245(.dina(n3436), .dinb(n3434), .dout(n3437));
  jxor g03246(.dina(n3437), .dinb(n3433), .dout(n3438));
  jand g03247(.dina(n3365), .dinb(n3362), .dout(n3439));
  jand g03248(.dina(n3366), .dinb(n3357), .dout(n3440));
  jor  g03249(.dina(n3440), .dinb(n3439), .dout(n3441));
  jand g03250(.dina(n3335), .dinb(n3334), .dout(n3442));
  jand g03251(.dina(\a[41] ), .dinb(\a[2] ), .dout(n3443));
  jand g03252(.dina(n3443), .dinb(n3079), .dout(n3444));
  jnot g03253(.din(n3444), .dout(n3445));
  jand g03254(.dina(\a[41] ), .dinb(\a[0] ), .dout(n3446));
  jand g03255(.dina(\a[39] ), .dinb(\a[2] ), .dout(n3447));
  jor  g03256(.dina(n3447), .dinb(n3446), .dout(n3448));
  jand g03257(.dina(n3448), .dinb(n3445), .dout(n3449));
  jxor g03258(.dina(n3449), .dinb(n3442), .dout(n3450));
  jxor g03259(.dina(n3450), .dinb(n3254), .dout(n3451));
  jnot g03260(.din(n3451), .dout(n3452));
  jand g03261(.dina(\a[38] ), .dinb(\a[3] ), .dout(n3453));
  jnot g03262(.din(n3453), .dout(n3454));
  jand g03263(.dina(\a[28] ), .dinb(\a[26] ), .dout(n3455));
  jand g03264(.dina(n3455), .dinb(n727), .dout(n3456));
  jnot g03265(.din(n3456), .dout(n3457));
  jand g03266(.dina(\a[28] ), .dinb(\a[13] ), .dout(n3458));
  jand g03267(.dina(\a[26] ), .dinb(\a[15] ), .dout(n3459));
  jor  g03268(.dina(n3459), .dinb(n3458), .dout(n3460));
  jand g03269(.dina(n3460), .dinb(n3457), .dout(n3461));
  jxor g03270(.dina(n3461), .dinb(n3454), .dout(n3462));
  jxor g03271(.dina(n3462), .dinb(n3452), .dout(n3463));
  jxor g03272(.dina(n3463), .dinb(n3441), .dout(n3464));
  jxor g03273(.dina(n3464), .dinb(n3438), .dout(n3465));
  jand g03274(.dina(n3367), .dinb(n3352), .dout(n3466));
  jand g03275(.dina(n3368), .dinb(n3349), .dout(n3467));
  jor  g03276(.dina(n3467), .dinb(n3466), .dout(n3468));
  jand g03277(.dina(n3336), .dinb(n3081), .dout(n3469));
  jand g03278(.dina(n3340), .dinb(n3337), .dout(n3470));
  jor  g03279(.dina(n3470), .dinb(n3469), .dout(n3471));
  jand g03280(.dina(\a[36] ), .dinb(\a[5] ), .dout(n3472));
  jand g03281(.dina(\a[35] ), .dinb(\a[6] ), .dout(n3473));
  jand g03282(.dina(\a[30] ), .dinb(\a[11] ), .dout(n3474));
  jor  g03283(.dina(n3474), .dinb(n3473), .dout(n3475));
  jand g03284(.dina(\a[35] ), .dinb(\a[30] ), .dout(n3476));
  jand g03285(.dina(n3476), .dinb(n725), .dout(n3477));
  jnot g03286(.din(n3477), .dout(n3478));
  jand g03287(.dina(n3478), .dinb(n3475), .dout(n3479));
  jxor g03288(.dina(n3479), .dinb(n3472), .dout(n3480));
  jand g03289(.dina(\a[33] ), .dinb(\a[8] ), .dout(n3481));
  jand g03290(.dina(\a[22] ), .dinb(\a[19] ), .dout(n3482));
  jxor g03291(.dina(n3482), .dinb(n1490), .dout(n3483));
  jxor g03292(.dina(n3483), .dinb(n3481), .dout(n3484));
  jxor g03293(.dina(n3484), .dinb(n3480), .dout(n3485));
  jxor g03294(.dina(n3485), .dinb(n3471), .dout(n3486));
  jand g03295(.dina(n3332), .dinb(n3329), .dout(n3487));
  jand g03296(.dina(n3341), .dinb(n3333), .dout(n3488));
  jor  g03297(.dina(n3488), .dinb(n3487), .dout(n3489));
  jxor g03298(.dina(n3489), .dinb(n3486), .dout(n3490));
  jand g03299(.dina(\a[31] ), .dinb(\a[10] ), .dout(n3491));
  jand g03300(.dina(\a[34] ), .dinb(\a[32] ), .dout(n3492));
  jand g03301(.dina(n3492), .dinb(n684), .dout(n3493));
  jnot g03302(.din(n3493), .dout(n3494));
  jand g03303(.dina(n3269), .dinb(n453), .dout(n3495));
  jand g03304(.dina(\a[34] ), .dinb(\a[7] ), .dout(n3496));
  jand g03305(.dina(n3496), .dinb(n3491), .dout(n3497));
  jor  g03306(.dina(n3497), .dinb(n3495), .dout(n3498));
  jand g03307(.dina(n3498), .dinb(n3494), .dout(n3499));
  jnot g03308(.din(n3499), .dout(n3500));
  jand g03309(.dina(n3500), .dinb(n3491), .dout(n3501));
  jor  g03310(.dina(n3498), .dinb(n3493), .dout(n3502));
  jnot g03311(.din(n3502), .dout(n3503));
  jand g03312(.dina(\a[32] ), .dinb(\a[9] ), .dout(n3504));
  jor  g03313(.dina(n3504), .dinb(n3496), .dout(n3505));
  jand g03314(.dina(n3505), .dinb(n3503), .dout(n3506));
  jor  g03315(.dina(n3506), .dinb(n3501), .dout(n3507));
  jand g03316(.dina(\a[27] ), .dinb(\a[14] ), .dout(n3508));
  jand g03317(.dina(\a[37] ), .dinb(\a[4] ), .dout(n3509));
  jand g03318(.dina(\a[29] ), .dinb(\a[12] ), .dout(n3510));
  jxor g03319(.dina(n3510), .dinb(n3509), .dout(n3511));
  jxor g03320(.dina(n3511), .dinb(n3508), .dout(n3512));
  jand g03321(.dina(\a[25] ), .dinb(\a[16] ), .dout(n3513));
  jand g03322(.dina(n1942), .dinb(n1107), .dout(n3514));
  jnot g03323(.din(n3514), .dout(n3515));
  jand g03324(.dina(\a[24] ), .dinb(\a[17] ), .dout(n3516));
  jand g03325(.dina(\a[23] ), .dinb(\a[18] ), .dout(n3517));
  jor  g03326(.dina(n3517), .dinb(n3516), .dout(n3518));
  jand g03327(.dina(n3518), .dinb(n3515), .dout(n3519));
  jxor g03328(.dina(n3519), .dinb(n3513), .dout(n3520));
  jxor g03329(.dina(n3520), .dinb(n3512), .dout(n3521));
  jxor g03330(.dina(n3521), .dinb(n3507), .dout(n3522));
  jxor g03331(.dina(n3522), .dinb(n3490), .dout(n3523));
  jxor g03332(.dina(n3523), .dinb(n3468), .dout(n3524));
  jxor g03333(.dina(n3524), .dinb(n3465), .dout(n3525));
  jxor g03334(.dina(n3525), .dinb(n3424), .dout(n3526));
  jxor g03335(.dina(n3526), .dinb(n3386), .dout(n3527));
  jnot g03336(.din(n3375), .dout(n3528));
  jor  g03337(.dina(n3381), .dinb(n3377), .dout(n3529));
  jand g03338(.dina(n3529), .dinb(n3528), .dout(n3530));
  jxor g03339(.dina(n3530), .dinb(n3527), .dout(\asquared[42] ));
  jand g03340(.dina(n3423), .dinb(n3420), .dout(n3532));
  jand g03341(.dina(n3525), .dinb(n3424), .dout(n3533));
  jor  g03342(.dina(n3533), .dinb(n3532), .dout(n3534));
  jand g03343(.dina(n3523), .dinb(n3468), .dout(n3535));
  jand g03344(.dina(n3524), .dinb(n3465), .dout(n3536));
  jor  g03345(.dina(n3536), .dinb(n3535), .dout(n3537));
  jand g03346(.dina(n3463), .dinb(n3441), .dout(n3538));
  jand g03347(.dina(n3464), .dinb(n3438), .dout(n3539));
  jor  g03348(.dina(n3539), .dinb(n3538), .dout(n3540));
  jand g03349(.dina(n3399), .dinb(n3396), .dout(n3541));
  jand g03350(.dina(n3400), .dinb(n3394), .dout(n3542));
  jor  g03351(.dina(n3542), .dinb(n3541), .dout(n3543));
  jnot g03352(.din(n3543), .dout(n3544));
  jand g03353(.dina(n3450), .dinb(n3254), .dout(n3545));
  jnot g03354(.din(n3545), .dout(n3546));
  jor  g03355(.dina(n3462), .dinb(n3452), .dout(n3547));
  jand g03356(.dina(n3547), .dinb(n3546), .dout(n3548));
  jxor g03357(.dina(n3548), .dinb(n3544), .dout(n3549));
  jand g03358(.dina(n3520), .dinb(n3512), .dout(n3550));
  jand g03359(.dina(n3521), .dinb(n3507), .dout(n3551));
  jor  g03360(.dina(n3551), .dinb(n3550), .dout(n3552));
  jxor g03361(.dina(n3552), .dinb(n3549), .dout(n3553));
  jand g03362(.dina(n3489), .dinb(n3486), .dout(n3554));
  jand g03363(.dina(n3522), .dinb(n3490), .dout(n3555));
  jor  g03364(.dina(n3555), .dinb(n3554), .dout(n3556));
  jxor g03365(.dina(n3556), .dinb(n3553), .dout(n3557));
  jxor g03366(.dina(n3557), .dinb(n3540), .dout(n3558));
  jxor g03367(.dina(n3558), .dinb(n3537), .dout(n3559));
  jand g03368(.dina(n3415), .dinb(n3412), .dout(n3560));
  jand g03369(.dina(n3416), .dinb(n3301), .dout(n3561));
  jor  g03370(.dina(n3561), .dinb(n3560), .dout(n3562));
  jand g03371(.dina(\a[29] ), .dinb(\a[13] ), .dout(n3563));
  jand g03372(.dina(\a[30] ), .dinb(\a[12] ), .dout(n3564));
  jand g03373(.dina(\a[37] ), .dinb(\a[5] ), .dout(n3565));
  jand g03374(.dina(n3565), .dinb(n3564), .dout(n3566));
  jnot g03375(.din(n3566), .dout(n3567));
  jand g03376(.dina(n3294), .dinb(n899), .dout(n3568));
  jand g03377(.dina(n3565), .dinb(n3563), .dout(n3569));
  jor  g03378(.dina(n3569), .dinb(n3568), .dout(n3570));
  jand g03379(.dina(n3570), .dinb(n3567), .dout(n3571));
  jnot g03380(.din(n3571), .dout(n3572));
  jand g03381(.dina(n3572), .dinb(n3563), .dout(n3573));
  jor  g03382(.dina(n3570), .dinb(n3566), .dout(n3574));
  jnot g03383(.din(n3574), .dout(n3575));
  jor  g03384(.dina(n3565), .dinb(n3564), .dout(n3576));
  jand g03385(.dina(n3576), .dinb(n3575), .dout(n3577));
  jor  g03386(.dina(n3577), .dinb(n3573), .dout(n3578));
  jand g03387(.dina(\a[42] ), .dinb(\a[0] ), .dout(n3579));
  jxor g03388(.dina(n3579), .dinb(n3408), .dout(n3580));
  jand g03389(.dina(\a[22] ), .dinb(\a[20] ), .dout(n3581));
  jand g03390(.dina(\a[41] ), .dinb(\a[1] ), .dout(n3582));
  jxor g03391(.dina(n3582), .dinb(n3581), .dout(n3583));
  jxor g03392(.dina(n3583), .dinb(n3580), .dout(n3584));
  jxor g03393(.dina(n3584), .dinb(n3578), .dout(n3585));
  jxor g03394(.dina(n3585), .dinb(n3562), .dout(n3586));
  jnot g03395(.din(n3586), .dout(n3587));
  jor  g03396(.dina(n3406), .dinb(n3402), .dout(n3588));
  jand g03397(.dina(n3417), .dinb(n3407), .dout(n3589));
  jnot g03398(.din(n3589), .dout(n3590));
  jand g03399(.dina(n3590), .dinb(n3588), .dout(n3591));
  jxor g03400(.dina(n3591), .dinb(n3587), .dout(n3592));
  jand g03401(.dina(n3479), .dinb(n3472), .dout(n3593));
  jor  g03402(.dina(n3593), .dinb(n3477), .dout(n3594));
  jand g03403(.dina(n3510), .dinb(n3509), .dout(n3595));
  jand g03404(.dina(n3511), .dinb(n3508), .dout(n3596));
  jor  g03405(.dina(n3596), .dinb(n3595), .dout(n3597));
  jor  g03406(.dina(n3482), .dinb(n1490), .dout(n3598));
  jand g03407(.dina(n3482), .dinb(n1490), .dout(n3599));
  jor  g03408(.dina(n3599), .dinb(n3481), .dout(n3600));
  jand g03409(.dina(n3600), .dinb(n3598), .dout(n3601));
  jxor g03410(.dina(n3601), .dinb(n3597), .dout(n3602));
  jxor g03411(.dina(n3602), .dinb(n3594), .dout(n3603));
  jand g03412(.dina(n3484), .dinb(n3480), .dout(n3604));
  jand g03413(.dina(n3485), .dinb(n3471), .dout(n3605));
  jor  g03414(.dina(n3605), .dinb(n3604), .dout(n3606));
  jxor g03415(.dina(n3606), .dinb(n3603), .dout(n3607));
  jand g03416(.dina(n3457), .dinb(n3454), .dout(n3608));
  jnot g03417(.din(n3608), .dout(n3609));
  jand g03418(.dina(n3609), .dinb(n3460), .dout(n3610));
  jor  g03419(.dina(n3514), .dinb(n3513), .dout(n3611));
  jand g03420(.dina(n3611), .dinb(n3518), .dout(n3612));
  jxor g03421(.dina(n3612), .dinb(n3610), .dout(n3613));
  jand g03422(.dina(n3449), .dinb(n3442), .dout(n3614));
  jor  g03423(.dina(n3614), .dinb(n3444), .dout(n3615));
  jxor g03424(.dina(n3615), .dinb(n3613), .dout(n3616));
  jxor g03425(.dina(n3616), .dinb(n3607), .dout(n3617));
  jxor g03426(.dina(n3617), .dinb(n3592), .dout(n3618));
  jand g03427(.dina(n3418), .dinb(n3392), .dout(n3619));
  jand g03428(.dina(n3419), .dinb(n3389), .dout(n3620));
  jor  g03429(.dina(n3620), .dinb(n3619), .dout(n3621));
  jand g03430(.dina(n3431), .dinb(n3427), .dout(n3622));
  jnot g03431(.din(n3622), .dout(n3623));
  jor  g03432(.dina(n3437), .dinb(n3433), .dout(n3624));
  jand g03433(.dina(n3624), .dinb(n3623), .dout(n3625));
  jnot g03434(.din(n3625), .dout(n3626));
  jand g03435(.dina(\a[36] ), .dinb(\a[6] ), .dout(n3627));
  jand g03436(.dina(\a[35] ), .dinb(\a[7] ), .dout(n3628));
  jand g03437(.dina(\a[31] ), .dinb(\a[11] ), .dout(n3629));
  jxor g03438(.dina(n3629), .dinb(n3628), .dout(n3630));
  jxor g03439(.dina(n3630), .dinb(n3627), .dout(n3631));
  jxor g03440(.dina(n3631), .dinb(n3502), .dout(n3632));
  jand g03441(.dina(\a[32] ), .dinb(\a[10] ), .dout(n3633));
  jand g03442(.dina(\a[34] ), .dinb(\a[33] ), .dout(n3634));
  jand g03443(.dina(n3634), .dinb(n395), .dout(n3635));
  jnot g03444(.din(n3635), .dout(n3636));
  jand g03445(.dina(\a[34] ), .dinb(\a[8] ), .dout(n3637));
  jand g03446(.dina(\a[33] ), .dinb(\a[9] ), .dout(n3638));
  jor  g03447(.dina(n3638), .dinb(n3637), .dout(n3639));
  jand g03448(.dina(n3639), .dinb(n3636), .dout(n3640));
  jxor g03449(.dina(n3640), .dinb(n3633), .dout(n3641));
  jxor g03450(.dina(n3641), .dinb(n3632), .dout(n3642));
  jxor g03451(.dina(n3642), .dinb(n3626), .dout(n3643));
  jand g03452(.dina(\a[27] ), .dinb(\a[15] ), .dout(n3644));
  jand g03453(.dina(\a[28] ), .dinb(\a[14] ), .dout(n3645));
  jand g03454(.dina(\a[38] ), .dinb(\a[4] ), .dout(n3646));
  jand g03455(.dina(n3646), .dinb(n3645), .dout(n3647));
  jnot g03456(.din(n3647), .dout(n3648));
  jand g03457(.dina(n2042), .dinb(n976), .dout(n3649));
  jand g03458(.dina(n3646), .dinb(n3644), .dout(n3650));
  jor  g03459(.dina(n3650), .dinb(n3649), .dout(n3651));
  jand g03460(.dina(n3651), .dinb(n3648), .dout(n3652));
  jnot g03461(.din(n3652), .dout(n3653));
  jand g03462(.dina(n3653), .dinb(n3644), .dout(n3654));
  jor  g03463(.dina(n3651), .dinb(n3647), .dout(n3655));
  jnot g03464(.din(n3655), .dout(n3656));
  jor  g03465(.dina(n3646), .dinb(n3645), .dout(n3657));
  jand g03466(.dina(n3657), .dinb(n3656), .dout(n3658));
  jor  g03467(.dina(n3658), .dinb(n3654), .dout(n3659));
  jand g03468(.dina(\a[39] ), .dinb(\a[3] ), .dout(n3660));
  jand g03469(.dina(\a[26] ), .dinb(\a[16] ), .dout(n3661));
  jand g03470(.dina(n3661), .dinb(n3660), .dout(n3662));
  jnot g03471(.din(n3662), .dout(n3663));
  jand g03472(.dina(n3661), .dinb(n3261), .dout(n3664));
  jand g03473(.dina(\a[40] ), .dinb(\a[39] ), .dout(n3665));
  jand g03474(.dina(n3665), .dinb(n248), .dout(n3666));
  jor  g03475(.dina(n3666), .dinb(n3664), .dout(n3667));
  jnot g03476(.din(n3667), .dout(n3668));
  jand g03477(.dina(n3668), .dinb(n3663), .dout(n3669));
  jor  g03478(.dina(n3661), .dinb(n3660), .dout(n3670));
  jand g03479(.dina(n3670), .dinb(n3669), .dout(n3671));
  jand g03480(.dina(n3667), .dinb(n3663), .dout(n3672));
  jnot g03481(.din(n3672), .dout(n3673));
  jand g03482(.dina(n3673), .dinb(n3261), .dout(n3674));
  jor  g03483(.dina(n3674), .dinb(n3671), .dout(n3675));
  jand g03484(.dina(\a[25] ), .dinb(\a[17] ), .dout(n3676));
  jnot g03485(.din(n3676), .dout(n3677));
  jand g03486(.dina(n1942), .dinb(n1024), .dout(n3678));
  jnot g03487(.din(n3678), .dout(n3679));
  jand g03488(.dina(\a[23] ), .dinb(\a[19] ), .dout(n3680));
  jand g03489(.dina(\a[24] ), .dinb(\a[18] ), .dout(n3681));
  jor  g03490(.dina(n3681), .dinb(n3680), .dout(n3682));
  jand g03491(.dina(n3682), .dinb(n3679), .dout(n3683));
  jxor g03492(.dina(n3683), .dinb(n3677), .dout(n3684));
  jnot g03493(.din(n3684), .dout(n3685));
  jxor g03494(.dina(n3685), .dinb(n3675), .dout(n3686));
  jxor g03495(.dina(n3686), .dinb(n3659), .dout(n3687));
  jxor g03496(.dina(n3687), .dinb(n3643), .dout(n3688));
  jxor g03497(.dina(n3688), .dinb(n3621), .dout(n3689));
  jxor g03498(.dina(n3689), .dinb(n3618), .dout(n3690));
  jxor g03499(.dina(n3690), .dinb(n3559), .dout(n3691));
  jand g03500(.dina(n3691), .dinb(n3534), .dout(n3692));
  jor  g03501(.dina(n3691), .dinb(n3534), .dout(n3693));
  jnot g03502(.din(n3693), .dout(n3694));
  jor  g03503(.dina(n3694), .dinb(n3692), .dout(n3695));
  jand g03504(.dina(n3526), .dinb(n3385), .dout(n3696));
  jnot g03505(.din(n3696), .dout(n3697));
  jnot g03506(.din(n3526), .dout(n3698));
  jand g03507(.dina(n3698), .dinb(n3386), .dout(n3699));
  jor  g03508(.dina(n3530), .dinb(n3699), .dout(n3700));
  jand g03509(.dina(n3700), .dinb(n3697), .dout(n3701));
  jxor g03510(.dina(n3701), .dinb(n3695), .dout(\asquared[43] ));
  jand g03511(.dina(n3558), .dinb(n3537), .dout(n3703));
  jand g03512(.dina(n3690), .dinb(n3559), .dout(n3704));
  jor  g03513(.dina(n3704), .dinb(n3703), .dout(n3705));
  jand g03514(.dina(n3556), .dinb(n3553), .dout(n3706));
  jand g03515(.dina(n3557), .dinb(n3540), .dout(n3707));
  jor  g03516(.dina(n3707), .dinb(n3706), .dout(n3708));
  jor  g03517(.dina(n3548), .dinb(n3544), .dout(n3709));
  jand g03518(.dina(n3552), .dinb(n3549), .dout(n3710));
  jnot g03519(.din(n3710), .dout(n3711));
  jand g03520(.dina(n3711), .dinb(n3709), .dout(n3712));
  jnot g03521(.din(n3712), .dout(n3713));
  jand g03522(.dina(\a[40] ), .dinb(\a[3] ), .dout(n3714));
  jand g03523(.dina(\a[43] ), .dinb(\a[0] ), .dout(n3715));
  jand g03524(.dina(n3715), .dinb(n3714), .dout(n3716));
  jnot g03525(.din(n3716), .dout(n3717));
  jand g03526(.dina(n3665), .dinb(n265), .dout(n3718));
  jand g03527(.dina(\a[39] ), .dinb(\a[4] ), .dout(n3719));
  jand g03528(.dina(n3719), .dinb(n3715), .dout(n3720));
  jor  g03529(.dina(n3720), .dinb(n3718), .dout(n3721));
  jnot g03530(.din(n3721), .dout(n3722));
  jand g03531(.dina(n3722), .dinb(n3717), .dout(n3723));
  jor  g03532(.dina(n3715), .dinb(n3714), .dout(n3724));
  jand g03533(.dina(n3724), .dinb(n3723), .dout(n3725));
  jand g03534(.dina(n3721), .dinb(n3717), .dout(n3726));
  jnot g03535(.din(n3726), .dout(n3727));
  jand g03536(.dina(n3727), .dinb(n3719), .dout(n3728));
  jor  g03537(.dina(n3728), .dinb(n3725), .dout(n3729));
  jand g03538(.dina(\a[29] ), .dinb(\a[14] ), .dout(n3730));
  jnot g03539(.din(n3730), .dout(n3731));
  jand g03540(.dina(n2042), .dinb(n829), .dout(n3732));
  jnot g03541(.din(n3732), .dout(n3733));
  jand g03542(.dina(\a[28] ), .dinb(\a[15] ), .dout(n3734));
  jand g03543(.dina(\a[27] ), .dinb(\a[16] ), .dout(n3735));
  jor  g03544(.dina(n3735), .dinb(n3734), .dout(n3736));
  jand g03545(.dina(n3736), .dinb(n3733), .dout(n3737));
  jxor g03546(.dina(n3737), .dinb(n3731), .dout(n3738));
  jnot g03547(.din(n3738), .dout(n3739));
  jxor g03548(.dina(n3739), .dinb(n3729), .dout(n3740));
  jnot g03549(.din(n3740), .dout(n3741));
  jand g03550(.dina(\a[26] ), .dinb(\a[17] ), .dout(n3742));
  jnot g03551(.din(n3742), .dout(n3743));
  jand g03552(.dina(n1648), .dinb(n1024), .dout(n3744));
  jnot g03553(.din(n3744), .dout(n3745));
  jand g03554(.dina(\a[24] ), .dinb(\a[19] ), .dout(n3746));
  jand g03555(.dina(\a[25] ), .dinb(\a[18] ), .dout(n3747));
  jor  g03556(.dina(n3747), .dinb(n3746), .dout(n3748));
  jand g03557(.dina(n3748), .dinb(n3745), .dout(n3749));
  jxor g03558(.dina(n3749), .dinb(n3743), .dout(n3750));
  jxor g03559(.dina(n3750), .dinb(n3741), .dout(n3751));
  jand g03560(.dina(\a[35] ), .dinb(\a[33] ), .dout(n3752));
  jand g03561(.dina(n3752), .dinb(n436), .dout(n3753));
  jnot g03562(.din(n3753), .dout(n3754));
  jand g03563(.dina(n3243), .dinb(n499), .dout(n3755));
  jand g03564(.dina(\a[33] ), .dinb(\a[10] ), .dout(n3756));
  jand g03565(.dina(\a[36] ), .dinb(\a[7] ), .dout(n3757));
  jand g03566(.dina(n3757), .dinb(n3756), .dout(n3758));
  jor  g03567(.dina(n3758), .dinb(n3755), .dout(n3759));
  jnot g03568(.din(n3759), .dout(n3760));
  jand g03569(.dina(n3760), .dinb(n3754), .dout(n3761));
  jand g03570(.dina(\a[35] ), .dinb(\a[8] ), .dout(n3762));
  jor  g03571(.dina(n3762), .dinb(n3756), .dout(n3763));
  jand g03572(.dina(n3763), .dinb(n3761), .dout(n3764));
  jand g03573(.dina(n3759), .dinb(n3754), .dout(n3765));
  jnot g03574(.din(n3765), .dout(n3766));
  jand g03575(.dina(n3766), .dinb(n3757), .dout(n3767));
  jor  g03576(.dina(n3767), .dinb(n3764), .dout(n3768));
  jand g03577(.dina(\a[34] ), .dinb(\a[9] ), .dout(n3769));
  jnot g03578(.din(n3769), .dout(n3770));
  jand g03579(.dina(n1658), .dinb(n1490), .dout(n3771));
  jnot g03580(.din(n3771), .dout(n3772));
  jand g03581(.dina(\a[23] ), .dinb(\a[20] ), .dout(n3773));
  jor  g03582(.dina(n3773), .dinb(n1376), .dout(n3774));
  jand g03583(.dina(n3774), .dinb(n3772), .dout(n3775));
  jxor g03584(.dina(n3775), .dinb(n3770), .dout(n3776));
  jnot g03585(.din(n3776), .dout(n3777));
  jxor g03586(.dina(n3777), .dinb(n3768), .dout(n3778));
  jand g03587(.dina(\a[38] ), .dinb(\a[5] ), .dout(n3779));
  jand g03588(.dina(\a[30] ), .dinb(\a[13] ), .dout(n3780));
  jxor g03589(.dina(n3780), .dinb(n3779), .dout(n3781));
  jxor g03590(.dina(n3781), .dinb(n3443), .dout(n3782));
  jxor g03591(.dina(n3782), .dinb(n3778), .dout(n3783));
  jxor g03592(.dina(n3783), .dinb(n3751), .dout(n3784));
  jxor g03593(.dina(n3784), .dinb(n3713), .dout(n3785));
  jxor g03594(.dina(n3785), .dinb(n3708), .dout(n3786));
  jand g03595(.dina(n3584), .dinb(n3578), .dout(n3787));
  jand g03596(.dina(n3585), .dinb(n3562), .dout(n3788));
  jor  g03597(.dina(n3788), .dinb(n3787), .dout(n3789));
  jand g03598(.dina(n3629), .dinb(n3628), .dout(n3790));
  jand g03599(.dina(n3630), .dinb(n3627), .dout(n3791));
  jor  g03600(.dina(n3791), .dinb(n3790), .dout(n3792));
  jxor g03601(.dina(n3792), .dinb(n3655), .dout(n3793));
  jand g03602(.dina(n3679), .dinb(n3677), .dout(n3794));
  jnot g03603(.din(n3794), .dout(n3795));
  jand g03604(.dina(n3795), .dinb(n3682), .dout(n3796));
  jxor g03605(.dina(n3796), .dinb(n3793), .dout(n3797));
  jxor g03606(.dina(n3669), .dinb(n3575), .dout(n3798));
  jand g03607(.dina(n3579), .dinb(n3408), .dout(n3799));
  jand g03608(.dina(n3583), .dinb(n3580), .dout(n3800));
  jor  g03609(.dina(n3800), .dinb(n3799), .dout(n3801));
  jxor g03610(.dina(n3801), .dinb(n3798), .dout(n3802));
  jxor g03611(.dina(n3802), .dinb(n3797), .dout(n3803));
  jxor g03612(.dina(n3803), .dinb(n3789), .dout(n3804));
  jand g03613(.dina(n3612), .dinb(n3610), .dout(n3805));
  jand g03614(.dina(n3615), .dinb(n3613), .dout(n3806));
  jor  g03615(.dina(n3806), .dinb(n3805), .dout(n3807));
  jand g03616(.dina(n3601), .dinb(n3597), .dout(n3808));
  jand g03617(.dina(n3602), .dinb(n3594), .dout(n3809));
  jor  g03618(.dina(n3809), .dinb(n3808), .dout(n3810));
  jand g03619(.dina(\a[31] ), .dinb(\a[12] ), .dout(n3811));
  jand g03620(.dina(n3269), .dinb(n555), .dout(n3812));
  jand g03621(.dina(\a[37] ), .dinb(\a[6] ), .dout(n3813));
  jand g03622(.dina(n3813), .dinb(n3811), .dout(n3814));
  jor  g03623(.dina(n3814), .dinb(n3812), .dout(n3815));
  jand g03624(.dina(\a[32] ), .dinb(\a[11] ), .dout(n3816));
  jand g03625(.dina(n3816), .dinb(n3813), .dout(n3817));
  jnot g03626(.din(n3817), .dout(n3818));
  jand g03627(.dina(n3818), .dinb(n3815), .dout(n3819));
  jnot g03628(.din(n3819), .dout(n3820));
  jand g03629(.dina(n3820), .dinb(n3811), .dout(n3821));
  jor  g03630(.dina(n3817), .dinb(n3815), .dout(n3822));
  jnot g03631(.din(n3822), .dout(n3823));
  jor  g03632(.dina(n3816), .dinb(n3813), .dout(n3824));
  jand g03633(.dina(n3824), .dinb(n3823), .dout(n3825));
  jor  g03634(.dina(n3825), .dinb(n3821), .dout(n3826));
  jxor g03635(.dina(n3826), .dinb(n3810), .dout(n3827));
  jxor g03636(.dina(n3827), .dinb(n3807), .dout(n3828));
  jand g03637(.dina(n3606), .dinb(n3603), .dout(n3829));
  jand g03638(.dina(n3616), .dinb(n3607), .dout(n3830));
  jor  g03639(.dina(n3830), .dinb(n3829), .dout(n3831));
  jxor g03640(.dina(n3831), .dinb(n3828), .dout(n3832));
  jxor g03641(.dina(n3832), .dinb(n3804), .dout(n3833));
  jxor g03642(.dina(n3833), .dinb(n3786), .dout(n3834));
  jand g03643(.dina(n3688), .dinb(n3621), .dout(n3835));
  jand g03644(.dina(n3689), .dinb(n3618), .dout(n3836));
  jor  g03645(.dina(n3836), .dinb(n3835), .dout(n3837));
  jor  g03646(.dina(n3591), .dinb(n3587), .dout(n3838));
  jand g03647(.dina(n3617), .dinb(n3592), .dout(n3839));
  jnot g03648(.din(n3839), .dout(n3840));
  jand g03649(.dina(n3840), .dinb(n3838), .dout(n3841));
  jnot g03650(.din(n3841), .dout(n3842));
  jand g03651(.dina(n3642), .dinb(n3626), .dout(n3843));
  jand g03652(.dina(n3687), .dinb(n3643), .dout(n3844));
  jor  g03653(.dina(n3844), .dinb(n3843), .dout(n3845));
  jand g03654(.dina(n3685), .dinb(n3675), .dout(n3846));
  jand g03655(.dina(n3686), .dinb(n3659), .dout(n3847));
  jor  g03656(.dina(n3847), .dinb(n3846), .dout(n3848));
  jand g03657(.dina(n3631), .dinb(n3502), .dout(n3849));
  jand g03658(.dina(n3641), .dinb(n3632), .dout(n3850));
  jor  g03659(.dina(n3850), .dinb(n3849), .dout(n3851));
  jand g03660(.dina(n3639), .dinb(n3633), .dout(n3852));
  jor  g03661(.dina(n3852), .dinb(n3635), .dout(n3853));
  jand g03662(.dina(\a[42] ), .dinb(\a[1] ), .dout(n3854));
  jnot g03663(.din(\a[22] ), .dout(n3855));
  jand g03664(.dina(n3582), .dinb(n3581), .dout(n3856));
  jor  g03665(.dina(n3856), .dinb(n3855), .dout(n3857));
  jxor g03666(.dina(n3857), .dinb(n3854), .dout(n3858));
  jnot g03667(.din(n3858), .dout(n3859));
  jxor g03668(.dina(n3859), .dinb(n3853), .dout(n3860));
  jxor g03669(.dina(n3860), .dinb(n3851), .dout(n3861));
  jxor g03670(.dina(n3861), .dinb(n3848), .dout(n3862));
  jxor g03671(.dina(n3862), .dinb(n3845), .dout(n3863));
  jxor g03672(.dina(n3863), .dinb(n3842), .dout(n3864));
  jxor g03673(.dina(n3864), .dinb(n3837), .dout(n3865));
  jxor g03674(.dina(n3865), .dinb(n3834), .dout(n3866));
  jand g03675(.dina(n3866), .dinb(n3705), .dout(n3867));
  jor  g03676(.dina(n3866), .dinb(n3705), .dout(n3868));
  jnot g03677(.din(n3868), .dout(n3869));
  jor  g03678(.dina(n3869), .dinb(n3867), .dout(n3870));
  jnot g03679(.din(n3692), .dout(n3871));
  jor  g03680(.dina(n3701), .dinb(n3694), .dout(n3872));
  jand g03681(.dina(n3872), .dinb(n3871), .dout(n3873));
  jxor g03682(.dina(n3873), .dinb(n3870), .dout(\asquared[44] ));
  jand g03683(.dina(n3864), .dinb(n3837), .dout(n3875));
  jand g03684(.dina(n3865), .dinb(n3834), .dout(n3876));
  jor  g03685(.dina(n3876), .dinb(n3875), .dout(n3877));
  jand g03686(.dina(n3785), .dinb(n3708), .dout(n3878));
  jand g03687(.dina(n3833), .dinb(n3786), .dout(n3879));
  jor  g03688(.dina(n3879), .dinb(n3878), .dout(n3880));
  jand g03689(.dina(n3831), .dinb(n3828), .dout(n3881));
  jand g03690(.dina(n3832), .dinb(n3804), .dout(n3882));
  jor  g03691(.dina(n3882), .dinb(n3881), .dout(n3883));
  jand g03692(.dina(n3783), .dinb(n3751), .dout(n3884));
  jand g03693(.dina(n3784), .dinb(n3713), .dout(n3885));
  jor  g03694(.dina(n3885), .dinb(n3884), .dout(n3886));
  jnot g03695(.din(n3723), .dout(n3887));
  jand g03696(.dina(n3780), .dinb(n3779), .dout(n3888));
  jand g03697(.dina(n3781), .dinb(n3443), .dout(n3889));
  jor  g03698(.dina(n3889), .dinb(n3888), .dout(n3890));
  jxor g03699(.dina(n3890), .dinb(n3887), .dout(n3891));
  jand g03700(.dina(n3745), .dinb(n3743), .dout(n3892));
  jnot g03701(.din(n3892), .dout(n3893));
  jand g03702(.dina(n3893), .dinb(n3748), .dout(n3894));
  jxor g03703(.dina(n3894), .dinb(n3891), .dout(n3895));
  jand g03704(.dina(n3777), .dinb(n3768), .dout(n3896));
  jand g03705(.dina(n3782), .dinb(n3778), .dout(n3897));
  jor  g03706(.dina(n3897), .dinb(n3896), .dout(n3898));
  jnot g03707(.din(n3898), .dout(n3899));
  jand g03708(.dina(n3739), .dinb(n3729), .dout(n3900));
  jnot g03709(.din(n3900), .dout(n3901));
  jor  g03710(.dina(n3750), .dinb(n3741), .dout(n3902));
  jand g03711(.dina(n3902), .dinb(n3901), .dout(n3903));
  jxor g03712(.dina(n3903), .dinb(n3899), .dout(n3904));
  jxor g03713(.dina(n3904), .dinb(n3895), .dout(n3905));
  jxor g03714(.dina(n3905), .dinb(n3886), .dout(n3906));
  jxor g03715(.dina(n3906), .dinb(n3883), .dout(n3907));
  jxor g03716(.dina(n3907), .dinb(n3880), .dout(n3908));
  jand g03717(.dina(n3862), .dinb(n3845), .dout(n3909));
  jand g03718(.dina(n3863), .dinb(n3842), .dout(n3910));
  jor  g03719(.dina(n3910), .dinb(n3909), .dout(n3911));
  jand g03720(.dina(n3860), .dinb(n3851), .dout(n3912));
  jand g03721(.dina(n3861), .dinb(n3848), .dout(n3913));
  jor  g03722(.dina(n3913), .dinb(n3912), .dout(n3914));
  jand g03723(.dina(\a[30] ), .dinb(\a[14] ), .dout(n3915));
  jand g03724(.dina(\a[40] ), .dinb(\a[4] ), .dout(n3916));
  jand g03725(.dina(n3916), .dinb(n3915), .dout(n3917));
  jnot g03726(.din(n3917), .dout(n3918));
  jand g03727(.dina(\a[28] ), .dinb(\a[16] ), .dout(n3919));
  jand g03728(.dina(n3919), .dinb(n3916), .dout(n3920));
  jand g03729(.dina(n2810), .dinb(n1874), .dout(n3921));
  jor  g03730(.dina(n3921), .dinb(n3920), .dout(n3922));
  jnot g03731(.din(n3922), .dout(n3923));
  jand g03732(.dina(n3923), .dinb(n3918), .dout(n3924));
  jor  g03733(.dina(n3916), .dinb(n3915), .dout(n3925));
  jand g03734(.dina(n3925), .dinb(n3924), .dout(n3926));
  jand g03735(.dina(n3922), .dinb(n3918), .dout(n3927));
  jnot g03736(.din(n3927), .dout(n3928));
  jand g03737(.dina(n3928), .dinb(n3919), .dout(n3929));
  jor  g03738(.dina(n3929), .dinb(n3926), .dout(n3930));
  jand g03739(.dina(\a[36] ), .dinb(\a[8] ), .dout(n3931));
  jnot g03740(.din(n3931), .dout(n3932));
  jand g03741(.dina(n2845), .dinb(n453), .dout(n3933));
  jnot g03742(.din(n3933), .dout(n3934));
  jand g03743(.dina(\a[34] ), .dinb(\a[10] ), .dout(n3935));
  jand g03744(.dina(\a[35] ), .dinb(\a[9] ), .dout(n3936));
  jor  g03745(.dina(n3936), .dinb(n3935), .dout(n3937));
  jand g03746(.dina(n3937), .dinb(n3934), .dout(n3938));
  jxor g03747(.dina(n3938), .dinb(n3932), .dout(n3939));
  jnot g03748(.din(n3939), .dout(n3940));
  jxor g03749(.dina(n3940), .dinb(n3930), .dout(n3941));
  jnot g03750(.din(n3941), .dout(n3942));
  jand g03751(.dina(\a[39] ), .dinb(\a[5] ), .dout(n3943));
  jnot g03752(.din(n3943), .dout(n3944));
  jand g03753(.dina(n3269), .dinb(n899), .dout(n3945));
  jnot g03754(.din(n3945), .dout(n3946));
  jand g03755(.dina(\a[32] ), .dinb(\a[12] ), .dout(n3947));
  jand g03756(.dina(\a[31] ), .dinb(\a[13] ), .dout(n3948));
  jor  g03757(.dina(n3948), .dinb(n3947), .dout(n3949));
  jand g03758(.dina(n3949), .dinb(n3946), .dout(n3950));
  jxor g03759(.dina(n3950), .dinb(n3944), .dout(n3951));
  jxor g03760(.dina(n3951), .dinb(n3942), .dout(n3952));
  jand g03761(.dina(\a[41] ), .dinb(\a[3] ), .dout(n3953));
  jand g03762(.dina(\a[29] ), .dinb(\a[15] ), .dout(n3954));
  jand g03763(.dina(\a[27] ), .dinb(\a[17] ), .dout(n3955));
  jor  g03764(.dina(n3955), .dinb(n3954), .dout(n3956));
  jand g03765(.dina(n2536), .dinb(n878), .dout(n3957));
  jnot g03766(.din(n3957), .dout(n3958));
  jand g03767(.dina(n3958), .dinb(n3956), .dout(n3959));
  jxor g03768(.dina(n3959), .dinb(n3953), .dout(n3960));
  jnot g03769(.din(n3960), .dout(n3961));
  jand g03770(.dina(\a[26] ), .dinb(\a[18] ), .dout(n3962));
  jnot g03771(.din(n3962), .dout(n3963));
  jand g03772(.dina(n1648), .dinb(n1287), .dout(n3964));
  jnot g03773(.din(n3964), .dout(n3965));
  jand g03774(.dina(\a[25] ), .dinb(\a[19] ), .dout(n3966));
  jand g03775(.dina(\a[24] ), .dinb(\a[20] ), .dout(n3967));
  jor  g03776(.dina(n3967), .dinb(n3966), .dout(n3968));
  jand g03777(.dina(n3968), .dinb(n3965), .dout(n3969));
  jxor g03778(.dina(n3969), .dinb(n3963), .dout(n3970));
  jxor g03779(.dina(n3970), .dinb(n3961), .dout(n3971));
  jnot g03780(.din(n3971), .dout(n3972));
  jand g03781(.dina(\a[38] ), .dinb(\a[6] ), .dout(n3973));
  jnot g03782(.din(n3973), .dout(n3974));
  jand g03783(.dina(\a[37] ), .dinb(\a[7] ), .dout(n3975));
  jand g03784(.dina(\a[33] ), .dinb(\a[11] ), .dout(n3976));
  jxor g03785(.dina(n3976), .dinb(n3975), .dout(n3977));
  jxor g03786(.dina(n3977), .dinb(n3974), .dout(n3978));
  jxor g03787(.dina(n3978), .dinb(n3972), .dout(n3979));
  jxor g03788(.dina(n3979), .dinb(n3952), .dout(n3980));
  jxor g03789(.dina(n3980), .dinb(n3914), .dout(n3981));
  jxor g03790(.dina(n3981), .dinb(n3911), .dout(n3982));
  jand g03791(.dina(n3826), .dinb(n3810), .dout(n3983));
  jand g03792(.dina(n3827), .dinb(n3807), .dout(n3984));
  jor  g03793(.dina(n3984), .dinb(n3983), .dout(n3985));
  jnot g03794(.din(n3761), .dout(n3986));
  jand g03795(.dina(\a[23] ), .dinb(\a[21] ), .dout(n3987));
  jand g03796(.dina(\a[43] ), .dinb(\a[1] ), .dout(n3988));
  jxor g03797(.dina(n3988), .dinb(n3987), .dout(n3989));
  jand g03798(.dina(n3772), .dinb(n3770), .dout(n3990));
  jnot g03799(.din(n3990), .dout(n3991));
  jand g03800(.dina(n3991), .dinb(n3774), .dout(n3992));
  jxor g03801(.dina(n3992), .dinb(n3989), .dout(n3993));
  jxor g03802(.dina(n3993), .dinb(n3986), .dout(n3994));
  jand g03803(.dina(n3733), .dinb(n3731), .dout(n3995));
  jnot g03804(.din(n3995), .dout(n3996));
  jand g03805(.dina(n3996), .dinb(n3736), .dout(n3997));
  jxor g03806(.dina(n3997), .dinb(n3822), .dout(n3998));
  jand g03807(.dina(n1238), .dinb(\a[42] ), .dout(n3999));
  jand g03808(.dina(\a[44] ), .dinb(\a[2] ), .dout(n4000));
  jand g03809(.dina(n4000), .dinb(n3579), .dout(n4001));
  jnot g03810(.din(n4001), .dout(n4002));
  jand g03811(.dina(\a[44] ), .dinb(\a[0] ), .dout(n4003));
  jand g03812(.dina(\a[42] ), .dinb(\a[2] ), .dout(n4004));
  jor  g03813(.dina(n4004), .dinb(n4003), .dout(n4005));
  jand g03814(.dina(n4005), .dinb(n4002), .dout(n4006));
  jxor g03815(.dina(n4006), .dinb(n3999), .dout(n4007));
  jxor g03816(.dina(n4007), .dinb(n3998), .dout(n4008));
  jxor g03817(.dina(n4008), .dinb(n3994), .dout(n4009));
  jxor g03818(.dina(n4009), .dinb(n3985), .dout(n4010));
  jand g03819(.dina(n3802), .dinb(n3797), .dout(n4011));
  jand g03820(.dina(n3803), .dinb(n3789), .dout(n4012));
  jor  g03821(.dina(n4012), .dinb(n4011), .dout(n4013));
  jnot g03822(.din(n3669), .dout(n4014));
  jand g03823(.dina(n4014), .dinb(n3574), .dout(n4015));
  jand g03824(.dina(n3801), .dinb(n3798), .dout(n4016));
  jor  g03825(.dina(n4016), .dinb(n4015), .dout(n4017));
  jand g03826(.dina(n3859), .dinb(n3853), .dout(n4018));
  jnot g03827(.din(\a[42] ), .dout(n4019));
  jand g03828(.dina(n3856), .dinb(n4019), .dout(n4020));
  jor  g03829(.dina(n4020), .dinb(n4018), .dout(n4021));
  jxor g03830(.dina(n4021), .dinb(n4017), .dout(n4022));
  jand g03831(.dina(n3792), .dinb(n3655), .dout(n4023));
  jand g03832(.dina(n3796), .dinb(n3793), .dout(n4024));
  jor  g03833(.dina(n4024), .dinb(n4023), .dout(n4025));
  jxor g03834(.dina(n4025), .dinb(n4022), .dout(n4026));
  jxor g03835(.dina(n4026), .dinb(n4013), .dout(n4027));
  jxor g03836(.dina(n4027), .dinb(n4010), .dout(n4028));
  jxor g03837(.dina(n4028), .dinb(n3982), .dout(n4029));
  jxor g03838(.dina(n4029), .dinb(n3908), .dout(n4030));
  jand g03839(.dina(n4030), .dinb(n3877), .dout(n4031));
  jor  g03840(.dina(n4030), .dinb(n3877), .dout(n4032));
  jnot g03841(.din(n4032), .dout(n4033));
  jor  g03842(.dina(n4033), .dinb(n4031), .dout(n4034));
  jnot g03843(.din(n3867), .dout(n4035));
  jor  g03844(.dina(n3873), .dinb(n3869), .dout(n4036));
  jand g03845(.dina(n4036), .dinb(n4035), .dout(n4037));
  jxor g03846(.dina(n4037), .dinb(n4034), .dout(\asquared[45] ));
  jand g03847(.dina(n3907), .dinb(n3880), .dout(n4039));
  jand g03848(.dina(n4029), .dinb(n3908), .dout(n4040));
  jor  g03849(.dina(n4040), .dinb(n4039), .dout(n4041));
  jand g03850(.dina(n3981), .dinb(n3911), .dout(n4042));
  jand g03851(.dina(n4028), .dinb(n3982), .dout(n4043));
  jor  g03852(.dina(n4043), .dinb(n4042), .dout(n4044));
  jand g03853(.dina(n3979), .dinb(n3952), .dout(n4045));
  jand g03854(.dina(n3980), .dinb(n3914), .dout(n4046));
  jor  g03855(.dina(n4046), .dinb(n4045), .dout(n4047));
  jand g03856(.dina(n4026), .dinb(n4013), .dout(n4048));
  jand g03857(.dina(n4027), .dinb(n4010), .dout(n4049));
  jor  g03858(.dina(n4049), .dinb(n4048), .dout(n4050));
  jxor g03859(.dina(n4050), .dinb(n4047), .dout(n4051));
  jand g03860(.dina(n3959), .dinb(n3953), .dout(n4052));
  jor  g03861(.dina(n4052), .dinb(n3957), .dout(n4053));
  jand g03862(.dina(n4006), .dinb(n3999), .dout(n4054));
  jor  g03863(.dina(n4054), .dinb(n4001), .dout(n4055));
  jxor g03864(.dina(n4055), .dinb(n4053), .dout(n4056));
  jand g03865(.dina(n3965), .dinb(n3963), .dout(n4057));
  jnot g03866(.din(n4057), .dout(n4058));
  jand g03867(.dina(n4058), .dinb(n3968), .dout(n4059));
  jxor g03868(.dina(n4059), .dinb(n4056), .dout(n4060));
  jand g03869(.dina(n4021), .dinb(n4017), .dout(n4061));
  jand g03870(.dina(n4025), .dinb(n4022), .dout(n4062));
  jor  g03871(.dina(n4062), .dinb(n4061), .dout(n4063));
  jxor g03872(.dina(n4063), .dinb(n4060), .dout(n4064));
  jand g03873(.dina(\a[34] ), .dinb(\a[11] ), .dout(n4065));
  jand g03874(.dina(\a[39] ), .dinb(\a[6] ), .dout(n4066));
  jor  g03875(.dina(n4066), .dinb(n4065), .dout(n4067));
  jand g03876(.dina(\a[39] ), .dinb(\a[34] ), .dout(n4068));
  jand g03877(.dina(n4068), .dinb(n725), .dout(n4069));
  jnot g03878(.din(n4069), .dout(n4070));
  jand g03879(.dina(\a[33] ), .dinb(\a[12] ), .dout(n4071));
  jand g03880(.dina(n4071), .dinb(n4066), .dout(n4072));
  jand g03881(.dina(n3634), .dinb(n555), .dout(n4073));
  jor  g03882(.dina(n4073), .dinb(n4072), .dout(n4074));
  jnot g03883(.din(n4074), .dout(n4075));
  jand g03884(.dina(n4075), .dinb(n4070), .dout(n4076));
  jand g03885(.dina(n4076), .dinb(n4067), .dout(n4077));
  jand g03886(.dina(n4074), .dinb(n4070), .dout(n4078));
  jnot g03887(.din(n4078), .dout(n4079));
  jand g03888(.dina(n4079), .dinb(n4071), .dout(n4080));
  jor  g03889(.dina(n4080), .dinb(n4077), .dout(n4081));
  jand g03890(.dina(\a[30] ), .dinb(\a[15] ), .dout(n4082));
  jnot g03891(.din(n4082), .dout(n4083));
  jand g03892(.dina(n2653), .dinb(n937), .dout(n4084));
  jnot g03893(.din(n4084), .dout(n4085));
  jand g03894(.dina(\a[28] ), .dinb(\a[17] ), .dout(n4086));
  jand g03895(.dina(\a[29] ), .dinb(\a[16] ), .dout(n4087));
  jor  g03896(.dina(n4087), .dinb(n4086), .dout(n4088));
  jand g03897(.dina(n4088), .dinb(n4085), .dout(n4089));
  jxor g03898(.dina(n4089), .dinb(n4083), .dout(n4090));
  jnot g03899(.din(n4090), .dout(n4091));
  jxor g03900(.dina(n4091), .dinb(n4081), .dout(n4092));
  jand g03901(.dina(n1277), .dinb(\a[44] ), .dout(n4093));
  jnot g03902(.din(n4093), .dout(n4094));
  jand g03903(.dina(\a[44] ), .dinb(\a[1] ), .dout(n4095));
  jor  g03904(.dina(n4095), .dinb(\a[23] ), .dout(n4096));
  jand g03905(.dina(n4096), .dinb(n4094), .dout(n4097));
  jand g03906(.dina(n3988), .dinb(n3987), .dout(n4098));
  jand g03907(.dina(\a[42] ), .dinb(\a[3] ), .dout(n4099));
  jxor g03908(.dina(n4099), .dinb(n4098), .dout(n4100));
  jxor g03909(.dina(n4100), .dinb(n4097), .dout(n4101));
  jxor g03910(.dina(n4101), .dinb(n4092), .dout(n4102));
  jxor g03911(.dina(n4102), .dinb(n4064), .dout(n4103));
  jxor g03912(.dina(n4103), .dinb(n4051), .dout(n4104));
  jxor g03913(.dina(n4104), .dinb(n4044), .dout(n4105));
  jand g03914(.dina(n3905), .dinb(n3886), .dout(n4106));
  jand g03915(.dina(n3906), .dinb(n3883), .dout(n4107));
  jor  g03916(.dina(n4107), .dinb(n4106), .dout(n4108));
  jor  g03917(.dina(n3903), .dinb(n3899), .dout(n4109));
  jand g03918(.dina(n3904), .dinb(n3895), .dout(n4110));
  jnot g03919(.din(n4110), .dout(n4111));
  jand g03920(.dina(n4111), .dinb(n4109), .dout(n4112));
  jnot g03921(.din(n4112), .dout(n4113));
  jand g03922(.dina(\a[45] ), .dinb(\a[0] ), .dout(n4114));
  jand g03923(.dina(\a[43] ), .dinb(\a[41] ), .dout(n4115));
  jand g03924(.dina(n4115), .dinb(n245), .dout(n4116));
  jnot g03925(.din(n4116), .dout(n4117));
  jand g03926(.dina(\a[43] ), .dinb(\a[2] ), .dout(n4118));
  jand g03927(.dina(\a[41] ), .dinb(\a[4] ), .dout(n4119));
  jor  g03928(.dina(n4119), .dinb(n4118), .dout(n4120));
  jand g03929(.dina(n4120), .dinb(n4117), .dout(n4121));
  jxor g03930(.dina(n4121), .dinb(n4114), .dout(n4122));
  jnot g03931(.din(n4122), .dout(n4123));
  jand g03932(.dina(\a[38] ), .dinb(\a[7] ), .dout(n4124));
  jnot g03933(.din(n4124), .dout(n4125));
  jand g03934(.dina(n3138), .dinb(n395), .dout(n4126));
  jnot g03935(.din(n4126), .dout(n4127));
  jand g03936(.dina(\a[37] ), .dinb(\a[8] ), .dout(n4128));
  jand g03937(.dina(\a[36] ), .dinb(\a[9] ), .dout(n4129));
  jor  g03938(.dina(n4129), .dinb(n4128), .dout(n4130));
  jand g03939(.dina(n4130), .dinb(n4127), .dout(n4131));
  jxor g03940(.dina(n4131), .dinb(n4125), .dout(n4132));
  jxor g03941(.dina(n4132), .dinb(n4123), .dout(n4133));
  jnot g03942(.din(n4133), .dout(n4134));
  jand g03943(.dina(\a[35] ), .dinb(\a[10] ), .dout(n4135));
  jnot g03944(.din(n4135), .dout(n4136));
  jand g03945(.dina(n1942), .dinb(n1376), .dout(n4137));
  jnot g03946(.din(n4137), .dout(n4138));
  jand g03947(.dina(\a[24] ), .dinb(\a[21] ), .dout(n4139));
  jor  g03948(.dina(n4139), .dinb(n1658), .dout(n4140));
  jand g03949(.dina(n4140), .dinb(n4138), .dout(n4141));
  jxor g03950(.dina(n4141), .dinb(n4136), .dout(n4142));
  jxor g03951(.dina(n4142), .dinb(n4134), .dout(n4143));
  jand g03952(.dina(\a[32] ), .dinb(\a[13] ), .dout(n4144));
  jand g03953(.dina(\a[40] ), .dinb(\a[5] ), .dout(n4145));
  jand g03954(.dina(n4145), .dinb(n4144), .dout(n4146));
  jnot g03955(.din(n4146), .dout(n4147));
  jand g03956(.dina(n3269), .dinb(n675), .dout(n4148));
  jand g03957(.dina(\a[31] ), .dinb(\a[14] ), .dout(n4149));
  jand g03958(.dina(n4149), .dinb(n4145), .dout(n4150));
  jor  g03959(.dina(n4150), .dinb(n4148), .dout(n4151));
  jnot g03960(.din(n4151), .dout(n4152));
  jand g03961(.dina(n4152), .dinb(n4147), .dout(n4153));
  jor  g03962(.dina(n4145), .dinb(n4144), .dout(n4154));
  jand g03963(.dina(n4154), .dinb(n4153), .dout(n4155));
  jand g03964(.dina(n4151), .dinb(n4147), .dout(n4156));
  jnot g03965(.din(n4156), .dout(n4157));
  jand g03966(.dina(n4157), .dinb(n4149), .dout(n4158));
  jor  g03967(.dina(n4158), .dinb(n4155), .dout(n4159));
  jand g03968(.dina(n3934), .dinb(n3932), .dout(n4160));
  jnot g03969(.din(n4160), .dout(n4161));
  jand g03970(.dina(n4161), .dinb(n3937), .dout(n4162));
  jand g03971(.dina(\a[27] ), .dinb(\a[18] ), .dout(n4163));
  jand g03972(.dina(n2128), .dinb(n1287), .dout(n4164));
  jnot g03973(.din(n4164), .dout(n4165));
  jand g03974(.dina(\a[26] ), .dinb(\a[19] ), .dout(n4166));
  jor  g03975(.dina(n4166), .dinb(n1581), .dout(n4167));
  jand g03976(.dina(n4167), .dinb(n4165), .dout(n4168));
  jxor g03977(.dina(n4168), .dinb(n4163), .dout(n4169));
  jxor g03978(.dina(n4169), .dinb(n4162), .dout(n4170));
  jxor g03979(.dina(n4170), .dinb(n4159), .dout(n4171));
  jxor g03980(.dina(n4171), .dinb(n4143), .dout(n4172));
  jxor g03981(.dina(n4172), .dinb(n4113), .dout(n4173));
  jxor g03982(.dina(n4173), .dinb(n4108), .dout(n4174));
  jand g03983(.dina(n3997), .dinb(n3822), .dout(n4175));
  jand g03984(.dina(n4007), .dinb(n3998), .dout(n4176));
  jor  g03985(.dina(n4176), .dinb(n4175), .dout(n4177));
  jand g03986(.dina(n3890), .dinb(n3887), .dout(n4178));
  jand g03987(.dina(n3894), .dinb(n3891), .dout(n4179));
  jor  g03988(.dina(n4179), .dinb(n4178), .dout(n4180));
  jxor g03989(.dina(n4180), .dinb(n4177), .dout(n4181));
  jand g03990(.dina(n3992), .dinb(n3989), .dout(n4182));
  jand g03991(.dina(n3993), .dinb(n3986), .dout(n4183));
  jor  g03992(.dina(n4183), .dinb(n4182), .dout(n4184));
  jxor g03993(.dina(n4184), .dinb(n4181), .dout(n4185));
  jand g03994(.dina(n4008), .dinb(n3994), .dout(n4186));
  jand g03995(.dina(n4009), .dinb(n3985), .dout(n4187));
  jor  g03996(.dina(n4187), .dinb(n4186), .dout(n4188));
  jxor g03997(.dina(n4188), .dinb(n4185), .dout(n4189));
  jnot g03998(.din(n3924), .dout(n4190));
  jor  g03999(.dina(n3976), .dinb(n3975), .dout(n4191));
  jand g04000(.dina(n3976), .dinb(n3975), .dout(n4192));
  jor  g04001(.dina(n4192), .dinb(n3973), .dout(n4193));
  jand g04002(.dina(n4193), .dinb(n4191), .dout(n4194));
  jxor g04003(.dina(n4194), .dinb(n4190), .dout(n4195));
  jand g04004(.dina(n3946), .dinb(n3944), .dout(n4196));
  jnot g04005(.din(n4196), .dout(n4197));
  jand g04006(.dina(n4197), .dinb(n3949), .dout(n4198));
  jxor g04007(.dina(n4198), .dinb(n4195), .dout(n4199));
  jand g04008(.dina(n3940), .dinb(n3930), .dout(n4200));
  jnot g04009(.din(n4200), .dout(n4201));
  jor  g04010(.dina(n3951), .dinb(n3942), .dout(n4202));
  jand g04011(.dina(n4202), .dinb(n4201), .dout(n4203));
  jor  g04012(.dina(n3970), .dinb(n3961), .dout(n4204));
  jor  g04013(.dina(n3978), .dinb(n3972), .dout(n4205));
  jand g04014(.dina(n4205), .dinb(n4204), .dout(n4206));
  jxor g04015(.dina(n4206), .dinb(n4203), .dout(n4207));
  jxor g04016(.dina(n4207), .dinb(n4199), .dout(n4208));
  jxor g04017(.dina(n4208), .dinb(n4189), .dout(n4209));
  jxor g04018(.dina(n4209), .dinb(n4174), .dout(n4210));
  jxor g04019(.dina(n4210), .dinb(n4105), .dout(n4211));
  jand g04020(.dina(n4211), .dinb(n4041), .dout(n4212));
  jor  g04021(.dina(n4211), .dinb(n4041), .dout(n4213));
  jnot g04022(.din(n4213), .dout(n4214));
  jor  g04023(.dina(n4214), .dinb(n4212), .dout(n4215));
  jnot g04024(.din(n4031), .dout(n4216));
  jor  g04025(.dina(n4037), .dinb(n4033), .dout(n4217));
  jand g04026(.dina(n4217), .dinb(n4216), .dout(n4218));
  jxor g04027(.dina(n4218), .dinb(n4215), .dout(\asquared[46] ));
  jand g04028(.dina(n4104), .dinb(n4044), .dout(n4220));
  jand g04029(.dina(n4210), .dinb(n4105), .dout(n4221));
  jor  g04030(.dina(n4221), .dinb(n4220), .dout(n4222));
  jand g04031(.dina(n4173), .dinb(n4108), .dout(n4223));
  jand g04032(.dina(n4209), .dinb(n4174), .dout(n4224));
  jor  g04033(.dina(n4224), .dinb(n4223), .dout(n4225));
  jand g04034(.dina(n4188), .dinb(n4185), .dout(n4226));
  jand g04035(.dina(n4208), .dinb(n4189), .dout(n4227));
  jor  g04036(.dina(n4227), .dinb(n4226), .dout(n4228));
  jand g04037(.dina(n4171), .dinb(n4143), .dout(n4229));
  jand g04038(.dina(n4172), .dinb(n4113), .dout(n4230));
  jor  g04039(.dina(n4230), .dinb(n4229), .dout(n4231));
  jxor g04040(.dina(n4231), .dinb(n4228), .dout(n4232));
  jand g04041(.dina(n4194), .dinb(n4190), .dout(n4233));
  jand g04042(.dina(n4198), .dinb(n4195), .dout(n4234));
  jor  g04043(.dina(n4234), .dinb(n4233), .dout(n4235));
  jand g04044(.dina(\a[41] ), .dinb(\a[5] ), .dout(n4236));
  jand g04045(.dina(\a[31] ), .dinb(\a[15] ), .dout(n4237));
  jor  g04046(.dina(n4237), .dinb(n4236), .dout(n4238));
  jand g04047(.dina(\a[41] ), .dinb(\a[31] ), .dout(n4239));
  jand g04048(.dina(n4239), .dinb(n981), .dout(n4240));
  jnot g04049(.din(n4240), .dout(n4241));
  jand g04050(.dina(n4241), .dinb(n4238), .dout(n4242));
  jxor g04051(.dina(n4242), .dinb(n4000), .dout(n4243));
  jand g04052(.dina(n2671), .dinb(n675), .dout(n4244));
  jand g04053(.dina(\a[32] ), .dinb(\a[14] ), .dout(n4245));
  jand g04054(.dina(\a[40] ), .dinb(\a[6] ), .dout(n4246));
  jand g04055(.dina(n4246), .dinb(n4245), .dout(n4247));
  jor  g04056(.dina(n4247), .dinb(n4244), .dout(n4248));
  jand g04057(.dina(\a[33] ), .dinb(\a[13] ), .dout(n4249));
  jand g04058(.dina(n4249), .dinb(n4246), .dout(n4250));
  jnot g04059(.din(n4250), .dout(n4251));
  jand g04060(.dina(n4251), .dinb(n4248), .dout(n4252));
  jnot g04061(.din(n4252), .dout(n4253));
  jxor g04062(.dina(n4249), .dinb(n4246), .dout(n4254));
  jor  g04063(.dina(n4254), .dinb(n4245), .dout(n4255));
  jand g04064(.dina(n4255), .dinb(n4253), .dout(n4256));
  jxor g04065(.dina(n4256), .dinb(n4243), .dout(n4257));
  jxor g04066(.dina(n4257), .dinb(n4235), .dout(n4258));
  jnot g04067(.din(n4076), .dout(n4259));
  jand g04068(.dina(n4167), .dinb(n4163), .dout(n4260));
  jor  g04069(.dina(n4260), .dinb(n4164), .dout(n4261));
  jand g04070(.dina(n4085), .dinb(n4083), .dout(n4262));
  jnot g04071(.din(n4262), .dout(n4263));
  jand g04072(.dina(n4263), .dinb(n4088), .dout(n4264));
  jxor g04073(.dina(n4264), .dinb(n4261), .dout(n4265));
  jxor g04074(.dina(n4265), .dinb(n4259), .dout(n4266));
  jand g04075(.dina(n4180), .dinb(n4177), .dout(n4267));
  jand g04076(.dina(n4184), .dinb(n4181), .dout(n4268));
  jor  g04077(.dina(n4268), .dinb(n4267), .dout(n4269));
  jxor g04078(.dina(n4269), .dinb(n4266), .dout(n4270));
  jxor g04079(.dina(n4270), .dinb(n4258), .dout(n4271));
  jxor g04080(.dina(n4271), .dinb(n4232), .dout(n4272));
  jxor g04081(.dina(n4272), .dinb(n4225), .dout(n4273));
  jxor g04082(.dina(n4273), .dinb(n4222), .dout(n4274));
  jand g04083(.dina(n4050), .dinb(n4047), .dout(n4275));
  jand g04084(.dina(n4103), .dinb(n4051), .dout(n4276));
  jor  g04085(.dina(n4276), .dinb(n4275), .dout(n4277));
  jor  g04086(.dina(n4206), .dinb(n4203), .dout(n4278));
  jand g04087(.dina(n4207), .dinb(n4199), .dout(n4279));
  jnot g04088(.din(n4279), .dout(n4280));
  jand g04089(.dina(n4280), .dinb(n4278), .dout(n4281));
  jnot g04090(.din(n4281), .dout(n4282));
  jor  g04091(.dina(n4099), .dinb(n4098), .dout(n4283));
  jand g04092(.dina(n4099), .dinb(n4098), .dout(n4284));
  jor  g04093(.dina(n4284), .dinb(n4097), .dout(n4285));
  jand g04094(.dina(n4285), .dinb(n4283), .dout(n4286));
  jnot g04095(.din(n4286), .dout(n4287));
  jand g04096(.dina(\a[30] ), .dinb(\a[16] ), .dout(n4288));
  jnot g04097(.din(n4288), .dout(n4289));
  jand g04098(.dina(n2653), .dinb(n1107), .dout(n4290));
  jnot g04099(.din(n4290), .dout(n4291));
  jand g04100(.dina(\a[29] ), .dinb(\a[17] ), .dout(n4292));
  jand g04101(.dina(\a[28] ), .dinb(\a[18] ), .dout(n4293));
  jor  g04102(.dina(n4293), .dinb(n4292), .dout(n4294));
  jand g04103(.dina(n4294), .dinb(n4291), .dout(n4295));
  jxor g04104(.dina(n4295), .dinb(n4289), .dout(n4296));
  jxor g04105(.dina(n4296), .dinb(n4287), .dout(n4297));
  jnot g04106(.din(n4297), .dout(n4298));
  jand g04107(.dina(\a[34] ), .dinb(\a[12] ), .dout(n4299));
  jnot g04108(.din(n4299), .dout(n4300));
  jand g04109(.dina(\a[39] ), .dinb(\a[8] ), .dout(n4301));
  jand g04110(.dina(n4301), .dinb(n4124), .dout(n4302));
  jnot g04111(.din(n4302), .dout(n4303));
  jand g04112(.dina(\a[39] ), .dinb(\a[7] ), .dout(n4304));
  jand g04113(.dina(\a[38] ), .dinb(\a[8] ), .dout(n4305));
  jor  g04114(.dina(n4305), .dinb(n4304), .dout(n4306));
  jand g04115(.dina(n4306), .dinb(n4303), .dout(n4307));
  jxor g04116(.dina(n4307), .dinb(n4300), .dout(n4308));
  jxor g04117(.dina(n4308), .dinb(n4298), .dout(n4309));
  jand g04118(.dina(\a[46] ), .dinb(\a[0] ), .dout(n4310));
  jnot g04119(.din(n4310), .dout(n4311));
  jand g04120(.dina(\a[42] ), .dinb(\a[4] ), .dout(n4312));
  jnot g04121(.din(n4312), .dout(n4313));
  jand g04122(.dina(n4313), .dinb(n4311), .dout(n4314));
  jand g04123(.dina(n4312), .dinb(n4310), .dout(n4315));
  jnot g04124(.din(n4315), .dout(n4316));
  jand g04125(.dina(\a[43] ), .dinb(\a[42] ), .dout(n4317));
  jand g04126(.dina(n4317), .dinb(n265), .dout(n4318));
  jand g04127(.dina(\a[43] ), .dinb(\a[3] ), .dout(n4319));
  jand g04128(.dina(n4319), .dinb(n4310), .dout(n4320));
  jor  g04129(.dina(n4320), .dinb(n4318), .dout(n4321));
  jnot g04130(.din(n4321), .dout(n4322));
  jand g04131(.dina(n4322), .dinb(n4316), .dout(n4323));
  jnot g04132(.din(n4323), .dout(n4324));
  jor  g04133(.dina(n4324), .dinb(n4314), .dout(n4325));
  jand g04134(.dina(n4321), .dinb(n4316), .dout(n4326));
  jnot g04135(.din(n4326), .dout(n4327));
  jand g04136(.dina(n4327), .dinb(n4319), .dout(n4328));
  jnot g04137(.din(n4328), .dout(n4329));
  jand g04138(.dina(n4329), .dinb(n4325), .dout(n4330));
  jand g04139(.dina(\a[37] ), .dinb(\a[9] ), .dout(n4331));
  jnot g04140(.din(n4331), .dout(n4332));
  jand g04141(.dina(n3243), .dinb(n655), .dout(n4333));
  jnot g04142(.din(n4333), .dout(n4334));
  jand g04143(.dina(\a[36] ), .dinb(\a[10] ), .dout(n4335));
  jand g04144(.dina(\a[35] ), .dinb(\a[11] ), .dout(n4336));
  jor  g04145(.dina(n4336), .dinb(n4335), .dout(n4337));
  jand g04146(.dina(n4337), .dinb(n4334), .dout(n4338));
  jxor g04147(.dina(n4338), .dinb(n4332), .dout(n4339));
  jxor g04148(.dina(n4339), .dinb(n4330), .dout(n4340));
  jnot g04149(.din(n4340), .dout(n4341));
  jand g04150(.dina(\a[27] ), .dinb(\a[19] ), .dout(n4342));
  jnot g04151(.din(n4342), .dout(n4343));
  jand g04152(.dina(n2128), .dinb(n1490), .dout(n4344));
  jnot g04153(.din(n4344), .dout(n4345));
  jand g04154(.dina(\a[26] ), .dinb(\a[20] ), .dout(n4346));
  jand g04155(.dina(\a[25] ), .dinb(\a[21] ), .dout(n4347));
  jor  g04156(.dina(n4347), .dinb(n4346), .dout(n4348));
  jand g04157(.dina(n4348), .dinb(n4345), .dout(n4349));
  jxor g04158(.dina(n4349), .dinb(n4343), .dout(n4350));
  jxor g04159(.dina(n4350), .dinb(n4341), .dout(n4351));
  jxor g04160(.dina(n4351), .dinb(n4309), .dout(n4352));
  jxor g04161(.dina(n4352), .dinb(n4282), .dout(n4353));
  jxor g04162(.dina(n4353), .dinb(n4277), .dout(n4354));
  jand g04163(.dina(n4169), .dinb(n4162), .dout(n4355));
  jand g04164(.dina(n4170), .dinb(n4159), .dout(n4356));
  jor  g04165(.dina(n4356), .dinb(n4355), .dout(n4357));
  jor  g04166(.dina(n4132), .dinb(n4123), .dout(n4358));
  jor  g04167(.dina(n4142), .dinb(n4134), .dout(n4359));
  jand g04168(.dina(n4359), .dinb(n4358), .dout(n4360));
  jnot g04169(.din(n4360), .dout(n4361));
  jxor g04170(.dina(n4361), .dinb(n4357), .dout(n4362));
  jand g04171(.dina(n4091), .dinb(n4081), .dout(n4363));
  jand g04172(.dina(n4101), .dinb(n4092), .dout(n4364));
  jor  g04173(.dina(n4364), .dinb(n4363), .dout(n4365));
  jxor g04174(.dina(n4365), .dinb(n4362), .dout(n4366));
  jand g04175(.dina(n4063), .dinb(n4060), .dout(n4367));
  jand g04176(.dina(n4102), .dinb(n4064), .dout(n4368));
  jor  g04177(.dina(n4368), .dinb(n4367), .dout(n4369));
  jnot g04178(.din(n4153), .dout(n4370));
  jand g04179(.dina(n4121), .dinb(n4114), .dout(n4371));
  jor  g04180(.dina(n4371), .dinb(n4116), .dout(n4372));
  jxor g04181(.dina(n4372), .dinb(n4370), .dout(n4373));
  jand g04182(.dina(n4127), .dinb(n4125), .dout(n4374));
  jnot g04183(.din(n4374), .dout(n4375));
  jand g04184(.dina(n4375), .dinb(n4130), .dout(n4376));
  jxor g04185(.dina(n4376), .dinb(n4373), .dout(n4377));
  jand g04186(.dina(n4055), .dinb(n4053), .dout(n4378));
  jand g04187(.dina(n4059), .dinb(n4056), .dout(n4379));
  jor  g04188(.dina(n4379), .dinb(n4378), .dout(n4380));
  jand g04189(.dina(\a[45] ), .dinb(\a[1] ), .dout(n4381));
  jxor g04190(.dina(n4381), .dinb(n1814), .dout(n4382));
  jxor g04191(.dina(n4382), .dinb(n4093), .dout(n4383));
  jand g04192(.dina(n4138), .dinb(n4136), .dout(n4384));
  jnot g04193(.din(n4384), .dout(n4385));
  jand g04194(.dina(n4385), .dinb(n4140), .dout(n4386));
  jxor g04195(.dina(n4386), .dinb(n4383), .dout(n4387));
  jxor g04196(.dina(n4387), .dinb(n4380), .dout(n4388));
  jxor g04197(.dina(n4388), .dinb(n4377), .dout(n4389));
  jxor g04198(.dina(n4389), .dinb(n4369), .dout(n4390));
  jxor g04199(.dina(n4390), .dinb(n4366), .dout(n4391));
  jxor g04200(.dina(n4391), .dinb(n4354), .dout(n4392));
  jnot g04201(.din(n4392), .dout(n4393));
  jxor g04202(.dina(n4393), .dinb(n4274), .dout(n4394));
  jnot g04203(.din(n4212), .dout(n4395));
  jor  g04204(.dina(n4218), .dinb(n4214), .dout(n4396));
  jand g04205(.dina(n4396), .dinb(n4395), .dout(n4397));
  jxor g04206(.dina(n4397), .dinb(n4394), .dout(\asquared[47] ));
  jand g04207(.dina(n4272), .dinb(n4225), .dout(n4399));
  jand g04208(.dina(n4273), .dinb(n4222), .dout(n4400));
  jor  g04209(.dina(n4400), .dinb(n4399), .dout(n4401));
  jand g04210(.dina(n4231), .dinb(n4228), .dout(n4402));
  jand g04211(.dina(n4271), .dinb(n4232), .dout(n4403));
  jor  g04212(.dina(n4403), .dinb(n4402), .dout(n4404));
  jand g04213(.dina(n4389), .dinb(n4369), .dout(n4405));
  jand g04214(.dina(n4390), .dinb(n4366), .dout(n4406));
  jor  g04215(.dina(n4406), .dinb(n4405), .dout(n4407));
  jxor g04216(.dina(n4407), .dinb(n4404), .dout(n4408));
  jand g04217(.dina(n4242), .dinb(n4000), .dout(n4409));
  jor  g04218(.dina(n4409), .dinb(n4240), .dout(n4410));
  jand g04219(.dina(n4345), .dinb(n4343), .dout(n4411));
  jnot g04220(.din(n4411), .dout(n4412));
  jand g04221(.dina(n4412), .dinb(n4348), .dout(n4413));
  jxor g04222(.dina(n4413), .dinb(n4410), .dout(n4414));
  jxor g04223(.dina(n4414), .dinb(n4324), .dout(n4415));
  jnot g04224(.din(n4415), .dout(n4416));
  jor  g04225(.dina(n4339), .dinb(n4330), .dout(n4417));
  jor  g04226(.dina(n4350), .dinb(n4341), .dout(n4418));
  jand g04227(.dina(n4418), .dinb(n4417), .dout(n4419));
  jxor g04228(.dina(n4419), .dinb(n4416), .dout(n4420));
  jand g04229(.dina(n4256), .dinb(n4243), .dout(n4421));
  jand g04230(.dina(n4257), .dinb(n4235), .dout(n4422));
  jor  g04231(.dina(n4422), .dinb(n4421), .dout(n4423));
  jxor g04232(.dina(n4423), .dinb(n4420), .dout(n4424));
  jand g04233(.dina(n4351), .dinb(n4309), .dout(n4425));
  jand g04234(.dina(n4352), .dinb(n4282), .dout(n4426));
  jor  g04235(.dina(n4426), .dinb(n4425), .dout(n4427));
  jand g04236(.dina(n4269), .dinb(n4266), .dout(n4428));
  jand g04237(.dina(n4270), .dinb(n4258), .dout(n4429));
  jor  g04238(.dina(n4429), .dinb(n4428), .dout(n4430));
  jxor g04239(.dina(n4430), .dinb(n4427), .dout(n4431));
  jxor g04240(.dina(n4431), .dinb(n4424), .dout(n4432));
  jxor g04241(.dina(n4432), .dinb(n4408), .dout(n4433));
  jand g04242(.dina(n4353), .dinb(n4277), .dout(n4434));
  jand g04243(.dina(n4391), .dinb(n4354), .dout(n4435));
  jor  g04244(.dina(n4435), .dinb(n4434), .dout(n4436));
  jand g04245(.dina(n4264), .dinb(n4261), .dout(n4437));
  jand g04246(.dina(n4265), .dinb(n4259), .dout(n4438));
  jor  g04247(.dina(n4438), .dinb(n4437), .dout(n4439));
  jand g04248(.dina(n4382), .dinb(n4093), .dout(n4440));
  jand g04249(.dina(n4386), .dinb(n4383), .dout(n4441));
  jor  g04250(.dina(n4441), .dinb(n4440), .dout(n4442));
  jand g04251(.dina(\a[34] ), .dinb(\a[13] ), .dout(n4443));
  jand g04252(.dina(\a[40] ), .dinb(\a[7] ), .dout(n4444));
  jand g04253(.dina(\a[35] ), .dinb(\a[12] ), .dout(n4445));
  jxor g04254(.dina(n4445), .dinb(n4444), .dout(n4446));
  jxor g04255(.dina(n4446), .dinb(n4443), .dout(n4447));
  jxor g04256(.dina(n4447), .dinb(n4442), .dout(n4448));
  jxor g04257(.dina(n4448), .dinb(n4439), .dout(n4449));
  jand g04258(.dina(n4387), .dinb(n4380), .dout(n4450));
  jand g04259(.dina(n4388), .dinb(n4377), .dout(n4451));
  jor  g04260(.dina(n4451), .dinb(n4450), .dout(n4452));
  jxor g04261(.dina(n4452), .dinb(n4449), .dout(n4453));
  jand g04262(.dina(n4361), .dinb(n4357), .dout(n4454));
  jand g04263(.dina(n4365), .dinb(n4362), .dout(n4455));
  jor  g04264(.dina(n4455), .dinb(n4454), .dout(n4456));
  jxor g04265(.dina(n4456), .dinb(n4453), .dout(n4457));
  jand g04266(.dina(n4381), .dinb(n1814), .dout(n4458));
  jand g04267(.dina(\a[47] ), .dinb(\a[0] ), .dout(n4459));
  jand g04268(.dina(\a[45] ), .dinb(\a[2] ), .dout(n4460));
  jor  g04269(.dina(n4460), .dinb(n4459), .dout(n4461));
  jand g04270(.dina(\a[47] ), .dinb(\a[2] ), .dout(n4462));
  jand g04271(.dina(n4462), .dinb(n4114), .dout(n4463));
  jnot g04272(.din(n4463), .dout(n4464));
  jand g04273(.dina(n4464), .dinb(n4461), .dout(n4465));
  jxor g04274(.dina(n4465), .dinb(n4458), .dout(n4466));
  jand g04275(.dina(\a[31] ), .dinb(\a[16] ), .dout(n4467));
  jand g04276(.dina(n3294), .dinb(n1107), .dout(n4468));
  jnot g04277(.din(n4468), .dout(n4469));
  jand g04278(.dina(\a[30] ), .dinb(\a[17] ), .dout(n4470));
  jand g04279(.dina(\a[29] ), .dinb(\a[18] ), .dout(n4471));
  jor  g04280(.dina(n4471), .dinb(n4470), .dout(n4472));
  jand g04281(.dina(n4472), .dinb(n4469), .dout(n4473));
  jxor g04282(.dina(n4473), .dinb(n4467), .dout(n4474));
  jxor g04283(.dina(n4474), .dinb(n4466), .dout(n4475));
  jnot g04284(.din(n4475), .dout(n4476));
  jand g04285(.dina(\a[28] ), .dinb(\a[19] ), .dout(n4477));
  jnot g04286(.din(n4477), .dout(n4478));
  jand g04287(.dina(n1927), .dinb(n1490), .dout(n4479));
  jnot g04288(.din(n4479), .dout(n4480));
  jand g04289(.dina(\a[27] ), .dinb(\a[20] ), .dout(n4481));
  jor  g04290(.dina(n4481), .dinb(n1834), .dout(n4482));
  jand g04291(.dina(n4482), .dinb(n4480), .dout(n4483));
  jxor g04292(.dina(n4483), .dinb(n4478), .dout(n4484));
  jxor g04293(.dina(n4484), .dinb(n4476), .dout(n4485));
  jor  g04294(.dina(n4250), .dinb(n4248), .dout(n4486));
  jand g04295(.dina(n4291), .dinb(n4289), .dout(n4487));
  jnot g04296(.din(n4487), .dout(n4488));
  jand g04297(.dina(n4488), .dinb(n4294), .dout(n4489));
  jxor g04298(.dina(n4489), .dinb(n4486), .dout(n4490));
  jand g04299(.dina(\a[44] ), .dinb(\a[3] ), .dout(n4491));
  jand g04300(.dina(\a[43] ), .dinb(\a[32] ), .dout(n4492));
  jand g04301(.dina(n4492), .dinb(n887), .dout(n4493));
  jnot g04302(.din(n4493), .dout(n4494));
  jand g04303(.dina(\a[44] ), .dinb(\a[43] ), .dout(n4495));
  jand g04304(.dina(n4495), .dinb(n265), .dout(n4496));
  jand g04305(.dina(\a[32] ), .dinb(\a[15] ), .dout(n4497));
  jand g04306(.dina(n4497), .dinb(n4491), .dout(n4498));
  jor  g04307(.dina(n4498), .dinb(n4496), .dout(n4499));
  jand g04308(.dina(n4499), .dinb(n4494), .dout(n4500));
  jnot g04309(.din(n4500), .dout(n4501));
  jand g04310(.dina(n4501), .dinb(n4491), .dout(n4502));
  jor  g04311(.dina(n4499), .dinb(n4493), .dout(n4503));
  jnot g04312(.din(n4503), .dout(n4504));
  jand g04313(.dina(\a[43] ), .dinb(\a[4] ), .dout(n4505));
  jor  g04314(.dina(n4505), .dinb(n4497), .dout(n4506));
  jand g04315(.dina(n4506), .dinb(n4504), .dout(n4507));
  jor  g04316(.dina(n4507), .dinb(n4502), .dout(n4508));
  jxor g04317(.dina(n4508), .dinb(n4490), .dout(n4509));
  jand g04318(.dina(\a[42] ), .dinb(\a[5] ), .dout(n4510));
  jand g04319(.dina(\a[41] ), .dinb(\a[33] ), .dout(n4511));
  jand g04320(.dina(n4511), .dinb(n990), .dout(n4512));
  jnot g04321(.din(n4512), .dout(n4513));
  jand g04322(.dina(\a[42] ), .dinb(\a[41] ), .dout(n4514));
  jand g04323(.dina(n4514), .dinb(n339), .dout(n4515));
  jand g04324(.dina(\a[33] ), .dinb(\a[14] ), .dout(n4516));
  jand g04325(.dina(n4516), .dinb(n4510), .dout(n4517));
  jor  g04326(.dina(n4517), .dinb(n4515), .dout(n4518));
  jand g04327(.dina(n4518), .dinb(n4513), .dout(n4519));
  jnot g04328(.din(n4519), .dout(n4520));
  jand g04329(.dina(n4520), .dinb(n4510), .dout(n4521));
  jand g04330(.dina(\a[41] ), .dinb(\a[6] ), .dout(n4522));
  jor  g04331(.dina(n4522), .dinb(n4516), .dout(n4523));
  jor  g04332(.dina(n4518), .dinb(n4512), .dout(n4524));
  jnot g04333(.din(n4524), .dout(n4525));
  jand g04334(.dina(n4525), .dinb(n4523), .dout(n4526));
  jor  g04335(.dina(n4526), .dinb(n4521), .dout(n4527));
  jand g04336(.dina(\a[38] ), .dinb(\a[36] ), .dout(n4528));
  jand g04337(.dina(n4528), .dinb(n959), .dout(n4529));
  jnot g04338(.din(n4529), .dout(n4530));
  jand g04339(.dina(\a[39] ), .dinb(\a[9] ), .dout(n4531));
  jand g04340(.dina(n4531), .dinb(n4305), .dout(n4532));
  jand g04341(.dina(\a[36] ), .dinb(\a[11] ), .dout(n4533));
  jand g04342(.dina(n4533), .dinb(n4301), .dout(n4534));
  jor  g04343(.dina(n4534), .dinb(n4532), .dout(n4535));
  jnot g04344(.din(n4535), .dout(n4536));
  jand g04345(.dina(n4536), .dinb(n4530), .dout(n4537));
  jand g04346(.dina(\a[38] ), .dinb(\a[9] ), .dout(n4538));
  jor  g04347(.dina(n4538), .dinb(n4533), .dout(n4539));
  jand g04348(.dina(n4539), .dinb(n4537), .dout(n4540));
  jand g04349(.dina(n4535), .dinb(n4530), .dout(n4541));
  jnot g04350(.din(n4541), .dout(n4542));
  jand g04351(.dina(n4542), .dinb(n4301), .dout(n4543));
  jor  g04352(.dina(n4543), .dinb(n4540), .dout(n4544));
  jand g04353(.dina(\a[37] ), .dinb(\a[10] ), .dout(n4545));
  jnot g04354(.din(n4545), .dout(n4546));
  jand g04355(.dina(n1658), .dinb(n1648), .dout(n4547));
  jnot g04356(.din(n4547), .dout(n4548));
  jand g04357(.dina(\a[25] ), .dinb(\a[22] ), .dout(n4549));
  jor  g04358(.dina(n4549), .dinb(n1942), .dout(n4550));
  jand g04359(.dina(n4550), .dinb(n4548), .dout(n4551));
  jxor g04360(.dina(n4551), .dinb(n4546), .dout(n4552));
  jnot g04361(.din(n4552), .dout(n4553));
  jxor g04362(.dina(n4553), .dinb(n4544), .dout(n4554));
  jxor g04363(.dina(n4554), .dinb(n4527), .dout(n4555));
  jxor g04364(.dina(n4555), .dinb(n4509), .dout(n4556));
  jxor g04365(.dina(n4556), .dinb(n4485), .dout(n4557));
  jor  g04366(.dina(n4296), .dinb(n4287), .dout(n4558));
  jor  g04367(.dina(n4308), .dinb(n4298), .dout(n4559));
  jand g04368(.dina(n4559), .dinb(n4558), .dout(n4560));
  jnot g04369(.din(n4560), .dout(n4561));
  jand g04370(.dina(n4372), .dinb(n4370), .dout(n4562));
  jand g04371(.dina(n4376), .dinb(n4373), .dout(n4563));
  jor  g04372(.dina(n4563), .dinb(n4562), .dout(n4564));
  jxor g04373(.dina(n4564), .dinb(n4561), .dout(n4565));
  jand g04374(.dina(\a[46] ), .dinb(\a[1] ), .dout(n4566));
  jor  g04375(.dina(n4566), .dinb(\a[24] ), .dout(n4567));
  jand g04376(.dina(n1386), .dinb(\a[46] ), .dout(n4568));
  jnot g04377(.din(n4568), .dout(n4569));
  jand g04378(.dina(n4569), .dinb(n4567), .dout(n4570));
  jand g04379(.dina(n4334), .dinb(n4332), .dout(n4571));
  jnot g04380(.din(n4571), .dout(n4572));
  jand g04381(.dina(n4572), .dinb(n4337), .dout(n4573));
  jxor g04382(.dina(n4573), .dinb(n4570), .dout(n4574));
  jand g04383(.dina(n4303), .dinb(n4300), .dout(n4575));
  jnot g04384(.din(n4575), .dout(n4576));
  jand g04385(.dina(n4576), .dinb(n4306), .dout(n4577));
  jxor g04386(.dina(n4577), .dinb(n4574), .dout(n4578));
  jxor g04387(.dina(n4578), .dinb(n4565), .dout(n4579));
  jxor g04388(.dina(n4579), .dinb(n4557), .dout(n4580));
  jxor g04389(.dina(n4580), .dinb(n4457), .dout(n4581));
  jxor g04390(.dina(n4581), .dinb(n4436), .dout(n4582));
  jxor g04391(.dina(n4582), .dinb(n4433), .dout(n4583));
  jand g04392(.dina(n4583), .dinb(n4401), .dout(n4584));
  jor  g04393(.dina(n4583), .dinb(n4401), .dout(n4585));
  jnot g04394(.din(n4585), .dout(n4586));
  jor  g04395(.dina(n4586), .dinb(n4584), .dout(n4587));
  jand g04396(.dina(n4392), .dinb(n4274), .dout(n4588));
  jnot g04397(.din(n4588), .dout(n4589));
  jnot g04398(.din(n4274), .dout(n4590));
  jand g04399(.dina(n4393), .dinb(n4590), .dout(n4591));
  jor  g04400(.dina(n4397), .dinb(n4591), .dout(n4592));
  jand g04401(.dina(n4592), .dinb(n4589), .dout(n4593));
  jxor g04402(.dina(n4593), .dinb(n4587), .dout(\asquared[48] ));
  jand g04403(.dina(n4581), .dinb(n4436), .dout(n4595));
  jand g04404(.dina(n4582), .dinb(n4433), .dout(n4596));
  jor  g04405(.dina(n4596), .dinb(n4595), .dout(n4597));
  jnot g04406(.din(n4597), .dout(n4598));
  jand g04407(.dina(n4407), .dinb(n4404), .dout(n4599));
  jand g04408(.dina(n4432), .dinb(n4408), .dout(n4600));
  jor  g04409(.dina(n4600), .dinb(n4599), .dout(n4601));
  jand g04410(.dina(n4430), .dinb(n4427), .dout(n4602));
  jand g04411(.dina(n4431), .dinb(n4424), .dout(n4603));
  jor  g04412(.dina(n4603), .dinb(n4602), .dout(n4604));
  jand g04413(.dina(n4452), .dinb(n4449), .dout(n4605));
  jand g04414(.dina(n4456), .dinb(n4453), .dout(n4606));
  jor  g04415(.dina(n4606), .dinb(n4605), .dout(n4607));
  jand g04416(.dina(n4447), .dinb(n4442), .dout(n4608));
  jand g04417(.dina(n4448), .dinb(n4439), .dout(n4609));
  jor  g04418(.dina(n4609), .dinb(n4608), .dout(n4610));
  jand g04419(.dina(\a[35] ), .dinb(\a[13] ), .dout(n4611));
  jand g04420(.dina(\a[42] ), .dinb(\a[6] ), .dout(n4612));
  jand g04421(.dina(n4612), .dinb(n4611), .dout(n4613));
  jnot g04422(.din(n4613), .dout(n4614));
  jand g04423(.dina(n2845), .dinb(n675), .dout(n4615));
  jand g04424(.dina(\a[34] ), .dinb(\a[14] ), .dout(n4616));
  jand g04425(.dina(n4616), .dinb(n4612), .dout(n4617));
  jor  g04426(.dina(n4617), .dinb(n4615), .dout(n4618));
  jnot g04427(.din(n4618), .dout(n4619));
  jand g04428(.dina(n4619), .dinb(n4614), .dout(n4620));
  jor  g04429(.dina(n4612), .dinb(n4611), .dout(n4621));
  jand g04430(.dina(n4621), .dinb(n4620), .dout(n4622));
  jand g04431(.dina(n4618), .dinb(n4614), .dout(n4623));
  jnot g04432(.din(n4623), .dout(n4624));
  jand g04433(.dina(n4624), .dinb(n4616), .dout(n4625));
  jor  g04434(.dina(n4625), .dinb(n4622), .dout(n4626));
  jand g04435(.dina(\a[41] ), .dinb(\a[7] ), .dout(n4627));
  jand g04436(.dina(\a[40] ), .dinb(\a[8] ), .dout(n4628));
  jand g04437(.dina(\a[36] ), .dinb(\a[12] ), .dout(n4629));
  jand g04438(.dina(n4629), .dinb(n4628), .dout(n4630));
  jnot g04439(.din(n4630), .dout(n4631));
  jand g04440(.dina(\a[41] ), .dinb(\a[40] ), .dout(n4632));
  jand g04441(.dina(n4632), .dinb(n499), .dout(n4633));
  jand g04442(.dina(n4629), .dinb(n4627), .dout(n4634));
  jor  g04443(.dina(n4634), .dinb(n4633), .dout(n4635));
  jand g04444(.dina(n4635), .dinb(n4631), .dout(n4636));
  jnot g04445(.din(n4636), .dout(n4637));
  jand g04446(.dina(n4637), .dinb(n4627), .dout(n4638));
  jor  g04447(.dina(n4629), .dinb(n4628), .dout(n4639));
  jor  g04448(.dina(n4635), .dinb(n4630), .dout(n4640));
  jnot g04449(.din(n4640), .dout(n4641));
  jand g04450(.dina(n4641), .dinb(n4639), .dout(n4642));
  jor  g04451(.dina(n4642), .dinb(n4638), .dout(n4643));
  jxor g04452(.dina(n4643), .dinb(n4626), .dout(n4644));
  jnot g04453(.din(n4531), .dout(n4645));
  jand g04454(.dina(\a[38] ), .dinb(\a[11] ), .dout(n4646));
  jand g04455(.dina(n4646), .dinb(n4545), .dout(n4647));
  jnot g04456(.din(n4647), .dout(n4648));
  jand g04457(.dina(\a[37] ), .dinb(\a[11] ), .dout(n4649));
  jand g04458(.dina(\a[38] ), .dinb(\a[10] ), .dout(n4650));
  jor  g04459(.dina(n4650), .dinb(n4649), .dout(n4651));
  jand g04460(.dina(n4651), .dinb(n4648), .dout(n4652));
  jxor g04461(.dina(n4652), .dinb(n4645), .dout(n4653));
  jnot g04462(.din(n4653), .dout(n4654));
  jxor g04463(.dina(n4654), .dinb(n4644), .dout(n4655));
  jxor g04464(.dina(n4655), .dinb(n4610), .dout(n4656));
  jand g04465(.dina(\a[44] ), .dinb(\a[4] ), .dout(n4657));
  jand g04466(.dina(\a[43] ), .dinb(\a[33] ), .dout(n4658));
  jand g04467(.dina(n4658), .dinb(n981), .dout(n4659));
  jnot g04468(.din(n4659), .dout(n4660));
  jand g04469(.dina(\a[43] ), .dinb(\a[5] ), .dout(n4661));
  jand g04470(.dina(\a[33] ), .dinb(\a[15] ), .dout(n4662));
  jor  g04471(.dina(n4662), .dinb(n4661), .dout(n4663));
  jand g04472(.dina(n4663), .dinb(n4660), .dout(n4664));
  jxor g04473(.dina(n4664), .dinb(n4657), .dout(n4665));
  jnot g04474(.din(n4665), .dout(n4666));
  jand g04475(.dina(\a[28] ), .dinb(\a[20] ), .dout(n4667));
  jnot g04476(.din(n4667), .dout(n4668));
  jand g04477(.dina(n1927), .dinb(n1376), .dout(n4669));
  jnot g04478(.din(n4669), .dout(n4670));
  jand g04479(.dina(\a[26] ), .dinb(\a[22] ), .dout(n4671));
  jand g04480(.dina(\a[27] ), .dinb(\a[21] ), .dout(n4672));
  jor  g04481(.dina(n4672), .dinb(n4671), .dout(n4673));
  jand g04482(.dina(n4673), .dinb(n4670), .dout(n4674));
  jxor g04483(.dina(n4674), .dinb(n4668), .dout(n4675));
  jxor g04484(.dina(n4675), .dinb(n4666), .dout(n4676));
  jand g04485(.dina(\a[31] ), .dinb(\a[17] ), .dout(n4677));
  jand g04486(.dina(n3294), .dinb(n1024), .dout(n4678));
  jnot g04487(.din(n4678), .dout(n4679));
  jand g04488(.dina(\a[30] ), .dinb(\a[18] ), .dout(n4680));
  jand g04489(.dina(\a[29] ), .dinb(\a[19] ), .dout(n4681));
  jor  g04490(.dina(n4681), .dinb(n4680), .dout(n4682));
  jand g04491(.dina(n4682), .dinb(n4679), .dout(n4683));
  jxor g04492(.dina(n4683), .dinb(n4677), .dout(n4684));
  jxor g04493(.dina(n4684), .dinb(n4676), .dout(n4685));
  jxor g04494(.dina(n4685), .dinb(n4656), .dout(n4686));
  jxor g04495(.dina(n4686), .dinb(n4607), .dout(n4687));
  jxor g04496(.dina(n4687), .dinb(n4604), .dout(n4688));
  jxor g04497(.dina(n4688), .dinb(n4601), .dout(n4689));
  jnot g04498(.din(n4537), .dout(n4690));
  jand g04499(.dina(n4480), .dinb(n4478), .dout(n4691));
  jnot g04500(.din(n4691), .dout(n4692));
  jand g04501(.dina(n4692), .dinb(n4482), .dout(n4693));
  jxor g04502(.dina(n4693), .dinb(n4690), .dout(n4694));
  jxor g04503(.dina(n4694), .dinb(n4524), .dout(n4695));
  jand g04504(.dina(n4553), .dinb(n4544), .dout(n4696));
  jand g04505(.dina(n4554), .dinb(n4527), .dout(n4697));
  jor  g04506(.dina(n4697), .dinb(n4696), .dout(n4698));
  jxor g04507(.dina(n4698), .dinb(n4695), .dout(n4699));
  jand g04508(.dina(n4548), .dinb(n4546), .dout(n4700));
  jnot g04509(.din(n4700), .dout(n4701));
  jand g04510(.dina(n4701), .dinb(n4550), .dout(n4702));
  jor  g04511(.dina(n4445), .dinb(n4444), .dout(n4703));
  jand g04512(.dina(n4445), .dinb(n4444), .dout(n4704));
  jor  g04513(.dina(n4704), .dinb(n4443), .dout(n4705));
  jand g04514(.dina(n4705), .dinb(n4703), .dout(n4706));
  jxor g04515(.dina(n4706), .dinb(n4702), .dout(n4707));
  jand g04516(.dina(\a[46] ), .dinb(\a[2] ), .dout(n4708));
  jnot g04517(.din(n4708), .dout(n4709));
  jand g04518(.dina(\a[45] ), .dinb(\a[3] ), .dout(n4710));
  jand g04519(.dina(\a[32] ), .dinb(\a[16] ), .dout(n4711));
  jxor g04520(.dina(n4711), .dinb(n4710), .dout(n4712));
  jxor g04521(.dina(n4712), .dinb(n4709), .dout(n4713));
  jnot g04522(.din(n4713), .dout(n4714));
  jxor g04523(.dina(n4714), .dinb(n4707), .dout(n4715));
  jxor g04524(.dina(n4715), .dinb(n4699), .dout(n4716));
  jand g04525(.dina(n4555), .dinb(n4509), .dout(n4717));
  jand g04526(.dina(n4556), .dinb(n4485), .dout(n4718));
  jor  g04527(.dina(n4718), .dinb(n4717), .dout(n4719));
  jxor g04528(.dina(n4719), .dinb(n4716), .dout(n4720));
  jand g04529(.dina(n4465), .dinb(n4458), .dout(n4721));
  jor  g04530(.dina(n4721), .dinb(n4463), .dout(n4722));
  jor  g04531(.dina(n4468), .dinb(n4467), .dout(n4723));
  jand g04532(.dina(n4723), .dinb(n4472), .dout(n4724));
  jxor g04533(.dina(n4724), .dinb(n4503), .dout(n4725));
  jxor g04534(.dina(n4725), .dinb(n4722), .dout(n4726));
  jand g04535(.dina(n4573), .dinb(n4570), .dout(n4727));
  jand g04536(.dina(n4577), .dinb(n4574), .dout(n4728));
  jor  g04537(.dina(n4728), .dinb(n4727), .dout(n4729));
  jnot g04538(.din(n4729), .dout(n4730));
  jand g04539(.dina(n4474), .dinb(n4466), .dout(n4731));
  jnot g04540(.din(n4731), .dout(n4732));
  jor  g04541(.dina(n4484), .dinb(n4476), .dout(n4733));
  jand g04542(.dina(n4733), .dinb(n4732), .dout(n4734));
  jxor g04543(.dina(n4734), .dinb(n4730), .dout(n4735));
  jxor g04544(.dina(n4735), .dinb(n4726), .dout(n4736));
  jxor g04545(.dina(n4736), .dinb(n4720), .dout(n4737));
  jand g04546(.dina(n4579), .dinb(n4557), .dout(n4738));
  jand g04547(.dina(n4580), .dinb(n4457), .dout(n4739));
  jor  g04548(.dina(n4739), .dinb(n4738), .dout(n4740));
  jor  g04549(.dina(n4419), .dinb(n4416), .dout(n4741));
  jand g04550(.dina(n4423), .dinb(n4420), .dout(n4742));
  jnot g04551(.din(n4742), .dout(n4743));
  jand g04552(.dina(n4743), .dinb(n4741), .dout(n4744));
  jnot g04553(.din(n4744), .dout(n4745));
  jand g04554(.dina(n4564), .dinb(n4561), .dout(n4746));
  jand g04555(.dina(n4578), .dinb(n4565), .dout(n4747));
  jor  g04556(.dina(n4747), .dinb(n4746), .dout(n4748));
  jxor g04557(.dina(n4748), .dinb(n4745), .dout(n4749));
  jand g04558(.dina(n4413), .dinb(n4410), .dout(n4750));
  jand g04559(.dina(n4414), .dinb(n4324), .dout(n4751));
  jor  g04560(.dina(n4751), .dinb(n4750), .dout(n4752));
  jand g04561(.dina(\a[48] ), .dinb(\a[0] ), .dout(n4753));
  jxor g04562(.dina(n4753), .dinb(n4568), .dout(n4754));
  jand g04563(.dina(\a[25] ), .dinb(\a[23] ), .dout(n4755));
  jand g04564(.dina(\a[47] ), .dinb(\a[1] ), .dout(n4756));
  jxor g04565(.dina(n4756), .dinb(n4755), .dout(n4757));
  jxor g04566(.dina(n4757), .dinb(n4754), .dout(n4758));
  jxor g04567(.dina(n4758), .dinb(n4752), .dout(n4759));
  jand g04568(.dina(n4489), .dinb(n4486), .dout(n4760));
  jand g04569(.dina(n4508), .dinb(n4490), .dout(n4761));
  jor  g04570(.dina(n4761), .dinb(n4760), .dout(n4762));
  jxor g04571(.dina(n4762), .dinb(n4759), .dout(n4763));
  jxor g04572(.dina(n4763), .dinb(n4749), .dout(n4764));
  jxor g04573(.dina(n4764), .dinb(n4740), .dout(n4765));
  jxor g04574(.dina(n4765), .dinb(n4737), .dout(n4766));
  jxor g04575(.dina(n4766), .dinb(n4689), .dout(n4767));
  jxor g04576(.dina(n4767), .dinb(n4598), .dout(n4768));
  jnot g04577(.din(n4584), .dout(n4769));
  jor  g04578(.dina(n4593), .dinb(n4586), .dout(n4770));
  jand g04579(.dina(n4770), .dinb(n4769), .dout(n4771));
  jxor g04580(.dina(n4771), .dinb(n4768), .dout(\asquared[49] ));
  jand g04581(.dina(n4764), .dinb(n4740), .dout(n4773));
  jand g04582(.dina(n4765), .dinb(n4737), .dout(n4774));
  jor  g04583(.dina(n4774), .dinb(n4773), .dout(n4775));
  jand g04584(.dina(n4719), .dinb(n4716), .dout(n4776));
  jand g04585(.dina(n4736), .dinb(n4720), .dout(n4777));
  jor  g04586(.dina(n4777), .dinb(n4776), .dout(n4778));
  jand g04587(.dina(n4748), .dinb(n4745), .dout(n4779));
  jand g04588(.dina(n4763), .dinb(n4749), .dout(n4780));
  jor  g04589(.dina(n4780), .dinb(n4779), .dout(n4781));
  jand g04590(.dina(\a[34] ), .dinb(\a[15] ), .dout(n4782));
  jand g04591(.dina(\a[43] ), .dinb(\a[35] ), .dout(n4783));
  jand g04592(.dina(n4783), .dinb(n990), .dout(n4784));
  jnot g04593(.din(n4784), .dout(n4785));
  jand g04594(.dina(\a[43] ), .dinb(\a[6] ), .dout(n4786));
  jand g04595(.dina(n4786), .dinb(n4782), .dout(n4787));
  jand g04596(.dina(n2845), .dinb(n976), .dout(n4788));
  jor  g04597(.dina(n4788), .dinb(n4787), .dout(n4789));
  jand g04598(.dina(n4789), .dinb(n4785), .dout(n4790));
  jnot g04599(.din(n4790), .dout(n4791));
  jand g04600(.dina(n4791), .dinb(n4782), .dout(n4792));
  jand g04601(.dina(\a[35] ), .dinb(\a[14] ), .dout(n4793));
  jor  g04602(.dina(n4793), .dinb(n4786), .dout(n4794));
  jor  g04603(.dina(n4789), .dinb(n4784), .dout(n4795));
  jnot g04604(.din(n4795), .dout(n4796));
  jand g04605(.dina(n4796), .dinb(n4794), .dout(n4797));
  jor  g04606(.dina(n4797), .dinb(n4792), .dout(n4798));
  jand g04607(.dina(\a[36] ), .dinb(\a[13] ), .dout(n4799));
  jand g04608(.dina(\a[42] ), .dinb(\a[7] ), .dout(n4800));
  jand g04609(.dina(\a[41] ), .dinb(\a[8] ), .dout(n4801));
  jor  g04610(.dina(n4801), .dinb(n4800), .dout(n4802));
  jand g04611(.dina(n4514), .dinb(n499), .dout(n4803));
  jnot g04612(.din(n4803), .dout(n4804));
  jand g04613(.dina(n4804), .dinb(n4802), .dout(n4805));
  jxor g04614(.dina(n4805), .dinb(n4799), .dout(n4806));
  jand g04615(.dina(\a[26] ), .dinb(\a[23] ), .dout(n4807));
  jxor g04616(.dina(n4807), .dinb(n1648), .dout(n4808));
  jxor g04617(.dina(n4808), .dinb(n4646), .dout(n4809));
  jxor g04618(.dina(n4809), .dinb(n4806), .dout(n4810));
  jxor g04619(.dina(n4810), .dinb(n4798), .dout(n4811));
  jand g04620(.dina(\a[45] ), .dinb(\a[44] ), .dout(n4812));
  jand g04621(.dina(n4812), .dinb(n242), .dout(n4813));
  jnot g04622(.din(n4813), .dout(n4814));
  jand g04623(.dina(n222), .dinb(\a[44] ), .dout(n4815));
  jand g04624(.dina(n4815), .dinb(\a[49] ), .dout(n4816));
  jand g04625(.dina(\a[45] ), .dinb(\a[4] ), .dout(n4817));
  jand g04626(.dina(\a[49] ), .dinb(\a[0] ), .dout(n4818));
  jand g04627(.dina(n4818), .dinb(n4817), .dout(n4819));
  jor  g04628(.dina(n4819), .dinb(n4816), .dout(n4820));
  jnot g04629(.din(n4820), .dout(n4821));
  jand g04630(.dina(n4821), .dinb(n4814), .dout(n4822));
  jand g04631(.dina(\a[44] ), .dinb(\a[5] ), .dout(n4823));
  jor  g04632(.dina(n4823), .dinb(n4817), .dout(n4824));
  jand g04633(.dina(n4824), .dinb(n4822), .dout(n4825));
  jand g04634(.dina(n4820), .dinb(n4814), .dout(n4826));
  jnot g04635(.din(n4826), .dout(n4827));
  jand g04636(.dina(n4827), .dinb(n4818), .dout(n4828));
  jor  g04637(.dina(n4828), .dinb(n4825), .dout(n4829));
  jand g04638(.dina(n4753), .dinb(n4568), .dout(n4830));
  jand g04639(.dina(n4757), .dinb(n4754), .dout(n4831));
  jor  g04640(.dina(n4831), .dinb(n4830), .dout(n4832));
  jxor g04641(.dina(n4832), .dinb(n4829), .dout(n4833));
  jand g04642(.dina(\a[33] ), .dinb(\a[16] ), .dout(n4834));
  jand g04643(.dina(n3269), .dinb(n1107), .dout(n4835));
  jnot g04644(.din(n4835), .dout(n4836));
  jand g04645(.dina(\a[32] ), .dinb(\a[17] ), .dout(n4837));
  jand g04646(.dina(\a[31] ), .dinb(\a[18] ), .dout(n4838));
  jor  g04647(.dina(n4838), .dinb(n4837), .dout(n4839));
  jand g04648(.dina(n4839), .dinb(n4836), .dout(n4840));
  jxor g04649(.dina(n4840), .dinb(n4834), .dout(n4841));
  jxor g04650(.dina(n4841), .dinb(n4833), .dout(n4842));
  jand g04651(.dina(\a[27] ), .dinb(\a[22] ), .dout(n4843));
  jand g04652(.dina(\a[46] ), .dinb(\a[3] ), .dout(n4844));
  jor  g04653(.dina(n4844), .dinb(n4462), .dout(n4845));
  jand g04654(.dina(\a[47] ), .dinb(\a[3] ), .dout(n4846));
  jand g04655(.dina(n4846), .dinb(n4708), .dout(n4847));
  jnot g04656(.din(n4847), .dout(n4848));
  jand g04657(.dina(n4848), .dinb(n4845), .dout(n4849));
  jxor g04658(.dina(n4849), .dinb(n4843), .dout(n4850));
  jnot g04659(.din(n4850), .dout(n4851));
  jand g04660(.dina(\a[30] ), .dinb(\a[19] ), .dout(n4852));
  jnot g04661(.din(n4852), .dout(n4853));
  jand g04662(.dina(n2653), .dinb(n1490), .dout(n4854));
  jnot g04663(.din(n4854), .dout(n4855));
  jand g04664(.dina(\a[28] ), .dinb(\a[21] ), .dout(n4856));
  jand g04665(.dina(\a[29] ), .dinb(\a[20] ), .dout(n4857));
  jor  g04666(.dina(n4857), .dinb(n4856), .dout(n4858));
  jand g04667(.dina(n4858), .dinb(n4855), .dout(n4859));
  jxor g04668(.dina(n4859), .dinb(n4853), .dout(n4860));
  jxor g04669(.dina(n4860), .dinb(n4851), .dout(n4861));
  jnot g04670(.din(n4861), .dout(n4862));
  jand g04671(.dina(\a[40] ), .dinb(\a[9] ), .dout(n4863));
  jnot g04672(.din(n4863), .dout(n4864));
  jand g04673(.dina(\a[39] ), .dinb(\a[37] ), .dout(n4865));
  jand g04674(.dina(n4865), .dinb(n1151), .dout(n4866));
  jnot g04675(.din(n4866), .dout(n4867));
  jand g04676(.dina(\a[37] ), .dinb(\a[12] ), .dout(n4868));
  jand g04677(.dina(\a[39] ), .dinb(\a[10] ), .dout(n4869));
  jor  g04678(.dina(n4869), .dinb(n4868), .dout(n4870));
  jand g04679(.dina(n4870), .dinb(n4867), .dout(n4871));
  jxor g04680(.dina(n4871), .dinb(n4864), .dout(n4872));
  jxor g04681(.dina(n4872), .dinb(n4862), .dout(n4873));
  jxor g04682(.dina(n4873), .dinb(n4842), .dout(n4874));
  jxor g04683(.dina(n4874), .dinb(n4811), .dout(n4875));
  jxor g04684(.dina(n4875), .dinb(n4781), .dout(n4876));
  jxor g04685(.dina(n4876), .dinb(n4778), .dout(n4877));
  jxor g04686(.dina(n4877), .dinb(n4775), .dout(n4878));
  jnot g04687(.din(n4620), .dout(n4879));
  jor  g04688(.dina(n4678), .dinb(n4677), .dout(n4880));
  jand g04689(.dina(n4880), .dinb(n4682), .dout(n4881));
  jxor g04690(.dina(n4881), .dinb(n4879), .dout(n4882));
  jxor g04691(.dina(n4882), .dinb(n4640), .dout(n4883));
  jnot g04692(.din(n4883), .dout(n4884));
  jor  g04693(.dina(n4675), .dinb(n4666), .dout(n4885));
  jand g04694(.dina(n4684), .dinb(n4676), .dout(n4886));
  jnot g04695(.din(n4886), .dout(n4887));
  jand g04696(.dina(n4887), .dinb(n4885), .dout(n4888));
  jxor g04697(.dina(n4888), .dinb(n4884), .dout(n4889));
  jand g04698(.dina(n4758), .dinb(n4752), .dout(n4890));
  jand g04699(.dina(n4762), .dinb(n4759), .dout(n4891));
  jor  g04700(.dina(n4891), .dinb(n4890), .dout(n4892));
  jxor g04701(.dina(n4892), .dinb(n4889), .dout(n4893));
  jand g04702(.dina(n4655), .dinb(n4610), .dout(n4894));
  jand g04703(.dina(n4685), .dinb(n4656), .dout(n4895));
  jor  g04704(.dina(n4895), .dinb(n4894), .dout(n4896));
  jxor g04705(.dina(n4896), .dinb(n4893), .dout(n4897));
  jand g04706(.dina(n4664), .dinb(n4657), .dout(n4898));
  jor  g04707(.dina(n4898), .dinb(n4659), .dout(n4899));
  jor  g04708(.dina(n4711), .dinb(n4710), .dout(n4900));
  jand g04709(.dina(n4711), .dinb(n4710), .dout(n4901));
  jor  g04710(.dina(n4901), .dinb(n4708), .dout(n4902));
  jand g04711(.dina(n4902), .dinb(n4900), .dout(n4903));
  jxor g04712(.dina(n4903), .dinb(n4899), .dout(n4904));
  jand g04713(.dina(n4670), .dinb(n4668), .dout(n4905));
  jnot g04714(.din(n4905), .dout(n4906));
  jand g04715(.dina(n4906), .dinb(n4673), .dout(n4907));
  jxor g04716(.dina(n4907), .dinb(n4904), .dout(n4908));
  jand g04717(.dina(n4643), .dinb(n4626), .dout(n4909));
  jand g04718(.dina(n4654), .dinb(n4644), .dout(n4910));
  jor  g04719(.dina(n4910), .dinb(n4909), .dout(n4911));
  jand g04720(.dina(\a[48] ), .dinb(\a[1] ), .dout(n4912));
  jnot g04721(.din(\a[25] ), .dout(n4913));
  jand g04722(.dina(n4756), .dinb(n4755), .dout(n4914));
  jor  g04723(.dina(n4914), .dinb(n4913), .dout(n4915));
  jxor g04724(.dina(n4915), .dinb(n4912), .dout(n4916));
  jnot g04725(.din(n4916), .dout(n4917));
  jand g04726(.dina(n4648), .dinb(n4645), .dout(n4918));
  jnot g04727(.din(n4918), .dout(n4919));
  jand g04728(.dina(n4919), .dinb(n4651), .dout(n4920));
  jxor g04729(.dina(n4920), .dinb(n4917), .dout(n4921));
  jxor g04730(.dina(n4921), .dinb(n4911), .dout(n4922));
  jxor g04731(.dina(n4922), .dinb(n4908), .dout(n4923));
  jxor g04732(.dina(n4923), .dinb(n4897), .dout(n4924));
  jand g04733(.dina(n4686), .dinb(n4607), .dout(n4925));
  jand g04734(.dina(n4687), .dinb(n4604), .dout(n4926));
  jor  g04735(.dina(n4926), .dinb(n4925), .dout(n4927));
  jand g04736(.dina(n4693), .dinb(n4690), .dout(n4928));
  jand g04737(.dina(n4694), .dinb(n4524), .dout(n4929));
  jor  g04738(.dina(n4929), .dinb(n4928), .dout(n4930));
  jand g04739(.dina(n4706), .dinb(n4702), .dout(n4931));
  jand g04740(.dina(n4714), .dinb(n4707), .dout(n4932));
  jor  g04741(.dina(n4932), .dinb(n4931), .dout(n4933));
  jxor g04742(.dina(n4933), .dinb(n4930), .dout(n4934));
  jand g04743(.dina(n4724), .dinb(n4503), .dout(n4935));
  jand g04744(.dina(n4725), .dinb(n4722), .dout(n4936));
  jor  g04745(.dina(n4936), .dinb(n4935), .dout(n4937));
  jxor g04746(.dina(n4937), .dinb(n4934), .dout(n4938));
  jand g04747(.dina(n4698), .dinb(n4695), .dout(n4939));
  jand g04748(.dina(n4715), .dinb(n4699), .dout(n4940));
  jor  g04749(.dina(n4940), .dinb(n4939), .dout(n4941));
  jnot g04750(.din(n4941), .dout(n4942));
  jor  g04751(.dina(n4734), .dinb(n4730), .dout(n4943));
  jand g04752(.dina(n4735), .dinb(n4726), .dout(n4944));
  jnot g04753(.din(n4944), .dout(n4945));
  jand g04754(.dina(n4945), .dinb(n4943), .dout(n4946));
  jxor g04755(.dina(n4946), .dinb(n4942), .dout(n4947));
  jxor g04756(.dina(n4947), .dinb(n4938), .dout(n4948));
  jxor g04757(.dina(n4948), .dinb(n4927), .dout(n4949));
  jxor g04758(.dina(n4949), .dinb(n4924), .dout(n4950));
  jxor g04759(.dina(n4950), .dinb(n4878), .dout(n4951));
  jnot g04760(.din(n4951), .dout(n4952));
  jand g04761(.dina(n4688), .dinb(n4601), .dout(n4953));
  jand g04762(.dina(n4766), .dinb(n4689), .dout(n4954));
  jor  g04763(.dina(n4954), .dinb(n4953), .dout(n4955));
  jxor g04764(.dina(n4955), .dinb(n4952), .dout(n4956));
  jand g04765(.dina(n4767), .dinb(n4597), .dout(n4957));
  jnot g04766(.din(n4957), .dout(n4958));
  jnot g04767(.din(n4767), .dout(n4959));
  jand g04768(.dina(n4959), .dinb(n4598), .dout(n4960));
  jor  g04769(.dina(n4771), .dinb(n4960), .dout(n4961));
  jand g04770(.dina(n4961), .dinb(n4958), .dout(n4962));
  jxor g04771(.dina(n4962), .dinb(n4956), .dout(\asquared[50] ));
  jand g04772(.dina(n4877), .dinb(n4775), .dout(n4964));
  jand g04773(.dina(n4950), .dinb(n4878), .dout(n4965));
  jor  g04774(.dina(n4965), .dinb(n4964), .dout(n4966));
  jnot g04775(.din(n4966), .dout(n4967));
  jand g04776(.dina(n4948), .dinb(n4927), .dout(n4968));
  jand g04777(.dina(n4949), .dinb(n4924), .dout(n4969));
  jor  g04778(.dina(n4969), .dinb(n4968), .dout(n4970));
  jand g04779(.dina(n4896), .dinb(n4893), .dout(n4971));
  jand g04780(.dina(n4923), .dinb(n4897), .dout(n4972));
  jor  g04781(.dina(n4972), .dinb(n4971), .dout(n4973));
  jor  g04782(.dina(n4946), .dinb(n4942), .dout(n4974));
  jand g04783(.dina(n4947), .dinb(n4938), .dout(n4975));
  jnot g04784(.din(n4975), .dout(n4976));
  jand g04785(.dina(n4976), .dinb(n4974), .dout(n4977));
  jnot g04786(.din(n4977), .dout(n4978));
  jand g04787(.dina(n4920), .dinb(n4917), .dout(n4979));
  jnot g04788(.din(\a[48] ), .dout(n4980));
  jand g04789(.dina(n4914), .dinb(n4980), .dout(n4981));
  jor  g04790(.dina(n4981), .dinb(n4979), .dout(n4982));
  jand g04791(.dina(\a[45] ), .dinb(\a[35] ), .dout(n4983));
  jand g04792(.dina(n4983), .dinb(n981), .dout(n4984));
  jnot g04793(.din(n4984), .dout(n4985));
  jand g04794(.dina(\a[45] ), .dinb(\a[5] ), .dout(n4986));
  jand g04795(.dina(\a[34] ), .dinb(\a[16] ), .dout(n4987));
  jand g04796(.dina(n4987), .dinb(n4986), .dout(n4988));
  jand g04797(.dina(n2845), .dinb(n829), .dout(n4989));
  jor  g04798(.dina(n4989), .dinb(n4988), .dout(n4990));
  jnot g04799(.din(n4990), .dout(n4991));
  jand g04800(.dina(n4991), .dinb(n4985), .dout(n4992));
  jand g04801(.dina(\a[35] ), .dinb(\a[15] ), .dout(n4993));
  jor  g04802(.dina(n4993), .dinb(n4986), .dout(n4994));
  jand g04803(.dina(n4994), .dinb(n4992), .dout(n4995));
  jand g04804(.dina(n4990), .dinb(n4985), .dout(n4996));
  jnot g04805(.din(n4996), .dout(n4997));
  jand g04806(.dina(n4997), .dinb(n4987), .dout(n4998));
  jor  g04807(.dina(n4998), .dinb(n4995), .dout(n4999));
  jand g04808(.dina(\a[28] ), .dinb(\a[22] ), .dout(n5000));
  jand g04809(.dina(\a[32] ), .dinb(\a[18] ), .dout(n5001));
  jand g04810(.dina(\a[27] ), .dinb(\a[23] ), .dout(n5002));
  jxor g04811(.dina(n5002), .dinb(n5001), .dout(n5003));
  jxor g04812(.dina(n5003), .dinb(n5000), .dout(n5004));
  jxor g04813(.dina(n5004), .dinb(n4999), .dout(n5005));
  jxor g04814(.dina(n5005), .dinb(n4982), .dout(n5006));
  jand g04815(.dina(\a[46] ), .dinb(\a[33] ), .dout(n5007));
  jand g04816(.dina(n5007), .dinb(n1044), .dout(n5008));
  jnot g04817(.din(n5008), .dout(n5009));
  jand g04818(.dina(\a[47] ), .dinb(\a[4] ), .dout(n5010));
  jand g04819(.dina(n5010), .dinb(n4844), .dout(n5011));
  jand g04820(.dina(\a[33] ), .dinb(\a[17] ), .dout(n5012));
  jand g04821(.dina(n5012), .dinb(n4846), .dout(n5013));
  jor  g04822(.dina(n5013), .dinb(n5011), .dout(n5014));
  jand g04823(.dina(n5014), .dinb(n5009), .dout(n5015));
  jnot g04824(.din(n5015), .dout(n5016));
  jand g04825(.dina(n5016), .dinb(n4846), .dout(n5017));
  jor  g04826(.dina(n5014), .dinb(n5008), .dout(n5018));
  jnot g04827(.din(n5018), .dout(n5019));
  jand g04828(.dina(\a[46] ), .dinb(\a[4] ), .dout(n5020));
  jor  g04829(.dina(n5020), .dinb(n5012), .dout(n5021));
  jand g04830(.dina(n5021), .dinb(n5019), .dout(n5022));
  jor  g04831(.dina(n5022), .dinb(n5017), .dout(n5023));
  jand g04832(.dina(n1446), .dinb(\a[48] ), .dout(n5024));
  jand g04833(.dina(\a[50] ), .dinb(\a[0] ), .dout(n5025));
  jand g04834(.dina(\a[48] ), .dinb(\a[2] ), .dout(n5026));
  jor  g04835(.dina(n5026), .dinb(n5025), .dout(n5027));
  jand g04836(.dina(\a[50] ), .dinb(\a[2] ), .dout(n5028));
  jand g04837(.dina(n5028), .dinb(n4753), .dout(n5029));
  jnot g04838(.din(n5029), .dout(n5030));
  jand g04839(.dina(n5030), .dinb(n5027), .dout(n5031));
  jxor g04840(.dina(n5031), .dinb(n5024), .dout(n5032));
  jxor g04841(.dina(n5032), .dinb(n5023), .dout(n5033));
  jnot g04842(.din(n5033), .dout(n5034));
  jand g04843(.dina(\a[31] ), .dinb(\a[19] ), .dout(n5035));
  jnot g04844(.din(n5035), .dout(n5036));
  jand g04845(.dina(n3294), .dinb(n1490), .dout(n5037));
  jnot g04846(.din(n5037), .dout(n5038));
  jand g04847(.dina(\a[30] ), .dinb(\a[20] ), .dout(n5039));
  jand g04848(.dina(\a[29] ), .dinb(\a[21] ), .dout(n5040));
  jor  g04849(.dina(n5040), .dinb(n5039), .dout(n5041));
  jand g04850(.dina(n5041), .dinb(n5038), .dout(n5042));
  jxor g04851(.dina(n5042), .dinb(n5036), .dout(n5043));
  jxor g04852(.dina(n5043), .dinb(n5034), .dout(n5044));
  jand g04853(.dina(\a[42] ), .dinb(\a[8] ), .dout(n5045));
  jand g04854(.dina(\a[41] ), .dinb(\a[37] ), .dout(n5046));
  jand g04855(.dina(n5046), .dinb(n479), .dout(n5047));
  jnot g04856(.din(n5047), .dout(n5048));
  jand g04857(.dina(n4514), .dinb(n395), .dout(n5049));
  jand g04858(.dina(\a[37] ), .dinb(\a[13] ), .dout(n5050));
  jand g04859(.dina(n5050), .dinb(n5045), .dout(n5051));
  jor  g04860(.dina(n5051), .dinb(n5049), .dout(n5052));
  jand g04861(.dina(n5052), .dinb(n5048), .dout(n5053));
  jnot g04862(.din(n5053), .dout(n5054));
  jand g04863(.dina(n5054), .dinb(n5045), .dout(n5055));
  jor  g04864(.dina(n5052), .dinb(n5047), .dout(n5056));
  jnot g04865(.din(n5056), .dout(n5057));
  jand g04866(.dina(\a[41] ), .dinb(\a[9] ), .dout(n5058));
  jor  g04867(.dina(n5058), .dinb(n5050), .dout(n5059));
  jand g04868(.dina(n5059), .dinb(n5057), .dout(n5060));
  jor  g04869(.dina(n5060), .dinb(n5055), .dout(n5061));
  jand g04870(.dina(\a[44] ), .dinb(\a[6] ), .dout(n5062));
  jand g04871(.dina(\a[43] ), .dinb(\a[7] ), .dout(n5063));
  jand g04872(.dina(\a[36] ), .dinb(\a[14] ), .dout(n5064));
  jxor g04873(.dina(n5064), .dinb(n5063), .dout(n5065));
  jxor g04874(.dina(n5065), .dinb(n5062), .dout(n5066));
  jxor g04875(.dina(n5066), .dinb(n5061), .dout(n5067));
  jnot g04876(.din(n5067), .dout(n5068));
  jand g04877(.dina(\a[38] ), .dinb(\a[12] ), .dout(n5069));
  jnot g04878(.din(n5069), .dout(n5070));
  jand g04879(.dina(n3665), .dinb(n655), .dout(n5071));
  jnot g04880(.din(n5071), .dout(n5072));
  jand g04881(.dina(\a[39] ), .dinb(\a[11] ), .dout(n5073));
  jand g04882(.dina(\a[40] ), .dinb(\a[10] ), .dout(n5074));
  jor  g04883(.dina(n5074), .dinb(n5073), .dout(n5075));
  jand g04884(.dina(n5075), .dinb(n5072), .dout(n5076));
  jxor g04885(.dina(n5076), .dinb(n5070), .dout(n5077));
  jxor g04886(.dina(n5077), .dinb(n5068), .dout(n5078));
  jxor g04887(.dina(n5078), .dinb(n5044), .dout(n5079));
  jxor g04888(.dina(n5079), .dinb(n5006), .dout(n5080));
  jxor g04889(.dina(n5080), .dinb(n4978), .dout(n5081));
  jxor g04890(.dina(n5081), .dinb(n4973), .dout(n5082));
  jxor g04891(.dina(n5082), .dinb(n4970), .dout(n5083));
  jand g04892(.dina(n4875), .dinb(n4781), .dout(n5084));
  jand g04893(.dina(n4876), .dinb(n4778), .dout(n5085));
  jor  g04894(.dina(n5085), .dinb(n5084), .dout(n5086));
  jor  g04895(.dina(n4888), .dinb(n4884), .dout(n5087));
  jand g04896(.dina(n4892), .dinb(n4889), .dout(n5088));
  jnot g04897(.din(n5088), .dout(n5089));
  jand g04898(.dina(n5089), .dinb(n5087), .dout(n5090));
  jnot g04899(.din(n5090), .dout(n5091));
  jand g04900(.dina(n4921), .dinb(n4911), .dout(n5092));
  jand g04901(.dina(n4922), .dinb(n4908), .dout(n5093));
  jor  g04902(.dina(n5093), .dinb(n5092), .dout(n5094));
  jxor g04903(.dina(n5094), .dinb(n5091), .dout(n5095));
  jand g04904(.dina(n4881), .dinb(n4879), .dout(n5096));
  jand g04905(.dina(n4882), .dinb(n4640), .dout(n5097));
  jor  g04906(.dina(n5097), .dinb(n5096), .dout(n5098));
  jand g04907(.dina(n4903), .dinb(n4899), .dout(n5099));
  jand g04908(.dina(n4907), .dinb(n4904), .dout(n5100));
  jor  g04909(.dina(n5100), .dinb(n5099), .dout(n5101));
  jxor g04910(.dina(n5101), .dinb(n5098), .dout(n5102));
  jnot g04911(.din(n4822), .dout(n5103));
  jand g04912(.dina(n4849), .dinb(n4843), .dout(n5104));
  jor  g04913(.dina(n5104), .dinb(n4847), .dout(n5105));
  jxor g04914(.dina(n5105), .dinb(n5103), .dout(n5106));
  jxor g04915(.dina(n5106), .dinb(n4795), .dout(n5107));
  jxor g04916(.dina(n5107), .dinb(n5102), .dout(n5108));
  jxor g04917(.dina(n5108), .dinb(n5095), .dout(n5109));
  jxor g04918(.dina(n5109), .dinb(n5086), .dout(n5110));
  jor  g04919(.dina(n4860), .dinb(n4851), .dout(n5111));
  jor  g04920(.dina(n4872), .dinb(n4862), .dout(n5112));
  jand g04921(.dina(n5112), .dinb(n5111), .dout(n5113));
  jnot g04922(.din(n5113), .dout(n5114));
  jand g04923(.dina(n4832), .dinb(n4829), .dout(n5115));
  jand g04924(.dina(n4841), .dinb(n4833), .dout(n5116));
  jor  g04925(.dina(n5116), .dinb(n5115), .dout(n5117));
  jxor g04926(.dina(n5117), .dinb(n5114), .dout(n5118));
  jand g04927(.dina(n4807), .dinb(n1648), .dout(n5119));
  jand g04928(.dina(n4808), .dinb(n4646), .dout(n5120));
  jor  g04929(.dina(n5120), .dinb(n5119), .dout(n5121));
  jand g04930(.dina(\a[49] ), .dinb(\a[1] ), .dout(n5122));
  jxor g04931(.dina(n5122), .dinb(n2022), .dout(n5123));
  jxor g04932(.dina(n5123), .dinb(n5121), .dout(n5124));
  jand g04933(.dina(n4867), .dinb(n4864), .dout(n5125));
  jnot g04934(.din(n5125), .dout(n5126));
  jand g04935(.dina(n5126), .dinb(n4870), .dout(n5127));
  jxor g04936(.dina(n5127), .dinb(n5124), .dout(n5128));
  jxor g04937(.dina(n5128), .dinb(n5118), .dout(n5129));
  jand g04938(.dina(n4805), .dinb(n4799), .dout(n5130));
  jor  g04939(.dina(n5130), .dinb(n4803), .dout(n5131));
  jor  g04940(.dina(n4835), .dinb(n4834), .dout(n5132));
  jand g04941(.dina(n5132), .dinb(n4839), .dout(n5133));
  jand g04942(.dina(n4855), .dinb(n4853), .dout(n5134));
  jnot g04943(.din(n5134), .dout(n5135));
  jand g04944(.dina(n5135), .dinb(n4858), .dout(n5136));
  jxor g04945(.dina(n5136), .dinb(n5133), .dout(n5137));
  jxor g04946(.dina(n5137), .dinb(n5131), .dout(n5138));
  jand g04947(.dina(n4809), .dinb(n4806), .dout(n5139));
  jand g04948(.dina(n4810), .dinb(n4798), .dout(n5140));
  jor  g04949(.dina(n5140), .dinb(n5139), .dout(n5141));
  jxor g04950(.dina(n5141), .dinb(n5138), .dout(n5142));
  jand g04951(.dina(n4933), .dinb(n4930), .dout(n5143));
  jand g04952(.dina(n4937), .dinb(n4934), .dout(n5144));
  jor  g04953(.dina(n5144), .dinb(n5143), .dout(n5145));
  jxor g04954(.dina(n5145), .dinb(n5142), .dout(n5146));
  jand g04955(.dina(n4873), .dinb(n4842), .dout(n5147));
  jand g04956(.dina(n4874), .dinb(n4811), .dout(n5148));
  jor  g04957(.dina(n5148), .dinb(n5147), .dout(n5149));
  jxor g04958(.dina(n5149), .dinb(n5146), .dout(n5150));
  jxor g04959(.dina(n5150), .dinb(n5129), .dout(n5151));
  jxor g04960(.dina(n5151), .dinb(n5110), .dout(n5152));
  jxor g04961(.dina(n5152), .dinb(n5083), .dout(n5153));
  jxor g04962(.dina(n5153), .dinb(n4967), .dout(n5154));
  jand g04963(.dina(n4955), .dinb(n4951), .dout(n5155));
  jnot g04964(.din(n5155), .dout(n5156));
  jnot g04965(.din(n4955), .dout(n5157));
  jand g04966(.dina(n5157), .dinb(n4952), .dout(n5158));
  jor  g04967(.dina(n4962), .dinb(n5158), .dout(n5159));
  jand g04968(.dina(n5159), .dinb(n5156), .dout(n5160));
  jxor g04969(.dina(n5160), .dinb(n5154), .dout(\asquared[51] ));
  jand g04970(.dina(n5082), .dinb(n4970), .dout(n5162));
  jand g04971(.dina(n5152), .dinb(n5083), .dout(n5163));
  jor  g04972(.dina(n5163), .dinb(n5162), .dout(n5164));
  jand g04973(.dina(n5109), .dinb(n5086), .dout(n5165));
  jand g04974(.dina(n5151), .dinb(n5110), .dout(n5166));
  jor  g04975(.dina(n5166), .dinb(n5165), .dout(n5167));
  jand g04976(.dina(n5149), .dinb(n5146), .dout(n5168));
  jand g04977(.dina(n5150), .dinb(n5129), .dout(n5169));
  jor  g04978(.dina(n5169), .dinb(n5168), .dout(n5170));
  jand g04979(.dina(n5094), .dinb(n5091), .dout(n5171));
  jand g04980(.dina(n5108), .dinb(n5095), .dout(n5172));
  jor  g04981(.dina(n5172), .dinb(n5171), .dout(n5173));
  jand g04982(.dina(n5136), .dinb(n5133), .dout(n5174));
  jand g04983(.dina(n5137), .dinb(n5131), .dout(n5175));
  jor  g04984(.dina(n5175), .dinb(n5174), .dout(n5176));
  jand g04985(.dina(n5122), .dinb(n2022), .dout(n5177));
  jand g04986(.dina(\a[51] ), .dinb(\a[0] ), .dout(n5178));
  jxor g04987(.dina(n5178), .dinb(n5177), .dout(n5179));
  jand g04988(.dina(\a[50] ), .dinb(\a[1] ), .dout(n5180));
  jxor g04989(.dina(n5180), .dinb(\a[26] ), .dout(n5181));
  jxor g04990(.dina(n5181), .dinb(n5179), .dout(n5182));
  jnot g04991(.din(n5182), .dout(n5183));
  jand g04992(.dina(\a[34] ), .dinb(\a[17] ), .dout(n5184));
  jnot g04993(.din(n5184), .dout(n5185));
  jand g04994(.dina(n3269), .dinb(n1287), .dout(n5186));
  jnot g04995(.din(n5186), .dout(n5187));
  jand g04996(.dina(\a[31] ), .dinb(\a[20] ), .dout(n5188));
  jand g04997(.dina(\a[32] ), .dinb(\a[19] ), .dout(n5189));
  jor  g04998(.dina(n5189), .dinb(n5188), .dout(n5190));
  jand g04999(.dina(n5190), .dinb(n5187), .dout(n5191));
  jxor g05000(.dina(n5191), .dinb(n5185), .dout(n5192));
  jxor g05001(.dina(n5192), .dinb(n5183), .dout(n5193));
  jxor g05002(.dina(n5193), .dinb(n5176), .dout(n5194));
  jand g05003(.dina(\a[36] ), .dinb(\a[15] ), .dout(n5195));
  jand g05004(.dina(\a[45] ), .dinb(\a[37] ), .dout(n5196));
  jand g05005(.dina(n5196), .dinb(n990), .dout(n5197));
  jnot g05006(.din(n5197), .dout(n5198));
  jand g05007(.dina(\a[45] ), .dinb(\a[6] ), .dout(n5199));
  jand g05008(.dina(n5199), .dinb(n5195), .dout(n5200));
  jand g05009(.dina(n3138), .dinb(n976), .dout(n5201));
  jor  g05010(.dina(n5201), .dinb(n5200), .dout(n5202));
  jand g05011(.dina(n5202), .dinb(n5198), .dout(n5203));
  jnot g05012(.din(n5203), .dout(n5204));
  jand g05013(.dina(n5204), .dinb(n5195), .dout(n5205));
  jand g05014(.dina(\a[37] ), .dinb(\a[14] ), .dout(n5206));
  jor  g05015(.dina(n5206), .dinb(n5199), .dout(n5207));
  jor  g05016(.dina(n5202), .dinb(n5197), .dout(n5208));
  jnot g05017(.din(n5208), .dout(n5209));
  jand g05018(.dina(n5209), .dinb(n5207), .dout(n5210));
  jor  g05019(.dina(n5210), .dinb(n5205), .dout(n5211));
  jand g05020(.dina(\a[33] ), .dinb(\a[18] ), .dout(n5212));
  jand g05021(.dina(\a[46] ), .dinb(\a[5] ), .dout(n5213));
  jand g05022(.dina(\a[35] ), .dinb(\a[16] ), .dout(n5214));
  jxor g05023(.dina(n5214), .dinb(n5213), .dout(n5215));
  jxor g05024(.dina(n5215), .dinb(n5212), .dout(n5216));
  jnot g05025(.din(n5216), .dout(n5217));
  jand g05026(.dina(\a[30] ), .dinb(\a[21] ), .dout(n5218));
  jnot g05027(.din(n5218), .dout(n5219));
  jand g05028(.dina(n2653), .dinb(n1658), .dout(n5220));
  jnot g05029(.din(n5220), .dout(n5221));
  jand g05030(.dina(\a[29] ), .dinb(\a[22] ), .dout(n5222));
  jand g05031(.dina(\a[28] ), .dinb(\a[23] ), .dout(n5223));
  jor  g05032(.dina(n5223), .dinb(n5222), .dout(n5224));
  jand g05033(.dina(n5224), .dinb(n5221), .dout(n5225));
  jxor g05034(.dina(n5225), .dinb(n5219), .dout(n5226));
  jxor g05035(.dina(n5226), .dinb(n5217), .dout(n5227));
  jxor g05036(.dina(n5227), .dinb(n5211), .dout(n5228));
  jand g05037(.dina(\a[43] ), .dinb(\a[8] ), .dout(n5229));
  jand g05038(.dina(\a[38] ), .dinb(\a[13] ), .dout(n5230));
  jand g05039(.dina(n5230), .dinb(n5229), .dout(n5231));
  jnot g05040(.din(n5231), .dout(n5232));
  jand g05041(.dina(n4495), .dinb(n499), .dout(n5233));
  jand g05042(.dina(\a[44] ), .dinb(\a[7] ), .dout(n5234));
  jand g05043(.dina(n5234), .dinb(n5230), .dout(n5235));
  jor  g05044(.dina(n5235), .dinb(n5233), .dout(n5236));
  jnot g05045(.din(n5236), .dout(n5237));
  jand g05046(.dina(n5237), .dinb(n5232), .dout(n5238));
  jor  g05047(.dina(n5230), .dinb(n5229), .dout(n5239));
  jand g05048(.dina(n5239), .dinb(n5238), .dout(n5240));
  jand g05049(.dina(n5236), .dinb(n5232), .dout(n5241));
  jnot g05050(.din(n5241), .dout(n5242));
  jand g05051(.dina(n5242), .dinb(n5234), .dout(n5243));
  jor  g05052(.dina(n5243), .dinb(n5240), .dout(n5244));
  jand g05053(.dina(\a[42] ), .dinb(\a[9] ), .dout(n5245));
  jand g05054(.dina(\a[41] ), .dinb(\a[39] ), .dout(n5246));
  jand g05055(.dina(n5246), .dinb(n1151), .dout(n5247));
  jnot g05056(.din(n5247), .dout(n5248));
  jand g05057(.dina(\a[39] ), .dinb(\a[12] ), .dout(n5249));
  jand g05058(.dina(n5249), .dinb(n5245), .dout(n5250));
  jand g05059(.dina(n4514), .dinb(n453), .dout(n5251));
  jor  g05060(.dina(n5251), .dinb(n5250), .dout(n5252));
  jand g05061(.dina(n5252), .dinb(n5248), .dout(n5253));
  jnot g05062(.din(n5253), .dout(n5254));
  jand g05063(.dina(n5254), .dinb(n5245), .dout(n5255));
  jor  g05064(.dina(n5252), .dinb(n5247), .dout(n5256));
  jnot g05065(.din(n5256), .dout(n5257));
  jand g05066(.dina(\a[41] ), .dinb(\a[10] ), .dout(n5258));
  jor  g05067(.dina(n5258), .dinb(n5249), .dout(n5259));
  jand g05068(.dina(n5259), .dinb(n5257), .dout(n5260));
  jor  g05069(.dina(n5260), .dinb(n5255), .dout(n5261));
  jxor g05070(.dina(n5261), .dinb(n5244), .dout(n5262));
  jand g05071(.dina(\a[40] ), .dinb(\a[11] ), .dout(n5263));
  jnot g05072(.din(n5263), .dout(n5264));
  jand g05073(.dina(n1927), .dinb(n1648), .dout(n5265));
  jnot g05074(.din(n5265), .dout(n5266));
  jand g05075(.dina(\a[27] ), .dinb(\a[24] ), .dout(n5267));
  jor  g05076(.dina(n5267), .dinb(n2128), .dout(n5268));
  jand g05077(.dina(n5268), .dinb(n5266), .dout(n5269));
  jxor g05078(.dina(n5269), .dinb(n5264), .dout(n5270));
  jnot g05079(.din(n5270), .dout(n5271));
  jxor g05080(.dina(n5271), .dinb(n5262), .dout(n5272));
  jxor g05081(.dina(n5272), .dinb(n5228), .dout(n5273));
  jxor g05082(.dina(n5273), .dinb(n5194), .dout(n5274));
  jxor g05083(.dina(n5274), .dinb(n5173), .dout(n5275));
  jxor g05084(.dina(n5275), .dinb(n5170), .dout(n5276));
  jxor g05085(.dina(n5276), .dinb(n5167), .dout(n5277));
  jand g05086(.dina(n5080), .dinb(n4978), .dout(n5278));
  jand g05087(.dina(n5081), .dinb(n4973), .dout(n5279));
  jor  g05088(.dina(n5279), .dinb(n5278), .dout(n5280));
  jand g05089(.dina(n5141), .dinb(n5138), .dout(n5281));
  jand g05090(.dina(n5145), .dinb(n5142), .dout(n5282));
  jor  g05091(.dina(n5282), .dinb(n5281), .dout(n5283));
  jand g05092(.dina(n5117), .dinb(n5114), .dout(n5284));
  jand g05093(.dina(n5128), .dinb(n5118), .dout(n5285));
  jor  g05094(.dina(n5285), .dinb(n5284), .dout(n5286));
  jxor g05095(.dina(n5286), .dinb(n5283), .dout(n5287));
  jand g05096(.dina(n5105), .dinb(n5103), .dout(n5288));
  jand g05097(.dina(n5106), .dinb(n4795), .dout(n5289));
  jor  g05098(.dina(n5289), .dinb(n5288), .dout(n5290));
  jand g05099(.dina(n5123), .dinb(n5121), .dout(n5291));
  jand g05100(.dina(n5127), .dinb(n5124), .dout(n5292));
  jor  g05101(.dina(n5292), .dinb(n5291), .dout(n5293));
  jxor g05102(.dina(n5293), .dinb(n5290), .dout(n5294));
  jnot g05103(.din(n5294), .dout(n5295));
  jand g05104(.dina(n5032), .dinb(n5023), .dout(n5296));
  jnot g05105(.din(n5296), .dout(n5297));
  jor  g05106(.dina(n5043), .dinb(n5034), .dout(n5298));
  jand g05107(.dina(n5298), .dinb(n5297), .dout(n5299));
  jxor g05108(.dina(n5299), .dinb(n5295), .dout(n5300));
  jxor g05109(.dina(n5300), .dinb(n5287), .dout(n5301));
  jxor g05110(.dina(n5301), .dinb(n5280), .dout(n5302));
  jand g05111(.dina(n5078), .dinb(n5044), .dout(n5303));
  jand g05112(.dina(n5079), .dinb(n5006), .dout(n5304));
  jor  g05113(.dina(n5304), .dinb(n5303), .dout(n5305));
  jand g05114(.dina(n5004), .dinb(n4999), .dout(n5306));
  jand g05115(.dina(n5005), .dinb(n4982), .dout(n5307));
  jor  g05116(.dina(n5307), .dinb(n5306), .dout(n5308));
  jnot g05117(.din(n4992), .dout(n5309));
  jand g05118(.dina(n5072), .dinb(n5070), .dout(n5310));
  jnot g05119(.din(n5310), .dout(n5311));
  jand g05120(.dina(n5311), .dinb(n5075), .dout(n5312));
  jxor g05121(.dina(n5312), .dinb(n5309), .dout(n5313));
  jand g05122(.dina(\a[49] ), .dinb(\a[2] ), .dout(n5314));
  jnot g05123(.din(n5314), .dout(n5315));
  jand g05124(.dina(\a[48] ), .dinb(\a[47] ), .dout(n5316));
  jand g05125(.dina(n5316), .dinb(n265), .dout(n5317));
  jnot g05126(.din(n5317), .dout(n5318));
  jand g05127(.dina(\a[48] ), .dinb(\a[3] ), .dout(n5319));
  jor  g05128(.dina(n5319), .dinb(n5010), .dout(n5320));
  jand g05129(.dina(n5320), .dinb(n5318), .dout(n5321));
  jxor g05130(.dina(n5321), .dinb(n5315), .dout(n5322));
  jnot g05131(.din(n5322), .dout(n5323));
  jxor g05132(.dina(n5323), .dinb(n5313), .dout(n5324));
  jxor g05133(.dina(n5324), .dinb(n5308), .dout(n5325));
  jand g05134(.dina(n5101), .dinb(n5098), .dout(n5326));
  jand g05135(.dina(n5107), .dinb(n5102), .dout(n5327));
  jor  g05136(.dina(n5327), .dinb(n5326), .dout(n5328));
  jxor g05137(.dina(n5328), .dinb(n5325), .dout(n5329));
  jxor g05138(.dina(n5329), .dinb(n5305), .dout(n5330));
  jand g05139(.dina(n5064), .dinb(n5063), .dout(n5331));
  jand g05140(.dina(n5065), .dinb(n5062), .dout(n5332));
  jor  g05141(.dina(n5332), .dinb(n5331), .dout(n5333));
  jxor g05142(.dina(n5333), .dinb(n5056), .dout(n5334));
  jor  g05143(.dina(n5002), .dinb(n5001), .dout(n5335));
  jand g05144(.dina(n5002), .dinb(n5001), .dout(n5336));
  jor  g05145(.dina(n5336), .dinb(n5000), .dout(n5337));
  jand g05146(.dina(n5337), .dinb(n5335), .dout(n5338));
  jxor g05147(.dina(n5338), .dinb(n5334), .dout(n5339));
  jnot g05148(.din(n5339), .dout(n5340));
  jand g05149(.dina(n5066), .dinb(n5061), .dout(n5341));
  jnot g05150(.din(n5341), .dout(n5342));
  jor  g05151(.dina(n5077), .dinb(n5068), .dout(n5343));
  jand g05152(.dina(n5343), .dinb(n5342), .dout(n5344));
  jxor g05153(.dina(n5344), .dinb(n5340), .dout(n5345));
  jand g05154(.dina(n5031), .dinb(n5024), .dout(n5346));
  jor  g05155(.dina(n5346), .dinb(n5029), .dout(n5347));
  jand g05156(.dina(n5038), .dinb(n5036), .dout(n5348));
  jnot g05157(.din(n5348), .dout(n5349));
  jand g05158(.dina(n5349), .dinb(n5041), .dout(n5350));
  jxor g05159(.dina(n5350), .dinb(n5018), .dout(n5351));
  jxor g05160(.dina(n5351), .dinb(n5347), .dout(n5352));
  jxor g05161(.dina(n5352), .dinb(n5345), .dout(n5353));
  jxor g05162(.dina(n5353), .dinb(n5330), .dout(n5354));
  jxor g05163(.dina(n5354), .dinb(n5302), .dout(n5355));
  jxor g05164(.dina(n5355), .dinb(n5277), .dout(n5356));
  jand g05165(.dina(n5356), .dinb(n5164), .dout(n5357));
  jor  g05166(.dina(n5356), .dinb(n5164), .dout(n5358));
  jnot g05167(.din(n5358), .dout(n5359));
  jor  g05168(.dina(n5359), .dinb(n5357), .dout(n5360));
  jand g05169(.dina(n5153), .dinb(n4966), .dout(n5361));
  jnot g05170(.din(n5361), .dout(n5362));
  jnot g05171(.din(n5153), .dout(n5363));
  jand g05172(.dina(n5363), .dinb(n4967), .dout(n5364));
  jor  g05173(.dina(n5160), .dinb(n5364), .dout(n5365));
  jand g05174(.dina(n5365), .dinb(n5362), .dout(n5366));
  jxor g05175(.dina(n5366), .dinb(n5360), .dout(\asquared[52] ));
  jand g05176(.dina(n5276), .dinb(n5167), .dout(n5368));
  jand g05177(.dina(n5355), .dinb(n5277), .dout(n5369));
  jor  g05178(.dina(n5369), .dinb(n5368), .dout(n5370));
  jand g05179(.dina(n5329), .dinb(n5305), .dout(n5371));
  jand g05180(.dina(n5353), .dinb(n5330), .dout(n5372));
  jor  g05181(.dina(n5372), .dinb(n5371), .dout(n5373));
  jand g05182(.dina(n5286), .dinb(n5283), .dout(n5374));
  jand g05183(.dina(n5300), .dinb(n5287), .dout(n5375));
  jor  g05184(.dina(n5375), .dinb(n5374), .dout(n5376));
  jor  g05185(.dina(n5344), .dinb(n5340), .dout(n5377));
  jand g05186(.dina(n5352), .dinb(n5345), .dout(n5378));
  jnot g05187(.din(n5378), .dout(n5379));
  jand g05188(.dina(n5379), .dinb(n5377), .dout(n5380));
  jnot g05189(.din(n5380), .dout(n5381));
  jand g05190(.dina(\a[46] ), .dinb(\a[36] ), .dout(n5382));
  jand g05191(.dina(n5382), .dinb(n1131), .dout(n5383));
  jnot g05192(.din(n5383), .dout(n5384));
  jand g05193(.dina(\a[47] ), .dinb(\a[6] ), .dout(n5385));
  jand g05194(.dina(n5385), .dinb(n5213), .dout(n5386));
  jand g05195(.dina(\a[36] ), .dinb(\a[16] ), .dout(n5387));
  jand g05196(.dina(\a[47] ), .dinb(\a[5] ), .dout(n5388));
  jand g05197(.dina(n5388), .dinb(n5387), .dout(n5389));
  jor  g05198(.dina(n5389), .dinb(n5386), .dout(n5390));
  jnot g05199(.din(n5390), .dout(n5391));
  jand g05200(.dina(n5391), .dinb(n5384), .dout(n5392));
  jand g05201(.dina(\a[46] ), .dinb(\a[6] ), .dout(n5393));
  jor  g05202(.dina(n5393), .dinb(n5387), .dout(n5394));
  jand g05203(.dina(n5394), .dinb(n5392), .dout(n5395));
  jand g05204(.dina(n5390), .dinb(n5384), .dout(n5396));
  jnot g05205(.din(n5396), .dout(n5397));
  jand g05206(.dina(n5397), .dinb(n5388), .dout(n5398));
  jor  g05207(.dina(n5398), .dinb(n5395), .dout(n5399));
  jand g05208(.dina(\a[42] ), .dinb(\a[10] ), .dout(n5400));
  jnot g05209(.din(n5400), .dout(n5401));
  jand g05210(.dina(n4632), .dinb(n555), .dout(n5402));
  jnot g05211(.din(n5402), .dout(n5403));
  jand g05212(.dina(\a[40] ), .dinb(\a[12] ), .dout(n5404));
  jand g05213(.dina(\a[41] ), .dinb(\a[11] ), .dout(n5405));
  jor  g05214(.dina(n5405), .dinb(n5404), .dout(n5406));
  jand g05215(.dina(n5406), .dinb(n5403), .dout(n5407));
  jxor g05216(.dina(n5407), .dinb(n5401), .dout(n5408));
  jnot g05217(.din(n5408), .dout(n5409));
  jxor g05218(.dina(n5409), .dinb(n5399), .dout(n5410));
  jnot g05219(.din(n5410), .dout(n5411));
  jand g05220(.dina(\a[37] ), .dinb(\a[15] ), .dout(n5412));
  jnot g05221(.din(n5412), .dout(n5413));
  jand g05222(.dina(n4812), .dinb(n499), .dout(n5414));
  jnot g05223(.din(n5414), .dout(n5415));
  jand g05224(.dina(\a[45] ), .dinb(\a[7] ), .dout(n5416));
  jand g05225(.dina(\a[44] ), .dinb(\a[8] ), .dout(n5417));
  jor  g05226(.dina(n5417), .dinb(n5416), .dout(n5418));
  jand g05227(.dina(n5418), .dinb(n5415), .dout(n5419));
  jxor g05228(.dina(n5419), .dinb(n5413), .dout(n5420));
  jxor g05229(.dina(n5420), .dinb(n5411), .dout(n5421));
  jand g05230(.dina(\a[38] ), .dinb(\a[14] ), .dout(n5422));
  jand g05231(.dina(\a[39] ), .dinb(\a[13] ), .dout(n5423));
  jand g05232(.dina(\a[43] ), .dinb(\a[9] ), .dout(n5424));
  jand g05233(.dina(n5424), .dinb(n5423), .dout(n5425));
  jnot g05234(.din(n5425), .dout(n5426));
  jand g05235(.dina(n5424), .dinb(n5422), .dout(n5427));
  jand g05236(.dina(\a[39] ), .dinb(\a[14] ), .dout(n5428));
  jand g05237(.dina(n5428), .dinb(n5230), .dout(n5429));
  jor  g05238(.dina(n5429), .dinb(n5427), .dout(n5430));
  jand g05239(.dina(n5430), .dinb(n5426), .dout(n5431));
  jnot g05240(.din(n5431), .dout(n5432));
  jand g05241(.dina(n5432), .dinb(n5422), .dout(n5433));
  jor  g05242(.dina(n5430), .dinb(n5425), .dout(n5434));
  jnot g05243(.din(n5434), .dout(n5435));
  jor  g05244(.dina(n5424), .dinb(n5423), .dout(n5436));
  jand g05245(.dina(n5436), .dinb(n5435), .dout(n5437));
  jor  g05246(.dina(n5437), .dinb(n5433), .dout(n5438));
  jand g05247(.dina(\a[34] ), .dinb(\a[18] ), .dout(n5439));
  jand g05248(.dina(n3269), .dinb(n1490), .dout(n5440));
  jnot g05249(.din(n5440), .dout(n5441));
  jand g05250(.dina(\a[31] ), .dinb(\a[21] ), .dout(n5442));
  jand g05251(.dina(\a[32] ), .dinb(\a[20] ), .dout(n5443));
  jor  g05252(.dina(n5443), .dinb(n5442), .dout(n5444));
  jand g05253(.dina(n5444), .dinb(n5441), .dout(n5445));
  jxor g05254(.dina(n5445), .dinb(n5439), .dout(n5446));
  jnot g05255(.din(n5446), .dout(n5447));
  jand g05256(.dina(\a[30] ), .dinb(\a[22] ), .dout(n5448));
  jnot g05257(.din(n5448), .dout(n5449));
  jand g05258(.dina(n2653), .dinb(n1942), .dout(n5450));
  jnot g05259(.din(n5450), .dout(n5451));
  jand g05260(.dina(\a[29] ), .dinb(\a[23] ), .dout(n5452));
  jand g05261(.dina(\a[28] ), .dinb(\a[24] ), .dout(n5453));
  jor  g05262(.dina(n5453), .dinb(n5452), .dout(n5454));
  jand g05263(.dina(n5454), .dinb(n5451), .dout(n5455));
  jxor g05264(.dina(n5455), .dinb(n5449), .dout(n5456));
  jxor g05265(.dina(n5456), .dinb(n5447), .dout(n5457));
  jxor g05266(.dina(n5457), .dinb(n5438), .dout(n5458));
  jxor g05267(.dina(n5458), .dinb(n5421), .dout(n5459));
  jxor g05268(.dina(n5459), .dinb(n5381), .dout(n5460));
  jxor g05269(.dina(n5460), .dinb(n5376), .dout(n5461));
  jxor g05270(.dina(n5461), .dinb(n5373), .dout(n5462));
  jand g05271(.dina(n5301), .dinb(n5280), .dout(n5463));
  jand g05272(.dina(n5354), .dinb(n5302), .dout(n5464));
  jor  g05273(.dina(n5464), .dinb(n5463), .dout(n5465));
  jxor g05274(.dina(n5465), .dinb(n5462), .dout(n5466));
  jand g05275(.dina(n5274), .dinb(n5173), .dout(n5467));
  jand g05276(.dina(n5275), .dinb(n5170), .dout(n5468));
  jor  g05277(.dina(n5468), .dinb(n5467), .dout(n5469));
  jand g05278(.dina(n5333), .dinb(n5056), .dout(n5470));
  jand g05279(.dina(n5338), .dinb(n5334), .dout(n5471));
  jor  g05280(.dina(n5471), .dinb(n5470), .dout(n5472));
  jand g05281(.dina(n5350), .dinb(n5018), .dout(n5473));
  jand g05282(.dina(n5351), .dinb(n5347), .dout(n5474));
  jor  g05283(.dina(n5474), .dinb(n5473), .dout(n5475));
  jand g05284(.dina(\a[33] ), .dinb(\a[19] ), .dout(n5476));
  jand g05285(.dina(\a[50] ), .dinb(\a[3] ), .dout(n5477));
  jand g05286(.dina(n5477), .dinb(n5314), .dout(n5478));
  jnot g05287(.din(n5478), .dout(n5479));
  jand g05288(.dina(\a[49] ), .dinb(\a[3] ), .dout(n5480));
  jor  g05289(.dina(n5480), .dinb(n5028), .dout(n5481));
  jand g05290(.dina(n5481), .dinb(n5479), .dout(n5482));
  jxor g05291(.dina(n5482), .dinb(n5476), .dout(n5483));
  jxor g05292(.dina(n5483), .dinb(n5475), .dout(n5484));
  jxor g05293(.dina(n5484), .dinb(n5472), .dout(n5485));
  jand g05294(.dina(n5324), .dinb(n5308), .dout(n5486));
  jand g05295(.dina(n5328), .dinb(n5325), .dout(n5487));
  jor  g05296(.dina(n5487), .dinb(n5486), .dout(n5488));
  jxor g05297(.dina(n5488), .dinb(n5485), .dout(n5489));
  jand g05298(.dina(n5261), .dinb(n5244), .dout(n5490));
  jand g05299(.dina(n5271), .dinb(n5262), .dout(n5491));
  jor  g05300(.dina(n5491), .dinb(n5490), .dout(n5492));
  jand g05301(.dina(n5312), .dinb(n5309), .dout(n5493));
  jand g05302(.dina(n5323), .dinb(n5313), .dout(n5494));
  jor  g05303(.dina(n5494), .dinb(n5493), .dout(n5495));
  jand g05304(.dina(n5180), .dinb(\a[26] ), .dout(n5496));
  jand g05305(.dina(\a[51] ), .dinb(\a[1] ), .dout(n5497));
  jxor g05306(.dina(n5497), .dinb(n2259), .dout(n5498));
  jxor g05307(.dina(n5498), .dinb(n5496), .dout(n5499));
  jand g05308(.dina(n5266), .dinb(n5264), .dout(n5500));
  jnot g05309(.din(n5500), .dout(n5501));
  jand g05310(.dina(n5501), .dinb(n5268), .dout(n5502));
  jxor g05311(.dina(n5502), .dinb(n5499), .dout(n5503));
  jxor g05312(.dina(n5503), .dinb(n5495), .dout(n5504));
  jxor g05313(.dina(n5504), .dinb(n5492), .dout(n5505));
  jxor g05314(.dina(n5505), .dinb(n5489), .dout(n5506));
  jxor g05315(.dina(n5506), .dinb(n5469), .dout(n5507));
  jor  g05316(.dina(n5192), .dinb(n5183), .dout(n5508));
  jand g05317(.dina(n5193), .dinb(n5176), .dout(n5509));
  jnot g05318(.din(n5509), .dout(n5510));
  jand g05319(.dina(n5510), .dinb(n5508), .dout(n5511));
  jnot g05320(.din(n5511), .dout(n5512));
  jand g05321(.dina(n5178), .dinb(n5177), .dout(n5513));
  jand g05322(.dina(n5181), .dinb(n5179), .dout(n5514));
  jor  g05323(.dina(n5514), .dinb(n5513), .dout(n5515));
  jxor g05324(.dina(n5515), .dinb(n5256), .dout(n5516));
  jand g05325(.dina(\a[48] ), .dinb(\a[4] ), .dout(n5517));
  jand g05326(.dina(\a[35] ), .dinb(\a[17] ), .dout(n5518));
  jand g05327(.dina(n5518), .dinb(n5517), .dout(n5519));
  jnot g05328(.din(n5519), .dout(n5520));
  jand g05329(.dina(n711), .dinb(\a[35] ), .dout(n5521));
  jand g05330(.dina(n5521), .dinb(\a[52] ), .dout(n5522));
  jand g05331(.dina(\a[52] ), .dinb(\a[0] ), .dout(n5523));
  jand g05332(.dina(n5523), .dinb(n5517), .dout(n5524));
  jor  g05333(.dina(n5524), .dinb(n5522), .dout(n5525));
  jnot g05334(.din(n5525), .dout(n5526));
  jand g05335(.dina(n5526), .dinb(n5520), .dout(n5527));
  jor  g05336(.dina(n5518), .dinb(n5517), .dout(n5528));
  jand g05337(.dina(n5528), .dinb(n5527), .dout(n5529));
  jand g05338(.dina(n5525), .dinb(n5520), .dout(n5530));
  jnot g05339(.din(n5530), .dout(n5531));
  jand g05340(.dina(n5531), .dinb(n5523), .dout(n5532));
  jor  g05341(.dina(n5532), .dinb(n5529), .dout(n5533));
  jxor g05342(.dina(n5533), .dinb(n5516), .dout(n5534));
  jxor g05343(.dina(n5534), .dinb(n5512), .dout(n5535));
  jnot g05344(.din(n5535), .dout(n5536));
  jand g05345(.dina(n5293), .dinb(n5290), .dout(n5537));
  jnot g05346(.din(n5537), .dout(n5538));
  jor  g05347(.dina(n5299), .dinb(n5295), .dout(n5539));
  jand g05348(.dina(n5539), .dinb(n5538), .dout(n5540));
  jxor g05349(.dina(n5540), .dinb(n5536), .dout(n5541));
  jand g05350(.dina(n5272), .dinb(n5228), .dout(n5542));
  jand g05351(.dina(n5273), .dinb(n5194), .dout(n5543));
  jor  g05352(.dina(n5543), .dinb(n5542), .dout(n5544));
  jnot g05353(.din(n5238), .dout(n5545));
  jand g05354(.dina(n5214), .dinb(n5213), .dout(n5546));
  jand g05355(.dina(n5215), .dinb(n5212), .dout(n5547));
  jor  g05356(.dina(n5547), .dinb(n5546), .dout(n5548));
  jxor g05357(.dina(n5548), .dinb(n5545), .dout(n5549));
  jand g05358(.dina(n5221), .dinb(n5219), .dout(n5550));
  jnot g05359(.din(n5550), .dout(n5551));
  jand g05360(.dina(n5551), .dinb(n5224), .dout(n5552));
  jxor g05361(.dina(n5552), .dinb(n5549), .dout(n5553));
  jand g05362(.dina(n5187), .dinb(n5185), .dout(n5554));
  jnot g05363(.din(n5554), .dout(n5555));
  jand g05364(.dina(n5555), .dinb(n5190), .dout(n5556));
  jand g05365(.dina(n5318), .dinb(n5315), .dout(n5557));
  jnot g05366(.din(n5557), .dout(n5558));
  jand g05367(.dina(n5558), .dinb(n5320), .dout(n5559));
  jxor g05368(.dina(n5559), .dinb(n5556), .dout(n5560));
  jxor g05369(.dina(n5560), .dinb(n5208), .dout(n5561));
  jnot g05370(.din(n5561), .dout(n5562));
  jor  g05371(.dina(n5226), .dinb(n5217), .dout(n5563));
  jand g05372(.dina(n5227), .dinb(n5211), .dout(n5564));
  jnot g05373(.din(n5564), .dout(n5565));
  jand g05374(.dina(n5565), .dinb(n5563), .dout(n5566));
  jxor g05375(.dina(n5566), .dinb(n5562), .dout(n5567));
  jxor g05376(.dina(n5567), .dinb(n5553), .dout(n5568));
  jxor g05377(.dina(n5568), .dinb(n5544), .dout(n5569));
  jxor g05378(.dina(n5569), .dinb(n5541), .dout(n5570));
  jxor g05379(.dina(n5570), .dinb(n5507), .dout(n5571));
  jxor g05380(.dina(n5571), .dinb(n5466), .dout(n5572));
  jnot g05381(.din(n5572), .dout(n5573));
  jxor g05382(.dina(n5573), .dinb(n5370), .dout(n5574));
  jnot g05383(.din(n5357), .dout(n5575));
  jor  g05384(.dina(n5366), .dinb(n5359), .dout(n5576));
  jand g05385(.dina(n5576), .dinb(n5575), .dout(n5577));
  jxor g05386(.dina(n5577), .dinb(n5574), .dout(\asquared[53] ));
  jand g05387(.dina(n5465), .dinb(n5462), .dout(n5579));
  jand g05388(.dina(n5571), .dinb(n5466), .dout(n5580));
  jor  g05389(.dina(n5580), .dinb(n5579), .dout(n5581));
  jand g05390(.dina(n5506), .dinb(n5469), .dout(n5582));
  jand g05391(.dina(n5570), .dinb(n5507), .dout(n5583));
  jor  g05392(.dina(n5583), .dinb(n5582), .dout(n5584));
  jand g05393(.dina(n5568), .dinb(n5544), .dout(n5585));
  jand g05394(.dina(n5569), .dinb(n5541), .dout(n5586));
  jor  g05395(.dina(n5586), .dinb(n5585), .dout(n5587));
  jand g05396(.dina(n5483), .dinb(n5475), .dout(n5588));
  jand g05397(.dina(n5484), .dinb(n5472), .dout(n5589));
  jor  g05398(.dina(n5589), .dinb(n5588), .dout(n5590));
  jand g05399(.dina(n5497), .dinb(n2259), .dout(n5591));
  jand g05400(.dina(\a[51] ), .dinb(\a[2] ), .dout(n5592));
  jor  g05401(.dina(n5592), .dinb(n5477), .dout(n5593));
  jand g05402(.dina(\a[51] ), .dinb(\a[50] ), .dout(n5594));
  jand g05403(.dina(n5594), .dinb(n248), .dout(n5595));
  jnot g05404(.din(n5595), .dout(n5596));
  jand g05405(.dina(n5596), .dinb(n5593), .dout(n5597));
  jxor g05406(.dina(n5597), .dinb(n5591), .dout(n5598));
  jand g05407(.dina(\a[49] ), .dinb(\a[4] ), .dout(n5599));
  jand g05408(.dina(n3243), .dinb(n1107), .dout(n5600));
  jnot g05409(.din(n5600), .dout(n5601));
  jand g05410(.dina(\a[36] ), .dinb(\a[17] ), .dout(n5602));
  jand g05411(.dina(\a[35] ), .dinb(\a[18] ), .dout(n5603));
  jor  g05412(.dina(n5603), .dinb(n5602), .dout(n5604));
  jand g05413(.dina(n5604), .dinb(n5601), .dout(n5605));
  jxor g05414(.dina(n5605), .dinb(n5599), .dout(n5606));
  jxor g05415(.dina(n5606), .dinb(n5598), .dout(n5607));
  jnot g05416(.din(n5607), .dout(n5608));
  jand g05417(.dina(\a[34] ), .dinb(\a[19] ), .dout(n5609));
  jnot g05418(.din(n5609), .dout(n5610));
  jand g05419(.dina(n2671), .dinb(n1490), .dout(n5611));
  jnot g05420(.din(n5611), .dout(n5612));
  jand g05421(.dina(\a[33] ), .dinb(\a[20] ), .dout(n5613));
  jand g05422(.dina(\a[32] ), .dinb(\a[21] ), .dout(n5614));
  jor  g05423(.dina(n5614), .dinb(n5613), .dout(n5615));
  jand g05424(.dina(n5615), .dinb(n5612), .dout(n5616));
  jxor g05425(.dina(n5616), .dinb(n5610), .dout(n5617));
  jxor g05426(.dina(n5617), .dinb(n5608), .dout(n5618));
  jxor g05427(.dina(n5618), .dinb(n5590), .dout(n5619));
  jand g05428(.dina(\a[46] ), .dinb(\a[7] ), .dout(n5620));
  jand g05429(.dina(\a[38] ), .dinb(\a[15] ), .dout(n5621));
  jand g05430(.dina(n5621), .dinb(n5620), .dout(n5622));
  jnot g05431(.din(n5622), .dout(n5623));
  jand g05432(.dina(\a[47] ), .dinb(\a[7] ), .dout(n5624));
  jand g05433(.dina(n5624), .dinb(n5393), .dout(n5625));
  jand g05434(.dina(n5621), .dinb(n5385), .dout(n5626));
  jor  g05435(.dina(n5626), .dinb(n5625), .dout(n5627));
  jnot g05436(.din(n5627), .dout(n5628));
  jand g05437(.dina(n5628), .dinb(n5623), .dout(n5629));
  jor  g05438(.dina(n5621), .dinb(n5620), .dout(n5630));
  jand g05439(.dina(n5630), .dinb(n5629), .dout(n5631));
  jand g05440(.dina(n5627), .dinb(n5623), .dout(n5632));
  jnot g05441(.din(n5632), .dout(n5633));
  jand g05442(.dina(n5633), .dinb(n5385), .dout(n5634));
  jor  g05443(.dina(n5634), .dinb(n5631), .dout(n5635));
  jand g05444(.dina(\a[44] ), .dinb(\a[9] ), .dout(n5636));
  jand g05445(.dina(n5636), .dinb(n5428), .dout(n5637));
  jnot g05446(.din(n5637), .dout(n5638));
  jand g05447(.dina(n4812), .dinb(n395), .dout(n5639));
  jand g05448(.dina(\a[45] ), .dinb(\a[8] ), .dout(n5640));
  jand g05449(.dina(n5640), .dinb(n5428), .dout(n5641));
  jor  g05450(.dina(n5641), .dinb(n5639), .dout(n5642));
  jnot g05451(.din(n5642), .dout(n5643));
  jand g05452(.dina(n5643), .dinb(n5638), .dout(n5644));
  jor  g05453(.dina(n5636), .dinb(n5428), .dout(n5645));
  jand g05454(.dina(n5645), .dinb(n5644), .dout(n5646));
  jand g05455(.dina(n5642), .dinb(n5638), .dout(n5647));
  jnot g05456(.din(n5647), .dout(n5648));
  jand g05457(.dina(n5648), .dinb(n5640), .dout(n5649));
  jor  g05458(.dina(n5649), .dinb(n5646), .dout(n5650));
  jxor g05459(.dina(n5650), .dinb(n5635), .dout(n5651));
  jand g05460(.dina(\a[53] ), .dinb(\a[0] ), .dout(n5652));
  jand g05461(.dina(\a[48] ), .dinb(\a[5] ), .dout(n5653));
  jand g05462(.dina(\a[37] ), .dinb(\a[16] ), .dout(n5654));
  jxor g05463(.dina(n5654), .dinb(n5653), .dout(n5655));
  jxor g05464(.dina(n5655), .dinb(n5652), .dout(n5656));
  jxor g05465(.dina(n5656), .dinb(n5651), .dout(n5657));
  jxor g05466(.dina(n5657), .dinb(n5619), .dout(n5658));
  jand g05467(.dina(n5503), .dinb(n5495), .dout(n5659));
  jand g05468(.dina(n5504), .dinb(n5492), .dout(n5660));
  jor  g05469(.dina(n5660), .dinb(n5659), .dout(n5661));
  jand g05470(.dina(\a[43] ), .dinb(\a[10] ), .dout(n5662));
  jand g05471(.dina(\a[41] ), .dinb(\a[12] ), .dout(n5663));
  jor  g05472(.dina(n5663), .dinb(n5662), .dout(n5664));
  jand g05473(.dina(n4115), .dinb(n1151), .dout(n5665));
  jnot g05474(.din(n5665), .dout(n5666));
  jand g05475(.dina(\a[40] ), .dinb(\a[13] ), .dout(n5667));
  jand g05476(.dina(n5667), .dinb(n5662), .dout(n5668));
  jand g05477(.dina(n4632), .dinb(n899), .dout(n5669));
  jor  g05478(.dina(n5669), .dinb(n5668), .dout(n5670));
  jnot g05479(.din(n5670), .dout(n5671));
  jand g05480(.dina(n5671), .dinb(n5666), .dout(n5672));
  jand g05481(.dina(n5672), .dinb(n5664), .dout(n5673));
  jand g05482(.dina(n5670), .dinb(n5666), .dout(n5674));
  jnot g05483(.din(n5674), .dout(n5675));
  jand g05484(.dina(n5675), .dinb(n5667), .dout(n5676));
  jor  g05485(.dina(n5676), .dinb(n5673), .dout(n5677));
  jnot g05486(.din(n1989), .dout(n5678));
  jand g05487(.dina(n3294), .dinb(n1942), .dout(n5679));
  jnot g05488(.din(n5679), .dout(n5680));
  jand g05489(.dina(\a[29] ), .dinb(\a[24] ), .dout(n5681));
  jand g05490(.dina(\a[30] ), .dinb(\a[23] ), .dout(n5682));
  jor  g05491(.dina(n5682), .dinb(n5681), .dout(n5683));
  jand g05492(.dina(n5683), .dinb(n5680), .dout(n5684));
  jxor g05493(.dina(n5684), .dinb(n5678), .dout(n5685));
  jnot g05494(.din(n5685), .dout(n5686));
  jxor g05495(.dina(n5686), .dinb(n5677), .dout(n5687));
  jnot g05496(.din(n5687), .dout(n5688));
  jand g05497(.dina(\a[42] ), .dinb(\a[11] ), .dout(n5689));
  jnot g05498(.din(n5689), .dout(n5690));
  jand g05499(.dina(n2128), .dinb(n2042), .dout(n5691));
  jnot g05500(.din(n5691), .dout(n5692));
  jand g05501(.dina(\a[28] ), .dinb(\a[25] ), .dout(n5693));
  jor  g05502(.dina(n5693), .dinb(n1927), .dout(n5694));
  jand g05503(.dina(n5694), .dinb(n5692), .dout(n5695));
  jxor g05504(.dina(n5695), .dinb(n5690), .dout(n5696));
  jxor g05505(.dina(n5696), .dinb(n5688), .dout(n5697));
  jxor g05506(.dina(n5697), .dinb(n5661), .dout(n5698));
  jnot g05507(.din(n5698), .dout(n5699));
  jor  g05508(.dina(n5566), .dinb(n5562), .dout(n5700));
  jand g05509(.dina(n5567), .dinb(n5553), .dout(n5701));
  jnot g05510(.din(n5701), .dout(n5702));
  jand g05511(.dina(n5702), .dinb(n5700), .dout(n5703));
  jxor g05512(.dina(n5703), .dinb(n5699), .dout(n5704));
  jxor g05513(.dina(n5704), .dinb(n5658), .dout(n5705));
  jxor g05514(.dina(n5705), .dinb(n5587), .dout(n5706));
  jxor g05515(.dina(n5706), .dinb(n5584), .dout(n5707));
  jand g05516(.dina(n5488), .dinb(n5485), .dout(n5708));
  jand g05517(.dina(n5505), .dinb(n5489), .dout(n5709));
  jor  g05518(.dina(n5709), .dinb(n5708), .dout(n5710));
  jnot g05519(.din(n5527), .dout(n5711));
  jand g05520(.dina(n5481), .dinb(n5476), .dout(n5712));
  jor  g05521(.dina(n5712), .dinb(n5478), .dout(n5713));
  jxor g05522(.dina(n5713), .dinb(n5711), .dout(n5714));
  jand g05523(.dina(n5451), .dinb(n5449), .dout(n5715));
  jnot g05524(.din(n5715), .dout(n5716));
  jand g05525(.dina(n5716), .dinb(n5454), .dout(n5717));
  jxor g05526(.dina(n5717), .dinb(n5714), .dout(n5718));
  jor  g05527(.dina(n5456), .dinb(n5447), .dout(n5719));
  jand g05528(.dina(n5457), .dinb(n5438), .dout(n5720));
  jnot g05529(.din(n5720), .dout(n5721));
  jand g05530(.dina(n5721), .dinb(n5719), .dout(n5722));
  jnot g05531(.din(n5722), .dout(n5723));
  jand g05532(.dina(n5515), .dinb(n5256), .dout(n5724));
  jand g05533(.dina(n5533), .dinb(n5516), .dout(n5725));
  jor  g05534(.dina(n5725), .dinb(n5724), .dout(n5726));
  jxor g05535(.dina(n5726), .dinb(n5723), .dout(n5727));
  jxor g05536(.dina(n5727), .dinb(n5718), .dout(n5728));
  jnot g05537(.din(n5392), .dout(n5729));
  jand g05538(.dina(n5445), .dinb(n5439), .dout(n5730));
  jor  g05539(.dina(n5730), .dinb(n5440), .dout(n5731));
  jxor g05540(.dina(n5731), .dinb(n5729), .dout(n5732));
  jand g05541(.dina(n5415), .dinb(n5413), .dout(n5733));
  jnot g05542(.din(n5733), .dout(n5734));
  jand g05543(.dina(n5734), .dinb(n5418), .dout(n5735));
  jxor g05544(.dina(n5735), .dinb(n5732), .dout(n5736));
  jand g05545(.dina(n5409), .dinb(n5399), .dout(n5737));
  jnot g05546(.din(n5737), .dout(n5738));
  jor  g05547(.dina(n5420), .dinb(n5411), .dout(n5739));
  jand g05548(.dina(n5739), .dinb(n5738), .dout(n5740));
  jnot g05549(.din(n5740), .dout(n5741));
  jand g05550(.dina(n1677), .dinb(\a[52] ), .dout(n5742));
  jnot g05551(.din(n5742), .dout(n5743));
  jand g05552(.dina(\a[52] ), .dinb(\a[1] ), .dout(n5744));
  jor  g05553(.dina(n5744), .dinb(\a[27] ), .dout(n5745));
  jand g05554(.dina(n5745), .dinb(n5743), .dout(n5746));
  jand g05555(.dina(n5403), .dinb(n5401), .dout(n5747));
  jnot g05556(.din(n5747), .dout(n5748));
  jand g05557(.dina(n5748), .dinb(n5406), .dout(n5749));
  jxor g05558(.dina(n5749), .dinb(n5746), .dout(n5750));
  jxor g05559(.dina(n5750), .dinb(n5434), .dout(n5751));
  jxor g05560(.dina(n5751), .dinb(n5741), .dout(n5752));
  jxor g05561(.dina(n5752), .dinb(n5736), .dout(n5753));
  jxor g05562(.dina(n5753), .dinb(n5728), .dout(n5754));
  jxor g05563(.dina(n5754), .dinb(n5710), .dout(n5755));
  jand g05564(.dina(n5458), .dinb(n5421), .dout(n5756));
  jand g05565(.dina(n5459), .dinb(n5381), .dout(n5757));
  jor  g05566(.dina(n5757), .dinb(n5756), .dout(n5758));
  jand g05567(.dina(n5548), .dinb(n5545), .dout(n5759));
  jand g05568(.dina(n5552), .dinb(n5549), .dout(n5760));
  jor  g05569(.dina(n5760), .dinb(n5759), .dout(n5761));
  jand g05570(.dina(n5498), .dinb(n5496), .dout(n5762));
  jand g05571(.dina(n5502), .dinb(n5499), .dout(n5763));
  jor  g05572(.dina(n5763), .dinb(n5762), .dout(n5764));
  jxor g05573(.dina(n5764), .dinb(n5761), .dout(n5765));
  jand g05574(.dina(n5559), .dinb(n5556), .dout(n5766));
  jand g05575(.dina(n5560), .dinb(n5208), .dout(n5767));
  jor  g05576(.dina(n5767), .dinb(n5766), .dout(n5768));
  jxor g05577(.dina(n5768), .dinb(n5765), .dout(n5769));
  jnot g05578(.din(n5769), .dout(n5770));
  jand g05579(.dina(n5534), .dinb(n5512), .dout(n5771));
  jnot g05580(.din(n5771), .dout(n5772));
  jor  g05581(.dina(n5540), .dinb(n5536), .dout(n5773));
  jand g05582(.dina(n5773), .dinb(n5772), .dout(n5774));
  jxor g05583(.dina(n5774), .dinb(n5770), .dout(n5775));
  jxor g05584(.dina(n5775), .dinb(n5758), .dout(n5776));
  jand g05585(.dina(n5460), .dinb(n5376), .dout(n5777));
  jand g05586(.dina(n5461), .dinb(n5373), .dout(n5778));
  jor  g05587(.dina(n5778), .dinb(n5777), .dout(n5779));
  jxor g05588(.dina(n5779), .dinb(n5776), .dout(n5780));
  jxor g05589(.dina(n5780), .dinb(n5755), .dout(n5781));
  jxor g05590(.dina(n5781), .dinb(n5707), .dout(n5782));
  jand g05591(.dina(n5782), .dinb(n5581), .dout(n5783));
  jor  g05592(.dina(n5782), .dinb(n5581), .dout(n5784));
  jnot g05593(.din(n5784), .dout(n5785));
  jor  g05594(.dina(n5785), .dinb(n5783), .dout(n5786));
  jand g05595(.dina(n5572), .dinb(n5370), .dout(n5787));
  jnot g05596(.din(n5787), .dout(n5788));
  jnot g05597(.din(n5370), .dout(n5789));
  jand g05598(.dina(n5573), .dinb(n5789), .dout(n5790));
  jor  g05599(.dina(n5577), .dinb(n5790), .dout(n5791));
  jand g05600(.dina(n5791), .dinb(n5788), .dout(n5792));
  jxor g05601(.dina(n5792), .dinb(n5786), .dout(\asquared[54] ));
  jand g05602(.dina(n5706), .dinb(n5584), .dout(n5794));
  jand g05603(.dina(n5781), .dinb(n5707), .dout(n5795));
  jor  g05604(.dina(n5795), .dinb(n5794), .dout(n5796));
  jand g05605(.dina(n5779), .dinb(n5776), .dout(n5797));
  jand g05606(.dina(n5780), .dinb(n5755), .dout(n5798));
  jor  g05607(.dina(n5798), .dinb(n5797), .dout(n5799));
  jand g05608(.dina(n5753), .dinb(n5728), .dout(n5800));
  jand g05609(.dina(n5754), .dinb(n5710), .dout(n5801));
  jor  g05610(.dina(n5801), .dinb(n5800), .dout(n5802));
  jnot g05611(.din(n5802), .dout(n5803));
  jor  g05612(.dina(n5774), .dinb(n5770), .dout(n5804));
  jand g05613(.dina(n5775), .dinb(n5758), .dout(n5805));
  jnot g05614(.din(n5805), .dout(n5806));
  jand g05615(.dina(n5806), .dinb(n5804), .dout(n5807));
  jxor g05616(.dina(n5807), .dinb(n5803), .dout(n5808));
  jand g05617(.dina(n5751), .dinb(n5741), .dout(n5809));
  jand g05618(.dina(n5752), .dinb(n5736), .dout(n5810));
  jor  g05619(.dina(n5810), .dinb(n5809), .dout(n5811));
  jand g05620(.dina(n5726), .dinb(n5723), .dout(n5812));
  jand g05621(.dina(n5727), .dinb(n5718), .dout(n5813));
  jor  g05622(.dina(n5813), .dinb(n5812), .dout(n5814));
  jand g05623(.dina(\a[35] ), .dinb(\a[19] ), .dout(n5815));
  jand g05624(.dina(n2671), .dinb(n1376), .dout(n5816));
  jnot g05625(.din(n5816), .dout(n5817));
  jand g05626(.dina(\a[33] ), .dinb(\a[21] ), .dout(n5818));
  jand g05627(.dina(\a[32] ), .dinb(\a[22] ), .dout(n5819));
  jor  g05628(.dina(n5819), .dinb(n5818), .dout(n5820));
  jand g05629(.dina(n5820), .dinb(n5817), .dout(n5821));
  jxor g05630(.dina(n5821), .dinb(n5815), .dout(n5822));
  jnot g05631(.din(n5822), .dout(n5823));
  jand g05632(.dina(\a[31] ), .dinb(\a[23] ), .dout(n5824));
  jnot g05633(.din(n5824), .dout(n5825));
  jand g05634(.dina(n3294), .dinb(n1648), .dout(n5826));
  jnot g05635(.din(n5826), .dout(n5827));
  jand g05636(.dina(\a[29] ), .dinb(\a[25] ), .dout(n5828));
  jand g05637(.dina(\a[30] ), .dinb(\a[24] ), .dout(n5829));
  jor  g05638(.dina(n5829), .dinb(n5828), .dout(n5830));
  jand g05639(.dina(n5830), .dinb(n5827), .dout(n5831));
  jxor g05640(.dina(n5831), .dinb(n5825), .dout(n5832));
  jxor g05641(.dina(n5832), .dinb(n5823), .dout(n5833));
  jand g05642(.dina(\a[54] ), .dinb(\a[0] ), .dout(n5834));
  jxor g05643(.dina(n5834), .dinb(n5742), .dout(n5835));
  jand g05644(.dina(\a[53] ), .dinb(\a[1] ), .dout(n5836));
  jxor g05645(.dina(n5836), .dinb(n3455), .dout(n5837));
  jxor g05646(.dina(n5837), .dinb(n5835), .dout(n5838));
  jxor g05647(.dina(n5838), .dinb(n5833), .dout(n5839));
  jxor g05648(.dina(n5839), .dinb(n5814), .dout(n5840));
  jxor g05649(.dina(n5840), .dinb(n5811), .dout(n5841));
  jxor g05650(.dina(n5841), .dinb(n5808), .dout(n5842));
  jxor g05651(.dina(n5842), .dinb(n5799), .dout(n5843));
  jand g05652(.dina(n5704), .dinb(n5658), .dout(n5844));
  jand g05653(.dina(n5705), .dinb(n5587), .dout(n5845));
  jor  g05654(.dina(n5845), .dinb(n5844), .dout(n5846));
  jand g05655(.dina(n5731), .dinb(n5729), .dout(n5847));
  jand g05656(.dina(n5735), .dinb(n5732), .dout(n5848));
  jor  g05657(.dina(n5848), .dinb(n5847), .dout(n5849));
  jand g05658(.dina(n5713), .dinb(n5711), .dout(n5850));
  jand g05659(.dina(n5717), .dinb(n5714), .dout(n5851));
  jor  g05660(.dina(n5851), .dinb(n5850), .dout(n5852));
  jxor g05661(.dina(n5852), .dinb(n5849), .dout(n5853));
  jand g05662(.dina(n5749), .dinb(n5746), .dout(n5854));
  jand g05663(.dina(n5750), .dinb(n5434), .dout(n5855));
  jor  g05664(.dina(n5855), .dinb(n5854), .dout(n5856));
  jxor g05665(.dina(n5856), .dinb(n5853), .dout(n5857));
  jand g05666(.dina(n5618), .dinb(n5590), .dout(n5858));
  jand g05667(.dina(n5657), .dinb(n5619), .dout(n5859));
  jor  g05668(.dina(n5859), .dinb(n5858), .dout(n5860));
  jxor g05669(.dina(n5860), .dinb(n5857), .dout(n5861));
  jnot g05670(.din(n5629), .dout(n5862));
  jor  g05671(.dina(n5654), .dinb(n5653), .dout(n5863));
  jand g05672(.dina(n5654), .dinb(n5653), .dout(n5864));
  jor  g05673(.dina(n5864), .dinb(n5652), .dout(n5865));
  jand g05674(.dina(n5865), .dinb(n5863), .dout(n5866));
  jxor g05675(.dina(n5866), .dinb(n5862), .dout(n5867));
  jand g05676(.dina(n5692), .dinb(n5690), .dout(n5868));
  jnot g05677(.din(n5868), .dout(n5869));
  jand g05678(.dina(n5869), .dinb(n5694), .dout(n5870));
  jxor g05679(.dina(n5870), .dinb(n5867), .dout(n5871));
  jand g05680(.dina(n5604), .dinb(n5599), .dout(n5872));
  jor  g05681(.dina(n5872), .dinb(n5600), .dout(n5873));
  jand g05682(.dina(n5612), .dinb(n5610), .dout(n5874));
  jnot g05683(.din(n5874), .dout(n5875));
  jand g05684(.dina(n5875), .dinb(n5615), .dout(n5876));
  jxor g05685(.dina(n5876), .dinb(n5873), .dout(n5877));
  jand g05686(.dina(n5680), .dinb(n5678), .dout(n5878));
  jnot g05687(.din(n5878), .dout(n5879));
  jand g05688(.dina(n5879), .dinb(n5683), .dout(n5880));
  jxor g05689(.dina(n5880), .dinb(n5877), .dout(n5881));
  jand g05690(.dina(n5650), .dinb(n5635), .dout(n5882));
  jand g05691(.dina(n5656), .dinb(n5651), .dout(n5883));
  jor  g05692(.dina(n5883), .dinb(n5882), .dout(n5884));
  jxor g05693(.dina(n5884), .dinb(n5881), .dout(n5885));
  jxor g05694(.dina(n5885), .dinb(n5871), .dout(n5886));
  jxor g05695(.dina(n5886), .dinb(n5861), .dout(n5887));
  jxor g05696(.dina(n5887), .dinb(n5846), .dout(n5888));
  jand g05697(.dina(n5764), .dinb(n5761), .dout(n5889));
  jand g05698(.dina(n5768), .dinb(n5765), .dout(n5890));
  jor  g05699(.dina(n5890), .dinb(n5889), .dout(n5891));
  jand g05700(.dina(\a[37] ), .dinb(\a[17] ), .dout(n5892));
  jand g05701(.dina(\a[48] ), .dinb(\a[38] ), .dout(n5893));
  jand g05702(.dina(n5893), .dinb(n1131), .dout(n5894));
  jnot g05703(.din(n5894), .dout(n5895));
  jand g05704(.dina(\a[48] ), .dinb(\a[6] ), .dout(n5896));
  jand g05705(.dina(n5896), .dinb(n5892), .dout(n5897));
  jand g05706(.dina(\a[38] ), .dinb(\a[17] ), .dout(n5898));
  jand g05707(.dina(n5898), .dinb(n5654), .dout(n5899));
  jor  g05708(.dina(n5899), .dinb(n5897), .dout(n5900));
  jand g05709(.dina(n5900), .dinb(n5895), .dout(n5901));
  jnot g05710(.din(n5901), .dout(n5902));
  jand g05711(.dina(n5902), .dinb(n5892), .dout(n5903));
  jand g05712(.dina(\a[38] ), .dinb(\a[16] ), .dout(n5904));
  jor  g05713(.dina(n5904), .dinb(n5896), .dout(n5905));
  jor  g05714(.dina(n5900), .dinb(n5894), .dout(n5906));
  jnot g05715(.din(n5906), .dout(n5907));
  jand g05716(.dina(n5907), .dinb(n5905), .dout(n5908));
  jor  g05717(.dina(n5908), .dinb(n5903), .dout(n5909));
  jand g05718(.dina(\a[36] ), .dinb(\a[18] ), .dout(n5910));
  jand g05719(.dina(\a[49] ), .dinb(\a[5] ), .dout(n5911));
  jand g05720(.dina(n5911), .dinb(n5910), .dout(n5912));
  jnot g05721(.din(n5912), .dout(n5913));
  jand g05722(.dina(\a[34] ), .dinb(\a[20] ), .dout(n5914));
  jand g05723(.dina(n5914), .dinb(n5911), .dout(n5915));
  jand g05724(.dina(\a[36] ), .dinb(\a[34] ), .dout(n5916));
  jand g05725(.dina(n5916), .dinb(n1181), .dout(n5917));
  jor  g05726(.dina(n5917), .dinb(n5915), .dout(n5918));
  jand g05727(.dina(n5918), .dinb(n5913), .dout(n5919));
  jnot g05728(.din(n5919), .dout(n5920));
  jxor g05729(.dina(n5911), .dinb(n5910), .dout(n5921));
  jor  g05730(.dina(n5921), .dinb(n5914), .dout(n5922));
  jand g05731(.dina(n5922), .dinb(n5920), .dout(n5923));
  jand g05732(.dina(\a[41] ), .dinb(\a[13] ), .dout(n5924));
  jnot g05733(.din(n5924), .dout(n5925));
  jand g05734(.dina(n4317), .dinb(n555), .dout(n5926));
  jnot g05735(.din(n5926), .dout(n5927));
  jand g05736(.dina(\a[43] ), .dinb(\a[11] ), .dout(n5928));
  jand g05737(.dina(\a[42] ), .dinb(\a[12] ), .dout(n5929));
  jor  g05738(.dina(n5929), .dinb(n5928), .dout(n5930));
  jand g05739(.dina(n5930), .dinb(n5927), .dout(n5931));
  jxor g05740(.dina(n5931), .dinb(n5925), .dout(n5932));
  jnot g05741(.din(n5932), .dout(n5933));
  jxor g05742(.dina(n5933), .dinb(n5923), .dout(n5934));
  jxor g05743(.dina(n5934), .dinb(n5909), .dout(n5935));
  jxor g05744(.dina(n5935), .dinb(n5891), .dout(n5936));
  jand g05745(.dina(\a[45] ), .dinb(\a[9] ), .dout(n5937));
  jand g05746(.dina(\a[44] ), .dinb(\a[10] ), .dout(n5938));
  jand g05747(.dina(\a[40] ), .dinb(\a[14] ), .dout(n5939));
  jand g05748(.dina(n5939), .dinb(n5938), .dout(n5940));
  jnot g05749(.din(n5940), .dout(n5941));
  jand g05750(.dina(n4812), .dinb(n453), .dout(n5942));
  jand g05751(.dina(n5939), .dinb(n5937), .dout(n5943));
  jor  g05752(.dina(n5943), .dinb(n5942), .dout(n5944));
  jand g05753(.dina(n5944), .dinb(n5941), .dout(n5945));
  jnot g05754(.din(n5945), .dout(n5946));
  jand g05755(.dina(n5946), .dinb(n5937), .dout(n5947));
  jor  g05756(.dina(n5944), .dinb(n5940), .dout(n5948));
  jnot g05757(.din(n5948), .dout(n5949));
  jor  g05758(.dina(n5939), .dinb(n5938), .dout(n5950));
  jand g05759(.dina(n5950), .dinb(n5949), .dout(n5951));
  jor  g05760(.dina(n5951), .dinb(n5947), .dout(n5952));
  jand g05761(.dina(\a[39] ), .dinb(\a[15] ), .dout(n5953));
  jand g05762(.dina(n5953), .dinb(n5624), .dout(n5954));
  jand g05763(.dina(\a[47] ), .dinb(\a[8] ), .dout(n5955));
  jand g05764(.dina(n5955), .dinb(n5620), .dout(n5956));
  jor  g05765(.dina(n5956), .dinb(n5954), .dout(n5957));
  jand g05766(.dina(\a[46] ), .dinb(\a[8] ), .dout(n5958));
  jand g05767(.dina(n5958), .dinb(n5953), .dout(n5959));
  jnot g05768(.din(n5959), .dout(n5960));
  jand g05769(.dina(n5960), .dinb(n5957), .dout(n5961));
  jnot g05770(.din(n5961), .dout(n5962));
  jand g05771(.dina(n5962), .dinb(n5624), .dout(n5963));
  jor  g05772(.dina(n5959), .dinb(n5957), .dout(n5964));
  jnot g05773(.din(n5964), .dout(n5965));
  jor  g05774(.dina(n5958), .dinb(n5953), .dout(n5966));
  jand g05775(.dina(n5966), .dinb(n5965), .dout(n5967));
  jor  g05776(.dina(n5967), .dinb(n5963), .dout(n5968));
  jand g05777(.dina(\a[52] ), .dinb(\a[2] ), .dout(n5969));
  jand g05778(.dina(n5594), .dinb(n265), .dout(n5970));
  jnot g05779(.din(n5970), .dout(n5971));
  jand g05780(.dina(\a[51] ), .dinb(\a[3] ), .dout(n5972));
  jand g05781(.dina(\a[50] ), .dinb(\a[4] ), .dout(n5973));
  jor  g05782(.dina(n5973), .dinb(n5972), .dout(n5974));
  jand g05783(.dina(n5974), .dinb(n5971), .dout(n5975));
  jxor g05784(.dina(n5975), .dinb(n5969), .dout(n5976));
  jxor g05785(.dina(n5976), .dinb(n5968), .dout(n5977));
  jxor g05786(.dina(n5977), .dinb(n5952), .dout(n5978));
  jxor g05787(.dina(n5978), .dinb(n5936), .dout(n5979));
  jand g05788(.dina(n5697), .dinb(n5661), .dout(n5980));
  jnot g05789(.din(n5980), .dout(n5981));
  jor  g05790(.dina(n5703), .dinb(n5699), .dout(n5982));
  jand g05791(.dina(n5982), .dinb(n5981), .dout(n5983));
  jnot g05792(.din(n5983), .dout(n5984));
  jnot g05793(.din(n5672), .dout(n5985));
  jnot g05794(.din(n5644), .dout(n5986));
  jand g05795(.dina(n5597), .dinb(n5591), .dout(n5987));
  jor  g05796(.dina(n5987), .dinb(n5595), .dout(n5988));
  jxor g05797(.dina(n5988), .dinb(n5986), .dout(n5989));
  jxor g05798(.dina(n5989), .dinb(n5985), .dout(n5990));
  jand g05799(.dina(n5686), .dinb(n5677), .dout(n5991));
  jnot g05800(.din(n5991), .dout(n5992));
  jor  g05801(.dina(n5696), .dinb(n5688), .dout(n5993));
  jand g05802(.dina(n5993), .dinb(n5992), .dout(n5994));
  jand g05803(.dina(n5606), .dinb(n5598), .dout(n5995));
  jnot g05804(.din(n5995), .dout(n5996));
  jor  g05805(.dina(n5617), .dinb(n5608), .dout(n5997));
  jand g05806(.dina(n5997), .dinb(n5996), .dout(n5998));
  jxor g05807(.dina(n5998), .dinb(n5994), .dout(n5999));
  jxor g05808(.dina(n5999), .dinb(n5990), .dout(n6000));
  jxor g05809(.dina(n6000), .dinb(n5984), .dout(n6001));
  jxor g05810(.dina(n6001), .dinb(n5979), .dout(n6002));
  jxor g05811(.dina(n6002), .dinb(n5888), .dout(n6003));
  jxor g05812(.dina(n6003), .dinb(n5843), .dout(n6004));
  jand g05813(.dina(n6004), .dinb(n5796), .dout(n6005));
  jor  g05814(.dina(n6004), .dinb(n5796), .dout(n6006));
  jnot g05815(.din(n6006), .dout(n6007));
  jor  g05816(.dina(n6007), .dinb(n6005), .dout(n6008));
  jnot g05817(.din(n5783), .dout(n6009));
  jor  g05818(.dina(n5792), .dinb(n5785), .dout(n6010));
  jand g05819(.dina(n6010), .dinb(n6009), .dout(n6011));
  jxor g05820(.dina(n6011), .dinb(n6008), .dout(\asquared[55] ));
  jand g05821(.dina(n5842), .dinb(n5799), .dout(n6013));
  jand g05822(.dina(n6003), .dinb(n5843), .dout(n6014));
  jor  g05823(.dina(n6014), .dinb(n6013), .dout(n6015));
  jor  g05824(.dina(n5807), .dinb(n5803), .dout(n6016));
  jand g05825(.dina(n5841), .dinb(n5808), .dout(n6017));
  jnot g05826(.din(n6017), .dout(n6018));
  jand g05827(.dina(n6018), .dinb(n6016), .dout(n6019));
  jnot g05828(.din(n6019), .dout(n6020));
  jand g05829(.dina(n5935), .dinb(n5891), .dout(n6021));
  jand g05830(.dina(n5978), .dinb(n5936), .dout(n6022));
  jor  g05831(.dina(n6022), .dinb(n6021), .dout(n6023));
  jand g05832(.dina(n5866), .dinb(n5862), .dout(n6024));
  jand g05833(.dina(n5870), .dinb(n5867), .dout(n6025));
  jor  g05834(.dina(n6025), .dinb(n6024), .dout(n6026));
  jand g05835(.dina(n5988), .dinb(n5986), .dout(n6027));
  jand g05836(.dina(n5989), .dinb(n5985), .dout(n6028));
  jor  g05837(.dina(n6028), .dinb(n6027), .dout(n6029));
  jxor g05838(.dina(n6029), .dinb(n6026), .dout(n6030));
  jand g05839(.dina(n5836), .dinb(n3455), .dout(n6031));
  jnot g05840(.din(n6031), .dout(n6032));
  jand g05841(.dina(n1803), .dinb(\a[54] ), .dout(n6033));
  jand g05842(.dina(n6033), .dinb(n6032), .dout(n6034));
  jnot g05843(.din(n6034), .dout(n6035));
  jand g05844(.dina(\a[54] ), .dinb(\a[1] ), .dout(n6036));
  jand g05845(.dina(n6032), .dinb(\a[28] ), .dout(n6037));
  jor  g05846(.dina(n6037), .dinb(n6036), .dout(n6038));
  jand g05847(.dina(n6038), .dinb(n6035), .dout(n6039));
  jand g05848(.dina(n5927), .dinb(n5925), .dout(n6040));
  jnot g05849(.din(n6040), .dout(n6041));
  jand g05850(.dina(n6041), .dinb(n5930), .dout(n6042));
  jxor g05851(.dina(n6042), .dinb(n6039), .dout(n6043));
  jxor g05852(.dina(n6043), .dinb(n6030), .dout(n6044));
  jxor g05853(.dina(n6044), .dinb(n6023), .dout(n6045));
  jor  g05854(.dina(n5918), .dinb(n5912), .dout(n6046));
  jand g05855(.dina(n5975), .dinb(n5969), .dout(n6047));
  jor  g05856(.dina(n6047), .dinb(n5970), .dout(n6048));
  jxor g05857(.dina(n6048), .dinb(n5948), .dout(n6049));
  jxor g05858(.dina(n6049), .dinb(n6046), .dout(n6050));
  jnot g05859(.din(n6050), .dout(n6051));
  jor  g05860(.dina(n5832), .dinb(n5823), .dout(n6052));
  jand g05861(.dina(n5838), .dinb(n5833), .dout(n6053));
  jnot g05862(.din(n6053), .dout(n6054));
  jand g05863(.dina(n6054), .dinb(n6052), .dout(n6055));
  jxor g05864(.dina(n6055), .dinb(n6051), .dout(n6056));
  jand g05865(.dina(n5834), .dinb(n5742), .dout(n6057));
  jand g05866(.dina(n5837), .dinb(n5835), .dout(n6058));
  jor  g05867(.dina(n6058), .dinb(n6057), .dout(n6059));
  jxor g05868(.dina(n6059), .dinb(n5964), .dout(n6060));
  jnot g05869(.din(n6060), .dout(n6061));
  jand g05870(.dina(\a[50] ), .dinb(\a[5] ), .dout(n6062));
  jnot g05871(.din(n6062), .dout(n6063));
  jand g05872(.dina(n3138), .dinb(n1024), .dout(n6064));
  jnot g05873(.din(n6064), .dout(n6065));
  jand g05874(.dina(\a[37] ), .dinb(\a[18] ), .dout(n6066));
  jand g05875(.dina(\a[36] ), .dinb(\a[19] ), .dout(n6067));
  jor  g05876(.dina(n6067), .dinb(n6066), .dout(n6068));
  jand g05877(.dina(n6068), .dinb(n6065), .dout(n6069));
  jxor g05878(.dina(n6069), .dinb(n6063), .dout(n6070));
  jxor g05879(.dina(n6070), .dinb(n6061), .dout(n6071));
  jxor g05880(.dina(n6071), .dinb(n6056), .dout(n6072));
  jxor g05881(.dina(n6072), .dinb(n6045), .dout(n6073));
  jxor g05882(.dina(n6073), .dinb(n6020), .dout(n6074));
  jand g05883(.dina(n5839), .dinb(n5814), .dout(n6075));
  jand g05884(.dina(n5840), .dinb(n5811), .dout(n6076));
  jor  g05885(.dina(n6076), .dinb(n6075), .dout(n6077));
  jand g05886(.dina(n5821), .dinb(n5815), .dout(n6078));
  jor  g05887(.dina(n6078), .dinb(n5816), .dout(n6079));
  jand g05888(.dina(n5827), .dinb(n5825), .dout(n6080));
  jnot g05889(.din(n6080), .dout(n6081));
  jand g05890(.dina(n6081), .dinb(n5830), .dout(n6082));
  jxor g05891(.dina(n6082), .dinb(n6079), .dout(n6083));
  jxor g05892(.dina(n6083), .dinb(n5906), .dout(n6084));
  jand g05893(.dina(n5933), .dinb(n5923), .dout(n6085));
  jand g05894(.dina(n5934), .dinb(n5909), .dout(n6086));
  jor  g05895(.dina(n6086), .dinb(n6085), .dout(n6087));
  jand g05896(.dina(n5976), .dinb(n5968), .dout(n6088));
  jand g05897(.dina(n5977), .dinb(n5952), .dout(n6089));
  jor  g05898(.dina(n6089), .dinb(n6088), .dout(n6090));
  jxor g05899(.dina(n6090), .dinb(n6087), .dout(n6091));
  jxor g05900(.dina(n6091), .dinb(n6084), .dout(n6092));
  jxor g05901(.dina(n6092), .dinb(n6077), .dout(n6093));
  jand g05902(.dina(n5852), .dinb(n5849), .dout(n6094));
  jand g05903(.dina(n5856), .dinb(n5853), .dout(n6095));
  jor  g05904(.dina(n6095), .dinb(n6094), .dout(n6096));
  jand g05905(.dina(\a[44] ), .dinb(\a[42] ), .dout(n6097));
  jand g05906(.dina(n6097), .dinb(n816), .dout(n6098));
  jnot g05907(.din(n6098), .dout(n6099));
  jand g05908(.dina(n4812), .dinb(n655), .dout(n6100));
  jand g05909(.dina(\a[42] ), .dinb(\a[13] ), .dout(n6101));
  jand g05910(.dina(\a[45] ), .dinb(\a[10] ), .dout(n6102));
  jand g05911(.dina(n6102), .dinb(n6101), .dout(n6103));
  jor  g05912(.dina(n6103), .dinb(n6100), .dout(n6104));
  jnot g05913(.din(n6104), .dout(n6105));
  jand g05914(.dina(n6105), .dinb(n6099), .dout(n6106));
  jand g05915(.dina(\a[44] ), .dinb(\a[11] ), .dout(n6107));
  jor  g05916(.dina(n6107), .dinb(n6101), .dout(n6108));
  jand g05917(.dina(n6108), .dinb(n6106), .dout(n6109));
  jand g05918(.dina(n6104), .dinb(n6099), .dout(n6110));
  jnot g05919(.din(n6110), .dout(n6111));
  jand g05920(.dina(n6111), .dinb(n6102), .dout(n6112));
  jor  g05921(.dina(n6112), .dinb(n6109), .dout(n6113));
  jand g05922(.dina(\a[43] ), .dinb(\a[12] ), .dout(n6114));
  jand g05923(.dina(\a[29] ), .dinb(\a[26] ), .dout(n6115));
  jxor g05924(.dina(n6115), .dinb(n2042), .dout(n6116));
  jxor g05925(.dina(n6116), .dinb(n6114), .dout(n6117));
  jxor g05926(.dina(n6117), .dinb(n6113), .dout(n6118));
  jnot g05927(.din(n6118), .dout(n6119));
  jand g05928(.dina(\a[39] ), .dinb(\a[16] ), .dout(n6120));
  jnot g05929(.din(n6120), .dout(n6121));
  jand g05930(.dina(n5316), .dinb(n499), .dout(n6122));
  jnot g05931(.din(n6122), .dout(n6123));
  jand g05932(.dina(\a[48] ), .dinb(\a[7] ), .dout(n6124));
  jor  g05933(.dina(n6124), .dinb(n5955), .dout(n6125));
  jand g05934(.dina(n6125), .dinb(n6123), .dout(n6126));
  jxor g05935(.dina(n6126), .dinb(n6121), .dout(n6127));
  jxor g05936(.dina(n6127), .dinb(n6119), .dout(n6128));
  jxor g05937(.dina(n6128), .dinb(n6096), .dout(n6129));
  jand g05938(.dina(\a[53] ), .dinb(\a[51] ), .dout(n6130));
  jand g05939(.dina(n6130), .dinb(n245), .dout(n6131));
  jand g05940(.dina(n212), .dinb(\a[51] ), .dout(n6132));
  jand g05941(.dina(\a[53] ), .dinb(\a[2] ), .dout(n6133));
  jand g05942(.dina(n6133), .dinb(\a[0] ), .dout(n6134));
  jor  g05943(.dina(n6134), .dinb(n6132), .dout(n6135));
  jand g05944(.dina(n6135), .dinb(\a[55] ), .dout(n6136));
  jor  g05945(.dina(n6136), .dinb(n6131), .dout(n6137));
  jnot g05946(.din(n6137), .dout(n6138));
  jand g05947(.dina(\a[51] ), .dinb(\a[4] ), .dout(n6139));
  jor  g05948(.dina(n6139), .dinb(n6133), .dout(n6140));
  jand g05949(.dina(n6140), .dinb(n6138), .dout(n6141));
  jnot g05950(.din(n6141), .dout(n6142));
  jnot g05951(.din(\a[55] ), .dout(n6143));
  jnot g05952(.din(n6131), .dout(n6144));
  jand g05953(.dina(n6135), .dinb(n6144), .dout(n6145));
  jor  g05954(.dina(n6145), .dinb(n6143), .dout(n6146));
  jor  g05955(.dina(n6146), .dinb(n193), .dout(n6147));
  jand g05956(.dina(n6147), .dinb(n6142), .dout(n6148));
  jand g05957(.dina(\a[35] ), .dinb(\a[20] ), .dout(n6149));
  jnot g05958(.din(n6149), .dout(n6150));
  jand g05959(.dina(n3634), .dinb(n1376), .dout(n6151));
  jnot g05960(.din(n6151), .dout(n6152));
  jand g05961(.dina(\a[34] ), .dinb(\a[21] ), .dout(n6153));
  jor  g05962(.dina(n6153), .dinb(n2248), .dout(n6154));
  jand g05963(.dina(n6154), .dinb(n6152), .dout(n6155));
  jxor g05964(.dina(n6155), .dinb(n6150), .dout(n6156));
  jxor g05965(.dina(n6156), .dinb(n6148), .dout(n6157));
  jnot g05966(.din(n6157), .dout(n6158));
  jand g05967(.dina(\a[32] ), .dinb(\a[23] ), .dout(n6159));
  jnot g05968(.din(n6159), .dout(n6160));
  jand g05969(.dina(n2440), .dinb(n1648), .dout(n6161));
  jnot g05970(.din(n6161), .dout(n6162));
  jand g05971(.dina(\a[31] ), .dinb(\a[24] ), .dout(n6163));
  jand g05972(.dina(\a[30] ), .dinb(\a[25] ), .dout(n6164));
  jor  g05973(.dina(n6164), .dinb(n6163), .dout(n6165));
  jand g05974(.dina(n6165), .dinb(n6162), .dout(n6166));
  jxor g05975(.dina(n6166), .dinb(n6160), .dout(n6167));
  jxor g05976(.dina(n6167), .dinb(n6158), .dout(n6168));
  jxor g05977(.dina(n6168), .dinb(n6129), .dout(n6169));
  jxor g05978(.dina(n6169), .dinb(n6093), .dout(n6170));
  jxor g05979(.dina(n6170), .dinb(n6074), .dout(n6171));
  jand g05980(.dina(n5887), .dinb(n5846), .dout(n6172));
  jand g05981(.dina(n6002), .dinb(n5888), .dout(n6173));
  jor  g05982(.dina(n6173), .dinb(n6172), .dout(n6174));
  jand g05983(.dina(n6000), .dinb(n5984), .dout(n6175));
  jand g05984(.dina(n6001), .dinb(n5979), .dout(n6176));
  jor  g05985(.dina(n6176), .dinb(n6175), .dout(n6177));
  jand g05986(.dina(n5860), .dinb(n5857), .dout(n6178));
  jand g05987(.dina(n5886), .dinb(n5861), .dout(n6179));
  jor  g05988(.dina(n6179), .dinb(n6178), .dout(n6180));
  jand g05989(.dina(n5884), .dinb(n5881), .dout(n6181));
  jand g05990(.dina(n5885), .dinb(n5871), .dout(n6182));
  jor  g05991(.dina(n6182), .dinb(n6181), .dout(n6183));
  jand g05992(.dina(n5876), .dinb(n5873), .dout(n6184));
  jand g05993(.dina(n5880), .dinb(n5877), .dout(n6185));
  jor  g05994(.dina(n6185), .dinb(n6184), .dout(n6186));
  jand g05995(.dina(\a[52] ), .dinb(\a[3] ), .dout(n6187));
  jand g05996(.dina(\a[49] ), .dinb(\a[6] ), .dout(n6188));
  jxor g05997(.dina(n6188), .dinb(n5898), .dout(n6189));
  jxor g05998(.dina(n6189), .dinb(n6187), .dout(n6190));
  jand g05999(.dina(\a[40] ), .dinb(\a[15] ), .dout(n6191));
  jand g06000(.dina(\a[46] ), .dinb(\a[9] ), .dout(n6192));
  jand g06001(.dina(\a[41] ), .dinb(\a[14] ), .dout(n6193));
  jxor g06002(.dina(n6193), .dinb(n6192), .dout(n6194));
  jxor g06003(.dina(n6194), .dinb(n6191), .dout(n6195));
  jxor g06004(.dina(n6195), .dinb(n6190), .dout(n6196));
  jxor g06005(.dina(n6196), .dinb(n6186), .dout(n6197));
  jnot g06006(.din(n6197), .dout(n6198));
  jor  g06007(.dina(n5998), .dinb(n5994), .dout(n6199));
  jand g06008(.dina(n5999), .dinb(n5990), .dout(n6200));
  jnot g06009(.din(n6200), .dout(n6201));
  jand g06010(.dina(n6201), .dinb(n6199), .dout(n6202));
  jxor g06011(.dina(n6202), .dinb(n6198), .dout(n6203));
  jxor g06012(.dina(n6203), .dinb(n6183), .dout(n6204));
  jxor g06013(.dina(n6204), .dinb(n6180), .dout(n6205));
  jxor g06014(.dina(n6205), .dinb(n6177), .dout(n6206));
  jxor g06015(.dina(n6206), .dinb(n6174), .dout(n6207));
  jxor g06016(.dina(n6207), .dinb(n6171), .dout(n6208));
  jand g06017(.dina(n6208), .dinb(n6015), .dout(n6209));
  jor  g06018(.dina(n6208), .dinb(n6015), .dout(n6210));
  jnot g06019(.din(n6210), .dout(n6211));
  jor  g06020(.dina(n6211), .dinb(n6209), .dout(n6212));
  jnot g06021(.din(n6005), .dout(n6213));
  jor  g06022(.dina(n6011), .dinb(n6007), .dout(n6214));
  jand g06023(.dina(n6214), .dinb(n6213), .dout(n6215));
  jxor g06024(.dina(n6215), .dinb(n6212), .dout(\asquared[56] ));
  jand g06025(.dina(n6206), .dinb(n6174), .dout(n6217));
  jand g06026(.dina(n6207), .dinb(n6171), .dout(n6218));
  jor  g06027(.dina(n6218), .dinb(n6217), .dout(n6219));
  jand g06028(.dina(\a[49] ), .dinb(\a[7] ), .dout(n6220));
  jnot g06029(.din(n6220), .dout(n6221));
  jand g06030(.dina(\a[39] ), .dinb(\a[17] ), .dout(n6222));
  jnot g06031(.din(n6222), .dout(n6223));
  jand g06032(.dina(n6223), .dinb(n6221), .dout(n6224));
  jand g06033(.dina(n6222), .dinb(n6220), .dout(n6225));
  jnot g06034(.din(n6225), .dout(n6226));
  jand g06035(.dina(\a[50] ), .dinb(\a[7] ), .dout(n6227));
  jand g06036(.dina(n6227), .dinb(n6188), .dout(n6228));
  jand g06037(.dina(\a[50] ), .dinb(\a[6] ), .dout(n6229));
  jand g06038(.dina(n6229), .dinb(n6222), .dout(n6230));
  jor  g06039(.dina(n6230), .dinb(n6228), .dout(n6231));
  jnot g06040(.din(n6231), .dout(n6232));
  jand g06041(.dina(n6232), .dinb(n6226), .dout(n6233));
  jnot g06042(.din(n6233), .dout(n6234));
  jor  g06043(.dina(n6234), .dinb(n6224), .dout(n6235));
  jand g06044(.dina(n6231), .dinb(n6226), .dout(n6236));
  jnot g06045(.din(n6236), .dout(n6237));
  jand g06046(.dina(n6237), .dinb(n6229), .dout(n6238));
  jnot g06047(.din(n6238), .dout(n6239));
  jand g06048(.dina(n6239), .dinb(n6235), .dout(n6240));
  jand g06049(.dina(\a[45] ), .dinb(\a[11] ), .dout(n6241));
  jnot g06050(.din(n6241), .dout(n6242));
  jand g06051(.dina(n4495), .dinb(n899), .dout(n6243));
  jnot g06052(.din(n6243), .dout(n6244));
  jand g06053(.dina(\a[43] ), .dinb(\a[13] ), .dout(n6245));
  jand g06054(.dina(\a[44] ), .dinb(\a[12] ), .dout(n6246));
  jor  g06055(.dina(n6246), .dinb(n6245), .dout(n6247));
  jand g06056(.dina(n6247), .dinb(n6244), .dout(n6248));
  jxor g06057(.dina(n6248), .dinb(n6242), .dout(n6249));
  jxor g06058(.dina(n6249), .dinb(n6240), .dout(n6250));
  jand g06059(.dina(\a[40] ), .dinb(\a[16] ), .dout(n6251));
  jand g06060(.dina(\a[48] ), .dinb(\a[8] ), .dout(n6252));
  jand g06061(.dina(\a[41] ), .dinb(\a[15] ), .dout(n6253));
  jxor g06062(.dina(n6253), .dinb(n6252), .dout(n6254));
  jxor g06063(.dina(n6254), .dinb(n6251), .dout(n6255));
  jxor g06064(.dina(n6255), .dinb(n6250), .dout(n6256));
  jand g06065(.dina(\a[47] ), .dinb(\a[9] ), .dout(n6257));
  jand g06066(.dina(\a[46] ), .dinb(\a[10] ), .dout(n6258));
  jand g06067(.dina(\a[42] ), .dinb(\a[14] ), .dout(n6259));
  jand g06068(.dina(n6259), .dinb(n6258), .dout(n6260));
  jnot g06069(.din(n6260), .dout(n6261));
  jand g06070(.dina(\a[47] ), .dinb(\a[10] ), .dout(n6262));
  jand g06071(.dina(n6262), .dinb(n6192), .dout(n6263));
  jand g06072(.dina(n6259), .dinb(n6257), .dout(n6264));
  jor  g06073(.dina(n6264), .dinb(n6263), .dout(n6265));
  jand g06074(.dina(n6265), .dinb(n6261), .dout(n6266));
  jnot g06075(.din(n6266), .dout(n6267));
  jand g06076(.dina(n6267), .dinb(n6257), .dout(n6268));
  jor  g06077(.dina(n6265), .dinb(n6260), .dout(n6269));
  jnot g06078(.din(n6269), .dout(n6270));
  jor  g06079(.dina(n6259), .dinb(n6258), .dout(n6271));
  jand g06080(.dina(n6271), .dinb(n6270), .dout(n6272));
  jor  g06081(.dina(n6272), .dinb(n6268), .dout(n6273));
  jand g06082(.dina(\a[36] ), .dinb(\a[20] ), .dout(n6274));
  jand g06083(.dina(n3634), .dinb(n1658), .dout(n6275));
  jnot g06084(.din(n6275), .dout(n6276));
  jand g06085(.dina(\a[34] ), .dinb(\a[22] ), .dout(n6277));
  jand g06086(.dina(\a[33] ), .dinb(\a[23] ), .dout(n6278));
  jor  g06087(.dina(n6278), .dinb(n6277), .dout(n6279));
  jand g06088(.dina(n6279), .dinb(n6276), .dout(n6280));
  jxor g06089(.dina(n6280), .dinb(n6274), .dout(n6281));
  jnot g06090(.din(n6281), .dout(n6282));
  jand g06091(.dina(\a[32] ), .dinb(\a[24] ), .dout(n6283));
  jnot g06092(.din(n6283), .dout(n6284));
  jand g06093(.dina(n2440), .dinb(n2128), .dout(n6285));
  jnot g06094(.din(n6285), .dout(n6286));
  jand g06095(.dina(\a[31] ), .dinb(\a[25] ), .dout(n6287));
  jand g06096(.dina(\a[30] ), .dinb(\a[26] ), .dout(n6288));
  jor  g06097(.dina(n6288), .dinb(n6287), .dout(n6289));
  jand g06098(.dina(n6289), .dinb(n6286), .dout(n6290));
  jxor g06099(.dina(n6290), .dinb(n6284), .dout(n6291));
  jxor g06100(.dina(n6291), .dinb(n6282), .dout(n6292));
  jxor g06101(.dina(n6292), .dinb(n6273), .dout(n6293));
  jxor g06102(.dina(n6293), .dinb(n6256), .dout(n6294));
  jand g06103(.dina(\a[56] ), .dinb(\a[2] ), .dout(n6295));
  jand g06104(.dina(n6295), .dinb(n5834), .dout(n6296));
  jnot g06105(.din(n6296), .dout(n6297));
  jand g06106(.dina(\a[56] ), .dinb(\a[0] ), .dout(n6298));
  jand g06107(.dina(\a[54] ), .dinb(\a[2] ), .dout(n6299));
  jor  g06108(.dina(n6299), .dinb(n6298), .dout(n6300));
  jand g06109(.dina(n6300), .dinb(n6297), .dout(n6301));
  jxor g06110(.dina(n6301), .dinb(n6033), .dout(n6302));
  jand g06111(.dina(n6123), .dinb(n6121), .dout(n6303));
  jnot g06112(.din(n6303), .dout(n6304));
  jand g06113(.dina(n6304), .dinb(n6125), .dout(n6305));
  jxor g06114(.dina(n6305), .dinb(n6302), .dout(n6306));
  jnot g06115(.din(n6306), .dout(n6307));
  jand g06116(.dina(\a[53] ), .dinb(\a[3] ), .dout(n6308));
  jnot g06117(.din(n6308), .dout(n6309));
  jand g06118(.dina(\a[52] ), .dinb(\a[4] ), .dout(n6310));
  jand g06119(.dina(\a[37] ), .dinb(\a[19] ), .dout(n6311));
  jxor g06120(.dina(n6311), .dinb(n6310), .dout(n6312));
  jxor g06121(.dina(n6312), .dinb(n6309), .dout(n6313));
  jxor g06122(.dina(n6313), .dinb(n6307), .dout(n6314));
  jxor g06123(.dina(n6314), .dinb(n6294), .dout(n6315));
  jor  g06124(.dina(n6202), .dinb(n6198), .dout(n6316));
  jand g06125(.dina(n6203), .dinb(n6183), .dout(n6317));
  jnot g06126(.din(n6317), .dout(n6318));
  jand g06127(.dina(n6318), .dinb(n6316), .dout(n6319));
  jnot g06128(.din(n6319), .dout(n6320));
  jand g06129(.dina(n6188), .dinb(n5898), .dout(n6321));
  jand g06130(.dina(n6189), .dinb(n6187), .dout(n6322));
  jor  g06131(.dina(n6322), .dinb(n6321), .dout(n6323));
  jand g06132(.dina(n6162), .dinb(n6160), .dout(n6324));
  jnot g06133(.din(n6324), .dout(n6325));
  jand g06134(.dina(n6325), .dinb(n6165), .dout(n6326));
  jand g06135(.dina(n6152), .dinb(n6150), .dout(n6327));
  jnot g06136(.din(n6327), .dout(n6328));
  jand g06137(.dina(n6328), .dinb(n6154), .dout(n6329));
  jxor g06138(.dina(n6329), .dinb(n6326), .dout(n6330));
  jxor g06139(.dina(n6330), .dinb(n6323), .dout(n6331));
  jand g06140(.dina(n6117), .dinb(n6113), .dout(n6332));
  jnot g06141(.din(n6332), .dout(n6333));
  jor  g06142(.dina(n6127), .dinb(n6119), .dout(n6334));
  jand g06143(.dina(n6334), .dinb(n6333), .dout(n6335));
  jnot g06144(.din(n6335), .dout(n6336));
  jnot g06145(.din(n6106), .dout(n6337));
  jand g06146(.dina(n6115), .dinb(n2042), .dout(n6338));
  jand g06147(.dina(n6116), .dinb(n6114), .dout(n6339));
  jor  g06148(.dina(n6339), .dinb(n6338), .dout(n6340));
  jand g06149(.dina(\a[55] ), .dinb(\a[1] ), .dout(n6341));
  jxor g06150(.dina(n6341), .dinb(n2536), .dout(n6342));
  jxor g06151(.dina(n6342), .dinb(n6340), .dout(n6343));
  jxor g06152(.dina(n6343), .dinb(n6337), .dout(n6344));
  jxor g06153(.dina(n6344), .dinb(n6336), .dout(n6345));
  jxor g06154(.dina(n6345), .dinb(n6331), .dout(n6346));
  jxor g06155(.dina(n6346), .dinb(n6320), .dout(n6347));
  jxor g06156(.dina(n6347), .dinb(n6315), .dout(n6348));
  jand g06157(.dina(n6204), .dinb(n6180), .dout(n6349));
  jand g06158(.dina(n6205), .dinb(n6177), .dout(n6350));
  jor  g06159(.dina(n6350), .dinb(n6349), .dout(n6351));
  jand g06160(.dina(n6065), .dinb(n6063), .dout(n6352));
  jnot g06161(.din(n6352), .dout(n6353));
  jand g06162(.dina(n6353), .dinb(n6068), .dout(n6354));
  jxor g06163(.dina(n6354), .dinb(n6137), .dout(n6355));
  jor  g06164(.dina(n6193), .dinb(n6192), .dout(n6356));
  jand g06165(.dina(n6193), .dinb(n6192), .dout(n6357));
  jor  g06166(.dina(n6357), .dinb(n6191), .dout(n6358));
  jand g06167(.dina(n6358), .dinb(n6356), .dout(n6359));
  jxor g06168(.dina(n6359), .dinb(n6355), .dout(n6360));
  jand g06169(.dina(n6195), .dinb(n6190), .dout(n6361));
  jand g06170(.dina(n6196), .dinb(n6186), .dout(n6362));
  jor  g06171(.dina(n6362), .dinb(n6361), .dout(n6363));
  jxor g06172(.dina(n6363), .dinb(n6360), .dout(n6364));
  jand g06173(.dina(n6029), .dinb(n6026), .dout(n6365));
  jand g06174(.dina(n6043), .dinb(n6030), .dout(n6366));
  jor  g06175(.dina(n6366), .dinb(n6365), .dout(n6367));
  jxor g06176(.dina(n6367), .dinb(n6364), .dout(n6368));
  jand g06177(.dina(n6082), .dinb(n6079), .dout(n6369));
  jand g06178(.dina(n6083), .dinb(n5906), .dout(n6370));
  jor  g06179(.dina(n6370), .dinb(n6369), .dout(n6371));
  jnot g06180(.din(n6371), .dout(n6372));
  jand g06181(.dina(n6059), .dinb(n5964), .dout(n6373));
  jnot g06182(.din(n6373), .dout(n6374));
  jor  g06183(.dina(n6070), .dinb(n6061), .dout(n6375));
  jand g06184(.dina(n6375), .dinb(n6374), .dout(n6376));
  jxor g06185(.dina(n6376), .dinb(n6372), .dout(n6377));
  jnot g06186(.din(n6377), .dout(n6378));
  jor  g06187(.dina(n6156), .dinb(n6148), .dout(n6379));
  jor  g06188(.dina(n6167), .dinb(n6158), .dout(n6380));
  jand g06189(.dina(n6380), .dinb(n6379), .dout(n6381));
  jxor g06190(.dina(n6381), .dinb(n6378), .dout(n6382));
  jand g06191(.dina(n6128), .dinb(n6096), .dout(n6383));
  jand g06192(.dina(n6168), .dinb(n6129), .dout(n6384));
  jor  g06193(.dina(n6384), .dinb(n6383), .dout(n6385));
  jxor g06194(.dina(n6385), .dinb(n6382), .dout(n6386));
  jxor g06195(.dina(n6386), .dinb(n6368), .dout(n6387));
  jxor g06196(.dina(n6387), .dinb(n6351), .dout(n6388));
  jxor g06197(.dina(n6388), .dinb(n6348), .dout(n6389));
  jor  g06198(.dina(n6055), .dinb(n6051), .dout(n6390));
  jand g06199(.dina(n6071), .dinb(n6056), .dout(n6391));
  jnot g06200(.din(n6391), .dout(n6392));
  jand g06201(.dina(n6392), .dinb(n6390), .dout(n6393));
  jnot g06202(.din(n6393), .dout(n6394));
  jand g06203(.dina(n6048), .dinb(n5948), .dout(n6395));
  jand g06204(.dina(n6049), .dinb(n6046), .dout(n6396));
  jor  g06205(.dina(n6396), .dinb(n6395), .dout(n6397));
  jand g06206(.dina(n6042), .dinb(n6039), .dout(n6398));
  jnot g06207(.din(\a[54] ), .dout(n6399));
  jand g06208(.dina(n6031), .dinb(n6399), .dout(n6400));
  jor  g06209(.dina(n6400), .dinb(n6398), .dout(n6401));
  jand g06210(.dina(\a[35] ), .dinb(\a[21] ), .dout(n6402));
  jnot g06211(.din(n6402), .dout(n6403));
  jand g06212(.dina(\a[51] ), .dinb(\a[38] ), .dout(n6404));
  jand g06213(.dina(n6404), .dinb(n1185), .dout(n6405));
  jnot g06214(.din(n6405), .dout(n6406));
  jand g06215(.dina(\a[51] ), .dinb(\a[5] ), .dout(n6407));
  jand g06216(.dina(\a[38] ), .dinb(\a[18] ), .dout(n6408));
  jor  g06217(.dina(n6408), .dinb(n6407), .dout(n6409));
  jand g06218(.dina(n6409), .dinb(n6406), .dout(n6410));
  jxor g06219(.dina(n6410), .dinb(n6403), .dout(n6411));
  jnot g06220(.din(n6411), .dout(n6412));
  jxor g06221(.dina(n6412), .dinb(n6401), .dout(n6413));
  jxor g06222(.dina(n6413), .dinb(n6397), .dout(n6414));
  jand g06223(.dina(n6090), .dinb(n6087), .dout(n6415));
  jand g06224(.dina(n6091), .dinb(n6084), .dout(n6416));
  jor  g06225(.dina(n6416), .dinb(n6415), .dout(n6417));
  jxor g06226(.dina(n6417), .dinb(n6414), .dout(n6418));
  jxor g06227(.dina(n6418), .dinb(n6394), .dout(n6419));
  jand g06228(.dina(n6044), .dinb(n6023), .dout(n6420));
  jand g06229(.dina(n6072), .dinb(n6045), .dout(n6421));
  jor  g06230(.dina(n6421), .dinb(n6420), .dout(n6422));
  jxor g06231(.dina(n6422), .dinb(n6419), .dout(n6423));
  jand g06232(.dina(n6092), .dinb(n6077), .dout(n6424));
  jand g06233(.dina(n6169), .dinb(n6093), .dout(n6425));
  jor  g06234(.dina(n6425), .dinb(n6424), .dout(n6426));
  jxor g06235(.dina(n6426), .dinb(n6423), .dout(n6427));
  jand g06236(.dina(n6073), .dinb(n6020), .dout(n6428));
  jand g06237(.dina(n6170), .dinb(n6074), .dout(n6429));
  jor  g06238(.dina(n6429), .dinb(n6428), .dout(n6430));
  jxor g06239(.dina(n6430), .dinb(n6427), .dout(n6431));
  jxor g06240(.dina(n6431), .dinb(n6389), .dout(n6432));
  jand g06241(.dina(n6432), .dinb(n6219), .dout(n6433));
  jor  g06242(.dina(n6432), .dinb(n6219), .dout(n6434));
  jnot g06243(.din(n6434), .dout(n6435));
  jor  g06244(.dina(n6435), .dinb(n6433), .dout(n6436));
  jnot g06245(.din(n6209), .dout(n6437));
  jor  g06246(.dina(n6215), .dinb(n6211), .dout(n6438));
  jand g06247(.dina(n6438), .dinb(n6437), .dout(n6439));
  jxor g06248(.dina(n6439), .dinb(n6436), .dout(\asquared[57] ));
  jand g06249(.dina(n6430), .dinb(n6427), .dout(n6441));
  jand g06250(.dina(n6431), .dinb(n6389), .dout(n6442));
  jor  g06251(.dina(n6442), .dinb(n6441), .dout(n6443));
  jand g06252(.dina(n6422), .dinb(n6419), .dout(n6444));
  jand g06253(.dina(n6426), .dinb(n6423), .dout(n6445));
  jor  g06254(.dina(n6445), .dinb(n6444), .dout(n6446));
  jand g06255(.dina(n6342), .dinb(n6340), .dout(n6447));
  jand g06256(.dina(n6343), .dinb(n6337), .dout(n6448));
  jor  g06257(.dina(n6448), .dinb(n6447), .dout(n6449));
  jnot g06258(.din(n6449), .dout(n6450));
  jand g06259(.dina(n6305), .dinb(n6302), .dout(n6451));
  jnot g06260(.din(n6451), .dout(n6452));
  jor  g06261(.dina(n6313), .dinb(n6307), .dout(n6453));
  jand g06262(.dina(n6453), .dinb(n6452), .dout(n6454));
  jxor g06263(.dina(n6454), .dinb(n6450), .dout(n6455));
  jnot g06264(.din(n6455), .dout(n6456));
  jor  g06265(.dina(n6291), .dinb(n6282), .dout(n6457));
  jand g06266(.dina(n6292), .dinb(n6273), .dout(n6458));
  jnot g06267(.din(n6458), .dout(n6459));
  jand g06268(.dina(n6459), .dinb(n6457), .dout(n6460));
  jxor g06269(.dina(n6460), .dinb(n6456), .dout(n6461));
  jand g06270(.dina(n6293), .dinb(n6256), .dout(n6462));
  jand g06271(.dina(n6314), .dinb(n6294), .dout(n6463));
  jor  g06272(.dina(n6463), .dinb(n6462), .dout(n6464));
  jxor g06273(.dina(n6464), .dinb(n6461), .dout(n6465));
  jor  g06274(.dina(n6249), .dinb(n6240), .dout(n6466));
  jand g06275(.dina(n6255), .dinb(n6250), .dout(n6467));
  jnot g06276(.din(n6467), .dout(n6468));
  jand g06277(.dina(n6468), .dinb(n6466), .dout(n6469));
  jnot g06278(.din(n6469), .dout(n6470));
  jand g06279(.dina(n6253), .dinb(n6252), .dout(n6471));
  jand g06280(.dina(n6254), .dinb(n6251), .dout(n6472));
  jor  g06281(.dina(n6472), .dinb(n6471), .dout(n6473));
  jand g06282(.dina(n6286), .dinb(n6284), .dout(n6474));
  jnot g06283(.din(n6474), .dout(n6475));
  jand g06284(.dina(n6475), .dinb(n6289), .dout(n6476));
  jxor g06285(.dina(n6476), .dinb(n6473), .dout(n6477));
  jxor g06286(.dina(n6477), .dinb(n6234), .dout(n6478));
  jand g06287(.dina(n6280), .dinb(n6274), .dout(n6479));
  jor  g06288(.dina(n6479), .dinb(n6275), .dout(n6480));
  jor  g06289(.dina(n6311), .dinb(n6310), .dout(n6481));
  jand g06290(.dina(n6311), .dinb(n6310), .dout(n6482));
  jor  g06291(.dina(n6482), .dinb(n6308), .dout(n6483));
  jand g06292(.dina(n6483), .dinb(n6481), .dout(n6484));
  jxor g06293(.dina(n6484), .dinb(n6480), .dout(n6485));
  jand g06294(.dina(n6301), .dinb(n6033), .dout(n6486));
  jor  g06295(.dina(n6486), .dinb(n6296), .dout(n6487));
  jxor g06296(.dina(n6487), .dinb(n6485), .dout(n6488));
  jxor g06297(.dina(n6488), .dinb(n6478), .dout(n6489));
  jxor g06298(.dina(n6489), .dinb(n6470), .dout(n6490));
  jxor g06299(.dina(n6490), .dinb(n6465), .dout(n6491));
  jxor g06300(.dina(n6491), .dinb(n6446), .dout(n6492));
  jor  g06301(.dina(n6376), .dinb(n6372), .dout(n6493));
  jor  g06302(.dina(n6381), .dinb(n6378), .dout(n6494));
  jand g06303(.dina(n6494), .dinb(n6493), .dout(n6495));
  jnot g06304(.din(n6495), .dout(n6496));
  jand g06305(.dina(\a[54] ), .dinb(\a[3] ), .dout(n6497));
  jand g06306(.dina(\a[55] ), .dinb(\a[53] ), .dout(n6498));
  jand g06307(.dina(n6498), .dinb(n245), .dout(n6499));
  jnot g06308(.din(n6499), .dout(n6500));
  jand g06309(.dina(\a[55] ), .dinb(\a[2] ), .dout(n6501));
  jand g06310(.dina(\a[53] ), .dinb(\a[4] ), .dout(n6502));
  jor  g06311(.dina(n6502), .dinb(n6501), .dout(n6503));
  jand g06312(.dina(n6503), .dinb(n6500), .dout(n6504));
  jxor g06313(.dina(n6504), .dinb(n6497), .dout(n6505));
  jnot g06314(.din(n6505), .dout(n6506));
  jand g06315(.dina(\a[52] ), .dinb(\a[5] ), .dout(n6507));
  jnot g06316(.din(n6507), .dout(n6508));
  jand g06317(.dina(\a[38] ), .dinb(\a[20] ), .dout(n6509));
  jand g06318(.dina(n6509), .dinb(n6311), .dout(n6510));
  jnot g06319(.din(n6510), .dout(n6511));
  jand g06320(.dina(\a[37] ), .dinb(\a[20] ), .dout(n6512));
  jand g06321(.dina(\a[38] ), .dinb(\a[19] ), .dout(n6513));
  jor  g06322(.dina(n6513), .dinb(n6512), .dout(n6514));
  jand g06323(.dina(n6514), .dinb(n6511), .dout(n6515));
  jxor g06324(.dina(n6515), .dinb(n6508), .dout(n6516));
  jxor g06325(.dina(n6516), .dinb(n6506), .dout(n6517));
  jnot g06326(.din(n6517), .dout(n6518));
  jand g06327(.dina(\a[42] ), .dinb(\a[15] ), .dout(n6519));
  jnot g06328(.din(n6519), .dout(n6520));
  jand g06329(.dina(n5316), .dinb(n453), .dout(n6521));
  jnot g06330(.din(n6521), .dout(n6522));
  jand g06331(.dina(\a[48] ), .dinb(\a[9] ), .dout(n6523));
  jor  g06332(.dina(n6523), .dinb(n6262), .dout(n6524));
  jand g06333(.dina(n6524), .dinb(n6522), .dout(n6525));
  jxor g06334(.dina(n6525), .dinb(n6520), .dout(n6526));
  jxor g06335(.dina(n6526), .dinb(n6518), .dout(n6527));
  jand g06336(.dina(\a[44] ), .dinb(\a[13] ), .dout(n6528));
  jand g06337(.dina(\a[46] ), .dinb(\a[11] ), .dout(n6529));
  jor  g06338(.dina(n6529), .dinb(n6528), .dout(n6530));
  jand g06339(.dina(\a[46] ), .dinb(\a[44] ), .dout(n6531));
  jand g06340(.dina(n6531), .dinb(n816), .dout(n6532));
  jnot g06341(.din(n6532), .dout(n6533));
  jand g06342(.dina(n4495), .dinb(n675), .dout(n6534));
  jand g06343(.dina(\a[43] ), .dinb(\a[14] ), .dout(n6535));
  jand g06344(.dina(n6535), .dinb(n6529), .dout(n6536));
  jor  g06345(.dina(n6536), .dinb(n6534), .dout(n6537));
  jnot g06346(.din(n6537), .dout(n6538));
  jand g06347(.dina(n6538), .dinb(n6533), .dout(n6539));
  jand g06348(.dina(n6539), .dinb(n6530), .dout(n6540));
  jand g06349(.dina(n6537), .dinb(n6533), .dout(n6541));
  jnot g06350(.din(n6541), .dout(n6542));
  jand g06351(.dina(n6542), .dinb(n6535), .dout(n6543));
  jor  g06352(.dina(n6543), .dinb(n6540), .dout(n6544));
  jand g06353(.dina(\a[45] ), .dinb(\a[12] ), .dout(n6545));
  jnot g06354(.din(n6545), .dout(n6546));
  jand g06355(.dina(n3294), .dinb(n2042), .dout(n6547));
  jnot g06356(.din(n6547), .dout(n6548));
  jand g06357(.dina(\a[30] ), .dinb(\a[27] ), .dout(n6549));
  jor  g06358(.dina(n6549), .dinb(n2653), .dout(n6550));
  jand g06359(.dina(n6550), .dinb(n6548), .dout(n6551));
  jxor g06360(.dina(n6551), .dinb(n6546), .dout(n6552));
  jnot g06361(.din(n6552), .dout(n6553));
  jxor g06362(.dina(n6553), .dinb(n6544), .dout(n6554));
  jand g06363(.dina(\a[39] ), .dinb(\a[18] ), .dout(n6555));
  jand g06364(.dina(\a[51] ), .dinb(\a[6] ), .dout(n6556));
  jand g06365(.dina(\a[40] ), .dinb(\a[17] ), .dout(n6557));
  jxor g06366(.dina(n6557), .dinb(n6556), .dout(n6558));
  jxor g06367(.dina(n6558), .dinb(n6555), .dout(n6559));
  jxor g06368(.dina(n6559), .dinb(n6554), .dout(n6560));
  jxor g06369(.dina(n6560), .dinb(n6527), .dout(n6561));
  jxor g06370(.dina(n6561), .dinb(n6496), .dout(n6562));
  jand g06371(.dina(n6417), .dinb(n6414), .dout(n6563));
  jand g06372(.dina(n6418), .dinb(n6394), .dout(n6564));
  jor  g06373(.dina(n6564), .dinb(n6563), .dout(n6565));
  jand g06374(.dina(n6406), .dinb(n6403), .dout(n6566));
  jnot g06375(.din(n6566), .dout(n6567));
  jand g06376(.dina(n6567), .dinb(n6409), .dout(n6568));
  jxor g06377(.dina(n6568), .dinb(n6269), .dout(n6569));
  jand g06378(.dina(n6244), .dinb(n6242), .dout(n6570));
  jnot g06379(.din(n6570), .dout(n6571));
  jand g06380(.dina(n6571), .dinb(n6247), .dout(n6572));
  jxor g06381(.dina(n6572), .dinb(n6569), .dout(n6573));
  jand g06382(.dina(n6412), .dinb(n6401), .dout(n6574));
  jand g06383(.dina(n6413), .dinb(n6397), .dout(n6575));
  jor  g06384(.dina(n6575), .dinb(n6574), .dout(n6576));
  jxor g06385(.dina(n6576), .dinb(n6573), .dout(n6577));
  jand g06386(.dina(\a[49] ), .dinb(\a[8] ), .dout(n6578));
  jand g06387(.dina(\a[41] ), .dinb(\a[16] ), .dout(n6579));
  jand g06388(.dina(n6579), .dinb(n6578), .dout(n6580));
  jnot g06389(.din(n6580), .dout(n6581));
  jand g06390(.dina(\a[50] ), .dinb(\a[8] ), .dout(n6582));
  jand g06391(.dina(n6582), .dinb(n6220), .dout(n6583));
  jand g06392(.dina(n6579), .dinb(n6227), .dout(n6584));
  jor  g06393(.dina(n6584), .dinb(n6583), .dout(n6585));
  jnot g06394(.din(n6585), .dout(n6586));
  jand g06395(.dina(n6586), .dinb(n6581), .dout(n6587));
  jor  g06396(.dina(n6579), .dinb(n6578), .dout(n6588));
  jand g06397(.dina(n6588), .dinb(n6587), .dout(n6589));
  jand g06398(.dina(n6585), .dinb(n6581), .dout(n6590));
  jnot g06399(.din(n6590), .dout(n6591));
  jand g06400(.dina(n6591), .dinb(n6227), .dout(n6592));
  jor  g06401(.dina(n6592), .dinb(n6589), .dout(n6593));
  jand g06402(.dina(\a[36] ), .dinb(\a[21] ), .dout(n6594));
  jnot g06403(.din(n6594), .dout(n6595));
  jand g06404(.dina(n2845), .dinb(n1658), .dout(n6596));
  jnot g06405(.din(n6596), .dout(n6597));
  jand g06406(.dina(\a[35] ), .dinb(\a[22] ), .dout(n6598));
  jand g06407(.dina(\a[34] ), .dinb(\a[23] ), .dout(n6599));
  jor  g06408(.dina(n6599), .dinb(n6598), .dout(n6600));
  jand g06409(.dina(n6600), .dinb(n6597), .dout(n6601));
  jxor g06410(.dina(n6601), .dinb(n6595), .dout(n6602));
  jnot g06411(.din(n6602), .dout(n6603));
  jxor g06412(.dina(n6603), .dinb(n6593), .dout(n6604));
  jnot g06413(.din(n6604), .dout(n6605));
  jand g06414(.dina(\a[33] ), .dinb(\a[24] ), .dout(n6606));
  jnot g06415(.din(n6606), .dout(n6607));
  jand g06416(.dina(n3269), .dinb(n2128), .dout(n6608));
  jnot g06417(.din(n6608), .dout(n6609));
  jand g06418(.dina(\a[31] ), .dinb(\a[26] ), .dout(n6610));
  jand g06419(.dina(\a[32] ), .dinb(\a[25] ), .dout(n6611));
  jor  g06420(.dina(n6611), .dinb(n6610), .dout(n6612));
  jand g06421(.dina(n6612), .dinb(n6609), .dout(n6613));
  jxor g06422(.dina(n6613), .dinb(n6607), .dout(n6614));
  jxor g06423(.dina(n6614), .dinb(n6605), .dout(n6615));
  jxor g06424(.dina(n6615), .dinb(n6577), .dout(n6616));
  jxor g06425(.dina(n6616), .dinb(n6565), .dout(n6617));
  jxor g06426(.dina(n6617), .dinb(n6562), .dout(n6618));
  jxor g06427(.dina(n6618), .dinb(n6492), .dout(n6619));
  jand g06428(.dina(n6387), .dinb(n6351), .dout(n6620));
  jand g06429(.dina(n6388), .dinb(n6348), .dout(n6621));
  jor  g06430(.dina(n6621), .dinb(n6620), .dout(n6622));
  jand g06431(.dina(n6346), .dinb(n6320), .dout(n6623));
  jand g06432(.dina(n6347), .dinb(n6315), .dout(n6624));
  jor  g06433(.dina(n6624), .dinb(n6623), .dout(n6625));
  jand g06434(.dina(n6385), .dinb(n6382), .dout(n6626));
  jand g06435(.dina(n6386), .dinb(n6368), .dout(n6627));
  jor  g06436(.dina(n6627), .dinb(n6626), .dout(n6628));
  jand g06437(.dina(n6363), .dinb(n6360), .dout(n6629));
  jand g06438(.dina(n6367), .dinb(n6364), .dout(n6630));
  jor  g06439(.dina(n6630), .dinb(n6629), .dout(n6631));
  jand g06440(.dina(n6344), .dinb(n6336), .dout(n6632));
  jand g06441(.dina(n6345), .dinb(n6331), .dout(n6633));
  jor  g06442(.dina(n6633), .dinb(n6632), .dout(n6634));
  jxor g06443(.dina(n6634), .dinb(n6631), .dout(n6635));
  jand g06444(.dina(n6329), .dinb(n6326), .dout(n6636));
  jand g06445(.dina(n6330), .dinb(n6323), .dout(n6637));
  jor  g06446(.dina(n6637), .dinb(n6636), .dout(n6638));
  jand g06447(.dina(n6341), .dinb(n2536), .dout(n6639));
  jand g06448(.dina(\a[57] ), .dinb(\a[0] ), .dout(n6640));
  jxor g06449(.dina(n6640), .dinb(n6639), .dout(n6641));
  jand g06450(.dina(\a[56] ), .dinb(\a[1] ), .dout(n6642));
  jxor g06451(.dina(n6642), .dinb(\a[29] ), .dout(n6643));
  jxor g06452(.dina(n6643), .dinb(n6641), .dout(n6644));
  jxor g06453(.dina(n6644), .dinb(n6638), .dout(n6645));
  jand g06454(.dina(n6354), .dinb(n6137), .dout(n6646));
  jand g06455(.dina(n6359), .dinb(n6355), .dout(n6647));
  jor  g06456(.dina(n6647), .dinb(n6646), .dout(n6648));
  jxor g06457(.dina(n6648), .dinb(n6645), .dout(n6649));
  jxor g06458(.dina(n6649), .dinb(n6635), .dout(n6650));
  jxor g06459(.dina(n6650), .dinb(n6628), .dout(n6651));
  jxor g06460(.dina(n6651), .dinb(n6625), .dout(n6652));
  jxor g06461(.dina(n6652), .dinb(n6622), .dout(n6653));
  jxor g06462(.dina(n6653), .dinb(n6619), .dout(n6654));
  jand g06463(.dina(n6654), .dinb(n6443), .dout(n6655));
  jor  g06464(.dina(n6654), .dinb(n6443), .dout(n6656));
  jnot g06465(.din(n6656), .dout(n6657));
  jor  g06466(.dina(n6657), .dinb(n6655), .dout(n6658));
  jnot g06467(.din(n6433), .dout(n6659));
  jor  g06468(.dina(n6439), .dinb(n6435), .dout(n6660));
  jand g06469(.dina(n6660), .dinb(n6659), .dout(n6661));
  jxor g06470(.dina(n6661), .dinb(n6658), .dout(\asquared[58] ));
  jand g06471(.dina(n6652), .dinb(n6622), .dout(n6663));
  jand g06472(.dina(n6653), .dinb(n6619), .dout(n6664));
  jor  g06473(.dina(n6664), .dinb(n6663), .dout(n6665));
  jand g06474(.dina(n6491), .dinb(n6446), .dout(n6666));
  jand g06475(.dina(n6618), .dinb(n6492), .dout(n6667));
  jor  g06476(.dina(n6667), .dinb(n6666), .dout(n6668));
  jand g06477(.dina(n6464), .dinb(n6461), .dout(n6669));
  jand g06478(.dina(n6490), .dinb(n6465), .dout(n6670));
  jor  g06479(.dina(n6670), .dinb(n6669), .dout(n6671));
  jand g06480(.dina(n6576), .dinb(n6573), .dout(n6672));
  jand g06481(.dina(n6615), .dinb(n6577), .dout(n6673));
  jor  g06482(.dina(n6673), .dinb(n6672), .dout(n6674));
  jand g06483(.dina(n6568), .dinb(n6269), .dout(n6675));
  jand g06484(.dina(n6572), .dinb(n6569), .dout(n6676));
  jor  g06485(.dina(n6676), .dinb(n6675), .dout(n6677));
  jand g06486(.dina(n6484), .dinb(n6480), .dout(n6678));
  jand g06487(.dina(n6487), .dinb(n6485), .dout(n6679));
  jor  g06488(.dina(n6679), .dinb(n6678), .dout(n6680));
  jxor g06489(.dina(n6680), .dinb(n6677), .dout(n6681));
  jand g06490(.dina(n6476), .dinb(n6473), .dout(n6682));
  jand g06491(.dina(n6477), .dinb(n6234), .dout(n6683));
  jor  g06492(.dina(n6683), .dinb(n6682), .dout(n6684));
  jxor g06493(.dina(n6684), .dinb(n6681), .dout(n6685));
  jand g06494(.dina(n6488), .dinb(n6478), .dout(n6686));
  jand g06495(.dina(n6489), .dinb(n6470), .dout(n6687));
  jor  g06496(.dina(n6687), .dinb(n6686), .dout(n6688));
  jxor g06497(.dina(n6688), .dinb(n6685), .dout(n6689));
  jxor g06498(.dina(n6689), .dinb(n6674), .dout(n6690));
  jxor g06499(.dina(n6690), .dinb(n6671), .dout(n6691));
  jand g06500(.dina(n6616), .dinb(n6565), .dout(n6692));
  jand g06501(.dina(n6617), .dinb(n6562), .dout(n6693));
  jor  g06502(.dina(n6693), .dinb(n6692), .dout(n6694));
  jxor g06503(.dina(n6694), .dinb(n6691), .dout(n6695));
  jxor g06504(.dina(n6695), .dinb(n6668), .dout(n6696));
  jand g06505(.dina(n6650), .dinb(n6628), .dout(n6697));
  jand g06506(.dina(n6651), .dinb(n6625), .dout(n6698));
  jor  g06507(.dina(n6698), .dinb(n6697), .dout(n6699));
  jand g06508(.dina(n6560), .dinb(n6527), .dout(n6700));
  jand g06509(.dina(n6561), .dinb(n6496), .dout(n6701));
  jor  g06510(.dina(n6701), .dinb(n6700), .dout(n6702));
  jand g06511(.dina(n6553), .dinb(n6544), .dout(n6703));
  jand g06512(.dina(n6559), .dinb(n6554), .dout(n6704));
  jor  g06513(.dina(n6704), .dinb(n6703), .dout(n6705));
  jor  g06514(.dina(n6516), .dinb(n6506), .dout(n6706));
  jor  g06515(.dina(n6526), .dinb(n6518), .dout(n6707));
  jand g06516(.dina(n6707), .dinb(n6706), .dout(n6708));
  jnot g06517(.din(n6708), .dout(n6709));
  jand g06518(.dina(n6642), .dinb(\a[29] ), .dout(n6710));
  jand g06519(.dina(\a[57] ), .dinb(\a[1] ), .dout(n6711));
  jxor g06520(.dina(n6711), .dinb(n2810), .dout(n6712));
  jxor g06521(.dina(n6712), .dinb(n6710), .dout(n6713));
  jand g06522(.dina(n6548), .dinb(n6546), .dout(n6714));
  jnot g06523(.din(n6714), .dout(n6715));
  jand g06524(.dina(n6715), .dinb(n6550), .dout(n6716));
  jxor g06525(.dina(n6716), .dinb(n6713), .dout(n6717));
  jxor g06526(.dina(n6717), .dinb(n6709), .dout(n6718));
  jxor g06527(.dina(n6718), .dinb(n6705), .dout(n6719));
  jxor g06528(.dina(n6719), .dinb(n6702), .dout(n6720));
  jand g06529(.dina(n6603), .dinb(n6593), .dout(n6721));
  jnot g06530(.din(n6721), .dout(n6722));
  jor  g06531(.dina(n6614), .dinb(n6605), .dout(n6723));
  jand g06532(.dina(n6723), .dinb(n6722), .dout(n6724));
  jnot g06533(.din(n6724), .dout(n6725));
  jand g06534(.dina(n6522), .dinb(n6520), .dout(n6726));
  jnot g06535(.din(n6726), .dout(n6727));
  jand g06536(.dina(n6727), .dinb(n6524), .dout(n6728));
  jand g06537(.dina(n6609), .dinb(n6607), .dout(n6729));
  jnot g06538(.din(n6729), .dout(n6730));
  jand g06539(.dina(n6730), .dinb(n6612), .dout(n6731));
  jxor g06540(.dina(n6731), .dinb(n6728), .dout(n6732));
  jand g06541(.dina(n6597), .dinb(n6595), .dout(n6733));
  jnot g06542(.din(n6733), .dout(n6734));
  jand g06543(.dina(n6734), .dinb(n6600), .dout(n6735));
  jxor g06544(.dina(n6735), .dinb(n6732), .dout(n6736));
  jnot g06545(.din(n6539), .dout(n6737));
  jand g06546(.dina(n6504), .dinb(n6497), .dout(n6738));
  jor  g06547(.dina(n6738), .dinb(n6499), .dout(n6739));
  jand g06548(.dina(n6511), .dinb(n6508), .dout(n6740));
  jnot g06549(.din(n6740), .dout(n6741));
  jand g06550(.dina(n6741), .dinb(n6514), .dout(n6742));
  jxor g06551(.dina(n6742), .dinb(n6739), .dout(n6743));
  jxor g06552(.dina(n6743), .dinb(n6737), .dout(n6744));
  jxor g06553(.dina(n6744), .dinb(n6736), .dout(n6745));
  jxor g06554(.dina(n6745), .dinb(n6725), .dout(n6746));
  jxor g06555(.dina(n6746), .dinb(n6720), .dout(n6747));
  jxor g06556(.dina(n6747), .dinb(n6699), .dout(n6748));
  jor  g06557(.dina(n6454), .dinb(n6450), .dout(n6749));
  jor  g06558(.dina(n6460), .dinb(n6456), .dout(n6750));
  jand g06559(.dina(n6750), .dinb(n6749), .dout(n6751));
  jnot g06560(.din(n6751), .dout(n6752));
  jand g06561(.dina(\a[41] ), .dinb(\a[17] ), .dout(n6753));
  jand g06562(.dina(\a[49] ), .dinb(\a[42] ), .dout(n6754));
  jand g06563(.dina(n6754), .dinb(n1367), .dout(n6755));
  jnot g06564(.din(n6755), .dout(n6756));
  jand g06565(.dina(n4514), .dinb(n937), .dout(n6757));
  jand g06566(.dina(\a[49] ), .dinb(\a[9] ), .dout(n6758));
  jand g06567(.dina(n6758), .dinb(n6753), .dout(n6759));
  jor  g06568(.dina(n6759), .dinb(n6757), .dout(n6760));
  jand g06569(.dina(n6760), .dinb(n6756), .dout(n6761));
  jnot g06570(.din(n6761), .dout(n6762));
  jand g06571(.dina(n6762), .dinb(n6753), .dout(n6763));
  jand g06572(.dina(\a[42] ), .dinb(\a[16] ), .dout(n6764));
  jor  g06573(.dina(n6764), .dinb(n6758), .dout(n6765));
  jor  g06574(.dina(n6760), .dinb(n6755), .dout(n6766));
  jnot g06575(.din(n6766), .dout(n6767));
  jand g06576(.dina(n6767), .dinb(n6765), .dout(n6768));
  jor  g06577(.dina(n6768), .dinb(n6763), .dout(n6769));
  jand g06578(.dina(\a[58] ), .dinb(\a[0] ), .dout(n6770));
  jand g06579(.dina(\a[54] ), .dinb(\a[4] ), .dout(n6771));
  jxor g06580(.dina(n6771), .dinb(n6770), .dout(n6772));
  jxor g06581(.dina(n6772), .dinb(n6295), .dout(n6773));
  jand g06582(.dina(\a[53] ), .dinb(\a[5] ), .dout(n6774));
  jand g06583(.dina(\a[38] ), .dinb(\a[21] ), .dout(n6775));
  jand g06584(.dina(n6775), .dinb(n6512), .dout(n6776));
  jnot g06585(.din(n6776), .dout(n6777));
  jand g06586(.dina(\a[37] ), .dinb(\a[21] ), .dout(n6778));
  jor  g06587(.dina(n6778), .dinb(n6509), .dout(n6779));
  jand g06588(.dina(n6779), .dinb(n6777), .dout(n6780));
  jxor g06589(.dina(n6780), .dinb(n6774), .dout(n6781));
  jxor g06590(.dina(n6781), .dinb(n6773), .dout(n6782));
  jxor g06591(.dina(n6782), .dinb(n6769), .dout(n6783));
  jand g06592(.dina(\a[40] ), .dinb(\a[18] ), .dout(n6784));
  jand g06593(.dina(\a[51] ), .dinb(\a[7] ), .dout(n6785));
  jor  g06594(.dina(n6785), .dinb(n6582), .dout(n6786));
  jand g06595(.dina(n5594), .dinb(n499), .dout(n6787));
  jnot g06596(.din(n6787), .dout(n6788));
  jand g06597(.dina(n6788), .dinb(n6786), .dout(n6789));
  jxor g06598(.dina(n6789), .dinb(n6784), .dout(n6790));
  jand g06599(.dina(\a[36] ), .dinb(\a[22] ), .dout(n6791));
  jand g06600(.dina(n2845), .dinb(n1942), .dout(n6792));
  jnot g06601(.din(n6792), .dout(n6793));
  jand g06602(.dina(\a[35] ), .dinb(\a[23] ), .dout(n6794));
  jand g06603(.dina(\a[34] ), .dinb(\a[24] ), .dout(n6795));
  jor  g06604(.dina(n6795), .dinb(n6794), .dout(n6796));
  jand g06605(.dina(n6796), .dinb(n6793), .dout(n6797));
  jxor g06606(.dina(n6797), .dinb(n6791), .dout(n6798));
  jxor g06607(.dina(n6798), .dinb(n6790), .dout(n6799));
  jnot g06608(.din(n6799), .dout(n6800));
  jnot g06609(.din(n2824), .dout(n6801));
  jand g06610(.dina(n3269), .dinb(n1927), .dout(n6802));
  jnot g06611(.din(n6802), .dout(n6803));
  jand g06612(.dina(\a[31] ), .dinb(\a[27] ), .dout(n6804));
  jand g06613(.dina(\a[32] ), .dinb(\a[26] ), .dout(n6805));
  jor  g06614(.dina(n6805), .dinb(n6804), .dout(n6806));
  jand g06615(.dina(n6806), .dinb(n6803), .dout(n6807));
  jxor g06616(.dina(n6807), .dinb(n6801), .dout(n6808));
  jxor g06617(.dina(n6808), .dinb(n6800), .dout(n6809));
  jxor g06618(.dina(n6809), .dinb(n6783), .dout(n6810));
  jxor g06619(.dina(n6810), .dinb(n6752), .dout(n6811));
  jand g06620(.dina(n6634), .dinb(n6631), .dout(n6812));
  jand g06621(.dina(n6649), .dinb(n6635), .dout(n6813));
  jor  g06622(.dina(n6813), .dinb(n6812), .dout(n6814));
  jnot g06623(.din(n6587), .dout(n6815));
  jand g06624(.dina(n6557), .dinb(n6556), .dout(n6816));
  jand g06625(.dina(n6558), .dinb(n6555), .dout(n6817));
  jor  g06626(.dina(n6817), .dinb(n6816), .dout(n6818));
  jxor g06627(.dina(n6818), .dinb(n6815), .dout(n6819));
  jand g06628(.dina(n6640), .dinb(n6639), .dout(n6820));
  jand g06629(.dina(n6643), .dinb(n6641), .dout(n6821));
  jor  g06630(.dina(n6821), .dinb(n6820), .dout(n6822));
  jxor g06631(.dina(n6822), .dinb(n6819), .dout(n6823));
  jand g06632(.dina(n6644), .dinb(n6638), .dout(n6824));
  jand g06633(.dina(n6648), .dinb(n6645), .dout(n6825));
  jor  g06634(.dina(n6825), .dinb(n6824), .dout(n6826));
  jxor g06635(.dina(n6826), .dinb(n6823), .dout(n6827));
  jand g06636(.dina(\a[47] ), .dinb(\a[43] ), .dout(n6828));
  jand g06637(.dina(n6828), .dinb(n1469), .dout(n6829));
  jnot g06638(.din(n6829), .dout(n6830));
  jand g06639(.dina(n5316), .dinb(n655), .dout(n6831));
  jand g06640(.dina(\a[43] ), .dinb(\a[15] ), .dout(n6832));
  jand g06641(.dina(\a[48] ), .dinb(\a[10] ), .dout(n6833));
  jand g06642(.dina(n6833), .dinb(n6832), .dout(n6834));
  jor  g06643(.dina(n6834), .dinb(n6831), .dout(n6835));
  jnot g06644(.din(n6835), .dout(n6836));
  jand g06645(.dina(n6836), .dinb(n6830), .dout(n6837));
  jand g06646(.dina(\a[47] ), .dinb(\a[11] ), .dout(n6838));
  jor  g06647(.dina(n6838), .dinb(n6832), .dout(n6839));
  jand g06648(.dina(n6839), .dinb(n6837), .dout(n6840));
  jand g06649(.dina(n6835), .dinb(n6830), .dout(n6841));
  jnot g06650(.din(n6841), .dout(n6842));
  jand g06651(.dina(n6842), .dinb(n6833), .dout(n6843));
  jor  g06652(.dina(n6843), .dinb(n6840), .dout(n6844));
  jand g06653(.dina(\a[44] ), .dinb(\a[14] ), .dout(n6845));
  jnot g06654(.din(n6845), .dout(n6846));
  jand g06655(.dina(\a[46] ), .dinb(\a[13] ), .dout(n6847));
  jand g06656(.dina(n6847), .dinb(n6545), .dout(n6848));
  jnot g06657(.din(n6848), .dout(n6849));
  jand g06658(.dina(\a[45] ), .dinb(\a[13] ), .dout(n6850));
  jand g06659(.dina(\a[46] ), .dinb(\a[12] ), .dout(n6851));
  jor  g06660(.dina(n6851), .dinb(n6850), .dout(n6852));
  jand g06661(.dina(n6852), .dinb(n6849), .dout(n6853));
  jxor g06662(.dina(n6853), .dinb(n6846), .dout(n6854));
  jnot g06663(.din(n6854), .dout(n6855));
  jxor g06664(.dina(n6855), .dinb(n6844), .dout(n6856));
  jand g06665(.dina(\a[55] ), .dinb(\a[3] ), .dout(n6857));
  jand g06666(.dina(\a[52] ), .dinb(\a[6] ), .dout(n6858));
  jand g06667(.dina(\a[39] ), .dinb(\a[19] ), .dout(n6859));
  jxor g06668(.dina(n6859), .dinb(n6858), .dout(n6860));
  jxor g06669(.dina(n6860), .dinb(n6857), .dout(n6861));
  jxor g06670(.dina(n6861), .dinb(n6856), .dout(n6862));
  jxor g06671(.dina(n6862), .dinb(n6827), .dout(n6863));
  jxor g06672(.dina(n6863), .dinb(n6814), .dout(n6864));
  jxor g06673(.dina(n6864), .dinb(n6811), .dout(n6865));
  jxor g06674(.dina(n6865), .dinb(n6748), .dout(n6866));
  jxor g06675(.dina(n6866), .dinb(n6696), .dout(n6867));
  jand g06676(.dina(n6867), .dinb(n6665), .dout(n6868));
  jor  g06677(.dina(n6867), .dinb(n6665), .dout(n6869));
  jnot g06678(.din(n6869), .dout(n6870));
  jor  g06679(.dina(n6870), .dinb(n6868), .dout(n6871));
  jnot g06680(.din(n6655), .dout(n6872));
  jor  g06681(.dina(n6661), .dinb(n6657), .dout(n6873));
  jand g06682(.dina(n6873), .dinb(n6872), .dout(n6874));
  jxor g06683(.dina(n6874), .dinb(n6871), .dout(\asquared[59] ));
  jand g06684(.dina(n6747), .dinb(n6699), .dout(n6876));
  jand g06685(.dina(n6865), .dinb(n6748), .dout(n6877));
  jor  g06686(.dina(n6877), .dinb(n6876), .dout(n6878));
  jand g06687(.dina(n6863), .dinb(n6814), .dout(n6879));
  jand g06688(.dina(n6864), .dinb(n6811), .dout(n6880));
  jor  g06689(.dina(n6880), .dinb(n6879), .dout(n6881));
  jand g06690(.dina(n6719), .dinb(n6702), .dout(n6882));
  jand g06691(.dina(n6746), .dinb(n6720), .dout(n6883));
  jor  g06692(.dina(n6883), .dinb(n6882), .dout(n6884));
  jand g06693(.dina(n6826), .dinb(n6823), .dout(n6885));
  jand g06694(.dina(n6862), .dinb(n6827), .dout(n6886));
  jor  g06695(.dina(n6886), .dinb(n6885), .dout(n6887));
  jand g06696(.dina(n6818), .dinb(n6815), .dout(n6888));
  jand g06697(.dina(n6822), .dinb(n6819), .dout(n6889));
  jor  g06698(.dina(n6889), .dinb(n6888), .dout(n6890));
  jand g06699(.dina(n6742), .dinb(n6739), .dout(n6891));
  jand g06700(.dina(n6743), .dinb(n6737), .dout(n6892));
  jor  g06701(.dina(n6892), .dinb(n6891), .dout(n6893));
  jxor g06702(.dina(n6893), .dinb(n6890), .dout(n6894));
  jand g06703(.dina(n6731), .dinb(n6728), .dout(n6895));
  jand g06704(.dina(n6735), .dinb(n6732), .dout(n6896));
  jor  g06705(.dina(n6896), .dinb(n6895), .dout(n6897));
  jxor g06706(.dina(n6897), .dinb(n6894), .dout(n6898));
  jand g06707(.dina(n6744), .dinb(n6736), .dout(n6899));
  jand g06708(.dina(n6745), .dinb(n6725), .dout(n6900));
  jor  g06709(.dina(n6900), .dinb(n6899), .dout(n6901));
  jxor g06710(.dina(n6901), .dinb(n6898), .dout(n6902));
  jxor g06711(.dina(n6902), .dinb(n6887), .dout(n6903));
  jxor g06712(.dina(n6903), .dinb(n6884), .dout(n6904));
  jxor g06713(.dina(n6904), .dinb(n6881), .dout(n6905));
  jxor g06714(.dina(n6905), .dinb(n6878), .dout(n6906));
  jand g06715(.dina(n6690), .dinb(n6671), .dout(n6907));
  jand g06716(.dina(n6694), .dinb(n6691), .dout(n6908));
  jor  g06717(.dina(n6908), .dinb(n6907), .dout(n6909));
  jand g06718(.dina(n6855), .dinb(n6844), .dout(n6910));
  jand g06719(.dina(n6861), .dinb(n6856), .dout(n6911));
  jor  g06720(.dina(n6911), .dinb(n6910), .dout(n6912));
  jnot g06721(.din(n6912), .dout(n6913));
  jand g06722(.dina(n6798), .dinb(n6790), .dout(n6914));
  jnot g06723(.din(n6914), .dout(n6915));
  jor  g06724(.dina(n6808), .dinb(n6800), .dout(n6916));
  jand g06725(.dina(n6916), .dinb(n6915), .dout(n6917));
  jxor g06726(.dina(n6917), .dinb(n6913), .dout(n6918));
  jand g06727(.dina(n6781), .dinb(n6773), .dout(n6919));
  jand g06728(.dina(n6782), .dinb(n6769), .dout(n6920));
  jor  g06729(.dina(n6920), .dinb(n6919), .dout(n6921));
  jxor g06730(.dina(n6921), .dinb(n6918), .dout(n6922));
  jand g06731(.dina(n6809), .dinb(n6783), .dout(n6923));
  jand g06732(.dina(n6810), .dinb(n6752), .dout(n6924));
  jor  g06733(.dina(n6924), .dinb(n6923), .dout(n6925));
  jand g06734(.dina(n6771), .dinb(n6770), .dout(n6926));
  jand g06735(.dina(n6772), .dinb(n6295), .dout(n6927));
  jor  g06736(.dina(n6927), .dinb(n6926), .dout(n6928));
  jand g06737(.dina(n6859), .dinb(n6858), .dout(n6929));
  jand g06738(.dina(n6860), .dinb(n6857), .dout(n6930));
  jor  g06739(.dina(n6930), .dinb(n6929), .dout(n6931));
  jxor g06740(.dina(n6931), .dinb(n6928), .dout(n6932));
  jxor g06741(.dina(n6932), .dinb(n6766), .dout(n6933));
  jand g06742(.dina(n6789), .dinb(n6784), .dout(n6934));
  jor  g06743(.dina(n6934), .dinb(n6787), .dout(n6935));
  jand g06744(.dina(n6779), .dinb(n6774), .dout(n6936));
  jor  g06745(.dina(n6936), .dinb(n6776), .dout(n6937));
  jor  g06746(.dina(n6792), .dinb(n6791), .dout(n6938));
  jand g06747(.dina(n6938), .dinb(n6796), .dout(n6939));
  jxor g06748(.dina(n6939), .dinb(n6937), .dout(n6940));
  jxor g06749(.dina(n6940), .dinb(n6935), .dout(n6941));
  jnot g06750(.din(n6837), .dout(n6942));
  jand g06751(.dina(n2064), .dinb(\a[58] ), .dout(n6943));
  jnot g06752(.din(n6943), .dout(n6944));
  jand g06753(.dina(\a[58] ), .dinb(\a[1] ), .dout(n6945));
  jor  g06754(.dina(n6945), .dinb(\a[30] ), .dout(n6946));
  jand g06755(.dina(n6946), .dinb(n6944), .dout(n6947));
  jand g06756(.dina(n6849), .dinb(n6846), .dout(n6948));
  jnot g06757(.din(n6948), .dout(n6949));
  jand g06758(.dina(n6949), .dinb(n6852), .dout(n6950));
  jxor g06759(.dina(n6950), .dinb(n6947), .dout(n6951));
  jxor g06760(.dina(n6951), .dinb(n6942), .dout(n6952));
  jxor g06761(.dina(n6952), .dinb(n6941), .dout(n6953));
  jxor g06762(.dina(n6953), .dinb(n6933), .dout(n6954));
  jxor g06763(.dina(n6954), .dinb(n6925), .dout(n6955));
  jxor g06764(.dina(n6955), .dinb(n6922), .dout(n6956));
  jxor g06765(.dina(n6956), .dinb(n6909), .dout(n6957));
  jand g06766(.dina(n6688), .dinb(n6685), .dout(n6958));
  jand g06767(.dina(n6689), .dinb(n6674), .dout(n6959));
  jor  g06768(.dina(n6959), .dinb(n6958), .dout(n6960));
  jand g06769(.dina(n6717), .dinb(n6709), .dout(n6961));
  jand g06770(.dina(n6718), .dinb(n6705), .dout(n6962));
  jor  g06771(.dina(n6962), .dinb(n6961), .dout(n6963));
  jand g06772(.dina(\a[55] ), .dinb(\a[4] ), .dout(n6964));
  jand g06773(.dina(\a[55] ), .dinb(\a[5] ), .dout(n6965));
  jand g06774(.dina(n6965), .dinb(n6771), .dout(n6966));
  jand g06775(.dina(\a[40] ), .dinb(\a[19] ), .dout(n6967));
  jand g06776(.dina(n6967), .dinb(n6964), .dout(n6968));
  jor  g06777(.dina(n6968), .dinb(n6966), .dout(n6969));
  jand g06778(.dina(\a[54] ), .dinb(\a[5] ), .dout(n6970));
  jand g06779(.dina(n6970), .dinb(n6967), .dout(n6971));
  jnot g06780(.din(n6971), .dout(n6972));
  jand g06781(.dina(n6972), .dinb(n6969), .dout(n6973));
  jnot g06782(.din(n6973), .dout(n6974));
  jand g06783(.dina(n6974), .dinb(n6964), .dout(n6975));
  jor  g06784(.dina(n6971), .dinb(n6969), .dout(n6976));
  jnot g06785(.din(n6976), .dout(n6977));
  jor  g06786(.dina(n6970), .dinb(n6967), .dout(n6978));
  jand g06787(.dina(n6978), .dinb(n6977), .dout(n6979));
  jor  g06788(.dina(n6979), .dinb(n6975), .dout(n6980));
  jand g06789(.dina(n6711), .dinb(n2810), .dout(n6981));
  jand g06790(.dina(\a[57] ), .dinb(\a[2] ), .dout(n6982));
  jand g06791(.dina(\a[56] ), .dinb(\a[3] ), .dout(n6983));
  jor  g06792(.dina(n6983), .dinb(n6982), .dout(n6984));
  jand g06793(.dina(\a[57] ), .dinb(\a[3] ), .dout(n6985));
  jand g06794(.dina(n6985), .dinb(n6295), .dout(n6986));
  jnot g06795(.din(n6986), .dout(n6987));
  jand g06796(.dina(n6987), .dinb(n6984), .dout(n6988));
  jxor g06797(.dina(n6988), .dinb(n6981), .dout(n6989));
  jand g06798(.dina(n6803), .dinb(n6801), .dout(n6990));
  jnot g06799(.din(n6990), .dout(n6991));
  jand g06800(.dina(n6991), .dinb(n6806), .dout(n6992));
  jxor g06801(.dina(n6992), .dinb(n6989), .dout(n6993));
  jxor g06802(.dina(n6993), .dinb(n6980), .dout(n6994));
  jand g06803(.dina(\a[48] ), .dinb(\a[11] ), .dout(n6995));
  jand g06804(.dina(\a[47] ), .dinb(\a[45] ), .dout(n6996));
  jand g06805(.dina(n6996), .dinb(n979), .dout(n6997));
  jnot g06806(.din(n6997), .dout(n6998));
  jand g06807(.dina(\a[47] ), .dinb(\a[12] ), .dout(n6999));
  jand g06808(.dina(\a[45] ), .dinb(\a[14] ), .dout(n7000));
  jor  g06809(.dina(n7000), .dinb(n6999), .dout(n7001));
  jand g06810(.dina(n7001), .dinb(n6998), .dout(n7002));
  jxor g06811(.dina(n7002), .dinb(n6995), .dout(n7003));
  jand g06812(.dina(\a[31] ), .dinb(\a[28] ), .dout(n7004));
  jxor g06813(.dina(n7004), .dinb(n3294), .dout(n7005));
  jxor g06814(.dina(n7005), .dinb(n6847), .dout(n7006));
  jxor g06815(.dina(n7006), .dinb(n7003), .dout(n7007));
  jnot g06816(.din(n7007), .dout(n7008));
  jand g06817(.dina(\a[51] ), .dinb(\a[8] ), .dout(n7009));
  jnot g06818(.din(n7009), .dout(n7010));
  jand g06819(.dina(n4317), .dinb(n937), .dout(n7011));
  jnot g06820(.din(n7011), .dout(n7012));
  jand g06821(.dina(\a[43] ), .dinb(\a[16] ), .dout(n7013));
  jand g06822(.dina(\a[42] ), .dinb(\a[17] ), .dout(n7014));
  jor  g06823(.dina(n7014), .dinb(n7013), .dout(n7015));
  jand g06824(.dina(n7015), .dinb(n7012), .dout(n7016));
  jxor g06825(.dina(n7016), .dinb(n7010), .dout(n7017));
  jxor g06826(.dina(n7017), .dinb(n7008), .dout(n7018));
  jxor g06827(.dina(n7018), .dinb(n6994), .dout(n7019));
  jxor g06828(.dina(n7019), .dinb(n6963), .dout(n7020));
  jxor g06829(.dina(n7020), .dinb(n6960), .dout(n7021));
  jand g06830(.dina(n6712), .dinb(n6710), .dout(n7022));
  jand g06831(.dina(n6716), .dinb(n6713), .dout(n7023));
  jor  g06832(.dina(n7023), .dinb(n7022), .dout(n7024));
  jand g06833(.dina(\a[53] ), .dinb(\a[6] ), .dout(n7025));
  jand g06834(.dina(\a[52] ), .dinb(\a[7] ), .dout(n7026));
  jand g06835(.dina(\a[41] ), .dinb(\a[18] ), .dout(n7027));
  jxor g06836(.dina(n7027), .dinb(n7026), .dout(n7028));
  jxor g06837(.dina(n7028), .dinb(n7025), .dout(n7029));
  jnot g06838(.din(n7029), .dout(n7030));
  jand g06839(.dina(\a[50] ), .dinb(\a[9] ), .dout(n7031));
  jnot g06840(.din(n7031), .dout(n7032));
  jand g06841(.dina(\a[49] ), .dinb(\a[44] ), .dout(n7033));
  jand g06842(.dina(n7033), .dinb(n1354), .dout(n7034));
  jnot g06843(.din(n7034), .dout(n7035));
  jand g06844(.dina(\a[44] ), .dinb(\a[15] ), .dout(n7036));
  jand g06845(.dina(\a[49] ), .dinb(\a[10] ), .dout(n7037));
  jor  g06846(.dina(n7037), .dinb(n7036), .dout(n7038));
  jand g06847(.dina(n7038), .dinb(n7035), .dout(n7039));
  jxor g06848(.dina(n7039), .dinb(n7032), .dout(n7040));
  jxor g06849(.dina(n7040), .dinb(n7030), .dout(n7041));
  jxor g06850(.dina(n7041), .dinb(n7024), .dout(n7042));
  jand g06851(.dina(n6680), .dinb(n6677), .dout(n7043));
  jand g06852(.dina(n6684), .dinb(n6681), .dout(n7044));
  jor  g06853(.dina(n7044), .dinb(n7043), .dout(n7045));
  jxor g06854(.dina(n7045), .dinb(n7042), .dout(n7046));
  jand g06855(.dina(\a[33] ), .dinb(\a[26] ), .dout(n7047));
  jand g06856(.dina(\a[59] ), .dinb(\a[32] ), .dout(n7048));
  jand g06857(.dina(n7048), .dinb(n1551), .dout(n7049));
  jnot g06858(.din(n7049), .dout(n7050));
  jand g06859(.dina(n2671), .dinb(n1927), .dout(n7051));
  jand g06860(.dina(\a[59] ), .dinb(\a[0] ), .dout(n7052));
  jand g06861(.dina(n7052), .dinb(n7047), .dout(n7053));
  jor  g06862(.dina(n7053), .dinb(n7051), .dout(n7054));
  jand g06863(.dina(n7054), .dinb(n7050), .dout(n7055));
  jnot g06864(.din(n7055), .dout(n7056));
  jand g06865(.dina(n7056), .dinb(n7047), .dout(n7057));
  jor  g06866(.dina(n7054), .dinb(n7049), .dout(n7058));
  jnot g06867(.din(n7058), .dout(n7059));
  jand g06868(.dina(\a[32] ), .dinb(\a[27] ), .dout(n7060));
  jor  g06869(.dina(n7060), .dinb(n7052), .dout(n7061));
  jand g06870(.dina(n7061), .dinb(n7059), .dout(n7062));
  jor  g06871(.dina(n7062), .dinb(n7057), .dout(n7063));
  jand g06872(.dina(\a[39] ), .dinb(\a[20] ), .dout(n7064));
  jand g06873(.dina(\a[38] ), .dinb(\a[22] ), .dout(n7065));
  jand g06874(.dina(n7065), .dinb(n6778), .dout(n7066));
  jnot g06875(.din(n7066), .dout(n7067));
  jand g06876(.dina(\a[37] ), .dinb(\a[22] ), .dout(n7068));
  jor  g06877(.dina(n7068), .dinb(n6775), .dout(n7069));
  jand g06878(.dina(n7069), .dinb(n7067), .dout(n7070));
  jxor g06879(.dina(n7070), .dinb(n7064), .dout(n7071));
  jand g06880(.dina(\a[36] ), .dinb(\a[23] ), .dout(n7072));
  jand g06881(.dina(n2845), .dinb(n1648), .dout(n7073));
  jnot g06882(.din(n7073), .dout(n7074));
  jand g06883(.dina(\a[35] ), .dinb(\a[24] ), .dout(n7075));
  jand g06884(.dina(\a[34] ), .dinb(\a[25] ), .dout(n7076));
  jor  g06885(.dina(n7076), .dinb(n7075), .dout(n7077));
  jand g06886(.dina(n7077), .dinb(n7074), .dout(n7078));
  jxor g06887(.dina(n7078), .dinb(n7072), .dout(n7079));
  jxor g06888(.dina(n7079), .dinb(n7071), .dout(n7080));
  jxor g06889(.dina(n7080), .dinb(n7063), .dout(n7081));
  jxor g06890(.dina(n7081), .dinb(n7046), .dout(n7082));
  jxor g06891(.dina(n7082), .dinb(n7021), .dout(n7083));
  jxor g06892(.dina(n7083), .dinb(n6957), .dout(n7084));
  jxor g06893(.dina(n7084), .dinb(n6906), .dout(n7085));
  jand g06894(.dina(n6695), .dinb(n6668), .dout(n7086));
  jand g06895(.dina(n6866), .dinb(n6696), .dout(n7087));
  jor  g06896(.dina(n7087), .dinb(n7086), .dout(n7088));
  jnot g06897(.din(n7088), .dout(n7089));
  jxor g06898(.dina(n7089), .dinb(n7085), .dout(n7090));
  jnot g06899(.din(n6868), .dout(n7091));
  jor  g06900(.dina(n6874), .dinb(n6870), .dout(n7092));
  jand g06901(.dina(n7092), .dinb(n7091), .dout(n7093));
  jxor g06902(.dina(n7093), .dinb(n7090), .dout(\asquared[60] ));
  jand g06903(.dina(n6905), .dinb(n6878), .dout(n7095));
  jand g06904(.dina(n7084), .dinb(n6906), .dout(n7096));
  jor  g06905(.dina(n7096), .dinb(n7095), .dout(n7097));
  jand g06906(.dina(n6956), .dinb(n6909), .dout(n7098));
  jand g06907(.dina(n7083), .dinb(n6957), .dout(n7099));
  jor  g06908(.dina(n7099), .dinb(n7098), .dout(n7100));
  jand g06909(.dina(n7020), .dinb(n6960), .dout(n7101));
  jand g06910(.dina(n7082), .dinb(n7021), .dout(n7102));
  jor  g06911(.dina(n7102), .dinb(n7101), .dout(n7103));
  jand g06912(.dina(n6954), .dinb(n6925), .dout(n7104));
  jand g06913(.dina(n6955), .dinb(n6922), .dout(n7105));
  jor  g06914(.dina(n7105), .dinb(n7104), .dout(n7106));
  jand g06915(.dina(n6939), .dinb(n6937), .dout(n7107));
  jand g06916(.dina(n6940), .dinb(n6935), .dout(n7108));
  jor  g06917(.dina(n7108), .dinb(n7107), .dout(n7109));
  jand g06918(.dina(n6931), .dinb(n6928), .dout(n7110));
  jand g06919(.dina(n6932), .dinb(n6766), .dout(n7111));
  jor  g06920(.dina(n7111), .dinb(n7110), .dout(n7112));
  jxor g06921(.dina(n7112), .dinb(n7109), .dout(n7113));
  jand g06922(.dina(n6992), .dinb(n6989), .dout(n7114));
  jand g06923(.dina(n6993), .dinb(n6980), .dout(n7115));
  jor  g06924(.dina(n7115), .dinb(n7114), .dout(n7116));
  jxor g06925(.dina(n7116), .dinb(n7113), .dout(n7117));
  jnot g06926(.din(n7117), .dout(n7118));
  jor  g06927(.dina(n6917), .dinb(n6913), .dout(n7119));
  jand g06928(.dina(n6921), .dinb(n6918), .dout(n7120));
  jnot g06929(.din(n7120), .dout(n7121));
  jand g06930(.dina(n7121), .dinb(n7119), .dout(n7122));
  jxor g06931(.dina(n7122), .dinb(n7118), .dout(n7123));
  jand g06932(.dina(n7045), .dinb(n7042), .dout(n7124));
  jand g06933(.dina(n7081), .dinb(n7046), .dout(n7125));
  jor  g06934(.dina(n7125), .dinb(n7124), .dout(n7126));
  jxor g06935(.dina(n7126), .dinb(n7123), .dout(n7127));
  jxor g06936(.dina(n7127), .dinb(n7106), .dout(n7128));
  jxor g06937(.dina(n7128), .dinb(n7103), .dout(n7129));
  jxor g06938(.dina(n7129), .dinb(n7100), .dout(n7130));
  jand g06939(.dina(n6952), .dinb(n6941), .dout(n7131));
  jand g06940(.dina(n6953), .dinb(n6933), .dout(n7132));
  jor  g06941(.dina(n7132), .dinb(n7131), .dout(n7133));
  jand g06942(.dina(n6950), .dinb(n6947), .dout(n7134));
  jand g06943(.dina(n6951), .dinb(n6942), .dout(n7135));
  jor  g06944(.dina(n7135), .dinb(n7134), .dout(n7136));
  jand g06945(.dina(\a[33] ), .dinb(\a[27] ), .dout(n7137));
  jand g06946(.dina(n2671), .dinb(n2042), .dout(n7138));
  jand g06947(.dina(\a[37] ), .dinb(\a[23] ), .dout(n7139));
  jand g06948(.dina(n7139), .dinb(n7137), .dout(n7140));
  jor  g06949(.dina(n7140), .dinb(n7138), .dout(n7141));
  jand g06950(.dina(\a[32] ), .dinb(\a[28] ), .dout(n7142));
  jand g06951(.dina(n7142), .dinb(n7139), .dout(n7143));
  jnot g06952(.din(n7143), .dout(n7144));
  jand g06953(.dina(n7144), .dinb(n7141), .dout(n7145));
  jnot g06954(.din(n7145), .dout(n7146));
  jand g06955(.dina(n7146), .dinb(n7137), .dout(n7147));
  jor  g06956(.dina(n7143), .dinb(n7141), .dout(n7148));
  jnot g06957(.din(n7148), .dout(n7149));
  jor  g06958(.dina(n7142), .dinb(n7139), .dout(n7150));
  jand g06959(.dina(n7150), .dinb(n7149), .dout(n7151));
  jor  g06960(.dina(n7151), .dinb(n7147), .dout(n7152));
  jand g06961(.dina(\a[60] ), .dinb(\a[0] ), .dout(n7153));
  jxor g06962(.dina(n7153), .dinb(n6943), .dout(n7154));
  jand g06963(.dina(\a[31] ), .dinb(\a[29] ), .dout(n7155));
  jand g06964(.dina(\a[59] ), .dinb(\a[1] ), .dout(n7156));
  jxor g06965(.dina(n7156), .dinb(n7155), .dout(n7157));
  jxor g06966(.dina(n7157), .dinb(n7154), .dout(n7158));
  jxor g06967(.dina(n7158), .dinb(n7152), .dout(n7159));
  jxor g06968(.dina(n7159), .dinb(n7136), .dout(n7160));
  jand g06969(.dina(\a[52] ), .dinb(\a[8] ), .dout(n7161));
  jand g06970(.dina(\a[42] ), .dinb(\a[18] ), .dout(n7162));
  jand g06971(.dina(n7162), .dinb(n7161), .dout(n7163));
  jnot g06972(.din(n7163), .dout(n7164));
  jand g06973(.dina(\a[53] ), .dinb(\a[52] ), .dout(n7165));
  jand g06974(.dina(n7165), .dinb(n499), .dout(n7166));
  jand g06975(.dina(\a[53] ), .dinb(\a[7] ), .dout(n7167));
  jand g06976(.dina(n7167), .dinb(n7162), .dout(n7168));
  jor  g06977(.dina(n7168), .dinb(n7166), .dout(n7169));
  jnot g06978(.din(n7169), .dout(n7170));
  jand g06979(.dina(n7170), .dinb(n7164), .dout(n7171));
  jor  g06980(.dina(n7162), .dinb(n7161), .dout(n7172));
  jand g06981(.dina(n7172), .dinb(n7171), .dout(n7173));
  jand g06982(.dina(n7169), .dinb(n7164), .dout(n7174));
  jnot g06983(.din(n7174), .dout(n7175));
  jand g06984(.dina(n7175), .dinb(n7167), .dout(n7176));
  jor  g06985(.dina(n7176), .dinb(n7173), .dout(n7177));
  jand g06986(.dina(\a[46] ), .dinb(\a[14] ), .dout(n7178));
  jnot g06987(.din(n7178), .dout(n7179));
  jand g06988(.dina(n5316), .dinb(n899), .dout(n7180));
  jnot g06989(.din(n7180), .dout(n7181));
  jand g06990(.dina(\a[48] ), .dinb(\a[12] ), .dout(n7182));
  jand g06991(.dina(\a[47] ), .dinb(\a[13] ), .dout(n7183));
  jor  g06992(.dina(n7183), .dinb(n7182), .dout(n7184));
  jand g06993(.dina(n7184), .dinb(n7181), .dout(n7185));
  jxor g06994(.dina(n7185), .dinb(n7179), .dout(n7186));
  jnot g06995(.din(n7186), .dout(n7187));
  jxor g06996(.dina(n7187), .dinb(n7177), .dout(n7188));
  jand g06997(.dina(\a[54] ), .dinb(\a[6] ), .dout(n7189));
  jand g06998(.dina(\a[41] ), .dinb(\a[19] ), .dout(n7190));
  jxor g06999(.dina(n7190), .dinb(n7189), .dout(n7191));
  jxor g07000(.dina(n7191), .dinb(n6965), .dout(n7192));
  jxor g07001(.dina(n7192), .dinb(n7188), .dout(n7193));
  jxor g07002(.dina(n7193), .dinb(n7160), .dout(n7194));
  jxor g07003(.dina(n7194), .dinb(n7133), .dout(n7195));
  jand g07004(.dina(n6901), .dinb(n6898), .dout(n7196));
  jand g07005(.dina(n6902), .dinb(n6887), .dout(n7197));
  jor  g07006(.dina(n7197), .dinb(n7196), .dout(n7198));
  jand g07007(.dina(n6893), .dinb(n6890), .dout(n7199));
  jand g07008(.dina(n6897), .dinb(n6894), .dout(n7200));
  jor  g07009(.dina(n7200), .dinb(n7199), .dout(n7201));
  jand g07010(.dina(\a[58] ), .dinb(\a[2] ), .dout(n7202));
  jand g07011(.dina(\a[57] ), .dinb(\a[4] ), .dout(n7203));
  jand g07012(.dina(n7203), .dinb(n6983), .dout(n7204));
  jnot g07013(.din(n7204), .dout(n7205));
  jand g07014(.dina(\a[56] ), .dinb(\a[4] ), .dout(n7206));
  jor  g07015(.dina(n7206), .dinb(n6985), .dout(n7207));
  jand g07016(.dina(n7207), .dinb(n7205), .dout(n7208));
  jxor g07017(.dina(n7208), .dinb(n7202), .dout(n7209));
  jnot g07018(.din(n7209), .dout(n7210));
  jand g07019(.dina(\a[40] ), .dinb(\a[20] ), .dout(n7211));
  jnot g07020(.din(n7211), .dout(n7212));
  jand g07021(.dina(\a[39] ), .dinb(\a[22] ), .dout(n7213));
  jand g07022(.dina(n7213), .dinb(n6775), .dout(n7214));
  jnot g07023(.din(n7214), .dout(n7215));
  jand g07024(.dina(\a[39] ), .dinb(\a[21] ), .dout(n7216));
  jor  g07025(.dina(n7216), .dinb(n7065), .dout(n7217));
  jand g07026(.dina(n7217), .dinb(n7215), .dout(n7218));
  jxor g07027(.dina(n7218), .dinb(n7212), .dout(n7219));
  jxor g07028(.dina(n7219), .dinb(n7210), .dout(n7220));
  jnot g07029(.din(n7220), .dout(n7221));
  jand g07030(.dina(\a[36] ), .dinb(\a[24] ), .dout(n7222));
  jnot g07031(.din(n7222), .dout(n7223));
  jand g07032(.dina(n2845), .dinb(n2128), .dout(n7224));
  jnot g07033(.din(n7224), .dout(n7225));
  jand g07034(.dina(\a[34] ), .dinb(\a[26] ), .dout(n7226));
  jand g07035(.dina(\a[35] ), .dinb(\a[25] ), .dout(n7227));
  jor  g07036(.dina(n7227), .dinb(n7226), .dout(n7228));
  jand g07037(.dina(n7228), .dinb(n7225), .dout(n7229));
  jxor g07038(.dina(n7229), .dinb(n7223), .dout(n7230));
  jxor g07039(.dina(n7230), .dinb(n7221), .dout(n7231));
  jxor g07040(.dina(n7231), .dinb(n7201), .dout(n7232));
  jand g07041(.dina(n7002), .dinb(n6995), .dout(n7233));
  jor  g07042(.dina(n7233), .dinb(n6997), .dout(n7234));
  jand g07043(.dina(\a[43] ), .dinb(\a[17] ), .dout(n7235));
  jand g07044(.dina(\a[51] ), .dinb(\a[44] ), .dout(n7236));
  jand g07045(.dina(n7236), .dinb(n1367), .dout(n7237));
  jnot g07046(.din(n7237), .dout(n7238));
  jand g07047(.dina(n4495), .dinb(n937), .dout(n7239));
  jand g07048(.dina(\a[51] ), .dinb(\a[9] ), .dout(n7240));
  jand g07049(.dina(n7240), .dinb(n7235), .dout(n7241));
  jor  g07050(.dina(n7241), .dinb(n7239), .dout(n7242));
  jand g07051(.dina(n7242), .dinb(n7238), .dout(n7243));
  jnot g07052(.din(n7243), .dout(n7244));
  jand g07053(.dina(n7244), .dinb(n7235), .dout(n7245));
  jor  g07054(.dina(n7242), .dinb(n7237), .dout(n7246));
  jnot g07055(.din(n7246), .dout(n7247));
  jand g07056(.dina(\a[44] ), .dinb(\a[16] ), .dout(n7248));
  jor  g07057(.dina(n7248), .dinb(n7240), .dout(n7249));
  jand g07058(.dina(n7249), .dinb(n7247), .dout(n7250));
  jor  g07059(.dina(n7250), .dinb(n7245), .dout(n7251));
  jxor g07060(.dina(n7251), .dinb(n7234), .dout(n7252));
  jnot g07061(.din(n7252), .dout(n7253));
  jand g07062(.dina(\a[50] ), .dinb(\a[10] ), .dout(n7254));
  jand g07063(.dina(\a[49] ), .dinb(\a[45] ), .dout(n7255));
  jand g07064(.dina(n7255), .dinb(n1469), .dout(n7256));
  jand g07065(.dina(\a[49] ), .dinb(\a[11] ), .dout(n7257));
  jnot g07066(.din(n7257), .dout(n7258));
  jand g07067(.dina(\a[45] ), .dinb(\a[15] ), .dout(n7259));
  jnot g07068(.din(n7259), .dout(n7260));
  jand g07069(.dina(n7260), .dinb(n7258), .dout(n7261));
  jor  g07070(.dina(n7261), .dinb(n7256), .dout(n7262));
  jxor g07071(.dina(n7262), .dinb(n7254), .dout(n7263));
  jxor g07072(.dina(n7263), .dinb(n7253), .dout(n7264));
  jxor g07073(.dina(n7264), .dinb(n7232), .dout(n7265));
  jxor g07074(.dina(n7265), .dinb(n7198), .dout(n7266));
  jxor g07075(.dina(n7266), .dinb(n7195), .dout(n7267));
  jand g07076(.dina(n6903), .dinb(n6884), .dout(n7268));
  jand g07077(.dina(n6904), .dinb(n6881), .dout(n7269));
  jor  g07078(.dina(n7269), .dinb(n7268), .dout(n7270));
  jand g07079(.dina(n7004), .dinb(n3294), .dout(n7271));
  jand g07080(.dina(n7005), .dinb(n6847), .dout(n7272));
  jor  g07081(.dina(n7272), .dinb(n7271), .dout(n7273));
  jand g07082(.dina(n7027), .dinb(n7026), .dout(n7274));
  jand g07083(.dina(n7028), .dinb(n7025), .dout(n7275));
  jor  g07084(.dina(n7275), .dinb(n7274), .dout(n7276));
  jand g07085(.dina(n7012), .dinb(n7010), .dout(n7277));
  jnot g07086(.din(n7277), .dout(n7278));
  jand g07087(.dina(n7278), .dinb(n7015), .dout(n7279));
  jxor g07088(.dina(n7279), .dinb(n7276), .dout(n7280));
  jxor g07089(.dina(n7280), .dinb(n7273), .dout(n7281));
  jand g07090(.dina(n7079), .dinb(n7071), .dout(n7282));
  jand g07091(.dina(n7080), .dinb(n7063), .dout(n7283));
  jor  g07092(.dina(n7283), .dinb(n7282), .dout(n7284));
  jxor g07093(.dina(n7284), .dinb(n7281), .dout(n7285));
  jnot g07094(.din(n7285), .dout(n7286));
  jand g07095(.dina(n7006), .dinb(n7003), .dout(n7287));
  jnot g07096(.din(n7287), .dout(n7288));
  jor  g07097(.dina(n7017), .dinb(n7008), .dout(n7289));
  jand g07098(.dina(n7289), .dinb(n7288), .dout(n7290));
  jxor g07099(.dina(n7290), .dinb(n7286), .dout(n7291));
  jand g07100(.dina(n7018), .dinb(n6994), .dout(n7292));
  jand g07101(.dina(n7019), .dinb(n6963), .dout(n7293));
  jor  g07102(.dina(n7293), .dinb(n7292), .dout(n7294));
  jor  g07103(.dina(n7040), .dinb(n7030), .dout(n7295));
  jand g07104(.dina(n7041), .dinb(n7024), .dout(n7296));
  jnot g07105(.din(n7296), .dout(n7297));
  jand g07106(.dina(n7297), .dinb(n7295), .dout(n7298));
  jnot g07107(.din(n7298), .dout(n7299));
  jand g07108(.dina(n7070), .dinb(n7064), .dout(n7300));
  jor  g07109(.dina(n7300), .dinb(n7066), .dout(n7301));
  jxor g07110(.dina(n7301), .dinb(n6976), .dout(n7302));
  jor  g07111(.dina(n7073), .dinb(n7072), .dout(n7303));
  jand g07112(.dina(n7303), .dinb(n7077), .dout(n7304));
  jxor g07113(.dina(n7304), .dinb(n7302), .dout(n7305));
  jand g07114(.dina(n6988), .dinb(n6981), .dout(n7306));
  jor  g07115(.dina(n7306), .dinb(n6986), .dout(n7307));
  jxor g07116(.dina(n7307), .dinb(n7058), .dout(n7308));
  jand g07117(.dina(n7035), .dinb(n7032), .dout(n7309));
  jnot g07118(.din(n7309), .dout(n7310));
  jand g07119(.dina(n7310), .dinb(n7038), .dout(n7311));
  jxor g07120(.dina(n7311), .dinb(n7308), .dout(n7312));
  jxor g07121(.dina(n7312), .dinb(n7305), .dout(n7313));
  jxor g07122(.dina(n7313), .dinb(n7299), .dout(n7314));
  jxor g07123(.dina(n7314), .dinb(n7294), .dout(n7315));
  jxor g07124(.dina(n7315), .dinb(n7291), .dout(n7316));
  jxor g07125(.dina(n7316), .dinb(n7270), .dout(n7317));
  jxor g07126(.dina(n7317), .dinb(n7267), .dout(n7318));
  jxor g07127(.dina(n7318), .dinb(n7130), .dout(n7319));
  jnot g07128(.din(n7319), .dout(n7320));
  jxor g07129(.dina(n7320), .dinb(n7097), .dout(n7321));
  jand g07130(.dina(n7088), .dinb(n7085), .dout(n7322));
  jnot g07131(.din(n7322), .dout(n7323));
  jnot g07132(.din(n7085), .dout(n7324));
  jand g07133(.dina(n7089), .dinb(n7324), .dout(n7325));
  jor  g07134(.dina(n7093), .dinb(n7325), .dout(n7326));
  jand g07135(.dina(n7326), .dinb(n7323), .dout(n7327));
  jxor g07136(.dina(n7327), .dinb(n7321), .dout(\asquared[61] ));
  jand g07137(.dina(n7129), .dinb(n7100), .dout(n7329));
  jand g07138(.dina(n7318), .dinb(n7130), .dout(n7330));
  jor  g07139(.dina(n7330), .dinb(n7329), .dout(n7331));
  jand g07140(.dina(n7127), .dinb(n7106), .dout(n7332));
  jand g07141(.dina(n7128), .dinb(n7103), .dout(n7333));
  jor  g07142(.dina(n7333), .dinb(n7332), .dout(n7334));
  jnot g07143(.din(n7334), .dout(n7335));
  jand g07144(.dina(n7193), .dinb(n7160), .dout(n7336));
  jand g07145(.dina(n7194), .dinb(n7133), .dout(n7337));
  jor  g07146(.dina(n7337), .dinb(n7336), .dout(n7338));
  jxor g07147(.dina(n7247), .dinb(n7171), .dout(n7339));
  jand g07148(.dina(n7153), .dinb(n6943), .dout(n7340));
  jand g07149(.dina(n7157), .dinb(n7154), .dout(n7341));
  jor  g07150(.dina(n7341), .dinb(n7340), .dout(n7342));
  jxor g07151(.dina(n7342), .dinb(n7339), .dout(n7343));
  jand g07152(.dina(n7187), .dinb(n7177), .dout(n7344));
  jand g07153(.dina(n7192), .dinb(n7188), .dout(n7345));
  jor  g07154(.dina(n7345), .dinb(n7344), .dout(n7346));
  jxor g07155(.dina(n7346), .dinb(n7343), .dout(n7347));
  jand g07156(.dina(n7158), .dinb(n7152), .dout(n7348));
  jand g07157(.dina(n7159), .dinb(n7136), .dout(n7349));
  jor  g07158(.dina(n7349), .dinb(n7348), .dout(n7350));
  jxor g07159(.dina(n7350), .dinb(n7347), .dout(n7351));
  jor  g07160(.dina(n7219), .dinb(n7210), .dout(n7352));
  jor  g07161(.dina(n7230), .dinb(n7221), .dout(n7353));
  jand g07162(.dina(n7353), .dinb(n7352), .dout(n7354));
  jnot g07163(.din(n7354), .dout(n7355));
  jand g07164(.dina(n7225), .dinb(n7223), .dout(n7356));
  jnot g07165(.din(n7356), .dout(n7357));
  jand g07166(.dina(n7357), .dinb(n7228), .dout(n7358));
  jxor g07167(.dina(n7358), .dinb(n7148), .dout(n7359));
  jand g07168(.dina(n7215), .dinb(n7212), .dout(n7360));
  jnot g07169(.din(n7360), .dout(n7361));
  jand g07170(.dina(n7361), .dinb(n7217), .dout(n7362));
  jxor g07171(.dina(n7362), .dinb(n7359), .dout(n7363));
  jand g07172(.dina(n7190), .dinb(n7189), .dout(n7364));
  jand g07173(.dina(n7191), .dinb(n6965), .dout(n7365));
  jor  g07174(.dina(n7365), .dinb(n7364), .dout(n7366));
  jand g07175(.dina(n7208), .dinb(n7202), .dout(n7367));
  jor  g07176(.dina(n7367), .dinb(n7204), .dout(n7368));
  jxor g07177(.dina(n7368), .dinb(n7366), .dout(n7369));
  jnot g07178(.din(n7254), .dout(n7370));
  jnot g07179(.din(n7256), .dout(n7371));
  jand g07180(.dina(n7371), .dinb(n7370), .dout(n7372));
  jor  g07181(.dina(n7372), .dinb(n7261), .dout(n7373));
  jnot g07182(.din(n7373), .dout(n7374));
  jxor g07183(.dina(n7374), .dinb(n7369), .dout(n7375));
  jxor g07184(.dina(n7375), .dinb(n7363), .dout(n7376));
  jxor g07185(.dina(n7376), .dinb(n7355), .dout(n7377));
  jnot g07186(.din(n7377), .dout(n7378));
  jxor g07187(.dina(n7378), .dinb(n7351), .dout(n7379));
  jxor g07188(.dina(n7379), .dinb(n7338), .dout(n7380));
  jxor g07189(.dina(n7380), .dinb(n7335), .dout(n7381));
  jand g07190(.dina(n7314), .dinb(n7294), .dout(n7382));
  jand g07191(.dina(n7315), .dinb(n7291), .dout(n7383));
  jor  g07192(.dina(n7383), .dinb(n7382), .dout(n7384));
  jor  g07193(.dina(n7122), .dinb(n7118), .dout(n7385));
  jand g07194(.dina(n7126), .dinb(n7123), .dout(n7386));
  jnot g07195(.din(n7386), .dout(n7387));
  jand g07196(.dina(n7387), .dinb(n7385), .dout(n7388));
  jnot g07197(.din(n7388), .dout(n7389));
  jand g07198(.dina(n7112), .dinb(n7109), .dout(n7390));
  jand g07199(.dina(n7116), .dinb(n7113), .dout(n7391));
  jor  g07200(.dina(n7391), .dinb(n7390), .dout(n7392));
  jand g07201(.dina(\a[51] ), .dinb(\a[46] ), .dout(n7393));
  jand g07202(.dina(n7393), .dinb(n1354), .dout(n7394));
  jnot g07203(.din(n7394), .dout(n7395));
  jand g07204(.dina(\a[46] ), .dinb(\a[16] ), .dout(n7396));
  jand g07205(.dina(n7396), .dinb(n7259), .dout(n7397));
  jand g07206(.dina(\a[51] ), .dinb(\a[10] ), .dout(n7398));
  jand g07207(.dina(\a[45] ), .dinb(\a[16] ), .dout(n7399));
  jand g07208(.dina(n7399), .dinb(n7398), .dout(n7400));
  jor  g07209(.dina(n7400), .dinb(n7397), .dout(n7401));
  jnot g07210(.din(n7401), .dout(n7402));
  jand g07211(.dina(n7402), .dinb(n7395), .dout(n7403));
  jand g07212(.dina(\a[46] ), .dinb(\a[15] ), .dout(n7404));
  jor  g07213(.dina(n7404), .dinb(n7398), .dout(n7405));
  jand g07214(.dina(n7405), .dinb(n7403), .dout(n7406));
  jand g07215(.dina(n7401), .dinb(n7395), .dout(n7407));
  jnot g07216(.din(n7407), .dout(n7408));
  jand g07217(.dina(n7408), .dinb(n7399), .dout(n7409));
  jor  g07218(.dina(n7409), .dinb(n7406), .dout(n7410));
  jand g07219(.dina(\a[50] ), .dinb(\a[11] ), .dout(n7411));
  jand g07220(.dina(\a[49] ), .dinb(\a[47] ), .dout(n7412));
  jand g07221(.dina(n7412), .dinb(n979), .dout(n7413));
  jnot g07222(.din(n7413), .dout(n7414));
  jand g07223(.dina(\a[47] ), .dinb(\a[14] ), .dout(n7415));
  jand g07224(.dina(n7415), .dinb(n7411), .dout(n7416));
  jand g07225(.dina(\a[50] ), .dinb(\a[12] ), .dout(n7417));
  jand g07226(.dina(n7417), .dinb(n7257), .dout(n7418));
  jor  g07227(.dina(n7418), .dinb(n7416), .dout(n7419));
  jand g07228(.dina(n7419), .dinb(n7414), .dout(n7420));
  jnot g07229(.din(n7420), .dout(n7421));
  jand g07230(.dina(n7421), .dinb(n7411), .dout(n7422));
  jor  g07231(.dina(n7419), .dinb(n7413), .dout(n7423));
  jnot g07232(.din(n7423), .dout(n7424));
  jand g07233(.dina(\a[49] ), .dinb(\a[12] ), .dout(n7425));
  jor  g07234(.dina(n7425), .dinb(n7415), .dout(n7426));
  jand g07235(.dina(n7426), .dinb(n7424), .dout(n7427));
  jor  g07236(.dina(n7427), .dinb(n7422), .dout(n7428));
  jxor g07237(.dina(n7428), .dinb(n7410), .dout(n7429));
  jand g07238(.dina(\a[48] ), .dinb(\a[13] ), .dout(n7430));
  jnot g07239(.din(n7430), .dout(n7431));
  jand g07240(.dina(n3294), .dinb(n3269), .dout(n7432));
  jnot g07241(.din(n7432), .dout(n7433));
  jand g07242(.dina(\a[32] ), .dinb(\a[29] ), .dout(n7434));
  jor  g07243(.dina(n7434), .dinb(n2440), .dout(n7435));
  jand g07244(.dina(n7435), .dinb(n7433), .dout(n7436));
  jxor g07245(.dina(n7436), .dinb(n7431), .dout(n7437));
  jnot g07246(.din(n7437), .dout(n7438));
  jxor g07247(.dina(n7438), .dinb(n7429), .dout(n7439));
  jxor g07248(.dina(n7439), .dinb(n7392), .dout(n7440));
  jand g07249(.dina(\a[59] ), .dinb(\a[2] ), .dout(n7441));
  jand g07250(.dina(\a[56] ), .dinb(\a[5] ), .dout(n7442));
  jand g07251(.dina(n7442), .dinb(n7441), .dout(n7443));
  jnot g07252(.din(n7443), .dout(n7444));
  jand g07253(.dina(\a[61] ), .dinb(\a[2] ), .dout(n7445));
  jand g07254(.dina(n7445), .dinb(n7052), .dout(n7446));
  jand g07255(.dina(\a[61] ), .dinb(\a[0] ), .dout(n7447));
  jand g07256(.dina(n7447), .dinb(n7442), .dout(n7448));
  jor  g07257(.dina(n7448), .dinb(n7446), .dout(n7449));
  jnot g07258(.din(n7449), .dout(n7450));
  jand g07259(.dina(n7450), .dinb(n7444), .dout(n7451));
  jor  g07260(.dina(n7442), .dinb(n7441), .dout(n7452));
  jand g07261(.dina(n7452), .dinb(n7451), .dout(n7453));
  jand g07262(.dina(n7449), .dinb(n7444), .dout(n7454));
  jnot g07263(.din(n7454), .dout(n7455));
  jand g07264(.dina(n7455), .dinb(n7447), .dout(n7456));
  jor  g07265(.dina(n7456), .dinb(n7453), .dout(n7457));
  jand g07266(.dina(\a[55] ), .dinb(\a[6] ), .dout(n7458));
  jnot g07267(.din(n7458), .dout(n7459));
  jand g07268(.dina(n4632), .dinb(n1490), .dout(n7460));
  jnot g07269(.din(n7460), .dout(n7461));
  jand g07270(.dina(\a[41] ), .dinb(\a[20] ), .dout(n7462));
  jand g07271(.dina(\a[40] ), .dinb(\a[21] ), .dout(n7463));
  jor  g07272(.dina(n7463), .dinb(n7462), .dout(n7464));
  jand g07273(.dina(n7464), .dinb(n7461), .dout(n7465));
  jxor g07274(.dina(n7465), .dinb(n7459), .dout(n7466));
  jnot g07275(.din(n7466), .dout(n7467));
  jxor g07276(.dina(n7467), .dinb(n7457), .dout(n7468));
  jnot g07277(.din(n7468), .dout(n7469));
  jnot g07278(.din(n7213), .dout(n7470));
  jand g07279(.dina(n3138), .dinb(n1648), .dout(n7471));
  jnot g07280(.din(n7471), .dout(n7472));
  jand g07281(.dina(\a[37] ), .dinb(\a[24] ), .dout(n7473));
  jand g07282(.dina(\a[36] ), .dinb(\a[25] ), .dout(n7474));
  jor  g07283(.dina(n7474), .dinb(n7473), .dout(n7475));
  jand g07284(.dina(n7475), .dinb(n7472), .dout(n7476));
  jxor g07285(.dina(n7476), .dinb(n7470), .dout(n7477));
  jxor g07286(.dina(n7477), .dinb(n7469), .dout(n7478));
  jxor g07287(.dina(n7478), .dinb(n7440), .dout(n7479));
  jxor g07288(.dina(n7479), .dinb(n7389), .dout(n7480));
  jxor g07289(.dina(n7480), .dinb(n7384), .dout(n7481));
  jxor g07290(.dina(n7481), .dinb(n7381), .dout(n7482));
  jand g07291(.dina(n7316), .dinb(n7270), .dout(n7483));
  jand g07292(.dina(n7317), .dinb(n7267), .dout(n7484));
  jor  g07293(.dina(n7484), .dinb(n7483), .dout(n7485));
  jand g07294(.dina(n7265), .dinb(n7198), .dout(n7486));
  jand g07295(.dina(n7266), .dinb(n7195), .dout(n7487));
  jor  g07296(.dina(n7487), .dinb(n7486), .dout(n7488));
  jand g07297(.dina(n7231), .dinb(n7201), .dout(n7489));
  jand g07298(.dina(n7264), .dinb(n7232), .dout(n7490));
  jor  g07299(.dina(n7490), .dinb(n7489), .dout(n7491));
  jand g07300(.dina(n7251), .dinb(n7234), .dout(n7492));
  jnot g07301(.din(n7492), .dout(n7493));
  jor  g07302(.dina(n7263), .dinb(n7253), .dout(n7494));
  jand g07303(.dina(n7494), .dinb(n7493), .dout(n7495));
  jnot g07304(.din(n7495), .dout(n7496));
  jand g07305(.dina(n7301), .dinb(n6976), .dout(n7497));
  jand g07306(.dina(n7304), .dinb(n7302), .dout(n7498));
  jor  g07307(.dina(n7498), .dinb(n7497), .dout(n7499));
  jand g07308(.dina(\a[60] ), .dinb(\a[1] ), .dout(n7500));
  jnot g07309(.din(n7500), .dout(n7501));
  jnot g07310(.din(\a[31] ), .dout(n7502));
  jand g07311(.dina(n7156), .dinb(n7155), .dout(n7503));
  jor  g07312(.dina(n7503), .dinb(n7502), .dout(n7504));
  jxor g07313(.dina(n7504), .dinb(n7501), .dout(n7505));
  jand g07314(.dina(n7181), .dinb(n7179), .dout(n7506));
  jnot g07315(.din(n7506), .dout(n7507));
  jand g07316(.dina(n7507), .dinb(n7184), .dout(n7508));
  jxor g07317(.dina(n7508), .dinb(n7505), .dout(n7509));
  jxor g07318(.dina(n7509), .dinb(n7499), .dout(n7510));
  jxor g07319(.dina(n7510), .dinb(n7496), .dout(n7511));
  jand g07320(.dina(n7307), .dinb(n7058), .dout(n7512));
  jand g07321(.dina(n7311), .dinb(n7308), .dout(n7513));
  jor  g07322(.dina(n7513), .dinb(n7512), .dout(n7514));
  jand g07323(.dina(n7279), .dinb(n7276), .dout(n7515));
  jand g07324(.dina(n7280), .dinb(n7273), .dout(n7516));
  jor  g07325(.dina(n7516), .dinb(n7515), .dout(n7517));
  jand g07326(.dina(\a[38] ), .dinb(\a[23] ), .dout(n7518));
  jand g07327(.dina(\a[58] ), .dinb(\a[57] ), .dout(n7519));
  jand g07328(.dina(n7519), .dinb(n265), .dout(n7520));
  jnot g07329(.din(n7520), .dout(n7521));
  jand g07330(.dina(\a[58] ), .dinb(\a[3] ), .dout(n7522));
  jor  g07331(.dina(n7522), .dinb(n7203), .dout(n7523));
  jand g07332(.dina(n7523), .dinb(n7521), .dout(n7524));
  jxor g07333(.dina(n7524), .dinb(n7518), .dout(n7525));
  jxor g07334(.dina(n7525), .dinb(n7517), .dout(n7526));
  jxor g07335(.dina(n7526), .dinb(n7514), .dout(n7527));
  jxor g07336(.dina(n7527), .dinb(n7511), .dout(n7528));
  jxor g07337(.dina(n7528), .dinb(n7491), .dout(n7529));
  jand g07338(.dina(n7284), .dinb(n7281), .dout(n7530));
  jnot g07339(.din(n7530), .dout(n7531));
  jor  g07340(.dina(n7290), .dinb(n7286), .dout(n7532));
  jand g07341(.dina(n7532), .dinb(n7531), .dout(n7533));
  jnot g07342(.din(n7533), .dout(n7534));
  jand g07343(.dina(n7312), .dinb(n7305), .dout(n7535));
  jand g07344(.dina(n7313), .dinb(n7299), .dout(n7536));
  jor  g07345(.dina(n7536), .dinb(n7535), .dout(n7537));
  jand g07346(.dina(\a[43] ), .dinb(\a[18] ), .dout(n7538));
  jand g07347(.dina(\a[52] ), .dinb(\a[44] ), .dout(n7539));
  jand g07348(.dina(n7539), .dinb(n1465), .dout(n7540));
  jnot g07349(.din(n7540), .dout(n7541));
  jand g07350(.dina(\a[52] ), .dinb(\a[9] ), .dout(n7542));
  jand g07351(.dina(n7542), .dinb(n7538), .dout(n7543));
  jand g07352(.dina(n4495), .dinb(n1107), .dout(n7544));
  jor  g07353(.dina(n7544), .dinb(n7543), .dout(n7545));
  jand g07354(.dina(n7545), .dinb(n7541), .dout(n7546));
  jnot g07355(.din(n7546), .dout(n7547));
  jand g07356(.dina(n7547), .dinb(n7538), .dout(n7548));
  jor  g07357(.dina(n7545), .dinb(n7540), .dout(n7549));
  jnot g07358(.din(n7549), .dout(n7550));
  jand g07359(.dina(\a[44] ), .dinb(\a[17] ), .dout(n7551));
  jor  g07360(.dina(n7551), .dinb(n7542), .dout(n7552));
  jand g07361(.dina(n7552), .dinb(n7550), .dout(n7553));
  jor  g07362(.dina(n7553), .dinb(n7548), .dout(n7554));
  jand g07363(.dina(\a[42] ), .dinb(\a[19] ), .dout(n7555));
  jand g07364(.dina(\a[54] ), .dinb(\a[7] ), .dout(n7556));
  jand g07365(.dina(\a[53] ), .dinb(\a[8] ), .dout(n7557));
  jor  g07366(.dina(n7557), .dinb(n7556), .dout(n7558));
  jand g07367(.dina(\a[54] ), .dinb(\a[53] ), .dout(n7559));
  jand g07368(.dina(n7559), .dinb(n499), .dout(n7560));
  jnot g07369(.din(n7560), .dout(n7561));
  jand g07370(.dina(n7561), .dinb(n7558), .dout(n7562));
  jxor g07371(.dina(n7562), .dinb(n7555), .dout(n7563));
  jxor g07372(.dina(n7563), .dinb(n7554), .dout(n7564));
  jnot g07373(.din(n7564), .dout(n7565));
  jand g07374(.dina(\a[35] ), .dinb(\a[26] ), .dout(n7566));
  jnot g07375(.din(n7566), .dout(n7567));
  jand g07376(.dina(n3634), .dinb(n2042), .dout(n7568));
  jnot g07377(.din(n7568), .dout(n7569));
  jand g07378(.dina(\a[33] ), .dinb(\a[28] ), .dout(n7570));
  jor  g07379(.dina(n7570), .dinb(n3009), .dout(n7571));
  jand g07380(.dina(n7571), .dinb(n7569), .dout(n7572));
  jxor g07381(.dina(n7572), .dinb(n7567), .dout(n7573));
  jxor g07382(.dina(n7573), .dinb(n7565), .dout(n7574));
  jxor g07383(.dina(n7574), .dinb(n7537), .dout(n7575));
  jxor g07384(.dina(n7575), .dinb(n7534), .dout(n7576));
  jxor g07385(.dina(n7576), .dinb(n7529), .dout(n7577));
  jxor g07386(.dina(n7577), .dinb(n7488), .dout(n7578));
  jxor g07387(.dina(n7578), .dinb(n7485), .dout(n7579));
  jxor g07388(.dina(n7579), .dinb(n7482), .dout(n7580));
  jand g07389(.dina(n7580), .dinb(n7331), .dout(n7581));
  jor  g07390(.dina(n7580), .dinb(n7331), .dout(n7582));
  jnot g07391(.din(n7582), .dout(n7583));
  jor  g07392(.dina(n7583), .dinb(n7581), .dout(n7584));
  jand g07393(.dina(n7319), .dinb(n7097), .dout(n7585));
  jnot g07394(.din(n7585), .dout(n7586));
  jnot g07395(.din(n7097), .dout(n7587));
  jand g07396(.dina(n7320), .dinb(n7587), .dout(n7588));
  jor  g07397(.dina(n7327), .dinb(n7588), .dout(n7589));
  jand g07398(.dina(n7589), .dinb(n7586), .dout(n7590));
  jxor g07399(.dina(n7590), .dinb(n7584), .dout(\asquared[62] ));
  jand g07400(.dina(n7578), .dinb(n7485), .dout(n7592));
  jand g07401(.dina(n7579), .dinb(n7482), .dout(n7593));
  jor  g07402(.dina(n7593), .dinb(n7592), .dout(n7594));
  jand g07403(.dina(n7576), .dinb(n7529), .dout(n7595));
  jand g07404(.dina(n7577), .dinb(n7488), .dout(n7596));
  jor  g07405(.dina(n7596), .dinb(n7595), .dout(n7597));
  jand g07406(.dina(n7563), .dinb(n7554), .dout(n7598));
  jnot g07407(.din(n7598), .dout(n7599));
  jor  g07408(.dina(n7573), .dinb(n7565), .dout(n7600));
  jand g07409(.dina(n7600), .dinb(n7599), .dout(n7601));
  jnot g07410(.din(n7601), .dout(n7602));
  jxor g07411(.dina(n7550), .dinb(n7403), .dout(n7603));
  jand g07412(.dina(\a[59] ), .dinb(\a[3] ), .dout(n7604));
  jand g07413(.dina(n7519), .dinb(n242), .dout(n7605));
  jnot g07414(.din(n7605), .dout(n7606));
  jand g07415(.dina(\a[58] ), .dinb(\a[4] ), .dout(n7607));
  jand g07416(.dina(\a[57] ), .dinb(\a[5] ), .dout(n7608));
  jor  g07417(.dina(n7608), .dinb(n7607), .dout(n7609));
  jand g07418(.dina(n7609), .dinb(n7606), .dout(n7610));
  jxor g07419(.dina(n7610), .dinb(n7604), .dout(n7611));
  jxor g07420(.dina(n7611), .dinb(n7603), .dout(n7612));
  jxor g07421(.dina(n7612), .dinb(n7602), .dout(n7613));
  jand g07422(.dina(n7525), .dinb(n7517), .dout(n7614));
  jand g07423(.dina(n7526), .dinb(n7514), .dout(n7615));
  jor  g07424(.dina(n7615), .dinb(n7614), .dout(n7616));
  jxor g07425(.dina(n7616), .dinb(n7613), .dout(n7617));
  jnot g07426(.din(n7171), .dout(n7618));
  jand g07427(.dina(n7246), .dinb(n7618), .dout(n7619));
  jand g07428(.dina(n7342), .dinb(n7339), .dout(n7620));
  jor  g07429(.dina(n7620), .dinb(n7619), .dout(n7621));
  jand g07430(.dina(n7508), .dinb(n7505), .dout(n7622));
  jand g07431(.dina(n7501), .dinb(n7503), .dout(n7623));
  jor  g07432(.dina(n7623), .dinb(n7622), .dout(n7624));
  jxor g07433(.dina(n7624), .dinb(n7621), .dout(n7625));
  jand g07434(.dina(n7358), .dinb(n7148), .dout(n7626));
  jand g07435(.dina(n7362), .dinb(n7359), .dout(n7627));
  jor  g07436(.dina(n7627), .dinb(n7626), .dout(n7628));
  jxor g07437(.dina(n7628), .dinb(n7625), .dout(n7629));
  jand g07438(.dina(n7439), .dinb(n7392), .dout(n7630));
  jand g07439(.dina(n7478), .dinb(n7440), .dout(n7631));
  jor  g07440(.dina(n7631), .dinb(n7630), .dout(n7632));
  jxor g07441(.dina(n7632), .dinb(n7629), .dout(n7633));
  jxor g07442(.dina(n7633), .dinb(n7617), .dout(n7634));
  jxor g07443(.dina(n7634), .dinb(n7597), .dout(n7635));
  jand g07444(.dina(n7527), .dinb(n7511), .dout(n7636));
  jand g07445(.dina(n7528), .dinb(n7491), .dout(n7637));
  jor  g07446(.dina(n7637), .dinb(n7636), .dout(n7638));
  jand g07447(.dina(\a[54] ), .dinb(\a[8] ), .dout(n7639));
  jnot g07448(.din(n7639), .dout(n7640));
  jand g07449(.dina(\a[44] ), .dinb(\a[18] ), .dout(n7641));
  jnot g07450(.din(n7641), .dout(n7642));
  jand g07451(.dina(n7642), .dinb(n7640), .dout(n7643));
  jand g07452(.dina(n7641), .dinb(n7639), .dout(n7644));
  jnot g07453(.din(n7644), .dout(n7645));
  jand g07454(.dina(n4495), .dinb(n1024), .dout(n7646));
  jand g07455(.dina(\a[43] ), .dinb(\a[19] ), .dout(n7647));
  jand g07456(.dina(n7647), .dinb(n7639), .dout(n7648));
  jor  g07457(.dina(n7648), .dinb(n7646), .dout(n7649));
  jnot g07458(.din(n7649), .dout(n7650));
  jand g07459(.dina(n7650), .dinb(n7645), .dout(n7651));
  jnot g07460(.din(n7651), .dout(n7652));
  jor  g07461(.dina(n7652), .dinb(n7643), .dout(n7653));
  jand g07462(.dina(n7649), .dinb(n7645), .dout(n7654));
  jnot g07463(.din(n7654), .dout(n7655));
  jand g07464(.dina(n7655), .dinb(n7647), .dout(n7656));
  jnot g07465(.din(n7656), .dout(n7657));
  jand g07466(.dina(n7657), .dinb(n7653), .dout(n7658));
  jand g07467(.dina(\a[35] ), .dinb(\a[27] ), .dout(n7659));
  jnot g07468(.din(n7659), .dout(n7660));
  jand g07469(.dina(n3634), .dinb(n2653), .dout(n7661));
  jnot g07470(.din(n7661), .dout(n7662));
  jand g07471(.dina(\a[34] ), .dinb(\a[28] ), .dout(n7663));
  jand g07472(.dina(\a[33] ), .dinb(\a[29] ), .dout(n7664));
  jor  g07473(.dina(n7664), .dinb(n7663), .dout(n7665));
  jand g07474(.dina(n7665), .dinb(n7662), .dout(n7666));
  jxor g07475(.dina(n7666), .dinb(n7660), .dout(n7667));
  jxor g07476(.dina(n7667), .dinb(n7658), .dout(n7668));
  jnot g07477(.din(n7668), .dout(n7669));
  jand g07478(.dina(\a[40] ), .dinb(\a[22] ), .dout(n7670));
  jnot g07479(.din(n7670), .dout(n7671));
  jand g07480(.dina(\a[39] ), .dinb(\a[24] ), .dout(n7672));
  jand g07481(.dina(n7672), .dinb(n7518), .dout(n7673));
  jnot g07482(.din(n7673), .dout(n7674));
  jand g07483(.dina(\a[39] ), .dinb(\a[23] ), .dout(n7675));
  jand g07484(.dina(\a[38] ), .dinb(\a[24] ), .dout(n7676));
  jor  g07485(.dina(n7676), .dinb(n7675), .dout(n7677));
  jand g07486(.dina(n7677), .dinb(n7674), .dout(n7678));
  jxor g07487(.dina(n7678), .dinb(n7671), .dout(n7679));
  jxor g07488(.dina(n7679), .dinb(n7669), .dout(n7680));
  jand g07489(.dina(\a[53] ), .dinb(\a[9] ), .dout(n7681));
  jand g07490(.dina(\a[52] ), .dinb(\a[45] ), .dout(n7682));
  jand g07491(.dina(n7682), .dinb(n1601), .dout(n7683));
  jnot g07492(.din(n7683), .dout(n7684));
  jand g07493(.dina(n7165), .dinb(n453), .dout(n7685));
  jand g07494(.dina(\a[45] ), .dinb(\a[17] ), .dout(n7686));
  jand g07495(.dina(n7686), .dinb(n7681), .dout(n7687));
  jor  g07496(.dina(n7687), .dinb(n7685), .dout(n7688));
  jand g07497(.dina(n7688), .dinb(n7684), .dout(n7689));
  jnot g07498(.din(n7689), .dout(n7690));
  jand g07499(.dina(n7690), .dinb(n7681), .dout(n7691));
  jor  g07500(.dina(n7688), .dinb(n7683), .dout(n7692));
  jnot g07501(.din(n7692), .dout(n7693));
  jand g07502(.dina(\a[52] ), .dinb(\a[10] ), .dout(n7694));
  jor  g07503(.dina(n7694), .dinb(n7686), .dout(n7695));
  jand g07504(.dina(n7695), .dinb(n7693), .dout(n7696));
  jor  g07505(.dina(n7696), .dinb(n7691), .dout(n7697));
  jand g07506(.dina(n7500), .dinb(\a[31] ), .dout(n7698));
  jand g07507(.dina(\a[62] ), .dinb(\a[0] ), .dout(n7699));
  jand g07508(.dina(\a[60] ), .dinb(\a[2] ), .dout(n7700));
  jor  g07509(.dina(n7700), .dinb(n7699), .dout(n7701));
  jand g07510(.dina(\a[62] ), .dinb(\a[2] ), .dout(n7702));
  jand g07511(.dina(n7702), .dinb(n7153), .dout(n7703));
  jnot g07512(.din(n7703), .dout(n7704));
  jand g07513(.dina(n7704), .dinb(n7701), .dout(n7705));
  jxor g07514(.dina(n7705), .dinb(n7698), .dout(n7706));
  jnot g07515(.din(n7706), .dout(n7707));
  jand g07516(.dina(\a[41] ), .dinb(\a[21] ), .dout(n7708));
  jnot g07517(.din(n7708), .dout(n7709));
  jand g07518(.dina(n3138), .dinb(n2128), .dout(n7710));
  jnot g07519(.din(n7710), .dout(n7711));
  jand g07520(.dina(\a[36] ), .dinb(\a[26] ), .dout(n7712));
  jand g07521(.dina(\a[37] ), .dinb(\a[25] ), .dout(n7713));
  jor  g07522(.dina(n7713), .dinb(n7712), .dout(n7714));
  jand g07523(.dina(n7714), .dinb(n7711), .dout(n7715));
  jxor g07524(.dina(n7715), .dinb(n7709), .dout(n7716));
  jxor g07525(.dina(n7716), .dinb(n7707), .dout(n7717));
  jxor g07526(.dina(n7717), .dinb(n7697), .dout(n7718));
  jand g07527(.dina(\a[51] ), .dinb(\a[47] ), .dout(n7719));
  jand g07528(.dina(n7719), .dinb(n1469), .dout(n7720));
  jnot g07529(.din(n7720), .dout(n7721));
  jand g07530(.dina(\a[51] ), .dinb(\a[11] ), .dout(n7722));
  jand g07531(.dina(\a[47] ), .dinb(\a[15] ), .dout(n7723));
  jor  g07532(.dina(n7723), .dinb(n7722), .dout(n7724));
  jand g07533(.dina(n7724), .dinb(n7721), .dout(n7725));
  jxor g07534(.dina(n7725), .dinb(n7396), .dout(n7726));
  jnot g07535(.din(n7726), .dout(n7727));
  jnot g07536(.din(n7417), .dout(n7728));
  jand g07537(.dina(\a[49] ), .dinb(\a[48] ), .dout(n7729));
  jand g07538(.dina(n7729), .dinb(n675), .dout(n7730));
  jnot g07539(.din(n7730), .dout(n7731));
  jand g07540(.dina(\a[49] ), .dinb(\a[13] ), .dout(n7732));
  jand g07541(.dina(\a[48] ), .dinb(\a[14] ), .dout(n7733));
  jor  g07542(.dina(n7733), .dinb(n7732), .dout(n7734));
  jand g07543(.dina(n7734), .dinb(n7731), .dout(n7735));
  jxor g07544(.dina(n7735), .dinb(n7728), .dout(n7736));
  jxor g07545(.dina(n7736), .dinb(n7727), .dout(n7737));
  jand g07546(.dina(\a[42] ), .dinb(\a[20] ), .dout(n7738));
  jand g07547(.dina(\a[56] ), .dinb(\a[7] ), .dout(n7739));
  jand g07548(.dina(n7739), .dinb(n7458), .dout(n7740));
  jnot g07549(.din(n7740), .dout(n7741));
  jand g07550(.dina(\a[56] ), .dinb(\a[6] ), .dout(n7742));
  jand g07551(.dina(\a[55] ), .dinb(\a[7] ), .dout(n7743));
  jor  g07552(.dina(n7743), .dinb(n7742), .dout(n7744));
  jand g07553(.dina(n7744), .dinb(n7741), .dout(n7745));
  jxor g07554(.dina(n7745), .dinb(n7738), .dout(n7746));
  jxor g07555(.dina(n7746), .dinb(n7737), .dout(n7747));
  jxor g07556(.dina(n7747), .dinb(n7718), .dout(n7748));
  jxor g07557(.dina(n7748), .dinb(n7680), .dout(n7749));
  jxor g07558(.dina(n7749), .dinb(n7638), .dout(n7750));
  jnot g07559(.din(n7351), .dout(n7751));
  jand g07560(.dina(n7378), .dinb(n7751), .dout(n7752));
  jnot g07561(.din(n7752), .dout(n7753));
  jand g07562(.dina(n7377), .dinb(n7351), .dout(n7754));
  jor  g07563(.dina(n7754), .dinb(n7338), .dout(n7755));
  jand g07564(.dina(n7755), .dinb(n7753), .dout(n7756));
  jxor g07565(.dina(n7756), .dinb(n7750), .dout(n7757));
  jxor g07566(.dina(n7757), .dinb(n7635), .dout(n7758));
  jor  g07567(.dina(n7380), .dinb(n7335), .dout(n7759));
  jand g07568(.dina(n7481), .dinb(n7381), .dout(n7760));
  jnot g07569(.din(n7760), .dout(n7761));
  jand g07570(.dina(n7761), .dinb(n7759), .dout(n7762));
  jnot g07571(.din(n7762), .dout(n7763));
  jand g07572(.dina(n7574), .dinb(n7537), .dout(n7764));
  jand g07573(.dina(n7575), .dinb(n7534), .dout(n7765));
  jor  g07574(.dina(n7765), .dinb(n7764), .dout(n7766));
  jand g07575(.dina(n7368), .dinb(n7366), .dout(n7767));
  jand g07576(.dina(n7374), .dinb(n7369), .dout(n7768));
  jor  g07577(.dina(n7768), .dinb(n7767), .dout(n7769));
  jnot g07578(.din(n7769), .dout(n7770));
  jand g07579(.dina(n7467), .dinb(n7457), .dout(n7771));
  jnot g07580(.din(n7771), .dout(n7772));
  jor  g07581(.dina(n7477), .dinb(n7469), .dout(n7773));
  jand g07582(.dina(n7773), .dinb(n7772), .dout(n7774));
  jxor g07583(.dina(n7774), .dinb(n7770), .dout(n7775));
  jand g07584(.dina(n7428), .dinb(n7410), .dout(n7776));
  jand g07585(.dina(n7438), .dinb(n7429), .dout(n7777));
  jor  g07586(.dina(n7777), .dinb(n7776), .dout(n7778));
  jxor g07587(.dina(n7778), .dinb(n7775), .dout(n7779));
  jand g07588(.dina(n7562), .dinb(n7555), .dout(n7780));
  jor  g07589(.dina(n7780), .dinb(n7560), .dout(n7781));
  jnot g07590(.din(n7451), .dout(n7782));
  jand g07591(.dina(n7461), .dinb(n7459), .dout(n7783));
  jnot g07592(.din(n7783), .dout(n7784));
  jand g07593(.dina(n7784), .dinb(n7464), .dout(n7785));
  jxor g07594(.dina(n7785), .dinb(n7782), .dout(n7786));
  jxor g07595(.dina(n7786), .dinb(n7781), .dout(n7787));
  jor  g07596(.dina(n7520), .dinb(n7518), .dout(n7788));
  jand g07597(.dina(n7788), .dinb(n7523), .dout(n7789));
  jand g07598(.dina(n7569), .dinb(n7567), .dout(n7790));
  jnot g07599(.din(n7790), .dout(n7791));
  jand g07600(.dina(n7791), .dinb(n7571), .dout(n7792));
  jxor g07601(.dina(n7792), .dinb(n7789), .dout(n7793));
  jand g07602(.dina(n7472), .dinb(n7470), .dout(n7794));
  jnot g07603(.din(n7794), .dout(n7795));
  jand g07604(.dina(n7795), .dinb(n7475), .dout(n7796));
  jxor g07605(.dina(n7796), .dinb(n7793), .dout(n7797));
  jand g07606(.dina(\a[61] ), .dinb(\a[1] ), .dout(n7798));
  jxor g07607(.dina(n7798), .dinb(n3118), .dout(n7799));
  jand g07608(.dina(n7433), .dinb(n7431), .dout(n7800));
  jnot g07609(.din(n7800), .dout(n7801));
  jand g07610(.dina(n7801), .dinb(n7435), .dout(n7802));
  jxor g07611(.dina(n7802), .dinb(n7799), .dout(n7803));
  jxor g07612(.dina(n7803), .dinb(n7423), .dout(n7804));
  jxor g07613(.dina(n7804), .dinb(n7797), .dout(n7805));
  jxor g07614(.dina(n7805), .dinb(n7787), .dout(n7806));
  jxor g07615(.dina(n7806), .dinb(n7779), .dout(n7807));
  jxor g07616(.dina(n7807), .dinb(n7766), .dout(n7808));
  jand g07617(.dina(n7375), .dinb(n7363), .dout(n7809));
  jand g07618(.dina(n7376), .dinb(n7355), .dout(n7810));
  jor  g07619(.dina(n7810), .dinb(n7809), .dout(n7811));
  jand g07620(.dina(n7509), .dinb(n7499), .dout(n7812));
  jand g07621(.dina(n7510), .dinb(n7496), .dout(n7813));
  jor  g07622(.dina(n7813), .dinb(n7812), .dout(n7814));
  jxor g07623(.dina(n7814), .dinb(n7811), .dout(n7815));
  jand g07624(.dina(n7346), .dinb(n7343), .dout(n7816));
  jand g07625(.dina(n7350), .dinb(n7347), .dout(n7817));
  jor  g07626(.dina(n7817), .dinb(n7816), .dout(n7818));
  jxor g07627(.dina(n7818), .dinb(n7815), .dout(n7819));
  jand g07628(.dina(n7479), .dinb(n7389), .dout(n7820));
  jand g07629(.dina(n7480), .dinb(n7384), .dout(n7821));
  jor  g07630(.dina(n7821), .dinb(n7820), .dout(n7822));
  jxor g07631(.dina(n7822), .dinb(n7819), .dout(n7823));
  jxor g07632(.dina(n7823), .dinb(n7808), .dout(n7824));
  jxor g07633(.dina(n7824), .dinb(n7763), .dout(n7825));
  jxor g07634(.dina(n7825), .dinb(n7758), .dout(n7826));
  jand g07635(.dina(n7826), .dinb(n7594), .dout(n7827));
  jor  g07636(.dina(n7826), .dinb(n7594), .dout(n7828));
  jnot g07637(.din(n7828), .dout(n7829));
  jor  g07638(.dina(n7829), .dinb(n7827), .dout(n7830));
  jnot g07639(.din(n7581), .dout(n7831));
  jor  g07640(.dina(n7590), .dinb(n7583), .dout(n7832));
  jand g07641(.dina(n7832), .dinb(n7831), .dout(n7833));
  jxor g07642(.dina(n7833), .dinb(n7830), .dout(\asquared[63] ));
  jand g07643(.dina(n7824), .dinb(n7763), .dout(n7835));
  jand g07644(.dina(n7825), .dinb(n7758), .dout(n7836));
  jor  g07645(.dina(n7836), .dinb(n7835), .dout(n7837));
  jand g07646(.dina(n7634), .dinb(n7597), .dout(n7838));
  jand g07647(.dina(n7757), .dinb(n7635), .dout(n7839));
  jor  g07648(.dina(n7839), .dinb(n7838), .dout(n7840));
  jand g07649(.dina(n7749), .dinb(n7638), .dout(n7841));
  jand g07650(.dina(n7756), .dinb(n7750), .dout(n7842));
  jor  g07651(.dina(n7842), .dinb(n7841), .dout(n7843));
  jand g07652(.dina(n7804), .dinb(n7797), .dout(n7844));
  jand g07653(.dina(n7805), .dinb(n7787), .dout(n7845));
  jor  g07654(.dina(n7845), .dinb(n7844), .dout(n7846));
  jnot g07655(.din(n7846), .dout(n7847));
  jor  g07656(.dina(n7774), .dinb(n7770), .dout(n7848));
  jand g07657(.dina(n7778), .dinb(n7775), .dout(n7849));
  jnot g07658(.din(n7849), .dout(n7850));
  jand g07659(.dina(n7850), .dinb(n7848), .dout(n7851));
  jxor g07660(.dina(n7851), .dinb(n7847), .dout(n7852));
  jand g07661(.dina(n7612), .dinb(n7602), .dout(n7853));
  jand g07662(.dina(n7616), .dinb(n7613), .dout(n7854));
  jor  g07663(.dina(n7854), .dinb(n7853), .dout(n7855));
  jxor g07664(.dina(n7855), .dinb(n7852), .dout(n7856));
  jnot g07665(.din(n7403), .dout(n7857));
  jand g07666(.dina(n7549), .dinb(n7857), .dout(n7858));
  jand g07667(.dina(n7611), .dinb(n7603), .dout(n7859));
  jor  g07668(.dina(n7859), .dinb(n7858), .dout(n7860));
  jand g07669(.dina(n7792), .dinb(n7789), .dout(n7861));
  jand g07670(.dina(n7796), .dinb(n7793), .dout(n7862));
  jor  g07671(.dina(n7862), .dinb(n7861), .dout(n7863));
  jxor g07672(.dina(n7863), .dinb(n7860), .dout(n7864));
  jand g07673(.dina(n7802), .dinb(n7799), .dout(n7865));
  jand g07674(.dina(n7803), .dinb(n7423), .dout(n7866));
  jor  g07675(.dina(n7866), .dinb(n7865), .dout(n7867));
  jxor g07676(.dina(n7867), .dinb(n7864), .dout(n7868));
  jand g07677(.dina(n7747), .dinb(n7718), .dout(n7869));
  jand g07678(.dina(n7748), .dinb(n7680), .dout(n7870));
  jor  g07679(.dina(n7870), .dinb(n7869), .dout(n7871));
  jxor g07680(.dina(n7871), .dinb(n7868), .dout(n7872));
  jand g07681(.dina(n7674), .dinb(n7671), .dout(n7873));
  jnot g07682(.din(n7873), .dout(n7874));
  jand g07683(.dina(n7874), .dinb(n7677), .dout(n7875));
  jor  g07684(.dina(n7740), .dinb(n7738), .dout(n7876));
  jand g07685(.dina(n7876), .dinb(n7744), .dout(n7877));
  jxor g07686(.dina(n7877), .dinb(n7875), .dout(n7878));
  jand g07687(.dina(n7731), .dinb(n7728), .dout(n7879));
  jnot g07688(.din(n7879), .dout(n7880));
  jand g07689(.dina(n7880), .dinb(n7734), .dout(n7881));
  jxor g07690(.dina(n7881), .dinb(n7878), .dout(n7882));
  jand g07691(.dina(n7705), .dinb(n7698), .dout(n7883));
  jor  g07692(.dina(n7883), .dinb(n7703), .dout(n7884));
  jnot g07693(.din(n7604), .dout(n7885));
  jand g07694(.dina(n7606), .dinb(n7885), .dout(n7886));
  jnot g07695(.din(n7886), .dout(n7887));
  jand g07696(.dina(n7887), .dinb(n7609), .dout(n7888));
  jand g07697(.dina(n7711), .dinb(n7709), .dout(n7889));
  jnot g07698(.din(n7889), .dout(n7890));
  jand g07699(.dina(n7890), .dinb(n7714), .dout(n7891));
  jxor g07700(.dina(n7891), .dinb(n7888), .dout(n7892));
  jxor g07701(.dina(n7892), .dinb(n7884), .dout(n7893));
  jand g07702(.dina(n7785), .dinb(n7782), .dout(n7894));
  jand g07703(.dina(n7786), .dinb(n7781), .dout(n7895));
  jor  g07704(.dina(n7895), .dinb(n7894), .dout(n7896));
  jxor g07705(.dina(n7896), .dinb(n7893), .dout(n7897));
  jxor g07706(.dina(n7897), .dinb(n7882), .dout(n7898));
  jxor g07707(.dina(n7898), .dinb(n7872), .dout(n7899));
  jxor g07708(.dina(n7899), .dinb(n7856), .dout(n7900));
  jxor g07709(.dina(n7900), .dinb(n7843), .dout(n7901));
  jxor g07710(.dina(n7901), .dinb(n7840), .dout(n7902));
  jand g07711(.dina(n7822), .dinb(n7819), .dout(n7903));
  jand g07712(.dina(n7823), .dinb(n7808), .dout(n7904));
  jor  g07713(.dina(n7904), .dinb(n7903), .dout(n7905));
  jand g07714(.dina(n7814), .dinb(n7811), .dout(n7906));
  jand g07715(.dina(n7818), .dinb(n7815), .dout(n7907));
  jor  g07716(.dina(n7907), .dinb(n7906), .dout(n7908));
  jand g07717(.dina(n7662), .dinb(n7660), .dout(n7909));
  jnot g07718(.din(n7909), .dout(n7910));
  jand g07719(.dina(n7910), .dinb(n7665), .dout(n7911));
  jxor g07720(.dina(n7911), .dinb(n7692), .dout(n7912));
  jxor g07721(.dina(n7912), .dinb(n7652), .dout(n7913));
  jnot g07722(.din(n7913), .dout(n7914));
  jor  g07723(.dina(n7667), .dinb(n7658), .dout(n7915));
  jor  g07724(.dina(n7679), .dinb(n7669), .dout(n7916));
  jand g07725(.dina(n7916), .dinb(n7915), .dout(n7917));
  jxor g07726(.dina(n7917), .dinb(n7914), .dout(n7918));
  jnot g07727(.din(n7918), .dout(n7919));
  jor  g07728(.dina(n7736), .dinb(n7727), .dout(n7920));
  jand g07729(.dina(n7746), .dinb(n7737), .dout(n7921));
  jnot g07730(.din(n7921), .dout(n7922));
  jand g07731(.dina(n7922), .dinb(n7920), .dout(n7923));
  jxor g07732(.dina(n7923), .dinb(n7919), .dout(n7924));
  jand g07733(.dina(n7624), .dinb(n7621), .dout(n7925));
  jand g07734(.dina(n7628), .dinb(n7625), .dout(n7926));
  jor  g07735(.dina(n7926), .dinb(n7925), .dout(n7927));
  jnot g07736(.din(n7927), .dout(n7928));
  jor  g07737(.dina(n7716), .dinb(n7707), .dout(n7929));
  jand g07738(.dina(n7717), .dinb(n7697), .dout(n7930));
  jnot g07739(.din(n7930), .dout(n7931));
  jand g07740(.dina(n7931), .dinb(n7929), .dout(n7932));
  jxor g07741(.dina(n7932), .dinb(n7928), .dout(n7933));
  jand g07742(.dina(\a[38] ), .dinb(\a[26] ), .dout(n7934));
  jand g07743(.dina(n7934), .dinb(n7713), .dout(n7935));
  jnot g07744(.din(n7935), .dout(n7936));
  jand g07745(.dina(\a[37] ), .dinb(\a[26] ), .dout(n7937));
  jand g07746(.dina(\a[38] ), .dinb(\a[25] ), .dout(n7938));
  jor  g07747(.dina(n7938), .dinb(n7937), .dout(n7939));
  jand g07748(.dina(n7939), .dinb(n7936), .dout(n7940));
  jxor g07749(.dina(n7940), .dinb(n7672), .dout(n7941));
  jnot g07750(.din(n7941), .dout(n7942));
  jand g07751(.dina(\a[36] ), .dinb(\a[27] ), .dout(n7943));
  jnot g07752(.din(n7943), .dout(n7944));
  jand g07753(.dina(n2845), .dinb(n2653), .dout(n7945));
  jnot g07754(.din(n7945), .dout(n7946));
  jand g07755(.dina(\a[35] ), .dinb(\a[28] ), .dout(n7947));
  jor  g07756(.dina(n7947), .dinb(n3183), .dout(n7948));
  jand g07757(.dina(n7948), .dinb(n7946), .dout(n7949));
  jxor g07758(.dina(n7949), .dinb(n7944), .dout(n7950));
  jxor g07759(.dina(n7950), .dinb(n7942), .dout(n7951));
  jand g07760(.dina(n2296), .dinb(\a[62] ), .dout(n7952));
  jnot g07761(.din(n7952), .dout(n7953));
  jand g07762(.dina(n7953), .dinb(\a[32] ), .dout(n7954));
  jand g07763(.dina(\a[62] ), .dinb(\a[32] ), .dout(n7955));
  jnot g07764(.din(n7955), .dout(n7956));
  jand g07765(.dina(n7956), .dinb(\a[1] ), .dout(n7957));
  jand g07766(.dina(n7957), .dinb(\a[62] ), .dout(n7958));
  jor  g07767(.dina(n7958), .dinb(n7954), .dout(n7959));
  jand g07768(.dina(n7798), .dinb(n3118), .dout(n7960));
  jand g07769(.dina(\a[63] ), .dinb(\a[0] ), .dout(n7961));
  jxor g07770(.dina(n7961), .dinb(n7960), .dout(n7962));
  jxor g07771(.dina(n7962), .dinb(n7959), .dout(n7963));
  jxor g07772(.dina(n7963), .dinb(n7951), .dout(n7964));
  jxor g07773(.dina(n7964), .dinb(n7933), .dout(n7965));
  jxor g07774(.dina(n7965), .dinb(n7924), .dout(n7966));
  jxor g07775(.dina(n7966), .dinb(n7908), .dout(n7967));
  jxor g07776(.dina(n7967), .dinb(n7905), .dout(n7968));
  jand g07777(.dina(n7806), .dinb(n7779), .dout(n7969));
  jand g07778(.dina(n7807), .dinb(n7766), .dout(n7970));
  jor  g07779(.dina(n7970), .dinb(n7969), .dout(n7971));
  jand g07780(.dina(n7632), .dinb(n7629), .dout(n7972));
  jand g07781(.dina(n7633), .dinb(n7617), .dout(n7973));
  jor  g07782(.dina(n7973), .dinb(n7972), .dout(n7974));
  jand g07783(.dina(\a[48] ), .dinb(\a[15] ), .dout(n7975));
  jand g07784(.dina(n5594), .dinb(n899), .dout(n7976));
  jnot g07785(.din(n7976), .dout(n7977));
  jand g07786(.dina(\a[50] ), .dinb(\a[48] ), .dout(n7978));
  jand g07787(.dina(n7978), .dinb(n727), .dout(n7979));
  jand g07788(.dina(\a[51] ), .dinb(\a[12] ), .dout(n7980));
  jand g07789(.dina(n7980), .dinb(n7975), .dout(n7981));
  jor  g07790(.dina(n7981), .dinb(n7979), .dout(n7982));
  jand g07791(.dina(n7982), .dinb(n7977), .dout(n7983));
  jnot g07792(.din(n7983), .dout(n7984));
  jand g07793(.dina(n7984), .dinb(n7975), .dout(n7985));
  jor  g07794(.dina(n7982), .dinb(n7976), .dout(n7986));
  jnot g07795(.din(n7986), .dout(n7987));
  jand g07796(.dina(\a[50] ), .dinb(\a[13] ), .dout(n7988));
  jor  g07797(.dina(n7988), .dinb(n7980), .dout(n7989));
  jand g07798(.dina(n7989), .dinb(n7987), .dout(n7990));
  jor  g07799(.dina(n7990), .dinb(n7985), .dout(n7991));
  jand g07800(.dina(\a[54] ), .dinb(\a[46] ), .dout(n7992));
  jand g07801(.dina(n7992), .dinb(n1465), .dout(n7993));
  jnot g07802(.din(n7993), .dout(n7994));
  jand g07803(.dina(\a[54] ), .dinb(\a[9] ), .dout(n7995));
  jand g07804(.dina(\a[45] ), .dinb(\a[18] ), .dout(n7996));
  jand g07805(.dina(n7996), .dinb(n7995), .dout(n7997));
  jand g07806(.dina(\a[46] ), .dinb(\a[18] ), .dout(n7998));
  jand g07807(.dina(n7998), .dinb(n7686), .dout(n7999));
  jor  g07808(.dina(n7999), .dinb(n7997), .dout(n8000));
  jnot g07809(.din(n8000), .dout(n8001));
  jand g07810(.dina(n8001), .dinb(n7994), .dout(n8002));
  jand g07811(.dina(\a[46] ), .dinb(\a[17] ), .dout(n8003));
  jor  g07812(.dina(n8003), .dinb(n7995), .dout(n8004));
  jand g07813(.dina(n8004), .dinb(n8002), .dout(n8005));
  jnot g07814(.din(n8005), .dout(n8006));
  jnot g07815(.din(n7996), .dout(n8007));
  jand g07816(.dina(n8000), .dinb(n7994), .dout(n8008));
  jor  g07817(.dina(n8008), .dinb(n8007), .dout(n8009));
  jand g07818(.dina(n8009), .dinb(n8006), .dout(n8010));
  jnot g07819(.din(n8010), .dout(n8011));
  jand g07820(.dina(\a[53] ), .dinb(\a[10] ), .dout(n8012));
  jand g07821(.dina(\a[52] ), .dinb(\a[47] ), .dout(n8013));
  jand g07822(.dina(n8013), .dinb(n1580), .dout(n8014));
  jnot g07823(.din(n8014), .dout(n8015));
  jand g07824(.dina(n7165), .dinb(n655), .dout(n8016));
  jand g07825(.dina(\a[47] ), .dinb(\a[16] ), .dout(n8017));
  jand g07826(.dina(n8017), .dinb(n8012), .dout(n8018));
  jor  g07827(.dina(n8018), .dinb(n8016), .dout(n8019));
  jand g07828(.dina(n8019), .dinb(n8015), .dout(n8020));
  jnot g07829(.din(n8020), .dout(n8021));
  jand g07830(.dina(n8021), .dinb(n8012), .dout(n8022));
  jand g07831(.dina(\a[52] ), .dinb(\a[11] ), .dout(n8023));
  jor  g07832(.dina(n8023), .dinb(n8017), .dout(n8024));
  jor  g07833(.dina(n8019), .dinb(n8014), .dout(n8025));
  jnot g07834(.din(n8025), .dout(n8026));
  jand g07835(.dina(n8026), .dinb(n8024), .dout(n8027));
  jor  g07836(.dina(n8027), .dinb(n8022), .dout(n8028));
  jxor g07837(.dina(n8028), .dinb(n8011), .dout(n8029));
  jxor g07838(.dina(n8029), .dinb(n7991), .dout(n8030));
  jand g07839(.dina(n7725), .dinb(n7396), .dout(n8031));
  jor  g07840(.dina(n8031), .dinb(n7720), .dout(n8032));
  jnot g07841(.din(n8032), .dout(n8033));
  jnot g07842(.din(n7445), .dout(n8034));
  jand g07843(.dina(\a[60] ), .dinb(\a[4] ), .dout(n8035));
  jand g07844(.dina(n8035), .dinb(n7604), .dout(n8036));
  jnot g07845(.din(n8036), .dout(n8037));
  jand g07846(.dina(\a[60] ), .dinb(\a[3] ), .dout(n8038));
  jand g07847(.dina(\a[59] ), .dinb(\a[4] ), .dout(n8039));
  jor  g07848(.dina(n8039), .dinb(n8038), .dout(n8040));
  jand g07849(.dina(n8040), .dinb(n8037), .dout(n8041));
  jxor g07850(.dina(n8041), .dinb(n8034), .dout(n8042));
  jxor g07851(.dina(n8042), .dinb(n8033), .dout(n8043));
  jnot g07852(.din(n8043), .dout(n8044));
  jand g07853(.dina(\a[58] ), .dinb(\a[5] ), .dout(n8045));
  jnot g07854(.din(n8045), .dout(n8046));
  jand g07855(.dina(n4514), .dinb(n1376), .dout(n8047));
  jnot g07856(.din(n8047), .dout(n8048));
  jand g07857(.dina(\a[41] ), .dinb(\a[22] ), .dout(n8049));
  jand g07858(.dina(\a[42] ), .dinb(\a[21] ), .dout(n8050));
  jor  g07859(.dina(n8050), .dinb(n8049), .dout(n8051));
  jand g07860(.dina(n8051), .dinb(n8048), .dout(n8052));
  jxor g07861(.dina(n8052), .dinb(n8046), .dout(n8053));
  jxor g07862(.dina(n8053), .dinb(n8044), .dout(n8054));
  jand g07863(.dina(\a[40] ), .dinb(\a[23] ), .dout(n8055));
  jand g07864(.dina(\a[57] ), .dinb(\a[6] ), .dout(n8056));
  jand g07865(.dina(\a[43] ), .dinb(\a[20] ), .dout(n8057));
  jxor g07866(.dina(n8057), .dinb(n8056), .dout(n8058));
  jxor g07867(.dina(n8058), .dinb(n8055), .dout(n8059));
  jand g07868(.dina(\a[49] ), .dinb(\a[14] ), .dout(n8060));
  jand g07869(.dina(\a[33] ), .dinb(\a[30] ), .dout(n8061));
  jxor g07870(.dina(n8061), .dinb(n3269), .dout(n8062));
  jxor g07871(.dina(n8062), .dinb(n8060), .dout(n8063));
  jxor g07872(.dina(n8063), .dinb(n8059), .dout(n8064));
  jnot g07873(.din(n8064), .dout(n8065));
  jnot g07874(.din(n7739), .dout(n8066));
  jand g07875(.dina(\a[55] ), .dinb(\a[44] ), .dout(n8067));
  jand g07876(.dina(n8067), .dinb(n1597), .dout(n8068));
  jnot g07877(.din(n8068), .dout(n8069));
  jand g07878(.dina(\a[55] ), .dinb(\a[8] ), .dout(n8070));
  jand g07879(.dina(\a[44] ), .dinb(\a[19] ), .dout(n8071));
  jor  g07880(.dina(n8071), .dinb(n8070), .dout(n8072));
  jand g07881(.dina(n8072), .dinb(n8069), .dout(n8073));
  jxor g07882(.dina(n8073), .dinb(n8066), .dout(n8074));
  jxor g07883(.dina(n8074), .dinb(n8065), .dout(n8075));
  jxor g07884(.dina(n8075), .dinb(n8054), .dout(n8076));
  jxor g07885(.dina(n8076), .dinb(n8030), .dout(n8077));
  jxor g07886(.dina(n8077), .dinb(n7974), .dout(n8078));
  jxor g07887(.dina(n8078), .dinb(n7971), .dout(n8079));
  jxor g07888(.dina(n8079), .dinb(n7968), .dout(n8080));
  jxor g07889(.dina(n8080), .dinb(n7902), .dout(n8081));
  jnot g07890(.din(n8081), .dout(n8082));
  jxor g07891(.dina(n8082), .dinb(n7837), .dout(n8083));
  jnot g07892(.din(n7827), .dout(n8084));
  jor  g07893(.dina(n7833), .dinb(n7829), .dout(n8085));
  jand g07894(.dina(n8085), .dinb(n8084), .dout(n8086));
  jxor g07895(.dina(n8086), .dinb(n8083), .dout(\asquared[64] ));
  jand g07896(.dina(n7899), .dinb(n7856), .dout(n8088));
  jand g07897(.dina(n7900), .dinb(n7843), .dout(n8089));
  jor  g07898(.dina(n8089), .dinb(n8088), .dout(n8090));
  jand g07899(.dina(n7940), .dinb(n7672), .dout(n8091));
  jor  g07900(.dina(n8091), .dinb(n7935), .dout(n8092));
  jxor g07901(.dina(n8092), .dinb(n7986), .dout(n8093));
  jxor g07902(.dina(n8093), .dinb(n8025), .dout(n8094));
  jnot g07903(.din(n8094), .dout(n8095));
  jand g07904(.dina(n8063), .dinb(n8059), .dout(n8096));
  jnot g07905(.din(n8096), .dout(n8097));
  jor  g07906(.dina(n8074), .dinb(n8065), .dout(n8098));
  jand g07907(.dina(n8098), .dinb(n8097), .dout(n8099));
  jxor g07908(.dina(n8099), .dinb(n8095), .dout(n8100));
  jand g07909(.dina(n8028), .dinb(n8011), .dout(n8101));
  jand g07910(.dina(n8029), .dinb(n7991), .dout(n8102));
  jor  g07911(.dina(n8102), .dinb(n8101), .dout(n8103));
  jxor g07912(.dina(n8103), .dinb(n8100), .dout(n8104));
  jnot g07913(.din(n8104), .dout(n8105));
  jor  g07914(.dina(n7851), .dinb(n7847), .dout(n8106));
  jand g07915(.dina(n7855), .dinb(n7852), .dout(n8107));
  jnot g07916(.din(n8107), .dout(n8108));
  jand g07917(.dina(n8108), .dinb(n8106), .dout(n8109));
  jxor g07918(.dina(n8109), .dinb(n8105), .dout(n8110));
  jand g07919(.dina(n7863), .dinb(n7860), .dout(n8111));
  jand g07920(.dina(n7867), .dinb(n7864), .dout(n8112));
  jor  g07921(.dina(n8112), .dinb(n8111), .dout(n8113));
  jor  g07922(.dina(n8042), .dinb(n8033), .dout(n8114));
  jor  g07923(.dina(n8053), .dinb(n8044), .dout(n8115));
  jand g07924(.dina(n8115), .dinb(n8114), .dout(n8116));
  jnot g07925(.din(n8116), .dout(n8117));
  jxor g07926(.dina(n8117), .dinb(n8113), .dout(n8118));
  jor  g07927(.dina(n8061), .dinb(n3269), .dout(n8119));
  jand g07928(.dina(n8061), .dinb(n3269), .dout(n8120));
  jor  g07929(.dina(n8120), .dinb(n8060), .dout(n8121));
  jand g07930(.dina(n8121), .dinb(n8119), .dout(n8122));
  jnot g07931(.din(\a[63] ), .dout(n8123));
  jand g07932(.dina(n7953), .dinb(n8123), .dout(n8124));
  jnot g07933(.din(n8124), .dout(n8125));
  jor  g07934(.dina(n7957), .dinb(n8123), .dout(n8126));
  jand g07935(.dina(n8126), .dinb(n8125), .dout(n8127));
  jxor g07936(.dina(n8127), .dinb(n8122), .dout(n8128));
  jand g07937(.dina(\a[55] ), .dinb(\a[9] ), .dout(n8129));
  jand g07938(.dina(\a[54] ), .dinb(\a[10] ), .dout(n8130));
  jand g07939(.dina(\a[49] ), .dinb(\a[15] ), .dout(n8131));
  jxor g07940(.dina(n8131), .dinb(n8130), .dout(n8132));
  jxor g07941(.dina(n8132), .dinb(n8129), .dout(n8133));
  jnot g07942(.din(n8133), .dout(n8134));
  jand g07943(.dina(\a[51] ), .dinb(\a[13] ), .dout(n8135));
  jnot g07944(.din(n8135), .dout(n8136));
  jand g07945(.dina(n7165), .dinb(n555), .dout(n8137));
  jnot g07946(.din(n8137), .dout(n8138));
  jand g07947(.dina(\a[53] ), .dinb(\a[11] ), .dout(n8139));
  jand g07948(.dina(\a[52] ), .dinb(\a[12] ), .dout(n8140));
  jor  g07949(.dina(n8140), .dinb(n8139), .dout(n8141));
  jand g07950(.dina(n8141), .dinb(n8138), .dout(n8142));
  jxor g07951(.dina(n8142), .dinb(n8136), .dout(n8143));
  jxor g07952(.dina(n8143), .dinb(n8134), .dout(n8144));
  jxor g07953(.dina(n8144), .dinb(n8128), .dout(n8145));
  jxor g07954(.dina(n8145), .dinb(n8118), .dout(n8146));
  jxor g07955(.dina(n8146), .dinb(n8110), .dout(n8147));
  jxor g07956(.dina(n8147), .dinb(n8090), .dout(n8148));
  jand g07957(.dina(n7871), .dinb(n7868), .dout(n8149));
  jand g07958(.dina(n7898), .dinb(n7872), .dout(n8150));
  jor  g07959(.dina(n8150), .dinb(n8149), .dout(n8151));
  jand g07960(.dina(\a[47] ), .dinb(\a[17] ), .dout(n8152));
  jnot g07961(.din(n8152), .dout(n8153));
  jand g07962(.dina(\a[57] ), .dinb(\a[7] ), .dout(n8154));
  jnot g07963(.din(n8154), .dout(n8155));
  jand g07964(.dina(n8155), .dinb(n8153), .dout(n8156));
  jand g07965(.dina(n8154), .dinb(n8152), .dout(n8157));
  jnot g07966(.din(n8157), .dout(n8158));
  jand g07967(.dina(\a[58] ), .dinb(\a[6] ), .dout(n8159));
  jand g07968(.dina(n8159), .dinb(n8152), .dout(n8160));
  jand g07969(.dina(n7519), .dinb(n410), .dout(n8161));
  jor  g07970(.dina(n8161), .dinb(n8160), .dout(n8162));
  jnot g07971(.din(n8162), .dout(n8163));
  jand g07972(.dina(n8163), .dinb(n8158), .dout(n8164));
  jnot g07973(.din(n8164), .dout(n8165));
  jor  g07974(.dina(n8165), .dinb(n8156), .dout(n8166));
  jnot g07975(.din(n8159), .dout(n8167));
  jand g07976(.dina(n8162), .dinb(n8158), .dout(n8168));
  jor  g07977(.dina(n8168), .dinb(n8167), .dout(n8169));
  jand g07978(.dina(n8169), .dinb(n8166), .dout(n8170));
  jand g07979(.dina(\a[44] ), .dinb(\a[20] ), .dout(n8171));
  jnot g07980(.din(n8171), .dout(n8172));
  jand g07981(.dina(n4317), .dinb(n1376), .dout(n8173));
  jnot g07982(.din(n8173), .dout(n8174));
  jand g07983(.dina(\a[43] ), .dinb(\a[21] ), .dout(n8175));
  jand g07984(.dina(\a[42] ), .dinb(\a[22] ), .dout(n8176));
  jor  g07985(.dina(n8176), .dinb(n8175), .dout(n8177));
  jand g07986(.dina(n8177), .dinb(n8174), .dout(n8178));
  jxor g07987(.dina(n8178), .dinb(n8172), .dout(n8179));
  jxor g07988(.dina(n8179), .dinb(n8170), .dout(n8180));
  jnot g07989(.din(n8180), .dout(n8181));
  jand g07990(.dina(\a[41] ), .dinb(\a[23] ), .dout(n8182));
  jnot g07991(.din(n8182), .dout(n8183));
  jand g07992(.dina(n3665), .dinb(n1648), .dout(n8184));
  jnot g07993(.din(n8184), .dout(n8185));
  jand g07994(.dina(\a[40] ), .dinb(\a[24] ), .dout(n8186));
  jand g07995(.dina(\a[39] ), .dinb(\a[25] ), .dout(n8187));
  jor  g07996(.dina(n8187), .dinb(n8186), .dout(n8188));
  jand g07997(.dina(n8188), .dinb(n8185), .dout(n8189));
  jxor g07998(.dina(n8189), .dinb(n8183), .dout(n8190));
  jxor g07999(.dina(n8190), .dinb(n8181), .dout(n8191));
  jand g08000(.dina(n7961), .dinb(n7960), .dout(n8192));
  jand g08001(.dina(n7962), .dinb(n7959), .dout(n8193));
  jor  g08002(.dina(n8193), .dinb(n8192), .dout(n8194));
  jand g08003(.dina(\a[59] ), .dinb(\a[5] ), .dout(n8195));
  jand g08004(.dina(\a[46] ), .dinb(\a[19] ), .dout(n8196));
  jand g08005(.dina(n8196), .dinb(n7996), .dout(n8197));
  jnot g08006(.din(n8197), .dout(n8198));
  jand g08007(.dina(\a[45] ), .dinb(\a[19] ), .dout(n8199));
  jor  g08008(.dina(n8199), .dinb(n7998), .dout(n8200));
  jand g08009(.dina(n8200), .dinb(n8198), .dout(n8201));
  jxor g08010(.dina(n8201), .dinb(n8195), .dout(n8202));
  jxor g08011(.dina(n8202), .dinb(n8194), .dout(n8203));
  jand g08012(.dina(\a[61] ), .dinb(\a[4] ), .dout(n8204));
  jand g08013(.dina(n8204), .dinb(n8038), .dout(n8205));
  jnot g08014(.din(n8205), .dout(n8206));
  jand g08015(.dina(\a[61] ), .dinb(\a[3] ), .dout(n8207));
  jor  g08016(.dina(n8207), .dinb(n8035), .dout(n8208));
  jand g08017(.dina(n8208), .dinb(n8206), .dout(n8209));
  jxor g08018(.dina(n8209), .dinb(n7702), .dout(n8210));
  jxor g08019(.dina(n8210), .dinb(n8203), .dout(n8211));
  jand g08020(.dina(\a[48] ), .dinb(\a[16] ), .dout(n8212));
  jand g08021(.dina(\a[56] ), .dinb(\a[8] ), .dout(n8213));
  jor  g08022(.dina(n8213), .dinb(n8212), .dout(n8214));
  jand g08023(.dina(\a[56] ), .dinb(\a[48] ), .dout(n8215));
  jand g08024(.dina(n8215), .dinb(n1297), .dout(n8216));
  jnot g08025(.din(n8216), .dout(n8217));
  jand g08026(.dina(n8217), .dinb(n8214), .dout(n8218));
  jxor g08027(.dina(n8218), .dinb(n7934), .dout(n8219));
  jnot g08028(.din(n8219), .dout(n8220));
  jand g08029(.dina(\a[37] ), .dinb(\a[27] ), .dout(n8221));
  jnot g08030(.din(n8221), .dout(n8222));
  jand g08031(.dina(n3243), .dinb(n2653), .dout(n8223));
  jnot g08032(.din(n8223), .dout(n8224));
  jand g08033(.dina(\a[36] ), .dinb(\a[28] ), .dout(n8225));
  jand g08034(.dina(\a[35] ), .dinb(\a[29] ), .dout(n8226));
  jor  g08035(.dina(n8226), .dinb(n8225), .dout(n8227));
  jand g08036(.dina(n8227), .dinb(n8224), .dout(n8228));
  jxor g08037(.dina(n8228), .dinb(n8222), .dout(n8229));
  jxor g08038(.dina(n8229), .dinb(n8220), .dout(n8230));
  jnot g08039(.din(n8230), .dout(n8231));
  jand g08040(.dina(\a[50] ), .dinb(\a[14] ), .dout(n8232));
  jnot g08041(.din(n8232), .dout(n8233));
  jand g08042(.dina(n3634), .dinb(n2440), .dout(n8234));
  jnot g08043(.din(n8234), .dout(n8235));
  jand g08044(.dina(\a[34] ), .dinb(\a[30] ), .dout(n8236));
  jand g08045(.dina(\a[33] ), .dinb(\a[31] ), .dout(n8237));
  jor  g08046(.dina(n8237), .dinb(n8236), .dout(n8238));
  jand g08047(.dina(n8238), .dinb(n8235), .dout(n8239));
  jxor g08048(.dina(n8239), .dinb(n8233), .dout(n8240));
  jxor g08049(.dina(n8240), .dinb(n8231), .dout(n8241));
  jxor g08050(.dina(n8241), .dinb(n8211), .dout(n8242));
  jxor g08051(.dina(n8242), .dinb(n8191), .dout(n8243));
  jxor g08052(.dina(n8243), .dinb(n8151), .dout(n8244));
  jand g08053(.dina(n7877), .dinb(n7875), .dout(n8245));
  jand g08054(.dina(n7881), .dinb(n7878), .dout(n8246));
  jor  g08055(.dina(n8246), .dinb(n8245), .dout(n8247));
  jand g08056(.dina(n7911), .dinb(n7692), .dout(n8248));
  jand g08057(.dina(n7912), .dinb(n7652), .dout(n8249));
  jor  g08058(.dina(n8249), .dinb(n8248), .dout(n8250));
  jxor g08059(.dina(n8250), .dinb(n8247), .dout(n8251));
  jand g08060(.dina(n7891), .dinb(n7888), .dout(n8252));
  jand g08061(.dina(n7892), .dinb(n7884), .dout(n8253));
  jor  g08062(.dina(n8253), .dinb(n8252), .dout(n8254));
  jxor g08063(.dina(n8254), .dinb(n8251), .dout(n8255));
  jor  g08064(.dina(n7917), .dinb(n7914), .dout(n8256));
  jor  g08065(.dina(n7923), .dinb(n7919), .dout(n8257));
  jand g08066(.dina(n8257), .dinb(n8256), .dout(n8258));
  jnot g08067(.din(n8258), .dout(n8259));
  jand g08068(.dina(n7896), .dinb(n7893), .dout(n8260));
  jand g08069(.dina(n7897), .dinb(n7882), .dout(n8261));
  jor  g08070(.dina(n8261), .dinb(n8260), .dout(n8262));
  jxor g08071(.dina(n8262), .dinb(n8259), .dout(n8263));
  jxor g08072(.dina(n8263), .dinb(n8255), .dout(n8264));
  jxor g08073(.dina(n8264), .dinb(n8244), .dout(n8265));
  jxor g08074(.dina(n8265), .dinb(n8148), .dout(n8266));
  jand g08075(.dina(n7967), .dinb(n7905), .dout(n8267));
  jand g08076(.dina(n8079), .dinb(n7968), .dout(n8268));
  jor  g08077(.dina(n8268), .dinb(n8267), .dout(n8269));
  jand g08078(.dina(n8077), .dinb(n7974), .dout(n8270));
  jand g08079(.dina(n8078), .dinb(n7971), .dout(n8271));
  jor  g08080(.dina(n8271), .dinb(n8270), .dout(n8272));
  jand g08081(.dina(n7965), .dinb(n7924), .dout(n8273));
  jand g08082(.dina(n7966), .dinb(n7908), .dout(n8274));
  jor  g08083(.dina(n8274), .dinb(n8273), .dout(n8275));
  jand g08084(.dina(n8075), .dinb(n8054), .dout(n8276));
  jand g08085(.dina(n8076), .dinb(n8030), .dout(n8277));
  jor  g08086(.dina(n8277), .dinb(n8276), .dout(n8278));
  jnot g08087(.din(n8278), .dout(n8279));
  jor  g08088(.dina(n7932), .dinb(n7928), .dout(n8280));
  jand g08089(.dina(n7964), .dinb(n7933), .dout(n8281));
  jnot g08090(.din(n8281), .dout(n8282));
  jand g08091(.dina(n8282), .dinb(n8280), .dout(n8283));
  jxor g08092(.dina(n8283), .dinb(n8279), .dout(n8284));
  jor  g08093(.dina(n7950), .dinb(n7942), .dout(n8285));
  jand g08094(.dina(n7963), .dinb(n7951), .dout(n8286));
  jnot g08095(.din(n8286), .dout(n8287));
  jand g08096(.dina(n8287), .dinb(n8285), .dout(n8288));
  jnot g08097(.din(n8288), .dout(n8289));
  jnot g08098(.din(n8002), .dout(n8290));
  jand g08099(.dina(n8057), .dinb(n8056), .dout(n8291));
  jand g08100(.dina(n8058), .dinb(n8055), .dout(n8292));
  jor  g08101(.dina(n8292), .dinb(n8291), .dout(n8293));
  jxor g08102(.dina(n8293), .dinb(n8290), .dout(n8294));
  jand g08103(.dina(n7946), .dinb(n7944), .dout(n8295));
  jnot g08104(.din(n8295), .dout(n8296));
  jand g08105(.dina(n8296), .dinb(n7948), .dout(n8297));
  jxor g08106(.dina(n8297), .dinb(n8294), .dout(n8298));
  jand g08107(.dina(n8048), .dinb(n8046), .dout(n8299));
  jnot g08108(.din(n8299), .dout(n8300));
  jand g08109(.dina(n8300), .dinb(n8051), .dout(n8301));
  jand g08110(.dina(n8037), .dinb(n8034), .dout(n8302));
  jnot g08111(.din(n8302), .dout(n8303));
  jand g08112(.dina(n8303), .dinb(n8040), .dout(n8304));
  jxor g08113(.dina(n8304), .dinb(n8301), .dout(n8305));
  jand g08114(.dina(n8069), .dinb(n8066), .dout(n8306));
  jnot g08115(.din(n8306), .dout(n8307));
  jand g08116(.dina(n8307), .dinb(n8072), .dout(n8308));
  jxor g08117(.dina(n8308), .dinb(n8305), .dout(n8309));
  jxor g08118(.dina(n8309), .dinb(n8298), .dout(n8310));
  jxor g08119(.dina(n8310), .dinb(n8289), .dout(n8311));
  jxor g08120(.dina(n8311), .dinb(n8284), .dout(n8312));
  jxor g08121(.dina(n8312), .dinb(n8275), .dout(n8313));
  jxor g08122(.dina(n8313), .dinb(n8272), .dout(n8314));
  jxor g08123(.dina(n8314), .dinb(n8269), .dout(n8315));
  jxor g08124(.dina(n8315), .dinb(n8266), .dout(n8316));
  jand g08125(.dina(n7901), .dinb(n7840), .dout(n8317));
  jand g08126(.dina(n8080), .dinb(n7902), .dout(n8318));
  jor  g08127(.dina(n8318), .dinb(n8317), .dout(n8319));
  jnot g08128(.din(n8319), .dout(n8320));
  jxor g08129(.dina(n8320), .dinb(n8316), .dout(n8321));
  jand g08130(.dina(n8081), .dinb(n7837), .dout(n8322));
  jnot g08131(.din(n8322), .dout(n8323));
  jnot g08132(.din(n7837), .dout(n8324));
  jand g08133(.dina(n8082), .dinb(n8324), .dout(n8325));
  jor  g08134(.dina(n8086), .dinb(n8325), .dout(n8326));
  jand g08135(.dina(n8326), .dinb(n8323), .dout(n8327));
  jxor g08136(.dina(n8327), .dinb(n8321), .dout(\asquared[65] ));
  jand g08137(.dina(n8314), .dinb(n8269), .dout(n8329));
  jand g08138(.dina(n8315), .dinb(n8266), .dout(n8330));
  jor  g08139(.dina(n8330), .dinb(n8329), .dout(n8331));
  jand g08140(.dina(n8147), .dinb(n8090), .dout(n8332));
  jand g08141(.dina(n8265), .dinb(n8148), .dout(n8333));
  jor  g08142(.dina(n8333), .dinb(n8332), .dout(n8334));
  jand g08143(.dina(n8243), .dinb(n8151), .dout(n8335));
  jand g08144(.dina(n8264), .dinb(n8244), .dout(n8336));
  jor  g08145(.dina(n8336), .dinb(n8335), .dout(n8337));
  jor  g08146(.dina(n8109), .dinb(n8105), .dout(n8338));
  jand g08147(.dina(n8146), .dinb(n8110), .dout(n8339));
  jnot g08148(.din(n8339), .dout(n8340));
  jand g08149(.dina(n8340), .dinb(n8338), .dout(n8341));
  jnot g08150(.din(n8341), .dout(n8342));
  jand g08151(.dina(n8241), .dinb(n8211), .dout(n8343));
  jand g08152(.dina(n8242), .dinb(n8191), .dout(n8344));
  jor  g08153(.dina(n8344), .dinb(n8343), .dout(n8345));
  jand g08154(.dina(n8117), .dinb(n8113), .dout(n8346));
  jand g08155(.dina(n8145), .dinb(n8118), .dout(n8347));
  jor  g08156(.dina(n8347), .dinb(n8346), .dout(n8348));
  jxor g08157(.dina(n8348), .dinb(n8345), .dout(n8349));
  jor  g08158(.dina(n8143), .dinb(n8134), .dout(n8350));
  jand g08159(.dina(n8144), .dinb(n8128), .dout(n8351));
  jnot g08160(.din(n8351), .dout(n8352));
  jand g08161(.dina(n8352), .dinb(n8350), .dout(n8353));
  jnot g08162(.din(n8353), .dout(n8354));
  jand g08163(.dina(n8131), .dinb(n8130), .dout(n8355));
  jand g08164(.dina(n8132), .dinb(n8129), .dout(n8356));
  jor  g08165(.dina(n8356), .dinb(n8355), .dout(n8357));
  jand g08166(.dina(n8185), .dinb(n8183), .dout(n8358));
  jnot g08167(.din(n8358), .dout(n8359));
  jand g08168(.dina(n8359), .dinb(n8188), .dout(n8360));
  jxor g08169(.dina(n8360), .dinb(n8357), .dout(n8361));
  jxor g08170(.dina(n8361), .dinb(n8165), .dout(n8362));
  jand g08171(.dina(n8218), .dinb(n7934), .dout(n8363));
  jor  g08172(.dina(n8363), .dinb(n8216), .dout(n8364));
  jand g08173(.dina(n8208), .dinb(n7702), .dout(n8365));
  jor  g08174(.dina(n8365), .dinb(n8205), .dout(n8366));
  jand g08175(.dina(n8201), .dinb(n8195), .dout(n8367));
  jor  g08176(.dina(n8367), .dinb(n8197), .dout(n8368));
  jxor g08177(.dina(n8368), .dinb(n8366), .dout(n8369));
  jxor g08178(.dina(n8369), .dinb(n8364), .dout(n8370));
  jxor g08179(.dina(n8370), .dinb(n8362), .dout(n8371));
  jxor g08180(.dina(n8371), .dinb(n8354), .dout(n8372));
  jxor g08181(.dina(n8372), .dinb(n8349), .dout(n8373));
  jxor g08182(.dina(n8373), .dinb(n8342), .dout(n8374));
  jxor g08183(.dina(n8374), .dinb(n8337), .dout(n8375));
  jxor g08184(.dina(n8375), .dinb(n8334), .dout(n8376));
  jand g08185(.dina(n8312), .dinb(n8275), .dout(n8377));
  jand g08186(.dina(n8313), .dinb(n8272), .dout(n8378));
  jor  g08187(.dina(n8378), .dinb(n8377), .dout(n8379));
  jand g08188(.dina(n8250), .dinb(n8247), .dout(n8380));
  jand g08189(.dina(n8254), .dinb(n8251), .dout(n8381));
  jor  g08190(.dina(n8381), .dinb(n8380), .dout(n8382));
  jand g08191(.dina(n8202), .dinb(n8194), .dout(n8383));
  jand g08192(.dina(n8210), .dinb(n8203), .dout(n8384));
  jor  g08193(.dina(n8384), .dinb(n8383), .dout(n8385));
  jxor g08194(.dina(n8385), .dinb(n8382), .dout(n8386));
  jand g08195(.dina(\a[63] ), .dinb(\a[61] ), .dout(n8387));
  jand g08196(.dina(n8387), .dinb(n245), .dout(n8388));
  jnot g08197(.din(n8388), .dout(n8389));
  jand g08198(.dina(\a[63] ), .dinb(\a[2] ), .dout(n8390));
  jor  g08199(.dina(n8390), .dinb(n8204), .dout(n8391));
  jand g08200(.dina(n8391), .dinb(n8389), .dout(n8392));
  jand g08201(.dina(n8235), .dinb(n8233), .dout(n8393));
  jnot g08202(.din(n8393), .dout(n8394));
  jand g08203(.dina(n8394), .dinb(n8238), .dout(n8395));
  jxor g08204(.dina(n8395), .dinb(n8392), .dout(n8396));
  jand g08205(.dina(\a[52] ), .dinb(\a[13] ), .dout(n8397));
  jand g08206(.dina(\a[47] ), .dinb(\a[18] ), .dout(n8398));
  jand g08207(.dina(n8398), .dinb(n8397), .dout(n8399));
  jnot g08208(.din(n8399), .dout(n8400));
  jand g08209(.dina(n7165), .dinb(n899), .dout(n8401));
  jand g08210(.dina(\a[53] ), .dinb(\a[12] ), .dout(n8402));
  jand g08211(.dina(n8402), .dinb(n8398), .dout(n8403));
  jor  g08212(.dina(n8403), .dinb(n8401), .dout(n8404));
  jnot g08213(.din(n8404), .dout(n8405));
  jand g08214(.dina(n8405), .dinb(n8400), .dout(n8406));
  jor  g08215(.dina(n8398), .dinb(n8397), .dout(n8407));
  jand g08216(.dina(n8407), .dinb(n8406), .dout(n8408));
  jand g08217(.dina(n8404), .dinb(n8400), .dout(n8409));
  jnot g08218(.din(n8409), .dout(n8410));
  jand g08219(.dina(n8410), .dinb(n8402), .dout(n8411));
  jor  g08220(.dina(n8411), .dinb(n8408), .dout(n8412));
  jand g08221(.dina(\a[49] ), .dinb(\a[16] ), .dout(n8413));
  jnot g08222(.din(n8413), .dout(n8414));
  jand g08223(.dina(n5594), .dinb(n976), .dout(n8415));
  jnot g08224(.din(n8415), .dout(n8416));
  jand g08225(.dina(\a[51] ), .dinb(\a[14] ), .dout(n8417));
  jand g08226(.dina(\a[50] ), .dinb(\a[15] ), .dout(n8418));
  jor  g08227(.dina(n8418), .dinb(n8417), .dout(n8419));
  jand g08228(.dina(n8419), .dinb(n8416), .dout(n8420));
  jxor g08229(.dina(n8420), .dinb(n8414), .dout(n8421));
  jnot g08230(.din(n8421), .dout(n8422));
  jxor g08231(.dina(n8422), .dinb(n8412), .dout(n8423));
  jxor g08232(.dina(n8423), .dinb(n8396), .dout(n8424));
  jxor g08233(.dina(n8424), .dinb(n8386), .dout(n8425));
  jand g08234(.dina(n8174), .dinb(n8172), .dout(n8426));
  jnot g08235(.din(n8426), .dout(n8427));
  jand g08236(.dina(n8427), .dinb(n8177), .dout(n8428));
  jand g08237(.dina(n8224), .dinb(n8222), .dout(n8429));
  jnot g08238(.din(n8429), .dout(n8430));
  jand g08239(.dina(n8430), .dinb(n8227), .dout(n8431));
  jxor g08240(.dina(n8431), .dinb(n8428), .dout(n8432));
  jand g08241(.dina(n8138), .dinb(n8136), .dout(n8433));
  jnot g08242(.din(n8433), .dout(n8434));
  jand g08243(.dina(n8434), .dinb(n8141), .dout(n8435));
  jxor g08244(.dina(n8435), .dinb(n8432), .dout(n8436));
  jnot g08245(.din(n8436), .dout(n8437));
  jor  g08246(.dina(n8229), .dinb(n8220), .dout(n8438));
  jor  g08247(.dina(n8240), .dinb(n8231), .dout(n8439));
  jand g08248(.dina(n8439), .dinb(n8438), .dout(n8440));
  jxor g08249(.dina(n8440), .dinb(n8437), .dout(n8441));
  jnot g08250(.din(n8441), .dout(n8442));
  jor  g08251(.dina(n8179), .dinb(n8170), .dout(n8443));
  jor  g08252(.dina(n8190), .dinb(n8181), .dout(n8444));
  jand g08253(.dina(n8444), .dinb(n8443), .dout(n8445));
  jxor g08254(.dina(n8445), .dinb(n8442), .dout(n8446));
  jand g08255(.dina(n8262), .dinb(n8259), .dout(n8447));
  jand g08256(.dina(n8263), .dinb(n8255), .dout(n8448));
  jor  g08257(.dina(n8448), .dinb(n8447), .dout(n8449));
  jxor g08258(.dina(n8449), .dinb(n8446), .dout(n8450));
  jxor g08259(.dina(n8450), .dinb(n8425), .dout(n8451));
  jxor g08260(.dina(n8451), .dinb(n8379), .dout(n8452));
  jand g08261(.dina(n8092), .dinb(n7986), .dout(n8453));
  jand g08262(.dina(n8093), .dinb(n8025), .dout(n8454));
  jor  g08263(.dina(n8454), .dinb(n8453), .dout(n8455));
  jand g08264(.dina(n8293), .dinb(n8290), .dout(n8456));
  jand g08265(.dina(n8297), .dinb(n8294), .dout(n8457));
  jor  g08266(.dina(n8457), .dinb(n8456), .dout(n8458));
  jxor g08267(.dina(n8458), .dinb(n8455), .dout(n8459));
  jand g08268(.dina(n8304), .dinb(n8301), .dout(n8460));
  jand g08269(.dina(n8308), .dinb(n8305), .dout(n8461));
  jor  g08270(.dina(n8461), .dinb(n8460), .dout(n8462));
  jxor g08271(.dina(n8462), .dinb(n8459), .dout(n8463));
  jand g08272(.dina(n8309), .dinb(n8298), .dout(n8464));
  jand g08273(.dina(n8310), .dinb(n8289), .dout(n8465));
  jor  g08274(.dina(n8465), .dinb(n8464), .dout(n8466));
  jor  g08275(.dina(n8099), .dinb(n8095), .dout(n8467));
  jand g08276(.dina(n8103), .dinb(n8100), .dout(n8468));
  jnot g08277(.din(n8468), .dout(n8469));
  jand g08278(.dina(n8469), .dinb(n8467), .dout(n8470));
  jnot g08279(.din(n8470), .dout(n8471));
  jxor g08280(.dina(n8471), .dinb(n8466), .dout(n8472));
  jxor g08281(.dina(n8472), .dinb(n8463), .dout(n8473));
  jor  g08282(.dina(n8283), .dinb(n8279), .dout(n8474));
  jand g08283(.dina(n8311), .dinb(n8284), .dout(n8475));
  jnot g08284(.din(n8475), .dout(n8476));
  jand g08285(.dina(n8476), .dinb(n8474), .dout(n8477));
  jnot g08286(.din(n8477), .dout(n8478));
  jand g08287(.dina(\a[55] ), .dinb(\a[10] ), .dout(n8479));
  jand g08288(.dina(\a[45] ), .dinb(\a[20] ), .dout(n8480));
  jand g08289(.dina(n8480), .dinb(n8479), .dout(n8481));
  jnot g08290(.din(n8481), .dout(n8482));
  jand g08291(.dina(\a[56] ), .dinb(\a[9] ), .dout(n8483));
  jand g08292(.dina(n8483), .dinb(n8480), .dout(n8484));
  jand g08293(.dina(\a[56] ), .dinb(\a[10] ), .dout(n8485));
  jand g08294(.dina(n8485), .dinb(n8129), .dout(n8486));
  jor  g08295(.dina(n8486), .dinb(n8484), .dout(n8487));
  jnot g08296(.din(n8487), .dout(n8488));
  jand g08297(.dina(n8488), .dinb(n8482), .dout(n8489));
  jor  g08298(.dina(n8480), .dinb(n8479), .dout(n8490));
  jand g08299(.dina(n8490), .dinb(n8489), .dout(n8491));
  jand g08300(.dina(n8487), .dinb(n8482), .dout(n8492));
  jnot g08301(.din(n8492), .dout(n8493));
  jand g08302(.dina(n8493), .dinb(n8483), .dout(n8494));
  jor  g08303(.dina(n8494), .dinb(n8491), .dout(n8495));
  jand g08304(.dina(\a[42] ), .dinb(\a[23] ), .dout(n8496));
  jnot g08305(.din(n8496), .dout(n8497));
  jand g08306(.dina(n4632), .dinb(n1648), .dout(n8498));
  jnot g08307(.din(n8498), .dout(n8499));
  jand g08308(.dina(\a[41] ), .dinb(\a[24] ), .dout(n8500));
  jand g08309(.dina(\a[40] ), .dinb(\a[25] ), .dout(n8501));
  jor  g08310(.dina(n8501), .dinb(n8500), .dout(n8502));
  jand g08311(.dina(n8502), .dinb(n8499), .dout(n8503));
  jxor g08312(.dina(n8503), .dinb(n8497), .dout(n8504));
  jnot g08313(.din(n8504), .dout(n8505));
  jxor g08314(.dina(n8505), .dinb(n8495), .dout(n8506));
  jnot g08315(.din(n8506), .dout(n8507));
  jand g08316(.dina(\a[39] ), .dinb(\a[26] ), .dout(n8508));
  jnot g08317(.din(n8508), .dout(n8509));
  jand g08318(.dina(\a[38] ), .dinb(\a[28] ), .dout(n8510));
  jand g08319(.dina(n8510), .dinb(n8221), .dout(n8511));
  jnot g08320(.din(n8511), .dout(n8512));
  jand g08321(.dina(\a[38] ), .dinb(\a[27] ), .dout(n8513));
  jand g08322(.dina(\a[37] ), .dinb(\a[28] ), .dout(n8514));
  jor  g08323(.dina(n8514), .dinb(n8513), .dout(n8515));
  jand g08324(.dina(n8515), .dinb(n8512), .dout(n8516));
  jxor g08325(.dina(n8516), .dinb(n8509), .dout(n8517));
  jxor g08326(.dina(n8517), .dinb(n8507), .dout(n8518));
  jand g08327(.dina(n8127), .dinb(n8122), .dout(n8519));
  jand g08328(.dina(n7952), .dinb(\a[63] ), .dout(n8520));
  jor  g08329(.dina(n8520), .dinb(n8519), .dout(n8521));
  jand g08330(.dina(\a[57] ), .dinb(\a[8] ), .dout(n8522));
  jand g08331(.dina(n4495), .dinb(n1376), .dout(n8523));
  jnot g08332(.din(n8523), .dout(n8524));
  jand g08333(.dina(\a[44] ), .dinb(\a[21] ), .dout(n8525));
  jand g08334(.dina(\a[43] ), .dinb(\a[22] ), .dout(n8526));
  jor  g08335(.dina(n8526), .dinb(n8525), .dout(n8527));
  jand g08336(.dina(n8527), .dinb(n8524), .dout(n8528));
  jxor g08337(.dina(n8528), .dinb(n8522), .dout(n8529));
  jxor g08338(.dina(n8529), .dinb(n8521), .dout(n8530));
  jnot g08339(.din(n8530), .dout(n8531));
  jand g08340(.dina(\a[60] ), .dinb(\a[5] ), .dout(n8532));
  jnot g08341(.din(n8532), .dout(n8533));
  jand g08342(.dina(\a[59] ), .dinb(\a[7] ), .dout(n8534));
  jand g08343(.dina(n8534), .dinb(n8159), .dout(n8535));
  jnot g08344(.din(n8535), .dout(n8536));
  jand g08345(.dina(\a[59] ), .dinb(\a[6] ), .dout(n8537));
  jand g08346(.dina(\a[58] ), .dinb(\a[7] ), .dout(n8538));
  jor  g08347(.dina(n8538), .dinb(n8537), .dout(n8539));
  jand g08348(.dina(n8539), .dinb(n8536), .dout(n8540));
  jxor g08349(.dina(n8540), .dinb(n8533), .dout(n8541));
  jxor g08350(.dina(n8541), .dinb(n8531), .dout(n8542));
  jand g08351(.dina(n3634), .dinb(n3269), .dout(n8543));
  jnot g08352(.din(n8543), .dout(n8544));
  jand g08353(.dina(n3476), .dinb(n2671), .dout(n8545));
  jand g08354(.dina(n2845), .dinb(n2440), .dout(n8546));
  jor  g08355(.dina(n8546), .dinb(n8545), .dout(n8547));
  jand g08356(.dina(n8547), .dinb(n8544), .dout(n8548));
  jnot g08357(.din(n8548), .dout(n8549));
  jand g08358(.dina(n8549), .dinb(n3476), .dout(n8550));
  jor  g08359(.dina(n8547), .dinb(n8543), .dout(n8551));
  jnot g08360(.din(n8551), .dout(n8552));
  jand g08361(.dina(\a[34] ), .dinb(\a[31] ), .dout(n8553));
  jor  g08362(.dina(n8553), .dinb(n2671), .dout(n8554));
  jand g08363(.dina(n8554), .dinb(n8552), .dout(n8555));
  jor  g08364(.dina(n8555), .dinb(n8550), .dout(n8556));
  jand g08365(.dina(\a[36] ), .dinb(\a[29] ), .dout(n8557));
  jand g08366(.dina(\a[54] ), .dinb(\a[11] ), .dout(n8558));
  jxor g08367(.dina(n8558), .dinb(n8196), .dout(n8559));
  jxor g08368(.dina(n8559), .dinb(n8557), .dout(n8560));
  jxor g08369(.dina(n8560), .dinb(n8556), .dout(n8561));
  jand g08370(.dina(\a[48] ), .dinb(\a[17] ), .dout(n8562));
  jand g08371(.dina(\a[62] ), .dinb(\a[3] ), .dout(n8563));
  jxor g08372(.dina(n8563), .dinb(\a[33] ), .dout(n8564));
  jxor g08373(.dina(n8564), .dinb(n8562), .dout(n8565));
  jxor g08374(.dina(n8565), .dinb(n8561), .dout(n8566));
  jxor g08375(.dina(n8566), .dinb(n8542), .dout(n8567));
  jxor g08376(.dina(n8567), .dinb(n8518), .dout(n8568));
  jxor g08377(.dina(n8568), .dinb(n8478), .dout(n8569));
  jxor g08378(.dina(n8569), .dinb(n8473), .dout(n8570));
  jxor g08379(.dina(n8570), .dinb(n8452), .dout(n8571));
  jxor g08380(.dina(n8571), .dinb(n8376), .dout(n8572));
  jand g08381(.dina(n8572), .dinb(n8331), .dout(n8573));
  jor  g08382(.dina(n8572), .dinb(n8331), .dout(n8574));
  jnot g08383(.din(n8574), .dout(n8575));
  jor  g08384(.dina(n8575), .dinb(n8573), .dout(n8576));
  jand g08385(.dina(n8319), .dinb(n8316), .dout(n8577));
  jnot g08386(.din(n8577), .dout(n8578));
  jnot g08387(.din(n8316), .dout(n8579));
  jand g08388(.dina(n8320), .dinb(n8579), .dout(n8580));
  jor  g08389(.dina(n8327), .dinb(n8580), .dout(n8581));
  jand g08390(.dina(n8581), .dinb(n8578), .dout(n8582));
  jxor g08391(.dina(n8582), .dinb(n8576), .dout(\asquared[66] ));
  jand g08392(.dina(n8375), .dinb(n8334), .dout(n8584));
  jand g08393(.dina(n8571), .dinb(n8376), .dout(n8585));
  jor  g08394(.dina(n8585), .dinb(n8584), .dout(n8586));
  jand g08395(.dina(n8451), .dinb(n8379), .dout(n8587));
  jand g08396(.dina(n8570), .dinb(n8452), .dout(n8588));
  jor  g08397(.dina(n8588), .dinb(n8587), .dout(n8589));
  jand g08398(.dina(n8471), .dinb(n8466), .dout(n8590));
  jand g08399(.dina(n8472), .dinb(n8463), .dout(n8591));
  jor  g08400(.dina(n8591), .dinb(n8590), .dout(n8592));
  jand g08401(.dina(n8458), .dinb(n8455), .dout(n8593));
  jand g08402(.dina(n8462), .dinb(n8459), .dout(n8594));
  jor  g08403(.dina(n8594), .dinb(n8593), .dout(n8595));
  jand g08404(.dina(n8422), .dinb(n8412), .dout(n8596));
  jand g08405(.dina(n8423), .dinb(n8396), .dout(n8597));
  jor  g08406(.dina(n8597), .dinb(n8596), .dout(n8598));
  jand g08407(.dina(n8395), .dinb(n8392), .dout(n8599));
  jor  g08408(.dina(n8599), .dinb(n8388), .dout(n8600));
  jand g08409(.dina(n8512), .dinb(n8509), .dout(n8601));
  jnot g08410(.din(n8601), .dout(n8602));
  jand g08411(.dina(n8602), .dinb(n8515), .dout(n8603));
  jxor g08412(.dina(n8603), .dinb(n8600), .dout(n8604));
  jnot g08413(.din(n8604), .dout(n8605));
  jand g08414(.dina(\a[60] ), .dinb(\a[6] ), .dout(n8606));
  jnot g08415(.din(n8606), .dout(n8607));
  jand g08416(.dina(\a[59] ), .dinb(\a[8] ), .dout(n8608));
  jand g08417(.dina(n8608), .dinb(n8538), .dout(n8609));
  jnot g08418(.din(n8609), .dout(n8610));
  jand g08419(.dina(\a[58] ), .dinb(\a[8] ), .dout(n8611));
  jor  g08420(.dina(n8611), .dinb(n8534), .dout(n8612));
  jand g08421(.dina(n8612), .dinb(n8610), .dout(n8613));
  jxor g08422(.dina(n8613), .dinb(n8607), .dout(n8614));
  jxor g08423(.dina(n8614), .dinb(n8605), .dout(n8615));
  jxor g08424(.dina(n8615), .dinb(n8598), .dout(n8616));
  jxor g08425(.dina(n8616), .dinb(n8595), .dout(n8617));
  jand g08426(.dina(n8563), .dinb(\a[33] ), .dout(n8618));
  jand g08427(.dina(n8564), .dinb(n8562), .dout(n8619));
  jor  g08428(.dina(n8619), .dinb(n8618), .dout(n8620));
  jxor g08429(.dina(n8620), .dinb(n8551), .dout(n8621));
  jand g08430(.dina(n8416), .dinb(n8414), .dout(n8622));
  jnot g08431(.din(n8622), .dout(n8623));
  jand g08432(.dina(n8623), .dinb(n8419), .dout(n8624));
  jxor g08433(.dina(n8624), .dinb(n8621), .dout(n8625));
  jand g08434(.dina(n8558), .dinb(n8196), .dout(n8626));
  jand g08435(.dina(n8559), .dinb(n8557), .dout(n8627));
  jor  g08436(.dina(n8627), .dinb(n8626), .dout(n8628));
  jand g08437(.dina(n8536), .dinb(n8533), .dout(n8629));
  jnot g08438(.din(n8629), .dout(n8630));
  jand g08439(.dina(n8630), .dinb(n8539), .dout(n8631));
  jor  g08440(.dina(n8523), .dinb(n8522), .dout(n8632));
  jand g08441(.dina(n8632), .dinb(n8527), .dout(n8633));
  jxor g08442(.dina(n8633), .dinb(n8631), .dout(n8634));
  jxor g08443(.dina(n8634), .dinb(n8628), .dout(n8635));
  jand g08444(.dina(n8560), .dinb(n8556), .dout(n8636));
  jand g08445(.dina(n8565), .dinb(n8561), .dout(n8637));
  jor  g08446(.dina(n8637), .dinb(n8636), .dout(n8638));
  jxor g08447(.dina(n8638), .dinb(n8635), .dout(n8639));
  jxor g08448(.dina(n8639), .dinb(n8625), .dout(n8640));
  jxor g08449(.dina(n8640), .dinb(n8617), .dout(n8641));
  jxor g08450(.dina(n8641), .dinb(n8592), .dout(n8642));
  jand g08451(.dina(n8449), .dinb(n8446), .dout(n8643));
  jand g08452(.dina(n8450), .dinb(n8425), .dout(n8644));
  jor  g08453(.dina(n8644), .dinb(n8643), .dout(n8645));
  jxor g08454(.dina(n8489), .dinb(n8406), .dout(n8646));
  jand g08455(.dina(n8499), .dinb(n8497), .dout(n8647));
  jnot g08456(.din(n8647), .dout(n8648));
  jand g08457(.dina(n8648), .dinb(n8502), .dout(n8649));
  jxor g08458(.dina(n8649), .dinb(n8646), .dout(n8650));
  jnot g08459(.din(n8650), .dout(n8651));
  jand g08460(.dina(n8529), .dinb(n8521), .dout(n8652));
  jnot g08461(.din(n8652), .dout(n8653));
  jor  g08462(.dina(n8541), .dinb(n8531), .dout(n8654));
  jand g08463(.dina(n8654), .dinb(n8653), .dout(n8655));
  jxor g08464(.dina(n8655), .dinb(n8651), .dout(n8656));
  jnot g08465(.din(n8656), .dout(n8657));
  jand g08466(.dina(n8505), .dinb(n8495), .dout(n8658));
  jnot g08467(.din(n8658), .dout(n8659));
  jor  g08468(.dina(n8517), .dinb(n8507), .dout(n8660));
  jand g08469(.dina(n8660), .dinb(n8659), .dout(n8661));
  jxor g08470(.dina(n8661), .dinb(n8657), .dout(n8662));
  jand g08471(.dina(n8566), .dinb(n8542), .dout(n8663));
  jand g08472(.dina(n8567), .dinb(n8518), .dout(n8664));
  jor  g08473(.dina(n8664), .dinb(n8663), .dout(n8665));
  jand g08474(.dina(n8385), .dinb(n8382), .dout(n8666));
  jand g08475(.dina(n8424), .dinb(n8386), .dout(n8667));
  jor  g08476(.dina(n8667), .dinb(n8666), .dout(n8668));
  jxor g08477(.dina(n8668), .dinb(n8665), .dout(n8669));
  jxor g08478(.dina(n8669), .dinb(n8662), .dout(n8670));
  jxor g08479(.dina(n8670), .dinb(n8645), .dout(n8671));
  jxor g08480(.dina(n8671), .dinb(n8642), .dout(n8672));
  jxor g08481(.dina(n8672), .dinb(n8589), .dout(n8673));
  jand g08482(.dina(n8373), .dinb(n8342), .dout(n8674));
  jand g08483(.dina(n8374), .dinb(n8337), .dout(n8675));
  jor  g08484(.dina(n8675), .dinb(n8674), .dout(n8676));
  jand g08485(.dina(n8568), .dinb(n8478), .dout(n8677));
  jand g08486(.dina(n8569), .dinb(n8473), .dout(n8678));
  jor  g08487(.dina(n8678), .dinb(n8677), .dout(n8679));
  jxor g08488(.dina(n8679), .dinb(n8676), .dout(n8680));
  jand g08489(.dina(n8348), .dinb(n8345), .dout(n8681));
  jand g08490(.dina(n8372), .dinb(n8349), .dout(n8682));
  jor  g08491(.dina(n8682), .dinb(n8681), .dout(n8683));
  jand g08492(.dina(\a[55] ), .dinb(\a[11] ), .dout(n8684));
  jand g08493(.dina(\a[54] ), .dinb(\a[12] ), .dout(n8685));
  jand g08494(.dina(\a[47] ), .dinb(\a[19] ), .dout(n8686));
  jand g08495(.dina(n8686), .dinb(n8685), .dout(n8687));
  jnot g08496(.din(n8687), .dout(n8688));
  jand g08497(.dina(\a[55] ), .dinb(\a[12] ), .dout(n8689));
  jand g08498(.dina(n8689), .dinb(n8558), .dout(n8690));
  jand g08499(.dina(n8686), .dinb(n8684), .dout(n8691));
  jor  g08500(.dina(n8691), .dinb(n8690), .dout(n8692));
  jand g08501(.dina(n8692), .dinb(n8688), .dout(n8693));
  jnot g08502(.din(n8693), .dout(n8694));
  jand g08503(.dina(n8694), .dinb(n8684), .dout(n8695));
  jor  g08504(.dina(n8692), .dinb(n8687), .dout(n8696));
  jnot g08505(.din(n8696), .dout(n8697));
  jor  g08506(.dina(n8686), .dinb(n8685), .dout(n8698));
  jand g08507(.dina(n8698), .dinb(n8697), .dout(n8699));
  jor  g08508(.dina(n8699), .dinb(n8695), .dout(n8700));
  jand g08509(.dina(\a[63] ), .dinb(\a[3] ), .dout(n8701));
  jand g08510(.dina(\a[62] ), .dinb(\a[61] ), .dout(n8702));
  jand g08511(.dina(n8702), .dinb(n242), .dout(n8703));
  jnot g08512(.din(n8703), .dout(n8704));
  jand g08513(.dina(\a[61] ), .dinb(\a[5] ), .dout(n8705));
  jand g08514(.dina(\a[62] ), .dinb(\a[4] ), .dout(n8706));
  jor  g08515(.dina(n8706), .dinb(n8705), .dout(n8707));
  jand g08516(.dina(n8707), .dinb(n8704), .dout(n8708));
  jxor g08517(.dina(n8708), .dinb(n8701), .dout(n8709));
  jnot g08518(.din(n8709), .dout(n8710));
  jand g08519(.dina(\a[39] ), .dinb(\a[27] ), .dout(n8711));
  jnot g08520(.din(n8711), .dout(n8712));
  jand g08521(.dina(\a[38] ), .dinb(\a[29] ), .dout(n8713));
  jand g08522(.dina(n8713), .dinb(n8514), .dout(n8714));
  jnot g08523(.din(n8714), .dout(n8715));
  jand g08524(.dina(\a[37] ), .dinb(\a[29] ), .dout(n8716));
  jor  g08525(.dina(n8716), .dinb(n8510), .dout(n8717));
  jand g08526(.dina(n8717), .dinb(n8715), .dout(n8718));
  jxor g08527(.dina(n8718), .dinb(n8712), .dout(n8719));
  jxor g08528(.dina(n8719), .dinb(n8710), .dout(n8720));
  jxor g08529(.dina(n8720), .dinb(n8700), .dout(n8721));
  jand g08530(.dina(\a[43] ), .dinb(\a[23] ), .dout(n8722));
  jand g08531(.dina(\a[57] ), .dinb(\a[9] ), .dout(n8723));
  jand g08532(.dina(\a[42] ), .dinb(\a[24] ), .dout(n8724));
  jxor g08533(.dina(n8724), .dinb(n8723), .dout(n8725));
  jxor g08534(.dina(n8725), .dinb(n8722), .dout(n8726));
  jnot g08535(.din(n8726), .dout(n8727));
  jand g08536(.dina(\a[46] ), .dinb(\a[20] ), .dout(n8728));
  jnot g08537(.din(n8728), .dout(n8729));
  jand g08538(.dina(n4812), .dinb(n1376), .dout(n8730));
  jnot g08539(.din(n8730), .dout(n8731));
  jand g08540(.dina(\a[45] ), .dinb(\a[21] ), .dout(n8732));
  jand g08541(.dina(\a[44] ), .dinb(\a[22] ), .dout(n8733));
  jor  g08542(.dina(n8733), .dinb(n8732), .dout(n8734));
  jand g08543(.dina(n8734), .dinb(n8731), .dout(n8735));
  jxor g08544(.dina(n8735), .dinb(n8729), .dout(n8736));
  jxor g08545(.dina(n8736), .dinb(n8727), .dout(n8737));
  jnot g08546(.din(n8737), .dout(n8738));
  jnot g08547(.din(n8485), .dout(n8739));
  jand g08548(.dina(n4632), .dinb(n2128), .dout(n8740));
  jnot g08549(.din(n8740), .dout(n8741));
  jand g08550(.dina(\a[40] ), .dinb(\a[26] ), .dout(n8742));
  jand g08551(.dina(\a[41] ), .dinb(\a[25] ), .dout(n8743));
  jor  g08552(.dina(n8743), .dinb(n8742), .dout(n8744));
  jand g08553(.dina(n8744), .dinb(n8741), .dout(n8745));
  jxor g08554(.dina(n8745), .dinb(n8739), .dout(n8746));
  jxor g08555(.dina(n8746), .dinb(n8738), .dout(n8747));
  jand g08556(.dina(\a[48] ), .dinb(\a[18] ), .dout(n8748));
  jand g08557(.dina(\a[53] ), .dinb(\a[13] ), .dout(n8749));
  jand g08558(.dina(\a[51] ), .dinb(\a[15] ), .dout(n8750));
  jor  g08559(.dina(n8750), .dinb(n8749), .dout(n8751));
  jand g08560(.dina(n6130), .dinb(n727), .dout(n8752));
  jnot g08561(.din(n8752), .dout(n8753));
  jand g08562(.dina(n8753), .dinb(n8751), .dout(n8754));
  jxor g08563(.dina(n8754), .dinb(n8748), .dout(n8755));
  jnot g08564(.din(n8755), .dout(n8756));
  jand g08565(.dina(\a[52] ), .dinb(\a[14] ), .dout(n8757));
  jnot g08566(.din(n8757), .dout(n8758));
  jand g08567(.dina(n3243), .dinb(n2440), .dout(n8759));
  jnot g08568(.din(n8759), .dout(n8760));
  jand g08569(.dina(\a[35] ), .dinb(\a[31] ), .dout(n8761));
  jand g08570(.dina(\a[36] ), .dinb(\a[30] ), .dout(n8762));
  jor  g08571(.dina(n8762), .dinb(n8761), .dout(n8763));
  jand g08572(.dina(n8763), .dinb(n8760), .dout(n8764));
  jxor g08573(.dina(n8764), .dinb(n8758), .dout(n8765));
  jxor g08574(.dina(n8765), .dinb(n8756), .dout(n8766));
  jnot g08575(.din(n8766), .dout(n8767));
  jnot g08576(.din(n3492), .dout(n8768));
  jand g08577(.dina(\a[50] ), .dinb(\a[17] ), .dout(n8769));
  jand g08578(.dina(n8769), .dinb(n8413), .dout(n8770));
  jnot g08579(.din(n8770), .dout(n8771));
  jand g08580(.dina(\a[49] ), .dinb(\a[17] ), .dout(n8772));
  jand g08581(.dina(\a[50] ), .dinb(\a[16] ), .dout(n8773));
  jor  g08582(.dina(n8773), .dinb(n8772), .dout(n8774));
  jand g08583(.dina(n8774), .dinb(n8771), .dout(n8775));
  jxor g08584(.dina(n8775), .dinb(n8768), .dout(n8776));
  jxor g08585(.dina(n8776), .dinb(n8767), .dout(n8777));
  jxor g08586(.dina(n8777), .dinb(n8747), .dout(n8778));
  jxor g08587(.dina(n8778), .dinb(n8721), .dout(n8779));
  jxor g08588(.dina(n8779), .dinb(n8683), .dout(n8780));
  jand g08589(.dina(n8360), .dinb(n8357), .dout(n8781));
  jand g08590(.dina(n8361), .dinb(n8165), .dout(n8782));
  jor  g08591(.dina(n8782), .dinb(n8781), .dout(n8783));
  jand g08592(.dina(n8368), .dinb(n8366), .dout(n8784));
  jand g08593(.dina(n8369), .dinb(n8364), .dout(n8785));
  jor  g08594(.dina(n8785), .dinb(n8784), .dout(n8786));
  jxor g08595(.dina(n8786), .dinb(n8783), .dout(n8787));
  jand g08596(.dina(n8431), .dinb(n8428), .dout(n8788));
  jand g08597(.dina(n8435), .dinb(n8432), .dout(n8789));
  jor  g08598(.dina(n8789), .dinb(n8788), .dout(n8790));
  jxor g08599(.dina(n8790), .dinb(n8787), .dout(n8791));
  jand g08600(.dina(n8370), .dinb(n8362), .dout(n8792));
  jand g08601(.dina(n8371), .dinb(n8354), .dout(n8793));
  jor  g08602(.dina(n8793), .dinb(n8792), .dout(n8794));
  jnot g08603(.din(n8794), .dout(n8795));
  jor  g08604(.dina(n8440), .dinb(n8437), .dout(n8796));
  jor  g08605(.dina(n8445), .dinb(n8442), .dout(n8797));
  jand g08606(.dina(n8797), .dinb(n8796), .dout(n8798));
  jxor g08607(.dina(n8798), .dinb(n8795), .dout(n8799));
  jxor g08608(.dina(n8799), .dinb(n8791), .dout(n8800));
  jxor g08609(.dina(n8800), .dinb(n8780), .dout(n8801));
  jxor g08610(.dina(n8801), .dinb(n8680), .dout(n8802));
  jxor g08611(.dina(n8802), .dinb(n8673), .dout(n8803));
  jand g08612(.dina(n8803), .dinb(n8586), .dout(n8804));
  jor  g08613(.dina(n8803), .dinb(n8586), .dout(n8805));
  jnot g08614(.din(n8805), .dout(n8806));
  jor  g08615(.dina(n8806), .dinb(n8804), .dout(n8807));
  jnot g08616(.din(n8573), .dout(n8808));
  jor  g08617(.dina(n8582), .dinb(n8575), .dout(n8809));
  jand g08618(.dina(n8809), .dinb(n8808), .dout(n8810));
  jxor g08619(.dina(n8810), .dinb(n8807), .dout(\asquared[67] ));
  jand g08620(.dina(n8672), .dinb(n8589), .dout(n8812));
  jand g08621(.dina(n8802), .dinb(n8673), .dout(n8813));
  jor  g08622(.dina(n8813), .dinb(n8812), .dout(n8814));
  jand g08623(.dina(n8679), .dinb(n8676), .dout(n8815));
  jand g08624(.dina(n8801), .dinb(n8680), .dout(n8816));
  jor  g08625(.dina(n8816), .dinb(n8815), .dout(n8817));
  jand g08626(.dina(n8640), .dinb(n8617), .dout(n8818));
  jand g08627(.dina(n8641), .dinb(n8592), .dout(n8819));
  jor  g08628(.dina(n8819), .dinb(n8818), .dout(n8820));
  jor  g08629(.dina(n8798), .dinb(n8795), .dout(n8821));
  jand g08630(.dina(n8799), .dinb(n8791), .dout(n8822));
  jnot g08631(.din(n8822), .dout(n8823));
  jand g08632(.dina(n8823), .dinb(n8821), .dout(n8824));
  jnot g08633(.din(n8824), .dout(n8825));
  jor  g08634(.dina(n8736), .dinb(n8727), .dout(n8826));
  jor  g08635(.dina(n8746), .dinb(n8738), .dout(n8827));
  jand g08636(.dina(n8827), .dinb(n8826), .dout(n8828));
  jand g08637(.dina(n8603), .dinb(n8600), .dout(n8829));
  jnot g08638(.din(n8829), .dout(n8830));
  jor  g08639(.dina(n8614), .dinb(n8605), .dout(n8831));
  jand g08640(.dina(n8831), .dinb(n8830), .dout(n8832));
  jxor g08641(.dina(n8832), .dinb(n8828), .dout(n8833));
  jnot g08642(.din(n8833), .dout(n8834));
  jor  g08643(.dina(n8719), .dinb(n8710), .dout(n8835));
  jand g08644(.dina(n8720), .dinb(n8700), .dout(n8836));
  jnot g08645(.din(n8836), .dout(n8837));
  jand g08646(.dina(n8837), .dinb(n8835), .dout(n8838));
  jxor g08647(.dina(n8838), .dinb(n8834), .dout(n8839));
  jand g08648(.dina(n8708), .dinb(n8701), .dout(n8840));
  jor  g08649(.dina(n8840), .dinb(n8703), .dout(n8841));
  jand g08650(.dina(n8610), .dinb(n8607), .dout(n8842));
  jnot g08651(.din(n8842), .dout(n8843));
  jand g08652(.dina(n8843), .dinb(n8612), .dout(n8844));
  jxor g08653(.dina(n8844), .dinb(n8841), .dout(n8845));
  jand g08654(.dina(n8715), .dinb(n8712), .dout(n8846));
  jnot g08655(.din(n8846), .dout(n8847));
  jand g08656(.dina(n8847), .dinb(n8717), .dout(n8848));
  jxor g08657(.dina(n8848), .dinb(n8845), .dout(n8849));
  jand g08658(.dina(n8724), .dinb(n8723), .dout(n8850));
  jand g08659(.dina(n8725), .dinb(n8722), .dout(n8851));
  jor  g08660(.dina(n8851), .dinb(n8850), .dout(n8852));
  jand g08661(.dina(n8741), .dinb(n8739), .dout(n8853));
  jnot g08662(.din(n8853), .dout(n8854));
  jand g08663(.dina(n8854), .dinb(n8744), .dout(n8855));
  jxor g08664(.dina(n8855), .dinb(n8852), .dout(n8856));
  jand g08665(.dina(n8731), .dinb(n8729), .dout(n8857));
  jnot g08666(.din(n8857), .dout(n8858));
  jand g08667(.dina(n8858), .dinb(n8734), .dout(n8859));
  jxor g08668(.dina(n8859), .dinb(n8856), .dout(n8860));
  jand g08669(.dina(\a[61] ), .dinb(\a[6] ), .dout(n8861));
  jand g08670(.dina(n8771), .dinb(n8768), .dout(n8862));
  jnot g08671(.din(n8862), .dout(n8863));
  jand g08672(.dina(n8863), .dinb(n8774), .dout(n8864));
  jxor g08673(.dina(n8864), .dinb(n8861), .dout(n8865));
  jand g08674(.dina(n8760), .dinb(n8758), .dout(n8866));
  jnot g08675(.din(n8866), .dout(n8867));
  jand g08676(.dina(n8867), .dinb(n8763), .dout(n8868));
  jxor g08677(.dina(n8868), .dinb(n8865), .dout(n8869));
  jxor g08678(.dina(n8869), .dinb(n8860), .dout(n8870));
  jxor g08679(.dina(n8870), .dinb(n8849), .dout(n8871));
  jxor g08680(.dina(n8871), .dinb(n8839), .dout(n8872));
  jxor g08681(.dina(n8872), .dinb(n8825), .dout(n8873));
  jxor g08682(.dina(n8873), .dinb(n8820), .dout(n8874));
  jor  g08683(.dina(n8765), .dinb(n8756), .dout(n8875));
  jor  g08684(.dina(n8776), .dinb(n8767), .dout(n8876));
  jand g08685(.dina(n8876), .dinb(n8875), .dout(n8877));
  jnot g08686(.din(n8877), .dout(n8878));
  jand g08687(.dina(n8754), .dinb(n8748), .dout(n8879));
  jor  g08688(.dina(n8879), .dinb(n8752), .dout(n8880));
  jxor g08689(.dina(n8880), .dinb(n8696), .dout(n8881));
  jand g08690(.dina(\a[57] ), .dinb(\a[10] ), .dout(n8882));
  jand g08691(.dina(\a[56] ), .dinb(\a[11] ), .dout(n8883));
  jand g08692(.dina(\a[47] ), .dinb(\a[20] ), .dout(n8884));
  jand g08693(.dina(n8884), .dinb(n8883), .dout(n8885));
  jnot g08694(.din(n8885), .dout(n8886));
  jand g08695(.dina(\a[57] ), .dinb(\a[11] ), .dout(n8887));
  jand g08696(.dina(n8887), .dinb(n8485), .dout(n8888));
  jand g08697(.dina(n8884), .dinb(n8882), .dout(n8889));
  jor  g08698(.dina(n8889), .dinb(n8888), .dout(n8890));
  jand g08699(.dina(n8890), .dinb(n8886), .dout(n8891));
  jnot g08700(.din(n8891), .dout(n8892));
  jand g08701(.dina(n8892), .dinb(n8882), .dout(n8893));
  jor  g08702(.dina(n8890), .dinb(n8885), .dout(n8894));
  jnot g08703(.din(n8894), .dout(n8895));
  jor  g08704(.dina(n8884), .dinb(n8883), .dout(n8896));
  jand g08705(.dina(n8896), .dinb(n8895), .dout(n8897));
  jor  g08706(.dina(n8897), .dinb(n8893), .dout(n8898));
  jxor g08707(.dina(n8898), .dinb(n8881), .dout(n8899));
  jxor g08708(.dina(n8899), .dinb(n8878), .dout(n8900));
  jand g08709(.dina(n8786), .dinb(n8783), .dout(n8901));
  jand g08710(.dina(n8790), .dinb(n8787), .dout(n8902));
  jor  g08711(.dina(n8902), .dinb(n8901), .dout(n8903));
  jxor g08712(.dina(n8903), .dinb(n8900), .dout(n8904));
  jand g08713(.dina(n8777), .dinb(n8747), .dout(n8905));
  jand g08714(.dina(n8778), .dinb(n8721), .dout(n8906));
  jor  g08715(.dina(n8906), .dinb(n8905), .dout(n8907));
  jand g08716(.dina(n8615), .dinb(n8598), .dout(n8908));
  jand g08717(.dina(n8616), .dinb(n8595), .dout(n8909));
  jor  g08718(.dina(n8909), .dinb(n8908), .dout(n8910));
  jxor g08719(.dina(n8910), .dinb(n8907), .dout(n8911));
  jxor g08720(.dina(n8911), .dinb(n8904), .dout(n8912));
  jxor g08721(.dina(n8912), .dinb(n8874), .dout(n8913));
  jxor g08722(.dina(n8913), .dinb(n8817), .dout(n8914));
  jand g08723(.dina(n8670), .dinb(n8645), .dout(n8915));
  jand g08724(.dina(n8671), .dinb(n8642), .dout(n8916));
  jor  g08725(.dina(n8916), .dinb(n8915), .dout(n8917));
  jand g08726(.dina(n8779), .dinb(n8683), .dout(n8918));
  jand g08727(.dina(n8800), .dinb(n8780), .dout(n8919));
  jor  g08728(.dina(n8919), .dinb(n8918), .dout(n8920));
  jxor g08729(.dina(n8920), .dinb(n8917), .dout(n8921));
  jand g08730(.dina(n8668), .dinb(n8665), .dout(n8922));
  jand g08731(.dina(n8669), .dinb(n8662), .dout(n8923));
  jor  g08732(.dina(n8923), .dinb(n8922), .dout(n8924));
  jand g08733(.dina(\a[42] ), .dinb(\a[25] ), .dout(n8925));
  jand g08734(.dina(n4514), .dinb(n2128), .dout(n8926));
  jand g08735(.dina(\a[46] ), .dinb(\a[21] ), .dout(n8927));
  jand g08736(.dina(n8927), .dinb(n8925), .dout(n8928));
  jor  g08737(.dina(n8928), .dinb(n8926), .dout(n8929));
  jand g08738(.dina(\a[41] ), .dinb(\a[26] ), .dout(n8930));
  jand g08739(.dina(n8930), .dinb(n8927), .dout(n8931));
  jnot g08740(.din(n8931), .dout(n8932));
  jand g08741(.dina(n8932), .dinb(n8929), .dout(n8933));
  jnot g08742(.din(n8933), .dout(n8934));
  jand g08743(.dina(n8934), .dinb(n8925), .dout(n8935));
  jor  g08744(.dina(n8931), .dinb(n8929), .dout(n8936));
  jnot g08745(.din(n8936), .dout(n8937));
  jor  g08746(.dina(n8930), .dinb(n8927), .dout(n8938));
  jand g08747(.dina(n8938), .dinb(n8937), .dout(n8939));
  jor  g08748(.dina(n8939), .dinb(n8935), .dout(n8940));
  jand g08749(.dina(\a[48] ), .dinb(\a[19] ), .dout(n8941));
  jand g08750(.dina(\a[53] ), .dinb(\a[14] ), .dout(n8942));
  jxor g08751(.dina(n8942), .dinb(n8769), .dout(n8943));
  jxor g08752(.dina(n8943), .dinb(n8941), .dout(n8944));
  jxor g08753(.dina(n8944), .dinb(n8940), .dout(n8945));
  jnot g08754(.din(n8945), .dout(n8946));
  jand g08755(.dina(\a[63] ), .dinb(\a[4] ), .dout(n8947));
  jnot g08756(.din(n8947), .dout(n8948));
  jand g08757(.dina(n3665), .dinb(n2042), .dout(n8949));
  jnot g08758(.din(n8949), .dout(n8950));
  jand g08759(.dina(\a[40] ), .dinb(\a[27] ), .dout(n8951));
  jand g08760(.dina(\a[39] ), .dinb(\a[28] ), .dout(n8952));
  jor  g08761(.dina(n8952), .dinb(n8951), .dout(n8953));
  jand g08762(.dina(n8953), .dinb(n8950), .dout(n8954));
  jxor g08763(.dina(n8954), .dinb(n8948), .dout(n8955));
  jxor g08764(.dina(n8955), .dinb(n8946), .dout(n8956));
  jand g08765(.dina(\a[36] ), .dinb(\a[31] ), .dout(n8957));
  jand g08766(.dina(n2845), .dinb(n2671), .dout(n8958));
  jnot g08767(.din(n8958), .dout(n8959));
  jand g08768(.dina(n8957), .dinb(n3634), .dout(n8960));
  jand g08769(.dina(n3269), .dinb(n3243), .dout(n8961));
  jor  g08770(.dina(n8961), .dinb(n8960), .dout(n8962));
  jand g08771(.dina(n8962), .dinb(n8959), .dout(n8963));
  jnot g08772(.din(n8963), .dout(n8964));
  jand g08773(.dina(n8964), .dinb(n8957), .dout(n8965));
  jor  g08774(.dina(n8962), .dinb(n8958), .dout(n8966));
  jnot g08775(.din(n8966), .dout(n8967));
  jand g08776(.dina(\a[35] ), .dinb(\a[32] ), .dout(n8968));
  jor  g08777(.dina(n8968), .dinb(n3634), .dout(n8969));
  jand g08778(.dina(n8969), .dinb(n8967), .dout(n8970));
  jor  g08779(.dina(n8970), .dinb(n8965), .dout(n8971));
  jand g08780(.dina(\a[49] ), .dinb(\a[18] ), .dout(n8972));
  jnot g08781(.din(\a[34] ), .dout(n8973));
  jand g08782(.dina(\a[62] ), .dinb(\a[5] ), .dout(n8974));
  jnot g08783(.din(n8974), .dout(n8975));
  jand g08784(.dina(n8975), .dinb(n8973), .dout(n8976));
  jand g08785(.dina(n3186), .dinb(\a[62] ), .dout(n8977));
  jor  g08786(.dina(n8977), .dinb(n8976), .dout(n8978));
  jnot g08787(.din(n8978), .dout(n8979));
  jxor g08788(.dina(n8979), .dinb(n8972), .dout(n8980));
  jxor g08789(.dina(n8980), .dinb(n8971), .dout(n8981));
  jnot g08790(.din(n8981), .dout(n8982));
  jnot g08791(.din(n8713), .dout(n8983));
  jand g08792(.dina(\a[55] ), .dinb(\a[13] ), .dout(n8984));
  jand g08793(.dina(n8984), .dinb(n8685), .dout(n8985));
  jnot g08794(.din(n8985), .dout(n8986));
  jand g08795(.dina(\a[54] ), .dinb(\a[13] ), .dout(n8987));
  jor  g08796(.dina(n8987), .dinb(n8689), .dout(n8988));
  jand g08797(.dina(n8988), .dinb(n8986), .dout(n8989));
  jxor g08798(.dina(n8989), .dinb(n8983), .dout(n8990));
  jxor g08799(.dina(n8990), .dinb(n8982), .dout(n8991));
  jand g08800(.dina(\a[60] ), .dinb(\a[7] ), .dout(n8992));
  jand g08801(.dina(\a[58] ), .dinb(\a[9] ), .dout(n8993));
  jor  g08802(.dina(n8993), .dinb(n8608), .dout(n8994));
  jand g08803(.dina(\a[59] ), .dinb(\a[9] ), .dout(n8995));
  jand g08804(.dina(n8995), .dinb(n8611), .dout(n8996));
  jnot g08805(.din(n8996), .dout(n8997));
  jand g08806(.dina(n8997), .dinb(n8994), .dout(n8998));
  jxor g08807(.dina(n8998), .dinb(n8992), .dout(n8999));
  jnot g08808(.din(n8999), .dout(n9000));
  jand g08809(.dina(\a[45] ), .dinb(\a[22] ), .dout(n9001));
  jnot g08810(.din(n9001), .dout(n9002));
  jand g08811(.dina(n4495), .dinb(n1942), .dout(n9003));
  jnot g08812(.din(n9003), .dout(n9004));
  jand g08813(.dina(\a[44] ), .dinb(\a[23] ), .dout(n9005));
  jand g08814(.dina(\a[43] ), .dinb(\a[24] ), .dout(n9006));
  jor  g08815(.dina(n9006), .dinb(n9005), .dout(n9007));
  jand g08816(.dina(n9007), .dinb(n9004), .dout(n9008));
  jxor g08817(.dina(n9008), .dinb(n9002), .dout(n9009));
  jxor g08818(.dina(n9009), .dinb(n9000), .dout(n9010));
  jand g08819(.dina(\a[52] ), .dinb(\a[15] ), .dout(n9011));
  jand g08820(.dina(\a[37] ), .dinb(\a[30] ), .dout(n9012));
  jand g08821(.dina(\a[51] ), .dinb(\a[16] ), .dout(n9013));
  jxor g08822(.dina(n9013), .dinb(n9012), .dout(n9014));
  jxor g08823(.dina(n9014), .dinb(n9011), .dout(n9015));
  jxor g08824(.dina(n9015), .dinb(n9010), .dout(n9016));
  jxor g08825(.dina(n9016), .dinb(n8991), .dout(n9017));
  jxor g08826(.dina(n9017), .dinb(n8956), .dout(n9018));
  jxor g08827(.dina(n9018), .dinb(n8924), .dout(n9019));
  jand g08828(.dina(n8633), .dinb(n8631), .dout(n9020));
  jand g08829(.dina(n8634), .dinb(n8628), .dout(n9021));
  jor  g08830(.dina(n9021), .dinb(n9020), .dout(n9022));
  jnot g08831(.din(n8406), .dout(n9023));
  jnot g08832(.din(n8489), .dout(n9024));
  jand g08833(.dina(n9024), .dinb(n9023), .dout(n9025));
  jand g08834(.dina(n8649), .dinb(n8646), .dout(n9026));
  jor  g08835(.dina(n9026), .dinb(n9025), .dout(n9027));
  jxor g08836(.dina(n9027), .dinb(n9022), .dout(n9028));
  jand g08837(.dina(n8620), .dinb(n8551), .dout(n9029));
  jand g08838(.dina(n8624), .dinb(n8621), .dout(n9030));
  jor  g08839(.dina(n9030), .dinb(n9029), .dout(n9031));
  jxor g08840(.dina(n9031), .dinb(n9028), .dout(n9032));
  jand g08841(.dina(n8638), .dinb(n8635), .dout(n9033));
  jand g08842(.dina(n8639), .dinb(n8625), .dout(n9034));
  jor  g08843(.dina(n9034), .dinb(n9033), .dout(n9035));
  jnot g08844(.din(n9035), .dout(n9036));
  jor  g08845(.dina(n8655), .dinb(n8651), .dout(n9037));
  jor  g08846(.dina(n8661), .dinb(n8657), .dout(n9038));
  jand g08847(.dina(n9038), .dinb(n9037), .dout(n9039));
  jxor g08848(.dina(n9039), .dinb(n9036), .dout(n9040));
  jxor g08849(.dina(n9040), .dinb(n9032), .dout(n9041));
  jxor g08850(.dina(n9041), .dinb(n9019), .dout(n9042));
  jxor g08851(.dina(n9042), .dinb(n8921), .dout(n9043));
  jxor g08852(.dina(n9043), .dinb(n8914), .dout(n9044));
  jand g08853(.dina(n9044), .dinb(n8814), .dout(n9045));
  jor  g08854(.dina(n9044), .dinb(n8814), .dout(n9046));
  jnot g08855(.din(n9046), .dout(n9047));
  jor  g08856(.dina(n9047), .dinb(n9045), .dout(n9048));
  jnot g08857(.din(n8804), .dout(n9049));
  jor  g08858(.dina(n8810), .dinb(n8806), .dout(n9050));
  jand g08859(.dina(n9050), .dinb(n9049), .dout(n9051));
  jxor g08860(.dina(n9051), .dinb(n9048), .dout(\asquared[68] ));
  jand g08861(.dina(n8913), .dinb(n8817), .dout(n9053));
  jand g08862(.dina(n9043), .dinb(n8914), .dout(n9054));
  jor  g08863(.dina(n9054), .dinb(n9053), .dout(n9055));
  jand g08864(.dina(n8873), .dinb(n8820), .dout(n9056));
  jand g08865(.dina(n8912), .dinb(n8874), .dout(n9057));
  jor  g08866(.dina(n9057), .dinb(n9056), .dout(n9058));
  jand g08867(.dina(n9018), .dinb(n8924), .dout(n9059));
  jand g08868(.dina(n9041), .dinb(n9019), .dout(n9060));
  jor  g08869(.dina(n9060), .dinb(n9059), .dout(n9061));
  jand g08870(.dina(n8910), .dinb(n8907), .dout(n9062));
  jand g08871(.dina(n8911), .dinb(n8904), .dout(n9063));
  jor  g08872(.dina(n9063), .dinb(n9062), .dout(n9064));
  jand g08873(.dina(n8869), .dinb(n8860), .dout(n9065));
  jand g08874(.dina(n8870), .dinb(n8849), .dout(n9066));
  jor  g08875(.dina(n9066), .dinb(n9065), .dout(n9067));
  jnot g08876(.din(n9067), .dout(n9068));
  jor  g08877(.dina(n8832), .dinb(n8828), .dout(n9069));
  jor  g08878(.dina(n8838), .dinb(n8834), .dout(n9070));
  jand g08879(.dina(n9070), .dinb(n9069), .dout(n9071));
  jxor g08880(.dina(n9071), .dinb(n9068), .dout(n9072));
  jand g08881(.dina(n8899), .dinb(n8878), .dout(n9073));
  jand g08882(.dina(n8903), .dinb(n8900), .dout(n9074));
  jor  g08883(.dina(n9074), .dinb(n9073), .dout(n9075));
  jxor g08884(.dina(n9075), .dinb(n9072), .dout(n9076));
  jand g08885(.dina(n7519), .dinb(n655), .dout(n9077));
  jnot g08886(.din(n9077), .dout(n9078));
  jand g08887(.dina(\a[58] ), .dinb(\a[10] ), .dout(n9079));
  jor  g08888(.dina(n9079), .dinb(n8887), .dout(n9080));
  jand g08889(.dina(n9080), .dinb(n9078), .dout(n9081));
  jxor g08890(.dina(n9081), .dinb(n8995), .dout(n9082));
  jnot g08891(.din(n9082), .dout(n9083));
  jand g08892(.dina(\a[41] ), .dinb(\a[27] ), .dout(n9084));
  jnot g08893(.din(n9084), .dout(n9085));
  jand g08894(.dina(n3665), .dinb(n2653), .dout(n9086));
  jnot g08895(.din(n9086), .dout(n9087));
  jand g08896(.dina(\a[40] ), .dinb(\a[28] ), .dout(n9088));
  jand g08897(.dina(\a[39] ), .dinb(\a[29] ), .dout(n9089));
  jor  g08898(.dina(n9089), .dinb(n9088), .dout(n9090));
  jand g08899(.dina(n9090), .dinb(n9087), .dout(n9091));
  jxor g08900(.dina(n9091), .dinb(n9085), .dout(n9092));
  jxor g08901(.dina(n9092), .dinb(n9083), .dout(n9093));
  jand g08902(.dina(\a[47] ), .dinb(\a[21] ), .dout(n9094));
  jand g08903(.dina(\a[63] ), .dinb(\a[6] ), .dout(n9095));
  jand g08904(.dina(n9095), .dinb(n8974), .dout(n9096));
  jnot g08905(.din(n9096), .dout(n9097));
  jand g08906(.dina(\a[63] ), .dinb(\a[5] ), .dout(n9098));
  jand g08907(.dina(\a[62] ), .dinb(\a[6] ), .dout(n9099));
  jor  g08908(.dina(n9099), .dinb(n9098), .dout(n9100));
  jand g08909(.dina(n9100), .dinb(n9097), .dout(n9101));
  jxor g08910(.dina(n9101), .dinb(n9094), .dout(n9102));
  jxor g08911(.dina(n9102), .dinb(n9093), .dout(n9103));
  jand g08912(.dina(\a[56] ), .dinb(\a[12] ), .dout(n9104));
  jnot g08913(.din(n9104), .dout(n9105));
  jand g08914(.dina(\a[51] ), .dinb(\a[17] ), .dout(n9106));
  jand g08915(.dina(n9106), .dinb(n9104), .dout(n9107));
  jand g08916(.dina(\a[56] ), .dinb(\a[13] ), .dout(n9108));
  jand g08917(.dina(n9108), .dinb(n8689), .dout(n9109));
  jor  g08918(.dina(n9109), .dinb(n9107), .dout(n9110));
  jand g08919(.dina(n9106), .dinb(n8984), .dout(n9111));
  jnot g08920(.din(n9111), .dout(n9112));
  jand g08921(.dina(n9112), .dinb(n9110), .dout(n9113));
  jor  g08922(.dina(n9113), .dinb(n9105), .dout(n9114));
  jor  g08923(.dina(n9111), .dinb(n9110), .dout(n9115));
  jnot g08924(.din(n9115), .dout(n9116));
  jor  g08925(.dina(n9106), .dinb(n8984), .dout(n9117));
  jand g08926(.dina(n9117), .dinb(n9116), .dout(n9118));
  jnot g08927(.din(n9118), .dout(n9119));
  jand g08928(.dina(n9119), .dinb(n9114), .dout(n9120));
  jand g08929(.dina(\a[50] ), .dinb(\a[18] ), .dout(n9121));
  jand g08930(.dina(\a[49] ), .dinb(\a[19] ), .dout(n9122));
  jor  g08931(.dina(n9122), .dinb(n9121), .dout(n9123));
  jand g08932(.dina(\a[50] ), .dinb(\a[19] ), .dout(n9124));
  jand g08933(.dina(n9124), .dinb(n8972), .dout(n9125));
  jnot g08934(.din(n9125), .dout(n9126));
  jand g08935(.dina(n9126), .dinb(n9123), .dout(n9127));
  jxor g08936(.dina(n9127), .dinb(n3752), .dout(n9128));
  jnot g08937(.din(n9128), .dout(n9129));
  jand g08938(.dina(\a[38] ), .dinb(\a[30] ), .dout(n9130));
  jnot g08939(.din(n9130), .dout(n9131));
  jand g08940(.dina(n3269), .dinb(n3138), .dout(n9132));
  jnot g08941(.din(n9132), .dout(n9133));
  jand g08942(.dina(\a[37] ), .dinb(\a[31] ), .dout(n9134));
  jand g08943(.dina(\a[36] ), .dinb(\a[32] ), .dout(n9135));
  jor  g08944(.dina(n9135), .dinb(n9134), .dout(n9136));
  jand g08945(.dina(n9136), .dinb(n9133), .dout(n9137));
  jxor g08946(.dina(n9137), .dinb(n9131), .dout(n9138));
  jxor g08947(.dina(n9138), .dinb(n9129), .dout(n9139));
  jnot g08948(.din(n9139), .dout(n9140));
  jxor g08949(.dina(n9140), .dinb(n9120), .dout(n9141));
  jand g08950(.dina(\a[54] ), .dinb(\a[14] ), .dout(n9142));
  jand g08951(.dina(\a[53] ), .dinb(\a[15] ), .dout(n9143));
  jand g08952(.dina(\a[52] ), .dinb(\a[16] ), .dout(n9144));
  jor  g08953(.dina(n9144), .dinb(n9143), .dout(n9145));
  jand g08954(.dina(n7165), .dinb(n829), .dout(n9146));
  jnot g08955(.din(n9146), .dout(n9147));
  jand g08956(.dina(n9147), .dinb(n9145), .dout(n9148));
  jxor g08957(.dina(n9148), .dinb(n9142), .dout(n9149));
  jnot g08958(.din(n9149), .dout(n9150));
  jand g08959(.dina(\a[48] ), .dinb(\a[20] ), .dout(n9151));
  jnot g08960(.din(n9151), .dout(n9152));
  jand g08961(.dina(\a[46] ), .dinb(\a[23] ), .dout(n9153));
  jand g08962(.dina(n9153), .dinb(n9001), .dout(n9154));
  jnot g08963(.din(n9154), .dout(n9155));
  jand g08964(.dina(\a[45] ), .dinb(\a[23] ), .dout(n9156));
  jand g08965(.dina(\a[46] ), .dinb(\a[22] ), .dout(n9157));
  jor  g08966(.dina(n9157), .dinb(n9156), .dout(n9158));
  jand g08967(.dina(n9158), .dinb(n9155), .dout(n9159));
  jxor g08968(.dina(n9159), .dinb(n9152), .dout(n9160));
  jxor g08969(.dina(n9160), .dinb(n9150), .dout(n9161));
  jnot g08970(.din(n9161), .dout(n9162));
  jand g08971(.dina(\a[44] ), .dinb(\a[24] ), .dout(n9163));
  jnot g08972(.din(n9163), .dout(n9164));
  jand g08973(.dina(n4317), .dinb(n2128), .dout(n9165));
  jnot g08974(.din(n9165), .dout(n9166));
  jand g08975(.dina(\a[43] ), .dinb(\a[25] ), .dout(n9167));
  jand g08976(.dina(\a[42] ), .dinb(\a[26] ), .dout(n9168));
  jor  g08977(.dina(n9168), .dinb(n9167), .dout(n9169));
  jand g08978(.dina(n9169), .dinb(n9166), .dout(n9170));
  jxor g08979(.dina(n9170), .dinb(n9164), .dout(n9171));
  jxor g08980(.dina(n9171), .dinb(n9162), .dout(n9172));
  jxor g08981(.dina(n9172), .dinb(n9141), .dout(n9173));
  jxor g08982(.dina(n9173), .dinb(n9103), .dout(n9174));
  jxor g08983(.dina(n9174), .dinb(n9076), .dout(n9175));
  jxor g08984(.dina(n9175), .dinb(n9064), .dout(n9176));
  jxor g08985(.dina(n9176), .dinb(n9061), .dout(n9177));
  jxor g08986(.dina(n9177), .dinb(n9058), .dout(n9178));
  jand g08987(.dina(n8920), .dinb(n8917), .dout(n9179));
  jand g08988(.dina(n9042), .dinb(n8921), .dout(n9180));
  jor  g08989(.dina(n9180), .dinb(n9179), .dout(n9181));
  jor  g08990(.dina(n9039), .dinb(n9036), .dout(n9182));
  jand g08991(.dina(n9040), .dinb(n9032), .dout(n9183));
  jnot g08992(.din(n9183), .dout(n9184));
  jand g08993(.dina(n9184), .dinb(n9182), .dout(n9185));
  jnot g08994(.din(n9185), .dout(n9186));
  jand g08995(.dina(n8942), .dinb(n8769), .dout(n9187));
  jand g08996(.dina(n8943), .dinb(n8941), .dout(n9188));
  jor  g08997(.dina(n9188), .dinb(n9187), .dout(n9189));
  jxor g08998(.dina(n9189), .dinb(n8936), .dout(n9190));
  jand g08999(.dina(n8986), .dinb(n8983), .dout(n9191));
  jnot g09000(.din(n9191), .dout(n9192));
  jand g09001(.dina(n9192), .dinb(n8988), .dout(n9193));
  jxor g09002(.dina(n9193), .dinb(n9190), .dout(n9194));
  jand g09003(.dina(n8944), .dinb(n8940), .dout(n9195));
  jnot g09004(.din(n9195), .dout(n9196));
  jor  g09005(.dina(n8955), .dinb(n8946), .dout(n9197));
  jand g09006(.dina(n9197), .dinb(n9196), .dout(n9198));
  jand g09007(.dina(n8980), .dinb(n8971), .dout(n9199));
  jnot g09008(.din(n9199), .dout(n9200));
  jor  g09009(.dina(n8990), .dinb(n8982), .dout(n9201));
  jand g09010(.dina(n9201), .dinb(n9200), .dout(n9202));
  jxor g09011(.dina(n9202), .dinb(n9198), .dout(n9203));
  jxor g09012(.dina(n9203), .dinb(n9194), .dout(n9204));
  jand g09013(.dina(n9027), .dinb(n9022), .dout(n9205));
  jand g09014(.dina(n9031), .dinb(n9028), .dout(n9206));
  jor  g09015(.dina(n9206), .dinb(n9205), .dout(n9207));
  jand g09016(.dina(n8998), .dinb(n8992), .dout(n9208));
  jor  g09017(.dina(n9208), .dinb(n8996), .dout(n9209));
  jand g09018(.dina(n9004), .dinb(n9002), .dout(n9210));
  jnot g09019(.din(n9210), .dout(n9211));
  jand g09020(.dina(n9211), .dinb(n9007), .dout(n9212));
  jxor g09021(.dina(n9212), .dinb(n8894), .dout(n9213));
  jxor g09022(.dina(n9213), .dinb(n9209), .dout(n9214));
  jand g09023(.dina(n9013), .dinb(n9012), .dout(n9215));
  jand g09024(.dina(n9014), .dinb(n9011), .dout(n9216));
  jor  g09025(.dina(n9216), .dinb(n9215), .dout(n9217));
  jand g09026(.dina(n8950), .dinb(n8948), .dout(n9218));
  jnot g09027(.din(n9218), .dout(n9219));
  jand g09028(.dina(n9219), .dinb(n8953), .dout(n9220));
  jxor g09029(.dina(n9220), .dinb(n8966), .dout(n9221));
  jxor g09030(.dina(n9221), .dinb(n9217), .dout(n9222));
  jxor g09031(.dina(n9222), .dinb(n9214), .dout(n9223));
  jxor g09032(.dina(n9223), .dinb(n9207), .dout(n9224));
  jxor g09033(.dina(n9224), .dinb(n9204), .dout(n9225));
  jxor g09034(.dina(n9225), .dinb(n9186), .dout(n9226));
  jand g09035(.dina(n8871), .dinb(n8839), .dout(n9227));
  jand g09036(.dina(n8872), .dinb(n8825), .dout(n9228));
  jor  g09037(.dina(n9228), .dinb(n9227), .dout(n9229));
  jand g09038(.dina(n9016), .dinb(n8991), .dout(n9230));
  jand g09039(.dina(n9017), .dinb(n8956), .dout(n9231));
  jor  g09040(.dina(n9231), .dinb(n9230), .dout(n9232));
  jand g09041(.dina(n8880), .dinb(n8696), .dout(n9233));
  jand g09042(.dina(n8898), .dinb(n8881), .dout(n9234));
  jor  g09043(.dina(n9234), .dinb(n9233), .dout(n9235));
  jand g09044(.dina(n8855), .dinb(n8852), .dout(n9236));
  jand g09045(.dina(n8859), .dinb(n8856), .dout(n9237));
  jor  g09046(.dina(n9237), .dinb(n9236), .dout(n9238));
  jxor g09047(.dina(n9238), .dinb(n9235), .dout(n9239));
  jnot g09048(.din(n9239), .dout(n9240));
  jor  g09049(.dina(n9009), .dinb(n9000), .dout(n9241));
  jand g09050(.dina(n9015), .dinb(n9010), .dout(n9242));
  jnot g09051(.din(n9242), .dout(n9243));
  jand g09052(.dina(n9243), .dinb(n9241), .dout(n9244));
  jxor g09053(.dina(n9244), .dinb(n9240), .dout(n9245));
  jand g09054(.dina(n8864), .dinb(n8861), .dout(n9246));
  jand g09055(.dina(n8868), .dinb(n8865), .dout(n9247));
  jor  g09056(.dina(n9247), .dinb(n9246), .dout(n9248));
  jand g09057(.dina(n8979), .dinb(n8972), .dout(n9249));
  jor  g09058(.dina(n9249), .dinb(n8977), .dout(n9250));
  jand g09059(.dina(\a[61] ), .dinb(\a[8] ), .dout(n9251));
  jand g09060(.dina(n9251), .dinb(n8992), .dout(n9252));
  jnot g09061(.din(n9252), .dout(n9253));
  jand g09062(.dina(\a[61] ), .dinb(\a[7] ), .dout(n9254));
  jand g09063(.dina(\a[60] ), .dinb(\a[8] ), .dout(n9255));
  jor  g09064(.dina(n9255), .dinb(n9254), .dout(n9256));
  jand g09065(.dina(n9256), .dinb(n9253), .dout(n9257));
  jxor g09066(.dina(n9257), .dinb(n9250), .dout(n9258));
  jxor g09067(.dina(n9258), .dinb(n9248), .dout(n9259));
  jand g09068(.dina(n8844), .dinb(n8841), .dout(n9260));
  jand g09069(.dina(n8848), .dinb(n8845), .dout(n9261));
  jor  g09070(.dina(n9261), .dinb(n9260), .dout(n9262));
  jxor g09071(.dina(n9262), .dinb(n9259), .dout(n9263));
  jxor g09072(.dina(n9263), .dinb(n9245), .dout(n9264));
  jxor g09073(.dina(n9264), .dinb(n9232), .dout(n9265));
  jxor g09074(.dina(n9265), .dinb(n9229), .dout(n9266));
  jxor g09075(.dina(n9266), .dinb(n9226), .dout(n9267));
  jxor g09076(.dina(n9267), .dinb(n9181), .dout(n9268));
  jxor g09077(.dina(n9268), .dinb(n9178), .dout(n9269));
  jnot g09078(.din(n9269), .dout(n9270));
  jxor g09079(.dina(n9270), .dinb(n9055), .dout(n9271));
  jnot g09080(.din(n9045), .dout(n9272));
  jor  g09081(.dina(n9051), .dinb(n9047), .dout(n9273));
  jand g09082(.dina(n9273), .dinb(n9272), .dout(n9274));
  jxor g09083(.dina(n9274), .dinb(n9271), .dout(\asquared[69] ));
  jand g09084(.dina(n9267), .dinb(n9181), .dout(n9276));
  jand g09085(.dina(n9268), .dinb(n9178), .dout(n9277));
  jor  g09086(.dina(n9277), .dinb(n9276), .dout(n9278));
  jand g09087(.dina(n9176), .dinb(n9061), .dout(n9279));
  jand g09088(.dina(n9177), .dinb(n9058), .dout(n9280));
  jor  g09089(.dina(n9280), .dinb(n9279), .dout(n9281));
  jand g09090(.dina(n9224), .dinb(n9204), .dout(n9282));
  jand g09091(.dina(n9225), .dinb(n9186), .dout(n9283));
  jor  g09092(.dina(n9283), .dinb(n9282), .dout(n9284));
  jand g09093(.dina(n9172), .dinb(n9141), .dout(n9285));
  jand g09094(.dina(n9173), .dinb(n9103), .dout(n9286));
  jor  g09095(.dina(n9286), .dinb(n9285), .dout(n9287));
  jand g09096(.dina(n9222), .dinb(n9214), .dout(n9288));
  jand g09097(.dina(n9223), .dinb(n9207), .dout(n9289));
  jor  g09098(.dina(n9289), .dinb(n9288), .dout(n9290));
  jand g09099(.dina(n9166), .dinb(n9164), .dout(n9291));
  jnot g09100(.din(n9291), .dout(n9292));
  jand g09101(.dina(n9292), .dinb(n9169), .dout(n9293));
  jxor g09102(.dina(n9293), .dinb(n9115), .dout(n9294));
  jand g09103(.dina(n9087), .dinb(n9085), .dout(n9295));
  jnot g09104(.din(n9295), .dout(n9296));
  jand g09105(.dina(n9296), .dinb(n9090), .dout(n9297));
  jxor g09106(.dina(n9297), .dinb(n9294), .dout(n9298));
  jand g09107(.dina(n9220), .dinb(n8966), .dout(n9299));
  jand g09108(.dina(n9221), .dinb(n9217), .dout(n9300));
  jor  g09109(.dina(n9300), .dinb(n9299), .dout(n9301));
  jand g09110(.dina(n9189), .dinb(n8936), .dout(n9302));
  jand g09111(.dina(n9193), .dinb(n9190), .dout(n9303));
  jor  g09112(.dina(n9303), .dinb(n9302), .dout(n9304));
  jxor g09113(.dina(n9304), .dinb(n9301), .dout(n9305));
  jxor g09114(.dina(n9305), .dinb(n9298), .dout(n9306));
  jxor g09115(.dina(n9306), .dinb(n9290), .dout(n9307));
  jxor g09116(.dina(n9307), .dinb(n9287), .dout(n9308));
  jxor g09117(.dina(n9308), .dinb(n9284), .dout(n9309));
  jor  g09118(.dina(n9071), .dinb(n9068), .dout(n9310));
  jand g09119(.dina(n9075), .dinb(n9072), .dout(n9311));
  jnot g09120(.din(n9311), .dout(n9312));
  jand g09121(.dina(n9312), .dinb(n9310), .dout(n9313));
  jnot g09122(.din(n9313), .dout(n9314));
  jor  g09123(.dina(n9138), .dinb(n9129), .dout(n9315));
  jor  g09124(.dina(n9140), .dinb(n9120), .dout(n9316));
  jand g09125(.dina(n9316), .dinb(n9315), .dout(n9317));
  jor  g09126(.dina(n9160), .dinb(n9150), .dout(n9318));
  jor  g09127(.dina(n9171), .dinb(n9162), .dout(n9319));
  jand g09128(.dina(n9319), .dinb(n9318), .dout(n9320));
  jxor g09129(.dina(n9320), .dinb(n9317), .dout(n9321));
  jand g09130(.dina(n9258), .dinb(n9248), .dout(n9322));
  jand g09131(.dina(n9262), .dinb(n9259), .dout(n9323));
  jor  g09132(.dina(n9323), .dinb(n9322), .dout(n9324));
  jxor g09133(.dina(n9324), .dinb(n9321), .dout(n9325));
  jand g09134(.dina(n9081), .dinb(n8995), .dout(n9326));
  jor  g09135(.dina(n9326), .dinb(n9077), .dout(n9327));
  jor  g09136(.dina(n9096), .dinb(n9094), .dout(n9328));
  jand g09137(.dina(n9328), .dinb(n9100), .dout(n9329));
  jxor g09138(.dina(n9329), .dinb(n9327), .dout(n9330));
  jand g09139(.dina(n9155), .dinb(n9152), .dout(n9331));
  jnot g09140(.din(n9331), .dout(n9332));
  jand g09141(.dina(n9332), .dinb(n9158), .dout(n9333));
  jxor g09142(.dina(n9333), .dinb(n9330), .dout(n9334));
  jand g09143(.dina(n9148), .dinb(n9142), .dout(n9335));
  jor  g09144(.dina(n9335), .dinb(n9146), .dout(n9336));
  jand g09145(.dina(n9127), .dinb(n3752), .dout(n9337));
  jor  g09146(.dina(n9337), .dinb(n9125), .dout(n9338));
  jand g09147(.dina(n9133), .dinb(n9131), .dout(n9339));
  jnot g09148(.din(n9339), .dout(n9340));
  jand g09149(.dina(n9340), .dinb(n9136), .dout(n9341));
  jxor g09150(.dina(n9341), .dinb(n9338), .dout(n9342));
  jxor g09151(.dina(n9342), .dinb(n9336), .dout(n9343));
  jnot g09152(.din(n9343), .dout(n9344));
  jor  g09153(.dina(n9092), .dinb(n9083), .dout(n9345));
  jand g09154(.dina(n9102), .dinb(n9093), .dout(n9346));
  jnot g09155(.din(n9346), .dout(n9347));
  jand g09156(.dina(n9347), .dinb(n9345), .dout(n9348));
  jxor g09157(.dina(n9348), .dinb(n9344), .dout(n9349));
  jxor g09158(.dina(n9349), .dinb(n9334), .dout(n9350));
  jxor g09159(.dina(n9350), .dinb(n9325), .dout(n9351));
  jxor g09160(.dina(n9351), .dinb(n9314), .dout(n9352));
  jxor g09161(.dina(n9352), .dinb(n9309), .dout(n9353));
  jxor g09162(.dina(n9353), .dinb(n9281), .dout(n9354));
  jand g09163(.dina(n9265), .dinb(n9229), .dout(n9355));
  jand g09164(.dina(n9266), .dinb(n9226), .dout(n9356));
  jor  g09165(.dina(n9356), .dinb(n9355), .dout(n9357));
  jand g09166(.dina(n9174), .dinb(n9076), .dout(n9358));
  jand g09167(.dina(n9175), .dinb(n9064), .dout(n9359));
  jor  g09168(.dina(n9359), .dinb(n9358), .dout(n9360));
  jxor g09169(.dina(n9360), .dinb(n9357), .dout(n9361));
  jand g09170(.dina(n9263), .dinb(n9245), .dout(n9362));
  jand g09171(.dina(n9264), .dinb(n9232), .dout(n9363));
  jor  g09172(.dina(n9363), .dinb(n9362), .dout(n9364));
  jor  g09173(.dina(n9202), .dinb(n9198), .dout(n9365));
  jand g09174(.dina(n9203), .dinb(n9194), .dout(n9366));
  jnot g09175(.din(n9366), .dout(n9367));
  jand g09176(.dina(n9367), .dinb(n9365), .dout(n9368));
  jnot g09177(.din(n9368), .dout(n9369));
  jand g09178(.dina(n9212), .dinb(n8894), .dout(n9370));
  jand g09179(.dina(n9213), .dinb(n9209), .dout(n9371));
  jor  g09180(.dina(n9371), .dinb(n9370), .dout(n9372));
  jand g09181(.dina(\a[52] ), .dinb(\a[18] ), .dout(n9373));
  jand g09182(.dina(n9373), .dinb(n9106), .dout(n9374));
  jnot g09183(.din(n9374), .dout(n9375));
  jand g09184(.dina(\a[52] ), .dinb(\a[17] ), .dout(n9376));
  jand g09185(.dina(\a[51] ), .dinb(\a[18] ), .dout(n9377));
  jor  g09186(.dina(n9377), .dinb(n9376), .dout(n9378));
  jand g09187(.dina(n9378), .dinb(n9375), .dout(n9379));
  jxor g09188(.dina(n9379), .dinb(n9124), .dout(n9380));
  jand g09189(.dina(\a[41] ), .dinb(\a[28] ), .dout(n9381));
  jand g09190(.dina(n3665), .dinb(n3294), .dout(n9382));
  jnot g09191(.din(n9382), .dout(n9383));
  jand g09192(.dina(\a[40] ), .dinb(\a[29] ), .dout(n9384));
  jand g09193(.dina(\a[39] ), .dinb(\a[30] ), .dout(n9385));
  jor  g09194(.dina(n9385), .dinb(n9384), .dout(n9386));
  jand g09195(.dina(n9386), .dinb(n9383), .dout(n9387));
  jxor g09196(.dina(n9387), .dinb(n9381), .dout(n9388));
  jxor g09197(.dina(n9388), .dinb(n9380), .dout(n9389));
  jxor g09198(.dina(n9389), .dinb(n9372), .dout(n9390));
  jand g09199(.dina(\a[54] ), .dinb(\a[15] ), .dout(n9391));
  jand g09200(.dina(n7559), .dinb(n829), .dout(n9392));
  jand g09201(.dina(\a[49] ), .dinb(\a[20] ), .dout(n9393));
  jand g09202(.dina(n9393), .dinb(n9391), .dout(n9394));
  jor  g09203(.dina(n9394), .dinb(n9392), .dout(n9395));
  jand g09204(.dina(\a[53] ), .dinb(\a[16] ), .dout(n9396));
  jand g09205(.dina(n9396), .dinb(n9393), .dout(n9397));
  jnot g09206(.din(n9397), .dout(n9398));
  jand g09207(.dina(n9398), .dinb(n9395), .dout(n9399));
  jnot g09208(.din(n9399), .dout(n9400));
  jand g09209(.dina(n9400), .dinb(n9391), .dout(n9401));
  jor  g09210(.dina(n9397), .dinb(n9395), .dout(n9402));
  jnot g09211(.din(n9402), .dout(n9403));
  jor  g09212(.dina(n9396), .dinb(n9393), .dout(n9404));
  jand g09213(.dina(n9404), .dinb(n9403), .dout(n9405));
  jor  g09214(.dina(n9405), .dinb(n9401), .dout(n9406));
  jand g09215(.dina(\a[62] ), .dinb(\a[7] ), .dout(n9407));
  jand g09216(.dina(\a[35] ), .dinb(n8973), .dout(n9408));
  jxor g09217(.dina(n9408), .dinb(n9407), .dout(n9409));
  jnot g09218(.din(n9409), .dout(n9410));
  jand g09219(.dina(\a[38] ), .dinb(\a[31] ), .dout(n9411));
  jnot g09220(.din(n9411), .dout(n9412));
  jand g09221(.dina(n3138), .dinb(n2671), .dout(n9413));
  jnot g09222(.din(n9413), .dout(n9414));
  jand g09223(.dina(\a[36] ), .dinb(\a[33] ), .dout(n9415));
  jand g09224(.dina(\a[37] ), .dinb(\a[32] ), .dout(n9416));
  jor  g09225(.dina(n9416), .dinb(n9415), .dout(n9417));
  jand g09226(.dina(n9417), .dinb(n9414), .dout(n9418));
  jxor g09227(.dina(n9418), .dinb(n9412), .dout(n9419));
  jxor g09228(.dina(n9419), .dinb(n9410), .dout(n9420));
  jxor g09229(.dina(n9420), .dinb(n9406), .dout(n9421));
  jxor g09230(.dina(n9421), .dinb(n9390), .dout(n9422));
  jxor g09231(.dina(n9422), .dinb(n9369), .dout(n9423));
  jxor g09232(.dina(n9423), .dinb(n9364), .dout(n9424));
  jand g09233(.dina(n9238), .dinb(n9235), .dout(n9425));
  jnot g09234(.din(n9425), .dout(n9426));
  jor  g09235(.dina(n9244), .dinb(n9240), .dout(n9427));
  jand g09236(.dina(n9427), .dinb(n9426), .dout(n9428));
  jnot g09237(.din(n9428), .dout(n9429));
  jand g09238(.dina(\a[60] ), .dinb(\a[10] ), .dout(n9430));
  jand g09239(.dina(n9430), .dinb(n8995), .dout(n9431));
  jnot g09240(.din(n9431), .dout(n9432));
  jand g09241(.dina(\a[60] ), .dinb(\a[9] ), .dout(n9433));
  jand g09242(.dina(\a[59] ), .dinb(\a[10] ), .dout(n9434));
  jor  g09243(.dina(n9434), .dinb(n9433), .dout(n9435));
  jand g09244(.dina(n9435), .dinb(n9432), .dout(n9436));
  jxor g09245(.dina(n9436), .dinb(n9251), .dout(n9437));
  jnot g09246(.din(n9437), .dout(n9438));
  jnot g09247(.din(n9153), .dout(n9439));
  jand g09248(.dina(n4812), .dinb(n1648), .dout(n9440));
  jnot g09249(.din(n9440), .dout(n9441));
  jand g09250(.dina(\a[45] ), .dinb(\a[24] ), .dout(n9442));
  jand g09251(.dina(\a[44] ), .dinb(\a[25] ), .dout(n9443));
  jor  g09252(.dina(n9443), .dinb(n9442), .dout(n9444));
  jand g09253(.dina(n9444), .dinb(n9441), .dout(n9445));
  jxor g09254(.dina(n9445), .dinb(n9439), .dout(n9446));
  jxor g09255(.dina(n9446), .dinb(n9438), .dout(n9447));
  jnot g09256(.din(n9447), .dout(n9448));
  jnot g09257(.din(n9095), .dout(n9449));
  jand g09258(.dina(n4317), .dinb(n1927), .dout(n9450));
  jnot g09259(.din(n9450), .dout(n9451));
  jand g09260(.dina(\a[43] ), .dinb(\a[26] ), .dout(n9452));
  jand g09261(.dina(\a[42] ), .dinb(\a[27] ), .dout(n9453));
  jor  g09262(.dina(n9453), .dinb(n9452), .dout(n9454));
  jand g09263(.dina(n9454), .dinb(n9451), .dout(n9455));
  jxor g09264(.dina(n9455), .dinb(n9449), .dout(n9456));
  jxor g09265(.dina(n9456), .dinb(n9448), .dout(n9457));
  jxor g09266(.dina(n9457), .dinb(n9429), .dout(n9458));
  jand g09267(.dina(n9257), .dinb(n9250), .dout(n9459));
  jor  g09268(.dina(n9459), .dinb(n9252), .dout(n9460));
  jand g09269(.dina(\a[58] ), .dinb(\a[11] ), .dout(n9461));
  jand g09270(.dina(\a[57] ), .dinb(\a[13] ), .dout(n9462));
  jand g09271(.dina(n9462), .dinb(n9104), .dout(n9463));
  jnot g09272(.din(n9463), .dout(n9464));
  jand g09273(.dina(\a[57] ), .dinb(\a[12] ), .dout(n9465));
  jor  g09274(.dina(n9465), .dinb(n9108), .dout(n9466));
  jand g09275(.dina(n9466), .dinb(n9464), .dout(n9467));
  jxor g09276(.dina(n9467), .dinb(n9461), .dout(n9468));
  jxor g09277(.dina(n9468), .dinb(n9460), .dout(n9469));
  jnot g09278(.din(n9469), .dout(n9470));
  jand g09279(.dina(\a[55] ), .dinb(\a[14] ), .dout(n9471));
  jnot g09280(.din(n9471), .dout(n9472));
  jand g09281(.dina(n5316), .dinb(n1376), .dout(n9473));
  jnot g09282(.din(n9473), .dout(n9474));
  jand g09283(.dina(\a[48] ), .dinb(\a[21] ), .dout(n9475));
  jand g09284(.dina(\a[47] ), .dinb(\a[22] ), .dout(n9476));
  jor  g09285(.dina(n9476), .dinb(n9475), .dout(n9477));
  jand g09286(.dina(n9477), .dinb(n9474), .dout(n9478));
  jxor g09287(.dina(n9478), .dinb(n9472), .dout(n9479));
  jxor g09288(.dina(n9479), .dinb(n9470), .dout(n9480));
  jxor g09289(.dina(n9480), .dinb(n9458), .dout(n9481));
  jxor g09290(.dina(n9481), .dinb(n9424), .dout(n9482));
  jxor g09291(.dina(n9482), .dinb(n9361), .dout(n9483));
  jxor g09292(.dina(n9483), .dinb(n9354), .dout(n9484));
  jand g09293(.dina(n9484), .dinb(n9278), .dout(n9485));
  jor  g09294(.dina(n9484), .dinb(n9278), .dout(n9486));
  jnot g09295(.din(n9486), .dout(n9487));
  jor  g09296(.dina(n9487), .dinb(n9485), .dout(n9488));
  jand g09297(.dina(n9269), .dinb(n9055), .dout(n9489));
  jnot g09298(.din(n9489), .dout(n9490));
  jnot g09299(.din(n9055), .dout(n9491));
  jand g09300(.dina(n9270), .dinb(n9491), .dout(n9492));
  jor  g09301(.dina(n9274), .dinb(n9492), .dout(n9493));
  jand g09302(.dina(n9493), .dinb(n9490), .dout(n9494));
  jxor g09303(.dina(n9494), .dinb(n9488), .dout(\asquared[70] ));
  jand g09304(.dina(n9353), .dinb(n9281), .dout(n9496));
  jand g09305(.dina(n9483), .dinb(n9354), .dout(n9497));
  jor  g09306(.dina(n9497), .dinb(n9496), .dout(n9498));
  jnot g09307(.din(n9498), .dout(n9499));
  jand g09308(.dina(n9308), .dinb(n9284), .dout(n9500));
  jand g09309(.dina(n9352), .dinb(n9309), .dout(n9501));
  jor  g09310(.dina(n9501), .dinb(n9500), .dout(n9502));
  jand g09311(.dina(n9388), .dinb(n9380), .dout(n9503));
  jand g09312(.dina(n9389), .dinb(n9372), .dout(n9504));
  jor  g09313(.dina(n9504), .dinb(n9503), .dout(n9505));
  jor  g09314(.dina(n9382), .dinb(n9381), .dout(n9506));
  jand g09315(.dina(n9506), .dinb(n9386), .dout(n9507));
  jand g09316(.dina(n9451), .dinb(n9449), .dout(n9508));
  jnot g09317(.din(n9508), .dout(n9509));
  jand g09318(.dina(n9509), .dinb(n9454), .dout(n9510));
  jxor g09319(.dina(n9510), .dinb(n9507), .dout(n9511));
  jand g09320(.dina(n9441), .dinb(n9439), .dout(n9512));
  jnot g09321(.din(n9512), .dout(n9513));
  jand g09322(.dina(n9513), .dinb(n9444), .dout(n9514));
  jxor g09323(.dina(n9514), .dinb(n9511), .dout(n9515));
  jand g09324(.dina(\a[62] ), .dinb(\a[8] ), .dout(n9516));
  jor  g09325(.dina(n9407), .dinb(\a[34] ), .dout(n9517));
  jand g09326(.dina(n9517), .dinb(\a[35] ), .dout(n9518));
  jxor g09327(.dina(n9518), .dinb(n9516), .dout(n9519));
  jand g09328(.dina(n9414), .dinb(n9412), .dout(n9520));
  jnot g09329(.din(n9520), .dout(n9521));
  jand g09330(.dina(n9521), .dinb(n9417), .dout(n9522));
  jxor g09331(.dina(n9522), .dinb(n9519), .dout(n9523));
  jxor g09332(.dina(n9523), .dinb(n9515), .dout(n9524));
  jxor g09333(.dina(n9524), .dinb(n9505), .dout(n9525));
  jand g09334(.dina(n9421), .dinb(n9390), .dout(n9526));
  jand g09335(.dina(n9422), .dinb(n9369), .dout(n9527));
  jor  g09336(.dina(n9527), .dinb(n9526), .dout(n9528));
  jor  g09337(.dina(n9446), .dinb(n9438), .dout(n9529));
  jor  g09338(.dina(n9456), .dinb(n9448), .dout(n9530));
  jand g09339(.dina(n9530), .dinb(n9529), .dout(n9531));
  jand g09340(.dina(n9468), .dinb(n9460), .dout(n9532));
  jnot g09341(.din(n9532), .dout(n9533));
  jor  g09342(.dina(n9479), .dinb(n9470), .dout(n9534));
  jand g09343(.dina(n9534), .dinb(n9533), .dout(n9535));
  jxor g09344(.dina(n9535), .dinb(n9531), .dout(n9536));
  jnot g09345(.din(n9536), .dout(n9537));
  jor  g09346(.dina(n9419), .dinb(n9410), .dout(n9538));
  jand g09347(.dina(n9420), .dinb(n9406), .dout(n9539));
  jnot g09348(.din(n9539), .dout(n9540));
  jand g09349(.dina(n9540), .dinb(n9538), .dout(n9541));
  jxor g09350(.dina(n9541), .dinb(n9537), .dout(n9542));
  jxor g09351(.dina(n9542), .dinb(n9528), .dout(n9543));
  jxor g09352(.dina(n9543), .dinb(n9525), .dout(n9544));
  jxor g09353(.dina(n9544), .dinb(n9502), .dout(n9545));
  jand g09354(.dina(n9306), .dinb(n9290), .dout(n9546));
  jand g09355(.dina(n9307), .dinb(n9287), .dout(n9547));
  jor  g09356(.dina(n9547), .dinb(n9546), .dout(n9548));
  jand g09357(.dina(n9304), .dinb(n9301), .dout(n9549));
  jand g09358(.dina(n9305), .dinb(n9298), .dout(n9550));
  jor  g09359(.dina(n9550), .dinb(n9549), .dout(n9551));
  jand g09360(.dina(n9379), .dinb(n9124), .dout(n9552));
  jor  g09361(.dina(n9552), .dinb(n9374), .dout(n9553));
  jxor g09362(.dina(n9553), .dinb(n9402), .dout(n9554));
  jnot g09363(.din(n9554), .dout(n9555));
  jand g09364(.dina(\a[38] ), .dinb(\a[32] ), .dout(n9556));
  jand g09365(.dina(n3634), .dinb(n3138), .dout(n9557));
  jnot g09366(.din(n9557), .dout(n9558));
  jand g09367(.dina(\a[38] ), .dinb(\a[33] ), .dout(n9559));
  jand g09368(.dina(n9559), .dinb(n9416), .dout(n9560));
  jand g09369(.dina(n9556), .dinb(n5916), .dout(n9561));
  jor  g09370(.dina(n9561), .dinb(n9560), .dout(n9562));
  jand g09371(.dina(n9562), .dinb(n9558), .dout(n9563));
  jnot g09372(.din(n9563), .dout(n9564));
  jand g09373(.dina(n9564), .dinb(n9556), .dout(n9565));
  jnot g09374(.din(n9565), .dout(n9566));
  jor  g09375(.dina(n9562), .dinb(n9557), .dout(n9567));
  jnot g09376(.din(n5916), .dout(n9568));
  jand g09377(.dina(\a[37] ), .dinb(\a[33] ), .dout(n9569));
  jnot g09378(.din(n9569), .dout(n9570));
  jand g09379(.dina(n9570), .dinb(n9568), .dout(n9571));
  jor  g09380(.dina(n9571), .dinb(n9567), .dout(n9572));
  jand g09381(.dina(n9572), .dinb(n9566), .dout(n9573));
  jxor g09382(.dina(n9573), .dinb(n9555), .dout(n9574));
  jxor g09383(.dina(n9574), .dinb(n9551), .dout(n9575));
  jand g09384(.dina(\a[58] ), .dinb(\a[12] ), .dout(n9576));
  jnot g09385(.din(n9576), .dout(n9577));
  jand g09386(.dina(\a[46] ), .dinb(\a[24] ), .dout(n9578));
  jand g09387(.dina(n9578), .dinb(n9462), .dout(n9579));
  jnot g09388(.din(n9579), .dout(n9580));
  jand g09389(.dina(n7519), .dinb(n899), .dout(n9581));
  jand g09390(.dina(n9578), .dinb(n9576), .dout(n9582));
  jor  g09391(.dina(n9582), .dinb(n9581), .dout(n9583));
  jand g09392(.dina(n9583), .dinb(n9580), .dout(n9584));
  jor  g09393(.dina(n9584), .dinb(n9577), .dout(n9585));
  jor  g09394(.dina(n9583), .dinb(n9579), .dout(n9586));
  jnot g09395(.din(n9586), .dout(n9587));
  jor  g09396(.dina(n9578), .dinb(n9462), .dout(n9588));
  jand g09397(.dina(n9588), .dinb(n9587), .dout(n9589));
  jnot g09398(.din(n9589), .dout(n9590));
  jand g09399(.dina(n9590), .dinb(n9585), .dout(n9591));
  jand g09400(.dina(\a[61] ), .dinb(\a[9] ), .dout(n9592));
  jand g09401(.dina(\a[60] ), .dinb(\a[11] ), .dout(n9593));
  jand g09402(.dina(n9593), .dinb(n9434), .dout(n9594));
  jnot g09403(.din(n9594), .dout(n9595));
  jand g09404(.dina(\a[59] ), .dinb(\a[11] ), .dout(n9596));
  jor  g09405(.dina(n9596), .dinb(n9430), .dout(n9597));
  jand g09406(.dina(n9597), .dinb(n9595), .dout(n9598));
  jxor g09407(.dina(n9598), .dinb(n9592), .dout(n9599));
  jnot g09408(.din(n9599), .dout(n9600));
  jnot g09409(.din(n9373), .dout(n9601));
  jand g09410(.dina(n7559), .dinb(n937), .dout(n9602));
  jnot g09411(.din(n9602), .dout(n9603));
  jand g09412(.dina(\a[53] ), .dinb(\a[17] ), .dout(n9604));
  jand g09413(.dina(\a[54] ), .dinb(\a[16] ), .dout(n9605));
  jor  g09414(.dina(n9605), .dinb(n9604), .dout(n9606));
  jand g09415(.dina(n9606), .dinb(n9603), .dout(n9607));
  jxor g09416(.dina(n9607), .dinb(n9601), .dout(n9608));
  jxor g09417(.dina(n9608), .dinb(n9600), .dout(n9609));
  jnot g09418(.din(n9609), .dout(n9610));
  jxor g09419(.dina(n9610), .dinb(n9591), .dout(n9611));
  jxor g09420(.dina(n9611), .dinb(n9575), .dout(n9612));
  jxor g09421(.dina(n9612), .dinb(n9548), .dout(n9613));
  jor  g09422(.dina(n9348), .dinb(n9344), .dout(n9614));
  jand g09423(.dina(n9349), .dinb(n9334), .dout(n9615));
  jnot g09424(.din(n9615), .dout(n9616));
  jand g09425(.dina(n9616), .dinb(n9614), .dout(n9617));
  jnot g09426(.din(n9617), .dout(n9618));
  jand g09427(.dina(n9341), .dinb(n9338), .dout(n9619));
  jand g09428(.dina(n9342), .dinb(n9336), .dout(n9620));
  jor  g09429(.dina(n9620), .dinb(n9619), .dout(n9621));
  jand g09430(.dina(\a[42] ), .dinb(\a[28] ), .dout(n9622));
  jand g09431(.dina(\a[63] ), .dinb(\a[7] ), .dout(n9623));
  jand g09432(.dina(\a[47] ), .dinb(\a[23] ), .dout(n9624));
  jxor g09433(.dina(n9624), .dinb(n9623), .dout(n9625));
  jxor g09434(.dina(n9625), .dinb(n9622), .dout(n9626));
  jnot g09435(.din(n9626), .dout(n9627));
  jand g09436(.dina(\a[41] ), .dinb(\a[29] ), .dout(n9628));
  jnot g09437(.din(n9628), .dout(n9629));
  jand g09438(.dina(n3665), .dinb(n2440), .dout(n9630));
  jnot g09439(.din(n9630), .dout(n9631));
  jand g09440(.dina(\a[40] ), .dinb(\a[30] ), .dout(n9632));
  jand g09441(.dina(\a[39] ), .dinb(\a[31] ), .dout(n9633));
  jor  g09442(.dina(n9633), .dinb(n9632), .dout(n9634));
  jand g09443(.dina(n9634), .dinb(n9631), .dout(n9635));
  jxor g09444(.dina(n9635), .dinb(n9629), .dout(n9636));
  jxor g09445(.dina(n9636), .dinb(n9627), .dout(n9637));
  jxor g09446(.dina(n9637), .dinb(n9621), .dout(n9638));
  jand g09447(.dina(\a[48] ), .dinb(\a[22] ), .dout(n9639));
  jand g09448(.dina(\a[56] ), .dinb(\a[14] ), .dout(n9640));
  jand g09449(.dina(\a[55] ), .dinb(\a[15] ), .dout(n9641));
  jor  g09450(.dina(n9641), .dinb(n9640), .dout(n9642));
  jand g09451(.dina(\a[56] ), .dinb(\a[15] ), .dout(n9643));
  jand g09452(.dina(n9643), .dinb(n9471), .dout(n9644));
  jnot g09453(.din(n9644), .dout(n9645));
  jand g09454(.dina(n9645), .dinb(n9642), .dout(n9646));
  jxor g09455(.dina(n9646), .dinb(n9639), .dout(n9647));
  jnot g09456(.din(n9647), .dout(n9648));
  jand g09457(.dina(\a[45] ), .dinb(\a[25] ), .dout(n9649));
  jnot g09458(.din(n9649), .dout(n9650));
  jand g09459(.dina(n4495), .dinb(n1927), .dout(n9651));
  jnot g09460(.din(n9651), .dout(n9652));
  jand g09461(.dina(\a[44] ), .dinb(\a[26] ), .dout(n9653));
  jand g09462(.dina(\a[43] ), .dinb(\a[27] ), .dout(n9654));
  jor  g09463(.dina(n9654), .dinb(n9653), .dout(n9655));
  jand g09464(.dina(n9655), .dinb(n9652), .dout(n9656));
  jxor g09465(.dina(n9656), .dinb(n9650), .dout(n9657));
  jxor g09466(.dina(n9657), .dinb(n9648), .dout(n9658));
  jnot g09467(.din(n9658), .dout(n9659));
  jand g09468(.dina(\a[49] ), .dinb(\a[21] ), .dout(n9660));
  jnot g09469(.din(n9660), .dout(n9661));
  jand g09470(.dina(n5594), .dinb(n1287), .dout(n9662));
  jnot g09471(.din(n9662), .dout(n9663));
  jand g09472(.dina(\a[51] ), .dinb(\a[19] ), .dout(n9664));
  jand g09473(.dina(\a[50] ), .dinb(\a[20] ), .dout(n9665));
  jor  g09474(.dina(n9665), .dinb(n9664), .dout(n9666));
  jand g09475(.dina(n9666), .dinb(n9663), .dout(n9667));
  jxor g09476(.dina(n9667), .dinb(n9661), .dout(n9668));
  jxor g09477(.dina(n9668), .dinb(n9659), .dout(n9669));
  jxor g09478(.dina(n9669), .dinb(n9638), .dout(n9670));
  jxor g09479(.dina(n9670), .dinb(n9618), .dout(n9671));
  jxor g09480(.dina(n9671), .dinb(n9613), .dout(n9672));
  jxor g09481(.dina(n9672), .dinb(n9545), .dout(n9673));
  jand g09482(.dina(n9423), .dinb(n9364), .dout(n9674));
  jand g09483(.dina(n9481), .dinb(n9424), .dout(n9675));
  jor  g09484(.dina(n9675), .dinb(n9674), .dout(n9676));
  jand g09485(.dina(n9350), .dinb(n9325), .dout(n9677));
  jand g09486(.dina(n9351), .dinb(n9314), .dout(n9678));
  jor  g09487(.dina(n9678), .dinb(n9677), .dout(n9679));
  jand g09488(.dina(n9457), .dinb(n9429), .dout(n9680));
  jand g09489(.dina(n9480), .dinb(n9458), .dout(n9681));
  jor  g09490(.dina(n9681), .dinb(n9680), .dout(n9682));
  jor  g09491(.dina(n9320), .dinb(n9317), .dout(n9683));
  jand g09492(.dina(n9324), .dinb(n9321), .dout(n9684));
  jnot g09493(.din(n9684), .dout(n9685));
  jand g09494(.dina(n9685), .dinb(n9683), .dout(n9686));
  jnot g09495(.din(n9686), .dout(n9687));
  jand g09496(.dina(n9436), .dinb(n9251), .dout(n9688));
  jor  g09497(.dina(n9688), .dinb(n9431), .dout(n9689));
  jor  g09498(.dina(n9463), .dinb(n9461), .dout(n9690));
  jand g09499(.dina(n9690), .dinb(n9466), .dout(n9691));
  jxor g09500(.dina(n9691), .dinb(n9689), .dout(n9692));
  jand g09501(.dina(n9474), .dinb(n9472), .dout(n9693));
  jnot g09502(.din(n9693), .dout(n9694));
  jand g09503(.dina(n9694), .dinb(n9477), .dout(n9695));
  jxor g09504(.dina(n9695), .dinb(n9692), .dout(n9696));
  jand g09505(.dina(n9329), .dinb(n9327), .dout(n9697));
  jand g09506(.dina(n9333), .dinb(n9330), .dout(n9698));
  jor  g09507(.dina(n9698), .dinb(n9697), .dout(n9699));
  jand g09508(.dina(n9293), .dinb(n9115), .dout(n9700));
  jand g09509(.dina(n9297), .dinb(n9294), .dout(n9701));
  jor  g09510(.dina(n9701), .dinb(n9700), .dout(n9702));
  jxor g09511(.dina(n9702), .dinb(n9699), .dout(n9703));
  jxor g09512(.dina(n9703), .dinb(n9696), .dout(n9704));
  jxor g09513(.dina(n9704), .dinb(n9687), .dout(n9705));
  jxor g09514(.dina(n9705), .dinb(n9682), .dout(n9706));
  jxor g09515(.dina(n9706), .dinb(n9679), .dout(n9707));
  jxor g09516(.dina(n9707), .dinb(n9676), .dout(n9708));
  jand g09517(.dina(n9360), .dinb(n9357), .dout(n9709));
  jand g09518(.dina(n9482), .dinb(n9361), .dout(n9710));
  jor  g09519(.dina(n9710), .dinb(n9709), .dout(n9711));
  jxor g09520(.dina(n9711), .dinb(n9708), .dout(n9712));
  jxor g09521(.dina(n9712), .dinb(n9673), .dout(n9713));
  jxor g09522(.dina(n9713), .dinb(n9499), .dout(n9714));
  jnot g09523(.din(n9485), .dout(n9715));
  jor  g09524(.dina(n9494), .dinb(n9487), .dout(n9716));
  jand g09525(.dina(n9716), .dinb(n9715), .dout(n9717));
  jxor g09526(.dina(n9717), .dinb(n9714), .dout(\asquared[71] ));
  jand g09527(.dina(n9711), .dinb(n9708), .dout(n9719));
  jand g09528(.dina(n9712), .dinb(n9673), .dout(n9720));
  jor  g09529(.dina(n9720), .dinb(n9719), .dout(n9721));
  jnot g09530(.din(n9721), .dout(n9722));
  jand g09531(.dina(n9612), .dinb(n9548), .dout(n9723));
  jand g09532(.dina(n9671), .dinb(n9613), .dout(n9724));
  jor  g09533(.dina(n9724), .dinb(n9723), .dout(n9725));
  jand g09534(.dina(n9518), .dinb(n9516), .dout(n9726));
  jand g09535(.dina(n9522), .dinb(n9519), .dout(n9727));
  jor  g09536(.dina(n9727), .dinb(n9726), .dout(n9728));
  jnot g09537(.din(n9728), .dout(n9729));
  jand g09538(.dina(n9553), .dinb(n9402), .dout(n9730));
  jnot g09539(.din(n9730), .dout(n9731));
  jor  g09540(.dina(n9573), .dinb(n9555), .dout(n9732));
  jand g09541(.dina(n9732), .dinb(n9731), .dout(n9733));
  jxor g09542(.dina(n9733), .dinb(n9729), .dout(n9734));
  jand g09543(.dina(n9510), .dinb(n9507), .dout(n9735));
  jand g09544(.dina(n9514), .dinb(n9511), .dout(n9736));
  jor  g09545(.dina(n9736), .dinb(n9735), .dout(n9737));
  jxor g09546(.dina(n9737), .dinb(n9734), .dout(n9738));
  jand g09547(.dina(n9523), .dinb(n9515), .dout(n9739));
  jand g09548(.dina(n9524), .dinb(n9505), .dout(n9740));
  jor  g09549(.dina(n9740), .dinb(n9739), .dout(n9741));
  jxor g09550(.dina(n9741), .dinb(n9738), .dout(n9742));
  jand g09551(.dina(n9574), .dinb(n9551), .dout(n9743));
  jand g09552(.dina(n9611), .dinb(n9575), .dout(n9744));
  jor  g09553(.dina(n9744), .dinb(n9743), .dout(n9745));
  jxor g09554(.dina(n9745), .dinb(n9742), .dout(n9746));
  jand g09555(.dina(n9542), .dinb(n9528), .dout(n9747));
  jand g09556(.dina(n9543), .dinb(n9525), .dout(n9748));
  jor  g09557(.dina(n9748), .dinb(n9747), .dout(n9749));
  jxor g09558(.dina(n9749), .dinb(n9746), .dout(n9750));
  jxor g09559(.dina(n9750), .dinb(n9725), .dout(n9751));
  jand g09560(.dina(n9544), .dinb(n9502), .dout(n9752));
  jand g09561(.dina(n9672), .dinb(n9545), .dout(n9753));
  jor  g09562(.dina(n9753), .dinb(n9752), .dout(n9754));
  jxor g09563(.dina(n9754), .dinb(n9751), .dout(n9755));
  jand g09564(.dina(n9706), .dinb(n9679), .dout(n9756));
  jand g09565(.dina(n9707), .dinb(n9676), .dout(n9757));
  jor  g09566(.dina(n9757), .dinb(n9756), .dout(n9758));
  jand g09567(.dina(n9669), .dinb(n9638), .dout(n9759));
  jand g09568(.dina(n9670), .dinb(n9618), .dout(n9760));
  jor  g09569(.dina(n9760), .dinb(n9759), .dout(n9761));
  jor  g09570(.dina(n9608), .dinb(n9600), .dout(n9762));
  jor  g09571(.dina(n9610), .dinb(n9591), .dout(n9763));
  jand g09572(.dina(n9763), .dinb(n9762), .dout(n9764));
  jnot g09573(.din(n9764), .dout(n9765));
  jand g09574(.dina(n9691), .dinb(n9689), .dout(n9766));
  jand g09575(.dina(n9695), .dinb(n9692), .dout(n9767));
  jor  g09576(.dina(n9767), .dinb(n9766), .dout(n9768));
  jxor g09577(.dina(n9768), .dinb(n9765), .dout(n9769));
  jnot g09578(.din(n9769), .dout(n9770));
  jor  g09579(.dina(n9657), .dinb(n9648), .dout(n9771));
  jor  g09580(.dina(n9668), .dinb(n9659), .dout(n9772));
  jand g09581(.dina(n9772), .dinb(n9771), .dout(n9773));
  jxor g09582(.dina(n9773), .dinb(n9770), .dout(n9774));
  jxor g09583(.dina(n9774), .dinb(n9761), .dout(n9775));
  jor  g09584(.dina(n9636), .dinb(n9627), .dout(n9776));
  jand g09585(.dina(n9637), .dinb(n9621), .dout(n9777));
  jnot g09586(.din(n9777), .dout(n9778));
  jand g09587(.dina(n9778), .dinb(n9776), .dout(n9779));
  jnot g09588(.din(n9779), .dout(n9780));
  jand g09589(.dina(n9598), .dinb(n9592), .dout(n9781));
  jor  g09590(.dina(n9781), .dinb(n9594), .dout(n9782));
  jxor g09591(.dina(n9782), .dinb(n9586), .dout(n9783));
  jand g09592(.dina(n9652), .dinb(n9650), .dout(n9784));
  jnot g09593(.din(n9784), .dout(n9785));
  jand g09594(.dina(n9785), .dinb(n9655), .dout(n9786));
  jxor g09595(.dina(n9786), .dinb(n9783), .dout(n9787));
  jand g09596(.dina(n9624), .dinb(n9623), .dout(n9788));
  jand g09597(.dina(n9625), .dinb(n9622), .dout(n9789));
  jor  g09598(.dina(n9789), .dinb(n9788), .dout(n9790));
  jand g09599(.dina(n9646), .dinb(n9639), .dout(n9791));
  jor  g09600(.dina(n9791), .dinb(n9644), .dout(n9792));
  jand g09601(.dina(n9631), .dinb(n9629), .dout(n9793));
  jnot g09602(.din(n9793), .dout(n9794));
  jand g09603(.dina(n9794), .dinb(n9634), .dout(n9795));
  jxor g09604(.dina(n9795), .dinb(n9792), .dout(n9796));
  jxor g09605(.dina(n9796), .dinb(n9790), .dout(n9797));
  jxor g09606(.dina(n9797), .dinb(n9787), .dout(n9798));
  jxor g09607(.dina(n9798), .dinb(n9780), .dout(n9799));
  jxor g09608(.dina(n9799), .dinb(n9775), .dout(n9800));
  jxor g09609(.dina(n9800), .dinb(n9758), .dout(n9801));
  jand g09610(.dina(n9704), .dinb(n9687), .dout(n9802));
  jand g09611(.dina(n9705), .dinb(n9682), .dout(n9803));
  jor  g09612(.dina(n9803), .dinb(n9802), .dout(n9804));
  jand g09613(.dina(n9702), .dinb(n9699), .dout(n9805));
  jand g09614(.dina(n9703), .dinb(n9696), .dout(n9806));
  jor  g09615(.dina(n9806), .dinb(n9805), .dout(n9807));
  jand g09616(.dina(n9603), .dinb(n9601), .dout(n9808));
  jnot g09617(.din(n9808), .dout(n9809));
  jand g09618(.dina(n9809), .dinb(n9606), .dout(n9810));
  jxor g09619(.dina(n9810), .dinb(n9567), .dout(n9811));
  jnot g09620(.din(n9593), .dout(n9812));
  jand g09621(.dina(n8387), .dinb(n436), .dout(n9813));
  jnot g09622(.din(n9813), .dout(n9814));
  jand g09623(.dina(\a[63] ), .dinb(\a[8] ), .dout(n9815));
  jand g09624(.dina(\a[61] ), .dinb(\a[10] ), .dout(n9816));
  jor  g09625(.dina(n9816), .dinb(n9815), .dout(n9817));
  jand g09626(.dina(n9817), .dinb(n9814), .dout(n9818));
  jxor g09627(.dina(n9818), .dinb(n9812), .dout(n9819));
  jnot g09628(.din(n9819), .dout(n9820));
  jxor g09629(.dina(n9820), .dinb(n9811), .dout(n9821));
  jxor g09630(.dina(n9821), .dinb(n9807), .dout(n9822));
  jnot g09631(.din(n9559), .dout(n9823));
  jand g09632(.dina(\a[37] ), .dinb(\a[34] ), .dout(n9824));
  jand g09633(.dina(n9824), .dinb(n3243), .dout(n9825));
  jnot g09634(.din(n9825), .dout(n9826));
  jand g09635(.dina(n9559), .dinb(n3243), .dout(n9827));
  jand g09636(.dina(\a[38] ), .dinb(\a[34] ), .dout(n9828));
  jand g09637(.dina(n9828), .dinb(n9569), .dout(n9829));
  jor  g09638(.dina(n9829), .dinb(n9827), .dout(n9830));
  jand g09639(.dina(n9830), .dinb(n9826), .dout(n9831));
  jor  g09640(.dina(n9831), .dinb(n9823), .dout(n9832));
  jor  g09641(.dina(n9830), .dinb(n9825), .dout(n9833));
  jnot g09642(.din(n9833), .dout(n9834));
  jor  g09643(.dina(n9824), .dinb(n3243), .dout(n9835));
  jand g09644(.dina(n9835), .dinb(n9834), .dout(n9836));
  jnot g09645(.din(n9836), .dout(n9837));
  jand g09646(.dina(n9837), .dinb(n9832), .dout(n9838));
  jand g09647(.dina(\a[49] ), .dinb(\a[22] ), .dout(n9839));
  jand g09648(.dina(\a[62] ), .dinb(\a[9] ), .dout(n9840));
  jor  g09649(.dina(n9840), .dinb(\a[36] ), .dout(n9841));
  jand g09650(.dina(n4129), .dinb(\a[62] ), .dout(n9842));
  jnot g09651(.din(n9842), .dout(n9843));
  jand g09652(.dina(n9843), .dinb(n9841), .dout(n9844));
  jxor g09653(.dina(n9844), .dinb(n9839), .dout(n9845));
  jnot g09654(.din(n9845), .dout(n9846));
  jand g09655(.dina(\a[50] ), .dinb(\a[21] ), .dout(n9847));
  jnot g09656(.din(n9847), .dout(n9848));
  jand g09657(.dina(\a[52] ), .dinb(\a[20] ), .dout(n9849));
  jand g09658(.dina(n9849), .dinb(n9664), .dout(n9850));
  jnot g09659(.din(n9850), .dout(n9851));
  jand g09660(.dina(\a[52] ), .dinb(\a[19] ), .dout(n9852));
  jand g09661(.dina(\a[51] ), .dinb(\a[20] ), .dout(n9853));
  jor  g09662(.dina(n9853), .dinb(n9852), .dout(n9854));
  jand g09663(.dina(n9854), .dinb(n9851), .dout(n9855));
  jxor g09664(.dina(n9855), .dinb(n9848), .dout(n9856));
  jxor g09665(.dina(n9856), .dinb(n9846), .dout(n9857));
  jnot g09666(.din(n9857), .dout(n9858));
  jxor g09667(.dina(n9858), .dinb(n9838), .dout(n9859));
  jxor g09668(.dina(n9859), .dinb(n9822), .dout(n9860));
  jxor g09669(.dina(n9860), .dinb(n9804), .dout(n9861));
  jor  g09670(.dina(n9535), .dinb(n9531), .dout(n9862));
  jor  g09671(.dina(n9541), .dinb(n9537), .dout(n9863));
  jand g09672(.dina(n9863), .dinb(n9862), .dout(n9864));
  jnot g09673(.din(n9864), .dout(n9865));
  jand g09674(.dina(\a[44] ), .dinb(\a[27] ), .dout(n9866));
  jand g09675(.dina(n4317), .dinb(n2653), .dout(n9867));
  jnot g09676(.din(n9867), .dout(n9868));
  jand g09677(.dina(\a[43] ), .dinb(\a[28] ), .dout(n9869));
  jand g09678(.dina(\a[42] ), .dinb(\a[29] ), .dout(n9870));
  jor  g09679(.dina(n9870), .dinb(n9869), .dout(n9871));
  jand g09680(.dina(n9871), .dinb(n9868), .dout(n9872));
  jxor g09681(.dina(n9872), .dinb(n9866), .dout(n9873));
  jnot g09682(.din(n9873), .dout(n9874));
  jand g09683(.dina(\a[41] ), .dinb(\a[30] ), .dout(n9875));
  jnot g09684(.din(n9875), .dout(n9876));
  jand g09685(.dina(n3665), .dinb(n3269), .dout(n9877));
  jnot g09686(.din(n9877), .dout(n9878));
  jand g09687(.dina(\a[40] ), .dinb(\a[31] ), .dout(n9879));
  jand g09688(.dina(\a[39] ), .dinb(\a[32] ), .dout(n9880));
  jor  g09689(.dina(n9880), .dinb(n9879), .dout(n9881));
  jand g09690(.dina(n9881), .dinb(n9878), .dout(n9882));
  jxor g09691(.dina(n9882), .dinb(n9876), .dout(n9883));
  jxor g09692(.dina(n9883), .dinb(n9874), .dout(n9884));
  jand g09693(.dina(\a[48] ), .dinb(\a[23] ), .dout(n9885));
  jand g09694(.dina(n7559), .dinb(n1107), .dout(n9886));
  jnot g09695(.din(n9886), .dout(n9887));
  jand g09696(.dina(\a[53] ), .dinb(\a[18] ), .dout(n9888));
  jand g09697(.dina(\a[54] ), .dinb(\a[17] ), .dout(n9889));
  jor  g09698(.dina(n9889), .dinb(n9888), .dout(n9890));
  jand g09699(.dina(n9890), .dinb(n9887), .dout(n9891));
  jxor g09700(.dina(n9891), .dinb(n9885), .dout(n9892));
  jxor g09701(.dina(n9892), .dinb(n9884), .dout(n9893));
  jand g09702(.dina(\a[59] ), .dinb(\a[13] ), .dout(n9894));
  jand g09703(.dina(n9894), .dinb(n9576), .dout(n9895));
  jnot g09704(.din(n9895), .dout(n9896));
  jand g09705(.dina(\a[59] ), .dinb(\a[12] ), .dout(n9897));
  jand g09706(.dina(\a[58] ), .dinb(\a[13] ), .dout(n9898));
  jor  g09707(.dina(n9898), .dinb(n9897), .dout(n9899));
  jand g09708(.dina(n9899), .dinb(n9896), .dout(n9900));
  jand g09709(.dina(n9663), .dinb(n9661), .dout(n9901));
  jnot g09710(.din(n9901), .dout(n9902));
  jand g09711(.dina(n9902), .dinb(n9666), .dout(n9903));
  jxor g09712(.dina(n9903), .dinb(n9900), .dout(n9904));
  jand g09713(.dina(\a[57] ), .dinb(\a[14] ), .dout(n9905));
  jand g09714(.dina(\a[56] ), .dinb(\a[16] ), .dout(n9906));
  jand g09715(.dina(n9906), .dinb(n9641), .dout(n9907));
  jnot g09716(.din(n9907), .dout(n9908));
  jand g09717(.dina(\a[55] ), .dinb(\a[16] ), .dout(n9909));
  jor  g09718(.dina(n9909), .dinb(n9643), .dout(n9910));
  jand g09719(.dina(n9910), .dinb(n9908), .dout(n9911));
  jxor g09720(.dina(n9911), .dinb(n9905), .dout(n9912));
  jnot g09721(.din(n9912), .dout(n9913));
  jand g09722(.dina(\a[47] ), .dinb(\a[24] ), .dout(n9914));
  jnot g09723(.din(n9914), .dout(n9915));
  jand g09724(.dina(\a[46] ), .dinb(\a[26] ), .dout(n9916));
  jand g09725(.dina(n9916), .dinb(n9649), .dout(n9917));
  jnot g09726(.din(n9917), .dout(n9918));
  jand g09727(.dina(\a[46] ), .dinb(\a[25] ), .dout(n9919));
  jand g09728(.dina(\a[45] ), .dinb(\a[26] ), .dout(n9920));
  jor  g09729(.dina(n9920), .dinb(n9919), .dout(n9921));
  jand g09730(.dina(n9921), .dinb(n9918), .dout(n9922));
  jxor g09731(.dina(n9922), .dinb(n9915), .dout(n9923));
  jxor g09732(.dina(n9923), .dinb(n9913), .dout(n9924));
  jxor g09733(.dina(n9924), .dinb(n9904), .dout(n9925));
  jxor g09734(.dina(n9925), .dinb(n9893), .dout(n9926));
  jxor g09735(.dina(n9926), .dinb(n9865), .dout(n9927));
  jxor g09736(.dina(n9927), .dinb(n9861), .dout(n9928));
  jxor g09737(.dina(n9928), .dinb(n9801), .dout(n9929));
  jxor g09738(.dina(n9929), .dinb(n9755), .dout(n9930));
  jxor g09739(.dina(n9930), .dinb(n9722), .dout(n9931));
  jand g09740(.dina(n9713), .dinb(n9498), .dout(n9932));
  jnot g09741(.din(n9932), .dout(n9933));
  jnot g09742(.din(n9713), .dout(n9934));
  jand g09743(.dina(n9934), .dinb(n9499), .dout(n9935));
  jor  g09744(.dina(n9717), .dinb(n9935), .dout(n9936));
  jand g09745(.dina(n9936), .dinb(n9933), .dout(n9937));
  jxor g09746(.dina(n9937), .dinb(n9931), .dout(\asquared[72] ));
  jand g09747(.dina(n9860), .dinb(n9804), .dout(n9939));
  jand g09748(.dina(n9927), .dinb(n9861), .dout(n9940));
  jor  g09749(.dina(n9940), .dinb(n9939), .dout(n9941));
  jand g09750(.dina(n9797), .dinb(n9787), .dout(n9942));
  jand g09751(.dina(n9798), .dinb(n9780), .dout(n9943));
  jor  g09752(.dina(n9943), .dinb(n9942), .dout(n9944));
  jand g09753(.dina(n9795), .dinb(n9792), .dout(n9945));
  jand g09754(.dina(n9796), .dinb(n9790), .dout(n9946));
  jor  g09755(.dina(n9946), .dinb(n9945), .dout(n9947));
  jand g09756(.dina(n9810), .dinb(n9567), .dout(n9948));
  jand g09757(.dina(n9820), .dinb(n9811), .dout(n9949));
  jor  g09758(.dina(n9949), .dinb(n9948), .dout(n9950));
  jand g09759(.dina(\a[43] ), .dinb(\a[29] ), .dout(n9951));
  jand g09760(.dina(n4514), .dinb(n2440), .dout(n9952));
  jnot g09761(.din(n9952), .dout(n9953));
  jand g09762(.dina(\a[42] ), .dinb(\a[30] ), .dout(n9954));
  jor  g09763(.dina(n9954), .dinb(n4239), .dout(n9955));
  jand g09764(.dina(n9955), .dinb(n9953), .dout(n9956));
  jxor g09765(.dina(n9956), .dinb(n9951), .dout(n9957));
  jxor g09766(.dina(n9957), .dinb(n9950), .dout(n9958));
  jxor g09767(.dina(n9958), .dinb(n9947), .dout(n9959));
  jxor g09768(.dina(n9959), .dinb(n9944), .dout(n9960));
  jand g09769(.dina(n9821), .dinb(n9807), .dout(n9961));
  jand g09770(.dina(n9859), .dinb(n9822), .dout(n9962));
  jor  g09771(.dina(n9962), .dinb(n9961), .dout(n9963));
  jxor g09772(.dina(n9963), .dinb(n9960), .dout(n9964));
  jand g09773(.dina(n9774), .dinb(n9761), .dout(n9965));
  jand g09774(.dina(n9799), .dinb(n9775), .dout(n9966));
  jor  g09775(.dina(n9966), .dinb(n9965), .dout(n9967));
  jxor g09776(.dina(n9967), .dinb(n9964), .dout(n9968));
  jxor g09777(.dina(n9968), .dinb(n9941), .dout(n9969));
  jand g09778(.dina(n9800), .dinb(n9758), .dout(n9970));
  jand g09779(.dina(n9928), .dinb(n9801), .dout(n9971));
  jor  g09780(.dina(n9971), .dinb(n9970), .dout(n9972));
  jxor g09781(.dina(n9972), .dinb(n9969), .dout(n9973));
  jand g09782(.dina(n9749), .dinb(n9746), .dout(n9974));
  jand g09783(.dina(n9750), .dinb(n9725), .dout(n9975));
  jor  g09784(.dina(n9975), .dinb(n9974), .dout(n9976));
  jor  g09785(.dina(n9883), .dinb(n9874), .dout(n9977));
  jand g09786(.dina(n9892), .dinb(n9884), .dout(n9978));
  jnot g09787(.din(n9978), .dout(n9979));
  jand g09788(.dina(n9979), .dinb(n9977), .dout(n9980));
  jnot g09789(.din(n9980), .dout(n9981));
  jand g09790(.dina(n9782), .dinb(n9586), .dout(n9982));
  jand g09791(.dina(n9786), .dinb(n9783), .dout(n9983));
  jor  g09792(.dina(n9983), .dinb(n9982), .dout(n9984));
  jxor g09793(.dina(n9984), .dinb(n9981), .dout(n9985));
  jnot g09794(.din(n9985), .dout(n9986));
  jor  g09795(.dina(n9856), .dinb(n9846), .dout(n9987));
  jor  g09796(.dina(n9858), .dinb(n9838), .dout(n9988));
  jand g09797(.dina(n9988), .dinb(n9987), .dout(n9989));
  jxor g09798(.dina(n9989), .dinb(n9986), .dout(n9990));
  jand g09799(.dina(n9925), .dinb(n9893), .dout(n9991));
  jand g09800(.dina(n9926), .dinb(n9865), .dout(n9992));
  jor  g09801(.dina(n9992), .dinb(n9991), .dout(n9993));
  jxor g09802(.dina(n9993), .dinb(n9990), .dout(n9994));
  jor  g09803(.dina(n9923), .dinb(n9913), .dout(n9995));
  jand g09804(.dina(n9924), .dinb(n9904), .dout(n9996));
  jnot g09805(.din(n9996), .dout(n9997));
  jand g09806(.dina(n9997), .dinb(n9995), .dout(n9998));
  jnot g09807(.din(n9998), .dout(n9999));
  jand g09808(.dina(n9872), .dinb(n9866), .dout(n10000));
  jor  g09809(.dina(n10000), .dinb(n9867), .dout(n10001));
  jor  g09810(.dina(n9886), .dinb(n9885), .dout(n10002));
  jand g09811(.dina(n10002), .dinb(n9890), .dout(n10003));
  jxor g09812(.dina(n10003), .dinb(n10001), .dout(n10004));
  jand g09813(.dina(n9878), .dinb(n9876), .dout(n10005));
  jnot g09814(.din(n10005), .dout(n10006));
  jand g09815(.dina(n10006), .dinb(n9881), .dout(n10007));
  jxor g09816(.dina(n10007), .dinb(n10004), .dout(n10008));
  jand g09817(.dina(n9844), .dinb(n9839), .dout(n10009));
  jor  g09818(.dina(n10009), .dinb(n9842), .dout(n10010));
  jxor g09819(.dina(n10010), .dinb(n9833), .dout(n10011));
  jand g09820(.dina(n9851), .dinb(n9848), .dout(n10012));
  jnot g09821(.din(n10012), .dout(n10013));
  jand g09822(.dina(n10013), .dinb(n9854), .dout(n10014));
  jxor g09823(.dina(n10014), .dinb(n10011), .dout(n10015));
  jxor g09824(.dina(n10015), .dinb(n10008), .dout(n10016));
  jxor g09825(.dina(n10016), .dinb(n9999), .dout(n10017));
  jxor g09826(.dina(n10017), .dinb(n9994), .dout(n10018));
  jxor g09827(.dina(n10018), .dinb(n9976), .dout(n10019));
  jand g09828(.dina(n9768), .dinb(n9765), .dout(n10020));
  jnot g09829(.din(n10020), .dout(n10021));
  jor  g09830(.dina(n9773), .dinb(n9770), .dout(n10022));
  jand g09831(.dina(n10022), .dinb(n10021), .dout(n10023));
  jnot g09832(.din(n10023), .dout(n10024));
  jand g09833(.dina(n9903), .dinb(n9900), .dout(n10025));
  jor  g09834(.dina(n10025), .dinb(n9895), .dout(n10026));
  jand g09835(.dina(\a[60] ), .dinb(\a[12] ), .dout(n10027));
  jnot g09836(.din(n10027), .dout(n10028));
  jand g09837(.dina(n5316), .dinb(n1648), .dout(n10029));
  jnot g09838(.din(n10029), .dout(n10030));
  jand g09839(.dina(\a[47] ), .dinb(\a[25] ), .dout(n10031));
  jand g09840(.dina(\a[48] ), .dinb(\a[24] ), .dout(n10032));
  jor  g09841(.dina(n10032), .dinb(n10031), .dout(n10033));
  jand g09842(.dina(n10033), .dinb(n10030), .dout(n10034));
  jxor g09843(.dina(n10034), .dinb(n10028), .dout(n10035));
  jnot g09844(.din(n10035), .dout(n10036));
  jxor g09845(.dina(n10036), .dinb(n10026), .dout(n10037));
  jand g09846(.dina(\a[63] ), .dinb(\a[9] ), .dout(n10038));
  jand g09847(.dina(n8702), .dinb(n655), .dout(n10039));
  jnot g09848(.din(n10039), .dout(n10040));
  jand g09849(.dina(\a[62] ), .dinb(\a[10] ), .dout(n10041));
  jand g09850(.dina(\a[61] ), .dinb(\a[11] ), .dout(n10042));
  jor  g09851(.dina(n10042), .dinb(n10041), .dout(n10043));
  jand g09852(.dina(n10043), .dinb(n10040), .dout(n10044));
  jxor g09853(.dina(n10044), .dinb(n10038), .dout(n10045));
  jxor g09854(.dina(n10045), .dinb(n10037), .dout(n10046));
  jand g09855(.dina(\a[55] ), .dinb(\a[17] ), .dout(n10047));
  jand g09856(.dina(\a[54] ), .dinb(\a[52] ), .dout(n10048));
  jand g09857(.dina(n10048), .dinb(n1181), .dout(n10049));
  jnot g09858(.din(n10049), .dout(n10050));
  jand g09859(.dina(\a[55] ), .dinb(\a[18] ), .dout(n10051));
  jand g09860(.dina(n10051), .dinb(n9889), .dout(n10052));
  jand g09861(.dina(n10047), .dinb(n9849), .dout(n10053));
  jor  g09862(.dina(n10053), .dinb(n10052), .dout(n10054));
  jand g09863(.dina(n10054), .dinb(n10050), .dout(n10055));
  jnot g09864(.din(n10055), .dout(n10056));
  jand g09865(.dina(n10056), .dinb(n10047), .dout(n10057));
  jand g09866(.dina(\a[54] ), .dinb(\a[18] ), .dout(n10058));
  jor  g09867(.dina(n10058), .dinb(n9849), .dout(n10059));
  jor  g09868(.dina(n10054), .dinb(n10049), .dout(n10060));
  jnot g09869(.din(n10060), .dout(n10061));
  jand g09870(.dina(n10061), .dinb(n10059), .dout(n10062));
  jor  g09871(.dina(n10062), .dinb(n10057), .dout(n10063));
  jand g09872(.dina(\a[40] ), .dinb(\a[32] ), .dout(n10064));
  jand g09873(.dina(\a[49] ), .dinb(\a[23] ), .dout(n10065));
  jxor g09874(.dina(n10065), .dinb(n9906), .dout(n10066));
  jxor g09875(.dina(n10066), .dinb(n10064), .dout(n10067));
  jnot g09876(.din(n10067), .dout(n10068));
  jand g09877(.dina(\a[37] ), .dinb(\a[35] ), .dout(n10069));
  jnot g09878(.din(n10069), .dout(n10070));
  jand g09879(.dina(n5594), .dinb(n1376), .dout(n10071));
  jnot g09880(.din(n10071), .dout(n10072));
  jand g09881(.dina(\a[51] ), .dinb(\a[21] ), .dout(n10073));
  jand g09882(.dina(\a[50] ), .dinb(\a[22] ), .dout(n10074));
  jor  g09883(.dina(n10074), .dinb(n10073), .dout(n10075));
  jand g09884(.dina(n10075), .dinb(n10072), .dout(n10076));
  jxor g09885(.dina(n10076), .dinb(n10070), .dout(n10077));
  jxor g09886(.dina(n10077), .dinb(n10068), .dout(n10078));
  jxor g09887(.dina(n10078), .dinb(n10063), .dout(n10079));
  jxor g09888(.dina(n10079), .dinb(n10046), .dout(n10080));
  jxor g09889(.dina(n10080), .dinb(n10024), .dout(n10081));
  jand g09890(.dina(n9741), .dinb(n9738), .dout(n10082));
  jand g09891(.dina(n9745), .dinb(n9742), .dout(n10083));
  jor  g09892(.dina(n10083), .dinb(n10082), .dout(n10084));
  jand g09893(.dina(n9911), .dinb(n9905), .dout(n10085));
  jor  g09894(.dina(n10085), .dinb(n9907), .dout(n10086));
  jand g09895(.dina(n9918), .dinb(n9915), .dout(n10087));
  jnot g09896(.din(n10087), .dout(n10088));
  jand g09897(.dina(n10088), .dinb(n9921), .dout(n10089));
  jxor g09898(.dina(n10089), .dinb(n10086), .dout(n10090));
  jand g09899(.dina(n9814), .dinb(n9812), .dout(n10091));
  jnot g09900(.din(n10091), .dout(n10092));
  jand g09901(.dina(n10092), .dinb(n9817), .dout(n10093));
  jxor g09902(.dina(n10093), .dinb(n10090), .dout(n10094));
  jnot g09903(.din(n10094), .dout(n10095));
  jor  g09904(.dina(n9733), .dinb(n9729), .dout(n10096));
  jand g09905(.dina(n9737), .dinb(n9734), .dout(n10097));
  jnot g09906(.din(n10097), .dout(n10098));
  jand g09907(.dina(n10098), .dinb(n10096), .dout(n10099));
  jxor g09908(.dina(n10099), .dinb(n10095), .dout(n10100));
  jand g09909(.dina(n7519), .dinb(n976), .dout(n10101));
  jnot g09910(.din(n10101), .dout(n10102));
  jand g09911(.dina(\a[58] ), .dinb(\a[14] ), .dout(n10103));
  jand g09912(.dina(\a[57] ), .dinb(\a[15] ), .dout(n10104));
  jor  g09913(.dina(n10104), .dinb(n10103), .dout(n10105));
  jand g09914(.dina(n10105), .dinb(n10102), .dout(n10106));
  jxor g09915(.dina(n10106), .dinb(n9894), .dout(n10107));
  jand g09916(.dina(n4812), .dinb(n2042), .dout(n10108));
  jnot g09917(.din(n10108), .dout(n10109));
  jand g09918(.dina(\a[45] ), .dinb(\a[27] ), .dout(n10110));
  jand g09919(.dina(\a[44] ), .dinb(\a[28] ), .dout(n10111));
  jor  g09920(.dina(n10111), .dinb(n10110), .dout(n10112));
  jand g09921(.dina(n10112), .dinb(n10109), .dout(n10113));
  jxor g09922(.dina(n10113), .dinb(n9916), .dout(n10114));
  jxor g09923(.dina(n10114), .dinb(n10107), .dout(n10115));
  jnot g09924(.din(n10115), .dout(n10116));
  jand g09925(.dina(\a[53] ), .dinb(\a[19] ), .dout(n10117));
  jnot g09926(.din(n10117), .dout(n10118));
  jand g09927(.dina(n9559), .dinb(n4068), .dout(n10119));
  jnot g09928(.din(n10119), .dout(n10120));
  jand g09929(.dina(\a[39] ), .dinb(\a[33] ), .dout(n10121));
  jor  g09930(.dina(n10121), .dinb(n9828), .dout(n10122));
  jand g09931(.dina(n10122), .dinb(n10120), .dout(n10123));
  jxor g09932(.dina(n10123), .dinb(n10118), .dout(n10124));
  jxor g09933(.dina(n10124), .dinb(n10116), .dout(n10125));
  jxor g09934(.dina(n10125), .dinb(n10100), .dout(n10126));
  jxor g09935(.dina(n10126), .dinb(n10084), .dout(n10127));
  jxor g09936(.dina(n10127), .dinb(n10081), .dout(n10128));
  jxor g09937(.dina(n10128), .dinb(n10019), .dout(n10129));
  jxor g09938(.dina(n10129), .dinb(n9973), .dout(n10130));
  jnot g09939(.din(n10130), .dout(n10131));
  jand g09940(.dina(n9754), .dinb(n9751), .dout(n10132));
  jand g09941(.dina(n9929), .dinb(n9755), .dout(n10133));
  jor  g09942(.dina(n10133), .dinb(n10132), .dout(n10134));
  jxor g09943(.dina(n10134), .dinb(n10131), .dout(n10135));
  jand g09944(.dina(n9930), .dinb(n9721), .dout(n10136));
  jnot g09945(.din(n10136), .dout(n10137));
  jnot g09946(.din(n9930), .dout(n10138));
  jand g09947(.dina(n10138), .dinb(n9722), .dout(n10139));
  jor  g09948(.dina(n9937), .dinb(n10139), .dout(n10140));
  jand g09949(.dina(n10140), .dinb(n10137), .dout(n10141));
  jxor g09950(.dina(n10141), .dinb(n10135), .dout(\asquared[73] ));
  jand g09951(.dina(n9972), .dinb(n9969), .dout(n10143));
  jand g09952(.dina(n10129), .dinb(n9973), .dout(n10144));
  jor  g09953(.dina(n10144), .dinb(n10143), .dout(n10145));
  jand g09954(.dina(n10018), .dinb(n9976), .dout(n10146));
  jand g09955(.dina(n10128), .dinb(n10019), .dout(n10147));
  jor  g09956(.dina(n10147), .dinb(n10146), .dout(n10148));
  jand g09957(.dina(n10126), .dinb(n10084), .dout(n10149));
  jand g09958(.dina(n10127), .dinb(n10081), .dout(n10150));
  jor  g09959(.dina(n10150), .dinb(n10149), .dout(n10151));
  jand g09960(.dina(n9993), .dinb(n9990), .dout(n10152));
  jand g09961(.dina(n10017), .dinb(n9994), .dout(n10153));
  jor  g09962(.dina(n10153), .dinb(n10152), .dout(n10154));
  jor  g09963(.dina(n10099), .dinb(n10095), .dout(n10155));
  jand g09964(.dina(n10125), .dinb(n10100), .dout(n10156));
  jnot g09965(.din(n10156), .dout(n10157));
  jand g09966(.dina(n10157), .dinb(n10155), .dout(n10158));
  jnot g09967(.din(n10158), .dout(n10159));
  jand g09968(.dina(n10003), .dinb(n10001), .dout(n10160));
  jand g09969(.dina(n10007), .dinb(n10004), .dout(n10161));
  jor  g09970(.dina(n10161), .dinb(n10160), .dout(n10162));
  jand g09971(.dina(n10089), .dinb(n10086), .dout(n10163));
  jand g09972(.dina(n10093), .dinb(n10090), .dout(n10164));
  jor  g09973(.dina(n10164), .dinb(n10163), .dout(n10165));
  jnot g09974(.din(n10165), .dout(n10166));
  jand g09975(.dina(\a[42] ), .dinb(\a[31] ), .dout(n10167));
  jnot g09976(.din(n10167), .dout(n10168));
  jand g09977(.dina(n4632), .dinb(n2671), .dout(n10169));
  jnot g09978(.din(n10169), .dout(n10170));
  jand g09979(.dina(\a[40] ), .dinb(\a[33] ), .dout(n10171));
  jand g09980(.dina(\a[41] ), .dinb(\a[32] ), .dout(n10172));
  jor  g09981(.dina(n10172), .dinb(n10171), .dout(n10173));
  jand g09982(.dina(n10173), .dinb(n10170), .dout(n10174));
  jxor g09983(.dina(n10174), .dinb(n10168), .dout(n10175));
  jxor g09984(.dina(n10175), .dinb(n10166), .dout(n10176));
  jxor g09985(.dina(n10176), .dinb(n10162), .dout(n10177));
  jand g09986(.dina(n10015), .dinb(n10008), .dout(n10178));
  jand g09987(.dina(n10016), .dinb(n9999), .dout(n10179));
  jor  g09988(.dina(n10179), .dinb(n10178), .dout(n10180));
  jxor g09989(.dina(n10180), .dinb(n10177), .dout(n10181));
  jxor g09990(.dina(n10181), .dinb(n10159), .dout(n10182));
  jxor g09991(.dina(n10182), .dinb(n10154), .dout(n10183));
  jxor g09992(.dina(n10183), .dinb(n10151), .dout(n10184));
  jxor g09993(.dina(n10184), .dinb(n10148), .dout(n10185));
  jand g09994(.dina(n9967), .dinb(n9964), .dout(n10186));
  jand g09995(.dina(n9968), .dinb(n9941), .dout(n10187));
  jor  g09996(.dina(n10187), .dinb(n10186), .dout(n10188));
  jand g09997(.dina(n10036), .dinb(n10026), .dout(n10189));
  jand g09998(.dina(n10045), .dinb(n10037), .dout(n10190));
  jor  g09999(.dina(n10190), .dinb(n10189), .dout(n10191));
  jand g10000(.dina(n10010), .dinb(n9833), .dout(n10192));
  jand g10001(.dina(n10014), .dinb(n10011), .dout(n10193));
  jor  g10002(.dina(n10193), .dinb(n10192), .dout(n10194));
  jxor g10003(.dina(n10194), .dinb(n10191), .dout(n10195));
  jnot g10004(.din(n10195), .dout(n10196));
  jand g10005(.dina(n10114), .dinb(n10107), .dout(n10197));
  jnot g10006(.din(n10197), .dout(n10198));
  jor  g10007(.dina(n10124), .dinb(n10116), .dout(n10199));
  jand g10008(.dina(n10199), .dinb(n10198), .dout(n10200));
  jxor g10009(.dina(n10200), .dinb(n10196), .dout(n10201));
  jand g10010(.dina(n10079), .dinb(n10046), .dout(n10202));
  jand g10011(.dina(n10080), .dinb(n10024), .dout(n10203));
  jor  g10012(.dina(n10203), .dinb(n10202), .dout(n10204));
  jxor g10013(.dina(n10204), .dinb(n10201), .dout(n10205));
  jor  g10014(.dina(n10077), .dinb(n10068), .dout(n10206));
  jand g10015(.dina(n10078), .dinb(n10063), .dout(n10207));
  jnot g10016(.din(n10207), .dout(n10208));
  jand g10017(.dina(n10208), .dinb(n10206), .dout(n10209));
  jnot g10018(.din(n10209), .dout(n10210));
  jand g10019(.dina(\a[60] ), .dinb(\a[13] ), .dout(n10211));
  jand g10020(.dina(n10072), .dinb(n10070), .dout(n10212));
  jnot g10021(.din(n10212), .dout(n10213));
  jand g10022(.dina(n10213), .dinb(n10075), .dout(n10214));
  jxor g10023(.dina(n10214), .dinb(n10211), .dout(n10215));
  jand g10024(.dina(n10120), .dinb(n10118), .dout(n10216));
  jnot g10025(.din(n10216), .dout(n10217));
  jand g10026(.dina(n10217), .dinb(n10122), .dout(n10218));
  jxor g10027(.dina(n10218), .dinb(n10215), .dout(n10219));
  jand g10028(.dina(n10044), .dinb(n10038), .dout(n10220));
  jor  g10029(.dina(n10220), .dinb(n10039), .dout(n10221));
  jand g10030(.dina(n10030), .dinb(n10028), .dout(n10222));
  jnot g10031(.din(n10222), .dout(n10223));
  jand g10032(.dina(n10223), .dinb(n10033), .dout(n10224));
  jxor g10033(.dina(n10224), .dinb(n10221), .dout(n10225));
  jxor g10034(.dina(n10225), .dinb(n10060), .dout(n10226));
  jxor g10035(.dina(n10226), .dinb(n10219), .dout(n10227));
  jxor g10036(.dina(n10227), .dinb(n10210), .dout(n10228));
  jxor g10037(.dina(n10228), .dinb(n10205), .dout(n10229));
  jxor g10038(.dina(n10229), .dinb(n10188), .dout(n10230));
  jand g10039(.dina(n9984), .dinb(n9981), .dout(n10231));
  jnot g10040(.din(n10231), .dout(n10232));
  jor  g10041(.dina(n9989), .dinb(n9986), .dout(n10233));
  jand g10042(.dina(n10233), .dinb(n10232), .dout(n10234));
  jnot g10043(.din(n10234), .dout(n10235));
  jand g10044(.dina(\a[50] ), .dinb(\a[23] ), .dout(n10236));
  jand g10045(.dina(\a[62] ), .dinb(\a[11] ), .dout(n10237));
  jor  g10046(.dina(n10237), .dinb(\a[37] ), .dout(n10238));
  jand g10047(.dina(n4649), .dinb(\a[62] ), .dout(n10239));
  jnot g10048(.din(n10239), .dout(n10240));
  jand g10049(.dina(n10240), .dinb(n10238), .dout(n10241));
  jxor g10050(.dina(n10241), .dinb(n10236), .dout(n10242));
  jnot g10051(.din(n10242), .dout(n10243));
  jnot g10052(.din(n10051), .dout(n10244));
  jand g10053(.dina(\a[54] ), .dinb(\a[49] ), .dout(n10245));
  jand g10054(.dina(n10245), .dinb(n3746), .dout(n10246));
  jnot g10055(.din(n10246), .dout(n10247));
  jand g10056(.dina(\a[54] ), .dinb(\a[19] ), .dout(n10248));
  jand g10057(.dina(\a[49] ), .dinb(\a[24] ), .dout(n10249));
  jor  g10058(.dina(n10249), .dinb(n10248), .dout(n10250));
  jand g10059(.dina(n10250), .dinb(n10247), .dout(n10251));
  jxor g10060(.dina(n10251), .dinb(n10244), .dout(n10252));
  jxor g10061(.dina(n10252), .dinb(n10243), .dout(n10253));
  jand g10062(.dina(\a[51] ), .dinb(\a[22] ), .dout(n10254));
  jand g10063(.dina(n7165), .dinb(n1490), .dout(n10255));
  jnot g10064(.din(n10255), .dout(n10256));
  jand g10065(.dina(\a[53] ), .dinb(\a[20] ), .dout(n10257));
  jand g10066(.dina(\a[52] ), .dinb(\a[21] ), .dout(n10258));
  jor  g10067(.dina(n10258), .dinb(n10257), .dout(n10259));
  jand g10068(.dina(n10259), .dinb(n10256), .dout(n10260));
  jxor g10069(.dina(n10260), .dinb(n10254), .dout(n10261));
  jxor g10070(.dina(n10261), .dinb(n10253), .dout(n10262));
  jand g10071(.dina(n10065), .dinb(n9906), .dout(n10263));
  jand g10072(.dina(n10066), .dinb(n10064), .dout(n10264));
  jor  g10073(.dina(n10264), .dinb(n10263), .dout(n10265));
  jand g10074(.dina(\a[56] ), .dinb(\a[17] ), .dout(n10266));
  jand g10075(.dina(\a[47] ), .dinb(\a[27] ), .dout(n10267));
  jand g10076(.dina(n10267), .dinb(n9916), .dout(n10268));
  jnot g10077(.din(n10268), .dout(n10269));
  jand g10078(.dina(\a[47] ), .dinb(\a[26] ), .dout(n10270));
  jand g10079(.dina(\a[46] ), .dinb(\a[27] ), .dout(n10271));
  jor  g10080(.dina(n10271), .dinb(n10270), .dout(n10272));
  jand g10081(.dina(n10272), .dinb(n10269), .dout(n10273));
  jxor g10082(.dina(n10273), .dinb(n10266), .dout(n10274));
  jxor g10083(.dina(n10274), .dinb(n10265), .dout(n10275));
  jand g10084(.dina(\a[59] ), .dinb(\a[14] ), .dout(n10276));
  jand g10085(.dina(\a[58] ), .dinb(\a[15] ), .dout(n10277));
  jand g10086(.dina(\a[57] ), .dinb(\a[16] ), .dout(n10278));
  jor  g10087(.dina(n10278), .dinb(n10277), .dout(n10279));
  jand g10088(.dina(n7519), .dinb(n829), .dout(n10280));
  jnot g10089(.din(n10280), .dout(n10281));
  jand g10090(.dina(n10281), .dinb(n10279), .dout(n10282));
  jxor g10091(.dina(n10282), .dinb(n10276), .dout(n10283));
  jxor g10092(.dina(n10283), .dinb(n10275), .dout(n10284));
  jxor g10093(.dina(n10284), .dinb(n10262), .dout(n10285));
  jxor g10094(.dina(n10285), .dinb(n10235), .dout(n10286));
  jand g10095(.dina(n9959), .dinb(n9944), .dout(n10287));
  jand g10096(.dina(n9963), .dinb(n9960), .dout(n10288));
  jor  g10097(.dina(n10288), .dinb(n10287), .dout(n10289));
  jand g10098(.dina(n9955), .dinb(n9951), .dout(n10290));
  jor  g10099(.dina(n10290), .dinb(n9952), .dout(n10291));
  jand g10100(.dina(n10106), .dinb(n9894), .dout(n10292));
  jor  g10101(.dina(n10292), .dinb(n10101), .dout(n10293));
  jor  g10102(.dina(n10108), .dinb(n9916), .dout(n10294));
  jand g10103(.dina(n10294), .dinb(n10112), .dout(n10295));
  jxor g10104(.dina(n10295), .dinb(n10293), .dout(n10296));
  jxor g10105(.dina(n10296), .dinb(n10291), .dout(n10297));
  jand g10106(.dina(n9957), .dinb(n9950), .dout(n10298));
  jand g10107(.dina(n9958), .dinb(n9947), .dout(n10299));
  jor  g10108(.dina(n10299), .dinb(n10298), .dout(n10300));
  jxor g10109(.dina(n10300), .dinb(n10297), .dout(n10301));
  jand g10110(.dina(n10069), .dinb(n4528), .dout(n10302));
  jnot g10111(.din(n10302), .dout(n10303));
  jand g10112(.dina(n4068), .dinb(n3138), .dout(n10304));
  jand g10113(.dina(\a[39] ), .dinb(\a[35] ), .dout(n10305));
  jand g10114(.dina(n10305), .dinb(n9828), .dout(n10306));
  jor  g10115(.dina(n10306), .dinb(n10304), .dout(n10307));
  jand g10116(.dina(n10307), .dinb(n10303), .dout(n10308));
  jnot g10117(.din(n10308), .dout(n10309));
  jand g10118(.dina(n10309), .dinb(n4068), .dout(n10310));
  jor  g10119(.dina(n10307), .dinb(n10302), .dout(n10311));
  jnot g10120(.din(n10311), .dout(n10312));
  jand g10121(.dina(\a[38] ), .dinb(\a[35] ), .dout(n10313));
  jor  g10122(.dina(n10313), .dinb(n3138), .dout(n10314));
  jand g10123(.dina(n10314), .dinb(n10312), .dout(n10315));
  jor  g10124(.dina(n10315), .dinb(n10310), .dout(n10316));
  jand g10125(.dina(\a[48] ), .dinb(\a[25] ), .dout(n10317));
  jand g10126(.dina(\a[63] ), .dinb(\a[10] ), .dout(n10318));
  jand g10127(.dina(\a[61] ), .dinb(\a[12] ), .dout(n10319));
  jor  g10128(.dina(n10319), .dinb(n10318), .dout(n10320));
  jand g10129(.dina(n8387), .dinb(n1151), .dout(n10321));
  jnot g10130(.din(n10321), .dout(n10322));
  jand g10131(.dina(n10322), .dinb(n10320), .dout(n10323));
  jxor g10132(.dina(n10323), .dinb(n10317), .dout(n10324));
  jand g10133(.dina(\a[45] ), .dinb(\a[28] ), .dout(n10325));
  jand g10134(.dina(n4495), .dinb(n3294), .dout(n10326));
  jnot g10135(.din(n10326), .dout(n10327));
  jand g10136(.dina(\a[44] ), .dinb(\a[29] ), .dout(n10328));
  jand g10137(.dina(\a[43] ), .dinb(\a[30] ), .dout(n10329));
  jor  g10138(.dina(n10329), .dinb(n10328), .dout(n10330));
  jand g10139(.dina(n10330), .dinb(n10327), .dout(n10331));
  jxor g10140(.dina(n10331), .dinb(n10325), .dout(n10332));
  jxor g10141(.dina(n10332), .dinb(n10324), .dout(n10333));
  jxor g10142(.dina(n10333), .dinb(n10316), .dout(n10334));
  jxor g10143(.dina(n10334), .dinb(n10301), .dout(n10335));
  jxor g10144(.dina(n10335), .dinb(n10289), .dout(n10336));
  jxor g10145(.dina(n10336), .dinb(n10286), .dout(n10337));
  jxor g10146(.dina(n10337), .dinb(n10230), .dout(n10338));
  jxor g10147(.dina(n10338), .dinb(n10185), .dout(n10339));
  jnot g10148(.din(n10339), .dout(n10340));
  jxor g10149(.dina(n10340), .dinb(n10145), .dout(n10341));
  jand g10150(.dina(n10134), .dinb(n10130), .dout(n10342));
  jnot g10151(.din(n10342), .dout(n10343));
  jnot g10152(.din(n10134), .dout(n10344));
  jand g10153(.dina(n10344), .dinb(n10131), .dout(n10345));
  jor  g10154(.dina(n10141), .dinb(n10345), .dout(n10346));
  jand g10155(.dina(n10346), .dinb(n10343), .dout(n10347));
  jxor g10156(.dina(n10347), .dinb(n10341), .dout(\asquared[74] ));
  jand g10157(.dina(n10184), .dinb(n10148), .dout(n10349));
  jand g10158(.dina(n10338), .dinb(n10185), .dout(n10350));
  jor  g10159(.dina(n10350), .dinb(n10349), .dout(n10351));
  jand g10160(.dina(n10229), .dinb(n10188), .dout(n10352));
  jand g10161(.dina(n10337), .dinb(n10230), .dout(n10353));
  jor  g10162(.dina(n10353), .dinb(n10352), .dout(n10354));
  jand g10163(.dina(n10335), .dinb(n10289), .dout(n10355));
  jand g10164(.dina(n10336), .dinb(n10286), .dout(n10356));
  jor  g10165(.dina(n10356), .dinb(n10355), .dout(n10357));
  jand g10166(.dina(n10204), .dinb(n10201), .dout(n10358));
  jand g10167(.dina(n10228), .dinb(n10205), .dout(n10359));
  jor  g10168(.dina(n10359), .dinb(n10358), .dout(n10360));
  jand g10169(.dina(n10224), .dinb(n10221), .dout(n10361));
  jand g10170(.dina(n10225), .dinb(n10060), .dout(n10362));
  jor  g10171(.dina(n10362), .dinb(n10361), .dout(n10363));
  jand g10172(.dina(n10214), .dinb(n10211), .dout(n10364));
  jand g10173(.dina(n10218), .dinb(n10215), .dout(n10365));
  jor  g10174(.dina(n10365), .dinb(n10364), .dout(n10366));
  jxor g10175(.dina(n10366), .dinb(n10363), .dout(n10367));
  jand g10176(.dina(n10274), .dinb(n10265), .dout(n10368));
  jand g10177(.dina(n10283), .dinb(n10275), .dout(n10369));
  jor  g10178(.dina(n10369), .dinb(n10368), .dout(n10370));
  jxor g10179(.dina(n10370), .dinb(n10367), .dout(n10371));
  jand g10180(.dina(n10226), .dinb(n10219), .dout(n10372));
  jand g10181(.dina(n10227), .dinb(n10210), .dout(n10373));
  jor  g10182(.dina(n10373), .dinb(n10372), .dout(n10374));
  jnot g10183(.din(n10374), .dout(n10375));
  jand g10184(.dina(n10194), .dinb(n10191), .dout(n10376));
  jnot g10185(.din(n10376), .dout(n10377));
  jor  g10186(.dina(n10200), .dinb(n10196), .dout(n10378));
  jand g10187(.dina(n10378), .dinb(n10377), .dout(n10379));
  jxor g10188(.dina(n10379), .dinb(n10375), .dout(n10380));
  jxor g10189(.dina(n10380), .dinb(n10371), .dout(n10381));
  jxor g10190(.dina(n10381), .dinb(n10360), .dout(n10382));
  jxor g10191(.dina(n10382), .dinb(n10357), .dout(n10383));
  jxor g10192(.dina(n10383), .dinb(n10354), .dout(n10384));
  jand g10193(.dina(n10182), .dinb(n10154), .dout(n10385));
  jand g10194(.dina(n10183), .dinb(n10151), .dout(n10386));
  jor  g10195(.dina(n10386), .dinb(n10385), .dout(n10387));
  jor  g10196(.dina(n10252), .dinb(n10243), .dout(n10388));
  jand g10197(.dina(n10261), .dinb(n10253), .dout(n10389));
  jnot g10198(.din(n10389), .dout(n10390));
  jand g10199(.dina(n10390), .dinb(n10388), .dout(n10391));
  jnot g10200(.din(n10391), .dout(n10392));
  jand g10201(.dina(n10170), .dinb(n10168), .dout(n10393));
  jnot g10202(.din(n10393), .dout(n10394));
  jand g10203(.dina(n10394), .dinb(n10173), .dout(n10395));
  jxor g10204(.dina(n10395), .dinb(n10311), .dout(n10396));
  jand g10205(.dina(\a[60] ), .dinb(\a[14] ), .dout(n10397));
  jnot g10206(.din(n10397), .dout(n10398));
  jand g10207(.dina(\a[59] ), .dinb(\a[16] ), .dout(n10399));
  jand g10208(.dina(n10399), .dinb(n10277), .dout(n10400));
  jnot g10209(.din(n10400), .dout(n10401));
  jand g10210(.dina(\a[59] ), .dinb(\a[15] ), .dout(n10402));
  jand g10211(.dina(\a[58] ), .dinb(\a[16] ), .dout(n10403));
  jor  g10212(.dina(n10403), .dinb(n10402), .dout(n10404));
  jand g10213(.dina(n10404), .dinb(n10401), .dout(n10405));
  jxor g10214(.dina(n10405), .dinb(n10398), .dout(n10406));
  jnot g10215(.din(n10406), .dout(n10407));
  jxor g10216(.dina(n10407), .dinb(n10396), .dout(n10408));
  jxor g10217(.dina(n10408), .dinb(n10392), .dout(n10409));
  jnot g10218(.din(n10409), .dout(n10410));
  jor  g10219(.dina(n10175), .dinb(n10166), .dout(n10411));
  jand g10220(.dina(n10176), .dinb(n10162), .dout(n10412));
  jnot g10221(.din(n10412), .dout(n10413));
  jand g10222(.dina(n10413), .dinb(n10411), .dout(n10414));
  jxor g10223(.dina(n10414), .dinb(n10410), .dout(n10415));
  jand g10224(.dina(n10284), .dinb(n10262), .dout(n10416));
  jand g10225(.dina(n10285), .dinb(n10235), .dout(n10417));
  jor  g10226(.dina(n10417), .dinb(n10416), .dout(n10418));
  jand g10227(.dina(n10300), .dinb(n10297), .dout(n10419));
  jand g10228(.dina(n10334), .dinb(n10301), .dout(n10420));
  jor  g10229(.dina(n10420), .dinb(n10419), .dout(n10421));
  jxor g10230(.dina(n10421), .dinb(n10418), .dout(n10422));
  jxor g10231(.dina(n10422), .dinb(n10415), .dout(n10423));
  jxor g10232(.dina(n10423), .dinb(n10387), .dout(n10424));
  jand g10233(.dina(n10180), .dinb(n10177), .dout(n10425));
  jand g10234(.dina(n10181), .dinb(n10159), .dout(n10426));
  jor  g10235(.dina(n10426), .dinb(n10425), .dout(n10427));
  jand g10236(.dina(n10282), .dinb(n10276), .dout(n10428));
  jor  g10237(.dina(n10428), .dinb(n10280), .dout(n10429));
  jand g10238(.dina(n10272), .dinb(n10266), .dout(n10430));
  jor  g10239(.dina(n10430), .dinb(n10268), .dout(n10431));
  jor  g10240(.dina(n10326), .dinb(n10325), .dout(n10432));
  jand g10241(.dina(n10432), .dinb(n10330), .dout(n10433));
  jxor g10242(.dina(n10433), .dinb(n10431), .dout(n10434));
  jxor g10243(.dina(n10434), .dinb(n10429), .dout(n10435));
  jand g10244(.dina(n10323), .dinb(n10317), .dout(n10436));
  jor  g10245(.dina(n10436), .dinb(n10321), .dout(n10437));
  jand g10246(.dina(n10259), .dinb(n10254), .dout(n10438));
  jor  g10247(.dina(n10438), .dinb(n10255), .dout(n10439));
  jand g10248(.dina(n10247), .dinb(n10244), .dout(n10440));
  jnot g10249(.din(n10440), .dout(n10441));
  jand g10250(.dina(n10441), .dinb(n10250), .dout(n10442));
  jxor g10251(.dina(n10442), .dinb(n10439), .dout(n10443));
  jxor g10252(.dina(n10443), .dinb(n10437), .dout(n10444));
  jand g10253(.dina(n10332), .dinb(n10324), .dout(n10445));
  jand g10254(.dina(n10333), .dinb(n10316), .dout(n10446));
  jor  g10255(.dina(n10446), .dinb(n10445), .dout(n10447));
  jxor g10256(.dina(n10447), .dinb(n10444), .dout(n10448));
  jxor g10257(.dina(n10448), .dinb(n10435), .dout(n10449));
  jxor g10258(.dina(n10449), .dinb(n10427), .dout(n10450));
  jand g10259(.dina(n10295), .dinb(n10293), .dout(n10451));
  jand g10260(.dina(n10296), .dinb(n10291), .dout(n10452));
  jor  g10261(.dina(n10452), .dinb(n10451), .dout(n10453));
  jand g10262(.dina(\a[45] ), .dinb(\a[29] ), .dout(n10454));
  jand g10263(.dina(\a[44] ), .dinb(\a[30] ), .dout(n10455));
  jand g10264(.dina(\a[57] ), .dinb(\a[17] ), .dout(n10456));
  jand g10265(.dina(n10456), .dinb(n10455), .dout(n10457));
  jnot g10266(.din(n10457), .dout(n10458));
  jand g10267(.dina(n4812), .dinb(n3294), .dout(n10459));
  jand g10268(.dina(n10456), .dinb(n10454), .dout(n10460));
  jor  g10269(.dina(n10460), .dinb(n10459), .dout(n10461));
  jand g10270(.dina(n10461), .dinb(n10458), .dout(n10462));
  jnot g10271(.din(n10462), .dout(n10463));
  jand g10272(.dina(n10463), .dinb(n10454), .dout(n10464));
  jor  g10273(.dina(n10461), .dinb(n10457), .dout(n10465));
  jnot g10274(.din(n10465), .dout(n10466));
  jor  g10275(.dina(n10456), .dinb(n10455), .dout(n10467));
  jand g10276(.dina(n10467), .dinb(n10466), .dout(n10468));
  jor  g10277(.dina(n10468), .dinb(n10464), .dout(n10469));
  jand g10278(.dina(n10241), .dinb(n10236), .dout(n10470));
  jor  g10279(.dina(n10470), .dinb(n10239), .dout(n10471));
  jand g10280(.dina(n8702), .dinb(n899), .dout(n10472));
  jnot g10281(.din(n10472), .dout(n10473));
  jand g10282(.dina(\a[62] ), .dinb(\a[12] ), .dout(n10474));
  jand g10283(.dina(\a[61] ), .dinb(\a[13] ), .dout(n10475));
  jor  g10284(.dina(n10475), .dinb(n10474), .dout(n10476));
  jand g10285(.dina(n10476), .dinb(n10473), .dout(n10477));
  jxor g10286(.dina(n10477), .dinb(n10471), .dout(n10478));
  jxor g10287(.dina(n10478), .dinb(n10469), .dout(n10479));
  jxor g10288(.dina(n10479), .dinb(n10453), .dout(n10480));
  jand g10289(.dina(\a[63] ), .dinb(\a[11] ), .dout(n10481));
  jand g10290(.dina(\a[43] ), .dinb(\a[31] ), .dout(n10482));
  jand g10291(.dina(\a[42] ), .dinb(\a[32] ), .dout(n10483));
  jor  g10292(.dina(n10483), .dinb(n10482), .dout(n10484));
  jand g10293(.dina(n4317), .dinb(n3269), .dout(n10485));
  jnot g10294(.din(n10485), .dout(n10486));
  jand g10295(.dina(n10486), .dinb(n10484), .dout(n10487));
  jxor g10296(.dina(n10487), .dinb(n10481), .dout(n10488));
  jand g10297(.dina(\a[56] ), .dinb(\a[18] ), .dout(n10489));
  jand g10298(.dina(\a[49] ), .dinb(\a[25] ), .dout(n10490));
  jxor g10299(.dina(n10490), .dinb(n10489), .dout(n10491));
  jxor g10300(.dina(n10491), .dinb(n4511), .dout(n10492));
  jxor g10301(.dina(n10492), .dinb(n10488), .dout(n10493));
  jnot g10302(.din(n10493), .dout(n10494));
  jand g10303(.dina(\a[48] ), .dinb(\a[26] ), .dout(n10495));
  jnot g10304(.din(n10495), .dout(n10496));
  jand g10305(.dina(\a[47] ), .dinb(\a[28] ), .dout(n10497));
  jand g10306(.dina(n10497), .dinb(n10271), .dout(n10498));
  jnot g10307(.din(n10498), .dout(n10499));
  jand g10308(.dina(\a[46] ), .dinb(\a[28] ), .dout(n10500));
  jor  g10309(.dina(n10500), .dinb(n10267), .dout(n10501));
  jand g10310(.dina(n10501), .dinb(n10499), .dout(n10502));
  jxor g10311(.dina(n10502), .dinb(n10496), .dout(n10503));
  jxor g10312(.dina(n10503), .dinb(n10494), .dout(n10504));
  jand g10313(.dina(\a[52] ), .dinb(\a[22] ), .dout(n10505));
  jand g10314(.dina(\a[55] ), .dinb(\a[19] ), .dout(n10506));
  jand g10315(.dina(\a[53] ), .dinb(\a[21] ), .dout(n10507));
  jor  g10316(.dina(n10507), .dinb(n10506), .dout(n10508));
  jand g10317(.dina(n6498), .dinb(n3334), .dout(n10509));
  jnot g10318(.din(n10509), .dout(n10510));
  jand g10319(.dina(n10510), .dinb(n10508), .dout(n10511));
  jxor g10320(.dina(n10511), .dinb(n10505), .dout(n10512));
  jnot g10321(.din(n10512), .dout(n10513));
  jand g10322(.dina(\a[54] ), .dinb(\a[20] ), .dout(n10514));
  jnot g10323(.din(n10514), .dout(n10515));
  jand g10324(.dina(n3665), .dinb(n2845), .dout(n10516));
  jnot g10325(.din(n10516), .dout(n10517));
  jand g10326(.dina(\a[40] ), .dinb(\a[34] ), .dout(n10518));
  jor  g10327(.dina(n10518), .dinb(n10305), .dout(n10519));
  jand g10328(.dina(n10519), .dinb(n10517), .dout(n10520));
  jxor g10329(.dina(n10520), .dinb(n10515), .dout(n10521));
  jxor g10330(.dina(n10521), .dinb(n10513), .dout(n10522));
  jnot g10331(.din(n10522), .dout(n10523));
  jnot g10332(.din(n4528), .dout(n10524));
  jand g10333(.dina(n5594), .dinb(n1942), .dout(n10525));
  jnot g10334(.din(n10525), .dout(n10526));
  jand g10335(.dina(\a[51] ), .dinb(\a[23] ), .dout(n10527));
  jand g10336(.dina(\a[50] ), .dinb(\a[24] ), .dout(n10528));
  jor  g10337(.dina(n10528), .dinb(n10527), .dout(n10529));
  jand g10338(.dina(n10529), .dinb(n10526), .dout(n10530));
  jxor g10339(.dina(n10530), .dinb(n10524), .dout(n10531));
  jxor g10340(.dina(n10531), .dinb(n10523), .dout(n10532));
  jxor g10341(.dina(n10532), .dinb(n10504), .dout(n10533));
  jxor g10342(.dina(n10533), .dinb(n10480), .dout(n10534));
  jxor g10343(.dina(n10534), .dinb(n10450), .dout(n10535));
  jxor g10344(.dina(n10535), .dinb(n10424), .dout(n10536));
  jxor g10345(.dina(n10536), .dinb(n10384), .dout(n10537));
  jnot g10346(.din(n10537), .dout(n10538));
  jxor g10347(.dina(n10538), .dinb(n10351), .dout(n10539));
  jand g10348(.dina(n10339), .dinb(n10145), .dout(n10540));
  jnot g10349(.din(n10540), .dout(n10541));
  jnot g10350(.din(n10145), .dout(n10542));
  jand g10351(.dina(n10340), .dinb(n10542), .dout(n10543));
  jor  g10352(.dina(n10347), .dinb(n10543), .dout(n10544));
  jand g10353(.dina(n10544), .dinb(n10541), .dout(n10545));
  jxor g10354(.dina(n10545), .dinb(n10539), .dout(\asquared[75] ));
  jand g10355(.dina(n10383), .dinb(n10354), .dout(n10547));
  jand g10356(.dina(n10536), .dinb(n10384), .dout(n10548));
  jor  g10357(.dina(n10548), .dinb(n10547), .dout(n10549));
  jand g10358(.dina(n10381), .dinb(n10360), .dout(n10550));
  jand g10359(.dina(n10382), .dinb(n10357), .dout(n10551));
  jor  g10360(.dina(n10551), .dinb(n10550), .dout(n10552));
  jand g10361(.dina(n10395), .dinb(n10311), .dout(n10553));
  jand g10362(.dina(n10407), .dinb(n10396), .dout(n10554));
  jor  g10363(.dina(n10554), .dinb(n10553), .dout(n10555));
  jand g10364(.dina(n10442), .dinb(n10439), .dout(n10556));
  jand g10365(.dina(n10443), .dinb(n10437), .dout(n10557));
  jor  g10366(.dina(n10557), .dinb(n10556), .dout(n10558));
  jxor g10367(.dina(n10558), .dinb(n10555), .dout(n10559));
  jand g10368(.dina(n10433), .dinb(n10431), .dout(n10560));
  jand g10369(.dina(n10434), .dinb(n10429), .dout(n10561));
  jor  g10370(.dina(n10561), .dinb(n10560), .dout(n10562));
  jxor g10371(.dina(n10562), .dinb(n10559), .dout(n10563));
  jand g10372(.dina(n10532), .dinb(n10504), .dout(n10564));
  jand g10373(.dina(n10533), .dinb(n10480), .dout(n10565));
  jor  g10374(.dina(n10565), .dinb(n10564), .dout(n10566));
  jxor g10375(.dina(n10566), .dinb(n10563), .dout(n10567));
  jand g10376(.dina(n10478), .dinb(n10469), .dout(n10568));
  jand g10377(.dina(n10479), .dinb(n10453), .dout(n10569));
  jor  g10378(.dina(n10569), .dinb(n10568), .dout(n10570));
  jand g10379(.dina(n10511), .dinb(n10505), .dout(n10571));
  jor  g10380(.dina(n10571), .dinb(n10509), .dout(n10572));
  jand g10381(.dina(n10526), .dinb(n10524), .dout(n10573));
  jnot g10382(.din(n10573), .dout(n10574));
  jand g10383(.dina(n10574), .dinb(n10529), .dout(n10575));
  jand g10384(.dina(n10517), .dinb(n10515), .dout(n10576));
  jnot g10385(.din(n10576), .dout(n10577));
  jand g10386(.dina(n10577), .dinb(n10519), .dout(n10578));
  jxor g10387(.dina(n10578), .dinb(n10575), .dout(n10579));
  jxor g10388(.dina(n10579), .dinb(n10572), .dout(n10580));
  jand g10389(.dina(n10487), .dinb(n10481), .dout(n10581));
  jor  g10390(.dina(n10581), .dinb(n10485), .dout(n10582));
  jand g10391(.dina(n10490), .dinb(n10489), .dout(n10583));
  jand g10392(.dina(n10491), .dinb(n4511), .dout(n10584));
  jor  g10393(.dina(n10584), .dinb(n10583), .dout(n10585));
  jxor g10394(.dina(n10585), .dinb(n10582), .dout(n10586));
  jand g10395(.dina(n10477), .dinb(n10471), .dout(n10587));
  jor  g10396(.dina(n10587), .dinb(n10472), .dout(n10588));
  jxor g10397(.dina(n10588), .dinb(n10586), .dout(n10589));
  jxor g10398(.dina(n10589), .dinb(n10580), .dout(n10590));
  jxor g10399(.dina(n10590), .dinb(n10570), .dout(n10591));
  jxor g10400(.dina(n10591), .dinb(n10567), .dout(n10592));
  jxor g10401(.dina(n10592), .dinb(n10552), .dout(n10593));
  jor  g10402(.dina(n10379), .dinb(n10375), .dout(n10594));
  jand g10403(.dina(n10380), .dinb(n10371), .dout(n10595));
  jnot g10404(.din(n10595), .dout(n10596));
  jand g10405(.dina(n10596), .dinb(n10594), .dout(n10597));
  jnot g10406(.din(n10597), .dout(n10598));
  jand g10407(.dina(n10499), .dinb(n10496), .dout(n10599));
  jnot g10408(.din(n10599), .dout(n10600));
  jand g10409(.dina(n10600), .dinb(n10501), .dout(n10601));
  jxor g10410(.dina(n10601), .dinb(n10465), .dout(n10602));
  jand g10411(.dina(n10401), .dinb(n10398), .dout(n10603));
  jnot g10412(.din(n10603), .dout(n10604));
  jand g10413(.dina(n10604), .dinb(n10404), .dout(n10605));
  jxor g10414(.dina(n10605), .dinb(n10602), .dout(n10606));
  jor  g10415(.dina(n10521), .dinb(n10513), .dout(n10607));
  jor  g10416(.dina(n10531), .dinb(n10523), .dout(n10608));
  jand g10417(.dina(n10608), .dinb(n10607), .dout(n10609));
  jand g10418(.dina(n10492), .dinb(n10488), .dout(n10610));
  jnot g10419(.din(n10610), .dout(n10611));
  jor  g10420(.dina(n10503), .dinb(n10494), .dout(n10612));
  jand g10421(.dina(n10612), .dinb(n10611), .dout(n10613));
  jxor g10422(.dina(n10613), .dinb(n10609), .dout(n10614));
  jxor g10423(.dina(n10614), .dinb(n10606), .dout(n10615));
  jxor g10424(.dina(n10615), .dinb(n10598), .dout(n10616));
  jand g10425(.dina(n10366), .dinb(n10363), .dout(n10617));
  jand g10426(.dina(n10370), .dinb(n10367), .dout(n10618));
  jor  g10427(.dina(n10618), .dinb(n10617), .dout(n10619));
  jand g10428(.dina(\a[45] ), .dinb(\a[30] ), .dout(n10620));
  jand g10429(.dina(\a[63] ), .dinb(\a[12] ), .dout(n10621));
  jand g10430(.dina(\a[56] ), .dinb(\a[19] ), .dout(n10622));
  jxor g10431(.dina(n10622), .dinb(n10621), .dout(n10623));
  jxor g10432(.dina(n10623), .dinb(n10620), .dout(n10624));
  jnot g10433(.din(n10624), .dout(n10625));
  jand g10434(.dina(\a[52] ), .dinb(\a[23] ), .dout(n10626));
  jnot g10435(.din(n10626), .dout(n10627));
  jand g10436(.dina(n3665), .dinb(n3243), .dout(n10628));
  jnot g10437(.din(n10628), .dout(n10629));
  jand g10438(.dina(\a[40] ), .dinb(\a[35] ), .dout(n10630));
  jand g10439(.dina(\a[39] ), .dinb(\a[36] ), .dout(n10631));
  jor  g10440(.dina(n10631), .dinb(n10630), .dout(n10632));
  jand g10441(.dina(n10632), .dinb(n10629), .dout(n10633));
  jxor g10442(.dina(n10633), .dinb(n10627), .dout(n10634));
  jxor g10443(.dina(n10634), .dinb(n10625), .dout(n10635));
  jnot g10444(.din(n10635), .dout(n10636));
  jand g10445(.dina(\a[62] ), .dinb(\a[13] ), .dout(n10637));
  jnot g10446(.din(n10637), .dout(n10638));
  jand g10447(.dina(\a[38] ), .dinb(n2837), .dout(n10639));
  jxor g10448(.dina(n10639), .dinb(n10638), .dout(n10640));
  jxor g10449(.dina(n10640), .dinb(n10636), .dout(n10641));
  jxor g10450(.dina(n10641), .dinb(n10619), .dout(n10642));
  jand g10451(.dina(\a[58] ), .dinb(\a[17] ), .dout(n10643));
  jand g10452(.dina(\a[57] ), .dinb(\a[49] ), .dout(n10644));
  jand g10453(.dina(n10644), .dinb(n3962), .dout(n10645));
  jnot g10454(.din(n10645), .dout(n10646));
  jand g10455(.dina(\a[49] ), .dinb(\a[26] ), .dout(n10647));
  jand g10456(.dina(n10647), .dinb(n10643), .dout(n10648));
  jand g10457(.dina(n7519), .dinb(n1107), .dout(n10649));
  jor  g10458(.dina(n10649), .dinb(n10648), .dout(n10650));
  jand g10459(.dina(n10650), .dinb(n10646), .dout(n10651));
  jnot g10460(.din(n10651), .dout(n10652));
  jand g10461(.dina(n10652), .dinb(n10643), .dout(n10653));
  jor  g10462(.dina(n10650), .dinb(n10645), .dout(n10654));
  jnot g10463(.din(n10654), .dout(n10655));
  jand g10464(.dina(\a[57] ), .dinb(\a[18] ), .dout(n10656));
  jor  g10465(.dina(n10656), .dinb(n10647), .dout(n10657));
  jand g10466(.dina(n10657), .dinb(n10655), .dout(n10658));
  jor  g10467(.dina(n10658), .dinb(n10653), .dout(n10659));
  jand g10468(.dina(\a[61] ), .dinb(\a[14] ), .dout(n10660));
  jand g10469(.dina(\a[60] ), .dinb(\a[16] ), .dout(n10661));
  jand g10470(.dina(n10661), .dinb(n10402), .dout(n10662));
  jnot g10471(.din(n10662), .dout(n10663));
  jand g10472(.dina(\a[60] ), .dinb(\a[15] ), .dout(n10664));
  jor  g10473(.dina(n10664), .dinb(n10399), .dout(n10665));
  jand g10474(.dina(n10665), .dinb(n10663), .dout(n10666));
  jxor g10475(.dina(n10666), .dinb(n10660), .dout(n10667));
  jxor g10476(.dina(n10667), .dinb(n10659), .dout(n10668));
  jnot g10477(.din(n10668), .dout(n10669));
  jand g10478(.dina(\a[48] ), .dinb(\a[27] ), .dout(n10670));
  jnot g10479(.din(n10670), .dout(n10671));
  jand g10480(.dina(\a[47] ), .dinb(\a[29] ), .dout(n10672));
  jand g10481(.dina(n10672), .dinb(n10500), .dout(n10673));
  jnot g10482(.din(n10673), .dout(n10674));
  jand g10483(.dina(\a[46] ), .dinb(\a[29] ), .dout(n10675));
  jor  g10484(.dina(n10675), .dinb(n10497), .dout(n10676));
  jand g10485(.dina(n10676), .dinb(n10674), .dout(n10677));
  jxor g10486(.dina(n10677), .dinb(n10671), .dout(n10678));
  jxor g10487(.dina(n10678), .dinb(n10669), .dout(n10679));
  jxor g10488(.dina(n10679), .dinb(n10642), .dout(n10680));
  jxor g10489(.dina(n10680), .dinb(n10616), .dout(n10681));
  jxor g10490(.dina(n10681), .dinb(n10593), .dout(n10682));
  jand g10491(.dina(n10449), .dinb(n10427), .dout(n10683));
  jand g10492(.dina(n10534), .dinb(n10450), .dout(n10684));
  jor  g10493(.dina(n10684), .dinb(n10683), .dout(n10685));
  jand g10494(.dina(n10421), .dinb(n10418), .dout(n10686));
  jand g10495(.dina(n10422), .dinb(n10415), .dout(n10687));
  jor  g10496(.dina(n10687), .dinb(n10686), .dout(n10688));
  jand g10497(.dina(n10408), .dinb(n10392), .dout(n10689));
  jnot g10498(.din(n10689), .dout(n10690));
  jor  g10499(.dina(n10414), .dinb(n10410), .dout(n10691));
  jand g10500(.dina(n10691), .dinb(n10690), .dout(n10692));
  jnot g10501(.din(n10692), .dout(n10693));
  jand g10502(.dina(n10447), .dinb(n10444), .dout(n10694));
  jand g10503(.dina(n10448), .dinb(n10435), .dout(n10695));
  jor  g10504(.dina(n10695), .dinb(n10694), .dout(n10696));
  jand g10505(.dina(\a[54] ), .dinb(\a[21] ), .dout(n10697));
  jnot g10506(.din(n10697), .dout(n10698));
  jand g10507(.dina(n6130), .dinb(n1814), .dout(n10699));
  jnot g10508(.din(n10699), .dout(n10700));
  jand g10509(.dina(n7559), .dinb(n1376), .dout(n10701));
  jand g10510(.dina(\a[51] ), .dinb(\a[24] ), .dout(n10702));
  jand g10511(.dina(n10702), .dinb(n10697), .dout(n10703));
  jor  g10512(.dina(n10703), .dinb(n10701), .dout(n10704));
  jand g10513(.dina(n10704), .dinb(n10700), .dout(n10705));
  jor  g10514(.dina(n10705), .dinb(n10698), .dout(n10706));
  jor  g10515(.dina(n10704), .dinb(n10699), .dout(n10707));
  jnot g10516(.din(n10707), .dout(n10708));
  jand g10517(.dina(\a[53] ), .dinb(\a[22] ), .dout(n10709));
  jor  g10518(.dina(n10709), .dinb(n10702), .dout(n10710));
  jand g10519(.dina(n10710), .dinb(n10708), .dout(n10711));
  jnot g10520(.din(n10711), .dout(n10712));
  jand g10521(.dina(n10712), .dinb(n10706), .dout(n10713));
  jand g10522(.dina(\a[41] ), .dinb(\a[34] ), .dout(n10714));
  jand g10523(.dina(\a[55] ), .dinb(\a[20] ), .dout(n10715));
  jand g10524(.dina(\a[50] ), .dinb(\a[25] ), .dout(n10716));
  jxor g10525(.dina(n10716), .dinb(n10715), .dout(n10717));
  jxor g10526(.dina(n10717), .dinb(n10714), .dout(n10718));
  jnot g10527(.din(n10718), .dout(n10719));
  jand g10528(.dina(\a[44] ), .dinb(\a[31] ), .dout(n10720));
  jnot g10529(.din(n10720), .dout(n10721));
  jand g10530(.dina(n4317), .dinb(n2671), .dout(n10722));
  jnot g10531(.din(n10722), .dout(n10723));
  jand g10532(.dina(\a[42] ), .dinb(\a[33] ), .dout(n10724));
  jor  g10533(.dina(n10724), .dinb(n4492), .dout(n10725));
  jand g10534(.dina(n10725), .dinb(n10723), .dout(n10726));
  jxor g10535(.dina(n10726), .dinb(n10721), .dout(n10727));
  jxor g10536(.dina(n10727), .dinb(n10719), .dout(n10728));
  jnot g10537(.din(n10728), .dout(n10729));
  jxor g10538(.dina(n10729), .dinb(n10713), .dout(n10730));
  jxor g10539(.dina(n10730), .dinb(n10696), .dout(n10731));
  jxor g10540(.dina(n10731), .dinb(n10693), .dout(n10732));
  jxor g10541(.dina(n10732), .dinb(n10688), .dout(n10733));
  jxor g10542(.dina(n10733), .dinb(n10685), .dout(n10734));
  jand g10543(.dina(n10423), .dinb(n10387), .dout(n10735));
  jand g10544(.dina(n10535), .dinb(n10424), .dout(n10736));
  jor  g10545(.dina(n10736), .dinb(n10735), .dout(n10737));
  jxor g10546(.dina(n10737), .dinb(n10734), .dout(n10738));
  jxor g10547(.dina(n10738), .dinb(n10682), .dout(n10739));
  jand g10548(.dina(n10739), .dinb(n10549), .dout(n10740));
  jor  g10549(.dina(n10739), .dinb(n10549), .dout(n10741));
  jnot g10550(.din(n10741), .dout(n10742));
  jor  g10551(.dina(n10742), .dinb(n10740), .dout(n10743));
  jand g10552(.dina(n10537), .dinb(n10351), .dout(n10744));
  jnot g10553(.din(n10744), .dout(n10745));
  jnot g10554(.din(n10351), .dout(n10746));
  jand g10555(.dina(n10538), .dinb(n10746), .dout(n10747));
  jor  g10556(.dina(n10545), .dinb(n10747), .dout(n10748));
  jand g10557(.dina(n10748), .dinb(n10745), .dout(n10749));
  jxor g10558(.dina(n10749), .dinb(n10743), .dout(\asquared[76] ));
  jand g10559(.dina(n10737), .dinb(n10734), .dout(n10751));
  jand g10560(.dina(n10738), .dinb(n10682), .dout(n10752));
  jor  g10561(.dina(n10752), .dinb(n10751), .dout(n10753));
  jand g10562(.dina(n10592), .dinb(n10552), .dout(n10754));
  jand g10563(.dina(n10681), .dinb(n10593), .dout(n10755));
  jor  g10564(.dina(n10755), .dinb(n10754), .dout(n10756));
  jand g10565(.dina(n10615), .dinb(n10598), .dout(n10757));
  jand g10566(.dina(n10680), .dinb(n10616), .dout(n10758));
  jor  g10567(.dina(n10758), .dinb(n10757), .dout(n10759));
  jand g10568(.dina(n10566), .dinb(n10563), .dout(n10760));
  jand g10569(.dina(n10591), .dinb(n10567), .dout(n10761));
  jor  g10570(.dina(n10761), .dinb(n10760), .dout(n10762));
  jand g10571(.dina(n10589), .dinb(n10580), .dout(n10763));
  jand g10572(.dina(n10590), .dinb(n10570), .dout(n10764));
  jor  g10573(.dina(n10764), .dinb(n10763), .dout(n10765));
  jor  g10574(.dina(n10613), .dinb(n10609), .dout(n10766));
  jand g10575(.dina(n10614), .dinb(n10606), .dout(n10767));
  jnot g10576(.din(n10767), .dout(n10768));
  jand g10577(.dina(n10768), .dinb(n10766), .dout(n10769));
  jnot g10578(.din(n10769), .dout(n10770));
  jand g10579(.dina(\a[63] ), .dinb(\a[13] ), .dout(n10771));
  jand g10580(.dina(\a[44] ), .dinb(\a[32] ), .dout(n10772));
  jand g10581(.dina(\a[45] ), .dinb(\a[31] ), .dout(n10773));
  jor  g10582(.dina(n10773), .dinb(n10772), .dout(n10774));
  jand g10583(.dina(n4812), .dinb(n3269), .dout(n10775));
  jnot g10584(.din(n10775), .dout(n10776));
  jand g10585(.dina(n10776), .dinb(n10774), .dout(n10777));
  jxor g10586(.dina(n10777), .dinb(n10771), .dout(n10778));
  jand g10587(.dina(\a[57] ), .dinb(\a[19] ), .dout(n10779));
  jand g10588(.dina(\a[53] ), .dinb(\a[23] ), .dout(n10780));
  jxor g10589(.dina(n10780), .dinb(n10779), .dout(n10781));
  jxor g10590(.dina(n10781), .dinb(n4658), .dout(n10782));
  jxor g10591(.dina(n10782), .dinb(n10778), .dout(n10783));
  jnot g10592(.din(n10783), .dout(n10784));
  jand g10593(.dina(\a[56] ), .dinb(\a[20] ), .dout(n10785));
  jnot g10594(.din(n10785), .dout(n10786));
  jand g10595(.dina(\a[55] ), .dinb(\a[22] ), .dout(n10787));
  jand g10596(.dina(n10787), .dinb(n10697), .dout(n10788));
  jnot g10597(.din(n10788), .dout(n10789));
  jand g10598(.dina(\a[55] ), .dinb(\a[21] ), .dout(n10790));
  jand g10599(.dina(\a[54] ), .dinb(\a[22] ), .dout(n10791));
  jor  g10600(.dina(n10791), .dinb(n10790), .dout(n10792));
  jand g10601(.dina(n10792), .dinb(n10789), .dout(n10793));
  jxor g10602(.dina(n10793), .dinb(n10786), .dout(n10794));
  jxor g10603(.dina(n10794), .dinb(n10784), .dout(n10795));
  jxor g10604(.dina(n10795), .dinb(n10770), .dout(n10796));
  jxor g10605(.dina(n10796), .dinb(n10765), .dout(n10797));
  jxor g10606(.dina(n10797), .dinb(n10762), .dout(n10798));
  jxor g10607(.dina(n10798), .dinb(n10759), .dout(n10799));
  jxor g10608(.dina(n10799), .dinb(n10756), .dout(n10800));
  jand g10609(.dina(n10732), .dinb(n10688), .dout(n10801));
  jand g10610(.dina(n10733), .dinb(n10685), .dout(n10802));
  jor  g10611(.dina(n10802), .dinb(n10801), .dout(n10803));
  jand g10612(.dina(n10585), .dinb(n10582), .dout(n10804));
  jand g10613(.dina(n10588), .dinb(n10586), .dout(n10805));
  jor  g10614(.dina(n10805), .dinb(n10804), .dout(n10806));
  jand g10615(.dina(n10601), .dinb(n10465), .dout(n10807));
  jand g10616(.dina(n10605), .dinb(n10602), .dout(n10808));
  jor  g10617(.dina(n10808), .dinb(n10807), .dout(n10809));
  jxor g10618(.dina(n10809), .dinb(n10806), .dout(n10810));
  jand g10619(.dina(n10578), .dinb(n10575), .dout(n10811));
  jand g10620(.dina(n10579), .dinb(n10572), .dout(n10812));
  jor  g10621(.dina(n10812), .dinb(n10811), .dout(n10813));
  jxor g10622(.dina(n10813), .dinb(n10810), .dout(n10814));
  jand g10623(.dina(n10641), .dinb(n10619), .dout(n10815));
  jand g10624(.dina(n10679), .dinb(n10642), .dout(n10816));
  jor  g10625(.dina(n10816), .dinb(n10815), .dout(n10817));
  jxor g10626(.dina(n10817), .dinb(n10814), .dout(n10818));
  jand g10627(.dina(n10622), .dinb(n10621), .dout(n10819));
  jand g10628(.dina(n10623), .dinb(n10620), .dout(n10820));
  jor  g10629(.dina(n10820), .dinb(n10819), .dout(n10821));
  jand g10630(.dina(n10716), .dinb(n10715), .dout(n10822));
  jand g10631(.dina(n10717), .dinb(n10714), .dout(n10823));
  jor  g10632(.dina(n10823), .dinb(n10822), .dout(n10824));
  jand g10633(.dina(n10674), .dinb(n10671), .dout(n10825));
  jnot g10634(.din(n10825), .dout(n10826));
  jand g10635(.dina(n10826), .dinb(n10676), .dout(n10827));
  jxor g10636(.dina(n10827), .dinb(n10824), .dout(n10828));
  jxor g10637(.dina(n10828), .dinb(n10821), .dout(n10829));
  jor  g10638(.dina(n10727), .dinb(n10719), .dout(n10830));
  jor  g10639(.dina(n10729), .dinb(n10713), .dout(n10831));
  jand g10640(.dina(n10831), .dinb(n10830), .dout(n10832));
  jand g10641(.dina(\a[62] ), .dinb(\a[14] ), .dout(n10833));
  jnot g10642(.din(\a[38] ), .dout(n10834));
  jand g10643(.dina(n10638), .dinb(n2837), .dout(n10835));
  jor  g10644(.dina(n10835), .dinb(n10834), .dout(n10836));
  jnot g10645(.din(n10836), .dout(n10837));
  jxor g10646(.dina(n10837), .dinb(n10833), .dout(n10838));
  jand g10647(.dina(n10629), .dinb(n10627), .dout(n10839));
  jnot g10648(.din(n10839), .dout(n10840));
  jand g10649(.dina(n10840), .dinb(n10632), .dout(n10841));
  jxor g10650(.dina(n10841), .dinb(n10838), .dout(n10842));
  jnot g10651(.din(n10842), .dout(n10843));
  jxor g10652(.dina(n10843), .dinb(n10832), .dout(n10844));
  jxor g10653(.dina(n10844), .dinb(n10829), .dout(n10845));
  jxor g10654(.dina(n10845), .dinb(n10818), .dout(n10846));
  jxor g10655(.dina(n10846), .dinb(n10803), .dout(n10847));
  jand g10656(.dina(n10730), .dinb(n10696), .dout(n10848));
  jand g10657(.dina(n10731), .dinb(n10693), .dout(n10849));
  jor  g10658(.dina(n10849), .dinb(n10848), .dout(n10850));
  jand g10659(.dina(n10666), .dinb(n10660), .dout(n10851));
  jor  g10660(.dina(n10851), .dinb(n10662), .dout(n10852));
  jxor g10661(.dina(n10852), .dinb(n10654), .dout(n10853));
  jand g10662(.dina(n10723), .dinb(n10721), .dout(n10854));
  jnot g10663(.din(n10854), .dout(n10855));
  jand g10664(.dina(n10855), .dinb(n10725), .dout(n10856));
  jxor g10665(.dina(n10856), .dinb(n10853), .dout(n10857));
  jand g10666(.dina(n10667), .dinb(n10659), .dout(n10858));
  jnot g10667(.din(n10858), .dout(n10859));
  jor  g10668(.dina(n10678), .dinb(n10669), .dout(n10860));
  jand g10669(.dina(n10860), .dinb(n10859), .dout(n10861));
  jor  g10670(.dina(n10634), .dinb(n10625), .dout(n10862));
  jor  g10671(.dina(n10640), .dinb(n10636), .dout(n10863));
  jand g10672(.dina(n10863), .dinb(n10862), .dout(n10864));
  jxor g10673(.dina(n10864), .dinb(n10861), .dout(n10865));
  jxor g10674(.dina(n10865), .dinb(n10857), .dout(n10866));
  jxor g10675(.dina(n10866), .dinb(n10850), .dout(n10867));
  jand g10676(.dina(n10558), .dinb(n10555), .dout(n10868));
  jand g10677(.dina(n10562), .dinb(n10559), .dout(n10869));
  jor  g10678(.dina(n10869), .dinb(n10868), .dout(n10870));
  jand g10679(.dina(\a[48] ), .dinb(\a[28] ), .dout(n10871));
  jand g10680(.dina(\a[47] ), .dinb(\a[30] ), .dout(n10872));
  jand g10681(.dina(n10872), .dinb(n10675), .dout(n10873));
  jnot g10682(.din(n10873), .dout(n10874));
  jand g10683(.dina(\a[46] ), .dinb(\a[30] ), .dout(n10875));
  jor  g10684(.dina(n10875), .dinb(n10672), .dout(n10876));
  jand g10685(.dina(n10876), .dinb(n10874), .dout(n10877));
  jxor g10686(.dina(n10877), .dinb(n10871), .dout(n10878));
  jnot g10687(.din(n10878), .dout(n10879));
  jand g10688(.dina(\a[42] ), .dinb(\a[34] ), .dout(n10880));
  jnot g10689(.din(n10880), .dout(n10881));
  jand g10690(.dina(n4632), .dinb(n3243), .dout(n10882));
  jnot g10691(.din(n10882), .dout(n10883));
  jand g10692(.dina(\a[40] ), .dinb(\a[36] ), .dout(n10884));
  jand g10693(.dina(\a[41] ), .dinb(\a[35] ), .dout(n10885));
  jor  g10694(.dina(n10885), .dinb(n10884), .dout(n10886));
  jand g10695(.dina(n10886), .dinb(n10883), .dout(n10887));
  jxor g10696(.dina(n10887), .dinb(n10881), .dout(n10888));
  jxor g10697(.dina(n10888), .dinb(n10879), .dout(n10889));
  jnot g10698(.din(n10889), .dout(n10890));
  jnot g10699(.din(n4865), .dout(n10891));
  jand g10700(.dina(\a[52] ), .dinb(\a[25] ), .dout(n10892));
  jand g10701(.dina(n10892), .dinb(n10702), .dout(n10893));
  jnot g10702(.din(n10893), .dout(n10894));
  jand g10703(.dina(\a[52] ), .dinb(\a[24] ), .dout(n10895));
  jand g10704(.dina(\a[51] ), .dinb(\a[25] ), .dout(n10896));
  jor  g10705(.dina(n10896), .dinb(n10895), .dout(n10897));
  jand g10706(.dina(n10897), .dinb(n10894), .dout(n10898));
  jxor g10707(.dina(n10898), .dinb(n10891), .dout(n10899));
  jxor g10708(.dina(n10899), .dinb(n10890), .dout(n10900));
  jxor g10709(.dina(n10900), .dinb(n10870), .dout(n10901));
  jand g10710(.dina(\a[61] ), .dinb(\a[15] ), .dout(n10902));
  jnot g10711(.din(n10902), .dout(n10903));
  jand g10712(.dina(\a[60] ), .dinb(\a[17] ), .dout(n10904));
  jand g10713(.dina(n10904), .dinb(n10399), .dout(n10905));
  jnot g10714(.din(n10905), .dout(n10906));
  jand g10715(.dina(\a[59] ), .dinb(\a[17] ), .dout(n10907));
  jor  g10716(.dina(n10907), .dinb(n10661), .dout(n10908));
  jand g10717(.dina(n10908), .dinb(n10906), .dout(n10909));
  jxor g10718(.dina(n10909), .dinb(n10903), .dout(n10910));
  jxor g10719(.dina(n10910), .dinb(n10708), .dout(n10911));
  jand g10720(.dina(\a[58] ), .dinb(\a[18] ), .dout(n10912));
  jand g10721(.dina(\a[50] ), .dinb(\a[27] ), .dout(n10913));
  jand g10722(.dina(n10913), .dinb(n10647), .dout(n10914));
  jnot g10723(.din(n10914), .dout(n10915));
  jand g10724(.dina(\a[50] ), .dinb(\a[26] ), .dout(n10916));
  jand g10725(.dina(\a[49] ), .dinb(\a[27] ), .dout(n10917));
  jor  g10726(.dina(n10917), .dinb(n10916), .dout(n10918));
  jand g10727(.dina(n10918), .dinb(n10915), .dout(n10919));
  jxor g10728(.dina(n10919), .dinb(n10912), .dout(n10920));
  jxor g10729(.dina(n10920), .dinb(n10911), .dout(n10921));
  jxor g10730(.dina(n10921), .dinb(n10901), .dout(n10922));
  jxor g10731(.dina(n10922), .dinb(n10867), .dout(n10923));
  jxor g10732(.dina(n10923), .dinb(n10847), .dout(n10924));
  jxor g10733(.dina(n10924), .dinb(n10800), .dout(n10925));
  jand g10734(.dina(n10925), .dinb(n10753), .dout(n10926));
  jor  g10735(.dina(n10925), .dinb(n10753), .dout(n10927));
  jnot g10736(.din(n10927), .dout(n10928));
  jor  g10737(.dina(n10928), .dinb(n10926), .dout(n10929));
  jnot g10738(.din(n10740), .dout(n10930));
  jor  g10739(.dina(n10749), .dinb(n10742), .dout(n10931));
  jand g10740(.dina(n10931), .dinb(n10930), .dout(n10932));
  jxor g10741(.dina(n10932), .dinb(n10929), .dout(\asquared[77] ));
  jand g10742(.dina(n10799), .dinb(n10756), .dout(n10934));
  jand g10743(.dina(n10924), .dinb(n10800), .dout(n10935));
  jor  g10744(.dina(n10935), .dinb(n10934), .dout(n10936));
  jand g10745(.dina(n10846), .dinb(n10803), .dout(n10937));
  jand g10746(.dina(n10923), .dinb(n10847), .dout(n10938));
  jor  g10747(.dina(n10938), .dinb(n10937), .dout(n10939));
  jand g10748(.dina(n10866), .dinb(n10850), .dout(n10940));
  jand g10749(.dina(n10922), .dinb(n10867), .dout(n10941));
  jor  g10750(.dina(n10941), .dinb(n10940), .dout(n10942));
  jand g10751(.dina(n10817), .dinb(n10814), .dout(n10943));
  jand g10752(.dina(n10845), .dinb(n10818), .dout(n10944));
  jor  g10753(.dina(n10944), .dinb(n10943), .dout(n10945));
  jor  g10754(.dina(n10843), .dinb(n10832), .dout(n10946));
  jand g10755(.dina(n10844), .dinb(n10829), .dout(n10947));
  jnot g10756(.din(n10947), .dout(n10948));
  jand g10757(.dina(n10948), .dinb(n10946), .dout(n10949));
  jnot g10758(.din(n10949), .dout(n10950));
  jor  g10759(.dina(n10864), .dinb(n10861), .dout(n10951));
  jand g10760(.dina(n10865), .dinb(n10857), .dout(n10952));
  jnot g10761(.din(n10952), .dout(n10953));
  jand g10762(.dina(n10953), .dinb(n10951), .dout(n10954));
  jnot g10763(.din(n10954), .dout(n10955));
  jand g10764(.dina(\a[43] ), .dinb(\a[34] ), .dout(n10956));
  jand g10765(.dina(\a[51] ), .dinb(\a[26] ), .dout(n10957));
  jxor g10766(.dina(n10957), .dinb(n10787), .dout(n10958));
  jxor g10767(.dina(n10958), .dinb(n10956), .dout(n10959));
  jnot g10768(.din(n10959), .dout(n10960));
  jnot g10769(.din(n10892), .dout(n10961));
  jand g10770(.dina(n7559), .dinb(n1942), .dout(n10962));
  jnot g10771(.din(n10962), .dout(n10963));
  jand g10772(.dina(\a[54] ), .dinb(\a[23] ), .dout(n10964));
  jand g10773(.dina(\a[53] ), .dinb(\a[24] ), .dout(n10965));
  jor  g10774(.dina(n10965), .dinb(n10964), .dout(n10966));
  jand g10775(.dina(n10966), .dinb(n10963), .dout(n10967));
  jxor g10776(.dina(n10967), .dinb(n10961), .dout(n10968));
  jxor g10777(.dina(n10968), .dinb(n10960), .dout(n10969));
  jnot g10778(.din(n10969), .dout(n10970));
  jand g10779(.dina(\a[61] ), .dinb(\a[16] ), .dout(n10971));
  jnot g10780(.din(n10971), .dout(n10972));
  jand g10781(.dina(n4812), .dinb(n2671), .dout(n10973));
  jnot g10782(.din(n10973), .dout(n10974));
  jand g10783(.dina(\a[45] ), .dinb(\a[32] ), .dout(n10975));
  jand g10784(.dina(\a[44] ), .dinb(\a[33] ), .dout(n10976));
  jor  g10785(.dina(n10976), .dinb(n10975), .dout(n10977));
  jand g10786(.dina(n10977), .dinb(n10974), .dout(n10978));
  jxor g10787(.dina(n10978), .dinb(n10972), .dout(n10979));
  jxor g10788(.dina(n10979), .dinb(n10970), .dout(n10980));
  jxor g10789(.dina(n10980), .dinb(n10955), .dout(n10981));
  jxor g10790(.dina(n10981), .dinb(n10950), .dout(n10982));
  jxor g10791(.dina(n10982), .dinb(n10945), .dout(n10983));
  jxor g10792(.dina(n10983), .dinb(n10942), .dout(n10984));
  jxor g10793(.dina(n10984), .dinb(n10939), .dout(n10985));
  jand g10794(.dina(n10797), .dinb(n10762), .dout(n10986));
  jand g10795(.dina(n10798), .dinb(n10759), .dout(n10987));
  jor  g10796(.dina(n10987), .dinb(n10986), .dout(n10988));
  jand g10797(.dina(n10852), .dinb(n10654), .dout(n10989));
  jand g10798(.dina(n10856), .dinb(n10853), .dout(n10990));
  jor  g10799(.dina(n10990), .dinb(n10989), .dout(n10991));
  jand g10800(.dina(\a[60] ), .dinb(\a[18] ), .dout(n10992));
  jand g10801(.dina(n10992), .dinb(n10907), .dout(n10993));
  jnot g10802(.din(n10993), .dout(n10994));
  jand g10803(.dina(\a[59] ), .dinb(\a[18] ), .dout(n10995));
  jor  g10804(.dina(n10995), .dinb(n10904), .dout(n10996));
  jand g10805(.dina(n10996), .dinb(n10994), .dout(n10997));
  jand g10806(.dina(n10894), .dinb(n10891), .dout(n10998));
  jnot g10807(.din(n10998), .dout(n10999));
  jand g10808(.dina(n10999), .dinb(n10897), .dout(n11000));
  jxor g10809(.dina(n11000), .dinb(n10997), .dout(n11001));
  jxor g10810(.dina(n11001), .dinb(n10991), .dout(n11002));
  jand g10811(.dina(n10827), .dinb(n10824), .dout(n11003));
  jand g10812(.dina(n10828), .dinb(n10821), .dout(n11004));
  jor  g10813(.dina(n11004), .dinb(n11003), .dout(n11005));
  jxor g10814(.dina(n11005), .dinb(n11002), .dout(n11006));
  jand g10815(.dina(n10900), .dinb(n10870), .dout(n11007));
  jand g10816(.dina(n10921), .dinb(n10901), .dout(n11008));
  jor  g10817(.dina(n11008), .dinb(n11007), .dout(n11009));
  jxor g10818(.dina(n11009), .dinb(n11006), .dout(n11010));
  jand g10819(.dina(n10777), .dinb(n10771), .dout(n11011));
  jor  g10820(.dina(n11011), .dinb(n10775), .dout(n11012));
  jand g10821(.dina(n10877), .dinb(n10871), .dout(n11013));
  jor  g10822(.dina(n11013), .dinb(n10873), .dout(n11014));
  jand g10823(.dina(n10789), .dinb(n10786), .dout(n11015));
  jnot g10824(.din(n11015), .dout(n11016));
  jand g10825(.dina(n11016), .dinb(n10792), .dout(n11017));
  jxor g10826(.dina(n11017), .dinb(n11014), .dout(n11018));
  jxor g10827(.dina(n11018), .dinb(n11012), .dout(n11019));
  jand g10828(.dina(n10780), .dinb(n10779), .dout(n11020));
  jand g10829(.dina(n10781), .dinb(n4658), .dout(n11021));
  jor  g10830(.dina(n11021), .dinb(n11020), .dout(n11022));
  jand g10831(.dina(n10918), .dinb(n10912), .dout(n11023));
  jor  g10832(.dina(n11023), .dinb(n10914), .dout(n11024));
  jand g10833(.dina(n10906), .dinb(n10903), .dout(n11025));
  jnot g10834(.din(n11025), .dout(n11026));
  jand g10835(.dina(n11026), .dinb(n10908), .dout(n11027));
  jxor g10836(.dina(n11027), .dinb(n11024), .dout(n11028));
  jxor g10837(.dina(n11028), .dinb(n11022), .dout(n11029));
  jnot g10838(.din(n11029), .dout(n11030));
  jand g10839(.dina(n10782), .dinb(n10778), .dout(n11031));
  jnot g10840(.din(n11031), .dout(n11032));
  jor  g10841(.dina(n10794), .dinb(n10784), .dout(n11033));
  jand g10842(.dina(n11033), .dinb(n11032), .dout(n11034));
  jxor g10843(.dina(n11034), .dinb(n11030), .dout(n11035));
  jxor g10844(.dina(n11035), .dinb(n11019), .dout(n11036));
  jxor g10845(.dina(n11036), .dinb(n11010), .dout(n11037));
  jxor g10846(.dina(n11037), .dinb(n10988), .dout(n11038));
  jand g10847(.dina(n10837), .dinb(n10833), .dout(n11039));
  jand g10848(.dina(n10841), .dinb(n10838), .dout(n11040));
  jor  g10849(.dina(n11040), .dinb(n11039), .dout(n11041));
  jnot g10850(.din(n11041), .dout(n11042));
  jor  g10851(.dina(n10910), .dinb(n10708), .dout(n11043));
  jand g10852(.dina(n10920), .dinb(n10911), .dout(n11044));
  jnot g10853(.din(n11044), .dout(n11045));
  jand g10854(.dina(n11045), .dinb(n11043), .dout(n11046));
  jxor g10855(.dina(n11046), .dinb(n11042), .dout(n11047));
  jnot g10856(.din(n11047), .dout(n11048));
  jor  g10857(.dina(n10888), .dinb(n10879), .dout(n11049));
  jor  g10858(.dina(n10899), .dinb(n10890), .dout(n11050));
  jand g10859(.dina(n11050), .dinb(n11049), .dout(n11051));
  jxor g10860(.dina(n11051), .dinb(n11048), .dout(n11052));
  jand g10861(.dina(n10795), .dinb(n10770), .dout(n11053));
  jand g10862(.dina(n10796), .dinb(n10765), .dout(n11054));
  jor  g10863(.dina(n11054), .dinb(n11053), .dout(n11055));
  jxor g10864(.dina(n11055), .dinb(n11052), .dout(n11056));
  jand g10865(.dina(n10809), .dinb(n10806), .dout(n11057));
  jand g10866(.dina(n10813), .dinb(n10810), .dout(n11058));
  jor  g10867(.dina(n11058), .dinb(n11057), .dout(n11059));
  jand g10868(.dina(\a[46] ), .dinb(\a[31] ), .dout(n11060));
  jand g10869(.dina(\a[63] ), .dinb(\a[14] ), .dout(n11061));
  jand g10870(.dina(n11061), .dinb(n11060), .dout(n11062));
  jnot g10871(.din(n11062), .dout(n11063));
  jand g10872(.dina(\a[47] ), .dinb(\a[31] ), .dout(n11064));
  jand g10873(.dina(n11064), .dinb(n10875), .dout(n11065));
  jand g10874(.dina(n11061), .dinb(n10872), .dout(n11066));
  jor  g10875(.dina(n11066), .dinb(n11065), .dout(n11067));
  jnot g10876(.din(n11067), .dout(n11068));
  jand g10877(.dina(n11068), .dinb(n11063), .dout(n11069));
  jor  g10878(.dina(n11061), .dinb(n11060), .dout(n11070));
  jand g10879(.dina(n11070), .dinb(n11069), .dout(n11071));
  jand g10880(.dina(n11067), .dinb(n11063), .dout(n11072));
  jnot g10881(.din(n11072), .dout(n11073));
  jand g10882(.dina(n11073), .dinb(n10872), .dout(n11074));
  jor  g10883(.dina(n11074), .dinb(n11071), .dout(n11075));
  jand g10884(.dina(\a[42] ), .dinb(\a[35] ), .dout(n11076));
  jnot g10885(.din(n11076), .dout(n11077));
  jand g10886(.dina(n4632), .dinb(n3138), .dout(n11078));
  jnot g10887(.din(n11078), .dout(n11079));
  jand g10888(.dina(\a[41] ), .dinb(\a[36] ), .dout(n11080));
  jand g10889(.dina(\a[40] ), .dinb(\a[37] ), .dout(n11081));
  jor  g10890(.dina(n11081), .dinb(n11080), .dout(n11082));
  jand g10891(.dina(n11082), .dinb(n11079), .dout(n11083));
  jxor g10892(.dina(n11083), .dinb(n11077), .dout(n11084));
  jnot g10893(.din(n11084), .dout(n11085));
  jxor g10894(.dina(n11085), .dinb(n11075), .dout(n11086));
  jnot g10895(.din(n11086), .dout(n11087));
  jand g10896(.dina(\a[62] ), .dinb(\a[15] ), .dout(n11088));
  jnot g10897(.din(n11088), .dout(n11089));
  jand g10898(.dina(\a[39] ), .dinb(n10834), .dout(n11090));
  jxor g10899(.dina(n11090), .dinb(n11089), .dout(n11091));
  jxor g10900(.dina(n11091), .dinb(n11087), .dout(n11092));
  jxor g10901(.dina(n11092), .dinb(n11059), .dout(n11093));
  jand g10902(.dina(n10883), .dinb(n10881), .dout(n11094));
  jnot g10903(.din(n11094), .dout(n11095));
  jand g10904(.dina(n11095), .dinb(n10886), .dout(n11096));
  jnot g10905(.din(n11096), .dout(n11097));
  jand g10906(.dina(\a[58] ), .dinb(\a[19] ), .dout(n11098));
  jnot g10907(.din(n11098), .dout(n11099));
  jand g10908(.dina(\a[57] ), .dinb(\a[21] ), .dout(n11100));
  jand g10909(.dina(n11100), .dinb(n10785), .dout(n11101));
  jnot g10910(.din(n11101), .dout(n11102));
  jand g10911(.dina(\a[57] ), .dinb(\a[20] ), .dout(n11103));
  jand g10912(.dina(\a[56] ), .dinb(\a[21] ), .dout(n11104));
  jor  g10913(.dina(n11104), .dinb(n11103), .dout(n11105));
  jand g10914(.dina(n11105), .dinb(n11102), .dout(n11106));
  jxor g10915(.dina(n11106), .dinb(n11099), .dout(n11107));
  jxor g10916(.dina(n11107), .dinb(n11097), .dout(n11108));
  jnot g10917(.din(n11108), .dout(n11109));
  jnot g10918(.din(n10913), .dout(n11110));
  jand g10919(.dina(n7729), .dinb(n2653), .dout(n11111));
  jnot g10920(.din(n11111), .dout(n11112));
  jand g10921(.dina(\a[49] ), .dinb(\a[28] ), .dout(n11113));
  jand g10922(.dina(\a[48] ), .dinb(\a[29] ), .dout(n11114));
  jor  g10923(.dina(n11114), .dinb(n11113), .dout(n11115));
  jand g10924(.dina(n11115), .dinb(n11112), .dout(n11116));
  jxor g10925(.dina(n11116), .dinb(n11110), .dout(n11117));
  jxor g10926(.dina(n11117), .dinb(n11109), .dout(n11118));
  jxor g10927(.dina(n11118), .dinb(n11093), .dout(n11119));
  jxor g10928(.dina(n11119), .dinb(n11056), .dout(n11120));
  jxor g10929(.dina(n11120), .dinb(n11038), .dout(n11121));
  jxor g10930(.dina(n11121), .dinb(n10985), .dout(n11122));
  jand g10931(.dina(n11122), .dinb(n10936), .dout(n11123));
  jor  g10932(.dina(n11122), .dinb(n10936), .dout(n11124));
  jnot g10933(.din(n11124), .dout(n11125));
  jor  g10934(.dina(n11125), .dinb(n11123), .dout(n11126));
  jnot g10935(.din(n10926), .dout(n11127));
  jor  g10936(.dina(n10932), .dinb(n10928), .dout(n11128));
  jand g10937(.dina(n11128), .dinb(n11127), .dout(n11129));
  jxor g10938(.dina(n11129), .dinb(n11126), .dout(\asquared[78] ));
  jand g10939(.dina(n10984), .dinb(n10939), .dout(n11131));
  jand g10940(.dina(n11121), .dinb(n10985), .dout(n11132));
  jor  g10941(.dina(n11132), .dinb(n11131), .dout(n11133));
  jand g10942(.dina(n11055), .dinb(n11052), .dout(n11134));
  jand g10943(.dina(n11119), .dinb(n11056), .dout(n11135));
  jor  g10944(.dina(n11135), .dinb(n11134), .dout(n11136));
  jand g10945(.dina(n11009), .dinb(n11006), .dout(n11137));
  jand g10946(.dina(n11036), .dinb(n11010), .dout(n11138));
  jor  g10947(.dina(n11138), .dinb(n11137), .dout(n11139));
  jor  g10948(.dina(n11046), .dinb(n11042), .dout(n11140));
  jor  g10949(.dina(n11051), .dinb(n11048), .dout(n11141));
  jand g10950(.dina(n11141), .dinb(n11140), .dout(n11142));
  jnot g10951(.din(n11142), .dout(n11143));
  jand g10952(.dina(\a[59] ), .dinb(\a[57] ), .dout(n11144));
  jand g10953(.dina(n11144), .dinb(n3334), .dout(n11145));
  jnot g10954(.din(n11145), .dout(n11146));
  jand g10955(.dina(\a[59] ), .dinb(\a[19] ), .dout(n11147));
  jor  g10956(.dina(n11147), .dinb(n11100), .dout(n11148));
  jand g10957(.dina(n11148), .dinb(n11146), .dout(n11149));
  jxor g10958(.dina(n11149), .dinb(n10992), .dout(n11150));
  jand g10959(.dina(\a[51] ), .dinb(\a[27] ), .dout(n11151));
  jand g10960(.dina(\a[50] ), .dinb(\a[29] ), .dout(n11152));
  jand g10961(.dina(n11152), .dinb(n11113), .dout(n11153));
  jnot g10962(.din(n11153), .dout(n11154));
  jand g10963(.dina(\a[50] ), .dinb(\a[28] ), .dout(n11155));
  jand g10964(.dina(\a[49] ), .dinb(\a[29] ), .dout(n11156));
  jor  g10965(.dina(n11156), .dinb(n11155), .dout(n11157));
  jand g10966(.dina(n11157), .dinb(n11154), .dout(n11158));
  jxor g10967(.dina(n11158), .dinb(n11151), .dout(n11159));
  jxor g10968(.dina(n11159), .dinb(n11150), .dout(n11160));
  jnot g10969(.din(n11160), .dout(n11161));
  jand g10970(.dina(\a[63] ), .dinb(\a[15] ), .dout(n11162));
  jnot g10971(.din(n11162), .dout(n11163));
  jand g10972(.dina(n8702), .dinb(n937), .dout(n11164));
  jnot g10973(.din(n11164), .dout(n11165));
  jand g10974(.dina(\a[62] ), .dinb(\a[16] ), .dout(n11166));
  jand g10975(.dina(\a[61] ), .dinb(\a[17] ), .dout(n11167));
  jor  g10976(.dina(n11167), .dinb(n11166), .dout(n11168));
  jand g10977(.dina(n11168), .dinb(n11165), .dout(n11169));
  jxor g10978(.dina(n11169), .dinb(n11163), .dout(n11170));
  jxor g10979(.dina(n11170), .dinb(n11161), .dout(n11171));
  jand g10980(.dina(\a[58] ), .dinb(\a[20] ), .dout(n11172));
  jand g10981(.dina(\a[48] ), .dinb(\a[30] ), .dout(n11173));
  jor  g10982(.dina(n11173), .dinb(n11064), .dout(n11174));
  jand g10983(.dina(n5316), .dinb(n2440), .dout(n11175));
  jnot g10984(.din(n11175), .dout(n11176));
  jand g10985(.dina(n11176), .dinb(n11174), .dout(n11177));
  jxor g10986(.dina(n11177), .dinb(n11172), .dout(n11178));
  jand g10987(.dina(\a[46] ), .dinb(\a[32] ), .dout(n11179));
  jand g10988(.dina(\a[45] ), .dinb(\a[33] ), .dout(n11180));
  jand g10989(.dina(\a[44] ), .dinb(\a[34] ), .dout(n11181));
  jor  g10990(.dina(n11181), .dinb(n11180), .dout(n11182));
  jand g10991(.dina(n4812), .dinb(n3634), .dout(n11183));
  jnot g10992(.din(n11183), .dout(n11184));
  jand g10993(.dina(n11184), .dinb(n11182), .dout(n11185));
  jxor g10994(.dina(n11185), .dinb(n11179), .dout(n11186));
  jxor g10995(.dina(n11186), .dinb(n11178), .dout(n11187));
  jnot g10996(.din(n11187), .dout(n11188));
  jand g10997(.dina(\a[53] ), .dinb(\a[25] ), .dout(n11189));
  jnot g10998(.din(n11189), .dout(n11190));
  jand g10999(.dina(\a[56] ), .dinb(\a[54] ), .dout(n11191));
  jand g11000(.dina(n11191), .dinb(n1814), .dout(n11192));
  jnot g11001(.din(n11192), .dout(n11193));
  jand g11002(.dina(\a[54] ), .dinb(\a[24] ), .dout(n11194));
  jand g11003(.dina(\a[56] ), .dinb(\a[22] ), .dout(n11195));
  jor  g11004(.dina(n11195), .dinb(n11194), .dout(n11196));
  jand g11005(.dina(n11196), .dinb(n11193), .dout(n11197));
  jxor g11006(.dina(n11197), .dinb(n11190), .dout(n11198));
  jxor g11007(.dina(n11198), .dinb(n11188), .dout(n11199));
  jxor g11008(.dina(n11199), .dinb(n11171), .dout(n11200));
  jxor g11009(.dina(n11200), .dinb(n11143), .dout(n11201));
  jxor g11010(.dina(n11201), .dinb(n11139), .dout(n11202));
  jxor g11011(.dina(n11202), .dinb(n11136), .dout(n11203));
  jand g11012(.dina(n11037), .dinb(n10988), .dout(n11204));
  jand g11013(.dina(n11120), .dinb(n11038), .dout(n11205));
  jor  g11014(.dina(n11205), .dinb(n11204), .dout(n11206));
  jxor g11015(.dina(n11206), .dinb(n11203), .dout(n11207));
  jand g11016(.dina(n10982), .dinb(n10945), .dout(n11208));
  jand g11017(.dina(n10983), .dinb(n10942), .dout(n11209));
  jor  g11018(.dina(n11209), .dinb(n11208), .dout(n11210));
  jor  g11019(.dina(n11107), .dinb(n11097), .dout(n11211));
  jor  g11020(.dina(n11117), .dinb(n11109), .dout(n11212));
  jand g11021(.dina(n11212), .dinb(n11211), .dout(n11213));
  jand g11022(.dina(n11085), .dinb(n11075), .dout(n11214));
  jnot g11023(.din(n11214), .dout(n11215));
  jor  g11024(.dina(n11091), .dinb(n11087), .dout(n11216));
  jand g11025(.dina(n11216), .dinb(n11215), .dout(n11217));
  jxor g11026(.dina(n11217), .dinb(n11213), .dout(n11218));
  jnot g11027(.din(n11218), .dout(n11219));
  jor  g11028(.dina(n10968), .dinb(n10960), .dout(n11220));
  jor  g11029(.dina(n10979), .dinb(n10970), .dout(n11221));
  jand g11030(.dina(n11221), .dinb(n11220), .dout(n11222));
  jxor g11031(.dina(n11222), .dinb(n11219), .dout(n11223));
  jnot g11032(.din(n11223), .dout(n11224));
  jor  g11033(.dina(n11034), .dinb(n11030), .dout(n11225));
  jand g11034(.dina(n11035), .dinb(n11019), .dout(n11226));
  jnot g11035(.din(n11226), .dout(n11227));
  jand g11036(.dina(n11227), .dinb(n11225), .dout(n11228));
  jxor g11037(.dina(n11228), .dinb(n11224), .dout(n11229));
  jnot g11038(.din(\a[39] ), .dout(n11230));
  jand g11039(.dina(n11089), .dinb(n10834), .dout(n11231));
  jor  g11040(.dina(n11231), .dinb(n11230), .dout(n11232));
  jnot g11041(.din(n11232), .dout(n11233));
  jand g11042(.dina(n11079), .dinb(n11077), .dout(n11234));
  jnot g11043(.din(n11234), .dout(n11235));
  jand g11044(.dina(n11235), .dinb(n11082), .dout(n11236));
  jxor g11045(.dina(n11236), .dinb(n11233), .dout(n11237));
  jand g11046(.dina(n10963), .dinb(n10961), .dout(n11238));
  jnot g11047(.din(n11238), .dout(n11239));
  jand g11048(.dina(n11239), .dinb(n10966), .dout(n11240));
  jxor g11049(.dina(n11240), .dinb(n11237), .dout(n11241));
  jnot g11050(.din(n11069), .dout(n11242));
  jand g11051(.dina(n11112), .dinb(n11110), .dout(n11243));
  jnot g11052(.din(n11243), .dout(n11244));
  jand g11053(.dina(n11244), .dinb(n11115), .dout(n11245));
  jxor g11054(.dina(n11245), .dinb(n11242), .dout(n11246));
  jand g11055(.dina(n10974), .dinb(n10972), .dout(n11247));
  jnot g11056(.din(n11247), .dout(n11248));
  jand g11057(.dina(n11248), .dinb(n10977), .dout(n11249));
  jxor g11058(.dina(n11249), .dinb(n11246), .dout(n11250));
  jand g11059(.dina(n11027), .dinb(n11024), .dout(n11251));
  jand g11060(.dina(n11028), .dinb(n11022), .dout(n11252));
  jor  g11061(.dina(n11252), .dinb(n11251), .dout(n11253));
  jxor g11062(.dina(n11253), .dinb(n11250), .dout(n11254));
  jxor g11063(.dina(n11254), .dinb(n11241), .dout(n11255));
  jxor g11064(.dina(n11255), .dinb(n11229), .dout(n11256));
  jxor g11065(.dina(n11256), .dinb(n11210), .dout(n11257));
  jand g11066(.dina(n11017), .dinb(n11014), .dout(n11258));
  jand g11067(.dina(n11018), .dinb(n11012), .dout(n11259));
  jor  g11068(.dina(n11259), .dinb(n11258), .dout(n11260));
  jnot g11069(.din(n5046), .dout(n11261));
  jand g11070(.dina(\a[40] ), .dinb(\a[38] ), .dout(n11262));
  jand g11071(.dina(\a[52] ), .dinb(\a[26] ), .dout(n11263));
  jand g11072(.dina(n11263), .dinb(n11262), .dout(n11264));
  jnot g11073(.din(n11264), .dout(n11265));
  jand g11074(.dina(n11263), .dinb(n5046), .dout(n11266));
  jand g11075(.dina(\a[41] ), .dinb(\a[38] ), .dout(n11267));
  jand g11076(.dina(n11267), .dinb(n11081), .dout(n11268));
  jor  g11077(.dina(n11268), .dinb(n11266), .dout(n11269));
  jand g11078(.dina(n11269), .dinb(n11265), .dout(n11270));
  jor  g11079(.dina(n11270), .dinb(n11261), .dout(n11271));
  jor  g11080(.dina(n11269), .dinb(n11264), .dout(n11272));
  jnot g11081(.din(n11262), .dout(n11273));
  jnot g11082(.din(n11263), .dout(n11274));
  jand g11083(.dina(n11274), .dinb(n11273), .dout(n11275));
  jor  g11084(.dina(n11275), .dinb(n11272), .dout(n11276));
  jand g11085(.dina(n11276), .dinb(n11271), .dout(n11277));
  jand g11086(.dina(\a[55] ), .dinb(\a[23] ), .dout(n11278));
  jand g11087(.dina(\a[42] ), .dinb(\a[36] ), .dout(n11279));
  jor  g11088(.dina(n11279), .dinb(n4783), .dout(n11280));
  jand g11089(.dina(n4317), .dinb(n3243), .dout(n11281));
  jnot g11090(.din(n11281), .dout(n11282));
  jand g11091(.dina(n11282), .dinb(n11280), .dout(n11283));
  jxor g11092(.dina(n11283), .dinb(n11278), .dout(n11284));
  jnot g11093(.din(n11284), .dout(n11285));
  jxor g11094(.dina(n11285), .dinb(n11277), .dout(n11286));
  jxor g11095(.dina(n11286), .dinb(n11260), .dout(n11287));
  jand g11096(.dina(n10957), .dinb(n10787), .dout(n11288));
  jand g11097(.dina(n10958), .dinb(n10956), .dout(n11289));
  jor  g11098(.dina(n11289), .dinb(n11288), .dout(n11290));
  jand g11099(.dina(n11102), .dinb(n11099), .dout(n11291));
  jnot g11100(.din(n11291), .dout(n11292));
  jand g11101(.dina(n11292), .dinb(n11105), .dout(n11293));
  jxor g11102(.dina(n11293), .dinb(n11290), .dout(n11294));
  jand g11103(.dina(n11000), .dinb(n10997), .dout(n11295));
  jor  g11104(.dina(n11295), .dinb(n10993), .dout(n11296));
  jxor g11105(.dina(n11296), .dinb(n11294), .dout(n11297));
  jand g11106(.dina(n11001), .dinb(n10991), .dout(n11298));
  jand g11107(.dina(n11005), .dinb(n11002), .dout(n11299));
  jor  g11108(.dina(n11299), .dinb(n11298), .dout(n11300));
  jxor g11109(.dina(n11300), .dinb(n11297), .dout(n11301));
  jxor g11110(.dina(n11301), .dinb(n11287), .dout(n11302));
  jand g11111(.dina(n10980), .dinb(n10955), .dout(n11303));
  jand g11112(.dina(n10981), .dinb(n10950), .dout(n11304));
  jor  g11113(.dina(n11304), .dinb(n11303), .dout(n11305));
  jand g11114(.dina(n11092), .dinb(n11059), .dout(n11306));
  jand g11115(.dina(n11118), .dinb(n11093), .dout(n11307));
  jor  g11116(.dina(n11307), .dinb(n11306), .dout(n11308));
  jxor g11117(.dina(n11308), .dinb(n11305), .dout(n11309));
  jxor g11118(.dina(n11309), .dinb(n11302), .dout(n11310));
  jxor g11119(.dina(n11310), .dinb(n11257), .dout(n11311));
  jxor g11120(.dina(n11311), .dinb(n11207), .dout(n11312));
  jand g11121(.dina(n11312), .dinb(n11133), .dout(n11313));
  jor  g11122(.dina(n11312), .dinb(n11133), .dout(n11314));
  jnot g11123(.din(n11314), .dout(n11315));
  jor  g11124(.dina(n11315), .dinb(n11313), .dout(n11316));
  jnot g11125(.din(n11123), .dout(n11317));
  jor  g11126(.dina(n11129), .dinb(n11125), .dout(n11318));
  jand g11127(.dina(n11318), .dinb(n11317), .dout(n11319));
  jxor g11128(.dina(n11319), .dinb(n11316), .dout(\asquared[79] ));
  jand g11129(.dina(n11206), .dinb(n11203), .dout(n11321));
  jand g11130(.dina(n11311), .dinb(n11207), .dout(n11322));
  jor  g11131(.dina(n11322), .dinb(n11321), .dout(n11323));
  jand g11132(.dina(n11308), .dinb(n11305), .dout(n11324));
  jand g11133(.dina(n11309), .dinb(n11302), .dout(n11325));
  jor  g11134(.dina(n11325), .dinb(n11324), .dout(n11326));
  jand g11135(.dina(n11199), .dinb(n11171), .dout(n11327));
  jand g11136(.dina(n11200), .dinb(n11143), .dout(n11328));
  jor  g11137(.dina(n11328), .dinb(n11327), .dout(n11329));
  jand g11138(.dina(n11149), .dinb(n10992), .dout(n11330));
  jor  g11139(.dina(n11330), .dinb(n11145), .dout(n11331));
  jand g11140(.dina(n11157), .dinb(n11151), .dout(n11332));
  jor  g11141(.dina(n11332), .dinb(n11153), .dout(n11333));
  jxor g11142(.dina(n11333), .dinb(n11331), .dout(n11334));
  jand g11143(.dina(n11193), .dinb(n11190), .dout(n11335));
  jnot g11144(.din(n11335), .dout(n11336));
  jand g11145(.dina(n11336), .dinb(n11196), .dout(n11337));
  jxor g11146(.dina(n11337), .dinb(n11334), .dout(n11338));
  jnot g11147(.din(n11338), .dout(n11339));
  jor  g11148(.dina(n11285), .dinb(n11277), .dout(n11340));
  jand g11149(.dina(n11286), .dinb(n11260), .dout(n11341));
  jnot g11150(.din(n11341), .dout(n11342));
  jand g11151(.dina(n11342), .dinb(n11340), .dout(n11343));
  jxor g11152(.dina(n11343), .dinb(n11339), .dout(n11344));
  jand g11153(.dina(n11293), .dinb(n11290), .dout(n11345));
  jand g11154(.dina(n11296), .dinb(n11294), .dout(n11346));
  jor  g11155(.dina(n11346), .dinb(n11345), .dout(n11347));
  jand g11156(.dina(\a[63] ), .dinb(\a[16] ), .dout(n11348));
  jand g11157(.dina(\a[45] ), .dinb(\a[34] ), .dout(n11349));
  jand g11158(.dina(\a[44] ), .dinb(\a[35] ), .dout(n11350));
  jor  g11159(.dina(n11350), .dinb(n11349), .dout(n11351));
  jand g11160(.dina(n4812), .dinb(n2845), .dout(n11352));
  jnot g11161(.din(n11352), .dout(n11353));
  jand g11162(.dina(n11353), .dinb(n11351), .dout(n11354));
  jxor g11163(.dina(n11354), .dinb(n11348), .dout(n11355));
  jand g11164(.dina(\a[43] ), .dinb(\a[36] ), .dout(n11356));
  jand g11165(.dina(\a[56] ), .dinb(\a[23] ), .dout(n11357));
  jand g11166(.dina(\a[52] ), .dinb(\a[27] ), .dout(n11358));
  jxor g11167(.dina(n11358), .dinb(n11357), .dout(n11359));
  jxor g11168(.dina(n11359), .dinb(n11356), .dout(n11360));
  jxor g11169(.dina(n11360), .dinb(n11355), .dout(n11361));
  jxor g11170(.dina(n11361), .dinb(n11347), .dout(n11362));
  jxor g11171(.dina(n11362), .dinb(n11344), .dout(n11363));
  jxor g11172(.dina(n11363), .dinb(n11329), .dout(n11364));
  jand g11173(.dina(n11186), .dinb(n11178), .dout(n11365));
  jnot g11174(.din(n11365), .dout(n11366));
  jor  g11175(.dina(n11198), .dinb(n11188), .dout(n11367));
  jand g11176(.dina(n11367), .dinb(n11366), .dout(n11368));
  jnot g11177(.din(n11368), .dout(n11369));
  jand g11178(.dina(n11283), .dinb(n11278), .dout(n11370));
  jor  g11179(.dina(n11370), .dinb(n11281), .dout(n11371));
  jand g11180(.dina(\a[61] ), .dinb(\a[18] ), .dout(n11372));
  jxor g11181(.dina(n11372), .dinb(n11272), .dout(n11373));
  jxor g11182(.dina(n11373), .dinb(n11371), .dout(n11374));
  jand g11183(.dina(n11185), .dinb(n11179), .dout(n11375));
  jor  g11184(.dina(n11375), .dinb(n11183), .dout(n11376));
  jand g11185(.dina(n11177), .dinb(n11172), .dout(n11377));
  jor  g11186(.dina(n11377), .dinb(n11175), .dout(n11378));
  jand g11187(.dina(n11165), .dinb(n11163), .dout(n11379));
  jnot g11188(.din(n11379), .dout(n11380));
  jand g11189(.dina(n11380), .dinb(n11168), .dout(n11381));
  jxor g11190(.dina(n11381), .dinb(n11378), .dout(n11382));
  jxor g11191(.dina(n11382), .dinb(n11376), .dout(n11383));
  jxor g11192(.dina(n11383), .dinb(n11374), .dout(n11384));
  jxor g11193(.dina(n11384), .dinb(n11369), .dout(n11385));
  jxor g11194(.dina(n11385), .dinb(n11364), .dout(n11386));
  jxor g11195(.dina(n11386), .dinb(n11326), .dout(n11387));
  jand g11196(.dina(n11201), .dinb(n11139), .dout(n11388));
  jand g11197(.dina(n11202), .dinb(n11136), .dout(n11389));
  jor  g11198(.dina(n11389), .dinb(n11388), .dout(n11390));
  jxor g11199(.dina(n11390), .dinb(n11387), .dout(n11391));
  jor  g11200(.dina(n11228), .dinb(n11224), .dout(n11392));
  jand g11201(.dina(n11255), .dinb(n11229), .dout(n11393));
  jnot g11202(.din(n11393), .dout(n11394));
  jand g11203(.dina(n11394), .dinb(n11392), .dout(n11395));
  jnot g11204(.din(n11395), .dout(n11396));
  jand g11205(.dina(n11253), .dinb(n11250), .dout(n11397));
  jand g11206(.dina(n11254), .dinb(n11241), .dout(n11398));
  jor  g11207(.dina(n11398), .dinb(n11397), .dout(n11399));
  jand g11208(.dina(\a[42] ), .dinb(\a[37] ), .dout(n11400));
  jnot g11209(.din(n11400), .dout(n11401));
  jand g11210(.dina(n11262), .dinb(n5246), .dout(n11402));
  jnot g11211(.din(n11402), .dout(n11403));
  jand g11212(.dina(n11400), .dinb(n3665), .dout(n11404));
  jand g11213(.dina(\a[42] ), .dinb(\a[38] ), .dout(n11405));
  jand g11214(.dina(n11405), .dinb(n5046), .dout(n11406));
  jor  g11215(.dina(n11406), .dinb(n11404), .dout(n11407));
  jand g11216(.dina(n11407), .dinb(n11403), .dout(n11408));
  jor  g11217(.dina(n11408), .dinb(n11401), .dout(n11409));
  jor  g11218(.dina(n11407), .dinb(n11402), .dout(n11410));
  jnot g11219(.din(n11410), .dout(n11411));
  jor  g11220(.dina(n11267), .dinb(n3665), .dout(n11412));
  jand g11221(.dina(n11412), .dinb(n11411), .dout(n11413));
  jnot g11222(.din(n11413), .dout(n11414));
  jand g11223(.dina(n11414), .dinb(n11409), .dout(n11415));
  jand g11224(.dina(\a[55] ), .dinb(\a[24] ), .dout(n11416));
  jand g11225(.dina(n7559), .dinb(n2128), .dout(n11417));
  jnot g11226(.din(n11417), .dout(n11418));
  jand g11227(.dina(\a[54] ), .dinb(\a[25] ), .dout(n11419));
  jand g11228(.dina(\a[53] ), .dinb(\a[26] ), .dout(n11420));
  jor  g11229(.dina(n11420), .dinb(n11419), .dout(n11421));
  jand g11230(.dina(n11421), .dinb(n11418), .dout(n11422));
  jxor g11231(.dina(n11422), .dinb(n11416), .dout(n11423));
  jnot g11232(.din(n11423), .dout(n11424));
  jxor g11233(.dina(n11424), .dinb(n11415), .dout(n11425));
  jand g11234(.dina(\a[51] ), .dinb(\a[28] ), .dout(n11426));
  jand g11235(.dina(n6557), .dinb(\a[62] ), .dout(n11427));
  jnot g11236(.din(n11427), .dout(n11428));
  jand g11237(.dina(\a[62] ), .dinb(\a[17] ), .dout(n11429));
  jor  g11238(.dina(n11429), .dinb(\a[40] ), .dout(n11430));
  jand g11239(.dina(n11430), .dinb(n11428), .dout(n11431));
  jxor g11240(.dina(n11431), .dinb(n11426), .dout(n11432));
  jxor g11241(.dina(n11432), .dinb(n11425), .dout(n11433));
  jand g11242(.dina(\a[60] ), .dinb(\a[19] ), .dout(n11434));
  jand g11243(.dina(\a[59] ), .dinb(\a[21] ), .dout(n11435));
  jand g11244(.dina(n11435), .dinb(n11172), .dout(n11436));
  jnot g11245(.din(n11436), .dout(n11437));
  jand g11246(.dina(\a[59] ), .dinb(\a[20] ), .dout(n11438));
  jand g11247(.dina(\a[58] ), .dinb(\a[21] ), .dout(n11439));
  jor  g11248(.dina(n11439), .dinb(n11438), .dout(n11440));
  jand g11249(.dina(n11440), .dinb(n11437), .dout(n11441));
  jxor g11250(.dina(n11441), .dinb(n11434), .dout(n11442));
  jand g11251(.dina(\a[57] ), .dinb(\a[22] ), .dout(n11443));
  jand g11252(.dina(\a[50] ), .dinb(\a[30] ), .dout(n11444));
  jand g11253(.dina(n11444), .dinb(n11156), .dout(n11445));
  jnot g11254(.din(n11445), .dout(n11446));
  jand g11255(.dina(\a[49] ), .dinb(\a[30] ), .dout(n11447));
  jor  g11256(.dina(n11447), .dinb(n11152), .dout(n11448));
  jand g11257(.dina(n11448), .dinb(n11446), .dout(n11449));
  jxor g11258(.dina(n11449), .dinb(n11443), .dout(n11450));
  jxor g11259(.dina(n11450), .dinb(n11442), .dout(n11451));
  jnot g11260(.din(n11451), .dout(n11452));
  jand g11261(.dina(\a[48] ), .dinb(\a[31] ), .dout(n11453));
  jnot g11262(.din(n11453), .dout(n11454));
  jand g11263(.dina(\a[47] ), .dinb(\a[33] ), .dout(n11455));
  jand g11264(.dina(n11455), .dinb(n11179), .dout(n11456));
  jnot g11265(.din(n11456), .dout(n11457));
  jand g11266(.dina(\a[47] ), .dinb(\a[32] ), .dout(n11458));
  jor  g11267(.dina(n11458), .dinb(n5007), .dout(n11459));
  jand g11268(.dina(n11459), .dinb(n11457), .dout(n11460));
  jxor g11269(.dina(n11460), .dinb(n11454), .dout(n11461));
  jxor g11270(.dina(n11461), .dinb(n11452), .dout(n11462));
  jxor g11271(.dina(n11462), .dinb(n11433), .dout(n11463));
  jxor g11272(.dina(n11463), .dinb(n11399), .dout(n11464));
  jxor g11273(.dina(n11464), .dinb(n11396), .dout(n11465));
  jand g11274(.dina(n11245), .dinb(n11242), .dout(n11466));
  jand g11275(.dina(n11249), .dinb(n11246), .dout(n11467));
  jor  g11276(.dina(n11467), .dinb(n11466), .dout(n11468));
  jand g11277(.dina(n11236), .dinb(n11233), .dout(n11469));
  jand g11278(.dina(n11240), .dinb(n11237), .dout(n11470));
  jor  g11279(.dina(n11470), .dinb(n11469), .dout(n11471));
  jxor g11280(.dina(n11471), .dinb(n11468), .dout(n11472));
  jnot g11281(.din(n11472), .dout(n11473));
  jand g11282(.dina(n11159), .dinb(n11150), .dout(n11474));
  jnot g11283(.din(n11474), .dout(n11475));
  jor  g11284(.dina(n11170), .dinb(n11161), .dout(n11476));
  jand g11285(.dina(n11476), .dinb(n11475), .dout(n11477));
  jxor g11286(.dina(n11477), .dinb(n11473), .dout(n11478));
  jnot g11287(.din(n11478), .dout(n11479));
  jor  g11288(.dina(n11217), .dinb(n11213), .dout(n11480));
  jor  g11289(.dina(n11222), .dinb(n11219), .dout(n11481));
  jand g11290(.dina(n11481), .dinb(n11480), .dout(n11482));
  jxor g11291(.dina(n11482), .dinb(n11479), .dout(n11483));
  jand g11292(.dina(n11300), .dinb(n11297), .dout(n11484));
  jand g11293(.dina(n11301), .dinb(n11287), .dout(n11485));
  jor  g11294(.dina(n11485), .dinb(n11484), .dout(n11486));
  jxor g11295(.dina(n11486), .dinb(n11483), .dout(n11487));
  jxor g11296(.dina(n11487), .dinb(n11465), .dout(n11488));
  jand g11297(.dina(n11256), .dinb(n11210), .dout(n11489));
  jand g11298(.dina(n11310), .dinb(n11257), .dout(n11490));
  jor  g11299(.dina(n11490), .dinb(n11489), .dout(n11491));
  jxor g11300(.dina(n11491), .dinb(n11488), .dout(n11492));
  jxor g11301(.dina(n11492), .dinb(n11391), .dout(n11493));
  jand g11302(.dina(n11493), .dinb(n11323), .dout(n11494));
  jor  g11303(.dina(n11493), .dinb(n11323), .dout(n11495));
  jnot g11304(.din(n11495), .dout(n11496));
  jor  g11305(.dina(n11496), .dinb(n11494), .dout(n11497));
  jnot g11306(.din(n11313), .dout(n11498));
  jor  g11307(.dina(n11319), .dinb(n11315), .dout(n11499));
  jand g11308(.dina(n11499), .dinb(n11498), .dout(n11500));
  jxor g11309(.dina(n11500), .dinb(n11497), .dout(\asquared[80] ));
  jand g11310(.dina(n11491), .dinb(n11488), .dout(n11502));
  jand g11311(.dina(n11492), .dinb(n11391), .dout(n11503));
  jor  g11312(.dina(n11503), .dinb(n11502), .dout(n11504));
  jand g11313(.dina(n11386), .dinb(n11326), .dout(n11505));
  jand g11314(.dina(n11390), .dinb(n11387), .dout(n11506));
  jor  g11315(.dina(n11506), .dinb(n11505), .dout(n11507));
  jand g11316(.dina(n11363), .dinb(n11329), .dout(n11508));
  jand g11317(.dina(n11385), .dinb(n11364), .dout(n11509));
  jor  g11318(.dina(n11509), .dinb(n11508), .dout(n11510));
  jor  g11319(.dina(n11482), .dinb(n11479), .dout(n11511));
  jand g11320(.dina(n11486), .dinb(n11483), .dout(n11512));
  jnot g11321(.din(n11512), .dout(n11513));
  jand g11322(.dina(n11513), .dinb(n11511), .dout(n11514));
  jnot g11323(.din(n11514), .dout(n11515));
  jand g11324(.dina(\a[59] ), .dinb(\a[22] ), .dout(n11516));
  jand g11325(.dina(n11516), .dinb(n11439), .dout(n11517));
  jnot g11326(.din(n11517), .dout(n11518));
  jand g11327(.dina(\a[58] ), .dinb(\a[22] ), .dout(n11519));
  jor  g11328(.dina(n11519), .dinb(n11435), .dout(n11520));
  jand g11329(.dina(n11520), .dinb(n11518), .dout(n11521));
  jand g11330(.dina(\a[60] ), .dinb(\a[20] ), .dout(n11522));
  jxor g11331(.dina(n11522), .dinb(n11521), .dout(n11523));
  jxor g11332(.dina(n11523), .dinb(n11410), .dout(n11524));
  jnot g11333(.din(n11524), .dout(n11525));
  jnot g11334(.din(n11444), .dout(n11526));
  jand g11335(.dina(n7729), .dinb(n3269), .dout(n11527));
  jnot g11336(.din(n11527), .dout(n11528));
  jand g11337(.dina(\a[49] ), .dinb(\a[31] ), .dout(n11529));
  jand g11338(.dina(\a[48] ), .dinb(\a[32] ), .dout(n11530));
  jor  g11339(.dina(n11530), .dinb(n11529), .dout(n11531));
  jand g11340(.dina(n11531), .dinb(n11528), .dout(n11532));
  jxor g11341(.dina(n11532), .dinb(n11526), .dout(n11533));
  jxor g11342(.dina(n11533), .dinb(n11525), .dout(n11534));
  jand g11343(.dina(\a[57] ), .dinb(\a[23] ), .dout(n11535));
  jand g11344(.dina(\a[56] ), .dinb(\a[24] ), .dout(n11536));
  jand g11345(.dina(\a[54] ), .dinb(\a[26] ), .dout(n11537));
  jor  g11346(.dina(n11537), .dinb(n11536), .dout(n11538));
  jand g11347(.dina(n11191), .dinb(n2022), .dout(n11539));
  jnot g11348(.din(n11539), .dout(n11540));
  jand g11349(.dina(n11540), .dinb(n11538), .dout(n11541));
  jxor g11350(.dina(n11541), .dinb(n11535), .dout(n11542));
  jnot g11351(.din(n11542), .dout(n11543));
  jand g11352(.dina(\a[55] ), .dinb(\a[25] ), .dout(n11544));
  jnot g11353(.din(n11544), .dout(n11545));
  jand g11354(.dina(\a[43] ), .dinb(\a[38] ), .dout(n11546));
  jand g11355(.dina(n11546), .dinb(n11400), .dout(n11547));
  jnot g11356(.din(n11547), .dout(n11548));
  jand g11357(.dina(\a[43] ), .dinb(\a[37] ), .dout(n11549));
  jor  g11358(.dina(n11549), .dinb(n11405), .dout(n11550));
  jand g11359(.dina(n11550), .dinb(n11548), .dout(n11551));
  jxor g11360(.dina(n11551), .dinb(n11545), .dout(n11552));
  jxor g11361(.dina(n11552), .dinb(n11543), .dout(n11553));
  jnot g11362(.din(n11553), .dout(n11554));
  jnot g11363(.din(n5246), .dout(n11555));
  jand g11364(.dina(n7165), .dinb(n2042), .dout(n11556));
  jnot g11365(.din(n11556), .dout(n11557));
  jand g11366(.dina(\a[53] ), .dinb(\a[27] ), .dout(n11558));
  jand g11367(.dina(\a[52] ), .dinb(\a[28] ), .dout(n11559));
  jor  g11368(.dina(n11559), .dinb(n11558), .dout(n11560));
  jand g11369(.dina(n11560), .dinb(n11557), .dout(n11561));
  jxor g11370(.dina(n11561), .dinb(n11555), .dout(n11562));
  jxor g11371(.dina(n11562), .dinb(n11554), .dout(n11563));
  jxor g11372(.dina(n11563), .dinb(n11534), .dout(n11564));
  jand g11373(.dina(\a[63] ), .dinb(\a[17] ), .dout(n11565));
  jand g11374(.dina(\a[51] ), .dinb(\a[29] ), .dout(n11566));
  jxor g11375(.dina(n11566), .dinb(n11565), .dout(n11567));
  jxor g11376(.dina(n11567), .dinb(n11455), .dout(n11568));
  jnot g11377(.din(n11568), .dout(n11569));
  jand g11378(.dina(\a[46] ), .dinb(\a[34] ), .dout(n11570));
  jnot g11379(.din(n11570), .dout(n11571));
  jand g11380(.dina(n4812), .dinb(n3243), .dout(n11572));
  jnot g11381(.din(n11572), .dout(n11573));
  jand g11382(.dina(\a[44] ), .dinb(\a[36] ), .dout(n11574));
  jor  g11383(.dina(n11574), .dinb(n4983), .dout(n11575));
  jand g11384(.dina(n11575), .dinb(n11573), .dout(n11576));
  jxor g11385(.dina(n11576), .dinb(n11571), .dout(n11577));
  jxor g11386(.dina(n11577), .dinb(n11569), .dout(n11578));
  jand g11387(.dina(n8702), .dinb(n1024), .dout(n11579));
  jnot g11388(.din(n11579), .dout(n11580));
  jand g11389(.dina(\a[62] ), .dinb(\a[18] ), .dout(n11581));
  jand g11390(.dina(\a[61] ), .dinb(\a[19] ), .dout(n11582));
  jor  g11391(.dina(n11582), .dinb(n11581), .dout(n11583));
  jand g11392(.dina(n11583), .dinb(n11580), .dout(n11584));
  jor  g11393(.dina(n11427), .dinb(n11426), .dout(n11585));
  jand g11394(.dina(n11585), .dinb(n11430), .dout(n11586));
  jxor g11395(.dina(n11586), .dinb(n11584), .dout(n11587));
  jxor g11396(.dina(n11587), .dinb(n11578), .dout(n11588));
  jxor g11397(.dina(n11588), .dinb(n11564), .dout(n11589));
  jxor g11398(.dina(n11589), .dinb(n11515), .dout(n11590));
  jxor g11399(.dina(n11590), .dinb(n11510), .dout(n11591));
  jxor g11400(.dina(n11591), .dinb(n11507), .dout(n11592));
  jand g11401(.dina(n11464), .dinb(n11396), .dout(n11593));
  jand g11402(.dina(n11487), .dinb(n11465), .dout(n11594));
  jor  g11403(.dina(n11594), .dinb(n11593), .dout(n11595));
  jand g11404(.dina(n11462), .dinb(n11433), .dout(n11596));
  jand g11405(.dina(n11463), .dinb(n11399), .dout(n11597));
  jor  g11406(.dina(n11597), .dinb(n11596), .dout(n11598));
  jand g11407(.dina(n11358), .dinb(n11357), .dout(n11599));
  jand g11408(.dina(n11359), .dinb(n11356), .dout(n11600));
  jor  g11409(.dina(n11600), .dinb(n11599), .dout(n11601));
  jand g11410(.dina(n11354), .dinb(n11348), .dout(n11602));
  jor  g11411(.dina(n11602), .dinb(n11352), .dout(n11603));
  jand g11412(.dina(n11422), .dinb(n11416), .dout(n11604));
  jor  g11413(.dina(n11604), .dinb(n11417), .dout(n11605));
  jxor g11414(.dina(n11605), .dinb(n11603), .dout(n11606));
  jxor g11415(.dina(n11606), .dinb(n11601), .dout(n11607));
  jand g11416(.dina(n11360), .dinb(n11355), .dout(n11608));
  jand g11417(.dina(n11361), .dinb(n11347), .dout(n11609));
  jor  g11418(.dina(n11609), .dinb(n11608), .dout(n11610));
  jxor g11419(.dina(n11610), .dinb(n11607), .dout(n11611));
  jnot g11420(.din(n11611), .dout(n11612));
  jand g11421(.dina(n11471), .dinb(n11468), .dout(n11613));
  jnot g11422(.din(n11613), .dout(n11614));
  jor  g11423(.dina(n11477), .dinb(n11473), .dout(n11615));
  jand g11424(.dina(n11615), .dinb(n11614), .dout(n11616));
  jxor g11425(.dina(n11616), .dinb(n11612), .dout(n11617));
  jxor g11426(.dina(n11617), .dinb(n11598), .dout(n11618));
  jand g11427(.dina(n11441), .dinb(n11434), .dout(n11619));
  jor  g11428(.dina(n11619), .dinb(n11436), .dout(n11620));
  jor  g11429(.dina(n11445), .dinb(n11443), .dout(n11621));
  jand g11430(.dina(n11621), .dinb(n11448), .dout(n11622));
  jxor g11431(.dina(n11622), .dinb(n11620), .dout(n11623));
  jand g11432(.dina(n11457), .dinb(n11454), .dout(n11624));
  jnot g11433(.din(n11624), .dout(n11625));
  jand g11434(.dina(n11625), .dinb(n11459), .dout(n11626));
  jxor g11435(.dina(n11626), .dinb(n11623), .dout(n11627));
  jor  g11436(.dina(n11424), .dinb(n11415), .dout(n11628));
  jand g11437(.dina(n11432), .dinb(n11425), .dout(n11629));
  jnot g11438(.din(n11629), .dout(n11630));
  jand g11439(.dina(n11630), .dinb(n11628), .dout(n11631));
  jand g11440(.dina(n11450), .dinb(n11442), .dout(n11632));
  jnot g11441(.din(n11632), .dout(n11633));
  jor  g11442(.dina(n11461), .dinb(n11452), .dout(n11634));
  jand g11443(.dina(n11634), .dinb(n11633), .dout(n11635));
  jxor g11444(.dina(n11635), .dinb(n11631), .dout(n11636));
  jxor g11445(.dina(n11636), .dinb(n11627), .dout(n11637));
  jxor g11446(.dina(n11637), .dinb(n11618), .dout(n11638));
  jand g11447(.dina(n11333), .dinb(n11331), .dout(n11639));
  jand g11448(.dina(n11337), .dinb(n11334), .dout(n11640));
  jor  g11449(.dina(n11640), .dinb(n11639), .dout(n11641));
  jand g11450(.dina(n11381), .dinb(n11378), .dout(n11642));
  jand g11451(.dina(n11382), .dinb(n11376), .dout(n11643));
  jor  g11452(.dina(n11643), .dinb(n11642), .dout(n11644));
  jxor g11453(.dina(n11644), .dinb(n11641), .dout(n11645));
  jand g11454(.dina(n11372), .dinb(n11272), .dout(n11646));
  jand g11455(.dina(n11373), .dinb(n11371), .dout(n11647));
  jor  g11456(.dina(n11647), .dinb(n11646), .dout(n11648));
  jxor g11457(.dina(n11648), .dinb(n11645), .dout(n11649));
  jor  g11458(.dina(n11343), .dinb(n11339), .dout(n11650));
  jand g11459(.dina(n11362), .dinb(n11344), .dout(n11651));
  jnot g11460(.din(n11651), .dout(n11652));
  jand g11461(.dina(n11652), .dinb(n11650), .dout(n11653));
  jnot g11462(.din(n11653), .dout(n11654));
  jand g11463(.dina(n11383), .dinb(n11374), .dout(n11655));
  jand g11464(.dina(n11384), .dinb(n11369), .dout(n11656));
  jor  g11465(.dina(n11656), .dinb(n11655), .dout(n11657));
  jxor g11466(.dina(n11657), .dinb(n11654), .dout(n11658));
  jxor g11467(.dina(n11658), .dinb(n11649), .dout(n11659));
  jxor g11468(.dina(n11659), .dinb(n11638), .dout(n11660));
  jxor g11469(.dina(n11660), .dinb(n11595), .dout(n11661));
  jxor g11470(.dina(n11661), .dinb(n11592), .dout(n11662));
  jnot g11471(.din(n11662), .dout(n11663));
  jxor g11472(.dina(n11663), .dinb(n11504), .dout(n11664));
  jnot g11473(.din(n11494), .dout(n11665));
  jor  g11474(.dina(n11500), .dinb(n11496), .dout(n11666));
  jand g11475(.dina(n11666), .dinb(n11665), .dout(n11667));
  jxor g11476(.dina(n11667), .dinb(n11664), .dout(\asquared[81] ));
  jand g11477(.dina(n11591), .dinb(n11507), .dout(n11669));
  jand g11478(.dina(n11661), .dinb(n11592), .dout(n11670));
  jor  g11479(.dina(n11670), .dinb(n11669), .dout(n11671));
  jand g11480(.dina(n11659), .dinb(n11638), .dout(n11672));
  jand g11481(.dina(n11660), .dinb(n11595), .dout(n11673));
  jor  g11482(.dina(n11673), .dinb(n11672), .dout(n11674));
  jand g11483(.dina(n11617), .dinb(n11598), .dout(n11675));
  jand g11484(.dina(n11637), .dinb(n11618), .dout(n11676));
  jor  g11485(.dina(n11676), .dinb(n11675), .dout(n11677));
  jand g11486(.dina(n11657), .dinb(n11654), .dout(n11678));
  jand g11487(.dina(n11658), .dinb(n11649), .dout(n11679));
  jor  g11488(.dina(n11679), .dinb(n11678), .dout(n11680));
  jand g11489(.dina(n11644), .dinb(n11641), .dout(n11681));
  jand g11490(.dina(n11648), .dinb(n11645), .dout(n11682));
  jor  g11491(.dina(n11682), .dinb(n11681), .dout(n11683));
  jand g11492(.dina(\a[62] ), .dinb(\a[19] ), .dout(n11684));
  jnot g11493(.din(\a[40] ), .dout(n11685));
  jand g11494(.dina(\a[41] ), .dinb(n11685), .dout(n11686));
  jxor g11495(.dina(n11686), .dinb(n11684), .dout(n11687));
  jand g11496(.dina(\a[58] ), .dinb(\a[56] ), .dout(n11688));
  jand g11497(.dina(n11688), .dinb(n4755), .dout(n11689));
  jnot g11498(.din(n11689), .dout(n11690));
  jand g11499(.dina(\a[56] ), .dinb(\a[25] ), .dout(n11691));
  jand g11500(.dina(\a[58] ), .dinb(\a[23] ), .dout(n11692));
  jor  g11501(.dina(n11692), .dinb(n11691), .dout(n11693));
  jand g11502(.dina(n11693), .dinb(n11690), .dout(n11694));
  jxor g11503(.dina(n11694), .dinb(n11516), .dout(n11695));
  jxor g11504(.dina(n11695), .dinb(n11687), .dout(n11696));
  jand g11505(.dina(\a[57] ), .dinb(\a[24] ), .dout(n11697));
  jand g11506(.dina(n5316), .dinb(n3634), .dout(n11698));
  jnot g11507(.din(n11698), .dout(n11699));
  jand g11508(.dina(\a[48] ), .dinb(\a[33] ), .dout(n11700));
  jand g11509(.dina(\a[47] ), .dinb(\a[34] ), .dout(n11701));
  jor  g11510(.dina(n11701), .dinb(n11700), .dout(n11702));
  jand g11511(.dina(n11702), .dinb(n11699), .dout(n11703));
  jxor g11512(.dina(n11703), .dinb(n11697), .dout(n11704));
  jxor g11513(.dina(n11704), .dinb(n11696), .dout(n11705));
  jxor g11514(.dina(n11705), .dinb(n11683), .dout(n11706));
  jand g11515(.dina(\a[53] ), .dinb(\a[28] ), .dout(n11707));
  jand g11516(.dina(\a[52] ), .dinb(\a[29] ), .dout(n11708));
  jor  g11517(.dina(n11708), .dinb(n11707), .dout(n11709));
  jand g11518(.dina(n7165), .dinb(n2653), .dout(n11710));
  jnot g11519(.din(n11710), .dout(n11711));
  jand g11520(.dina(n11263), .dinb(\a[29] ), .dout(n11712));
  jand g11521(.dina(n11712), .dinb(\a[55] ), .dout(n11713));
  jand g11522(.dina(\a[55] ), .dinb(\a[26] ), .dout(n11714));
  jand g11523(.dina(n11714), .dinb(n11707), .dout(n11715));
  jor  g11524(.dina(n11715), .dinb(n11713), .dout(n11716));
  jnot g11525(.din(n11716), .dout(n11717));
  jand g11526(.dina(n11717), .dinb(n11711), .dout(n11718));
  jand g11527(.dina(n11718), .dinb(n11709), .dout(n11719));
  jand g11528(.dina(n11716), .dinb(n11711), .dout(n11720));
  jnot g11529(.din(n11720), .dout(n11721));
  jand g11530(.dina(n11721), .dinb(n11714), .dout(n11722));
  jor  g11531(.dina(n11722), .dinb(n11719), .dout(n11723));
  jand g11532(.dina(\a[46] ), .dinb(\a[35] ), .dout(n11724));
  jnot g11533(.din(n11724), .dout(n11725));
  jand g11534(.dina(n4812), .dinb(n3138), .dout(n11726));
  jnot g11535(.din(n11726), .dout(n11727));
  jand g11536(.dina(n5382), .dinb(n4983), .dout(n11728));
  jand g11537(.dina(\a[44] ), .dinb(\a[37] ), .dout(n11729));
  jand g11538(.dina(n11729), .dinb(n11724), .dout(n11730));
  jor  g11539(.dina(n11730), .dinb(n11728), .dout(n11731));
  jand g11540(.dina(n11731), .dinb(n11727), .dout(n11732));
  jor  g11541(.dina(n11732), .dinb(n11725), .dout(n11733));
  jand g11542(.dina(\a[45] ), .dinb(\a[36] ), .dout(n11734));
  jor  g11543(.dina(n11734), .dinb(n11729), .dout(n11735));
  jor  g11544(.dina(n11731), .dinb(n11726), .dout(n11736));
  jnot g11545(.din(n11736), .dout(n11737));
  jand g11546(.dina(n11737), .dinb(n11735), .dout(n11738));
  jnot g11547(.din(n11738), .dout(n11739));
  jand g11548(.dina(n11739), .dinb(n11733), .dout(n11740));
  jand g11549(.dina(\a[63] ), .dinb(\a[18] ), .dout(n11741));
  jand g11550(.dina(\a[61] ), .dinb(\a[21] ), .dout(n11742));
  jand g11551(.dina(n11742), .dinb(n11522), .dout(n11743));
  jnot g11552(.din(n11743), .dout(n11744));
  jand g11553(.dina(\a[61] ), .dinb(\a[20] ), .dout(n11745));
  jand g11554(.dina(\a[60] ), .dinb(\a[21] ), .dout(n11746));
  jor  g11555(.dina(n11746), .dinb(n11745), .dout(n11747));
  jand g11556(.dina(n11747), .dinb(n11744), .dout(n11748));
  jxor g11557(.dina(n11748), .dinb(n11741), .dout(n11749));
  jnot g11558(.din(n11749), .dout(n11750));
  jxor g11559(.dina(n11750), .dinb(n11740), .dout(n11751));
  jxor g11560(.dina(n11751), .dinb(n11723), .dout(n11752));
  jxor g11561(.dina(n11752), .dinb(n11706), .dout(n11753));
  jxor g11562(.dina(n11753), .dinb(n11680), .dout(n11754));
  jxor g11563(.dina(n11754), .dinb(n11677), .dout(n11755));
  jxor g11564(.dina(n11755), .dinb(n11674), .dout(n11756));
  jand g11565(.dina(n11563), .dinb(n11534), .dout(n11757));
  jand g11566(.dina(n11588), .dinb(n11564), .dout(n11758));
  jor  g11567(.dina(n11758), .dinb(n11757), .dout(n11759));
  jand g11568(.dina(n11566), .dinb(n11565), .dout(n11760));
  jand g11569(.dina(n11567), .dinb(n11455), .dout(n11761));
  jor  g11570(.dina(n11761), .dinb(n11760), .dout(n11762));
  jand g11571(.dina(n11528), .dinb(n11526), .dout(n11763));
  jnot g11572(.din(n11763), .dout(n11764));
  jand g11573(.dina(n11764), .dinb(n11531), .dout(n11765));
  jxor g11574(.dina(n11765), .dinb(n11762), .dout(n11766));
  jand g11575(.dina(n11522), .dinb(n11521), .dout(n11767));
  jor  g11576(.dina(n11767), .dinb(n11517), .dout(n11768));
  jxor g11577(.dina(n11768), .dinb(n11766), .dout(n11769));
  jnot g11578(.din(n11769), .dout(n11770));
  jor  g11579(.dina(n11577), .dinb(n11569), .dout(n11771));
  jand g11580(.dina(n11587), .dinb(n11578), .dout(n11772));
  jnot g11581(.din(n11772), .dout(n11773));
  jand g11582(.dina(n11773), .dinb(n11771), .dout(n11774));
  jxor g11583(.dina(n11774), .dinb(n11770), .dout(n11775));
  jand g11584(.dina(n11586), .dinb(n11584), .dout(n11776));
  jor  g11585(.dina(n11776), .dinb(n11579), .dout(n11777));
  jand g11586(.dina(n11573), .dinb(n11571), .dout(n11778));
  jnot g11587(.din(n11778), .dout(n11779));
  jand g11588(.dina(n11779), .dinb(n11575), .dout(n11780));
  jxor g11589(.dina(n11780), .dinb(n11777), .dout(n11781));
  jnot g11590(.din(n11781), .dout(n11782));
  jand g11591(.dina(\a[51] ), .dinb(\a[30] ), .dout(n11783));
  jnot g11592(.din(n11783), .dout(n11784));
  jand g11593(.dina(\a[50] ), .dinb(\a[32] ), .dout(n11785));
  jand g11594(.dina(n11785), .dinb(n11529), .dout(n11786));
  jnot g11595(.din(n11786), .dout(n11787));
  jand g11596(.dina(\a[50] ), .dinb(\a[31] ), .dout(n11788));
  jand g11597(.dina(\a[49] ), .dinb(\a[32] ), .dout(n11789));
  jor  g11598(.dina(n11789), .dinb(n11788), .dout(n11790));
  jand g11599(.dina(n11790), .dinb(n11787), .dout(n11791));
  jxor g11600(.dina(n11791), .dinb(n11784), .dout(n11792));
  jxor g11601(.dina(n11792), .dinb(n11782), .dout(n11793));
  jxor g11602(.dina(n11793), .dinb(n11775), .dout(n11794));
  jxor g11603(.dina(n11794), .dinb(n11759), .dout(n11795));
  jand g11604(.dina(n11541), .dinb(n11535), .dout(n11796));
  jor  g11605(.dina(n11796), .dinb(n11539), .dout(n11797));
  jand g11606(.dina(n11557), .dinb(n11555), .dout(n11798));
  jnot g11607(.din(n11798), .dout(n11799));
  jand g11608(.dina(n11799), .dinb(n11560), .dout(n11800));
  jand g11609(.dina(n11548), .dinb(n11545), .dout(n11801));
  jnot g11610(.din(n11801), .dout(n11802));
  jand g11611(.dina(n11802), .dinb(n11550), .dout(n11803));
  jxor g11612(.dina(n11803), .dinb(n11800), .dout(n11804));
  jxor g11613(.dina(n11804), .dinb(n11797), .dout(n11805));
  jor  g11614(.dina(n11552), .dinb(n11543), .dout(n11806));
  jor  g11615(.dina(n11562), .dinb(n11554), .dout(n11807));
  jand g11616(.dina(n11807), .dinb(n11806), .dout(n11808));
  jand g11617(.dina(n11523), .dinb(n11410), .dout(n11809));
  jnot g11618(.din(n11809), .dout(n11810));
  jor  g11619(.dina(n11533), .dinb(n11525), .dout(n11811));
  jand g11620(.dina(n11811), .dinb(n11810), .dout(n11812));
  jxor g11621(.dina(n11812), .dinb(n11808), .dout(n11813));
  jxor g11622(.dina(n11813), .dinb(n11805), .dout(n11814));
  jxor g11623(.dina(n11814), .dinb(n11795), .dout(n11815));
  jand g11624(.dina(n11589), .dinb(n11515), .dout(n11816));
  jand g11625(.dina(n11590), .dinb(n11510), .dout(n11817));
  jor  g11626(.dina(n11817), .dinb(n11816), .dout(n11818));
  jand g11627(.dina(n11605), .dinb(n11603), .dout(n11819));
  jand g11628(.dina(n11606), .dinb(n11601), .dout(n11820));
  jor  g11629(.dina(n11820), .dinb(n11819), .dout(n11821));
  jand g11630(.dina(n11622), .dinb(n11620), .dout(n11822));
  jand g11631(.dina(n11626), .dinb(n11623), .dout(n11823));
  jor  g11632(.dina(n11823), .dinb(n11822), .dout(n11824));
  jnot g11633(.din(n11824), .dout(n11825));
  jand g11634(.dina(\a[54] ), .dinb(\a[27] ), .dout(n11826));
  jnot g11635(.din(n11826), .dout(n11827));
  jand g11636(.dina(\a[43] ), .dinb(\a[39] ), .dout(n11828));
  jand g11637(.dina(n11828), .dinb(n11405), .dout(n11829));
  jnot g11638(.din(n11829), .dout(n11830));
  jand g11639(.dina(\a[42] ), .dinb(\a[39] ), .dout(n11831));
  jor  g11640(.dina(n11831), .dinb(n11546), .dout(n11832));
  jand g11641(.dina(n11832), .dinb(n11830), .dout(n11833));
  jxor g11642(.dina(n11833), .dinb(n11827), .dout(n11834));
  jxor g11643(.dina(n11834), .dinb(n11825), .dout(n11835));
  jxor g11644(.dina(n11835), .dinb(n11821), .dout(n11836));
  jand g11645(.dina(n11610), .dinb(n11607), .dout(n11837));
  jnot g11646(.din(n11837), .dout(n11838));
  jor  g11647(.dina(n11616), .dinb(n11612), .dout(n11839));
  jand g11648(.dina(n11839), .dinb(n11838), .dout(n11840));
  jor  g11649(.dina(n11635), .dinb(n11631), .dout(n11841));
  jand g11650(.dina(n11636), .dinb(n11627), .dout(n11842));
  jnot g11651(.din(n11842), .dout(n11843));
  jand g11652(.dina(n11843), .dinb(n11841), .dout(n11844));
  jxor g11653(.dina(n11844), .dinb(n11840), .dout(n11845));
  jxor g11654(.dina(n11845), .dinb(n11836), .dout(n11846));
  jxor g11655(.dina(n11846), .dinb(n11818), .dout(n11847));
  jxor g11656(.dina(n11847), .dinb(n11815), .dout(n11848));
  jxor g11657(.dina(n11848), .dinb(n11756), .dout(n11849));
  jand g11658(.dina(n11849), .dinb(n11671), .dout(n11850));
  jor  g11659(.dina(n11849), .dinb(n11671), .dout(n11851));
  jnot g11660(.din(n11851), .dout(n11852));
  jor  g11661(.dina(n11852), .dinb(n11850), .dout(n11853));
  jand g11662(.dina(n11662), .dinb(n11504), .dout(n11854));
  jnot g11663(.din(n11854), .dout(n11855));
  jnot g11664(.din(n11504), .dout(n11856));
  jand g11665(.dina(n11663), .dinb(n11856), .dout(n11857));
  jor  g11666(.dina(n11667), .dinb(n11857), .dout(n11858));
  jand g11667(.dina(n11858), .dinb(n11855), .dout(n11859));
  jxor g11668(.dina(n11859), .dinb(n11853), .dout(\asquared[82] ));
  jand g11669(.dina(n11755), .dinb(n11674), .dout(n11861));
  jand g11670(.dina(n11848), .dinb(n11756), .dout(n11862));
  jor  g11671(.dina(n11862), .dinb(n11861), .dout(n11863));
  jand g11672(.dina(n11846), .dinb(n11818), .dout(n11864));
  jand g11673(.dina(n11847), .dinb(n11815), .dout(n11865));
  jor  g11674(.dina(n11865), .dinb(n11864), .dout(n11866));
  jand g11675(.dina(n11794), .dinb(n11759), .dout(n11867));
  jand g11676(.dina(n11814), .dinb(n11795), .dout(n11868));
  jor  g11677(.dina(n11868), .dinb(n11867), .dout(n11869));
  jor  g11678(.dina(n11844), .dinb(n11840), .dout(n11870));
  jand g11679(.dina(n11845), .dinb(n11836), .dout(n11871));
  jnot g11680(.din(n11871), .dout(n11872));
  jand g11681(.dina(n11872), .dinb(n11870), .dout(n11873));
  jnot g11682(.din(n11873), .dout(n11874));
  jor  g11683(.dina(n11834), .dinb(n11825), .dout(n11875));
  jand g11684(.dina(n11835), .dinb(n11821), .dout(n11876));
  jnot g11685(.din(n11876), .dout(n11877));
  jand g11686(.dina(n11877), .dinb(n11875), .dout(n11878));
  jnot g11687(.din(n11878), .dout(n11879));
  jand g11688(.dina(\a[62] ), .dinb(\a[20] ), .dout(n11880));
  jand g11689(.dina(\a[51] ), .dinb(\a[31] ), .dout(n11881));
  jxor g11690(.dina(n11881), .dinb(n11742), .dout(n11882));
  jxor g11691(.dina(n11882), .dinb(n11880), .dout(n11883));
  jand g11692(.dina(n7729), .dinb(n3634), .dout(n11884));
  jnot g11693(.din(n11884), .dout(n11885));
  jand g11694(.dina(\a[49] ), .dinb(\a[33] ), .dout(n11886));
  jand g11695(.dina(\a[48] ), .dinb(\a[34] ), .dout(n11887));
  jor  g11696(.dina(n11887), .dinb(n11886), .dout(n11888));
  jand g11697(.dina(n11888), .dinb(n11885), .dout(n11889));
  jxor g11698(.dina(n11889), .dinb(n11785), .dout(n11890));
  jxor g11699(.dina(n11890), .dinb(n11883), .dout(n11891));
  jnot g11700(.din(n11891), .dout(n11892));
  jand g11701(.dina(\a[60] ), .dinb(\a[22] ), .dout(n11893));
  jnot g11702(.din(n11893), .dout(n11894));
  jand g11703(.dina(\a[59] ), .dinb(\a[24] ), .dout(n11895));
  jand g11704(.dina(n11895), .dinb(n11692), .dout(n11896));
  jnot g11705(.din(n11896), .dout(n11897));
  jand g11706(.dina(\a[58] ), .dinb(\a[24] ), .dout(n11898));
  jand g11707(.dina(\a[59] ), .dinb(\a[23] ), .dout(n11899));
  jor  g11708(.dina(n11899), .dinb(n11898), .dout(n11900));
  jand g11709(.dina(n11900), .dinb(n11897), .dout(n11901));
  jxor g11710(.dina(n11901), .dinb(n11894), .dout(n11902));
  jxor g11711(.dina(n11902), .dinb(n11892), .dout(n11903));
  jxor g11712(.dina(n11903), .dinb(n11879), .dout(n11904));
  jand g11713(.dina(\a[47] ), .dinb(\a[35] ), .dout(n11905));
  jand g11714(.dina(\a[46] ), .dinb(\a[37] ), .dout(n11906));
  jand g11715(.dina(n11906), .dinb(n11734), .dout(n11907));
  jnot g11716(.din(n11907), .dout(n11908));
  jand g11717(.dina(n11905), .dinb(n5196), .dout(n11909));
  jand g11718(.dina(\a[47] ), .dinb(\a[36] ), .dout(n11910));
  jand g11719(.dina(n11910), .dinb(n11724), .dout(n11911));
  jor  g11720(.dina(n11911), .dinb(n11909), .dout(n11912));
  jand g11721(.dina(n11912), .dinb(n11908), .dout(n11913));
  jnot g11722(.din(n11913), .dout(n11914));
  jand g11723(.dina(n11914), .dinb(n11905), .dout(n11915));
  jor  g11724(.dina(n11912), .dinb(n11907), .dout(n11916));
  jnot g11725(.din(n11916), .dout(n11917));
  jor  g11726(.dina(n5382), .dinb(n5196), .dout(n11918));
  jand g11727(.dina(n11918), .dinb(n11917), .dout(n11919));
  jor  g11728(.dina(n11919), .dinb(n11915), .dout(n11920));
  jand g11729(.dina(\a[56] ), .dinb(\a[26] ), .dout(n11921));
  jand g11730(.dina(\a[44] ), .dinb(\a[38] ), .dout(n11922));
  jor  g11731(.dina(n11922), .dinb(n11828), .dout(n11923));
  jand g11732(.dina(\a[44] ), .dinb(\a[39] ), .dout(n11924));
  jand g11733(.dina(n11924), .dinb(n11546), .dout(n11925));
  jnot g11734(.din(n11925), .dout(n11926));
  jand g11735(.dina(n11926), .dinb(n11923), .dout(n11927));
  jxor g11736(.dina(n11927), .dinb(n11921), .dout(n11928));
  jand g11737(.dina(\a[42] ), .dinb(\a[40] ), .dout(n11929));
  jand g11738(.dina(n7165), .dinb(n3294), .dout(n11930));
  jnot g11739(.din(n11930), .dout(n11931));
  jand g11740(.dina(\a[53] ), .dinb(\a[29] ), .dout(n11932));
  jand g11741(.dina(\a[52] ), .dinb(\a[30] ), .dout(n11933));
  jor  g11742(.dina(n11933), .dinb(n11932), .dout(n11934));
  jand g11743(.dina(n11934), .dinb(n11931), .dout(n11935));
  jxor g11744(.dina(n11935), .dinb(n11929), .dout(n11936));
  jxor g11745(.dina(n11936), .dinb(n11928), .dout(n11937));
  jxor g11746(.dina(n11937), .dinb(n11920), .dout(n11938));
  jxor g11747(.dina(n11938), .dinb(n11904), .dout(n11939));
  jxor g11748(.dina(n11939), .dinb(n11874), .dout(n11940));
  jxor g11749(.dina(n11940), .dinb(n11869), .dout(n11941));
  jxor g11750(.dina(n11941), .dinb(n11866), .dout(n11942));
  jand g11751(.dina(n11705), .dinb(n11683), .dout(n11943));
  jand g11752(.dina(n11752), .dinb(n11706), .dout(n11944));
  jor  g11753(.dina(n11944), .dinb(n11943), .dout(n11945));
  jnot g11754(.din(n11718), .dout(n11946));
  jand g11755(.dina(n11702), .dinb(n11697), .dout(n11947));
  jor  g11756(.dina(n11947), .dinb(n11698), .dout(n11948));
  jand g11757(.dina(n11787), .dinb(n11784), .dout(n11949));
  jnot g11758(.din(n11949), .dout(n11950));
  jand g11759(.dina(n11950), .dinb(n11790), .dout(n11951));
  jxor g11760(.dina(n11951), .dinb(n11948), .dout(n11952));
  jxor g11761(.dina(n11952), .dinb(n11946), .dout(n11953));
  jand g11762(.dina(n11748), .dinb(n11741), .dout(n11954));
  jor  g11763(.dina(n11954), .dinb(n11743), .dout(n11955));
  jor  g11764(.dina(n11689), .dinb(n11516), .dout(n11956));
  jand g11765(.dina(n11956), .dinb(n11693), .dout(n11957));
  jxor g11766(.dina(n11957), .dinb(n11955), .dout(n11958));
  jxor g11767(.dina(n11958), .dinb(n11736), .dout(n11959));
  jnot g11768(.din(n11959), .dout(n11960));
  jor  g11769(.dina(n11750), .dinb(n11740), .dout(n11961));
  jand g11770(.dina(n11751), .dinb(n11723), .dout(n11962));
  jnot g11771(.din(n11962), .dout(n11963));
  jand g11772(.dina(n11963), .dinb(n11961), .dout(n11964));
  jxor g11773(.dina(n11964), .dinb(n11960), .dout(n11965));
  jxor g11774(.dina(n11965), .dinb(n11953), .dout(n11966));
  jxor g11775(.dina(n11966), .dinb(n11945), .dout(n11967));
  jand g11776(.dina(n11780), .dinb(n11777), .dout(n11968));
  jnot g11777(.din(n11968), .dout(n11969));
  jor  g11778(.dina(n11792), .dinb(n11782), .dout(n11970));
  jand g11779(.dina(n11970), .dinb(n11969), .dout(n11971));
  jnot g11780(.din(n11971), .dout(n11972));
  jand g11781(.dina(n11695), .dinb(n11687), .dout(n11973));
  jand g11782(.dina(n11704), .dinb(n11696), .dout(n11974));
  jor  g11783(.dina(n11974), .dinb(n11973), .dout(n11975));
  jxor g11784(.dina(n11975), .dinb(n11972), .dout(n11976));
  jand g11785(.dina(\a[63] ), .dinb(\a[19] ), .dout(n11977));
  jor  g11786(.dina(n11684), .dinb(\a[40] ), .dout(n11978));
  jand g11787(.dina(n11978), .dinb(\a[41] ), .dout(n11979));
  jxor g11788(.dina(n11979), .dinb(n11977), .dout(n11980));
  jand g11789(.dina(n11830), .dinb(n11827), .dout(n11981));
  jnot g11790(.din(n11981), .dout(n11982));
  jand g11791(.dina(n11982), .dinb(n11832), .dout(n11983));
  jxor g11792(.dina(n11983), .dinb(n11980), .dout(n11984));
  jxor g11793(.dina(n11984), .dinb(n11976), .dout(n11985));
  jxor g11794(.dina(n11985), .dinb(n11967), .dout(n11986));
  jand g11795(.dina(n11753), .dinb(n11680), .dout(n11987));
  jand g11796(.dina(n11754), .dinb(n11677), .dout(n11988));
  jor  g11797(.dina(n11988), .dinb(n11987), .dout(n11989));
  jand g11798(.dina(n11803), .dinb(n11800), .dout(n11990));
  jand g11799(.dina(n11804), .dinb(n11797), .dout(n11991));
  jor  g11800(.dina(n11991), .dinb(n11990), .dout(n11992));
  jand g11801(.dina(n11765), .dinb(n11762), .dout(n11993));
  jand g11802(.dina(n11768), .dinb(n11766), .dout(n11994));
  jor  g11803(.dina(n11994), .dinb(n11993), .dout(n11995));
  jand g11804(.dina(\a[54] ), .dinb(\a[28] ), .dout(n11996));
  jand g11805(.dina(\a[57] ), .dinb(\a[55] ), .dout(n11997));
  jand g11806(.dina(n11997), .dinb(n2259), .dout(n11998));
  jnot g11807(.din(n11998), .dout(n11999));
  jand g11808(.dina(\a[55] ), .dinb(\a[28] ), .dout(n12000));
  jand g11809(.dina(n12000), .dinb(n11826), .dout(n12001));
  jand g11810(.dina(\a[57] ), .dinb(\a[25] ), .dout(n12002));
  jand g11811(.dina(n12002), .dinb(n11996), .dout(n12003));
  jor  g11812(.dina(n12003), .dinb(n12001), .dout(n12004));
  jand g11813(.dina(n12004), .dinb(n11999), .dout(n12005));
  jnot g11814(.din(n12005), .dout(n12006));
  jand g11815(.dina(n12006), .dinb(n11996), .dout(n12007));
  jand g11816(.dina(\a[55] ), .dinb(\a[27] ), .dout(n12008));
  jor  g11817(.dina(n12008), .dinb(n12002), .dout(n12009));
  jor  g11818(.dina(n12004), .dinb(n11998), .dout(n12010));
  jnot g11819(.din(n12010), .dout(n12011));
  jand g11820(.dina(n12011), .dinb(n12009), .dout(n12012));
  jor  g11821(.dina(n12012), .dinb(n12007), .dout(n12013));
  jxor g11822(.dina(n12013), .dinb(n11995), .dout(n12014));
  jxor g11823(.dina(n12014), .dinb(n11992), .dout(n12015));
  jor  g11824(.dina(n11774), .dinb(n11770), .dout(n12016));
  jand g11825(.dina(n11793), .dinb(n11775), .dout(n12017));
  jnot g11826(.din(n12017), .dout(n12018));
  jand g11827(.dina(n12018), .dinb(n12016), .dout(n12019));
  jor  g11828(.dina(n11812), .dinb(n11808), .dout(n12020));
  jand g11829(.dina(n11813), .dinb(n11805), .dout(n12021));
  jnot g11830(.din(n12021), .dout(n12022));
  jand g11831(.dina(n12022), .dinb(n12020), .dout(n12023));
  jxor g11832(.dina(n12023), .dinb(n12019), .dout(n12024));
  jxor g11833(.dina(n12024), .dinb(n12015), .dout(n12025));
  jxor g11834(.dina(n12025), .dinb(n11989), .dout(n12026));
  jxor g11835(.dina(n12026), .dinb(n11986), .dout(n12027));
  jxor g11836(.dina(n12027), .dinb(n11942), .dout(n12028));
  jand g11837(.dina(n12028), .dinb(n11863), .dout(n12029));
  jor  g11838(.dina(n12028), .dinb(n11863), .dout(n12030));
  jnot g11839(.din(n12030), .dout(n12031));
  jor  g11840(.dina(n12031), .dinb(n12029), .dout(n12032));
  jnot g11841(.din(n11850), .dout(n12033));
  jor  g11842(.dina(n11859), .dinb(n11852), .dout(n12034));
  jand g11843(.dina(n12034), .dinb(n12033), .dout(n12035));
  jxor g11844(.dina(n12035), .dinb(n12032), .dout(\asquared[83] ));
  jand g11845(.dina(n11941), .dinb(n11866), .dout(n12037));
  jand g11846(.dina(n12027), .dinb(n11942), .dout(n12038));
  jor  g11847(.dina(n12038), .dinb(n12037), .dout(n12039));
  jand g11848(.dina(n12025), .dinb(n11989), .dout(n12040));
  jand g11849(.dina(n12026), .dinb(n11986), .dout(n12041));
  jor  g11850(.dina(n12041), .dinb(n12040), .dout(n12042));
  jand g11851(.dina(n11966), .dinb(n11945), .dout(n12043));
  jand g11852(.dina(n11985), .dinb(n11967), .dout(n12044));
  jor  g11853(.dina(n12044), .dinb(n12043), .dout(n12045));
  jor  g11854(.dina(n12023), .dinb(n12019), .dout(n12046));
  jand g11855(.dina(n12024), .dinb(n12015), .dout(n12047));
  jnot g11856(.din(n12047), .dout(n12048));
  jand g11857(.dina(n12048), .dinb(n12046), .dout(n12049));
  jnot g11858(.din(n12049), .dout(n12050));
  jand g11859(.dina(n12013), .dinb(n11995), .dout(n12051));
  jand g11860(.dina(n12014), .dinb(n11992), .dout(n12052));
  jor  g11861(.dina(n12052), .dinb(n12051), .dout(n12053));
  jand g11862(.dina(\a[62] ), .dinb(\a[21] ), .dout(n12054));
  jnot g11863(.din(\a[41] ), .dout(n12055));
  jand g11864(.dina(\a[42] ), .dinb(n12055), .dout(n12056));
  jxor g11865(.dina(n12056), .dinb(n12054), .dout(n12057));
  jnot g11866(.din(n12057), .dout(n12058));
  jand g11867(.dina(\a[54] ), .dinb(\a[29] ), .dout(n12059));
  jnot g11868(.din(n12059), .dout(n12060));
  jand g11869(.dina(n4495), .dinb(n3665), .dout(n12061));
  jnot g11870(.din(n12061), .dout(n12062));
  jand g11871(.dina(\a[43] ), .dinb(\a[40] ), .dout(n12063));
  jor  g11872(.dina(n12063), .dinb(n11924), .dout(n12064));
  jand g11873(.dina(n12064), .dinb(n12062), .dout(n12065));
  jxor g11874(.dina(n12065), .dinb(n12060), .dout(n12066));
  jxor g11875(.dina(n12066), .dinb(n12058), .dout(n12067));
  jnot g11876(.din(n12067), .dout(n12068));
  jand g11877(.dina(\a[50] ), .dinb(\a[33] ), .dout(n12069));
  jnot g11878(.din(n12069), .dout(n12070));
  jand g11879(.dina(n7729), .dinb(n2845), .dout(n12071));
  jnot g11880(.din(n12071), .dout(n12072));
  jand g11881(.dina(\a[48] ), .dinb(\a[35] ), .dout(n12073));
  jand g11882(.dina(\a[49] ), .dinb(\a[34] ), .dout(n12074));
  jor  g11883(.dina(n12074), .dinb(n12073), .dout(n12075));
  jand g11884(.dina(n12075), .dinb(n12072), .dout(n12076));
  jxor g11885(.dina(n12076), .dinb(n12070), .dout(n12077));
  jxor g11886(.dina(n12077), .dinb(n12068), .dout(n12078));
  jxor g11887(.dina(n12078), .dinb(n12053), .dout(n12079));
  jand g11888(.dina(\a[57] ), .dinb(\a[26] ), .dout(n12080));
  jand g11889(.dina(\a[51] ), .dinb(\a[32] ), .dout(n12081));
  jor  g11890(.dina(n12081), .dinb(n12080), .dout(n12082));
  jand g11891(.dina(\a[57] ), .dinb(\a[51] ), .dout(n12083));
  jand g11892(.dina(n12083), .dinb(n6805), .dout(n12084));
  jnot g11893(.din(n12084), .dout(n12085));
  jand g11894(.dina(n7519), .dinb(n2128), .dout(n12086));
  jand g11895(.dina(\a[58] ), .dinb(\a[25] ), .dout(n12087));
  jand g11896(.dina(n12087), .dinb(n12081), .dout(n12088));
  jor  g11897(.dina(n12088), .dinb(n12086), .dout(n12089));
  jnot g11898(.din(n12089), .dout(n12090));
  jand g11899(.dina(n12090), .dinb(n12085), .dout(n12091));
  jand g11900(.dina(n12091), .dinb(n12082), .dout(n12092));
  jand g11901(.dina(n12089), .dinb(n12085), .dout(n12093));
  jnot g11902(.din(n12093), .dout(n12094));
  jand g11903(.dina(n12094), .dinb(n12087), .dout(n12095));
  jor  g11904(.dina(n12095), .dinb(n12092), .dout(n12096));
  jnot g11905(.din(n11910), .dout(n12097));
  jand g11906(.dina(\a[46] ), .dinb(\a[38] ), .dout(n12098));
  jand g11907(.dina(n12098), .dinb(n5196), .dout(n12099));
  jnot g11908(.din(n12099), .dout(n12100));
  jand g11909(.dina(\a[45] ), .dinb(\a[38] ), .dout(n12101));
  jor  g11910(.dina(n12101), .dinb(n11906), .dout(n12102));
  jand g11911(.dina(n12102), .dinb(n12100), .dout(n12103));
  jxor g11912(.dina(n12103), .dinb(n12097), .dout(n12104));
  jnot g11913(.din(n12104), .dout(n12105));
  jxor g11914(.dina(n12105), .dinb(n12096), .dout(n12106));
  jnot g11915(.din(n12106), .dout(n12107));
  jand g11916(.dina(\a[56] ), .dinb(\a[27] ), .dout(n12108));
  jnot g11917(.din(n12108), .dout(n12109));
  jand g11918(.dina(n8387), .dinb(n3581), .dout(n12110));
  jnot g11919(.din(n12110), .dout(n12111));
  jand g11920(.dina(\a[63] ), .dinb(\a[20] ), .dout(n12112));
  jand g11921(.dina(\a[61] ), .dinb(\a[22] ), .dout(n12113));
  jor  g11922(.dina(n12113), .dinb(n12112), .dout(n12114));
  jand g11923(.dina(n12114), .dinb(n12111), .dout(n12115));
  jxor g11924(.dina(n12115), .dinb(n12109), .dout(n12116));
  jxor g11925(.dina(n12116), .dinb(n12107), .dout(n12117));
  jxor g11926(.dina(n12117), .dinb(n12079), .dout(n12118));
  jxor g11927(.dina(n12118), .dinb(n12050), .dout(n12119));
  jxor g11928(.dina(n12119), .dinb(n12045), .dout(n12120));
  jxor g11929(.dina(n12120), .dinb(n12042), .dout(n12121));
  jand g11930(.dina(n11939), .dinb(n11874), .dout(n12122));
  jand g11931(.dina(n11940), .dinb(n11869), .dout(n12123));
  jor  g11932(.dina(n12123), .dinb(n12122), .dout(n12124));
  jand g11933(.dina(n11951), .dinb(n11948), .dout(n12125));
  jand g11934(.dina(n11952), .dinb(n11946), .dout(n12126));
  jor  g11935(.dina(n12126), .dinb(n12125), .dout(n12127));
  jand g11936(.dina(n11957), .dinb(n11955), .dout(n12128));
  jand g11937(.dina(n11958), .dinb(n11736), .dout(n12129));
  jor  g11938(.dina(n12129), .dinb(n12128), .dout(n12130));
  jxor g11939(.dina(n12130), .dinb(n12127), .dout(n12131));
  jnot g11940(.din(n12131), .dout(n12132));
  jand g11941(.dina(n11890), .dinb(n11883), .dout(n12133));
  jnot g11942(.din(n12133), .dout(n12134));
  jor  g11943(.dina(n11902), .dinb(n11892), .dout(n12135));
  jand g11944(.dina(n12135), .dinb(n12134), .dout(n12136));
  jxor g11945(.dina(n12136), .dinb(n12132), .dout(n12137));
  jand g11946(.dina(n11979), .dinb(n11977), .dout(n12138));
  jand g11947(.dina(n11983), .dinb(n11980), .dout(n12139));
  jor  g11948(.dina(n12139), .dinb(n12138), .dout(n12140));
  jand g11949(.dina(\a[52] ), .dinb(\a[31] ), .dout(n12141));
  jand g11950(.dina(n6498), .dinb(n2810), .dout(n12142));
  jnot g11951(.din(n12142), .dout(n12143));
  jand g11952(.dina(n7165), .dinb(n2440), .dout(n12144));
  jand g11953(.dina(n12141), .dinb(n12000), .dout(n12145));
  jor  g11954(.dina(n12145), .dinb(n12144), .dout(n12146));
  jand g11955(.dina(n12146), .dinb(n12143), .dout(n12147));
  jnot g11956(.din(n12147), .dout(n12148));
  jand g11957(.dina(n12148), .dinb(n12141), .dout(n12149));
  jand g11958(.dina(\a[53] ), .dinb(\a[30] ), .dout(n12150));
  jor  g11959(.dina(n12150), .dinb(n12000), .dout(n12151));
  jor  g11960(.dina(n12146), .dinb(n12142), .dout(n12152));
  jnot g11961(.din(n12152), .dout(n12153));
  jand g11962(.dina(n12153), .dinb(n12151), .dout(n12154));
  jor  g11963(.dina(n12154), .dinb(n12149), .dout(n12155));
  jand g11964(.dina(\a[60] ), .dinb(\a[24] ), .dout(n12156));
  jand g11965(.dina(n12156), .dinb(n11899), .dout(n12157));
  jnot g11966(.din(n12157), .dout(n12158));
  jand g11967(.dina(\a[60] ), .dinb(\a[23] ), .dout(n12159));
  jor  g11968(.dina(n12159), .dinb(n11895), .dout(n12160));
  jand g11969(.dina(n12160), .dinb(n12158), .dout(n12161));
  jor  g11970(.dina(n11930), .dinb(n11929), .dout(n12162));
  jand g11971(.dina(n12162), .dinb(n11934), .dout(n12163));
  jxor g11972(.dina(n12163), .dinb(n12161), .dout(n12164));
  jxor g11973(.dina(n12164), .dinb(n12155), .dout(n12165));
  jxor g11974(.dina(n12165), .dinb(n12140), .dout(n12166));
  jand g11975(.dina(n11975), .dinb(n11972), .dout(n12167));
  jand g11976(.dina(n11984), .dinb(n11976), .dout(n12168));
  jor  g11977(.dina(n12168), .dinb(n12167), .dout(n12169));
  jxor g11978(.dina(n12169), .dinb(n12166), .dout(n12170));
  jxor g11979(.dina(n12170), .dinb(n12137), .dout(n12171));
  jxor g11980(.dina(n12171), .dinb(n12124), .dout(n12172));
  jand g11981(.dina(n11927), .dinb(n11921), .dout(n12173));
  jor  g11982(.dina(n12173), .dinb(n11925), .dout(n12174));
  jand g11983(.dina(n11897), .dinb(n11894), .dout(n12175));
  jnot g11984(.din(n12175), .dout(n12176));
  jand g11985(.dina(n12176), .dinb(n11900), .dout(n12177));
  jxor g11986(.dina(n12177), .dinb(n11916), .dout(n12178));
  jxor g11987(.dina(n12178), .dinb(n12174), .dout(n12179));
  jand g11988(.dina(n11881), .dinb(n11742), .dout(n12180));
  jand g11989(.dina(n11882), .dinb(n11880), .dout(n12181));
  jor  g11990(.dina(n12181), .dinb(n12180), .dout(n12182));
  jor  g11991(.dina(n11884), .dinb(n11785), .dout(n12183));
  jand g11992(.dina(n12183), .dinb(n11888), .dout(n12184));
  jxor g11993(.dina(n12184), .dinb(n12182), .dout(n12185));
  jxor g11994(.dina(n12185), .dinb(n12010), .dout(n12186));
  jand g11995(.dina(n11936), .dinb(n11928), .dout(n12187));
  jand g11996(.dina(n11937), .dinb(n11920), .dout(n12188));
  jor  g11997(.dina(n12188), .dinb(n12187), .dout(n12189));
  jxor g11998(.dina(n12189), .dinb(n12186), .dout(n12190));
  jxor g11999(.dina(n12190), .dinb(n12179), .dout(n12191));
  jand g12000(.dina(n11903), .dinb(n11879), .dout(n12192));
  jand g12001(.dina(n11938), .dinb(n11904), .dout(n12193));
  jor  g12002(.dina(n12193), .dinb(n12192), .dout(n12194));
  jnot g12003(.din(n12194), .dout(n12195));
  jor  g12004(.dina(n11964), .dinb(n11960), .dout(n12196));
  jand g12005(.dina(n11965), .dinb(n11953), .dout(n12197));
  jnot g12006(.din(n12197), .dout(n12198));
  jand g12007(.dina(n12198), .dinb(n12196), .dout(n12199));
  jxor g12008(.dina(n12199), .dinb(n12195), .dout(n12200));
  jxor g12009(.dina(n12200), .dinb(n12191), .dout(n12201));
  jxor g12010(.dina(n12201), .dinb(n12172), .dout(n12202));
  jxor g12011(.dina(n12202), .dinb(n12121), .dout(n12203));
  jand g12012(.dina(n12203), .dinb(n12039), .dout(n12204));
  jor  g12013(.dina(n12203), .dinb(n12039), .dout(n12205));
  jnot g12014(.din(n12205), .dout(n12206));
  jor  g12015(.dina(n12206), .dinb(n12204), .dout(n12207));
  jnot g12016(.din(n12029), .dout(n12208));
  jor  g12017(.dina(n12035), .dinb(n12031), .dout(n12209));
  jand g12018(.dina(n12209), .dinb(n12208), .dout(n12210));
  jxor g12019(.dina(n12210), .dinb(n12207), .dout(\asquared[84] ));
  jand g12020(.dina(n12120), .dinb(n12042), .dout(n12212));
  jand g12021(.dina(n12202), .dinb(n12121), .dout(n12213));
  jor  g12022(.dina(n12213), .dinb(n12212), .dout(n12214));
  jand g12023(.dina(n12171), .dinb(n12124), .dout(n12215));
  jand g12024(.dina(n12201), .dinb(n12172), .dout(n12216));
  jor  g12025(.dina(n12216), .dinb(n12215), .dout(n12217));
  jand g12026(.dina(n12164), .dinb(n12155), .dout(n12218));
  jand g12027(.dina(n12165), .dinb(n12140), .dout(n12219));
  jor  g12028(.dina(n12219), .dinb(n12218), .dout(n12220));
  jand g12029(.dina(n12163), .dinb(n12161), .dout(n12221));
  jor  g12030(.dina(n12221), .dinb(n12157), .dout(n12222));
  jand g12031(.dina(n12111), .dinb(n12109), .dout(n12223));
  jnot g12032(.din(n12223), .dout(n12224));
  jand g12033(.dina(n12224), .dinb(n12114), .dout(n12225));
  jxor g12034(.dina(n12225), .dinb(n12222), .dout(n12226));
  jand g12035(.dina(\a[58] ), .dinb(\a[26] ), .dout(n12227));
  jand g12036(.dina(n7165), .dinb(n3269), .dout(n12228));
  jnot g12037(.din(n12228), .dout(n12229));
  jand g12038(.dina(\a[53] ), .dinb(\a[31] ), .dout(n12230));
  jand g12039(.dina(\a[52] ), .dinb(\a[32] ), .dout(n12231));
  jor  g12040(.dina(n12231), .dinb(n12230), .dout(n12232));
  jand g12041(.dina(n12232), .dinb(n12229), .dout(n12233));
  jxor g12042(.dina(n12233), .dinb(n12227), .dout(n12234));
  jxor g12043(.dina(n12234), .dinb(n12226), .dout(n12235));
  jxor g12044(.dina(n12235), .dinb(n12220), .dout(n12236));
  jnot g12045(.din(n12236), .dout(n12237));
  jand g12046(.dina(n12130), .dinb(n12127), .dout(n12238));
  jnot g12047(.din(n12238), .dout(n12239));
  jor  g12048(.dina(n12136), .dinb(n12132), .dout(n12240));
  jand g12049(.dina(n12240), .dinb(n12239), .dout(n12241));
  jxor g12050(.dina(n12241), .dinb(n12237), .dout(n12242));
  jand g12051(.dina(n12169), .dinb(n12166), .dout(n12243));
  jand g12052(.dina(n12170), .dinb(n12137), .dout(n12244));
  jor  g12053(.dina(n12244), .dinb(n12243), .dout(n12245));
  jxor g12054(.dina(n12245), .dinb(n12242), .dout(n12246));
  jnot g12055(.din(n12091), .dout(n12247));
  jand g12056(.dina(n12072), .dinb(n12070), .dout(n12248));
  jnot g12057(.din(n12248), .dout(n12249));
  jand g12058(.dina(n12249), .dinb(n12075), .dout(n12250));
  jand g12059(.dina(n12100), .dinb(n12097), .dout(n12251));
  jnot g12060(.din(n12251), .dout(n12252));
  jand g12061(.dina(n12252), .dinb(n12102), .dout(n12253));
  jxor g12062(.dina(n12253), .dinb(n12250), .dout(n12254));
  jxor g12063(.dina(n12254), .dinb(n12247), .dout(n12255));
  jand g12064(.dina(n12177), .dinb(n11916), .dout(n12256));
  jand g12065(.dina(n12178), .dinb(n12174), .dout(n12257));
  jor  g12066(.dina(n12257), .dinb(n12256), .dout(n12258));
  jand g12067(.dina(n12184), .dinb(n12182), .dout(n12259));
  jand g12068(.dina(n12185), .dinb(n12010), .dout(n12260));
  jor  g12069(.dina(n12260), .dinb(n12259), .dout(n12261));
  jxor g12070(.dina(n12261), .dinb(n12258), .dout(n12262));
  jxor g12071(.dina(n12262), .dinb(n12255), .dout(n12263));
  jand g12072(.dina(\a[63] ), .dinb(\a[21] ), .dout(n12264));
  jand g12073(.dina(n8702), .dinb(n1658), .dout(n12265));
  jnot g12074(.din(n12265), .dout(n12266));
  jand g12075(.dina(\a[62] ), .dinb(\a[22] ), .dout(n12267));
  jand g12076(.dina(\a[61] ), .dinb(\a[23] ), .dout(n12268));
  jor  g12077(.dina(n12268), .dinb(n12267), .dout(n12269));
  jand g12078(.dina(n12269), .dinb(n12266), .dout(n12270));
  jxor g12079(.dina(n12270), .dinb(n12264), .dout(n12271));
  jnot g12080(.din(n12271), .dout(n12272));
  jand g12081(.dina(\a[51] ), .dinb(\a[33] ), .dout(n12273));
  jnot g12082(.din(n12273), .dout(n12274));
  jand g12083(.dina(\a[60] ), .dinb(\a[25] ), .dout(n12275));
  jand g12084(.dina(n12275), .dinb(n11895), .dout(n12276));
  jnot g12085(.din(n12276), .dout(n12277));
  jand g12086(.dina(\a[59] ), .dinb(\a[25] ), .dout(n12278));
  jor  g12087(.dina(n12278), .dinb(n12156), .dout(n12279));
  jand g12088(.dina(n12279), .dinb(n12277), .dout(n12280));
  jxor g12089(.dina(n12280), .dinb(n12274), .dout(n12281));
  jxor g12090(.dina(n12281), .dinb(n12272), .dout(n12282));
  jnot g12091(.din(n12282), .dout(n12283));
  jand g12092(.dina(\a[50] ), .dinb(\a[34] ), .dout(n12284));
  jnot g12093(.din(n12284), .dout(n12285));
  jand g12094(.dina(n7729), .dinb(n3243), .dout(n12286));
  jnot g12095(.din(n12286), .dout(n12287));
  jand g12096(.dina(\a[49] ), .dinb(\a[35] ), .dout(n12288));
  jand g12097(.dina(\a[48] ), .dinb(\a[36] ), .dout(n12289));
  jor  g12098(.dina(n12289), .dinb(n12288), .dout(n12290));
  jand g12099(.dina(n12290), .dinb(n12287), .dout(n12291));
  jxor g12100(.dina(n12291), .dinb(n12285), .dout(n12292));
  jxor g12101(.dina(n12292), .dinb(n12283), .dout(n12293));
  jnot g12102(.din(n12098), .dout(n12294));
  jand g12103(.dina(\a[55] ), .dinb(\a[29] ), .dout(n12295));
  jnot g12104(.din(n12295), .dout(n12296));
  jand g12105(.dina(n12296), .dinb(n12294), .dout(n12297));
  jand g12106(.dina(n12295), .dinb(n12098), .dout(n12298));
  jnot g12107(.din(n12298), .dout(n12299));
  jand g12108(.dina(\a[56] ), .dinb(\a[29] ), .dout(n12300));
  jand g12109(.dina(n12300), .dinb(n12000), .dout(n12301));
  jand g12110(.dina(\a[56] ), .dinb(\a[28] ), .dout(n12302));
  jand g12111(.dina(n12302), .dinb(n12098), .dout(n12303));
  jor  g12112(.dina(n12303), .dinb(n12301), .dout(n12304));
  jnot g12113(.din(n12304), .dout(n12305));
  jand g12114(.dina(n12305), .dinb(n12299), .dout(n12306));
  jnot g12115(.din(n12306), .dout(n12307));
  jor  g12116(.dina(n12307), .dinb(n12297), .dout(n12308));
  jand g12117(.dina(n12304), .dinb(n12299), .dout(n12309));
  jnot g12118(.din(n12309), .dout(n12310));
  jand g12119(.dina(n12310), .dinb(n12302), .dout(n12311));
  jnot g12120(.din(n12311), .dout(n12312));
  jand g12121(.dina(n12312), .dinb(n12308), .dout(n12313));
  jand g12122(.dina(\a[45] ), .dinb(\a[39] ), .dout(n12314));
  jnot g12123(.din(n12314), .dout(n12315));
  jand g12124(.dina(n4632), .dinb(n4495), .dout(n12316));
  jnot g12125(.din(n12316), .dout(n12317));
  jand g12126(.dina(\a[44] ), .dinb(\a[40] ), .dout(n12318));
  jor  g12127(.dina(n12318), .dinb(n4115), .dout(n12319));
  jand g12128(.dina(n12319), .dinb(n12317), .dout(n12320));
  jxor g12129(.dina(n12320), .dinb(n12315), .dout(n12321));
  jxor g12130(.dina(n12321), .dinb(n12313), .dout(n12322));
  jnot g12131(.din(n12322), .dout(n12323));
  jand g12132(.dina(\a[47] ), .dinb(\a[37] ), .dout(n12324));
  jnot g12133(.din(n12324), .dout(n12325));
  jand g12134(.dina(\a[57] ), .dinb(\a[27] ), .dout(n12326));
  jand g12135(.dina(\a[54] ), .dinb(\a[30] ), .dout(n12327));
  jxor g12136(.dina(n12327), .dinb(n12326), .dout(n12328));
  jxor g12137(.dina(n12328), .dinb(n12325), .dout(n12329));
  jxor g12138(.dina(n12329), .dinb(n12323), .dout(n12330));
  jxor g12139(.dina(n12330), .dinb(n12293), .dout(n12331));
  jxor g12140(.dina(n12331), .dinb(n12263), .dout(n12332));
  jxor g12141(.dina(n12332), .dinb(n12246), .dout(n12333));
  jxor g12142(.dina(n12333), .dinb(n12217), .dout(n12334));
  jand g12143(.dina(n12118), .dinb(n12050), .dout(n12335));
  jand g12144(.dina(n12119), .dinb(n12045), .dout(n12336));
  jor  g12145(.dina(n12336), .dinb(n12335), .dout(n12337));
  jnot g12146(.din(n12337), .dout(n12338));
  jor  g12147(.dina(n12199), .dinb(n12195), .dout(n12339));
  jand g12148(.dina(n12200), .dinb(n12191), .dout(n12340));
  jnot g12149(.din(n12340), .dout(n12341));
  jand g12150(.dina(n12341), .dinb(n12339), .dout(n12342));
  jxor g12151(.dina(n12342), .dinb(n12338), .dout(n12343));
  jand g12152(.dina(n12062), .dinb(n12060), .dout(n12344));
  jnot g12153(.din(n12344), .dout(n12345));
  jand g12154(.dina(n12345), .dinb(n12064), .dout(n12346));
  jor  g12155(.dina(n12054), .dinb(\a[41] ), .dout(n12347));
  jand g12156(.dina(n12347), .dinb(\a[42] ), .dout(n12348));
  jxor g12157(.dina(n12348), .dinb(n12346), .dout(n12349));
  jxor g12158(.dina(n12349), .dinb(n12152), .dout(n12350));
  jand g12159(.dina(n12105), .dinb(n12096), .dout(n12351));
  jnot g12160(.din(n12351), .dout(n12352));
  jor  g12161(.dina(n12116), .dinb(n12107), .dout(n12353));
  jand g12162(.dina(n12353), .dinb(n12352), .dout(n12354));
  jor  g12163(.dina(n12066), .dinb(n12058), .dout(n12355));
  jor  g12164(.dina(n12077), .dinb(n12068), .dout(n12356));
  jand g12165(.dina(n12356), .dinb(n12355), .dout(n12357));
  jxor g12166(.dina(n12357), .dinb(n12354), .dout(n12358));
  jxor g12167(.dina(n12358), .dinb(n12350), .dout(n12359));
  jand g12168(.dina(n12078), .dinb(n12053), .dout(n12360));
  jand g12169(.dina(n12117), .dinb(n12079), .dout(n12361));
  jor  g12170(.dina(n12361), .dinb(n12360), .dout(n12362));
  jand g12171(.dina(n12189), .dinb(n12186), .dout(n12363));
  jand g12172(.dina(n12190), .dinb(n12179), .dout(n12364));
  jor  g12173(.dina(n12364), .dinb(n12363), .dout(n12365));
  jxor g12174(.dina(n12365), .dinb(n12362), .dout(n12366));
  jxor g12175(.dina(n12366), .dinb(n12359), .dout(n12367));
  jxor g12176(.dina(n12367), .dinb(n12343), .dout(n12368));
  jxor g12177(.dina(n12368), .dinb(n12334), .dout(n12369));
  jand g12178(.dina(n12369), .dinb(n12214), .dout(n12370));
  jor  g12179(.dina(n12369), .dinb(n12214), .dout(n12371));
  jnot g12180(.din(n12371), .dout(n12372));
  jor  g12181(.dina(n12372), .dinb(n12370), .dout(n12373));
  jnot g12182(.din(n12204), .dout(n12374));
  jor  g12183(.dina(n12210), .dinb(n12206), .dout(n12375));
  jand g12184(.dina(n12375), .dinb(n12374), .dout(n12376));
  jxor g12185(.dina(n12376), .dinb(n12373), .dout(\asquared[85] ));
  jand g12186(.dina(n12333), .dinb(n12217), .dout(n12378));
  jand g12187(.dina(n12368), .dinb(n12334), .dout(n12379));
  jor  g12188(.dina(n12379), .dinb(n12378), .dout(n12380));
  jand g12189(.dina(n12365), .dinb(n12362), .dout(n12381));
  jand g12190(.dina(n12366), .dinb(n12359), .dout(n12382));
  jor  g12191(.dina(n12382), .dinb(n12381), .dout(n12383));
  jand g12192(.dina(n12253), .dinb(n12250), .dout(n12384));
  jand g12193(.dina(n12254), .dinb(n12247), .dout(n12385));
  jor  g12194(.dina(n12385), .dinb(n12384), .dout(n12386));
  jand g12195(.dina(n12348), .dinb(n12346), .dout(n12387));
  jand g12196(.dina(n12349), .dinb(n12152), .dout(n12388));
  jor  g12197(.dina(n12388), .dinb(n12387), .dout(n12389));
  jxor g12198(.dina(n12389), .dinb(n12386), .dout(n12390));
  jand g12199(.dina(n12225), .dinb(n12222), .dout(n12391));
  jand g12200(.dina(n12234), .dinb(n12226), .dout(n12392));
  jor  g12201(.dina(n12392), .dinb(n12391), .dout(n12393));
  jxor g12202(.dina(n12393), .dinb(n12390), .dout(n12394));
  jnot g12203(.din(n12394), .dout(n12395));
  jand g12204(.dina(n12235), .dinb(n12220), .dout(n12396));
  jnot g12205(.din(n12396), .dout(n12397));
  jor  g12206(.dina(n12241), .dinb(n12237), .dout(n12398));
  jand g12207(.dina(n12398), .dinb(n12397), .dout(n12399));
  jxor g12208(.dina(n12399), .dinb(n12395), .dout(n12400));
  jand g12209(.dina(n12330), .dinb(n12293), .dout(n12401));
  jand g12210(.dina(n12331), .dinb(n12263), .dout(n12402));
  jor  g12211(.dina(n12402), .dinb(n12401), .dout(n12403));
  jxor g12212(.dina(n12403), .dinb(n12400), .dout(n12404));
  jxor g12213(.dina(n12404), .dinb(n12383), .dout(n12405));
  jand g12214(.dina(n12245), .dinb(n12242), .dout(n12406));
  jand g12215(.dina(n12332), .dinb(n12246), .dout(n12407));
  jor  g12216(.dina(n12407), .dinb(n12406), .dout(n12408));
  jxor g12217(.dina(n12408), .dinb(n12405), .dout(n12409));
  jor  g12218(.dina(n12342), .dinb(n12338), .dout(n12410));
  jand g12219(.dina(n12367), .dinb(n12343), .dout(n12411));
  jnot g12220(.din(n12411), .dout(n12412));
  jand g12221(.dina(n12412), .dinb(n12410), .dout(n12413));
  jnot g12222(.din(n12413), .dout(n12414));
  jor  g12223(.dina(n12357), .dinb(n12354), .dout(n12415));
  jand g12224(.dina(n12358), .dinb(n12350), .dout(n12416));
  jnot g12225(.din(n12416), .dout(n12417));
  jand g12226(.dina(n12417), .dinb(n12415), .dout(n12418));
  jnot g12227(.din(n12418), .dout(n12419));
  jand g12228(.dina(\a[50] ), .dinb(\a[35] ), .dout(n12420));
  jand g12229(.dina(\a[63] ), .dinb(\a[22] ), .dout(n12421));
  jand g12230(.dina(\a[57] ), .dinb(\a[28] ), .dout(n12422));
  jxor g12231(.dina(n12422), .dinb(n12421), .dout(n12423));
  jxor g12232(.dina(n12423), .dinb(n12420), .dout(n12424));
  jnot g12233(.din(n12424), .dout(n12425));
  jand g12234(.dina(\a[53] ), .dinb(\a[32] ), .dout(n12426));
  jnot g12235(.din(n12426), .dout(n12427));
  jand g12236(.dina(\a[52] ), .dinb(\a[34] ), .dout(n12428));
  jand g12237(.dina(n12428), .dinb(n12273), .dout(n12429));
  jnot g12238(.din(n12429), .dout(n12430));
  jand g12239(.dina(\a[52] ), .dinb(\a[33] ), .dout(n12431));
  jand g12240(.dina(\a[51] ), .dinb(\a[34] ), .dout(n12432));
  jor  g12241(.dina(n12432), .dinb(n12431), .dout(n12433));
  jand g12242(.dina(n12433), .dinb(n12430), .dout(n12434));
  jxor g12243(.dina(n12434), .dinb(n12427), .dout(n12435));
  jxor g12244(.dina(n12435), .dinb(n12425), .dout(n12436));
  jnot g12245(.din(n12436), .dout(n12437));
  jand g12246(.dina(\a[46] ), .dinb(\a[39] ), .dout(n12438));
  jnot g12247(.din(n12438), .dout(n12439));
  jand g12248(.dina(n4812), .dinb(n4632), .dout(n12440));
  jnot g12249(.din(n12440), .dout(n12441));
  jand g12250(.dina(\a[45] ), .dinb(\a[40] ), .dout(n12442));
  jand g12251(.dina(\a[44] ), .dinb(\a[41] ), .dout(n12443));
  jor  g12252(.dina(n12443), .dinb(n12442), .dout(n12444));
  jand g12253(.dina(n12444), .dinb(n12441), .dout(n12445));
  jxor g12254(.dina(n12445), .dinb(n12439), .dout(n12446));
  jxor g12255(.dina(n12446), .dinb(n12437), .dout(n12447));
  jand g12256(.dina(\a[62] ), .dinb(\a[23] ), .dout(n12448));
  jand g12257(.dina(\a[43] ), .dinb(n4019), .dout(n12449));
  jxor g12258(.dina(n12449), .dinb(n12448), .dout(n12450));
  jnot g12259(.din(n12450), .dout(n12451));
  jand g12260(.dina(\a[49] ), .dinb(\a[36] ), .dout(n12452));
  jnot g12261(.din(n12452), .dout(n12453));
  jand g12262(.dina(n12324), .dinb(n5893), .dout(n12454));
  jnot g12263(.din(n12454), .dout(n12455));
  jand g12264(.dina(\a[47] ), .dinb(\a[38] ), .dout(n12456));
  jand g12265(.dina(\a[48] ), .dinb(\a[37] ), .dout(n12457));
  jor  g12266(.dina(n12457), .dinb(n12456), .dout(n12458));
  jand g12267(.dina(n12458), .dinb(n12455), .dout(n12459));
  jxor g12268(.dina(n12459), .dinb(n12453), .dout(n12460));
  jxor g12269(.dina(n12460), .dinb(n12451), .dout(n12461));
  jnot g12270(.din(n12461), .dout(n12462));
  jnot g12271(.din(n12300), .dout(n12463));
  jand g12272(.dina(\a[55] ), .dinb(\a[31] ), .dout(n12464));
  jand g12273(.dina(n12464), .dinb(n12327), .dout(n12465));
  jnot g12274(.din(n12465), .dout(n12466));
  jand g12275(.dina(\a[55] ), .dinb(\a[30] ), .dout(n12467));
  jand g12276(.dina(\a[54] ), .dinb(\a[31] ), .dout(n12468));
  jor  g12277(.dina(n12468), .dinb(n12467), .dout(n12469));
  jand g12278(.dina(n12469), .dinb(n12466), .dout(n12470));
  jxor g12279(.dina(n12470), .dinb(n12463), .dout(n12471));
  jxor g12280(.dina(n12471), .dinb(n12462), .dout(n12472));
  jxor g12281(.dina(n12472), .dinb(n12447), .dout(n12473));
  jxor g12282(.dina(n12473), .dinb(n12419), .dout(n12474));
  jand g12283(.dina(n12270), .dinb(n12264), .dout(n12475));
  jor  g12284(.dina(n12475), .dinb(n12265), .dout(n12476));
  jand g12285(.dina(n12287), .dinb(n12285), .dout(n12477));
  jnot g12286(.din(n12477), .dout(n12478));
  jand g12287(.dina(n12478), .dinb(n12290), .dout(n12479));
  jxor g12288(.dina(n12479), .dinb(n12476), .dout(n12480));
  jand g12289(.dina(n12277), .dinb(n12274), .dout(n12481));
  jnot g12290(.din(n12481), .dout(n12482));
  jand g12291(.dina(n12482), .dinb(n12279), .dout(n12483));
  jxor g12292(.dina(n12483), .dinb(n12480), .dout(n12484));
  jor  g12293(.dina(n12321), .dinb(n12313), .dout(n12485));
  jor  g12294(.dina(n12329), .dinb(n12323), .dout(n12486));
  jand g12295(.dina(n12486), .dinb(n12485), .dout(n12487));
  jor  g12296(.dina(n12281), .dinb(n12272), .dout(n12488));
  jor  g12297(.dina(n12292), .dinb(n12283), .dout(n12489));
  jand g12298(.dina(n12489), .dinb(n12488), .dout(n12490));
  jxor g12299(.dina(n12490), .dinb(n12487), .dout(n12491));
  jxor g12300(.dina(n12491), .dinb(n12484), .dout(n12492));
  jand g12301(.dina(n12261), .dinb(n12258), .dout(n12493));
  jand g12302(.dina(n12262), .dinb(n12255), .dout(n12494));
  jor  g12303(.dina(n12494), .dinb(n12493), .dout(n12495));
  jand g12304(.dina(\a[61] ), .dinb(\a[24] ), .dout(n12496));
  jand g12305(.dina(n12317), .dinb(n12315), .dout(n12497));
  jnot g12306(.din(n12497), .dout(n12498));
  jand g12307(.dina(n12498), .dinb(n12319), .dout(n12499));
  jxor g12308(.dina(n12499), .dinb(n12496), .dout(n12500));
  jxor g12309(.dina(n12500), .dinb(n12307), .dout(n12501));
  jand g12310(.dina(n12232), .dinb(n12227), .dout(n12502));
  jor  g12311(.dina(n12502), .dinb(n12228), .dout(n12503));
  jor  g12312(.dina(n12327), .dinb(n12326), .dout(n12504));
  jand g12313(.dina(n12327), .dinb(n12326), .dout(n12505));
  jor  g12314(.dina(n12505), .dinb(n12324), .dout(n12506));
  jand g12315(.dina(n12506), .dinb(n12504), .dout(n12507));
  jxor g12316(.dina(n12507), .dinb(n12503), .dout(n12508));
  jand g12317(.dina(\a[59] ), .dinb(\a[27] ), .dout(n12509));
  jand g12318(.dina(n12509), .dinb(n12227), .dout(n12510));
  jnot g12319(.din(n12510), .dout(n12511));
  jand g12320(.dina(\a[59] ), .dinb(\a[26] ), .dout(n12512));
  jand g12321(.dina(\a[58] ), .dinb(\a[27] ), .dout(n12513));
  jor  g12322(.dina(n12513), .dinb(n12512), .dout(n12514));
  jand g12323(.dina(n12514), .dinb(n12511), .dout(n12515));
  jxor g12324(.dina(n12515), .dinb(n12275), .dout(n12516));
  jxor g12325(.dina(n12516), .dinb(n12508), .dout(n12517));
  jxor g12326(.dina(n12517), .dinb(n12501), .dout(n12518));
  jxor g12327(.dina(n12518), .dinb(n12495), .dout(n12519));
  jxor g12328(.dina(n12519), .dinb(n12492), .dout(n12520));
  jxor g12329(.dina(n12520), .dinb(n12474), .dout(n12521));
  jxor g12330(.dina(n12521), .dinb(n12414), .dout(n12522));
  jxor g12331(.dina(n12522), .dinb(n12409), .dout(n12523));
  jand g12332(.dina(n12523), .dinb(n12380), .dout(n12524));
  jor  g12333(.dina(n12523), .dinb(n12380), .dout(n12525));
  jnot g12334(.din(n12525), .dout(n12526));
  jor  g12335(.dina(n12526), .dinb(n12524), .dout(n12527));
  jnot g12336(.din(n12370), .dout(n12528));
  jor  g12337(.dina(n12376), .dinb(n12372), .dout(n12529));
  jand g12338(.dina(n12529), .dinb(n12528), .dout(n12530));
  jxor g12339(.dina(n12530), .dinb(n12527), .dout(\asquared[86] ));
  jand g12340(.dina(n12521), .dinb(n12414), .dout(n12532));
  jand g12341(.dina(n12522), .dinb(n12409), .dout(n12533));
  jor  g12342(.dina(n12533), .dinb(n12532), .dout(n12534));
  jand g12343(.dina(n12519), .dinb(n12492), .dout(n12535));
  jand g12344(.dina(n12520), .dinb(n12474), .dout(n12536));
  jor  g12345(.dina(n12536), .dinb(n12535), .dout(n12537));
  jnot g12346(.din(n12537), .dout(n12538));
  jor  g12347(.dina(n12399), .dinb(n12395), .dout(n12539));
  jand g12348(.dina(n12403), .dinb(n12400), .dout(n12540));
  jnot g12349(.din(n12540), .dout(n12541));
  jand g12350(.dina(n12541), .dinb(n12539), .dout(n12542));
  jxor g12351(.dina(n12542), .dinb(n12538), .dout(n12543));
  jand g12352(.dina(n12517), .dinb(n12501), .dout(n12544));
  jand g12353(.dina(n12518), .dinb(n12495), .dout(n12545));
  jor  g12354(.dina(n12545), .dinb(n12544), .dout(n12546));
  jand g12355(.dina(n12499), .dinb(n12496), .dout(n12547));
  jand g12356(.dina(n12500), .dinb(n12307), .dout(n12548));
  jor  g12357(.dina(n12548), .dinb(n12547), .dout(n12549));
  jand g12358(.dina(n8702), .dinb(n1648), .dout(n12550));
  jnot g12359(.din(n12550), .dout(n12551));
  jand g12360(.dina(\a[62] ), .dinb(\a[24] ), .dout(n12552));
  jand g12361(.dina(\a[61] ), .dinb(\a[25] ), .dout(n12553));
  jor  g12362(.dina(n12553), .dinb(n12552), .dout(n12554));
  jand g12363(.dina(n12554), .dinb(n12551), .dout(n12555));
  jor  g12364(.dina(n12448), .dinb(\a[42] ), .dout(n12556));
  jand g12365(.dina(n12556), .dinb(\a[43] ), .dout(n12557));
  jxor g12366(.dina(n12557), .dinb(n12555), .dout(n12558));
  jxor g12367(.dina(n12558), .dinb(n12549), .dout(n12559));
  jand g12368(.dina(n12479), .dinb(n12476), .dout(n12560));
  jand g12369(.dina(n12483), .dinb(n12480), .dout(n12561));
  jor  g12370(.dina(n12561), .dinb(n12560), .dout(n12562));
  jxor g12371(.dina(n12562), .dinb(n12559), .dout(n12563));
  jxor g12372(.dina(n12563), .dinb(n12546), .dout(n12564));
  jand g12373(.dina(n12472), .dinb(n12447), .dout(n12565));
  jand g12374(.dina(n12473), .dinb(n12419), .dout(n12566));
  jor  g12375(.dina(n12566), .dinb(n12565), .dout(n12567));
  jxor g12376(.dina(n12567), .dinb(n12564), .dout(n12568));
  jxor g12377(.dina(n12568), .dinb(n12543), .dout(n12569));
  jand g12378(.dina(n12404), .dinb(n12383), .dout(n12570));
  jand g12379(.dina(n12408), .dinb(n12405), .dout(n12571));
  jor  g12380(.dina(n12571), .dinb(n12570), .dout(n12572));
  jand g12381(.dina(n12507), .dinb(n12503), .dout(n12573));
  jand g12382(.dina(n12516), .dinb(n12508), .dout(n12574));
  jor  g12383(.dina(n12574), .dinb(n12573), .dout(n12575));
  jnot g12384(.din(n12575), .dout(n12576));
  jor  g12385(.dina(n12435), .dinb(n12425), .dout(n12577));
  jor  g12386(.dina(n12446), .dinb(n12437), .dout(n12578));
  jand g12387(.dina(n12578), .dinb(n12577), .dout(n12579));
  jxor g12388(.dina(n12579), .dinb(n12576), .dout(n12580));
  jnot g12389(.din(n12580), .dout(n12581));
  jor  g12390(.dina(n12460), .dinb(n12451), .dout(n12582));
  jor  g12391(.dina(n12471), .dinb(n12462), .dout(n12583));
  jand g12392(.dina(n12583), .dinb(n12582), .dout(n12584));
  jxor g12393(.dina(n12584), .dinb(n12581), .dout(n12585));
  jand g12394(.dina(n12389), .dinb(n12386), .dout(n12586));
  jand g12395(.dina(n12393), .dinb(n12390), .dout(n12587));
  jor  g12396(.dina(n12587), .dinb(n12586), .dout(n12588));
  jand g12397(.dina(n12441), .dinb(n12439), .dout(n12589));
  jnot g12398(.din(n12589), .dout(n12590));
  jand g12399(.dina(n12590), .dinb(n12444), .dout(n12591));
  jand g12400(.dina(n12466), .dinb(n12463), .dout(n12592));
  jnot g12401(.din(n12592), .dout(n12593));
  jand g12402(.dina(n12593), .dinb(n12469), .dout(n12594));
  jxor g12403(.dina(n12594), .dinb(n12591), .dout(n12595));
  jand g12404(.dina(n12455), .dinb(n12453), .dout(n12596));
  jnot g12405(.din(n12596), .dout(n12597));
  jand g12406(.dina(n12597), .dinb(n12458), .dout(n12598));
  jxor g12407(.dina(n12598), .dinb(n12595), .dout(n12599));
  jand g12408(.dina(n12422), .dinb(n12421), .dout(n12600));
  jand g12409(.dina(n12423), .dinb(n12420), .dout(n12601));
  jor  g12410(.dina(n12601), .dinb(n12600), .dout(n12602));
  jand g12411(.dina(n12514), .dinb(n12275), .dout(n12603));
  jor  g12412(.dina(n12603), .dinb(n12510), .dout(n12604));
  jand g12413(.dina(n12430), .dinb(n12427), .dout(n12605));
  jnot g12414(.din(n12605), .dout(n12606));
  jand g12415(.dina(n12606), .dinb(n12433), .dout(n12607));
  jxor g12416(.dina(n12607), .dinb(n12604), .dout(n12608));
  jxor g12417(.dina(n12608), .dinb(n12602), .dout(n12609));
  jxor g12418(.dina(n12609), .dinb(n12599), .dout(n12610));
  jxor g12419(.dina(n12610), .dinb(n12588), .dout(n12611));
  jxor g12420(.dina(n12611), .dinb(n12585), .dout(n12612));
  jor  g12421(.dina(n12490), .dinb(n12487), .dout(n12613));
  jand g12422(.dina(n12491), .dinb(n12484), .dout(n12614));
  jnot g12423(.din(n12614), .dout(n12615));
  jand g12424(.dina(n12615), .dinb(n12613), .dout(n12616));
  jnot g12425(.din(n12616), .dout(n12617));
  jand g12426(.dina(\a[45] ), .dinb(\a[41] ), .dout(n12618));
  jnot g12427(.din(n12618), .dout(n12619));
  jand g12428(.dina(\a[54] ), .dinb(\a[32] ), .dout(n12620));
  jand g12429(.dina(n12620), .dinb(n6097), .dout(n12621));
  jnot g12430(.din(n12621), .dout(n12622));
  jand g12431(.dina(n12620), .dinb(n12618), .dout(n12623));
  jand g12432(.dina(n4812), .dinb(n4514), .dout(n12624));
  jor  g12433(.dina(n12624), .dinb(n12623), .dout(n12625));
  jand g12434(.dina(n12625), .dinb(n12622), .dout(n12626));
  jor  g12435(.dina(n12626), .dinb(n12619), .dout(n12627));
  jor  g12436(.dina(n12625), .dinb(n12621), .dout(n12628));
  jnot g12437(.din(n12628), .dout(n12629));
  jor  g12438(.dina(n12620), .dinb(n6097), .dout(n12630));
  jand g12439(.dina(n12630), .dinb(n12629), .dout(n12631));
  jnot g12440(.din(n12631), .dout(n12632));
  jand g12441(.dina(n12632), .dinb(n12627), .dout(n12633));
  jand g12442(.dina(\a[60] ), .dinb(\a[26] ), .dout(n12634));
  jand g12443(.dina(\a[59] ), .dinb(\a[28] ), .dout(n12635));
  jand g12444(.dina(n12635), .dinb(n12513), .dout(n12636));
  jnot g12445(.din(n12636), .dout(n12637));
  jand g12446(.dina(\a[58] ), .dinb(\a[28] ), .dout(n12638));
  jor  g12447(.dina(n12638), .dinb(n12509), .dout(n12639));
  jand g12448(.dina(n12639), .dinb(n12637), .dout(n12640));
  jxor g12449(.dina(n12640), .dinb(n12634), .dout(n12641));
  jnot g12450(.din(n12641), .dout(n12642));
  jxor g12451(.dina(n12642), .dinb(n12633), .dout(n12643));
  jnot g12452(.din(n12643), .dout(n12644));
  jand g12453(.dina(\a[56] ), .dinb(\a[30] ), .dout(n12645));
  jnot g12454(.din(n12645), .dout(n12646));
  jand g12455(.dina(\a[47] ), .dinb(\a[40] ), .dout(n12647));
  jand g12456(.dina(n12647), .dinb(n12438), .dout(n12648));
  jnot g12457(.din(n12648), .dout(n12649));
  jand g12458(.dina(\a[47] ), .dinb(\a[39] ), .dout(n12650));
  jand g12459(.dina(\a[46] ), .dinb(\a[40] ), .dout(n12651));
  jor  g12460(.dina(n12651), .dinb(n12650), .dout(n12652));
  jand g12461(.dina(n12652), .dinb(n12649), .dout(n12653));
  jxor g12462(.dina(n12653), .dinb(n12646), .dout(n12654));
  jxor g12463(.dina(n12654), .dinb(n12644), .dout(n12655));
  jand g12464(.dina(\a[63] ), .dinb(\a[23] ), .dout(n12656));
  jand g12465(.dina(\a[50] ), .dinb(\a[36] ), .dout(n12657));
  jand g12466(.dina(\a[49] ), .dinb(\a[37] ), .dout(n12658));
  jor  g12467(.dina(n12658), .dinb(n12657), .dout(n12659));
  jand g12468(.dina(\a[50] ), .dinb(\a[37] ), .dout(n12660));
  jand g12469(.dina(n12660), .dinb(n12452), .dout(n12661));
  jnot g12470(.din(n12661), .dout(n12662));
  jand g12471(.dina(n12662), .dinb(n12659), .dout(n12663));
  jxor g12472(.dina(n12663), .dinb(n12656), .dout(n12664));
  jand g12473(.dina(\a[53] ), .dinb(\a[33] ), .dout(n12665));
  jand g12474(.dina(\a[52] ), .dinb(\a[35] ), .dout(n12666));
  jand g12475(.dina(n12666), .dinb(n12432), .dout(n12667));
  jnot g12476(.din(n12667), .dout(n12668));
  jand g12477(.dina(\a[51] ), .dinb(\a[35] ), .dout(n12669));
  jor  g12478(.dina(n12669), .dinb(n12428), .dout(n12670));
  jand g12479(.dina(n12670), .dinb(n12668), .dout(n12671));
  jxor g12480(.dina(n12671), .dinb(n12665), .dout(n12672));
  jxor g12481(.dina(n12672), .dinb(n12664), .dout(n12673));
  jand g12482(.dina(n11997), .dinb(n7155), .dout(n12674));
  jnot g12483(.din(n12674), .dout(n12675));
  jand g12484(.dina(\a[57] ), .dinb(\a[29] ), .dout(n12676));
  jor  g12485(.dina(n12676), .dinb(n12464), .dout(n12677));
  jand g12486(.dina(n12677), .dinb(n12675), .dout(n12678));
  jxor g12487(.dina(n12678), .dinb(n5893), .dout(n12679));
  jxor g12488(.dina(n12679), .dinb(n12673), .dout(n12680));
  jxor g12489(.dina(n12680), .dinb(n12655), .dout(n12681));
  jxor g12490(.dina(n12681), .dinb(n12617), .dout(n12682));
  jxor g12491(.dina(n12682), .dinb(n12612), .dout(n12683));
  jxor g12492(.dina(n12683), .dinb(n12572), .dout(n12684));
  jxor g12493(.dina(n12684), .dinb(n12569), .dout(n12685));
  jnot g12494(.din(n12685), .dout(n12686));
  jxor g12495(.dina(n12686), .dinb(n12534), .dout(n12687));
  jnot g12496(.din(n12524), .dout(n12688));
  jor  g12497(.dina(n12530), .dinb(n12526), .dout(n12689));
  jand g12498(.dina(n12689), .dinb(n12688), .dout(n12690));
  jxor g12499(.dina(n12690), .dinb(n12687), .dout(\asquared[87] ));
  jand g12500(.dina(n12683), .dinb(n12572), .dout(n12692));
  jand g12501(.dina(n12684), .dinb(n12569), .dout(n12693));
  jor  g12502(.dina(n12693), .dinb(n12692), .dout(n12694));
  jnot g12503(.din(n12694), .dout(n12695));
  jand g12504(.dina(n12680), .dinb(n12655), .dout(n12696));
  jand g12505(.dina(n12681), .dinb(n12617), .dout(n12697));
  jor  g12506(.dina(n12697), .dinb(n12696), .dout(n12698));
  jand g12507(.dina(n12594), .dinb(n12591), .dout(n12699));
  jand g12508(.dina(n12598), .dinb(n12595), .dout(n12700));
  jor  g12509(.dina(n12700), .dinb(n12699), .dout(n12701));
  jand g12510(.dina(n12672), .dinb(n12664), .dout(n12702));
  jand g12511(.dina(n12679), .dinb(n12673), .dout(n12703));
  jor  g12512(.dina(n12703), .dinb(n12702), .dout(n12704));
  jxor g12513(.dina(n12704), .dinb(n12701), .dout(n12705));
  jnot g12514(.din(n12705), .dout(n12706));
  jor  g12515(.dina(n12642), .dinb(n12633), .dout(n12707));
  jor  g12516(.dina(n12654), .dinb(n12644), .dout(n12708));
  jand g12517(.dina(n12708), .dinb(n12707), .dout(n12709));
  jxor g12518(.dina(n12709), .dinb(n12706), .dout(n12710));
  jxor g12519(.dina(n12710), .dinb(n12698), .dout(n12711));
  jand g12520(.dina(n12563), .dinb(n12546), .dout(n12712));
  jand g12521(.dina(n12567), .dinb(n12564), .dout(n12713));
  jor  g12522(.dina(n12713), .dinb(n12712), .dout(n12714));
  jxor g12523(.dina(n12714), .dinb(n12711), .dout(n12715));
  jnot g12524(.din(n12715), .dout(n12716));
  jor  g12525(.dina(n12542), .dinb(n12538), .dout(n12717));
  jand g12526(.dina(n12568), .dinb(n12543), .dout(n12718));
  jnot g12527(.din(n12718), .dout(n12719));
  jand g12528(.dina(n12719), .dinb(n12717), .dout(n12720));
  jxor g12529(.dina(n12720), .dinb(n12716), .dout(n12721));
  jand g12530(.dina(n12611), .dinb(n12585), .dout(n12722));
  jand g12531(.dina(n12682), .dinb(n12612), .dout(n12723));
  jor  g12532(.dina(n12723), .dinb(n12722), .dout(n12724));
  jand g12533(.dina(n12607), .dinb(n12604), .dout(n12725));
  jand g12534(.dina(n12608), .dinb(n12602), .dout(n12726));
  jor  g12535(.dina(n12726), .dinb(n12725), .dout(n12727));
  jand g12536(.dina(\a[62] ), .dinb(\a[25] ), .dout(n12728));
  jnot g12537(.din(\a[43] ), .dout(n12729));
  jand g12538(.dina(\a[44] ), .dinb(n12729), .dout(n12730));
  jxor g12539(.dina(n12730), .dinb(n12728), .dout(n12731));
  jnot g12540(.din(n12731), .dout(n12732));
  jnot g12541(.din(n12647), .dout(n12733));
  jand g12542(.dina(n11191), .dinb(n8237), .dout(n12734));
  jnot g12543(.din(n12734), .dout(n12735));
  jand g12544(.dina(\a[56] ), .dinb(\a[31] ), .dout(n12736));
  jand g12545(.dina(\a[54] ), .dinb(\a[33] ), .dout(n12737));
  jor  g12546(.dina(n12737), .dinb(n12736), .dout(n12738));
  jand g12547(.dina(n12738), .dinb(n12735), .dout(n12739));
  jxor g12548(.dina(n12739), .dinb(n12733), .dout(n12740));
  jxor g12549(.dina(n12740), .dinb(n12732), .dout(n12741));
  jxor g12550(.dina(n12741), .dinb(n12727), .dout(n12742));
  jand g12551(.dina(\a[63] ), .dinb(\a[24] ), .dout(n12743));
  jand g12552(.dina(\a[61] ), .dinb(\a[27] ), .dout(n12744));
  jand g12553(.dina(n12744), .dinb(n12634), .dout(n12745));
  jnot g12554(.din(n12745), .dout(n12746));
  jand g12555(.dina(\a[61] ), .dinb(\a[26] ), .dout(n12747));
  jand g12556(.dina(\a[60] ), .dinb(\a[27] ), .dout(n12748));
  jor  g12557(.dina(n12748), .dinb(n12747), .dout(n12749));
  jand g12558(.dina(n12749), .dinb(n12746), .dout(n12750));
  jxor g12559(.dina(n12750), .dinb(n12743), .dout(n12751));
  jnot g12560(.din(n12751), .dout(n12752));
  jnot g12561(.din(n12660), .dout(n12753));
  jand g12562(.dina(\a[49] ), .dinb(\a[39] ), .dout(n12754));
  jand g12563(.dina(n12754), .dinb(n5893), .dout(n12755));
  jnot g12564(.din(n12755), .dout(n12756));
  jand g12565(.dina(\a[49] ), .dinb(\a[38] ), .dout(n12757));
  jand g12566(.dina(\a[48] ), .dinb(\a[39] ), .dout(n12758));
  jor  g12567(.dina(n12758), .dinb(n12757), .dout(n12759));
  jand g12568(.dina(n12759), .dinb(n12756), .dout(n12760));
  jxor g12569(.dina(n12760), .dinb(n12753), .dout(n12761));
  jxor g12570(.dina(n12761), .dinb(n12752), .dout(n12762));
  jnot g12571(.din(n12762), .dout(n12763));
  jand g12572(.dina(\a[55] ), .dinb(\a[32] ), .dout(n12764));
  jnot g12573(.din(n12764), .dout(n12765));
  jand g12574(.dina(\a[46] ), .dinb(\a[42] ), .dout(n12766));
  jand g12575(.dina(n12766), .dinb(n12618), .dout(n12767));
  jnot g12576(.din(n12767), .dout(n12768));
  jand g12577(.dina(\a[45] ), .dinb(\a[42] ), .dout(n12769));
  jand g12578(.dina(\a[46] ), .dinb(\a[41] ), .dout(n12770));
  jor  g12579(.dina(n12770), .dinb(n12769), .dout(n12771));
  jand g12580(.dina(n12771), .dinb(n12768), .dout(n12772));
  jxor g12581(.dina(n12772), .dinb(n12765), .dout(n12773));
  jxor g12582(.dina(n12773), .dinb(n12763), .dout(n12774));
  jxor g12583(.dina(n12774), .dinb(n12742), .dout(n12775));
  jand g12584(.dina(\a[52] ), .dinb(\a[36] ), .dout(n12776));
  jand g12585(.dina(n12776), .dinb(n12669), .dout(n12777));
  jand g12586(.dina(\a[58] ), .dinb(\a[29] ), .dout(n12778));
  jand g12587(.dina(n12778), .dinb(n12666), .dout(n12779));
  jor  g12588(.dina(n12779), .dinb(n12777), .dout(n12780));
  jand g12589(.dina(\a[51] ), .dinb(\a[36] ), .dout(n12781));
  jand g12590(.dina(n12781), .dinb(n12778), .dout(n12782));
  jnot g12591(.din(n12782), .dout(n12783));
  jand g12592(.dina(n12783), .dinb(n12780), .dout(n12784));
  jnot g12593(.din(n12784), .dout(n12785));
  jand g12594(.dina(n12785), .dinb(n12666), .dout(n12786));
  jor  g12595(.dina(n12782), .dinb(n12780), .dout(n12787));
  jnot g12596(.din(n12787), .dout(n12788));
  jor  g12597(.dina(n12781), .dinb(n12778), .dout(n12789));
  jand g12598(.dina(n12789), .dinb(n12788), .dout(n12790));
  jor  g12599(.dina(n12790), .dinb(n12786), .dout(n12791));
  jand g12600(.dina(\a[57] ), .dinb(\a[30] ), .dout(n12792));
  jand g12601(.dina(\a[53] ), .dinb(\a[34] ), .dout(n12793));
  jand g12602(.dina(n12793), .dinb(n12792), .dout(n12794));
  jnot g12603(.din(n12794), .dout(n12795));
  jand g12604(.dina(n11144), .dinb(n2810), .dout(n12796));
  jand g12605(.dina(n12793), .dinb(n12635), .dout(n12797));
  jor  g12606(.dina(n12797), .dinb(n12796), .dout(n12798));
  jand g12607(.dina(n12798), .dinb(n12795), .dout(n12799));
  jnot g12608(.din(n12799), .dout(n12800));
  jand g12609(.dina(n12800), .dinb(n12635), .dout(n12801));
  jor  g12610(.dina(n12798), .dinb(n12794), .dout(n12802));
  jnot g12611(.din(n12802), .dout(n12803));
  jor  g12612(.dina(n12793), .dinb(n12792), .dout(n12804));
  jand g12613(.dina(n12804), .dinb(n12803), .dout(n12805));
  jor  g12614(.dina(n12805), .dinb(n12801), .dout(n12806));
  jand g12615(.dina(n12557), .dinb(n12555), .dout(n12807));
  jor  g12616(.dina(n12807), .dinb(n12550), .dout(n12808));
  jxor g12617(.dina(n12808), .dinb(n12806), .dout(n12809));
  jxor g12618(.dina(n12809), .dinb(n12791), .dout(n12810));
  jxor g12619(.dina(n12810), .dinb(n12775), .dout(n12811));
  jxor g12620(.dina(n12811), .dinb(n12724), .dout(n12812));
  jand g12621(.dina(n12609), .dinb(n12599), .dout(n12813));
  jand g12622(.dina(n12610), .dinb(n12588), .dout(n12814));
  jor  g12623(.dina(n12814), .dinb(n12813), .dout(n12815));
  jnot g12624(.din(n12815), .dout(n12816));
  jor  g12625(.dina(n12579), .dinb(n12576), .dout(n12817));
  jor  g12626(.dina(n12584), .dinb(n12581), .dout(n12818));
  jand g12627(.dina(n12818), .dinb(n12817), .dout(n12819));
  jxor g12628(.dina(n12819), .dinb(n12816), .dout(n12820));
  jand g12629(.dina(n12558), .dinb(n12549), .dout(n12821));
  jand g12630(.dina(n12562), .dinb(n12559), .dout(n12822));
  jor  g12631(.dina(n12822), .dinb(n12821), .dout(n12823));
  jand g12632(.dina(n12677), .dinb(n5893), .dout(n12824));
  jor  g12633(.dina(n12824), .dinb(n12674), .dout(n12825));
  jand g12634(.dina(n12649), .dinb(n12646), .dout(n12826));
  jnot g12635(.din(n12826), .dout(n12827));
  jand g12636(.dina(n12827), .dinb(n12652), .dout(n12828));
  jxor g12637(.dina(n12828), .dinb(n12628), .dout(n12829));
  jxor g12638(.dina(n12829), .dinb(n12825), .dout(n12830));
  jand g12639(.dina(n12663), .dinb(n12656), .dout(n12831));
  jor  g12640(.dina(n12831), .dinb(n12661), .dout(n12832));
  jand g12641(.dina(n12640), .dinb(n12634), .dout(n12833));
  jor  g12642(.dina(n12833), .dinb(n12636), .dout(n12834));
  jor  g12643(.dina(n12667), .dinb(n12665), .dout(n12835));
  jand g12644(.dina(n12835), .dinb(n12670), .dout(n12836));
  jxor g12645(.dina(n12836), .dinb(n12834), .dout(n12837));
  jxor g12646(.dina(n12837), .dinb(n12832), .dout(n12838));
  jxor g12647(.dina(n12838), .dinb(n12830), .dout(n12839));
  jxor g12648(.dina(n12839), .dinb(n12823), .dout(n12840));
  jxor g12649(.dina(n12840), .dinb(n12820), .dout(n12841));
  jxor g12650(.dina(n12841), .dinb(n12812), .dout(n12842));
  jxor g12651(.dina(n12842), .dinb(n12721), .dout(n12843));
  jxor g12652(.dina(n12843), .dinb(n12695), .dout(n12844));
  jand g12653(.dina(n12685), .dinb(n12534), .dout(n12845));
  jnot g12654(.din(n12845), .dout(n12846));
  jnot g12655(.din(n12534), .dout(n12847));
  jand g12656(.dina(n12686), .dinb(n12847), .dout(n12848));
  jor  g12657(.dina(n12690), .dinb(n12848), .dout(n12849));
  jand g12658(.dina(n12849), .dinb(n12846), .dout(n12850));
  jxor g12659(.dina(n12850), .dinb(n12844), .dout(\asquared[88] ));
  jor  g12660(.dina(n12720), .dinb(n12716), .dout(n12852));
  jand g12661(.dina(n12842), .dinb(n12721), .dout(n12853));
  jnot g12662(.din(n12853), .dout(n12854));
  jand g12663(.dina(n12854), .dinb(n12852), .dout(n12855));
  jand g12664(.dina(n12811), .dinb(n12724), .dout(n12856));
  jand g12665(.dina(n12841), .dinb(n12812), .dout(n12857));
  jor  g12666(.dina(n12857), .dinb(n12856), .dout(n12858));
  jor  g12667(.dina(n12819), .dinb(n12816), .dout(n12859));
  jand g12668(.dina(n12840), .dinb(n12820), .dout(n12860));
  jnot g12669(.din(n12860), .dout(n12861));
  jand g12670(.dina(n12861), .dinb(n12859), .dout(n12862));
  jnot g12671(.din(n12862), .dout(n12863));
  jand g12672(.dina(n12836), .dinb(n12834), .dout(n12864));
  jand g12673(.dina(n12837), .dinb(n12832), .dout(n12865));
  jor  g12674(.dina(n12865), .dinb(n12864), .dout(n12866));
  jand g12675(.dina(n12808), .dinb(n12806), .dout(n12867));
  jand g12676(.dina(n12809), .dinb(n12791), .dout(n12868));
  jor  g12677(.dina(n12868), .dinb(n12867), .dout(n12869));
  jxor g12678(.dina(n12869), .dinb(n12866), .dout(n12870));
  jnot g12679(.din(n12870), .dout(n12871));
  jor  g12680(.dina(n12761), .dinb(n12752), .dout(n12872));
  jor  g12681(.dina(n12773), .dinb(n12763), .dout(n12873));
  jand g12682(.dina(n12873), .dinb(n12872), .dout(n12874));
  jxor g12683(.dina(n12874), .dinb(n12871), .dout(n12875));
  jand g12684(.dina(n12774), .dinb(n12742), .dout(n12876));
  jand g12685(.dina(n12810), .dinb(n12775), .dout(n12877));
  jor  g12686(.dina(n12877), .dinb(n12876), .dout(n12878));
  jxor g12687(.dina(n12878), .dinb(n12875), .dout(n12879));
  jxor g12688(.dina(n12879), .dinb(n12863), .dout(n12880));
  jxor g12689(.dina(n12880), .dinb(n12858), .dout(n12881));
  jand g12690(.dina(n12838), .dinb(n12830), .dout(n12882));
  jand g12691(.dina(n12839), .dinb(n12823), .dout(n12883));
  jor  g12692(.dina(n12883), .dinb(n12882), .dout(n12884));
  jnot g12693(.din(n12884), .dout(n12885));
  jand g12694(.dina(n12704), .dinb(n12701), .dout(n12886));
  jnot g12695(.din(n12886), .dout(n12887));
  jor  g12696(.dina(n12709), .dinb(n12706), .dout(n12888));
  jand g12697(.dina(n12888), .dinb(n12887), .dout(n12889));
  jxor g12698(.dina(n12889), .dinb(n12885), .dout(n12890));
  jand g12699(.dina(n12750), .dinb(n12743), .dout(n12891));
  jor  g12700(.dina(n12891), .dinb(n12745), .dout(n12892));
  jxor g12701(.dina(n12892), .dinb(n12802), .dout(n12893));
  jand g12702(.dina(n12756), .dinb(n12753), .dout(n12894));
  jnot g12703(.din(n12894), .dout(n12895));
  jand g12704(.dina(n12895), .dinb(n12759), .dout(n12896));
  jxor g12705(.dina(n12896), .dinb(n12893), .dout(n12897));
  jor  g12706(.dina(n12740), .dinb(n12732), .dout(n12898));
  jand g12707(.dina(n12741), .dinb(n12727), .dout(n12899));
  jnot g12708(.din(n12899), .dout(n12900));
  jand g12709(.dina(n12900), .dinb(n12898), .dout(n12901));
  jnot g12710(.din(n12901), .dout(n12902));
  jand g12711(.dina(n12735), .dinb(n12733), .dout(n12903));
  jnot g12712(.din(n12903), .dout(n12904));
  jand g12713(.dina(n12904), .dinb(n12738), .dout(n12905));
  jxor g12714(.dina(n12905), .dinb(n12787), .dout(n12906));
  jand g12715(.dina(\a[45] ), .dinb(\a[43] ), .dout(n12907));
  jnot g12716(.din(n12907), .dout(n12908));
  jand g12717(.dina(\a[55] ), .dinb(\a[34] ), .dout(n12909));
  jand g12718(.dina(n12909), .dinb(n12737), .dout(n12910));
  jnot g12719(.din(n12910), .dout(n12911));
  jand g12720(.dina(\a[55] ), .dinb(\a[33] ), .dout(n12912));
  jand g12721(.dina(\a[54] ), .dinb(\a[34] ), .dout(n12913));
  jor  g12722(.dina(n12913), .dinb(n12912), .dout(n12914));
  jand g12723(.dina(n12914), .dinb(n12911), .dout(n12915));
  jxor g12724(.dina(n12915), .dinb(n12908), .dout(n12916));
  jnot g12725(.din(n12916), .dout(n12917));
  jxor g12726(.dina(n12917), .dinb(n12906), .dout(n12918));
  jxor g12727(.dina(n12918), .dinb(n12902), .dout(n12919));
  jxor g12728(.dina(n12919), .dinb(n12897), .dout(n12920));
  jxor g12729(.dina(n12920), .dinb(n12890), .dout(n12921));
  jand g12730(.dina(n12710), .dinb(n12698), .dout(n12922));
  jand g12731(.dina(n12714), .dinb(n12711), .dout(n12923));
  jor  g12732(.dina(n12923), .dinb(n12922), .dout(n12924));
  jand g12733(.dina(n12828), .dinb(n12628), .dout(n12925));
  jand g12734(.dina(n12829), .dinb(n12825), .dout(n12926));
  jor  g12735(.dina(n12926), .dinb(n12925), .dout(n12927));
  jand g12736(.dina(\a[59] ), .dinb(\a[29] ), .dout(n12928));
  jand g12737(.dina(\a[50] ), .dinb(\a[38] ), .dout(n12929));
  jor  g12738(.dina(n12929), .dinb(n12754), .dout(n12930));
  jand g12739(.dina(\a[50] ), .dinb(\a[39] ), .dout(n12931));
  jand g12740(.dina(n12931), .dinb(n12757), .dout(n12932));
  jnot g12741(.din(n12932), .dout(n12933));
  jand g12742(.dina(n12933), .dinb(n12930), .dout(n12934));
  jxor g12743(.dina(n12934), .dinb(n12928), .dout(n12935));
  jnot g12744(.din(n12935), .dout(n12936));
  jand g12745(.dina(\a[48] ), .dinb(\a[40] ), .dout(n12937));
  jnot g12746(.din(n12937), .dout(n12938));
  jand g12747(.dina(n11688), .dinb(n3118), .dout(n12939));
  jnot g12748(.din(n12939), .dout(n12940));
  jand g12749(.dina(\a[58] ), .dinb(\a[30] ), .dout(n12941));
  jand g12750(.dina(\a[56] ), .dinb(\a[32] ), .dout(n12942));
  jor  g12751(.dina(n12942), .dinb(n12941), .dout(n12943));
  jand g12752(.dina(n12943), .dinb(n12940), .dout(n12944));
  jxor g12753(.dina(n12944), .dinb(n12938), .dout(n12945));
  jxor g12754(.dina(n12945), .dinb(n12936), .dout(n12946));
  jxor g12755(.dina(n12946), .dinb(n12927), .dout(n12947));
  jand g12756(.dina(\a[63] ), .dinb(\a[25] ), .dout(n12948));
  jor  g12757(.dina(n12728), .dinb(\a[43] ), .dout(n12949));
  jand g12758(.dina(n12949), .dinb(\a[44] ), .dout(n12950));
  jxor g12759(.dina(n12950), .dinb(n12948), .dout(n12951));
  jand g12760(.dina(n12768), .dinb(n12765), .dout(n12952));
  jnot g12761(.din(n12952), .dout(n12953));
  jand g12762(.dina(n12953), .dinb(n12771), .dout(n12954));
  jxor g12763(.dina(n12954), .dinb(n12951), .dout(n12955));
  jxor g12764(.dina(n12955), .dinb(n12947), .dout(n12956));
  jand g12765(.dina(\a[62] ), .dinb(\a[26] ), .dout(n12957));
  jand g12766(.dina(\a[61] ), .dinb(\a[28] ), .dout(n12958));
  jand g12767(.dina(n12958), .dinb(n12748), .dout(n12959));
  jnot g12768(.din(n12959), .dout(n12960));
  jand g12769(.dina(\a[60] ), .dinb(\a[28] ), .dout(n12961));
  jor  g12770(.dina(n12961), .dinb(n12744), .dout(n12962));
  jand g12771(.dina(n12962), .dinb(n12960), .dout(n12963));
  jxor g12772(.dina(n12963), .dinb(n12957), .dout(n12964));
  jnot g12773(.din(n12964), .dout(n12965));
  jand g12774(.dina(\a[57] ), .dinb(\a[31] ), .dout(n12966));
  jnot g12775(.din(n12966), .dout(n12967));
  jand g12776(.dina(\a[47] ), .dinb(\a[42] ), .dout(n12968));
  jand g12777(.dina(n12968), .dinb(n12770), .dout(n12969));
  jnot g12778(.din(n12969), .dout(n12970));
  jand g12779(.dina(\a[47] ), .dinb(\a[41] ), .dout(n12971));
  jor  g12780(.dina(n12971), .dinb(n12766), .dout(n12972));
  jand g12781(.dina(n12972), .dinb(n12970), .dout(n12973));
  jxor g12782(.dina(n12973), .dinb(n12967), .dout(n12974));
  jxor g12783(.dina(n12974), .dinb(n12965), .dout(n12975));
  jnot g12784(.din(n12975), .dout(n12976));
  jand g12785(.dina(\a[53] ), .dinb(\a[35] ), .dout(n12977));
  jnot g12786(.din(n12977), .dout(n12978));
  jand g12787(.dina(\a[52] ), .dinb(\a[37] ), .dout(n12979));
  jand g12788(.dina(n12979), .dinb(n12781), .dout(n12980));
  jnot g12789(.din(n12980), .dout(n12981));
  jand g12790(.dina(\a[51] ), .dinb(\a[37] ), .dout(n12982));
  jor  g12791(.dina(n12982), .dinb(n12776), .dout(n12983));
  jand g12792(.dina(n12983), .dinb(n12981), .dout(n12984));
  jxor g12793(.dina(n12984), .dinb(n12978), .dout(n12985));
  jxor g12794(.dina(n12985), .dinb(n12976), .dout(n12986));
  jxor g12795(.dina(n12986), .dinb(n12956), .dout(n12987));
  jxor g12796(.dina(n12987), .dinb(n12924), .dout(n12988));
  jxor g12797(.dina(n12988), .dinb(n12921), .dout(n12989));
  jxor g12798(.dina(n12989), .dinb(n12881), .dout(n12990));
  jxor g12799(.dina(n12990), .dinb(n12855), .dout(n12991));
  jand g12800(.dina(n12843), .dinb(n12694), .dout(n12992));
  jnot g12801(.din(n12992), .dout(n12993));
  jnot g12802(.din(n12843), .dout(n12994));
  jand g12803(.dina(n12994), .dinb(n12695), .dout(n12995));
  jor  g12804(.dina(n12850), .dinb(n12995), .dout(n12996));
  jand g12805(.dina(n12996), .dinb(n12993), .dout(n12997));
  jxor g12806(.dina(n12997), .dinb(n12991), .dout(\asquared[89] ));
  jand g12807(.dina(n12880), .dinb(n12858), .dout(n12999));
  jand g12808(.dina(n12989), .dinb(n12881), .dout(n13000));
  jor  g12809(.dina(n13000), .dinb(n12999), .dout(n13001));
  jand g12810(.dina(n12892), .dinb(n12802), .dout(n13002));
  jand g12811(.dina(n12896), .dinb(n12893), .dout(n13003));
  jor  g12812(.dina(n13003), .dinb(n13002), .dout(n13004));
  jand g12813(.dina(n12950), .dinb(n12948), .dout(n13005));
  jand g12814(.dina(n12954), .dinb(n12951), .dout(n13006));
  jor  g12815(.dina(n13006), .dinb(n13005), .dout(n13007));
  jxor g12816(.dina(n13007), .dinb(n13004), .dout(n13008));
  jand g12817(.dina(n12905), .dinb(n12787), .dout(n13009));
  jand g12818(.dina(n12917), .dinb(n12906), .dout(n13010));
  jor  g12819(.dina(n13010), .dinb(n13009), .dout(n13011));
  jxor g12820(.dina(n13011), .dinb(n13008), .dout(n13012));
  jnot g12821(.din(n13012), .dout(n13013));
  jand g12822(.dina(n12869), .dinb(n12866), .dout(n13014));
  jnot g12823(.din(n13014), .dout(n13015));
  jor  g12824(.dina(n12874), .dinb(n12871), .dout(n13016));
  jand g12825(.dina(n13016), .dinb(n13015), .dout(n13017));
  jxor g12826(.dina(n13017), .dinb(n13013), .dout(n13018));
  jand g12827(.dina(n12918), .dinb(n12902), .dout(n13019));
  jand g12828(.dina(n12919), .dinb(n12897), .dout(n13020));
  jor  g12829(.dina(n13020), .dinb(n13019), .dout(n13021));
  jxor g12830(.dina(n13021), .dinb(n13018), .dout(n13022));
  jand g12831(.dina(n12878), .dinb(n12875), .dout(n13023));
  jand g12832(.dina(n12879), .dinb(n12863), .dout(n13024));
  jor  g12833(.dina(n13024), .dinb(n13023), .dout(n13025));
  jand g12834(.dina(\a[48] ), .dinb(\a[41] ), .dout(n13026));
  jand g12835(.dina(\a[56] ), .dinb(\a[33] ), .dout(n13027));
  jand g12836(.dina(\a[54] ), .dinb(\a[35] ), .dout(n13028));
  jor  g12837(.dina(n13028), .dinb(n13027), .dout(n13029));
  jand g12838(.dina(n11191), .dinb(n3752), .dout(n13030));
  jnot g12839(.din(n13030), .dout(n13031));
  jand g12840(.dina(n13031), .dinb(n13029), .dout(n13032));
  jxor g12841(.dina(n13032), .dinb(n13026), .dout(n13033));
  jnot g12842(.din(n13033), .dout(n13034));
  jand g12843(.dina(\a[53] ), .dinb(\a[36] ), .dout(n13035));
  jnot g12844(.din(n13035), .dout(n13036));
  jand g12845(.dina(\a[52] ), .dinb(\a[38] ), .dout(n13037));
  jand g12846(.dina(n13037), .dinb(n12982), .dout(n13038));
  jnot g12847(.din(n13038), .dout(n13039));
  jor  g12848(.dina(n12979), .dinb(n6404), .dout(n13040));
  jand g12849(.dina(n13040), .dinb(n13039), .dout(n13041));
  jxor g12850(.dina(n13041), .dinb(n13036), .dout(n13042));
  jxor g12851(.dina(n13042), .dinb(n13034), .dout(n13043));
  jnot g12852(.din(n13043), .dout(n13044));
  jand g12853(.dina(\a[59] ), .dinb(\a[30] ), .dout(n13045));
  jnot g12854(.din(n13045), .dout(n13046));
  jand g12855(.dina(n7519), .dinb(n3269), .dout(n13047));
  jnot g12856(.din(n13047), .dout(n13048));
  jand g12857(.dina(\a[58] ), .dinb(\a[31] ), .dout(n13049));
  jand g12858(.dina(\a[57] ), .dinb(\a[32] ), .dout(n13050));
  jor  g12859(.dina(n13050), .dinb(n13049), .dout(n13051));
  jand g12860(.dina(n13051), .dinb(n13048), .dout(n13052));
  jxor g12861(.dina(n13052), .dinb(n13046), .dout(n13053));
  jxor g12862(.dina(n13053), .dinb(n13044), .dout(n13054));
  jand g12863(.dina(n12963), .dinb(n12957), .dout(n13055));
  jor  g12864(.dina(n13055), .dinb(n12959), .dout(n13056));
  jand g12865(.dina(n12981), .dinb(n12978), .dout(n13057));
  jnot g12866(.din(n13057), .dout(n13058));
  jand g12867(.dina(n13058), .dinb(n12983), .dout(n13059));
  jxor g12868(.dina(n13059), .dinb(n13056), .dout(n13060));
  jand g12869(.dina(n12940), .dinb(n12938), .dout(n13061));
  jnot g12870(.din(n13061), .dout(n13062));
  jand g12871(.dina(n13062), .dinb(n12943), .dout(n13063));
  jxor g12872(.dina(n13063), .dinb(n13060), .dout(n13064));
  jand g12873(.dina(\a[62] ), .dinb(\a[27] ), .dout(n13065));
  jnot g12874(.din(\a[44] ), .dout(n13066));
  jand g12875(.dina(\a[45] ), .dinb(n13066), .dout(n13067));
  jxor g12876(.dina(n13067), .dinb(n13065), .dout(n13068));
  jnot g12877(.din(n13068), .dout(n13069));
  jnot g12878(.din(n12909), .dout(n13070));
  jand g12879(.dina(n12766), .dinb(n6828), .dout(n13071));
  jnot g12880(.din(n13071), .dout(n13072));
  jand g12881(.dina(\a[46] ), .dinb(\a[43] ), .dout(n13073));
  jor  g12882(.dina(n13073), .dinb(n12968), .dout(n13074));
  jand g12883(.dina(n13074), .dinb(n13072), .dout(n13075));
  jxor g12884(.dina(n13075), .dinb(n13070), .dout(n13076));
  jxor g12885(.dina(n13076), .dinb(n13069), .dout(n13077));
  jand g12886(.dina(\a[61] ), .dinb(\a[29] ), .dout(n13078));
  jand g12887(.dina(n13078), .dinb(n12961), .dout(n13079));
  jnot g12888(.din(n13079), .dout(n13080));
  jand g12889(.dina(\a[60] ), .dinb(\a[29] ), .dout(n13081));
  jor  g12890(.dina(n13081), .dinb(n12958), .dout(n13082));
  jand g12891(.dina(n13082), .dinb(n13080), .dout(n13083));
  jand g12892(.dina(n12911), .dinb(n12908), .dout(n13084));
  jnot g12893(.din(n13084), .dout(n13085));
  jand g12894(.dina(n13085), .dinb(n12914), .dout(n13086));
  jxor g12895(.dina(n13086), .dinb(n13083), .dout(n13087));
  jxor g12896(.dina(n13087), .dinb(n13077), .dout(n13088));
  jxor g12897(.dina(n13088), .dinb(n13064), .dout(n13089));
  jxor g12898(.dina(n13089), .dinb(n13054), .dout(n13090));
  jxor g12899(.dina(n13090), .dinb(n13025), .dout(n13091));
  jxor g12900(.dina(n13091), .dinb(n13022), .dout(n13092));
  jor  g12901(.dina(n12889), .dinb(n12885), .dout(n13093));
  jand g12902(.dina(n12920), .dinb(n12890), .dout(n13094));
  jnot g12903(.din(n13094), .dout(n13095));
  jand g12904(.dina(n13095), .dinb(n13093), .dout(n13096));
  jnot g12905(.din(n13096), .dout(n13097));
  jand g12906(.dina(n12955), .dinb(n12947), .dout(n13098));
  jand g12907(.dina(n12986), .dinb(n12956), .dout(n13099));
  jor  g12908(.dina(n13099), .dinb(n13098), .dout(n13100));
  jor  g12909(.dina(n12945), .dinb(n12936), .dout(n13101));
  jand g12910(.dina(n12946), .dinb(n12927), .dout(n13102));
  jnot g12911(.din(n13102), .dout(n13103));
  jand g12912(.dina(n13103), .dinb(n13101), .dout(n13104));
  jor  g12913(.dina(n12974), .dinb(n12965), .dout(n13105));
  jor  g12914(.dina(n12985), .dinb(n12976), .dout(n13106));
  jand g12915(.dina(n13106), .dinb(n13105), .dout(n13107));
  jxor g12916(.dina(n13107), .dinb(n13104), .dout(n13108));
  jand g12917(.dina(n12934), .dinb(n12928), .dout(n13109));
  jor  g12918(.dina(n13109), .dinb(n12932), .dout(n13110));
  jand g12919(.dina(n12970), .dinb(n12967), .dout(n13111));
  jnot g12920(.din(n13111), .dout(n13112));
  jand g12921(.dina(n13112), .dinb(n12972), .dout(n13113));
  jxor g12922(.dina(n13113), .dinb(n13110), .dout(n13114));
  jnot g12923(.din(n13114), .dout(n13115));
  jand g12924(.dina(\a[63] ), .dinb(\a[26] ), .dout(n13116));
  jnot g12925(.din(n13116), .dout(n13117));
  jand g12926(.dina(\a[49] ), .dinb(\a[40] ), .dout(n13118));
  jor  g12927(.dina(n13118), .dinb(n12931), .dout(n13119));
  jand g12928(.dina(\a[50] ), .dinb(\a[40] ), .dout(n13120));
  jand g12929(.dina(n13120), .dinb(n12754), .dout(n13121));
  jnot g12930(.din(n13121), .dout(n13122));
  jand g12931(.dina(n13122), .dinb(n13119), .dout(n13123));
  jxor g12932(.dina(n13123), .dinb(n13117), .dout(n13124));
  jxor g12933(.dina(n13124), .dinb(n13115), .dout(n13125));
  jxor g12934(.dina(n13125), .dinb(n13108), .dout(n13126));
  jxor g12935(.dina(n13126), .dinb(n13100), .dout(n13127));
  jxor g12936(.dina(n13127), .dinb(n13097), .dout(n13128));
  jand g12937(.dina(n12987), .dinb(n12924), .dout(n13129));
  jand g12938(.dina(n12988), .dinb(n12921), .dout(n13130));
  jor  g12939(.dina(n13130), .dinb(n13129), .dout(n13131));
  jxor g12940(.dina(n13131), .dinb(n13128), .dout(n13132));
  jxor g12941(.dina(n13132), .dinb(n13092), .dout(n13133));
  jand g12942(.dina(n13133), .dinb(n13001), .dout(n13134));
  jor  g12943(.dina(n13133), .dinb(n13001), .dout(n13135));
  jnot g12944(.din(n13135), .dout(n13136));
  jor  g12945(.dina(n13136), .dinb(n13134), .dout(n13137));
  jnot g12946(.din(n12990), .dout(n13138));
  jor  g12947(.dina(n13138), .dinb(n12855), .dout(n13139));
  jand g12948(.dina(n13138), .dinb(n12855), .dout(n13140));
  jor  g12949(.dina(n12997), .dinb(n13140), .dout(n13141));
  jand g12950(.dina(n13141), .dinb(n13139), .dout(n13142));
  jxor g12951(.dina(n13142), .dinb(n13137), .dout(\asquared[90] ));
  jand g12952(.dina(n13131), .dinb(n13128), .dout(n13144));
  jand g12953(.dina(n13132), .dinb(n13092), .dout(n13145));
  jor  g12954(.dina(n13145), .dinb(n13144), .dout(n13146));
  jor  g12955(.dina(n13017), .dinb(n13013), .dout(n13147));
  jand g12956(.dina(n13021), .dinb(n13018), .dout(n13148));
  jnot g12957(.din(n13148), .dout(n13149));
  jand g12958(.dina(n13149), .dinb(n13147), .dout(n13150));
  jnot g12959(.din(n13150), .dout(n13151));
  jand g12960(.dina(n13088), .dinb(n13064), .dout(n13152));
  jand g12961(.dina(n13089), .dinb(n13054), .dout(n13153));
  jor  g12962(.dina(n13153), .dinb(n13152), .dout(n13154));
  jand g12963(.dina(n13032), .dinb(n13026), .dout(n13155));
  jor  g12964(.dina(n13155), .dinb(n13030), .dout(n13156));
  jand g12965(.dina(n13072), .dinb(n13070), .dout(n13157));
  jnot g12966(.din(n13157), .dout(n13158));
  jand g12967(.dina(n13158), .dinb(n13074), .dout(n13159));
  jor  g12968(.dina(n13065), .dinb(\a[44] ), .dout(n13160));
  jand g12969(.dina(n13160), .dinb(\a[45] ), .dout(n13161));
  jxor g12970(.dina(n13161), .dinb(n13159), .dout(n13162));
  jxor g12971(.dina(n13162), .dinb(n13156), .dout(n13163));
  jor  g12972(.dina(n13076), .dinb(n13069), .dout(n13164));
  jand g12973(.dina(n13087), .dinb(n13077), .dout(n13165));
  jnot g12974(.din(n13165), .dout(n13166));
  jand g12975(.dina(n13166), .dinb(n13164), .dout(n13167));
  jor  g12976(.dina(n13042), .dinb(n13034), .dout(n13168));
  jor  g12977(.dina(n13053), .dinb(n13044), .dout(n13169));
  jand g12978(.dina(n13169), .dinb(n13168), .dout(n13170));
  jxor g12979(.dina(n13170), .dinb(n13167), .dout(n13171));
  jxor g12980(.dina(n13171), .dinb(n13163), .dout(n13172));
  jxor g12981(.dina(n13172), .dinb(n13154), .dout(n13173));
  jxor g12982(.dina(n13173), .dinb(n13151), .dout(n13174));
  jand g12983(.dina(n13090), .dinb(n13025), .dout(n13175));
  jand g12984(.dina(n13091), .dinb(n13022), .dout(n13176));
  jor  g12985(.dina(n13176), .dinb(n13175), .dout(n13177));
  jxor g12986(.dina(n13177), .dinb(n13174), .dout(n13178));
  jand g12987(.dina(n13126), .dinb(n13100), .dout(n13179));
  jand g12988(.dina(n13127), .dinb(n13097), .dout(n13180));
  jor  g12989(.dina(n13180), .dinb(n13179), .dout(n13181));
  jand g12990(.dina(n13048), .dinb(n13046), .dout(n13182));
  jnot g12991(.din(n13182), .dout(n13183));
  jand g12992(.dina(n13183), .dinb(n13051), .dout(n13184));
  jand g12993(.dina(n13039), .dinb(n13036), .dout(n13185));
  jnot g12994(.din(n13185), .dout(n13186));
  jand g12995(.dina(n13186), .dinb(n13040), .dout(n13187));
  jxor g12996(.dina(n13187), .dinb(n13184), .dout(n13188));
  jand g12997(.dina(n13122), .dinb(n13117), .dout(n13189));
  jnot g12998(.din(n13189), .dout(n13190));
  jand g12999(.dina(n13190), .dinb(n13119), .dout(n13191));
  jxor g13000(.dina(n13191), .dinb(n13188), .dout(n13192));
  jand g13001(.dina(n13007), .dinb(n13004), .dout(n13193));
  jand g13002(.dina(n13011), .dinb(n13008), .dout(n13194));
  jor  g13003(.dina(n13194), .dinb(n13193), .dout(n13195));
  jxor g13004(.dina(n13195), .dinb(n13192), .dout(n13196));
  jand g13005(.dina(\a[55] ), .dinb(\a[35] ), .dout(n13197));
  jand g13006(.dina(\a[57] ), .dinb(\a[33] ), .dout(n13198));
  jand g13007(.dina(\a[56] ), .dinb(\a[34] ), .dout(n13199));
  jor  g13008(.dina(n13199), .dinb(n13198), .dout(n13200));
  jand g13009(.dina(\a[57] ), .dinb(\a[34] ), .dout(n13201));
  jand g13010(.dina(n13201), .dinb(n13027), .dout(n13202));
  jnot g13011(.din(n13202), .dout(n13203));
  jand g13012(.dina(n13203), .dinb(n13200), .dout(n13204));
  jxor g13013(.dina(n13204), .dinb(n13197), .dout(n13205));
  jnot g13014(.din(n13205), .dout(n13206));
  jand g13015(.dina(\a[54] ), .dinb(\a[36] ), .dout(n13207));
  jnot g13016(.din(n13207), .dout(n13208));
  jand g13017(.dina(\a[53] ), .dinb(\a[38] ), .dout(n13209));
  jand g13018(.dina(n13209), .dinb(n12979), .dout(n13210));
  jnot g13019(.din(n13210), .dout(n13211));
  jand g13020(.dina(\a[53] ), .dinb(\a[37] ), .dout(n13212));
  jor  g13021(.dina(n13212), .dinb(n13037), .dout(n13213));
  jand g13022(.dina(n13213), .dinb(n13211), .dout(n13214));
  jxor g13023(.dina(n13214), .dinb(n13208), .dout(n13215));
  jxor g13024(.dina(n13215), .dinb(n13206), .dout(n13216));
  jnot g13025(.din(n13216), .dout(n13217));
  jand g13026(.dina(\a[48] ), .dinb(\a[42] ), .dout(n13218));
  jnot g13027(.din(n13218), .dout(n13219));
  jand g13028(.dina(\a[47] ), .dinb(\a[44] ), .dout(n13220));
  jand g13029(.dina(n13220), .dinb(n13073), .dout(n13221));
  jnot g13030(.din(n13221), .dout(n13222));
  jor  g13031(.dina(n6828), .dinb(n6531), .dout(n13223));
  jand g13032(.dina(n13223), .dinb(n13222), .dout(n13224));
  jxor g13033(.dina(n13224), .dinb(n13219), .dout(n13225));
  jxor g13034(.dina(n13225), .dinb(n13217), .dout(n13226));
  jxor g13035(.dina(n13226), .dinb(n13196), .dout(n13227));
  jxor g13036(.dina(n13227), .dinb(n13181), .dout(n13228));
  jnot g13037(.din(n13104), .dout(n13229));
  jnot g13038(.din(n13107), .dout(n13230));
  jand g13039(.dina(n13230), .dinb(n13229), .dout(n13231));
  jand g13040(.dina(n13125), .dinb(n13108), .dout(n13232));
  jor  g13041(.dina(n13232), .dinb(n13231), .dout(n13233));
  jand g13042(.dina(n13113), .dinb(n13110), .dout(n13234));
  jnot g13043(.din(n13234), .dout(n13235));
  jor  g13044(.dina(n13124), .dinb(n13115), .dout(n13236));
  jand g13045(.dina(n13236), .dinb(n13235), .dout(n13237));
  jnot g13046(.din(n13237), .dout(n13238));
  jand g13047(.dina(n13059), .dinb(n13056), .dout(n13239));
  jand g13048(.dina(n13063), .dinb(n13060), .dout(n13240));
  jor  g13049(.dina(n13240), .dinb(n13239), .dout(n13241));
  jnot g13050(.din(n13241), .dout(n13242));
  jand g13051(.dina(\a[51] ), .dinb(\a[39] ), .dout(n13243));
  jnot g13052(.din(n13243), .dout(n13244));
  jand g13053(.dina(\a[50] ), .dinb(\a[41] ), .dout(n13245));
  jand g13054(.dina(n13245), .dinb(n13118), .dout(n13246));
  jnot g13055(.din(n13246), .dout(n13247));
  jand g13056(.dina(\a[49] ), .dinb(\a[41] ), .dout(n13248));
  jor  g13057(.dina(n13248), .dinb(n13120), .dout(n13249));
  jand g13058(.dina(n13249), .dinb(n13247), .dout(n13250));
  jxor g13059(.dina(n13250), .dinb(n13244), .dout(n13251));
  jxor g13060(.dina(n13251), .dinb(n13242), .dout(n13252));
  jxor g13061(.dina(n13252), .dinb(n13238), .dout(n13253));
  jand g13062(.dina(n13086), .dinb(n13083), .dout(n13254));
  jor  g13063(.dina(n13254), .dinb(n13079), .dout(n13255));
  jand g13064(.dina(n13049), .dinb(n7048), .dout(n13256));
  jnot g13065(.din(n13256), .dout(n13257));
  jand g13066(.dina(\a[59] ), .dinb(\a[31] ), .dout(n13258));
  jand g13067(.dina(\a[58] ), .dinb(\a[32] ), .dout(n13259));
  jor  g13068(.dina(n13259), .dinb(n13258), .dout(n13260));
  jand g13069(.dina(n13260), .dinb(n13257), .dout(n13261));
  jand g13070(.dina(\a[60] ), .dinb(\a[30] ), .dout(n13262));
  jxor g13071(.dina(n13262), .dinb(n13261), .dout(n13263));
  jxor g13072(.dina(n13263), .dinb(n13255), .dout(n13264));
  jand g13073(.dina(\a[63] ), .dinb(\a[27] ), .dout(n13265));
  jand g13074(.dina(n8702), .dinb(n2653), .dout(n13266));
  jnot g13075(.din(n13266), .dout(n13267));
  jand g13076(.dina(\a[62] ), .dinb(\a[28] ), .dout(n13268));
  jor  g13077(.dina(n13268), .dinb(n13078), .dout(n13269));
  jand g13078(.dina(n13269), .dinb(n13267), .dout(n13270));
  jxor g13079(.dina(n13270), .dinb(n13265), .dout(n13271));
  jxor g13080(.dina(n13271), .dinb(n13264), .dout(n13272));
  jxor g13081(.dina(n13272), .dinb(n13253), .dout(n13273));
  jxor g13082(.dina(n13273), .dinb(n13233), .dout(n13274));
  jxor g13083(.dina(n13274), .dinb(n13228), .dout(n13275));
  jxor g13084(.dina(n13275), .dinb(n13178), .dout(n13276));
  jnot g13085(.din(n13276), .dout(n13277));
  jxor g13086(.dina(n13277), .dinb(n13146), .dout(n13278));
  jnot g13087(.din(n13134), .dout(n13279));
  jor  g13088(.dina(n13142), .dinb(n13136), .dout(n13280));
  jand g13089(.dina(n13280), .dinb(n13279), .dout(n13281));
  jxor g13090(.dina(n13281), .dinb(n13278), .dout(\asquared[91] ));
  jand g13091(.dina(n13177), .dinb(n13174), .dout(n13283));
  jand g13092(.dina(n13275), .dinb(n13178), .dout(n13284));
  jor  g13093(.dina(n13284), .dinb(n13283), .dout(n13285));
  jand g13094(.dina(n13270), .dinb(n13265), .dout(n13286));
  jor  g13095(.dina(n13286), .dinb(n13266), .dout(n13287));
  jand g13096(.dina(n13211), .dinb(n13208), .dout(n13288));
  jnot g13097(.din(n13288), .dout(n13289));
  jand g13098(.dina(n13289), .dinb(n13213), .dout(n13290));
  jxor g13099(.dina(n13290), .dinb(n13287), .dout(n13291));
  jand g13100(.dina(n13262), .dinb(n13261), .dout(n13292));
  jor  g13101(.dina(n13292), .dinb(n13256), .dout(n13293));
  jxor g13102(.dina(n13293), .dinb(n13291), .dout(n13294));
  jnot g13103(.din(n13294), .dout(n13295));
  jor  g13104(.dina(n13251), .dinb(n13242), .dout(n13296));
  jand g13105(.dina(n13252), .dinb(n13238), .dout(n13297));
  jnot g13106(.din(n13297), .dout(n13298));
  jand g13107(.dina(n13298), .dinb(n13296), .dout(n13299));
  jxor g13108(.dina(n13299), .dinb(n13295), .dout(n13300));
  jand g13109(.dina(\a[63] ), .dinb(\a[28] ), .dout(n13301));
  jand g13110(.dina(\a[51] ), .dinb(\a[40] ), .dout(n13302));
  jor  g13111(.dina(n13302), .dinb(n13245), .dout(n13303));
  jand g13112(.dina(n5594), .dinb(n4632), .dout(n13304));
  jnot g13113(.din(n13304), .dout(n13305));
  jand g13114(.dina(n13305), .dinb(n13303), .dout(n13306));
  jxor g13115(.dina(n13306), .dinb(n13301), .dout(n13307));
  jnot g13116(.din(n13307), .dout(n13308));
  jand g13117(.dina(\a[56] ), .dinb(\a[35] ), .dout(n13309));
  jnot g13118(.din(n13309), .dout(n13310));
  jand g13119(.dina(n5316), .dinb(n4495), .dout(n13311));
  jnot g13120(.din(n13311), .dout(n13312));
  jand g13121(.dina(\a[48] ), .dinb(\a[43] ), .dout(n13313));
  jor  g13122(.dina(n13313), .dinb(n13220), .dout(n13314));
  jand g13123(.dina(n13314), .dinb(n13312), .dout(n13315));
  jxor g13124(.dina(n13315), .dinb(n13310), .dout(n13316));
  jxor g13125(.dina(n13316), .dinb(n13308), .dout(n13317));
  jnot g13126(.din(n13317), .dout(n13318));
  jand g13127(.dina(\a[62] ), .dinb(\a[29] ), .dout(n13319));
  jnot g13128(.din(n13319), .dout(n13320));
  jnot g13129(.din(\a[45] ), .dout(n13321));
  jand g13130(.dina(\a[46] ), .dinb(n13321), .dout(n13322));
  jxor g13131(.dina(n13322), .dinb(n13320), .dout(n13323));
  jxor g13132(.dina(n13323), .dinb(n13318), .dout(n13324));
  jxor g13133(.dina(n13324), .dinb(n13300), .dout(n13325));
  jand g13134(.dina(n13172), .dinb(n13154), .dout(n13326));
  jand g13135(.dina(n13173), .dinb(n13151), .dout(n13327));
  jor  g13136(.dina(n13327), .dinb(n13326), .dout(n13328));
  jxor g13137(.dina(n13328), .dinb(n13325), .dout(n13329));
  jand g13138(.dina(n13187), .dinb(n13184), .dout(n13330));
  jand g13139(.dina(n13191), .dinb(n13188), .dout(n13331));
  jor  g13140(.dina(n13331), .dinb(n13330), .dout(n13332));
  jand g13141(.dina(n13161), .dinb(n13159), .dout(n13333));
  jand g13142(.dina(n13162), .dinb(n13156), .dout(n13334));
  jor  g13143(.dina(n13334), .dinb(n13333), .dout(n13335));
  jnot g13144(.din(n13335), .dout(n13336));
  jnot g13145(.din(n6754), .dout(n13337));
  jand g13146(.dina(n11997), .dinb(n5916), .dout(n13338));
  jnot g13147(.din(n13338), .dout(n13339));
  jand g13148(.dina(\a[55] ), .dinb(\a[36] ), .dout(n13340));
  jor  g13149(.dina(n13340), .dinb(n13201), .dout(n13341));
  jand g13150(.dina(n13341), .dinb(n13339), .dout(n13342));
  jxor g13151(.dina(n13342), .dinb(n13337), .dout(n13343));
  jxor g13152(.dina(n13343), .dinb(n13336), .dout(n13344));
  jxor g13153(.dina(n13344), .dinb(n13332), .dout(n13345));
  jor  g13154(.dina(n13170), .dinb(n13167), .dout(n13346));
  jand g13155(.dina(n13171), .dinb(n13163), .dout(n13347));
  jnot g13156(.din(n13347), .dout(n13348));
  jand g13157(.dina(n13348), .dinb(n13346), .dout(n13349));
  jnot g13158(.din(n13349), .dout(n13350));
  jand g13159(.dina(n13247), .dinb(n13244), .dout(n13351));
  jnot g13160(.din(n13351), .dout(n13352));
  jand g13161(.dina(n13352), .dinb(n13249), .dout(n13353));
  jnot g13162(.din(n13353), .dout(n13354));
  jand g13163(.dina(\a[54] ), .dinb(\a[37] ), .dout(n13355));
  jnot g13164(.din(n13355), .dout(n13356));
  jand g13165(.dina(\a[53] ), .dinb(\a[39] ), .dout(n13357));
  jand g13166(.dina(n13357), .dinb(n13037), .dout(n13358));
  jnot g13167(.din(n13358), .dout(n13359));
  jand g13168(.dina(\a[52] ), .dinb(\a[39] ), .dout(n13360));
  jor  g13169(.dina(n13360), .dinb(n13209), .dout(n13361));
  jand g13170(.dina(n13361), .dinb(n13359), .dout(n13362));
  jxor g13171(.dina(n13362), .dinb(n13356), .dout(n13363));
  jxor g13172(.dina(n13363), .dinb(n13354), .dout(n13364));
  jand g13173(.dina(\a[60] ), .dinb(\a[31] ), .dout(n13365));
  jand g13174(.dina(\a[59] ), .dinb(\a[33] ), .dout(n13366));
  jand g13175(.dina(n13366), .dinb(n13259), .dout(n13367));
  jnot g13176(.din(n13367), .dout(n13368));
  jand g13177(.dina(\a[58] ), .dinb(\a[33] ), .dout(n13369));
  jor  g13178(.dina(n13369), .dinb(n7048), .dout(n13370));
  jand g13179(.dina(n13370), .dinb(n13368), .dout(n13371));
  jxor g13180(.dina(n13371), .dinb(n13365), .dout(n13372));
  jxor g13181(.dina(n13372), .dinb(n13364), .dout(n13373));
  jxor g13182(.dina(n13373), .dinb(n13350), .dout(n13374));
  jxor g13183(.dina(n13374), .dinb(n13345), .dout(n13375));
  jxor g13184(.dina(n13375), .dinb(n13329), .dout(n13376));
  jand g13185(.dina(n13227), .dinb(n13181), .dout(n13377));
  jand g13186(.dina(n13274), .dinb(n13228), .dout(n13378));
  jor  g13187(.dina(n13378), .dinb(n13377), .dout(n13379));
  jand g13188(.dina(n13272), .dinb(n13253), .dout(n13380));
  jand g13189(.dina(n13273), .dinb(n13233), .dout(n13381));
  jor  g13190(.dina(n13381), .dinb(n13380), .dout(n13382));
  jand g13191(.dina(n13195), .dinb(n13192), .dout(n13383));
  jand g13192(.dina(n13226), .dinb(n13196), .dout(n13384));
  jor  g13193(.dina(n13384), .dinb(n13383), .dout(n13385));
  jand g13194(.dina(n13204), .dinb(n13197), .dout(n13386));
  jor  g13195(.dina(n13386), .dinb(n13202), .dout(n13387));
  jand g13196(.dina(\a[61] ), .dinb(\a[30] ), .dout(n13388));
  jand g13197(.dina(n13222), .dinb(n13219), .dout(n13389));
  jnot g13198(.din(n13389), .dout(n13390));
  jand g13199(.dina(n13390), .dinb(n13223), .dout(n13391));
  jxor g13200(.dina(n13391), .dinb(n13388), .dout(n13392));
  jxor g13201(.dina(n13392), .dinb(n13387), .dout(n13393));
  jand g13202(.dina(n13263), .dinb(n13255), .dout(n13394));
  jand g13203(.dina(n13271), .dinb(n13264), .dout(n13395));
  jor  g13204(.dina(n13395), .dinb(n13394), .dout(n13396));
  jnot g13205(.din(n13396), .dout(n13397));
  jor  g13206(.dina(n13215), .dinb(n13206), .dout(n13398));
  jor  g13207(.dina(n13225), .dinb(n13217), .dout(n13399));
  jand g13208(.dina(n13399), .dinb(n13398), .dout(n13400));
  jxor g13209(.dina(n13400), .dinb(n13397), .dout(n13401));
  jxor g13210(.dina(n13401), .dinb(n13393), .dout(n13402));
  jxor g13211(.dina(n13402), .dinb(n13385), .dout(n13403));
  jxor g13212(.dina(n13403), .dinb(n13382), .dout(n13404));
  jxor g13213(.dina(n13404), .dinb(n13379), .dout(n13405));
  jxor g13214(.dina(n13405), .dinb(n13376), .dout(n13406));
  jand g13215(.dina(n13406), .dinb(n13285), .dout(n13407));
  jor  g13216(.dina(n13406), .dinb(n13285), .dout(n13408));
  jnot g13217(.din(n13408), .dout(n13409));
  jor  g13218(.dina(n13409), .dinb(n13407), .dout(n13410));
  jand g13219(.dina(n13276), .dinb(n13146), .dout(n13411));
  jnot g13220(.din(n13411), .dout(n13412));
  jnot g13221(.din(n13146), .dout(n13413));
  jand g13222(.dina(n13277), .dinb(n13413), .dout(n13414));
  jor  g13223(.dina(n13281), .dinb(n13414), .dout(n13415));
  jand g13224(.dina(n13415), .dinb(n13412), .dout(n13416));
  jxor g13225(.dina(n13416), .dinb(n13410), .dout(\asquared[92] ));
  jand g13226(.dina(n13402), .dinb(n13385), .dout(n13418));
  jand g13227(.dina(n13403), .dinb(n13382), .dout(n13419));
  jor  g13228(.dina(n13419), .dinb(n13418), .dout(n13420));
  jand g13229(.dina(n13373), .dinb(n13350), .dout(n13421));
  jand g13230(.dina(n13374), .dinb(n13345), .dout(n13422));
  jor  g13231(.dina(n13422), .dinb(n13421), .dout(n13423));
  jor  g13232(.dina(n13400), .dinb(n13397), .dout(n13424));
  jand g13233(.dina(n13401), .dinb(n13393), .dout(n13425));
  jnot g13234(.din(n13425), .dout(n13426));
  jand g13235(.dina(n13426), .dinb(n13424), .dout(n13427));
  jnot g13236(.din(n13427), .dout(n13428));
  jand g13237(.dina(n13391), .dinb(n13388), .dout(n13429));
  jand g13238(.dina(n13392), .dinb(n13387), .dout(n13430));
  jor  g13239(.dina(n13430), .dinb(n13429), .dout(n13431));
  jand g13240(.dina(n8702), .dinb(n2440), .dout(n13432));
  jnot g13241(.din(n13432), .dout(n13433));
  jand g13242(.dina(\a[62] ), .dinb(\a[30] ), .dout(n13434));
  jand g13243(.dina(\a[61] ), .dinb(\a[31] ), .dout(n13435));
  jor  g13244(.dina(n13435), .dinb(n13434), .dout(n13436));
  jand g13245(.dina(n13436), .dinb(n13433), .dout(n13437));
  jnot g13246(.din(\a[46] ), .dout(n13438));
  jand g13247(.dina(n13320), .dinb(n13321), .dout(n13439));
  jor  g13248(.dina(n13439), .dinb(n13438), .dout(n13440));
  jnot g13249(.din(n13440), .dout(n13441));
  jxor g13250(.dina(n13441), .dinb(n13437), .dout(n13442));
  jnot g13251(.din(n13442), .dout(n13443));
  jnot g13252(.din(n13357), .dout(n13444));
  jand g13253(.dina(\a[52] ), .dinb(\a[41] ), .dout(n13445));
  jand g13254(.dina(n13445), .dinb(n13302), .dout(n13446));
  jnot g13255(.din(n13446), .dout(n13447));
  jand g13256(.dina(\a[52] ), .dinb(\a[40] ), .dout(n13448));
  jand g13257(.dina(\a[51] ), .dinb(\a[41] ), .dout(n13449));
  jor  g13258(.dina(n13449), .dinb(n13448), .dout(n13450));
  jand g13259(.dina(n13450), .dinb(n13447), .dout(n13451));
  jxor g13260(.dina(n13451), .dinb(n13444), .dout(n13452));
  jxor g13261(.dina(n13452), .dinb(n13443), .dout(n13453));
  jxor g13262(.dina(n13453), .dinb(n13431), .dout(n13454));
  jand g13263(.dina(\a[57] ), .dinb(\a[35] ), .dout(n13455));
  jand g13264(.dina(\a[50] ), .dinb(\a[42] ), .dout(n13456));
  jand g13265(.dina(n13456), .dinb(n13455), .dout(n13457));
  jnot g13266(.din(n13457), .dout(n13458));
  jand g13267(.dina(\a[58] ), .dinb(\a[34] ), .dout(n13459));
  jand g13268(.dina(n13459), .dinb(n13456), .dout(n13460));
  jand g13269(.dina(n7519), .dinb(n2845), .dout(n13461));
  jor  g13270(.dina(n13461), .dinb(n13460), .dout(n13462));
  jnot g13271(.din(n13462), .dout(n13463));
  jand g13272(.dina(n13463), .dinb(n13458), .dout(n13464));
  jor  g13273(.dina(n13456), .dinb(n13455), .dout(n13465));
  jand g13274(.dina(n13465), .dinb(n13464), .dout(n13466));
  jand g13275(.dina(n13462), .dinb(n13458), .dout(n13467));
  jnot g13276(.din(n13467), .dout(n13468));
  jand g13277(.dina(n13468), .dinb(n13459), .dout(n13469));
  jor  g13278(.dina(n13469), .dinb(n13466), .dout(n13470));
  jand g13279(.dina(\a[49] ), .dinb(\a[43] ), .dout(n13471));
  jnot g13280(.din(n13471), .dout(n13472));
  jand g13281(.dina(n5316), .dinb(n4812), .dout(n13473));
  jnot g13282(.din(n13473), .dout(n13474));
  jand g13283(.dina(\a[48] ), .dinb(\a[44] ), .dout(n13475));
  jor  g13284(.dina(n13475), .dinb(n6996), .dout(n13476));
  jand g13285(.dina(n13476), .dinb(n13474), .dout(n13477));
  jxor g13286(.dina(n13477), .dinb(n13472), .dout(n13478));
  jnot g13287(.din(n13478), .dout(n13479));
  jxor g13288(.dina(n13479), .dinb(n13470), .dout(n13480));
  jand g13289(.dina(\a[56] ), .dinb(\a[36] ), .dout(n13481));
  jand g13290(.dina(\a[63] ), .dinb(\a[29] ), .dout(n13482));
  jxor g13291(.dina(n13482), .dinb(n13366), .dout(n13483));
  jxor g13292(.dina(n13483), .dinb(n13481), .dout(n13484));
  jxor g13293(.dina(n13484), .dinb(n13480), .dout(n13485));
  jxor g13294(.dina(n13485), .dinb(n13454), .dout(n13486));
  jxor g13295(.dina(n13486), .dinb(n13428), .dout(n13487));
  jxor g13296(.dina(n13487), .dinb(n13423), .dout(n13488));
  jxor g13297(.dina(n13488), .dinb(n13420), .dout(n13489));
  jand g13298(.dina(n13328), .dinb(n13325), .dout(n13490));
  jand g13299(.dina(n13375), .dinb(n13329), .dout(n13491));
  jor  g13300(.dina(n13491), .dinb(n13490), .dout(n13492));
  jor  g13301(.dina(n13363), .dinb(n13354), .dout(n13493));
  jand g13302(.dina(n13372), .dinb(n13364), .dout(n13494));
  jnot g13303(.din(n13494), .dout(n13495));
  jand g13304(.dina(n13495), .dinb(n13493), .dout(n13496));
  jnot g13305(.din(n13496), .dout(n13497));
  jand g13306(.dina(n13290), .dinb(n13287), .dout(n13498));
  jand g13307(.dina(n13293), .dinb(n13291), .dout(n13499));
  jor  g13308(.dina(n13499), .dinb(n13498), .dout(n13500));
  jxor g13309(.dina(n13500), .dinb(n13497), .dout(n13501));
  jnot g13310(.din(n13501), .dout(n13502));
  jor  g13311(.dina(n13316), .dinb(n13308), .dout(n13503));
  jor  g13312(.dina(n13323), .dinb(n13318), .dout(n13504));
  jand g13313(.dina(n13504), .dinb(n13503), .dout(n13505));
  jxor g13314(.dina(n13505), .dinb(n13502), .dout(n13506));
  jor  g13315(.dina(n13299), .dinb(n13295), .dout(n13507));
  jand g13316(.dina(n13324), .dinb(n13300), .dout(n13508));
  jnot g13317(.din(n13508), .dout(n13509));
  jand g13318(.dina(n13509), .dinb(n13507), .dout(n13510));
  jnot g13319(.din(n13510), .dout(n13511));
  jor  g13320(.dina(n13343), .dinb(n13336), .dout(n13512));
  jand g13321(.dina(n13344), .dinb(n13332), .dout(n13513));
  jnot g13322(.din(n13513), .dout(n13514));
  jand g13323(.dina(n13514), .dinb(n13512), .dout(n13515));
  jnot g13324(.din(n13515), .dout(n13516));
  jand g13325(.dina(n13306), .dinb(n13301), .dout(n13517));
  jor  g13326(.dina(n13517), .dinb(n13304), .dout(n13518));
  jand g13327(.dina(n13371), .dinb(n13365), .dout(n13519));
  jor  g13328(.dina(n13519), .dinb(n13367), .dout(n13520));
  jand g13329(.dina(n13359), .dinb(n13356), .dout(n13521));
  jnot g13330(.din(n13521), .dout(n13522));
  jand g13331(.dina(n13522), .dinb(n13361), .dout(n13523));
  jxor g13332(.dina(n13523), .dinb(n13520), .dout(n13524));
  jxor g13333(.dina(n13524), .dinb(n13518), .dout(n13525));
  jand g13334(.dina(n13312), .dinb(n13310), .dout(n13526));
  jnot g13335(.din(n13526), .dout(n13527));
  jand g13336(.dina(n13527), .dinb(n13314), .dout(n13528));
  jand g13337(.dina(n13339), .dinb(n13337), .dout(n13529));
  jnot g13338(.din(n13529), .dout(n13530));
  jand g13339(.dina(n13530), .dinb(n13341), .dout(n13531));
  jxor g13340(.dina(n13531), .dinb(n13528), .dout(n13532));
  jand g13341(.dina(\a[60] ), .dinb(\a[32] ), .dout(n13533));
  jand g13342(.dina(\a[55] ), .dinb(\a[38] ), .dout(n13534));
  jand g13343(.dina(n13534), .dinb(n13355), .dout(n13535));
  jnot g13344(.din(n13535), .dout(n13536));
  jand g13345(.dina(\a[55] ), .dinb(\a[37] ), .dout(n13537));
  jand g13346(.dina(\a[54] ), .dinb(\a[38] ), .dout(n13538));
  jor  g13347(.dina(n13538), .dinb(n13537), .dout(n13539));
  jand g13348(.dina(n13539), .dinb(n13536), .dout(n13540));
  jxor g13349(.dina(n13540), .dinb(n13533), .dout(n13541));
  jxor g13350(.dina(n13541), .dinb(n13532), .dout(n13542));
  jxor g13351(.dina(n13542), .dinb(n13525), .dout(n13543));
  jxor g13352(.dina(n13543), .dinb(n13516), .dout(n13544));
  jxor g13353(.dina(n13544), .dinb(n13511), .dout(n13545));
  jxor g13354(.dina(n13545), .dinb(n13506), .dout(n13546));
  jxor g13355(.dina(n13546), .dinb(n13492), .dout(n13547));
  jxor g13356(.dina(n13547), .dinb(n13489), .dout(n13548));
  jnot g13357(.din(n13548), .dout(n13549));
  jand g13358(.dina(n13404), .dinb(n13379), .dout(n13550));
  jand g13359(.dina(n13405), .dinb(n13376), .dout(n13551));
  jor  g13360(.dina(n13551), .dinb(n13550), .dout(n13552));
  jxor g13361(.dina(n13552), .dinb(n13549), .dout(n13553));
  jnot g13362(.din(n13407), .dout(n13554));
  jor  g13363(.dina(n13416), .dinb(n13409), .dout(n13555));
  jand g13364(.dina(n13555), .dinb(n13554), .dout(n13556));
  jxor g13365(.dina(n13556), .dinb(n13553), .dout(\asquared[93] ));
  jand g13366(.dina(n13546), .dinb(n13492), .dout(n13558));
  jand g13367(.dina(n13547), .dinb(n13489), .dout(n13559));
  jor  g13368(.dina(n13559), .dinb(n13558), .dout(n13560));
  jand g13369(.dina(n13487), .dinb(n13423), .dout(n13561));
  jand g13370(.dina(n13488), .dinb(n13420), .dout(n13562));
  jor  g13371(.dina(n13562), .dinb(n13561), .dout(n13563));
  jand g13372(.dina(n13531), .dinb(n13528), .dout(n13564));
  jand g13373(.dina(n13541), .dinb(n13532), .dout(n13565));
  jor  g13374(.dina(n13565), .dinb(n13564), .dout(n13566));
  jand g13375(.dina(n13523), .dinb(n13520), .dout(n13567));
  jand g13376(.dina(n13524), .dinb(n13518), .dout(n13568));
  jor  g13377(.dina(n13568), .dinb(n13567), .dout(n13569));
  jxor g13378(.dina(n13569), .dinb(n13566), .dout(n13570));
  jand g13379(.dina(n13479), .dinb(n13470), .dout(n13571));
  jand g13380(.dina(n13484), .dinb(n13480), .dout(n13572));
  jor  g13381(.dina(n13572), .dinb(n13571), .dout(n13573));
  jxor g13382(.dina(n13573), .dinb(n13570), .dout(n13574));
  jand g13383(.dina(n13542), .dinb(n13525), .dout(n13575));
  jand g13384(.dina(n13543), .dinb(n13516), .dout(n13576));
  jor  g13385(.dina(n13576), .dinb(n13575), .dout(n13577));
  jxor g13386(.dina(n13577), .dinb(n13574), .dout(n13578));
  jor  g13387(.dina(n13452), .dinb(n13443), .dout(n13579));
  jand g13388(.dina(n13453), .dinb(n13431), .dout(n13580));
  jnot g13389(.din(n13580), .dout(n13581));
  jand g13390(.dina(n13581), .dinb(n13579), .dout(n13582));
  jnot g13391(.din(n13582), .dout(n13583));
  jnot g13392(.din(n13464), .dout(n13584));
  jand g13393(.dina(n13474), .dinb(n13472), .dout(n13585));
  jnot g13394(.din(n13585), .dout(n13586));
  jand g13395(.dina(n13586), .dinb(n13476), .dout(n13587));
  jxor g13396(.dina(n13587), .dinb(n13584), .dout(n13588));
  jand g13397(.dina(n13447), .dinb(n13444), .dout(n13589));
  jnot g13398(.din(n13589), .dout(n13590));
  jand g13399(.dina(n13590), .dinb(n13450), .dout(n13591));
  jxor g13400(.dina(n13591), .dinb(n13588), .dout(n13592));
  jand g13401(.dina(n13482), .dinb(n13366), .dout(n13593));
  jand g13402(.dina(n13483), .dinb(n13481), .dout(n13594));
  jor  g13403(.dina(n13594), .dinb(n13593), .dout(n13595));
  jnot g13404(.din(n13533), .dout(n13596));
  jand g13405(.dina(n13536), .dinb(n13596), .dout(n13597));
  jnot g13406(.din(n13597), .dout(n13598));
  jand g13407(.dina(n13598), .dinb(n13539), .dout(n13599));
  jxor g13408(.dina(n13599), .dinb(n13595), .dout(n13600));
  jand g13409(.dina(n13441), .dinb(n13437), .dout(n13601));
  jor  g13410(.dina(n13601), .dinb(n13432), .dout(n13602));
  jxor g13411(.dina(n13602), .dinb(n13600), .dout(n13603));
  jxor g13412(.dina(n13603), .dinb(n13592), .dout(n13604));
  jxor g13413(.dina(n13604), .dinb(n13583), .dout(n13605));
  jxor g13414(.dina(n13605), .dinb(n13578), .dout(n13606));
  jxor g13415(.dina(n13606), .dinb(n13563), .dout(n13607));
  jand g13416(.dina(n13544), .dinb(n13511), .dout(n13608));
  jand g13417(.dina(n13545), .dinb(n13506), .dout(n13609));
  jor  g13418(.dina(n13609), .dinb(n13608), .dout(n13610));
  jand g13419(.dina(n13485), .dinb(n13454), .dout(n13611));
  jand g13420(.dina(n13486), .dinb(n13428), .dout(n13612));
  jor  g13421(.dina(n13612), .dinb(n13611), .dout(n13613));
  jand g13422(.dina(n13500), .dinb(n13497), .dout(n13614));
  jnot g13423(.din(n13614), .dout(n13615));
  jor  g13424(.dina(n13505), .dinb(n13502), .dout(n13616));
  jand g13425(.dina(n13616), .dinb(n13615), .dout(n13617));
  jnot g13426(.din(n13617), .dout(n13618));
  jand g13427(.dina(\a[58] ), .dinb(\a[35] ), .dout(n13619));
  jand g13428(.dina(\a[57] ), .dinb(\a[54] ), .dout(n13620));
  jand g13429(.dina(n13620), .dinb(n10631), .dout(n13621));
  jnot g13430(.din(n13621), .dout(n13622));
  jand g13431(.dina(n7519), .dinb(n3243), .dout(n13623));
  jand g13432(.dina(\a[54] ), .dinb(\a[39] ), .dout(n13624));
  jand g13433(.dina(n13624), .dinb(n13619), .dout(n13625));
  jor  g13434(.dina(n13625), .dinb(n13623), .dout(n13626));
  jand g13435(.dina(n13626), .dinb(n13622), .dout(n13627));
  jnot g13436(.din(n13627), .dout(n13628));
  jand g13437(.dina(n13628), .dinb(n13619), .dout(n13629));
  jor  g13438(.dina(n13626), .dinb(n13621), .dout(n13630));
  jnot g13439(.din(n13630), .dout(n13631));
  jand g13440(.dina(\a[57] ), .dinb(\a[36] ), .dout(n13632));
  jor  g13441(.dina(n13632), .dinb(n13624), .dout(n13633));
  jand g13442(.dina(n13633), .dinb(n13631), .dout(n13634));
  jor  g13443(.dina(n13634), .dinb(n13629), .dout(n13635));
  jand g13444(.dina(\a[63] ), .dinb(\a[30] ), .dout(n13636));
  jand g13445(.dina(\a[61] ), .dinb(\a[33] ), .dout(n13637));
  jand g13446(.dina(n13637), .dinb(n13533), .dout(n13638));
  jnot g13447(.din(n13638), .dout(n13639));
  jand g13448(.dina(\a[61] ), .dinb(\a[32] ), .dout(n13640));
  jand g13449(.dina(\a[60] ), .dinb(\a[33] ), .dout(n13641));
  jor  g13450(.dina(n13641), .dinb(n13640), .dout(n13642));
  jand g13451(.dina(n13642), .dinb(n13639), .dout(n13643));
  jxor g13452(.dina(n13643), .dinb(n13636), .dout(n13644));
  jxor g13453(.dina(n13644), .dinb(n13635), .dout(n13645));
  jnot g13454(.din(n13645), .dout(n13646));
  jand g13455(.dina(\a[59] ), .dinb(\a[34] ), .dout(n13647));
  jnot g13456(.din(n13647), .dout(n13648));
  jand g13457(.dina(n7165), .dinb(n4632), .dout(n13649));
  jnot g13458(.din(n13649), .dout(n13650));
  jand g13459(.dina(\a[53] ), .dinb(\a[40] ), .dout(n13651));
  jor  g13460(.dina(n13651), .dinb(n13445), .dout(n13652));
  jand g13461(.dina(n13652), .dinb(n13650), .dout(n13653));
  jxor g13462(.dina(n13653), .dinb(n13648), .dout(n13654));
  jxor g13463(.dina(n13654), .dinb(n13646), .dout(n13655));
  jand g13464(.dina(\a[56] ), .dinb(\a[37] ), .dout(n13656));
  jand g13465(.dina(\a[48] ), .dinb(\a[45] ), .dout(n13657));
  jxor g13466(.dina(n13657), .dinb(n13534), .dout(n13658));
  jxor g13467(.dina(n13658), .dinb(n13656), .dout(n13659));
  jnot g13468(.din(n13659), .dout(n13660));
  jand g13469(.dina(\a[51] ), .dinb(\a[42] ), .dout(n13661));
  jnot g13470(.din(n13661), .dout(n13662));
  jand g13471(.dina(\a[50] ), .dinb(\a[44] ), .dout(n13663));
  jand g13472(.dina(n13663), .dinb(n13471), .dout(n13664));
  jnot g13473(.din(n13664), .dout(n13665));
  jand g13474(.dina(\a[50] ), .dinb(\a[43] ), .dout(n13666));
  jor  g13475(.dina(n13666), .dinb(n7033), .dout(n13667));
  jand g13476(.dina(n13667), .dinb(n13665), .dout(n13668));
  jxor g13477(.dina(n13668), .dinb(n13662), .dout(n13669));
  jxor g13478(.dina(n13669), .dinb(n13660), .dout(n13670));
  jnot g13479(.din(n13670), .dout(n13671));
  jand g13480(.dina(\a[62] ), .dinb(\a[31] ), .dout(n13672));
  jnot g13481(.din(n13672), .dout(n13673));
  jand g13482(.dina(\a[47] ), .dinb(n13438), .dout(n13674));
  jxor g13483(.dina(n13674), .dinb(n13673), .dout(n13675));
  jxor g13484(.dina(n13675), .dinb(n13671), .dout(n13676));
  jxor g13485(.dina(n13676), .dinb(n13655), .dout(n13677));
  jxor g13486(.dina(n13677), .dinb(n13618), .dout(n13678));
  jxor g13487(.dina(n13678), .dinb(n13613), .dout(n13679));
  jxor g13488(.dina(n13679), .dinb(n13610), .dout(n13680));
  jxor g13489(.dina(n13680), .dinb(n13607), .dout(n13681));
  jand g13490(.dina(n13681), .dinb(n13560), .dout(n13682));
  jor  g13491(.dina(n13681), .dinb(n13560), .dout(n13683));
  jnot g13492(.din(n13683), .dout(n13684));
  jor  g13493(.dina(n13684), .dinb(n13682), .dout(n13685));
  jand g13494(.dina(n13552), .dinb(n13548), .dout(n13686));
  jnot g13495(.din(n13686), .dout(n13687));
  jnot g13496(.din(n13552), .dout(n13688));
  jand g13497(.dina(n13688), .dinb(n13549), .dout(n13689));
  jor  g13498(.dina(n13556), .dinb(n13689), .dout(n13690));
  jand g13499(.dina(n13690), .dinb(n13687), .dout(n13691));
  jxor g13500(.dina(n13691), .dinb(n13685), .dout(\asquared[94] ));
  jand g13501(.dina(n13678), .dinb(n13613), .dout(n13693));
  jand g13502(.dina(n13679), .dinb(n13610), .dout(n13694));
  jor  g13503(.dina(n13694), .dinb(n13693), .dout(n13695));
  jand g13504(.dina(n13676), .dinb(n13655), .dout(n13696));
  jand g13505(.dina(n13677), .dinb(n13618), .dout(n13697));
  jor  g13506(.dina(n13697), .dinb(n13696), .dout(n13698));
  jand g13507(.dina(n13599), .dinb(n13595), .dout(n13699));
  jand g13508(.dina(n13602), .dinb(n13600), .dout(n13700));
  jor  g13509(.dina(n13700), .dinb(n13699), .dout(n13701));
  jand g13510(.dina(n13587), .dinb(n13584), .dout(n13702));
  jand g13511(.dina(n13591), .dinb(n13588), .dout(n13703));
  jor  g13512(.dina(n13703), .dinb(n13702), .dout(n13704));
  jxor g13513(.dina(n13704), .dinb(n13701), .dout(n13705));
  jnot g13514(.din(n13705), .dout(n13706));
  jand g13515(.dina(n13644), .dinb(n13635), .dout(n13707));
  jnot g13516(.din(n13707), .dout(n13708));
  jor  g13517(.dina(n13654), .dinb(n13646), .dout(n13709));
  jand g13518(.dina(n13709), .dinb(n13708), .dout(n13710));
  jxor g13519(.dina(n13710), .dinb(n13706), .dout(n13711));
  jand g13520(.dina(n13603), .dinb(n13592), .dout(n13712));
  jand g13521(.dina(n13604), .dinb(n13583), .dout(n13713));
  jor  g13522(.dina(n13713), .dinb(n13712), .dout(n13714));
  jxor g13523(.dina(n13714), .dinb(n13711), .dout(n13715));
  jxor g13524(.dina(n13715), .dinb(n13698), .dout(n13716));
  jxor g13525(.dina(n13716), .dinb(n13695), .dout(n13717));
  jand g13526(.dina(n13577), .dinb(n13574), .dout(n13718));
  jand g13527(.dina(n13605), .dinb(n13578), .dout(n13719));
  jor  g13528(.dina(n13719), .dinb(n13718), .dout(n13720));
  jand g13529(.dina(n13657), .dinb(n13534), .dout(n13721));
  jand g13530(.dina(n13658), .dinb(n13656), .dout(n13722));
  jor  g13531(.dina(n13722), .dinb(n13721), .dout(n13723));
  jand g13532(.dina(\a[63] ), .dinb(\a[31] ), .dout(n13724));
  jnot g13533(.din(\a[47] ), .dout(n13725));
  jand g13534(.dina(n13673), .dinb(n13438), .dout(n13726));
  jor  g13535(.dina(n13726), .dinb(n13725), .dout(n13727));
  jnot g13536(.din(n13727), .dout(n13728));
  jxor g13537(.dina(n13728), .dinb(n13724), .dout(n13729));
  jxor g13538(.dina(n13729), .dinb(n13723), .dout(n13730));
  jnot g13539(.din(n13730), .dout(n13731));
  jor  g13540(.dina(n13669), .dinb(n13660), .dout(n13732));
  jor  g13541(.dina(n13675), .dinb(n13671), .dout(n13733));
  jand g13542(.dina(n13733), .dinb(n13732), .dout(n13734));
  jxor g13543(.dina(n13734), .dinb(n13731), .dout(n13735));
  jand g13544(.dina(n13643), .dinb(n13636), .dout(n13736));
  jor  g13545(.dina(n13736), .dinb(n13638), .dout(n13737));
  jxor g13546(.dina(n13737), .dinb(n13630), .dout(n13738));
  jand g13547(.dina(n13650), .dinb(n13648), .dout(n13739));
  jnot g13548(.din(n13739), .dout(n13740));
  jand g13549(.dina(n13740), .dinb(n13652), .dout(n13741));
  jxor g13550(.dina(n13741), .dinb(n13738), .dout(n13742));
  jxor g13551(.dina(n13742), .dinb(n13735), .dout(n13743));
  jxor g13552(.dina(n13743), .dinb(n13720), .dout(n13744));
  jand g13553(.dina(n13569), .dinb(n13566), .dout(n13745));
  jand g13554(.dina(n13573), .dinb(n13570), .dout(n13746));
  jor  g13555(.dina(n13746), .dinb(n13745), .dout(n13747));
  jnot g13556(.din(n7255), .dout(n13748));
  jand g13557(.dina(\a[56] ), .dinb(\a[38] ), .dout(n13749));
  jand g13558(.dina(n13749), .dinb(n7255), .dout(n13750));
  jand g13559(.dina(\a[49] ), .dinb(\a[46] ), .dout(n13751));
  jand g13560(.dina(n13751), .dinb(n13657), .dout(n13752));
  jor  g13561(.dina(n13752), .dinb(n13750), .dout(n13753));
  jand g13562(.dina(\a[48] ), .dinb(\a[46] ), .dout(n13754));
  jand g13563(.dina(n13754), .dinb(n13749), .dout(n13755));
  jnot g13564(.din(n13755), .dout(n13756));
  jand g13565(.dina(n13756), .dinb(n13753), .dout(n13757));
  jor  g13566(.dina(n13757), .dinb(n13748), .dout(n13758));
  jor  g13567(.dina(n13755), .dinb(n13753), .dout(n13759));
  jnot g13568(.din(n13759), .dout(n13760));
  jor  g13569(.dina(n13754), .dinb(n13749), .dout(n13761));
  jand g13570(.dina(n13761), .dinb(n13760), .dout(n13762));
  jnot g13571(.din(n13762), .dout(n13763));
  jand g13572(.dina(n13763), .dinb(n13758), .dout(n13764));
  jand g13573(.dina(\a[58] ), .dinb(\a[36] ), .dout(n13765));
  jand g13574(.dina(\a[51] ), .dinb(\a[43] ), .dout(n13766));
  jor  g13575(.dina(n13766), .dinb(n13663), .dout(n13767));
  jand g13576(.dina(n5594), .dinb(n4495), .dout(n13768));
  jnot g13577(.din(n13768), .dout(n13769));
  jand g13578(.dina(n13769), .dinb(n13767), .dout(n13770));
  jxor g13579(.dina(n13770), .dinb(n13765), .dout(n13771));
  jnot g13580(.din(n13771), .dout(n13772));
  jand g13581(.dina(\a[54] ), .dinb(\a[40] ), .dout(n13773));
  jnot g13582(.din(n13773), .dout(n13774));
  jand g13583(.dina(n7165), .dinb(n4514), .dout(n13775));
  jnot g13584(.din(n13775), .dout(n13776));
  jand g13585(.dina(\a[52] ), .dinb(\a[42] ), .dout(n13777));
  jand g13586(.dina(\a[53] ), .dinb(\a[41] ), .dout(n13778));
  jor  g13587(.dina(n13778), .dinb(n13777), .dout(n13779));
  jand g13588(.dina(n13779), .dinb(n13776), .dout(n13780));
  jxor g13589(.dina(n13780), .dinb(n13774), .dout(n13781));
  jxor g13590(.dina(n13781), .dinb(n13772), .dout(n13782));
  jnot g13591(.din(n13782), .dout(n13783));
  jxor g13592(.dina(n13783), .dinb(n13764), .dout(n13784));
  jxor g13593(.dina(n13784), .dinb(n13747), .dout(n13785));
  jand g13594(.dina(n13665), .dinb(n13662), .dout(n13786));
  jnot g13595(.din(n13786), .dout(n13787));
  jand g13596(.dina(n13787), .dinb(n13667), .dout(n13788));
  jnot g13597(.din(n13788), .dout(n13789));
  jand g13598(.dina(\a[61] ), .dinb(\a[59] ), .dout(n13790));
  jand g13599(.dina(n13790), .dinb(n3752), .dout(n13791));
  jnot g13600(.din(n13791), .dout(n13792));
  jand g13601(.dina(\a[59] ), .dinb(\a[35] ), .dout(n13793));
  jor  g13602(.dina(n13793), .dinb(n13637), .dout(n13794));
  jand g13603(.dina(n13794), .dinb(n13792), .dout(n13795));
  jxor g13604(.dina(n13795), .dinb(n7956), .dout(n13796));
  jxor g13605(.dina(n13796), .dinb(n13789), .dout(n13797));
  jand g13606(.dina(\a[57] ), .dinb(\a[37] ), .dout(n13798));
  jand g13607(.dina(\a[60] ), .dinb(\a[34] ), .dout(n13799));
  jand g13608(.dina(\a[55] ), .dinb(\a[39] ), .dout(n13800));
  jxor g13609(.dina(n13800), .dinb(n13799), .dout(n13801));
  jxor g13610(.dina(n13801), .dinb(n13798), .dout(n13802));
  jxor g13611(.dina(n13802), .dinb(n13797), .dout(n13803));
  jxor g13612(.dina(n13803), .dinb(n13785), .dout(n13804));
  jxor g13613(.dina(n13804), .dinb(n13744), .dout(n13805));
  jxor g13614(.dina(n13805), .dinb(n13717), .dout(n13806));
  jand g13615(.dina(n13606), .dinb(n13563), .dout(n13807));
  jand g13616(.dina(n13680), .dinb(n13607), .dout(n13808));
  jor  g13617(.dina(n13808), .dinb(n13807), .dout(n13809));
  jnot g13618(.din(n13809), .dout(n13810));
  jxor g13619(.dina(n13810), .dinb(n13806), .dout(n13811));
  jnot g13620(.din(n13682), .dout(n13812));
  jor  g13621(.dina(n13691), .dinb(n13684), .dout(n13813));
  jand g13622(.dina(n13813), .dinb(n13812), .dout(n13814));
  jxor g13623(.dina(n13814), .dinb(n13811), .dout(\asquared[95] ));
  jand g13624(.dina(n13716), .dinb(n13695), .dout(n13816));
  jand g13625(.dina(n13805), .dinb(n13717), .dout(n13817));
  jor  g13626(.dina(n13817), .dinb(n13816), .dout(n13818));
  jand g13627(.dina(n13743), .dinb(n13720), .dout(n13819));
  jand g13628(.dina(n13804), .dinb(n13744), .dout(n13820));
  jor  g13629(.dina(n13820), .dinb(n13819), .dout(n13821));
  jand g13630(.dina(n13784), .dinb(n13747), .dout(n13822));
  jand g13631(.dina(n13803), .dinb(n13785), .dout(n13823));
  jor  g13632(.dina(n13823), .dinb(n13822), .dout(n13824));
  jand g13633(.dina(n13728), .dinb(n13724), .dout(n13825));
  jand g13634(.dina(n13729), .dinb(n13723), .dout(n13826));
  jor  g13635(.dina(n13826), .dinb(n13825), .dout(n13827));
  jand g13636(.dina(\a[60] ), .dinb(\a[36] ), .dout(n13828));
  jand g13637(.dina(n13828), .dinb(n13793), .dout(n13829));
  jnot g13638(.din(n13829), .dout(n13830));
  jand g13639(.dina(\a[60] ), .dinb(\a[35] ), .dout(n13831));
  jand g13640(.dina(\a[59] ), .dinb(\a[36] ), .dout(n13832));
  jor  g13641(.dina(n13832), .dinb(n13831), .dout(n13833));
  jand g13642(.dina(n13833), .dinb(n13830), .dout(n13834));
  jxor g13643(.dina(n13834), .dinb(n13759), .dout(n13835));
  jxor g13644(.dina(n13835), .dinb(n13827), .dout(n13836));
  jand g13645(.dina(n13737), .dinb(n13630), .dout(n13837));
  jand g13646(.dina(n13741), .dinb(n13738), .dout(n13838));
  jor  g13647(.dina(n13838), .dinb(n13837), .dout(n13839));
  jxor g13648(.dina(n13839), .dinb(n13836), .dout(n13840));
  jnot g13649(.din(n13840), .dout(n13841));
  jor  g13650(.dina(n13734), .dinb(n13731), .dout(n13842));
  jand g13651(.dina(n13742), .dinb(n13735), .dout(n13843));
  jnot g13652(.din(n13843), .dout(n13844));
  jand g13653(.dina(n13844), .dinb(n13842), .dout(n13845));
  jxor g13654(.dina(n13845), .dinb(n13841), .dout(n13846));
  jxor g13655(.dina(n13846), .dinb(n13824), .dout(n13847));
  jxor g13656(.dina(n13847), .dinb(n13821), .dout(n13848));
  jand g13657(.dina(n13714), .dinb(n13711), .dout(n13849));
  jand g13658(.dina(n13715), .dinb(n13698), .dout(n13850));
  jor  g13659(.dina(n13850), .dinb(n13849), .dout(n13851));
  jand g13660(.dina(n13800), .dinb(n13799), .dout(n13852));
  jand g13661(.dina(n13801), .dinb(n13798), .dout(n13853));
  jor  g13662(.dina(n13853), .dinb(n13852), .dout(n13854));
  jand g13663(.dina(n13792), .dinb(n7956), .dout(n13855));
  jnot g13664(.din(n13855), .dout(n13856));
  jand g13665(.dina(n13856), .dinb(n13794), .dout(n13857));
  jxor g13666(.dina(n13857), .dinb(n13854), .dout(n13858));
  jand g13667(.dina(n13776), .dinb(n13774), .dout(n13859));
  jnot g13668(.din(n13859), .dout(n13860));
  jand g13669(.dina(n13860), .dinb(n13779), .dout(n13861));
  jxor g13670(.dina(n13861), .dinb(n13858), .dout(n13862));
  jor  g13671(.dina(n13781), .dinb(n13772), .dout(n13863));
  jor  g13672(.dina(n13783), .dinb(n13764), .dout(n13864));
  jand g13673(.dina(n13864), .dinb(n13863), .dout(n13865));
  jor  g13674(.dina(n13796), .dinb(n13789), .dout(n13866));
  jand g13675(.dina(n13802), .dinb(n13797), .dout(n13867));
  jnot g13676(.din(n13867), .dout(n13868));
  jand g13677(.dina(n13868), .dinb(n13866), .dout(n13869));
  jxor g13678(.dina(n13869), .dinb(n13865), .dout(n13870));
  jxor g13679(.dina(n13870), .dinb(n13862), .dout(n13871));
  jxor g13680(.dina(n13871), .dinb(n13851), .dout(n13872));
  jand g13681(.dina(n13704), .dinb(n13701), .dout(n13873));
  jnot g13682(.din(n13873), .dout(n13874));
  jor  g13683(.dina(n13710), .dinb(n13706), .dout(n13875));
  jand g13684(.dina(n13875), .dinb(n13874), .dout(n13876));
  jnot g13685(.din(n13876), .dout(n13877));
  jand g13686(.dina(\a[62] ), .dinb(\a[33] ), .dout(n13878));
  jand g13687(.dina(\a[48] ), .dinb(n13725), .dout(n13879));
  jxor g13688(.dina(n13879), .dinb(n13878), .dout(n13880));
  jand g13689(.dina(\a[56] ), .dinb(\a[39] ), .dout(n13881));
  jnot g13690(.din(n13881), .dout(n13882));
  jand g13691(.dina(\a[50] ), .dinb(\a[46] ), .dout(n13883));
  jand g13692(.dina(n13883), .dinb(n7255), .dout(n13884));
  jnot g13693(.din(n13751), .dout(n13885));
  jand g13694(.dina(\a[50] ), .dinb(\a[45] ), .dout(n13886));
  jnot g13695(.din(n13886), .dout(n13887));
  jand g13696(.dina(n13887), .dinb(n13885), .dout(n13888));
  jor  g13697(.dina(n13888), .dinb(n13884), .dout(n13889));
  jxor g13698(.dina(n13889), .dinb(n13882), .dout(n13890));
  jxor g13699(.dina(n13890), .dinb(n13880), .dout(n13891));
  jand g13700(.dina(\a[53] ), .dinb(\a[42] ), .dout(n13892));
  jand g13701(.dina(n13766), .dinb(n7539), .dout(n13893));
  jnot g13702(.din(n13893), .dout(n13894));
  jand g13703(.dina(\a[52] ), .dinb(\a[43] ), .dout(n13895));
  jor  g13704(.dina(n13895), .dinb(n7236), .dout(n13896));
  jand g13705(.dina(n13896), .dinb(n13894), .dout(n13897));
  jxor g13706(.dina(n13897), .dinb(n13892), .dout(n13898));
  jxor g13707(.dina(n13898), .dinb(n13891), .dout(n13899));
  jxor g13708(.dina(n13899), .dinb(n13877), .dout(n13900));
  jand g13709(.dina(n13770), .dinb(n13765), .dout(n13901));
  jor  g13710(.dina(n13901), .dinb(n13768), .dout(n13902));
  jnot g13711(.din(n13902), .dout(n13903));
  jand g13712(.dina(\a[58] ), .dinb(\a[37] ), .dout(n13904));
  jnot g13713(.din(n13904), .dout(n13905));
  jand g13714(.dina(n11997), .dinb(n11262), .dout(n13906));
  jnot g13715(.din(n13906), .dout(n13907));
  jand g13716(.dina(\a[55] ), .dinb(\a[40] ), .dout(n13908));
  jand g13717(.dina(\a[57] ), .dinb(\a[38] ), .dout(n13909));
  jor  g13718(.dina(n13909), .dinb(n13908), .dout(n13910));
  jand g13719(.dina(n13910), .dinb(n13907), .dout(n13911));
  jxor g13720(.dina(n13911), .dinb(n13905), .dout(n13912));
  jxor g13721(.dina(n13912), .dinb(n13903), .dout(n13913));
  jand g13722(.dina(\a[54] ), .dinb(\a[41] ), .dout(n13914));
  jand g13723(.dina(\a[63] ), .dinb(\a[32] ), .dout(n13915));
  jand g13724(.dina(\a[61] ), .dinb(\a[34] ), .dout(n13916));
  jor  g13725(.dina(n13916), .dinb(n13915), .dout(n13917));
  jand g13726(.dina(n8387), .dinb(n3492), .dout(n13918));
  jnot g13727(.din(n13918), .dout(n13919));
  jand g13728(.dina(n13919), .dinb(n13917), .dout(n13920));
  jxor g13729(.dina(n13920), .dinb(n13914), .dout(n13921));
  jxor g13730(.dina(n13921), .dinb(n13913), .dout(n13922));
  jxor g13731(.dina(n13922), .dinb(n13900), .dout(n13923));
  jxor g13732(.dina(n13923), .dinb(n13872), .dout(n13924));
  jxor g13733(.dina(n13924), .dinb(n13848), .dout(n13925));
  jand g13734(.dina(n13925), .dinb(n13818), .dout(n13926));
  jor  g13735(.dina(n13925), .dinb(n13818), .dout(n13927));
  jnot g13736(.din(n13927), .dout(n13928));
  jor  g13737(.dina(n13928), .dinb(n13926), .dout(n13929));
  jand g13738(.dina(n13809), .dinb(n13806), .dout(n13930));
  jnot g13739(.din(n13930), .dout(n13931));
  jnot g13740(.din(n13806), .dout(n13932));
  jand g13741(.dina(n13810), .dinb(n13932), .dout(n13933));
  jor  g13742(.dina(n13814), .dinb(n13933), .dout(n13934));
  jand g13743(.dina(n13934), .dinb(n13931), .dout(n13935));
  jxor g13744(.dina(n13935), .dinb(n13929), .dout(\asquared[96] ));
  jand g13745(.dina(n13847), .dinb(n13821), .dout(n13937));
  jand g13746(.dina(n13924), .dinb(n13848), .dout(n13938));
  jor  g13747(.dina(n13938), .dinb(n13937), .dout(n13939));
  jnot g13748(.din(n13939), .dout(n13940));
  jor  g13749(.dina(n13845), .dinb(n13841), .dout(n13941));
  jand g13750(.dina(n13846), .dinb(n13824), .dout(n13942));
  jnot g13751(.din(n13942), .dout(n13943));
  jand g13752(.dina(n13943), .dinb(n13941), .dout(n13944));
  jnot g13753(.din(n13944), .dout(n13945));
  jnot g13754(.din(n13888), .dout(n13946));
  jor  g13755(.dina(n13884), .dinb(n13881), .dout(n13947));
  jand g13756(.dina(n13947), .dinb(n13946), .dout(n13948));
  jor  g13757(.dina(n13878), .dinb(\a[47] ), .dout(n13949));
  jand g13758(.dina(n13949), .dinb(\a[48] ), .dout(n13950));
  jxor g13759(.dina(n13950), .dinb(n13948), .dout(n13951));
  jor  g13760(.dina(n13893), .dinb(n13892), .dout(n13952));
  jand g13761(.dina(n13952), .dinb(n13896), .dout(n13953));
  jxor g13762(.dina(n13953), .dinb(n13951), .dout(n13954));
  jor  g13763(.dina(n13912), .dinb(n13903), .dout(n13955));
  jand g13764(.dina(n13921), .dinb(n13913), .dout(n13956));
  jnot g13765(.din(n13956), .dout(n13957));
  jand g13766(.dina(n13957), .dinb(n13955), .dout(n13958));
  jnot g13767(.din(n13958), .dout(n13959));
  jand g13768(.dina(n13890), .dinb(n13880), .dout(n13960));
  jand g13769(.dina(n13898), .dinb(n13891), .dout(n13961));
  jor  g13770(.dina(n13961), .dinb(n13960), .dout(n13962));
  jxor g13771(.dina(n13962), .dinb(n13959), .dout(n13963));
  jxor g13772(.dina(n13963), .dinb(n13954), .dout(n13964));
  jxor g13773(.dina(n13964), .dinb(n13945), .dout(n13965));
  jand g13774(.dina(n13857), .dinb(n13854), .dout(n13966));
  jand g13775(.dina(n13861), .dinb(n13858), .dout(n13967));
  jor  g13776(.dina(n13967), .dinb(n13966), .dout(n13968));
  jand g13777(.dina(\a[55] ), .dinb(\a[41] ), .dout(n13969));
  jnot g13778(.din(n13969), .dout(n13970));
  jand g13779(.dina(n7559), .dinb(n4317), .dout(n13971));
  jnot g13780(.din(n13971), .dout(n13972));
  jand g13781(.dina(\a[53] ), .dinb(\a[43] ), .dout(n13973));
  jand g13782(.dina(n13973), .dinb(n13969), .dout(n13974));
  jand g13783(.dina(\a[55] ), .dinb(\a[42] ), .dout(n13975));
  jand g13784(.dina(n13975), .dinb(n13914), .dout(n13976));
  jor  g13785(.dina(n13976), .dinb(n13974), .dout(n13977));
  jand g13786(.dina(n13977), .dinb(n13972), .dout(n13978));
  jor  g13787(.dina(n13978), .dinb(n13970), .dout(n13979));
  jand g13788(.dina(\a[54] ), .dinb(\a[42] ), .dout(n13980));
  jor  g13789(.dina(n13980), .dinb(n13973), .dout(n13981));
  jor  g13790(.dina(n13977), .dinb(n13971), .dout(n13982));
  jnot g13791(.din(n13982), .dout(n13983));
  jand g13792(.dina(n13983), .dinb(n13981), .dout(n13984));
  jnot g13793(.din(n13984), .dout(n13985));
  jand g13794(.dina(n13985), .dinb(n13979), .dout(n13986));
  jand g13795(.dina(\a[63] ), .dinb(\a[33] ), .dout(n13987));
  jand g13796(.dina(n8702), .dinb(n2845), .dout(n13988));
  jnot g13797(.din(n13988), .dout(n13989));
  jand g13798(.dina(\a[62] ), .dinb(\a[34] ), .dout(n13990));
  jand g13799(.dina(\a[61] ), .dinb(\a[35] ), .dout(n13991));
  jor  g13800(.dina(n13991), .dinb(n13990), .dout(n13992));
  jand g13801(.dina(n13992), .dinb(n13989), .dout(n13993));
  jxor g13802(.dina(n13993), .dinb(n13987), .dout(n13994));
  jnot g13803(.din(n13994), .dout(n13995));
  jxor g13804(.dina(n13995), .dinb(n13986), .dout(n13996));
  jxor g13805(.dina(n13996), .dinb(n13968), .dout(n13997));
  jand g13806(.dina(n13920), .dinb(n13914), .dout(n13998));
  jor  g13807(.dina(n13998), .dinb(n13918), .dout(n13999));
  jand g13808(.dina(n13907), .dinb(n13905), .dout(n14000));
  jnot g13809(.din(n14000), .dout(n14001));
  jand g13810(.dina(n14001), .dinb(n13910), .dout(n14002));
  jxor g13811(.dina(n14002), .dinb(n13999), .dout(n14003));
  jand g13812(.dina(n13834), .dinb(n13759), .dout(n14004));
  jor  g13813(.dina(n14004), .dinb(n13829), .dout(n14005));
  jxor g13814(.dina(n14005), .dinb(n14003), .dout(n14006));
  jand g13815(.dina(n13835), .dinb(n13827), .dout(n14007));
  jand g13816(.dina(n13839), .dinb(n13836), .dout(n14008));
  jor  g13817(.dina(n14008), .dinb(n14007), .dout(n14009));
  jxor g13818(.dina(n14009), .dinb(n14006), .dout(n14010));
  jxor g13819(.dina(n14010), .dinb(n13997), .dout(n14011));
  jxor g13820(.dina(n14011), .dinb(n13965), .dout(n14012));
  jand g13821(.dina(n13871), .dinb(n13851), .dout(n14013));
  jand g13822(.dina(n13923), .dinb(n13872), .dout(n14014));
  jor  g13823(.dina(n14014), .dinb(n14013), .dout(n14015));
  jand g13824(.dina(n13899), .dinb(n13877), .dout(n14016));
  jand g13825(.dina(n13922), .dinb(n13900), .dout(n14017));
  jor  g13826(.dina(n14017), .dinb(n14016), .dout(n14018));
  jor  g13827(.dina(n13869), .dinb(n13865), .dout(n14019));
  jand g13828(.dina(n13870), .dinb(n13862), .dout(n14020));
  jnot g13829(.din(n14020), .dout(n14021));
  jand g13830(.dina(n14021), .dinb(n14019), .dout(n14022));
  jnot g13831(.din(n14022), .dout(n14023));
  jand g13832(.dina(\a[51] ), .dinb(\a[45] ), .dout(n14024));
  jand g13833(.dina(\a[50] ), .dinb(\a[47] ), .dout(n14025));
  jand g13834(.dina(n14025), .dinb(n13751), .dout(n14026));
  jnot g13835(.din(n14026), .dout(n14027));
  jand g13836(.dina(n14024), .dinb(n7412), .dout(n14028));
  jand g13837(.dina(n13886), .dinb(n7393), .dout(n14029));
  jor  g13838(.dina(n14029), .dinb(n14028), .dout(n14030));
  jand g13839(.dina(n14030), .dinb(n14027), .dout(n14031));
  jnot g13840(.din(n14031), .dout(n14032));
  jand g13841(.dina(n14032), .dinb(n14024), .dout(n14033));
  jor  g13842(.dina(n14030), .dinb(n14026), .dout(n14034));
  jnot g13843(.din(n14034), .dout(n14035));
  jor  g13844(.dina(n13883), .dinb(n7412), .dout(n14036));
  jand g13845(.dina(n14036), .dinb(n14035), .dout(n14037));
  jor  g13846(.dina(n14037), .dinb(n14033), .dout(n14038));
  jand g13847(.dina(\a[59] ), .dinb(\a[56] ), .dout(n14039));
  jand g13848(.dina(n14039), .dinb(n11081), .dout(n14040));
  jnot g13849(.din(n14040), .dout(n14041));
  jand g13850(.dina(\a[60] ), .dinb(\a[37] ), .dout(n14042));
  jand g13851(.dina(n14042), .dinb(n13832), .dout(n14043));
  jand g13852(.dina(\a[56] ), .dinb(\a[40] ), .dout(n14044));
  jand g13853(.dina(n14044), .dinb(n13828), .dout(n14045));
  jor  g13854(.dina(n14045), .dinb(n14043), .dout(n14046));
  jnot g13855(.din(n14046), .dout(n14047));
  jand g13856(.dina(n14047), .dinb(n14041), .dout(n14048));
  jand g13857(.dina(\a[59] ), .dinb(\a[37] ), .dout(n14049));
  jor  g13858(.dina(n14049), .dinb(n14044), .dout(n14050));
  jand g13859(.dina(n14050), .dinb(n14048), .dout(n14051));
  jand g13860(.dina(n14046), .dinb(n14041), .dout(n14052));
  jnot g13861(.din(n14052), .dout(n14053));
  jand g13862(.dina(n14053), .dinb(n13828), .dout(n14054));
  jor  g13863(.dina(n14054), .dinb(n14051), .dout(n14055));
  jnot g13864(.din(n7539), .dout(n14056));
  jand g13865(.dina(\a[58] ), .dinb(\a[39] ), .dout(n14057));
  jand g13866(.dina(n14057), .dinb(n13909), .dout(n14058));
  jnot g13867(.din(n14058), .dout(n14059));
  jand g13868(.dina(\a[58] ), .dinb(\a[38] ), .dout(n14060));
  jand g13869(.dina(\a[57] ), .dinb(\a[39] ), .dout(n14061));
  jor  g13870(.dina(n14061), .dinb(n14060), .dout(n14062));
  jand g13871(.dina(n14062), .dinb(n14059), .dout(n14063));
  jxor g13872(.dina(n14063), .dinb(n14056), .dout(n14064));
  jnot g13873(.din(n14064), .dout(n14065));
  jxor g13874(.dina(n14065), .dinb(n14055), .dout(n14066));
  jxor g13875(.dina(n14066), .dinb(n14038), .dout(n14067));
  jxor g13876(.dina(n14067), .dinb(n14023), .dout(n14068));
  jxor g13877(.dina(n14068), .dinb(n14018), .dout(n14069));
  jxor g13878(.dina(n14069), .dinb(n14015), .dout(n14070));
  jxor g13879(.dina(n14070), .dinb(n14012), .dout(n14071));
  jxor g13880(.dina(n14071), .dinb(n13940), .dout(n14072));
  jnot g13881(.din(n13926), .dout(n14073));
  jor  g13882(.dina(n13935), .dinb(n13928), .dout(n14074));
  jand g13883(.dina(n14074), .dinb(n14073), .dout(n14075));
  jxor g13884(.dina(n14075), .dinb(n14072), .dout(\asquared[97] ));
  jand g13885(.dina(n14069), .dinb(n14015), .dout(n14077));
  jand g13886(.dina(n14070), .dinb(n14012), .dout(n14078));
  jor  g13887(.dina(n14078), .dinb(n14077), .dout(n14079));
  jand g13888(.dina(n14067), .dinb(n14023), .dout(n14080));
  jand g13889(.dina(n14068), .dinb(n14018), .dout(n14081));
  jor  g13890(.dina(n14081), .dinb(n14080), .dout(n14082));
  jand g13891(.dina(\a[61] ), .dinb(\a[36] ), .dout(n14083));
  jxor g13892(.dina(n14083), .dinb(n14034), .dout(n14084));
  jand g13893(.dina(n14059), .dinb(n14056), .dout(n14085));
  jnot g13894(.din(n14085), .dout(n14086));
  jand g13895(.dina(n14086), .dinb(n14062), .dout(n14087));
  jxor g13896(.dina(n14087), .dinb(n14084), .dout(n14088));
  jand g13897(.dina(n14065), .dinb(n14055), .dout(n14089));
  jand g13898(.dina(n14066), .dinb(n14038), .dout(n14090));
  jor  g13899(.dina(n14090), .dinb(n14089), .dout(n14091));
  jand g13900(.dina(n14002), .dinb(n13999), .dout(n14092));
  jand g13901(.dina(n14005), .dinb(n14003), .dout(n14093));
  jor  g13902(.dina(n14093), .dinb(n14092), .dout(n14094));
  jxor g13903(.dina(n14094), .dinb(n14091), .dout(n14095));
  jxor g13904(.dina(n14095), .dinb(n14088), .dout(n14096));
  jand g13905(.dina(n13950), .dinb(n13948), .dout(n14097));
  jand g13906(.dina(n13953), .dinb(n13951), .dout(n14098));
  jor  g13907(.dina(n14098), .dinb(n14097), .dout(n14099));
  jand g13908(.dina(\a[62] ), .dinb(\a[35] ), .dout(n14100));
  jand g13909(.dina(\a[49] ), .dinb(n4980), .dout(n14101));
  jxor g13910(.dina(n14101), .dinb(n14100), .dout(n14102));
  jnot g13911(.din(n14102), .dout(n14103));
  jand g13912(.dina(\a[57] ), .dinb(\a[40] ), .dout(n14104));
  jnot g13913(.din(n14104), .dout(n14105));
  jand g13914(.dina(n13883), .dinb(n7719), .dout(n14106));
  jnot g13915(.din(n14106), .dout(n14107));
  jor  g13916(.dina(n14025), .dinb(n7393), .dout(n14108));
  jand g13917(.dina(n14108), .dinb(n14107), .dout(n14109));
  jxor g13918(.dina(n14109), .dinb(n14105), .dout(n14110));
  jxor g13919(.dina(n14110), .dinb(n14103), .dout(n14111));
  jxor g13920(.dina(n14111), .dinb(n14099), .dout(n14112));
  jnot g13921(.din(n14048), .dout(n14113));
  jand g13922(.dina(n13993), .dinb(n13987), .dout(n14114));
  jor  g13923(.dina(n14114), .dinb(n13988), .dout(n14115));
  jxor g13924(.dina(n14115), .dinb(n14113), .dout(n14116));
  jxor g13925(.dina(n14116), .dinb(n13982), .dout(n14117));
  jor  g13926(.dina(n13995), .dinb(n13986), .dout(n14118));
  jand g13927(.dina(n13996), .dinb(n13968), .dout(n14119));
  jnot g13928(.din(n14119), .dout(n14120));
  jand g13929(.dina(n14120), .dinb(n14118), .dout(n14121));
  jnot g13930(.din(n14121), .dout(n14122));
  jxor g13931(.dina(n14122), .dinb(n14117), .dout(n14123));
  jxor g13932(.dina(n14123), .dinb(n14112), .dout(n14124));
  jxor g13933(.dina(n14124), .dinb(n14096), .dout(n14125));
  jxor g13934(.dina(n14125), .dinb(n14082), .dout(n14126));
  jand g13935(.dina(n13964), .dinb(n13945), .dout(n14127));
  jand g13936(.dina(n14011), .dinb(n13965), .dout(n14128));
  jor  g13937(.dina(n14128), .dinb(n14127), .dout(n14129));
  jand g13938(.dina(n14009), .dinb(n14006), .dout(n14130));
  jand g13939(.dina(n14010), .dinb(n13997), .dout(n14131));
  jor  g13940(.dina(n14131), .dinb(n14130), .dout(n14132));
  jand g13941(.dina(n13962), .dinb(n13959), .dout(n14133));
  jand g13942(.dina(n13963), .dinb(n13954), .dout(n14134));
  jor  g13943(.dina(n14134), .dinb(n14133), .dout(n14135));
  jand g13944(.dina(\a[63] ), .dinb(\a[34] ), .dout(n14136));
  jand g13945(.dina(n14136), .dinb(n13975), .dout(n14137));
  jnot g13946(.din(n14137), .dout(n14138));
  jand g13947(.dina(\a[56] ), .dinb(\a[42] ), .dout(n14139));
  jand g13948(.dina(n14139), .dinb(n13969), .dout(n14140));
  jand g13949(.dina(\a[56] ), .dinb(\a[41] ), .dout(n14141));
  jand g13950(.dina(n14141), .dinb(n14136), .dout(n14142));
  jor  g13951(.dina(n14142), .dinb(n14140), .dout(n14143));
  jand g13952(.dina(n14143), .dinb(n14138), .dout(n14144));
  jnot g13953(.din(n14144), .dout(n14145));
  jxor g13954(.dina(n14136), .dinb(n13975), .dout(n14146));
  jor  g13955(.dina(n14146), .dinb(n14141), .dout(n14147));
  jand g13956(.dina(n14147), .dinb(n14145), .dout(n14148));
  jnot g13957(.din(n14042), .dout(n14149));
  jand g13958(.dina(\a[59] ), .dinb(\a[39] ), .dout(n14150));
  jand g13959(.dina(n14150), .dinb(n14060), .dout(n14151));
  jnot g13960(.din(n14151), .dout(n14152));
  jand g13961(.dina(\a[59] ), .dinb(\a[38] ), .dout(n14153));
  jor  g13962(.dina(n14153), .dinb(n14057), .dout(n14154));
  jand g13963(.dina(n14154), .dinb(n14152), .dout(n14155));
  jxor g13964(.dina(n14155), .dinb(n14149), .dout(n14156));
  jnot g13965(.din(n14156), .dout(n14157));
  jxor g13966(.dina(n14157), .dinb(n14148), .dout(n14158));
  jnot g13967(.din(n14158), .dout(n14159));
  jand g13968(.dina(\a[54] ), .dinb(\a[43] ), .dout(n14160));
  jnot g13969(.din(n14160), .dout(n14161));
  jand g13970(.dina(n7165), .dinb(n4812), .dout(n14162));
  jnot g13971(.din(n14162), .dout(n14163));
  jand g13972(.dina(\a[53] ), .dinb(\a[44] ), .dout(n14164));
  jor  g13973(.dina(n14164), .dinb(n7682), .dout(n14165));
  jand g13974(.dina(n14165), .dinb(n14163), .dout(n14166));
  jxor g13975(.dina(n14166), .dinb(n14161), .dout(n14167));
  jxor g13976(.dina(n14167), .dinb(n14159), .dout(n14168));
  jxor g13977(.dina(n14168), .dinb(n14135), .dout(n14169));
  jxor g13978(.dina(n14169), .dinb(n14132), .dout(n14170));
  jxor g13979(.dina(n14170), .dinb(n14129), .dout(n14171));
  jxor g13980(.dina(n14171), .dinb(n14126), .dout(n14172));
  jand g13981(.dina(n14172), .dinb(n14079), .dout(n14173));
  jor  g13982(.dina(n14172), .dinb(n14079), .dout(n14174));
  jnot g13983(.din(n14174), .dout(n14175));
  jor  g13984(.dina(n14175), .dinb(n14173), .dout(n14176));
  jand g13985(.dina(n14071), .dinb(n13939), .dout(n14177));
  jnot g13986(.din(n14177), .dout(n14178));
  jnot g13987(.din(n14071), .dout(n14179));
  jand g13988(.dina(n14179), .dinb(n13940), .dout(n14180));
  jor  g13989(.dina(n14075), .dinb(n14180), .dout(n14181));
  jand g13990(.dina(n14181), .dinb(n14178), .dout(n14182));
  jxor g13991(.dina(n14182), .dinb(n14176), .dout(\asquared[98] ));
  jand g13992(.dina(n14170), .dinb(n14129), .dout(n14184));
  jand g13993(.dina(n14171), .dinb(n14126), .dout(n14185));
  jor  g13994(.dina(n14185), .dinb(n14184), .dout(n14186));
  jand g13995(.dina(n14124), .dinb(n14096), .dout(n14187));
  jand g13996(.dina(n14125), .dinb(n14082), .dout(n14188));
  jor  g13997(.dina(n14188), .dinb(n14187), .dout(n14189));
  jand g13998(.dina(n14122), .dinb(n14117), .dout(n14190));
  jand g13999(.dina(n14123), .dinb(n14112), .dout(n14191));
  jor  g14000(.dina(n14191), .dinb(n14190), .dout(n14192));
  jand g14001(.dina(n14094), .dinb(n14091), .dout(n14193));
  jand g14002(.dina(n14095), .dinb(n14088), .dout(n14194));
  jor  g14003(.dina(n14194), .dinb(n14193), .dout(n14195));
  jand g14004(.dina(n14160), .dinb(n8067), .dout(n14196));
  jnot g14005(.din(n14196), .dout(n14197));
  jand g14006(.dina(\a[54] ), .dinb(\a[44] ), .dout(n14198));
  jand g14007(.dina(\a[55] ), .dinb(\a[43] ), .dout(n14199));
  jor  g14008(.dina(n14199), .dinb(n14198), .dout(n14200));
  jand g14009(.dina(n14200), .dinb(n14197), .dout(n14201));
  jand g14010(.dina(\a[63] ), .dinb(\a[35] ), .dout(n14202));
  jxor g14011(.dina(n14202), .dinb(n14201), .dout(n14203));
  jand g14012(.dina(n14107), .dinb(n14105), .dout(n14204));
  jnot g14013(.din(n14204), .dout(n14205));
  jand g14014(.dina(n14205), .dinb(n14108), .dout(n14206));
  jxor g14015(.dina(n14206), .dinb(n14203), .dout(n14207));
  jnot g14016(.din(n14207), .dout(n14208));
  jand g14017(.dina(\a[60] ), .dinb(\a[38] ), .dout(n14209));
  jnot g14018(.din(n14209), .dout(n14210));
  jand g14019(.dina(\a[57] ), .dinb(\a[42] ), .dout(n14211));
  jand g14020(.dina(n14211), .dinb(n14141), .dout(n14212));
  jnot g14021(.din(n14212), .dout(n14213));
  jand g14022(.dina(\a[57] ), .dinb(\a[41] ), .dout(n14214));
  jor  g14023(.dina(n14214), .dinb(n14139), .dout(n14215));
  jand g14024(.dina(n14215), .dinb(n14213), .dout(n14216));
  jxor g14025(.dina(n14216), .dinb(n14210), .dout(n14217));
  jxor g14026(.dina(n14217), .dinb(n14208), .dout(n14218));
  jxor g14027(.dina(n14218), .dinb(n14195), .dout(n14219));
  jxor g14028(.dina(n14219), .dinb(n14192), .dout(n14220));
  jxor g14029(.dina(n14220), .dinb(n14189), .dout(n14221));
  jand g14030(.dina(n14168), .dinb(n14135), .dout(n14222));
  jand g14031(.dina(n14169), .dinb(n14132), .dout(n14223));
  jor  g14032(.dina(n14223), .dinb(n14222), .dout(n14224));
  jand g14033(.dina(n14115), .dinb(n14113), .dout(n14225));
  jand g14034(.dina(n14116), .dinb(n13982), .dout(n14226));
  jor  g14035(.dina(n14226), .dinb(n14225), .dout(n14227));
  jand g14036(.dina(n14083), .dinb(n14034), .dout(n14228));
  jand g14037(.dina(n14087), .dinb(n14084), .dout(n14229));
  jor  g14038(.dina(n14229), .dinb(n14228), .dout(n14230));
  jxor g14039(.dina(n14230), .dinb(n14227), .dout(n14231));
  jnot g14040(.din(n14231), .dout(n14232));
  jand g14041(.dina(n14157), .dinb(n14148), .dout(n14233));
  jnot g14042(.din(n14233), .dout(n14234));
  jor  g14043(.dina(n14167), .dinb(n14159), .dout(n14235));
  jand g14044(.dina(n14235), .dinb(n14234), .dout(n14236));
  jxor g14045(.dina(n14236), .dinb(n14232), .dout(n14237));
  jor  g14046(.dina(n14143), .dinb(n14137), .dout(n14238));
  jand g14047(.dina(n14152), .dinb(n14149), .dout(n14239));
  jnot g14048(.din(n14239), .dout(n14240));
  jand g14049(.dina(n14240), .dinb(n14154), .dout(n14241));
  jxor g14050(.dina(n14241), .dinb(n14238), .dout(n14242));
  jand g14051(.dina(n14163), .dinb(n14161), .dout(n14243));
  jnot g14052(.din(n14243), .dout(n14244));
  jand g14053(.dina(n14244), .dinb(n14165), .dout(n14245));
  jxor g14054(.dina(n14245), .dinb(n14242), .dout(n14246));
  jnot g14055(.din(n14246), .dout(n14247));
  jor  g14056(.dina(n14110), .dinb(n14103), .dout(n14248));
  jand g14057(.dina(n14111), .dinb(n14099), .dout(n14249));
  jnot g14058(.din(n14249), .dout(n14250));
  jand g14059(.dina(n14250), .dinb(n14248), .dout(n14251));
  jxor g14060(.dina(n14251), .dinb(n14247), .dout(n14252));
  jand g14061(.dina(n8702), .dinb(n3138), .dout(n14253));
  jnot g14062(.din(n14253), .dout(n14254));
  jand g14063(.dina(\a[62] ), .dinb(\a[36] ), .dout(n14255));
  jand g14064(.dina(\a[61] ), .dinb(\a[37] ), .dout(n14256));
  jor  g14065(.dina(n14256), .dinb(n14255), .dout(n14257));
  jand g14066(.dina(n14257), .dinb(n14254), .dout(n14258));
  jor  g14067(.dina(n14100), .dinb(\a[48] ), .dout(n14259));
  jand g14068(.dina(n14259), .dinb(\a[49] ), .dout(n14260));
  jxor g14069(.dina(n14260), .dinb(n14258), .dout(n14261));
  jand g14070(.dina(\a[52] ), .dinb(\a[46] ), .dout(n14262));
  jnot g14071(.din(n14262), .dout(n14263));
  jand g14072(.dina(n5594), .dinb(n5316), .dout(n14264));
  jnot g14073(.din(n14264), .dout(n14265));
  jand g14074(.dina(n8013), .dinb(n7393), .dout(n14266));
  jand g14075(.dina(n14262), .dinb(n7978), .dout(n14267));
  jor  g14076(.dina(n14267), .dinb(n14266), .dout(n14268));
  jand g14077(.dina(n14268), .dinb(n14265), .dout(n14269));
  jor  g14078(.dina(n14269), .dinb(n14263), .dout(n14270));
  jor  g14079(.dina(n14268), .dinb(n14264), .dout(n14271));
  jnot g14080(.din(n14271), .dout(n14272));
  jor  g14081(.dina(n7978), .dinb(n7719), .dout(n14273));
  jand g14082(.dina(n14273), .dinb(n14272), .dout(n14274));
  jnot g14083(.din(n14274), .dout(n14275));
  jand g14084(.dina(n14275), .dinb(n14270), .dout(n14276));
  jand g14085(.dina(\a[53] ), .dinb(\a[45] ), .dout(n14277));
  jand g14086(.dina(\a[58] ), .dinb(\a[40] ), .dout(n14278));
  jor  g14087(.dina(n14278), .dinb(n14150), .dout(n14279));
  jand g14088(.dina(\a[59] ), .dinb(\a[40] ), .dout(n14280));
  jand g14089(.dina(n14280), .dinb(n14057), .dout(n14281));
  jnot g14090(.din(n14281), .dout(n14282));
  jand g14091(.dina(n14282), .dinb(n14279), .dout(n14283));
  jxor g14092(.dina(n14283), .dinb(n14277), .dout(n14284));
  jnot g14093(.din(n14284), .dout(n14285));
  jxor g14094(.dina(n14285), .dinb(n14276), .dout(n14286));
  jxor g14095(.dina(n14286), .dinb(n14261), .dout(n14287));
  jxor g14096(.dina(n14287), .dinb(n14252), .dout(n14288));
  jxor g14097(.dina(n14288), .dinb(n14237), .dout(n14289));
  jxor g14098(.dina(n14289), .dinb(n14224), .dout(n14290));
  jxor g14099(.dina(n14290), .dinb(n14221), .dout(n14291));
  jnot g14100(.din(n14291), .dout(n14292));
  jxor g14101(.dina(n14292), .dinb(n14186), .dout(n14293));
  jnot g14102(.din(n14173), .dout(n14294));
  jor  g14103(.dina(n14182), .dinb(n14175), .dout(n14295));
  jand g14104(.dina(n14295), .dinb(n14294), .dout(n14296));
  jxor g14105(.dina(n14296), .dinb(n14293), .dout(\asquared[99] ));
  jand g14106(.dina(n14220), .dinb(n14189), .dout(n14298));
  jand g14107(.dina(n14290), .dinb(n14221), .dout(n14299));
  jor  g14108(.dina(n14299), .dinb(n14298), .dout(n14300));
  jand g14109(.dina(n14218), .dinb(n14195), .dout(n14301));
  jand g14110(.dina(n14219), .dinb(n14192), .dout(n14302));
  jor  g14111(.dina(n14302), .dinb(n14301), .dout(n14303));
  jand g14112(.dina(n14206), .dinb(n14203), .dout(n14304));
  jnot g14113(.din(n14304), .dout(n14305));
  jor  g14114(.dina(n14217), .dinb(n14208), .dout(n14306));
  jand g14115(.dina(n14306), .dinb(n14305), .dout(n14307));
  jnot g14116(.din(n14307), .dout(n14308));
  jand g14117(.dina(n14241), .dinb(n14238), .dout(n14309));
  jand g14118(.dina(n14245), .dinb(n14242), .dout(n14310));
  jor  g14119(.dina(n14310), .dinb(n14309), .dout(n14311));
  jand g14120(.dina(\a[62] ), .dinb(\a[37] ), .dout(n14312));
  jnot g14121(.din(n14312), .dout(n14313));
  jnot g14122(.din(\a[49] ), .dout(n14314));
  jand g14123(.dina(\a[50] ), .dinb(n14314), .dout(n14315));
  jxor g14124(.dina(n14315), .dinb(n14313), .dout(n14316));
  jnot g14125(.din(n14316), .dout(n14317));
  jxor g14126(.dina(n14317), .dinb(n14311), .dout(n14318));
  jxor g14127(.dina(n14318), .dinb(n14308), .dout(n14319));
  jand g14128(.dina(n14283), .dinb(n14277), .dout(n14320));
  jor  g14129(.dina(n14320), .dinb(n14281), .dout(n14321));
  jxor g14130(.dina(n14321), .dinb(n14271), .dout(n14322));
  jand g14131(.dina(n14202), .dinb(n14201), .dout(n14323));
  jor  g14132(.dina(n14323), .dinb(n14196), .dout(n14324));
  jxor g14133(.dina(n14324), .dinb(n14322), .dout(n14325));
  jnot g14134(.din(n14325), .dout(n14326));
  jor  g14135(.dina(n14285), .dinb(n14276), .dout(n14327));
  jand g14136(.dina(n14286), .dinb(n14261), .dout(n14328));
  jnot g14137(.din(n14328), .dout(n14329));
  jand g14138(.dina(n14329), .dinb(n14327), .dout(n14330));
  jxor g14139(.dina(n14330), .dinb(n14326), .dout(n14331));
  jand g14140(.dina(n14260), .dinb(n14258), .dout(n14332));
  jor  g14141(.dina(n14332), .dinb(n14253), .dout(n14333));
  jand g14142(.dina(n14213), .dinb(n14210), .dout(n14334));
  jnot g14143(.din(n14334), .dout(n14335));
  jand g14144(.dina(n14335), .dinb(n14215), .dout(n14336));
  jxor g14145(.dina(n14336), .dinb(n14333), .dout(n14337));
  jnot g14146(.din(n14337), .dout(n14338));
  jand g14147(.dina(\a[63] ), .dinb(\a[36] ), .dout(n14339));
  jand g14148(.dina(\a[61] ), .dinb(\a[39] ), .dout(n14340));
  jand g14149(.dina(n14340), .dinb(n14209), .dout(n14341));
  jand g14150(.dina(\a[61] ), .dinb(\a[38] ), .dout(n14342));
  jnot g14151(.din(n14342), .dout(n14343));
  jand g14152(.dina(\a[60] ), .dinb(\a[39] ), .dout(n14344));
  jnot g14153(.din(n14344), .dout(n14345));
  jand g14154(.dina(n14345), .dinb(n14343), .dout(n14346));
  jor  g14155(.dina(n14346), .dinb(n14341), .dout(n14347));
  jxor g14156(.dina(n14347), .dinb(n14339), .dout(n14348));
  jxor g14157(.dina(n14348), .dinb(n14338), .dout(n14349));
  jxor g14158(.dina(n14349), .dinb(n14331), .dout(n14350));
  jxor g14159(.dina(n14350), .dinb(n14319), .dout(n14351));
  jxor g14160(.dina(n14351), .dinb(n14303), .dout(n14352));
  jand g14161(.dina(n14288), .dinb(n14237), .dout(n14353));
  jand g14162(.dina(n14289), .dinb(n14224), .dout(n14354));
  jor  g14163(.dina(n14354), .dinb(n14353), .dout(n14355));
  jand g14164(.dina(n14230), .dinb(n14227), .dout(n14356));
  jnot g14165(.din(n14356), .dout(n14357));
  jor  g14166(.dina(n14236), .dinb(n14232), .dout(n14358));
  jand g14167(.dina(n14358), .dinb(n14357), .dout(n14359));
  jnot g14168(.din(n14359), .dout(n14360));
  jnot g14169(.din(n8067), .dout(n14361));
  jand g14170(.dina(\a[58] ), .dinb(\a[41] ), .dout(n14362));
  jnot g14171(.din(n14362), .dout(n14363));
  jand g14172(.dina(n14363), .dinb(n14361), .dout(n14364));
  jand g14173(.dina(n14362), .dinb(n8067), .dout(n14365));
  jnot g14174(.din(n14365), .dout(n14366));
  jand g14175(.dina(\a[59] ), .dinb(\a[41] ), .dout(n14367));
  jand g14176(.dina(n14367), .dinb(n14278), .dout(n14368));
  jand g14177(.dina(n14280), .dinb(n8067), .dout(n14369));
  jor  g14178(.dina(n14369), .dinb(n14368), .dout(n14370));
  jnot g14179(.din(n14370), .dout(n14371));
  jand g14180(.dina(n14371), .dinb(n14366), .dout(n14372));
  jnot g14181(.din(n14372), .dout(n14373));
  jor  g14182(.dina(n14373), .dinb(n14364), .dout(n14374));
  jand g14183(.dina(n14370), .dinb(n14366), .dout(n14375));
  jnot g14184(.din(n14375), .dout(n14376));
  jand g14185(.dina(n14376), .dinb(n14280), .dout(n14377));
  jnot g14186(.din(n14377), .dout(n14378));
  jand g14187(.dina(n14378), .dinb(n14374), .dout(n14379));
  jand g14188(.dina(\a[54] ), .dinb(\a[45] ), .dout(n14380));
  jnot g14189(.din(n14380), .dout(n14381));
  jand g14190(.dina(\a[53] ), .dinb(\a[47] ), .dout(n14382));
  jand g14191(.dina(n14382), .dinb(n14262), .dout(n14383));
  jnot g14192(.din(n14383), .dout(n14384));
  jand g14193(.dina(\a[53] ), .dinb(\a[46] ), .dout(n14385));
  jor  g14194(.dina(n14385), .dinb(n8013), .dout(n14386));
  jand g14195(.dina(n14386), .dinb(n14384), .dout(n14387));
  jxor g14196(.dina(n14387), .dinb(n14381), .dout(n14388));
  jxor g14197(.dina(n14388), .dinb(n14379), .dout(n14389));
  jnot g14198(.din(n14389), .dout(n14390));
  jand g14199(.dina(\a[51] ), .dinb(\a[48] ), .dout(n14391));
  jnot g14200(.din(n14391), .dout(n14392));
  jand g14201(.dina(\a[57] ), .dinb(\a[43] ), .dout(n14393));
  jand g14202(.dina(n14393), .dinb(n14139), .dout(n14394));
  jnot g14203(.din(n14394), .dout(n14395));
  jand g14204(.dina(\a[56] ), .dinb(\a[43] ), .dout(n14396));
  jor  g14205(.dina(n14396), .dinb(n14211), .dout(n14397));
  jand g14206(.dina(n14397), .dinb(n14395), .dout(n14398));
  jxor g14207(.dina(n14398), .dinb(n14392), .dout(n14399));
  jxor g14208(.dina(n14399), .dinb(n14390), .dout(n14400));
  jxor g14209(.dina(n14400), .dinb(n14360), .dout(n14401));
  jnot g14210(.din(n14401), .dout(n14402));
  jor  g14211(.dina(n14251), .dinb(n14247), .dout(n14403));
  jand g14212(.dina(n14287), .dinb(n14252), .dout(n14404));
  jnot g14213(.din(n14404), .dout(n14405));
  jand g14214(.dina(n14405), .dinb(n14403), .dout(n14406));
  jxor g14215(.dina(n14406), .dinb(n14402), .dout(n14407));
  jxor g14216(.dina(n14407), .dinb(n14355), .dout(n14408));
  jxor g14217(.dina(n14408), .dinb(n14352), .dout(n14409));
  jand g14218(.dina(n14409), .dinb(n14300), .dout(n14410));
  jor  g14219(.dina(n14409), .dinb(n14300), .dout(n14411));
  jnot g14220(.din(n14411), .dout(n14412));
  jor  g14221(.dina(n14412), .dinb(n14410), .dout(n14413));
  jand g14222(.dina(n14291), .dinb(n14186), .dout(n14414));
  jnot g14223(.din(n14414), .dout(n14415));
  jnot g14224(.din(n14186), .dout(n14416));
  jand g14225(.dina(n14292), .dinb(n14416), .dout(n14417));
  jor  g14226(.dina(n14296), .dinb(n14417), .dout(n14418));
  jand g14227(.dina(n14418), .dinb(n14415), .dout(n14419));
  jxor g14228(.dina(n14419), .dinb(n14413), .dout(\asquared[100] ));
  jand g14229(.dina(n14407), .dinb(n14355), .dout(n14421));
  jand g14230(.dina(n14408), .dinb(n14352), .dout(n14422));
  jor  g14231(.dina(n14422), .dinb(n14421), .dout(n14423));
  jand g14232(.dina(n14336), .dinb(n14333), .dout(n14424));
  jnot g14233(.din(n14424), .dout(n14425));
  jor  g14234(.dina(n14348), .dinb(n14338), .dout(n14426));
  jand g14235(.dina(n14426), .dinb(n14425), .dout(n14427));
  jnot g14236(.din(n14427), .dout(n14428));
  jand g14237(.dina(n14321), .dinb(n14271), .dout(n14429));
  jand g14238(.dina(n14324), .dinb(n14322), .dout(n14430));
  jor  g14239(.dina(n14430), .dinb(n14429), .dout(n14431));
  jnot g14240(.din(n14431), .dout(n14432));
  jnot g14241(.din(n14382), .dout(n14433));
  jand g14242(.dina(\a[52] ), .dinb(\a[49] ), .dout(n14434));
  jand g14243(.dina(n14434), .dinb(n14391), .dout(n14435));
  jnot g14244(.din(n14435), .dout(n14436));
  jand g14245(.dina(\a[51] ), .dinb(\a[49] ), .dout(n14437));
  jand g14246(.dina(\a[52] ), .dinb(\a[48] ), .dout(n14438));
  jor  g14247(.dina(n14438), .dinb(n14437), .dout(n14439));
  jand g14248(.dina(n14439), .dinb(n14436), .dout(n14440));
  jxor g14249(.dina(n14440), .dinb(n14433), .dout(n14441));
  jxor g14250(.dina(n14441), .dinb(n14432), .dout(n14442));
  jxor g14251(.dina(n14442), .dinb(n14428), .dout(n14443));
  jnot g14252(.din(n14443), .dout(n14444));
  jand g14253(.dina(n14400), .dinb(n14360), .dout(n14445));
  jnot g14254(.din(n14445), .dout(n14446));
  jor  g14255(.dina(n14406), .dinb(n14402), .dout(n14447));
  jand g14256(.dina(n14447), .dinb(n14446), .dout(n14448));
  jxor g14257(.dina(n14448), .dinb(n14444), .dout(n14449));
  jnot g14258(.din(n14339), .dout(n14450));
  jnot g14259(.din(n14341), .dout(n14451));
  jand g14260(.dina(n14451), .dinb(n14450), .dout(n14452));
  jor  g14261(.dina(n14452), .dinb(n14346), .dout(n14453));
  jnot g14262(.din(n14453), .dout(n14454));
  jand g14263(.dina(n14384), .dinb(n14381), .dout(n14455));
  jnot g14264(.din(n14455), .dout(n14456));
  jand g14265(.dina(n14456), .dinb(n14386), .dout(n14457));
  jxor g14266(.dina(n14457), .dinb(n14454), .dout(n14458));
  jxor g14267(.dina(n14458), .dinb(n14373), .dout(n14459));
  jnot g14268(.din(n14459), .dout(n14460));
  jor  g14269(.dina(n14388), .dinb(n14379), .dout(n14461));
  jor  g14270(.dina(n14399), .dinb(n14390), .dout(n14462));
  jand g14271(.dina(n14462), .dinb(n14461), .dout(n14463));
  jxor g14272(.dina(n14463), .dinb(n14460), .dout(n14464));
  jand g14273(.dina(\a[63] ), .dinb(\a[37] ), .dout(n14465));
  jnot g14274(.din(\a[50] ), .dout(n14466));
  jand g14275(.dina(n14313), .dinb(n14314), .dout(n14467));
  jor  g14276(.dina(n14467), .dinb(n14466), .dout(n14468));
  jnot g14277(.din(n14468), .dout(n14469));
  jxor g14278(.dina(n14469), .dinb(n14465), .dout(n14470));
  jand g14279(.dina(n14395), .dinb(n14392), .dout(n14471));
  jnot g14280(.din(n14471), .dout(n14472));
  jand g14281(.dina(n14472), .dinb(n14397), .dout(n14473));
  jxor g14282(.dina(n14473), .dinb(n14470), .dout(n14474));
  jxor g14283(.dina(n14474), .dinb(n14464), .dout(n14475));
  jxor g14284(.dina(n14475), .dinb(n14449), .dout(n14476));
  jand g14285(.dina(n14350), .dinb(n14319), .dout(n14477));
  jand g14286(.dina(n14351), .dinb(n14303), .dout(n14478));
  jor  g14287(.dina(n14478), .dinb(n14477), .dout(n14479));
  jand g14288(.dina(n14317), .dinb(n14311), .dout(n14480));
  jand g14289(.dina(n14318), .dinb(n14308), .dout(n14481));
  jor  g14290(.dina(n14481), .dinb(n14480), .dout(n14482));
  jand g14291(.dina(\a[61] ), .dinb(\a[40] ), .dout(n14483));
  jand g14292(.dina(n14483), .dinb(n14344), .dout(n14484));
  jnot g14293(.din(n14484), .dout(n14485));
  jand g14294(.dina(\a[60] ), .dinb(\a[40] ), .dout(n14486));
  jand g14295(.dina(\a[62] ), .dinb(\a[38] ), .dout(n14487));
  jand g14296(.dina(n14487), .dinb(n14486), .dout(n14488));
  jand g14297(.dina(\a[62] ), .dinb(\a[39] ), .dout(n14489));
  jand g14298(.dina(n14489), .dinb(n14342), .dout(n14490));
  jor  g14299(.dina(n14490), .dinb(n14488), .dout(n14491));
  jnot g14300(.din(n14491), .dout(n14492));
  jand g14301(.dina(n14492), .dinb(n14485), .dout(n14493));
  jor  g14302(.dina(n14486), .dinb(n14340), .dout(n14494));
  jand g14303(.dina(n14494), .dinb(n14493), .dout(n14495));
  jand g14304(.dina(n14491), .dinb(n14485), .dout(n14496));
  jnot g14305(.din(n14496), .dout(n14497));
  jand g14306(.dina(n14497), .dinb(n14487), .dout(n14498));
  jor  g14307(.dina(n14498), .dinb(n14495), .dout(n14499));
  jnot g14308(.din(n14393), .dout(n14500));
  jand g14309(.dina(\a[56] ), .dinb(\a[45] ), .dout(n14501));
  jand g14310(.dina(n14501), .dinb(n8067), .dout(n14502));
  jnot g14311(.din(n14502), .dout(n14503));
  jand g14312(.dina(\a[55] ), .dinb(\a[45] ), .dout(n14504));
  jand g14313(.dina(\a[56] ), .dinb(\a[44] ), .dout(n14505));
  jor  g14314(.dina(n14505), .dinb(n14504), .dout(n14506));
  jand g14315(.dina(n14506), .dinb(n14503), .dout(n14507));
  jxor g14316(.dina(n14507), .dinb(n14500), .dout(n14508));
  jnot g14317(.din(n14508), .dout(n14509));
  jxor g14318(.dina(n14509), .dinb(n14499), .dout(n14510));
  jnot g14319(.din(n14510), .dout(n14511));
  jnot g14320(.din(n7992), .dout(n14512));
  jand g14321(.dina(\a[59] ), .dinb(\a[42] ), .dout(n14513));
  jand g14322(.dina(n14513), .dinb(n14362), .dout(n14514));
  jnot g14323(.din(n14514), .dout(n14515));
  jand g14324(.dina(\a[58] ), .dinb(\a[42] ), .dout(n14516));
  jor  g14325(.dina(n14516), .dinb(n14367), .dout(n14517));
  jand g14326(.dina(n14517), .dinb(n14515), .dout(n14518));
  jxor g14327(.dina(n14518), .dinb(n14512), .dout(n14519));
  jxor g14328(.dina(n14519), .dinb(n14511), .dout(n14520));
  jxor g14329(.dina(n14520), .dinb(n14482), .dout(n14521));
  jnot g14330(.din(n14521), .dout(n14522));
  jor  g14331(.dina(n14330), .dinb(n14326), .dout(n14523));
  jand g14332(.dina(n14349), .dinb(n14331), .dout(n14524));
  jnot g14333(.din(n14524), .dout(n14525));
  jand g14334(.dina(n14525), .dinb(n14523), .dout(n14526));
  jxor g14335(.dina(n14526), .dinb(n14522), .dout(n14527));
  jxor g14336(.dina(n14527), .dinb(n14479), .dout(n14528));
  jxor g14337(.dina(n14528), .dinb(n14476), .dout(n14529));
  jand g14338(.dina(n14529), .dinb(n14423), .dout(n14530));
  jor  g14339(.dina(n14529), .dinb(n14423), .dout(n14531));
  jnot g14340(.din(n14531), .dout(n14532));
  jor  g14341(.dina(n14532), .dinb(n14530), .dout(n14533));
  jnot g14342(.din(n14410), .dout(n14534));
  jor  g14343(.dina(n14419), .dinb(n14412), .dout(n14535));
  jand g14344(.dina(n14535), .dinb(n14534), .dout(n14536));
  jxor g14345(.dina(n14536), .dinb(n14533), .dout(\asquared[101] ));
  jand g14346(.dina(n14527), .dinb(n14479), .dout(n14538));
  jand g14347(.dina(n14528), .dinb(n14476), .dout(n14539));
  jor  g14348(.dina(n14539), .dinb(n14538), .dout(n14540));
  jor  g14349(.dina(n14448), .dinb(n14444), .dout(n14541));
  jand g14350(.dina(n14475), .dinb(n14449), .dout(n14542));
  jnot g14351(.din(n14542), .dout(n14543));
  jand g14352(.dina(n14543), .dinb(n14541), .dout(n14544));
  jnot g14353(.din(n14544), .dout(n14545));
  jor  g14354(.dina(n14441), .dinb(n14432), .dout(n14546));
  jand g14355(.dina(n14442), .dinb(n14428), .dout(n14547));
  jnot g14356(.din(n14547), .dout(n14548));
  jand g14357(.dina(n14548), .dinb(n14546), .dout(n14549));
  jnot g14358(.din(n14549), .dout(n14550));
  jand g14359(.dina(\a[53] ), .dinb(\a[48] ), .dout(n14551));
  jand g14360(.dina(\a[57] ), .dinb(\a[44] ), .dout(n14552));
  jand g14361(.dina(n14552), .dinb(n14434), .dout(n14553));
  jnot g14362(.din(n14553), .dout(n14554));
  jand g14363(.dina(n7729), .dinb(n7165), .dout(n14555));
  jand g14364(.dina(n14552), .dinb(n14551), .dout(n14556));
  jor  g14365(.dina(n14556), .dinb(n14555), .dout(n14557));
  jand g14366(.dina(n14557), .dinb(n14554), .dout(n14558));
  jnot g14367(.din(n14558), .dout(n14559));
  jand g14368(.dina(n14559), .dinb(n14551), .dout(n14560));
  jor  g14369(.dina(n14557), .dinb(n14553), .dout(n14561));
  jnot g14370(.din(n14561), .dout(n14562));
  jor  g14371(.dina(n14552), .dinb(n14434), .dout(n14563));
  jand g14372(.dina(n14563), .dinb(n14562), .dout(n14564));
  jor  g14373(.dina(n14564), .dinb(n14560), .dout(n14565));
  jand g14374(.dina(\a[63] ), .dinb(\a[38] ), .dout(n14566));
  jand g14375(.dina(\a[54] ), .dinb(\a[47] ), .dout(n14567));
  jand g14376(.dina(\a[55] ), .dinb(\a[46] ), .dout(n14568));
  jor  g14377(.dina(n14568), .dinb(n14567), .dout(n14569));
  jand g14378(.dina(\a[55] ), .dinb(\a[47] ), .dout(n14570));
  jand g14379(.dina(n14570), .dinb(n7992), .dout(n14571));
  jnot g14380(.din(n14571), .dout(n14572));
  jand g14381(.dina(n14572), .dinb(n14569), .dout(n14573));
  jxor g14382(.dina(n14573), .dinb(n14566), .dout(n14574));
  jnot g14383(.din(n14574), .dout(n14575));
  jnot g14384(.din(n14513), .dout(n14576));
  jand g14385(.dina(n12907), .dinb(n11688), .dout(n14577));
  jnot g14386(.din(n14577), .dout(n14578));
  jand g14387(.dina(\a[58] ), .dinb(\a[43] ), .dout(n14579));
  jor  g14388(.dina(n14579), .dinb(n14501), .dout(n14580));
  jand g14389(.dina(n14580), .dinb(n14578), .dout(n14581));
  jxor g14390(.dina(n14581), .dinb(n14576), .dout(n14582));
  jxor g14391(.dina(n14582), .dinb(n14575), .dout(n14583));
  jxor g14392(.dina(n14583), .dinb(n14565), .dout(n14584));
  jxor g14393(.dina(n14584), .dinb(n14550), .dout(n14585));
  jand g14394(.dina(n14469), .dinb(n14465), .dout(n14586));
  jand g14395(.dina(n14473), .dinb(n14470), .dout(n14587));
  jor  g14396(.dina(n14587), .dinb(n14586), .dout(n14588));
  jand g14397(.dina(\a[61] ), .dinb(\a[41] ), .dout(n14589));
  jand g14398(.dina(n14589), .dinb(n14486), .dout(n14590));
  jnot g14399(.din(n14590), .dout(n14591));
  jand g14400(.dina(\a[60] ), .dinb(\a[41] ), .dout(n14592));
  jor  g14401(.dina(n14592), .dinb(n14483), .dout(n14593));
  jand g14402(.dina(n14593), .dinb(n14591), .dout(n14594));
  jand g14403(.dina(n14436), .dinb(n14433), .dout(n14595));
  jnot g14404(.din(n14595), .dout(n14596));
  jand g14405(.dina(n14596), .dinb(n14439), .dout(n14597));
  jxor g14406(.dina(n14597), .dinb(n14594), .dout(n14598));
  jand g14407(.dina(\a[51] ), .dinb(n14466), .dout(n14599));
  jxor g14408(.dina(n14599), .dinb(n14489), .dout(n14600));
  jxor g14409(.dina(n14600), .dinb(n14598), .dout(n14601));
  jxor g14410(.dina(n14601), .dinb(n14588), .dout(n14602));
  jxor g14411(.dina(n14602), .dinb(n14585), .dout(n14603));
  jxor g14412(.dina(n14603), .dinb(n14545), .dout(n14604));
  jnot g14413(.din(n14493), .dout(n14605));
  jand g14414(.dina(n14515), .dinb(n14512), .dout(n14606));
  jnot g14415(.din(n14606), .dout(n14607));
  jand g14416(.dina(n14607), .dinb(n14517), .dout(n14608));
  jxor g14417(.dina(n14608), .dinb(n14605), .dout(n14609));
  jand g14418(.dina(n14503), .dinb(n14500), .dout(n14610));
  jnot g14419(.din(n14610), .dout(n14611));
  jand g14420(.dina(n14611), .dinb(n14506), .dout(n14612));
  jxor g14421(.dina(n14612), .dinb(n14609), .dout(n14613));
  jand g14422(.dina(n14509), .dinb(n14499), .dout(n14614));
  jnot g14423(.din(n14614), .dout(n14615));
  jor  g14424(.dina(n14519), .dinb(n14511), .dout(n14616));
  jand g14425(.dina(n14616), .dinb(n14615), .dout(n14617));
  jnot g14426(.din(n14617), .dout(n14618));
  jand g14427(.dina(n14457), .dinb(n14454), .dout(n14619));
  jand g14428(.dina(n14458), .dinb(n14373), .dout(n14620));
  jor  g14429(.dina(n14620), .dinb(n14619), .dout(n14621));
  jxor g14430(.dina(n14621), .dinb(n14618), .dout(n14622));
  jxor g14431(.dina(n14622), .dinb(n14613), .dout(n14623));
  jand g14432(.dina(n14520), .dinb(n14482), .dout(n14624));
  jnot g14433(.din(n14624), .dout(n14625));
  jor  g14434(.dina(n14526), .dinb(n14522), .dout(n14626));
  jand g14435(.dina(n14626), .dinb(n14625), .dout(n14627));
  jor  g14436(.dina(n14463), .dinb(n14460), .dout(n14628));
  jand g14437(.dina(n14474), .dinb(n14464), .dout(n14629));
  jnot g14438(.din(n14629), .dout(n14630));
  jand g14439(.dina(n14630), .dinb(n14628), .dout(n14631));
  jxor g14440(.dina(n14631), .dinb(n14627), .dout(n14632));
  jxor g14441(.dina(n14632), .dinb(n14623), .dout(n14633));
  jxor g14442(.dina(n14633), .dinb(n14604), .dout(n14634));
  jand g14443(.dina(n14634), .dinb(n14540), .dout(n14635));
  jor  g14444(.dina(n14634), .dinb(n14540), .dout(n14636));
  jnot g14445(.din(n14636), .dout(n14637));
  jor  g14446(.dina(n14637), .dinb(n14635), .dout(n14638));
  jnot g14447(.din(n14530), .dout(n14639));
  jor  g14448(.dina(n14536), .dinb(n14532), .dout(n14640));
  jand g14449(.dina(n14640), .dinb(n14639), .dout(n14641));
  jxor g14450(.dina(n14641), .dinb(n14638), .dout(\asquared[102] ));
  jand g14451(.dina(n14603), .dinb(n14545), .dout(n14643));
  jand g14452(.dina(n14633), .dinb(n14604), .dout(n14644));
  jor  g14453(.dina(n14644), .dinb(n14643), .dout(n14645));
  jor  g14454(.dina(n14631), .dinb(n14627), .dout(n14646));
  jand g14455(.dina(n14632), .dinb(n14623), .dout(n14647));
  jnot g14456(.din(n14647), .dout(n14648));
  jand g14457(.dina(n14648), .dinb(n14646), .dout(n14649));
  jnot g14458(.din(n14649), .dout(n14650));
  jand g14459(.dina(n14600), .dinb(n14598), .dout(n14651));
  jand g14460(.dina(n14601), .dinb(n14588), .dout(n14652));
  jor  g14461(.dina(n14652), .dinb(n14651), .dout(n14653));
  jand g14462(.dina(n14597), .dinb(n14594), .dout(n14654));
  jor  g14463(.dina(n14654), .dinb(n14590), .dout(n14655));
  jand g14464(.dina(n14578), .dinb(n14576), .dout(n14656));
  jnot g14465(.din(n14656), .dout(n14657));
  jand g14466(.dina(n14657), .dinb(n14580), .dout(n14658));
  jxor g14467(.dina(n14658), .dinb(n14655), .dout(n14659));
  jnot g14468(.din(n14659), .dout(n14660));
  jand g14469(.dina(\a[63] ), .dinb(\a[39] ), .dout(n14661));
  jnot g14470(.din(n14661), .dout(n14662));
  jand g14471(.dina(\a[61] ), .dinb(\a[42] ), .dout(n14663));
  jand g14472(.dina(n14663), .dinb(n14592), .dout(n14664));
  jnot g14473(.din(n14664), .dout(n14665));
  jand g14474(.dina(\a[60] ), .dinb(\a[42] ), .dout(n14666));
  jor  g14475(.dina(n14666), .dinb(n14589), .dout(n14667));
  jand g14476(.dina(n14667), .dinb(n14665), .dout(n14668));
  jxor g14477(.dina(n14668), .dinb(n14662), .dout(n14669));
  jxor g14478(.dina(n14669), .dinb(n14660), .dout(n14670));
  jxor g14479(.dina(n14670), .dinb(n14653), .dout(n14671));
  jand g14480(.dina(\a[62] ), .dinb(\a[40] ), .dout(n14672));
  jand g14481(.dina(\a[59] ), .dinb(\a[43] ), .dout(n14673));
  jand g14482(.dina(\a[58] ), .dinb(\a[44] ), .dout(n14674));
  jor  g14483(.dina(n14674), .dinb(n14673), .dout(n14675));
  jand g14484(.dina(\a[59] ), .dinb(\a[44] ), .dout(n14676));
  jand g14485(.dina(n14676), .dinb(n14579), .dout(n14677));
  jnot g14486(.din(n14677), .dout(n14678));
  jand g14487(.dina(n14678), .dinb(n14675), .dout(n14679));
  jxor g14488(.dina(n14679), .dinb(n14672), .dout(n14680));
  jnot g14489(.din(n14680), .dout(n14681));
  jand g14490(.dina(\a[57] ), .dinb(\a[45] ), .dout(n14682));
  jnot g14491(.din(n14682), .dout(n14683));
  jand g14492(.dina(\a[56] ), .dinb(\a[47] ), .dout(n14684));
  jand g14493(.dina(n14684), .dinb(n14568), .dout(n14685));
  jnot g14494(.din(n14685), .dout(n14686));
  jand g14495(.dina(\a[56] ), .dinb(\a[46] ), .dout(n14687));
  jor  g14496(.dina(n14687), .dinb(n14570), .dout(n14688));
  jand g14497(.dina(n14688), .dinb(n14686), .dout(n14689));
  jxor g14498(.dina(n14689), .dinb(n14683), .dout(n14690));
  jxor g14499(.dina(n14690), .dinb(n14681), .dout(n14691));
  jnot g14500(.din(n14691), .dout(n14692));
  jand g14501(.dina(\a[54] ), .dinb(\a[48] ), .dout(n14693));
  jnot g14502(.din(n14693), .dout(n14694));
  jand g14503(.dina(\a[53] ), .dinb(\a[50] ), .dout(n14695));
  jand g14504(.dina(n14695), .dinb(n14434), .dout(n14696));
  jnot g14505(.din(n14696), .dout(n14697));
  jand g14506(.dina(\a[53] ), .dinb(\a[49] ), .dout(n14698));
  jand g14507(.dina(\a[52] ), .dinb(\a[50] ), .dout(n14699));
  jor  g14508(.dina(n14699), .dinb(n14698), .dout(n14700));
  jand g14509(.dina(n14700), .dinb(n14697), .dout(n14701));
  jxor g14510(.dina(n14701), .dinb(n14694), .dout(n14702));
  jxor g14511(.dina(n14702), .dinb(n14692), .dout(n14703));
  jxor g14512(.dina(n14703), .dinb(n14671), .dout(n14704));
  jxor g14513(.dina(n14704), .dinb(n14650), .dout(n14705));
  jand g14514(.dina(n14573), .dinb(n14566), .dout(n14706));
  jor  g14515(.dina(n14706), .dinb(n14571), .dout(n14707));
  jor  g14516(.dina(n14489), .dinb(\a[50] ), .dout(n14708));
  jand g14517(.dina(n14708), .dinb(\a[51] ), .dout(n14709));
  jxor g14518(.dina(n14709), .dinb(n14561), .dout(n14710));
  jxor g14519(.dina(n14710), .dinb(n14707), .dout(n14711));
  jand g14520(.dina(n14608), .dinb(n14605), .dout(n14712));
  jand g14521(.dina(n14612), .dinb(n14609), .dout(n14713));
  jor  g14522(.dina(n14713), .dinb(n14712), .dout(n14714));
  jxor g14523(.dina(n14714), .dinb(n14711), .dout(n14715));
  jnot g14524(.din(n14715), .dout(n14716));
  jor  g14525(.dina(n14582), .dinb(n14575), .dout(n14717));
  jand g14526(.dina(n14583), .dinb(n14565), .dout(n14718));
  jnot g14527(.din(n14718), .dout(n14719));
  jand g14528(.dina(n14719), .dinb(n14717), .dout(n14720));
  jxor g14529(.dina(n14720), .dinb(n14716), .dout(n14721));
  jand g14530(.dina(n14584), .dinb(n14550), .dout(n14722));
  jand g14531(.dina(n14602), .dinb(n14585), .dout(n14723));
  jor  g14532(.dina(n14723), .dinb(n14722), .dout(n14724));
  jand g14533(.dina(n14621), .dinb(n14618), .dout(n14725));
  jand g14534(.dina(n14622), .dinb(n14613), .dout(n14726));
  jor  g14535(.dina(n14726), .dinb(n14725), .dout(n14727));
  jxor g14536(.dina(n14727), .dinb(n14724), .dout(n14728));
  jxor g14537(.dina(n14728), .dinb(n14721), .dout(n14729));
  jxor g14538(.dina(n14729), .dinb(n14705), .dout(n14730));
  jnot g14539(.din(n14730), .dout(n14731));
  jxor g14540(.dina(n14731), .dinb(n14645), .dout(n14732));
  jnot g14541(.din(n14635), .dout(n14733));
  jor  g14542(.dina(n14641), .dinb(n14637), .dout(n14734));
  jand g14543(.dina(n14734), .dinb(n14733), .dout(n14735));
  jxor g14544(.dina(n14735), .dinb(n14732), .dout(\asquared[103] ));
  jand g14545(.dina(n14704), .dinb(n14650), .dout(n14737));
  jand g14546(.dina(n14729), .dinb(n14705), .dout(n14738));
  jor  g14547(.dina(n14738), .dinb(n14737), .dout(n14739));
  jand g14548(.dina(n14658), .dinb(n14655), .dout(n14740));
  jnot g14549(.din(n14740), .dout(n14741));
  jor  g14550(.dina(n14669), .dinb(n14660), .dout(n14742));
  jand g14551(.dina(n14742), .dinb(n14741), .dout(n14743));
  jnot g14552(.din(n14743), .dout(n14744));
  jand g14553(.dina(n14709), .dinb(n14561), .dout(n14745));
  jand g14554(.dina(n14710), .dinb(n14707), .dout(n14746));
  jor  g14555(.dina(n14746), .dinb(n14745), .dout(n14747));
  jxor g14556(.dina(n14747), .dinb(n14744), .dout(n14748));
  jnot g14557(.din(n14748), .dout(n14749));
  jor  g14558(.dina(n14690), .dinb(n14681), .dout(n14750));
  jor  g14559(.dina(n14702), .dinb(n14692), .dout(n14751));
  jand g14560(.dina(n14751), .dinb(n14750), .dout(n14752));
  jxor g14561(.dina(n14752), .dinb(n14749), .dout(n14753));
  jand g14562(.dina(n14670), .dinb(n14653), .dout(n14754));
  jand g14563(.dina(n14703), .dinb(n14671), .dout(n14755));
  jor  g14564(.dina(n14755), .dinb(n14754), .dout(n14756));
  jnot g14565(.din(n14756), .dout(n14757));
  jand g14566(.dina(n14714), .dinb(n14711), .dout(n14758));
  jnot g14567(.din(n14758), .dout(n14759));
  jor  g14568(.dina(n14720), .dinb(n14716), .dout(n14760));
  jand g14569(.dina(n14760), .dinb(n14759), .dout(n14761));
  jxor g14570(.dina(n14761), .dinb(n14757), .dout(n14762));
  jxor g14571(.dina(n14762), .dinb(n14753), .dout(n14763));
  jand g14572(.dina(n14727), .dinb(n14724), .dout(n14764));
  jand g14573(.dina(n14728), .dinb(n14721), .dout(n14765));
  jor  g14574(.dina(n14765), .dinb(n14764), .dout(n14766));
  jand g14575(.dina(\a[63] ), .dinb(\a[40] ), .dout(n14767));
  jand g14576(.dina(n14697), .dinb(n14694), .dout(n14768));
  jnot g14577(.din(n14768), .dout(n14769));
  jand g14578(.dina(n14769), .dinb(n14700), .dout(n14770));
  jxor g14579(.dina(n14770), .dinb(n14767), .dout(n14771));
  jand g14580(.dina(n14686), .dinb(n14683), .dout(n14772));
  jnot g14581(.din(n14772), .dout(n14773));
  jand g14582(.dina(n14773), .dinb(n14688), .dout(n14774));
  jxor g14583(.dina(n14774), .dinb(n14771), .dout(n14775));
  jand g14584(.dina(n14679), .dinb(n14672), .dout(n14776));
  jor  g14585(.dina(n14776), .dinb(n14677), .dout(n14777));
  jand g14586(.dina(n14665), .dinb(n14662), .dout(n14778));
  jnot g14587(.din(n14778), .dout(n14779));
  jand g14588(.dina(n14779), .dinb(n14667), .dout(n14780));
  jxor g14589(.dina(n14780), .dinb(n14777), .dout(n14781));
  jand g14590(.dina(\a[59] ), .dinb(\a[45] ), .dout(n14782));
  jand g14591(.dina(n14782), .dinb(n14674), .dout(n14783));
  jnot g14592(.din(n14783), .dout(n14784));
  jand g14593(.dina(n13790), .dinb(n6097), .dout(n14785));
  jand g14594(.dina(\a[58] ), .dinb(\a[45] ), .dout(n14786));
  jand g14595(.dina(n14786), .dinb(n14663), .dout(n14787));
  jor  g14596(.dina(n14787), .dinb(n14785), .dout(n14788));
  jand g14597(.dina(n14788), .dinb(n14784), .dout(n14789));
  jnot g14598(.din(n14789), .dout(n14790));
  jand g14599(.dina(n14790), .dinb(n14663), .dout(n14791));
  jor  g14600(.dina(n14786), .dinb(n14676), .dout(n14792));
  jor  g14601(.dina(n14788), .dinb(n14783), .dout(n14793));
  jnot g14602(.din(n14793), .dout(n14794));
  jand g14603(.dina(n14794), .dinb(n14792), .dout(n14795));
  jor  g14604(.dina(n14795), .dinb(n14791), .dout(n14796));
  jxor g14605(.dina(n14796), .dinb(n14781), .dout(n14797));
  jxor g14606(.dina(n14797), .dinb(n14775), .dout(n14798));
  jand g14607(.dina(\a[60] ), .dinb(\a[43] ), .dout(n14799));
  jnot g14608(.din(n14684), .dout(n14800));
  jand g14609(.dina(\a[57] ), .dinb(\a[46] ), .dout(n14801));
  jnot g14610(.din(n14801), .dout(n14802));
  jand g14611(.dina(n14802), .dinb(n14800), .dout(n14803));
  jand g14612(.dina(\a[57] ), .dinb(\a[47] ), .dout(n14804));
  jand g14613(.dina(n14804), .dinb(n14687), .dout(n14805));
  jor  g14614(.dina(n14805), .dinb(n14803), .dout(n14806));
  jnot g14615(.din(n14806), .dout(n14807));
  jxor g14616(.dina(n14807), .dinb(n14799), .dout(n14808));
  jnot g14617(.din(n14808), .dout(n14809));
  jand g14618(.dina(\a[55] ), .dinb(\a[48] ), .dout(n14810));
  jnot g14619(.din(n14810), .dout(n14811));
  jand g14620(.dina(\a[54] ), .dinb(\a[50] ), .dout(n14812));
  jand g14621(.dina(n14812), .dinb(n14698), .dout(n14813));
  jnot g14622(.din(n14813), .dout(n14814));
  jor  g14623(.dina(n14695), .dinb(n10245), .dout(n14815));
  jand g14624(.dina(n14815), .dinb(n14814), .dout(n14816));
  jxor g14625(.dina(n14816), .dinb(n14811), .dout(n14817));
  jxor g14626(.dina(n14817), .dinb(n14809), .dout(n14818));
  jnot g14627(.din(n14818), .dout(n14819));
  jand g14628(.dina(\a[62] ), .dinb(\a[41] ), .dout(n14820));
  jnot g14629(.din(n14820), .dout(n14821));
  jnot g14630(.din(\a[51] ), .dout(n14822));
  jand g14631(.dina(\a[52] ), .dinb(n14822), .dout(n14823));
  jxor g14632(.dina(n14823), .dinb(n14821), .dout(n14824));
  jxor g14633(.dina(n14824), .dinb(n14819), .dout(n14825));
  jxor g14634(.dina(n14825), .dinb(n14798), .dout(n14826));
  jxor g14635(.dina(n14826), .dinb(n14766), .dout(n14827));
  jxor g14636(.dina(n14827), .dinb(n14763), .dout(n14828));
  jand g14637(.dina(n14828), .dinb(n14739), .dout(n14829));
  jor  g14638(.dina(n14828), .dinb(n14739), .dout(n14830));
  jnot g14639(.din(n14830), .dout(n14831));
  jor  g14640(.dina(n14831), .dinb(n14829), .dout(n14832));
  jand g14641(.dina(n14730), .dinb(n14645), .dout(n14833));
  jnot g14642(.din(n14833), .dout(n14834));
  jnot g14643(.din(n14645), .dout(n14835));
  jand g14644(.dina(n14731), .dinb(n14835), .dout(n14836));
  jor  g14645(.dina(n14735), .dinb(n14836), .dout(n14837));
  jand g14646(.dina(n14837), .dinb(n14834), .dout(n14838));
  jxor g14647(.dina(n14838), .dinb(n14832), .dout(\asquared[104] ));
  jand g14648(.dina(n14826), .dinb(n14766), .dout(n14840));
  jand g14649(.dina(n14827), .dinb(n14763), .dout(n14841));
  jor  g14650(.dina(n14841), .dinb(n14840), .dout(n14842));
  jand g14651(.dina(n14797), .dinb(n14775), .dout(n14843));
  jand g14652(.dina(n14825), .dinb(n14798), .dout(n14844));
  jor  g14653(.dina(n14844), .dinb(n14843), .dout(n14845));
  jnot g14654(.din(n14845), .dout(n14846));
  jand g14655(.dina(n14747), .dinb(n14744), .dout(n14847));
  jnot g14656(.din(n14847), .dout(n14848));
  jor  g14657(.dina(n14752), .dinb(n14749), .dout(n14849));
  jand g14658(.dina(n14849), .dinb(n14848), .dout(n14850));
  jxor g14659(.dina(n14850), .dinb(n14846), .dout(n14851));
  jand g14660(.dina(n14770), .dinb(n14767), .dout(n14852));
  jand g14661(.dina(n14774), .dinb(n14771), .dout(n14853));
  jor  g14662(.dina(n14853), .dinb(n14852), .dout(n14854));
  jand g14663(.dina(\a[63] ), .dinb(\a[42] ), .dout(n14855));
  jand g14664(.dina(n14855), .dinb(n14820), .dout(n14856));
  jnot g14665(.din(n14856), .dout(n14857));
  jand g14666(.dina(\a[62] ), .dinb(\a[42] ), .dout(n14858));
  jand g14667(.dina(\a[63] ), .dinb(\a[41] ), .dout(n14859));
  jor  g14668(.dina(n14859), .dinb(n14858), .dout(n14860));
  jand g14669(.dina(n14860), .dinb(n14857), .dout(n14861));
  jnot g14670(.din(\a[52] ), .dout(n14862));
  jand g14671(.dina(n14821), .dinb(n14822), .dout(n14863));
  jor  g14672(.dina(n14863), .dinb(n14862), .dout(n14864));
  jnot g14673(.din(n14864), .dout(n14865));
  jxor g14674(.dina(n14865), .dinb(n14861), .dout(n14866));
  jxor g14675(.dina(n14866), .dinb(n14854), .dout(n14867));
  jand g14676(.dina(n14780), .dinb(n14777), .dout(n14868));
  jand g14677(.dina(n14796), .dinb(n14781), .dout(n14869));
  jor  g14678(.dina(n14869), .dinb(n14868), .dout(n14870));
  jxor g14679(.dina(n14870), .dinb(n14867), .dout(n14871));
  jxor g14680(.dina(n14871), .dinb(n14851), .dout(n14872));
  jor  g14681(.dina(n14761), .dinb(n14757), .dout(n14873));
  jand g14682(.dina(n14762), .dinb(n14753), .dout(n14874));
  jnot g14683(.din(n14874), .dout(n14875));
  jand g14684(.dina(n14875), .dinb(n14873), .dout(n14876));
  jnot g14685(.din(n14876), .dout(n14877));
  jand g14686(.dina(n14807), .dinb(n14799), .dout(n14878));
  jor  g14687(.dina(n14878), .dinb(n14805), .dout(n14879));
  jand g14688(.dina(n14814), .dinb(n14811), .dout(n14880));
  jnot g14689(.din(n14880), .dout(n14881));
  jand g14690(.dina(n14881), .dinb(n14815), .dout(n14882));
  jxor g14691(.dina(n14882), .dinb(n14879), .dout(n14883));
  jxor g14692(.dina(n14883), .dinb(n14793), .dout(n14884));
  jnot g14693(.din(n14884), .dout(n14885));
  jor  g14694(.dina(n14817), .dinb(n14809), .dout(n14886));
  jor  g14695(.dina(n14824), .dinb(n14819), .dout(n14887));
  jand g14696(.dina(n14887), .dinb(n14886), .dout(n14888));
  jxor g14697(.dina(n14888), .dinb(n14885), .dout(n14889));
  jand g14698(.dina(\a[55] ), .dinb(\a[49] ), .dout(n14890));
  jand g14699(.dina(n7559), .dinb(n5594), .dout(n14891));
  jnot g14700(.din(n14891), .dout(n14892));
  jand g14701(.dina(n14890), .dinb(n6130), .dout(n14893));
  jand g14702(.dina(\a[55] ), .dinb(\a[50] ), .dout(n14894));
  jand g14703(.dina(n14894), .dinb(n10245), .dout(n14895));
  jor  g14704(.dina(n14895), .dinb(n14893), .dout(n14896));
  jand g14705(.dina(n14896), .dinb(n14892), .dout(n14897));
  jnot g14706(.din(n14897), .dout(n14898));
  jand g14707(.dina(n14898), .dinb(n14890), .dout(n14899));
  jor  g14708(.dina(n14896), .dinb(n14891), .dout(n14900));
  jnot g14709(.din(n14900), .dout(n14901));
  jor  g14710(.dina(n14812), .dinb(n6130), .dout(n14902));
  jand g14711(.dina(n14902), .dinb(n14901), .dout(n14903));
  jor  g14712(.dina(n14903), .dinb(n14899), .dout(n14904));
  jand g14713(.dina(\a[58] ), .dinb(\a[46] ), .dout(n14905));
  jand g14714(.dina(\a[57] ), .dinb(\a[48] ), .dout(n14906));
  jand g14715(.dina(n14906), .dinb(n14684), .dout(n14907));
  jnot g14716(.din(n14907), .dout(n14908));
  jand g14717(.dina(\a[58] ), .dinb(\a[47] ), .dout(n14909));
  jand g14718(.dina(n14909), .dinb(n14801), .dout(n14910));
  jand g14719(.dina(n14905), .dinb(n8215), .dout(n14911));
  jor  g14720(.dina(n14911), .dinb(n14910), .dout(n14912));
  jand g14721(.dina(n14912), .dinb(n14908), .dout(n14913));
  jnot g14722(.din(n14913), .dout(n14914));
  jand g14723(.dina(n14914), .dinb(n14905), .dout(n14915));
  jor  g14724(.dina(n14912), .dinb(n14907), .dout(n14916));
  jnot g14725(.din(n14916), .dout(n14917));
  jor  g14726(.dina(n14804), .dinb(n8215), .dout(n14918));
  jand g14727(.dina(n14918), .dinb(n14917), .dout(n14919));
  jor  g14728(.dina(n14919), .dinb(n14915), .dout(n14920));
  jand g14729(.dina(\a[60] ), .dinb(\a[44] ), .dout(n14921));
  jand g14730(.dina(\a[61] ), .dinb(\a[43] ), .dout(n14922));
  jor  g14731(.dina(n14922), .dinb(n14782), .dout(n14923));
  jand g14732(.dina(n13790), .dinb(n12907), .dout(n14924));
  jnot g14733(.din(n14924), .dout(n14925));
  jand g14734(.dina(n14925), .dinb(n14923), .dout(n14926));
  jxor g14735(.dina(n14926), .dinb(n14921), .dout(n14927));
  jxor g14736(.dina(n14927), .dinb(n14920), .dout(n14928));
  jxor g14737(.dina(n14928), .dinb(n14904), .dout(n14929));
  jxor g14738(.dina(n14929), .dinb(n14889), .dout(n14930));
  jxor g14739(.dina(n14930), .dinb(n14877), .dout(n14931));
  jxor g14740(.dina(n14931), .dinb(n14872), .dout(n14932));
  jand g14741(.dina(n14932), .dinb(n14842), .dout(n14933));
  jor  g14742(.dina(n14932), .dinb(n14842), .dout(n14934));
  jnot g14743(.din(n14934), .dout(n14935));
  jor  g14744(.dina(n14935), .dinb(n14933), .dout(n14936));
  jnot g14745(.din(n14829), .dout(n14937));
  jor  g14746(.dina(n14838), .dinb(n14831), .dout(n14938));
  jand g14747(.dina(n14938), .dinb(n14937), .dout(n14939));
  jxor g14748(.dina(n14939), .dinb(n14936), .dout(\asquared[105] ));
  jand g14749(.dina(n14926), .dinb(n14921), .dout(n14941));
  jor  g14750(.dina(n14941), .dinb(n14924), .dout(n14942));
  jxor g14751(.dina(n14916), .dinb(n14900), .dout(n14943));
  jxor g14752(.dina(n14943), .dinb(n14942), .dout(n14944));
  jand g14753(.dina(n14927), .dinb(n14920), .dout(n14945));
  jand g14754(.dina(n14928), .dinb(n14904), .dout(n14946));
  jor  g14755(.dina(n14946), .dinb(n14945), .dout(n14947));
  jxor g14756(.dina(n14947), .dinb(n14944), .dout(n14948));
  jand g14757(.dina(n14866), .dinb(n14854), .dout(n14949));
  jand g14758(.dina(n14870), .dinb(n14867), .dout(n14950));
  jor  g14759(.dina(n14950), .dinb(n14949), .dout(n14951));
  jxor g14760(.dina(n14951), .dinb(n14948), .dout(n14952));
  jnot g14761(.din(n14952), .dout(n14953));
  jor  g14762(.dina(n14850), .dinb(n14846), .dout(n14954));
  jand g14763(.dina(n14871), .dinb(n14851), .dout(n14955));
  jnot g14764(.din(n14955), .dout(n14956));
  jand g14765(.dina(n14956), .dinb(n14954), .dout(n14957));
  jxor g14766(.dina(n14957), .dinb(n14953), .dout(n14958));
  jor  g14767(.dina(n14888), .dinb(n14885), .dout(n14959));
  jand g14768(.dina(n14929), .dinb(n14889), .dout(n14960));
  jnot g14769(.din(n14960), .dout(n14961));
  jand g14770(.dina(n14961), .dinb(n14959), .dout(n14962));
  jnot g14771(.din(n14962), .dout(n14963));
  jand g14772(.dina(n14882), .dinb(n14879), .dout(n14964));
  jand g14773(.dina(n14883), .dinb(n14793), .dout(n14965));
  jor  g14774(.dina(n14965), .dinb(n14964), .dout(n14966));
  jand g14775(.dina(\a[62] ), .dinb(\a[43] ), .dout(n14967));
  jand g14776(.dina(\a[53] ), .dinb(n14862), .dout(n14968));
  jxor g14777(.dina(n14968), .dinb(n14967), .dout(n14969));
  jnot g14778(.din(n14969), .dout(n14970));
  jand g14779(.dina(\a[56] ), .dinb(\a[49] ), .dout(n14971));
  jnot g14780(.din(n14971), .dout(n14972));
  jand g14781(.dina(\a[55] ), .dinb(\a[51] ), .dout(n14973));
  jand g14782(.dina(n14973), .dinb(n14812), .dout(n14974));
  jnot g14783(.din(n14974), .dout(n14975));
  jand g14784(.dina(\a[54] ), .dinb(\a[51] ), .dout(n14976));
  jor  g14785(.dina(n14976), .dinb(n14894), .dout(n14977));
  jand g14786(.dina(n14977), .dinb(n14975), .dout(n14978));
  jxor g14787(.dina(n14978), .dinb(n14972), .dout(n14979));
  jxor g14788(.dina(n14979), .dinb(n14970), .dout(n14980));
  jxor g14789(.dina(n14980), .dinb(n14966), .dout(n14981));
  jand g14790(.dina(n14865), .dinb(n14861), .dout(n14982));
  jor  g14791(.dina(n14982), .dinb(n14856), .dout(n14983));
  jnot g14792(.din(n14983), .dout(n14984));
  jnot g14793(.din(n14855), .dout(n14985));
  jand g14794(.dina(\a[61] ), .dinb(\a[45] ), .dout(n14986));
  jand g14795(.dina(n14986), .dinb(n14921), .dout(n14987));
  jnot g14796(.din(n14987), .dout(n14988));
  jand g14797(.dina(\a[61] ), .dinb(\a[44] ), .dout(n14989));
  jand g14798(.dina(\a[60] ), .dinb(\a[45] ), .dout(n14990));
  jor  g14799(.dina(n14990), .dinb(n14989), .dout(n14991));
  jand g14800(.dina(n14991), .dinb(n14988), .dout(n14992));
  jxor g14801(.dina(n14992), .dinb(n14985), .dout(n14993));
  jxor g14802(.dina(n14993), .dinb(n14984), .dout(n14994));
  jnot g14803(.din(n14994), .dout(n14995));
  jand g14804(.dina(\a[59] ), .dinb(\a[46] ), .dout(n14996));
  jnot g14805(.din(n14996), .dout(n14997));
  jand g14806(.dina(n7519), .dinb(n5316), .dout(n14998));
  jnot g14807(.din(n14998), .dout(n14999));
  jor  g14808(.dina(n14909), .dinb(n14906), .dout(n15000));
  jand g14809(.dina(n15000), .dinb(n14999), .dout(n15001));
  jxor g14810(.dina(n15001), .dinb(n14997), .dout(n15002));
  jxor g14811(.dina(n15002), .dinb(n14995), .dout(n15003));
  jxor g14812(.dina(n15003), .dinb(n14981), .dout(n15004));
  jxor g14813(.dina(n15004), .dinb(n14963), .dout(n15005));
  jxor g14814(.dina(n15005), .dinb(n14958), .dout(n15006));
  jand g14815(.dina(n14930), .dinb(n14877), .dout(n15007));
  jand g14816(.dina(n14931), .dinb(n14872), .dout(n15008));
  jor  g14817(.dina(n15008), .dinb(n15007), .dout(n15009));
  jnot g14818(.din(n15009), .dout(n15010));
  jxor g14819(.dina(n15010), .dinb(n15006), .dout(n15011));
  jnot g14820(.din(n14933), .dout(n15012));
  jor  g14821(.dina(n14939), .dinb(n14935), .dout(n15013));
  jand g14822(.dina(n15013), .dinb(n15012), .dout(n15014));
  jxor g14823(.dina(n15014), .dinb(n15011), .dout(\asquared[106] ));
  jor  g14824(.dina(n14957), .dinb(n14953), .dout(n15016));
  jand g14825(.dina(n15005), .dinb(n14958), .dout(n15017));
  jnot g14826(.din(n15017), .dout(n15018));
  jand g14827(.dina(n15018), .dinb(n15016), .dout(n15019));
  jand g14828(.dina(\a[63] ), .dinb(\a[43] ), .dout(n15020));
  jor  g14829(.dina(n14967), .dinb(\a[52] ), .dout(n15021));
  jand g14830(.dina(n15021), .dinb(\a[53] ), .dout(n15022));
  jxor g14831(.dina(n15022), .dinb(n15020), .dout(n15023));
  jand g14832(.dina(n14975), .dinb(n14972), .dout(n15024));
  jnot g14833(.din(n15024), .dout(n15025));
  jand g14834(.dina(n15025), .dinb(n14977), .dout(n15026));
  jxor g14835(.dina(n15026), .dinb(n15023), .dout(n15027));
  jnot g14836(.din(n15027), .dout(n15028));
  jor  g14837(.dina(n14993), .dinb(n14984), .dout(n15029));
  jor  g14838(.dina(n15002), .dinb(n14995), .dout(n15030));
  jand g14839(.dina(n15030), .dinb(n15029), .dout(n15031));
  jxor g14840(.dina(n15031), .dinb(n15028), .dout(n15032));
  jnot g14841(.din(n15032), .dout(n15033));
  jor  g14842(.dina(n14979), .dinb(n14970), .dout(n15034));
  jand g14843(.dina(n14980), .dinb(n14966), .dout(n15035));
  jnot g14844(.din(n15035), .dout(n15036));
  jand g14845(.dina(n15036), .dinb(n15034), .dout(n15037));
  jxor g14846(.dina(n15037), .dinb(n15033), .dout(n15038));
  jand g14847(.dina(n15003), .dinb(n14981), .dout(n15039));
  jand g14848(.dina(n15004), .dinb(n14963), .dout(n15040));
  jor  g14849(.dina(n15040), .dinb(n15039), .dout(n15041));
  jxor g14850(.dina(n15041), .dinb(n15038), .dout(n15042));
  jand g14851(.dina(n14947), .dinb(n14944), .dout(n15043));
  jand g14852(.dina(n14951), .dinb(n14948), .dout(n15044));
  jor  g14853(.dina(n15044), .dinb(n15043), .dout(n15045));
  jand g14854(.dina(n14916), .dinb(n14900), .dout(n15046));
  jand g14855(.dina(n14943), .dinb(n14942), .dout(n15047));
  jor  g14856(.dina(n15047), .dinb(n15046), .dout(n15048));
  jand g14857(.dina(\a[59] ), .dinb(\a[47] ), .dout(n15049));
  jand g14858(.dina(n7729), .dinb(n7519), .dout(n15050));
  jnot g14859(.din(n15050), .dout(n15051));
  jand g14860(.dina(\a[58] ), .dinb(\a[48] ), .dout(n15052));
  jor  g14861(.dina(n15052), .dinb(n10644), .dout(n15053));
  jand g14862(.dina(n15053), .dinb(n15051), .dout(n15054));
  jxor g14863(.dina(n15054), .dinb(n15049), .dout(n15055));
  jnot g14864(.din(n15055), .dout(n15056));
  jand g14865(.dina(\a[56] ), .dinb(\a[50] ), .dout(n15057));
  jnot g14866(.din(n15057), .dout(n15058));
  jand g14867(.dina(\a[55] ), .dinb(\a[52] ), .dout(n15059));
  jand g14868(.dina(n15059), .dinb(n14976), .dout(n15060));
  jnot g14869(.din(n15060), .dout(n15061));
  jor  g14870(.dina(n14973), .dinb(n10048), .dout(n15062));
  jand g14871(.dina(n15062), .dinb(n15061), .dout(n15063));
  jxor g14872(.dina(n15063), .dinb(n15058), .dout(n15064));
  jxor g14873(.dina(n15064), .dinb(n15056), .dout(n15065));
  jxor g14874(.dina(n15065), .dinb(n15048), .dout(n15066));
  jand g14875(.dina(n14999), .dinb(n14997), .dout(n15067));
  jnot g14876(.din(n15067), .dout(n15068));
  jand g14877(.dina(n15068), .dinb(n15000), .dout(n15069));
  jand g14878(.dina(n14988), .dinb(n14985), .dout(n15070));
  jnot g14879(.din(n15070), .dout(n15071));
  jand g14880(.dina(n15071), .dinb(n14991), .dout(n15072));
  jxor g14881(.dina(n15072), .dinb(n15069), .dout(n15073));
  jand g14882(.dina(\a[62] ), .dinb(\a[44] ), .dout(n15074));
  jand g14883(.dina(\a[61] ), .dinb(\a[46] ), .dout(n15075));
  jand g14884(.dina(n15075), .dinb(n14990), .dout(n15076));
  jnot g14885(.din(n15076), .dout(n15077));
  jand g14886(.dina(n8702), .dinb(n4812), .dout(n15078));
  jand g14887(.dina(\a[60] ), .dinb(\a[46] ), .dout(n15079));
  jand g14888(.dina(n15079), .dinb(n15074), .dout(n15080));
  jor  g14889(.dina(n15080), .dinb(n15078), .dout(n15081));
  jand g14890(.dina(n15081), .dinb(n15077), .dout(n15082));
  jnot g14891(.din(n15082), .dout(n15083));
  jand g14892(.dina(n15083), .dinb(n15074), .dout(n15084));
  jor  g14893(.dina(n15081), .dinb(n15076), .dout(n15085));
  jnot g14894(.din(n15085), .dout(n15086));
  jor  g14895(.dina(n15079), .dinb(n14986), .dout(n15087));
  jand g14896(.dina(n15087), .dinb(n15086), .dout(n15088));
  jor  g14897(.dina(n15088), .dinb(n15084), .dout(n15089));
  jxor g14898(.dina(n15089), .dinb(n15073), .dout(n15090));
  jxor g14899(.dina(n15090), .dinb(n15066), .dout(n15091));
  jxor g14900(.dina(n15091), .dinb(n15045), .dout(n15092));
  jxor g14901(.dina(n15092), .dinb(n15042), .dout(n15093));
  jxor g14902(.dina(n15093), .dinb(n15019), .dout(n15094));
  jand g14903(.dina(n15009), .dinb(n15006), .dout(n15095));
  jnot g14904(.din(n15095), .dout(n15096));
  jnot g14905(.din(n15006), .dout(n15097));
  jand g14906(.dina(n15010), .dinb(n15097), .dout(n15098));
  jor  g14907(.dina(n15014), .dinb(n15098), .dout(n15099));
  jand g14908(.dina(n15099), .dinb(n15096), .dout(n15100));
  jxor g14909(.dina(n15100), .dinb(n15094), .dout(\asquared[107] ));
  jand g14910(.dina(n15041), .dinb(n15038), .dout(n15102));
  jand g14911(.dina(n15092), .dinb(n15042), .dout(n15103));
  jor  g14912(.dina(n15103), .dinb(n15102), .dout(n15104));
  jor  g14913(.dina(n15031), .dinb(n15028), .dout(n15105));
  jor  g14914(.dina(n15037), .dinb(n15033), .dout(n15106));
  jand g14915(.dina(n15106), .dinb(n15105), .dout(n15107));
  jnot g14916(.din(n15107), .dout(n15108));
  jand g14917(.dina(n15054), .dinb(n15049), .dout(n15109));
  jor  g14918(.dina(n15109), .dinb(n15050), .dout(n15110));
  jxor g14919(.dina(n15110), .dinb(n15085), .dout(n15111));
  jnot g14920(.din(n15111), .dout(n15112));
  jand g14921(.dina(\a[59] ), .dinb(\a[48] ), .dout(n15113));
  jnot g14922(.din(n15113), .dout(n15114));
  jand g14923(.dina(\a[63] ), .dinb(\a[58] ), .dout(n15115));
  jand g14924(.dina(n15115), .dinb(n7033), .dout(n15116));
  jnot g14925(.din(n15116), .dout(n15117));
  jand g14926(.dina(\a[58] ), .dinb(\a[49] ), .dout(n15118));
  jand g14927(.dina(\a[63] ), .dinb(\a[44] ), .dout(n15119));
  jor  g14928(.dina(n15119), .dinb(n15118), .dout(n15120));
  jand g14929(.dina(n15120), .dinb(n15117), .dout(n15121));
  jxor g14930(.dina(n15121), .dinb(n15114), .dout(n15122));
  jxor g14931(.dina(n15122), .dinb(n15112), .dout(n15123));
  jand g14932(.dina(\a[62] ), .dinb(\a[45] ), .dout(n15124));
  jnot g14933(.din(\a[53] ), .dout(n15125));
  jand g14934(.dina(\a[54] ), .dinb(n15125), .dout(n15126));
  jxor g14935(.dina(n15126), .dinb(n15124), .dout(n15127));
  jnot g14936(.din(n15127), .dout(n15128));
  jand g14937(.dina(\a[57] ), .dinb(\a[50] ), .dout(n15129));
  jnot g14938(.din(n15129), .dout(n15130));
  jand g14939(.dina(\a[56] ), .dinb(\a[52] ), .dout(n15131));
  jand g14940(.dina(n15131), .dinb(n14973), .dout(n15132));
  jnot g14941(.din(n15132), .dout(n15133));
  jand g14942(.dina(\a[56] ), .dinb(\a[51] ), .dout(n15134));
  jor  g14943(.dina(n15134), .dinb(n15059), .dout(n15135));
  jand g14944(.dina(n15135), .dinb(n15133), .dout(n15136));
  jxor g14945(.dina(n15136), .dinb(n15130), .dout(n15137));
  jxor g14946(.dina(n15137), .dinb(n15128), .dout(n15138));
  jand g14947(.dina(\a[61] ), .dinb(\a[47] ), .dout(n15139));
  jand g14948(.dina(n15139), .dinb(n15079), .dout(n15140));
  jnot g14949(.din(n15140), .dout(n15141));
  jand g14950(.dina(\a[60] ), .dinb(\a[47] ), .dout(n15142));
  jor  g14951(.dina(n15142), .dinb(n15075), .dout(n15143));
  jand g14952(.dina(n15143), .dinb(n15141), .dout(n15144));
  jand g14953(.dina(n15061), .dinb(n15058), .dout(n15145));
  jnot g14954(.din(n15145), .dout(n15146));
  jand g14955(.dina(n15146), .dinb(n15062), .dout(n15147));
  jxor g14956(.dina(n15147), .dinb(n15144), .dout(n15148));
  jxor g14957(.dina(n15148), .dinb(n15138), .dout(n15149));
  jxor g14958(.dina(n15149), .dinb(n15123), .dout(n15150));
  jxor g14959(.dina(n15150), .dinb(n15108), .dout(n15151));
  jand g14960(.dina(n15090), .dinb(n15066), .dout(n15152));
  jand g14961(.dina(n15091), .dinb(n15045), .dout(n15153));
  jor  g14962(.dina(n15153), .dinb(n15152), .dout(n15154));
  jand g14963(.dina(n15072), .dinb(n15069), .dout(n15155));
  jand g14964(.dina(n15089), .dinb(n15073), .dout(n15156));
  jor  g14965(.dina(n15156), .dinb(n15155), .dout(n15157));
  jand g14966(.dina(n15022), .dinb(n15020), .dout(n15158));
  jand g14967(.dina(n15026), .dinb(n15023), .dout(n15159));
  jor  g14968(.dina(n15159), .dinb(n15158), .dout(n15160));
  jxor g14969(.dina(n15160), .dinb(n15157), .dout(n15161));
  jnot g14970(.din(n15161), .dout(n15162));
  jor  g14971(.dina(n15064), .dinb(n15056), .dout(n15163));
  jand g14972(.dina(n15065), .dinb(n15048), .dout(n15164));
  jnot g14973(.din(n15164), .dout(n15165));
  jand g14974(.dina(n15165), .dinb(n15163), .dout(n15166));
  jxor g14975(.dina(n15166), .dinb(n15162), .dout(n15167));
  jxor g14976(.dina(n15167), .dinb(n15154), .dout(n15168));
  jxor g14977(.dina(n15168), .dinb(n15151), .dout(n15169));
  jnot g14978(.din(n15169), .dout(n15170));
  jxor g14979(.dina(n15170), .dinb(n15104), .dout(n15171));
  jnot g14980(.din(n15019), .dout(n15172));
  jand g14981(.dina(n15093), .dinb(n15172), .dout(n15173));
  jnot g14982(.din(n15173), .dout(n15174));
  jor  g14983(.dina(n15093), .dinb(n15172), .dout(n15175));
  jnot g14984(.din(n15175), .dout(n15176));
  jor  g14985(.dina(n15100), .dinb(n15176), .dout(n15177));
  jand g14986(.dina(n15177), .dinb(n15174), .dout(n15178));
  jxor g14987(.dina(n15178), .dinb(n15171), .dout(\asquared[108] ));
  jand g14988(.dina(n15167), .dinb(n15154), .dout(n15180));
  jand g14989(.dina(n15168), .dinb(n15151), .dout(n15181));
  jor  g14990(.dina(n15181), .dinb(n15180), .dout(n15182));
  jnot g14991(.din(n15182), .dout(n15183));
  jand g14992(.dina(n15149), .dinb(n15123), .dout(n15184));
  jand g14993(.dina(n15150), .dinb(n15108), .dout(n15185));
  jor  g14994(.dina(n15185), .dinb(n15184), .dout(n15186));
  jor  g14995(.dina(n15137), .dinb(n15128), .dout(n15187));
  jand g14996(.dina(n15148), .dinb(n15138), .dout(n15188));
  jnot g14997(.din(n15188), .dout(n15189));
  jand g14998(.dina(n15189), .dinb(n15187), .dout(n15190));
  jnot g14999(.din(n15190), .dout(n15191));
  jand g15000(.dina(n15110), .dinb(n15085), .dout(n15192));
  jnot g15001(.din(n15192), .dout(n15193));
  jor  g15002(.dina(n15122), .dinb(n15112), .dout(n15194));
  jand g15003(.dina(n15194), .dinb(n15193), .dout(n15195));
  jnot g15004(.din(n12083), .dout(n15196));
  jand g15005(.dina(\a[56] ), .dinb(\a[53] ), .dout(n15197));
  jand g15006(.dina(n15197), .dinb(n15059), .dout(n15198));
  jnot g15007(.din(n15198), .dout(n15199));
  jor  g15008(.dina(n15131), .dinb(n6498), .dout(n15200));
  jand g15009(.dina(n15200), .dinb(n15199), .dout(n15201));
  jxor g15010(.dina(n15201), .dinb(n15196), .dout(n15202));
  jxor g15011(.dina(n15202), .dinb(n15195), .dout(n15203));
  jxor g15012(.dina(n15203), .dinb(n15191), .dout(n15204));
  jxor g15013(.dina(n15204), .dinb(n15186), .dout(n15205));
  jand g15014(.dina(n15133), .dinb(n15130), .dout(n15206));
  jnot g15015(.din(n15206), .dout(n15207));
  jand g15016(.dina(n15207), .dinb(n15135), .dout(n15208));
  jor  g15017(.dina(n15124), .dinb(\a[53] ), .dout(n15209));
  jand g15018(.dina(n15209), .dinb(\a[54] ), .dout(n15210));
  jxor g15019(.dina(n15210), .dinb(n15208), .dout(n15211));
  jand g15020(.dina(n15117), .dinb(n15114), .dout(n15212));
  jnot g15021(.din(n15212), .dout(n15213));
  jand g15022(.dina(n15213), .dinb(n15120), .dout(n15214));
  jxor g15023(.dina(n15214), .dinb(n15211), .dout(n15215));
  jnot g15024(.din(n15215), .dout(n15216));
  jand g15025(.dina(n15160), .dinb(n15157), .dout(n15217));
  jnot g15026(.din(n15217), .dout(n15218));
  jor  g15027(.dina(n15166), .dinb(n15162), .dout(n15219));
  jand g15028(.dina(n15219), .dinb(n15218), .dout(n15220));
  jxor g15029(.dina(n15220), .dinb(n15216), .dout(n15221));
  jand g15030(.dina(n15147), .dinb(n15144), .dout(n15222));
  jor  g15031(.dina(n15222), .dinb(n15140), .dout(n15223));
  jand g15032(.dina(\a[63] ), .dinb(\a[45] ), .dout(n15224));
  jnot g15033(.din(n15224), .dout(n15225));
  jand g15034(.dina(\a[62] ), .dinb(\a[47] ), .dout(n15226));
  jand g15035(.dina(n15226), .dinb(n15075), .dout(n15227));
  jnot g15036(.din(n15227), .dout(n15228));
  jand g15037(.dina(\a[62] ), .dinb(\a[46] ), .dout(n15229));
  jor  g15038(.dina(n15229), .dinb(n15139), .dout(n15230));
  jand g15039(.dina(n15230), .dinb(n15228), .dout(n15231));
  jxor g15040(.dina(n15231), .dinb(n15225), .dout(n15232));
  jnot g15041(.din(n15232), .dout(n15233));
  jxor g15042(.dina(n15233), .dinb(n15223), .dout(n15234));
  jnot g15043(.din(n15234), .dout(n15235));
  jand g15044(.dina(\a[60] ), .dinb(\a[48] ), .dout(n15236));
  jnot g15045(.din(n15236), .dout(n15237));
  jand g15046(.dina(\a[59] ), .dinb(\a[50] ), .dout(n15238));
  jand g15047(.dina(n15238), .dinb(n15118), .dout(n15239));
  jnot g15048(.din(n15239), .dout(n15240));
  jand g15049(.dina(\a[58] ), .dinb(\a[50] ), .dout(n15241));
  jand g15050(.dina(\a[59] ), .dinb(\a[49] ), .dout(n15242));
  jor  g15051(.dina(n15242), .dinb(n15241), .dout(n15243));
  jand g15052(.dina(n15243), .dinb(n15240), .dout(n15244));
  jxor g15053(.dina(n15244), .dinb(n15237), .dout(n15245));
  jxor g15054(.dina(n15245), .dinb(n15235), .dout(n15246));
  jxor g15055(.dina(n15246), .dinb(n15221), .dout(n15247));
  jxor g15056(.dina(n15247), .dinb(n15205), .dout(n15248));
  jxor g15057(.dina(n15248), .dinb(n15183), .dout(n15249));
  jand g15058(.dina(n15169), .dinb(n15104), .dout(n15250));
  jnot g15059(.din(n15250), .dout(n15251));
  jnot g15060(.din(n15104), .dout(n15252));
  jand g15061(.dina(n15170), .dinb(n15252), .dout(n15253));
  jor  g15062(.dina(n15178), .dinb(n15253), .dout(n15254));
  jand g15063(.dina(n15254), .dinb(n15251), .dout(n15255));
  jxor g15064(.dina(n15255), .dinb(n15249), .dout(\asquared[109] ));
  jand g15065(.dina(n15204), .dinb(n15186), .dout(n15257));
  jand g15066(.dina(n15247), .dinb(n15205), .dout(n15258));
  jor  g15067(.dina(n15258), .dinb(n15257), .dout(n15259));
  jand g15068(.dina(n15233), .dinb(n15223), .dout(n15260));
  jnot g15069(.din(n15260), .dout(n15261));
  jor  g15070(.dina(n15245), .dinb(n15235), .dout(n15262));
  jand g15071(.dina(n15262), .dinb(n15261), .dout(n15263));
  jnot g15072(.din(n15263), .dout(n15264));
  jand g15073(.dina(n15210), .dinb(n15208), .dout(n15265));
  jand g15074(.dina(n15214), .dinb(n15211), .dout(n15266));
  jor  g15075(.dina(n15266), .dinb(n15265), .dout(n15267));
  jnot g15076(.din(n15267), .dout(n15268));
  jnot g15077(.din(n15226), .dout(n15269));
  jand g15078(.dina(\a[55] ), .dinb(n6399), .dout(n15270));
  jxor g15079(.dina(n15270), .dinb(n15269), .dout(n15271));
  jxor g15080(.dina(n15271), .dinb(n15268), .dout(n15272));
  jxor g15081(.dina(n15272), .dinb(n15264), .dout(n15273));
  jnot g15082(.din(n15273), .dout(n15274));
  jor  g15083(.dina(n15220), .dinb(n15216), .dout(n15275));
  jand g15084(.dina(n15246), .dinb(n15221), .dout(n15276));
  jnot g15085(.din(n15276), .dout(n15277));
  jand g15086(.dina(n15277), .dinb(n15275), .dout(n15278));
  jxor g15087(.dina(n15278), .dinb(n15274), .dout(n15279));
  jand g15088(.dina(\a[63] ), .dinb(\a[46] ), .dout(n15280));
  jand g15089(.dina(n15199), .dinb(n15196), .dout(n15281));
  jnot g15090(.din(n15281), .dout(n15282));
  jand g15091(.dina(n15282), .dinb(n15200), .dout(n15283));
  jxor g15092(.dina(n15283), .dinb(n15280), .dout(n15284));
  jand g15093(.dina(n15240), .dinb(n15237), .dout(n15285));
  jnot g15094(.din(n15285), .dout(n15286));
  jand g15095(.dina(n15286), .dinb(n15243), .dout(n15287));
  jxor g15096(.dina(n15287), .dinb(n15284), .dout(n15288));
  jnot g15097(.din(n15288), .dout(n15289));
  jor  g15098(.dina(n15202), .dinb(n15195), .dout(n15290));
  jand g15099(.dina(n15203), .dinb(n15191), .dout(n15291));
  jnot g15100(.din(n15291), .dout(n15292));
  jand g15101(.dina(n15292), .dinb(n15290), .dout(n15293));
  jxor g15102(.dina(n15293), .dinb(n15289), .dout(n15294));
  jand g15103(.dina(n15228), .dinb(n15225), .dout(n15295));
  jnot g15104(.din(n15295), .dout(n15296));
  jand g15105(.dina(n15296), .dinb(n15230), .dout(n15297));
  jand g15106(.dina(\a[61] ), .dinb(\a[48] ), .dout(n15298));
  jand g15107(.dina(\a[60] ), .dinb(\a[50] ), .dout(n15299));
  jand g15108(.dina(n15299), .dinb(n15242), .dout(n15300));
  jnot g15109(.din(n15300), .dout(n15301));
  jand g15110(.dina(\a[60] ), .dinb(\a[49] ), .dout(n15302));
  jor  g15111(.dina(n15302), .dinb(n15238), .dout(n15303));
  jand g15112(.dina(n15303), .dinb(n15301), .dout(n15304));
  jxor g15113(.dina(n15304), .dinb(n15298), .dout(n15305));
  jxor g15114(.dina(n15305), .dinb(n15297), .dout(n15306));
  jnot g15115(.din(n15306), .dout(n15307));
  jand g15116(.dina(\a[58] ), .dinb(\a[51] ), .dout(n15308));
  jnot g15117(.din(n15308), .dout(n15309));
  jand g15118(.dina(\a[57] ), .dinb(\a[53] ), .dout(n15310));
  jand g15119(.dina(n15310), .dinb(n15131), .dout(n15311));
  jnot g15120(.din(n15311), .dout(n15312));
  jand g15121(.dina(\a[57] ), .dinb(\a[52] ), .dout(n15313));
  jor  g15122(.dina(n15313), .dinb(n15197), .dout(n15314));
  jand g15123(.dina(n15314), .dinb(n15312), .dout(n15315));
  jxor g15124(.dina(n15315), .dinb(n15309), .dout(n15316));
  jxor g15125(.dina(n15316), .dinb(n15307), .dout(n15317));
  jxor g15126(.dina(n15317), .dinb(n15294), .dout(n15318));
  jxor g15127(.dina(n15318), .dinb(n15279), .dout(n15319));
  jand g15128(.dina(n15319), .dinb(n15259), .dout(n15320));
  jor  g15129(.dina(n15319), .dinb(n15259), .dout(n15321));
  jnot g15130(.din(n15321), .dout(n15322));
  jor  g15131(.dina(n15322), .dinb(n15320), .dout(n15323));
  jand g15132(.dina(n15248), .dinb(n15182), .dout(n15324));
  jnot g15133(.din(n15324), .dout(n15325));
  jnot g15134(.din(n15248), .dout(n15326));
  jand g15135(.dina(n15326), .dinb(n15183), .dout(n15327));
  jor  g15136(.dina(n15255), .dinb(n15327), .dout(n15328));
  jand g15137(.dina(n15328), .dinb(n15325), .dout(n15329));
  jxor g15138(.dina(n15329), .dinb(n15323), .dout(\asquared[110] ));
  jor  g15139(.dina(n15278), .dinb(n15274), .dout(n15331));
  jand g15140(.dina(n15318), .dinb(n15279), .dout(n15332));
  jnot g15141(.din(n15332), .dout(n15333));
  jand g15142(.dina(n15333), .dinb(n15331), .dout(n15334));
  jand g15143(.dina(n15305), .dinb(n15297), .dout(n15335));
  jnot g15144(.din(n15335), .dout(n15336));
  jor  g15145(.dina(n15316), .dinb(n15307), .dout(n15337));
  jand g15146(.dina(n15337), .dinb(n15336), .dout(n15338));
  jnot g15147(.din(n15338), .dout(n15339));
  jand g15148(.dina(n15312), .dinb(n15309), .dout(n15340));
  jnot g15149(.din(n15340), .dout(n15341));
  jand g15150(.dina(n15341), .dinb(n15314), .dout(n15342));
  jor  g15151(.dina(n15300), .dinb(n15298), .dout(n15343));
  jand g15152(.dina(n15343), .dinb(n15303), .dout(n15344));
  jxor g15153(.dina(n15344), .dinb(n15342), .dout(n15345));
  jand g15154(.dina(\a[61] ), .dinb(\a[49] ), .dout(n15346));
  jnot g15155(.din(n15346), .dout(n15347));
  jand g15156(.dina(\a[60] ), .dinb(\a[51] ), .dout(n15348));
  jand g15157(.dina(n15348), .dinb(n15238), .dout(n15349));
  jnot g15158(.din(n15349), .dout(n15350));
  jand g15159(.dina(\a[59] ), .dinb(\a[51] ), .dout(n15351));
  jor  g15160(.dina(n15351), .dinb(n15299), .dout(n15352));
  jand g15161(.dina(n15352), .dinb(n15350), .dout(n15353));
  jxor g15162(.dina(n15353), .dinb(n15347), .dout(n15354));
  jnot g15163(.din(n15354), .dout(n15355));
  jxor g15164(.dina(n15355), .dinb(n15345), .dout(n15356));
  jxor g15165(.dina(n15356), .dinb(n15339), .dout(n15357));
  jnot g15166(.din(n15357), .dout(n15358));
  jor  g15167(.dina(n15271), .dinb(n15268), .dout(n15359));
  jand g15168(.dina(n15272), .dinb(n15264), .dout(n15360));
  jnot g15169(.din(n15360), .dout(n15361));
  jand g15170(.dina(n15361), .dinb(n15359), .dout(n15362));
  jxor g15171(.dina(n15362), .dinb(n15358), .dout(n15363));
  jand g15172(.dina(n15283), .dinb(n15280), .dout(n15364));
  jand g15173(.dina(n15287), .dinb(n15284), .dout(n15365));
  jor  g15174(.dina(n15365), .dinb(n15364), .dout(n15366));
  jand g15175(.dina(\a[63] ), .dinb(\a[48] ), .dout(n15367));
  jand g15176(.dina(n15367), .dinb(n15226), .dout(n15368));
  jnot g15177(.din(n15368), .dout(n15369));
  jand g15178(.dina(\a[63] ), .dinb(\a[47] ), .dout(n15370));
  jand g15179(.dina(\a[62] ), .dinb(\a[48] ), .dout(n15371));
  jor  g15180(.dina(n15371), .dinb(n15370), .dout(n15372));
  jand g15181(.dina(n15372), .dinb(n15369), .dout(n15373));
  jand g15182(.dina(n15269), .dinb(n6399), .dout(n15374));
  jor  g15183(.dina(n15374), .dinb(n6143), .dout(n15375));
  jnot g15184(.din(n15375), .dout(n15376));
  jxor g15185(.dina(n15376), .dinb(n15373), .dout(n15377));
  jand g15186(.dina(\a[58] ), .dinb(\a[52] ), .dout(n15378));
  jand g15187(.dina(n15197), .dinb(n13620), .dout(n15379));
  jnot g15188(.din(n15379), .dout(n15380));
  jand g15189(.dina(n7519), .dinb(n7165), .dout(n15381));
  jand g15190(.dina(n15378), .dinb(n11191), .dout(n15382));
  jor  g15191(.dina(n15382), .dinb(n15381), .dout(n15383));
  jand g15192(.dina(n15383), .dinb(n15380), .dout(n15384));
  jnot g15193(.din(n15384), .dout(n15385));
  jand g15194(.dina(n15385), .dinb(n15378), .dout(n15386));
  jor  g15195(.dina(n15383), .dinb(n15379), .dout(n15387));
  jnot g15196(.din(n15387), .dout(n15388));
  jor  g15197(.dina(n15310), .dinb(n11191), .dout(n15389));
  jand g15198(.dina(n15389), .dinb(n15388), .dout(n15390));
  jor  g15199(.dina(n15390), .dinb(n15386), .dout(n15391));
  jxor g15200(.dina(n15391), .dinb(n15377), .dout(n15392));
  jxor g15201(.dina(n15392), .dinb(n15366), .dout(n15393));
  jnot g15202(.din(n15393), .dout(n15394));
  jor  g15203(.dina(n15293), .dinb(n15289), .dout(n15395));
  jand g15204(.dina(n15317), .dinb(n15294), .dout(n15396));
  jnot g15205(.din(n15396), .dout(n15397));
  jand g15206(.dina(n15397), .dinb(n15395), .dout(n15398));
  jxor g15207(.dina(n15398), .dinb(n15394), .dout(n15399));
  jxor g15208(.dina(n15399), .dinb(n15363), .dout(n15400));
  jxor g15209(.dina(n15400), .dinb(n15334), .dout(n15401));
  jnot g15210(.din(n15320), .dout(n15402));
  jor  g15211(.dina(n15329), .dinb(n15322), .dout(n15403));
  jand g15212(.dina(n15403), .dinb(n15402), .dout(n15404));
  jxor g15213(.dina(n15404), .dinb(n15401), .dout(\asquared[111] ));
  jor  g15214(.dina(n15398), .dinb(n15394), .dout(n15406));
  jand g15215(.dina(n15399), .dinb(n15363), .dout(n15407));
  jnot g15216(.din(n15407), .dout(n15408));
  jand g15217(.dina(n15408), .dinb(n15406), .dout(n15409));
  jand g15218(.dina(n15350), .dinb(n15347), .dout(n15410));
  jnot g15219(.din(n15410), .dout(n15411));
  jand g15220(.dina(n15411), .dinb(n15352), .dout(n15412));
  jxor g15221(.dina(n15412), .dinb(n15387), .dout(n15413));
  jand g15222(.dina(n15376), .dinb(n15373), .dout(n15414));
  jor  g15223(.dina(n15414), .dinb(n15368), .dout(n15415));
  jxor g15224(.dina(n15415), .dinb(n15413), .dout(n15416));
  jand g15225(.dina(n15344), .dinb(n15342), .dout(n15417));
  jand g15226(.dina(n15355), .dinb(n15345), .dout(n15418));
  jor  g15227(.dina(n15418), .dinb(n15417), .dout(n15419));
  jxor g15228(.dina(n15419), .dinb(n15416), .dout(n15420));
  jand g15229(.dina(n15391), .dinb(n15377), .dout(n15421));
  jand g15230(.dina(n15392), .dinb(n15366), .dout(n15422));
  jor  g15231(.dina(n15422), .dinb(n15421), .dout(n15423));
  jxor g15232(.dina(n15423), .dinb(n15420), .dout(n15424));
  jand g15233(.dina(n15356), .dinb(n15339), .dout(n15425));
  jnot g15234(.din(n15425), .dout(n15426));
  jor  g15235(.dina(n15362), .dinb(n15358), .dout(n15427));
  jand g15236(.dina(n15427), .dinb(n15426), .dout(n15428));
  jnot g15237(.din(n15428), .dout(n15429));
  jand g15238(.dina(\a[61] ), .dinb(\a[51] ), .dout(n15430));
  jand g15239(.dina(n15430), .dinb(n15299), .dout(n15431));
  jnot g15240(.din(n15431), .dout(n15432));
  jand g15241(.dina(\a[61] ), .dinb(\a[50] ), .dout(n15433));
  jor  g15242(.dina(n15433), .dinb(n15348), .dout(n15434));
  jand g15243(.dina(n15434), .dinb(n15432), .dout(n15435));
  jxor g15244(.dina(n15435), .dinb(n15367), .dout(n15436));
  jnot g15245(.din(n15436), .dout(n15437));
  jand g15246(.dina(\a[62] ), .dinb(\a[49] ), .dout(n15438));
  jnot g15247(.din(n15438), .dout(n15439));
  jand g15248(.dina(\a[56] ), .dinb(n6143), .dout(n15440));
  jxor g15249(.dina(n15440), .dinb(n15439), .dout(n15441));
  jxor g15250(.dina(n15441), .dinb(n15437), .dout(n15442));
  jnot g15251(.din(n15442), .dout(n15443));
  jand g15252(.dina(\a[59] ), .dinb(\a[52] ), .dout(n15444));
  jand g15253(.dina(n7559), .dinb(n7519), .dout(n15445));
  jnot g15254(.din(n13620), .dout(n15446));
  jand g15255(.dina(\a[58] ), .dinb(\a[53] ), .dout(n15447));
  jnot g15256(.din(n15447), .dout(n15448));
  jand g15257(.dina(n15448), .dinb(n15446), .dout(n15449));
  jor  g15258(.dina(n15449), .dinb(n15445), .dout(n15450));
  jxor g15259(.dina(n15450), .dinb(n15444), .dout(n15451));
  jxor g15260(.dina(n15451), .dinb(n15443), .dout(n15452));
  jxor g15261(.dina(n15452), .dinb(n15429), .dout(n15453));
  jxor g15262(.dina(n15453), .dinb(n15424), .dout(n15454));
  jxor g15263(.dina(n15454), .dinb(n15409), .dout(n15455));
  jnot g15264(.din(n15400), .dout(n15456));
  jor  g15265(.dina(n15456), .dinb(n15334), .dout(n15457));
  jand g15266(.dina(n15456), .dinb(n15334), .dout(n15458));
  jor  g15267(.dina(n15404), .dinb(n15458), .dout(n15459));
  jand g15268(.dina(n15459), .dinb(n15457), .dout(n15460));
  jxor g15269(.dina(n15460), .dinb(n15455), .dout(\asquared[112] ));
  jand g15270(.dina(n15452), .dinb(n15429), .dout(n15462));
  jand g15271(.dina(n15453), .dinb(n15424), .dout(n15463));
  jor  g15272(.dina(n15463), .dinb(n15462), .dout(n15464));
  jand g15273(.dina(n15419), .dinb(n15416), .dout(n15465));
  jand g15274(.dina(n15423), .dinb(n15420), .dout(n15466));
  jor  g15275(.dina(n15466), .dinb(n15465), .dout(n15467));
  jand g15276(.dina(\a[59] ), .dinb(\a[53] ), .dout(n15468));
  jand g15277(.dina(\a[58] ), .dinb(\a[55] ), .dout(n15469));
  jand g15278(.dina(n15469), .dinb(n13620), .dout(n15470));
  jnot g15279(.din(n15470), .dout(n15471));
  jand g15280(.dina(\a[59] ), .dinb(\a[54] ), .dout(n15472));
  jand g15281(.dina(n15472), .dinb(n15447), .dout(n15473));
  jand g15282(.dina(n15468), .dinb(n11997), .dout(n15474));
  jor  g15283(.dina(n15474), .dinb(n15473), .dout(n15475));
  jand g15284(.dina(n15475), .dinb(n15471), .dout(n15476));
  jnot g15285(.din(n15476), .dout(n15477));
  jand g15286(.dina(n15477), .dinb(n15468), .dout(n15478));
  jor  g15287(.dina(n15475), .dinb(n15470), .dout(n15479));
  jnot g15288(.din(n15479), .dout(n15480));
  jand g15289(.dina(\a[58] ), .dinb(\a[54] ), .dout(n15481));
  jor  g15290(.dina(n15481), .dinb(n11997), .dout(n15482));
  jand g15291(.dina(n15482), .dinb(n15480), .dout(n15483));
  jor  g15292(.dina(n15483), .dinb(n15478), .dout(n15484));
  jand g15293(.dina(n15435), .dinb(n15367), .dout(n15485));
  jor  g15294(.dina(n15485), .dinb(n15431), .dout(n15486));
  jand g15295(.dina(\a[63] ), .dinb(\a[49] ), .dout(n15487));
  jand g15296(.dina(\a[61] ), .dinb(\a[52] ), .dout(n15488));
  jand g15297(.dina(n15488), .dinb(n15348), .dout(n15489));
  jnot g15298(.din(n15489), .dout(n15490));
  jand g15299(.dina(\a[60] ), .dinb(\a[52] ), .dout(n15491));
  jor  g15300(.dina(n15491), .dinb(n15430), .dout(n15492));
  jand g15301(.dina(n15492), .dinb(n15490), .dout(n15493));
  jxor g15302(.dina(n15493), .dinb(n15487), .dout(n15494));
  jxor g15303(.dina(n15494), .dinb(n15486), .dout(n15495));
  jxor g15304(.dina(n15495), .dinb(n15484), .dout(n15496));
  jxor g15305(.dina(n15496), .dinb(n15467), .dout(n15497));
  jand g15306(.dina(\a[62] ), .dinb(\a[50] ), .dout(n15498));
  jnot g15307(.din(\a[56] ), .dout(n15499));
  jand g15308(.dina(n15439), .dinb(n6143), .dout(n15500));
  jor  g15309(.dina(n15500), .dinb(n15499), .dout(n15501));
  jnot g15310(.din(n15501), .dout(n15502));
  jxor g15311(.dina(n15502), .dinb(n15498), .dout(n15503));
  jnot g15312(.din(n15444), .dout(n15504));
  jnot g15313(.din(n15445), .dout(n15505));
  jand g15314(.dina(n15505), .dinb(n15504), .dout(n15506));
  jor  g15315(.dina(n15506), .dinb(n15449), .dout(n15507));
  jnot g15316(.din(n15507), .dout(n15508));
  jxor g15317(.dina(n15508), .dinb(n15503), .dout(n15509));
  jand g15318(.dina(n15412), .dinb(n15387), .dout(n15510));
  jand g15319(.dina(n15415), .dinb(n15413), .dout(n15511));
  jor  g15320(.dina(n15511), .dinb(n15510), .dout(n15512));
  jnot g15321(.din(n15512), .dout(n15513));
  jor  g15322(.dina(n15441), .dinb(n15437), .dout(n15514));
  jor  g15323(.dina(n15451), .dinb(n15443), .dout(n15515));
  jand g15324(.dina(n15515), .dinb(n15514), .dout(n15516));
  jxor g15325(.dina(n15516), .dinb(n15513), .dout(n15517));
  jxor g15326(.dina(n15517), .dinb(n15509), .dout(n15518));
  jxor g15327(.dina(n15518), .dinb(n15497), .dout(n15519));
  jnot g15328(.din(n15519), .dout(n15520));
  jxor g15329(.dina(n15520), .dinb(n15464), .dout(n15521));
  jnot g15330(.din(n15409), .dout(n15522));
  jand g15331(.dina(n15454), .dinb(n15522), .dout(n15523));
  jnot g15332(.din(n15523), .dout(n15524));
  jor  g15333(.dina(n15454), .dinb(n15522), .dout(n15525));
  jnot g15334(.din(n15525), .dout(n15526));
  jor  g15335(.dina(n15460), .dinb(n15526), .dout(n15527));
  jand g15336(.dina(n15527), .dinb(n15524), .dout(n15528));
  jxor g15337(.dina(n15528), .dinb(n15521), .dout(\asquared[113] ));
  jand g15338(.dina(n15496), .dinb(n15467), .dout(n15530));
  jand g15339(.dina(n15518), .dinb(n15497), .dout(n15531));
  jor  g15340(.dina(n15531), .dinb(n15530), .dout(n15532));
  jnot g15341(.din(n15532), .dout(n15533));
  jand g15342(.dina(n15502), .dinb(n15498), .dout(n15534));
  jand g15343(.dina(n15508), .dinb(n15503), .dout(n15535));
  jor  g15344(.dina(n15535), .dinb(n15534), .dout(n15536));
  jand g15345(.dina(\a[61] ), .dinb(\a[53] ), .dout(n15537));
  jand g15346(.dina(n15537), .dinb(n15491), .dout(n15538));
  jnot g15347(.din(n15538), .dout(n15539));
  jand g15348(.dina(\a[60] ), .dinb(\a[53] ), .dout(n15540));
  jor  g15349(.dina(n15540), .dinb(n15488), .dout(n15541));
  jand g15350(.dina(n15541), .dinb(n15539), .dout(n15542));
  jxor g15351(.dina(n15542), .dinb(n15479), .dout(n15543));
  jxor g15352(.dina(n15543), .dinb(n15536), .dout(n15544));
  jand g15353(.dina(n15494), .dinb(n15486), .dout(n15545));
  jand g15354(.dina(n15495), .dinb(n15484), .dout(n15546));
  jor  g15355(.dina(n15546), .dinb(n15545), .dout(n15547));
  jxor g15356(.dina(n15547), .dinb(n15544), .dout(n15548));
  jor  g15357(.dina(n15516), .dinb(n15513), .dout(n15549));
  jand g15358(.dina(n15517), .dinb(n15509), .dout(n15550));
  jnot g15359(.din(n15550), .dout(n15551));
  jand g15360(.dina(n15551), .dinb(n15549), .dout(n15552));
  jnot g15361(.din(n15552), .dout(n15553));
  jand g15362(.dina(n15492), .dinb(n15487), .dout(n15554));
  jor  g15363(.dina(n15554), .dinb(n15489), .dout(n15555));
  jnot g15364(.din(n15555), .dout(n15556));
  jand g15365(.dina(\a[63] ), .dinb(\a[50] ), .dout(n15557));
  jnot g15366(.din(n15557), .dout(n15558));
  jand g15367(.dina(\a[59] ), .dinb(\a[55] ), .dout(n15559));
  jand g15368(.dina(n15559), .dinb(n15481), .dout(n15560));
  jnot g15369(.din(n15560), .dout(n15561));
  jor  g15370(.dina(n15472), .dinb(n15469), .dout(n15562));
  jand g15371(.dina(n15562), .dinb(n15561), .dout(n15563));
  jxor g15372(.dina(n15563), .dinb(n15558), .dout(n15564));
  jxor g15373(.dina(n15564), .dinb(n15556), .dout(n15565));
  jnot g15374(.din(n15565), .dout(n15566));
  jand g15375(.dina(\a[62] ), .dinb(\a[51] ), .dout(n15567));
  jnot g15376(.din(n15567), .dout(n15568));
  jand g15377(.dina(\a[57] ), .dinb(n15499), .dout(n15569));
  jxor g15378(.dina(n15569), .dinb(n15568), .dout(n15570));
  jxor g15379(.dina(n15570), .dinb(n15566), .dout(n15571));
  jxor g15380(.dina(n15571), .dinb(n15553), .dout(n15572));
  jxor g15381(.dina(n15572), .dinb(n15548), .dout(n15573));
  jxor g15382(.dina(n15573), .dinb(n15533), .dout(n15574));
  jand g15383(.dina(n15519), .dinb(n15464), .dout(n15575));
  jnot g15384(.din(n15575), .dout(n15576));
  jnot g15385(.din(n15464), .dout(n15577));
  jand g15386(.dina(n15520), .dinb(n15577), .dout(n15578));
  jor  g15387(.dina(n15528), .dinb(n15578), .dout(n15579));
  jand g15388(.dina(n15579), .dinb(n15576), .dout(n15580));
  jxor g15389(.dina(n15580), .dinb(n15574), .dout(\asquared[114] ));
  jand g15390(.dina(n15571), .dinb(n15553), .dout(n15582));
  jand g15391(.dina(n15572), .dinb(n15548), .dout(n15583));
  jor  g15392(.dina(n15583), .dinb(n15582), .dout(n15584));
  jnot g15393(.din(\a[57] ), .dout(n15585));
  jand g15394(.dina(n15568), .dinb(n15499), .dout(n15586));
  jor  g15395(.dina(n15586), .dinb(n15585), .dout(n15587));
  jnot g15396(.din(n15587), .dout(n15588));
  jand g15397(.dina(n15561), .dinb(n15558), .dout(n15589));
  jnot g15398(.din(n15589), .dout(n15590));
  jand g15399(.dina(n15590), .dinb(n15562), .dout(n15591));
  jxor g15400(.dina(n15591), .dinb(n15588), .dout(n15592));
  jand g15401(.dina(n15542), .dinb(n15479), .dout(n15593));
  jor  g15402(.dina(n15593), .dinb(n15538), .dout(n15594));
  jxor g15403(.dina(n15594), .dinb(n15592), .dout(n15595));
  jand g15404(.dina(n15543), .dinb(n15536), .dout(n15596));
  jand g15405(.dina(n15547), .dinb(n15544), .dout(n15597));
  jor  g15406(.dina(n15597), .dinb(n15596), .dout(n15598));
  jxor g15407(.dina(n15598), .dinb(n15595), .dout(n15599));
  jor  g15408(.dina(n15564), .dinb(n15556), .dout(n15600));
  jor  g15409(.dina(n15570), .dinb(n15566), .dout(n15601));
  jand g15410(.dina(n15601), .dinb(n15600), .dout(n15602));
  jnot g15411(.din(n15602), .dout(n15603));
  jand g15412(.dina(\a[63] ), .dinb(\a[51] ), .dout(n15604));
  jand g15413(.dina(\a[62] ), .dinb(\a[52] ), .dout(n15605));
  jor  g15414(.dina(n15605), .dinb(n15537), .dout(n15606));
  jand g15415(.dina(n8702), .dinb(n7165), .dout(n15607));
  jnot g15416(.din(n15607), .dout(n15608));
  jand g15417(.dina(n15608), .dinb(n15606), .dout(n15609));
  jxor g15418(.dina(n15609), .dinb(n15604), .dout(n15610));
  jnot g15419(.din(n15610), .dout(n15611));
  jand g15420(.dina(\a[60] ), .dinb(\a[54] ), .dout(n15612));
  jand g15421(.dina(n15469), .dinb(n14039), .dout(n15613));
  jnot g15422(.din(n11688), .dout(n15614));
  jnot g15423(.din(n15559), .dout(n15615));
  jand g15424(.dina(n15615), .dinb(n15614), .dout(n15616));
  jor  g15425(.dina(n15616), .dinb(n15613), .dout(n15617));
  jxor g15426(.dina(n15617), .dinb(n15612), .dout(n15618));
  jxor g15427(.dina(n15618), .dinb(n15611), .dout(n15619));
  jxor g15428(.dina(n15619), .dinb(n15603), .dout(n15620));
  jxor g15429(.dina(n15620), .dinb(n15599), .dout(n15621));
  jnot g15430(.din(n15621), .dout(n15622));
  jxor g15431(.dina(n15622), .dinb(n15584), .dout(n15623));
  jand g15432(.dina(n15573), .dinb(n15532), .dout(n15624));
  jnot g15433(.din(n15624), .dout(n15625));
  jnot g15434(.din(n15573), .dout(n15626));
  jand g15435(.dina(n15626), .dinb(n15533), .dout(n15627));
  jor  g15436(.dina(n15580), .dinb(n15627), .dout(n15628));
  jand g15437(.dina(n15628), .dinb(n15625), .dout(n15629));
  jxor g15438(.dina(n15629), .dinb(n15623), .dout(\asquared[115] ));
  jand g15439(.dina(n15598), .dinb(n15595), .dout(n15631));
  jand g15440(.dina(n15620), .dinb(n15599), .dout(n15632));
  jor  g15441(.dina(n15632), .dinb(n15631), .dout(n15633));
  jand g15442(.dina(n15591), .dinb(n15588), .dout(n15634));
  jand g15443(.dina(n15594), .dinb(n15592), .dout(n15635));
  jor  g15444(.dina(n15635), .dinb(n15634), .dout(n15636));
  jand g15445(.dina(\a[62] ), .dinb(\a[53] ), .dout(n15637));
  jand g15446(.dina(\a[58] ), .dinb(n15585), .dout(n15638));
  jxor g15447(.dina(n15638), .dinb(n15637), .dout(n15639));
  jnot g15448(.din(n15639), .dout(n15640));
  jand g15449(.dina(\a[61] ), .dinb(\a[54] ), .dout(n15641));
  jnot g15450(.din(n15641), .dout(n15642));
  jand g15451(.dina(\a[60] ), .dinb(\a[56] ), .dout(n15643));
  jand g15452(.dina(n15643), .dinb(n15559), .dout(n15644));
  jnot g15453(.din(n15644), .dout(n15645));
  jand g15454(.dina(\a[60] ), .dinb(\a[55] ), .dout(n15646));
  jor  g15455(.dina(n15646), .dinb(n14039), .dout(n15647));
  jand g15456(.dina(n15647), .dinb(n15645), .dout(n15648));
  jxor g15457(.dina(n15648), .dinb(n15642), .dout(n15649));
  jxor g15458(.dina(n15649), .dinb(n15640), .dout(n15650));
  jxor g15459(.dina(n15650), .dinb(n15636), .dout(n15651));
  jand g15460(.dina(n15609), .dinb(n15604), .dout(n15652));
  jor  g15461(.dina(n15652), .dinb(n15607), .dout(n15653));
  jand g15462(.dina(\a[63] ), .dinb(\a[52] ), .dout(n15654));
  jnot g15463(.din(n15612), .dout(n15655));
  jnot g15464(.din(n15613), .dout(n15656));
  jand g15465(.dina(n15656), .dinb(n15655), .dout(n15657));
  jor  g15466(.dina(n15657), .dinb(n15616), .dout(n15658));
  jnot g15467(.din(n15658), .dout(n15659));
  jxor g15468(.dina(n15659), .dinb(n15654), .dout(n15660));
  jxor g15469(.dina(n15660), .dinb(n15653), .dout(n15661));
  jnot g15470(.din(n15661), .dout(n15662));
  jor  g15471(.dina(n15618), .dinb(n15611), .dout(n15663));
  jand g15472(.dina(n15619), .dinb(n15603), .dout(n15664));
  jnot g15473(.din(n15664), .dout(n15665));
  jand g15474(.dina(n15665), .dinb(n15663), .dout(n15666));
  jxor g15475(.dina(n15666), .dinb(n15662), .dout(n15667));
  jxor g15476(.dina(n15667), .dinb(n15651), .dout(n15668));
  jand g15477(.dina(n15668), .dinb(n15633), .dout(n15669));
  jor  g15478(.dina(n15668), .dinb(n15633), .dout(n15670));
  jnot g15479(.din(n15670), .dout(n15671));
  jor  g15480(.dina(n15671), .dinb(n15669), .dout(n15672));
  jand g15481(.dina(n15621), .dinb(n15584), .dout(n15673));
  jnot g15482(.din(n15673), .dout(n15674));
  jnot g15483(.din(n15584), .dout(n15675));
  jand g15484(.dina(n15622), .dinb(n15675), .dout(n15676));
  jor  g15485(.dina(n15629), .dinb(n15676), .dout(n15677));
  jand g15486(.dina(n15677), .dinb(n15674), .dout(n15678));
  jxor g15487(.dina(n15678), .dinb(n15672), .dout(\asquared[116] ));
  jor  g15488(.dina(n15649), .dinb(n15640), .dout(n15680));
  jand g15489(.dina(n15650), .dinb(n15636), .dout(n15681));
  jnot g15490(.din(n15681), .dout(n15682));
  jand g15491(.dina(n15682), .dinb(n15680), .dout(n15683));
  jnot g15492(.din(n15683), .dout(n15684));
  jand g15493(.dina(n15659), .dinb(n15654), .dout(n15685));
  jand g15494(.dina(n15660), .dinb(n15653), .dout(n15686));
  jor  g15495(.dina(n15686), .dinb(n15685), .dout(n15687));
  jxor g15496(.dina(n15687), .dinb(n15684), .dout(n15688));
  jand g15497(.dina(\a[63] ), .dinb(\a[54] ), .dout(n15689));
  jand g15498(.dina(n15689), .dinb(n15637), .dout(n15690));
  jnot g15499(.din(n15690), .dout(n15691));
  jand g15500(.dina(\a[62] ), .dinb(\a[54] ), .dout(n15692));
  jand g15501(.dina(\a[63] ), .dinb(\a[53] ), .dout(n15693));
  jor  g15502(.dina(n15693), .dinb(n15692), .dout(n15694));
  jand g15503(.dina(n15694), .dinb(n15691), .dout(n15695));
  jor  g15504(.dina(n15637), .dinb(\a[57] ), .dout(n15696));
  jand g15505(.dina(n15696), .dinb(\a[58] ), .dout(n15697));
  jxor g15506(.dina(n15697), .dinb(n15695), .dout(n15698));
  jand g15507(.dina(n15645), .dinb(n15642), .dout(n15699));
  jnot g15508(.din(n15699), .dout(n15700));
  jand g15509(.dina(n15700), .dinb(n15647), .dout(n15701));
  jnot g15510(.din(n15701), .dout(n15702));
  jand g15511(.dina(\a[61] ), .dinb(\a[55] ), .dout(n15703));
  jnot g15512(.din(n15703), .dout(n15704));
  jand g15513(.dina(\a[60] ), .dinb(\a[57] ), .dout(n15705));
  jand g15514(.dina(n15705), .dinb(n14039), .dout(n15706));
  jnot g15515(.din(n15706), .dout(n15707));
  jor  g15516(.dina(n15643), .dinb(n11144), .dout(n15708));
  jand g15517(.dina(n15708), .dinb(n15707), .dout(n15709));
  jxor g15518(.dina(n15709), .dinb(n15704), .dout(n15710));
  jxor g15519(.dina(n15710), .dinb(n15702), .dout(n15711));
  jxor g15520(.dina(n15711), .dinb(n15698), .dout(n15712));
  jxor g15521(.dina(n15712), .dinb(n15688), .dout(n15713));
  jor  g15522(.dina(n15666), .dinb(n15662), .dout(n15714));
  jand g15523(.dina(n15667), .dinb(n15651), .dout(n15715));
  jnot g15524(.din(n15715), .dout(n15716));
  jand g15525(.dina(n15716), .dinb(n15714), .dout(n15717));
  jxor g15526(.dina(n15717), .dinb(n15713), .dout(n15718));
  jnot g15527(.din(n15669), .dout(n15719));
  jor  g15528(.dina(n15678), .dinb(n15671), .dout(n15720));
  jand g15529(.dina(n15720), .dinb(n15719), .dout(n15721));
  jxor g15530(.dina(n15721), .dinb(n15718), .dout(\asquared[117] ));
  jand g15531(.dina(n15687), .dinb(n15684), .dout(n15723));
  jand g15532(.dina(n15712), .dinb(n15688), .dout(n15724));
  jor  g15533(.dina(n15724), .dinb(n15723), .dout(n15725));
  jand g15534(.dina(n15697), .dinb(n15695), .dout(n15726));
  jor  g15535(.dina(n15726), .dinb(n15690), .dout(n15727));
  jand g15536(.dina(n15707), .dinb(n15704), .dout(n15728));
  jnot g15537(.din(n15728), .dout(n15729));
  jand g15538(.dina(n15729), .dinb(n15708), .dout(n15730));
  jxor g15539(.dina(n15730), .dinb(n15727), .dout(n15731));
  jnot g15540(.din(n15731), .dout(n15732));
  jand g15541(.dina(\a[61] ), .dinb(\a[57] ), .dout(n15733));
  jand g15542(.dina(n15733), .dinb(n15643), .dout(n15734));
  jnot g15543(.din(n15705), .dout(n15735));
  jand g15544(.dina(\a[61] ), .dinb(\a[56] ), .dout(n15736));
  jnot g15545(.din(n15736), .dout(n15737));
  jand g15546(.dina(n15737), .dinb(n15735), .dout(n15738));
  jor  g15547(.dina(n15738), .dinb(n15734), .dout(n15739));
  jxor g15548(.dina(n15739), .dinb(n15689), .dout(n15740));
  jxor g15549(.dina(n15740), .dinb(n15732), .dout(n15741));
  jor  g15550(.dina(n15710), .dinb(n15702), .dout(n15742));
  jand g15551(.dina(n15711), .dinb(n15698), .dout(n15743));
  jnot g15552(.din(n15743), .dout(n15744));
  jand g15553(.dina(n15744), .dinb(n15742), .dout(n15745));
  jand g15554(.dina(\a[62] ), .dinb(\a[55] ), .dout(n15746));
  jnot g15555(.din(n15746), .dout(n15747));
  jnot g15556(.din(\a[58] ), .dout(n15748));
  jand g15557(.dina(\a[59] ), .dinb(n15748), .dout(n15749));
  jxor g15558(.dina(n15749), .dinb(n15747), .dout(n15750));
  jxor g15559(.dina(n15750), .dinb(n15745), .dout(n15751));
  jxor g15560(.dina(n15751), .dinb(n15741), .dout(n15752));
  jand g15561(.dina(n15752), .dinb(n15725), .dout(n15753));
  jor  g15562(.dina(n15752), .dinb(n15725), .dout(n15754));
  jnot g15563(.din(n15754), .dout(n15755));
  jor  g15564(.dina(n15755), .dinb(n15753), .dout(n15756));
  jnot g15565(.din(n15713), .dout(n15757));
  jor  g15566(.dina(n15717), .dinb(n15757), .dout(n15758));
  jand g15567(.dina(n15717), .dinb(n15757), .dout(n15759));
  jor  g15568(.dina(n15721), .dinb(n15759), .dout(n15760));
  jand g15569(.dina(n15760), .dinb(n15758), .dout(n15761));
  jxor g15570(.dina(n15761), .dinb(n15756), .dout(\asquared[118] ));
  jand g15571(.dina(\a[63] ), .dinb(\a[55] ), .dout(n15763));
  jnot g15572(.din(\a[59] ), .dout(n15764));
  jand g15573(.dina(n15747), .dinb(n15748), .dout(n15765));
  jor  g15574(.dina(n15765), .dinb(n15764), .dout(n15766));
  jnot g15575(.din(n15766), .dout(n15767));
  jxor g15576(.dina(n15767), .dinb(n15763), .dout(n15768));
  jnot g15577(.din(n15689), .dout(n15769));
  jnot g15578(.din(n15734), .dout(n15770));
  jand g15579(.dina(n15770), .dinb(n15769), .dout(n15771));
  jor  g15580(.dina(n15771), .dinb(n15738), .dout(n15772));
  jnot g15581(.din(n15772), .dout(n15773));
  jxor g15582(.dina(n15773), .dinb(n15768), .dout(n15774));
  jand g15583(.dina(n15730), .dinb(n15727), .dout(n15775));
  jnot g15584(.din(n15775), .dout(n15776));
  jor  g15585(.dina(n15740), .dinb(n15732), .dout(n15777));
  jand g15586(.dina(n15777), .dinb(n15776), .dout(n15778));
  jnot g15587(.din(n15778), .dout(n15779));
  jand g15588(.dina(\a[62] ), .dinb(\a[56] ), .dout(n15780));
  jand g15589(.dina(\a[61] ), .dinb(\a[58] ), .dout(n15781));
  jand g15590(.dina(n15781), .dinb(n15705), .dout(n15782));
  jnot g15591(.din(n15782), .dout(n15783));
  jand g15592(.dina(\a[60] ), .dinb(\a[58] ), .dout(n15784));
  jand g15593(.dina(n15784), .dinb(n15780), .dout(n15785));
  jand g15594(.dina(\a[62] ), .dinb(\a[57] ), .dout(n15786));
  jand g15595(.dina(n15786), .dinb(n15736), .dout(n15787));
  jor  g15596(.dina(n15787), .dinb(n15785), .dout(n15788));
  jand g15597(.dina(n15788), .dinb(n15783), .dout(n15789));
  jnot g15598(.din(n15789), .dout(n15790));
  jand g15599(.dina(n15790), .dinb(n15780), .dout(n15791));
  jor  g15600(.dina(n15788), .dinb(n15782), .dout(n15792));
  jnot g15601(.din(n15792), .dout(n15793));
  jor  g15602(.dina(n15784), .dinb(n15733), .dout(n15794));
  jand g15603(.dina(n15794), .dinb(n15793), .dout(n15795));
  jor  g15604(.dina(n15795), .dinb(n15791), .dout(n15796));
  jxor g15605(.dina(n15796), .dinb(n15779), .dout(n15797));
  jxor g15606(.dina(n15797), .dinb(n15774), .dout(n15798));
  jor  g15607(.dina(n15750), .dinb(n15745), .dout(n15799));
  jand g15608(.dina(n15751), .dinb(n15741), .dout(n15800));
  jnot g15609(.din(n15800), .dout(n15801));
  jand g15610(.dina(n15801), .dinb(n15799), .dout(n15802));
  jxor g15611(.dina(n15802), .dinb(n15798), .dout(n15803));
  jnot g15612(.din(n15753), .dout(n15804));
  jor  g15613(.dina(n15761), .dinb(n15755), .dout(n15805));
  jand g15614(.dina(n15805), .dinb(n15804), .dout(n15806));
  jxor g15615(.dina(n15806), .dinb(n15803), .dout(\asquared[119] ));
  jand g15616(.dina(n15767), .dinb(n15763), .dout(n15808));
  jand g15617(.dina(n15773), .dinb(n15768), .dout(n15809));
  jor  g15618(.dina(n15809), .dinb(n15808), .dout(n15810));
  jand g15619(.dina(n11688), .dinb(n8387), .dout(n15811));
  jnot g15620(.din(n15811), .dout(n15812));
  jand g15621(.dina(\a[63] ), .dinb(\a[56] ), .dout(n15813));
  jor  g15622(.dina(n15813), .dinb(n15781), .dout(n15814));
  jand g15623(.dina(n15814), .dinb(n15812), .dout(n15815));
  jxor g15624(.dina(n15815), .dinb(n15792), .dout(n15816));
  jnot g15625(.din(n15816), .dout(n15817));
  jnot g15626(.din(n15786), .dout(n15818));
  jand g15627(.dina(\a[60] ), .dinb(n15764), .dout(n15819));
  jxor g15628(.dina(n15819), .dinb(n15818), .dout(n15820));
  jxor g15629(.dina(n15820), .dinb(n15817), .dout(n15821));
  jxor g15630(.dina(n15821), .dinb(n15810), .dout(n15822));
  jand g15631(.dina(n15796), .dinb(n15779), .dout(n15823));
  jand g15632(.dina(n15797), .dinb(n15774), .dout(n15824));
  jor  g15633(.dina(n15824), .dinb(n15823), .dout(n15825));
  jand g15634(.dina(n15825), .dinb(n15822), .dout(n15826));
  jor  g15635(.dina(n15825), .dinb(n15822), .dout(n15827));
  jnot g15636(.din(n15827), .dout(n15828));
  jor  g15637(.dina(n15828), .dinb(n15826), .dout(n15829));
  jnot g15638(.din(n15798), .dout(n15830));
  jor  g15639(.dina(n15802), .dinb(n15830), .dout(n15831));
  jand g15640(.dina(n15802), .dinb(n15830), .dout(n15832));
  jor  g15641(.dina(n15806), .dinb(n15832), .dout(n15833));
  jand g15642(.dina(n15833), .dinb(n15831), .dout(n15834));
  jxor g15643(.dina(n15834), .dinb(n15829), .dout(\asquared[120] ));
  jor  g15644(.dina(n15820), .dinb(n15817), .dout(n15836));
  jand g15645(.dina(n15821), .dinb(n15810), .dout(n15837));
  jnot g15646(.din(n15837), .dout(n15838));
  jand g15647(.dina(n15838), .dinb(n15836), .dout(n15839));
  jand g15648(.dina(n15815), .dinb(n15792), .dout(n15840));
  jor  g15649(.dina(n15840), .dinb(n15811), .dout(n15841));
  jnot g15650(.din(\a[60] ), .dout(n15842));
  jand g15651(.dina(n15818), .dinb(n15764), .dout(n15843));
  jor  g15652(.dina(n15843), .dinb(n15842), .dout(n15844));
  jnot g15653(.din(n15844), .dout(n15845));
  jxor g15654(.dina(n15845), .dinb(n15841), .dout(n15846));
  jnot g15655(.din(n15846), .dout(n15847));
  jand g15656(.dina(\a[63] ), .dinb(\a[57] ), .dout(n15848));
  jnot g15657(.din(n15848), .dout(n15849));
  jand g15658(.dina(\a[62] ), .dinb(\a[59] ), .dout(n15850));
  jand g15659(.dina(n15850), .dinb(n15781), .dout(n15851));
  jnot g15660(.din(n15851), .dout(n15852));
  jand g15661(.dina(\a[62] ), .dinb(\a[58] ), .dout(n15853));
  jor  g15662(.dina(n15853), .dinb(n13790), .dout(n15854));
  jand g15663(.dina(n15854), .dinb(n15852), .dout(n15855));
  jxor g15664(.dina(n15855), .dinb(n15849), .dout(n15856));
  jxor g15665(.dina(n15856), .dinb(n15847), .dout(n15857));
  jxor g15666(.dina(n15857), .dinb(n15839), .dout(n15858));
  jnot g15667(.din(n15826), .dout(n15859));
  jor  g15668(.dina(n15834), .dinb(n15828), .dout(n15860));
  jand g15669(.dina(n15860), .dinb(n15859), .dout(n15861));
  jxor g15670(.dina(n15861), .dinb(n15858), .dout(\asquared[121] ));
  jand g15671(.dina(n15852), .dinb(n15849), .dout(n15863));
  jnot g15672(.din(n15863), .dout(n15864));
  jand g15673(.dina(n15864), .dinb(n15854), .dout(n15865));
  jxor g15674(.dina(n15865), .dinb(n15115), .dout(n15866));
  jnot g15675(.din(n15866), .dout(n15867));
  jnot g15676(.din(n15850), .dout(n15868));
  jand g15677(.dina(\a[61] ), .dinb(n15842), .dout(n15869));
  jxor g15678(.dina(n15869), .dinb(n15868), .dout(n15870));
  jxor g15679(.dina(n15870), .dinb(n15867), .dout(n15871));
  jand g15680(.dina(n15845), .dinb(n15841), .dout(n15872));
  jnot g15681(.din(n15872), .dout(n15873));
  jor  g15682(.dina(n15856), .dinb(n15847), .dout(n15874));
  jand g15683(.dina(n15874), .dinb(n15873), .dout(n15875));
  jxor g15684(.dina(n15875), .dinb(n15871), .dout(n15876));
  jnot g15685(.din(n15839), .dout(n15877));
  jand g15686(.dina(n15857), .dinb(n15877), .dout(n15878));
  jnot g15687(.din(n15878), .dout(n15879));
  jnot g15688(.din(n15857), .dout(n15880));
  jand g15689(.dina(n15880), .dinb(n15839), .dout(n15881));
  jor  g15690(.dina(n15861), .dinb(n15881), .dout(n15882));
  jand g15691(.dina(n15882), .dinb(n15879), .dout(n15883));
  jxor g15692(.dina(n15883), .dinb(n15876), .dout(\asquared[122] ));
  jand g15693(.dina(n15865), .dinb(n15115), .dout(n15885));
  jnot g15694(.din(n15885), .dout(n15886));
  jor  g15695(.dina(n15870), .dinb(n15867), .dout(n15887));
  jand g15696(.dina(n15887), .dinb(n15886), .dout(n15888));
  jnot g15697(.din(\a[61] ), .dout(n15889));
  jand g15698(.dina(n15868), .dinb(n15842), .dout(n15890));
  jor  g15699(.dina(n15890), .dinb(n15889), .dout(n15891));
  jnot g15700(.din(n15891), .dout(n15892));
  jand g15701(.dina(\a[63] ), .dinb(\a[59] ), .dout(n15893));
  jand g15702(.dina(\a[62] ), .dinb(\a[60] ), .dout(n15894));
  jor  g15703(.dina(n15894), .dinb(n15893), .dout(n15895));
  jand g15704(.dina(\a[63] ), .dinb(\a[60] ), .dout(n15896));
  jand g15705(.dina(n15896), .dinb(n15850), .dout(n15897));
  jnot g15706(.din(n15897), .dout(n15898));
  jand g15707(.dina(n15898), .dinb(n15895), .dout(n15899));
  jxor g15708(.dina(n15899), .dinb(n15892), .dout(n15900));
  jxor g15709(.dina(n15900), .dinb(n15888), .dout(n15901));
  jnot g15710(.din(n15871), .dout(n15902));
  jor  g15711(.dina(n15875), .dinb(n15902), .dout(n15903));
  jand g15712(.dina(n15875), .dinb(n15902), .dout(n15904));
  jor  g15713(.dina(n15883), .dinb(n15904), .dout(n15905));
  jand g15714(.dina(n15905), .dinb(n15903), .dout(n15906));
  jxor g15715(.dina(n15906), .dinb(n15901), .dout(\asquared[123] ));
  jand g15716(.dina(n15895), .dinb(n15892), .dout(n15908));
  jor  g15717(.dina(n15908), .dinb(n15897), .dout(n15909));
  jand g15718(.dina(\a[62] ), .dinb(n15889), .dout(n15910));
  jxor g15719(.dina(n15910), .dinb(n15896), .dout(n15911));
  jnot g15720(.din(n15911), .dout(n15912));
  jxor g15721(.dina(n15912), .dinb(n15909), .dout(n15913));
  jnot g15722(.din(n15900), .dout(n15914));
  jor  g15723(.dina(n15914), .dinb(n15888), .dout(n15915));
  jand g15724(.dina(n15914), .dinb(n15888), .dout(n15916));
  jor  g15725(.dina(n15906), .dinb(n15916), .dout(n15917));
  jand g15726(.dina(n15917), .dinb(n15915), .dout(n15918));
  jxor g15727(.dina(n15918), .dinb(n15913), .dout(\asquared[124] ));
  jand g15728(.dina(n15911), .dinb(n15909), .dout(n15920));
  jnot g15729(.din(n15920), .dout(n15921));
  jnot g15730(.din(n15909), .dout(n15922));
  jand g15731(.dina(n15912), .dinb(n15922), .dout(n15923));
  jor  g15732(.dina(n15918), .dinb(n15923), .dout(n15924));
  jand g15733(.dina(n15924), .dinb(n15921), .dout(n15925));
  jand g15734(.dina(n15910), .dinb(n15896), .dout(n15926));
  jor  g15735(.dina(n15926), .dinb(n8387), .dout(n15927));
  jor  g15736(.dina(n15927), .dinb(n8702), .dout(n15928));
  jnot g15737(.din(n15928), .dout(n15929));
  jand g15738(.dina(n8387), .dinb(\a[62] ), .dout(n15930));
  jor  g15739(.dina(n15930), .dinb(n15929), .dout(n15931));
  jxor g15740(.dina(n15931), .dinb(n15925), .dout(\asquared[125] ));
  jnot g15741(.din(n15923), .dout(n15933));
  jnot g15742(.din(n15915), .dout(n15934));
  jnot g15743(.din(n15916), .dout(n15935));
  jnot g15744(.din(n15903), .dout(n15936));
  jnot g15745(.din(n15904), .dout(n15937));
  jnot g15746(.din(n15881), .dout(n15938));
  jnot g15747(.din(n15831), .dout(n15939));
  jnot g15748(.din(n15832), .dout(n15940));
  jnot g15749(.din(n15758), .dout(n15941));
  jnot g15750(.din(n15759), .dout(n15942));
  jnot g15751(.din(n15676), .dout(n15943));
  jnot g15752(.din(n15627), .dout(n15944));
  jnot g15753(.din(n15578), .dout(n15945));
  jnot g15754(.din(n15457), .dout(n15946));
  jnot g15755(.din(n15458), .dout(n15947));
  jnot g15756(.din(n15327), .dout(n15948));
  jnot g15757(.din(n15253), .dout(n15949));
  jnot g15758(.din(n15098), .dout(n15950));
  jnot g15759(.din(n14836), .dout(n15951));
  jnot g15760(.din(n14417), .dout(n15952));
  jnot g15761(.din(n14180), .dout(n15953));
  jnot g15762(.din(n13933), .dout(n15954));
  jnot g15763(.din(n13689), .dout(n15955));
  jnot g15764(.din(n13414), .dout(n15956));
  jnot g15765(.din(n13139), .dout(n15957));
  jnot g15766(.din(n13140), .dout(n15958));
  jnot g15767(.din(n12995), .dout(n15959));
  jnot g15768(.din(n12848), .dout(n15960));
  jnot g15769(.din(n11857), .dout(n15961));
  jnot g15770(.din(n10747), .dout(n15962));
  jnot g15771(.din(n10543), .dout(n15963));
  jnot g15772(.din(n10345), .dout(n15964));
  jnot g15773(.din(n10139), .dout(n15965));
  jnot g15774(.din(n9935), .dout(n15966));
  jnot g15775(.din(n9492), .dout(n15967));
  jnot g15776(.din(n8580), .dout(n15968));
  jnot g15777(.din(n8325), .dout(n15969));
  jnot g15778(.din(n7588), .dout(n15970));
  jnot g15779(.din(n7325), .dout(n15971));
  jnot g15780(.din(n5790), .dout(n15972));
  jnot g15781(.din(n5364), .dout(n15973));
  jnot g15782(.din(n5158), .dout(n15974));
  jnot g15783(.din(n4960), .dout(n15975));
  jnot g15784(.din(n4591), .dout(n15976));
  jnot g15785(.din(n3699), .dout(n15977));
  jnot g15786(.din(n2897), .dout(n15978));
  jnot g15787(.din(n2742), .dout(n15979));
  jnot g15788(.din(n2468), .dout(n15980));
  jnot g15789(.din(n1862), .dout(n15981));
  jnot g15790(.din(n1529), .dout(n15982));
  jnot g15791(.din(n1343), .dout(n15983));
  jnot g15792(.din(n1002), .dout(n15984));
  jnot g15793(.din(n589), .dout(n15985));
  jnot g15794(.din(n532), .dout(n15986));
  jnot g15795(.din(n472), .dout(n15987));
  jnot g15796(.din(n421), .dout(n15988));
  jnot g15797(.din(n321), .dout(n15989));
  jor  g15798(.dina(n228), .dinb(n218), .dout(n15990));
  jand g15799(.dina(n214), .dinb(n195), .dout(n15991));
  jor  g15800(.dina(n214), .dinb(n195), .dout(n15992));
  jand g15801(.dina(n15992), .dinb(n204), .dout(n15993));
  jor  g15802(.dina(n15993), .dinb(n15991), .dout(n15994));
  jand g15803(.dina(n15994), .dinb(n15990), .dout(n15995));
  jor  g15804(.dina(n15995), .dinb(n256), .dout(n15996));
  jand g15805(.dina(n15996), .dinb(n252), .dout(n15997));
  jor  g15806(.dina(n15997), .dinb(n254), .dout(n15998));
  jand g15807(.dina(n15998), .dinb(n15989), .dout(n15999));
  jor  g15808(.dina(n15999), .dinb(n318), .dout(n16000));
  jand g15809(.dina(n16000), .dinb(n314), .dout(n16001));
  jor  g15810(.dina(n16001), .dinb(n316), .dout(n16002));
  jand g15811(.dina(n16002), .dinb(n349), .dout(n16003));
  jor  g15812(.dina(n16003), .dinb(n348), .dout(n16004));
  jand g15813(.dina(n16004), .dinb(n15988), .dout(n16005));
  jor  g15814(.dina(n16005), .dinb(n418), .dout(n16006));
  jand g15815(.dina(n16006), .dinb(n15987), .dout(n16007));
  jor  g15816(.dina(n16007), .dinb(n469), .dout(n16008));
  jand g15817(.dina(n16008), .dinb(n15986), .dout(n16009));
  jor  g15818(.dina(n16009), .dinb(n529), .dout(n16010));
  jand g15819(.dina(n16010), .dinb(n15985), .dout(n16011));
  jor  g15820(.dina(n16011), .dinb(n586), .dout(n16012));
  jand g15821(.dina(n16012), .dinb(n583), .dout(n16013));
  jor  g15822(.dina(n16013), .dinb(n582), .dout(n16014));
  jand g15823(.dina(n16014), .dinb(n629), .dout(n16015));
  jor  g15824(.dina(n16015), .dinb(n628), .dout(n16016));
  jand g15825(.dina(n16016), .dinb(n696), .dout(n16017));
  jor  g15826(.dina(n16017), .dinb(n695), .dout(n16018));
  jand g15827(.dina(n16018), .dinb(n758), .dout(n16019));
  jor  g15828(.dina(n16019), .dinb(n757), .dout(n16020));
  jand g15829(.dina(n16020), .dinb(n843), .dout(n16021));
  jor  g15830(.dina(n16021), .dinb(n842), .dout(n16022));
  jand g15831(.dina(n16022), .dinb(n15984), .dout(n16023));
  jor  g15832(.dina(n16023), .dinb(n999), .dout(n16024));
  jand g15833(.dina(n16024), .dinb(n1082), .dout(n16025));
  jor  g15834(.dina(n16025), .dinb(n1080), .dout(n16026));
  jand g15835(.dina(n16026), .dinb(n1076), .dout(n16027));
  jor  g15836(.dina(n16027), .dinb(n1075), .dout(n16028));
  jand g15837(.dina(n16028), .dinb(n1164), .dout(n16029));
  jor  g15838(.dina(n16029), .dinb(n1163), .dout(n16030));
  jand g15839(.dina(n16030), .dinb(n15983), .dout(n16031));
  jor  g15840(.dina(n16031), .dinb(n1340), .dout(n16032));
  jand g15841(.dina(n16032), .dinb(n1337), .dout(n16033));
  jor  g15842(.dina(n16033), .dinb(n1336), .dout(n16034));
  jand g15843(.dina(n16034), .dinb(n15982), .dout(n16035));
  jor  g15844(.dina(n16035), .dinb(n1526), .dout(n16036));
  jand g15845(.dina(n16036), .dinb(n1523), .dout(n16037));
  jor  g15846(.dina(n16037), .dinb(n1522), .dout(n16038));
  jand g15847(.dina(n16038), .dinb(n1632), .dout(n16039));
  jor  g15848(.dina(n16039), .dinb(n1631), .dout(n16040));
  jand g15849(.dina(n16040), .dinb(n15981), .dout(n16041));
  jor  g15850(.dina(n16041), .dinb(n1859), .dout(n16042));
  jand g15851(.dina(n16042), .dinb(n1856), .dout(n16043));
  jor  g15852(.dina(n16043), .dinb(n1855), .dout(n16044));
  jand g15853(.dina(n16044), .dinb(n1971), .dout(n16045));
  jor  g15854(.dina(n16045), .dinb(n1970), .dout(n16046));
  jand g15855(.dina(n16046), .dinb(n2098), .dout(n16047));
  jor  g15856(.dina(n16047), .dinb(n2097), .dout(n16048));
  jand g15857(.dina(n16048), .dinb(n2209), .dout(n16049));
  jor  g15858(.dina(n16049), .dinb(n2208), .dout(n16050));
  jand g15859(.dina(n16050), .dinb(n15980), .dout(n16051));
  jor  g15860(.dina(n16051), .dinb(n2465), .dout(n16052));
  jand g15861(.dina(n16052), .dinb(n2462), .dout(n16053));
  jor  g15862(.dina(n16053), .dinb(n2461), .dout(n16054));
  jand g15863(.dina(n16054), .dinb(n15979), .dout(n16055));
  jor  g15864(.dina(n16055), .dinb(n2739), .dout(n16056));
  jand g15865(.dina(n16056), .dinb(n15978), .dout(n16057));
  jor  g15866(.dina(n16057), .dinb(n2894), .dout(n16058));
  jand g15867(.dina(n16058), .dinb(n2891), .dout(n16059));
  jor  g15868(.dina(n16059), .dinb(n2890), .dout(n16060));
  jand g15869(.dina(n16060), .dinb(n3059), .dout(n16061));
  jor  g15870(.dina(n16061), .dinb(n3058), .dout(n16062));
  jand g15871(.dina(n16062), .dinb(n3220), .dout(n16063));
  jor  g15872(.dina(n16063), .dinb(n3219), .dout(n16064));
  jand g15873(.dina(n16064), .dinb(n3376), .dout(n16065));
  jor  g15874(.dina(n16065), .dinb(n3375), .dout(n16066));
  jand g15875(.dina(n16066), .dinb(n15977), .dout(n16067));
  jor  g15876(.dina(n16067), .dinb(n3696), .dout(n16068));
  jand g15877(.dina(n16068), .dinb(n3693), .dout(n16069));
  jor  g15878(.dina(n16069), .dinb(n3692), .dout(n16070));
  jand g15879(.dina(n16070), .dinb(n3868), .dout(n16071));
  jor  g15880(.dina(n16071), .dinb(n3867), .dout(n16072));
  jand g15881(.dina(n16072), .dinb(n4032), .dout(n16073));
  jor  g15882(.dina(n16073), .dinb(n4031), .dout(n16074));
  jand g15883(.dina(n16074), .dinb(n4213), .dout(n16075));
  jor  g15884(.dina(n16075), .dinb(n4212), .dout(n16076));
  jand g15885(.dina(n16076), .dinb(n15976), .dout(n16077));
  jor  g15886(.dina(n16077), .dinb(n4588), .dout(n16078));
  jand g15887(.dina(n16078), .dinb(n4585), .dout(n16079));
  jor  g15888(.dina(n16079), .dinb(n4584), .dout(n16080));
  jand g15889(.dina(n16080), .dinb(n15975), .dout(n16081));
  jor  g15890(.dina(n16081), .dinb(n4957), .dout(n16082));
  jand g15891(.dina(n16082), .dinb(n15974), .dout(n16083));
  jor  g15892(.dina(n16083), .dinb(n5155), .dout(n16084));
  jand g15893(.dina(n16084), .dinb(n15973), .dout(n16085));
  jor  g15894(.dina(n16085), .dinb(n5361), .dout(n16086));
  jand g15895(.dina(n16086), .dinb(n5358), .dout(n16087));
  jor  g15896(.dina(n16087), .dinb(n5357), .dout(n16088));
  jand g15897(.dina(n16088), .dinb(n15972), .dout(n16089));
  jor  g15898(.dina(n16089), .dinb(n5787), .dout(n16090));
  jand g15899(.dina(n16090), .dinb(n5784), .dout(n16091));
  jor  g15900(.dina(n16091), .dinb(n5783), .dout(n16092));
  jand g15901(.dina(n16092), .dinb(n6006), .dout(n16093));
  jor  g15902(.dina(n16093), .dinb(n6005), .dout(n16094));
  jand g15903(.dina(n16094), .dinb(n6210), .dout(n16095));
  jor  g15904(.dina(n16095), .dinb(n6209), .dout(n16096));
  jand g15905(.dina(n16096), .dinb(n6434), .dout(n16097));
  jor  g15906(.dina(n16097), .dinb(n6433), .dout(n16098));
  jand g15907(.dina(n16098), .dinb(n6656), .dout(n16099));
  jor  g15908(.dina(n16099), .dinb(n6655), .dout(n16100));
  jand g15909(.dina(n16100), .dinb(n6869), .dout(n16101));
  jor  g15910(.dina(n16101), .dinb(n6868), .dout(n16102));
  jand g15911(.dina(n16102), .dinb(n15971), .dout(n16103));
  jor  g15912(.dina(n16103), .dinb(n7322), .dout(n16104));
  jand g15913(.dina(n16104), .dinb(n15970), .dout(n16105));
  jor  g15914(.dina(n16105), .dinb(n7585), .dout(n16106));
  jand g15915(.dina(n16106), .dinb(n7582), .dout(n16107));
  jor  g15916(.dina(n16107), .dinb(n7581), .dout(n16108));
  jand g15917(.dina(n16108), .dinb(n7828), .dout(n16109));
  jor  g15918(.dina(n16109), .dinb(n7827), .dout(n16110));
  jand g15919(.dina(n16110), .dinb(n15969), .dout(n16111));
  jor  g15920(.dina(n16111), .dinb(n8322), .dout(n16112));
  jand g15921(.dina(n16112), .dinb(n15968), .dout(n16113));
  jor  g15922(.dina(n16113), .dinb(n8577), .dout(n16114));
  jand g15923(.dina(n16114), .dinb(n8574), .dout(n16115));
  jor  g15924(.dina(n16115), .dinb(n8573), .dout(n16116));
  jand g15925(.dina(n16116), .dinb(n8805), .dout(n16117));
  jor  g15926(.dina(n16117), .dinb(n8804), .dout(n16118));
  jand g15927(.dina(n16118), .dinb(n9046), .dout(n16119));
  jor  g15928(.dina(n16119), .dinb(n9045), .dout(n16120));
  jand g15929(.dina(n16120), .dinb(n15967), .dout(n16121));
  jor  g15930(.dina(n16121), .dinb(n9489), .dout(n16122));
  jand g15931(.dina(n16122), .dinb(n9486), .dout(n16123));
  jor  g15932(.dina(n16123), .dinb(n9485), .dout(n16124));
  jand g15933(.dina(n16124), .dinb(n15966), .dout(n16125));
  jor  g15934(.dina(n16125), .dinb(n9932), .dout(n16126));
  jand g15935(.dina(n16126), .dinb(n15965), .dout(n16127));
  jor  g15936(.dina(n16127), .dinb(n10136), .dout(n16128));
  jand g15937(.dina(n16128), .dinb(n15964), .dout(n16129));
  jor  g15938(.dina(n16129), .dinb(n10342), .dout(n16130));
  jand g15939(.dina(n16130), .dinb(n15963), .dout(n16131));
  jor  g15940(.dina(n16131), .dinb(n10540), .dout(n16132));
  jand g15941(.dina(n16132), .dinb(n15962), .dout(n16133));
  jor  g15942(.dina(n16133), .dinb(n10744), .dout(n16134));
  jand g15943(.dina(n16134), .dinb(n10741), .dout(n16135));
  jor  g15944(.dina(n16135), .dinb(n10740), .dout(n16136));
  jand g15945(.dina(n16136), .dinb(n10927), .dout(n16137));
  jor  g15946(.dina(n16137), .dinb(n10926), .dout(n16138));
  jand g15947(.dina(n16138), .dinb(n11124), .dout(n16139));
  jor  g15948(.dina(n16139), .dinb(n11123), .dout(n16140));
  jand g15949(.dina(n16140), .dinb(n11314), .dout(n16141));
  jor  g15950(.dina(n16141), .dinb(n11313), .dout(n16142));
  jand g15951(.dina(n16142), .dinb(n11495), .dout(n16143));
  jor  g15952(.dina(n16143), .dinb(n11494), .dout(n16144));
  jand g15953(.dina(n16144), .dinb(n15961), .dout(n16145));
  jor  g15954(.dina(n16145), .dinb(n11854), .dout(n16146));
  jand g15955(.dina(n16146), .dinb(n11851), .dout(n16147));
  jor  g15956(.dina(n16147), .dinb(n11850), .dout(n16148));
  jand g15957(.dina(n16148), .dinb(n12030), .dout(n16149));
  jor  g15958(.dina(n16149), .dinb(n12029), .dout(n16150));
  jand g15959(.dina(n16150), .dinb(n12205), .dout(n16151));
  jor  g15960(.dina(n16151), .dinb(n12204), .dout(n16152));
  jand g15961(.dina(n16152), .dinb(n12371), .dout(n16153));
  jor  g15962(.dina(n16153), .dinb(n12370), .dout(n16154));
  jand g15963(.dina(n16154), .dinb(n12525), .dout(n16155));
  jor  g15964(.dina(n16155), .dinb(n12524), .dout(n16156));
  jand g15965(.dina(n16156), .dinb(n15960), .dout(n16157));
  jor  g15966(.dina(n16157), .dinb(n12845), .dout(n16158));
  jand g15967(.dina(n16158), .dinb(n15959), .dout(n16159));
  jor  g15968(.dina(n16159), .dinb(n12992), .dout(n16160));
  jand g15969(.dina(n16160), .dinb(n15958), .dout(n16161));
  jor  g15970(.dina(n16161), .dinb(n15957), .dout(n16162));
  jand g15971(.dina(n16162), .dinb(n13135), .dout(n16163));
  jor  g15972(.dina(n16163), .dinb(n13134), .dout(n16164));
  jand g15973(.dina(n16164), .dinb(n15956), .dout(n16165));
  jor  g15974(.dina(n16165), .dinb(n13411), .dout(n16166));
  jand g15975(.dina(n16166), .dinb(n13408), .dout(n16167));
  jor  g15976(.dina(n16167), .dinb(n13407), .dout(n16168));
  jand g15977(.dina(n16168), .dinb(n15955), .dout(n16169));
  jor  g15978(.dina(n16169), .dinb(n13686), .dout(n16170));
  jand g15979(.dina(n16170), .dinb(n13683), .dout(n16171));
  jor  g15980(.dina(n16171), .dinb(n13682), .dout(n16172));
  jand g15981(.dina(n16172), .dinb(n15954), .dout(n16173));
  jor  g15982(.dina(n16173), .dinb(n13930), .dout(n16174));
  jand g15983(.dina(n16174), .dinb(n13927), .dout(n16175));
  jor  g15984(.dina(n16175), .dinb(n13926), .dout(n16176));
  jand g15985(.dina(n16176), .dinb(n15953), .dout(n16177));
  jor  g15986(.dina(n16177), .dinb(n14177), .dout(n16178));
  jand g15987(.dina(n16178), .dinb(n14174), .dout(n16179));
  jor  g15988(.dina(n16179), .dinb(n14173), .dout(n16180));
  jand g15989(.dina(n16180), .dinb(n15952), .dout(n16181));
  jor  g15990(.dina(n16181), .dinb(n14414), .dout(n16182));
  jand g15991(.dina(n16182), .dinb(n14411), .dout(n16183));
  jor  g15992(.dina(n16183), .dinb(n14410), .dout(n16184));
  jand g15993(.dina(n16184), .dinb(n14531), .dout(n16185));
  jor  g15994(.dina(n16185), .dinb(n14530), .dout(n16186));
  jand g15995(.dina(n16186), .dinb(n14636), .dout(n16187));
  jor  g15996(.dina(n16187), .dinb(n14635), .dout(n16188));
  jand g15997(.dina(n16188), .dinb(n15951), .dout(n16189));
  jor  g15998(.dina(n16189), .dinb(n14833), .dout(n16190));
  jand g15999(.dina(n16190), .dinb(n14830), .dout(n16191));
  jor  g16000(.dina(n16191), .dinb(n14829), .dout(n16192));
  jand g16001(.dina(n16192), .dinb(n14934), .dout(n16193));
  jor  g16002(.dina(n16193), .dinb(n14933), .dout(n16194));
  jand g16003(.dina(n16194), .dinb(n15950), .dout(n16195));
  jor  g16004(.dina(n16195), .dinb(n15095), .dout(n16196));
  jand g16005(.dina(n16196), .dinb(n15175), .dout(n16197));
  jor  g16006(.dina(n16197), .dinb(n15173), .dout(n16198));
  jand g16007(.dina(n16198), .dinb(n15949), .dout(n16199));
  jor  g16008(.dina(n16199), .dinb(n15250), .dout(n16200));
  jand g16009(.dina(n16200), .dinb(n15948), .dout(n16201));
  jor  g16010(.dina(n16201), .dinb(n15324), .dout(n16202));
  jand g16011(.dina(n16202), .dinb(n15321), .dout(n16203));
  jor  g16012(.dina(n16203), .dinb(n15320), .dout(n16204));
  jand g16013(.dina(n16204), .dinb(n15947), .dout(n16205));
  jor  g16014(.dina(n16205), .dinb(n15946), .dout(n16206));
  jand g16015(.dina(n16206), .dinb(n15525), .dout(n16207));
  jor  g16016(.dina(n16207), .dinb(n15523), .dout(n16208));
  jand g16017(.dina(n16208), .dinb(n15945), .dout(n16209));
  jor  g16018(.dina(n16209), .dinb(n15575), .dout(n16210));
  jand g16019(.dina(n16210), .dinb(n15944), .dout(n16211));
  jor  g16020(.dina(n16211), .dinb(n15624), .dout(n16212));
  jand g16021(.dina(n16212), .dinb(n15943), .dout(n16213));
  jor  g16022(.dina(n16213), .dinb(n15673), .dout(n16214));
  jand g16023(.dina(n16214), .dinb(n15670), .dout(n16215));
  jor  g16024(.dina(n16215), .dinb(n15669), .dout(n16216));
  jand g16025(.dina(n16216), .dinb(n15942), .dout(n16217));
  jor  g16026(.dina(n16217), .dinb(n15941), .dout(n16218));
  jand g16027(.dina(n16218), .dinb(n15754), .dout(n16219));
  jor  g16028(.dina(n16219), .dinb(n15753), .dout(n16220));
  jand g16029(.dina(n16220), .dinb(n15940), .dout(n16221));
  jor  g16030(.dina(n16221), .dinb(n15939), .dout(n16222));
  jand g16031(.dina(n16222), .dinb(n15827), .dout(n16223));
  jor  g16032(.dina(n16223), .dinb(n15826), .dout(n16224));
  jand g16033(.dina(n16224), .dinb(n15938), .dout(n16225));
  jor  g16034(.dina(n16225), .dinb(n15878), .dout(n16226));
  jand g16035(.dina(n16226), .dinb(n15937), .dout(n16227));
  jor  g16036(.dina(n16227), .dinb(n15936), .dout(n16228));
  jand g16037(.dina(n16228), .dinb(n15935), .dout(n16229));
  jor  g16038(.dina(n16229), .dinb(n15934), .dout(n16230));
  jand g16039(.dina(n16230), .dinb(n15933), .dout(n16231));
  jor  g16040(.dina(n16231), .dinb(n15920), .dout(n16232));
  jand g16041(.dina(n15928), .dinb(n16232), .dout(n16233));
  jnot g16042(.din(n15910), .dout(n16234));
  jand g16043(.dina(n16234), .dinb(\a[63] ), .dout(n16235));
  jor  g16044(.dina(n16235), .dinb(n16233), .dout(n16236));
  jor  g16045(.dina(n15929), .dinb(n15925), .dout(n16237));
  jor  g16046(.dina(n8123), .dinb(\a[62] ), .dout(n16238));
  jor  g16047(.dina(n16238), .dinb(n16237), .dout(n16239));
  jand g16048(.dina(n16239), .dinb(n16236), .dout(\asquared[126] ));
  jor  g16049(.dina(n16233), .dinb(\a[62] ), .dout(n16241));
  jand g16050(.dina(n16241), .dinb(\a[63] ), .dout(\asquared[127] ));
  buf  g16051(.din(\a[0] ), .dout(\asquared[0] ));
endmodule


