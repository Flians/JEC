module rf_c6288(G511gat, G154gat, G222gat, G256gat, G375gat, G137gat, G52gat, G35gat, G171gat, G69gat, G18gat, G86gat, G409gat, G443gat, G188gat, G1gat, G120gat, G494gat, G477gat, G205gat, G307gat, G239gat, G273gat, G290gat, G358gat, G324gat, G528gat, G341gat, G392gat, G426gat, G103gat, G460gat, G6287gat, G6280gat, G5308gat, G4591gat, G2877gat, G4946gat, G3895gat, G3552gat, G6250gat, G3211gat, G2548gat, G6270gat, G1901gat, G6170gat, G1581gat, G4241gat, G545gat, G5672gat, G6160gat, G5971gat, G6123gat, G6200gat, G6288gat, G6150gat, G2223gat, G6260gat, G6180gat, G6190gat, G6220gat, G6230gat, G6210gat, G6240gat);
    input G511gat, G154gat, G222gat, G256gat, G375gat, G137gat, G52gat, G35gat, G171gat, G69gat, G18gat, G86gat, G409gat, G443gat, G188gat, G1gat, G120gat, G494gat, G477gat, G205gat, G307gat, G239gat, G273gat, G290gat, G358gat, G324gat, G528gat, G341gat, G392gat, G426gat, G103gat, G460gat;
    output G6287gat, G6280gat, G5308gat, G4591gat, G2877gat, G4946gat, G3895gat, G3552gat, G6250gat, G3211gat, G2548gat, G6270gat, G1901gat, G6170gat, G1581gat, G4241gat, G545gat, G5672gat, G6160gat, G5971gat, G6123gat, G6200gat, G6288gat, G6150gat, G2223gat, G6260gat, G6180gat, G6190gat, G6220gat, G6230gat, G6210gat, G6240gat;
    wire n67;
    wire n71;
    wire n75;
    wire n79;
    wire n83;
    wire n87;
    wire n90;
    wire n94;
    wire n98;
    wire n101;
    wire n104;
    wire n107;
    wire n111;
    wire n114;
    wire n117;
    wire n121;
    wire n125;
    wire n129;
    wire n133;
    wire n137;
    wire n141;
    wire n144;
    wire n148;
    wire n152;
    wire n156;
    wire n160;
    wire n163;
    wire n166;
    wire n170;
    wire n174;
    wire n178;
    wire n181;
    wire n185;
    wire n189;
    wire n193;
    wire n197;
    wire n201;
    wire n204;
    wire n208;
    wire n212;
    wire n216;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n242;
    wire n245;
    wire n249;
    wire n253;
    wire n257;
    wire n261;
    wire n264;
    wire n268;
    wire n271;
    wire n275;
    wire n279;
    wire n283;
    wire n287;
    wire n291;
    wire n295;
    wire n299;
    wire n303;
    wire n306;
    wire n310;
    wire n314;
    wire n318;
    wire n322;
    wire n325;
    wire n329;
    wire n333;
    wire n337;
    wire n340;
    wire n344;
    wire n348;
    wire n351;
    wire n355;
    wire n359;
    wire n363;
    wire n367;
    wire n371;
    wire n374;
    wire n377;
    wire n381;
    wire n385;
    wire n389;
    wire n393;
    wire n396;
    wire n400;
    wire n404;
    wire n408;
    wire n412;
    wire n416;
    wire n419;
    wire n422;
    wire n426;
    wire n430;
    wire n434;
    wire n438;
    wire n442;
    wire n445;
    wire n449;
    wire n453;
    wire n457;
    wire n461;
    wire n464;
    wire n468;
    wire n472;
    wire n476;
    wire n480;
    wire n484;
    wire n488;
    wire n492;
    wire n495;
    wire n499;
    wire n503;
    wire n507;
    wire n511;
    wire n515;
    wire n518;
    wire n521;
    wire n525;
    wire n529;
    wire n533;
    wire n537;
    wire n540;
    wire n544;
    wire n548;
    wire n552;
    wire n556;
    wire n560;
    wire n563;
    wire n567;
    wire n571;
    wire n575;
    wire n579;
    wire n582;
    wire n585;
    wire n589;
    wire n593;
    wire n597;
    wire n600;
    wire n604;
    wire n608;
    wire n612;
    wire n616;
    wire n619;
    wire n623;
    wire n627;
    wire n631;
    wire n635;
    wire n639;
    wire n643;
    wire n647;
    wire n651;
    wire n655;
    wire n658;
    wire n662;
    wire n666;
    wire n670;
    wire n674;
    wire n678;
    wire n681;
    wire n684;
    wire n688;
    wire n692;
    wire n696;
    wire n700;
    wire n703;
    wire n707;
    wire n711;
    wire n715;
    wire n719;
    wire n723;
    wire n726;
    wire n730;
    wire n734;
    wire n738;
    wire n742;
    wire n745;
    wire n749;
    wire n753;
    wire n757;
    wire n761;
    wire n764;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n782;
    wire n786;
    wire n790;
    wire n794;
    wire n798;
    wire n801;
    wire n805;
    wire n809;
    wire n813;
    wire n816;
    wire n820;
    wire n824;
    wire n828;
    wire n832;
    wire n836;
    wire n840;
    wire n844;
    wire n848;
    wire n851;
    wire n855;
    wire n859;
    wire n863;
    wire n867;
    wire n871;
    wire n874;
    wire n877;
    wire n881;
    wire n885;
    wire n889;
    wire n893;
    wire n896;
    wire n900;
    wire n904;
    wire n908;
    wire n912;
    wire n916;
    wire n919;
    wire n923;
    wire n927;
    wire n931;
    wire n935;
    wire n938;
    wire n942;
    wire n946;
    wire n950;
    wire n954;
    wire n957;
    wire n961;
    wire n965;
    wire n969;
    wire n973;
    wire n976;
    wire n979;
    wire n983;
    wire n987;
    wire n991;
    wire n994;
    wire n998;
    wire n1002;
    wire n1006;
    wire n1010;
    wire n1013;
    wire n1017;
    wire n1021;
    wire n1025;
    wire n1028;
    wire n1032;
    wire n1036;
    wire n1040;
    wire n1044;
    wire n1048;
    wire n1052;
    wire n1056;
    wire n1060;
    wire n1064;
    wire n1068;
    wire n1071;
    wire n1075;
    wire n1079;
    wire n1083;
    wire n1087;
    wire n1091;
    wire n1094;
    wire n1097;
    wire n1101;
    wire n1105;
    wire n1109;
    wire n1113;
    wire n1116;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1139;
    wire n1143;
    wire n1147;
    wire n1151;
    wire n1155;
    wire n1158;
    wire n1162;
    wire n1166;
    wire n1170;
    wire n1174;
    wire n1177;
    wire n1181;
    wire n1185;
    wire n1189;
    wire n1193;
    wire n1196;
    wire n1200;
    wire n1204;
    wire n1208;
    wire n1212;
    wire n1215;
    wire n1218;
    wire n1222;
    wire n1226;
    wire n1230;
    wire n1234;
    wire n1238;
    wire n1242;
    wire n1246;
    wire n1249;
    wire n1253;
    wire n1257;
    wire n1260;
    wire n1264;
    wire n1268;
    wire n1272;
    wire n1276;
    wire n1280;
    wire n1284;
    wire n1288;
    wire n1292;
    wire n1296;
    wire n1300;
    wire n1304;
    wire n1308;
    wire n1312;
    wire n1315;
    wire n1319;
    wire n1323;
    wire n1327;
    wire n1331;
    wire n1335;
    wire n1338;
    wire n1341;
    wire n1345;
    wire n1349;
    wire n1353;
    wire n1357;
    wire n1360;
    wire n1364;
    wire n1368;
    wire n1372;
    wire n1376;
    wire n1380;
    wire n1383;
    wire n1387;
    wire n1391;
    wire n1395;
    wire n1399;
    wire n1402;
    wire n1406;
    wire n1410;
    wire n1414;
    wire n1418;
    wire n1421;
    wire n1425;
    wire n1429;
    wire n1433;
    wire n1437;
    wire n1440;
    wire n1444;
    wire n1448;
    wire n1452;
    wire n1456;
    wire n1459;
    wire n1463;
    wire n1467;
    wire n1471;
    wire n1475;
    wire n1478;
    wire n1481;
    wire n1484;
    wire n1488;
    wire n1492;
    wire n1496;
    wire n1500;
    wire n1504;
    wire n1508;
    wire n1512;
    wire n1515;
    wire n1519;
    wire n1523;
    wire n1526;
    wire n1530;
    wire n1534;
    wire n1538;
    wire n1542;
    wire n1546;
    wire n1550;
    wire n1554;
    wire n1558;
    wire n1562;
    wire n1566;
    wire n1570;
    wire n1574;
    wire n1578;
    wire n1582;
    wire n1586;
    wire n1589;
    wire n1593;
    wire n1597;
    wire n1601;
    wire n1605;
    wire n1609;
    wire n1612;
    wire n1615;
    wire n1619;
    wire n1623;
    wire n1627;
    wire n1631;
    wire n1634;
    wire n1638;
    wire n1642;
    wire n1646;
    wire n1650;
    wire n1654;
    wire n1657;
    wire n1661;
    wire n1665;
    wire n1669;
    wire n1673;
    wire n1676;
    wire n1680;
    wire n1684;
    wire n1688;
    wire n1692;
    wire n1695;
    wire n1699;
    wire n1703;
    wire n1707;
    wire n1711;
    wire n1714;
    wire n1718;
    wire n1722;
    wire n1726;
    wire n1730;
    wire n1733;
    wire n1737;
    wire n1741;
    wire n1745;
    wire n1749;
    wire n1752;
    wire n1756;
    wire n1760;
    wire n1764;
    wire n1768;
    wire n1771;
    wire n1774;
    wire n1777;
    wire n1781;
    wire n1785;
    wire n1789;
    wire n1793;
    wire n1797;
    wire n1801;
    wire n1805;
    wire n1808;
    wire n1812;
    wire n1816;
    wire n1819;
    wire n1823;
    wire n1827;
    wire n1831;
    wire n1835;
    wire n1839;
    wire n1843;
    wire n1847;
    wire n1851;
    wire n1855;
    wire n1859;
    wire n1863;
    wire n1867;
    wire n1871;
    wire n1875;
    wire n1879;
    wire n1883;
    wire n1887;
    wire n1890;
    wire n1894;
    wire n1898;
    wire n1902;
    wire n1906;
    wire n1910;
    wire n1913;
    wire n1916;
    wire n1920;
    wire n1924;
    wire n1928;
    wire n1932;
    wire n1935;
    wire n1939;
    wire n1943;
    wire n1947;
    wire n1951;
    wire n1955;
    wire n1958;
    wire n1962;
    wire n1966;
    wire n1970;
    wire n1974;
    wire n1977;
    wire n1981;
    wire n1985;
    wire n1989;
    wire n1993;
    wire n1996;
    wire n2000;
    wire n2004;
    wire n2008;
    wire n2012;
    wire n2015;
    wire n2019;
    wire n2023;
    wire n2027;
    wire n2031;
    wire n2034;
    wire n2038;
    wire n2042;
    wire n2046;
    wire n2050;
    wire n2053;
    wire n2057;
    wire n2061;
    wire n2065;
    wire n2069;
    wire n2072;
    wire n2076;
    wire n2080;
    wire n2084;
    wire n2088;
    wire n2091;
    wire n2094;
    wire n2097;
    wire n2101;
    wire n2105;
    wire n2109;
    wire n2113;
    wire n2117;
    wire n2121;
    wire n2125;
    wire n2128;
    wire n2132;
    wire n2136;
    wire n2139;
    wire n2143;
    wire n2147;
    wire n2151;
    wire n2155;
    wire n2159;
    wire n2163;
    wire n2167;
    wire n2171;
    wire n2175;
    wire n2179;
    wire n2183;
    wire n2187;
    wire n2191;
    wire n2195;
    wire n2199;
    wire n2203;
    wire n2207;
    wire n2211;
    wire n2215;
    wire n2218;
    wire n2222;
    wire n2226;
    wire n2230;
    wire n2234;
    wire n2238;
    wire n2241;
    wire n2244;
    wire n2248;
    wire n2252;
    wire n2256;
    wire n2260;
    wire n2263;
    wire n2267;
    wire n2271;
    wire n2275;
    wire n2279;
    wire n2283;
    wire n2286;
    wire n2290;
    wire n2294;
    wire n2298;
    wire n2302;
    wire n2305;
    wire n2309;
    wire n2313;
    wire n2317;
    wire n2321;
    wire n2324;
    wire n2328;
    wire n2332;
    wire n2336;
    wire n2340;
    wire n2343;
    wire n2347;
    wire n2351;
    wire n2355;
    wire n2359;
    wire n2362;
    wire n2366;
    wire n2370;
    wire n2374;
    wire n2378;
    wire n2381;
    wire n2385;
    wire n2389;
    wire n2393;
    wire n2397;
    wire n2400;
    wire n2404;
    wire n2408;
    wire n2412;
    wire n2416;
    wire n2419;
    wire n2423;
    wire n2427;
    wire n2431;
    wire n2435;
    wire n2438;
    wire n2441;
    wire n2444;
    wire n2448;
    wire n2452;
    wire n2456;
    wire n2460;
    wire n2464;
    wire n2468;
    wire n2472;
    wire n2475;
    wire n2479;
    wire n2483;
    wire n2486;
    wire n2490;
    wire n2494;
    wire n2498;
    wire n2502;
    wire n2506;
    wire n2510;
    wire n2514;
    wire n2518;
    wire n2522;
    wire n2526;
    wire n2530;
    wire n2534;
    wire n2538;
    wire n2542;
    wire n2546;
    wire n2550;
    wire n2554;
    wire n2558;
    wire n2562;
    wire n2566;
    wire n2570;
    wire n2573;
    wire n2577;
    wire n2581;
    wire n2585;
    wire n2589;
    wire n2593;
    wire n2596;
    wire n2599;
    wire n2603;
    wire n2607;
    wire n2611;
    wire n2615;
    wire n2618;
    wire n2622;
    wire n2626;
    wire n2630;
    wire n2634;
    wire n2638;
    wire n2641;
    wire n2645;
    wire n2649;
    wire n2653;
    wire n2657;
    wire n2660;
    wire n2664;
    wire n2668;
    wire n2672;
    wire n2676;
    wire n2679;
    wire n2683;
    wire n2687;
    wire n2691;
    wire n2695;
    wire n2698;
    wire n2702;
    wire n2706;
    wire n2710;
    wire n2714;
    wire n2717;
    wire n2721;
    wire n2725;
    wire n2729;
    wire n2733;
    wire n2736;
    wire n2740;
    wire n2744;
    wire n2748;
    wire n2752;
    wire n2755;
    wire n2759;
    wire n2763;
    wire n2767;
    wire n2771;
    wire n2774;
    wire n2778;
    wire n2782;
    wire n2786;
    wire n2790;
    wire n2793;
    wire n2797;
    wire n2801;
    wire n2805;
    wire n2809;
    wire n2812;
    wire n2815;
    wire n2818;
    wire n2822;
    wire n2826;
    wire n2830;
    wire n2834;
    wire n2838;
    wire n2842;
    wire n2846;
    wire n2849;
    wire n2853;
    wire n2857;
    wire n2860;
    wire n2864;
    wire n2868;
    wire n2872;
    wire n2876;
    wire n2880;
    wire n2884;
    wire n2888;
    wire n2892;
    wire n2896;
    wire n2900;
    wire n2904;
    wire n2908;
    wire n2912;
    wire n2916;
    wire n2920;
    wire n2924;
    wire n2928;
    wire n2932;
    wire n2936;
    wire n2940;
    wire n2944;
    wire n2948;
    wire n2952;
    wire n2955;
    wire n2959;
    wire n2963;
    wire n2967;
    wire n2971;
    wire n2975;
    wire n2978;
    wire n2981;
    wire n2985;
    wire n2989;
    wire n2993;
    wire n2997;
    wire n3001;
    wire n3005;
    wire n3009;
    wire n3013;
    wire n3017;
    wire n3020;
    wire n3024;
    wire n3028;
    wire n3032;
    wire n3036;
    wire n3039;
    wire n3043;
    wire n3047;
    wire n3051;
    wire n3055;
    wire n3058;
    wire n3062;
    wire n3066;
    wire n3070;
    wire n3074;
    wire n3077;
    wire n3081;
    wire n3085;
    wire n3089;
    wire n3093;
    wire n3096;
    wire n3100;
    wire n3104;
    wire n3108;
    wire n3112;
    wire n3115;
    wire n3119;
    wire n3123;
    wire n3127;
    wire n3131;
    wire n3134;
    wire n3138;
    wire n3142;
    wire n3146;
    wire n3150;
    wire n3153;
    wire n3157;
    wire n3161;
    wire n3165;
    wire n3169;
    wire n3172;
    wire n3176;
    wire n3180;
    wire n3184;
    wire n3188;
    wire n3191;
    wire n3195;
    wire n3199;
    wire n3203;
    wire n3207;
    wire n3210;
    wire n3213;
    wire n3216;
    wire n3220;
    wire n3224;
    wire n3228;
    wire n3231;
    wire n3235;
    wire n3239;
    wire n3242;
    wire n3246;
    wire n3250;
    wire n3254;
    wire n3257;
    wire n3261;
    wire n3265;
    wire n3269;
    wire n3273;
    wire n3277;
    wire n3281;
    wire n3285;
    wire n3289;
    wire n3293;
    wire n3297;
    wire n3301;
    wire n3305;
    wire n3309;
    wire n3313;
    wire n3317;
    wire n3321;
    wire n3325;
    wire n3329;
    wire n3333;
    wire n3337;
    wire n3341;
    wire n3345;
    wire n3349;
    wire n3353;
    wire n3357;
    wire n3361;
    wire n3365;
    wire n3369;
    wire n3373;
    wire n3376;
    wire n3380;
    wire n3384;
    wire n3388;
    wire n3392;
    wire n3395;
    wire n3399;
    wire n3403;
    wire n3407;
    wire n3411;
    wire n3415;
    wire n3418;
    wire n3421;
    wire n3425;
    wire n3429;
    wire n3433;
    wire n3437;
    wire n3440;
    wire n3444;
    wire n3448;
    wire n3452;
    wire n3456;
    wire n3459;
    wire n3463;
    wire n3467;
    wire n3471;
    wire n3475;
    wire n3478;
    wire n3482;
    wire n3486;
    wire n3490;
    wire n3494;
    wire n3497;
    wire n3501;
    wire n3505;
    wire n3509;
    wire n3513;
    wire n3516;
    wire n3520;
    wire n3524;
    wire n3528;
    wire n3532;
    wire n3535;
    wire n3539;
    wire n3543;
    wire n3547;
    wire n3551;
    wire n3554;
    wire n3558;
    wire n3562;
    wire n3566;
    wire n3570;
    wire n3573;
    wire n3577;
    wire n3581;
    wire n3585;
    wire n3589;
    wire n3592;
    wire n3596;
    wire n3600;
    wire n3604;
    wire n3608;
    wire n3611;
    wire n3615;
    wire n3619;
    wire n3623;
    wire n3627;
    wire n3630;
    wire n3633;
    wire n3636;
    wire n3640;
    wire n3644;
    wire n3648;
    wire n3652;
    wire n3655;
    wire n3659;
    wire n3663;
    wire n3667;
    wire n3671;
    wire n3675;
    wire n3679;
    wire n3683;
    wire n3687;
    wire n3691;
    wire n3695;
    wire n3699;
    wire n3703;
    wire n3707;
    wire n3711;
    wire n3715;
    wire n3719;
    wire n3723;
    wire n3727;
    wire n3731;
    wire n3735;
    wire n3739;
    wire n3743;
    wire n3747;
    wire n3751;
    wire n3755;
    wire n3759;
    wire n3762;
    wire n3766;
    wire n3770;
    wire n3774;
    wire n3778;
    wire n3782;
    wire n3786;
    wire n3790;
    wire n3794;
    wire n3798;
    wire n3801;
    wire n3805;
    wire n3809;
    wire n3813;
    wire n3817;
    wire n3821;
    wire n3825;
    wire n3829;
    wire n3833;
    wire n3836;
    wire n3840;
    wire n3844;
    wire n3848;
    wire n3852;
    wire n3855;
    wire n3859;
    wire n3863;
    wire n3867;
    wire n3871;
    wire n3874;
    wire n3878;
    wire n3882;
    wire n3886;
    wire n3890;
    wire n3893;
    wire n3897;
    wire n3901;
    wire n3905;
    wire n3909;
    wire n3912;
    wire n3916;
    wire n3920;
    wire n3924;
    wire n3928;
    wire n3931;
    wire n3935;
    wire n3939;
    wire n3943;
    wire n3947;
    wire n3950;
    wire n3954;
    wire n3958;
    wire n3962;
    wire n3966;
    wire n3969;
    wire n3973;
    wire n3977;
    wire n3981;
    wire n3985;
    wire n3988;
    wire n3992;
    wire n3996;
    wire n4000;
    wire n4004;
    wire n4007;
    wire n4011;
    wire n4015;
    wire n4019;
    wire n4023;
    wire n4027;
    wire n4030;
    wire n4033;
    wire n4037;
    wire n4041;
    wire n4044;
    wire n4048;
    wire n4052;
    wire n4055;
    wire n4059;
    wire n4062;
    wire n4066;
    wire n4070;
    wire n4074;
    wire n4078;
    wire n4082;
    wire n4086;
    wire n4090;
    wire n4094;
    wire n4098;
    wire n4102;
    wire n4106;
    wire n4110;
    wire n4114;
    wire n4118;
    wire n4122;
    wire n4126;
    wire n4130;
    wire n4134;
    wire n4138;
    wire n4142;
    wire n4146;
    wire n4150;
    wire n4153;
    wire n4157;
    wire n4161;
    wire n4165;
    wire n4169;
    wire n4172;
    wire n4176;
    wire n4179;
    wire n4183;
    wire n4187;
    wire n4191;
    wire n4194;
    wire n4198;
    wire n4202;
    wire n4206;
    wire n4210;
    wire n4214;
    wire n4217;
    wire n4221;
    wire n4225;
    wire n4229;
    wire n4232;
    wire n4236;
    wire n4240;
    wire n4244;
    wire n4248;
    wire n4251;
    wire n4255;
    wire n4259;
    wire n4263;
    wire n4267;
    wire n4270;
    wire n4274;
    wire n4278;
    wire n4282;
    wire n4286;
    wire n4289;
    wire n4293;
    wire n4297;
    wire n4301;
    wire n4305;
    wire n4308;
    wire n4312;
    wire n4316;
    wire n4320;
    wire n4324;
    wire n4327;
    wire n4331;
    wire n4335;
    wire n4339;
    wire n4343;
    wire n4346;
    wire n4350;
    wire n4354;
    wire n4358;
    wire n4362;
    wire n4365;
    wire n4369;
    wire n4373;
    wire n4377;
    wire n4381;
    wire n4384;
    wire n4388;
    wire n4392;
    wire n4396;
    wire n4400;
    wire n4403;
    wire n4407;
    wire n4411;
    wire n4415;
    wire n4419;
    wire n4423;
    wire n4427;
    wire n4431;
    wire n4435;
    wire n4438;
    wire n4442;
    wire n4446;
    wire n4450;
    wire n4454;
    wire n4458;
    wire n4462;
    wire n4466;
    wire n4470;
    wire n4474;
    wire n4478;
    wire n4482;
    wire n4486;
    wire n4490;
    wire n4494;
    wire n4498;
    wire n4502;
    wire n4506;
    wire n4510;
    wire n4514;
    wire n4518;
    wire n4522;
    wire n4525;
    wire n4529;
    wire n4532;
    wire n4536;
    wire n4540;
    wire n4543;
    wire n4547;
    wire n4550;
    wire n4554;
    wire n4558;
    wire n4562;
    wire n4566;
    wire n4570;
    wire n4574;
    wire n4578;
    wire n4582;
    wire n4586;
    wire n4590;
    wire n4594;
    wire n4597;
    wire n4601;
    wire n4605;
    wire n4609;
    wire n4613;
    wire n4616;
    wire n4620;
    wire n4624;
    wire n4628;
    wire n4632;
    wire n4635;
    wire n4639;
    wire n4643;
    wire n4647;
    wire n4651;
    wire n4654;
    wire n4658;
    wire n4662;
    wire n4666;
    wire n4670;
    wire n4673;
    wire n4677;
    wire n4681;
    wire n4685;
    wire n4689;
    wire n4692;
    wire n4696;
    wire n4700;
    wire n4704;
    wire n4708;
    wire n4711;
    wire n4715;
    wire n4719;
    wire n4723;
    wire n4727;
    wire n4730;
    wire n4734;
    wire n4738;
    wire n4742;
    wire n4746;
    wire n4749;
    wire n4753;
    wire n4757;
    wire n4761;
    wire n4765;
    wire n4769;
    wire n4773;
    wire n4777;
    wire n4781;
    wire n4785;
    wire n4788;
    wire n4792;
    wire n4796;
    wire n4800;
    wire n4804;
    wire n4808;
    wire n4812;
    wire n4816;
    wire n4820;
    wire n4824;
    wire n4828;
    wire n4832;
    wire n4836;
    wire n4840;
    wire n4844;
    wire n4848;
    wire n4852;
    wire n4856;
    wire n4860;
    wire n4864;
    wire n4868;
    wire n4871;
    wire n4875;
    wire n4879;
    wire n4882;
    wire n4886;
    wire n4889;
    wire n4893;
    wire n4897;
    wire n4901;
    wire n4904;
    wire n4907;
    wire n4911;
    wire n4915;
    wire n4919;
    wire n4923;
    wire n4927;
    wire n4931;
    wire n4935;
    wire n4939;
    wire n4942;
    wire n4946;
    wire n4950;
    wire n4954;
    wire n4958;
    wire n4961;
    wire n4965;
    wire n4969;
    wire n4973;
    wire n4977;
    wire n4980;
    wire n4984;
    wire n4988;
    wire n4992;
    wire n4996;
    wire n4999;
    wire n5003;
    wire n5007;
    wire n5011;
    wire n5015;
    wire n5018;
    wire n5022;
    wire n5026;
    wire n5030;
    wire n5034;
    wire n5037;
    wire n5041;
    wire n5045;
    wire n5049;
    wire n5053;
    wire n5056;
    wire n5060;
    wire n5064;
    wire n5068;
    wire n5072;
    wire n5075;
    wire n5079;
    wire n5083;
    wire n5087;
    wire n5091;
    wire n5095;
    wire n5099;
    wire n5103;
    wire n5107;
    wire n5111;
    wire n5114;
    wire n5118;
    wire n5122;
    wire n5126;
    wire n5130;
    wire n5134;
    wire n5138;
    wire n5142;
    wire n5146;
    wire n5150;
    wire n5154;
    wire n5158;
    wire n5162;
    wire n5166;
    wire n5170;
    wire n5174;
    wire n5178;
    wire n5182;
    wire n5186;
    wire n5189;
    wire n5193;
    wire n5196;
    wire n5200;
    wire n5204;
    wire n5208;
    wire n5211;
    wire n5215;
    wire n5219;
    wire n5222;
    wire n5225;
    wire n5229;
    wire n5233;
    wire n5237;
    wire n5241;
    wire n5245;
    wire n5249;
    wire n5253;
    wire n5257;
    wire n5260;
    wire n5264;
    wire n5268;
    wire n5272;
    wire n5276;
    wire n5279;
    wire n5283;
    wire n5287;
    wire n5291;
    wire n5295;
    wire n5298;
    wire n5302;
    wire n5306;
    wire n5310;
    wire n5314;
    wire n5317;
    wire n5321;
    wire n5325;
    wire n5329;
    wire n5333;
    wire n5336;
    wire n5340;
    wire n5344;
    wire n5348;
    wire n5352;
    wire n5355;
    wire n5359;
    wire n5363;
    wire n5367;
    wire n5371;
    wire n5374;
    wire n5378;
    wire n5382;
    wire n5386;
    wire n5390;
    wire n5394;
    wire n5398;
    wire n5402;
    wire n5406;
    wire n5410;
    wire n5413;
    wire n5417;
    wire n5421;
    wire n5425;
    wire n5429;
    wire n5433;
    wire n5437;
    wire n5441;
    wire n5445;
    wire n5449;
    wire n5453;
    wire n5457;
    wire n5461;
    wire n5465;
    wire n5469;
    wire n5473;
    wire n5477;
    wire n5480;
    wire n5484;
    wire n5487;
    wire n5491;
    wire n5495;
    wire n5499;
    wire n5502;
    wire n5506;
    wire n5510;
    wire n5513;
    wire n5516;
    wire n5520;
    wire n5524;
    wire n5528;
    wire n5532;
    wire n5536;
    wire n5540;
    wire n5544;
    wire n5548;
    wire n5551;
    wire n5555;
    wire n5559;
    wire n5563;
    wire n5567;
    wire n5570;
    wire n5574;
    wire n5578;
    wire n5582;
    wire n5586;
    wire n5589;
    wire n5593;
    wire n5597;
    wire n5601;
    wire n5605;
    wire n5608;
    wire n5612;
    wire n5616;
    wire n5620;
    wire n5624;
    wire n5627;
    wire n5631;
    wire n5635;
    wire n5639;
    wire n5643;
    wire n5646;
    wire n5650;
    wire n5654;
    wire n5658;
    wire n5662;
    wire n5666;
    wire n5670;
    wire n5674;
    wire n5678;
    wire n5682;
    wire n5685;
    wire n5689;
    wire n5693;
    wire n5697;
    wire n5701;
    wire n5705;
    wire n5709;
    wire n5713;
    wire n5717;
    wire n5721;
    wire n5725;
    wire n5729;
    wire n5733;
    wire n5737;
    wire n5741;
    wire n5744;
    wire n5748;
    wire n5751;
    wire n5755;
    wire n5759;
    wire n5763;
    wire n5766;
    wire n5770;
    wire n5774;
    wire n5777;
    wire n5780;
    wire n5784;
    wire n5788;
    wire n5792;
    wire n5796;
    wire n5800;
    wire n5804;
    wire n5808;
    wire n5812;
    wire n5815;
    wire n5819;
    wire n5823;
    wire n5827;
    wire n5831;
    wire n5834;
    wire n5838;
    wire n5842;
    wire n5846;
    wire n5850;
    wire n5853;
    wire n5857;
    wire n5861;
    wire n5865;
    wire n5869;
    wire n5872;
    wire n5876;
    wire n5880;
    wire n5884;
    wire n5888;
    wire n5891;
    wire n5895;
    wire n5899;
    wire n5903;
    wire n5907;
    wire n5911;
    wire n5915;
    wire n5919;
    wire n5923;
    wire n5927;
    wire n5930;
    wire n5934;
    wire n5938;
    wire n5942;
    wire n5946;
    wire n5950;
    wire n5954;
    wire n5958;
    wire n5962;
    wire n5966;
    wire n5970;
    wire n5974;
    wire n5978;
    wire n5981;
    wire n5985;
    wire n5988;
    wire n5992;
    wire n5996;
    wire n6000;
    wire n6003;
    wire n6007;
    wire n6011;
    wire n6014;
    wire n6017;
    wire n6021;
    wire n6025;
    wire n6029;
    wire n6033;
    wire n6037;
    wire n6041;
    wire n6045;
    wire n6049;
    wire n6052;
    wire n6056;
    wire n6060;
    wire n6064;
    wire n6068;
    wire n6071;
    wire n6075;
    wire n6079;
    wire n6083;
    wire n6087;
    wire n6090;
    wire n6094;
    wire n6098;
    wire n6102;
    wire n6106;
    wire n6109;
    wire n6113;
    wire n6117;
    wire n6121;
    wire n6125;
    wire n6129;
    wire n6133;
    wire n6137;
    wire n6141;
    wire n6145;
    wire n6148;
    wire n6152;
    wire n6156;
    wire n6160;
    wire n6164;
    wire n6168;
    wire n6172;
    wire n6176;
    wire n6180;
    wire n6184;
    wire n6188;
    wire n6191;
    wire n6195;
    wire n6198;
    wire n6202;
    wire n6206;
    wire n6210;
    wire n6213;
    wire n6217;
    wire n6221;
    wire n6224;
    wire n6227;
    wire n6231;
    wire n6235;
    wire n6239;
    wire n6243;
    wire n6246;
    wire n6250;
    wire n6254;
    wire n6258;
    wire n6262;
    wire n6265;
    wire n6269;
    wire n6273;
    wire n6277;
    wire n6281;
    wire n6284;
    wire n6288;
    wire n6292;
    wire n6296;
    wire n6300;
    wire n6303;
    wire n6307;
    wire n6311;
    wire n6315;
    wire n6319;
    wire n6323;
    wire n6327;
    wire n6331;
    wire n6335;
    wire n6339;
    wire n6342;
    wire n6346;
    wire n6350;
    wire n6354;
    wire n6358;
    wire n6362;
    wire n6366;
    wire n6370;
    wire n6374;
    wire n6378;
    wire n6381;
    wire n6385;
    wire n6389;
    wire n6393;
    wire n6396;
    wire n6400;
    wire n6404;
    wire n6408;
    wire n6412;
    wire n6416;
    wire n6420;
    wire n6423;
    wire n6427;
    wire n6431;
    wire n6435;
    wire n6439;
    wire n6442;
    wire n6446;
    wire n6450;
    wire n6454;
    wire n6458;
    wire n6461;
    wire n6465;
    wire n6469;
    wire n6473;
    wire n6477;
    wire n6481;
    wire n6485;
    wire n6489;
    wire n6493;
    wire n6497;
    wire n6500;
    wire n6504;
    wire n6508;
    wire n6512;
    wire n6516;
    wire n6520;
    wire n6524;
    wire n6528;
    wire n6532;
    wire n6536;
    wire n6539;
    wire n6542;
    wire n6546;
    wire n6549;
    wire n6553;
    wire n6557;
    wire n6561;
    wire n6565;
    wire n6569;
    wire n6573;
    wire n6576;
    wire n6580;
    wire n6584;
    wire n6588;
    wire n6592;
    wire n6595;
    wire n6599;
    wire n6603;
    wire n6607;
    wire n6611;
    wire n6615;
    wire n6619;
    wire n6623;
    wire n6627;
    wire n6631;
    wire n6634;
    wire n6638;
    wire n6642;
    wire n6646;
    wire n6650;
    wire n6654;
    wire n6658;
    wire n6662;
    wire n6665;
    wire n6668;
    wire n6672;
    wire n6675;
    wire n6679;
    wire n6683;
    wire n6687;
    wire n6691;
    wire n6695;
    wire n6699;
    wire n6702;
    wire n6706;
    wire n6710;
    wire n6714;
    wire n6718;
    wire n6722;
    wire n6726;
    wire n6730;
    wire n6734;
    wire n6738;
    wire n6741;
    wire n6745;
    wire n6749;
    wire n6753;
    wire n6757;
    wire n6761;
    wire n6764;
    wire n6767;
    wire n6771;
    wire n6774;
    wire n6778;
    wire n6782;
    wire n6786;
    wire n6790;
    wire n6794;
    wire n6798;
    wire n6802;
    wire n6806;
    wire n6810;
    wire n6814;
    wire n6818;
    wire n6821;
    wire n6825;
    wire n6829;
    wire n6833;
    wire n6837;
    wire n6841;
    wire n6845;
    wire n6849;
    wire n6853;
    wire n6856;
    wire n6859;
    wire n6863;
    wire n6866;
    wire n6870;
    wire n6874;
    wire n6878;
    wire n6881;
    wire n6885;
    wire n6893;
    wire n10756;
    wire n10759;
    wire n10762;
    wire n10765;
    wire n10768;
    wire n10771;
    wire n10774;
    wire n10777;
    wire n10780;
    wire n10783;
    wire n10786;
    wire n10789;
    wire n10792;
    wire n10795;
    wire n10798;
    wire n10801;
    wire n10804;
    wire n10807;
    wire n10810;
    wire n10813;
    wire n10816;
    wire n10819;
    wire n10822;
    wire n10825;
    wire n10828;
    wire n10831;
    wire n10834;
    wire n10837;
    wire n10840;
    wire n10843;
    wire n10846;
    wire n10849;
    wire n10852;
    wire n10855;
    wire n10858;
    wire n10861;
    wire n10864;
    wire n10867;
    wire n10870;
    wire n10873;
    wire n10876;
    wire n10879;
    wire n10882;
    wire n10885;
    wire n10888;
    wire n10891;
    wire n10894;
    wire n10897;
    wire n10900;
    wire n10903;
    wire n10906;
    wire n10909;
    wire n10912;
    wire n10915;
    wire n10918;
    wire n10921;
    wire n10924;
    wire n10927;
    wire n10930;
    wire n10933;
    wire n10936;
    wire n10939;
    wire n10942;
    wire n10945;
    wire n10948;
    wire n10951;
    wire n10954;
    wire n10957;
    wire n10960;
    wire n10963;
    wire n10966;
    wire n10969;
    wire n10972;
    wire n10975;
    wire n10978;
    wire n10981;
    wire n10984;
    wire n10987;
    wire n10990;
    wire n10993;
    wire n10996;
    wire n10999;
    wire n11002;
    wire n11005;
    wire n11008;
    wire n11011;
    wire n11014;
    wire n11017;
    wire n11020;
    wire n11023;
    wire n11026;
    wire n11029;
    wire n11032;
    wire n11035;
    wire n11038;
    wire n11041;
    wire n11044;
    wire n11047;
    wire n11050;
    wire n11053;
    wire n11056;
    wire n11059;
    wire n11062;
    wire n11065;
    wire n11068;
    wire n11071;
    wire n11074;
    wire n11077;
    wire n11080;
    wire n11083;
    wire n11086;
    wire n11089;
    wire n11092;
    wire n11095;
    wire n11098;
    wire n11101;
    wire n11104;
    wire n11107;
    wire n11110;
    wire n11113;
    wire n11116;
    wire n11119;
    wire n11122;
    wire n11125;
    wire n11128;
    wire n11131;
    wire n11134;
    wire n11137;
    wire n11140;
    wire n11143;
    wire n11146;
    wire n11149;
    wire n11152;
    wire n11155;
    wire n11158;
    wire n11161;
    wire n11164;
    wire n11167;
    wire n11170;
    wire n11173;
    wire n11176;
    wire n11179;
    wire n11182;
    wire n11185;
    wire n11188;
    wire n11191;
    wire n11194;
    wire n11197;
    wire n11200;
    wire n11203;
    wire n11206;
    wire n11209;
    wire n11212;
    wire n11215;
    wire n11218;
    wire n11221;
    wire n11224;
    wire n11227;
    wire n11230;
    wire n11233;
    wire n11236;
    wire n11239;
    wire n11242;
    wire n11245;
    wire n11248;
    wire n11251;
    wire n11254;
    wire n11257;
    wire n11260;
    wire n11263;
    wire n11266;
    wire n11269;
    wire n11272;
    wire n11275;
    wire n11278;
    wire n11281;
    wire n11284;
    wire n11287;
    wire n11290;
    wire n11293;
    wire n11296;
    wire n11299;
    wire n11302;
    wire n11305;
    wire n11308;
    wire n11311;
    wire n11314;
    wire n11317;
    wire n11320;
    wire n11323;
    wire n11326;
    wire n11329;
    wire n11332;
    wire n11335;
    wire n11338;
    wire n11341;
    wire n11344;
    wire n11347;
    wire n11350;
    wire n11353;
    wire n11356;
    wire n11359;
    wire n11362;
    wire n11365;
    wire n11368;
    wire n11371;
    wire n11374;
    wire n11377;
    wire n11380;
    wire n11383;
    wire n11386;
    wire n11389;
    wire n11392;
    wire n11395;
    wire n11398;
    wire n11401;
    wire n11404;
    wire n11407;
    wire n11410;
    wire n11413;
    wire n11416;
    wire n11419;
    wire n11422;
    wire n11425;
    wire n11428;
    wire n11431;
    wire n11434;
    wire n11437;
    wire n11440;
    wire n11443;
    wire n11446;
    wire n11449;
    wire n11452;
    wire n11455;
    wire n11458;
    wire n11461;
    wire n11464;
    wire n11467;
    wire n11470;
    wire n11473;
    wire n11476;
    wire n11479;
    wire n11482;
    wire n11485;
    wire n11488;
    wire n11491;
    wire n11494;
    wire n11497;
    wire n11500;
    wire n11503;
    wire n11506;
    wire n11509;
    wire n11512;
    wire n11515;
    wire n11518;
    wire n11521;
    wire n11524;
    wire n11527;
    wire n11530;
    wire n11533;
    wire n11536;
    wire n11539;
    wire n11542;
    wire n11545;
    wire n11548;
    wire n11551;
    wire n11554;
    wire n11557;
    wire n11560;
    wire n11563;
    wire n11566;
    wire n11569;
    wire n11572;
    wire n11575;
    wire n11578;
    wire n11581;
    wire n11584;
    wire n11587;
    wire n11590;
    wire n11593;
    wire n11596;
    wire n11599;
    wire n11602;
    wire n11605;
    wire n11608;
    wire n11611;
    wire n11614;
    wire n11617;
    wire n11620;
    wire n11623;
    wire n11626;
    wire n11629;
    wire n11632;
    wire n11635;
    wire n11638;
    wire n11641;
    wire n11644;
    wire n11647;
    wire n11650;
    wire n11653;
    wire n11656;
    wire n11659;
    wire n11662;
    wire n11665;
    wire n11668;
    wire n11671;
    wire n11674;
    wire n11677;
    wire n11680;
    wire n11683;
    wire n11686;
    wire n11689;
    wire n11692;
    wire n11695;
    wire n11698;
    wire n11701;
    wire n11704;
    wire n11707;
    wire n11710;
    wire n11713;
    wire n11716;
    wire n11719;
    wire n11722;
    wire n11725;
    wire n11728;
    wire n11731;
    wire n11734;
    wire n11737;
    wire n11740;
    wire n11743;
    wire n11746;
    wire n11749;
    wire n11752;
    wire n11755;
    wire n11758;
    wire n11761;
    wire n11764;
    wire n11767;
    wire n11770;
    wire n11773;
    wire n11776;
    wire n11779;
    wire n11782;
    wire n11785;
    wire n11788;
    wire n11791;
    wire n11794;
    wire n11797;
    wire n11800;
    wire n11803;
    wire n11806;
    wire n11809;
    wire n11812;
    wire n11815;
    wire n11818;
    wire n11820;
    wire n11823;
    wire n11826;
    wire n11829;
    wire n11832;
    wire n11835;
    wire n11838;
    wire n11841;
    wire n11844;
    wire n11847;
    wire n11850;
    wire n11853;
    wire n11857;
    wire n11860;
    wire n11863;
    wire n11866;
    wire n11869;
    wire n11872;
    wire n11875;
    wire n11878;
    wire n11881;
    wire n11884;
    wire n11887;
    wire n11890;
    wire n11893;
    wire n11896;
    wire n11899;
    wire n11902;
    wire n11905;
    wire n11908;
    wire n11911;
    wire n11914;
    wire n11917;
    wire n11920;
    wire n11923;
    wire n11926;
    wire n11929;
    wire n11932;
    wire n11935;
    wire n11938;
    wire n11941;
    wire n11944;
    wire n11947;
    wire n11950;
    wire n11953;
    wire n11956;
    wire n11959;
    wire n11962;
    wire n11965;
    wire n11968;
    wire n11971;
    wire n11974;
    wire n11977;
    wire n11980;
    wire n11983;
    wire n11986;
    wire n11989;
    wire n11992;
    wire n11995;
    wire n11998;
    wire n12001;
    wire n12004;
    wire n12007;
    wire n12010;
    wire n12013;
    wire n12016;
    wire n12019;
    wire n12022;
    wire n12025;
    wire n12028;
    wire n12031;
    wire n12034;
    wire n12037;
    wire n12040;
    wire n12043;
    wire n12046;
    wire n12049;
    wire n12052;
    wire n12055;
    wire n12058;
    wire n12061;
    wire n12064;
    wire n12067;
    wire n12070;
    wire n12073;
    wire n12076;
    wire n12079;
    wire n12082;
    wire n12085;
    wire n12088;
    wire n12091;
    wire n12094;
    wire n12097;
    wire n12100;
    wire n12103;
    wire n12105;
    wire n12108;
    wire n12111;
    wire n12114;
    wire n12117;
    wire n12120;
    wire n12123;
    wire n12126;
    wire n12129;
    wire n12132;
    wire n12135;
    wire n12139;
    wire n12142;
    wire n12145;
    wire n12148;
    wire n12151;
    wire n12154;
    wire n12157;
    wire n12160;
    wire n12163;
    wire n12166;
    wire n12169;
    wire n12172;
    wire n12175;
    wire n12178;
    wire n12181;
    wire n12184;
    wire n12187;
    wire n12190;
    wire n12193;
    wire n12196;
    wire n12199;
    wire n12201;
    wire n12204;
    wire n12207;
    wire n12210;
    wire n12213;
    wire n12216;
    wire n12219;
    wire n12222;
    wire n12225;
    wire n12228;
    wire n12231;
    wire n12235;
    wire n12238;
    wire n12241;
    wire n12244;
    wire n12247;
    wire n12250;
    wire n12253;
    wire n12256;
    wire n12259;
    wire n12262;
    wire n12265;
    wire n12268;
    wire n12271;
    wire n12274;
    wire n12277;
    wire n12280;
    wire n12283;
    wire n12286;
    wire n12289;
    wire n12292;
    wire n12295;
    wire n12297;
    wire n12300;
    wire n12303;
    wire n12306;
    wire n12309;
    wire n12312;
    wire n12315;
    wire n12318;
    wire n12321;
    wire n12324;
    wire n12327;
    wire n12331;
    wire n12334;
    wire n12337;
    wire n12340;
    wire n12343;
    wire n12346;
    wire n12349;
    wire n12352;
    wire n12355;
    wire n12358;
    wire n12361;
    wire n12364;
    wire n12367;
    wire n12370;
    wire n12373;
    wire n12376;
    wire n12379;
    wire n12382;
    wire n12385;
    wire n12388;
    wire n12391;
    wire n12393;
    wire n12396;
    wire n12399;
    wire n12402;
    wire n12405;
    wire n12408;
    wire n12411;
    wire n12414;
    wire n12417;
    wire n12420;
    wire n12423;
    wire n12427;
    wire n12430;
    wire n12433;
    wire n12436;
    wire n12439;
    wire n12442;
    wire n12445;
    wire n12448;
    wire n12451;
    wire n12454;
    wire n12457;
    wire n12460;
    wire n12463;
    wire n12466;
    wire n12469;
    wire n12472;
    wire n12475;
    wire n12478;
    wire n12481;
    wire n12484;
    wire n12486;
    wire n12489;
    wire n12492;
    wire n12495;
    wire n12498;
    wire n12501;
    wire n12504;
    wire n12507;
    wire n12510;
    wire n12513;
    wire n12517;
    wire n12520;
    wire n12523;
    wire n12526;
    wire n12529;
    wire n12532;
    wire n12535;
    wire n12538;
    wire n12541;
    wire n12544;
    wire n12547;
    wire n12550;
    wire n12553;
    wire n12556;
    wire n12559;
    wire n12562;
    wire n12565;
    wire n12568;
    wire n12570;
    wire n12573;
    wire n12576;
    wire n12579;
    wire n12582;
    wire n12585;
    wire n12588;
    wire n12591;
    wire n12594;
    wire n12598;
    wire n12601;
    wire n12604;
    wire n12607;
    wire n12610;
    wire n12613;
    wire n12616;
    wire n12619;
    wire n12622;
    wire n12625;
    wire n12628;
    wire n12631;
    wire n12634;
    wire n12637;
    wire n12640;
    wire n12643;
    wire n12646;
    wire n12649;
    wire n12651;
    wire n12654;
    wire n12657;
    wire n12660;
    wire n12663;
    wire n12666;
    wire n12669;
    wire n12672;
    wire n12675;
    wire n12679;
    wire n12682;
    wire n12685;
    wire n12688;
    wire n12691;
    wire n12694;
    wire n12697;
    wire n12700;
    wire n12703;
    wire n12706;
    wire n12709;
    wire n12712;
    wire n12715;
    wire n12718;
    wire n12720;
    wire n12723;
    wire n12726;
    wire n12729;
    wire n12732;
    wire n12735;
    wire n12738;
    wire n12742;
    wire n12745;
    wire n12748;
    wire n12751;
    wire n12754;
    wire n12757;
    wire n12760;
    wire n12763;
    wire n12766;
    wire n12769;
    wire n12772;
    wire n12775;
    wire n12777;
    wire n12780;
    wire n12783;
    wire n12786;
    wire n12789;
    wire n12792;
    wire n12796;
    wire n12799;
    wire n12802;
    wire n12805;
    wire n12808;
    wire n12811;
    wire n12814;
    wire n12817;
    wire n12820;
    wire n12823;
    wire n12825;
    wire n12828;
    wire n12831;
    wire n12834;
    wire n12837;
    wire n12841;
    wire n12844;
    wire n12847;
    wire n12849;
    wire n12852;
    wire n12856;
    wire n12858;
    wire n12862;
    wire n12864;
    wire n12868;
    wire n12871;
    wire n12873;
    wire n12876;
    wire n12879;
    wire n12882;
    wire n12885;
    wire n12888;
    wire n12891;
    wire n12894;
    wire n12897;
    wire n12900;
    wire n12903;
    wire n12906;
    wire n12909;
    wire n12912;
    wire n12915;
    wire n12918;
    wire n12921;
    wire n12924;
    wire n12927;
    wire n12930;
    wire n12933;
    wire n12936;
    wire n12939;
    wire n12942;
    wire n12945;
    wire n12948;
    wire n12951;
    wire n12954;
    wire n12957;
    wire n12960;
    wire n12963;
    wire n12966;
    wire n12969;
    wire n12972;
    wire n12975;
    wire n12978;
    wire n12981;
    wire n12984;
    wire n12987;
    wire n12990;
    wire n12993;
    wire n12996;
    wire n12999;
    wire n13002;
    wire n13005;
    wire n13009;
    wire n13011;
    wire n13014;
    wire n13017;
    wire n13020;
    wire n13023;
    wire n13026;
    wire n13029;
    wire n13032;
    wire n13035;
    wire n13038;
    wire n13041;
    wire n13044;
    wire n13047;
    wire n13050;
    wire n13053;
    wire n13056;
    wire n13059;
    wire n13062;
    wire n13065;
    wire n13068;
    wire n13071;
    wire n13074;
    wire n13077;
    wire n13080;
    wire n13083;
    wire n13086;
    wire n13089;
    wire n13092;
    wire n13095;
    wire n13098;
    wire n13101;
    wire n13104;
    wire n13107;
    wire n13110;
    wire n13113;
    wire n13116;
    wire n13119;
    wire n13122;
    wire n13125;
    wire n13128;
    wire n13131;
    wire n13134;
    wire n13138;
    wire n13141;
    wire n13144;
    wire n13147;
    wire n13150;
    wire n13153;
    wire n13156;
    wire n13159;
    wire n13162;
    wire n13165;
    wire n13168;
    wire n13171;
    wire n13174;
    wire n13177;
    wire n13180;
    wire n13183;
    wire n13186;
    wire n13189;
    wire n13192;
    wire n13195;
    wire n13198;
    wire n13201;
    wire n13204;
    wire n13207;
    wire n13210;
    wire n13213;
    wire n13216;
    wire n13219;
    wire n13222;
    wire n13225;
    wire n13228;
    wire n13231;
    wire n13234;
    wire n13237;
    wire n13240;
    wire n13243;
    wire n13246;
    wire n13249;
    wire n13251;
    wire n13254;
    wire n13257;
    wire n13260;
    wire n13263;
    wire n13266;
    wire n13269;
    wire n13272;
    wire n13275;
    wire n13278;
    wire n13281;
    wire n13284;
    wire n13287;
    wire n13290;
    wire n13293;
    wire n13296;
    wire n13299;
    wire n13302;
    wire n13305;
    wire n13308;
    wire n13311;
    wire n13314;
    wire n13317;
    wire n13320;
    wire n13323;
    wire n13326;
    wire n13329;
    wire n13332;
    wire n13335;
    wire n13338;
    wire n13341;
    wire n13344;
    wire n13347;
    wire n13350;
    wire n13353;
    wire n13356;
    wire n13359;
    wire n13362;
    wire n13365;
    wire n13369;
    wire n13372;
    wire n13375;
    wire n13378;
    wire n13381;
    wire n13384;
    wire n13387;
    wire n13390;
    wire n13393;
    wire n13396;
    wire n13399;
    wire n13402;
    wire n13405;
    wire n13408;
    wire n13411;
    wire n13414;
    wire n13417;
    wire n13420;
    wire n13423;
    wire n13426;
    wire n13429;
    wire n13432;
    wire n13435;
    wire n13438;
    wire n13441;
    wire n13444;
    wire n13447;
    wire n13450;
    wire n13453;
    wire n13456;
    wire n13459;
    wire n13462;
    wire n13465;
    wire n13468;
    wire n13471;
    wire n13473;
    wire n13476;
    wire n13479;
    wire n13482;
    wire n13485;
    wire n13488;
    wire n13491;
    wire n13494;
    wire n13497;
    wire n13500;
    wire n13503;
    wire n13506;
    wire n13509;
    wire n13512;
    wire n13515;
    wire n13518;
    wire n13521;
    wire n13524;
    wire n13527;
    wire n13530;
    wire n13533;
    wire n13536;
    wire n13539;
    wire n13542;
    wire n13545;
    wire n13548;
    wire n13551;
    wire n13554;
    wire n13557;
    wire n13560;
    wire n13563;
    wire n13566;
    wire n13569;
    wire n13572;
    wire n13575;
    wire n13578;
    wire n13582;
    wire n13585;
    wire n13588;
    wire n13591;
    wire n13594;
    wire n13597;
    wire n13600;
    wire n13603;
    wire n13606;
    wire n13609;
    wire n13612;
    wire n13615;
    wire n13618;
    wire n13621;
    wire n13624;
    wire n13627;
    wire n13630;
    wire n13633;
    wire n13636;
    wire n13639;
    wire n13642;
    wire n13645;
    wire n13648;
    wire n13651;
    wire n13654;
    wire n13657;
    wire n13660;
    wire n13663;
    wire n13666;
    wire n13669;
    wire n13672;
    wire n13675;
    wire n13677;
    wire n13680;
    wire n13683;
    wire n13686;
    wire n13689;
    wire n13692;
    wire n13695;
    wire n13698;
    wire n13701;
    wire n13704;
    wire n13707;
    wire n13710;
    wire n13713;
    wire n13716;
    wire n13719;
    wire n13722;
    wire n13725;
    wire n13728;
    wire n13731;
    wire n13734;
    wire n13737;
    wire n13740;
    wire n13743;
    wire n13746;
    wire n13749;
    wire n13752;
    wire n13755;
    wire n13758;
    wire n13761;
    wire n13764;
    wire n13767;
    wire n13770;
    wire n13773;
    wire n13777;
    wire n13780;
    wire n13783;
    wire n13786;
    wire n13789;
    wire n13792;
    wire n13795;
    wire n13798;
    wire n13801;
    wire n13804;
    wire n13807;
    wire n13810;
    wire n13813;
    wire n13816;
    wire n13819;
    wire n13822;
    wire n13825;
    wire n13828;
    wire n13831;
    wire n13834;
    wire n13837;
    wire n13840;
    wire n13843;
    wire n13846;
    wire n13849;
    wire n13852;
    wire n13855;
    wire n13858;
    wire n13861;
    wire n13863;
    wire n13866;
    wire n13869;
    wire n13872;
    wire n13875;
    wire n13878;
    wire n13881;
    wire n13884;
    wire n13887;
    wire n13890;
    wire n13893;
    wire n13896;
    wire n13899;
    wire n13902;
    wire n13905;
    wire n13908;
    wire n13911;
    wire n13914;
    wire n13917;
    wire n13920;
    wire n13923;
    wire n13926;
    wire n13929;
    wire n13932;
    wire n13935;
    wire n13938;
    wire n13941;
    wire n13944;
    wire n13947;
    wire n13950;
    wire n13954;
    wire n13957;
    wire n13960;
    wire n13963;
    wire n13966;
    wire n13969;
    wire n13972;
    wire n13975;
    wire n13978;
    wire n13981;
    wire n13984;
    wire n13987;
    wire n13990;
    wire n13993;
    wire n13996;
    wire n13999;
    wire n14002;
    wire n14005;
    wire n14008;
    wire n14011;
    wire n14014;
    wire n14017;
    wire n14020;
    wire n14023;
    wire n14026;
    wire n14029;
    wire n14031;
    wire n14034;
    wire n14037;
    wire n14040;
    wire n14043;
    wire n14046;
    wire n14049;
    wire n14052;
    wire n14055;
    wire n14058;
    wire n14061;
    wire n14064;
    wire n14067;
    wire n14070;
    wire n14073;
    wire n14076;
    wire n14079;
    wire n14082;
    wire n14085;
    wire n14088;
    wire n14091;
    wire n14094;
    wire n14097;
    wire n14100;
    wire n14103;
    wire n14106;
    wire n14109;
    wire n14113;
    wire n14116;
    wire n14119;
    wire n14122;
    wire n14125;
    wire n14128;
    wire n14131;
    wire n14134;
    wire n14137;
    wire n14140;
    wire n14143;
    wire n14146;
    wire n14149;
    wire n14152;
    wire n14155;
    wire n14158;
    wire n14161;
    wire n14164;
    wire n14167;
    wire n14170;
    wire n14173;
    wire n14176;
    wire n14179;
    wire n14181;
    wire n14184;
    wire n14187;
    wire n14190;
    wire n14193;
    wire n14196;
    wire n14199;
    wire n14202;
    wire n14205;
    wire n14208;
    wire n14211;
    wire n14214;
    wire n14217;
    wire n14220;
    wire n14223;
    wire n14226;
    wire n14229;
    wire n14232;
    wire n14235;
    wire n14238;
    wire n14241;
    wire n14244;
    wire n14247;
    wire n14250;
    wire n14254;
    wire n14257;
    wire n14260;
    wire n14263;
    wire n14266;
    wire n14269;
    wire n14272;
    wire n14275;
    wire n14278;
    wire n14281;
    wire n14284;
    wire n14287;
    wire n14290;
    wire n14293;
    wire n14296;
    wire n14299;
    wire n14302;
    wire n14305;
    wire n14308;
    wire n14311;
    wire n14313;
    wire n14316;
    wire n14319;
    wire n14322;
    wire n14325;
    wire n14328;
    wire n14331;
    wire n14334;
    wire n14337;
    wire n14340;
    wire n14343;
    wire n14346;
    wire n14349;
    wire n14352;
    wire n14355;
    wire n14358;
    wire n14361;
    wire n14364;
    wire n14367;
    wire n14370;
    wire n14373;
    wire n14377;
    wire n14380;
    wire n14383;
    wire n14386;
    wire n14389;
    wire n14392;
    wire n14395;
    wire n14398;
    wire n14401;
    wire n14404;
    wire n14407;
    wire n14410;
    wire n14413;
    wire n14416;
    wire n14419;
    wire n14422;
    wire n14425;
    wire n14427;
    wire n14430;
    wire n14433;
    wire n14436;
    wire n14439;
    wire n14442;
    wire n14445;
    wire n14448;
    wire n14451;
    wire n14454;
    wire n14457;
    wire n14460;
    wire n14463;
    wire n14466;
    wire n14469;
    wire n14472;
    wire n14475;
    wire n14478;
    wire n14482;
    wire n14485;
    wire n14488;
    wire n14491;
    wire n14494;
    wire n14497;
    wire n14500;
    wire n14503;
    wire n14506;
    wire n14509;
    wire n14512;
    wire n14515;
    wire n14518;
    wire n14521;
    wire n14523;
    wire n14526;
    wire n14529;
    wire n14532;
    wire n14535;
    wire n14538;
    wire n14541;
    wire n14544;
    wire n14547;
    wire n14550;
    wire n14553;
    wire n14556;
    wire n14559;
    wire n14562;
    wire n14565;
    wire n14569;
    wire n14572;
    wire n14575;
    wire n14578;
    wire n14581;
    wire n14584;
    wire n14587;
    wire n14590;
    wire n14593;
    wire n14596;
    wire n14599;
    wire n14601;
    wire n14604;
    wire n14607;
    wire n14610;
    wire n14613;
    wire n14616;
    wire n14619;
    wire n14622;
    wire n14625;
    wire n14628;
    wire n14631;
    wire n14634;
    wire n14638;
    wire n14641;
    wire n14644;
    wire n14647;
    wire n14650;
    wire n14653;
    wire n14656;
    wire n14659;
    wire n14661;
    wire n14664;
    wire n14667;
    wire n14670;
    wire n14673;
    wire n14676;
    wire n14679;
    wire n14682;
    wire n14685;
    wire n14689;
    wire n14692;
    wire n14695;
    wire n14698;
    wire n14701;
    wire n14704;
    wire n14706;
    wire n14709;
    wire n14712;
    wire n14715;
    wire n14718;
    wire n14721;
    wire n14724;
    wire n14727;
    wire n14731;
    wire n14734;
    wire n14737;
    wire n14740;
    wire n14743;
    wire n14746;
    wire n14749;
    wire n14752;
    wire n14755;
    wire n14758;
    wire n14761;
    wire n14764;
    wire n14767;
    wire n14770;
    wire n14773;
    wire n14776;
    wire n14779;
    wire n14782;
    wire n14785;
    wire n14788;
    wire n14791;
    wire n14794;
    wire n14797;
    wire n14800;
    wire n14803;
    wire n14806;
    wire n14809;
    wire n14812;
    wire n14815;
    wire n14818;
    wire n14821;
    wire n14824;
    wire n14827;
    wire n14830;
    wire n14833;
    wire n14836;
    wire n14839;
    wire n14842;
    wire n14845;
    wire n14848;
    wire n14851;
    wire n14854;
    wire n14857;
    wire n14860;
    wire n14863;
    wire n14865;
    wire n14869;
    wire n14872;
    wire n14875;
    wire n14878;
    wire n14881;
    wire n14884;
    wire n14887;
    wire n14890;
    wire n14893;
    wire n14896;
    wire n14899;
    wire n14902;
    wire n14905;
    wire n14908;
    wire n14911;
    wire n14914;
    wire n14917;
    wire n14920;
    wire n14923;
    wire n14926;
    wire n14929;
    wire n14932;
    wire n14935;
    wire n14938;
    wire n14941;
    wire n14944;
    wire n14947;
    wire n14950;
    wire n14953;
    wire n14956;
    wire n14959;
    wire n14962;
    wire n14965;
    wire n14968;
    wire n14971;
    wire n14974;
    wire n14977;
    wire n14980;
    wire n14983;
    wire n14986;
    wire n14989;
    wire n14992;
    wire n14994;
    wire n14998;
    wire n15001;
    wire n15004;
    wire n15007;
    wire n15010;
    wire n15013;
    wire n15016;
    wire n15019;
    wire n15022;
    wire n15025;
    wire n15028;
    wire n15031;
    wire n15034;
    wire n15037;
    wire n15040;
    wire n15043;
    wire n15046;
    wire n15049;
    wire n15052;
    wire n15055;
    wire n15058;
    wire n15061;
    wire n15064;
    wire n15067;
    wire n15070;
    wire n15073;
    wire n15076;
    wire n15079;
    wire n15082;
    wire n15085;
    wire n15088;
    wire n15091;
    wire n15094;
    wire n15097;
    wire n15100;
    wire n15103;
    wire n15106;
    wire n15109;
    wire n15111;
    wire n15114;
    wire n15117;
    wire n15120;
    wire n15123;
    wire n15126;
    wire n15129;
    wire n15132;
    wire n15135;
    wire n15138;
    wire n15141;
    wire n15144;
    wire n15147;
    wire n15150;
    wire n15153;
    wire n15156;
    wire n15159;
    wire n15162;
    wire n15165;
    wire n15168;
    wire n15171;
    wire n15174;
    wire n15177;
    wire n15180;
    wire n15183;
    wire n15186;
    wire n15189;
    wire n15192;
    wire n15195;
    wire n15198;
    wire n15201;
    wire n15204;
    wire n15207;
    wire n15210;
    wire n15213;
    wire n15216;
    wire n15219;
    wire n15222;
    wire n15225;
    wire n15229;
    wire n15231;
    wire n15234;
    wire n15237;
    wire n15240;
    wire n15243;
    wire n15246;
    wire n15249;
    wire n15252;
    wire n15255;
    wire n15258;
    wire n15261;
    wire n15264;
    wire n15267;
    wire n15270;
    wire n15273;
    wire n15276;
    wire n15279;
    wire n15282;
    wire n15285;
    wire n15288;
    wire n15291;
    wire n15294;
    wire n15297;
    wire n15300;
    wire n15303;
    wire n15306;
    wire n15309;
    wire n15312;
    wire n15315;
    wire n15318;
    wire n15321;
    wire n15324;
    wire n15327;
    wire n15330;
    wire n15333;
    wire n15336;
    wire n15340;
    wire n15342;
    wire n15345;
    wire n15348;
    wire n15351;
    wire n15354;
    wire n15357;
    wire n15360;
    wire n15363;
    wire n15366;
    wire n15369;
    wire n15372;
    wire n15375;
    wire n15378;
    wire n15381;
    wire n15384;
    wire n15387;
    wire n15390;
    wire n15393;
    wire n15396;
    wire n15399;
    wire n15402;
    wire n15405;
    wire n15408;
    wire n15411;
    wire n15414;
    wire n15417;
    wire n15420;
    wire n15423;
    wire n15426;
    wire n15429;
    wire n15432;
    wire n15435;
    wire n15438;
    wire n15442;
    wire n15444;
    wire n15447;
    wire n15450;
    wire n15453;
    wire n15456;
    wire n15459;
    wire n15462;
    wire n15465;
    wire n15468;
    wire n15471;
    wire n15474;
    wire n15477;
    wire n15480;
    wire n15483;
    wire n15486;
    wire n15489;
    wire n15492;
    wire n15495;
    wire n15498;
    wire n15501;
    wire n15504;
    wire n15507;
    wire n15510;
    wire n15513;
    wire n15516;
    wire n15519;
    wire n15522;
    wire n15525;
    wire n15528;
    wire n15531;
    wire n15535;
    wire n15537;
    wire n15540;
    wire n15543;
    wire n15546;
    wire n15549;
    wire n15552;
    wire n15555;
    wire n15558;
    wire n15561;
    wire n15564;
    wire n15567;
    wire n15570;
    wire n15573;
    wire n15576;
    wire n15579;
    wire n15582;
    wire n15585;
    wire n15588;
    wire n15591;
    wire n15594;
    wire n15597;
    wire n15600;
    wire n15603;
    wire n15606;
    wire n15609;
    wire n15612;
    wire n15615;
    wire n15619;
    wire n15621;
    wire n15624;
    wire n15627;
    wire n15630;
    wire n15633;
    wire n15636;
    wire n15639;
    wire n15642;
    wire n15645;
    wire n15648;
    wire n15651;
    wire n15654;
    wire n15657;
    wire n15660;
    wire n15663;
    wire n15666;
    wire n15669;
    wire n15672;
    wire n15675;
    wire n15678;
    wire n15681;
    wire n15684;
    wire n15687;
    wire n15690;
    wire n15694;
    wire n15696;
    wire n15699;
    wire n15702;
    wire n15705;
    wire n15708;
    wire n15711;
    wire n15714;
    wire n15717;
    wire n15720;
    wire n15723;
    wire n15726;
    wire n15729;
    wire n15732;
    wire n15735;
    wire n15738;
    wire n15741;
    wire n15744;
    wire n15747;
    wire n15750;
    wire n15753;
    wire n15756;
    wire n15760;
    wire n15762;
    wire n15765;
    wire n15768;
    wire n15771;
    wire n15774;
    wire n15777;
    wire n15780;
    wire n15783;
    wire n15786;
    wire n15789;
    wire n15792;
    wire n15795;
    wire n15798;
    wire n15801;
    wire n15804;
    wire n15807;
    wire n15810;
    wire n15813;
    wire n15817;
    wire n15819;
    wire n15822;
    wire n15825;
    wire n15828;
    wire n15831;
    wire n15834;
    wire n15837;
    wire n15840;
    wire n15843;
    wire n15846;
    wire n15849;
    wire n15852;
    wire n15855;
    wire n15858;
    wire n15861;
    wire n15865;
    wire n15867;
    wire n15870;
    wire n15873;
    wire n15876;
    wire n15879;
    wire n15882;
    wire n15885;
    wire n15888;
    wire n15891;
    wire n15894;
    wire n15897;
    wire n15900;
    wire n15904;
    wire n15906;
    wire n15909;
    wire n15912;
    wire n15915;
    wire n15918;
    wire n15921;
    wire n15924;
    wire n15927;
    wire n15930;
    wire n15933;
    wire n15936;
    wire n15939;
    wire n15942;
    wire n15945;
    wire n15948;
    wire n15951;
    wire n15954;
    wire n15957;
    wire n15960;
    wire n15964;
    wire n15966;
    wire n15969;
    wire n15972;
    wire n15975;
    wire n15979;
    wire n15982;
    wire n15985;
    wire n15988;
    wire n15991;
    wire n15994;
    wire n15997;
    wire n16000;
    wire n16003;
    wire n16006;
    wire n16009;
    wire n16012;
    wire n16015;
    wire n16018;
    wire n16021;
    wire n16024;
    wire n16027;
    wire n16030;
    wire n16033;
    wire n16036;
    wire n16039;
    wire n16042;
    wire n16045;
    wire n16048;
    wire n16051;
    wire n16054;
    wire n16057;
    wire n16060;
    wire n16063;
    wire n16066;
    wire n16069;
    wire n16072;
    wire n16075;
    wire n16078;
    wire n16081;
    wire n16084;
    wire n16087;
    wire n16090;
    wire n16093;
    wire n16096;
    wire n16099;
    wire n16102;
    wire n16105;
    wire n16108;
    wire n16111;
    wire n16113;
    wire n16117;
    wire n16120;
    wire n16123;
    wire n16126;
    wire n16129;
    wire n16132;
    wire n16135;
    wire n16138;
    wire n16141;
    wire n16144;
    wire n16147;
    wire n16150;
    wire n16153;
    wire n16156;
    wire n16159;
    wire n16162;
    wire n16165;
    wire n16168;
    wire n16171;
    wire n16174;
    wire n16177;
    wire n16180;
    wire n16183;
    wire n16186;
    wire n16189;
    wire n16192;
    wire n16195;
    wire n16198;
    wire n16201;
    wire n16204;
    wire n16207;
    wire n16210;
    wire n16213;
    wire n16216;
    wire n16219;
    wire n16222;
    wire n16225;
    wire n16228;
    wire n16231;
    wire n16234;
    wire n16237;
    wire n16240;
    wire n16242;
    wire n16245;
    wire n16248;
    wire n16251;
    wire n16254;
    wire n16257;
    wire n16260;
    wire n16263;
    wire n16266;
    wire n16269;
    wire n16272;
    wire n16275;
    wire n16278;
    wire n16281;
    wire n16284;
    wire n16287;
    wire n16290;
    wire n16293;
    wire n16296;
    wire n16299;
    wire n16302;
    wire n16305;
    wire n16308;
    wire n16311;
    wire n16314;
    wire n16317;
    wire n16320;
    wire n16323;
    wire n16326;
    wire n16329;
    wire n16332;
    wire n16335;
    wire n16338;
    wire n16341;
    wire n16344;
    wire n16347;
    wire n16350;
    wire n16353;
    wire n16356;
    wire n16359;
    wire n16362;
    wire n16366;
    wire n16369;
    wire n16372;
    wire n16375;
    wire n16378;
    wire n16381;
    wire n16384;
    wire n16387;
    wire n16390;
    wire n16393;
    wire n16396;
    wire n16399;
    wire n16402;
    wire n16405;
    wire n16408;
    wire n16411;
    wire n16414;
    wire n16417;
    wire n16420;
    wire n16423;
    wire n16426;
    wire n16429;
    wire n16432;
    wire n16435;
    wire n16438;
    wire n16441;
    wire n16444;
    wire n16447;
    wire n16450;
    wire n16453;
    wire n16456;
    wire n16459;
    wire n16462;
    wire n16465;
    wire n16468;
    wire n16471;
    wire n16474;
    wire n16477;
    wire n16480;
    wire n16483;
    wire n16486;
    wire n16489;
    wire n16492;
    wire n16495;
    wire n16498;
    wire n16501;
    wire n16504;
    wire n16507;
    wire n16510;
    wire n16513;
    wire n16516;
    wire n16519;
    wire n16522;
    wire n16525;
    wire n16528;
    wire n16531;
    wire n16534;
    wire n16537;
    wire n16540;
    wire n16543;
    wire n16546;
    wire n16549;
    wire n16552;
    wire n16555;
    wire n16558;
    wire n16561;
    wire n16564;
    wire n16567;
    wire n16570;
    wire n16573;
    wire n16576;
    wire n16579;
    wire n16582;
    wire n16585;
    wire n16588;
    wire n16591;
    wire n16594;
    wire n16597;
    wire n16600;
    wire n16603;
    wire n16606;
    wire n16609;
    wire n16612;
    wire n16615;
    wire n16618;
    wire n16621;
    wire n16624;
    wire n16627;
    wire n16630;
    wire n16633;
    wire n16636;
    wire n16639;
    wire n16642;
    wire n16645;
    wire n16648;
    wire n16651;
    wire n16654;
    wire n16657;
    wire n16660;
    wire n16663;
    wire n16666;
    wire n16669;
    wire n16672;
    wire n16675;
    wire n16678;
    wire n16681;
    wire n16684;
    wire n16687;
    wire n16690;
    wire n16693;
    wire n16696;
    wire n16699;
    wire n16702;
    wire n16705;
    wire n16708;
    wire n16711;
    wire n16714;
    wire n16717;
    wire n16720;
    wire n16723;
    wire n16726;
    wire n16729;
    wire n16732;
    wire n16735;
    wire n16738;
    wire n16741;
    wire n16744;
    wire n16747;
    wire n16750;
    wire n16753;
    wire n16756;
    wire n16759;
    wire n16762;
    wire n16765;
    wire n16768;
    wire n16771;
    wire n16774;
    wire n16777;
    wire n16780;
    wire n16783;
    wire n16786;
    wire n16789;
    wire n16792;
    wire n16795;
    wire n16798;
    wire n16801;
    wire n16804;
    wire n16807;
    wire n16810;
    wire n16813;
    wire n16816;
    wire n16819;
    wire n16822;
    wire n16825;
    wire n16828;
    wire n16831;
    wire n16834;
    wire n16837;
    wire n16840;
    wire n16843;
    wire n16846;
    wire n16849;
    wire n16852;
    wire n16855;
    wire n16858;
    wire n16861;
    wire n16864;
    wire n16867;
    wire n16870;
    wire n16873;
    wire n16876;
    wire n16879;
    wire n16882;
    wire n16885;
    wire n16888;
    wire n16891;
    wire n16894;
    wire n16897;
    wire n16900;
    wire n16903;
    wire n16906;
    wire n16909;
    wire n16912;
    wire n16915;
    wire n16918;
    wire n16921;
    wire n16924;
    wire n16927;
    wire n16930;
    wire n16933;
    wire n16936;
    wire n16939;
    wire n16942;
    wire n16945;
    wire n16948;
    wire n16951;
    wire n16954;
    wire n16957;
    wire n16960;
    wire n16963;
    wire n16966;
    wire n16969;
    wire n16972;
    wire n16975;
    wire n16978;
    wire n16981;
    wire n16984;
    wire n16987;
    wire n16990;
    wire n16993;
    wire n16996;
    wire n16999;
    wire n17002;
    wire n17005;
    wire n17008;
    wire n17011;
    wire n17014;
    wire n17017;
    wire n17020;
    wire n17023;
    wire n17026;
    wire n17029;
    wire n17032;
    wire n17035;
    wire n17038;
    wire n17041;
    wire n17044;
    wire n17047;
    wire n17050;
    wire n17053;
    wire n17056;
    wire n17058;
    wire n17061;
    wire n17064;
    wire n17067;
    wire n17070;
    wire n17073;
    wire n17077;
    wire n17079;
    wire n17082;
    wire n17086;
    wire n17089;
    wire n17092;
    wire n17095;
    wire n17098;
    wire n17101;
    wire n17104;
    wire n17107;
    wire n17110;
    wire n17113;
    wire n17116;
    wire n17119;
    wire n17122;
    wire n17125;
    wire n17128;
    wire n17131;
    wire n17134;
    wire n17137;
    wire n17140;
    wire n17143;
    wire n17146;
    wire n17149;
    wire n17152;
    wire n17155;
    wire n17158;
    wire n17161;
    wire n17164;
    wire n17167;
    wire n17170;
    wire n17173;
    wire n17176;
    wire n17179;
    wire n17182;
    wire n17185;
    wire n17188;
    wire n17191;
    wire n17194;
    wire n17197;
    wire n17200;
    wire n17203;
    wire n17206;
    wire n17209;
    wire n17212;
    wire n17215;
    wire n17218;
    wire n17221;
    wire n17224;
    wire n17227;
    wire n17230;
    wire n17233;
    wire n17236;
    wire n17239;
    wire n17242;
    wire n17245;
    wire n17248;
    wire n17251;
    wire n17254;
    wire n17257;
    wire n17260;
    wire n17263;
    wire n17266;
    wire n17269;
    wire n17272;
    wire n17275;
    wire n17278;
    wire n17281;
    wire n17284;
    wire n17287;
    wire n17290;
    wire n17293;
    wire n17296;
    wire n17299;
    wire n17302;
    wire n17305;
    wire n17308;
    wire n17311;
    wire n17314;
    wire n17317;
    wire n17320;
    wire n17323;
    wire n17326;
    wire n17329;
    wire n17332;
    wire n17335;
    wire n17338;
    wire n17341;
    wire n17344;
    wire n17347;
    wire n17350;
    wire n17353;
    wire n17356;
    wire n17359;
    wire n17362;
    wire n17365;
    wire n17368;
    wire n17371;
    wire n17374;
    wire n17377;
    wire n17380;
    wire n17383;
    wire n17386;
    wire n17389;
    wire n17392;
    wire n17395;
    wire n17398;
    wire n17401;
    wire n17404;
    wire n17407;
    wire n17410;
    wire n17413;
    wire n17416;
    wire n17419;
    wire n17422;
    wire n17425;
    wire n17428;
    wire n17431;
    wire n17434;
    wire n17437;
    wire n17440;
    wire n17443;
    wire n17446;
    wire n17449;
    wire n17452;
    wire n17455;
    wire n17458;
    wire n17461;
    wire n17464;
    wire n17467;
    wire n17470;
    wire n17473;
    wire n17476;
    wire n17479;
    wire n17482;
    wire n17485;
    wire n17488;
    wire n17491;
    wire n17494;
    wire n17497;
    wire n17500;
    wire n17503;
    wire n17506;
    wire n17509;
    wire n17512;
    wire n17515;
    wire n17518;
    wire n17521;
    wire n17524;
    wire n17527;
    wire n17530;
    wire n17533;
    wire n17536;
    wire n17539;
    wire n17542;
    wire n17545;
    wire n17548;
    wire n17551;
    wire n17554;
    wire n17557;
    wire n17560;
    wire n17563;
    wire n17566;
    wire n17569;
    wire n17572;
    wire n17575;
    wire n17578;
    wire n17581;
    wire n17584;
    wire n17587;
    wire n17590;
    wire n17593;
    wire n17596;
    wire n17599;
    wire n17602;
    wire n17605;
    wire n17608;
    wire n17611;
    wire n17614;
    wire n17617;
    wire n17620;
    wire n17623;
    wire n17626;
    wire n17629;
    wire n17632;
    wire n17635;
    wire n17638;
    wire n17641;
    wire n17644;
    wire n17647;
    wire n17650;
    wire n17653;
    wire n17656;
    wire n17659;
    wire n17662;
    wire n17665;
    wire n17668;
    wire n17671;
    wire n17674;
    wire n17677;
    wire n17680;
    wire n17683;
    wire n17686;
    wire n17689;
    wire n17692;
    wire n17695;
    wire n17698;
    wire n17701;
    wire n17704;
    wire n17707;
    wire n17710;
    wire n17713;
    wire n17716;
    wire n17719;
    wire n17722;
    wire n17725;
    wire n17728;
    wire n17731;
    wire n17734;
    wire n17737;
    wire n17740;
    wire n17743;
    wire n17746;
    wire n17749;
    wire n17752;
    wire n17755;
    wire n17758;
    wire n17761;
    wire n17764;
    wire n17767;
    wire n17770;
    wire n17773;
    wire n17776;
    wire n17779;
    wire n17782;
    wire n17785;
    wire n17788;
    wire n17791;
    wire n17794;
    wire n17797;
    wire n17800;
    wire n17803;
    wire n17806;
    wire n17809;
    wire n17812;
    wire n17815;
    wire n17818;
    wire n17821;
    wire n17824;
    wire n17827;
    wire n17830;
    wire n17833;
    wire n17836;
    wire n17839;
    wire n17842;
    wire n17845;
    wire n17848;
    wire n17851;
    wire n17854;
    wire n17857;
    wire n17860;
    wire n17863;
    wire n17866;
    wire n17869;
    wire n17872;
    wire n17875;
    wire n17878;
    wire n17881;
    wire n17884;
    wire n17887;
    wire n17890;
    wire n17893;
    wire n17896;
    wire n17899;
    wire n17902;
    wire n17905;
    wire n17908;
    wire n17911;
    wire n17914;
    wire n17917;
    wire n17920;
    wire n17923;
    wire n17926;
    wire n17929;
    wire n17932;
    wire n17935;
    wire n17938;
    wire n17941;
    wire n17944;
    wire n17947;
    wire n17950;
    wire n17953;
    wire n17956;
    wire n17959;
    wire n17962;
    wire n17965;
    wire n17968;
    wire n17971;
    wire n17974;
    wire n17977;
    wire n17980;
    wire n17983;
    wire n17986;
    wire n17989;
    wire n17992;
    wire n17995;
    wire n17998;
    wire n18001;
    wire n18004;
    wire n18007;
    wire n18010;
    wire n18013;
    wire n18016;
    wire n18019;
    wire n18022;
    wire n18025;
    wire n18028;
    wire n18031;
    wire n18034;
    wire n18037;
    wire n18040;
    wire n18043;
    wire n18046;
    wire n18049;
    wire n18052;
    wire n18055;
    wire n18058;
    wire n18061;
    wire n18064;
    wire n18067;
    wire n18070;
    wire n18073;
    wire n18076;
    wire n18079;
    wire n18082;
    wire n18085;
    wire n18088;
    wire n18091;
    wire n18094;
    wire n18097;
    wire n18100;
    wire n18103;
    wire n18106;
    wire n18109;
    wire n18112;
    wire n18115;
    wire n18118;
    wire n18121;
    wire n18124;
    wire n18127;
    wire n18130;
    wire n18133;
    wire n18136;
    wire n18139;
    wire n18142;
    wire n18145;
    wire n18148;
    wire n18151;
    wire n18154;
    wire n18157;
    wire n18160;
    wire n18163;
    wire n18166;
    wire n18169;
    wire n18172;
    wire n18175;
    wire n18177;
    wire n18180;
    wire n18183;
    wire n18187;
    wire n18190;
    wire n18193;
    wire n18196;
    wire n18199;
    wire n18202;
    wire n18205;
    wire n18208;
    wire n18211;
    wire n18214;
    wire n18217;
    wire n18220;
    wire n18223;
    wire n18226;
    wire n18229;
    wire n18232;
    wire n18235;
    wire n18238;
    wire n18241;
    wire n18244;
    wire n18247;
    wire n18250;
    wire n18253;
    wire n18256;
    wire n18259;
    wire n18262;
    wire n18265;
    wire n18268;
    wire n18271;
    wire n18274;
    wire n18277;
    wire n18280;
    wire n18283;
    wire n18286;
    wire n18289;
    wire n18292;
    wire n18295;
    wire n18298;
    wire n18301;
    wire n18304;
    wire n18307;
    wire n18310;
    wire n18313;
    wire n18316;
    wire n18319;
    wire n18322;
    wire n18325;
    wire n18327;
    wire n18331;
    wire n18334;
    wire n18337;
    wire n18340;
    wire n18343;
    wire n18346;
    wire n18349;
    wire n18352;
    wire n18355;
    wire n18358;
    wire n18361;
    wire n18364;
    wire n18367;
    wire n18370;
    wire n18373;
    wire n18376;
    wire n18379;
    wire n18382;
    wire n18385;
    wire n18388;
    wire n18391;
    wire n18394;
    wire n18397;
    wire n18400;
    wire n18403;
    wire n18406;
    wire n18409;
    wire n18412;
    wire n18415;
    wire n18418;
    wire n18421;
    wire n18424;
    wire n18427;
    wire n18430;
    wire n18433;
    wire n18436;
    wire n18439;
    wire n18442;
    wire n18445;
    wire n18448;
    wire n18451;
    wire n18454;
    wire n18457;
    wire n18460;
    wire n18463;
    wire n18466;
    wire n18469;
    wire n18472;
    wire n18475;
    wire n18478;
    wire n18481;
    wire n18484;
    wire n18487;
    wire n18490;
    wire n18493;
    wire n18496;
    wire n18499;
    wire n18502;
    wire n18505;
    wire n18508;
    wire n18511;
    wire n18514;
    wire n18517;
    wire n18520;
    wire n18523;
    wire n18526;
    wire n18529;
    wire n18532;
    wire n18535;
    wire n18538;
    wire n18541;
    wire n18544;
    wire n18547;
    wire n18550;
    wire n18553;
    wire n18556;
    wire n18559;
    wire n18562;
    wire n18565;
    wire n18568;
    wire n18571;
    wire n18574;
    wire n18577;
    wire n18580;
    wire n18583;
    wire n18586;
    wire n18589;
    wire n18592;
    wire n18595;
    wire n18598;
    wire n18601;
    wire n18604;
    wire n18607;
    wire n18610;
    wire n18613;
    wire n18616;
    wire n18619;
    wire n18622;
    wire n18625;
    wire n18628;
    wire n18631;
    wire n18634;
    wire n18637;
    wire n18640;
    wire n18643;
    wire n18646;
    wire n18649;
    wire n18652;
    wire n18655;
    wire n18658;
    wire n18661;
    wire n18664;
    wire n18667;
    wire n18670;
    wire n18673;
    wire n18676;
    wire n18679;
    wire n18682;
    wire n18685;
    wire n18688;
    wire n18691;
    wire n18694;
    wire n18697;
    wire n18700;
    wire n18703;
    wire n18706;
    wire n18709;
    wire n18712;
    wire n18715;
    wire n18718;
    wire n18721;
    wire n18724;
    wire n18727;
    wire n18730;
    wire n18733;
    wire n18736;
    wire n18739;
    wire n18742;
    wire n18745;
    wire n18748;
    wire n18751;
    wire n18754;
    wire n18757;
    wire n18760;
    wire n18763;
    wire n18766;
    wire n18769;
    wire n18772;
    wire n18775;
    wire n18778;
    wire n18781;
    wire n18784;
    wire n18787;
    wire n18790;
    wire n18793;
    wire n18796;
    wire n18799;
    wire n18802;
    wire n18805;
    wire n18808;
    wire n18811;
    wire n18814;
    wire n18817;
    wire n18820;
    wire n18823;
    wire n18826;
    wire n18829;
    wire n18832;
    wire n18835;
    wire n18838;
    wire n18841;
    wire n18844;
    wire n18847;
    wire n18850;
    wire n18853;
    wire n18856;
    wire n18859;
    wire n18862;
    wire n18865;
    wire n18868;
    wire n18871;
    wire n18874;
    wire n18877;
    wire n18880;
    wire n18883;
    wire n18886;
    wire n18889;
    wire n18892;
    wire n18895;
    wire n18898;
    wire n18901;
    wire n18904;
    wire n18907;
    wire n18910;
    wire n18913;
    wire n18916;
    wire n18919;
    wire n18922;
    wire n18925;
    wire n18928;
    wire n18931;
    wire n18934;
    wire n18937;
    wire n18940;
    wire n18943;
    wire n18946;
    wire n18949;
    wire n18952;
    wire n18955;
    wire n18958;
    wire n18961;
    wire n18964;
    wire n18967;
    wire n18970;
    wire n18973;
    wire n18976;
    wire n18979;
    wire n18982;
    wire n18985;
    wire n18988;
    wire n18991;
    wire n18994;
    wire n18997;
    wire n19000;
    wire n19003;
    wire n19006;
    wire n19009;
    wire n19012;
    wire n19015;
    wire n19018;
    wire n19021;
    wire n19024;
    wire n19027;
    wire n19030;
    wire n19033;
    wire n19036;
    wire n19039;
    wire n19042;
    wire n19045;
    wire n19048;
    wire n19051;
    wire n19054;
    wire n19057;
    wire n19060;
    wire n19063;
    wire n19066;
    wire n19069;
    wire n19072;
    wire n19075;
    wire n19078;
    wire n19081;
    wire n19084;
    wire n19087;
    wire n19090;
    wire n19093;
    wire n19096;
    wire n19099;
    wire n19102;
    wire n19105;
    wire n19108;
    wire n19111;
    wire n19114;
    wire n19117;
    wire n19120;
    wire n19123;
    wire n19126;
    wire n19129;
    wire n19132;
    wire n19135;
    wire n19138;
    wire n19141;
    wire n19144;
    wire n19147;
    wire n19150;
    wire n19153;
    wire n19156;
    wire n19159;
    wire n19162;
    wire n19165;
    wire n19168;
    wire n19171;
    wire n19174;
    wire n19177;
    wire n19180;
    wire n19183;
    wire n19186;
    wire n19189;
    wire n19192;
    wire n19195;
    wire n19198;
    wire n19201;
    wire n19204;
    wire n19207;
    wire n19210;
    wire n19213;
    wire n19216;
    wire n19219;
    wire n19222;
    wire n19225;
    wire n19228;
    wire n19231;
    wire n19234;
    wire n19237;
    wire n19240;
    wire n19243;
    wire n19246;
    wire n19249;
    wire n19252;
    wire n19255;
    wire n19258;
    wire n19261;
    wire n19264;
    wire n19267;
    wire n19269;
    wire n19272;
    wire n19275;
    wire n19278;
    wire n19282;
    wire n19285;
    wire n19288;
    wire n19291;
    wire n19294;
    wire n19297;
    wire n19300;
    wire n19303;
    wire n19306;
    wire n19309;
    wire n19312;
    wire n19315;
    wire n19318;
    wire n19321;
    wire n19324;
    wire n19327;
    wire n19330;
    wire n19333;
    wire n19336;
    wire n19339;
    wire n19342;
    wire n19345;
    wire n19348;
    wire n19351;
    wire n19354;
    wire n19357;
    wire n19360;
    wire n19363;
    wire n19366;
    wire n19369;
    wire n19372;
    wire n19375;
    wire n19378;
    wire n19381;
    wire n19384;
    wire n19387;
    wire n19390;
    wire n19393;
    wire n19396;
    wire n19399;
    wire n19402;
    wire n19405;
    wire n19408;
    wire n19411;
    wire n19414;
    wire n19417;
    wire n19420;
    wire n19423;
    wire n19426;
    wire n19429;
    wire n19432;
    wire n19435;
    wire n19438;
    wire n19441;
    wire n19444;
    wire n19447;
    wire n19450;
    wire n19453;
    wire n19456;
    wire n19459;
    wire n19462;
    wire n19465;
    wire n19468;
    wire n19471;
    wire n19474;
    wire n19477;
    wire n19480;
    wire n19483;
    wire n19486;
    wire n19489;
    wire n19492;
    wire n19495;
    wire n19498;
    wire n19501;
    wire n19504;
    wire n19507;
    wire n19510;
    wire n19513;
    wire n19516;
    wire n19519;
    wire n19522;
    wire n19525;
    wire n19528;
    wire n19531;
    wire n19534;
    wire n19537;
    wire n19540;
    wire n19543;
    wire n19546;
    wire n19549;
    wire n19552;
    wire n19555;
    wire n19558;
    wire n19561;
    wire n19564;
    wire n19567;
    wire n19570;
    wire n19573;
    wire n19576;
    wire n19579;
    wire n19582;
    wire n19585;
    wire n19588;
    wire n19591;
    wire n19594;
    wire n19597;
    wire n19600;
    wire n19603;
    wire n19606;
    wire n19609;
    wire n19612;
    wire n19615;
    wire n19618;
    wire n19621;
    wire n19624;
    wire n19627;
    wire n19630;
    wire n19633;
    wire n19636;
    wire n19639;
    wire n19642;
    wire n19645;
    wire n19648;
    wire n19651;
    wire n19654;
    wire n19657;
    wire n19660;
    wire n19663;
    wire n19666;
    wire n19669;
    wire n19672;
    wire n19675;
    wire n19678;
    wire n19681;
    wire n19684;
    wire n19687;
    wire n19690;
    wire n19693;
    wire n19696;
    wire n19699;
    wire n19702;
    wire n19705;
    wire n19708;
    wire n19711;
    wire n19714;
    wire n19717;
    wire n19720;
    wire n19723;
    wire n19726;
    wire n19729;
    wire n19732;
    wire n19735;
    wire n19738;
    wire n19741;
    wire n19744;
    wire n19747;
    wire n19750;
    wire n19753;
    wire n19756;
    wire n19759;
    wire n19762;
    wire n19765;
    wire n19768;
    wire n19771;
    wire n19774;
    wire n19777;
    wire n19780;
    wire n19783;
    wire n19786;
    wire n19789;
    wire n19792;
    wire n19795;
    wire n19798;
    wire n19801;
    wire n19804;
    wire n19807;
    wire n19810;
    wire n19813;
    wire n19816;
    wire n19819;
    wire n19822;
    wire n19825;
    wire n19828;
    wire n19831;
    wire n19834;
    wire n19837;
    wire n19840;
    wire n19843;
    wire n19846;
    wire n19849;
    wire n19852;
    wire n19855;
    wire n19858;
    wire n19861;
    wire n19864;
    wire n19867;
    wire n19870;
    wire n19873;
    wire n19876;
    wire n19879;
    wire n19882;
    wire n19885;
    wire n19888;
    wire n19891;
    wire n19894;
    wire n19897;
    wire n19900;
    wire n19903;
    wire n19906;
    wire n19909;
    wire n19912;
    wire n19915;
    wire n19918;
    wire n19921;
    wire n19924;
    wire n19927;
    wire n19930;
    wire n19933;
    wire n19936;
    wire n19939;
    wire n19942;
    wire n19945;
    wire n19948;
    wire n19951;
    wire n19954;
    wire n19957;
    wire n19960;
    wire n19963;
    wire n19966;
    wire n19969;
    wire n19972;
    wire n19975;
    wire n19978;
    wire n19981;
    wire n19984;
    wire n19987;
    wire n19990;
    wire n19993;
    wire n19996;
    wire n19999;
    wire n20002;
    wire n20005;
    wire n20008;
    wire n20011;
    wire n20014;
    wire n20017;
    wire n20020;
    wire n20023;
    wire n20026;
    wire n20029;
    wire n20032;
    wire n20035;
    wire n20038;
    wire n20041;
    wire n20044;
    wire n20047;
    wire n20050;
    wire n20053;
    wire n20056;
    wire n20059;
    wire n20062;
    wire n20065;
    wire n20068;
    wire n20071;
    wire n20074;
    wire n20077;
    wire n20080;
    wire n20083;
    wire n20086;
    wire n20089;
    wire n20092;
    wire n20095;
    wire n20098;
    wire n20101;
    wire n20104;
    wire n20107;
    wire n20110;
    wire n20113;
    wire n20116;
    wire n20119;
    wire n20122;
    wire n20125;
    wire n20128;
    wire n20131;
    wire n20134;
    wire n20137;
    wire n20140;
    wire n20143;
    wire n20146;
    wire n20149;
    wire n20152;
    wire n20155;
    wire n20158;
    wire n20161;
    wire n20164;
    wire n20167;
    wire n20170;
    wire n20173;
    wire n20176;
    wire n20179;
    wire n20182;
    wire n20185;
    wire n20188;
    wire n20191;
    wire n20194;
    wire n20197;
    wire n20200;
    wire n20203;
    wire n20206;
    wire n20209;
    wire n20212;
    wire n20215;
    wire n20218;
    wire n20221;
    wire n20224;
    wire n20227;
    wire n20230;
    wire n20233;
    wire n20236;
    wire n20239;
    wire n20242;
    wire n20245;
    wire n20248;
    wire n20251;
    wire n20254;
    wire n20257;
    wire n20260;
    wire n20263;
    wire n20266;
    wire n20269;
    wire n20272;
    wire n20275;
    wire n20278;
    wire n20281;
    wire n20284;
    wire n20287;
    wire n20290;
    wire n20293;
    wire n20296;
    wire n20299;
    wire n20302;
    wire n20305;
    wire n20308;
    wire n20311;
    wire n20314;
    wire n20317;
    wire n20320;
    wire n20323;
    wire n20326;
    wire n20328;
    wire n20331;
    wire n20334;
    wire n20338;
    wire n20341;
    wire n20344;
    wire n20347;
    wire n20350;
    wire n20353;
    wire n20356;
    wire n20359;
    wire n20362;
    wire n20365;
    wire n20368;
    wire n20371;
    wire n20374;
    wire n20377;
    wire n20380;
    wire n20383;
    wire n20386;
    wire n20389;
    wire n20392;
    wire n20395;
    wire n20398;
    wire n20401;
    wire n20404;
    wire n20407;
    wire n20410;
    wire n20413;
    wire n20416;
    wire n20419;
    wire n20422;
    wire n20425;
    wire n20428;
    wire n20431;
    wire n20434;
    wire n20437;
    wire n20440;
    wire n20443;
    wire n20446;
    wire n20449;
    wire n20452;
    wire n20455;
    wire n20458;
    wire n20461;
    wire n20464;
    wire n20467;
    wire n20470;
    wire n20473;
    wire n20476;
    wire n20479;
    wire n20482;
    wire n20485;
    wire n20488;
    wire n20491;
    wire n20494;
    wire n20497;
    wire n20500;
    wire n20503;
    wire n20506;
    wire n20509;
    wire n20512;
    wire n20515;
    wire n20518;
    wire n20521;
    wire n20524;
    wire n20527;
    wire n20530;
    wire n20533;
    wire n20536;
    wire n20539;
    wire n20542;
    wire n20545;
    wire n20548;
    wire n20551;
    wire n20554;
    wire n20557;
    wire n20560;
    wire n20563;
    wire n20566;
    wire n20569;
    wire n20572;
    wire n20575;
    wire n20578;
    wire n20581;
    wire n20584;
    wire n20587;
    wire n20590;
    wire n20593;
    wire n20596;
    wire n20599;
    wire n20602;
    wire n20605;
    wire n20608;
    wire n20611;
    wire n20614;
    wire n20617;
    wire n20620;
    wire n20623;
    wire n20626;
    wire n20629;
    wire n20632;
    wire n20635;
    wire n20638;
    wire n20641;
    wire n20644;
    wire n20647;
    wire n20650;
    wire n20653;
    wire n20656;
    wire n20659;
    wire n20662;
    wire n20665;
    wire n20668;
    wire n20671;
    wire n20674;
    wire n20677;
    wire n20680;
    wire n20683;
    wire n20686;
    wire n20689;
    wire n20692;
    wire n20695;
    wire n20698;
    wire n20701;
    wire n20704;
    wire n20707;
    wire n20710;
    wire n20713;
    wire n20716;
    wire n20719;
    wire n20722;
    wire n20725;
    wire n20728;
    wire n20731;
    wire n20734;
    wire n20737;
    wire n20740;
    wire n20743;
    wire n20746;
    wire n20749;
    wire n20752;
    wire n20755;
    wire n20758;
    wire n20761;
    wire n20764;
    wire n20767;
    wire n20770;
    wire n20773;
    wire n20776;
    wire n20779;
    wire n20782;
    wire n20785;
    wire n20788;
    wire n20791;
    wire n20794;
    wire n20797;
    wire n20800;
    wire n20803;
    wire n20806;
    wire n20809;
    wire n20812;
    wire n20815;
    wire n20818;
    wire n20821;
    wire n20824;
    wire n20827;
    wire n20830;
    wire n20833;
    wire n20836;
    wire n20839;
    wire n20842;
    wire n20845;
    wire n20848;
    wire n20851;
    wire n20854;
    wire n20857;
    wire n20860;
    wire n20863;
    wire n20866;
    wire n20869;
    wire n20872;
    wire n20875;
    wire n20878;
    wire n20881;
    wire n20884;
    wire n20887;
    wire n20890;
    wire n20893;
    wire n20896;
    wire n20899;
    wire n20902;
    wire n20905;
    wire n20908;
    wire n20911;
    wire n20914;
    wire n20917;
    wire n20920;
    wire n20923;
    wire n20926;
    wire n20929;
    wire n20932;
    wire n20935;
    wire n20938;
    wire n20941;
    wire n20944;
    wire n20947;
    wire n20950;
    wire n20953;
    wire n20956;
    wire n20959;
    wire n20962;
    wire n20965;
    wire n20968;
    wire n20971;
    wire n20974;
    wire n20977;
    wire n20980;
    wire n20983;
    wire n20986;
    wire n20989;
    wire n20992;
    wire n20995;
    wire n20998;
    wire n21001;
    wire n21004;
    wire n21007;
    wire n21010;
    wire n21013;
    wire n21016;
    wire n21019;
    wire n21022;
    wire n21025;
    wire n21028;
    wire n21031;
    wire n21034;
    wire n21037;
    wire n21040;
    wire n21043;
    wire n21046;
    wire n21049;
    wire n21052;
    wire n21055;
    wire n21058;
    wire n21061;
    wire n21064;
    wire n21067;
    wire n21070;
    wire n21073;
    wire n21076;
    wire n21079;
    wire n21082;
    wire n21085;
    wire n21088;
    wire n21091;
    wire n21094;
    wire n21097;
    wire n21100;
    wire n21103;
    wire n21106;
    wire n21109;
    wire n21112;
    wire n21115;
    wire n21118;
    wire n21121;
    wire n21124;
    wire n21127;
    wire n21130;
    wire n21133;
    wire n21136;
    wire n21139;
    wire n21142;
    wire n21145;
    wire n21148;
    wire n21151;
    wire n21154;
    wire n21157;
    wire n21160;
    wire n21163;
    wire n21166;
    wire n21169;
    wire n21172;
    wire n21175;
    wire n21178;
    wire n21181;
    wire n21184;
    wire n21187;
    wire n21190;
    wire n21193;
    wire n21196;
    wire n21199;
    wire n21202;
    wire n21205;
    wire n21208;
    wire n21211;
    wire n21214;
    wire n21217;
    wire n21220;
    wire n21223;
    wire n21226;
    wire n21229;
    wire n21232;
    wire n21235;
    wire n21238;
    wire n21241;
    wire n21244;
    wire n21247;
    wire n21250;
    wire n21253;
    wire n21256;
    wire n21259;
    wire n21262;
    wire n21265;
    wire n21268;
    wire n21271;
    wire n21274;
    wire n21277;
    wire n21280;
    wire n21283;
    wire n21286;
    wire n21289;
    wire n21292;
    wire n21295;
    wire n21298;
    wire n21301;
    wire n21304;
    wire n21307;
    wire n21310;
    wire n21313;
    wire n21316;
    wire n21319;
    wire n21322;
    wire n21325;
    wire n21328;
    wire n21331;
    wire n21334;
    wire n21337;
    wire n21340;
    wire n21343;
    wire n21346;
    wire n21349;
    wire n21352;
    wire n21355;
    wire n21358;
    wire n21361;
    wire n21364;
    wire n21367;
    wire n21370;
    wire n21373;
    wire n21376;
    wire n21379;
    wire n21382;
    wire n21385;
    wire n21388;
    wire n21391;
    wire n21394;
    wire n21397;
    wire n21400;
    wire n21403;
    wire n21406;
    wire n21409;
    wire n21412;
    wire n21415;
    wire n21417;
    wire n21420;
    wire n21423;
    wire n21427;
    wire n21430;
    wire n21433;
    wire n21436;
    wire n21439;
    wire n21442;
    wire n21445;
    wire n21448;
    wire n21451;
    wire n21454;
    wire n21457;
    wire n21460;
    wire n21463;
    wire n21466;
    wire n21469;
    wire n21472;
    wire n21475;
    wire n21478;
    wire n21481;
    wire n21484;
    wire n21487;
    wire n21490;
    wire n21493;
    wire n21496;
    wire n21499;
    wire n21502;
    wire n21505;
    wire n21508;
    wire n21511;
    wire n21514;
    wire n21517;
    wire n21520;
    wire n21523;
    wire n21526;
    wire n21529;
    wire n21532;
    wire n21535;
    wire n21538;
    wire n21541;
    wire n21544;
    wire n21547;
    wire n21550;
    wire n21553;
    wire n21556;
    wire n21559;
    wire n21562;
    wire n21565;
    wire n21568;
    wire n21571;
    wire n21573;
    wire n21577;
    wire n21580;
    wire n21583;
    wire n21586;
    wire n21589;
    wire n21592;
    wire n21595;
    wire n21598;
    wire n21601;
    wire n21604;
    wire n21607;
    wire n21610;
    wire n21613;
    wire n21616;
    wire n21619;
    wire n21622;
    wire n21625;
    wire n21628;
    wire n21631;
    wire n21634;
    wire n21637;
    wire n21640;
    wire n21643;
    wire n21646;
    wire n21649;
    wire n21652;
    wire n21655;
    wire n21658;
    wire n21661;
    wire n21664;
    wire n21667;
    wire n21670;
    wire n21673;
    wire n21676;
    wire n21679;
    wire n21682;
    wire n21685;
    wire n21688;
    wire n21691;
    wire n21694;
    wire n21697;
    wire n21700;
    wire n21703;
    wire n21706;
    wire n21709;
    wire n21712;
    wire n21715;
    wire n21718;
    wire n21721;
    wire n21724;
    wire n21727;
    wire n21730;
    wire n21733;
    wire n21736;
    wire n21739;
    wire n21742;
    wire n21745;
    wire n21748;
    wire n21751;
    wire n21754;
    wire n21757;
    wire n21760;
    wire n21763;
    wire n21766;
    wire n21769;
    wire n21772;
    wire n21775;
    wire n21778;
    wire n21781;
    wire n21784;
    wire n21787;
    wire n21790;
    wire n21793;
    wire n21796;
    wire n21799;
    wire n21802;
    wire n21805;
    wire n21808;
    wire n21811;
    wire n21814;
    wire n21817;
    wire n21820;
    wire n21823;
    wire n21826;
    wire n21829;
    wire n21832;
    wire n21835;
    wire n21838;
    wire n21841;
    wire n21844;
    wire n21847;
    wire n21850;
    wire n21853;
    wire n21856;
    wire n21859;
    wire n21862;
    wire n21865;
    wire n21868;
    wire n21871;
    wire n21874;
    wire n21877;
    wire n21880;
    wire n21883;
    wire n21886;
    wire n21889;
    wire n21892;
    wire n21895;
    wire n21898;
    wire n21901;
    wire n21904;
    wire n21907;
    wire n21910;
    wire n21913;
    wire n21916;
    wire n21919;
    wire n21922;
    wire n21925;
    wire n21928;
    wire n21931;
    wire n21934;
    wire n21937;
    wire n21940;
    wire n21943;
    wire n21946;
    wire n21949;
    wire n21952;
    wire n21955;
    wire n21958;
    wire n21961;
    wire n21964;
    wire n21967;
    wire n21970;
    wire n21973;
    wire n21976;
    wire n21979;
    wire n21982;
    wire n21985;
    wire n21988;
    wire n21991;
    wire n21994;
    wire n21997;
    wire n22000;
    wire n22003;
    wire n22006;
    wire n22009;
    wire n22012;
    wire n22015;
    wire n22018;
    wire n22021;
    wire n22024;
    wire n22027;
    wire n22030;
    wire n22033;
    wire n22036;
    wire n22039;
    wire n22042;
    wire n22045;
    wire n22048;
    wire n22051;
    wire n22054;
    wire n22057;
    wire n22060;
    wire n22063;
    wire n22066;
    wire n22069;
    wire n22072;
    wire n22075;
    wire n22078;
    wire n22081;
    wire n22084;
    wire n22087;
    wire n22090;
    wire n22093;
    wire n22096;
    wire n22099;
    wire n22102;
    wire n22105;
    wire n22108;
    wire n22111;
    wire n22114;
    wire n22117;
    wire n22120;
    wire n22123;
    wire n22126;
    wire n22129;
    wire n22132;
    wire n22135;
    wire n22138;
    wire n22141;
    wire n22144;
    wire n22147;
    wire n22150;
    wire n22153;
    wire n22156;
    wire n22159;
    wire n22162;
    wire n22165;
    wire n22168;
    wire n22171;
    wire n22174;
    wire n22177;
    wire n22180;
    wire n22183;
    wire n22186;
    wire n22189;
    wire n22192;
    wire n22195;
    wire n22198;
    wire n22201;
    wire n22204;
    wire n22207;
    wire n22210;
    wire n22213;
    wire n22216;
    wire n22219;
    wire n22222;
    wire n22225;
    wire n22228;
    wire n22231;
    wire n22234;
    wire n22237;
    wire n22240;
    wire n22243;
    wire n22246;
    wire n22249;
    wire n22252;
    wire n22255;
    wire n22258;
    wire n22261;
    wire n22264;
    wire n22267;
    wire n22270;
    wire n22273;
    wire n22276;
    wire n22279;
    wire n22282;
    wire n22285;
    wire n22288;
    wire n22291;
    wire n22294;
    wire n22297;
    wire n22300;
    wire n22303;
    wire n22306;
    wire n22309;
    wire n22312;
    wire n22315;
    wire n22318;
    wire n22321;
    wire n22324;
    wire n22327;
    wire n22330;
    wire n22333;
    wire n22336;
    wire n22339;
    wire n22342;
    wire n22345;
    wire n22348;
    wire n22351;
    wire n22354;
    wire n22357;
    wire n22360;
    wire n22363;
    wire n22366;
    wire n22369;
    wire n22372;
    wire n22375;
    wire n22378;
    wire n22381;
    wire n22384;
    wire n22387;
    wire n22390;
    wire n22393;
    wire n22396;
    wire n22399;
    wire n22402;
    wire n22405;
    wire n22408;
    wire n22411;
    wire n22414;
    wire n22417;
    wire n22420;
    wire n22423;
    wire n22426;
    wire n22429;
    wire n22432;
    wire n22435;
    wire n22438;
    wire n22441;
    wire n22444;
    wire n22447;
    wire n22450;
    wire n22453;
    wire n22456;
    wire n22459;
    wire n22462;
    wire n22465;
    wire n22468;
    wire n22471;
    wire n22474;
    wire n22477;
    wire n22480;
    wire n22483;
    wire n22486;
    wire n22489;
    wire n22492;
    wire n22495;
    wire n22498;
    wire n22501;
    wire n22504;
    wire n22507;
    wire n22510;
    wire n22513;
    wire n22516;
    wire n22519;
    wire n22522;
    wire n22525;
    wire n22528;
    wire n22531;
    wire n22534;
    wire n22537;
    wire n22540;
    wire n22543;
    wire n22546;
    wire n22549;
    wire n22552;
    wire n22555;
    wire n22558;
    wire n22561;
    wire n22564;
    wire n22567;
    wire n22570;
    wire n22573;
    wire n22576;
    wire n22579;
    wire n22582;
    wire n22585;
    wire n22588;
    wire n22591;
    wire n22593;
    wire n22596;
    wire n22599;
    wire n22603;
    wire n22605;
    wire n22608;
    wire n22611;
    wire n22614;
    wire n22617;
    wire n22620;
    wire n22623;
    wire n22626;
    wire n22629;
    wire n22633;
    wire n22636;
    wire n22639;
    wire n22642;
    wire n22645;
    wire n22648;
    wire n22651;
    wire n22654;
    wire n22657;
    wire n22660;
    wire n22663;
    wire n22666;
    wire n22669;
    wire n22672;
    wire n22675;
    wire n22678;
    wire n22681;
    wire n22684;
    wire n22687;
    wire n22690;
    wire n22693;
    wire n22696;
    wire n22699;
    wire n22702;
    wire n22705;
    wire n22708;
    wire n22711;
    wire n22714;
    wire n22717;
    wire n22720;
    wire n22723;
    wire n22726;
    wire n22729;
    wire n22732;
    wire n22735;
    wire n22738;
    wire n22741;
    wire n22744;
    wire n22747;
    wire n22750;
    wire n22753;
    wire n22756;
    wire n22759;
    wire n22762;
    wire n22765;
    wire n22768;
    wire n22771;
    wire n22774;
    wire n22777;
    wire n22780;
    wire n22783;
    wire n22786;
    wire n22789;
    wire n22792;
    wire n22795;
    wire n22798;
    wire n22801;
    wire n22804;
    wire n22807;
    wire n22810;
    wire n22813;
    wire n22816;
    wire n22819;
    wire n22822;
    wire n22825;
    wire n22828;
    wire n22831;
    wire n22834;
    wire n22837;
    wire n22840;
    wire n22843;
    wire n22846;
    wire n22849;
    wire n22852;
    wire n22855;
    wire n22858;
    wire n22861;
    wire n22864;
    wire n22867;
    wire n22870;
    wire n22873;
    wire n22876;
    wire n22879;
    wire n22882;
    wire n22885;
    wire n22888;
    wire n22891;
    wire n22894;
    wire n22897;
    wire n22900;
    wire n22903;
    wire n22906;
    wire n22909;
    wire n22912;
    wire n22915;
    wire n22918;
    wire n22921;
    wire n22924;
    wire n22927;
    wire n22930;
    wire n22933;
    wire n22936;
    wire n22939;
    wire n22942;
    wire n22945;
    wire n22948;
    wire n22951;
    wire n22954;
    wire n22957;
    wire n22960;
    wire n22963;
    wire n22966;
    wire n22969;
    wire n22972;
    wire n22975;
    wire n22978;
    wire n22981;
    wire n22984;
    wire n22987;
    wire n22990;
    wire n22993;
    wire n22996;
    wire n22999;
    wire n23002;
    wire n23005;
    wire n23008;
    wire n23011;
    wire n23014;
    wire n23017;
    wire n23020;
    wire n23023;
    wire n23026;
    wire n23029;
    wire n23032;
    wire n23035;
    wire n23038;
    wire n23041;
    wire n23044;
    wire n23047;
    wire n23050;
    wire n23053;
    wire n23056;
    wire n23059;
    wire n23062;
    wire n23065;
    wire n23068;
    wire n23071;
    wire n23074;
    wire n23077;
    wire n23080;
    wire n23083;
    wire n23086;
    wire n23089;
    wire n23092;
    wire n23095;
    wire n23098;
    wire n23101;
    wire n23104;
    wire n23107;
    wire n23110;
    wire n23113;
    wire n23116;
    wire n23119;
    wire n23122;
    wire n23125;
    wire n23128;
    wire n23131;
    wire n23134;
    wire n23137;
    wire n23140;
    wire n23143;
    wire n23146;
    wire n23149;
    wire n23152;
    wire n23155;
    wire n23158;
    wire n23161;
    wire n23164;
    wire n23167;
    wire n23170;
    wire n23173;
    wire n23176;
    wire n23179;
    wire n23182;
    wire n23185;
    wire n23188;
    wire n23191;
    wire n23194;
    wire n23197;
    wire n23200;
    wire n23203;
    wire n23206;
    wire n23209;
    wire n23212;
    wire n23215;
    wire n23218;
    wire n23221;
    wire n23224;
    wire n23227;
    wire n23230;
    wire n23233;
    wire n23236;
    wire n23239;
    wire n23242;
    wire n23245;
    wire n23248;
    wire n23251;
    wire n23254;
    wire n23257;
    wire n23260;
    wire n23263;
    wire n23266;
    wire n23269;
    wire n23272;
    wire n23275;
    wire n23278;
    wire n23281;
    wire n23284;
    wire n23287;
    wire n23290;
    wire n23293;
    wire n23296;
    wire n23299;
    wire n23302;
    wire n23305;
    wire n23308;
    wire n23311;
    wire n23314;
    wire n23317;
    wire n23320;
    wire n23323;
    wire n23326;
    wire n23329;
    wire n23332;
    wire n23335;
    wire n23338;
    wire n23341;
    wire n23344;
    wire n23347;
    wire n23350;
    wire n23353;
    wire n23356;
    wire n23359;
    wire n23362;
    wire n23365;
    wire n23368;
    wire n23371;
    wire n23374;
    wire n23377;
    wire n23380;
    wire n23383;
    wire n23386;
    wire n23389;
    wire n23392;
    wire n23395;
    wire n23398;
    wire n23401;
    wire n23404;
    wire n23407;
    wire n23410;
    wire n23413;
    wire n23416;
    wire n23419;
    wire n23422;
    wire n23425;
    wire n23428;
    wire n23431;
    wire n23434;
    wire n23437;
    wire n23440;
    wire n23443;
    wire n23446;
    wire n23449;
    wire n23452;
    wire n23455;
    wire n23458;
    wire n23461;
    wire n23464;
    wire n23467;
    wire n23470;
    wire n23473;
    wire n23476;
    wire n23479;
    wire n23482;
    wire n23485;
    wire n23488;
    wire n23491;
    wire n23494;
    wire n23497;
    wire n23500;
    wire n23503;
    wire n23506;
    wire n23509;
    wire n23512;
    wire n23515;
    wire n23518;
    wire n23521;
    wire n23524;
    wire n23527;
    wire n23530;
    wire n23533;
    wire n23536;
    wire n23539;
    wire n23542;
    wire n23545;
    wire n23548;
    wire n23551;
    wire n23554;
    wire n23557;
    wire n23560;
    wire n23563;
    wire n23566;
    wire n23569;
    wire n23572;
    wire n23575;
    wire n23578;
    wire n23581;
    wire n23584;
    wire n23587;
    wire n23590;
    wire n23593;
    wire n23596;
    wire n23599;
    wire n23602;
    wire n23605;
    wire n23608;
    wire n23611;
    wire n23614;
    wire n23617;
    wire n23620;
    wire n23623;
    wire n23626;
    wire n23629;
    wire n23632;
    wire n23635;
    wire n23638;
    wire n23641;
    wire n23644;
    wire n23647;
    wire n23650;
    wire n23653;
    wire n23656;
    wire n23659;
    wire n23662;
    wire n23665;
    wire n23668;
    wire n23671;
    wire n23674;
    wire n23677;
    wire n23680;
    wire n23683;
    wire n23686;
    wire n23689;
    wire n23692;
    wire n23695;
    wire n23698;
    wire n23701;
    wire n23704;
    wire n23707;
    wire n23710;
    wire n23713;
    wire n23716;
    wire n23719;
    wire n23722;
    wire n23725;
    wire n23728;
    wire n23731;
    wire n23734;
    wire n23737;
    wire n23740;
    wire n23743;
    wire n23746;
    wire n23749;
    wire n23752;
    wire n23755;
    wire n23758;
    wire n23761;
    wire n23764;
    wire n23767;
    wire n23770;
    wire n23773;
    wire n23776;
    wire n23779;
    wire n23782;
    wire n23785;
    wire n23788;
    wire n23791;
    wire n23794;
    wire n23797;
    wire n23799;
    wire n23802;
    wire n23805;
    wire n23809;
    wire n23811;
    wire n23814;
    wire n23817;
    wire n23820;
    wire n23823;
    wire n23826;
    wire n23829;
    wire n23832;
    wire n23835;
    wire n23839;
    wire n23842;
    wire n23845;
    wire n23848;
    wire n23851;
    wire n23854;
    wire n23857;
    wire n23860;
    wire n23863;
    wire n23866;
    wire n23869;
    wire n23872;
    wire n23875;
    wire n23878;
    wire n23881;
    wire n23884;
    wire n23887;
    wire n23890;
    wire n23893;
    wire n23896;
    wire n23899;
    wire n23902;
    wire n23905;
    wire n23908;
    wire n23911;
    wire n23914;
    wire n23917;
    wire n23920;
    wire n23923;
    wire n23926;
    wire n23929;
    wire n23932;
    wire n23935;
    wire n23938;
    wire n23941;
    wire n23944;
    wire n23947;
    wire n23950;
    wire n23953;
    wire n23956;
    wire n23959;
    wire n23962;
    wire n23965;
    wire n23968;
    wire n23971;
    wire n23974;
    wire n23977;
    wire n23980;
    wire n23983;
    wire n23986;
    wire n23989;
    wire n23992;
    wire n23994;
    wire n23998;
    wire n24001;
    wire n24004;
    wire n24007;
    wire n24010;
    wire n24013;
    wire n24016;
    wire n24019;
    wire n24022;
    wire n24025;
    wire n24028;
    wire n24031;
    wire n24034;
    wire n24037;
    wire n24040;
    wire n24043;
    wire n24046;
    wire n24049;
    wire n24052;
    wire n24055;
    wire n24058;
    wire n24061;
    wire n24064;
    wire n24067;
    wire n24070;
    wire n24073;
    wire n24076;
    wire n24079;
    wire n24082;
    wire n24085;
    wire n24088;
    wire n24091;
    wire n24094;
    wire n24097;
    wire n24100;
    wire n24103;
    wire n24106;
    wire n24109;
    wire n24112;
    wire n24115;
    wire n24118;
    wire n24121;
    wire n24124;
    wire n24127;
    wire n24130;
    wire n24133;
    wire n24136;
    wire n24139;
    wire n24142;
    wire n24145;
    wire n24148;
    wire n24151;
    wire n24154;
    wire n24157;
    wire n24160;
    wire n24163;
    wire n24166;
    wire n24169;
    wire n24172;
    wire n24175;
    wire n24178;
    wire n24181;
    wire n24184;
    wire n24187;
    wire n24190;
    wire n24193;
    wire n24196;
    wire n24199;
    wire n24202;
    wire n24205;
    wire n24208;
    wire n24211;
    wire n24214;
    wire n24217;
    wire n24220;
    wire n24223;
    wire n24226;
    wire n24229;
    wire n24232;
    wire n24235;
    wire n24238;
    wire n24241;
    wire n24244;
    wire n24247;
    wire n24250;
    wire n24253;
    wire n24256;
    wire n24259;
    wire n24262;
    wire n24265;
    wire n24268;
    wire n24271;
    wire n24274;
    wire n24277;
    wire n24280;
    wire n24283;
    wire n24286;
    wire n24289;
    wire n24292;
    wire n24295;
    wire n24298;
    wire n24301;
    wire n24304;
    wire n24307;
    wire n24310;
    wire n24313;
    wire n24316;
    wire n24319;
    wire n24322;
    wire n24325;
    wire n24328;
    wire n24331;
    wire n24334;
    wire n24337;
    wire n24340;
    wire n24343;
    wire n24346;
    wire n24349;
    wire n24352;
    wire n24355;
    wire n24358;
    wire n24361;
    wire n24364;
    wire n24367;
    wire n24370;
    wire n24373;
    wire n24376;
    wire n24379;
    wire n24382;
    wire n24385;
    wire n24388;
    wire n24391;
    wire n24394;
    wire n24397;
    wire n24400;
    wire n24403;
    wire n24406;
    wire n24409;
    wire n24412;
    wire n24415;
    wire n24418;
    wire n24421;
    wire n24424;
    wire n24427;
    wire n24430;
    wire n24433;
    wire n24436;
    wire n24439;
    wire n24442;
    wire n24445;
    wire n24448;
    wire n24451;
    wire n24454;
    wire n24457;
    wire n24460;
    wire n24463;
    wire n24466;
    wire n24469;
    wire n24472;
    wire n24475;
    wire n24478;
    wire n24481;
    wire n24484;
    wire n24487;
    wire n24490;
    wire n24493;
    wire n24496;
    wire n24499;
    wire n24502;
    wire n24505;
    wire n24508;
    wire n24511;
    wire n24514;
    wire n24517;
    wire n24520;
    wire n24523;
    wire n24526;
    wire n24529;
    wire n24532;
    wire n24535;
    wire n24538;
    wire n24541;
    wire n24544;
    wire n24547;
    wire n24550;
    wire n24553;
    wire n24556;
    wire n24559;
    wire n24562;
    wire n24565;
    wire n24568;
    wire n24571;
    wire n24574;
    wire n24577;
    wire n24580;
    wire n24583;
    wire n24586;
    wire n24589;
    wire n24592;
    wire n24595;
    wire n24598;
    wire n24601;
    wire n24604;
    wire n24607;
    wire n24610;
    wire n24613;
    wire n24616;
    wire n24619;
    wire n24622;
    wire n24625;
    wire n24628;
    wire n24631;
    wire n24634;
    wire n24637;
    wire n24640;
    wire n24643;
    wire n24646;
    wire n24649;
    wire n24652;
    wire n24655;
    wire n24658;
    wire n24661;
    wire n24664;
    wire n24667;
    wire n24670;
    wire n24673;
    wire n24676;
    wire n24679;
    wire n24682;
    wire n24685;
    wire n24688;
    wire n24691;
    wire n24694;
    wire n24697;
    wire n24700;
    wire n24703;
    wire n24706;
    wire n24709;
    wire n24712;
    wire n24715;
    wire n24718;
    wire n24721;
    wire n24724;
    wire n24727;
    wire n24730;
    wire n24733;
    wire n24736;
    wire n24739;
    wire n24742;
    wire n24745;
    wire n24748;
    wire n24751;
    wire n24754;
    wire n24757;
    wire n24760;
    wire n24763;
    wire n24766;
    wire n24769;
    wire n24772;
    wire n24775;
    wire n24778;
    wire n24781;
    wire n24784;
    wire n24787;
    wire n24790;
    wire n24793;
    wire n24796;
    wire n24799;
    wire n24802;
    wire n24805;
    wire n24808;
    wire n24811;
    wire n24814;
    wire n24817;
    wire n24820;
    wire n24823;
    wire n24826;
    wire n24829;
    wire n24832;
    wire n24835;
    wire n24838;
    wire n24841;
    wire n24844;
    wire n24847;
    wire n24850;
    wire n24853;
    wire n24856;
    wire n24859;
    wire n24862;
    wire n24865;
    wire n24868;
    wire n24871;
    wire n24874;
    wire n24877;
    wire n24880;
    wire n24883;
    wire n24886;
    wire n24889;
    wire n24892;
    wire n24895;
    wire n24898;
    wire n24901;
    wire n24904;
    wire n24907;
    wire n24910;
    wire n24913;
    wire n24916;
    wire n24919;
    wire n24922;
    wire n24925;
    wire n24928;
    wire n24931;
    wire n24934;
    wire n24937;
    wire n24940;
    wire n24943;
    wire n24946;
    wire n24949;
    wire n24952;
    wire n24955;
    wire n24958;
    wire n24961;
    wire n24964;
    wire n24967;
    wire n24970;
    wire n24973;
    wire n24976;
    wire n24979;
    wire n24982;
    wire n24985;
    wire n24988;
    wire n24991;
    wire n24994;
    wire n24997;
    wire n25000;
    wire n25003;
    wire n25006;
    wire n25009;
    wire n25012;
    wire n25014;
    wire n25017;
    wire n25020;
    wire n25024;
    wire n25026;
    wire n25029;
    wire n25032;
    wire n25035;
    wire n25038;
    wire n25041;
    wire n25044;
    wire n25047;
    wire n25050;
    wire n25054;
    wire n25056;
    wire n25060;
    wire n25063;
    wire n25066;
    wire n25069;
    wire n25072;
    wire n25075;
    wire n25078;
    wire n25081;
    wire n25084;
    wire n25087;
    wire n25090;
    wire n25093;
    wire n25096;
    wire n25099;
    wire n25102;
    wire n25105;
    wire n25108;
    wire n25111;
    wire n25114;
    wire n25117;
    wire n25120;
    wire n25123;
    wire n25126;
    wire n25129;
    wire n25132;
    wire n25135;
    wire n25138;
    wire n25141;
    wire n25144;
    wire n25147;
    wire n25150;
    wire n25153;
    wire n25156;
    wire n25159;
    wire n25162;
    wire n25165;
    wire n25168;
    wire n25171;
    wire n25174;
    wire n25177;
    wire n25180;
    wire n25183;
    wire n25186;
    wire n25189;
    wire n25192;
    wire n25195;
    wire n25198;
    wire n25201;
    wire n25204;
    wire n25207;
    wire n25210;
    wire n25213;
    wire n25216;
    wire n25219;
    wire n25222;
    wire n25225;
    wire n25228;
    wire n25231;
    wire n25234;
    wire n25237;
    wire n25240;
    wire n25243;
    wire n25246;
    wire n25249;
    wire n25252;
    wire n25255;
    wire n25258;
    wire n25261;
    wire n25264;
    wire n25267;
    wire n25270;
    wire n25273;
    wire n25276;
    wire n25279;
    wire n25282;
    wire n25285;
    wire n25288;
    wire n25291;
    wire n25294;
    wire n25297;
    wire n25300;
    wire n25303;
    wire n25306;
    wire n25309;
    wire n25312;
    wire n25315;
    wire n25318;
    wire n25321;
    wire n25324;
    wire n25327;
    wire n25330;
    wire n25333;
    wire n25336;
    wire n25339;
    wire n25342;
    wire n25345;
    wire n25348;
    wire n25351;
    wire n25354;
    wire n25357;
    wire n25360;
    wire n25363;
    wire n25366;
    wire n25369;
    wire n25372;
    wire n25375;
    wire n25378;
    wire n25381;
    wire n25384;
    wire n25387;
    wire n25390;
    wire n25393;
    wire n25396;
    wire n25399;
    wire n25402;
    wire n25405;
    wire n25408;
    wire n25411;
    wire n25414;
    wire n25417;
    wire n25420;
    wire n25423;
    wire n25426;
    wire n25429;
    wire n25432;
    wire n25435;
    wire n25438;
    wire n25441;
    wire n25444;
    wire n25447;
    wire n25450;
    wire n25453;
    wire n25456;
    wire n25459;
    wire n25462;
    wire n25465;
    wire n25468;
    wire n25471;
    wire n25474;
    wire n25477;
    wire n25480;
    wire n25483;
    wire n25486;
    wire n25489;
    wire n25492;
    wire n25495;
    wire n25498;
    wire n25501;
    wire n25504;
    wire n25507;
    wire n25510;
    wire n25513;
    wire n25516;
    wire n25519;
    wire n25522;
    wire n25525;
    wire n25528;
    wire n25531;
    wire n25534;
    wire n25537;
    wire n25540;
    wire n25543;
    wire n25546;
    wire n25549;
    wire n25552;
    wire n25555;
    wire n25558;
    wire n25561;
    wire n25564;
    wire n25567;
    wire n25570;
    wire n25573;
    wire n25576;
    wire n25579;
    wire n25582;
    wire n25585;
    wire n25588;
    wire n25591;
    wire n25594;
    wire n25597;
    wire n25600;
    wire n25603;
    wire n25606;
    wire n25609;
    wire n25612;
    wire n25615;
    wire n25618;
    wire n25621;
    wire n25624;
    wire n25627;
    wire n25630;
    wire n25633;
    wire n25636;
    wire n25639;
    wire n25642;
    wire n25645;
    wire n25648;
    wire n25651;
    wire n25654;
    wire n25657;
    wire n25660;
    wire n25663;
    wire n25666;
    wire n25669;
    wire n25672;
    wire n25675;
    wire n25678;
    wire n25681;
    wire n25684;
    wire n25687;
    wire n25690;
    wire n25693;
    wire n25696;
    wire n25699;
    wire n25702;
    wire n25705;
    wire n25708;
    wire n25711;
    wire n25714;
    wire n25717;
    wire n25720;
    wire n25723;
    wire n25726;
    wire n25729;
    wire n25732;
    wire n25735;
    wire n25738;
    wire n25741;
    wire n25744;
    wire n25747;
    wire n25750;
    wire n25753;
    wire n25756;
    wire n25759;
    wire n25762;
    wire n25765;
    wire n25768;
    wire n25771;
    wire n25774;
    wire n25777;
    wire n25780;
    wire n25783;
    wire n25786;
    wire n25789;
    wire n25792;
    wire n25795;
    wire n25798;
    wire n25801;
    wire n25804;
    wire n25807;
    wire n25810;
    wire n25813;
    wire n25816;
    wire n25819;
    wire n25822;
    wire n25825;
    wire n25828;
    wire n25831;
    wire n25834;
    wire n25837;
    wire n25840;
    wire n25843;
    wire n25846;
    wire n25849;
    wire n25852;
    wire n25855;
    wire n25858;
    wire n25861;
    wire n25864;
    wire n25867;
    wire n25870;
    wire n25873;
    wire n25876;
    wire n25879;
    wire n25882;
    wire n25885;
    wire n25888;
    wire n25891;
    wire n25894;
    wire n25897;
    wire n25900;
    wire n25903;
    wire n25906;
    wire n25909;
    wire n25912;
    wire n25915;
    wire n25918;
    wire n25921;
    wire n25924;
    wire n25927;
    wire n25930;
    wire n25933;
    wire n25936;
    wire n25939;
    wire n25942;
    wire n25945;
    wire n25948;
    wire n25951;
    wire n25954;
    wire n25957;
    wire n25960;
    wire n25963;
    wire n25966;
    wire n25969;
    wire n25972;
    wire n25975;
    wire n25978;
    wire n25981;
    wire n25984;
    wire n25987;
    wire n25990;
    wire n25993;
    wire n25996;
    wire n25999;
    wire n26002;
    wire n26005;
    wire n26008;
    wire n26011;
    wire n26014;
    wire n26017;
    wire n26020;
    wire n26023;
    wire n26026;
    wire n26029;
    wire n26032;
    wire n26035;
    wire n26038;
    wire n26041;
    wire n26044;
    wire n26047;
    wire n26050;
    wire n26053;
    wire n26056;
    wire n26059;
    wire n26062;
    wire n26065;
    wire n26068;
    wire n26071;
    wire n26074;
    wire n26077;
    wire n26080;
    wire n26083;
    wire n26086;
    wire n26089;
    wire n26092;
    wire n26095;
    wire n26098;
    wire n26101;
    wire n26104;
    wire n26107;
    wire n26110;
    wire n26113;
    wire n26116;
    wire n26119;
    wire n26122;
    wire n26125;
    wire n26128;
    wire n26131;
    wire n26134;
    wire n26137;
    wire n26140;
    wire n26143;
    wire n26146;
    wire n26149;
    wire n26152;
    wire n26155;
    wire n26158;
    wire n26161;
    wire n26164;
    wire n26167;
    wire n26170;
    wire n26173;
    wire n26176;
    wire n26179;
    wire n26182;
    wire n26185;
    wire n26188;
    wire n26191;
    wire n26194;
    wire n26197;
    wire n26200;
    wire n26203;
    wire n26206;
    wire n26209;
    wire n26212;
    wire n26215;
    wire n26218;
    wire n26221;
    wire n26224;
    wire n26227;
    wire n26230;
    wire n26233;
    wire n26236;
    wire n26239;
    wire n26242;
    wire n26244;
    wire n26247;
    wire n26250;
    wire n26254;
    wire n26256;
    wire n26259;
    wire n26262;
    wire n26265;
    wire n26268;
    wire n26271;
    wire n26274;
    wire n26277;
    wire n26280;
    wire n26284;
    wire n26286;
    wire n26290;
    wire n26293;
    wire n26296;
    wire n26299;
    wire n26302;
    wire n26305;
    wire n26308;
    wire n26311;
    wire n26314;
    wire n26317;
    wire n26320;
    wire n26323;
    wire n26326;
    wire n26329;
    wire n26332;
    wire n26335;
    wire n26338;
    wire n26341;
    wire n26344;
    wire n26347;
    wire n26350;
    wire n26353;
    wire n26356;
    wire n26359;
    wire n26362;
    wire n26365;
    wire n26368;
    wire n26371;
    wire n26374;
    wire n26377;
    wire n26380;
    wire n26383;
    wire n26386;
    wire n26389;
    wire n26392;
    wire n26395;
    wire n26398;
    wire n26401;
    wire n26404;
    wire n26407;
    wire n26410;
    wire n26413;
    wire n26416;
    wire n26419;
    wire n26422;
    wire n26425;
    wire n26428;
    wire n26431;
    wire n26434;
    wire n26437;
    wire n26440;
    wire n26443;
    wire n26446;
    wire n26449;
    wire n26452;
    wire n26455;
    wire n26458;
    wire n26461;
    wire n26464;
    wire n26467;
    wire n26470;
    wire n26473;
    wire n26476;
    wire n26479;
    wire n26482;
    wire n26485;
    wire n26488;
    wire n26491;
    wire n26494;
    wire n26497;
    wire n26500;
    wire n26503;
    wire n26506;
    wire n26509;
    wire n26512;
    wire n26515;
    wire n26518;
    wire n26521;
    wire n26524;
    wire n26527;
    wire n26530;
    wire n26533;
    wire n26536;
    wire n26539;
    wire n26542;
    wire n26545;
    wire n26548;
    wire n26551;
    wire n26554;
    wire n26557;
    wire n26560;
    wire n26563;
    wire n26566;
    wire n26569;
    wire n26572;
    wire n26575;
    wire n26578;
    wire n26581;
    wire n26584;
    wire n26587;
    wire n26590;
    wire n26593;
    wire n26596;
    wire n26599;
    wire n26602;
    wire n26605;
    wire n26608;
    wire n26611;
    wire n26614;
    wire n26617;
    wire n26620;
    wire n26623;
    wire n26626;
    wire n26629;
    wire n26632;
    wire n26635;
    wire n26638;
    wire n26641;
    wire n26644;
    wire n26647;
    wire n26650;
    wire n26653;
    wire n26656;
    wire n26659;
    wire n26662;
    wire n26665;
    wire n26668;
    wire n26671;
    wire n26674;
    wire n26677;
    wire n26680;
    wire n26683;
    wire n26686;
    wire n26689;
    wire n26692;
    wire n26695;
    wire n26698;
    wire n26701;
    wire n26704;
    wire n26707;
    wire n26710;
    wire n26713;
    wire n26716;
    wire n26719;
    wire n26722;
    wire n26725;
    wire n26728;
    wire n26731;
    wire n26734;
    wire n26737;
    wire n26740;
    wire n26743;
    wire n26746;
    wire n26749;
    wire n26752;
    wire n26755;
    wire n26758;
    wire n26761;
    wire n26764;
    wire n26767;
    wire n26770;
    wire n26773;
    wire n26776;
    wire n26779;
    wire n26782;
    wire n26785;
    wire n26788;
    wire n26791;
    wire n26794;
    wire n26797;
    wire n26800;
    wire n26803;
    wire n26806;
    wire n26809;
    wire n26812;
    wire n26815;
    wire n26818;
    wire n26821;
    wire n26824;
    wire n26827;
    wire n26830;
    wire n26833;
    wire n26836;
    wire n26839;
    wire n26842;
    wire n26845;
    wire n26848;
    wire n26851;
    wire n26854;
    wire n26857;
    wire n26860;
    wire n26863;
    wire n26866;
    wire n26869;
    wire n26872;
    wire n26875;
    wire n26878;
    wire n26881;
    wire n26884;
    wire n26887;
    wire n26890;
    wire n26893;
    wire n26896;
    wire n26899;
    wire n26902;
    wire n26905;
    wire n26908;
    wire n26911;
    wire n26914;
    wire n26917;
    wire n26920;
    wire n26923;
    wire n26926;
    wire n26929;
    wire n26932;
    wire n26935;
    wire n26938;
    wire n26941;
    wire n26944;
    wire n26947;
    wire n26950;
    wire n26953;
    wire n26956;
    wire n26959;
    wire n26962;
    wire n26965;
    wire n26968;
    wire n26971;
    wire n26974;
    wire n26977;
    wire n26980;
    wire n26983;
    wire n26986;
    wire n26989;
    wire n26992;
    wire n26995;
    wire n26998;
    wire n27001;
    wire n27004;
    wire n27007;
    wire n27010;
    wire n27013;
    wire n27016;
    wire n27019;
    wire n27022;
    wire n27025;
    wire n27028;
    wire n27031;
    wire n27034;
    wire n27037;
    wire n27040;
    wire n27043;
    wire n27046;
    wire n27049;
    wire n27052;
    wire n27055;
    wire n27058;
    wire n27061;
    wire n27064;
    wire n27067;
    wire n27070;
    wire n27073;
    wire n27076;
    wire n27079;
    wire n27082;
    wire n27085;
    wire n27088;
    wire n27091;
    wire n27094;
    wire n27097;
    wire n27100;
    wire n27103;
    wire n27106;
    wire n27109;
    wire n27112;
    wire n27115;
    wire n27118;
    wire n27121;
    wire n27124;
    wire n27127;
    wire n27130;
    wire n27133;
    wire n27136;
    wire n27139;
    wire n27142;
    wire n27145;
    wire n27148;
    wire n27151;
    wire n27154;
    wire n27157;
    wire n27160;
    wire n27163;
    wire n27166;
    wire n27169;
    wire n27172;
    wire n27175;
    wire n27178;
    wire n27181;
    wire n27184;
    wire n27187;
    wire n27190;
    wire n27193;
    wire n27196;
    wire n27199;
    wire n27202;
    wire n27205;
    wire n27208;
    wire n27211;
    wire n27214;
    wire n27217;
    wire n27220;
    wire n27223;
    wire n27226;
    wire n27229;
    wire n27232;
    wire n27235;
    wire n27238;
    wire n27241;
    wire n27244;
    wire n27247;
    wire n27250;
    wire n27253;
    wire n27256;
    wire n27259;
    wire n27262;
    wire n27265;
    wire n27268;
    wire n27271;
    wire n27274;
    wire n27277;
    wire n27280;
    wire n27283;
    wire n27286;
    wire n27289;
    wire n27292;
    wire n27295;
    wire n27298;
    wire n27301;
    wire n27304;
    wire n27307;
    wire n27310;
    wire n27313;
    wire n27316;
    wire n27319;
    wire n27322;
    wire n27325;
    wire n27328;
    wire n27331;
    wire n27334;
    wire n27337;
    wire n27340;
    wire n27343;
    wire n27346;
    wire n27349;
    wire n27352;
    wire n27355;
    wire n27358;
    wire n27361;
    wire n27364;
    wire n27367;
    wire n27370;
    wire n27373;
    wire n27376;
    wire n27379;
    wire n27382;
    wire n27385;
    wire n27388;
    wire n27391;
    wire n27394;
    wire n27397;
    wire n27400;
    wire n27403;
    wire n27406;
    wire n27409;
    wire n27412;
    wire n27415;
    wire n27418;
    wire n27421;
    wire n27424;
    wire n27427;
    wire n27430;
    wire n27433;
    wire n27436;
    wire n27439;
    wire n27442;
    wire n27445;
    wire n27448;
    wire n27451;
    wire n27454;
    wire n27457;
    wire n27460;
    wire n27463;
    wire n27466;
    wire n27469;
    wire n27472;
    wire n27475;
    wire n27478;
    wire n27481;
    wire n27484;
    wire n27487;
    wire n27490;
    wire n27493;
    wire n27496;
    wire n27499;
    wire n27502;
    wire n27505;
    wire n27507;
    wire n27510;
    wire n27513;
    wire n27517;
    wire n27519;
    wire n27522;
    wire n27525;
    wire n27528;
    wire n27531;
    wire n27534;
    wire n27537;
    wire n27540;
    wire n27543;
    wire n27547;
    wire n27549;
    wire n27553;
    wire n27556;
    wire n27559;
    wire n27562;
    wire n27565;
    wire n27568;
    wire n27571;
    wire n27574;
    wire n27577;
    wire n27580;
    wire n27583;
    wire n27586;
    wire n27589;
    wire n27592;
    wire n27595;
    wire n27598;
    wire n27601;
    wire n27604;
    wire n27607;
    wire n27610;
    wire n27613;
    wire n27616;
    wire n27619;
    wire n27622;
    wire n27625;
    wire n27628;
    wire n27631;
    wire n27634;
    wire n27637;
    wire n27640;
    wire n27643;
    wire n27646;
    wire n27649;
    wire n27652;
    wire n27655;
    wire n27658;
    wire n27661;
    wire n27664;
    wire n27667;
    wire n27670;
    wire n27673;
    wire n27676;
    wire n27679;
    wire n27682;
    wire n27685;
    wire n27688;
    wire n27691;
    wire n27694;
    wire n27697;
    wire n27700;
    wire n27703;
    wire n27706;
    wire n27709;
    wire n27712;
    wire n27715;
    wire n27718;
    wire n27721;
    wire n27724;
    wire n27727;
    wire n27730;
    wire n27733;
    wire n27736;
    wire n27739;
    wire n27742;
    wire n27745;
    wire n27748;
    wire n27751;
    wire n27754;
    wire n27757;
    wire n27760;
    wire n27763;
    wire n27766;
    wire n27769;
    wire n27772;
    wire n27775;
    wire n27778;
    wire n27781;
    wire n27784;
    wire n27787;
    wire n27790;
    wire n27793;
    wire n27796;
    wire n27799;
    wire n27802;
    wire n27805;
    wire n27808;
    wire n27811;
    wire n27814;
    wire n27817;
    wire n27820;
    wire n27823;
    wire n27826;
    wire n27829;
    wire n27832;
    wire n27835;
    wire n27838;
    wire n27841;
    wire n27844;
    wire n27847;
    wire n27850;
    wire n27853;
    wire n27856;
    wire n27859;
    wire n27862;
    wire n27865;
    wire n27868;
    wire n27871;
    wire n27874;
    wire n27877;
    wire n27880;
    wire n27883;
    wire n27886;
    wire n27889;
    wire n27892;
    wire n27895;
    wire n27898;
    wire n27901;
    wire n27904;
    wire n27907;
    wire n27910;
    wire n27913;
    wire n27916;
    wire n27919;
    wire n27922;
    wire n27925;
    wire n27928;
    wire n27931;
    wire n27934;
    wire n27937;
    wire n27940;
    wire n27943;
    wire n27946;
    wire n27949;
    wire n27952;
    wire n27955;
    wire n27958;
    wire n27961;
    wire n27964;
    wire n27967;
    wire n27970;
    wire n27973;
    wire n27976;
    wire n27979;
    wire n27982;
    wire n27985;
    wire n27988;
    wire n27991;
    wire n27994;
    wire n27997;
    wire n28000;
    wire n28003;
    wire n28006;
    wire n28009;
    wire n28012;
    wire n28015;
    wire n28018;
    wire n28021;
    wire n28024;
    wire n28027;
    wire n28030;
    wire n28033;
    wire n28036;
    wire n28039;
    wire n28042;
    wire n28045;
    wire n28048;
    wire n28051;
    wire n28054;
    wire n28057;
    wire n28060;
    wire n28063;
    wire n28066;
    wire n28069;
    wire n28072;
    wire n28075;
    wire n28078;
    wire n28081;
    wire n28084;
    wire n28087;
    wire n28090;
    wire n28093;
    wire n28096;
    wire n28099;
    wire n28102;
    wire n28105;
    wire n28108;
    wire n28111;
    wire n28114;
    wire n28117;
    wire n28120;
    wire n28123;
    wire n28126;
    wire n28129;
    wire n28132;
    wire n28135;
    wire n28138;
    wire n28141;
    wire n28144;
    wire n28147;
    wire n28150;
    wire n28153;
    wire n28156;
    wire n28159;
    wire n28162;
    wire n28165;
    wire n28168;
    wire n28171;
    wire n28174;
    wire n28177;
    wire n28180;
    wire n28183;
    wire n28186;
    wire n28189;
    wire n28192;
    wire n28195;
    wire n28198;
    wire n28201;
    wire n28204;
    wire n28207;
    wire n28210;
    wire n28213;
    wire n28216;
    wire n28219;
    wire n28222;
    wire n28225;
    wire n28228;
    wire n28231;
    wire n28234;
    wire n28237;
    wire n28240;
    wire n28243;
    wire n28246;
    wire n28249;
    wire n28252;
    wire n28255;
    wire n28258;
    wire n28261;
    wire n28264;
    wire n28267;
    wire n28270;
    wire n28273;
    wire n28276;
    wire n28279;
    wire n28282;
    wire n28285;
    wire n28288;
    wire n28291;
    wire n28294;
    wire n28297;
    wire n28300;
    wire n28303;
    wire n28306;
    wire n28309;
    wire n28312;
    wire n28315;
    wire n28318;
    wire n28321;
    wire n28324;
    wire n28327;
    wire n28330;
    wire n28333;
    wire n28336;
    wire n28339;
    wire n28342;
    wire n28345;
    wire n28348;
    wire n28351;
    wire n28354;
    wire n28357;
    wire n28360;
    wire n28363;
    wire n28366;
    wire n28369;
    wire n28372;
    wire n28375;
    wire n28378;
    wire n28381;
    wire n28384;
    wire n28387;
    wire n28390;
    wire n28393;
    wire n28396;
    wire n28399;
    wire n28402;
    wire n28405;
    wire n28408;
    wire n28411;
    wire n28414;
    wire n28417;
    wire n28420;
    wire n28423;
    wire n28426;
    wire n28429;
    wire n28432;
    wire n28435;
    wire n28438;
    wire n28441;
    wire n28444;
    wire n28447;
    wire n28450;
    wire n28453;
    wire n28456;
    wire n28459;
    wire n28462;
    wire n28465;
    wire n28468;
    wire n28471;
    wire n28474;
    wire n28477;
    wire n28480;
    wire n28483;
    wire n28486;
    wire n28489;
    wire n28492;
    wire n28495;
    wire n28498;
    wire n28501;
    wire n28504;
    wire n28507;
    wire n28510;
    wire n28513;
    wire n28516;
    wire n28519;
    wire n28522;
    wire n28525;
    wire n28528;
    wire n28531;
    wire n28534;
    wire n28537;
    wire n28540;
    wire n28543;
    wire n28546;
    wire n28549;
    wire n28552;
    wire n28555;
    wire n28558;
    wire n28561;
    wire n28564;
    wire n28567;
    wire n28570;
    wire n28573;
    wire n28576;
    wire n28579;
    wire n28582;
    wire n28585;
    wire n28588;
    wire n28591;
    wire n28594;
    wire n28597;
    wire n28600;
    wire n28603;
    wire n28606;
    wire n28609;
    wire n28612;
    wire n28615;
    wire n28618;
    wire n28621;
    wire n28624;
    wire n28627;
    wire n28630;
    wire n28633;
    wire n28636;
    wire n28639;
    wire n28642;
    wire n28645;
    wire n28648;
    wire n28651;
    wire n28654;
    wire n28657;
    wire n28660;
    wire n28663;
    wire n28666;
    wire n28669;
    wire n28672;
    wire n28675;
    wire n28678;
    wire n28681;
    wire n28684;
    wire n28687;
    wire n28690;
    wire n28693;
    wire n28696;
    wire n28699;
    wire n28702;
    wire n28705;
    wire n28708;
    wire n28711;
    wire n28714;
    wire n28717;
    wire n28720;
    wire n28723;
    wire n28726;
    wire n28729;
    wire n28732;
    wire n28735;
    wire n28738;
    wire n28741;
    wire n28744;
    wire n28747;
    wire n28750;
    wire n28753;
    wire n28756;
    wire n28759;
    wire n28762;
    wire n28765;
    wire n28768;
    wire n28771;
    wire n28774;
    wire n28777;
    wire n28780;
    wire n28783;
    wire n28786;
    wire n28789;
    wire n28792;
    wire n28795;
    wire n28798;
    wire n28801;
    wire n28804;
    wire n28807;
    wire n28810;
    wire n28813;
    wire n28816;
    wire n28819;
    wire n28822;
    wire n28824;
    wire n28827;
    wire n28830;
    wire n28834;
    wire n28836;
    wire n28839;
    wire n28842;
    wire n28845;
    wire n28848;
    wire n28851;
    wire n28854;
    wire n28857;
    wire n28860;
    wire n28864;
    wire n28867;
    wire n28870;
    wire n28873;
    wire n28876;
    wire n28879;
    wire n28882;
    wire n28885;
    wire n28888;
    wire n28891;
    wire n28894;
    wire n28897;
    wire n28900;
    wire n28903;
    wire n28906;
    wire n28909;
    wire n28912;
    wire n28915;
    wire n28918;
    wire n28921;
    wire n28924;
    wire n28927;
    wire n28930;
    wire n28933;
    wire n28936;
    wire n28939;
    wire n28942;
    wire n28945;
    wire n28948;
    wire n28951;
    wire n28954;
    wire n28957;
    wire n28960;
    wire n28963;
    wire n28966;
    wire n28969;
    wire n28972;
    wire n28975;
    wire n28978;
    wire n28981;
    wire n28984;
    wire n28987;
    wire n28990;
    wire n28993;
    wire n28996;
    wire n28999;
    wire n29002;
    wire n29005;
    wire n29008;
    wire n29011;
    wire n29014;
    wire n29017;
    wire n29020;
    wire n29023;
    wire n29026;
    wire n29029;
    wire n29032;
    wire n29035;
    wire n29038;
    wire n29041;
    wire n29044;
    wire n29047;
    wire n29050;
    wire n29053;
    wire n29056;
    wire n29059;
    wire n29062;
    wire n29065;
    wire n29068;
    wire n29071;
    wire n29074;
    wire n29077;
    wire n29080;
    wire n29083;
    wire n29086;
    wire n29089;
    wire n29092;
    wire n29095;
    wire n29098;
    wire n29101;
    wire n29104;
    wire n29107;
    wire n29110;
    wire n29113;
    wire n29116;
    wire n29119;
    wire n29122;
    wire n29125;
    wire n29128;
    wire n29131;
    wire n29134;
    wire n29137;
    wire n29140;
    wire n29143;
    wire n29146;
    wire n29149;
    wire n29152;
    wire n29155;
    wire n29158;
    wire n29161;
    wire n29164;
    wire n29167;
    wire n29170;
    wire n29173;
    wire n29176;
    wire n29179;
    wire n29182;
    wire n29185;
    wire n29188;
    wire n29191;
    wire n29194;
    wire n29197;
    wire n29200;
    wire n29203;
    wire n29206;
    wire n29209;
    wire n29212;
    wire n29214;
    wire n29218;
    wire n29221;
    wire n29224;
    wire n29227;
    wire n29230;
    wire n29233;
    wire n29236;
    wire n29239;
    wire n29242;
    wire n29245;
    wire n29248;
    wire n29251;
    wire n29254;
    wire n29257;
    wire n29260;
    wire n29263;
    wire n29266;
    wire n29269;
    wire n29272;
    wire n29275;
    wire n29278;
    wire n29281;
    wire n29284;
    wire n29287;
    wire n29290;
    wire n29293;
    wire n29296;
    wire n29299;
    wire n29302;
    wire n29305;
    wire n29308;
    wire n29311;
    wire n29314;
    wire n29317;
    wire n29320;
    wire n29323;
    wire n29326;
    wire n29329;
    wire n29332;
    wire n29335;
    wire n29338;
    wire n29341;
    wire n29344;
    wire n29347;
    wire n29350;
    wire n29353;
    wire n29356;
    wire n29359;
    wire n29362;
    wire n29365;
    wire n29368;
    wire n29371;
    wire n29374;
    wire n29377;
    wire n29380;
    wire n29383;
    wire n29386;
    wire n29389;
    wire n29392;
    wire n29395;
    wire n29398;
    wire n29401;
    wire n29404;
    wire n29407;
    wire n29410;
    wire n29413;
    wire n29416;
    wire n29419;
    wire n29422;
    wire n29425;
    wire n29428;
    wire n29431;
    wire n29434;
    wire n29437;
    wire n29440;
    wire n29443;
    wire n29446;
    wire n29449;
    wire n29452;
    wire n29455;
    wire n29458;
    wire n29461;
    wire n29464;
    wire n29467;
    wire n29470;
    wire n29473;
    wire n29476;
    wire n29479;
    wire n29482;
    wire n29485;
    wire n29488;
    wire n29491;
    wire n29494;
    wire n29497;
    wire n29500;
    wire n29503;
    wire n29506;
    wire n29509;
    wire n29512;
    wire n29515;
    wire n29518;
    wire n29521;
    wire n29524;
    wire n29527;
    wire n29530;
    wire n29533;
    wire n29536;
    wire n29539;
    wire n29542;
    wire n29545;
    wire n29548;
    wire n29551;
    wire n29554;
    wire n29557;
    wire n29560;
    wire n29563;
    wire n29566;
    wire n29569;
    wire n29572;
    wire n29575;
    wire n29578;
    wire n29581;
    wire n29584;
    wire n29587;
    wire n29590;
    wire n29593;
    wire n29596;
    wire n29599;
    wire n29602;
    wire n29605;
    wire n29608;
    wire n29611;
    wire n29614;
    wire n29617;
    wire n29620;
    wire n29623;
    wire n29626;
    wire n29629;
    wire n29632;
    wire n29635;
    wire n29638;
    wire n29641;
    wire n29644;
    wire n29647;
    wire n29650;
    wire n29653;
    wire n29656;
    wire n29659;
    wire n29662;
    wire n29665;
    wire n29668;
    wire n29671;
    wire n29674;
    wire n29677;
    wire n29680;
    wire n29683;
    wire n29686;
    wire n29689;
    wire n29692;
    wire n29695;
    wire n29698;
    wire n29701;
    wire n29704;
    wire n29707;
    wire n29710;
    wire n29713;
    wire n29716;
    wire n29719;
    wire n29722;
    wire n29725;
    wire n29728;
    wire n29731;
    wire n29734;
    wire n29737;
    wire n29740;
    wire n29743;
    wire n29746;
    wire n29749;
    wire n29752;
    wire n29755;
    wire n29758;
    wire n29761;
    wire n29764;
    wire n29767;
    wire n29770;
    wire n29773;
    wire n29776;
    wire n29779;
    wire n29782;
    wire n29785;
    wire n29788;
    wire n29791;
    wire n29794;
    wire n29797;
    wire n29800;
    wire n29803;
    wire n29806;
    wire n29809;
    wire n29812;
    wire n29815;
    wire n29818;
    wire n29821;
    wire n29824;
    wire n29827;
    wire n29830;
    wire n29833;
    wire n29836;
    wire n29839;
    wire n29842;
    wire n29845;
    wire n29848;
    wire n29851;
    wire n29854;
    wire n29857;
    wire n29860;
    wire n29863;
    wire n29866;
    wire n29869;
    wire n29872;
    wire n29875;
    wire n29878;
    wire n29881;
    wire n29884;
    wire n29887;
    wire n29890;
    wire n29893;
    wire n29896;
    wire n29899;
    wire n29902;
    wire n29905;
    wire n29908;
    wire n29911;
    wire n29914;
    wire n29917;
    wire n29920;
    wire n29923;
    wire n29926;
    wire n29929;
    wire n29932;
    wire n29935;
    wire n29938;
    wire n29941;
    wire n29944;
    wire n29947;
    wire n29950;
    wire n29953;
    wire n29956;
    wire n29959;
    wire n29962;
    wire n29965;
    wire n29968;
    wire n29971;
    wire n29974;
    wire n29977;
    wire n29980;
    wire n29983;
    wire n29986;
    wire n29989;
    wire n29992;
    wire n29995;
    wire n29998;
    wire n30001;
    wire n30004;
    wire n30007;
    wire n30010;
    wire n30013;
    wire n30016;
    wire n30019;
    wire n30022;
    wire n30025;
    wire n30028;
    wire n30031;
    wire n30034;
    wire n30037;
    wire n30040;
    wire n30043;
    wire n30046;
    wire n30049;
    wire n30052;
    wire n30055;
    wire n30058;
    wire n30061;
    wire n30064;
    wire n30067;
    wire n30070;
    wire n30073;
    wire n30076;
    wire n30079;
    wire n30082;
    wire n30085;
    wire n30088;
    wire n30091;
    wire n30094;
    wire n30097;
    wire n30100;
    wire n30103;
    wire n30106;
    wire n30109;
    wire n30112;
    wire n30115;
    wire n30118;
    wire n30121;
    wire n30124;
    wire n30127;
    wire n30130;
    wire n30133;
    wire n30136;
    wire n30139;
    wire n30142;
    wire n30145;
    wire n30148;
    wire n30151;
    wire n30154;
    wire n30157;
    wire n30160;
    wire n30163;
    wire n30166;
    wire n30169;
    wire n30172;
    wire n30175;
    wire n30178;
    wire n30181;
    wire n30184;
    wire n30187;
    wire n30190;
    wire n30193;
    wire n30196;
    wire n30199;
    wire n30202;
    wire n30205;
    wire n30208;
    wire n30211;
    wire n30214;
    wire n30217;
    wire n30220;
    wire n30223;
    wire n30226;
    wire n30229;
    wire n30232;
    wire n30235;
    wire n30238;
    wire n30241;
    wire n30244;
    wire n30247;
    wire n30250;
    wire n30253;
    wire n30256;
    wire n30259;
    wire n30262;
    wire n30265;
    wire n30268;
    wire n30271;
    wire n30274;
    wire n30277;
    wire n30280;
    wire n30283;
    wire n30286;
    wire n30289;
    wire n30292;
    wire n30295;
    wire n30298;
    wire n30301;
    wire n30304;
    wire n30307;
    wire n30310;
    wire n30313;
    wire n30316;
    wire n30319;
    wire n30322;
    wire n30325;
    wire n30328;
    wire n30331;
    wire n30334;
    wire n30337;
    wire n30340;
    wire n30343;
    wire n30346;
    wire n30349;
    wire n30352;
    wire n30355;
    wire n30358;
    wire n30361;
    wire n30364;
    wire n30367;
    wire n30370;
    wire n30373;
    wire n30376;
    wire n30379;
    wire n30382;
    wire n30385;
    wire n30388;
    wire n30391;
    wire n30394;
    wire n30397;
    wire n30400;
    wire n30403;
    wire n30406;
    wire n30409;
    wire n30412;
    wire n30415;
    wire n30418;
    wire n30421;
    wire n30424;
    wire n30427;
    wire n30430;
    wire n30433;
    wire n30436;
    wire n30439;
    wire n30442;
    wire n30445;
    wire n30448;
    wire n30451;
    wire n30454;
    wire n30457;
    wire n30460;
    wire n30463;
    wire n30466;
    wire n30469;
    wire n30472;
    wire n30475;
    wire n30478;
    wire n30481;
    wire n30484;
    wire n30487;
    wire n30490;
    wire n30493;
    wire n30496;
    wire n30499;
    wire n30502;
    wire n30505;
    wire n30508;
    wire n30511;
    wire n30514;
    wire n30517;
    wire n30520;
    wire n30523;
    wire n30526;
    wire n30529;
    wire n30532;
    wire n30535;
    wire n30538;
    wire n30541;
    wire n30544;
    wire n30547;
    wire n30550;
    wire n30553;
    wire n30556;
    wire n30559;
    wire n30562;
    wire n30565;
    wire n30568;
    wire n30571;
    wire n30574;
    wire n30577;
    wire n30580;
    wire n30583;
    wire n30586;
    wire n30589;
    wire n30592;
    wire n30595;
    wire n30598;
    wire n30601;
    wire n30604;
    wire n30607;
    wire n30610;
    wire n30613;
    wire n30616;
    wire n30619;
    wire n30622;
    wire n30625;
    wire n30628;
    wire n30631;
    wire n30634;
    wire n30637;
    wire n30640;
    wire n30643;
    wire n30646;
    wire n30649;
    wire n30652;
    wire n30655;
    wire n30658;
    wire n30661;
    wire n30664;
    wire n30667;
    wire n30670;
    wire n30673;
    wire n30676;
    wire n30679;
    wire n30682;
    wire n30685;
    wire n30688;
    wire n30691;
    wire n30694;
    wire n30697;
    wire n30700;
    wire n30703;
    wire n30706;
    wire n30709;
    wire n30712;
    wire n30715;
    wire n30718;
    wire n30721;
    wire n30724;
    wire n30727;
    wire n30730;
    wire n30733;
    wire n30736;
    wire n30739;
    wire n30742;
    wire n30745;
    wire n30748;
    wire n30751;
    wire n30754;
    wire n30757;
    wire n30760;
    wire n30763;
    wire n30766;
    wire n30769;
    wire n30772;
    wire n30775;
    wire n30778;
    wire n30781;
    wire n30784;
    wire n30787;
    wire n30790;
    wire n30793;
    wire n30796;
    wire n30799;
    wire n30802;
    wire n30805;
    wire n30808;
    wire n30811;
    wire n30814;
    wire n30817;
    wire n30820;
    wire n30823;
    wire n30826;
    wire n30829;
    wire n30832;
    wire n30835;
    wire n30838;
    wire n30841;
    wire n30844;
    wire n30847;
    wire n30850;
    wire n30853;
    wire n30856;
    wire n30859;
    wire n30862;
    wire n30865;
    wire n30868;
    wire n30871;
    wire n30874;
    wire n30877;
    wire n30880;
    wire n30883;
    wire n30886;
    wire n30889;
    wire n30892;
    wire n30895;
    wire n30898;
    wire n30901;
    wire n30904;
    wire n30907;
    wire n30910;
    wire n30913;
    wire n30916;
    wire n30919;
    wire n30922;
    wire n30925;
    wire n30928;
    wire n30931;
    wire n30934;
    wire n30937;
    wire n30940;
    wire n30943;
    wire n30946;
    wire n30949;
    wire n30952;
    wire n30955;
    wire n30958;
    wire n30961;
    wire n30964;
    wire n30967;
    wire n30970;
    wire n30973;
    wire n30976;
    wire n30979;
    wire n30982;
    wire n30985;
    wire n30988;
    wire n30991;
    wire n30994;
    wire n30997;
    wire n31000;
    wire n31003;
    wire n31006;
    wire n31009;
    wire n31012;
    wire n31015;
    wire n31018;
    wire n31021;
    wire n31024;
    wire n31027;
    wire n31030;
    wire n31033;
    wire n31036;
    wire n31039;
    wire n31042;
    wire n31045;
    wire n31048;
    wire n31051;
    wire n31054;
    wire n31057;
    wire n31060;
    wire n31063;
    wire n31066;
    wire n31069;
    wire n31072;
    wire n31075;
    wire n31078;
    wire n31081;
    wire n31084;
    wire n31087;
    wire n31090;
    wire n31093;
    wire n31096;
    wire n31099;
    wire n31102;
    wire n31105;
    wire n31108;
    wire n31111;
    wire n31114;
    wire n31117;
    wire n31120;
    wire n31123;
    wire n31126;
    wire n31129;
    wire n31132;
    wire n31135;
    wire n31138;
    wire n31141;
    wire n31144;
    wire n31147;
    wire n31150;
    wire n31153;
    wire n31156;
    wire n31159;
    wire n31162;
    wire n31165;
    wire n31168;
    wire n31171;
    wire n31174;
    wire n31177;
    wire n31180;
    wire n31183;
    wire n31186;
    wire n31189;
    wire n31192;
    wire n31195;
    wire n31198;
    wire n31201;
    wire n31204;
    wire n31207;
    wire n31210;
    wire n31213;
    wire n31216;
    wire n31219;
    wire n31222;
    wire n31225;
    wire n31228;
    wire n31231;
    wire n31234;
    wire n31237;
    wire n31240;
    wire n31243;
    wire n31246;
    wire n31249;
    wire n31252;
    wire n31255;
    wire n31258;
    wire n31261;
    wire n31264;
    wire n31267;
    wire n31270;
    wire n31273;
    wire n31276;
    wire n31279;
    wire n31282;
    wire n31285;
    wire n31288;
    wire n31291;
    wire n31294;
    wire n31297;
    wire n31300;
    wire n31303;
    wire n31306;
    wire n31309;
    wire n31312;
    wire n31315;
    wire n31318;
    wire n31321;
    wire n31324;
    wire n31327;
    wire n31330;
    wire n31333;
    wire n31336;
    wire n31339;
    wire n31342;
    wire n31345;
    wire n31348;
    wire n31351;
    wire n31354;
    wire n31357;
    wire n31360;
    wire n31363;
    wire n31366;
    wire n31369;
    wire n31372;
    wire n31375;
    wire n31378;
    wire n31381;
    wire n31384;
    wire n31387;
    wire n31390;
    wire n31393;
    wire n31396;
    wire n31399;
    wire n31402;
    wire n31405;
    wire n31408;
    wire n31411;
    wire n31414;
    wire n31417;
    wire n31420;
    wire n31423;
    wire n31426;
    wire n31429;
    wire n31432;
    wire n31435;
    wire n31438;
    wire n31441;
    wire n31444;
    wire n31447;
    wire n31450;
    wire n31453;
    wire n31456;
    wire n31459;
    wire n31462;
    wire n31465;
    wire n31468;
    wire n31471;
    wire n31474;
    wire n31477;
    wire n31480;
    wire n31483;
    wire n31486;
    wire n31489;
    wire n31492;
    wire n31495;
    wire n31498;
    wire n31501;
    wire n31504;
    wire n31507;
    wire n31510;
    wire n31513;
    wire n31516;
    wire n31519;
    wire n31522;
    wire n31525;
    wire n31528;
    wire n31531;
    wire n31534;
    wire n31537;
    wire n31540;
    wire n31543;
    wire n31546;
    wire n31549;
    wire n31552;
    wire n31555;
    wire n31558;
    wire n31561;
    wire n31564;
    wire n31567;
    wire n31570;
    wire n31573;
    wire n31576;
    wire n31579;
    wire n31582;
    wire n31585;
    wire n31588;
    wire n31591;
    wire n31594;
    wire n31597;
    wire n31600;
    wire n31603;
    wire n31606;
    wire n31609;
    wire n31612;
    wire n31615;
    wire n31618;
    wire n31621;
    wire n31624;
    wire n31627;
    wire n31630;
    wire n31633;
    wire n31636;
    wire n31639;
    wire n31642;
    wire n31645;
    wire n31648;
    wire n31651;
    wire n31654;
    wire n31657;
    wire n31660;
    wire n31663;
    wire n31666;
    wire n31669;
    wire n31672;
    wire n31675;
    wire n31678;
    wire n31681;
    wire n31684;
    wire n31687;
    wire n31690;
    wire n31693;
    wire n31696;
    wire n31699;
    wire n31702;
    wire n31705;
    wire n31708;
    wire n31711;
    wire n31714;
    wire n31717;
    wire n31720;
    wire n31723;
    wire n31726;
    wire n31729;
    wire n31732;
    wire n31735;
    wire n31738;
    wire n31741;
    wire n31744;
    wire n31747;
    wire n31750;
    wire n31753;
    wire n31756;
    wire n31759;
    wire n31762;
    wire n31765;
    wire n31768;
    wire n31771;
    wire n31774;
    wire n31777;
    wire n31780;
    wire n31783;
    wire n31786;
    wire n31789;
    wire n31792;
    wire n31795;
    wire n31798;
    wire n31801;
    wire n31804;
    wire n31807;
    wire n31810;
    wire n31813;
    wire n31816;
    wire n31819;
    wire n31822;
    wire n31825;
    wire n31828;
    wire n31831;
    wire n31834;
    wire n31837;
    wire n31840;
    wire n31843;
    wire n31846;
    wire n31849;
    wire n31852;
    wire n31855;
    wire n31858;
    wire n31861;
    wire n31864;
    wire n31867;
    wire n31870;
    wire n31873;
    wire n31876;
    wire n31879;
    wire n31882;
    wire n31885;
    wire n31888;
    wire n31891;
    wire n31894;
    wire n31897;
    wire n31900;
    wire n31903;
    wire n31906;
    wire n31909;
    wire n31912;
    wire n31915;
    wire n31918;
    wire n31921;
    wire n31924;
    wire n31927;
    wire n31930;
    wire n31933;
    wire n31936;
    wire n31939;
    wire n31942;
    wire n31945;
    wire n31948;
    wire n31951;
    wire n31954;
    wire n31957;
    wire n31960;
    wire n31963;
    wire n31966;
    wire n31969;
    wire n31972;
    wire n31975;
    wire n31978;
    wire n31981;
    wire n31984;
    wire n31987;
    wire n31990;
    wire n31993;
    wire n31996;
    wire n31999;
    wire n32002;
    wire n32005;
    wire n32008;
    wire n32011;
    wire n32014;
    wire n32017;
    wire n32020;
    wire n32023;
    wire n32026;
    wire n32029;
    wire n32032;
    wire n32035;
    wire n32038;
    wire n32041;
    wire n32044;
    wire n32047;
    wire n32050;
    wire n32053;
    wire n32056;
    wire n32059;
    wire n32062;
    wire n32065;
    wire n32068;
    wire n32071;
    wire n32074;
    wire n32077;
    wire n32080;
    wire n32083;
    wire n32086;
    wire n32089;
    wire n32092;
    wire n32095;
    wire n32098;
    wire n32101;
    wire n32104;
    wire n32107;
    wire n32110;
    wire n32113;
    wire n32116;
    wire n32119;
    wire n32122;
    wire n32125;
    wire n32128;
    wire n32131;
    wire n32134;
    wire n32137;
    wire n32140;
    wire n32143;
    wire n32146;
    wire n32149;
    wire n32152;
    wire n32155;
    wire n32158;
    wire n32161;
    wire n32164;
    wire n32167;
    wire n32170;
    wire n32173;
    wire n32176;
    wire n32179;
    wire n32182;
    wire n32185;
    wire n32188;
    wire n32191;
    wire n32194;
    wire n32197;
    wire n32200;
    wire n32203;
    wire n32206;
    wire n32209;
    wire n32212;
    wire n32215;
    wire n32218;
    wire n32221;
    wire n32224;
    wire n32227;
    wire n32230;
    wire n32233;
    wire n32236;
    wire n32239;
    wire n32242;
    wire n32245;
    wire n32248;
    wire n32251;
    wire n32254;
    wire n32257;
    wire n32260;
    wire n32263;
    wire n32266;
    wire n32269;
    wire n32272;
    wire n32275;
    wire n32278;
    wire n32281;
    wire n32284;
    wire n32287;
    wire n32290;
    wire n32293;
    wire n32296;
    wire n32299;
    wire n32302;
    wire n32305;
    wire n32308;
    wire n32311;
    wire n32314;
    wire n32317;
    wire n32320;
    wire n32323;
    wire n32326;
    wire n32329;
    wire n32332;
    wire n32335;
    wire n32338;
    wire n32341;
    wire n32344;
    wire n32347;
    wire n32350;
    wire n32353;
    wire n32356;
    wire n32359;
    wire n32362;
    wire n32365;
    wire n32368;
    wire n32371;
    wire n32374;
    wire n32377;
    wire n32380;
    wire n32383;
    wire n32386;
    wire n32389;
    wire n32392;
    wire n32395;
    wire n32398;
    wire n32401;
    wire n32404;
    wire n32407;
    wire n32410;
    wire n32413;
    wire n32416;
    wire n32419;
    wire n32422;
    wire n32425;
    wire n32428;
    wire n32431;
    wire n32434;
    wire n32437;
    wire n32440;
    wire n32443;
    wire n32446;
    wire n32449;
    wire n32452;
    wire n32455;
    wire n32458;
    wire n32461;
    wire n32464;
    wire n32467;
    wire n32470;
    wire n32473;
    wire n32476;
    wire n32479;
    wire n32482;
    wire n32485;
    wire n32488;
    wire n32491;
    wire n32494;
    wire n32497;
    wire n32500;
    wire n32503;
    wire n32506;
    wire n32509;
    wire n32512;
    wire n32515;
    wire n32518;
    wire n32521;
    wire n32524;
    wire n32527;
    wire n32530;
    wire n32533;
    wire n32536;
    wire n32539;
    wire n32542;
    wire n32545;
    wire n32548;
    wire n32551;
    wire n32554;
    wire n32557;
    wire n32560;
    wire n32563;
    wire n32566;
    wire n32569;
    wire n32572;
    wire n32575;
    wire n32578;
    wire n32581;
    wire n32584;
    wire n32587;
    wire n32590;
    wire n32593;
    wire n32596;
    wire n32599;
    wire n32602;
    wire n32605;
    wire n32608;
    wire n32611;
    wire n32614;
    wire n32617;
    wire n32620;
    wire n32623;
    wire n32626;
    wire n32629;
    wire n32632;
    wire n32635;
    wire n32638;
    wire n32641;
    wire n32644;
    wire n32647;
    wire n32650;
    wire n32653;
    wire n32656;
    wire n32659;
    wire n32662;
    wire n32665;
    wire n32668;
    wire n32671;
    wire n32674;
    wire n32677;
    wire n32680;
    wire n32683;
    wire n32686;
    wire n32689;
    wire n32692;
    wire n32695;
    wire n32698;
    wire n32701;
    wire n32704;
    wire n32707;
    wire n32710;
    wire n32712;
    wire n32715;
    wire n32718;
    wire n32722;
    wire n32725;
    wire n32728;
    wire n32731;
    wire n32734;
    wire n32737;
    wire n32740;
    wire n32743;
    wire n32746;
    wire n32748;
    wire n32751;
    wire n32754;
    wire n32757;
    wire n32760;
    wire n32763;
    wire n32766;
    wire n32770;
    wire n32773;
    wire n32776;
    wire n32779;
    wire n32782;
    wire n32785;
    wire n32788;
    wire n32791;
    wire n32794;
    wire n32797;
    wire n32800;
    wire n32803;
    wire n32806;
    wire n32809;
    wire n32812;
    wire n32815;
    wire n32818;
    wire n32821;
    wire n32824;
    wire n32827;
    wire n32830;
    wire n32833;
    wire n32836;
    wire n32839;
    wire n32841;
    wire n32844;
    wire n32847;
    wire n32850;
    wire n32853;
    wire n32856;
    wire n32860;
    wire n32863;
    wire n32866;
    wire n32869;
    wire n32872;
    wire n32874;
    wire n32877;
    wire n32880;
    wire n32883;
    wire n32886;
    wire n32889;
    wire n32893;
    wire n32895;
    wire n32898;
    wire n32901;
    wire n32904;
    wire n32907;
    wire n32910;
    wire n32913;
    wire n32916;
    wire n32919;
    wire n32922;
    wire n32925;
    wire n32928;
    wire n32931;
    wire n32934;
    wire n32937;
    wire n32940;
    wire n32943;
    wire n32946;
    wire n32949;
    wire n32952;
    wire n32955;
    wire n32958;
    wire n32961;
    wire n32964;
    wire n32967;
    wire n32970;
    wire n32973;
    wire n32976;
    wire n32979;
    wire n32982;
    wire n32985;
    wire n32988;
    wire n32991;
    wire n32994;
    wire n32997;
    wire n33000;
    wire n33003;
    wire n33006;
    wire n33009;
    wire n33012;
    wire n33015;
    wire n33018;
    wire n33021;
    wire n33024;
    wire n33027;
    wire n33030;
    wire n33033;
    wire n33036;
    wire n33039;
    wire n33042;
    wire n33045;
    wire n33048;
    wire n33051;
    wire n33054;
    wire n33057;
    wire n33060;
    wire n33063;
    wire n33066;
    wire n33069;
    wire n33072;
    wire n33075;
    wire n33078;
    wire n33081;
    wire n33084;
    wire n33087;
    wire n33090;
    wire n33093;
    wire n33096;
    wire n33099;
    wire n33102;
    wire n33105;
    wire n33108;
    wire n33111;
    wire n33114;
    wire n33117;
    wire n33120;
    wire n33123;
    wire n33126;
    wire n33129;
    wire n33135;
    wire n33138;
    wire n33141;
    wire n33144;
    wire n33147;
    wire n33150;
    wire n33153;
    wire n33156;
    wire n33159;
    wire n33162;
    wire n33165;
    wire n33168;
    wire n33171;
    wire n33174;
    wire n33177;
    wire n33180;
    wire n33183;
    wire n33186;
    wire n33189;
    wire n33192;
    wire n33195;
    wire n33198;
    wire n33201;
    wire n33204;
    wire n33207;
    wire n33210;
    wire n33213;
    wire n33216;
    wire n33219;
    wire n33222;
    wire n33225;
    wire n33228;
    wire n33231;
    wire n33234;
    wire n33237;
    wire n33240;
    wire n33243;
    wire n33246;
    wire n33249;
    wire n33252;
    wire n33255;
    wire n33258;
    wire n33261;
    wire n33264;
    wire n33267;
    wire n33270;
    wire n33273;
    wire n33276;
    wire n33279;
    wire n33282;
    wire n33285;
    wire n33288;
    wire n33291;
    wire n33294;
    wire n33297;
    wire n33300;
    wire n33303;
    wire n33306;
    wire n33309;
    wire n33312;
    wire n33315;
    wire n33318;
    wire n33321;
    wire n33324;
    wire n33327;
    wire n33330;
    wire n33333;
    wire n33336;
    wire n33339;
    wire n33342;
    wire n33345;
    wire n33351;
    wire n33354;
    wire n33357;
    wire n33360;
    wire n33363;
    wire n33366;
    wire n33369;
    wire n33372;
    wire n33375;
    wire n33378;
    wire n33381;
    wire n33384;
    wire n33387;
    wire n33390;
    wire n33393;
    wire n33396;
    wire n33399;
    wire n33402;
    wire n33405;
    wire n33408;
    wire n33411;
    wire n33414;
    wire n33417;
    wire n33420;
    wire n33423;
    wire n33426;
    wire n33429;
    wire n33432;
    wire n33435;
    wire n33438;
    wire n33441;
    wire n33444;
    wire n33447;
    wire n33450;
    wire n33453;
    wire n33456;
    wire n33459;
    wire n33462;
    wire n33465;
    wire n33468;
    wire n33471;
    wire n33474;
    wire n33477;
    wire n33480;
    wire n33483;
    wire n33486;
    wire n33489;
    wire n33492;
    wire n33495;
    wire n33498;
    wire n33501;
    wire n33504;
    wire n33507;
    wire n33510;
    wire n33513;
    wire n33516;
    wire n33519;
    wire n33522;
    wire n33525;
    wire n33528;
    wire n33531;
    wire n33534;
    wire n33537;
    wire n33540;
    wire n33543;
    wire n33546;
    wire n33549;
    wire n33552;
    wire n33558;
    wire n33561;
    wire n33564;
    wire n33567;
    wire n33570;
    wire n33573;
    wire n33576;
    wire n33579;
    wire n33582;
    wire n33585;
    wire n33588;
    wire n33591;
    wire n33594;
    wire n33597;
    wire n33600;
    wire n33603;
    wire n33606;
    wire n33609;
    wire n33612;
    wire n33615;
    wire n33618;
    wire n33621;
    wire n33624;
    wire n33627;
    wire n33630;
    wire n33633;
    wire n33636;
    wire n33639;
    wire n33642;
    wire n33645;
    wire n33648;
    wire n33651;
    wire n33654;
    wire n33657;
    wire n33660;
    wire n33663;
    wire n33666;
    wire n33669;
    wire n33672;
    wire n33675;
    wire n33678;
    wire n33681;
    wire n33684;
    wire n33687;
    wire n33690;
    wire n33693;
    wire n33696;
    wire n33699;
    wire n33702;
    wire n33705;
    wire n33708;
    wire n33711;
    wire n33714;
    wire n33717;
    wire n33720;
    wire n33723;
    wire n33726;
    wire n33729;
    wire n33732;
    wire n33735;
    wire n33738;
    wire n33741;
    wire n33744;
    wire n33747;
    wire n33750;
    wire n33756;
    wire n33759;
    wire n33762;
    wire n33765;
    wire n33768;
    wire n33771;
    wire n33774;
    wire n33777;
    wire n33780;
    wire n33783;
    wire n33786;
    wire n33789;
    wire n33792;
    wire n33795;
    wire n33798;
    wire n33801;
    wire n33804;
    wire n33807;
    wire n33810;
    wire n33813;
    wire n33816;
    wire n33819;
    wire n33822;
    wire n33825;
    wire n33828;
    wire n33831;
    wire n33834;
    wire n33837;
    wire n33840;
    wire n33843;
    wire n33846;
    wire n33849;
    wire n33852;
    wire n33855;
    wire n33858;
    wire n33861;
    wire n33864;
    wire n33867;
    wire n33870;
    wire n33873;
    wire n33876;
    wire n33879;
    wire n33882;
    wire n33885;
    wire n33888;
    wire n33891;
    wire n33894;
    wire n33897;
    wire n33900;
    wire n33903;
    wire n33906;
    wire n33909;
    wire n33912;
    wire n33915;
    wire n33918;
    wire n33921;
    wire n33924;
    wire n33927;
    wire n33930;
    wire n33933;
    wire n33936;
    wire n33939;
    wire n33945;
    wire n33948;
    wire n33951;
    wire n33954;
    wire n33957;
    wire n33960;
    wire n33963;
    wire n33966;
    wire n33969;
    wire n33972;
    wire n33975;
    wire n33978;
    wire n33981;
    wire n33984;
    wire n33987;
    wire n33990;
    wire n33993;
    wire n33996;
    wire n33999;
    wire n34002;
    wire n34005;
    wire n34008;
    wire n34011;
    wire n34014;
    wire n34017;
    wire n34020;
    wire n34023;
    wire n34026;
    wire n34029;
    wire n34032;
    wire n34035;
    wire n34038;
    wire n34041;
    wire n34044;
    wire n34047;
    wire n34050;
    wire n34053;
    wire n34056;
    wire n34059;
    wire n34062;
    wire n34065;
    wire n34068;
    wire n34071;
    wire n34074;
    wire n34077;
    wire n34080;
    wire n34083;
    wire n34086;
    wire n34089;
    wire n34092;
    wire n34095;
    wire n34098;
    wire n34101;
    wire n34104;
    wire n34107;
    wire n34110;
    wire n34113;
    wire n34116;
    wire n34119;
    wire n34125;
    wire n34128;
    wire n34131;
    wire n34134;
    wire n34137;
    wire n34140;
    wire n34143;
    wire n34146;
    wire n34149;
    wire n34152;
    wire n34155;
    wire n34158;
    wire n34161;
    wire n34164;
    wire n34167;
    wire n34170;
    wire n34173;
    wire n34176;
    wire n34179;
    wire n34182;
    wire n34185;
    wire n34188;
    wire n34191;
    wire n34194;
    wire n34197;
    wire n34200;
    wire n34203;
    wire n34206;
    wire n34209;
    wire n34212;
    wire n34215;
    wire n34218;
    wire n34221;
    wire n34224;
    wire n34227;
    wire n34230;
    wire n34233;
    wire n34236;
    wire n34239;
    wire n34242;
    wire n34245;
    wire n34248;
    wire n34251;
    wire n34254;
    wire n34257;
    wire n34260;
    wire n34263;
    wire n34266;
    wire n34269;
    wire n34272;
    wire n34275;
    wire n34278;
    wire n34281;
    wire n34284;
    wire n34287;
    wire n34290;
    wire n34296;
    wire n34299;
    wire n34302;
    wire n34305;
    wire n34308;
    wire n34311;
    wire n34314;
    wire n34317;
    wire n34320;
    wire n34323;
    wire n34326;
    wire n34329;
    wire n34332;
    wire n34335;
    wire n34338;
    wire n34341;
    wire n34344;
    wire n34347;
    wire n34350;
    wire n34353;
    wire n34356;
    wire n34359;
    wire n34362;
    wire n34365;
    wire n34368;
    wire n34371;
    wire n34374;
    wire n34377;
    wire n34380;
    wire n34383;
    wire n34386;
    wire n34389;
    wire n34392;
    wire n34395;
    wire n34398;
    wire n34401;
    wire n34404;
    wire n34407;
    wire n34410;
    wire n34413;
    wire n34416;
    wire n34419;
    wire n34422;
    wire n34425;
    wire n34428;
    wire n34431;
    wire n34434;
    wire n34437;
    wire n34440;
    wire n34443;
    wire n34446;
    wire n34449;
    wire n34452;
    wire n34458;
    wire n34461;
    wire n34464;
    wire n34467;
    wire n34470;
    wire n34473;
    wire n34476;
    wire n34479;
    wire n34482;
    wire n34485;
    wire n34488;
    wire n34491;
    wire n34494;
    wire n34497;
    wire n34500;
    wire n34503;
    wire n34506;
    wire n34509;
    wire n34512;
    wire n34515;
    wire n34518;
    wire n34521;
    wire n34524;
    wire n34527;
    wire n34530;
    wire n34533;
    wire n34536;
    wire n34539;
    wire n34542;
    wire n34545;
    wire n34548;
    wire n34551;
    wire n34554;
    wire n34557;
    wire n34560;
    wire n34563;
    wire n34566;
    wire n34569;
    wire n34572;
    wire n34575;
    wire n34578;
    wire n34581;
    wire n34584;
    wire n34587;
    wire n34590;
    wire n34593;
    wire n34596;
    wire n34599;
    wire n34602;
    wire n34605;
    wire n34611;
    wire n34614;
    wire n34617;
    wire n34620;
    wire n34623;
    wire n34626;
    wire n34629;
    wire n34632;
    wire n34635;
    wire n34638;
    wire n34641;
    wire n34644;
    wire n34647;
    wire n34650;
    wire n34653;
    wire n34656;
    wire n34659;
    wire n34662;
    wire n34665;
    wire n34668;
    wire n34671;
    wire n34674;
    wire n34677;
    wire n34680;
    wire n34683;
    wire n34686;
    wire n34689;
    wire n34692;
    wire n34695;
    wire n34698;
    wire n34701;
    wire n34704;
    wire n34707;
    wire n34710;
    wire n34713;
    wire n34716;
    wire n34719;
    wire n34722;
    wire n34725;
    wire n34728;
    wire n34731;
    wire n34734;
    wire n34737;
    wire n34740;
    wire n34743;
    wire n34746;
    wire n34749;
    wire n34755;
    wire n34758;
    wire n34761;
    wire n34764;
    wire n34767;
    wire n34770;
    wire n34773;
    wire n34776;
    wire n34779;
    wire n34782;
    wire n34785;
    wire n34788;
    wire n34791;
    wire n34794;
    wire n34797;
    wire n34800;
    wire n34803;
    wire n34806;
    wire n34809;
    wire n34812;
    wire n34815;
    wire n34818;
    wire n34821;
    wire n34824;
    wire n34827;
    wire n34830;
    wire n34833;
    wire n34836;
    wire n34839;
    wire n34842;
    wire n34845;
    wire n34848;
    wire n34851;
    wire n34854;
    wire n34857;
    wire n34860;
    wire n34863;
    wire n34866;
    wire n34869;
    wire n34872;
    wire n34875;
    wire n34878;
    wire n34881;
    wire n34884;
    wire n34890;
    wire n34893;
    wire n34896;
    wire n34899;
    wire n34902;
    wire n34905;
    wire n34908;
    wire n34911;
    wire n34914;
    wire n34917;
    wire n34920;
    wire n34923;
    wire n34926;
    wire n34929;
    wire n34932;
    wire n34935;
    wire n34938;
    wire n34941;
    wire n34944;
    wire n34947;
    wire n34950;
    wire n34953;
    wire n34956;
    wire n34959;
    wire n34962;
    wire n34965;
    wire n34968;
    wire n34971;
    wire n34974;
    wire n34977;
    wire n34980;
    wire n34983;
    wire n34986;
    wire n34989;
    wire n34992;
    wire n34995;
    wire n34998;
    wire n35001;
    wire n35004;
    wire n35007;
    wire n35010;
    wire n35016;
    wire n35019;
    wire n35022;
    wire n35025;
    wire n35028;
    wire n35031;
    wire n35034;
    wire n35037;
    wire n35040;
    wire n35043;
    wire n35046;
    wire n35049;
    wire n35052;
    wire n35055;
    wire n35058;
    wire n35061;
    wire n35064;
    wire n35067;
    wire n35070;
    wire n35073;
    wire n35076;
    wire n35079;
    wire n35082;
    wire n35085;
    wire n35088;
    wire n35091;
    wire n35094;
    wire n35097;
    wire n35100;
    wire n35103;
    wire n35106;
    wire n35109;
    wire n35112;
    wire n35115;
    wire n35118;
    wire n35121;
    wire n35124;
    wire n35127;
    wire n35133;
    wire n35136;
    wire n35139;
    wire n35142;
    wire n35145;
    wire n35148;
    wire n35151;
    wire n35154;
    wire n35157;
    wire n35160;
    wire n35163;
    wire n35166;
    wire n35169;
    wire n35172;
    wire n35175;
    wire n35178;
    wire n35181;
    wire n35184;
    wire n35187;
    wire n35190;
    wire n35193;
    wire n35196;
    wire n35199;
    wire n35202;
    wire n35205;
    wire n35208;
    wire n35211;
    wire n35214;
    wire n35217;
    wire n35220;
    wire n35223;
    wire n35226;
    wire n35229;
    wire n35232;
    wire n35235;
    wire n35241;
    wire n35244;
    wire n35247;
    wire n35250;
    wire n35253;
    wire n35256;
    wire n35259;
    wire n35262;
    wire n35265;
    wire n35268;
    wire n35271;
    wire n35274;
    wire n35277;
    wire n35280;
    wire n35283;
    wire n35286;
    wire n35289;
    wire n35292;
    wire n35295;
    wire n35298;
    wire n35301;
    wire n35304;
    wire n35307;
    wire n35310;
    wire n35313;
    wire n35316;
    wire n35319;
    wire n35322;
    wire n35325;
    wire n35328;
    wire n35331;
    wire n35334;
    wire n35340;
    wire n35343;
    wire n35346;
    wire n35349;
    wire n35352;
    wire n35355;
    wire n35358;
    wire n35361;
    wire n35364;
    wire n35367;
    wire n35370;
    wire n35373;
    wire n35376;
    wire n35379;
    wire n35382;
    wire n35385;
    wire n35388;
    wire n35391;
    wire n35394;
    wire n35397;
    wire n35400;
    wire n35403;
    wire n35406;
    wire n35409;
    wire n35412;
    wire n35415;
    wire n35418;
    wire n35421;
    wire n35424;
    wire n35430;
    wire n35433;
    wire n35436;
    wire n35439;
    wire n35442;
    wire n35445;
    wire n35448;
    wire n35451;
    wire n35454;
    wire n35457;
    wire n35460;
    wire n35463;
    wire n35466;
    wire n35469;
    wire n35472;
    wire n35475;
    wire n35478;
    wire n35481;
    wire n35484;
    wire n35487;
    wire n35490;
    wire n35493;
    wire n35496;
    wire n35499;
    wire n35502;
    wire n35505;
    wire n35508;
    wire n35514;
    wire n35517;
    wire n35520;
    wire n35523;
    wire n35526;
    wire n35529;
    wire n35532;
    wire n35535;
    wire n35538;
    wire n35541;
    wire n35544;
    wire n35547;
    wire n35550;
    wire n35553;
    wire n35556;
    wire n35559;
    wire n35562;
    wire n35565;
    wire n35568;
    wire n35571;
    wire n35574;
    wire n35577;
    wire n35580;
    wire n35583;
    wire n35586;
    wire n35592;
    wire n35595;
    wire n35598;
    wire n35601;
    wire n35604;
    wire n35607;
    wire n35610;
    wire n35613;
    wire n35616;
    wire n35619;
    wire n35622;
    wire n35625;
    wire n35628;
    wire n35631;
    wire n35634;
    wire n35637;
    wire n35640;
    wire n35643;
    wire n35646;
    wire n35649;
    wire n35652;
    wire n35655;
    wire n35658;
    wire n35661;
    wire n35667;
    wire n35670;
    wire n35673;
    wire n35676;
    wire n35679;
    wire n35682;
    wire n35685;
    wire n35688;
    wire n35691;
    wire n35694;
    wire n35697;
    wire n35700;
    wire n35703;
    wire n35706;
    wire n35709;
    wire n35712;
    wire n35715;
    wire n35718;
    wire n35721;
    wire n35724;
    wire n35727;
    wire n35730;
    wire n35736;
    wire n35739;
    wire n35742;
    wire n35745;
    wire n35748;
    wire n35751;
    wire n35754;
    wire n35757;
    wire n35760;
    wire n35763;
    wire n35766;
    wire n35769;
    wire n35772;
    wire n35775;
    wire n35778;
    wire n35781;
    wire n35784;
    wire n35787;
    wire n35790;
    wire n35793;
    wire n35799;
    wire n35802;
    wire n35805;
    wire n35808;
    wire n35811;
    wire n35814;
    wire n35817;
    wire n35820;
    wire n35823;
    wire n35826;
    wire n35829;
    wire n35832;
    wire n35835;
    wire n35838;
    wire n35841;
    wire n35844;
    wire n35847;
    wire n35850;
    wire n35856;
    wire n35859;
    wire n35862;
    wire n35865;
    wire n35868;
    wire n35871;
    wire n35874;
    wire n35877;
    wire n35880;
    wire n35883;
    wire n35886;
    wire n35889;
    wire n35892;
    wire n35895;
    wire n35898;
    wire n35901;
    wire n35907;
    wire n35910;
    wire n35913;
    wire n35916;
    wire n35919;
    wire n35922;
    wire n35925;
    wire n35928;
    wire n35931;
    wire n35934;
    wire n35937;
    wire n35940;
    wire n35943;
    wire n35946;
    wire n35952;
    wire n35955;
    wire n35958;
    wire n35961;
    wire n35964;
    wire n35967;
    wire n35970;
    wire n35973;
    wire n35976;
    wire n35979;
    wire n35982;
    wire n35985;
    wire n35991;
    wire n35994;
    wire n35997;
    wire n36000;
    wire n36003;
    wire n36006;
    wire n36009;
    wire n36012;
    wire n36015;
    wire n36018;
    wire n36024;
    wire n36027;
    wire n36030;
    wire n36033;
    wire n36036;
    wire n36039;
    wire n36042;
    wire n36045;
    wire n36051;
    wire n36054;
    wire n36057;
    wire n36060;
    wire n36063;
    wire n36066;
    wire n36072;
    wire n36075;
    wire n36078;
    wire n36081;
    wire n36087;
    wire n36090;
    jand g0000(.dinb(G1gat), .dina(G273gat), .dout(n67));
    jxor g0001(.dinb(G18gat), .dina(G273gat), .dout(n71));
    jand g0002(.dinb(G1gat), .dina(G290gat), .dout(n75));
    jor g0003(.dinb(n71), .dina(n75), .dout(n79));
    jand g0004(.dinb(G18gat), .dina(G290gat), .dout(n83));
    jand g0005(.dinb(n67), .dina(n83), .dout(n87));
    jnot g0006(.din(n87), .dout(n90));
    jand g0007(.dinb(n10756), .dina(n90), .dout(n94));
    jand g0008(.dinb(G1gat), .dina(G307gat), .dout(n98));
    jnot g0009(.din(n98), .dout(n101));
    jdff g0010(.din(G18gat), .dout(n104));
    jnot g0011(.din(G290gat), .dout(n107));
    jor g0012(.dinb(n104), .dina(n107), .dout(n111));
    jnot g0013(.din(G35gat), .dout(n114));
    jnot g0014(.din(G273gat), .dout(n117));
    jor g0015(.dinb(n114), .dina(n117), .dout(n121));
    jand g0016(.dinb(n111), .dina(n121), .dout(n125));
    jand g0017(.dinb(G35gat), .dina(G290gat), .dout(n129));
    jand g0018(.dinb(n71), .dina(n129), .dout(n133));
    jor g0019(.dinb(n125), .dina(n15939), .dout(n137));
    jand g0020(.dinb(n14721), .dina(n137), .dout(n141));
    jnot g0021(.din(n133), .dout(n144));
    jand g0022(.dinb(n14724), .dina(n144), .dout(n148));
    jor g0023(.dinb(n141), .dina(n14704), .dout(n152));
    jxor g0024(.dinb(n10768), .dina(n152), .dout(n156));
    jand g0025(.dinb(G1gat), .dina(G324gat), .dout(n160));
    jnot g0026(.din(n160), .dout(n163));
    jnot g0027(.din(n141), .dout(n166));
    jor g0028(.dinb(n14706), .dina(n152), .dout(n170));
    jand g0029(.dinb(n14701), .dina(n170), .dout(n174));
    jand g0030(.dinb(G18gat), .dina(G307gat), .dout(n178));
    jnot g0031(.din(n178), .dout(n181));
    jand g0032(.dinb(G52gat), .dina(G273gat), .dout(n185));
    jor g0033(.dinb(n129), .dina(n185), .dout(n189));
    jand g0034(.dinb(G35gat), .dina(G273gat), .dout(n193));
    jand g0035(.dinb(G52gat), .dina(G290gat), .dout(n197));
    jand g0036(.dinb(n193), .dina(n197), .dout(n201));
    jnot g0037(.din(n201), .dout(n204));
    jand g0038(.dinb(n15964), .dina(n204), .dout(n208));
    jor g0039(.dinb(n15969), .dina(n208), .dout(n212));
    jand g0040(.dinb(n15966), .dina(n204), .dout(n216));
    jnot g0041(.din(n216), .dout(n219));
    jand g0042(.dinb(n212), .dina(n219), .dout(n223));
    jxor g0043(.dinb(n14698), .dina(n223), .dout(n227));
    jxor g0044(.dinb(n174), .dina(n14685), .dout(n231));
    jxor g0045(.dinb(n10789), .dina(n231), .dout(n235));
    jand g0046(.dinb(G1gat), .dina(G341gat), .dout(n239));
    jnot g0047(.din(n239), .dout(n242));
    jnot g0048(.din(n227), .dout(n245));
    jor g0049(.dinb(n174), .dina(n245), .dout(n249));
    jor g0050(.dinb(n14661), .dina(n231), .dout(n253));
    jand g0051(.dinb(n14659), .dina(n253), .dout(n257));
    jand g0052(.dinb(G18gat), .dina(G324gat), .dout(n261));
    jnot g0053(.din(n261), .dout(n264));
    jor g0054(.dinb(n114), .dina(n107), .dout(n268));
    jnot g0055(.din(G52gat), .dout(n271));
    jor g0056(.dinb(n271), .dina(n117), .dout(n275));
    jand g0057(.dinb(n268), .dina(n275), .dout(n279));
    jor g0058(.dinb(n279), .dina(n17064), .dout(n283));
    jand g0059(.dinb(n15936), .dina(n283), .dout(n287));
    jor g0060(.dinb(n287), .dina(n15933), .dout(n291));
    jor g0061(.dinb(n15942), .dina(n291), .dout(n295));
    jand g0062(.dinb(n15957), .dina(n295), .dout(n299));
    jand g0063(.dinb(G35gat), .dina(G307gat), .dout(n303));
    jnot g0064(.din(n303), .dout(n306));
    jand g0065(.dinb(G69gat), .dina(G273gat), .dout(n310));
    jor g0066(.dinb(n197), .dina(n310), .dout(n314));
    jand g0067(.dinb(G69gat), .dina(G290gat), .dout(n318));
    jand g0068(.dinb(n185), .dina(n318), .dout(n322));
    jnot g0069(.din(n322), .dout(n325));
    jand g0070(.dinb(n17058), .dina(n325), .dout(n329));
    jor g0071(.dinb(n17070), .dina(n329), .dout(n333));
    jand g0072(.dinb(n17067), .dina(n325), .dout(n337));
    jnot g0073(.din(n337), .dout(n340));
    jand g0074(.dinb(n333), .dina(n340), .dout(n344));
    jxor g0075(.dinb(n17056), .dina(n344), .dout(n348));
    jnot g0076(.din(n348), .dout(n351));
    jxor g0077(.dinb(n299), .dina(n351), .dout(n355));
    jxor g0078(.dinb(n14656), .dina(n355), .dout(n359));
    jxor g0079(.dinb(n257), .dina(n14634), .dout(n363));
    jxor g0080(.dinb(n10819), .dina(n363), .dout(n367));
    jand g0081(.dinb(G1gat), .dina(G358gat), .dout(n371));
    jnot g0082(.din(n371), .dout(n374));
    jnot g0083(.din(n359), .dout(n377));
    jor g0084(.dinb(n257), .dina(n377), .dout(n381));
    jor g0085(.dinb(n14601), .dina(n363), .dout(n385));
    jand g0086(.dinb(n14599), .dina(n385), .dout(n389));
    jand g0087(.dinb(G18gat), .dina(G341gat), .dout(n393));
    jnot g0088(.din(n393), .dout(n396));
    jor g0089(.dinb(n299), .dina(n351), .dout(n400));
    jxor g0090(.dinb(n299), .dina(n15930), .dout(n404));
    jor g0091(.dinb(n15906), .dina(n404), .dout(n408));
    jand g0092(.dinb(n15904), .dina(n408), .dout(n412));
    jand g0093(.dinb(G35gat), .dina(G324gat), .dout(n416));
    jnot g0094(.din(n416), .dout(n419));
    jnot g0095(.din(n314), .dout(n422));
    jor g0096(.dinb(n422), .dina(n18183), .dout(n426));
    jand g0097(.dinb(n17061), .dina(n426), .dout(n430));
    jand g0098(.dinb(n17056), .dina(n344), .dout(n434));
    jor g0099(.dinb(n17044), .dina(n434), .dout(n438));
    jand g0100(.dinb(G52gat), .dina(G307gat), .dout(n442));
    jnot g0101(.din(n442), .dout(n445));
    jand g0102(.dinb(G86gat), .dina(G273gat), .dout(n449));
    jor g0103(.dinb(n318), .dina(n449), .dout(n453));
    jand g0104(.dinb(G86gat), .dina(G290gat), .dout(n457));
    jand g0105(.dinb(n310), .dina(n457), .dout(n461));
    jnot g0106(.din(n461), .dout(n464));
    jand g0107(.dinb(n18175), .dina(n464), .dout(n468));
    jor g0108(.dinb(n18177), .dina(n468), .dout(n472));
    jor g0109(.dinb(n325), .dina(n19278), .dout(n476));
    jand g0110(.dinb(n472), .dina(n18160), .dout(n480));
    jxor g0111(.dinb(n18172), .dina(n480), .dout(n484));
    jxor g0112(.dinb(n438), .dina(n17038), .dout(n488));
    jxor g0113(.dinb(n17035), .dina(n488), .dout(n492));
    jnot g0114(.din(n492), .dout(n495));
    jxor g0115(.dinb(n412), .dina(n495), .dout(n499));
    jxor g0116(.dinb(n14596), .dina(n499), .dout(n503));
    jxor g0117(.dinb(n389), .dina(n14565), .dout(n507));
    jxor g0118(.dinb(n10858), .dina(n507), .dout(n511));
    jand g0119(.dinb(G1gat), .dina(G375gat), .dout(n515));
    jnot g0120(.din(n515), .dout(n518));
    jnot g0121(.din(n503), .dout(n521));
    jor g0122(.dinb(n389), .dina(n521), .dout(n525));
    jor g0123(.dinb(n14523), .dina(n507), .dout(n529));
    jand g0124(.dinb(n14521), .dina(n529), .dout(n533));
    jand g0125(.dinb(G18gat), .dina(G358gat), .dout(n537));
    jnot g0126(.din(n537), .dout(n540));
    jor g0127(.dinb(n412), .dina(n495), .dout(n544));
    jxor g0128(.dinb(n412), .dina(n15900), .dout(n548));
    jor g0129(.dinb(n15867), .dina(n548), .dout(n552));
    jand g0130(.dinb(n15865), .dina(n552), .dout(n556));
    jand g0131(.dinb(G35gat), .dina(G341gat), .dout(n560));
    jnot g0132(.din(n560), .dout(n563));
    jand g0133(.dinb(n438), .dina(n17038), .dout(n567));
    jand g0134(.dinb(n17035), .dina(n488), .dout(n571));
    jor g0135(.dinb(n17014), .dina(n571), .dout(n575));
    jand g0136(.dinb(G52gat), .dina(G324gat), .dout(n579));
    jnot g0137(.din(n579), .dout(n582));
    jnot g0138(.din(n472), .dout(n585));
    jand g0139(.dinb(n18172), .dina(n480), .dout(n589));
    jor g0140(.dinb(n18157), .dina(n589), .dout(n593));
    jand g0141(.dinb(G69gat), .dina(G307gat), .dout(n597));
    jnot g0142(.din(n597), .dout(n600));
    jand g0143(.dinb(G103gat), .dina(G273gat), .dout(n604));
    jor g0144(.dinb(n457), .dina(n604), .dout(n608));
    jand g0145(.dinb(G103gat), .dina(G290gat), .dout(n612));
    jand g0146(.dinb(n449), .dina(n612), .dout(n616));
    jnot g0147(.din(n616), .dout(n619));
    jand g0148(.dinb(n19267), .dina(n619), .dout(n623));
    jor g0149(.dinb(n19272), .dina(n623), .dout(n627));
    jor g0150(.dinb(n464), .dina(n19269), .dout(n631));
    jand g0151(.dinb(n627), .dina(n19252), .dout(n635));
    jxor g0152(.dinb(n19264), .dina(n635), .dout(n639));
    jxor g0153(.dinb(n593), .dina(n18154), .dout(n643));
    jxor g0154(.dinb(n18151), .dina(n643), .dout(n647));
    jxor g0155(.dinb(n575), .dina(n17011), .dout(n651));
    jxor g0156(.dinb(n17008), .dina(n651), .dout(n655));
    jnot g0157(.din(n655), .dout(n658));
    jxor g0158(.dinb(n556), .dina(n658), .dout(n662));
    jxor g0159(.dinb(n14518), .dina(n662), .dout(n666));
    jxor g0160(.dinb(n533), .dina(n14478), .dout(n670));
    jxor g0161(.dinb(n10906), .dina(n670), .dout(n674));
    jand g0162(.dinb(G1gat), .dina(G392gat), .dout(n678));
    jnot g0163(.din(n678), .dout(n681));
    jnot g0164(.din(n666), .dout(n684));
    jor g0165(.dinb(n533), .dina(n684), .dout(n688));
    jor g0166(.dinb(n14427), .dina(n670), .dout(n692));
    jand g0167(.dinb(n14425), .dina(n692), .dout(n696));
    jand g0168(.dinb(G18gat), .dina(G375gat), .dout(n700));
    jnot g0169(.din(n700), .dout(n703));
    jor g0170(.dinb(n556), .dina(n658), .dout(n707));
    jxor g0171(.dinb(n556), .dina(n15861), .dout(n711));
    jor g0172(.dinb(n15819), .dina(n711), .dout(n715));
    jand g0173(.dinb(n15817), .dina(n715), .dout(n719));
    jand g0174(.dinb(G35gat), .dina(G358gat), .dout(n723));
    jnot g0175(.din(n723), .dout(n726));
    jand g0176(.dinb(n575), .dina(n17011), .dout(n730));
    jand g0177(.dinb(n17008), .dina(n651), .dout(n734));
    jor g0178(.dinb(n16978), .dina(n734), .dout(n738));
    jand g0179(.dinb(G52gat), .dina(G341gat), .dout(n742));
    jnot g0180(.din(n742), .dout(n745));
    jand g0181(.dinb(n593), .dina(n18154), .dout(n749));
    jand g0182(.dinb(n18151), .dina(n643), .dout(n753));
    jor g0183(.dinb(n18130), .dina(n753), .dout(n757));
    jand g0184(.dinb(G69gat), .dina(G324gat), .dout(n761));
    jnot g0185(.din(n761), .dout(n764));
    jnot g0186(.din(n627), .dout(n767));
    jand g0187(.dinb(n19264), .dina(n635), .dout(n771));
    jor g0188(.dinb(n19249), .dina(n771), .dout(n775));
    jand g0189(.dinb(G86gat), .dina(G307gat), .dout(n779));
    jnot g0190(.din(n779), .dout(n782));
    jand g0191(.dinb(G120gat), .dina(G273gat), .dout(n786));
    jor g0192(.dinb(n612), .dina(n786), .dout(n790));
    jand g0193(.dinb(G120gat), .dina(G290gat), .dout(n794));
    jand g0194(.dinb(n604), .dina(n794), .dout(n798));
    jnot g0195(.din(n798), .dout(n801));
    jand g0196(.dinb(n20326), .dina(n801), .dout(n805));
    jor g0197(.dinb(n20331), .dina(n805), .dout(n809));
    jand g0198(.dinb(n20328), .dina(n801), .dout(n813));
    jnot g0199(.din(n813), .dout(n816));
    jand g0200(.dinb(n809), .dina(n816), .dout(n820));
    jxor g0201(.dinb(n20323), .dina(n820), .dout(n824));
    jxor g0202(.dinb(n775), .dina(n19246), .dout(n828));
    jxor g0203(.dinb(n19243), .dina(n828), .dout(n832));
    jxor g0204(.dinb(n757), .dina(n18127), .dout(n836));
    jxor g0205(.dinb(n18124), .dina(n836), .dout(n840));
    jxor g0206(.dinb(n738), .dina(n16975), .dout(n844));
    jxor g0207(.dinb(n16972), .dina(n844), .dout(n848));
    jnot g0208(.din(n848), .dout(n851));
    jxor g0209(.dinb(n719), .dina(n851), .dout(n855));
    jxor g0210(.dinb(n14422), .dina(n855), .dout(n859));
    jxor g0211(.dinb(n696), .dina(n14373), .dout(n863));
    jxor g0212(.dinb(n10963), .dina(n863), .dout(n867));
    jand g0213(.dinb(G1gat), .dina(G409gat), .dout(n871));
    jnot g0214(.din(n871), .dout(n874));
    jnot g0215(.din(n859), .dout(n877));
    jor g0216(.dinb(n696), .dina(n877), .dout(n881));
    jor g0217(.dinb(n14313), .dina(n863), .dout(n885));
    jand g0218(.dinb(n14311), .dina(n885), .dout(n889));
    jand g0219(.dinb(G18gat), .dina(G392gat), .dout(n893));
    jnot g0220(.din(n893), .dout(n896));
    jor g0221(.dinb(n719), .dina(n851), .dout(n900));
    jxor g0222(.dinb(n719), .dina(n15813), .dout(n904));
    jor g0223(.dinb(n15762), .dina(n904), .dout(n908));
    jand g0224(.dinb(n15760), .dina(n908), .dout(n912));
    jand g0225(.dinb(G35gat), .dina(G375gat), .dout(n916));
    jnot g0226(.din(n916), .dout(n919));
    jand g0227(.dinb(n738), .dina(n16975), .dout(n923));
    jand g0228(.dinb(n16972), .dina(n844), .dout(n927));
    jor g0229(.dinb(n16933), .dina(n927), .dout(n931));
    jand g0230(.dinb(G52gat), .dina(G358gat), .dout(n935));
    jnot g0231(.din(n935), .dout(n938));
    jand g0232(.dinb(n757), .dina(n18127), .dout(n942));
    jand g0233(.dinb(n18124), .dina(n836), .dout(n946));
    jor g0234(.dinb(n18094), .dina(n946), .dout(n950));
    jand g0235(.dinb(G69gat), .dina(G341gat), .dout(n954));
    jnot g0236(.din(n954), .dout(n957));
    jand g0237(.dinb(n775), .dina(n19246), .dout(n961));
    jand g0238(.dinb(n19243), .dina(n828), .dout(n965));
    jor g0239(.dinb(n19222), .dina(n965), .dout(n969));
    jand g0240(.dinb(G86gat), .dina(G324gat), .dout(n973));
    jnot g0241(.din(n973), .dout(n976));
    jnot g0242(.din(n809), .dout(n979));
    jand g0243(.dinb(n20323), .dina(n820), .dout(n983));
    jor g0244(.dinb(n20311), .dina(n983), .dout(n987));
    jand g0245(.dinb(G103gat), .dina(G307gat), .dout(n991));
    jnot g0246(.din(n991), .dout(n994));
    jand g0247(.dinb(G137gat), .dina(G273gat), .dout(n998));
    jor g0248(.dinb(n794), .dina(n998), .dout(n1002));
    jand g0249(.dinb(G137gat), .dina(G290gat), .dout(n1006));
    jand g0250(.dinb(n786), .dina(n1006), .dout(n1010));
    jnot g0251(.din(n1010), .dout(n1013));
    jand g0252(.dinb(n21415), .dina(n1013), .dout(n1017));
    jor g0253(.dinb(n21420), .dina(n1017), .dout(n1021));
    jand g0254(.dinb(n21417), .dina(n1013), .dout(n1025));
    jnot g0255(.din(n1025), .dout(n1028));
    jand g0256(.dinb(n1021), .dina(n1028), .dout(n1032));
    jxor g0257(.dinb(n21412), .dina(n1032), .dout(n1036));
    jxor g0258(.dinb(n987), .dina(n20308), .dout(n1040));
    jxor g0259(.dinb(n20305), .dina(n1040), .dout(n1044));
    jxor g0260(.dinb(n969), .dina(n19219), .dout(n1048));
    jxor g0261(.dinb(n19216), .dina(n1048), .dout(n1052));
    jxor g0262(.dinb(n950), .dina(n18091), .dout(n1056));
    jxor g0263(.dinb(n18088), .dina(n1056), .dout(n1060));
    jxor g0264(.dinb(n931), .dina(n16930), .dout(n1064));
    jxor g0265(.dinb(n16927), .dina(n1064), .dout(n1068));
    jnot g0266(.din(n1068), .dout(n1071));
    jxor g0267(.dinb(n912), .dina(n1071), .dout(n1075));
    jxor g0268(.dinb(n14308), .dina(n1075), .dout(n1079));
    jxor g0269(.dinb(n889), .dina(n14250), .dout(n1083));
    jxor g0270(.dinb(n11029), .dina(n1083), .dout(n1087));
    jand g0271(.dinb(G1gat), .dina(G426gat), .dout(n1091));
    jnot g0272(.din(n1091), .dout(n1094));
    jnot g0273(.din(n1079), .dout(n1097));
    jor g0274(.dinb(n889), .dina(n1097), .dout(n1101));
    jor g0275(.dinb(n14181), .dina(n1083), .dout(n1105));
    jand g0276(.dinb(n14179), .dina(n1105), .dout(n1109));
    jand g0277(.dinb(G18gat), .dina(G409gat), .dout(n1113));
    jnot g0278(.din(n1113), .dout(n1116));
    jor g0279(.dinb(n912), .dina(n1071), .dout(n1120));
    jxor g0280(.dinb(n912), .dina(n15756), .dout(n1124));
    jor g0281(.dinb(n15696), .dina(n1124), .dout(n1128));
    jand g0282(.dinb(n15694), .dina(n1128), .dout(n1132));
    jand g0283(.dinb(G35gat), .dina(G392gat), .dout(n1136));
    jnot g0284(.din(n1136), .dout(n1139));
    jand g0285(.dinb(n931), .dina(n16930), .dout(n1143));
    jand g0286(.dinb(n16927), .dina(n1064), .dout(n1147));
    jor g0287(.dinb(n16879), .dina(n1147), .dout(n1151));
    jand g0288(.dinb(G52gat), .dina(G375gat), .dout(n1155));
    jnot g0289(.din(n1155), .dout(n1158));
    jand g0290(.dinb(n950), .dina(n18091), .dout(n1162));
    jand g0291(.dinb(n18088), .dina(n1056), .dout(n1166));
    jor g0292(.dinb(n18049), .dina(n1166), .dout(n1170));
    jand g0293(.dinb(G69gat), .dina(G358gat), .dout(n1174));
    jnot g0294(.din(n1174), .dout(n1177));
    jand g0295(.dinb(n969), .dina(n19219), .dout(n1181));
    jand g0296(.dinb(n19216), .dina(n1048), .dout(n1185));
    jor g0297(.dinb(n19186), .dina(n1185), .dout(n1189));
    jand g0298(.dinb(G86gat), .dina(G341gat), .dout(n1193));
    jnot g0299(.din(n1193), .dout(n1196));
    jand g0300(.dinb(n987), .dina(n20308), .dout(n1200));
    jand g0301(.dinb(n20305), .dina(n1040), .dout(n1204));
    jor g0302(.dinb(n20284), .dina(n1204), .dout(n1208));
    jand g0303(.dinb(G103gat), .dina(G324gat), .dout(n1212));
    jnot g0304(.din(n1212), .dout(n1215));
    jnot g0305(.din(n1021), .dout(n1218));
    jand g0306(.dinb(n21412), .dina(n1032), .dout(n1222));
    jor g0307(.dinb(n21400), .dina(n1222), .dout(n1226));
    jand g0308(.dinb(G120gat), .dina(G307gat), .dout(n1230));
    jand g0309(.dinb(G154gat), .dina(G273gat), .dout(n1234));
    jor g0310(.dinb(n1006), .dina(n1234), .dout(n1238));
    jand g0311(.dinb(G154gat), .dina(G290gat), .dout(n1242));
    jand g0312(.dinb(n998), .dina(n1242), .dout(n1246));
    jnot g0313(.din(n1246), .dout(n1249));
    jand g0314(.dinb(n22603), .dina(n1249), .dout(n1253));
    jor g0315(.dinb(n22608), .dina(n1253), .dout(n1257));
    jnot g0316(.din(n1257), .dout(n1260));
    jand g0317(.dinb(n22605), .dina(n1249), .dout(n1264));
    jor g0318(.dinb(n1260), .dina(n22591), .dout(n1268));
    jxor g0319(.dinb(n22614), .dina(n1268), .dout(n1272));
    jxor g0320(.dinb(n1226), .dina(n1272), .dout(n1276));
    jxor g0321(.dinb(n21397), .dina(n1276), .dout(n1280));
    jxor g0322(.dinb(n1208), .dina(n20281), .dout(n1284));
    jxor g0323(.dinb(n20278), .dina(n1284), .dout(n1288));
    jxor g0324(.dinb(n1189), .dina(n19183), .dout(n1292));
    jxor g0325(.dinb(n19180), .dina(n1292), .dout(n1296));
    jxor g0326(.dinb(n1170), .dina(n18046), .dout(n1300));
    jxor g0327(.dinb(n18043), .dina(n1300), .dout(n1304));
    jxor g0328(.dinb(n1151), .dina(n16876), .dout(n1308));
    jxor g0329(.dinb(n16873), .dina(n1308), .dout(n1312));
    jnot g0330(.din(n1312), .dout(n1315));
    jxor g0331(.dinb(n1132), .dina(n1315), .dout(n1319));
    jxor g0332(.dinb(n14176), .dina(n1319), .dout(n1323));
    jxor g0333(.dinb(n1109), .dina(n14109), .dout(n1327));
    jxor g0334(.dinb(n11104), .dina(n1327), .dout(n1331));
    jand g0335(.dinb(G1gat), .dina(G443gat), .dout(n1335));
    jnot g0336(.din(n1335), .dout(n1338));
    jnot g0337(.din(n1323), .dout(n1341));
    jor g0338(.dinb(n1109), .dina(n1341), .dout(n1345));
    jor g0339(.dinb(n14031), .dina(n1327), .dout(n1349));
    jand g0340(.dinb(n14029), .dina(n1349), .dout(n1353));
    jand g0341(.dinb(G18gat), .dina(G426gat), .dout(n1357));
    jnot g0342(.din(n1357), .dout(n1360));
    jor g0343(.dinb(n1132), .dina(n1315), .dout(n1364));
    jxor g0344(.dinb(n1132), .dina(n15690), .dout(n1368));
    jor g0345(.dinb(n15621), .dina(n1368), .dout(n1372));
    jand g0346(.dinb(n15619), .dina(n1372), .dout(n1376));
    jand g0347(.dinb(G35gat), .dina(G409gat), .dout(n1380));
    jnot g0348(.din(n1380), .dout(n1383));
    jand g0349(.dinb(n1151), .dina(n16876), .dout(n1387));
    jand g0350(.dinb(n16873), .dina(n1308), .dout(n1391));
    jor g0351(.dinb(n16816), .dina(n1391), .dout(n1395));
    jand g0352(.dinb(G52gat), .dina(G392gat), .dout(n1399));
    jnot g0353(.din(n1399), .dout(n1402));
    jand g0354(.dinb(n1170), .dina(n18046), .dout(n1406));
    jand g0355(.dinb(n18043), .dina(n1300), .dout(n1410));
    jor g0356(.dinb(n17995), .dina(n1410), .dout(n1414));
    jand g0357(.dinb(G69gat), .dina(G375gat), .dout(n1418));
    jnot g0358(.din(n1418), .dout(n1421));
    jand g0359(.dinb(n1189), .dina(n19183), .dout(n1425));
    jand g0360(.dinb(n19180), .dina(n1292), .dout(n1429));
    jor g0361(.dinb(n19141), .dina(n1429), .dout(n1433));
    jand g0362(.dinb(G86gat), .dina(G358gat), .dout(n1437));
    jnot g0363(.din(n1437), .dout(n1440));
    jand g0364(.dinb(n1208), .dina(n20281), .dout(n1444));
    jand g0365(.dinb(n20278), .dina(n1284), .dout(n1448));
    jor g0366(.dinb(n20248), .dina(n1448), .dout(n1452));
    jand g0367(.dinb(G103gat), .dina(G341gat), .dout(n1456));
    jnot g0368(.din(n1456), .dout(n1459));
    jand g0369(.dinb(n1226), .dina(n1272), .dout(n1463));
    jand g0370(.dinb(n21397), .dina(n1276), .dout(n1467));
    jor g0371(.dinb(n21376), .dina(n1467), .dout(n1471));
    jand g0372(.dinb(G120gat), .dina(G324gat), .dout(n1475));
    jnot g0373(.din(n1475), .dout(n1478));
    jnot g0374(.din(n1230), .dout(n1481));
    jnot g0375(.din(n1268), .dout(n1484));
    jand g0376(.dinb(n22585), .dina(n1484), .dout(n1488));
    jor g0377(.dinb(n22593), .dina(n1488), .dout(n1492));
    jand g0378(.dinb(G137gat), .dina(G307gat), .dout(n1496));
    jand g0379(.dinb(G171gat), .dina(G273gat), .dout(n1500));
    jor g0380(.dinb(n1242), .dina(n1500), .dout(n1504));
    jand g0381(.dinb(G171gat), .dina(G290gat), .dout(n1508));
    jand g0382(.dinb(n1234), .dina(n1508), .dout(n1512));
    jnot g0383(.din(n1512), .dout(n1515));
    jand g0384(.dinb(n23809), .dina(n1515), .dout(n1519));
    jor g0385(.dinb(n23814), .dina(n1519), .dout(n1523));
    jnot g0386(.din(n1523), .dout(n1526));
    jand g0387(.dinb(n23811), .dina(n1515), .dout(n1530));
    jor g0388(.dinb(n1526), .dina(n23797), .dout(n1534));
    jxor g0389(.dinb(n23820), .dina(n1534), .dout(n1538));
    jxor g0390(.dinb(n1492), .dina(n22567), .dout(n1542));
    jxor g0391(.dinb(n22561), .dina(n1542), .dout(n1546));
    jxor g0392(.dinb(n21373), .dina(n1546), .dout(n1550));
    jxor g0393(.dinb(n21370), .dina(n1550), .dout(n1554));
    jxor g0394(.dinb(n1452), .dina(n1554), .dout(n1558));
    jxor g0395(.dinb(n20245), .dina(n1558), .dout(n1562));
    jxor g0396(.dinb(n1433), .dina(n19138), .dout(n1566));
    jxor g0397(.dinb(n19135), .dina(n1566), .dout(n1570));
    jxor g0398(.dinb(n1414), .dina(n17992), .dout(n1574));
    jxor g0399(.dinb(n17989), .dina(n1574), .dout(n1578));
    jxor g0400(.dinb(n1395), .dina(n16813), .dout(n1582));
    jxor g0401(.dinb(n16810), .dina(n1582), .dout(n1586));
    jnot g0402(.din(n1586), .dout(n1589));
    jxor g0403(.dinb(n1376), .dina(n1589), .dout(n1593));
    jxor g0404(.dinb(n14026), .dina(n1593), .dout(n1597));
    jxor g0405(.dinb(n1353), .dina(n13950), .dout(n1601));
    jxor g0406(.dinb(n11188), .dina(n1601), .dout(n1605));
    jand g0407(.dinb(G1gat), .dina(G460gat), .dout(n1609));
    jnot g0408(.din(n1609), .dout(n1612));
    jnot g0409(.din(n1597), .dout(n1615));
    jor g0410(.dinb(n1353), .dina(n1615), .dout(n1619));
    jor g0411(.dinb(n13863), .dina(n1601), .dout(n1623));
    jand g0412(.dinb(n13861), .dina(n1623), .dout(n1627));
    jand g0413(.dinb(G18gat), .dina(G443gat), .dout(n1631));
    jnot g0414(.din(n1631), .dout(n1634));
    jor g0415(.dinb(n1376), .dina(n1589), .dout(n1638));
    jxor g0416(.dinb(n1376), .dina(n15615), .dout(n1642));
    jor g0417(.dinb(n15537), .dina(n1642), .dout(n1646));
    jand g0418(.dinb(n15535), .dina(n1646), .dout(n1650));
    jand g0419(.dinb(G35gat), .dina(G426gat), .dout(n1654));
    jnot g0420(.din(n1654), .dout(n1657));
    jand g0421(.dinb(n1395), .dina(n16813), .dout(n1661));
    jand g0422(.dinb(n16810), .dina(n1582), .dout(n1665));
    jor g0423(.dinb(n16744), .dina(n1665), .dout(n1669));
    jand g0424(.dinb(G52gat), .dina(G409gat), .dout(n1673));
    jnot g0425(.din(n1673), .dout(n1676));
    jand g0426(.dinb(n1414), .dina(n17992), .dout(n1680));
    jand g0427(.dinb(n17989), .dina(n1574), .dout(n1684));
    jor g0428(.dinb(n17932), .dina(n1684), .dout(n1688));
    jand g0429(.dinb(G69gat), .dina(G392gat), .dout(n1692));
    jnot g0430(.din(n1692), .dout(n1695));
    jand g0431(.dinb(n1433), .dina(n19138), .dout(n1699));
    jand g0432(.dinb(n19135), .dina(n1566), .dout(n1703));
    jor g0433(.dinb(n19087), .dina(n1703), .dout(n1707));
    jand g0434(.dinb(G86gat), .dina(G375gat), .dout(n1711));
    jnot g0435(.din(n1711), .dout(n1714));
    jand g0436(.dinb(n1452), .dina(n1554), .dout(n1718));
    jand g0437(.dinb(n20245), .dina(n1558), .dout(n1722));
    jor g0438(.dinb(n20206), .dina(n1722), .dout(n1726));
    jand g0439(.dinb(G103gat), .dina(G358gat), .dout(n1730));
    jnot g0440(.din(n1730), .dout(n1733));
    jand g0441(.dinb(n21373), .dina(n1546), .dout(n1737));
    jand g0442(.dinb(n21370), .dina(n1550), .dout(n1741));
    jor g0443(.dinb(n21337), .dina(n1741), .dout(n1745));
    jand g0444(.dinb(G120gat), .dina(G341gat), .dout(n1749));
    jnot g0445(.din(n1749), .dout(n1752));
    jand g0446(.dinb(n1492), .dina(n22567), .dout(n1756));
    jand g0447(.dinb(n22561), .dina(n1542), .dout(n1760));
    jor g0448(.dinb(n22534), .dina(n1760), .dout(n1764));
    jand g0449(.dinb(G137gat), .dina(G324gat), .dout(n1768));
    jnot g0450(.din(n1768), .dout(n1771));
    jnot g0451(.din(n1496), .dout(n1774));
    jnot g0452(.din(n1534), .dout(n1777));
    jand g0453(.dinb(n23791), .dina(n1777), .dout(n1781));
    jor g0454(.dinb(n23799), .dina(n1781), .dout(n1785));
    jand g0455(.dinb(G154gat), .dina(G307gat), .dout(n1789));
    jand g0456(.dinb(G188gat), .dina(G273gat), .dout(n1793));
    jor g0457(.dinb(n1508), .dina(n1793), .dout(n1797));
    jand g0458(.dinb(G188gat), .dina(G290gat), .dout(n1801));
    jand g0459(.dinb(n1500), .dina(n1801), .dout(n1805));
    jnot g0460(.din(n1805), .dout(n1808));
    jand g0461(.dinb(n25024), .dina(n1808), .dout(n1812));
    jor g0462(.dinb(n25029), .dina(n1812), .dout(n1816));
    jnot g0463(.din(n1816), .dout(n1819));
    jand g0464(.dinb(n25026), .dina(n1808), .dout(n1823));
    jor g0465(.dinb(n1819), .dina(n25012), .dout(n1827));
    jxor g0466(.dinb(n25035), .dina(n1827), .dout(n1831));
    jxor g0467(.dinb(n1785), .dina(n23773), .dout(n1835));
    jxor g0468(.dinb(n23767), .dina(n1835), .dout(n1839));
    jxor g0469(.dinb(n1764), .dina(n22531), .dout(n1843));
    jxor g0470(.dinb(n22528), .dina(n1843), .dout(n1847));
    jxor g0471(.dinb(n1745), .dina(n1847), .dout(n1851));
    jxor g0472(.dinb(n21334), .dina(n1851), .dout(n1855));
    jxor g0473(.dinb(n1726), .dina(n1855), .dout(n1859));
    jxor g0474(.dinb(n20203), .dina(n1859), .dout(n1863));
    jxor g0475(.dinb(n1707), .dina(n19084), .dout(n1867));
    jxor g0476(.dinb(n19081), .dina(n1867), .dout(n1871));
    jxor g0477(.dinb(n1688), .dina(n17929), .dout(n1875));
    jxor g0478(.dinb(n17926), .dina(n1875), .dout(n1879));
    jxor g0479(.dinb(n1669), .dina(n16741), .dout(n1883));
    jxor g0480(.dinb(n16738), .dina(n1883), .dout(n1887));
    jnot g0481(.din(n1887), .dout(n1890));
    jxor g0482(.dinb(n1650), .dina(n1890), .dout(n1894));
    jxor g0483(.dinb(n13858), .dina(n1894), .dout(n1898));
    jxor g0484(.dinb(n1627), .dina(n13773), .dout(n1902));
    jxor g0485(.dinb(n11281), .dina(n1902), .dout(n1906));
    jand g0486(.dinb(G1gat), .dina(G477gat), .dout(n1910));
    jnot g0487(.din(n1910), .dout(n1913));
    jnot g0488(.din(n1898), .dout(n1916));
    jor g0489(.dinb(n1627), .dina(n1916), .dout(n1920));
    jor g0490(.dinb(n13677), .dina(n1902), .dout(n1924));
    jand g0491(.dinb(n13675), .dina(n1924), .dout(n1928));
    jand g0492(.dinb(G18gat), .dina(G460gat), .dout(n1932));
    jnot g0493(.din(n1932), .dout(n1935));
    jor g0494(.dinb(n1650), .dina(n1890), .dout(n1939));
    jxor g0495(.dinb(n1650), .dina(n15531), .dout(n1943));
    jor g0496(.dinb(n15444), .dina(n1943), .dout(n1947));
    jand g0497(.dinb(n15442), .dina(n1947), .dout(n1951));
    jand g0498(.dinb(G35gat), .dina(G443gat), .dout(n1955));
    jnot g0499(.din(n1955), .dout(n1958));
    jand g0500(.dinb(n1669), .dina(n16741), .dout(n1962));
    jand g0501(.dinb(n16738), .dina(n1883), .dout(n1966));
    jor g0502(.dinb(n16663), .dina(n1966), .dout(n1970));
    jand g0503(.dinb(G52gat), .dina(G426gat), .dout(n1974));
    jnot g0504(.din(n1974), .dout(n1977));
    jand g0505(.dinb(n1688), .dina(n17929), .dout(n1981));
    jand g0506(.dinb(n17926), .dina(n1875), .dout(n1985));
    jor g0507(.dinb(n17860), .dina(n1985), .dout(n1989));
    jand g0508(.dinb(G69gat), .dina(G409gat), .dout(n1993));
    jnot g0509(.din(n1993), .dout(n1996));
    jand g0510(.dinb(n1707), .dina(n19084), .dout(n2000));
    jand g0511(.dinb(n19081), .dina(n1867), .dout(n2004));
    jor g0512(.dinb(n19024), .dina(n2004), .dout(n2008));
    jand g0513(.dinb(G86gat), .dina(G392gat), .dout(n2012));
    jnot g0514(.din(n2012), .dout(n2015));
    jand g0515(.dinb(n1726), .dina(n1855), .dout(n2019));
    jand g0516(.dinb(n20203), .dina(n1859), .dout(n2023));
    jor g0517(.dinb(n20155), .dina(n2023), .dout(n2027));
    jand g0518(.dinb(G103gat), .dina(G375gat), .dout(n2031));
    jnot g0519(.din(n2031), .dout(n2034));
    jand g0520(.dinb(n1745), .dina(n1847), .dout(n2038));
    jand g0521(.dinb(n21334), .dina(n1851), .dout(n2042));
    jor g0522(.dinb(n21292), .dina(n2042), .dout(n2046));
    jand g0523(.dinb(G120gat), .dina(G358gat), .dout(n2050));
    jnot g0524(.din(n2050), .dout(n2053));
    jand g0525(.dinb(n1764), .dina(n22531), .dout(n2057));
    jand g0526(.dinb(n22528), .dina(n1843), .dout(n2061));
    jor g0527(.dinb(n22492), .dina(n2061), .dout(n2065));
    jand g0528(.dinb(G137gat), .dina(G341gat), .dout(n2069));
    jnot g0529(.din(n2069), .dout(n2072));
    jand g0530(.dinb(n1785), .dina(n23773), .dout(n2076));
    jand g0531(.dinb(n23767), .dina(n1835), .dout(n2080));
    jor g0532(.dinb(n23740), .dina(n2080), .dout(n2084));
    jand g0533(.dinb(G154gat), .dina(G324gat), .dout(n2088));
    jnot g0534(.din(n2088), .dout(n2091));
    jnot g0535(.din(n1789), .dout(n2094));
    jnot g0536(.din(n1827), .dout(n2097));
    jand g0537(.dinb(n25006), .dina(n2097), .dout(n2101));
    jor g0538(.dinb(n25014), .dina(n2101), .dout(n2105));
    jand g0539(.dinb(G171gat), .dina(G307gat), .dout(n2109));
    jand g0540(.dinb(G205gat), .dina(G273gat), .dout(n2113));
    jor g0541(.dinb(n1801), .dina(n2113), .dout(n2117));
    jand g0542(.dinb(G205gat), .dina(G290gat), .dout(n2121));
    jand g0543(.dinb(n1793), .dina(n2121), .dout(n2125));
    jnot g0544(.din(n2125), .dout(n2128));
    jand g0545(.dinb(n26254), .dina(n2128), .dout(n2132));
    jor g0546(.dinb(n26259), .dina(n2132), .dout(n2136));
    jnot g0547(.din(n2136), .dout(n2139));
    jand g0548(.dinb(n26256), .dina(n2128), .dout(n2143));
    jor g0549(.dinb(n2139), .dina(n26242), .dout(n2147));
    jxor g0550(.dinb(n26265), .dina(n2147), .dout(n2151));
    jxor g0551(.dinb(n2105), .dina(n24988), .dout(n2155));
    jxor g0552(.dinb(n24982), .dina(n2155), .dout(n2159));
    jxor g0553(.dinb(n2084), .dina(n23737), .dout(n2163));
    jxor g0554(.dinb(n23734), .dina(n2163), .dout(n2167));
    jxor g0555(.dinb(n2065), .dina(n22489), .dout(n2171));
    jxor g0556(.dinb(n22486), .dina(n2171), .dout(n2175));
    jxor g0557(.dinb(n2046), .dina(n2175), .dout(n2179));
    jxor g0558(.dinb(n21289), .dina(n2179), .dout(n2183));
    jxor g0559(.dinb(n2027), .dina(n2183), .dout(n2187));
    jxor g0560(.dinb(n20152), .dina(n2187), .dout(n2191));
    jxor g0561(.dinb(n2008), .dina(n19021), .dout(n2195));
    jxor g0562(.dinb(n19018), .dina(n2195), .dout(n2199));
    jxor g0563(.dinb(n1989), .dina(n17857), .dout(n2203));
    jxor g0564(.dinb(n17854), .dina(n2203), .dout(n2207));
    jxor g0565(.dinb(n1970), .dina(n16660), .dout(n2211));
    jxor g0566(.dinb(n16657), .dina(n2211), .dout(n2215));
    jnot g0567(.din(n2215), .dout(n2218));
    jxor g0568(.dinb(n1951), .dina(n2218), .dout(n2222));
    jxor g0569(.dinb(n13672), .dina(n2222), .dout(n2226));
    jxor g0570(.dinb(n1928), .dina(n13578), .dout(n2230));
    jxor g0571(.dinb(n11383), .dina(n2230), .dout(n2234));
    jand g0572(.dinb(G1gat), .dina(G494gat), .dout(n2238));
    jnot g0573(.din(n2238), .dout(n2241));
    jnot g0574(.din(n2226), .dout(n2244));
    jor g0575(.dinb(n1928), .dina(n2244), .dout(n2248));
    jor g0576(.dinb(n13473), .dina(n2230), .dout(n2252));
    jand g0577(.dinb(n13471), .dina(n2252), .dout(n2256));
    jand g0578(.dinb(G18gat), .dina(G477gat), .dout(n2260));
    jnot g0579(.din(n2260), .dout(n2263));
    jor g0580(.dinb(n1951), .dina(n2218), .dout(n2267));
    jxor g0581(.dinb(n1951), .dina(n15438), .dout(n2271));
    jor g0582(.dinb(n15342), .dina(n2271), .dout(n2275));
    jand g0583(.dinb(n15340), .dina(n2275), .dout(n2279));
    jand g0584(.dinb(G35gat), .dina(G460gat), .dout(n2283));
    jnot g0585(.din(n2283), .dout(n2286));
    jand g0586(.dinb(n1970), .dina(n16660), .dout(n2290));
    jand g0587(.dinb(n16657), .dina(n2211), .dout(n2294));
    jor g0588(.dinb(n16573), .dina(n2294), .dout(n2298));
    jand g0589(.dinb(G52gat), .dina(G443gat), .dout(n2302));
    jnot g0590(.din(n2302), .dout(n2305));
    jand g0591(.dinb(n1989), .dina(n17857), .dout(n2309));
    jand g0592(.dinb(n17854), .dina(n2203), .dout(n2313));
    jor g0593(.dinb(n17779), .dina(n2313), .dout(n2317));
    jand g0594(.dinb(G69gat), .dina(G426gat), .dout(n2321));
    jnot g0595(.din(n2321), .dout(n2324));
    jand g0596(.dinb(n2008), .dina(n19021), .dout(n2328));
    jand g0597(.dinb(n19018), .dina(n2195), .dout(n2332));
    jor g0598(.dinb(n18952), .dina(n2332), .dout(n2336));
    jand g0599(.dinb(G86gat), .dina(G409gat), .dout(n2340));
    jnot g0600(.din(n2340), .dout(n2343));
    jand g0601(.dinb(n2027), .dina(n2183), .dout(n2347));
    jand g0602(.dinb(n20152), .dina(n2187), .dout(n2351));
    jor g0603(.dinb(n20095), .dina(n2351), .dout(n2355));
    jand g0604(.dinb(G103gat), .dina(G392gat), .dout(n2359));
    jnot g0605(.din(n2359), .dout(n2362));
    jand g0606(.dinb(n2046), .dina(n2175), .dout(n2366));
    jand g0607(.dinb(n21289), .dina(n2179), .dout(n2370));
    jor g0608(.dinb(n21238), .dina(n2370), .dout(n2374));
    jand g0609(.dinb(G120gat), .dina(G375gat), .dout(n2378));
    jnot g0610(.din(n2378), .dout(n2381));
    jand g0611(.dinb(n2065), .dina(n22489), .dout(n2385));
    jand g0612(.dinb(n22486), .dina(n2171), .dout(n2389));
    jor g0613(.dinb(n22441), .dina(n2389), .dout(n2393));
    jand g0614(.dinb(G137gat), .dina(G358gat), .dout(n2397));
    jnot g0615(.din(n2397), .dout(n2400));
    jand g0616(.dinb(n2084), .dina(n23737), .dout(n2404));
    jand g0617(.dinb(n23734), .dina(n2163), .dout(n2408));
    jor g0618(.dinb(n23698), .dina(n2408), .dout(n2412));
    jand g0619(.dinb(G154gat), .dina(G341gat), .dout(n2416));
    jnot g0620(.din(n2416), .dout(n2419));
    jand g0621(.dinb(n2105), .dina(n24988), .dout(n2423));
    jand g0622(.dinb(n24982), .dina(n2155), .dout(n2427));
    jor g0623(.dinb(n24955), .dina(n2427), .dout(n2431));
    jand g0624(.dinb(G171gat), .dina(G324gat), .dout(n2435));
    jnot g0625(.din(n2435), .dout(n2438));
    jnot g0626(.din(n2109), .dout(n2441));
    jnot g0627(.din(n2147), .dout(n2444));
    jand g0628(.dinb(n26236), .dina(n2444), .dout(n2448));
    jor g0629(.dinb(n26244), .dina(n2448), .dout(n2452));
    jand g0630(.dinb(G188gat), .dina(G307gat), .dout(n2456));
    jand g0631(.dinb(G222gat), .dina(G273gat), .dout(n2460));
    jor g0632(.dinb(n2121), .dina(n2460), .dout(n2464));
    jand g0633(.dinb(G222gat), .dina(G290gat), .dout(n2468));
    jand g0634(.dinb(n2113), .dina(n2468), .dout(n2472));
    jnot g0635(.din(n2472), .dout(n2475));
    jand g0636(.dinb(n27517), .dina(n2475), .dout(n2479));
    jor g0637(.dinb(n27522), .dina(n2479), .dout(n2483));
    jnot g0638(.din(n2483), .dout(n2486));
    jand g0639(.dinb(n27519), .dina(n2475), .dout(n2490));
    jor g0640(.dinb(n2486), .dina(n27505), .dout(n2494));
    jxor g0641(.dinb(n27528), .dina(n2494), .dout(n2498));
    jxor g0642(.dinb(n2452), .dina(n26218), .dout(n2502));
    jxor g0643(.dinb(n26212), .dina(n2502), .dout(n2506));
    jxor g0644(.dinb(n2431), .dina(n24952), .dout(n2510));
    jxor g0645(.dinb(n24949), .dina(n2510), .dout(n2514));
    jxor g0646(.dinb(n2412), .dina(n23695), .dout(n2518));
    jxor g0647(.dinb(n23692), .dina(n2518), .dout(n2522));
    jxor g0648(.dinb(n2393), .dina(n22438), .dout(n2526));
    jxor g0649(.dinb(n22435), .dina(n2526), .dout(n2530));
    jxor g0650(.dinb(n2374), .dina(n2530), .dout(n2534));
    jxor g0651(.dinb(n21235), .dina(n2534), .dout(n2538));
    jxor g0652(.dinb(n2355), .dina(n2538), .dout(n2542));
    jxor g0653(.dinb(n20092), .dina(n2542), .dout(n2546));
    jxor g0654(.dinb(n2336), .dina(n18949), .dout(n2550));
    jxor g0655(.dinb(n18946), .dina(n2550), .dout(n2554));
    jxor g0656(.dinb(n2317), .dina(n17776), .dout(n2558));
    jxor g0657(.dinb(n17773), .dina(n2558), .dout(n2562));
    jxor g0658(.dinb(n2298), .dina(n16570), .dout(n2566));
    jxor g0659(.dinb(n16567), .dina(n2566), .dout(n2570));
    jnot g0660(.din(n2570), .dout(n2573));
    jxor g0661(.dinb(n2279), .dina(n2573), .dout(n2577));
    jxor g0662(.dinb(n13468), .dina(n2577), .dout(n2581));
    jxor g0663(.dinb(n2256), .dina(n13365), .dout(n2585));
    jxor g0664(.dinb(n11494), .dina(n2585), .dout(n2589));
    jand g0665(.dinb(G1gat), .dina(G511gat), .dout(n2593));
    jnot g0666(.din(n2593), .dout(n2596));
    jnot g0667(.din(n2581), .dout(n2599));
    jor g0668(.dinb(n2256), .dina(n2599), .dout(n2603));
    jor g0669(.dinb(n13251), .dina(n2585), .dout(n2607));
    jand g0670(.dinb(n13249), .dina(n2607), .dout(n2611));
    jand g0671(.dinb(G18gat), .dina(G494gat), .dout(n2615));
    jnot g0672(.din(n2615), .dout(n2618));
    jor g0673(.dinb(n2279), .dina(n2573), .dout(n2622));
    jxor g0674(.dinb(n2279), .dina(n15336), .dout(n2626));
    jor g0675(.dinb(n15231), .dina(n2626), .dout(n2630));
    jand g0676(.dinb(n15229), .dina(n2630), .dout(n2634));
    jand g0677(.dinb(G35gat), .dina(G477gat), .dout(n2638));
    jnot g0678(.din(n2638), .dout(n2641));
    jand g0679(.dinb(n2298), .dina(n16570), .dout(n2645));
    jand g0680(.dinb(n16567), .dina(n2566), .dout(n2649));
    jor g0681(.dinb(n16474), .dina(n2649), .dout(n2653));
    jand g0682(.dinb(G52gat), .dina(G460gat), .dout(n2657));
    jnot g0683(.din(n2657), .dout(n2660));
    jand g0684(.dinb(n2317), .dina(n17776), .dout(n2664));
    jand g0685(.dinb(n17773), .dina(n2558), .dout(n2668));
    jor g0686(.dinb(n17689), .dina(n2668), .dout(n2672));
    jand g0687(.dinb(G69gat), .dina(G443gat), .dout(n2676));
    jnot g0688(.din(n2676), .dout(n2679));
    jand g0689(.dinb(n2336), .dina(n18949), .dout(n2683));
    jand g0690(.dinb(n18946), .dina(n2550), .dout(n2687));
    jor g0691(.dinb(n18871), .dina(n2687), .dout(n2691));
    jand g0692(.dinb(G86gat), .dina(G426gat), .dout(n2695));
    jnot g0693(.din(n2695), .dout(n2698));
    jand g0694(.dinb(n2355), .dina(n2538), .dout(n2702));
    jand g0695(.dinb(n20092), .dina(n2542), .dout(n2706));
    jor g0696(.dinb(n20026), .dina(n2706), .dout(n2710));
    jand g0697(.dinb(G103gat), .dina(G409gat), .dout(n2714));
    jnot g0698(.din(n2714), .dout(n2717));
    jand g0699(.dinb(n2374), .dina(n2530), .dout(n2721));
    jand g0700(.dinb(n21235), .dina(n2534), .dout(n2725));
    jor g0701(.dinb(n21175), .dina(n2725), .dout(n2729));
    jand g0702(.dinb(G120gat), .dina(G392gat), .dout(n2733));
    jnot g0703(.din(n2733), .dout(n2736));
    jand g0704(.dinb(n2393), .dina(n22438), .dout(n2740));
    jand g0705(.dinb(n22435), .dina(n2526), .dout(n2744));
    jor g0706(.dinb(n22381), .dina(n2744), .dout(n2748));
    jand g0707(.dinb(G137gat), .dina(G375gat), .dout(n2752));
    jnot g0708(.din(n2752), .dout(n2755));
    jand g0709(.dinb(n2412), .dina(n23695), .dout(n2759));
    jand g0710(.dinb(n23692), .dina(n2518), .dout(n2763));
    jor g0711(.dinb(n23647), .dina(n2763), .dout(n2767));
    jand g0712(.dinb(G154gat), .dina(G358gat), .dout(n2771));
    jnot g0713(.din(n2771), .dout(n2774));
    jand g0714(.dinb(n2431), .dina(n24952), .dout(n2778));
    jand g0715(.dinb(n24949), .dina(n2510), .dout(n2782));
    jor g0716(.dinb(n24913), .dina(n2782), .dout(n2786));
    jand g0717(.dinb(G171gat), .dina(G341gat), .dout(n2790));
    jnot g0718(.din(n2790), .dout(n2793));
    jand g0719(.dinb(n2452), .dina(n26218), .dout(n2797));
    jand g0720(.dinb(n26212), .dina(n2502), .dout(n2801));
    jor g0721(.dinb(n26185), .dina(n2801), .dout(n2805));
    jand g0722(.dinb(G188gat), .dina(G324gat), .dout(n2809));
    jnot g0723(.din(n2809), .dout(n2812));
    jnot g0724(.din(n2456), .dout(n2815));
    jnot g0725(.din(n2494), .dout(n2818));
    jand g0726(.dinb(n27499), .dina(n2818), .dout(n2822));
    jor g0727(.dinb(n27507), .dina(n2822), .dout(n2826));
    jand g0728(.dinb(G205gat), .dina(G307gat), .dout(n2830));
    jand g0729(.dinb(G239gat), .dina(G273gat), .dout(n2834));
    jor g0730(.dinb(n2468), .dina(n2834), .dout(n2838));
    jand g0731(.dinb(G239gat), .dina(G290gat), .dout(n2842));
    jand g0732(.dinb(n2460), .dina(n2842), .dout(n2846));
    jnot g0733(.din(n2846), .dout(n2849));
    jand g0734(.dinb(n28834), .dina(n2849), .dout(n2853));
    jor g0735(.dinb(n28839), .dina(n2853), .dout(n2857));
    jnot g0736(.din(n2857), .dout(n2860));
    jand g0737(.dinb(n28836), .dina(n2849), .dout(n2864));
    jor g0738(.dinb(n2860), .dina(n28822), .dout(n2868));
    jxor g0739(.dinb(n28845), .dina(n2868), .dout(n2872));
    jxor g0740(.dinb(n2826), .dina(n27481), .dout(n2876));
    jxor g0741(.dinb(n27475), .dina(n2876), .dout(n2880));
    jxor g0742(.dinb(n2805), .dina(n26182), .dout(n2884));
    jxor g0743(.dinb(n26179), .dina(n2884), .dout(n2888));
    jxor g0744(.dinb(n2786), .dina(n24910), .dout(n2892));
    jxor g0745(.dinb(n24907), .dina(n2892), .dout(n2896));
    jxor g0746(.dinb(n2767), .dina(n23644), .dout(n2900));
    jxor g0747(.dinb(n23641), .dina(n2900), .dout(n2904));
    jxor g0748(.dinb(n2748), .dina(n22378), .dout(n2908));
    jxor g0749(.dinb(n22375), .dina(n2908), .dout(n2912));
    jxor g0750(.dinb(n2729), .dina(n2912), .dout(n2916));
    jxor g0751(.dinb(n21172), .dina(n2916), .dout(n2920));
    jxor g0752(.dinb(n2710), .dina(n2920), .dout(n2924));
    jxor g0753(.dinb(n20023), .dina(n2924), .dout(n2928));
    jxor g0754(.dinb(n2691), .dina(n18868), .dout(n2932));
    jxor g0755(.dinb(n18865), .dina(n2932), .dout(n2936));
    jxor g0756(.dinb(n2672), .dina(n17686), .dout(n2940));
    jxor g0757(.dinb(n17683), .dina(n2940), .dout(n2944));
    jxor g0758(.dinb(n2653), .dina(n16471), .dout(n2948));
    jxor g0759(.dinb(n16468), .dina(n2948), .dout(n2952));
    jnot g0760(.din(n2952), .dout(n2955));
    jxor g0761(.dinb(n2634), .dina(n2955), .dout(n2959));
    jxor g0762(.dinb(n13246), .dina(n2959), .dout(n2963));
    jxor g0763(.dinb(n2611), .dina(n13134), .dout(n2967));
    jxor g0764(.dinb(n11614), .dina(n2967), .dout(n2971));
    jand g0765(.dinb(G1gat), .dina(G528gat), .dout(n2975));
    jnot g0766(.din(n2975), .dout(n2978));
    jnot g0767(.din(n2963), .dout(n2981));
    jor g0768(.dinb(n2611), .dina(n2981), .dout(n2985));
    jor g0769(.dinb(n13011), .dina(n2967), .dout(n2989));
    jand g0770(.dinb(n13009), .dina(n2989), .dout(n2993));
    jand g0771(.dinb(G18gat), .dina(G511gat), .dout(n2997));
    jor g0772(.dinb(n2634), .dina(n2955), .dout(n3001));
    jxor g0773(.dinb(n2634), .dina(n15225), .dout(n3005));
    jor g0774(.dinb(n15111), .dina(n3005), .dout(n3009));
    jand g0775(.dinb(n15109), .dina(n3009), .dout(n3013));
    jand g0776(.dinb(G35gat), .dina(G494gat), .dout(n3017));
    jnot g0777(.din(n3017), .dout(n3020));
    jand g0778(.dinb(n2653), .dina(n16471), .dout(n3024));
    jand g0779(.dinb(n16468), .dina(n2948), .dout(n3028));
    jor g0780(.dinb(n16366), .dina(n3028), .dout(n3032));
    jand g0781(.dinb(G52gat), .dina(G477gat), .dout(n3036));
    jnot g0782(.din(n3036), .dout(n3039));
    jand g0783(.dinb(n2672), .dina(n17686), .dout(n3043));
    jand g0784(.dinb(n17683), .dina(n2940), .dout(n3047));
    jor g0785(.dinb(n17590), .dina(n3047), .dout(n3051));
    jand g0786(.dinb(G69gat), .dina(G460gat), .dout(n3055));
    jnot g0787(.din(n3055), .dout(n3058));
    jand g0788(.dinb(n2691), .dina(n18868), .dout(n3062));
    jand g0789(.dinb(n18865), .dina(n2932), .dout(n3066));
    jor g0790(.dinb(n18781), .dina(n3066), .dout(n3070));
    jand g0791(.dinb(G86gat), .dina(G443gat), .dout(n3074));
    jnot g0792(.din(n3074), .dout(n3077));
    jand g0793(.dinb(n2710), .dina(n2920), .dout(n3081));
    jand g0794(.dinb(n20023), .dina(n2924), .dout(n3085));
    jor g0795(.dinb(n19948), .dina(n3085), .dout(n3089));
    jand g0796(.dinb(G103gat), .dina(G426gat), .dout(n3093));
    jnot g0797(.din(n3093), .dout(n3096));
    jand g0798(.dinb(n2729), .dina(n2912), .dout(n3100));
    jand g0799(.dinb(n21172), .dina(n2916), .dout(n3104));
    jor g0800(.dinb(n21103), .dina(n3104), .dout(n3108));
    jand g0801(.dinb(G120gat), .dina(G409gat), .dout(n3112));
    jnot g0802(.din(n3112), .dout(n3115));
    jand g0803(.dinb(n2748), .dina(n22378), .dout(n3119));
    jand g0804(.dinb(n22375), .dina(n2908), .dout(n3123));
    jor g0805(.dinb(n22312), .dina(n3123), .dout(n3127));
    jand g0806(.dinb(G137gat), .dina(G392gat), .dout(n3131));
    jnot g0807(.din(n3131), .dout(n3134));
    jand g0808(.dinb(n2767), .dina(n23644), .dout(n3138));
    jand g0809(.dinb(n23641), .dina(n2900), .dout(n3142));
    jor g0810(.dinb(n23587), .dina(n3142), .dout(n3146));
    jand g0811(.dinb(G154gat), .dina(G375gat), .dout(n3150));
    jnot g0812(.din(n3150), .dout(n3153));
    jand g0813(.dinb(n2786), .dina(n24910), .dout(n3157));
    jand g0814(.dinb(n24907), .dina(n2892), .dout(n3161));
    jor g0815(.dinb(n24862), .dina(n3161), .dout(n3165));
    jand g0816(.dinb(G171gat), .dina(G358gat), .dout(n3169));
    jnot g0817(.din(n3169), .dout(n3172));
    jand g0818(.dinb(n2805), .dina(n26182), .dout(n3176));
    jand g0819(.dinb(n26179), .dina(n2884), .dout(n3180));
    jor g0820(.dinb(n26143), .dina(n3180), .dout(n3184));
    jand g0821(.dinb(G188gat), .dina(G341gat), .dout(n3188));
    jnot g0822(.din(n3188), .dout(n3191));
    jand g0823(.dinb(n2826), .dina(n27481), .dout(n3195));
    jand g0824(.dinb(n27475), .dina(n2876), .dout(n3199));
    jor g0825(.dinb(n27448), .dina(n3199), .dout(n3203));
    jand g0826(.dinb(G205gat), .dina(G324gat), .dout(n3207));
    jnot g0827(.din(n3207), .dout(n3210));
    jnot g0828(.din(n2830), .dout(n3213));
    jnot g0829(.din(n2868), .dout(n3216));
    jand g0830(.dinb(n28816), .dina(n3216), .dout(n3220));
    jor g0831(.dinb(n28824), .dina(n3220), .dout(n3224));
    jand g0832(.dinb(G222gat), .dina(G307gat), .dout(n3228));
    jnot g0833(.din(n2842), .dout(n3231));
    jand g0834(.dinb(G256gat), .dina(G273gat), .dout(n3235));
    jand g0835(.dinb(n3231), .dina(n32893), .dout(n3239));
    jnot g0836(.din(n3239), .dout(n3242));
    jor g0837(.dinb(n3231), .dina(n32893), .dout(n3246));
    jand g0838(.dinb(n2849), .dina(n3246), .dout(n3250));
    jand g0839(.dinb(n3242), .dina(n3250), .dout(n3254));
    jnot g0840(.din(n3246), .dout(n3257));
    jand g0841(.dinb(n32883), .dina(n3257), .dout(n3261));
    jor g0842(.dinb(n3254), .dina(n3261), .dout(n3265));
    jxor g0843(.dinb(n32895), .dina(n3265), .dout(n3269));
    jxor g0844(.dinb(n3224), .dina(n28798), .dout(n3273));
    jxor g0845(.dinb(n28789), .dina(n3273), .dout(n3277));
    jxor g0846(.dinb(n3203), .dina(n27445), .dout(n3281));
    jxor g0847(.dinb(n27442), .dina(n3281), .dout(n3285));
    jxor g0848(.dinb(n3184), .dina(n26140), .dout(n3289));
    jxor g0849(.dinb(n26137), .dina(n3289), .dout(n3293));
    jxor g0850(.dinb(n3165), .dina(n24859), .dout(n3297));
    jxor g0851(.dinb(n24856), .dina(n3297), .dout(n3301));
    jxor g0852(.dinb(n3146), .dina(n23584), .dout(n3305));
    jxor g0853(.dinb(n23581), .dina(n3305), .dout(n3309));
    jxor g0854(.dinb(n3127), .dina(n22309), .dout(n3313));
    jxor g0855(.dinb(n22306), .dina(n3313), .dout(n3317));
    jxor g0856(.dinb(n3108), .dina(n3317), .dout(n3321));
    jxor g0857(.dinb(n21100), .dina(n3321), .dout(n3325));
    jxor g0858(.dinb(n3089), .dina(n3325), .dout(n3329));
    jxor g0859(.dinb(n19945), .dina(n3329), .dout(n3333));
    jxor g0860(.dinb(n3070), .dina(n18778), .dout(n3337));
    jxor g0861(.dinb(n18775), .dina(n3337), .dout(n3341));
    jxor g0862(.dinb(n3051), .dina(n17587), .dout(n3345));
    jxor g0863(.dinb(n17584), .dina(n3345), .dout(n3349));
    jxor g0864(.dinb(n3032), .dina(n16362), .dout(n3353));
    jxor g0865(.dinb(n15106), .dina(n3353), .dout(n3357));
    jxor g0866(.dinb(n3013), .dina(n14994), .dout(n3361));
    jxor g0867(.dinb(n14992), .dina(n3361), .dout(n3365));
    jxor g0868(.dinb(n2993), .dina(n13005), .dout(n3369));
    jxor g0869(.dinb(n11743), .dina(n3369), .dout(n3373));
    jnot g0870(.din(n3365), .dout(n3376));
    jor g0871(.dinb(n2993), .dina(n3376), .dout(n3380));
    jor g0872(.dinb(n12873), .dina(n3369), .dout(n3384));
    jand g0873(.dinb(n12871), .dina(n3384), .dout(n3388));
    jand g0874(.dinb(G18gat), .dina(G528gat), .dout(n3392));
    jnot g0875(.din(n3357), .dout(n3395));
    jor g0876(.dinb(n3013), .dina(n3395), .dout(n3399));
    jor g0877(.dinb(n14992), .dina(n3361), .dout(n3403));
    jand g0878(.dinb(n14869), .dina(n3403), .dout(n3407));
    jand g0879(.dinb(G35gat), .dina(G511gat), .dout(n3411));
    jand g0880(.dinb(n3032), .dina(n16359), .dout(n3415));
    jnot g0881(.din(n3415), .dout(n3418));
    jnot g0882(.din(n3349), .dout(n3421));
    jxor g0883(.dinb(n3032), .dina(n3421), .dout(n3425));
    jor g0884(.dinb(n16245), .dina(n3425), .dout(n3429));
    jand g0885(.dinb(n3418), .dina(n3429), .dout(n3433));
    jand g0886(.dinb(G52gat), .dina(G494gat), .dout(n3437));
    jnot g0887(.din(n3437), .dout(n3440));
    jand g0888(.dinb(n3051), .dina(n17587), .dout(n3444));
    jand g0889(.dinb(n17584), .dina(n3345), .dout(n3448));
    jor g0890(.dinb(n17482), .dina(n3448), .dout(n3452));
    jand g0891(.dinb(G69gat), .dina(G477gat), .dout(n3456));
    jnot g0892(.din(n3456), .dout(n3459));
    jand g0893(.dinb(n3070), .dina(n18778), .dout(n3463));
    jand g0894(.dinb(n18775), .dina(n3337), .dout(n3467));
    jor g0895(.dinb(n18682), .dina(n3467), .dout(n3471));
    jand g0896(.dinb(G86gat), .dina(G460gat), .dout(n3475));
    jnot g0897(.din(n3475), .dout(n3478));
    jand g0898(.dinb(n3089), .dina(n3325), .dout(n3482));
    jand g0899(.dinb(n19945), .dina(n3329), .dout(n3486));
    jor g0900(.dinb(n19861), .dina(n3486), .dout(n3490));
    jand g0901(.dinb(G103gat), .dina(G443gat), .dout(n3494));
    jnot g0902(.din(n3494), .dout(n3497));
    jand g0903(.dinb(n3108), .dina(n3317), .dout(n3501));
    jand g0904(.dinb(n21100), .dina(n3321), .dout(n3505));
    jor g0905(.dinb(n21022), .dina(n3505), .dout(n3509));
    jand g0906(.dinb(G120gat), .dina(G426gat), .dout(n3513));
    jnot g0907(.din(n3513), .dout(n3516));
    jand g0908(.dinb(n3127), .dina(n22309), .dout(n3520));
    jand g0909(.dinb(n22306), .dina(n3313), .dout(n3524));
    jor g0910(.dinb(n22234), .dina(n3524), .dout(n3528));
    jand g0911(.dinb(G137gat), .dina(G409gat), .dout(n3532));
    jnot g0912(.din(n3532), .dout(n3535));
    jand g0913(.dinb(n3146), .dina(n23584), .dout(n3539));
    jand g0914(.dinb(n23581), .dina(n3305), .dout(n3543));
    jor g0915(.dinb(n23518), .dina(n3543), .dout(n3547));
    jand g0916(.dinb(G154gat), .dina(G392gat), .dout(n3551));
    jnot g0917(.din(n3551), .dout(n3554));
    jand g0918(.dinb(n3165), .dina(n24859), .dout(n3558));
    jand g0919(.dinb(n24856), .dina(n3297), .dout(n3562));
    jor g0920(.dinb(n24802), .dina(n3562), .dout(n3566));
    jand g0921(.dinb(G171gat), .dina(G375gat), .dout(n3570));
    jnot g0922(.din(n3570), .dout(n3573));
    jand g0923(.dinb(n3184), .dina(n26140), .dout(n3577));
    jand g0924(.dinb(n26137), .dina(n3289), .dout(n3581));
    jor g0925(.dinb(n26092), .dina(n3581), .dout(n3585));
    jand g0926(.dinb(G188gat), .dina(G358gat), .dout(n3589));
    jnot g0927(.din(n3589), .dout(n3592));
    jand g0928(.dinb(n3203), .dina(n27445), .dout(n3596));
    jand g0929(.dinb(n27442), .dina(n3281), .dout(n3600));
    jor g0930(.dinb(n27406), .dina(n3600), .dout(n3604));
    jand g0931(.dinb(G205gat), .dina(G341gat), .dout(n3608));
    jnot g0932(.din(n3608), .dout(n3611));
    jand g0933(.dinb(n3224), .dina(n28798), .dout(n3615));
    jand g0934(.dinb(n28789), .dina(n3273), .dout(n3619));
    jor g0935(.dinb(n28762), .dina(n3619), .dout(n3623));
    jand g0936(.dinb(G222gat), .dina(G324gat), .dout(n3627));
    jnot g0937(.din(n3627), .dout(n3630));
    jnot g0938(.din(n3228), .dout(n3633));
    jnot g0939(.din(n3265), .dout(n3636));
    jand g0940(.dinb(n32872), .dina(n3636), .dout(n3640));
    jor g0941(.dinb(n32874), .dina(n3640), .dout(n3644));
    jand g0942(.dinb(G239gat), .dina(G307gat), .dout(n3648));
    jand g0943(.dinb(G256gat), .dina(G290gat), .dout(n3652));
    jnot g0944(.din(n3652), .dout(n3655));
    jor g0945(.dinb(n32850), .dina(n3655), .dout(n3659));
    jxor g0946(.dinb(n32853), .dina(n3659), .dout(n3663));
    jxor g0947(.dinb(n3644), .dina(n32839), .dout(n3667));
    jxor g0948(.dinb(n32824), .dina(n3667), .dout(n3671));
    jxor g0949(.dinb(n3623), .dina(n28759), .dout(n3675));
    jxor g0950(.dinb(n28753), .dina(n3675), .dout(n3679));
    jxor g0951(.dinb(n3604), .dina(n27403), .dout(n3683));
    jxor g0952(.dinb(n27400), .dina(n3683), .dout(n3687));
    jxor g0953(.dinb(n3585), .dina(n26089), .dout(n3691));
    jxor g0954(.dinb(n26086), .dina(n3691), .dout(n3695));
    jxor g0955(.dinb(n3566), .dina(n24799), .dout(n3699));
    jxor g0956(.dinb(n24796), .dina(n3699), .dout(n3703));
    jxor g0957(.dinb(n3547), .dina(n23515), .dout(n3707));
    jxor g0958(.dinb(n23512), .dina(n3707), .dout(n3711));
    jxor g0959(.dinb(n3528), .dina(n22231), .dout(n3715));
    jxor g0960(.dinb(n22228), .dina(n3715), .dout(n3719));
    jxor g0961(.dinb(n3509), .dina(n3719), .dout(n3723));
    jxor g0962(.dinb(n21019), .dina(n3723), .dout(n3727));
    jxor g0963(.dinb(n3490), .dina(n3727), .dout(n3731));
    jxor g0964(.dinb(n19858), .dina(n3731), .dout(n3735));
    jxor g0965(.dinb(n3471), .dina(n18679), .dout(n3739));
    jxor g0966(.dinb(n18676), .dina(n3739), .dout(n3743));
    jxor g0967(.dinb(n3452), .dina(n17479), .dout(n3747));
    jxor g0968(.dinb(n17476), .dina(n3747), .dout(n3751));
    jxor g0969(.dinb(n3433), .dina(n16242), .dout(n3755));
    jxor g0970(.dinb(n16240), .dina(n3755), .dout(n3759));
    jnot g0971(.din(n3759), .dout(n3762));
    jxor g0972(.dinb(n3407), .dina(n3762), .dout(n3766));
    jxor g0973(.dinb(n14863), .dina(n3766), .dout(n3770));
    jxor g0974(.dinb(n3388), .dina(n12868), .dout(n3774));
    jand g0975(.dinb(n3388), .dina(n12868), .dout(n3778));
    jor g0976(.dinb(n3407), .dina(n3762), .dout(n3782));
    jxor g0977(.dinb(n3407), .dina(n14865), .dout(n3786));
    jor g0978(.dinb(n14863), .dina(n3786), .dout(n3790));
    jand g0979(.dinb(n14731), .dina(n3790), .dout(n3794));
    jand g0980(.dinb(G35gat), .dina(G528gat), .dout(n3798));
    jnot g0981(.din(n3751), .dout(n3801));
    jor g0982(.dinb(n3433), .dina(n3801), .dout(n3805));
    jor g0983(.dinb(n16240), .dina(n3755), .dout(n3809));
    jand g0984(.dinb(n16117), .dina(n3809), .dout(n3813));
    jand g0985(.dinb(G52gat), .dina(G511gat), .dout(n3817));
    jand g0986(.dinb(n3452), .dina(n17479), .dout(n3821));
    jand g0987(.dinb(n17476), .dina(n3747), .dout(n3825));
    jor g0988(.dinb(n17365), .dina(n3825), .dout(n3829));
    jand g0989(.dinb(G69gat), .dina(G494gat), .dout(n3833));
    jnot g0990(.din(n3833), .dout(n3836));
    jand g0991(.dinb(n3471), .dina(n18679), .dout(n3840));
    jand g0992(.dinb(n18676), .dina(n3739), .dout(n3844));
    jor g0993(.dinb(n18574), .dina(n3844), .dout(n3848));
    jand g0994(.dinb(G86gat), .dina(G477gat), .dout(n3852));
    jnot g0995(.din(n3852), .dout(n3855));
    jand g0996(.dinb(n3490), .dina(n3727), .dout(n3859));
    jand g0997(.dinb(n19858), .dina(n3731), .dout(n3863));
    jor g0998(.dinb(n19765), .dina(n3863), .dout(n3867));
    jand g0999(.dinb(G103gat), .dina(G460gat), .dout(n3871));
    jnot g1000(.din(n3871), .dout(n3874));
    jand g1001(.dinb(n3509), .dina(n3719), .dout(n3878));
    jand g1002(.dinb(n21019), .dina(n3723), .dout(n3882));
    jor g1003(.dinb(n20932), .dina(n3882), .dout(n3886));
    jand g1004(.dinb(G120gat), .dina(G443gat), .dout(n3890));
    jnot g1005(.din(n3890), .dout(n3893));
    jand g1006(.dinb(n3528), .dina(n22231), .dout(n3897));
    jand g1007(.dinb(n22228), .dina(n3715), .dout(n3901));
    jor g1008(.dinb(n22147), .dina(n3901), .dout(n3905));
    jand g1009(.dinb(G137gat), .dina(G426gat), .dout(n3909));
    jnot g1010(.din(n3909), .dout(n3912));
    jand g1011(.dinb(n3547), .dina(n23515), .dout(n3916));
    jand g1012(.dinb(n23512), .dina(n3707), .dout(n3920));
    jor g1013(.dinb(n23440), .dina(n3920), .dout(n3924));
    jand g1014(.dinb(G154gat), .dina(G409gat), .dout(n3928));
    jnot g1015(.din(n3928), .dout(n3931));
    jand g1016(.dinb(n3566), .dina(n24799), .dout(n3935));
    jand g1017(.dinb(n24796), .dina(n3699), .dout(n3939));
    jor g1018(.dinb(n24733), .dina(n3939), .dout(n3943));
    jand g1019(.dinb(G171gat), .dina(G392gat), .dout(n3947));
    jnot g1020(.din(n3947), .dout(n3950));
    jand g1021(.dinb(n3585), .dina(n26089), .dout(n3954));
    jand g1022(.dinb(n26086), .dina(n3691), .dout(n3958));
    jor g1023(.dinb(n26032), .dina(n3958), .dout(n3962));
    jand g1024(.dinb(G188gat), .dina(G375gat), .dout(n3966));
    jnot g1025(.din(n3966), .dout(n3969));
    jand g1026(.dinb(n3604), .dina(n27403), .dout(n3973));
    jand g1027(.dinb(n27400), .dina(n3683), .dout(n3977));
    jor g1028(.dinb(n27355), .dina(n3977), .dout(n3981));
    jand g1029(.dinb(G205gat), .dina(G358gat), .dout(n3985));
    jnot g1030(.din(n3985), .dout(n3988));
    jand g1031(.dinb(n3623), .dina(n28759), .dout(n3992));
    jand g1032(.dinb(n28753), .dina(n3675), .dout(n3996));
    jor g1033(.dinb(n28717), .dina(n3996), .dout(n4000));
    jand g1034(.dinb(G222gat), .dina(G341gat), .dout(n4004));
    jnot g1035(.din(n4004), .dout(n4007));
    jand g1036(.dinb(n3644), .dina(n32839), .dout(n4011));
    jand g1037(.dinb(n32824), .dina(n3667), .dout(n4015));
    jor g1038(.dinb(n32800), .dina(n4015), .dout(n4019));
    jand g1039(.dinb(G239gat), .dina(G324gat), .dout(n4023));
    jand g1040(.dinb(G256gat), .dina(G307gat), .dout(n4027));
    jnot g1041(.din(n3648), .dout(n4030));
    jnot g1042(.din(n3659), .dout(n4033));
    jand g1043(.dinb(n32746), .dina(n4033), .dout(n4037));
    jor g1044(.dinb(n32841), .dina(n4037), .dout(n4041));
    jnot g1045(.din(n4041), .dout(n4044));
    jor g1046(.dinb(n32740), .dina(n4044), .dout(n4048));
    jand g1047(.dinb(n32748), .dina(n4044), .dout(n4052));
    jnot g1048(.din(n4052), .dout(n4055));
    jand g1049(.dinb(n32722), .dina(n4055), .dout(n4059));
    jnot g1050(.din(n4059), .dout(n4062));
    jxor g1051(.dinb(n32797), .dina(n4062), .dout(n4066));
    jxor g1052(.dinb(n4019), .dina(n4066), .dout(n4070));
    jxor g1053(.dinb(n32710), .dina(n4070), .dout(n4074));
    jxor g1054(.dinb(n4000), .dina(n28714), .dout(n4078));
    jxor g1055(.dinb(n28708), .dina(n4078), .dout(n4082));
    jxor g1056(.dinb(n3981), .dina(n27352), .dout(n4086));
    jxor g1057(.dinb(n27349), .dina(n4086), .dout(n4090));
    jxor g1058(.dinb(n3962), .dina(n26029), .dout(n4094));
    jxor g1059(.dinb(n26026), .dina(n4094), .dout(n4098));
    jxor g1060(.dinb(n3943), .dina(n24730), .dout(n4102));
    jxor g1061(.dinb(n24727), .dina(n4102), .dout(n4106));
    jxor g1062(.dinb(n3924), .dina(n23437), .dout(n4110));
    jxor g1063(.dinb(n23434), .dina(n4110), .dout(n4114));
    jxor g1064(.dinb(n3905), .dina(n22144), .dout(n4118));
    jxor g1065(.dinb(n22141), .dina(n4118), .dout(n4122));
    jxor g1066(.dinb(n3886), .dina(n4122), .dout(n4126));
    jxor g1067(.dinb(n20929), .dina(n4126), .dout(n4130));
    jxor g1068(.dinb(n3867), .dina(n4130), .dout(n4134));
    jxor g1069(.dinb(n19762), .dina(n4134), .dout(n4138));
    jxor g1070(.dinb(n3848), .dina(n18571), .dout(n4142));
    jxor g1071(.dinb(n18568), .dina(n4142), .dout(n4146));
    jxor g1072(.dinb(n3829), .dina(n17362), .dout(n4150));
    jnot g1073(.din(n4150), .dout(n4153));
    jxor g1074(.dinb(n17359), .dina(n4153), .dout(n4157));
    jxor g1075(.dinb(n3813), .dina(n4157), .dout(n4161));
    jxor g1076(.dinb(n16111), .dina(n4161), .dout(n4165));
    jxor g1077(.dinb(n3794), .dina(n14727), .dout(n4169));
    jnot g1078(.din(n4169), .dout(n4172));
    jxor g1079(.dinb(n12864), .dina(n4172), .dout(n4176));
    jnot g1080(.din(n4165), .dout(n4179));
    jor g1081(.dinb(n3794), .dina(n4179), .dout(n4183));
    jor g1082(.dinb(n3778), .dina(n4169), .dout(n4187));
    jand g1083(.dinb(n12862), .dina(n4187), .dout(n4191));
    jnot g1084(.din(n4157), .dout(n4194));
    jor g1085(.dinb(n16113), .dina(n4194), .dout(n4198));
    jor g1086(.dinb(n16111), .dina(n4161), .dout(n4202));
    jand g1087(.dinb(n4198), .dina(n4202), .dout(n4206));
    jand g1088(.dinb(G52gat), .dina(G528gat), .dout(n4210));
    jand g1089(.dinb(n3829), .dina(n17362), .dout(n4214));
    jnot g1090(.din(n4214), .dout(n4217));
    jor g1091(.dinb(n17359), .dina(n4153), .dout(n4221));
    jand g1092(.dinb(n17233), .dina(n4221), .dout(n4225));
    jand g1093(.dinb(G69gat), .dina(G511gat), .dout(n4229));
    jnot g1094(.din(n4229), .dout(n4232));
    jand g1095(.dinb(n3848), .dina(n18571), .dout(n4236));
    jand g1096(.dinb(n18568), .dina(n4142), .dout(n4240));
    jor g1097(.dinb(n18457), .dina(n4240), .dout(n4244));
    jand g1098(.dinb(G86gat), .dina(G494gat), .dout(n4248));
    jnot g1099(.din(n4248), .dout(n4251));
    jand g1100(.dinb(n3867), .dina(n4130), .dout(n4255));
    jand g1101(.dinb(n19762), .dina(n4134), .dout(n4259));
    jor g1102(.dinb(n19660), .dina(n4259), .dout(n4263));
    jand g1103(.dinb(G103gat), .dina(G477gat), .dout(n4267));
    jnot g1104(.din(n4267), .dout(n4270));
    jand g1105(.dinb(n3886), .dina(n4122), .dout(n4274));
    jand g1106(.dinb(n20929), .dina(n4126), .dout(n4278));
    jor g1107(.dinb(n20833), .dina(n4278), .dout(n4282));
    jand g1108(.dinb(G120gat), .dina(G460gat), .dout(n4286));
    jnot g1109(.din(n4286), .dout(n4289));
    jand g1110(.dinb(n3905), .dina(n22144), .dout(n4293));
    jand g1111(.dinb(n22141), .dina(n4118), .dout(n4297));
    jor g1112(.dinb(n22051), .dina(n4297), .dout(n4301));
    jand g1113(.dinb(G137gat), .dina(G443gat), .dout(n4305));
    jnot g1114(.din(n4305), .dout(n4308));
    jand g1115(.dinb(n3924), .dina(n23437), .dout(n4312));
    jand g1116(.dinb(n23434), .dina(n4110), .dout(n4316));
    jor g1117(.dinb(n23353), .dina(n4316), .dout(n4320));
    jand g1118(.dinb(G154gat), .dina(G426gat), .dout(n4324));
    jnot g1119(.din(n4324), .dout(n4327));
    jand g1120(.dinb(n3943), .dina(n24730), .dout(n4331));
    jand g1121(.dinb(n24727), .dina(n4102), .dout(n4335));
    jor g1122(.dinb(n24655), .dina(n4335), .dout(n4339));
    jand g1123(.dinb(G171gat), .dina(G409gat), .dout(n4343));
    jnot g1124(.din(n4343), .dout(n4346));
    jand g1125(.dinb(n3962), .dina(n26029), .dout(n4350));
    jand g1126(.dinb(n26026), .dina(n4094), .dout(n4354));
    jor g1127(.dinb(n25963), .dina(n4354), .dout(n4358));
    jand g1128(.dinb(G188gat), .dina(G392gat), .dout(n4362));
    jnot g1129(.din(n4362), .dout(n4365));
    jand g1130(.dinb(n3981), .dina(n27352), .dout(n4369));
    jand g1131(.dinb(n27349), .dina(n4086), .dout(n4373));
    jor g1132(.dinb(n27295), .dina(n4373), .dout(n4377));
    jand g1133(.dinb(G205gat), .dina(G375gat), .dout(n4381));
    jnot g1134(.din(n4381), .dout(n4384));
    jand g1135(.dinb(n4000), .dina(n28714), .dout(n4388));
    jand g1136(.dinb(n28708), .dina(n4078), .dout(n4392));
    jor g1137(.dinb(n28663), .dina(n4392), .dout(n4396));
    jand g1138(.dinb(G222gat), .dina(G358gat), .dout(n4400));
    jnot g1139(.din(n4400), .dout(n4403));
    jand g1140(.dinb(n4019), .dina(n4066), .dout(n4407));
    jand g1141(.dinb(n32710), .dina(n4070), .dout(n4411));
    jor g1142(.dinb(n32677), .dina(n4411), .dout(n4415));
    jand g1143(.dinb(G239gat), .dina(G341gat), .dout(n4419));
    jand g1144(.dinb(G256gat), .dina(G324gat), .dout(n4423));
    jor g1145(.dinb(n32797), .dina(n4062), .dout(n4427));
    jand g1146(.dinb(n32712), .dina(n4427), .dout(n4431));
    jxor g1147(.dinb(n32629), .dina(n4431), .dout(n4435));
    jnot g1148(.din(n4435), .dout(n4438));
    jxor g1149(.dinb(n32671), .dina(n4438), .dout(n4442));
    jxor g1150(.dinb(n32674), .dina(n4442), .dout(n4446));
    jxor g1151(.dinb(n32593), .dina(n4446), .dout(n4450));
    jxor g1152(.dinb(n4396), .dina(n28660), .dout(n4454));
    jxor g1153(.dinb(n28657), .dina(n4454), .dout(n4458));
    jxor g1154(.dinb(n4377), .dina(n27292), .dout(n4462));
    jxor g1155(.dinb(n27289), .dina(n4462), .dout(n4466));
    jxor g1156(.dinb(n4358), .dina(n25960), .dout(n4470));
    jxor g1157(.dinb(n25957), .dina(n4470), .dout(n4474));
    jxor g1158(.dinb(n4339), .dina(n24652), .dout(n4478));
    jxor g1159(.dinb(n24649), .dina(n4478), .dout(n4482));
    jxor g1160(.dinb(n4320), .dina(n23350), .dout(n4486));
    jxor g1161(.dinb(n23347), .dina(n4486), .dout(n4490));
    jxor g1162(.dinb(n4301), .dina(n22048), .dout(n4494));
    jxor g1163(.dinb(n22045), .dina(n4494), .dout(n4498));
    jxor g1164(.dinb(n4282), .dina(n4498), .dout(n4502));
    jxor g1165(.dinb(n20830), .dina(n4502), .dout(n4506));
    jxor g1166(.dinb(n4263), .dina(n4506), .dout(n4510));
    jxor g1167(.dinb(n19657), .dina(n4510), .dout(n4514));
    jxor g1168(.dinb(n4244), .dina(n18454), .dout(n4518));
    jxor g1169(.dinb(n18451), .dina(n4518), .dout(n4522));
    jnot g1170(.din(n4522), .dout(n4525));
    jxor g1171(.dinb(n4225), .dina(n17230), .dout(n4529));
    jnot g1172(.din(n4529), .dout(n4532));
    jxor g1173(.dinb(n17227), .dina(n4532), .dout(n4536));
    jxor g1174(.dinb(n15979), .dina(n4536), .dout(n4540));
    jnot g1175(.din(n4540), .dout(n4543));
    jxor g1176(.dinb(n4191), .dina(n4543), .dout(n4547));
    jnot g1177(.din(n4536), .dout(n4550));
    jor g1178(.dinb(n15975), .dina(n4550), .dout(n4554));
    jor g1179(.dinb(n4191), .dina(n12858), .dout(n4558));
    jand g1180(.dinb(n12856), .dina(n4558), .dout(n4562));
    jor g1181(.dinb(n4225), .dina(n17230), .dout(n4566));
    jor g1182(.dinb(n17227), .dina(n4532), .dout(n4570));
    jand g1183(.dinb(n17089), .dina(n4570), .dout(n4574));
    jand g1184(.dinb(G69gat), .dina(G528gat), .dout(n4578));
    jand g1185(.dinb(n4244), .dina(n18454), .dout(n4582));
    jand g1186(.dinb(n18451), .dina(n4518), .dout(n4586));
    jor g1187(.dinb(n18331), .dina(n4586), .dout(n4590));
    jand g1188(.dinb(G86gat), .dina(G511gat), .dout(n4594));
    jnot g1189(.din(n4594), .dout(n4597));
    jand g1190(.dinb(n4263), .dina(n4506), .dout(n4601));
    jand g1191(.dinb(n19657), .dina(n4510), .dout(n4605));
    jor g1192(.dinb(n19546), .dina(n4605), .dout(n4609));
    jand g1193(.dinb(G103gat), .dina(G494gat), .dout(n4613));
    jnot g1194(.din(n4613), .dout(n4616));
    jand g1195(.dinb(n4282), .dina(n4498), .dout(n4620));
    jand g1196(.dinb(n20830), .dina(n4502), .dout(n4624));
    jor g1197(.dinb(n20725), .dina(n4624), .dout(n4628));
    jand g1198(.dinb(G120gat), .dina(G477gat), .dout(n4632));
    jnot g1199(.din(n4632), .dout(n4635));
    jand g1200(.dinb(n4301), .dina(n22048), .dout(n4639));
    jand g1201(.dinb(n22045), .dina(n4494), .dout(n4643));
    jor g1202(.dinb(n21946), .dina(n4643), .dout(n4647));
    jand g1203(.dinb(G137gat), .dina(G460gat), .dout(n4651));
    jnot g1204(.din(n4651), .dout(n4654));
    jand g1205(.dinb(n4320), .dina(n23350), .dout(n4658));
    jand g1206(.dinb(n23347), .dina(n4486), .dout(n4662));
    jor g1207(.dinb(n23257), .dina(n4662), .dout(n4666));
    jand g1208(.dinb(G154gat), .dina(G443gat), .dout(n4670));
    jnot g1209(.din(n4670), .dout(n4673));
    jand g1210(.dinb(n4339), .dina(n24652), .dout(n4677));
    jand g1211(.dinb(n24649), .dina(n4478), .dout(n4681));
    jor g1212(.dinb(n24568), .dina(n4681), .dout(n4685));
    jand g1213(.dinb(G171gat), .dina(G426gat), .dout(n4689));
    jnot g1214(.din(n4689), .dout(n4692));
    jand g1215(.dinb(n4358), .dina(n25960), .dout(n4696));
    jand g1216(.dinb(n25957), .dina(n4470), .dout(n4700));
    jor g1217(.dinb(n25885), .dina(n4700), .dout(n4704));
    jand g1218(.dinb(G188gat), .dina(G409gat), .dout(n4708));
    jnot g1219(.din(n4708), .dout(n4711));
    jand g1220(.dinb(n4377), .dina(n27292), .dout(n4715));
    jand g1221(.dinb(n27289), .dina(n4462), .dout(n4719));
    jor g1222(.dinb(n27226), .dina(n4719), .dout(n4723));
    jand g1223(.dinb(G205gat), .dina(G392gat), .dout(n4727));
    jnot g1224(.din(n4727), .dout(n4730));
    jand g1225(.dinb(n4396), .dina(n28660), .dout(n4734));
    jand g1226(.dinb(n28657), .dina(n4454), .dout(n4738));
    jor g1227(.dinb(n28603), .dina(n4738), .dout(n4742));
    jand g1228(.dinb(G222gat), .dina(G375gat), .dout(n4746));
    jnot g1229(.din(n4746), .dout(n4749));
    jand g1230(.dinb(n32674), .dina(n4442), .dout(n4753));
    jand g1231(.dinb(n32593), .dina(n4446), .dout(n4757));
    jor g1232(.dinb(n32548), .dina(n4757), .dout(n4761));
    jand g1233(.dinb(G239gat), .dina(G358gat), .dout(n4765));
    jand g1234(.dinb(G256gat), .dina(G341gat), .dout(n4769));
    jor g1235(.dinb(n32629), .dina(n4431), .dout(n4773));
    jor g1236(.dinb(n32671), .dina(n4438), .dout(n4777));
    jand g1237(.dinb(n32440), .dina(n4777), .dout(n4781));
    jxor g1238(.dinb(n32488), .dina(n4781), .dout(n4785));
    jnot g1239(.din(n4785), .dout(n4788));
    jxor g1240(.dinb(n32542), .dina(n4788), .dout(n4792));
    jxor g1241(.dinb(n32545), .dina(n4792), .dout(n4796));
    jxor g1242(.dinb(n32434), .dina(n4796), .dout(n4800));
    jxor g1243(.dinb(n4742), .dina(n4800), .dout(n4804));
    jxor g1244(.dinb(n28600), .dina(n4804), .dout(n4808));
    jxor g1245(.dinb(n4723), .dina(n27223), .dout(n4812));
    jxor g1246(.dinb(n27220), .dina(n4812), .dout(n4816));
    jxor g1247(.dinb(n4704), .dina(n25882), .dout(n4820));
    jxor g1248(.dinb(n25879), .dina(n4820), .dout(n4824));
    jxor g1249(.dinb(n4685), .dina(n24565), .dout(n4828));
    jxor g1250(.dinb(n24562), .dina(n4828), .dout(n4832));
    jxor g1251(.dinb(n4666), .dina(n23254), .dout(n4836));
    jxor g1252(.dinb(n23251), .dina(n4836), .dout(n4840));
    jxor g1253(.dinb(n4647), .dina(n21943), .dout(n4844));
    jxor g1254(.dinb(n21940), .dina(n4844), .dout(n4848));
    jxor g1255(.dinb(n4628), .dina(n4848), .dout(n4852));
    jxor g1256(.dinb(n20722), .dina(n4852), .dout(n4856));
    jxor g1257(.dinb(n4609), .dina(n4856), .dout(n4860));
    jxor g1258(.dinb(n19543), .dina(n4860), .dout(n4864));
    jxor g1259(.dinb(n4590), .dina(n18327), .dout(n4868));
    jnot g1260(.din(n4868), .dout(n4871));
    jxor g1261(.dinb(n18322), .dina(n4871), .dout(n4875));
    jxor g1262(.dinb(n4574), .dina(n17079), .dout(n4879));
    jnot g1263(.din(n4879), .dout(n4882));
    jxor g1264(.dinb(n4562), .dina(n11746), .dout(n4886));
    jnot g1265(.din(n4875), .dout(n4889));
    jor g1266(.dinb(n4574), .dina(n17077), .dout(n4893));
    jor g1267(.dinb(n4562), .dina(n12849), .dout(n4897));
    jand g1268(.dinb(n12847), .dina(n4897), .dout(n4901));
    jnot g1269(.din(n4590), .dout(n4904));
    jnot g1270(.din(n4864), .dout(n4907));
    jor g1271(.dinb(n4904), .dina(n18325), .dout(n4911));
    jor g1272(.dinb(n18322), .dina(n4871), .dout(n4915));
    jand g1273(.dinb(n18187), .dina(n4915), .dout(n4919));
    jand g1274(.dinb(G86gat), .dina(G528gat), .dout(n4923));
    jand g1275(.dinb(n4609), .dina(n4856), .dout(n4927));
    jand g1276(.dinb(n19543), .dina(n4860), .dout(n4931));
    jor g1277(.dinb(n19423), .dina(n4931), .dout(n4935));
    jand g1278(.dinb(G103gat), .dina(G511gat), .dout(n4939));
    jnot g1279(.din(n4939), .dout(n4942));
    jand g1280(.dinb(n4628), .dina(n4848), .dout(n4946));
    jand g1281(.dinb(n20722), .dina(n4852), .dout(n4950));
    jor g1282(.dinb(n20608), .dina(n4950), .dout(n4954));
    jand g1283(.dinb(G120gat), .dina(G494gat), .dout(n4958));
    jnot g1284(.din(n4958), .dout(n4961));
    jand g1285(.dinb(n4647), .dina(n21943), .dout(n4965));
    jand g1286(.dinb(n21940), .dina(n4844), .dout(n4969));
    jor g1287(.dinb(n21832), .dina(n4969), .dout(n4973));
    jand g1288(.dinb(G137gat), .dina(G477gat), .dout(n4977));
    jnot g1289(.din(n4977), .dout(n4980));
    jand g1290(.dinb(n4666), .dina(n23254), .dout(n4984));
    jand g1291(.dinb(n23251), .dina(n4836), .dout(n4988));
    jor g1292(.dinb(n23152), .dina(n4988), .dout(n4992));
    jand g1293(.dinb(G154gat), .dina(G460gat), .dout(n4996));
    jnot g1294(.din(n4996), .dout(n4999));
    jand g1295(.dinb(n4685), .dina(n24565), .dout(n5003));
    jand g1296(.dinb(n24562), .dina(n4828), .dout(n5007));
    jor g1297(.dinb(n24472), .dina(n5007), .dout(n5011));
    jand g1298(.dinb(G171gat), .dina(G443gat), .dout(n5015));
    jnot g1299(.din(n5015), .dout(n5018));
    jand g1300(.dinb(n4704), .dina(n25882), .dout(n5022));
    jand g1301(.dinb(n25879), .dina(n4820), .dout(n5026));
    jor g1302(.dinb(n25798), .dina(n5026), .dout(n5030));
    jand g1303(.dinb(G188gat), .dina(G426gat), .dout(n5034));
    jnot g1304(.din(n5034), .dout(n5037));
    jand g1305(.dinb(n4723), .dina(n27223), .dout(n5041));
    jand g1306(.dinb(n27220), .dina(n4812), .dout(n5045));
    jor g1307(.dinb(n27148), .dina(n5045), .dout(n5049));
    jand g1308(.dinb(G205gat), .dina(G409gat), .dout(n5053));
    jnot g1309(.din(n5053), .dout(n5056));
    jand g1310(.dinb(n4742), .dina(n4800), .dout(n5060));
    jand g1311(.dinb(n28600), .dina(n4804), .dout(n5064));
    jor g1312(.dinb(n28537), .dina(n5064), .dout(n5068));
    jand g1313(.dinb(G222gat), .dina(G392gat), .dout(n5072));
    jnot g1314(.din(n5072), .dout(n5075));
    jand g1315(.dinb(n32545), .dina(n4792), .dout(n5079));
    jand g1316(.dinb(n32434), .dina(n4796), .dout(n5083));
    jor g1317(.dinb(n32377), .dina(n5083), .dout(n5087));
    jand g1318(.dinb(G239gat), .dina(G375gat), .dout(n5091));
    jand g1319(.dinb(G256gat), .dina(G358gat), .dout(n5095));
    jor g1320(.dinb(n32488), .dina(n4781), .dout(n5099));
    jor g1321(.dinb(n32542), .dina(n4788), .dout(n5103));
    jand g1322(.dinb(n32245), .dina(n5103), .dout(n5107));
    jxor g1323(.dinb(n32305), .dina(n5107), .dout(n5111));
    jnot g1324(.din(n5111), .dout(n5114));
    jxor g1325(.dinb(n32371), .dina(n5114), .dout(n5118));
    jxor g1326(.dinb(n32374), .dina(n5118), .dout(n5122));
    jxor g1327(.dinb(n32239), .dina(n5122), .dout(n5126));
    jxor g1328(.dinb(n28534), .dina(n5126), .dout(n5130));
    jxor g1329(.dinb(n28531), .dina(n5130), .dout(n5134));
    jxor g1330(.dinb(n5049), .dina(n5134), .dout(n5138));
    jxor g1331(.dinb(n27145), .dina(n5138), .dout(n5142));
    jxor g1332(.dinb(n5030), .dina(n25795), .dout(n5146));
    jxor g1333(.dinb(n25792), .dina(n5146), .dout(n5150));
    jxor g1334(.dinb(n5011), .dina(n24469), .dout(n5154));
    jxor g1335(.dinb(n24466), .dina(n5154), .dout(n5158));
    jxor g1336(.dinb(n4992), .dina(n23149), .dout(n5162));
    jxor g1337(.dinb(n23146), .dina(n5162), .dout(n5166));
    jxor g1338(.dinb(n4973), .dina(n21829), .dout(n5170));
    jxor g1339(.dinb(n21826), .dina(n5170), .dout(n5174));
    jxor g1340(.dinb(n4954), .dina(n5174), .dout(n5178));
    jxor g1341(.dinb(n20605), .dina(n5178), .dout(n5182));
    jxor g1342(.dinb(n4935), .dina(n5182), .dout(n5186));
    jnot g1343(.din(n5186), .dout(n5189));
    jxor g1344(.dinb(n19420), .dina(n5189), .dout(n5193));
    jnot g1345(.din(n5193), .dout(n5196));
    jxor g1346(.dinb(n4919), .dina(n5196), .dout(n5200));
    jxor g1347(.dinb(n4901), .dina(n12825), .dout(n5204));
    jor g1348(.dinb(n4919), .dina(n5196), .dout(n5208));
    jnot g1349(.din(n5200), .dout(n5211));
    jor g1350(.dinb(n4901), .dina(n12823), .dout(n5215));
    jand g1351(.dinb(n12811), .dina(n5215), .dout(n5219));
    jnot g1352(.din(n4935), .dout(n5222));
    jnot g1353(.din(n5182), .dout(n5225));
    jor g1354(.dinb(n5222), .dina(n5225), .dout(n5229));
    jor g1355(.dinb(n19420), .dina(n5189), .dout(n5233));
    jand g1356(.dinb(n19285), .dina(n5233), .dout(n5237));
    jand g1357(.dinb(G103gat), .dina(G528gat), .dout(n5241));
    jand g1358(.dinb(n4954), .dina(n5174), .dout(n5245));
    jand g1359(.dinb(n20605), .dina(n5178), .dout(n5249));
    jor g1360(.dinb(n20482), .dina(n5249), .dout(n5253));
    jand g1361(.dinb(G120gat), .dina(G511gat), .dout(n5257));
    jnot g1362(.din(n5257), .dout(n5260));
    jand g1363(.dinb(n4973), .dina(n21829), .dout(n5264));
    jand g1364(.dinb(n21826), .dina(n5170), .dout(n5268));
    jor g1365(.dinb(n21709), .dina(n5268), .dout(n5272));
    jand g1366(.dinb(G137gat), .dina(G494gat), .dout(n5276));
    jnot g1367(.din(n5276), .dout(n5279));
    jand g1368(.dinb(n4992), .dina(n23149), .dout(n5283));
    jand g1369(.dinb(n23146), .dina(n5162), .dout(n5287));
    jor g1370(.dinb(n23038), .dina(n5287), .dout(n5291));
    jand g1371(.dinb(G154gat), .dina(G477gat), .dout(n5295));
    jnot g1372(.din(n5295), .dout(n5298));
    jand g1373(.dinb(n5011), .dina(n24469), .dout(n5302));
    jand g1374(.dinb(n24466), .dina(n5154), .dout(n5306));
    jor g1375(.dinb(n24367), .dina(n5306), .dout(n5310));
    jand g1376(.dinb(G171gat), .dina(G460gat), .dout(n5314));
    jnot g1377(.din(n5314), .dout(n5317));
    jand g1378(.dinb(n5030), .dina(n25795), .dout(n5321));
    jand g1379(.dinb(n25792), .dina(n5146), .dout(n5325));
    jor g1380(.dinb(n25702), .dina(n5325), .dout(n5329));
    jand g1381(.dinb(G188gat), .dina(G443gat), .dout(n5333));
    jnot g1382(.din(n5333), .dout(n5336));
    jand g1383(.dinb(n5049), .dina(n5134), .dout(n5340));
    jand g1384(.dinb(n27145), .dina(n5138), .dout(n5344));
    jor g1385(.dinb(n27064), .dina(n5344), .dout(n5348));
    jand g1386(.dinb(G205gat), .dina(G426gat), .dout(n5352));
    jnot g1387(.din(n5352), .dout(n5355));
    jand g1388(.dinb(n28534), .dina(n5126), .dout(n5359));
    jand g1389(.dinb(n28531), .dina(n5130), .dout(n5363));
    jor g1390(.dinb(n28456), .dina(n5363), .dout(n5367));
    jand g1391(.dinb(G222gat), .dina(G409gat), .dout(n5371));
    jnot g1392(.din(n5371), .dout(n5374));
    jand g1393(.dinb(n32374), .dina(n5118), .dout(n5378));
    jand g1394(.dinb(n32239), .dina(n5122), .dout(n5382));
    jor g1395(.dinb(n32170), .dina(n5382), .dout(n5386));
    jand g1396(.dinb(G239gat), .dina(G392gat), .dout(n5390));
    jand g1397(.dinb(G256gat), .dina(G375gat), .dout(n5394));
    jor g1398(.dinb(n32305), .dina(n5107), .dout(n5398));
    jor g1399(.dinb(n32371), .dina(n5114), .dout(n5402));
    jand g1400(.dinb(n32014), .dina(n5402), .dout(n5406));
    jxor g1401(.dinb(n32086), .dina(n5406), .dout(n5410));
    jnot g1402(.din(n5410), .dout(n5413));
    jxor g1403(.dinb(n32164), .dina(n5413), .dout(n5417));
    jxor g1404(.dinb(n32167), .dina(n5417), .dout(n5421));
    jxor g1405(.dinb(n32008), .dina(n5421), .dout(n5425));
    jxor g1406(.dinb(n28453), .dina(n5425), .dout(n5429));
    jxor g1407(.dinb(n28450), .dina(n5429), .dout(n5433));
    jxor g1408(.dinb(n27061), .dina(n5433), .dout(n5437));
    jxor g1409(.dinb(n27058), .dina(n5437), .dout(n5441));
    jxor g1410(.dinb(n5329), .dina(n5441), .dout(n5445));
    jxor g1411(.dinb(n25699), .dina(n5445), .dout(n5449));
    jxor g1412(.dinb(n5310), .dina(n24364), .dout(n5453));
    jxor g1413(.dinb(n24361), .dina(n5453), .dout(n5457));
    jxor g1414(.dinb(n5291), .dina(n23035), .dout(n5461));
    jxor g1415(.dinb(n23032), .dina(n5461), .dout(n5465));
    jxor g1416(.dinb(n5272), .dina(n21706), .dout(n5469));
    jxor g1417(.dinb(n21703), .dina(n5469), .dout(n5473));
    jxor g1418(.dinb(n5253), .dina(n5473), .dout(n5477));
    jnot g1419(.din(n5477), .dout(n5480));
    jxor g1420(.dinb(n20479), .dina(n5480), .dout(n5484));
    jnot g1421(.din(n5484), .dout(n5487));
    jxor g1422(.dinb(n19282), .dina(n5487), .dout(n5491));
    jxor g1423(.dinb(n5219), .dina(n12777), .dout(n5495));
    jor g1424(.dinb(n19282), .dina(n5487), .dout(n5499));
    jnot g1425(.din(n5491), .dout(n5502));
    jor g1426(.dinb(n5219), .dina(n12775), .dout(n5506));
    jand g1427(.dinb(n12760), .dina(n5506), .dout(n5510));
    jnot g1428(.din(n5253), .dout(n5513));
    jnot g1429(.din(n5473), .dout(n5516));
    jor g1430(.dinb(n5513), .dina(n5516), .dout(n5520));
    jor g1431(.dinb(n20479), .dina(n5480), .dout(n5524));
    jand g1432(.dinb(n20341), .dina(n5524), .dout(n5528));
    jand g1433(.dinb(G120gat), .dina(G528gat), .dout(n5532));
    jand g1434(.dinb(n5272), .dina(n21706), .dout(n5536));
    jand g1435(.dinb(n21703), .dina(n5469), .dout(n5540));
    jor g1436(.dinb(n21577), .dina(n5540), .dout(n5544));
    jand g1437(.dinb(G137gat), .dina(G511gat), .dout(n5548));
    jnot g1438(.din(n5548), .dout(n5551));
    jand g1439(.dinb(n5291), .dina(n23035), .dout(n5555));
    jand g1440(.dinb(n23032), .dina(n5461), .dout(n5559));
    jor g1441(.dinb(n22915), .dina(n5559), .dout(n5563));
    jand g1442(.dinb(G154gat), .dina(G494gat), .dout(n5567));
    jnot g1443(.din(n5567), .dout(n5570));
    jand g1444(.dinb(n5310), .dina(n24364), .dout(n5574));
    jand g1445(.dinb(n24361), .dina(n5453), .dout(n5578));
    jor g1446(.dinb(n24253), .dina(n5578), .dout(n5582));
    jand g1447(.dinb(G171gat), .dina(G477gat), .dout(n5586));
    jnot g1448(.din(n5586), .dout(n5589));
    jand g1449(.dinb(n5329), .dina(n5441), .dout(n5593));
    jand g1450(.dinb(n25699), .dina(n5445), .dout(n5597));
    jor g1451(.dinb(n25600), .dina(n5597), .dout(n5601));
    jand g1452(.dinb(G188gat), .dina(G460gat), .dout(n5605));
    jnot g1453(.din(n5605), .dout(n5608));
    jand g1454(.dinb(n27061), .dina(n5433), .dout(n5612));
    jand g1455(.dinb(n27058), .dina(n5437), .dout(n5616));
    jor g1456(.dinb(n26965), .dina(n5616), .dout(n5620));
    jand g1457(.dinb(G205gat), .dina(G443gat), .dout(n5624));
    jnot g1458(.din(n5624), .dout(n5627));
    jand g1459(.dinb(n28453), .dina(n5425), .dout(n5631));
    jand g1460(.dinb(n28450), .dina(n5429), .dout(n5635));
    jor g1461(.dinb(n28363), .dina(n5635), .dout(n5639));
    jand g1462(.dinb(G222gat), .dina(G426gat), .dout(n5643));
    jnot g1463(.din(n5643), .dout(n5646));
    jand g1464(.dinb(n32167), .dina(n5417), .dout(n5650));
    jand g1465(.dinb(n32008), .dina(n5421), .dout(n5654));
    jor g1466(.dinb(n31927), .dina(n5654), .dout(n5658));
    jand g1467(.dinb(G239gat), .dina(G409gat), .dout(n5662));
    jand g1468(.dinb(G256gat), .dina(G392gat), .dout(n5666));
    jor g1469(.dinb(n32086), .dina(n5406), .dout(n5670));
    jor g1470(.dinb(n32164), .dina(n5413), .dout(n5674));
    jand g1471(.dinb(n31747), .dina(n5674), .dout(n5678));
    jxor g1472(.dinb(n31831), .dina(n5678), .dout(n5682));
    jnot g1473(.din(n5682), .dout(n5685));
    jxor g1474(.dinb(n31921), .dina(n5685), .dout(n5689));
    jxor g1475(.dinb(n31924), .dina(n5689), .dout(n5693));
    jxor g1476(.dinb(n31741), .dina(n5693), .dout(n5697));
    jxor g1477(.dinb(n28360), .dina(n5697), .dout(n5701));
    jxor g1478(.dinb(n28357), .dina(n5701), .dout(n5705));
    jxor g1479(.dinb(n26962), .dina(n5705), .dout(n5709));
    jxor g1480(.dinb(n26959), .dina(n5709), .dout(n5713));
    jxor g1481(.dinb(n25597), .dina(n5713), .dout(n5717));
    jxor g1482(.dinb(n25594), .dina(n5717), .dout(n5721));
    jxor g1483(.dinb(n5582), .dina(n5721), .dout(n5725));
    jxor g1484(.dinb(n24250), .dina(n5725), .dout(n5729));
    jxor g1485(.dinb(n5563), .dina(n22912), .dout(n5733));
    jxor g1486(.dinb(n22909), .dina(n5733), .dout(n5737));
    jxor g1487(.dinb(n5544), .dina(n21573), .dout(n5741));
    jnot g1488(.din(n5741), .dout(n5744));
    jxor g1489(.dinb(n21568), .dina(n5744), .dout(n5748));
    jnot g1490(.din(n5748), .dout(n5751));
    jxor g1491(.dinb(n20338), .dina(n5751), .dout(n5755));
    jxor g1492(.dinb(n5510), .dina(n12720), .dout(n5759));
    jor g1493(.dinb(n20338), .dina(n5751), .dout(n5763));
    jnot g1494(.din(n5755), .dout(n5766));
    jor g1495(.dinb(n5510), .dina(n12718), .dout(n5770));
    jand g1496(.dinb(n12700), .dina(n5770), .dout(n5774));
    jnot g1497(.din(n5544), .dout(n5777));
    jnot g1498(.din(n5737), .dout(n5780));
    jor g1499(.dinb(n5777), .dina(n21571), .dout(n5784));
    jor g1500(.dinb(n21568), .dina(n5744), .dout(n5788));
    jand g1501(.dinb(n21427), .dina(n5788), .dout(n5792));
    jand g1502(.dinb(G137gat), .dina(G528gat), .dout(n5796));
    jand g1503(.dinb(n5563), .dina(n22912), .dout(n5800));
    jand g1504(.dinb(n22909), .dina(n5733), .dout(n5804));
    jor g1505(.dinb(n22783), .dina(n5804), .dout(n5808));
    jand g1506(.dinb(G154gat), .dina(G511gat), .dout(n5812));
    jnot g1507(.din(n5812), .dout(n5815));
    jand g1508(.dinb(n5582), .dina(n5721), .dout(n5819));
    jand g1509(.dinb(n24250), .dina(n5725), .dout(n5823));
    jor g1510(.dinb(n24133), .dina(n5823), .dout(n5827));
    jand g1511(.dinb(G171gat), .dina(G494gat), .dout(n5831));
    jnot g1512(.din(n5831), .dout(n5834));
    jand g1513(.dinb(n25597), .dina(n5713), .dout(n5838));
    jand g1514(.dinb(n25594), .dina(n5717), .dout(n5842));
    jor g1515(.dinb(n25483), .dina(n5842), .dout(n5846));
    jand g1516(.dinb(G188gat), .dina(G477gat), .dout(n5850));
    jnot g1517(.din(n5850), .dout(n5853));
    jand g1518(.dinb(n26962), .dina(n5705), .dout(n5857));
    jand g1519(.dinb(n26959), .dina(n5709), .dout(n5861));
    jor g1520(.dinb(n26854), .dina(n5861), .dout(n5865));
    jand g1521(.dinb(G205gat), .dina(G460gat), .dout(n5869));
    jnot g1522(.din(n5869), .dout(n5872));
    jand g1523(.dinb(n28360), .dina(n5697), .dout(n5876));
    jand g1524(.dinb(n28357), .dina(n5701), .dout(n5880));
    jor g1525(.dinb(n28258), .dina(n5880), .dout(n5884));
    jand g1526(.dinb(G222gat), .dina(G443gat), .dout(n5888));
    jnot g1527(.din(n5888), .dout(n5891));
    jand g1528(.dinb(n31924), .dina(n5689), .dout(n5895));
    jand g1529(.dinb(n31741), .dina(n5693), .dout(n5899));
    jor g1530(.dinb(n31648), .dina(n5899), .dout(n5903));
    jand g1531(.dinb(G239gat), .dina(G426gat), .dout(n5907));
    jand g1532(.dinb(G256gat), .dina(G409gat), .dout(n5911));
    jor g1533(.dinb(n31831), .dina(n5678), .dout(n5915));
    jor g1534(.dinb(n31921), .dina(n5685), .dout(n5919));
    jand g1535(.dinb(n31444), .dina(n5919), .dout(n5923));
    jxor g1536(.dinb(n31540), .dina(n5923), .dout(n5927));
    jnot g1537(.din(n5927), .dout(n5930));
    jxor g1538(.dinb(n31642), .dina(n5930), .dout(n5934));
    jxor g1539(.dinb(n31645), .dina(n5934), .dout(n5938));
    jxor g1540(.dinb(n31438), .dina(n5938), .dout(n5942));
    jxor g1541(.dinb(n28255), .dina(n5942), .dout(n5946));
    jxor g1542(.dinb(n28252), .dina(n5946), .dout(n5950));
    jxor g1543(.dinb(n26851), .dina(n5950), .dout(n5954));
    jxor g1544(.dinb(n26848), .dina(n5954), .dout(n5958));
    jxor g1545(.dinb(n25480), .dina(n5958), .dout(n5962));
    jxor g1546(.dinb(n25477), .dina(n5962), .dout(n5966));
    jxor g1547(.dinb(n24130), .dina(n5966), .dout(n5970));
    jxor g1548(.dinb(n24127), .dina(n5970), .dout(n5974));
    jxor g1549(.dinb(n5808), .dina(n5974), .dout(n5978));
    jnot g1550(.din(n5978), .dout(n5981));
    jxor g1551(.dinb(n22780), .dina(n5981), .dout(n5985));
    jnot g1552(.din(n5985), .dout(n5988));
    jxor g1553(.dinb(n5792), .dina(n5988), .dout(n5992));
    jxor g1554(.dinb(n5774), .dina(n12651), .dout(n5996));
    jor g1555(.dinb(n5792), .dina(n5988), .dout(n6000));
    jnot g1556(.din(n5992), .dout(n6003));
    jor g1557(.dinb(n5774), .dina(n12649), .dout(n6007));
    jand g1558(.dinb(n12625), .dina(n6007), .dout(n6011));
    jnot g1559(.din(n5808), .dout(n6014));
    jnot g1560(.din(n5974), .dout(n6017));
    jor g1561(.dinb(n6014), .dina(n6017), .dout(n6021));
    jor g1562(.dinb(n22780), .dina(n5981), .dout(n6025));
    jand g1563(.dinb(n22639), .dina(n6025), .dout(n6029));
    jand g1564(.dinb(G154gat), .dina(G528gat), .dout(n6033));
    jand g1565(.dinb(n24130), .dina(n5966), .dout(n6037));
    jand g1566(.dinb(n24127), .dina(n5970), .dout(n6041));
    jor g1567(.dinb(n23998), .dina(n6041), .dout(n6045));
    jand g1568(.dinb(G171gat), .dina(G511gat), .dout(n6049));
    jnot g1569(.din(n6049), .dout(n6052));
    jand g1570(.dinb(n25480), .dina(n5958), .dout(n6056));
    jand g1571(.dinb(n25477), .dina(n5962), .dout(n6060));
    jor g1572(.dinb(n25354), .dina(n6060), .dout(n6064));
    jand g1573(.dinb(G188gat), .dina(G494gat), .dout(n6068));
    jnot g1574(.din(n6068), .dout(n6071));
    jand g1575(.dinb(n26851), .dina(n5950), .dout(n6075));
    jand g1576(.dinb(n26848), .dina(n5954), .dout(n6079));
    jor g1577(.dinb(n26731), .dina(n6079), .dout(n6083));
    jand g1578(.dinb(G205gat), .dina(G477gat), .dout(n6087));
    jnot g1579(.din(n6087), .dout(n6090));
    jand g1580(.dinb(n28255), .dina(n5942), .dout(n6094));
    jand g1581(.dinb(n28252), .dina(n5946), .dout(n6098));
    jor g1582(.dinb(n28141), .dina(n6098), .dout(n6102));
    jand g1583(.dinb(G222gat), .dina(G460gat), .dout(n6106));
    jnot g1584(.din(n6106), .dout(n6109));
    jand g1585(.dinb(n31645), .dina(n5934), .dout(n6113));
    jand g1586(.dinb(n31438), .dina(n5938), .dout(n6117));
    jor g1587(.dinb(n31333), .dina(n6117), .dout(n6121));
    jand g1588(.dinb(G239gat), .dina(G443gat), .dout(n6125));
    jand g1589(.dinb(G256gat), .dina(G426gat), .dout(n6129));
    jor g1590(.dinb(n31540), .dina(n5923), .dout(n6133));
    jor g1591(.dinb(n31642), .dina(n5930), .dout(n6137));
    jand g1592(.dinb(n31105), .dina(n6137), .dout(n6141));
    jxor g1593(.dinb(n31213), .dina(n6141), .dout(n6145));
    jnot g1594(.din(n6145), .dout(n6148));
    jxor g1595(.dinb(n31327), .dina(n6148), .dout(n6152));
    jxor g1596(.dinb(n31330), .dina(n6152), .dout(n6156));
    jxor g1597(.dinb(n31099), .dina(n6156), .dout(n6160));
    jxor g1598(.dinb(n28138), .dina(n6160), .dout(n6164));
    jxor g1599(.dinb(n28135), .dina(n6164), .dout(n6168));
    jxor g1600(.dinb(n26728), .dina(n6168), .dout(n6172));
    jxor g1601(.dinb(n26725), .dina(n6172), .dout(n6176));
    jxor g1602(.dinb(n25351), .dina(n6176), .dout(n6180));
    jxor g1603(.dinb(n25348), .dina(n6180), .dout(n6184));
    jxor g1604(.dinb(n23994), .dina(n6184), .dout(n6188));
    jnot g1605(.din(n6188), .dout(n6191));
    jxor g1606(.dinb(n23989), .dina(n6191), .dout(n6195));
    jnot g1607(.din(n6195), .dout(n6198));
    jxor g1608(.dinb(n22636), .dina(n6198), .dout(n6202));
    jxor g1609(.dinb(n6011), .dina(n12570), .dout(n6206));
    jor g1610(.dinb(n22636), .dina(n6198), .dout(n6210));
    jnot g1611(.din(n6202), .dout(n6213));
    jor g1612(.dinb(n6011), .dina(n12568), .dout(n6217));
    jand g1613(.dinb(n12544), .dina(n6217), .dout(n6221));
    jnot g1614(.din(n6045), .dout(n6224));
    jnot g1615(.din(n6184), .dout(n6227));
    jor g1616(.dinb(n23992), .dina(n6227), .dout(n6231));
    jor g1617(.dinb(n23989), .dina(n6191), .dout(n6235));
    jand g1618(.dinb(n23842), .dina(n6235), .dout(n6239));
    jand g1619(.dinb(G171gat), .dina(G528gat), .dout(n6243));
    jnot g1620(.din(n6243), .dout(n6246));
    jand g1621(.dinb(n25351), .dina(n6176), .dout(n6250));
    jand g1622(.dinb(n25348), .dina(n6180), .dout(n6254));
    jor g1623(.dinb(n25213), .dina(n6254), .dout(n6258));
    jand g1624(.dinb(G188gat), .dina(G511gat), .dout(n6262));
    jnot g1625(.din(n6262), .dout(n6265));
    jand g1626(.dinb(n26728), .dina(n6168), .dout(n6269));
    jand g1627(.dinb(n26725), .dina(n6172), .dout(n6273));
    jor g1628(.dinb(n26596), .dina(n6273), .dout(n6277));
    jand g1629(.dinb(G205gat), .dina(G494gat), .dout(n6281));
    jnot g1630(.din(n6281), .dout(n6284));
    jand g1631(.dinb(n28138), .dina(n6160), .dout(n6288));
    jand g1632(.dinb(n28135), .dina(n6164), .dout(n6292));
    jor g1633(.dinb(n28012), .dina(n6292), .dout(n6296));
    jand g1634(.dinb(G222gat), .dina(G477gat), .dout(n6300));
    jnot g1635(.din(n6300), .dout(n6303));
    jand g1636(.dinb(n31330), .dina(n6152), .dout(n6307));
    jand g1637(.dinb(n31099), .dina(n6156), .dout(n6311));
    jor g1638(.dinb(n30982), .dina(n6311), .dout(n6315));
    jand g1639(.dinb(G239gat), .dina(G460gat), .dout(n6319));
    jand g1640(.dinb(G256gat), .dina(G443gat), .dout(n6323));
    jor g1641(.dinb(n31213), .dina(n6141), .dout(n6327));
    jor g1642(.dinb(n31327), .dina(n6148), .dout(n6331));
    jand g1643(.dinb(n30730), .dina(n6331), .dout(n6335));
    jxor g1644(.dinb(n30850), .dina(n6335), .dout(n6339));
    jnot g1645(.din(n6339), .dout(n6342));
    jxor g1646(.dinb(n30976), .dina(n6342), .dout(n6346));
    jxor g1647(.dinb(n30979), .dina(n6346), .dout(n6350));
    jxor g1648(.dinb(n30724), .dina(n6350), .dout(n6354));
    jxor g1649(.dinb(n28009), .dina(n6354), .dout(n6358));
    jxor g1650(.dinb(n28006), .dina(n6358), .dout(n6362));
    jxor g1651(.dinb(n26593), .dina(n6362), .dout(n6366));
    jxor g1652(.dinb(n26590), .dina(n6366), .dout(n6370));
    jxor g1653(.dinb(n25210), .dina(n6370), .dout(n6374));
    jxor g1654(.dinb(n25207), .dina(n6374), .dout(n6378));
    jnot g1655(.din(n6378), .dout(n6381));
    jxor g1656(.dinb(n23839), .dina(n6381), .dout(n6385));
    jxor g1657(.dinb(n6221), .dina(n12486), .dout(n6389));
    jor g1658(.dinb(n23839), .dina(n6381), .dout(n6393));
    jnot g1659(.din(n6385), .dout(n6396));
    jor g1660(.dinb(n6221), .dina(n12484), .dout(n6400));
    jand g1661(.dinb(n12457), .dina(n6400), .dout(n6404));
    jand g1662(.dinb(n25210), .dina(n6370), .dout(n6408));
    jand g1663(.dinb(n25207), .dina(n6374), .dout(n6412));
    jor g1664(.dinb(n25060), .dina(n6412), .dout(n6416));
    jand g1665(.dinb(G188gat), .dina(G528gat), .dout(n6420));
    jnot g1666(.din(n6420), .dout(n6423));
    jand g1667(.dinb(n26593), .dina(n6362), .dout(n6427));
    jand g1668(.dinb(n26590), .dina(n6366), .dout(n6431));
    jor g1669(.dinb(n26449), .dina(n6431), .dout(n6435));
    jand g1670(.dinb(G205gat), .dina(G511gat), .dout(n6439));
    jnot g1671(.din(n6439), .dout(n6442));
    jand g1672(.dinb(n28009), .dina(n6354), .dout(n6446));
    jand g1673(.dinb(n28006), .dina(n6358), .dout(n6450));
    jor g1674(.dinb(n27871), .dina(n6450), .dout(n6454));
    jand g1675(.dinb(G222gat), .dina(G494gat), .dout(n6458));
    jnot g1676(.din(n6458), .dout(n6461));
    jand g1677(.dinb(n30979), .dina(n6346), .dout(n6465));
    jand g1678(.dinb(n30724), .dina(n6350), .dout(n6469));
    jor g1679(.dinb(n30595), .dina(n6469), .dout(n6473));
    jand g1680(.dinb(G239gat), .dina(G477gat), .dout(n6477));
    jand g1681(.dinb(G256gat), .dina(G460gat), .dout(n6481));
    jor g1682(.dinb(n30850), .dina(n6335), .dout(n6485));
    jor g1683(.dinb(n30976), .dina(n6342), .dout(n6489));
    jand g1684(.dinb(n30319), .dina(n6489), .dout(n6493));
    jxor g1685(.dinb(n30451), .dina(n6493), .dout(n6497));
    jnot g1686(.din(n6497), .dout(n6500));
    jxor g1687(.dinb(n30589), .dina(n6500), .dout(n6504));
    jxor g1688(.dinb(n30592), .dina(n6504), .dout(n6508));
    jxor g1689(.dinb(n30313), .dina(n6508), .dout(n6512));
    jxor g1690(.dinb(n27868), .dina(n6512), .dout(n6516));
    jxor g1691(.dinb(n27865), .dina(n6516), .dout(n6520));
    jxor g1692(.dinb(n26446), .dina(n6520), .dout(n6524));
    jxor g1693(.dinb(n26443), .dina(n6524), .dout(n6528));
    jxor g1694(.dinb(n25056), .dina(n6528), .dout(n6532));
    jxor g1695(.dinb(n6404), .dina(n12393), .dout(n6536));
    jnot g1696(.din(n6416), .dout(n6539));
    jnot g1697(.din(n6528), .dout(n6542));
    jor g1698(.dinb(n25054), .dina(n6542), .dout(n6546));
    jnot g1699(.din(n6532), .dout(n6549));
    jor g1700(.dinb(n6404), .dina(n12391), .dout(n6553));
    jand g1701(.dinb(n12361), .dina(n6553), .dout(n6557));
    jand g1702(.dinb(n26446), .dina(n6520), .dout(n6561));
    jand g1703(.dinb(n26443), .dina(n6524), .dout(n6565));
    jor g1704(.dinb(n26290), .dina(n6565), .dout(n6569));
    jand g1705(.dinb(G205gat), .dina(G528gat), .dout(n6573));
    jnot g1706(.din(n6573), .dout(n6576));
    jand g1707(.dinb(n27868), .dina(n6512), .dout(n6580));
    jand g1708(.dinb(n27865), .dina(n6516), .dout(n6584));
    jor g1709(.dinb(n27718), .dina(n6584), .dout(n6588));
    jand g1710(.dinb(G222gat), .dina(G511gat), .dout(n6592));
    jnot g1711(.din(n6592), .dout(n6595));
    jand g1712(.dinb(n30592), .dina(n6504), .dout(n6599));
    jand g1713(.dinb(n30313), .dina(n6508), .dout(n6603));
    jor g1714(.dinb(n30172), .dina(n6603), .dout(n6607));
    jand g1715(.dinb(G239gat), .dina(G494gat), .dout(n6611));
    jand g1716(.dinb(G256gat), .dina(G477gat), .dout(n6615));
    jor g1717(.dinb(n30451), .dina(n6493), .dout(n6619));
    jor g1718(.dinb(n30589), .dina(n6500), .dout(n6623));
    jand g1719(.dinb(n29872), .dina(n6623), .dout(n6627));
    jxor g1720(.dinb(n30016), .dina(n6627), .dout(n6631));
    jnot g1721(.din(n6631), .dout(n6634));
    jxor g1722(.dinb(n30166), .dina(n6634), .dout(n6638));
    jxor g1723(.dinb(n30169), .dina(n6638), .dout(n6642));
    jxor g1724(.dinb(n29866), .dina(n6642), .dout(n6646));
    jxor g1725(.dinb(n27715), .dina(n6646), .dout(n6650));
    jxor g1726(.dinb(n27712), .dina(n6650), .dout(n6654));
    jxor g1727(.dinb(n26286), .dina(n6654), .dout(n6658));
    jxor g1728(.dinb(n6557), .dina(n12297), .dout(n6662));
    jnot g1729(.din(n6569), .dout(n6665));
    jnot g1730(.din(n6654), .dout(n6668));
    jor g1731(.dinb(n26284), .dina(n6668), .dout(n6672));
    jnot g1732(.din(n6658), .dout(n6675));
    jor g1733(.dinb(n6557), .dina(n12295), .dout(n6679));
    jand g1734(.dinb(n12265), .dina(n6679), .dout(n6683));
    jand g1735(.dinb(n27715), .dina(n6646), .dout(n6687));
    jand g1736(.dinb(n27712), .dina(n6650), .dout(n6691));
    jor g1737(.dinb(n27553), .dina(n6691), .dout(n6695));
    jand g1738(.dinb(G222gat), .dina(G528gat), .dout(n6699));
    jnot g1739(.din(n6699), .dout(n6702));
    jand g1740(.dinb(n30169), .dina(n6638), .dout(n6706));
    jand g1741(.dinb(n29866), .dina(n6642), .dout(n6710));
    jor g1742(.dinb(n29713), .dina(n6710), .dout(n6714));
    jand g1743(.dinb(G239gat), .dina(G511gat), .dout(n6718));
    jand g1744(.dinb(G256gat), .dina(G494gat), .dout(n6722));
    jor g1745(.dinb(n30016), .dina(n6627), .dout(n6726));
    jor g1746(.dinb(n30166), .dina(n6634), .dout(n6730));
    jand g1747(.dinb(n29389), .dina(n6730), .dout(n6734));
    jxor g1748(.dinb(n29545), .dina(n6734), .dout(n6738));
    jnot g1749(.din(n6738), .dout(n6741));
    jxor g1750(.dinb(n29707), .dina(n6741), .dout(n6745));
    jxor g1751(.dinb(n29710), .dina(n6745), .dout(n6749));
    jxor g1752(.dinb(n29383), .dina(n6749), .dout(n6753));
    jxor g1753(.dinb(n27549), .dina(n6753), .dout(n6757));
    jxor g1754(.dinb(n6683), .dina(n12201), .dout(n6761));
    jnot g1755(.din(n6695), .dout(n6764));
    jnot g1756(.din(n6753), .dout(n6767));
    jor g1757(.dinb(n27547), .dina(n6767), .dout(n6771));
    jnot g1758(.din(n6757), .dout(n6774));
    jor g1759(.dinb(n6683), .dina(n12199), .dout(n6778));
    jand g1760(.dinb(n12169), .dina(n6778), .dout(n6782));
    jand g1761(.dinb(n29710), .dina(n6745), .dout(n6786));
    jand g1762(.dinb(n29383), .dina(n6749), .dout(n6790));
    jor g1763(.dinb(n29218), .dina(n6790), .dout(n6794));
    jand g1764(.dinb(G239gat), .dina(G528gat), .dout(n6798));
    jand g1765(.dinb(G256gat), .dina(G511gat), .dout(n6802));
    jor g1766(.dinb(n29545), .dina(n6734), .dout(n6806));
    jor g1767(.dinb(n29707), .dina(n6741), .dout(n6810));
    jand g1768(.dinb(n28870), .dina(n6810), .dout(n6814));
    jxor g1769(.dinb(n29038), .dina(n6814), .dout(n6818));
    jnot g1770(.din(n6818), .dout(n6821));
    jxor g1771(.dinb(n29212), .dina(n6821), .dout(n6825));
    jxor g1772(.dinb(n29214), .dina(n6825), .dout(n6829));
    jxor g1773(.dinb(n6782), .dina(n12105), .dout(n6833));
    jand g1774(.dinb(G256gat), .dina(G528gat), .dout(n6837));
    jor g1775(.dinb(n29038), .dina(n6814), .dout(n6841));
    jor g1776(.dinb(n29212), .dina(n6821), .dout(n6845));
    jand g1777(.dinb(n11860), .dina(n6845), .dout(n6849));
    jor g1778(.dinb(n12040), .dina(n6849), .dout(n6853));
    jnot g1779(.din(n6794), .dout(n6856));
    jnot g1780(.din(n6825), .dout(n6859));
    jor g1781(.dinb(n28864), .dina(n6859), .dout(n6863));
    jnot g1782(.din(n6829), .dout(n6866));
    jor g1783(.dinb(n6782), .dina(n12103), .dout(n6870));
    jand g1784(.dinb(n12073), .dina(n6870), .dout(n6874));
    jxor g1785(.dinb(n12040), .dina(n6849), .dout(n6878));
    jnot g1786(.din(n6878), .dout(n6881));
    jor g1787(.dinb(n6874), .dina(n11818), .dout(n6885));
    jand g1788(.dinb(n11785), .dina(n6885), .dout(G6287gat));
    jxor g1789(.dinb(n6874), .dina(n11820), .dout(n6893));
    jdff dff_A_Sal8trTP1_2(.din(n6893), .dout(G6288gat));
    jdff dff_A_Axb5Z3Rn6_0(.din(n36090), .dout(G6280gat));
    jdff dff_A_PeO9O6Ih5_0(.din(n36087), .dout(n36090));
    jdff dff_A_8IBM46XT7_2(.din(n6833), .dout(n36087));
    jdff dff_A_MHHB6UYJ2_0(.din(n36081), .dout(G6270gat));
    jdff dff_A_6OgvdeOL1_0(.din(n36078), .dout(n36081));
    jdff dff_A_ifSQI7J07_0(.din(n36075), .dout(n36078));
    jdff dff_A_4TathcMT6_0(.din(n36072), .dout(n36075));
    jdff dff_A_WJUS03tP8_2(.din(n6761), .dout(n36072));
    jdff dff_A_VtpZWgPZ6_0(.din(n36066), .dout(G6260gat));
    jdff dff_A_C1glzCQw2_0(.din(n36063), .dout(n36066));
    jdff dff_A_QFPb4j7j6_0(.din(n36060), .dout(n36063));
    jdff dff_A_GG2KKa2p5_0(.din(n36057), .dout(n36060));
    jdff dff_A_W6uKVywC5_0(.din(n36054), .dout(n36057));
    jdff dff_A_C1CdSTLN7_0(.din(n36051), .dout(n36054));
    jdff dff_A_ItMjlGlT1_2(.din(n6662), .dout(n36051));
    jdff dff_A_he6AWlgo8_0(.din(n36045), .dout(G6250gat));
    jdff dff_A_pUDoKapv1_0(.din(n36042), .dout(n36045));
    jdff dff_A_S2fxXnOh9_0(.din(n36039), .dout(n36042));
    jdff dff_A_zWPEkxoE8_0(.din(n36036), .dout(n36039));
    jdff dff_A_dpmFDk4l4_0(.din(n36033), .dout(n36036));
    jdff dff_A_EGkVELoi0_0(.din(n36030), .dout(n36033));
    jdff dff_A_NaxIzPxG7_0(.din(n36027), .dout(n36030));
    jdff dff_A_4W1dVK516_0(.din(n36024), .dout(n36027));
    jdff dff_A_3iLVSEwm9_2(.din(n6536), .dout(n36024));
    jdff dff_A_v64lkwQT4_0(.din(n36018), .dout(G6240gat));
    jdff dff_A_O5HVrv8X7_0(.din(n36015), .dout(n36018));
    jdff dff_A_fwuPYOIa2_0(.din(n36012), .dout(n36015));
    jdff dff_A_PFx33hNw4_0(.din(n36009), .dout(n36012));
    jdff dff_A_dMe4vE8R8_0(.din(n36006), .dout(n36009));
    jdff dff_A_LK6wRUxT8_0(.din(n36003), .dout(n36006));
    jdff dff_A_S33jOICy7_0(.din(n36000), .dout(n36003));
    jdff dff_A_BovAFiDd6_0(.din(n35997), .dout(n36000));
    jdff dff_A_JL78wWS26_0(.din(n35994), .dout(n35997));
    jdff dff_A_Jd6PsPPu4_0(.din(n35991), .dout(n35994));
    jdff dff_A_hXEXHGJP4_2(.din(n6389), .dout(n35991));
    jdff dff_A_tVYZQ0xk2_0(.din(n35985), .dout(G6230gat));
    jdff dff_A_jemr7PEt7_0(.din(n35982), .dout(n35985));
    jdff dff_A_VxSjdbXL3_0(.din(n35979), .dout(n35982));
    jdff dff_A_B1mpiYQK7_0(.din(n35976), .dout(n35979));
    jdff dff_A_KMCrbG5i2_0(.din(n35973), .dout(n35976));
    jdff dff_A_C9lOJ36M2_0(.din(n35970), .dout(n35973));
    jdff dff_A_EDFDqcWu2_0(.din(n35967), .dout(n35970));
    jdff dff_A_EP4Nrif76_0(.din(n35964), .dout(n35967));
    jdff dff_A_CltQHqxN1_0(.din(n35961), .dout(n35964));
    jdff dff_A_QV3e7I3m6_0(.din(n35958), .dout(n35961));
    jdff dff_A_At2BKpWp7_0(.din(n35955), .dout(n35958));
    jdff dff_A_hboK2Rm15_0(.din(n35952), .dout(n35955));
    jdff dff_A_LmfDc3mX7_2(.din(n6206), .dout(n35952));
    jdff dff_A_zFU6cqn04_0(.din(n35946), .dout(G6220gat));
    jdff dff_A_FhgJ3KMa0_0(.din(n35943), .dout(n35946));
    jdff dff_A_ReOMoYRg9_0(.din(n35940), .dout(n35943));
    jdff dff_A_zvqnxQ0t7_0(.din(n35937), .dout(n35940));
    jdff dff_A_AidrJimb7_0(.din(n35934), .dout(n35937));
    jdff dff_A_TNemDBlJ5_0(.din(n35931), .dout(n35934));
    jdff dff_A_p3fTEORF6_0(.din(n35928), .dout(n35931));
    jdff dff_A_XiOyo2uX4_0(.din(n35925), .dout(n35928));
    jdff dff_A_csAyt3t46_0(.din(n35922), .dout(n35925));
    jdff dff_A_EvwOX0nf7_0(.din(n35919), .dout(n35922));
    jdff dff_A_h9JzAGb39_0(.din(n35916), .dout(n35919));
    jdff dff_A_93feg0hY2_0(.din(n35913), .dout(n35916));
    jdff dff_A_3phXYowu3_0(.din(n35910), .dout(n35913));
    jdff dff_A_Zvp8zY511_0(.din(n35907), .dout(n35910));
    jdff dff_A_bLrqy25k9_2(.din(n5996), .dout(n35907));
    jdff dff_A_q0ovqedw9_0(.din(n35901), .dout(G6210gat));
    jdff dff_A_Wqx6ig220_0(.din(n35898), .dout(n35901));
    jdff dff_A_LHDF6mO28_0(.din(n35895), .dout(n35898));
    jdff dff_A_ngYzzIIk4_0(.din(n35892), .dout(n35895));
    jdff dff_A_b9Imky7T9_0(.din(n35889), .dout(n35892));
    jdff dff_A_uTlf0yaM5_0(.din(n35886), .dout(n35889));
    jdff dff_A_KxfVw64E6_0(.din(n35883), .dout(n35886));
    jdff dff_A_Yq6pLs3I3_0(.din(n35880), .dout(n35883));
    jdff dff_A_fr2ZZxGV7_0(.din(n35877), .dout(n35880));
    jdff dff_A_xU2xglG99_0(.din(n35874), .dout(n35877));
    jdff dff_A_taIrpx5f3_0(.din(n35871), .dout(n35874));
    jdff dff_A_vYYr7qNX5_0(.din(n35868), .dout(n35871));
    jdff dff_A_6lpCmimB2_0(.din(n35865), .dout(n35868));
    jdff dff_A_XPescyqL8_0(.din(n35862), .dout(n35865));
    jdff dff_A_U1EP0ICI1_0(.din(n35859), .dout(n35862));
    jdff dff_A_xQeTjuds5_0(.din(n35856), .dout(n35859));
    jdff dff_A_IUYnNff39_2(.din(n5759), .dout(n35856));
    jdff dff_A_CwF0X3Qt5_0(.din(n35850), .dout(G6200gat));
    jdff dff_A_ryZ5pVjc1_0(.din(n35847), .dout(n35850));
    jdff dff_A_nNDroKgT3_0(.din(n35844), .dout(n35847));
    jdff dff_A_OS4F2H9T4_0(.din(n35841), .dout(n35844));
    jdff dff_A_JSEHANbP2_0(.din(n35838), .dout(n35841));
    jdff dff_A_RiKmipjv3_0(.din(n35835), .dout(n35838));
    jdff dff_A_Tfh6mXU79_0(.din(n35832), .dout(n35835));
    jdff dff_A_oTcZHgAl7_0(.din(n35829), .dout(n35832));
    jdff dff_A_gQCbsAhm6_0(.din(n35826), .dout(n35829));
    jdff dff_A_pzlp7gQm8_0(.din(n35823), .dout(n35826));
    jdff dff_A_4KyxBQfF9_0(.din(n35820), .dout(n35823));
    jdff dff_A_qQ7jFv5L9_0(.din(n35817), .dout(n35820));
    jdff dff_A_u2jthr0Z6_0(.din(n35814), .dout(n35817));
    jdff dff_A_nUyTD8ts3_0(.din(n35811), .dout(n35814));
    jdff dff_A_1vdIsrcS5_0(.din(n35808), .dout(n35811));
    jdff dff_A_QVEmwyc12_0(.din(n35805), .dout(n35808));
    jdff dff_A_aQIhDYMB0_0(.din(n35802), .dout(n35805));
    jdff dff_A_mGau4jRS5_0(.din(n35799), .dout(n35802));
    jdff dff_A_DbIDePej4_2(.din(n5495), .dout(n35799));
    jdff dff_A_4Tot9Ke45_0(.din(n35793), .dout(G6190gat));
    jdff dff_A_QDexrUex8_0(.din(n35790), .dout(n35793));
    jdff dff_A_ixdpxXyl9_0(.din(n35787), .dout(n35790));
    jdff dff_A_T6qWt4nx7_0(.din(n35784), .dout(n35787));
    jdff dff_A_bOQ97r6R4_0(.din(n35781), .dout(n35784));
    jdff dff_A_8jUGBtcG2_0(.din(n35778), .dout(n35781));
    jdff dff_A_kJMyCwVs3_0(.din(n35775), .dout(n35778));
    jdff dff_A_mHVkNbvH7_0(.din(n35772), .dout(n35775));
    jdff dff_A_CaEvomZQ3_0(.din(n35769), .dout(n35772));
    jdff dff_A_W7qz9fsH8_0(.din(n35766), .dout(n35769));
    jdff dff_A_bLdR2FXj9_0(.din(n35763), .dout(n35766));
    jdff dff_A_gTtrjauN9_0(.din(n35760), .dout(n35763));
    jdff dff_A_138kPFry8_0(.din(n35757), .dout(n35760));
    jdff dff_A_dWzIwmUM7_0(.din(n35754), .dout(n35757));
    jdff dff_A_UfmbiT5a1_0(.din(n35751), .dout(n35754));
    jdff dff_A_xjdaaH8o2_0(.din(n35748), .dout(n35751));
    jdff dff_A_W2hvF0zz0_0(.din(n35745), .dout(n35748));
    jdff dff_A_UiZcUW5a0_0(.din(n35742), .dout(n35745));
    jdff dff_A_YziWlVof8_0(.din(n35739), .dout(n35742));
    jdff dff_A_prtqAZc98_0(.din(n35736), .dout(n35739));
    jdff dff_A_0iZHqm6h1_2(.din(n5204), .dout(n35736));
    jdff dff_A_jIx7cOiV7_0(.din(n35730), .dout(G6180gat));
    jdff dff_A_2s2nWD7l1_0(.din(n35727), .dout(n35730));
    jdff dff_A_WwhykUhZ0_0(.din(n35724), .dout(n35727));
    jdff dff_A_FdyIXHAm7_0(.din(n35721), .dout(n35724));
    jdff dff_A_qHkWz9bX2_0(.din(n35718), .dout(n35721));
    jdff dff_A_IulUPpmL5_0(.din(n35715), .dout(n35718));
    jdff dff_A_Eo0iLPBH0_0(.din(n35712), .dout(n35715));
    jdff dff_A_LYPqDeu10_0(.din(n35709), .dout(n35712));
    jdff dff_A_gSEeBq5e7_0(.din(n35706), .dout(n35709));
    jdff dff_A_gGj8T90x1_0(.din(n35703), .dout(n35706));
    jdff dff_A_TwcTavwt2_0(.din(n35700), .dout(n35703));
    jdff dff_A_9t9c2ZSL7_0(.din(n35697), .dout(n35700));
    jdff dff_A_N4255XaA4_0(.din(n35694), .dout(n35697));
    jdff dff_A_DrbsFgqW9_0(.din(n35691), .dout(n35694));
    jdff dff_A_l0SLvcbN7_0(.din(n35688), .dout(n35691));
    jdff dff_A_gc57QrSY6_0(.din(n35685), .dout(n35688));
    jdff dff_A_qN60RfzG1_0(.din(n35682), .dout(n35685));
    jdff dff_A_XzSjgAJD4_0(.din(n35679), .dout(n35682));
    jdff dff_A_j61eup6U3_0(.din(n35676), .dout(n35679));
    jdff dff_A_mIRvBGgs2_0(.din(n35673), .dout(n35676));
    jdff dff_A_Vl6XXqKR4_0(.din(n35670), .dout(n35673));
    jdff dff_A_s8Lz3PP21_0(.din(n35667), .dout(n35670));
    jdff dff_A_XYc3sDAs5_2(.din(n4886), .dout(n35667));
    jdff dff_A_wJ6PBTgs4_0(.din(n35661), .dout(G6170gat));
    jdff dff_A_ytUpiMlJ5_0(.din(n35658), .dout(n35661));
    jdff dff_A_gM8cknpP4_0(.din(n35655), .dout(n35658));
    jdff dff_A_kFu9MVUT3_0(.din(n35652), .dout(n35655));
    jdff dff_A_LwNB3OKs1_0(.din(n35649), .dout(n35652));
    jdff dff_A_HvckR75J2_0(.din(n35646), .dout(n35649));
    jdff dff_A_oIOw8cGC7_0(.din(n35643), .dout(n35646));
    jdff dff_A_WEVIotbk2_0(.din(n35640), .dout(n35643));
    jdff dff_A_wK1dcayQ8_0(.din(n35637), .dout(n35640));
    jdff dff_A_ZPeyBSXX7_0(.din(n35634), .dout(n35637));
    jdff dff_A_vlDewE9B9_0(.din(n35631), .dout(n35634));
    jdff dff_A_tbZj41kF9_0(.din(n35628), .dout(n35631));
    jdff dff_A_ofAzioCB2_0(.din(n35625), .dout(n35628));
    jdff dff_A_j8rDyhVM4_0(.din(n35622), .dout(n35625));
    jdff dff_A_ISuhW5kz7_0(.din(n35619), .dout(n35622));
    jdff dff_A_jYnAtpYq3_0(.din(n35616), .dout(n35619));
    jdff dff_A_K9dQJapv8_0(.din(n35613), .dout(n35616));
    jdff dff_A_PFmNnG3k8_0(.din(n35610), .dout(n35613));
    jdff dff_A_DggnEZFj7_0(.din(n35607), .dout(n35610));
    jdff dff_A_RbZnFsIQ5_0(.din(n35604), .dout(n35607));
    jdff dff_A_uzrl6ITp3_0(.din(n35601), .dout(n35604));
    jdff dff_A_wX4PHBXr0_0(.din(n35598), .dout(n35601));
    jdff dff_A_Xouw1Ph47_0(.din(n35595), .dout(n35598));
    jdff dff_A_3LVBNeEx3_0(.din(n35592), .dout(n35595));
    jdff dff_A_obuUdNIl2_2(.din(n4547), .dout(n35592));
    jdff dff_A_K0VMRFxq2_0(.din(n35586), .dout(G6160gat));
    jdff dff_A_bPuLvC5u3_0(.din(n35583), .dout(n35586));
    jdff dff_A_VvnvkjsB7_0(.din(n35580), .dout(n35583));
    jdff dff_A_VrkgbPSv9_0(.din(n35577), .dout(n35580));
    jdff dff_A_9aIz1G115_0(.din(n35574), .dout(n35577));
    jdff dff_A_kiSBccT21_0(.din(n35571), .dout(n35574));
    jdff dff_A_aPx83fBB0_0(.din(n35568), .dout(n35571));
    jdff dff_A_tLXdZOYV8_0(.din(n35565), .dout(n35568));
    jdff dff_A_ChMB0Ynx5_0(.din(n35562), .dout(n35565));
    jdff dff_A_JYl2zW550_0(.din(n35559), .dout(n35562));
    jdff dff_A_diXooZ1c8_0(.din(n35556), .dout(n35559));
    jdff dff_A_XyVUbH8F1_0(.din(n35553), .dout(n35556));
    jdff dff_A_tCRfYsDX5_0(.din(n35550), .dout(n35553));
    jdff dff_A_KiciQbBH1_0(.din(n35547), .dout(n35550));
    jdff dff_A_NKLITBXP5_0(.din(n35544), .dout(n35547));
    jdff dff_A_NEEFFIV93_0(.din(n35541), .dout(n35544));
    jdff dff_A_oYaKYWwJ3_0(.din(n35538), .dout(n35541));
    jdff dff_A_mBkmDaAr7_0(.din(n35535), .dout(n35538));
    jdff dff_A_rYofgzWO9_0(.din(n35532), .dout(n35535));
    jdff dff_A_ryMO8kaz0_0(.din(n35529), .dout(n35532));
    jdff dff_A_OSQHFrAg1_0(.din(n35526), .dout(n35529));
    jdff dff_A_oppvS8j14_0(.din(n35523), .dout(n35526));
    jdff dff_A_LVL9bFe91_0(.din(n35520), .dout(n35523));
    jdff dff_A_4CLg10dh8_0(.din(n35517), .dout(n35520));
    jdff dff_A_FMBJe05O9_0(.din(n35514), .dout(n35517));
    jdff dff_A_fgq1tWlH0_2(.din(n4176), .dout(n35514));
    jdff dff_A_5SPcpRbO5_0(.din(n35508), .dout(G6150gat));
    jdff dff_A_kQnOLAU39_0(.din(n35505), .dout(n35508));
    jdff dff_A_Y7CuQ6JA8_0(.din(n35502), .dout(n35505));
    jdff dff_A_2l8yetws1_0(.din(n35499), .dout(n35502));
    jdff dff_A_Mig4cTnu4_0(.din(n35496), .dout(n35499));
    jdff dff_A_c2YqTHKU9_0(.din(n35493), .dout(n35496));
    jdff dff_A_mjBcYgBA6_0(.din(n35490), .dout(n35493));
    jdff dff_A_1gZyF6l89_0(.din(n35487), .dout(n35490));
    jdff dff_A_6tTqPnQr9_0(.din(n35484), .dout(n35487));
    jdff dff_A_BZaa3w2n4_0(.din(n35481), .dout(n35484));
    jdff dff_A_Po2kMWjL0_0(.din(n35478), .dout(n35481));
    jdff dff_A_8ywlq8QD5_0(.din(n35475), .dout(n35478));
    jdff dff_A_q04g2wjQ5_0(.din(n35472), .dout(n35475));
    jdff dff_A_w2Cxhf6o2_0(.din(n35469), .dout(n35472));
    jdff dff_A_gp0tKW2z2_0(.din(n35466), .dout(n35469));
    jdff dff_A_vSa1ery42_0(.din(n35463), .dout(n35466));
    jdff dff_A_YVwbXvNp5_0(.din(n35460), .dout(n35463));
    jdff dff_A_p3wQVyqS2_0(.din(n35457), .dout(n35460));
    jdff dff_A_v22zptni0_0(.din(n35454), .dout(n35457));
    jdff dff_A_ELBK5l5c3_0(.din(n35451), .dout(n35454));
    jdff dff_A_zwZK5P7g3_0(.din(n35448), .dout(n35451));
    jdff dff_A_OSRhVY1y6_0(.din(n35445), .dout(n35448));
    jdff dff_A_2pjyHanq4_0(.din(n35442), .dout(n35445));
    jdff dff_A_79cZBL3i4_0(.din(n35439), .dout(n35442));
    jdff dff_A_wzQDPlfJ8_0(.din(n35436), .dout(n35439));
    jdff dff_A_gJhzoAqT4_0(.din(n35433), .dout(n35436));
    jdff dff_A_dFa2grTs5_0(.din(n35430), .dout(n35433));
    jdff dff_A_GkoBMSiy7_2(.din(n3774), .dout(n35430));
    jdff dff_A_fvjl21Pj0_0(.din(n35424), .dout(G6123gat));
    jdff dff_A_slTLL1i85_0(.din(n35421), .dout(n35424));
    jdff dff_A_UG3LSBeI9_0(.din(n35418), .dout(n35421));
    jdff dff_A_ALOEaoHQ2_0(.din(n35415), .dout(n35418));
    jdff dff_A_RqIx8HCk4_0(.din(n35412), .dout(n35415));
    jdff dff_A_G9Hukp1N3_0(.din(n35409), .dout(n35412));
    jdff dff_A_wW8DdkE31_0(.din(n35406), .dout(n35409));
    jdff dff_A_RIzwbEFv3_0(.din(n35403), .dout(n35406));
    jdff dff_A_QPJq0wl87_0(.din(n35400), .dout(n35403));
    jdff dff_A_4uVDk40k9_0(.din(n35397), .dout(n35400));
    jdff dff_A_Mo48ahrG7_0(.din(n35394), .dout(n35397));
    jdff dff_A_wBb23zsF9_0(.din(n35391), .dout(n35394));
    jdff dff_A_4bLZjiLN2_0(.din(n35388), .dout(n35391));
    jdff dff_A_eUEtAQCo4_0(.din(n35385), .dout(n35388));
    jdff dff_A_O2DG3k1q4_0(.din(n35382), .dout(n35385));
    jdff dff_A_4c4B0fIt5_0(.din(n35379), .dout(n35382));
    jdff dff_A_jMGqfSc36_0(.din(n35376), .dout(n35379));
    jdff dff_A_ChGizsMB3_0(.din(n35373), .dout(n35376));
    jdff dff_A_ExpXmqPP2_0(.din(n35370), .dout(n35373));
    jdff dff_A_IjeC78Q92_0(.din(n35367), .dout(n35370));
    jdff dff_A_aWMd9Avm2_0(.din(n35364), .dout(n35367));
    jdff dff_A_sxEwDzW34_0(.din(n35361), .dout(n35364));
    jdff dff_A_XaxNQUaZ9_0(.din(n35358), .dout(n35361));
    jdff dff_A_xiSZTgnd1_0(.din(n35355), .dout(n35358));
    jdff dff_A_CkGOUhHZ3_0(.din(n35352), .dout(n35355));
    jdff dff_A_13jcXOoq3_0(.din(n35349), .dout(n35352));
    jdff dff_A_WFPPUgIw0_0(.din(n35346), .dout(n35349));
    jdff dff_A_YArGBafw5_0(.din(n35343), .dout(n35346));
    jdff dff_A_tTAugpDu8_0(.din(n35340), .dout(n35343));
    jdff dff_A_NtHJwKOW4_2(.din(n3373), .dout(n35340));
    jdff dff_A_7zApRyyX4_0(.din(n35334), .dout(G5971gat));
    jdff dff_A_BwrTxgv56_0(.din(n35331), .dout(n35334));
    jdff dff_A_fD7qzMXK6_0(.din(n35328), .dout(n35331));
    jdff dff_A_yhb5xtMo9_0(.din(n35325), .dout(n35328));
    jdff dff_A_hBHHZSBk0_0(.din(n35322), .dout(n35325));
    jdff dff_A_49v8goCE1_0(.din(n35319), .dout(n35322));
    jdff dff_A_Q7ZELAT24_0(.din(n35316), .dout(n35319));
    jdff dff_A_FxLDEICg3_0(.din(n35313), .dout(n35316));
    jdff dff_A_KIrgp2FT9_0(.din(n35310), .dout(n35313));
    jdff dff_A_6ri971VA8_0(.din(n35307), .dout(n35310));
    jdff dff_A_1MceHRts7_0(.din(n35304), .dout(n35307));
    jdff dff_A_TkTttgAE7_0(.din(n35301), .dout(n35304));
    jdff dff_A_tDwSXBuX8_0(.din(n35298), .dout(n35301));
    jdff dff_A_kNbLuFPy1_0(.din(n35295), .dout(n35298));
    jdff dff_A_fJ2ksThq7_0(.din(n35292), .dout(n35295));
    jdff dff_A_seMU5cwB7_0(.din(n35289), .dout(n35292));
    jdff dff_A_ctOe0XbO7_0(.din(n35286), .dout(n35289));
    jdff dff_A_QGzY2HHp8_0(.din(n35283), .dout(n35286));
    jdff dff_A_uO5GxKNN4_0(.din(n35280), .dout(n35283));
    jdff dff_A_3vS5ofQE4_0(.din(n35277), .dout(n35280));
    jdff dff_A_a6yGjMhT8_0(.din(n35274), .dout(n35277));
    jdff dff_A_4oxaVBo92_0(.din(n35271), .dout(n35274));
    jdff dff_A_DlEzE1mQ8_0(.din(n35268), .dout(n35271));
    jdff dff_A_64uUHRJo8_0(.din(n35265), .dout(n35268));
    jdff dff_A_uNvo4nFD0_0(.din(n35262), .dout(n35265));
    jdff dff_A_6luKBhuP9_0(.din(n35259), .dout(n35262));
    jdff dff_A_iSE9KQJO4_0(.din(n35256), .dout(n35259));
    jdff dff_A_dCcWln6m4_0(.din(n35253), .dout(n35256));
    jdff dff_A_UD61nGIn5_0(.din(n35250), .dout(n35253));
    jdff dff_A_noM0juy98_0(.din(n35247), .dout(n35250));
    jdff dff_A_ZoFID5zg1_0(.din(n35244), .dout(n35247));
    jdff dff_A_rnAfQz647_0(.din(n35241), .dout(n35244));
    jdff dff_A_ND5rrPHV5_2(.din(n2971), .dout(n35241));
    jdff dff_A_miMC25NO6_0(.din(n35235), .dout(G5672gat));
    jdff dff_A_ezVCfewI6_0(.din(n35232), .dout(n35235));
    jdff dff_A_lBGpUiJc3_0(.din(n35229), .dout(n35232));
    jdff dff_A_Vx8PwlVK2_0(.din(n35226), .dout(n35229));
    jdff dff_A_TiehvIPe1_0(.din(n35223), .dout(n35226));
    jdff dff_A_raTQam683_0(.din(n35220), .dout(n35223));
    jdff dff_A_Ltom9Con4_0(.din(n35217), .dout(n35220));
    jdff dff_A_r43YaIL49_0(.din(n35214), .dout(n35217));
    jdff dff_A_kBXQzIa09_0(.din(n35211), .dout(n35214));
    jdff dff_A_SVNBHzQj6_0(.din(n35208), .dout(n35211));
    jdff dff_A_F6jGdstK4_0(.din(n35205), .dout(n35208));
    jdff dff_A_lsm4iIuD7_0(.din(n35202), .dout(n35205));
    jdff dff_A_0XnJtovy0_0(.din(n35199), .dout(n35202));
    jdff dff_A_brPQUTpK2_0(.din(n35196), .dout(n35199));
    jdff dff_A_s2yProDA8_0(.din(n35193), .dout(n35196));
    jdff dff_A_ac4B31Zm5_0(.din(n35190), .dout(n35193));
    jdff dff_A_D50d9q789_0(.din(n35187), .dout(n35190));
    jdff dff_A_AiBYpJBN9_0(.din(n35184), .dout(n35187));
    jdff dff_A_NqdZPWQn1_0(.din(n35181), .dout(n35184));
    jdff dff_A_24sZSyuT2_0(.din(n35178), .dout(n35181));
    jdff dff_A_gqh9o9Uh4_0(.din(n35175), .dout(n35178));
    jdff dff_A_vKxdlqmx2_0(.din(n35172), .dout(n35175));
    jdff dff_A_8cLKzRYr0_0(.din(n35169), .dout(n35172));
    jdff dff_A_UINZN4gY4_0(.din(n35166), .dout(n35169));
    jdff dff_A_uzU0o8xR2_0(.din(n35163), .dout(n35166));
    jdff dff_A_hhlbElyG8_0(.din(n35160), .dout(n35163));
    jdff dff_A_2RppvQGd1_0(.din(n35157), .dout(n35160));
    jdff dff_A_LPRA2KEJ1_0(.din(n35154), .dout(n35157));
    jdff dff_A_AhKosuqg5_0(.din(n35151), .dout(n35154));
    jdff dff_A_9IUh5jR18_0(.din(n35148), .dout(n35151));
    jdff dff_A_hUJ43Mx16_0(.din(n35145), .dout(n35148));
    jdff dff_A_k3IAA0DQ1_0(.din(n35142), .dout(n35145));
    jdff dff_A_LEiV6ZbY0_0(.din(n35139), .dout(n35142));
    jdff dff_A_EeD76MjA9_0(.din(n35136), .dout(n35139));
    jdff dff_A_5mbaOIAJ7_0(.din(n35133), .dout(n35136));
    jdff dff_A_TEKx8qT56_2(.din(n2589), .dout(n35133));
    jdff dff_A_SCqH8zVk4_0(.din(n35127), .dout(G5308gat));
    jdff dff_A_LQ7uLL3z4_0(.din(n35124), .dout(n35127));
    jdff dff_A_xvKm44JZ0_0(.din(n35121), .dout(n35124));
    jdff dff_A_2AMhb9GJ6_0(.din(n35118), .dout(n35121));
    jdff dff_A_6Sybiw3c3_0(.din(n35115), .dout(n35118));
    jdff dff_A_wjoisF5K4_0(.din(n35112), .dout(n35115));
    jdff dff_A_1OqLBf1z9_0(.din(n35109), .dout(n35112));
    jdff dff_A_u3M4koVj4_0(.din(n35106), .dout(n35109));
    jdff dff_A_vROip8wM3_0(.din(n35103), .dout(n35106));
    jdff dff_A_Yh73tfam1_0(.din(n35100), .dout(n35103));
    jdff dff_A_Vb4wSG9j9_0(.din(n35097), .dout(n35100));
    jdff dff_A_3yAZ8lbo1_0(.din(n35094), .dout(n35097));
    jdff dff_A_Avkw0D2G0_0(.din(n35091), .dout(n35094));
    jdff dff_A_xDZBgepc1_0(.din(n35088), .dout(n35091));
    jdff dff_A_TUn1Bpxd1_0(.din(n35085), .dout(n35088));
    jdff dff_A_y09MRX6l3_0(.din(n35082), .dout(n35085));
    jdff dff_A_hxDU4T4v5_0(.din(n35079), .dout(n35082));
    jdff dff_A_R70apvjg6_0(.din(n35076), .dout(n35079));
    jdff dff_A_oJXbKlhp9_0(.din(n35073), .dout(n35076));
    jdff dff_A_cEGfUJgl3_0(.din(n35070), .dout(n35073));
    jdff dff_A_AUUizrVk3_0(.din(n35067), .dout(n35070));
    jdff dff_A_18ITMQEf6_0(.din(n35064), .dout(n35067));
    jdff dff_A_My7pE2MQ1_0(.din(n35061), .dout(n35064));
    jdff dff_A_LMHMNP2S0_0(.din(n35058), .dout(n35061));
    jdff dff_A_qFMdeTVf4_0(.din(n35055), .dout(n35058));
    jdff dff_A_AgMpUUJg0_0(.din(n35052), .dout(n35055));
    jdff dff_A_2fBCdJA41_0(.din(n35049), .dout(n35052));
    jdff dff_A_lWMirraW9_0(.din(n35046), .dout(n35049));
    jdff dff_A_TC6LzhCv1_0(.din(n35043), .dout(n35046));
    jdff dff_A_jgqmBM7u3_0(.din(n35040), .dout(n35043));
    jdff dff_A_p2BWwzJt9_0(.din(n35037), .dout(n35040));
    jdff dff_A_0Uc7yspJ2_0(.din(n35034), .dout(n35037));
    jdff dff_A_UKQhSSBv1_0(.din(n35031), .dout(n35034));
    jdff dff_A_6Zc0b0fZ8_0(.din(n35028), .dout(n35031));
    jdff dff_A_gxl8MQ4C1_0(.din(n35025), .dout(n35028));
    jdff dff_A_96qz8p685_0(.din(n35022), .dout(n35025));
    jdff dff_A_lSs1vlGz9_0(.din(n35019), .dout(n35022));
    jdff dff_A_rBGM1luv2_0(.din(n35016), .dout(n35019));
    jdff dff_A_7vyaZLbT9_2(.din(n2234), .dout(n35016));
    jdff dff_A_xgDN7rc03_0(.din(n35010), .dout(G4946gat));
    jdff dff_A_sGerDx5E0_0(.din(n35007), .dout(n35010));
    jdff dff_A_HbMaSnJb1_0(.din(n35004), .dout(n35007));
    jdff dff_A_jBG6z9Zz6_0(.din(n35001), .dout(n35004));
    jdff dff_A_dRqHU3vM2_0(.din(n34998), .dout(n35001));
    jdff dff_A_bc52apDh2_0(.din(n34995), .dout(n34998));
    jdff dff_A_kVagMUbd2_0(.din(n34992), .dout(n34995));
    jdff dff_A_BMI7anqQ5_0(.din(n34989), .dout(n34992));
    jdff dff_A_iMAxdH4P7_0(.din(n34986), .dout(n34989));
    jdff dff_A_YKM56Nk35_0(.din(n34983), .dout(n34986));
    jdff dff_A_9BaNkW873_0(.din(n34980), .dout(n34983));
    jdff dff_A_2GQKVBUa4_0(.din(n34977), .dout(n34980));
    jdff dff_A_2Bc3iSTU2_0(.din(n34974), .dout(n34977));
    jdff dff_A_9dQXlluI7_0(.din(n34971), .dout(n34974));
    jdff dff_A_PlGwnbl21_0(.din(n34968), .dout(n34971));
    jdff dff_A_5R1Urcqo2_0(.din(n34965), .dout(n34968));
    jdff dff_A_PhBFujKQ8_0(.din(n34962), .dout(n34965));
    jdff dff_A_TxihdmPS3_0(.din(n34959), .dout(n34962));
    jdff dff_A_38nBbQo59_0(.din(n34956), .dout(n34959));
    jdff dff_A_1FU2AFeo8_0(.din(n34953), .dout(n34956));
    jdff dff_A_hgW0cZ6R3_0(.din(n34950), .dout(n34953));
    jdff dff_A_0yEshw0C5_0(.din(n34947), .dout(n34950));
    jdff dff_A_AxWT3cyQ6_0(.din(n34944), .dout(n34947));
    jdff dff_A_HBs1nnTQ8_0(.din(n34941), .dout(n34944));
    jdff dff_A_bMRb5fEI9_0(.din(n34938), .dout(n34941));
    jdff dff_A_KvAm47Gq4_0(.din(n34935), .dout(n34938));
    jdff dff_A_BNP7UCab2_0(.din(n34932), .dout(n34935));
    jdff dff_A_CnZPTTrA1_0(.din(n34929), .dout(n34932));
    jdff dff_A_NiH8YMgt1_0(.din(n34926), .dout(n34929));
    jdff dff_A_DeGW5AQc1_0(.din(n34923), .dout(n34926));
    jdff dff_A_2kzbZG6l7_0(.din(n34920), .dout(n34923));
    jdff dff_A_EWuIz2Yi1_0(.din(n34917), .dout(n34920));
    jdff dff_A_AdqfIWAB0_0(.din(n34914), .dout(n34917));
    jdff dff_A_u2lVkaxh5_0(.din(n34911), .dout(n34914));
    jdff dff_A_HYP6mTaq8_0(.din(n34908), .dout(n34911));
    jdff dff_A_m8vhnz8X6_0(.din(n34905), .dout(n34908));
    jdff dff_A_4IEEwk6D1_0(.din(n34902), .dout(n34905));
    jdff dff_A_bXFsMF1j7_0(.din(n34899), .dout(n34902));
    jdff dff_A_4Z7Lme3u0_0(.din(n34896), .dout(n34899));
    jdff dff_A_8isAp7KB2_0(.din(n34893), .dout(n34896));
    jdff dff_A_4ZUMfstK2_0(.din(n34890), .dout(n34893));
    jdff dff_A_x2APV6JE4_2(.din(n1906), .dout(n34890));
    jdff dff_A_H8sTOo013_0(.din(n34884), .dout(G4591gat));
    jdff dff_A_vsJcTJdJ4_0(.din(n34881), .dout(n34884));
    jdff dff_A_YmCBS2ot5_0(.din(n34878), .dout(n34881));
    jdff dff_A_9jyakfJn9_0(.din(n34875), .dout(n34878));
    jdff dff_A_zsMZny7A9_0(.din(n34872), .dout(n34875));
    jdff dff_A_J86AyhRy1_0(.din(n34869), .dout(n34872));
    jdff dff_A_moRygh1K1_0(.din(n34866), .dout(n34869));
    jdff dff_A_Oa3dy7Jx0_0(.din(n34863), .dout(n34866));
    jdff dff_A_nhjQHZwh3_0(.din(n34860), .dout(n34863));
    jdff dff_A_o8iwBowI6_0(.din(n34857), .dout(n34860));
    jdff dff_A_MnTObEKb6_0(.din(n34854), .dout(n34857));
    jdff dff_A_85U7jzTf1_0(.din(n34851), .dout(n34854));
    jdff dff_A_6XOZBCHi0_0(.din(n34848), .dout(n34851));
    jdff dff_A_7XI49bBE6_0(.din(n34845), .dout(n34848));
    jdff dff_A_PuXQpVOz3_0(.din(n34842), .dout(n34845));
    jdff dff_A_QJEE8DWm4_0(.din(n34839), .dout(n34842));
    jdff dff_A_jNyxx1wT6_0(.din(n34836), .dout(n34839));
    jdff dff_A_3tX2e9C44_0(.din(n34833), .dout(n34836));
    jdff dff_A_hE0m3T3e9_0(.din(n34830), .dout(n34833));
    jdff dff_A_GoxV6nt89_0(.din(n34827), .dout(n34830));
    jdff dff_A_EPf5hEiT1_0(.din(n34824), .dout(n34827));
    jdff dff_A_PZD3Cajo7_0(.din(n34821), .dout(n34824));
    jdff dff_A_iuQwrsgM3_0(.din(n34818), .dout(n34821));
    jdff dff_A_GpRypKlf2_0(.din(n34815), .dout(n34818));
    jdff dff_A_0de3tUVL0_0(.din(n34812), .dout(n34815));
    jdff dff_A_Vy2WT7NC9_0(.din(n34809), .dout(n34812));
    jdff dff_A_TShY5e1Z7_0(.din(n34806), .dout(n34809));
    jdff dff_A_0JAzP6X92_0(.din(n34803), .dout(n34806));
    jdff dff_A_cTZlejHs1_0(.din(n34800), .dout(n34803));
    jdff dff_A_nGGdf9zh1_0(.din(n34797), .dout(n34800));
    jdff dff_A_xEF2irEO8_0(.din(n34794), .dout(n34797));
    jdff dff_A_MVtKYeAe9_0(.din(n34791), .dout(n34794));
    jdff dff_A_FB2kpki42_0(.din(n34788), .dout(n34791));
    jdff dff_A_LUg8UohJ2_0(.din(n34785), .dout(n34788));
    jdff dff_A_ngcDbCQN1_0(.din(n34782), .dout(n34785));
    jdff dff_A_KNsYc6qM1_0(.din(n34779), .dout(n34782));
    jdff dff_A_YpfIfAzr6_0(.din(n34776), .dout(n34779));
    jdff dff_A_9aQLkix55_0(.din(n34773), .dout(n34776));
    jdff dff_A_DUTLKYQL6_0(.din(n34770), .dout(n34773));
    jdff dff_A_Llfmmfo59_0(.din(n34767), .dout(n34770));
    jdff dff_A_Y84AA9ZC1_0(.din(n34764), .dout(n34767));
    jdff dff_A_q4LRSY5y5_0(.din(n34761), .dout(n34764));
    jdff dff_A_iiBkQspR7_0(.din(n34758), .dout(n34761));
    jdff dff_A_mR2Eva228_0(.din(n34755), .dout(n34758));
    jdff dff_A_Phb6U75D9_2(.din(n1605), .dout(n34755));
    jdff dff_A_UElGlsnx8_0(.din(n34749), .dout(G4241gat));
    jdff dff_A_TD0rCCw76_0(.din(n34746), .dout(n34749));
    jdff dff_A_kGMURzPc5_0(.din(n34743), .dout(n34746));
    jdff dff_A_BCvXb6co5_0(.din(n34740), .dout(n34743));
    jdff dff_A_d0TPnhfP7_0(.din(n34737), .dout(n34740));
    jdff dff_A_qc3faVvK6_0(.din(n34734), .dout(n34737));
    jdff dff_A_6c2Zg5Hw8_0(.din(n34731), .dout(n34734));
    jdff dff_A_SjRZRti05_0(.din(n34728), .dout(n34731));
    jdff dff_A_O50fT2260_0(.din(n34725), .dout(n34728));
    jdff dff_A_rIywPZc71_0(.din(n34722), .dout(n34725));
    jdff dff_A_PAynWK271_0(.din(n34719), .dout(n34722));
    jdff dff_A_C06t6JTJ2_0(.din(n34716), .dout(n34719));
    jdff dff_A_EsM5A4XG5_0(.din(n34713), .dout(n34716));
    jdff dff_A_UFeWtC3S0_0(.din(n34710), .dout(n34713));
    jdff dff_A_p3iF3YJn8_0(.din(n34707), .dout(n34710));
    jdff dff_A_YJElB5c46_0(.din(n34704), .dout(n34707));
    jdff dff_A_yfka91WD1_0(.din(n34701), .dout(n34704));
    jdff dff_A_w6tNTT3C9_0(.din(n34698), .dout(n34701));
    jdff dff_A_zsBQAZrm8_0(.din(n34695), .dout(n34698));
    jdff dff_A_EKThDx0b3_0(.din(n34692), .dout(n34695));
    jdff dff_A_gS7FByvC2_0(.din(n34689), .dout(n34692));
    jdff dff_A_ZWZPEdqW4_0(.din(n34686), .dout(n34689));
    jdff dff_A_VdZlvEUK6_0(.din(n34683), .dout(n34686));
    jdff dff_A_C4PI9ZpR7_0(.din(n34680), .dout(n34683));
    jdff dff_A_mPavfK0m8_0(.din(n34677), .dout(n34680));
    jdff dff_A_E2RjHl9D8_0(.din(n34674), .dout(n34677));
    jdff dff_A_kkd0xx6G5_0(.din(n34671), .dout(n34674));
    jdff dff_A_J6LhkjTI5_0(.din(n34668), .dout(n34671));
    jdff dff_A_kdfXz4xG5_0(.din(n34665), .dout(n34668));
    jdff dff_A_3U3ruLjg7_0(.din(n34662), .dout(n34665));
    jdff dff_A_v1cz1S526_0(.din(n34659), .dout(n34662));
    jdff dff_A_FjyxqxJR5_0(.din(n34656), .dout(n34659));
    jdff dff_A_JMBMXPot0_0(.din(n34653), .dout(n34656));
    jdff dff_A_TFdvfNZE4_0(.din(n34650), .dout(n34653));
    jdff dff_A_ewKztJgs5_0(.din(n34647), .dout(n34650));
    jdff dff_A_5rDcnqKM0_0(.din(n34644), .dout(n34647));
    jdff dff_A_SDwRpmoh6_0(.din(n34641), .dout(n34644));
    jdff dff_A_apc6Yn0R8_0(.din(n34638), .dout(n34641));
    jdff dff_A_EEAvtlMp8_0(.din(n34635), .dout(n34638));
    jdff dff_A_Ytk9gg1e7_0(.din(n34632), .dout(n34635));
    jdff dff_A_lNjD4OkO5_0(.din(n34629), .dout(n34632));
    jdff dff_A_ErXFPDHr2_0(.din(n34626), .dout(n34629));
    jdff dff_A_j0fwaono3_0(.din(n34623), .dout(n34626));
    jdff dff_A_RD4HbXrN3_0(.din(n34620), .dout(n34623));
    jdff dff_A_2Q16xPir4_0(.din(n34617), .dout(n34620));
    jdff dff_A_8wzFp3Rz4_0(.din(n34614), .dout(n34617));
    jdff dff_A_ucXRuTTy6_0(.din(n34611), .dout(n34614));
    jdff dff_A_mdcJ4ar90_2(.din(n1331), .dout(n34611));
    jdff dff_A_G853ioWQ5_0(.din(n34605), .dout(G3895gat));
    jdff dff_A_hZpcWkUB7_0(.din(n34602), .dout(n34605));
    jdff dff_A_WPod74vA5_0(.din(n34599), .dout(n34602));
    jdff dff_A_QGDy6GMk4_0(.din(n34596), .dout(n34599));
    jdff dff_A_5tWePsnQ5_0(.din(n34593), .dout(n34596));
    jdff dff_A_1I2yB0dQ3_0(.din(n34590), .dout(n34593));
    jdff dff_A_uUTRxxwB7_0(.din(n34587), .dout(n34590));
    jdff dff_A_d8ZKm9L55_0(.din(n34584), .dout(n34587));
    jdff dff_A_v1wARnUV7_0(.din(n34581), .dout(n34584));
    jdff dff_A_vGZPtRr95_0(.din(n34578), .dout(n34581));
    jdff dff_A_iWyeoXsu8_0(.din(n34575), .dout(n34578));
    jdff dff_A_GJiTmOg07_0(.din(n34572), .dout(n34575));
    jdff dff_A_8xKbKkRf2_0(.din(n34569), .dout(n34572));
    jdff dff_A_GCTuFQdP2_0(.din(n34566), .dout(n34569));
    jdff dff_A_97w0fdhi5_0(.din(n34563), .dout(n34566));
    jdff dff_A_UyEANOgG7_0(.din(n34560), .dout(n34563));
    jdff dff_A_PCqNBvVU8_0(.din(n34557), .dout(n34560));
    jdff dff_A_cHyQKoF31_0(.din(n34554), .dout(n34557));
    jdff dff_A_7SpiseeD3_0(.din(n34551), .dout(n34554));
    jdff dff_A_9LJ5SVdU0_0(.din(n34548), .dout(n34551));
    jdff dff_A_bMyFap6R8_0(.din(n34545), .dout(n34548));
    jdff dff_A_u5lQ2RIG2_0(.din(n34542), .dout(n34545));
    jdff dff_A_fVChj8QF5_0(.din(n34539), .dout(n34542));
    jdff dff_A_WO0q5qOl7_0(.din(n34536), .dout(n34539));
    jdff dff_A_uwXDEM0t8_0(.din(n34533), .dout(n34536));
    jdff dff_A_T1zyELv61_0(.din(n34530), .dout(n34533));
    jdff dff_A_FiLwcXha9_0(.din(n34527), .dout(n34530));
    jdff dff_A_jcMpPvlb7_0(.din(n34524), .dout(n34527));
    jdff dff_A_OxNPGvac0_0(.din(n34521), .dout(n34524));
    jdff dff_A_79dKQcCA6_0(.din(n34518), .dout(n34521));
    jdff dff_A_yzWhyFCM4_0(.din(n34515), .dout(n34518));
    jdff dff_A_6ljpBP196_0(.din(n34512), .dout(n34515));
    jdff dff_A_IIaFWszV3_0(.din(n34509), .dout(n34512));
    jdff dff_A_QSNsEGjp8_0(.din(n34506), .dout(n34509));
    jdff dff_A_Hx307nNz5_0(.din(n34503), .dout(n34506));
    jdff dff_A_MNG0GSFM8_0(.din(n34500), .dout(n34503));
    jdff dff_A_WIJih7lt7_0(.din(n34497), .dout(n34500));
    jdff dff_A_KWfWl4Vb3_0(.din(n34494), .dout(n34497));
    jdff dff_A_rnXu5VpJ8_0(.din(n34491), .dout(n34494));
    jdff dff_A_7wu4IHuK6_0(.din(n34488), .dout(n34491));
    jdff dff_A_Bblxg0SQ5_0(.din(n34485), .dout(n34488));
    jdff dff_A_mRhjIvPZ4_0(.din(n34482), .dout(n34485));
    jdff dff_A_vlL9DLbv4_0(.din(n34479), .dout(n34482));
    jdff dff_A_d3KWg11b4_0(.din(n34476), .dout(n34479));
    jdff dff_A_qAgfKp1R4_0(.din(n34473), .dout(n34476));
    jdff dff_A_5J3Q3rFA6_0(.din(n34470), .dout(n34473));
    jdff dff_A_5YmVidb34_0(.din(n34467), .dout(n34470));
    jdff dff_A_3vcoTw601_0(.din(n34464), .dout(n34467));
    jdff dff_A_JAUFx1H55_0(.din(n34461), .dout(n34464));
    jdff dff_A_gZhCNXNw1_0(.din(n34458), .dout(n34461));
    jdff dff_A_8gCK9mkA1_2(.din(n1087), .dout(n34458));
    jdff dff_A_E6Tczljx8_0(.din(n34452), .dout(G3552gat));
    jdff dff_A_XFF46Scq2_0(.din(n34449), .dout(n34452));
    jdff dff_A_e41qEz0N0_0(.din(n34446), .dout(n34449));
    jdff dff_A_tGZYoIwU7_0(.din(n34443), .dout(n34446));
    jdff dff_A_YDg62S291_0(.din(n34440), .dout(n34443));
    jdff dff_A_vBxmA6LB5_0(.din(n34437), .dout(n34440));
    jdff dff_A_PrqbpDdw6_0(.din(n34434), .dout(n34437));
    jdff dff_A_NWFLROeL9_0(.din(n34431), .dout(n34434));
    jdff dff_A_0CHITjur6_0(.din(n34428), .dout(n34431));
    jdff dff_A_DyDEiMTR9_0(.din(n34425), .dout(n34428));
    jdff dff_A_AABDCGJa1_0(.din(n34422), .dout(n34425));
    jdff dff_A_NEVy6wJg0_0(.din(n34419), .dout(n34422));
    jdff dff_A_0bmlHtoQ2_0(.din(n34416), .dout(n34419));
    jdff dff_A_Clh6yr2s4_0(.din(n34413), .dout(n34416));
    jdff dff_A_pwjGtfFN2_0(.din(n34410), .dout(n34413));
    jdff dff_A_5TP7WeBX6_0(.din(n34407), .dout(n34410));
    jdff dff_A_KpCWsgbB6_0(.din(n34404), .dout(n34407));
    jdff dff_A_nNAihJVP2_0(.din(n34401), .dout(n34404));
    jdff dff_A_rYLWwpsi5_0(.din(n34398), .dout(n34401));
    jdff dff_A_gUA9l13G5_0(.din(n34395), .dout(n34398));
    jdff dff_A_ZKRWuKQ48_0(.din(n34392), .dout(n34395));
    jdff dff_A_BglbO1Nb1_0(.din(n34389), .dout(n34392));
    jdff dff_A_bW12ClKR0_0(.din(n34386), .dout(n34389));
    jdff dff_A_9iXITTRO2_0(.din(n34383), .dout(n34386));
    jdff dff_A_oqXMtO5e1_0(.din(n34380), .dout(n34383));
    jdff dff_A_MbeVzEdF9_0(.din(n34377), .dout(n34380));
    jdff dff_A_9nAAV3iw0_0(.din(n34374), .dout(n34377));
    jdff dff_A_rfVEkmun7_0(.din(n34371), .dout(n34374));
    jdff dff_A_roPLPGKs4_0(.din(n34368), .dout(n34371));
    jdff dff_A_0yWtDODy3_0(.din(n34365), .dout(n34368));
    jdff dff_A_lecah2h29_0(.din(n34362), .dout(n34365));
    jdff dff_A_3mqbvP4W1_0(.din(n34359), .dout(n34362));
    jdff dff_A_AcMpOlLu9_0(.din(n34356), .dout(n34359));
    jdff dff_A_VHTLPc0a7_0(.din(n34353), .dout(n34356));
    jdff dff_A_AxcYoavu9_0(.din(n34350), .dout(n34353));
    jdff dff_A_BPh9lray7_0(.din(n34347), .dout(n34350));
    jdff dff_A_xgL3MgNv9_0(.din(n34344), .dout(n34347));
    jdff dff_A_R06KiJGO1_0(.din(n34341), .dout(n34344));
    jdff dff_A_IAEEHCxV1_0(.din(n34338), .dout(n34341));
    jdff dff_A_hmWynH6E1_0(.din(n34335), .dout(n34338));
    jdff dff_A_0Ej9uaVS9_0(.din(n34332), .dout(n34335));
    jdff dff_A_OU5mnSOI7_0(.din(n34329), .dout(n34332));
    jdff dff_A_vZkmqeXs2_0(.din(n34326), .dout(n34329));
    jdff dff_A_oijkPitJ0_0(.din(n34323), .dout(n34326));
    jdff dff_A_npqPB1Q28_0(.din(n34320), .dout(n34323));
    jdff dff_A_iWRwJXu99_0(.din(n34317), .dout(n34320));
    jdff dff_A_8teEXTp34_0(.din(n34314), .dout(n34317));
    jdff dff_A_n8Qrp2Vw8_0(.din(n34311), .dout(n34314));
    jdff dff_A_LOY1HQbs4_0(.din(n34308), .dout(n34311));
    jdff dff_A_Xxke3TNk9_0(.din(n34305), .dout(n34308));
    jdff dff_A_DQ4C7Sfr2_0(.din(n34302), .dout(n34305));
    jdff dff_A_ijtJorKs5_0(.din(n34299), .dout(n34302));
    jdff dff_A_k1paZK0Y2_0(.din(n34296), .dout(n34299));
    jdff dff_A_AWpHub178_2(.din(n867), .dout(n34296));
    jdff dff_A_yJ4EGLoz5_0(.din(n34290), .dout(G3211gat));
    jdff dff_A_1KEcECGy0_0(.din(n34287), .dout(n34290));
    jdff dff_A_XdntmXwb6_0(.din(n34284), .dout(n34287));
    jdff dff_A_2oBeUSdY0_0(.din(n34281), .dout(n34284));
    jdff dff_A_z29R41yA9_0(.din(n34278), .dout(n34281));
    jdff dff_A_XXBn1gv58_0(.din(n34275), .dout(n34278));
    jdff dff_A_qZ22fWx69_0(.din(n34272), .dout(n34275));
    jdff dff_A_BWCZocTP7_0(.din(n34269), .dout(n34272));
    jdff dff_A_DBTLQpSv1_0(.din(n34266), .dout(n34269));
    jdff dff_A_nagS59Gw5_0(.din(n34263), .dout(n34266));
    jdff dff_A_Y70DArRS4_0(.din(n34260), .dout(n34263));
    jdff dff_A_rPFu5ZpZ8_0(.din(n34257), .dout(n34260));
    jdff dff_A_KOXpkjoS4_0(.din(n34254), .dout(n34257));
    jdff dff_A_SuSjSHB70_0(.din(n34251), .dout(n34254));
    jdff dff_A_SPWjq15W3_0(.din(n34248), .dout(n34251));
    jdff dff_A_GD3P4vfF6_0(.din(n34245), .dout(n34248));
    jdff dff_A_MdjoMgUH1_0(.din(n34242), .dout(n34245));
    jdff dff_A_mGKEe4Tn7_0(.din(n34239), .dout(n34242));
    jdff dff_A_KQEBDqy60_0(.din(n34236), .dout(n34239));
    jdff dff_A_VVRS5WCw3_0(.din(n34233), .dout(n34236));
    jdff dff_A_V3mBh8Xe1_0(.din(n34230), .dout(n34233));
    jdff dff_A_h5UpJryP1_0(.din(n34227), .dout(n34230));
    jdff dff_A_urBqOGvO9_0(.din(n34224), .dout(n34227));
    jdff dff_A_lcAp889A4_0(.din(n34221), .dout(n34224));
    jdff dff_A_XhvDV9rF2_0(.din(n34218), .dout(n34221));
    jdff dff_A_P5Laq6MP6_0(.din(n34215), .dout(n34218));
    jdff dff_A_tZSNMhT42_0(.din(n34212), .dout(n34215));
    jdff dff_A_8aFoTaVN9_0(.din(n34209), .dout(n34212));
    jdff dff_A_TfhU36SW1_0(.din(n34206), .dout(n34209));
    jdff dff_A_IMY3fq3d2_0(.din(n34203), .dout(n34206));
    jdff dff_A_aWzaHUEc1_0(.din(n34200), .dout(n34203));
    jdff dff_A_4BGdnQu19_0(.din(n34197), .dout(n34200));
    jdff dff_A_cGlLDSgH2_0(.din(n34194), .dout(n34197));
    jdff dff_A_x75KIasX8_0(.din(n34191), .dout(n34194));
    jdff dff_A_Yf2eC9iE3_0(.din(n34188), .dout(n34191));
    jdff dff_A_QYU6znvH3_0(.din(n34185), .dout(n34188));
    jdff dff_A_wWCHn3aI2_0(.din(n34182), .dout(n34185));
    jdff dff_A_m3MsK69G3_0(.din(n34179), .dout(n34182));
    jdff dff_A_lv79t8RY6_0(.din(n34176), .dout(n34179));
    jdff dff_A_i55dgTbi1_0(.din(n34173), .dout(n34176));
    jdff dff_A_EIOYCWZT6_0(.din(n34170), .dout(n34173));
    jdff dff_A_dLTlhKMU5_0(.din(n34167), .dout(n34170));
    jdff dff_A_ET5BbgDx8_0(.din(n34164), .dout(n34167));
    jdff dff_A_z4swIlhP5_0(.din(n34161), .dout(n34164));
    jdff dff_A_RwzAJwkD4_0(.din(n34158), .dout(n34161));
    jdff dff_A_oZzv7tR73_0(.din(n34155), .dout(n34158));
    jdff dff_A_UIl9BgcD5_0(.din(n34152), .dout(n34155));
    jdff dff_A_SDcD5pXx9_0(.din(n34149), .dout(n34152));
    jdff dff_A_incpz5RR2_0(.din(n34146), .dout(n34149));
    jdff dff_A_d8LqlvIK9_0(.din(n34143), .dout(n34146));
    jdff dff_A_A4V818kf7_0(.din(n34140), .dout(n34143));
    jdff dff_A_zqHGa9GZ9_0(.din(n34137), .dout(n34140));
    jdff dff_A_Ixj4wH3s3_0(.din(n34134), .dout(n34137));
    jdff dff_A_sti6URCX3_0(.din(n34131), .dout(n34134));
    jdff dff_A_gbjDoEu50_0(.din(n34128), .dout(n34131));
    jdff dff_A_OeD4kmTb0_0(.din(n34125), .dout(n34128));
    jdff dff_A_3cNNDt623_2(.din(n674), .dout(n34125));
    jdff dff_A_XQpzOOFe4_0(.din(n34119), .dout(G2877gat));
    jdff dff_A_I9IweMtn6_0(.din(n34116), .dout(n34119));
    jdff dff_A_wn5HowOg8_0(.din(n34113), .dout(n34116));
    jdff dff_A_f4420IxB5_0(.din(n34110), .dout(n34113));
    jdff dff_A_fj6EaFpb0_0(.din(n34107), .dout(n34110));
    jdff dff_A_hsBftZC11_0(.din(n34104), .dout(n34107));
    jdff dff_A_3K3I5SLN9_0(.din(n34101), .dout(n34104));
    jdff dff_A_0kYKmnQE1_0(.din(n34098), .dout(n34101));
    jdff dff_A_hvHqZMJY9_0(.din(n34095), .dout(n34098));
    jdff dff_A_8MbgAvdt1_0(.din(n34092), .dout(n34095));
    jdff dff_A_jz5MI4T16_0(.din(n34089), .dout(n34092));
    jdff dff_A_IMUfPG2y2_0(.din(n34086), .dout(n34089));
    jdff dff_A_MD9CjD6p0_0(.din(n34083), .dout(n34086));
    jdff dff_A_xgSBFmNI2_0(.din(n34080), .dout(n34083));
    jdff dff_A_Np5uqXUX6_0(.din(n34077), .dout(n34080));
    jdff dff_A_bnRvhZUK2_0(.din(n34074), .dout(n34077));
    jdff dff_A_YIkkrbas4_0(.din(n34071), .dout(n34074));
    jdff dff_A_SH4AX4Fe8_0(.din(n34068), .dout(n34071));
    jdff dff_A_joOw27Ci1_0(.din(n34065), .dout(n34068));
    jdff dff_A_H0xHfJn59_0(.din(n34062), .dout(n34065));
    jdff dff_A_Rj33y8Qg2_0(.din(n34059), .dout(n34062));
    jdff dff_A_YKdDcgJM5_0(.din(n34056), .dout(n34059));
    jdff dff_A_uQOZSzyv7_0(.din(n34053), .dout(n34056));
    jdff dff_A_dn38EZaj9_0(.din(n34050), .dout(n34053));
    jdff dff_A_R9sSCIk98_0(.din(n34047), .dout(n34050));
    jdff dff_A_Czx8K6yD4_0(.din(n34044), .dout(n34047));
    jdff dff_A_XybjtclJ7_0(.din(n34041), .dout(n34044));
    jdff dff_A_19fCI6Zc0_0(.din(n34038), .dout(n34041));
    jdff dff_A_lpZGXu0y2_0(.din(n34035), .dout(n34038));
    jdff dff_A_qpsctrvC1_0(.din(n34032), .dout(n34035));
    jdff dff_A_BdxTEUHS9_0(.din(n34029), .dout(n34032));
    jdff dff_A_r8XYs8Hd3_0(.din(n34026), .dout(n34029));
    jdff dff_A_8Uat7pf94_0(.din(n34023), .dout(n34026));
    jdff dff_A_QxPjcjDw3_0(.din(n34020), .dout(n34023));
    jdff dff_A_O1DAztnV3_0(.din(n34017), .dout(n34020));
    jdff dff_A_QQyIJLSQ3_0(.din(n34014), .dout(n34017));
    jdff dff_A_RhKMlQyO5_0(.din(n34011), .dout(n34014));
    jdff dff_A_G3QlGVPr3_0(.din(n34008), .dout(n34011));
    jdff dff_A_awNIhsVs6_0(.din(n34005), .dout(n34008));
    jdff dff_A_3gSVC3rH2_0(.din(n34002), .dout(n34005));
    jdff dff_A_AxMvzLU83_0(.din(n33999), .dout(n34002));
    jdff dff_A_RAueuALN5_0(.din(n33996), .dout(n33999));
    jdff dff_A_yUimV0Bh9_0(.din(n33993), .dout(n33996));
    jdff dff_A_zDZVouRh0_0(.din(n33990), .dout(n33993));
    jdff dff_A_Mh1ZkqB01_0(.din(n33987), .dout(n33990));
    jdff dff_A_B9jwKtEi0_0(.din(n33984), .dout(n33987));
    jdff dff_A_TNghpsKr9_0(.din(n33981), .dout(n33984));
    jdff dff_A_tGrCqxOn3_0(.din(n33978), .dout(n33981));
    jdff dff_A_RDyDpIKL3_0(.din(n33975), .dout(n33978));
    jdff dff_A_J1woOXAB6_0(.din(n33972), .dout(n33975));
    jdff dff_A_fKVkzAPb6_0(.din(n33969), .dout(n33972));
    jdff dff_A_gqknKMfQ0_0(.din(n33966), .dout(n33969));
    jdff dff_A_aYXvXpA00_0(.din(n33963), .dout(n33966));
    jdff dff_A_i9vTsd9D9_0(.din(n33960), .dout(n33963));
    jdff dff_A_3c7oaCSD7_0(.din(n33957), .dout(n33960));
    jdff dff_A_Wgwibnsv3_0(.din(n33954), .dout(n33957));
    jdff dff_A_D8PKPrPK0_0(.din(n33951), .dout(n33954));
    jdff dff_A_lSRreIfz1_0(.din(n33948), .dout(n33951));
    jdff dff_A_FERBmCp34_0(.din(n33945), .dout(n33948));
    jdff dff_A_RUYPQsDY7_2(.din(n511), .dout(n33945));
    jdff dff_A_xu0HXtiL9_0(.din(n33939), .dout(G2548gat));
    jdff dff_A_nbpHtQDg8_0(.din(n33936), .dout(n33939));
    jdff dff_A_gkNXnR409_0(.din(n33933), .dout(n33936));
    jdff dff_A_KGlUjaKO8_0(.din(n33930), .dout(n33933));
    jdff dff_A_Ocxo46xu6_0(.din(n33927), .dout(n33930));
    jdff dff_A_qaoRYh0E1_0(.din(n33924), .dout(n33927));
    jdff dff_A_csHlvfVS8_0(.din(n33921), .dout(n33924));
    jdff dff_A_gArMwLcF2_0(.din(n33918), .dout(n33921));
    jdff dff_A_fR8LNZsj5_0(.din(n33915), .dout(n33918));
    jdff dff_A_09EW2rDW4_0(.din(n33912), .dout(n33915));
    jdff dff_A_qpXikVWH1_0(.din(n33909), .dout(n33912));
    jdff dff_A_8AIsEPAw5_0(.din(n33906), .dout(n33909));
    jdff dff_A_HnpzXgXD2_0(.din(n33903), .dout(n33906));
    jdff dff_A_S1jL8bHB9_0(.din(n33900), .dout(n33903));
    jdff dff_A_EPvQzi5F2_0(.din(n33897), .dout(n33900));
    jdff dff_A_xFfKk3BB7_0(.din(n33894), .dout(n33897));
    jdff dff_A_wR71dWOy1_0(.din(n33891), .dout(n33894));
    jdff dff_A_MYsLJGFR8_0(.din(n33888), .dout(n33891));
    jdff dff_A_W1ZfZD3z6_0(.din(n33885), .dout(n33888));
    jdff dff_A_v8EUxYoE6_0(.din(n33882), .dout(n33885));
    jdff dff_A_G4B3b3nI4_0(.din(n33879), .dout(n33882));
    jdff dff_A_cS8XrOzc9_0(.din(n33876), .dout(n33879));
    jdff dff_A_3pPmDxCy2_0(.din(n33873), .dout(n33876));
    jdff dff_A_R0kt95vW2_0(.din(n33870), .dout(n33873));
    jdff dff_A_io4ikEzF2_0(.din(n33867), .dout(n33870));
    jdff dff_A_ysW22CG84_0(.din(n33864), .dout(n33867));
    jdff dff_A_uYbfkqNb0_0(.din(n33861), .dout(n33864));
    jdff dff_A_Kqrr3aOs4_0(.din(n33858), .dout(n33861));
    jdff dff_A_EvxITJEX9_0(.din(n33855), .dout(n33858));
    jdff dff_A_Nk71cV790_0(.din(n33852), .dout(n33855));
    jdff dff_A_PY1Wxqvw7_0(.din(n33849), .dout(n33852));
    jdff dff_A_40sP0Bmi0_0(.din(n33846), .dout(n33849));
    jdff dff_A_LD930DMu4_0(.din(n33843), .dout(n33846));
    jdff dff_A_CFZpnAs40_0(.din(n33840), .dout(n33843));
    jdff dff_A_MvLXYLxv5_0(.din(n33837), .dout(n33840));
    jdff dff_A_FVKsp7M03_0(.din(n33834), .dout(n33837));
    jdff dff_A_dEmfk64u5_0(.din(n33831), .dout(n33834));
    jdff dff_A_wJOokmHS5_0(.din(n33828), .dout(n33831));
    jdff dff_A_QFUs9Ila8_0(.din(n33825), .dout(n33828));
    jdff dff_A_wZULdw2L9_0(.din(n33822), .dout(n33825));
    jdff dff_A_FbLdgRgn8_0(.din(n33819), .dout(n33822));
    jdff dff_A_Fl6TlHCf6_0(.din(n33816), .dout(n33819));
    jdff dff_A_QnVD2dQL5_0(.din(n33813), .dout(n33816));
    jdff dff_A_GBYgOpBd7_0(.din(n33810), .dout(n33813));
    jdff dff_A_AjK0qOSk1_0(.din(n33807), .dout(n33810));
    jdff dff_A_hJBYENos7_0(.din(n33804), .dout(n33807));
    jdff dff_A_AeEhZNnb2_0(.din(n33801), .dout(n33804));
    jdff dff_A_UGT5LskC9_0(.din(n33798), .dout(n33801));
    jdff dff_A_pnrcnN4J1_0(.din(n33795), .dout(n33798));
    jdff dff_A_CXGxDzkH2_0(.din(n33792), .dout(n33795));
    jdff dff_A_Ja78ZvCe2_0(.din(n33789), .dout(n33792));
    jdff dff_A_rOIcZZDu9_0(.din(n33786), .dout(n33789));
    jdff dff_A_tbpEb7BY9_0(.din(n33783), .dout(n33786));
    jdff dff_A_nyLnwlWy9_0(.din(n33780), .dout(n33783));
    jdff dff_A_APpQpcHi8_0(.din(n33777), .dout(n33780));
    jdff dff_A_6gqQAzuL4_0(.din(n33774), .dout(n33777));
    jdff dff_A_z0wpr7zP6_0(.din(n33771), .dout(n33774));
    jdff dff_A_Tcg6oiJu6_0(.din(n33768), .dout(n33771));
    jdff dff_A_nBUqx7vL4_0(.din(n33765), .dout(n33768));
    jdff dff_A_ZiAS5RSm0_0(.din(n33762), .dout(n33765));
    jdff dff_A_EdpmgK5y6_0(.din(n33759), .dout(n33762));
    jdff dff_A_AUDRS8GG1_0(.din(n33756), .dout(n33759));
    jdff dff_A_u59OK6MR6_2(.din(n367), .dout(n33756));
    jdff dff_A_49Gda4N82_0(.din(n33750), .dout(G2223gat));
    jdff dff_A_7E3bbe5x1_0(.din(n33747), .dout(n33750));
    jdff dff_A_jTlifDtK4_0(.din(n33744), .dout(n33747));
    jdff dff_A_deKqIOxp6_0(.din(n33741), .dout(n33744));
    jdff dff_A_G2CYWKhS2_0(.din(n33738), .dout(n33741));
    jdff dff_A_U61jtEFG5_0(.din(n33735), .dout(n33738));
    jdff dff_A_HkFVYLsx4_0(.din(n33732), .dout(n33735));
    jdff dff_A_dahJqzWt9_0(.din(n33729), .dout(n33732));
    jdff dff_A_CrKFiCqf1_0(.din(n33726), .dout(n33729));
    jdff dff_A_72m3X7Vd2_0(.din(n33723), .dout(n33726));
    jdff dff_A_K1YnwdvK1_0(.din(n33720), .dout(n33723));
    jdff dff_A_TvsniWpr4_0(.din(n33717), .dout(n33720));
    jdff dff_A_KCMgCse62_0(.din(n33714), .dout(n33717));
    jdff dff_A_u1mu6W740_0(.din(n33711), .dout(n33714));
    jdff dff_A_hVdqspZl2_0(.din(n33708), .dout(n33711));
    jdff dff_A_KHvpRFUN1_0(.din(n33705), .dout(n33708));
    jdff dff_A_lJ3FDdwu0_0(.din(n33702), .dout(n33705));
    jdff dff_A_fUn8xO5C3_0(.din(n33699), .dout(n33702));
    jdff dff_A_FslfGcvR1_0(.din(n33696), .dout(n33699));
    jdff dff_A_EOe5qfW22_0(.din(n33693), .dout(n33696));
    jdff dff_A_Q9mGDfoZ7_0(.din(n33690), .dout(n33693));
    jdff dff_A_aUujZGe54_0(.din(n33687), .dout(n33690));
    jdff dff_A_CuZuBnGt2_0(.din(n33684), .dout(n33687));
    jdff dff_A_q8X3NXYg4_0(.din(n33681), .dout(n33684));
    jdff dff_A_IXbyTuFa5_0(.din(n33678), .dout(n33681));
    jdff dff_A_yJZO6A449_0(.din(n33675), .dout(n33678));
    jdff dff_A_6kIevxMP0_0(.din(n33672), .dout(n33675));
    jdff dff_A_kJPi2ieZ8_0(.din(n33669), .dout(n33672));
    jdff dff_A_GwQLWlZ29_0(.din(n33666), .dout(n33669));
    jdff dff_A_Df4bkLAL2_0(.din(n33663), .dout(n33666));
    jdff dff_A_Tjw3eYba6_0(.din(n33660), .dout(n33663));
    jdff dff_A_NhVoXUf70_0(.din(n33657), .dout(n33660));
    jdff dff_A_WvDEKKvF0_0(.din(n33654), .dout(n33657));
    jdff dff_A_E6nEfCKl2_0(.din(n33651), .dout(n33654));
    jdff dff_A_TglgS7hl8_0(.din(n33648), .dout(n33651));
    jdff dff_A_ozZXWHbn6_0(.din(n33645), .dout(n33648));
    jdff dff_A_yZmlUCb06_0(.din(n33642), .dout(n33645));
    jdff dff_A_2QpKr6gk8_0(.din(n33639), .dout(n33642));
    jdff dff_A_zQgRC7OG7_0(.din(n33636), .dout(n33639));
    jdff dff_A_lBDkvRUu2_0(.din(n33633), .dout(n33636));
    jdff dff_A_xly4i3pr4_0(.din(n33630), .dout(n33633));
    jdff dff_A_DSpPYdNM5_0(.din(n33627), .dout(n33630));
    jdff dff_A_Gi9v8lA62_0(.din(n33624), .dout(n33627));
    jdff dff_A_gYj8Sm3I7_0(.din(n33621), .dout(n33624));
    jdff dff_A_Yg4WvvCX9_0(.din(n33618), .dout(n33621));
    jdff dff_A_OJlLLM5O7_0(.din(n33615), .dout(n33618));
    jdff dff_A_xzotiHdE6_0(.din(n33612), .dout(n33615));
    jdff dff_A_DHMaLv0r3_0(.din(n33609), .dout(n33612));
    jdff dff_A_wHt4zteD1_0(.din(n33606), .dout(n33609));
    jdff dff_A_ZIiaFsVb2_0(.din(n33603), .dout(n33606));
    jdff dff_A_kAcV4oxf0_0(.din(n33600), .dout(n33603));
    jdff dff_A_guS0juLC7_0(.din(n33597), .dout(n33600));
    jdff dff_A_l58SNuKq3_0(.din(n33594), .dout(n33597));
    jdff dff_A_c37TLJfK1_0(.din(n33591), .dout(n33594));
    jdff dff_A_188WxzeC5_0(.din(n33588), .dout(n33591));
    jdff dff_A_P9xwoMHP3_0(.din(n33585), .dout(n33588));
    jdff dff_A_C5iXU3DY6_0(.din(n33582), .dout(n33585));
    jdff dff_A_kWQRDeEs6_0(.din(n33579), .dout(n33582));
    jdff dff_A_dVLD3Ro47_0(.din(n33576), .dout(n33579));
    jdff dff_A_mwkUC4UP9_0(.din(n33573), .dout(n33576));
    jdff dff_A_dIuFx3vT5_0(.din(n33570), .dout(n33573));
    jdff dff_A_g6MFUHP52_0(.din(n33567), .dout(n33570));
    jdff dff_A_abpLbixo1_0(.din(n33564), .dout(n33567));
    jdff dff_A_GTMw07LJ7_0(.din(n33561), .dout(n33564));
    jdff dff_A_SC53etb39_0(.din(n33558), .dout(n33561));
    jdff dff_A_ihkYZoXx2_2(.din(n235), .dout(n33558));
    jdff dff_A_ZO8vVKK11_0(.din(n33552), .dout(G1901gat));
    jdff dff_A_QOUpQTe75_0(.din(n33549), .dout(n33552));
    jdff dff_A_UwY88ub12_0(.din(n33546), .dout(n33549));
    jdff dff_A_dA0i9buk1_0(.din(n33543), .dout(n33546));
    jdff dff_A_MYeHyNuP9_0(.din(n33540), .dout(n33543));
    jdff dff_A_1yl3Tr0K0_0(.din(n33537), .dout(n33540));
    jdff dff_A_1AMb7ab21_0(.din(n33534), .dout(n33537));
    jdff dff_A_KGNYuGTP1_0(.din(n33531), .dout(n33534));
    jdff dff_A_rYcqg5M32_0(.din(n33528), .dout(n33531));
    jdff dff_A_wCUZ1sVW6_0(.din(n33525), .dout(n33528));
    jdff dff_A_mBg5cCz30_0(.din(n33522), .dout(n33525));
    jdff dff_A_zVR9oK5w1_0(.din(n33519), .dout(n33522));
    jdff dff_A_KgoDcpQ35_0(.din(n33516), .dout(n33519));
    jdff dff_A_JFGtlC5t4_0(.din(n33513), .dout(n33516));
    jdff dff_A_8eNjoxBn4_0(.din(n33510), .dout(n33513));
    jdff dff_A_qqjCttYu8_0(.din(n33507), .dout(n33510));
    jdff dff_A_G2CKQlSS9_0(.din(n33504), .dout(n33507));
    jdff dff_A_NTln6Xsz8_0(.din(n33501), .dout(n33504));
    jdff dff_A_nD9hgrCF5_0(.din(n33498), .dout(n33501));
    jdff dff_A_ATBUR3tj3_0(.din(n33495), .dout(n33498));
    jdff dff_A_P5yrAl677_0(.din(n33492), .dout(n33495));
    jdff dff_A_pIIYnlCH7_0(.din(n33489), .dout(n33492));
    jdff dff_A_K11Uetar0_0(.din(n33486), .dout(n33489));
    jdff dff_A_Yqpxj6UB9_0(.din(n33483), .dout(n33486));
    jdff dff_A_Ia2f72Ci3_0(.din(n33480), .dout(n33483));
    jdff dff_A_tR05fWiy5_0(.din(n33477), .dout(n33480));
    jdff dff_A_wNigYBvw4_0(.din(n33474), .dout(n33477));
    jdff dff_A_9rqH1VZm4_0(.din(n33471), .dout(n33474));
    jdff dff_A_RYFMtx8M8_0(.din(n33468), .dout(n33471));
    jdff dff_A_qLjqvj5B3_0(.din(n33465), .dout(n33468));
    jdff dff_A_DWnq424u4_0(.din(n33462), .dout(n33465));
    jdff dff_A_rfogrGqH8_0(.din(n33459), .dout(n33462));
    jdff dff_A_0iddeGKK0_0(.din(n33456), .dout(n33459));
    jdff dff_A_YfxDWxVz7_0(.din(n33453), .dout(n33456));
    jdff dff_A_m6TfIlGV0_0(.din(n33450), .dout(n33453));
    jdff dff_A_8u57dXdM6_0(.din(n33447), .dout(n33450));
    jdff dff_A_cpQj61Q11_0(.din(n33444), .dout(n33447));
    jdff dff_A_cdoOIn1i1_0(.din(n33441), .dout(n33444));
    jdff dff_A_ZJOgWIsk0_0(.din(n33438), .dout(n33441));
    jdff dff_A_npB4fh242_0(.din(n33435), .dout(n33438));
    jdff dff_A_yWfJCSsM6_0(.din(n33432), .dout(n33435));
    jdff dff_A_Gox6RqJK1_0(.din(n33429), .dout(n33432));
    jdff dff_A_fJDhVgOz5_0(.din(n33426), .dout(n33429));
    jdff dff_A_sxyqDQwb0_0(.din(n33423), .dout(n33426));
    jdff dff_A_tPS7lwTn4_0(.din(n33420), .dout(n33423));
    jdff dff_A_B5EsmqgE8_0(.din(n33417), .dout(n33420));
    jdff dff_A_ue27BoMK0_0(.din(n33414), .dout(n33417));
    jdff dff_A_WSus9DQn2_0(.din(n33411), .dout(n33414));
    jdff dff_A_R6ur1G3R4_0(.din(n33408), .dout(n33411));
    jdff dff_A_X0r76xsS0_0(.din(n33405), .dout(n33408));
    jdff dff_A_LZmai8il1_0(.din(n33402), .dout(n33405));
    jdff dff_A_IsUssCpU0_0(.din(n33399), .dout(n33402));
    jdff dff_A_OsT9bsmP2_0(.din(n33396), .dout(n33399));
    jdff dff_A_GjzVWqgl2_0(.din(n33393), .dout(n33396));
    jdff dff_A_n6lkNNPd0_0(.din(n33390), .dout(n33393));
    jdff dff_A_J5JYw0Cg9_0(.din(n33387), .dout(n33390));
    jdff dff_A_fiuBGqNA6_0(.din(n33384), .dout(n33387));
    jdff dff_A_1ScT891b9_0(.din(n33381), .dout(n33384));
    jdff dff_A_itTsayCO6_0(.din(n33378), .dout(n33381));
    jdff dff_A_16J9Ltb47_0(.din(n33375), .dout(n33378));
    jdff dff_A_ee17YuJ77_0(.din(n33372), .dout(n33375));
    jdff dff_A_teGtxT7P7_0(.din(n33369), .dout(n33372));
    jdff dff_A_V99KVqkz2_0(.din(n33366), .dout(n33369));
    jdff dff_A_o8HRGzKQ7_0(.din(n33363), .dout(n33366));
    jdff dff_A_Dpyr2gKH1_0(.din(n33360), .dout(n33363));
    jdff dff_A_n57bBGQP3_0(.din(n33357), .dout(n33360));
    jdff dff_A_lC3t4jek6_0(.din(n33354), .dout(n33357));
    jdff dff_A_IKCfQeGD9_0(.din(n33351), .dout(n33354));
    jdff dff_A_bk66JIRc7_2(.din(n156), .dout(n33351));
    jdff dff_A_7LlMToQR5_0(.din(n33345), .dout(G1581gat));
    jdff dff_A_NoShJDYn0_0(.din(n33342), .dout(n33345));
    jdff dff_A_2Yd292y00_0(.din(n33339), .dout(n33342));
    jdff dff_A_UpFK9dU44_0(.din(n33336), .dout(n33339));
    jdff dff_A_BvEGz6x93_0(.din(n33333), .dout(n33336));
    jdff dff_A_TQU6YDac1_0(.din(n33330), .dout(n33333));
    jdff dff_A_KseXWj2U4_0(.din(n33327), .dout(n33330));
    jdff dff_A_JWJAKf7Q0_0(.din(n33324), .dout(n33327));
    jdff dff_A_FAYZJtDj5_0(.din(n33321), .dout(n33324));
    jdff dff_A_aligU5lK9_0(.din(n33318), .dout(n33321));
    jdff dff_A_Ulr0o6TO5_0(.din(n33315), .dout(n33318));
    jdff dff_A_RhiqKDrt0_0(.din(n33312), .dout(n33315));
    jdff dff_A_35XEmrYb4_0(.din(n33309), .dout(n33312));
    jdff dff_A_D1V1DfQ07_0(.din(n33306), .dout(n33309));
    jdff dff_A_U4GUl6kQ8_0(.din(n33303), .dout(n33306));
    jdff dff_A_7ZVKcPhK8_0(.din(n33300), .dout(n33303));
    jdff dff_A_NxZsVi9t8_0(.din(n33297), .dout(n33300));
    jdff dff_A_rY2wFcGx5_0(.din(n33294), .dout(n33297));
    jdff dff_A_BhZ3RtV71_0(.din(n33291), .dout(n33294));
    jdff dff_A_YerZPohO3_0(.din(n33288), .dout(n33291));
    jdff dff_A_1CBWRDSR3_0(.din(n33285), .dout(n33288));
    jdff dff_A_MXdsDW6I3_0(.din(n33282), .dout(n33285));
    jdff dff_A_7G07MALF0_0(.din(n33279), .dout(n33282));
    jdff dff_A_N8OZYB3v1_0(.din(n33276), .dout(n33279));
    jdff dff_A_khpJA9Vz3_0(.din(n33273), .dout(n33276));
    jdff dff_A_SF7FExQW6_0(.din(n33270), .dout(n33273));
    jdff dff_A_M8fUQQ3i5_0(.din(n33267), .dout(n33270));
    jdff dff_A_MHH2uqGI2_0(.din(n33264), .dout(n33267));
    jdff dff_A_05f6D0SG2_0(.din(n33261), .dout(n33264));
    jdff dff_A_agohsC0X8_0(.din(n33258), .dout(n33261));
    jdff dff_A_LpTzvMRc1_0(.din(n33255), .dout(n33258));
    jdff dff_A_Ct3URjSe1_0(.din(n33252), .dout(n33255));
    jdff dff_A_LFJqh0xF9_0(.din(n33249), .dout(n33252));
    jdff dff_A_kpY6t2RW1_0(.din(n33246), .dout(n33249));
    jdff dff_A_kpXii2qt5_0(.din(n33243), .dout(n33246));
    jdff dff_A_8yiAk4tD8_0(.din(n33240), .dout(n33243));
    jdff dff_A_xgRwYFbb3_0(.din(n33237), .dout(n33240));
    jdff dff_A_S0FYVG1S0_0(.din(n33234), .dout(n33237));
    jdff dff_A_JGeJVqJn3_0(.din(n33231), .dout(n33234));
    jdff dff_A_cdYbLOH19_0(.din(n33228), .dout(n33231));
    jdff dff_A_merzZsE68_0(.din(n33225), .dout(n33228));
    jdff dff_A_JkSPIyLB4_0(.din(n33222), .dout(n33225));
    jdff dff_A_OMTNsVM81_0(.din(n33219), .dout(n33222));
    jdff dff_A_FOjuWzTf0_0(.din(n33216), .dout(n33219));
    jdff dff_A_FKECd3dk6_0(.din(n33213), .dout(n33216));
    jdff dff_A_YcFPflsI3_0(.din(n33210), .dout(n33213));
    jdff dff_A_5ameRFIA4_0(.din(n33207), .dout(n33210));
    jdff dff_A_zxKvatpL2_0(.din(n33204), .dout(n33207));
    jdff dff_A_By7SmI832_0(.din(n33201), .dout(n33204));
    jdff dff_A_HxOUhU9n0_0(.din(n33198), .dout(n33201));
    jdff dff_A_6CjaYoLO1_0(.din(n33195), .dout(n33198));
    jdff dff_A_LVV36kZL1_0(.din(n33192), .dout(n33195));
    jdff dff_A_ktjbljTE0_0(.din(n33189), .dout(n33192));
    jdff dff_A_i9vzbcfc5_0(.din(n33186), .dout(n33189));
    jdff dff_A_jzfbyS4I7_0(.din(n33183), .dout(n33186));
    jdff dff_A_TTeC5tV14_0(.din(n33180), .dout(n33183));
    jdff dff_A_vfDdvrFO3_0(.din(n33177), .dout(n33180));
    jdff dff_A_p7puu2no7_0(.din(n33174), .dout(n33177));
    jdff dff_A_PFsb8Yf51_0(.din(n33171), .dout(n33174));
    jdff dff_A_W2yE3rvl0_0(.din(n33168), .dout(n33171));
    jdff dff_A_jDtwgd2i4_0(.din(n33165), .dout(n33168));
    jdff dff_A_fzAJolga8_0(.din(n33162), .dout(n33165));
    jdff dff_A_H3ssAJR90_0(.din(n33159), .dout(n33162));
    jdff dff_A_8B23OrgM6_0(.din(n33156), .dout(n33159));
    jdff dff_A_wGvRFbvr5_0(.din(n33153), .dout(n33156));
    jdff dff_A_or75KAGO6_0(.din(n33150), .dout(n33153));
    jdff dff_A_peI4Grcg6_0(.din(n33147), .dout(n33150));
    jdff dff_A_5RDbOpvM5_0(.din(n33144), .dout(n33147));
    jdff dff_A_SjmfjdMv9_0(.din(n33141), .dout(n33144));
    jdff dff_A_Kc8P7odh1_0(.din(n33138), .dout(n33141));
    jdff dff_A_p64RLqHA6_0(.din(n33135), .dout(n33138));
    jdff dff_A_YXiv6Yx23_2(.din(n94), .dout(n33135));
    jdff dff_A_P7Rt7lic5_0(.din(n33129), .dout(G545gat));
    jdff dff_A_98G6dCIX3_0(.din(n33126), .dout(n33129));
    jdff dff_A_aumP3CjT5_0(.din(n33123), .dout(n33126));
    jdff dff_A_VBKTxnU93_0(.din(n33120), .dout(n33123));
    jdff dff_A_cYf0crjQ1_0(.din(n33117), .dout(n33120));
    jdff dff_A_Giinq9195_0(.din(n33114), .dout(n33117));
    jdff dff_A_P4linBrj6_0(.din(n33111), .dout(n33114));
    jdff dff_A_irNDFiMt4_0(.din(n33108), .dout(n33111));
    jdff dff_A_NTuBIZC16_0(.din(n33105), .dout(n33108));
    jdff dff_A_qHIUtCQv8_0(.din(n33102), .dout(n33105));
    jdff dff_A_LM1FenCm6_0(.din(n33099), .dout(n33102));
    jdff dff_A_PWbMRYmD2_0(.din(n33096), .dout(n33099));
    jdff dff_A_jOaAEEDT2_0(.din(n33093), .dout(n33096));
    jdff dff_A_NPgZlsW65_0(.din(n33090), .dout(n33093));
    jdff dff_A_WAUmUw6U6_0(.din(n33087), .dout(n33090));
    jdff dff_A_kPG8ZVs28_0(.din(n33084), .dout(n33087));
    jdff dff_A_s78YTkNL7_0(.din(n33081), .dout(n33084));
    jdff dff_A_5gfEFDge0_0(.din(n33078), .dout(n33081));
    jdff dff_A_CgyGOVCN8_0(.din(n33075), .dout(n33078));
    jdff dff_A_dALT4q3n8_0(.din(n33072), .dout(n33075));
    jdff dff_A_OlYLz6wX1_0(.din(n33069), .dout(n33072));
    jdff dff_A_iYmAUuzm0_0(.din(n33066), .dout(n33069));
    jdff dff_A_lEDkFNI38_0(.din(n33063), .dout(n33066));
    jdff dff_A_slabGQfO5_0(.din(n33060), .dout(n33063));
    jdff dff_A_8qhQPsyN2_0(.din(n33057), .dout(n33060));
    jdff dff_A_TTH40hc38_0(.din(n33054), .dout(n33057));
    jdff dff_A_6Fb6qF1p2_0(.din(n33051), .dout(n33054));
    jdff dff_A_ZrwPCZx36_0(.din(n33048), .dout(n33051));
    jdff dff_A_LvmED0907_0(.din(n33045), .dout(n33048));
    jdff dff_A_qce9Ezw64_0(.din(n33042), .dout(n33045));
    jdff dff_A_98ErYpfl4_0(.din(n33039), .dout(n33042));
    jdff dff_A_ny7PYMA96_0(.din(n33036), .dout(n33039));
    jdff dff_A_AguR2ECu4_0(.din(n33033), .dout(n33036));
    jdff dff_A_2zk8f1AU5_0(.din(n33030), .dout(n33033));
    jdff dff_A_4MqFCvoH0_0(.din(n33027), .dout(n33030));
    jdff dff_A_nrufeGX17_0(.din(n33024), .dout(n33027));
    jdff dff_A_mLPPM5sn6_0(.din(n33021), .dout(n33024));
    jdff dff_A_548WKCsg9_0(.din(n33018), .dout(n33021));
    jdff dff_A_yJGhVhhl3_0(.din(n33015), .dout(n33018));
    jdff dff_A_mtZguglp8_0(.din(n33012), .dout(n33015));
    jdff dff_A_YN4nNPtx9_0(.din(n33009), .dout(n33012));
    jdff dff_A_hwq5kgka2_0(.din(n33006), .dout(n33009));
    jdff dff_A_AGJH553l7_0(.din(n33003), .dout(n33006));
    jdff dff_A_1D1Y6BUd5_0(.din(n33000), .dout(n33003));
    jdff dff_A_USQYQHf75_0(.din(n32997), .dout(n33000));
    jdff dff_A_1TftoEOW8_0(.din(n32994), .dout(n32997));
    jdff dff_A_6YgT5HmA5_0(.din(n32991), .dout(n32994));
    jdff dff_A_KdfBZQGv4_0(.din(n32988), .dout(n32991));
    jdff dff_A_UqtOzkKK3_0(.din(n32985), .dout(n32988));
    jdff dff_A_JcuAN9sZ9_0(.din(n32982), .dout(n32985));
    jdff dff_A_xu7skIGf8_0(.din(n32979), .dout(n32982));
    jdff dff_A_itn12WyD8_0(.din(n32976), .dout(n32979));
    jdff dff_A_J9yBLkpz7_0(.din(n32973), .dout(n32976));
    jdff dff_A_XYj3p9UF8_0(.din(n32970), .dout(n32973));
    jdff dff_A_NrivGG2h2_0(.din(n32967), .dout(n32970));
    jdff dff_A_bjAgsrpW0_0(.din(n32964), .dout(n32967));
    jdff dff_A_BHSr3EmJ0_0(.din(n32961), .dout(n32964));
    jdff dff_A_77ogvPP86_0(.din(n32958), .dout(n32961));
    jdff dff_A_9l1niQwx9_0(.din(n32955), .dout(n32958));
    jdff dff_A_4IMo6afp9_0(.din(n32952), .dout(n32955));
    jdff dff_A_7eGlORmV1_0(.din(n32949), .dout(n32952));
    jdff dff_A_AlYXZySL1_0(.din(n32946), .dout(n32949));
    jdff dff_A_sGgHrYJb0_0(.din(n32943), .dout(n32946));
    jdff dff_A_A30gUBkh9_0(.din(n32940), .dout(n32943));
    jdff dff_A_Qu8OTBtf4_0(.din(n32937), .dout(n32940));
    jdff dff_A_44kvQYtZ7_0(.din(n32934), .dout(n32937));
    jdff dff_A_fE7kvKyq3_0(.din(n32931), .dout(n32934));
    jdff dff_A_pr6bOVe40_0(.din(n32928), .dout(n32931));
    jdff dff_A_fGX7JfCv5_0(.din(n32925), .dout(n32928));
    jdff dff_A_BU4rTDgm3_0(.din(n32922), .dout(n32925));
    jdff dff_A_qNBEAGXc1_0(.din(n32919), .dout(n32922));
    jdff dff_A_GjJySaNj3_0(.din(n32916), .dout(n32919));
    jdff dff_A_a5FiIX6v2_0(.din(n32913), .dout(n32916));
    jdff dff_A_ZHjSjUI17_0(.din(n32910), .dout(n32913));
    jdff dff_A_rE4qmGgL3_1(.din(n67), .dout(n32910));
    jdff dff_A_AhwbHvEf1_1(.din(n3228), .dout(n32907));
    jdff dff_A_LFZNbteQ8_1(.din(n32907), .dout(n32904));
    jdff dff_A_PqR25d2d6_1(.din(n32904), .dout(n32901));
    jdff dff_A_z9GPjSto8_1(.din(n32901), .dout(n32898));
    jdff dff_A_HlqjyqD42_1(.din(n32898), .dout(n32895));
    jdff dff_B_lLac3uo07_2(.din(n3235), .dout(n32893));
    jdff dff_A_VCHMQp1s7_0(.din(n2460), .dout(n32889));
    jdff dff_A_0kBr7MwZ8_0(.din(n32889), .dout(n32886));
    jdff dff_A_f2OUeufa5_0(.din(n32886), .dout(n32883));
    jdff dff_A_uLByc2El7_0(.din(n3254), .dout(n32880));
    jdff dff_A_iPbA4AM20_0(.din(n32880), .dout(n32877));
    jdff dff_A_3tzYqdid4_0(.din(n32877), .dout(n32874));
    jdff dff_B_7ocKJlph9_1(.din(n32869), .dout(n32872));
    jdff dff_B_bvM5pOaO1_1(.din(n32866), .dout(n32869));
    jdff dff_B_YmpiVlK80_1(.din(n32863), .dout(n32866));
    jdff dff_B_KZLhzZXj0_1(.din(n32860), .dout(n32863));
    jdff dff_B_5oDqQnFC4_1(.din(n3633), .dout(n32860));
    jdff dff_A_DIA0lUDf8_1(.din(n3648), .dout(n32856));
    jdff dff_A_B5pqTIi46_1(.din(n32856), .dout(n32853));
    jdff dff_A_uVjBeraU8_0(.din(n2834), .dout(n32850));
    jdff dff_A_vaNofmMD7_0(.din(n3655), .dout(n32847));
    jdff dff_A_2ggyHQ8U6_0(.din(n32847), .dout(n32844));
    jdff dff_A_U1HcrelJ0_0(.din(n32844), .dout(n32841));
    jdff dff_B_rbubUt2i7_2(.din(n32836), .dout(n32839));
    jdff dff_B_Wp4tjeBe1_2(.din(n32833), .dout(n32836));
    jdff dff_B_m1RCkkPH9_2(.din(n32830), .dout(n32833));
    jdff dff_B_WbleH03o3_2(.din(n32827), .dout(n32830));
    jdff dff_B_aMxbGL8a2_2(.din(n3663), .dout(n32827));
    jdff dff_B_rvbvWtr08_2(.din(n32821), .dout(n32824));
    jdff dff_B_snnwlZP56_2(.din(n32818), .dout(n32821));
    jdff dff_B_JD0A8qP97_2(.din(n32815), .dout(n32818));
    jdff dff_B_jWFSNWq73_2(.din(n32812), .dout(n32815));
    jdff dff_B_y9DjVUcg0_2(.din(n32809), .dout(n32812));
    jdff dff_B_yV00sn1Q7_2(.din(n32806), .dout(n32809));
    jdff dff_B_UfPsd2bc2_2(.din(n32803), .dout(n32806));
    jdff dff_B_X1hBfCeL4_2(.din(n3630), .dout(n32803));
    jdff dff_B_cmfpmCl56_1(.din(n4011), .dout(n32800));
    jdff dff_B_cqFfBWP55_2(.din(n32794), .dout(n32797));
    jdff dff_B_pKyIMzVa8_2(.din(n32791), .dout(n32794));
    jdff dff_B_UC6AoPgJ6_2(.din(n32788), .dout(n32791));
    jdff dff_B_dq8Y05WN7_2(.din(n32785), .dout(n32788));
    jdff dff_B_1yeDeOyg8_2(.din(n32782), .dout(n32785));
    jdff dff_B_YNY4Uvzw2_2(.din(n32779), .dout(n32782));
    jdff dff_B_gZ8hmKrM8_2(.din(n32776), .dout(n32779));
    jdff dff_B_Ch6Yixrm2_2(.din(n32773), .dout(n32776));
    jdff dff_B_39TboRSy1_2(.din(n32770), .dout(n32773));
    jdff dff_B_RmMAyjat2_2(.din(n4023), .dout(n32770));
    jdff dff_A_TGokZRHD9_1(.din(G307gat), .dout(n32766));
    jdff dff_A_xXmrnfsi0_1(.din(n32766), .dout(n32763));
    jdff dff_A_vhJuOkKT5_1(.din(n32763), .dout(n32760));
    jdff dff_A_XdPmzeat0_1(.din(n32760), .dout(n32757));
    jdff dff_A_m2JdDYnS7_1(.din(n32757), .dout(n32754));
    jdff dff_A_4xiO9KTf8_1(.din(n32754), .dout(n32751));
    jdff dff_A_TZ6tGNyO8_1(.din(n32751), .dout(n32748));
    jdff dff_B_IWVdypPc3_1(.din(n32743), .dout(n32746));
    jdff dff_B_PQHk8nW76_1(.din(n4030), .dout(n32743));
    jdff dff_B_B5JNyJST3_1(.din(n32737), .dout(n32740));
    jdff dff_B_pfb2HwpJ1_1(.din(n32734), .dout(n32737));
    jdff dff_B_tLoMFTzR5_1(.din(n32731), .dout(n32734));
    jdff dff_B_vwTQ4LEh0_1(.din(n32728), .dout(n32731));
    jdff dff_B_mznpII4E5_1(.din(n32725), .dout(n32728));
    jdff dff_B_35JBD6cT9_1(.din(n4027), .dout(n32725));
    jdff dff_B_GDoq4Fl55_2(.din(n4048), .dout(n32722));
    jdff dff_A_f2e2Ey2h5_0(.din(n32722), .dout(n32718));
    jdff dff_A_AKZFsUKo0_0(.din(n32718), .dout(n32715));
    jdff dff_A_Ajg6pi0s7_0(.din(n32715), .dout(n32712));
    jdff dff_B_9lWhhvuT2_2(.din(n32707), .dout(n32710));
    jdff dff_B_lIu6VCdA5_2(.din(n32704), .dout(n32707));
    jdff dff_B_R5OmwPa20_2(.din(n32701), .dout(n32704));
    jdff dff_B_7IOOwjVc4_2(.din(n32698), .dout(n32701));
    jdff dff_B_gXurmGlr9_2(.din(n32695), .dout(n32698));
    jdff dff_B_TpDxDOgf3_2(.din(n32692), .dout(n32695));
    jdff dff_B_TI8ZuKjZ5_2(.din(n32689), .dout(n32692));
    jdff dff_B_o0zYhiyG4_2(.din(n32686), .dout(n32689));
    jdff dff_B_HzGCXw0e3_2(.din(n32683), .dout(n32686));
    jdff dff_B_tcQEwGcI6_2(.din(n32680), .dout(n32683));
    jdff dff_B_bStYKeD78_2(.din(n4007), .dout(n32680));
    jdff dff_B_ekLgpStc5_1(.din(n4407), .dout(n32677));
    jdff dff_B_ZnJx9fZ55_2(.din(n4415), .dout(n32674));
    jdff dff_B_y5rNK1No5_2(.din(n32668), .dout(n32671));
    jdff dff_B_5pvmsgAx2_2(.din(n32665), .dout(n32668));
    jdff dff_B_VSTZy9ar0_2(.din(n32662), .dout(n32665));
    jdff dff_B_uHG8XFyv3_2(.din(n32659), .dout(n32662));
    jdff dff_B_MW0mOvnW2_2(.din(n32656), .dout(n32659));
    jdff dff_B_9s7J8j272_2(.din(n32653), .dout(n32656));
    jdff dff_B_USPE4sBL7_2(.din(n32650), .dout(n32653));
    jdff dff_B_qEd7GUfv1_2(.din(n32647), .dout(n32650));
    jdff dff_B_EqXigxnl2_2(.din(n32644), .dout(n32647));
    jdff dff_B_YmJ0rA5v8_2(.din(n32641), .dout(n32644));
    jdff dff_B_wAlqMFZK2_2(.din(n32638), .dout(n32641));
    jdff dff_B_Cnh3ALpc1_2(.din(n32635), .dout(n32638));
    jdff dff_B_R7U1seq15_2(.din(n32632), .dout(n32635));
    jdff dff_B_wTSyRGBe8_2(.din(n4419), .dout(n32632));
    jdff dff_B_RqiMIXOz0_2(.din(n32626), .dout(n32629));
    jdff dff_B_fxYnfF0S9_2(.din(n32623), .dout(n32626));
    jdff dff_B_mES2Qmt23_2(.din(n32620), .dout(n32623));
    jdff dff_B_T2Q7Wbqm2_2(.din(n32617), .dout(n32620));
    jdff dff_B_QqvYuJ5h8_2(.din(n32614), .dout(n32617));
    jdff dff_B_5AdnHcnK5_2(.din(n32611), .dout(n32614));
    jdff dff_B_v2k9uez14_2(.din(n32608), .dout(n32611));
    jdff dff_B_0q3OCYoI2_2(.din(n32605), .dout(n32608));
    jdff dff_B_NT2Q9DQR8_2(.din(n32602), .dout(n32605));
    jdff dff_B_utpFtmHA2_2(.din(n32599), .dout(n32602));
    jdff dff_B_fG3DPFL78_2(.din(n32596), .dout(n32599));
    jdff dff_B_RntvHVY90_2(.din(n4423), .dout(n32596));
    jdff dff_B_B9IrkPD37_2(.din(n32590), .dout(n32593));
    jdff dff_B_6J2NyFim8_2(.din(n32587), .dout(n32590));
    jdff dff_B_xVlEOmrX7_2(.din(n32584), .dout(n32587));
    jdff dff_B_pgFTnIOK6_2(.din(n32581), .dout(n32584));
    jdff dff_B_BruesTkW2_2(.din(n32578), .dout(n32581));
    jdff dff_B_y4KSNL9q6_2(.din(n32575), .dout(n32578));
    jdff dff_B_EWB7lJfj3_2(.din(n32572), .dout(n32575));
    jdff dff_B_IM5IdGkX5_2(.din(n32569), .dout(n32572));
    jdff dff_B_kCVwGTK17_2(.din(n32566), .dout(n32569));
    jdff dff_B_EZjbtMY64_2(.din(n32563), .dout(n32566));
    jdff dff_B_cbUdpB1v5_2(.din(n32560), .dout(n32563));
    jdff dff_B_XiAMtTEU2_2(.din(n32557), .dout(n32560));
    jdff dff_B_Jqv4AdE23_2(.din(n32554), .dout(n32557));
    jdff dff_B_lOEFlTU39_2(.din(n32551), .dout(n32554));
    jdff dff_B_szCQqSSU2_2(.din(n4403), .dout(n32551));
    jdff dff_B_DZrKGAMs6_1(.din(n4753), .dout(n32548));
    jdff dff_B_MWaXlhv09_2(.din(n4761), .dout(n32545));
    jdff dff_B_HNwucoHX8_2(.din(n32539), .dout(n32542));
    jdff dff_B_IjKhdoj22_2(.din(n32536), .dout(n32539));
    jdff dff_B_pM6Mmx3n7_2(.din(n32533), .dout(n32536));
    jdff dff_B_yZAGZScQ3_2(.din(n32530), .dout(n32533));
    jdff dff_B_MSt4HiVG0_2(.din(n32527), .dout(n32530));
    jdff dff_B_Ws0GHVFN2_2(.din(n32524), .dout(n32527));
    jdff dff_B_73KwR9kl1_2(.din(n32521), .dout(n32524));
    jdff dff_B_oWCisUL88_2(.din(n32518), .dout(n32521));
    jdff dff_B_SbeIj4EA9_2(.din(n32515), .dout(n32518));
    jdff dff_B_RCXf0GSK9_2(.din(n32512), .dout(n32515));
    jdff dff_B_0kdqCHKs6_2(.din(n32509), .dout(n32512));
    jdff dff_B_NfJh0SOk3_2(.din(n32506), .dout(n32509));
    jdff dff_B_qFEL7Ce34_2(.din(n32503), .dout(n32506));
    jdff dff_B_HslQ4LMC2_2(.din(n32500), .dout(n32503));
    jdff dff_B_g23d2ye54_2(.din(n32497), .dout(n32500));
    jdff dff_B_ORLY9DPs0_1(.din(n79), .dout(n10756));
    jdff dff_B_oZHNDDvI5_1(.din(n101), .dout(n10759));
    jdff dff_B_Ij8bIAet5_1(.din(n10759), .dout(n10762));
    jdff dff_B_LNzalzae9_1(.din(n10762), .dout(n10765));
    jdff dff_B_G2992b235_1(.din(n10765), .dout(n10768));
    jdff dff_B_Y9xjsZpf4_1(.din(n163), .dout(n10771));
    jdff dff_B_cB49q0lG3_1(.din(n10771), .dout(n10774));
    jdff dff_B_w7BFs5Bb5_1(.din(n10774), .dout(n10777));
    jdff dff_B_gK2wT7JT1_1(.din(n10777), .dout(n10780));
    jdff dff_B_eri50NwL8_1(.din(n10780), .dout(n10783));
    jdff dff_B_sHtfu03p8_1(.din(n10783), .dout(n10786));
    jdff dff_B_YgdLPBYN7_1(.din(n10786), .dout(n10789));
    jdff dff_B_7odUktbF4_1(.din(n242), .dout(n10792));
    jdff dff_B_AIe7hqhN6_1(.din(n10792), .dout(n10795));
    jdff dff_B_LtMhjqtt0_1(.din(n10795), .dout(n10798));
    jdff dff_B_E8jnQa4e2_1(.din(n10798), .dout(n10801));
    jdff dff_B_k0vSFOZe6_1(.din(n10801), .dout(n10804));
    jdff dff_B_KTFb8unQ6_1(.din(n10804), .dout(n10807));
    jdff dff_B_JaqLzDzK5_1(.din(n10807), .dout(n10810));
    jdff dff_B_UaZUS7uq1_1(.din(n10810), .dout(n10813));
    jdff dff_B_Gw3gHxAU9_1(.din(n10813), .dout(n10816));
    jdff dff_B_M40SSfNW0_1(.din(n10816), .dout(n10819));
    jdff dff_B_k9xHOgEo2_1(.din(n374), .dout(n10822));
    jdff dff_B_EBqLY7Wb5_1(.din(n10822), .dout(n10825));
    jdff dff_B_r2MimJxL5_1(.din(n10825), .dout(n10828));
    jdff dff_B_IuaNMIbD0_1(.din(n10828), .dout(n10831));
    jdff dff_B_IX9gG3S53_1(.din(n10831), .dout(n10834));
    jdff dff_B_LRtb1ykq6_1(.din(n10834), .dout(n10837));
    jdff dff_B_JDdX9bxa1_1(.din(n10837), .dout(n10840));
    jdff dff_B_g2lSI0ru0_1(.din(n10840), .dout(n10843));
    jdff dff_B_QBhLXg9E7_1(.din(n10843), .dout(n10846));
    jdff dff_B_6ndOoDWP9_1(.din(n10846), .dout(n10849));
    jdff dff_B_xCeUiCs86_1(.din(n10849), .dout(n10852));
    jdff dff_B_oAZrojAF4_1(.din(n10852), .dout(n10855));
    jdff dff_B_Blu890lS8_1(.din(n10855), .dout(n10858));
    jdff dff_B_XmDg2Ir85_1(.din(n518), .dout(n10861));
    jdff dff_B_sWBqXna13_1(.din(n10861), .dout(n10864));
    jdff dff_B_eH6mOT2k8_1(.din(n10864), .dout(n10867));
    jdff dff_B_h6aemqzt4_1(.din(n10867), .dout(n10870));
    jdff dff_B_zCAitGh83_1(.din(n10870), .dout(n10873));
    jdff dff_B_yFASLsDr1_1(.din(n10873), .dout(n10876));
    jdff dff_B_IJSxLSEe1_1(.din(n10876), .dout(n10879));
    jdff dff_B_PFVS4DSZ5_1(.din(n10879), .dout(n10882));
    jdff dff_B_n6Xnw4qU0_1(.din(n10882), .dout(n10885));
    jdff dff_B_0AmiNKMU8_1(.din(n10885), .dout(n10888));
    jdff dff_B_dopvKpGm6_1(.din(n10888), .dout(n10891));
    jdff dff_B_rkGExKL76_1(.din(n10891), .dout(n10894));
    jdff dff_B_vaHARmQP2_1(.din(n10894), .dout(n10897));
    jdff dff_B_EOhZpgfC5_1(.din(n10897), .dout(n10900));
    jdff dff_B_1N97qTn32_1(.din(n10900), .dout(n10903));
    jdff dff_B_tADF5loM5_1(.din(n10903), .dout(n10906));
    jdff dff_B_oz165xF91_1(.din(n681), .dout(n10909));
    jdff dff_B_7xNgGFpp8_1(.din(n10909), .dout(n10912));
    jdff dff_B_tRx9jQr35_1(.din(n10912), .dout(n10915));
    jdff dff_B_Ryqjbisa9_1(.din(n10915), .dout(n10918));
    jdff dff_B_Y3zQrAZz4_1(.din(n10918), .dout(n10921));
    jdff dff_B_FqB3WI4q8_1(.din(n10921), .dout(n10924));
    jdff dff_B_to8w4a7x0_1(.din(n10924), .dout(n10927));
    jdff dff_B_OU0FYghf6_1(.din(n10927), .dout(n10930));
    jdff dff_B_H5DkQQS58_1(.din(n10930), .dout(n10933));
    jdff dff_B_0lzxZQvI1_1(.din(n10933), .dout(n10936));
    jdff dff_B_sGY503si0_1(.din(n10936), .dout(n10939));
    jdff dff_B_N40UKXNQ2_1(.din(n10939), .dout(n10942));
    jdff dff_B_hNRrtrSy6_1(.din(n10942), .dout(n10945));
    jdff dff_B_kCq1Pjjp4_1(.din(n10945), .dout(n10948));
    jdff dff_B_5hSiQmj88_1(.din(n10948), .dout(n10951));
    jdff dff_B_53B8NZmX8_1(.din(n10951), .dout(n10954));
    jdff dff_B_sVGJtqzn0_1(.din(n10954), .dout(n10957));
    jdff dff_B_R1c7Z2Ac4_1(.din(n10957), .dout(n10960));
    jdff dff_B_Rstyn61Z1_1(.din(n10960), .dout(n10963));
    jdff dff_B_VB1NPt8j4_1(.din(n874), .dout(n10966));
    jdff dff_B_ZXGd2pai9_1(.din(n10966), .dout(n10969));
    jdff dff_B_HpRRLtSh1_1(.din(n10969), .dout(n10972));
    jdff dff_B_BP6dCCub8_1(.din(n10972), .dout(n10975));
    jdff dff_B_7EYqV7Xu1_1(.din(n10975), .dout(n10978));
    jdff dff_B_W4LGGPQG0_1(.din(n10978), .dout(n10981));
    jdff dff_B_9mt1mbrt9_1(.din(n10981), .dout(n10984));
    jdff dff_B_MeN2bBFT2_1(.din(n10984), .dout(n10987));
    jdff dff_B_MNcptmay2_1(.din(n10987), .dout(n10990));
    jdff dff_B_80TRIpfk9_1(.din(n10990), .dout(n10993));
    jdff dff_B_YMAcT9ym8_1(.din(n10993), .dout(n10996));
    jdff dff_B_dnK0GQsU2_1(.din(n10996), .dout(n10999));
    jdff dff_B_Tpuf8Jvi6_1(.din(n10999), .dout(n11002));
    jdff dff_B_piRrKy2c2_1(.din(n11002), .dout(n11005));
    jdff dff_B_r4gZneIh8_1(.din(n11005), .dout(n11008));
    jdff dff_B_ZDLBo6Uh5_1(.din(n11008), .dout(n11011));
    jdff dff_B_WzugrBuw6_1(.din(n11011), .dout(n11014));
    jdff dff_B_vQoBen6M1_1(.din(n11014), .dout(n11017));
    jdff dff_B_ZqgtYdFw3_1(.din(n11017), .dout(n11020));
    jdff dff_B_Cq3OTBLI9_1(.din(n11020), .dout(n11023));
    jdff dff_B_By0i8jzb1_1(.din(n11023), .dout(n11026));
    jdff dff_B_sWvwVGJZ8_1(.din(n11026), .dout(n11029));
    jdff dff_B_VoQ6TS7b0_1(.din(n1094), .dout(n11032));
    jdff dff_B_Wle8A4Yf0_1(.din(n11032), .dout(n11035));
    jdff dff_B_UQQW8iTz5_1(.din(n11035), .dout(n11038));
    jdff dff_B_itdCWixZ0_1(.din(n11038), .dout(n11041));
    jdff dff_B_V5JRKZ0E7_1(.din(n11041), .dout(n11044));
    jdff dff_B_nuTxSf3V6_1(.din(n11044), .dout(n11047));
    jdff dff_B_NsCMPFEu6_1(.din(n11047), .dout(n11050));
    jdff dff_B_VTRLNAiW9_1(.din(n11050), .dout(n11053));
    jdff dff_B_MKOKdvzz0_1(.din(n11053), .dout(n11056));
    jdff dff_B_rLdClAAR1_1(.din(n11056), .dout(n11059));
    jdff dff_B_tjssuTd70_1(.din(n11059), .dout(n11062));
    jdff dff_B_OLX31m4k8_1(.din(n11062), .dout(n11065));
    jdff dff_B_aIeLOVwR2_1(.din(n11065), .dout(n11068));
    jdff dff_B_uC8AU9eC6_1(.din(n11068), .dout(n11071));
    jdff dff_B_IQ226zB29_1(.din(n11071), .dout(n11074));
    jdff dff_B_G9jovtSI4_1(.din(n11074), .dout(n11077));
    jdff dff_B_mmDSTvj04_1(.din(n11077), .dout(n11080));
    jdff dff_B_mDnqxGGm3_1(.din(n11080), .dout(n11083));
    jdff dff_B_BPQLcRlU0_1(.din(n11083), .dout(n11086));
    jdff dff_B_aiGt8Dic1_1(.din(n11086), .dout(n11089));
    jdff dff_B_s52Nu9LV3_1(.din(n11089), .dout(n11092));
    jdff dff_B_bSVOMIX40_1(.din(n11092), .dout(n11095));
    jdff dff_B_BJLX2naj7_1(.din(n11095), .dout(n11098));
    jdff dff_B_vcPR8CNy8_1(.din(n11098), .dout(n11101));
    jdff dff_B_EdoSg5X52_1(.din(n11101), .dout(n11104));
    jdff dff_B_4gsK11Xq9_1(.din(n1338), .dout(n11107));
    jdff dff_B_RiXaZqSO7_1(.din(n11107), .dout(n11110));
    jdff dff_B_YEdKv2G26_1(.din(n11110), .dout(n11113));
    jdff dff_B_MqDQFoRb5_1(.din(n11113), .dout(n11116));
    jdff dff_B_XAk9Ie3e6_1(.din(n11116), .dout(n11119));
    jdff dff_B_ZcCR1UC79_1(.din(n11119), .dout(n11122));
    jdff dff_B_RYAcUgtn8_1(.din(n11122), .dout(n11125));
    jdff dff_B_6U4SpEKA3_1(.din(n11125), .dout(n11128));
    jdff dff_B_1W6La1mW7_1(.din(n11128), .dout(n11131));
    jdff dff_B_U3NVz7Gm3_1(.din(n11131), .dout(n11134));
    jdff dff_B_uqQY5foB5_1(.din(n11134), .dout(n11137));
    jdff dff_B_f8Wxk0BQ4_1(.din(n11137), .dout(n11140));
    jdff dff_B_FdNtK8LV3_1(.din(n11140), .dout(n11143));
    jdff dff_B_nk4NLpLZ7_1(.din(n11143), .dout(n11146));
    jdff dff_B_uwf0iG056_1(.din(n11146), .dout(n11149));
    jdff dff_B_NfkAaFSp9_1(.din(n11149), .dout(n11152));
    jdff dff_B_FzXvi16b5_1(.din(n11152), .dout(n11155));
    jdff dff_B_ssy4zHjc9_1(.din(n11155), .dout(n11158));
    jdff dff_B_M4pUayoG1_1(.din(n11158), .dout(n11161));
    jdff dff_B_Cr8Iu6sw6_1(.din(n11161), .dout(n11164));
    jdff dff_B_y9oGrr659_1(.din(n11164), .dout(n11167));
    jdff dff_B_leFj1xjK8_1(.din(n11167), .dout(n11170));
    jdff dff_B_1SPpOoKH7_1(.din(n11170), .dout(n11173));
    jdff dff_B_yxOTRkff3_1(.din(n11173), .dout(n11176));
    jdff dff_B_NXBs2v549_1(.din(n11176), .dout(n11179));
    jdff dff_B_QxvYgTXT7_1(.din(n11179), .dout(n11182));
    jdff dff_B_7nDGrMEn4_1(.din(n11182), .dout(n11185));
    jdff dff_B_wgsWXVkt3_1(.din(n11185), .dout(n11188));
    jdff dff_B_Ng7TGNCt8_1(.din(n1612), .dout(n11191));
    jdff dff_B_eBBkXGyg4_1(.din(n11191), .dout(n11194));
    jdff dff_B_5oeXDePC1_1(.din(n11194), .dout(n11197));
    jdff dff_B_WNVXoER12_1(.din(n11197), .dout(n11200));
    jdff dff_B_Uh2Azmw13_1(.din(n11200), .dout(n11203));
    jdff dff_B_LB5rLVW66_1(.din(n11203), .dout(n11206));
    jdff dff_B_Q251MPaq6_1(.din(n11206), .dout(n11209));
    jdff dff_B_FxOmnJYt7_1(.din(n11209), .dout(n11212));
    jdff dff_B_b4tasGne0_1(.din(n11212), .dout(n11215));
    jdff dff_B_RQpEWAFG6_1(.din(n11215), .dout(n11218));
    jdff dff_B_udbH2LjQ4_1(.din(n11218), .dout(n11221));
    jdff dff_B_e6tXLClc7_1(.din(n11221), .dout(n11224));
    jdff dff_B_k5wDjoX28_1(.din(n11224), .dout(n11227));
    jdff dff_B_7n3OBNNV4_1(.din(n11227), .dout(n11230));
    jdff dff_B_AlWaHE5r6_1(.din(n11230), .dout(n11233));
    jdff dff_B_MuIFzA4v1_1(.din(n11233), .dout(n11236));
    jdff dff_B_xpKQQ4mf8_1(.din(n11236), .dout(n11239));
    jdff dff_B_TSMfxi0V4_1(.din(n11239), .dout(n11242));
    jdff dff_B_3Tyoumh72_1(.din(n11242), .dout(n11245));
    jdff dff_B_l8S7gwAd0_1(.din(n11245), .dout(n11248));
    jdff dff_B_teFzx1jm2_1(.din(n11248), .dout(n11251));
    jdff dff_B_Mb96YJlx9_1(.din(n11251), .dout(n11254));
    jdff dff_B_8r7Z6t1f5_1(.din(n11254), .dout(n11257));
    jdff dff_B_7Cm8J7323_1(.din(n11257), .dout(n11260));
    jdff dff_B_YO0GtC4U2_1(.din(n11260), .dout(n11263));
    jdff dff_B_L1iFFo4V1_1(.din(n11263), .dout(n11266));
    jdff dff_B_DPvSa2gd6_1(.din(n11266), .dout(n11269));
    jdff dff_B_NsC6prcU0_1(.din(n11269), .dout(n11272));
    jdff dff_B_7ROqNocH2_1(.din(n11272), .dout(n11275));
    jdff dff_B_QHokTbzR1_1(.din(n11275), .dout(n11278));
    jdff dff_B_g6Pg8PGz3_1(.din(n11278), .dout(n11281));
    jdff dff_B_o02MqCH97_1(.din(n1913), .dout(n11284));
    jdff dff_B_rzPZ16kv6_1(.din(n11284), .dout(n11287));
    jdff dff_B_MKEs9oF78_1(.din(n11287), .dout(n11290));
    jdff dff_B_NeRT2TyM7_1(.din(n11290), .dout(n11293));
    jdff dff_B_vjBECOxd6_1(.din(n11293), .dout(n11296));
    jdff dff_B_1i8tbPKA3_1(.din(n11296), .dout(n11299));
    jdff dff_B_843t3xRY4_1(.din(n11299), .dout(n11302));
    jdff dff_B_bdqLC7vo9_1(.din(n11302), .dout(n11305));
    jdff dff_B_TNcI5eRw5_1(.din(n11305), .dout(n11308));
    jdff dff_B_LwTHwz5h1_1(.din(n11308), .dout(n11311));
    jdff dff_B_ogKjg4TT7_1(.din(n11311), .dout(n11314));
    jdff dff_B_1tnGRLsd5_1(.din(n11314), .dout(n11317));
    jdff dff_B_VX77IbmL3_1(.din(n11317), .dout(n11320));
    jdff dff_B_OYPlSZWi4_1(.din(n11320), .dout(n11323));
    jdff dff_B_ZyFnTC5A9_1(.din(n11323), .dout(n11326));
    jdff dff_B_Bq9AfCGp8_1(.din(n11326), .dout(n11329));
    jdff dff_B_FBymBW7n1_1(.din(n11329), .dout(n11332));
    jdff dff_B_MBqbtgjv8_1(.din(n11332), .dout(n11335));
    jdff dff_B_atvdlYe82_1(.din(n11335), .dout(n11338));
    jdff dff_B_wuJiLk3f0_1(.din(n11338), .dout(n11341));
    jdff dff_B_f8wiba432_1(.din(n11341), .dout(n11344));
    jdff dff_B_iarYdNOs8_1(.din(n11344), .dout(n11347));
    jdff dff_B_SUNnvvs75_1(.din(n11347), .dout(n11350));
    jdff dff_B_p8pivOpx2_1(.din(n11350), .dout(n11353));
    jdff dff_B_WrnvBMAh0_1(.din(n11353), .dout(n11356));
    jdff dff_B_OMVFAJ2a6_1(.din(n11356), .dout(n11359));
    jdff dff_B_YElUZzDf9_1(.din(n11359), .dout(n11362));
    jdff dff_B_U1mmLwCZ0_1(.din(n11362), .dout(n11365));
    jdff dff_B_4oTRfwQr8_1(.din(n11365), .dout(n11368));
    jdff dff_B_dKRgVAHZ8_1(.din(n11368), .dout(n11371));
    jdff dff_B_UrxQXydp3_1(.din(n11371), .dout(n11374));
    jdff dff_B_5wtEYjLL2_1(.din(n11374), .dout(n11377));
    jdff dff_B_4lb9XoRh5_1(.din(n11377), .dout(n11380));
    jdff dff_B_I9nJ9Bc26_1(.din(n11380), .dout(n11383));
    jdff dff_B_ba7yHDor7_1(.din(n2241), .dout(n11386));
    jdff dff_B_1v9PejCt4_1(.din(n11386), .dout(n11389));
    jdff dff_B_E6K7aPBy9_1(.din(n11389), .dout(n11392));
    jdff dff_B_kjU0WIxU8_1(.din(n11392), .dout(n11395));
    jdff dff_B_m5VZ61L67_1(.din(n11395), .dout(n11398));
    jdff dff_B_hoJsCj2k7_1(.din(n11398), .dout(n11401));
    jdff dff_B_YNt5KqTj9_1(.din(n11401), .dout(n11404));
    jdff dff_B_KrtjcLqM4_1(.din(n11404), .dout(n11407));
    jdff dff_B_cjyca7w44_1(.din(n11407), .dout(n11410));
    jdff dff_B_LMGnYrWV7_1(.din(n11410), .dout(n11413));
    jdff dff_B_D0n8gG373_1(.din(n11413), .dout(n11416));
    jdff dff_B_xustH9JN0_1(.din(n11416), .dout(n11419));
    jdff dff_B_AdciMGAg0_1(.din(n11419), .dout(n11422));
    jdff dff_B_YgVZMix71_1(.din(n11422), .dout(n11425));
    jdff dff_B_2x8z9CsQ3_1(.din(n11425), .dout(n11428));
    jdff dff_B_3R5MpDEX5_1(.din(n11428), .dout(n11431));
    jdff dff_B_MAphkkXz6_1(.din(n11431), .dout(n11434));
    jdff dff_B_tBGD9mXy0_1(.din(n11434), .dout(n11437));
    jdff dff_B_nxywcEQT7_1(.din(n11437), .dout(n11440));
    jdff dff_B_43c16sot3_1(.din(n11440), .dout(n11443));
    jdff dff_B_YOI6Kdlw6_1(.din(n11443), .dout(n11446));
    jdff dff_B_4vog6DFp5_1(.din(n11446), .dout(n11449));
    jdff dff_B_HLRyeS8Z6_1(.din(n11449), .dout(n11452));
    jdff dff_B_YPLgVBAv6_1(.din(n11452), .dout(n11455));
    jdff dff_B_EnAH4Js65_1(.din(n11455), .dout(n11458));
    jdff dff_B_xvFx4mJ55_1(.din(n11458), .dout(n11461));
    jdff dff_B_TTSwfGcV1_1(.din(n11461), .dout(n11464));
    jdff dff_B_5a35RJUv5_1(.din(n11464), .dout(n11467));
    jdff dff_B_IkHbgszW1_1(.din(n11467), .dout(n11470));
    jdff dff_B_OHLiR9ce0_1(.din(n11470), .dout(n11473));
    jdff dff_B_aQJSDXwv1_1(.din(n11473), .dout(n11476));
    jdff dff_B_KEclRy8v4_1(.din(n11476), .dout(n11479));
    jdff dff_B_J6hTIKWU6_1(.din(n11479), .dout(n11482));
    jdff dff_B_1xGOBdgR8_1(.din(n11482), .dout(n11485));
    jdff dff_B_4I22MR9j5_1(.din(n11485), .dout(n11488));
    jdff dff_B_l9Znp2i90_1(.din(n11488), .dout(n11491));
    jdff dff_B_fX6XFwfv2_1(.din(n11491), .dout(n11494));
    jdff dff_B_bhERwpZM9_1(.din(n2596), .dout(n11497));
    jdff dff_B_vounQEKF0_1(.din(n11497), .dout(n11500));
    jdff dff_B_iEe7ZKqG0_1(.din(n11500), .dout(n11503));
    jdff dff_B_E0LBWgmp0_1(.din(n11503), .dout(n11506));
    jdff dff_B_fckmYLXb9_1(.din(n11506), .dout(n11509));
    jdff dff_B_ojD4jv0Q0_1(.din(n11509), .dout(n11512));
    jdff dff_B_0lII4XEZ5_1(.din(n11512), .dout(n11515));
    jdff dff_B_1yEjaGtF8_1(.din(n11515), .dout(n11518));
    jdff dff_B_16CiTP473_1(.din(n11518), .dout(n11521));
    jdff dff_B_GPpO06U95_1(.din(n11521), .dout(n11524));
    jdff dff_B_ywCLCs4H4_1(.din(n11524), .dout(n11527));
    jdff dff_B_cd6ipKFb5_1(.din(n11527), .dout(n11530));
    jdff dff_B_zxKrJ2Hg1_1(.din(n11530), .dout(n11533));
    jdff dff_B_4yU7EuX57_1(.din(n11533), .dout(n11536));
    jdff dff_B_TP0usAbO3_1(.din(n11536), .dout(n11539));
    jdff dff_B_sAXTRqGj2_1(.din(n11539), .dout(n11542));
    jdff dff_B_5ZVIeCy01_1(.din(n11542), .dout(n11545));
    jdff dff_B_gKeN94ss9_1(.din(n11545), .dout(n11548));
    jdff dff_B_mYQ91xFU0_1(.din(n11548), .dout(n11551));
    jdff dff_B_dqyaHDPz6_1(.din(n11551), .dout(n11554));
    jdff dff_B_83rQTowt2_1(.din(n11554), .dout(n11557));
    jdff dff_B_gGVYeCIU3_1(.din(n11557), .dout(n11560));
    jdff dff_B_qegBv0gk7_1(.din(n11560), .dout(n11563));
    jdff dff_B_ljCYe4Mi5_1(.din(n11563), .dout(n11566));
    jdff dff_B_eERNXww16_1(.din(n11566), .dout(n11569));
    jdff dff_B_1j0PqywI6_1(.din(n11569), .dout(n11572));
    jdff dff_B_Fp4hZQj24_1(.din(n11572), .dout(n11575));
    jdff dff_B_Bzd4Gd4G7_1(.din(n11575), .dout(n11578));
    jdff dff_B_IOkKtf9i2_1(.din(n11578), .dout(n11581));
    jdff dff_B_I0WggfyD7_1(.din(n11581), .dout(n11584));
    jdff dff_B_fonbVM4p5_1(.din(n11584), .dout(n11587));
    jdff dff_B_vaq0t36y3_1(.din(n11587), .dout(n11590));
    jdff dff_B_gorOyYwL1_1(.din(n11590), .dout(n11593));
    jdff dff_B_9aONanXf9_1(.din(n11593), .dout(n11596));
    jdff dff_B_VfrXnsV62_1(.din(n11596), .dout(n11599));
    jdff dff_B_Qvl9bDzk3_1(.din(n11599), .dout(n11602));
    jdff dff_B_A2DRuLiV4_1(.din(n11602), .dout(n11605));
    jdff dff_B_pjxF3ZmG0_1(.din(n11605), .dout(n11608));
    jdff dff_B_pCPX82E15_1(.din(n11608), .dout(n11611));
    jdff dff_B_P2cfAhMG6_1(.din(n11611), .dout(n11614));
    jdff dff_B_EcYzZ6w71_1(.din(n2978), .dout(n11617));
    jdff dff_B_wIr2XIFU7_1(.din(n11617), .dout(n11620));
    jdff dff_B_furpVV9k1_1(.din(n11620), .dout(n11623));
    jdff dff_B_QvHf1xwY0_1(.din(n11623), .dout(n11626));
    jdff dff_B_o4u3vI5k6_1(.din(n11626), .dout(n11629));
    jdff dff_B_kHPkxqTA9_1(.din(n11629), .dout(n11632));
    jdff dff_B_obd657vg8_1(.din(n11632), .dout(n11635));
    jdff dff_B_33mIoTbk8_1(.din(n11635), .dout(n11638));
    jdff dff_B_yxBmnghK9_1(.din(n11638), .dout(n11641));
    jdff dff_B_eXX13Pqf2_1(.din(n11641), .dout(n11644));
    jdff dff_B_0ueVHSbU3_1(.din(n11644), .dout(n11647));
    jdff dff_B_k8P4wljZ5_1(.din(n11647), .dout(n11650));
    jdff dff_B_xLEamzwr9_1(.din(n11650), .dout(n11653));
    jdff dff_B_zURI3Hdu6_1(.din(n11653), .dout(n11656));
    jdff dff_B_kYeKGal02_1(.din(n11656), .dout(n11659));
    jdff dff_B_wnEDff3J9_1(.din(n11659), .dout(n11662));
    jdff dff_B_vU0e0Ijl7_1(.din(n11662), .dout(n11665));
    jdff dff_B_TjK5C9pn3_1(.din(n11665), .dout(n11668));
    jdff dff_B_leCVotMu8_1(.din(n11668), .dout(n11671));
    jdff dff_B_Ocyxqbgr9_1(.din(n11671), .dout(n11674));
    jdff dff_B_3u7UaqNw8_1(.din(n11674), .dout(n11677));
    jdff dff_B_2SKH4sBb5_1(.din(n11677), .dout(n11680));
    jdff dff_B_xPcaFZLU2_1(.din(n11680), .dout(n11683));
    jdff dff_B_8S3jPgSq7_1(.din(n11683), .dout(n11686));
    jdff dff_B_vGd5woqt0_1(.din(n11686), .dout(n11689));
    jdff dff_B_ZTvQ8cOR8_1(.din(n11689), .dout(n11692));
    jdff dff_B_PirkwQWd4_1(.din(n11692), .dout(n11695));
    jdff dff_B_jpzYNZOM2_1(.din(n11695), .dout(n11698));
    jdff dff_B_Lg15YytX8_1(.din(n11698), .dout(n11701));
    jdff dff_B_C37td1dx7_1(.din(n11701), .dout(n11704));
    jdff dff_B_L6WtZiIo4_1(.din(n11704), .dout(n11707));
    jdff dff_B_n3S53RUV4_1(.din(n11707), .dout(n11710));
    jdff dff_B_hupLYL7c3_1(.din(n11710), .dout(n11713));
    jdff dff_B_gmBAj38L4_1(.din(n11713), .dout(n11716));
    jdff dff_B_qLJbvFUF3_1(.din(n11716), .dout(n11719));
    jdff dff_B_lMpFMA492_1(.din(n11719), .dout(n11722));
    jdff dff_B_DMuZ9GNp9_1(.din(n11722), .dout(n11725));
    jdff dff_B_eN08a2vV8_1(.din(n11725), .dout(n11728));
    jdff dff_B_TZVngQF69_1(.din(n11728), .dout(n11731));
    jdff dff_B_5aFT5H7H8_1(.din(n11731), .dout(n11734));
    jdff dff_B_AH6MrSp94_1(.din(n11734), .dout(n11737));
    jdff dff_B_fxHsrPUf6_1(.din(n11737), .dout(n11740));
    jdff dff_B_vYOXfILh7_1(.din(n11740), .dout(n11743));
    jdff dff_B_fMoeLlFX7_0(.din(n4882), .dout(n11746));
    jdff dff_B_sbFeo1EI5_1(.din(n6853), .dout(n11749));
    jdff dff_B_2INyUXAH4_1(.din(n11749), .dout(n11752));
    jdff dff_B_zTW8EAQk9_1(.din(n11752), .dout(n11755));
    jdff dff_B_kcolGlWG7_1(.din(n11755), .dout(n11758));
    jdff dff_B_bmKLUEvh2_1(.din(n11758), .dout(n11761));
    jdff dff_B_RwqUbpFi6_1(.din(n11761), .dout(n11764));
    jdff dff_B_ReuhXnQ20_1(.din(n11764), .dout(n11767));
    jdff dff_B_pAVLRkq43_1(.din(n11767), .dout(n11770));
    jdff dff_B_pihkHoxr6_1(.din(n11770), .dout(n11773));
    jdff dff_B_6xtnLTau1_1(.din(n11773), .dout(n11776));
    jdff dff_B_bna7xfMG2_1(.din(n11776), .dout(n11779));
    jdff dff_B_qeId6v1Q8_1(.din(n11779), .dout(n11782));
    jdff dff_B_tEIzL6Si8_1(.din(n11782), .dout(n11785));
    jdff dff_B_hQicRh9g9_0(.din(n6881), .dout(n11788));
    jdff dff_B_Zsh8d9J27_0(.din(n11788), .dout(n11791));
    jdff dff_B_EJ1uPLOd7_0(.din(n11791), .dout(n11794));
    jdff dff_B_49lDF8be5_0(.din(n11794), .dout(n11797));
    jdff dff_B_oubJSXAn0_0(.din(n11797), .dout(n11800));
    jdff dff_B_AgpVtZNU5_0(.din(n11800), .dout(n11803));
    jdff dff_B_aqxE7IaL6_0(.din(n11803), .dout(n11806));
    jdff dff_B_z2OGlrf04_0(.din(n11806), .dout(n11809));
    jdff dff_B_gMnJwXhg9_0(.din(n11809), .dout(n11812));
    jdff dff_B_MHn6vCaL1_0(.din(n11812), .dout(n11815));
    jdff dff_B_lO57ET7m6_0(.din(n11815), .dout(n11818));
    jdff dff_A_m0JjNuvI8_0(.din(n11823), .dout(n11820));
    jdff dff_A_XyLHhIko8_0(.din(n11826), .dout(n11823));
    jdff dff_A_YZyxKGH84_0(.din(n11829), .dout(n11826));
    jdff dff_A_zNE32iKI2_0(.din(n11832), .dout(n11829));
    jdff dff_A_J6oD1eTw0_0(.din(n11835), .dout(n11832));
    jdff dff_A_RzBZ9N197_0(.din(n11838), .dout(n11835));
    jdff dff_A_PbKFL8IP9_0(.din(n11841), .dout(n11838));
    jdff dff_A_w5ljE4UP8_0(.din(n11844), .dout(n11841));
    jdff dff_A_ldpsVJv72_0(.din(n11847), .dout(n11844));
    jdff dff_A_BIR0T2Er1_0(.din(n11850), .dout(n11847));
    jdff dff_A_UOZBiI5q7_0(.din(n11853), .dout(n11850));
    jdff dff_A_AfYw5laX3_0(.din(n6878), .dout(n11853));
    jdff dff_B_tWoZIzdD1_1(.din(n6841), .dout(n11857));
    jdff dff_B_l8E1hQ3o8_1(.din(n11857), .dout(n11860));
    jdff dff_B_iz9aTgB08_2(.din(n6837), .dout(n11863));
    jdff dff_B_bV3ZWcCp4_2(.din(n11863), .dout(n11866));
    jdff dff_B_qTkMv25N4_2(.din(n11866), .dout(n11869));
    jdff dff_B_qYKJNjHM8_2(.din(n11869), .dout(n11872));
    jdff dff_B_ZE0PLiXw4_2(.din(n11872), .dout(n11875));
    jdff dff_B_e7JmlJml1_2(.din(n11875), .dout(n11878));
    jdff dff_B_pSibLW3N1_2(.din(n11878), .dout(n11881));
    jdff dff_B_Xb5OxJb10_2(.din(n11881), .dout(n11884));
    jdff dff_B_2fv4WZuu7_2(.din(n11884), .dout(n11887));
    jdff dff_B_aU7SC2Mt6_2(.din(n11887), .dout(n11890));
    jdff dff_B_AMl8UHIt8_2(.din(n11890), .dout(n11893));
    jdff dff_B_zqxapdLY1_2(.din(n11893), .dout(n11896));
    jdff dff_B_r1kE9BxB6_2(.din(n11896), .dout(n11899));
    jdff dff_B_QatLuJBO0_2(.din(n11899), .dout(n11902));
    jdff dff_B_xgMpC9re1_2(.din(n11902), .dout(n11905));
    jdff dff_B_4XrfGHGV8_2(.din(n11905), .dout(n11908));
    jdff dff_B_tBJTXV7x1_2(.din(n11908), .dout(n11911));
    jdff dff_B_MR6tEHgC4_2(.din(n11911), .dout(n11914));
    jdff dff_B_e34WTH2O3_2(.din(n11914), .dout(n11917));
    jdff dff_B_hUnFkNs61_2(.din(n11917), .dout(n11920));
    jdff dff_B_RnZXvcQH5_2(.din(n11920), .dout(n11923));
    jdff dff_B_7ADFwLpP0_2(.din(n11923), .dout(n11926));
    jdff dff_B_wXScGgMg6_2(.din(n11926), .dout(n11929));
    jdff dff_B_A3sTDcJI9_2(.din(n11929), .dout(n11932));
    jdff dff_B_AUuzRjLB8_2(.din(n11932), .dout(n11935));
    jdff dff_B_3LPsbA4d6_2(.din(n11935), .dout(n11938));
    jdff dff_B_m28lmXxm5_2(.din(n11938), .dout(n11941));
    jdff dff_B_vGvo1yPu8_2(.din(n11941), .dout(n11944));
    jdff dff_B_orcXzQlX1_2(.din(n11944), .dout(n11947));
    jdff dff_B_TW4Lygyl1_2(.din(n11947), .dout(n11950));
    jdff dff_B_NehRVWgf9_2(.din(n11950), .dout(n11953));
    jdff dff_B_k6lnXCH26_2(.din(n11953), .dout(n11956));
    jdff dff_B_mtTvTe6Y9_2(.din(n11956), .dout(n11959));
    jdff dff_B_1Qyk3WNZ6_2(.din(n11959), .dout(n11962));
    jdff dff_B_CtmDnbP80_2(.din(n11962), .dout(n11965));
    jdff dff_B_3t6dei1P1_2(.din(n11965), .dout(n11968));
    jdff dff_B_7uNCo4D26_2(.din(n11968), .dout(n11971));
    jdff dff_B_T8ejGtNS7_2(.din(n11971), .dout(n11974));
    jdff dff_B_Yak9Udtk2_2(.din(n11974), .dout(n11977));
    jdff dff_B_R0LIlpBN7_2(.din(n11977), .dout(n11980));
    jdff dff_B_5SzAzHYS9_2(.din(n11980), .dout(n11983));
    jdff dff_B_ICHowvGj6_2(.din(n11983), .dout(n11986));
    jdff dff_B_J7UtQFDH1_2(.din(n11986), .dout(n11989));
    jdff dff_B_D6Ik5QjN1_2(.din(n11989), .dout(n11992));
    jdff dff_B_PMAbDxLz8_2(.din(n11992), .dout(n11995));
    jdff dff_B_ImRoXffv4_2(.din(n11995), .dout(n11998));
    jdff dff_B_Pftahw966_2(.din(n11998), .dout(n12001));
    jdff dff_B_lG50ej0b4_2(.din(n12001), .dout(n12004));
    jdff dff_B_r4AF2vQW2_2(.din(n12004), .dout(n12007));
    jdff dff_B_uBLBvLJo3_2(.din(n12007), .dout(n12010));
    jdff dff_B_fOJhEY0Y2_2(.din(n12010), .dout(n12013));
    jdff dff_B_ktcPXAgr7_2(.din(n12013), .dout(n12016));
    jdff dff_B_4OKefqFS1_2(.din(n12016), .dout(n12019));
    jdff dff_B_mF1Ktk8h2_2(.din(n12019), .dout(n12022));
    jdff dff_B_FhwPWVkg5_2(.din(n12022), .dout(n12025));
    jdff dff_B_ZRuRRZd25_2(.din(n12025), .dout(n12028));
    jdff dff_B_IgwhY4ht2_2(.din(n12028), .dout(n12031));
    jdff dff_B_rgzkUHGt0_2(.din(n12031), .dout(n12034));
    jdff dff_B_jAPfrKB49_2(.din(n12034), .dout(n12037));
    jdff dff_B_g4xoyXVp5_2(.din(n12037), .dout(n12040));
    jdff dff_B_YAyryhwi7_1(.din(n6863), .dout(n12043));
    jdff dff_B_n8wgVtZu5_1(.din(n12043), .dout(n12046));
    jdff dff_B_CEZXvmhg5_1(.din(n12046), .dout(n12049));
    jdff dff_B_iE86Ry8q4_1(.din(n12049), .dout(n12052));
    jdff dff_B_5Gr5F1uv0_1(.din(n12052), .dout(n12055));
    jdff dff_B_AjkQlkJc1_1(.din(n12055), .dout(n12058));
    jdff dff_B_lVVVOTHN7_1(.din(n12058), .dout(n12061));
    jdff dff_B_YjTJqmDs0_1(.din(n12061), .dout(n12064));
    jdff dff_B_OztWx61B7_1(.din(n12064), .dout(n12067));
    jdff dff_B_GCPIvll60_1(.din(n12067), .dout(n12070));
    jdff dff_B_wJhP7oj49_1(.din(n12070), .dout(n12073));
    jdff dff_B_EMOiCLTU2_0(.din(n6866), .dout(n12076));
    jdff dff_B_VZTT7cji8_0(.din(n12076), .dout(n12079));
    jdff dff_B_DC8U9q976_0(.din(n12079), .dout(n12082));
    jdff dff_B_3YqqsRiB0_0(.din(n12082), .dout(n12085));
    jdff dff_B_t7nv8bQi1_0(.din(n12085), .dout(n12088));
    jdff dff_B_I0yUCq319_0(.din(n12088), .dout(n12091));
    jdff dff_B_7Uv01WtP1_0(.din(n12091), .dout(n12094));
    jdff dff_B_LzStQ3BC8_0(.din(n12094), .dout(n12097));
    jdff dff_B_WmBNDTAf5_0(.din(n12097), .dout(n12100));
    jdff dff_B_4MdSaJGN5_0(.din(n12100), .dout(n12103));
    jdff dff_A_fmIwcrek3_1(.din(n12108), .dout(n12105));
    jdff dff_A_IdGKqR6F6_1(.din(n12111), .dout(n12108));
    jdff dff_A_xkn4FbBm7_1(.din(n12114), .dout(n12111));
    jdff dff_A_sJ43ChCR0_1(.din(n12117), .dout(n12114));
    jdff dff_A_Jnu1htZZ2_1(.din(n12120), .dout(n12117));
    jdff dff_A_2yfFXLks2_1(.din(n12123), .dout(n12120));
    jdff dff_A_ewtxhN3X2_1(.din(n12126), .dout(n12123));
    jdff dff_A_FQo0tz0n9_1(.din(n12129), .dout(n12126));
    jdff dff_A_TaYisTDI2_1(.din(n12132), .dout(n12129));
    jdff dff_A_JC7YBa092_1(.din(n12135), .dout(n12132));
    jdff dff_A_TxFnIYqv4_1(.din(n6829), .dout(n12135));
    jdff dff_B_q6Qq8Sg23_1(.din(n6771), .dout(n12139));
    jdff dff_B_Ay8glTj51_1(.din(n12139), .dout(n12142));
    jdff dff_B_b8Ma6md70_1(.din(n12142), .dout(n12145));
    jdff dff_B_aQi1gvLr0_1(.din(n12145), .dout(n12148));
    jdff dff_B_Ldv37RNC9_1(.din(n12148), .dout(n12151));
    jdff dff_B_4Nq2UBo37_1(.din(n12151), .dout(n12154));
    jdff dff_B_7vTiqso71_1(.din(n12154), .dout(n12157));
    jdff dff_B_gnm77Bmi3_1(.din(n12157), .dout(n12160));
    jdff dff_B_fO3h4D8N1_1(.din(n12160), .dout(n12163));
    jdff dff_B_OClDH2tm0_1(.din(n12163), .dout(n12166));
    jdff dff_B_V4tVImYF3_1(.din(n12166), .dout(n12169));
    jdff dff_B_m15yRGzY6_0(.din(n6774), .dout(n12172));
    jdff dff_B_UBlVmbjq0_0(.din(n12172), .dout(n12175));
    jdff dff_B_uNkVxzEa5_0(.din(n12175), .dout(n12178));
    jdff dff_B_KJL4lO9v3_0(.din(n12178), .dout(n12181));
    jdff dff_B_aPw0MuTd1_0(.din(n12181), .dout(n12184));
    jdff dff_B_rcNnLJ2S1_0(.din(n12184), .dout(n12187));
    jdff dff_B_j4djZjDh0_0(.din(n12187), .dout(n12190));
    jdff dff_B_82Yeytqs9_0(.din(n12190), .dout(n12193));
    jdff dff_B_qkz65yQF3_0(.din(n12193), .dout(n12196));
    jdff dff_B_k03xV37X7_0(.din(n12196), .dout(n12199));
    jdff dff_A_Yy2ZexX11_1(.din(n12204), .dout(n12201));
    jdff dff_A_6sBrAL3t7_1(.din(n12207), .dout(n12204));
    jdff dff_A_9BRfZH5s0_1(.din(n12210), .dout(n12207));
    jdff dff_A_L9cWyI3p3_1(.din(n12213), .dout(n12210));
    jdff dff_A_nIyoYqLH8_1(.din(n12216), .dout(n12213));
    jdff dff_A_dQdlcR7G4_1(.din(n12219), .dout(n12216));
    jdff dff_A_etzBS0ph8_1(.din(n12222), .dout(n12219));
    jdff dff_A_b1nMr4uH3_1(.din(n12225), .dout(n12222));
    jdff dff_A_LTxjtvaL4_1(.din(n12228), .dout(n12225));
    jdff dff_A_PfRSPYNF2_1(.din(n12231), .dout(n12228));
    jdff dff_A_axlC0KEc6_1(.din(n6757), .dout(n12231));
    jdff dff_B_kVPEUSYw5_1(.din(n6672), .dout(n12235));
    jdff dff_B_5l0iSaGZ3_1(.din(n12235), .dout(n12238));
    jdff dff_B_IIk8IVHM1_1(.din(n12238), .dout(n12241));
    jdff dff_B_OrVwB2EW5_1(.din(n12241), .dout(n12244));
    jdff dff_B_jC1WHUIe7_1(.din(n12244), .dout(n12247));
    jdff dff_B_JynPFKln8_1(.din(n12247), .dout(n12250));
    jdff dff_B_KvA4F5B44_1(.din(n12250), .dout(n12253));
    jdff dff_B_aYfYaXIp1_1(.din(n12253), .dout(n12256));
    jdff dff_B_1bzdDDi43_1(.din(n12256), .dout(n12259));
    jdff dff_B_IuZmrOTp9_1(.din(n12259), .dout(n12262));
    jdff dff_B_2lTowDer4_1(.din(n12262), .dout(n12265));
    jdff dff_B_C8qvizap8_0(.din(n6675), .dout(n12268));
    jdff dff_B_lBnjesKo5_0(.din(n12268), .dout(n12271));
    jdff dff_B_jz1RhArz6_0(.din(n12271), .dout(n12274));
    jdff dff_B_CuB6WOtN4_0(.din(n12274), .dout(n12277));
    jdff dff_B_zjvUSenK3_0(.din(n12277), .dout(n12280));
    jdff dff_B_23I54xxa7_0(.din(n12280), .dout(n12283));
    jdff dff_B_LPvYyFpm3_0(.din(n12283), .dout(n12286));
    jdff dff_B_C3nCA6dU3_0(.din(n12286), .dout(n12289));
    jdff dff_B_Y22ZQXVl8_0(.din(n12289), .dout(n12292));
    jdff dff_B_uo9daJrs0_0(.din(n12292), .dout(n12295));
    jdff dff_A_1wWc61pi3_1(.din(n12300), .dout(n12297));
    jdff dff_A_yQ3s8HxE3_1(.din(n12303), .dout(n12300));
    jdff dff_A_bZZlQ63Z6_1(.din(n12306), .dout(n12303));
    jdff dff_A_sJz3lPCI2_1(.din(n12309), .dout(n12306));
    jdff dff_A_AeVnl6g52_1(.din(n12312), .dout(n12309));
    jdff dff_A_ujEWTp711_1(.din(n12315), .dout(n12312));
    jdff dff_A_CjsMYCwH0_1(.din(n12318), .dout(n12315));
    jdff dff_A_3I90hbjW0_1(.din(n12321), .dout(n12318));
    jdff dff_A_P6IelWAb2_1(.din(n12324), .dout(n12321));
    jdff dff_A_6NepZbbQ7_1(.din(n12327), .dout(n12324));
    jdff dff_A_DbyttkQU3_1(.din(n6658), .dout(n12327));
    jdff dff_B_5IpxAz8Z3_1(.din(n6546), .dout(n12331));
    jdff dff_B_vmnqg6ss9_1(.din(n12331), .dout(n12334));
    jdff dff_B_a0HmcnQt4_1(.din(n12334), .dout(n12337));
    jdff dff_B_GDNd8PaH0_1(.din(n12337), .dout(n12340));
    jdff dff_B_Dx47z0606_1(.din(n12340), .dout(n12343));
    jdff dff_B_7y7VD2tk1_1(.din(n12343), .dout(n12346));
    jdff dff_B_RhgaHpNV8_1(.din(n12346), .dout(n12349));
    jdff dff_B_2eVIsDYU4_1(.din(n12349), .dout(n12352));
    jdff dff_B_LpGSaLql7_1(.din(n12352), .dout(n12355));
    jdff dff_B_B6zPzUqH3_1(.din(n12355), .dout(n12358));
    jdff dff_B_wn5H5gc59_1(.din(n12358), .dout(n12361));
    jdff dff_B_SNWo6Qzh0_0(.din(n6549), .dout(n12364));
    jdff dff_B_JCohFOdw7_0(.din(n12364), .dout(n12367));
    jdff dff_B_dBnURjkZ9_0(.din(n12367), .dout(n12370));
    jdff dff_B_KKfS702Q7_0(.din(n12370), .dout(n12373));
    jdff dff_B_SLl5u2BT3_0(.din(n12373), .dout(n12376));
    jdff dff_B_HcmqYFwf9_0(.din(n12376), .dout(n12379));
    jdff dff_B_6ZEM32JD3_0(.din(n12379), .dout(n12382));
    jdff dff_B_2mWIb39J0_0(.din(n12382), .dout(n12385));
    jdff dff_B_nnnlgVky2_0(.din(n12385), .dout(n12388));
    jdff dff_B_pS6Cq4dI7_0(.din(n12388), .dout(n12391));
    jdff dff_A_BL7JtSMX2_1(.din(n12396), .dout(n12393));
    jdff dff_A_gVAvQkw08_1(.din(n12399), .dout(n12396));
    jdff dff_A_OA5pJVT69_1(.din(n12402), .dout(n12399));
    jdff dff_A_19h8PTCo1_1(.din(n12405), .dout(n12402));
    jdff dff_A_L7S2zJkL2_1(.din(n12408), .dout(n12405));
    jdff dff_A_0knXNdyO8_1(.din(n12411), .dout(n12408));
    jdff dff_A_XLhx0YIo9_1(.din(n12414), .dout(n12411));
    jdff dff_A_DjUE5ZZc0_1(.din(n12417), .dout(n12414));
    jdff dff_A_8xz9VRPK9_1(.din(n12420), .dout(n12417));
    jdff dff_A_mHSJJKXo5_1(.din(n12423), .dout(n12420));
    jdff dff_A_RlkqRC6Q9_1(.din(n6532), .dout(n12423));
    jdff dff_B_v6IhuskW6_1(.din(n6393), .dout(n12427));
    jdff dff_B_63Mcjvni8_1(.din(n12427), .dout(n12430));
    jdff dff_B_wWKuo2wb4_1(.din(n12430), .dout(n12433));
    jdff dff_B_Bdhejcms1_1(.din(n12433), .dout(n12436));
    jdff dff_B_E5cBadYg7_1(.din(n12436), .dout(n12439));
    jdff dff_B_kvA1IVVx7_1(.din(n12439), .dout(n12442));
    jdff dff_B_KTiaSrYS3_1(.din(n12442), .dout(n12445));
    jdff dff_B_gdbnzCQD1_1(.din(n12445), .dout(n12448));
    jdff dff_B_YncGPHfT1_1(.din(n12448), .dout(n12451));
    jdff dff_B_g1SETCA08_1(.din(n12451), .dout(n12454));
    jdff dff_B_j8qeHvjW3_1(.din(n12454), .dout(n12457));
    jdff dff_B_NMCqCl6C4_0(.din(n6396), .dout(n12460));
    jdff dff_B_6NwIBqkQ4_0(.din(n12460), .dout(n12463));
    jdff dff_B_C65pYUIX2_0(.din(n12463), .dout(n12466));
    jdff dff_B_VrInQc6Q7_0(.din(n12466), .dout(n12469));
    jdff dff_B_qAXq7WAD6_0(.din(n12469), .dout(n12472));
    jdff dff_B_T8MwLudp5_0(.din(n12472), .dout(n12475));
    jdff dff_B_dDKNL7hr7_0(.din(n12475), .dout(n12478));
    jdff dff_B_NYILoQxo0_0(.din(n12478), .dout(n12481));
    jdff dff_B_plAUKf9m5_0(.din(n12481), .dout(n12484));
    jdff dff_A_JDqsIVPy3_1(.din(n12489), .dout(n12486));
    jdff dff_A_9Rl5Nb2Z0_1(.din(n12492), .dout(n12489));
    jdff dff_A_3yhR6Yn71_1(.din(n12495), .dout(n12492));
    jdff dff_A_FZKJHNdz8_1(.din(n12498), .dout(n12495));
    jdff dff_A_pe6LVOie1_1(.din(n12501), .dout(n12498));
    jdff dff_A_PRTjnTu04_1(.din(n12504), .dout(n12501));
    jdff dff_A_mwh0BfB78_1(.din(n12507), .dout(n12504));
    jdff dff_A_ho26mdp31_1(.din(n12510), .dout(n12507));
    jdff dff_A_G9YDQs7A9_1(.din(n12513), .dout(n12510));
    jdff dff_A_mHhCd8B79_1(.din(n6385), .dout(n12513));
    jdff dff_B_wn7ZCnbN9_1(.din(n6210), .dout(n12517));
    jdff dff_B_dn4JiUK64_1(.din(n12517), .dout(n12520));
    jdff dff_B_VUJCs6ZS0_1(.din(n12520), .dout(n12523));
    jdff dff_B_OrD85vZy6_1(.din(n12523), .dout(n12526));
    jdff dff_B_zEJMwPul2_1(.din(n12526), .dout(n12529));
    jdff dff_B_OWdu6gAX7_1(.din(n12529), .dout(n12532));
    jdff dff_B_w5AIDrQX9_1(.din(n12532), .dout(n12535));
    jdff dff_B_4mhNrqrI1_1(.din(n12535), .dout(n12538));
    jdff dff_B_OK4ySXev2_1(.din(n12538), .dout(n12541));
    jdff dff_B_J3ei1HvP0_1(.din(n12541), .dout(n12544));
    jdff dff_B_zqYyVafT0_0(.din(n6213), .dout(n12547));
    jdff dff_B_yFBrxJni0_0(.din(n12547), .dout(n12550));
    jdff dff_B_UQIfRW0B4_0(.din(n12550), .dout(n12553));
    jdff dff_B_73QqV5xQ9_0(.din(n12553), .dout(n12556));
    jdff dff_B_U7IAGtya2_0(.din(n12556), .dout(n12559));
    jdff dff_B_T6fUOHGE2_0(.din(n12559), .dout(n12562));
    jdff dff_B_Qh64Slzd2_0(.din(n12562), .dout(n12565));
    jdff dff_B_hwj8yCsY3_0(.din(n12565), .dout(n12568));
    jdff dff_A_PEMtf3vg5_1(.din(n12573), .dout(n12570));
    jdff dff_A_Cdu3USMO5_1(.din(n12576), .dout(n12573));
    jdff dff_A_zhX2MfbU8_1(.din(n12579), .dout(n12576));
    jdff dff_A_LFvGuECz9_1(.din(n12582), .dout(n12579));
    jdff dff_A_niCj6BqO6_1(.din(n12585), .dout(n12582));
    jdff dff_A_jxK1qrBp5_1(.din(n12588), .dout(n12585));
    jdff dff_A_eQCJCu5d0_1(.din(n12591), .dout(n12588));
    jdff dff_A_uuOsS5Nl6_1(.din(n12594), .dout(n12591));
    jdff dff_A_alqW54nR6_1(.din(n6202), .dout(n12594));
    jdff dff_B_hDIJRorC0_1(.din(n6000), .dout(n12598));
    jdff dff_B_XYhI3q5R6_1(.din(n12598), .dout(n12601));
    jdff dff_B_IT6zoV182_1(.din(n12601), .dout(n12604));
    jdff dff_B_91PgArA15_1(.din(n12604), .dout(n12607));
    jdff dff_B_hREdb58u6_1(.din(n12607), .dout(n12610));
    jdff dff_B_MWc4OmHJ5_1(.din(n12610), .dout(n12613));
    jdff dff_B_rK8WkAaj8_1(.din(n12613), .dout(n12616));
    jdff dff_B_BN5B8V2h3_1(.din(n12616), .dout(n12619));
    jdff dff_B_QPdpzU6K2_1(.din(n12619), .dout(n12622));
    jdff dff_B_LL8oMdvo3_1(.din(n12622), .dout(n12625));
    jdff dff_B_IYlB5aSd1_0(.din(n6003), .dout(n12628));
    jdff dff_B_ZTaSJ6TW1_0(.din(n12628), .dout(n12631));
    jdff dff_B_jdmB6ANR4_0(.din(n12631), .dout(n12634));
    jdff dff_B_3PQFhNu23_0(.din(n12634), .dout(n12637));
    jdff dff_B_Y0oZyQIu9_0(.din(n12637), .dout(n12640));
    jdff dff_B_N3LBxeXa8_0(.din(n12640), .dout(n12643));
    jdff dff_B_YGbr3H580_0(.din(n12643), .dout(n12646));
    jdff dff_B_UtgNrEWs9_0(.din(n12646), .dout(n12649));
    jdff dff_A_vqWjPbkR0_1(.din(n12654), .dout(n12651));
    jdff dff_A_fQ4eruGN5_1(.din(n12657), .dout(n12654));
    jdff dff_A_5M2X4v0J2_1(.din(n12660), .dout(n12657));
    jdff dff_A_2OamhUUX4_1(.din(n12663), .dout(n12660));
    jdff dff_A_iwFPN9Lb6_1(.din(n12666), .dout(n12663));
    jdff dff_A_OHdBHNXF9_1(.din(n12669), .dout(n12666));
    jdff dff_A_l60AQmtu6_1(.din(n12672), .dout(n12669));
    jdff dff_A_kro1kpmS6_1(.din(n12675), .dout(n12672));
    jdff dff_A_1K1g5fbW6_1(.din(n5992), .dout(n12675));
    jdff dff_B_qThZXVAS5_1(.din(n5763), .dout(n12679));
    jdff dff_B_4KsNT68r4_1(.din(n12679), .dout(n12682));
    jdff dff_B_m0321h2C0_1(.din(n12682), .dout(n12685));
    jdff dff_B_AtHV9SqQ6_1(.din(n12685), .dout(n12688));
    jdff dff_B_1taZFBdh8_1(.din(n12688), .dout(n12691));
    jdff dff_B_ZuRuUN8X6_1(.din(n12691), .dout(n12694));
    jdff dff_B_RNNhOt3S1_1(.din(n12694), .dout(n12697));
    jdff dff_B_PaiXs0mt7_1(.din(n12697), .dout(n12700));
    jdff dff_B_tH6DKS5D0_0(.din(n5766), .dout(n12703));
    jdff dff_B_wAzPyPXZ1_0(.din(n12703), .dout(n12706));
    jdff dff_B_453u6ucA1_0(.din(n12706), .dout(n12709));
    jdff dff_B_KBA9Z8uR9_0(.din(n12709), .dout(n12712));
    jdff dff_B_eK1Ui84y8_0(.din(n12712), .dout(n12715));
    jdff dff_B_qqrw33Vf4_0(.din(n12715), .dout(n12718));
    jdff dff_A_sBMcs55T8_1(.din(n12723), .dout(n12720));
    jdff dff_A_fyj4QY1o3_1(.din(n12726), .dout(n12723));
    jdff dff_A_oxyUvhSv3_1(.din(n12729), .dout(n12726));
    jdff dff_A_aaetnem01_1(.din(n12732), .dout(n12729));
    jdff dff_A_Bw5tnDwG9_1(.din(n12735), .dout(n12732));
    jdff dff_A_vFKT07tG1_1(.din(n12738), .dout(n12735));
    jdff dff_A_0GFTuX1r9_1(.din(n5755), .dout(n12738));
    jdff dff_B_89zGTgIV5_1(.din(n5499), .dout(n12742));
    jdff dff_B_tbNkuEda9_1(.din(n12742), .dout(n12745));
    jdff dff_B_Lf1hSQTd4_1(.din(n12745), .dout(n12748));
    jdff dff_B_B7Y8Xqzg5_1(.din(n12748), .dout(n12751));
    jdff dff_B_sipoZOv55_1(.din(n12751), .dout(n12754));
    jdff dff_B_I6yWBDMP5_1(.din(n12754), .dout(n12757));
    jdff dff_B_uM7kyvMl1_1(.din(n12757), .dout(n12760));
    jdff dff_B_BOAjz2Gm4_0(.din(n5502), .dout(n12763));
    jdff dff_B_NlqWlu6X0_0(.din(n12763), .dout(n12766));
    jdff dff_B_NBYt3pqa5_0(.din(n12766), .dout(n12769));
    jdff dff_B_WfTwraRJ8_0(.din(n12769), .dout(n12772));
    jdff dff_B_fW2lPW9w3_0(.din(n12772), .dout(n12775));
    jdff dff_A_YyE8LCpd2_1(.din(n12780), .dout(n12777));
    jdff dff_A_kyqDLJ360_1(.din(n12783), .dout(n12780));
    jdff dff_A_yVVeluAA9_1(.din(n12786), .dout(n12783));
    jdff dff_A_BK3FG69W3_1(.din(n12789), .dout(n12786));
    jdff dff_A_bd6lX0Qc8_1(.din(n12792), .dout(n12789));
    jdff dff_A_aEBeq1PX8_1(.din(n5491), .dout(n12792));
    jdff dff_B_7YPz0EEJ5_1(.din(n5208), .dout(n12796));
    jdff dff_B_vSqMAagr0_1(.din(n12796), .dout(n12799));
    jdff dff_B_g1EjlE8T9_1(.din(n12799), .dout(n12802));
    jdff dff_B_UukhTS6B9_1(.din(n12802), .dout(n12805));
    jdff dff_B_TnCH5q7Z6_1(.din(n12805), .dout(n12808));
    jdff dff_B_WWr6rpmz9_1(.din(n12808), .dout(n12811));
    jdff dff_B_fwtVPQSN3_0(.din(n5211), .dout(n12814));
    jdff dff_B_od5UusqG5_0(.din(n12814), .dout(n12817));
    jdff dff_B_L58Alc1U3_0(.din(n12817), .dout(n12820));
    jdff dff_B_RMHEEMGh8_0(.din(n12820), .dout(n12823));
    jdff dff_A_icapOvkN0_1(.din(n12828), .dout(n12825));
    jdff dff_A_Dh0iTn9n1_1(.din(n12831), .dout(n12828));
    jdff dff_A_00RSsezR6_1(.din(n12834), .dout(n12831));
    jdff dff_A_adH5Mp8P7_1(.din(n12837), .dout(n12834));
    jdff dff_A_VznJHwpx9_1(.din(n5200), .dout(n12837));
    jdff dff_B_EaACql833_1(.din(n4893), .dout(n12841));
    jdff dff_B_CNq2ygGW5_1(.din(n12841), .dout(n12844));
    jdff dff_B_3s0PRdKJ2_1(.din(n12844), .dout(n12847));
    jdff dff_A_MOiX7ir23_0(.din(n12852), .dout(n12849));
    jdff dff_A_K4ToNhLz9_0(.din(n4879), .dout(n12852));
    jdff dff_B_BFNl21zT8_1(.din(n4554), .dout(n12856));
    jdff dff_A_8LRjp0fZ3_0(.din(n4540), .dout(n12858));
    jdff dff_B_YxY9L11J6_1(.din(n4183), .dout(n12862));
    jdff dff_A_BLchi0CF4_1(.din(n3778), .dout(n12864));
    jdff dff_B_6NEy3HGz2_2(.din(n3770), .dout(n12868));
    jdff dff_B_uKVEnDbQ2_1(.din(n3380), .dout(n12871));
    jdff dff_A_6V7hrwzn6_0(.din(n12876), .dout(n12873));
    jdff dff_A_fNxtcm6l6_0(.din(n12879), .dout(n12876));
    jdff dff_A_6F0XgFpA4_0(.din(n12882), .dout(n12879));
    jdff dff_A_J44bVdcI7_0(.din(n12885), .dout(n12882));
    jdff dff_A_psvP85Nc8_0(.din(n12888), .dout(n12885));
    jdff dff_A_svKF7qMX4_0(.din(n12891), .dout(n12888));
    jdff dff_A_ceoaJjlg4_0(.din(n12894), .dout(n12891));
    jdff dff_A_uMh3wmh43_0(.din(n12897), .dout(n12894));
    jdff dff_A_W9TbWtlx1_0(.din(n12900), .dout(n12897));
    jdff dff_A_56uq5eD56_0(.din(n12903), .dout(n12900));
    jdff dff_A_pk7oJCgU3_0(.din(n12906), .dout(n12903));
    jdff dff_A_OWeYt4PU1_0(.din(n12909), .dout(n12906));
    jdff dff_A_BRlYgQwf5_0(.din(n12912), .dout(n12909));
    jdff dff_A_lXeA3x2S5_0(.din(n12915), .dout(n12912));
    jdff dff_A_izlyF6sL0_0(.din(n12918), .dout(n12915));
    jdff dff_A_8v87OChG1_0(.din(n12921), .dout(n12918));
    jdff dff_A_Q37cT2OV6_0(.din(n12924), .dout(n12921));
    jdff dff_A_8lR8qIBP6_0(.din(n12927), .dout(n12924));
    jdff dff_A_f2ymBBmN9_0(.din(n12930), .dout(n12927));
    jdff dff_A_uwxDyZH07_0(.din(n12933), .dout(n12930));
    jdff dff_A_TaJiwgA97_0(.din(n12936), .dout(n12933));
    jdff dff_A_JsTOEFvp2_0(.din(n12939), .dout(n12936));
    jdff dff_A_5XoUr31V9_0(.din(n12942), .dout(n12939));
    jdff dff_A_s2FCC40a3_0(.din(n12945), .dout(n12942));
    jdff dff_A_rCDjsYt57_0(.din(n12948), .dout(n12945));
    jdff dff_A_6XcoHjrL7_0(.din(n12951), .dout(n12948));
    jdff dff_A_plIe5c5R0_0(.din(n12954), .dout(n12951));
    jdff dff_A_lXIm4D0B8_0(.din(n12957), .dout(n12954));
    jdff dff_A_cjOmuz7j2_0(.din(n12960), .dout(n12957));
    jdff dff_A_MQJ1NTqI4_0(.din(n12963), .dout(n12960));
    jdff dff_A_6pA4xgLf6_0(.din(n12966), .dout(n12963));
    jdff dff_A_AVj3Kxvt1_0(.din(n12969), .dout(n12966));
    jdff dff_A_riwt5X847_0(.din(n12972), .dout(n12969));
    jdff dff_A_hQVe51HY8_0(.din(n12975), .dout(n12972));
    jdff dff_A_CT7W2dHd3_0(.din(n12978), .dout(n12975));
    jdff dff_A_lHUiqZYq7_0(.din(n12981), .dout(n12978));
    jdff dff_A_0DwLaxM29_0(.din(n12984), .dout(n12981));
    jdff dff_A_cvpYQpNF5_0(.din(n12987), .dout(n12984));
    jdff dff_A_K5Az5ea85_0(.din(n12990), .dout(n12987));
    jdff dff_A_9jw0b8U63_0(.din(n12993), .dout(n12990));
    jdff dff_A_UJ9I5hKy2_0(.din(n12996), .dout(n12993));
    jdff dff_A_0ZD60s2I6_0(.din(n12999), .dout(n12996));
    jdff dff_A_6Qm3LNbZ2_0(.din(n13002), .dout(n12999));
    jdff dff_A_4Cy19Jzl6_0(.din(n2975), .dout(n13002));
    jdff dff_A_nNe7f8Xx0_1(.din(n3365), .dout(n13005));
    jdff dff_B_cm5qEtPD6_1(.din(n2985), .dout(n13009));
    jdff dff_A_hpkQO7MK5_0(.din(n13014), .dout(n13011));
    jdff dff_A_S0gkK6by2_0(.din(n13017), .dout(n13014));
    jdff dff_A_wv30d5M87_0(.din(n13020), .dout(n13017));
    jdff dff_A_l5LiC6On9_0(.din(n13023), .dout(n13020));
    jdff dff_A_x8gfXW7k9_0(.din(n13026), .dout(n13023));
    jdff dff_A_sZ1guD3X8_0(.din(n13029), .dout(n13026));
    jdff dff_A_AMEnIHwt7_0(.din(n13032), .dout(n13029));
    jdff dff_A_XOlSkgMJ2_0(.din(n13035), .dout(n13032));
    jdff dff_A_BYrGcG2S3_0(.din(n13038), .dout(n13035));
    jdff dff_A_QEu5ft5c4_0(.din(n13041), .dout(n13038));
    jdff dff_A_4dHJ5FnO9_0(.din(n13044), .dout(n13041));
    jdff dff_A_0qZAWYTK7_0(.din(n13047), .dout(n13044));
    jdff dff_A_uF596t8g2_0(.din(n13050), .dout(n13047));
    jdff dff_A_ijqfPpKd9_0(.din(n13053), .dout(n13050));
    jdff dff_A_Ug3QQrpa5_0(.din(n13056), .dout(n13053));
    jdff dff_A_ZR61NCGG8_0(.din(n13059), .dout(n13056));
    jdff dff_A_v4Ozbc4b5_0(.din(n13062), .dout(n13059));
    jdff dff_A_WwPIPAVl7_0(.din(n13065), .dout(n13062));
    jdff dff_A_gb66Bs6G0_0(.din(n13068), .dout(n13065));
    jdff dff_A_uFyblmZr5_0(.din(n13071), .dout(n13068));
    jdff dff_A_jzHJH7ng6_0(.din(n13074), .dout(n13071));
    jdff dff_A_kvrYy2i36_0(.din(n13077), .dout(n13074));
    jdff dff_A_5bfFOKNy9_0(.din(n13080), .dout(n13077));
    jdff dff_A_YTXbspCj6_0(.din(n13083), .dout(n13080));
    jdff dff_A_QbgmQ9GR0_0(.din(n13086), .dout(n13083));
    jdff dff_A_DWtzE9Lg9_0(.din(n13089), .dout(n13086));
    jdff dff_A_rD2ES1qK5_0(.din(n13092), .dout(n13089));
    jdff dff_A_M8jWDMan9_0(.din(n13095), .dout(n13092));
    jdff dff_A_D9l9qJ8J3_0(.din(n13098), .dout(n13095));
    jdff dff_A_hd2BDvex8_0(.din(n13101), .dout(n13098));
    jdff dff_A_pQIeJ1yR6_0(.din(n13104), .dout(n13101));
    jdff dff_A_3nxdof6H0_0(.din(n13107), .dout(n13104));
    jdff dff_A_j3UuPga36_0(.din(n13110), .dout(n13107));
    jdff dff_A_jnYUxKz76_0(.din(n13113), .dout(n13110));
    jdff dff_A_s9qkdFRi6_0(.din(n13116), .dout(n13113));
    jdff dff_A_0Qx3SRCO8_0(.din(n13119), .dout(n13116));
    jdff dff_A_uknZAKxN2_0(.din(n13122), .dout(n13119));
    jdff dff_A_jIWh811E7_0(.din(n13125), .dout(n13122));
    jdff dff_A_CDbqx1dQ0_0(.din(n13128), .dout(n13125));
    jdff dff_A_zTPZjg254_0(.din(n13131), .dout(n13128));
    jdff dff_A_O44AF8rm8_0(.din(n2593), .dout(n13131));
    jdff dff_A_ve3QpJuC3_1(.din(n2963), .dout(n13134));
    jdff dff_B_L99dMJIv6_1(.din(n2618), .dout(n13138));
    jdff dff_B_KKp1gkxY3_1(.din(n13138), .dout(n13141));
    jdff dff_B_OprdLYLo0_1(.din(n13141), .dout(n13144));
    jdff dff_B_76Lwyahd0_1(.din(n13144), .dout(n13147));
    jdff dff_B_bwVhD8xL5_1(.din(n13147), .dout(n13150));
    jdff dff_B_c9FhlcRE6_1(.din(n13150), .dout(n13153));
    jdff dff_B_db3vdHwX2_1(.din(n13153), .dout(n13156));
    jdff dff_B_TzrojeaV2_1(.din(n13156), .dout(n13159));
    jdff dff_B_OdyuZ8aR4_1(.din(n13159), .dout(n13162));
    jdff dff_B_OtluU48w3_1(.din(n13162), .dout(n13165));
    jdff dff_B_1rwJXIys4_1(.din(n13165), .dout(n13168));
    jdff dff_B_yNTuvNMC9_1(.din(n13168), .dout(n13171));
    jdff dff_B_O7B3LFZ33_1(.din(n13171), .dout(n13174));
    jdff dff_B_Dt2BYe0z8_1(.din(n13174), .dout(n13177));
    jdff dff_B_bph5RScJ6_1(.din(n13177), .dout(n13180));
    jdff dff_B_srYuAKkj3_1(.din(n13180), .dout(n13183));
    jdff dff_B_22bIZSn63_1(.din(n13183), .dout(n13186));
    jdff dff_B_lYRTQzSs5_1(.din(n13186), .dout(n13189));
    jdff dff_B_hcq8z5Yw5_1(.din(n13189), .dout(n13192));
    jdff dff_B_5PdSpXBM8_1(.din(n13192), .dout(n13195));
    jdff dff_B_o3oBp1mo1_1(.din(n13195), .dout(n13198));
    jdff dff_B_eEfCfQXT7_1(.din(n13198), .dout(n13201));
    jdff dff_B_HTVDmjNe4_1(.din(n13201), .dout(n13204));
    jdff dff_B_bA9Iry2k2_1(.din(n13204), .dout(n13207));
    jdff dff_B_xcpF8nml9_1(.din(n13207), .dout(n13210));
    jdff dff_B_OyxFWTsp4_1(.din(n13210), .dout(n13213));
    jdff dff_B_qoWgq2Zp2_1(.din(n13213), .dout(n13216));
    jdff dff_B_u6EardZn0_1(.din(n13216), .dout(n13219));
    jdff dff_B_of8g8xc52_1(.din(n13219), .dout(n13222));
    jdff dff_B_Qasj3y822_1(.din(n13222), .dout(n13225));
    jdff dff_B_g0HV2ilx8_1(.din(n13225), .dout(n13228));
    jdff dff_B_A5sm3Avt5_1(.din(n13228), .dout(n13231));
    jdff dff_B_xuTN1zfU2_1(.din(n13231), .dout(n13234));
    jdff dff_B_0NtVP1NK5_1(.din(n13234), .dout(n13237));
    jdff dff_B_gZlEn6vm6_1(.din(n13237), .dout(n13240));
    jdff dff_B_VyAkWJzf9_1(.din(n13240), .dout(n13243));
    jdff dff_B_6piPLQWx6_1(.din(n13243), .dout(n13246));
    jdff dff_B_XehIwMva3_1(.din(n2603), .dout(n13249));
    jdff dff_A_dkFBMNyd3_0(.din(n13254), .dout(n13251));
    jdff dff_A_IYbI70kl3_0(.din(n13257), .dout(n13254));
    jdff dff_A_RV4KjewY1_0(.din(n13260), .dout(n13257));
    jdff dff_A_AD3xpUNw8_0(.din(n13263), .dout(n13260));
    jdff dff_A_pZk4GdOh0_0(.din(n13266), .dout(n13263));
    jdff dff_A_T0CF8oMq8_0(.din(n13269), .dout(n13266));
    jdff dff_A_eUxaKqhA6_0(.din(n13272), .dout(n13269));
    jdff dff_A_FHxmToAu5_0(.din(n13275), .dout(n13272));
    jdff dff_A_QsmErd6W4_0(.din(n13278), .dout(n13275));
    jdff dff_A_MnpNT35V7_0(.din(n13281), .dout(n13278));
    jdff dff_A_aQIKJJWY2_0(.din(n13284), .dout(n13281));
    jdff dff_A_51EP7Rqb8_0(.din(n13287), .dout(n13284));
    jdff dff_A_DPrAYKxd9_0(.din(n13290), .dout(n13287));
    jdff dff_A_BJjSs7Ka8_0(.din(n13293), .dout(n13290));
    jdff dff_A_6lMKKesw8_0(.din(n13296), .dout(n13293));
    jdff dff_A_oII8ASb93_0(.din(n13299), .dout(n13296));
    jdff dff_A_5vYfnKTv1_0(.din(n13302), .dout(n13299));
    jdff dff_A_TObYhCgW7_0(.din(n13305), .dout(n13302));
    jdff dff_A_0DYMsleC5_0(.din(n13308), .dout(n13305));
    jdff dff_A_fhKsflu15_0(.din(n13311), .dout(n13308));
    jdff dff_A_6DrtfXqu5_0(.din(n13314), .dout(n13311));
    jdff dff_A_yL4F9Vsb6_0(.din(n13317), .dout(n13314));
    jdff dff_A_waY3hmgA8_0(.din(n13320), .dout(n13317));
    jdff dff_A_KBExpihi0_0(.din(n13323), .dout(n13320));
    jdff dff_A_YskG4wLk4_0(.din(n13326), .dout(n13323));
    jdff dff_A_qpxTXPI91_0(.din(n13329), .dout(n13326));
    jdff dff_A_QwLV5MNt0_0(.din(n13332), .dout(n13329));
    jdff dff_A_xzuvi9cr1_0(.din(n13335), .dout(n13332));
    jdff dff_A_deE9DqQJ7_0(.din(n13338), .dout(n13335));
    jdff dff_A_KaBZbPk31_0(.din(n13341), .dout(n13338));
    jdff dff_A_OkqWzp1N0_0(.din(n13344), .dout(n13341));
    jdff dff_A_Ofu4lpNa4_0(.din(n13347), .dout(n13344));
    jdff dff_A_MQKVLyyw0_0(.din(n13350), .dout(n13347));
    jdff dff_A_I2smT1Jo3_0(.din(n13353), .dout(n13350));
    jdff dff_A_W7hnBpyI7_0(.din(n13356), .dout(n13353));
    jdff dff_A_bLF0rPgD2_0(.din(n13359), .dout(n13356));
    jdff dff_A_4iRi0tfL7_0(.din(n13362), .dout(n13359));
    jdff dff_A_MyPZGV0G3_0(.din(n2238), .dout(n13362));
    jdff dff_A_hATT4C2w2_1(.din(n2581), .dout(n13365));
    jdff dff_B_YKDZx7fy4_1(.din(n2263), .dout(n13369));
    jdff dff_B_30CAmLrj8_1(.din(n13369), .dout(n13372));
    jdff dff_B_0YaJDvfN2_1(.din(n13372), .dout(n13375));
    jdff dff_B_xYO3EXLV4_1(.din(n13375), .dout(n13378));
    jdff dff_B_YRhavu0M3_1(.din(n13378), .dout(n13381));
    jdff dff_B_gWiVubG23_1(.din(n13381), .dout(n13384));
    jdff dff_B_h6IxwEcD2_1(.din(n13384), .dout(n13387));
    jdff dff_B_o8F9vjcx2_1(.din(n13387), .dout(n13390));
    jdff dff_B_rd95D0NW5_1(.din(n13390), .dout(n13393));
    jdff dff_B_f2dDuNHD4_1(.din(n13393), .dout(n13396));
    jdff dff_B_6UVGXx0J7_1(.din(n13396), .dout(n13399));
    jdff dff_B_zzhPxBZM3_1(.din(n13399), .dout(n13402));
    jdff dff_B_Le6VQwOB4_1(.din(n13402), .dout(n13405));
    jdff dff_B_ViuBbaOd0_1(.din(n13405), .dout(n13408));
    jdff dff_B_8AZluf0v6_1(.din(n13408), .dout(n13411));
    jdff dff_B_JUi4qjU18_1(.din(n13411), .dout(n13414));
    jdff dff_B_JtZdrjT47_1(.din(n13414), .dout(n13417));
    jdff dff_B_B4lfhRrp4_1(.din(n13417), .dout(n13420));
    jdff dff_B_ebo5fi4h9_1(.din(n13420), .dout(n13423));
    jdff dff_B_Zr7omRJh7_1(.din(n13423), .dout(n13426));
    jdff dff_B_2K1G3JGf0_1(.din(n13426), .dout(n13429));
    jdff dff_B_UuRafueM8_1(.din(n13429), .dout(n13432));
    jdff dff_B_jkTLqjWb8_1(.din(n13432), .dout(n13435));
    jdff dff_B_hMUURlBV9_1(.din(n13435), .dout(n13438));
    jdff dff_B_WbWycBrW8_1(.din(n13438), .dout(n13441));
    jdff dff_B_ItSywzld8_1(.din(n13441), .dout(n13444));
    jdff dff_B_ItYAKeDP6_1(.din(n13444), .dout(n13447));
    jdff dff_B_ogltcAiF7_1(.din(n13447), .dout(n13450));
    jdff dff_B_sz1Trnej1_1(.din(n13450), .dout(n13453));
    jdff dff_B_Tqtrvtr68_1(.din(n13453), .dout(n13456));
    jdff dff_B_5KlUi48L2_1(.din(n13456), .dout(n13459));
    jdff dff_B_mFQJulWB4_1(.din(n13459), .dout(n13462));
    jdff dff_B_MA7cwNGm2_1(.din(n13462), .dout(n13465));
    jdff dff_B_gR0O5Ao48_1(.din(n13465), .dout(n13468));
    jdff dff_B_ycRlJSps1_1(.din(n2248), .dout(n13471));
    jdff dff_A_p7GUuktE2_0(.din(n13476), .dout(n13473));
    jdff dff_A_WHpTdWff5_0(.din(n13479), .dout(n13476));
    jdff dff_A_XCfgdy1a4_0(.din(n13482), .dout(n13479));
    jdff dff_A_DRj5AaGN2_0(.din(n13485), .dout(n13482));
    jdff dff_A_94I3XL4l4_0(.din(n13488), .dout(n13485));
    jdff dff_A_yy9zWcg31_0(.din(n13491), .dout(n13488));
    jdff dff_A_JeXyUzJI4_0(.din(n13494), .dout(n13491));
    jdff dff_A_p4iV8HMX0_0(.din(n13497), .dout(n13494));
    jdff dff_A_fPsliYym6_0(.din(n13500), .dout(n13497));
    jdff dff_A_ZKMmuNkq9_0(.din(n13503), .dout(n13500));
    jdff dff_A_gwudE4ZE6_0(.din(n13506), .dout(n13503));
    jdff dff_A_9io5mtJi6_0(.din(n13509), .dout(n13506));
    jdff dff_A_yYey6hKF0_0(.din(n13512), .dout(n13509));
    jdff dff_A_ZC2toaYY2_0(.din(n13515), .dout(n13512));
    jdff dff_A_I5CCOEl28_0(.din(n13518), .dout(n13515));
    jdff dff_A_Q1PIakiP2_0(.din(n13521), .dout(n13518));
    jdff dff_A_HoZCIjjc0_0(.din(n13524), .dout(n13521));
    jdff dff_A_gBioCk720_0(.din(n13527), .dout(n13524));
    jdff dff_A_fiU2mHFd9_0(.din(n13530), .dout(n13527));
    jdff dff_A_Gb6RctpV2_0(.din(n13533), .dout(n13530));
    jdff dff_A_A3rKjPti5_0(.din(n13536), .dout(n13533));
    jdff dff_A_8ueIGBPZ8_0(.din(n13539), .dout(n13536));
    jdff dff_A_MhypBxVz4_0(.din(n13542), .dout(n13539));
    jdff dff_A_PXkaP1gN3_0(.din(n13545), .dout(n13542));
    jdff dff_A_lTvnh4hg6_0(.din(n13548), .dout(n13545));
    jdff dff_A_401zNE1z2_0(.din(n13551), .dout(n13548));
    jdff dff_A_HiI0Rbrh6_0(.din(n13554), .dout(n13551));
    jdff dff_A_yB0SWjtR4_0(.din(n13557), .dout(n13554));
    jdff dff_A_BtnbUn9A9_0(.din(n13560), .dout(n13557));
    jdff dff_A_wYQVAkQO0_0(.din(n13563), .dout(n13560));
    jdff dff_A_CyWGjM0H9_0(.din(n13566), .dout(n13563));
    jdff dff_A_KQhmwlZn2_0(.din(n13569), .dout(n13566));
    jdff dff_A_3WzrqVap0_0(.din(n13572), .dout(n13569));
    jdff dff_A_AS5QDOLL6_0(.din(n13575), .dout(n13572));
    jdff dff_A_U6tTMT4n6_0(.din(n1910), .dout(n13575));
    jdff dff_A_aPxlJXc64_1(.din(n2226), .dout(n13578));
    jdff dff_B_iy31NKBE3_1(.din(n1935), .dout(n13582));
    jdff dff_B_RTB9HEF04_1(.din(n13582), .dout(n13585));
    jdff dff_B_I7c2d6g67_1(.din(n13585), .dout(n13588));
    jdff dff_B_gBizV6y55_1(.din(n13588), .dout(n13591));
    jdff dff_B_a2aYoDrQ9_1(.din(n13591), .dout(n13594));
    jdff dff_B_TBDvLm7N3_1(.din(n13594), .dout(n13597));
    jdff dff_B_IqOAo8VR3_1(.din(n13597), .dout(n13600));
    jdff dff_B_OSVZOmad4_1(.din(n13600), .dout(n13603));
    jdff dff_B_zCNee9JC4_1(.din(n13603), .dout(n13606));
    jdff dff_B_4ver7lNm3_1(.din(n13606), .dout(n13609));
    jdff dff_B_uiigXH6p4_1(.din(n13609), .dout(n13612));
    jdff dff_B_8VcGRPQe1_1(.din(n13612), .dout(n13615));
    jdff dff_B_Vxa46z4X8_1(.din(n13615), .dout(n13618));
    jdff dff_B_nnl1cWl62_1(.din(n13618), .dout(n13621));
    jdff dff_B_SEmewUDT4_1(.din(n13621), .dout(n13624));
    jdff dff_B_T4XHIcec4_1(.din(n13624), .dout(n13627));
    jdff dff_B_sKOzv35U8_1(.din(n13627), .dout(n13630));
    jdff dff_B_yEvHS9qk0_1(.din(n13630), .dout(n13633));
    jdff dff_B_Ips5b0QF2_1(.din(n13633), .dout(n13636));
    jdff dff_B_UWKtcUi81_1(.din(n13636), .dout(n13639));
    jdff dff_B_L4HA2sbK5_1(.din(n13639), .dout(n13642));
    jdff dff_B_YydlJqw35_1(.din(n13642), .dout(n13645));
    jdff dff_B_bZESkjES9_1(.din(n13645), .dout(n13648));
    jdff dff_B_5Uifv4636_1(.din(n13648), .dout(n13651));
    jdff dff_B_nyAcTbUx9_1(.din(n13651), .dout(n13654));
    jdff dff_B_quG33DA47_1(.din(n13654), .dout(n13657));
    jdff dff_B_DagU8vkE8_1(.din(n13657), .dout(n13660));
    jdff dff_B_NdnLBpy36_1(.din(n13660), .dout(n13663));
    jdff dff_B_qzLi7wxI0_1(.din(n13663), .dout(n13666));
    jdff dff_B_vFSrm8xK7_1(.din(n13666), .dout(n13669));
    jdff dff_B_fSmRDmHs5_1(.din(n13669), .dout(n13672));
    jdff dff_B_qOHS1r4z9_1(.din(n1920), .dout(n13675));
    jdff dff_A_25J1ABlK1_0(.din(n13680), .dout(n13677));
    jdff dff_A_dN3XHPRR1_0(.din(n13683), .dout(n13680));
    jdff dff_A_xhb7EiLO9_0(.din(n13686), .dout(n13683));
    jdff dff_A_fiM37NNF6_0(.din(n13689), .dout(n13686));
    jdff dff_A_Vt79zmtK1_0(.din(n13692), .dout(n13689));
    jdff dff_A_X86iegjD5_0(.din(n13695), .dout(n13692));
    jdff dff_A_1GqdSVGj9_0(.din(n13698), .dout(n13695));
    jdff dff_A_vNkKSNx74_0(.din(n13701), .dout(n13698));
    jdff dff_A_At5yY3qr4_0(.din(n13704), .dout(n13701));
    jdff dff_A_GGZLjlkr5_0(.din(n13707), .dout(n13704));
    jdff dff_A_JQnaDncF0_0(.din(n13710), .dout(n13707));
    jdff dff_A_gHGlTTdY7_0(.din(n13713), .dout(n13710));
    jdff dff_A_jEfy5eT24_0(.din(n13716), .dout(n13713));
    jdff dff_A_6IQDB7TZ7_0(.din(n13719), .dout(n13716));
    jdff dff_A_E7tr3AmN3_0(.din(n13722), .dout(n13719));
    jdff dff_A_hleiiF2t2_0(.din(n13725), .dout(n13722));
    jdff dff_A_eqLjgLOn4_0(.din(n13728), .dout(n13725));
    jdff dff_A_91W6l9NE5_0(.din(n13731), .dout(n13728));
    jdff dff_A_9e2Mw5bp3_0(.din(n13734), .dout(n13731));
    jdff dff_A_Bulf4hA77_0(.din(n13737), .dout(n13734));
    jdff dff_A_7HAxMaP98_0(.din(n13740), .dout(n13737));
    jdff dff_A_53WWlr557_0(.din(n13743), .dout(n13740));
    jdff dff_A_VJ9VPnRZ1_0(.din(n13746), .dout(n13743));
    jdff dff_A_1mR2f2WZ5_0(.din(n13749), .dout(n13746));
    jdff dff_A_pAYbq8Wm4_0(.din(n13752), .dout(n13749));
    jdff dff_A_vpfnu7Zo2_0(.din(n13755), .dout(n13752));
    jdff dff_A_8QmlS4kl5_0(.din(n13758), .dout(n13755));
    jdff dff_A_YVshM2O80_0(.din(n13761), .dout(n13758));
    jdff dff_A_BbvnutCV7_0(.din(n13764), .dout(n13761));
    jdff dff_A_9bNkaOUZ7_0(.din(n13767), .dout(n13764));
    jdff dff_A_3Z9gBS8J2_0(.din(n13770), .dout(n13767));
    jdff dff_A_QyYqNGcL2_0(.din(n1609), .dout(n13770));
    jdff dff_A_y52OnWIm4_1(.din(n1898), .dout(n13773));
    jdff dff_B_03OhajKk6_1(.din(n1634), .dout(n13777));
    jdff dff_B_78yyYrFy9_1(.din(n13777), .dout(n13780));
    jdff dff_B_gP9qIGun5_1(.din(n13780), .dout(n13783));
    jdff dff_B_a0D0ATka5_1(.din(n13783), .dout(n13786));
    jdff dff_B_r5GjRDuH9_1(.din(n13786), .dout(n13789));
    jdff dff_B_uyfJ7Mt46_1(.din(n13789), .dout(n13792));
    jdff dff_B_vEwSBPt70_1(.din(n13792), .dout(n13795));
    jdff dff_B_shnxaGXY8_1(.din(n13795), .dout(n13798));
    jdff dff_B_sjrSdDmm3_1(.din(n13798), .dout(n13801));
    jdff dff_B_WpSDGyFr8_1(.din(n13801), .dout(n13804));
    jdff dff_B_YSayJaUO7_1(.din(n13804), .dout(n13807));
    jdff dff_B_L1y1wUmA7_1(.din(n13807), .dout(n13810));
    jdff dff_B_DhnnIlKP4_1(.din(n13810), .dout(n13813));
    jdff dff_B_aPPAH2Ah1_1(.din(n13813), .dout(n13816));
    jdff dff_B_CbCL1So65_1(.din(n13816), .dout(n13819));
    jdff dff_B_tF0PQgSd6_1(.din(n13819), .dout(n13822));
    jdff dff_B_W1EZMm6m4_1(.din(n13822), .dout(n13825));
    jdff dff_B_HBH1vVDM0_1(.din(n13825), .dout(n13828));
    jdff dff_B_GobGod4P7_1(.din(n13828), .dout(n13831));
    jdff dff_B_lg1clGu56_1(.din(n13831), .dout(n13834));
    jdff dff_B_VGX2ImSY9_1(.din(n13834), .dout(n13837));
    jdff dff_B_old76uYA3_1(.din(n13837), .dout(n13840));
    jdff dff_B_WLCDqwmH1_1(.din(n13840), .dout(n13843));
    jdff dff_B_OiiVPp338_1(.din(n13843), .dout(n13846));
    jdff dff_B_TzjhTPpi6_1(.din(n13846), .dout(n13849));
    jdff dff_B_SMsTbFdw7_1(.din(n13849), .dout(n13852));
    jdff dff_B_rrKbl2Oz7_1(.din(n13852), .dout(n13855));
    jdff dff_B_9nDqJSLu7_1(.din(n13855), .dout(n13858));
    jdff dff_B_DQfbDQM90_1(.din(n1619), .dout(n13861));
    jdff dff_A_koecHf197_0(.din(n13866), .dout(n13863));
    jdff dff_A_88of4Y3H2_0(.din(n13869), .dout(n13866));
    jdff dff_A_zUKI2ipk6_0(.din(n13872), .dout(n13869));
    jdff dff_A_Mg1QMq1y0_0(.din(n13875), .dout(n13872));
    jdff dff_A_KO8gUpMt8_0(.din(n13878), .dout(n13875));
    jdff dff_A_bZyjf5QM0_0(.din(n13881), .dout(n13878));
    jdff dff_A_Jp87AN728_0(.din(n13884), .dout(n13881));
    jdff dff_A_Vw0XLAzK7_0(.din(n13887), .dout(n13884));
    jdff dff_A_j1sNWFGB9_0(.din(n13890), .dout(n13887));
    jdff dff_A_nX2OLA8t1_0(.din(n13893), .dout(n13890));
    jdff dff_A_3bBkmYjL4_0(.din(n13896), .dout(n13893));
    jdff dff_A_GeiHwEMD0_0(.din(n13899), .dout(n13896));
    jdff dff_A_WZnIHl6l9_0(.din(n13902), .dout(n13899));
    jdff dff_A_p5kFz4gF7_0(.din(n13905), .dout(n13902));
    jdff dff_A_sx8ig0DO6_0(.din(n13908), .dout(n13905));
    jdff dff_A_mYZKCLuz6_0(.din(n13911), .dout(n13908));
    jdff dff_A_1oFOzSW69_0(.din(n13914), .dout(n13911));
    jdff dff_A_uGPvtTVX7_0(.din(n13917), .dout(n13914));
    jdff dff_A_zZu1xyvL2_0(.din(n13920), .dout(n13917));
    jdff dff_A_VybmS4eT2_0(.din(n13923), .dout(n13920));
    jdff dff_A_j5yhgpTH9_0(.din(n13926), .dout(n13923));
    jdff dff_A_VW0iDvQY7_0(.din(n13929), .dout(n13926));
    jdff dff_A_lVUI89H38_0(.din(n13932), .dout(n13929));
    jdff dff_A_vcBEXZuq6_0(.din(n13935), .dout(n13932));
    jdff dff_A_QF69uTUZ8_0(.din(n13938), .dout(n13935));
    jdff dff_A_iaD0Ui6t2_0(.din(n13941), .dout(n13938));
    jdff dff_A_E4NDaTF07_0(.din(n13944), .dout(n13941));
    jdff dff_A_3CQsH5Ge1_0(.din(n13947), .dout(n13944));
    jdff dff_A_Bh1ZRL9E6_0(.din(n1335), .dout(n13947));
    jdff dff_A_CjzJvrro2_1(.din(n1597), .dout(n13950));
    jdff dff_B_jPf9d1437_1(.din(n1360), .dout(n13954));
    jdff dff_B_PMZhOHfG5_1(.din(n13954), .dout(n13957));
    jdff dff_B_7m5Ljs6L5_1(.din(n13957), .dout(n13960));
    jdff dff_B_91Eq0bsZ1_1(.din(n13960), .dout(n13963));
    jdff dff_B_caNJuHBv3_1(.din(n13963), .dout(n13966));
    jdff dff_B_uq5XLDR71_1(.din(n13966), .dout(n13969));
    jdff dff_B_7sdbKtDC6_1(.din(n13969), .dout(n13972));
    jdff dff_B_Hhdpf7DE2_1(.din(n13972), .dout(n13975));
    jdff dff_B_6UqegZxt9_1(.din(n13975), .dout(n13978));
    jdff dff_B_sU8svXl31_1(.din(n13978), .dout(n13981));
    jdff dff_B_Stgp5cb35_1(.din(n13981), .dout(n13984));
    jdff dff_B_qngqHhWW7_1(.din(n13984), .dout(n13987));
    jdff dff_B_tZVYjBeh0_1(.din(n13987), .dout(n13990));
    jdff dff_B_Ar81sFvH3_1(.din(n13990), .dout(n13993));
    jdff dff_B_3P3blIMd6_1(.din(n13993), .dout(n13996));
    jdff dff_B_tGnemvza7_1(.din(n13996), .dout(n13999));
    jdff dff_B_TSPrvUGD6_1(.din(n13999), .dout(n14002));
    jdff dff_B_FdpkVCvy7_1(.din(n14002), .dout(n14005));
    jdff dff_B_cLibVtUJ7_1(.din(n14005), .dout(n14008));
    jdff dff_B_hra5wWkj4_1(.din(n14008), .dout(n14011));
    jdff dff_B_L4Z2YD5P5_1(.din(n14011), .dout(n14014));
    jdff dff_B_zBbDLL0r2_1(.din(n14014), .dout(n14017));
    jdff dff_B_V8cBGbxW4_1(.din(n14017), .dout(n14020));
    jdff dff_B_cUpVF8kC7_1(.din(n14020), .dout(n14023));
    jdff dff_B_wop3Ppbk9_1(.din(n14023), .dout(n14026));
    jdff dff_B_ZBjdgUM75_1(.din(n1345), .dout(n14029));
    jdff dff_A_4yTvoOGG4_0(.din(n14034), .dout(n14031));
    jdff dff_A_f4aJ6Dam8_0(.din(n14037), .dout(n14034));
    jdff dff_A_lH0gg2iX6_0(.din(n14040), .dout(n14037));
    jdff dff_A_zUAKggiq6_0(.din(n14043), .dout(n14040));
    jdff dff_A_vNUFrGXP7_0(.din(n14046), .dout(n14043));
    jdff dff_A_UfxBdeRD1_0(.din(n14049), .dout(n14046));
    jdff dff_A_VdQzMsFY8_0(.din(n14052), .dout(n14049));
    jdff dff_A_GhDlmh643_0(.din(n14055), .dout(n14052));
    jdff dff_A_6B1Ba9kp1_0(.din(n14058), .dout(n14055));
    jdff dff_A_Orz0hikz5_0(.din(n14061), .dout(n14058));
    jdff dff_A_t472kEWT1_0(.din(n14064), .dout(n14061));
    jdff dff_A_r2bAcMBp7_0(.din(n14067), .dout(n14064));
    jdff dff_A_kuDJKgVV6_0(.din(n14070), .dout(n14067));
    jdff dff_A_4EAKvhJF0_0(.din(n14073), .dout(n14070));
    jdff dff_A_ScwgxVOV1_0(.din(n14076), .dout(n14073));
    jdff dff_A_xDNSVloW3_0(.din(n14079), .dout(n14076));
    jdff dff_A_mJ4UpHWR6_0(.din(n14082), .dout(n14079));
    jdff dff_A_FQBlAXKf7_0(.din(n14085), .dout(n14082));
    jdff dff_A_2rVn07hh8_0(.din(n14088), .dout(n14085));
    jdff dff_A_xaaj5BxM3_0(.din(n14091), .dout(n14088));
    jdff dff_A_ApncF34F8_0(.din(n14094), .dout(n14091));
    jdff dff_A_HfF4ygvD2_0(.din(n14097), .dout(n14094));
    jdff dff_A_TwrHOL4N2_0(.din(n14100), .dout(n14097));
    jdff dff_A_WBeW4mnR4_0(.din(n14103), .dout(n14100));
    jdff dff_A_f5dVDaYY7_0(.din(n14106), .dout(n14103));
    jdff dff_A_t8tAzgMp1_0(.din(n1091), .dout(n14106));
    jdff dff_A_CHZGfPAc5_1(.din(n1323), .dout(n14109));
    jdff dff_B_uPooh4ko2_1(.din(n1116), .dout(n14113));
    jdff dff_B_jB9bx6RJ4_1(.din(n14113), .dout(n14116));
    jdff dff_B_rEj5h7iN0_1(.din(n14116), .dout(n14119));
    jdff dff_B_y2Bpli1n5_1(.din(n14119), .dout(n14122));
    jdff dff_B_z1Cb8xDh4_1(.din(n14122), .dout(n14125));
    jdff dff_B_fg0i13d87_1(.din(n14125), .dout(n14128));
    jdff dff_B_KXGIOptQ6_1(.din(n14128), .dout(n14131));
    jdff dff_B_jcuzs3am8_1(.din(n14131), .dout(n14134));
    jdff dff_B_mSXkN6kp4_1(.din(n14134), .dout(n14137));
    jdff dff_B_noNM6B8J1_1(.din(n14137), .dout(n14140));
    jdff dff_B_O0RoGiIr8_1(.din(n14140), .dout(n14143));
    jdff dff_B_VDCUgvIi3_1(.din(n14143), .dout(n14146));
    jdff dff_B_GnCt8pN18_1(.din(n14146), .dout(n14149));
    jdff dff_B_V9ew3Jy92_1(.din(n14149), .dout(n14152));
    jdff dff_B_i0ViKzR78_1(.din(n14152), .dout(n14155));
    jdff dff_B_6ylNFGro7_1(.din(n14155), .dout(n14158));
    jdff dff_B_ACRkX0KM3_1(.din(n14158), .dout(n14161));
    jdff dff_B_LZbVOwwh8_1(.din(n14161), .dout(n14164));
    jdff dff_B_IH4X7iGM9_1(.din(n14164), .dout(n14167));
    jdff dff_B_yu6bXgS87_1(.din(n14167), .dout(n14170));
    jdff dff_B_k6SXAJtP2_1(.din(n14170), .dout(n14173));
    jdff dff_B_v1w7e7PW8_1(.din(n14173), .dout(n14176));
    jdff dff_B_AjWbN0rr3_1(.din(n1101), .dout(n14179));
    jdff dff_A_6PiLb6KC4_0(.din(n14184), .dout(n14181));
    jdff dff_A_Bb9UfAdB0_0(.din(n14187), .dout(n14184));
    jdff dff_A_HPwUAGCC3_0(.din(n14190), .dout(n14187));
    jdff dff_A_dFCAAs831_0(.din(n14193), .dout(n14190));
    jdff dff_A_Iy9sInHu9_0(.din(n14196), .dout(n14193));
    jdff dff_A_VclKgW8m9_0(.din(n14199), .dout(n14196));
    jdff dff_A_qI9EW8fy2_0(.din(n14202), .dout(n14199));
    jdff dff_A_xyJySTWb1_0(.din(n14205), .dout(n14202));
    jdff dff_A_JSmQBqyU7_0(.din(n14208), .dout(n14205));
    jdff dff_A_TtAhHQGa5_0(.din(n14211), .dout(n14208));
    jdff dff_A_RSrEA1wc2_0(.din(n14214), .dout(n14211));
    jdff dff_A_2eu7Rc9D6_0(.din(n14217), .dout(n14214));
    jdff dff_A_ke2CuF9w4_0(.din(n14220), .dout(n14217));
    jdff dff_A_DmWln3eR4_0(.din(n14223), .dout(n14220));
    jdff dff_A_JLIO5ySW8_0(.din(n14226), .dout(n14223));
    jdff dff_A_QR3vwlDf0_0(.din(n14229), .dout(n14226));
    jdff dff_A_lYlufg023_0(.din(n14232), .dout(n14229));
    jdff dff_A_k4nutc9v4_0(.din(n14235), .dout(n14232));
    jdff dff_A_vpDUgNWM4_0(.din(n14238), .dout(n14235));
    jdff dff_A_xMXRsrhP8_0(.din(n14241), .dout(n14238));
    jdff dff_A_naWIhevA7_0(.din(n14244), .dout(n14241));
    jdff dff_A_V1cu7Egm0_0(.din(n14247), .dout(n14244));
    jdff dff_A_eUbJdN5F3_0(.din(n871), .dout(n14247));
    jdff dff_A_peHk2qng5_1(.din(n1079), .dout(n14250));
    jdff dff_B_3jm1LoUs7_1(.din(n896), .dout(n14254));
    jdff dff_B_5OHO6uYD6_1(.din(n14254), .dout(n14257));
    jdff dff_B_YdpCmWmt5_1(.din(n14257), .dout(n14260));
    jdff dff_B_d2BgRoeI9_1(.din(n14260), .dout(n14263));
    jdff dff_B_XfRatf0y3_1(.din(n14263), .dout(n14266));
    jdff dff_B_zgYCR2wc2_1(.din(n14266), .dout(n14269));
    jdff dff_B_3nhwhcBJ4_1(.din(n14269), .dout(n14272));
    jdff dff_B_6ETBEvVU5_1(.din(n14272), .dout(n14275));
    jdff dff_B_JKJeDhBx4_1(.din(n14275), .dout(n14278));
    jdff dff_B_z2UOf6LZ5_1(.din(n14278), .dout(n14281));
    jdff dff_B_3Tk7LKh01_1(.din(n14281), .dout(n14284));
    jdff dff_B_5MH3Oeh13_1(.din(n14284), .dout(n14287));
    jdff dff_B_t99yLnjP3_1(.din(n14287), .dout(n14290));
    jdff dff_B_ECHD0jid6_1(.din(n14290), .dout(n14293));
    jdff dff_B_lksvYya75_1(.din(n14293), .dout(n14296));
    jdff dff_B_jqsJEwL29_1(.din(n14296), .dout(n14299));
    jdff dff_B_g0eg8jXV5_1(.din(n14299), .dout(n14302));
    jdff dff_B_umj1hFfn6_1(.din(n14302), .dout(n14305));
    jdff dff_B_U0LQCSR08_1(.din(n14305), .dout(n14308));
    jdff dff_B_pRSP3AEO9_1(.din(n881), .dout(n14311));
    jdff dff_A_9DNkYF7O1_0(.din(n14316), .dout(n14313));
    jdff dff_A_MTW7eLSF3_0(.din(n14319), .dout(n14316));
    jdff dff_A_XOaFlA969_0(.din(n14322), .dout(n14319));
    jdff dff_A_vW6bK1cy4_0(.din(n14325), .dout(n14322));
    jdff dff_A_Db1PgHsM6_0(.din(n14328), .dout(n14325));
    jdff dff_A_wXTeGHmP5_0(.din(n14331), .dout(n14328));
    jdff dff_A_57S724kv0_0(.din(n14334), .dout(n14331));
    jdff dff_A_cHuF6PXi2_0(.din(n14337), .dout(n14334));
    jdff dff_A_lIFHSSwv1_0(.din(n14340), .dout(n14337));
    jdff dff_A_UW6i24ke9_0(.din(n14343), .dout(n14340));
    jdff dff_A_hz9fPhRz7_0(.din(n14346), .dout(n14343));
    jdff dff_A_7RfluJ9C7_0(.din(n14349), .dout(n14346));
    jdff dff_A_2CBO0o5u6_0(.din(n14352), .dout(n14349));
    jdff dff_A_wPxwHqT10_0(.din(n14355), .dout(n14352));
    jdff dff_A_TQfBR9oN4_0(.din(n14358), .dout(n14355));
    jdff dff_A_WyQ6RYTx7_0(.din(n14361), .dout(n14358));
    jdff dff_A_eCWI2sTG8_0(.din(n14364), .dout(n14361));
    jdff dff_A_S0RWZkCc7_0(.din(n14367), .dout(n14364));
    jdff dff_A_5eQzsYTy1_0(.din(n14370), .dout(n14367));
    jdff dff_A_edGf9AFJ6_0(.din(n678), .dout(n14370));
    jdff dff_A_tZxpkrLk3_1(.din(n859), .dout(n14373));
    jdff dff_B_h6JbXv9q1_1(.din(n703), .dout(n14377));
    jdff dff_B_5pF6I5F77_1(.din(n14377), .dout(n14380));
    jdff dff_B_vVA7RSmo9_1(.din(n14380), .dout(n14383));
    jdff dff_B_mARE0DzF5_1(.din(n14383), .dout(n14386));
    jdff dff_B_jZnpDUjS2_1(.din(n14386), .dout(n14389));
    jdff dff_B_MBIWsY8n5_1(.din(n14389), .dout(n14392));
    jdff dff_B_JebC4doU8_1(.din(n14392), .dout(n14395));
    jdff dff_B_0k6QPpgW6_1(.din(n14395), .dout(n14398));
    jdff dff_B_0K1i2wLI0_1(.din(n14398), .dout(n14401));
    jdff dff_B_8ETZk4Mc5_1(.din(n14401), .dout(n14404));
    jdff dff_B_DqYHRLOG4_1(.din(n14404), .dout(n14407));
    jdff dff_B_VOnfjZ3w1_1(.din(n14407), .dout(n14410));
    jdff dff_B_k9OxSITD3_1(.din(n14410), .dout(n14413));
    jdff dff_B_CjOzhyUA6_1(.din(n14413), .dout(n14416));
    jdff dff_B_wpjKZvYm1_1(.din(n14416), .dout(n14419));
    jdff dff_B_txgUulhx8_1(.din(n14419), .dout(n14422));
    jdff dff_B_rd8mdpko9_1(.din(n688), .dout(n14425));
    jdff dff_A_jFTrrHOP4_0(.din(n14430), .dout(n14427));
    jdff dff_A_HnMp1a7O1_0(.din(n14433), .dout(n14430));
    jdff dff_A_QOFFq5fX4_0(.din(n14436), .dout(n14433));
    jdff dff_A_YsTdaKn61_0(.din(n14439), .dout(n14436));
    jdff dff_A_55FDEM2a4_0(.din(n14442), .dout(n14439));
    jdff dff_A_0MrTwIOG1_0(.din(n14445), .dout(n14442));
    jdff dff_A_wLDUqIBe9_0(.din(n14448), .dout(n14445));
    jdff dff_A_GCZtswWN6_0(.din(n14451), .dout(n14448));
    jdff dff_A_0h0x7GFn7_0(.din(n14454), .dout(n14451));
    jdff dff_A_kXcckj9G0_0(.din(n14457), .dout(n14454));
    jdff dff_A_qLW1G1338_0(.din(n14460), .dout(n14457));
    jdff dff_A_a3wbc89U7_0(.din(n14463), .dout(n14460));
    jdff dff_A_UoZYWiHc9_0(.din(n14466), .dout(n14463));
    jdff dff_A_HDQ0hPqB8_0(.din(n14469), .dout(n14466));
    jdff dff_A_SJPEAaCf7_0(.din(n14472), .dout(n14469));
    jdff dff_A_OV18yayR5_0(.din(n14475), .dout(n14472));
    jdff dff_A_Ond58uNP5_0(.din(n515), .dout(n14475));
    jdff dff_A_iWmMC9ts3_1(.din(n666), .dout(n14478));
    jdff dff_B_bbmCodpv9_1(.din(n540), .dout(n14482));
    jdff dff_B_T3DLMfQa1_1(.din(n14482), .dout(n14485));
    jdff dff_B_ZGze8S695_1(.din(n14485), .dout(n14488));
    jdff dff_B_KelZoE8Z9_1(.din(n14488), .dout(n14491));
    jdff dff_B_WZqPo0yc3_1(.din(n14491), .dout(n14494));
    jdff dff_B_u1qfyp3f0_1(.din(n14494), .dout(n14497));
    jdff dff_B_VZCzrF6J2_1(.din(n14497), .dout(n14500));
    jdff dff_B_ld2M7Io84_1(.din(n14500), .dout(n14503));
    jdff dff_B_ej3hterM9_1(.din(n14503), .dout(n14506));
    jdff dff_B_BNA27gul1_1(.din(n14506), .dout(n14509));
    jdff dff_B_1dBIy7716_1(.din(n14509), .dout(n14512));
    jdff dff_B_9B6EDUzt7_1(.din(n14512), .dout(n14515));
    jdff dff_B_AmcbYULr1_1(.din(n14515), .dout(n14518));
    jdff dff_B_AwKqnTL31_1(.din(n525), .dout(n14521));
    jdff dff_A_DJjqOhdm7_0(.din(n14526), .dout(n14523));
    jdff dff_A_YvHKOKcx4_0(.din(n14529), .dout(n14526));
    jdff dff_A_eVvSIuyt5_0(.din(n14532), .dout(n14529));
    jdff dff_A_TroSCxah7_0(.din(n14535), .dout(n14532));
    jdff dff_A_9WzLxNoc4_0(.din(n14538), .dout(n14535));
    jdff dff_A_0DsPOaC91_0(.din(n14541), .dout(n14538));
    jdff dff_A_SUaqs6Qk8_0(.din(n14544), .dout(n14541));
    jdff dff_A_vedmNpOY1_0(.din(n14547), .dout(n14544));
    jdff dff_A_hzU4Gapk7_0(.din(n14550), .dout(n14547));
    jdff dff_A_DU3UOxV42_0(.din(n14553), .dout(n14550));
    jdff dff_A_9hV77ayo2_0(.din(n14556), .dout(n14553));
    jdff dff_A_T6AGU7rH3_0(.din(n14559), .dout(n14556));
    jdff dff_A_CCzX6Ho66_0(.din(n14562), .dout(n14559));
    jdff dff_A_0h3CobnG1_0(.din(n371), .dout(n14562));
    jdff dff_A_kqbN4kqC7_1(.din(n503), .dout(n14565));
    jdff dff_B_WDHxITla2_1(.din(n396), .dout(n14569));
    jdff dff_B_YHInVKxR8_1(.din(n14569), .dout(n14572));
    jdff dff_B_zeOKIsAd7_1(.din(n14572), .dout(n14575));
    jdff dff_B_fdAkYsbd6_1(.din(n14575), .dout(n14578));
    jdff dff_B_rndcK6l50_1(.din(n14578), .dout(n14581));
    jdff dff_B_5Mq1T8Oi4_1(.din(n14581), .dout(n14584));
    jdff dff_B_nBl7lXVE3_1(.din(n14584), .dout(n14587));
    jdff dff_B_EdRrC5GC0_1(.din(n14587), .dout(n14590));
    jdff dff_B_0vCdFfoY2_1(.din(n14590), .dout(n14593));
    jdff dff_B_Y7QU2Ebk7_1(.din(n14593), .dout(n14596));
    jdff dff_B_TKqaCuwG8_1(.din(n381), .dout(n14599));
    jdff dff_A_8kpIdcK42_0(.din(n14604), .dout(n14601));
    jdff dff_A_8D7AhApE5_0(.din(n14607), .dout(n14604));
    jdff dff_A_h55Xr0L76_0(.din(n14610), .dout(n14607));
    jdff dff_A_BcyEWGfB6_0(.din(n14613), .dout(n14610));
    jdff dff_A_uo5N9op78_0(.din(n14616), .dout(n14613));
    jdff dff_A_22USeGXd2_0(.din(n14619), .dout(n14616));
    jdff dff_A_HducLP3S1_0(.din(n14622), .dout(n14619));
    jdff dff_A_NOebkhnB5_0(.din(n14625), .dout(n14622));
    jdff dff_A_zww6rqlG3_0(.din(n14628), .dout(n14625));
    jdff dff_A_r6DPxvsI5_0(.din(n14631), .dout(n14628));
    jdff dff_A_Tooep5n49_0(.din(n239), .dout(n14631));
    jdff dff_A_VpV1Wt6x7_1(.din(n359), .dout(n14634));
    jdff dff_B_FxJTXI7R9_1(.din(n264), .dout(n14638));
    jdff dff_B_y8vDRHA60_1(.din(n14638), .dout(n14641));
    jdff dff_B_63Slu4xQ8_1(.din(n14641), .dout(n14644));
    jdff dff_B_Rf2K9rdr8_1(.din(n14644), .dout(n14647));
    jdff dff_B_42yb08Af2_1(.din(n14647), .dout(n14650));
    jdff dff_B_19nrQdrO5_1(.din(n14650), .dout(n14653));
    jdff dff_B_tBHNWRrm0_1(.din(n14653), .dout(n14656));
    jdff dff_B_1qvD8ff13_1(.din(n249), .dout(n14659));
    jdff dff_A_dTyP0f7L8_0(.din(n14664), .dout(n14661));
    jdff dff_A_bV00JtyD4_0(.din(n14667), .dout(n14664));
    jdff dff_A_U1trpJOS5_0(.din(n14670), .dout(n14667));
    jdff dff_A_ePo85IVu4_0(.din(n14673), .dout(n14670));
    jdff dff_A_ruNAtg1E0_0(.din(n14676), .dout(n14673));
    jdff dff_A_aYd37mFd2_0(.din(n14679), .dout(n14676));
    jdff dff_A_BE4QZEcY8_0(.din(n14682), .dout(n14679));
    jdff dff_A_JUvwpQwb8_0(.din(n160), .dout(n14682));
    jdff dff_A_YXMU8p9c8_1(.din(n227), .dout(n14685));
    jdff dff_B_6LZmB3Gn3_1(.din(n181), .dout(n14689));
    jdff dff_B_012J1un06_1(.din(n14689), .dout(n14692));
    jdff dff_B_OxwRlb8w7_1(.din(n14692), .dout(n14695));
    jdff dff_B_jffWmVSl8_1(.din(n14695), .dout(n14698));
    jdff dff_B_GUp30YFz8_1(.din(n166), .dout(n14701));
    jdff dff_B_CNllXBTv4_0(.din(n148), .dout(n14704));
    jdff dff_A_gix6zsfO9_0(.din(n14709), .dout(n14706));
    jdff dff_A_IN8XLFiq7_0(.din(n14712), .dout(n14709));
    jdff dff_A_OgaaY1J50_0(.din(n14715), .dout(n14712));
    jdff dff_A_FLj6H75i3_0(.din(n14718), .dout(n14715));
    jdff dff_A_MuhjVLNl5_0(.din(n98), .dout(n14718));
    jdff dff_A_nYOTDYLC5_0(.din(n90), .dout(n14721));
    jdff dff_A_uhOhIG0A7_0(.din(n87), .dout(n14724));
    jdff dff_A_HyISg1en7_1(.din(n4165), .dout(n14727));
    jdff dff_B_oFoXuBJi1_1(.din(n3782), .dout(n14731));
    jdff dff_B_uu5s7mxV8_2(.din(n3392), .dout(n14734));
    jdff dff_B_RrcJzKsF4_2(.din(n14734), .dout(n14737));
    jdff dff_B_RM9G0PvZ0_2(.din(n14737), .dout(n14740));
    jdff dff_B_s4PasYeV7_2(.din(n14740), .dout(n14743));
    jdff dff_B_vxw4WpAf9_2(.din(n14743), .dout(n14746));
    jdff dff_B_CIWvcv9n0_2(.din(n14746), .dout(n14749));
    jdff dff_B_zrqvvdgs2_2(.din(n14749), .dout(n14752));
    jdff dff_B_ibP34pDL5_2(.din(n14752), .dout(n14755));
    jdff dff_B_KvdxSQg76_2(.din(n14755), .dout(n14758));
    jdff dff_B_qS1V03CX0_2(.din(n14758), .dout(n14761));
    jdff dff_B_Z0CElkhq4_2(.din(n14761), .dout(n14764));
    jdff dff_B_Z4oX2eZC2_2(.din(n14764), .dout(n14767));
    jdff dff_B_mmnzgVYX2_2(.din(n14767), .dout(n14770));
    jdff dff_B_nIFa6QTK4_2(.din(n14770), .dout(n14773));
    jdff dff_B_jmxhQi6B0_2(.din(n14773), .dout(n14776));
    jdff dff_B_TCn8qOCJ0_2(.din(n14776), .dout(n14779));
    jdff dff_B_5LFSMMoA6_2(.din(n14779), .dout(n14782));
    jdff dff_B_VltZJW6A5_2(.din(n14782), .dout(n14785));
    jdff dff_B_N1Y9uENj0_2(.din(n14785), .dout(n14788));
    jdff dff_B_sYSfSS3X1_2(.din(n14788), .dout(n14791));
    jdff dff_B_GgAsFdPT7_2(.din(n14791), .dout(n14794));
    jdff dff_B_wFhOb4C65_2(.din(n14794), .dout(n14797));
    jdff dff_B_ESdU0vGh2_2(.din(n14797), .dout(n14800));
    jdff dff_B_3V9cVasK4_2(.din(n14800), .dout(n14803));
    jdff dff_B_0cHK6SdN2_2(.din(n14803), .dout(n14806));
    jdff dff_B_5mXlmx2L3_2(.din(n14806), .dout(n14809));
    jdff dff_B_wGCg2bAy6_2(.din(n14809), .dout(n14812));
    jdff dff_B_RVQJ6Jm35_2(.din(n14812), .dout(n14815));
    jdff dff_B_ja9cWSXL8_2(.din(n14815), .dout(n14818));
    jdff dff_B_Se2B2VG83_2(.din(n14818), .dout(n14821));
    jdff dff_B_IiGk1jLN6_2(.din(n14821), .dout(n14824));
    jdff dff_B_4VFrOGka8_2(.din(n14824), .dout(n14827));
    jdff dff_B_zSN1oP7s0_2(.din(n14827), .dout(n14830));
    jdff dff_B_SzOasAmJ6_2(.din(n14830), .dout(n14833));
    jdff dff_B_Sn72WNp93_2(.din(n14833), .dout(n14836));
    jdff dff_B_aUPtDaFI0_2(.din(n14836), .dout(n14839));
    jdff dff_B_DJwCsm9G0_2(.din(n14839), .dout(n14842));
    jdff dff_B_iBTf6qWn7_2(.din(n14842), .dout(n14845));
    jdff dff_B_LSnm5eJl7_2(.din(n14845), .dout(n14848));
    jdff dff_B_pBlO0dTg7_2(.din(n14848), .dout(n14851));
    jdff dff_B_mtHqs9xD2_2(.din(n14851), .dout(n14854));
    jdff dff_B_bvKCUuvs3_2(.din(n14854), .dout(n14857));
    jdff dff_B_QGnr771I8_2(.din(n14857), .dout(n14860));
    jdff dff_B_OUTFygTT9_2(.din(n14860), .dout(n14863));
    jdff dff_A_8FZFsssn1_0(.din(n3759), .dout(n14865));
    jdff dff_B_YU9Fs9yY9_1(.din(n3399), .dout(n14869));
    jdff dff_B_Cmju4XkZ6_2(.din(n2997), .dout(n14872));
    jdff dff_B_XKJLECiX2_2(.din(n14872), .dout(n14875));
    jdff dff_B_9iJPZpOG0_2(.din(n14875), .dout(n14878));
    jdff dff_B_riD7Hhbp0_2(.din(n14878), .dout(n14881));
    jdff dff_B_MUBFnhlV8_2(.din(n14881), .dout(n14884));
    jdff dff_B_oWvVhCi61_2(.din(n14884), .dout(n14887));
    jdff dff_B_244JvJfI4_2(.din(n14887), .dout(n14890));
    jdff dff_B_smPeRvbF6_2(.din(n14890), .dout(n14893));
    jdff dff_B_144CYuEf9_2(.din(n14893), .dout(n14896));
    jdff dff_B_VUKIUUqr1_2(.din(n14896), .dout(n14899));
    jdff dff_B_89P51siD4_2(.din(n14899), .dout(n14902));
    jdff dff_B_53acqq0B2_2(.din(n14902), .dout(n14905));
    jdff dff_B_QZyI493c2_2(.din(n14905), .dout(n14908));
    jdff dff_B_ieQuILvB7_2(.din(n14908), .dout(n14911));
    jdff dff_B_9XVzMyIm3_2(.din(n14911), .dout(n14914));
    jdff dff_B_CBSWQztz5_2(.din(n14914), .dout(n14917));
    jdff dff_B_rLPlqZ4P8_2(.din(n14917), .dout(n14920));
    jdff dff_B_V0N7pwgU0_2(.din(n14920), .dout(n14923));
    jdff dff_B_mJkgIjw38_2(.din(n14923), .dout(n14926));
    jdff dff_B_7JTOvEP82_2(.din(n14926), .dout(n14929));
    jdff dff_B_PexFvD751_2(.din(n14929), .dout(n14932));
    jdff dff_B_cONiCm715_2(.din(n14932), .dout(n14935));
    jdff dff_B_1rjeMho76_2(.din(n14935), .dout(n14938));
    jdff dff_B_53CgxPdn7_2(.din(n14938), .dout(n14941));
    jdff dff_B_HFO9JKgM9_2(.din(n14941), .dout(n14944));
    jdff dff_B_gNeO94Sq5_2(.din(n14944), .dout(n14947));
    jdff dff_B_8ZKoRUde3_2(.din(n14947), .dout(n14950));
    jdff dff_B_Kce3qLiA4_2(.din(n14950), .dout(n14953));
    jdff dff_B_N0iyvKSp3_2(.din(n14953), .dout(n14956));
    jdff dff_B_7hRlI4ES7_2(.din(n14956), .dout(n14959));
    jdff dff_B_KpSFj8zI0_2(.din(n14959), .dout(n14962));
    jdff dff_B_hFDt0Kgj7_2(.din(n14962), .dout(n14965));
    jdff dff_B_uIG9bSch6_2(.din(n14965), .dout(n14968));
    jdff dff_B_MO1mBpfc0_2(.din(n14968), .dout(n14971));
    jdff dff_B_PpjVTIOw8_2(.din(n14971), .dout(n14974));
    jdff dff_B_5MoCXwDb0_2(.din(n14974), .dout(n14977));
    jdff dff_B_wR1jJcqr2_2(.din(n14977), .dout(n14980));
    jdff dff_B_exRrguur1_2(.din(n14980), .dout(n14983));
    jdff dff_B_wcFWD4uh4_2(.din(n14983), .dout(n14986));
    jdff dff_B_RRR1lM4Q7_2(.din(n14986), .dout(n14989));
    jdff dff_B_N6d7RHoj3_2(.din(n14989), .dout(n14992));
    jdff dff_A_hHU6UceV1_1(.din(n3357), .dout(n14994));
    jdff dff_B_fzzOmr8J1_1(.din(n3020), .dout(n14998));
    jdff dff_B_yIf3oAeV5_1(.din(n14998), .dout(n15001));
    jdff dff_B_n1ODXD237_1(.din(n15001), .dout(n15004));
    jdff dff_B_wsJVEs0y7_1(.din(n15004), .dout(n15007));
    jdff dff_B_E0fa8WJR7_1(.din(n15007), .dout(n15010));
    jdff dff_B_4P9o2Dp96_1(.din(n15010), .dout(n15013));
    jdff dff_B_xnWLgX6V4_1(.din(n15013), .dout(n15016));
    jdff dff_B_UY0riLX37_1(.din(n15016), .dout(n15019));
    jdff dff_B_3BS2JmOQ3_1(.din(n15019), .dout(n15022));
    jdff dff_B_GSLimxgR9_1(.din(n15022), .dout(n15025));
    jdff dff_B_xlxmilYB6_1(.din(n15025), .dout(n15028));
    jdff dff_B_g0smN5WD2_1(.din(n15028), .dout(n15031));
    jdff dff_B_pZCtFNNp6_1(.din(n15031), .dout(n15034));
    jdff dff_B_YwwKu8VX9_1(.din(n15034), .dout(n15037));
    jdff dff_B_reuRlGSb4_1(.din(n15037), .dout(n15040));
    jdff dff_B_LDMW8fnj0_1(.din(n15040), .dout(n15043));
    jdff dff_B_ldAQpglH3_1(.din(n15043), .dout(n15046));
    jdff dff_B_U8ofqQwm2_1(.din(n15046), .dout(n15049));
    jdff dff_B_rsk4C2hf8_1(.din(n15049), .dout(n15052));
    jdff dff_B_0kIq5otZ5_1(.din(n15052), .dout(n15055));
    jdff dff_B_KghDC9zd6_1(.din(n15055), .dout(n15058));
    jdff dff_B_mcbKVaae7_1(.din(n15058), .dout(n15061));
    jdff dff_B_3jhVv5In6_1(.din(n15061), .dout(n15064));
    jdff dff_B_b8eEDtjU1_1(.din(n15064), .dout(n15067));
    jdff dff_B_iqDhQZyc2_1(.din(n15067), .dout(n15070));
    jdff dff_B_8xbn7ygX3_1(.din(n15070), .dout(n15073));
    jdff dff_B_SOSxbKXV8_1(.din(n15073), .dout(n15076));
    jdff dff_B_FGd2q3r20_1(.din(n15076), .dout(n15079));
    jdff dff_B_MAUVOqBM6_1(.din(n15079), .dout(n15082));
    jdff dff_B_hzdiH5tC3_1(.din(n15082), .dout(n15085));
    jdff dff_B_wQDkuLSQ2_1(.din(n15085), .dout(n15088));
    jdff dff_B_gnZ80UEL4_1(.din(n15088), .dout(n15091));
    jdff dff_B_6RSExyqG0_1(.din(n15091), .dout(n15094));
    jdff dff_B_TEwbDJuc7_1(.din(n15094), .dout(n15097));
    jdff dff_B_xxvzGOjw8_1(.din(n15097), .dout(n15100));
    jdff dff_B_k2Occ9hC0_1(.din(n15100), .dout(n15103));
    jdff dff_B_VV2MIwFT6_1(.din(n15103), .dout(n15106));
    jdff dff_B_KpqY4Roc0_1(.din(n3001), .dout(n15109));
    jdff dff_A_0x7sXd5j0_0(.din(n15114), .dout(n15111));
    jdff dff_A_1t0KfLDD4_0(.din(n15117), .dout(n15114));
    jdff dff_A_c1C5p1y66_0(.din(n15120), .dout(n15117));
    jdff dff_A_OEpCSvpc2_0(.din(n15123), .dout(n15120));
    jdff dff_A_HboQAD2X9_0(.din(n15126), .dout(n15123));
    jdff dff_A_VSaBkZhR9_0(.din(n15129), .dout(n15126));
    jdff dff_A_tx41zBWz7_0(.din(n15132), .dout(n15129));
    jdff dff_A_ar4OMavj3_0(.din(n15135), .dout(n15132));
    jdff dff_A_3kyOvU4F9_0(.din(n15138), .dout(n15135));
    jdff dff_A_QqCw3m452_0(.din(n15141), .dout(n15138));
    jdff dff_A_2TVhhPhf6_0(.din(n15144), .dout(n15141));
    jdff dff_A_eQ9CyBdA7_0(.din(n15147), .dout(n15144));
    jdff dff_A_Q6Bpm4h13_0(.din(n15150), .dout(n15147));
    jdff dff_A_zz8k9yHb4_0(.din(n15153), .dout(n15150));
    jdff dff_A_itMEMbUa8_0(.din(n15156), .dout(n15153));
    jdff dff_A_gP9gCfzn7_0(.din(n15159), .dout(n15156));
    jdff dff_A_EPexjiHt3_0(.din(n15162), .dout(n15159));
    jdff dff_A_gpcO4scG3_0(.din(n15165), .dout(n15162));
    jdff dff_A_hISEMg0b2_0(.din(n15168), .dout(n15165));
    jdff dff_A_AErJsgPT6_0(.din(n15171), .dout(n15168));
    jdff dff_A_XnsgTuen7_0(.din(n15174), .dout(n15171));
    jdff dff_A_gSUsSpUM9_0(.din(n15177), .dout(n15174));
    jdff dff_A_xJh2KpoY8_0(.din(n15180), .dout(n15177));
    jdff dff_A_aqHw9f9o2_0(.din(n15183), .dout(n15180));
    jdff dff_A_Z1OQV4rR3_0(.din(n15186), .dout(n15183));
    jdff dff_A_aW88qQaB0_0(.din(n15189), .dout(n15186));
    jdff dff_A_dBKO5jgt7_0(.din(n15192), .dout(n15189));
    jdff dff_A_tvTL01T53_0(.din(n15195), .dout(n15192));
    jdff dff_A_0NIWXbRw4_0(.din(n15198), .dout(n15195));
    jdff dff_A_RF6jJ1qM4_0(.din(n15201), .dout(n15198));
    jdff dff_A_wpKf0Pax1_0(.din(n15204), .dout(n15201));
    jdff dff_A_cSGwaseN9_0(.din(n15207), .dout(n15204));
    jdff dff_A_IqWGRieV0_0(.din(n15210), .dout(n15207));
    jdff dff_A_MquVKvAs7_0(.din(n15213), .dout(n15210));
    jdff dff_A_iK6EvYbl7_0(.din(n15216), .dout(n15213));
    jdff dff_A_ojtGVxro0_0(.din(n15219), .dout(n15216));
    jdff dff_A_VdfbowkM1_0(.din(n15222), .dout(n15219));
    jdff dff_A_7YxzHdl95_0(.din(n2615), .dout(n15222));
    jdff dff_A_CZ2jEFdf6_0(.din(n2952), .dout(n15225));
    jdff dff_B_n1qofQ7N6_1(.din(n2622), .dout(n15229));
    jdff dff_A_To4CQYwR5_0(.din(n15234), .dout(n15231));
    jdff dff_A_ggh7op5Z7_0(.din(n15237), .dout(n15234));
    jdff dff_A_yxOIQ4lR2_0(.din(n15240), .dout(n15237));
    jdff dff_A_FrkpCw5a8_0(.din(n15243), .dout(n15240));
    jdff dff_A_JElZmtGa1_0(.din(n15246), .dout(n15243));
    jdff dff_A_3mFIzyLZ1_0(.din(n15249), .dout(n15246));
    jdff dff_A_3HmzR6yy1_0(.din(n15252), .dout(n15249));
    jdff dff_A_RlOVBzJF3_0(.din(n15255), .dout(n15252));
    jdff dff_A_eCWTqBit2_0(.din(n15258), .dout(n15255));
    jdff dff_A_smlIJURR8_0(.din(n15261), .dout(n15258));
    jdff dff_A_Aeraraba3_0(.din(n15264), .dout(n15261));
    jdff dff_A_WbXmNPCy1_0(.din(n15267), .dout(n15264));
    jdff dff_A_fzBGNR4C0_0(.din(n15270), .dout(n15267));
    jdff dff_A_pDscmNUD6_0(.din(n15273), .dout(n15270));
    jdff dff_A_1rabCNHB7_0(.din(n15276), .dout(n15273));
    jdff dff_A_tEb8e0M24_0(.din(n15279), .dout(n15276));
    jdff dff_A_EWJSBKE89_0(.din(n15282), .dout(n15279));
    jdff dff_A_GMdCjHzv1_0(.din(n15285), .dout(n15282));
    jdff dff_A_8DzFQCZx0_0(.din(n15288), .dout(n15285));
    jdff dff_A_5gg0W96i4_0(.din(n15291), .dout(n15288));
    jdff dff_A_mF2BH9hX5_0(.din(n15294), .dout(n15291));
    jdff dff_A_6qLITpxo1_0(.din(n15297), .dout(n15294));
    jdff dff_A_gvQuIHqD6_0(.din(n15300), .dout(n15297));
    jdff dff_A_np2AACK71_0(.din(n15303), .dout(n15300));
    jdff dff_A_dSSqv5el9_0(.din(n15306), .dout(n15303));
    jdff dff_A_6ZcnzBpi8_0(.din(n15309), .dout(n15306));
    jdff dff_A_9TJo8J1h8_0(.din(n15312), .dout(n15309));
    jdff dff_A_A3svwYQ96_0(.din(n15315), .dout(n15312));
    jdff dff_A_wgUbjRhB2_0(.din(n15318), .dout(n15315));
    jdff dff_A_7HSPdK1j0_0(.din(n15321), .dout(n15318));
    jdff dff_A_htXIfznG4_0(.din(n15324), .dout(n15321));
    jdff dff_A_WKGGiWb44_0(.din(n15327), .dout(n15324));
    jdff dff_A_XareqLXt0_0(.din(n15330), .dout(n15327));
    jdff dff_A_gM7V1X5D8_0(.din(n15333), .dout(n15330));
    jdff dff_A_1KDVfjr33_0(.din(n2260), .dout(n15333));
    jdff dff_A_OgeeSzwv6_0(.din(n2570), .dout(n15336));
    jdff dff_B_T0JlXUcf3_1(.din(n2267), .dout(n15340));
    jdff dff_A_1FBtlnJd4_0(.din(n15345), .dout(n15342));
    jdff dff_A_YRhvihQA6_0(.din(n15348), .dout(n15345));
    jdff dff_A_2u9NoB241_0(.din(n15351), .dout(n15348));
    jdff dff_A_qw0GAhjs9_0(.din(n15354), .dout(n15351));
    jdff dff_A_QDn77CaY5_0(.din(n15357), .dout(n15354));
    jdff dff_A_voPjoagP0_0(.din(n15360), .dout(n15357));
    jdff dff_A_FJAaoLIb1_0(.din(n15363), .dout(n15360));
    jdff dff_A_GLoNUQPe4_0(.din(n15366), .dout(n15363));
    jdff dff_A_hvLyiykL5_0(.din(n15369), .dout(n15366));
    jdff dff_A_6E27U3Vr7_0(.din(n15372), .dout(n15369));
    jdff dff_A_kZyClB2W3_0(.din(n15375), .dout(n15372));
    jdff dff_A_szql5YIY2_0(.din(n15378), .dout(n15375));
    jdff dff_A_dhUrHtm81_0(.din(n15381), .dout(n15378));
    jdff dff_A_uVzSUWcq3_0(.din(n15384), .dout(n15381));
    jdff dff_A_6OhY4Zcq0_0(.din(n15387), .dout(n15384));
    jdff dff_A_jlwv0Zhf6_0(.din(n15390), .dout(n15387));
    jdff dff_A_9AwAA0PN1_0(.din(n15393), .dout(n15390));
    jdff dff_A_jMPHnMES8_0(.din(n15396), .dout(n15393));
    jdff dff_A_STtMjR668_0(.din(n15399), .dout(n15396));
    jdff dff_A_i4fnA0FW5_0(.din(n15402), .dout(n15399));
    jdff dff_A_9ca1J4kT0_0(.din(n15405), .dout(n15402));
    jdff dff_A_4KZVR7Fb3_0(.din(n15408), .dout(n15405));
    jdff dff_A_OY8XUwl90_0(.din(n15411), .dout(n15408));
    jdff dff_A_qWRvH4Bx0_0(.din(n15414), .dout(n15411));
    jdff dff_A_Vp8wa24D0_0(.din(n15417), .dout(n15414));
    jdff dff_A_wVfnTa6n8_0(.din(n15420), .dout(n15417));
    jdff dff_A_ZVuLWI3g9_0(.din(n15423), .dout(n15420));
    jdff dff_A_ctXthAzv4_0(.din(n15426), .dout(n15423));
    jdff dff_A_iQzNwUYQ3_0(.din(n15429), .dout(n15426));
    jdff dff_A_pB3OO0pO7_0(.din(n15432), .dout(n15429));
    jdff dff_A_w2rvrd2E6_0(.din(n15435), .dout(n15432));
    jdff dff_A_4Sqb3nNa1_0(.din(n1932), .dout(n15435));
    jdff dff_A_5WYeOW9D8_0(.din(n2215), .dout(n15438));
    jdff dff_B_SpoUZEwd0_1(.din(n1939), .dout(n15442));
    jdff dff_A_BonLGtCS7_0(.din(n15447), .dout(n15444));
    jdff dff_A_qXCCAQEi7_0(.din(n15450), .dout(n15447));
    jdff dff_A_hvhrF0bn2_0(.din(n15453), .dout(n15450));
    jdff dff_A_hZ6uZVYi5_0(.din(n15456), .dout(n15453));
    jdff dff_A_FpERn6Cd7_0(.din(n15459), .dout(n15456));
    jdff dff_A_KEBm57gp9_0(.din(n15462), .dout(n15459));
    jdff dff_A_Ff4uTXqb2_0(.din(n15465), .dout(n15462));
    jdff dff_A_4KQt9KZB9_0(.din(n15468), .dout(n15465));
    jdff dff_A_aSzd3V5y7_0(.din(n15471), .dout(n15468));
    jdff dff_A_eQBooRoZ2_0(.din(n15474), .dout(n15471));
    jdff dff_A_9EjCucF43_0(.din(n15477), .dout(n15474));
    jdff dff_A_rnB0gZ014_0(.din(n15480), .dout(n15477));
    jdff dff_A_D8avDmqJ8_0(.din(n15483), .dout(n15480));
    jdff dff_A_zjAVnxuZ6_0(.din(n15486), .dout(n15483));
    jdff dff_A_QgM4FMme2_0(.din(n15489), .dout(n15486));
    jdff dff_A_6jVIJBg65_0(.din(n15492), .dout(n15489));
    jdff dff_A_iSLGsF3h3_0(.din(n15495), .dout(n15492));
    jdff dff_A_FHou2Rh10_0(.din(n15498), .dout(n15495));
    jdff dff_A_GQCklcge3_0(.din(n15501), .dout(n15498));
    jdff dff_A_oSYctBLT9_0(.din(n15504), .dout(n15501));
    jdff dff_A_jFsyfJ843_0(.din(n15507), .dout(n15504));
    jdff dff_A_eAmjjxs99_0(.din(n15510), .dout(n15507));
    jdff dff_A_Oa5q03m06_0(.din(n15513), .dout(n15510));
    jdff dff_A_slspMlqY1_0(.din(n15516), .dout(n15513));
    jdff dff_A_cSBYrpul6_0(.din(n15519), .dout(n15516));
    jdff dff_A_lzmXifd79_0(.din(n15522), .dout(n15519));
    jdff dff_A_InnUBaSo2_0(.din(n15525), .dout(n15522));
    jdff dff_A_E2J9lZA42_0(.din(n15528), .dout(n15525));
    jdff dff_A_UZ7DrGWN9_0(.din(n1631), .dout(n15528));
    jdff dff_A_8tiOknIL2_0(.din(n1887), .dout(n15531));
    jdff dff_B_wkFc1ith2_1(.din(n1638), .dout(n15535));
    jdff dff_A_Z0qkaj588_0(.din(n15540), .dout(n15537));
    jdff dff_A_Mgna3mO74_0(.din(n15543), .dout(n15540));
    jdff dff_A_0K0H1mcN6_0(.din(n15546), .dout(n15543));
    jdff dff_A_U8uKCunH7_0(.din(n15549), .dout(n15546));
    jdff dff_A_ZCcxNhSW5_0(.din(n15552), .dout(n15549));
    jdff dff_A_Vq4Igk4k9_0(.din(n15555), .dout(n15552));
    jdff dff_A_leSBSrue9_0(.din(n15558), .dout(n15555));
    jdff dff_A_a1D3WmsL1_0(.din(n15561), .dout(n15558));
    jdff dff_A_97FYEoeL1_0(.din(n15564), .dout(n15561));
    jdff dff_A_NeaUB9Zu6_0(.din(n15567), .dout(n15564));
    jdff dff_A_wLEdSDoS0_0(.din(n15570), .dout(n15567));
    jdff dff_A_AZ733hQx0_0(.din(n15573), .dout(n15570));
    jdff dff_A_owYA2bLA9_0(.din(n15576), .dout(n15573));
    jdff dff_A_h1BVIcgu9_0(.din(n15579), .dout(n15576));
    jdff dff_A_OKGD1lo05_0(.din(n15582), .dout(n15579));
    jdff dff_A_L2wyClKZ6_0(.din(n15585), .dout(n15582));
    jdff dff_A_1pTA4NV72_0(.din(n15588), .dout(n15585));
    jdff dff_A_sulAL0da8_0(.din(n15591), .dout(n15588));
    jdff dff_A_jKqVXPEE7_0(.din(n15594), .dout(n15591));
    jdff dff_A_5ZzBjgKr7_0(.din(n15597), .dout(n15594));
    jdff dff_A_fh5MXxQN3_0(.din(n15600), .dout(n15597));
    jdff dff_A_kCwfeBfB8_0(.din(n15603), .dout(n15600));
    jdff dff_A_Se7yCc9P7_0(.din(n15606), .dout(n15603));
    jdff dff_A_alDo3FBj1_0(.din(n15609), .dout(n15606));
    jdff dff_A_jw9LVS7v8_0(.din(n15612), .dout(n15609));
    jdff dff_A_pPk0ZHij9_0(.din(n1357), .dout(n15612));
    jdff dff_A_w7T9nth90_0(.din(n1586), .dout(n15615));
    jdff dff_B_cNZdpEw14_1(.din(n1364), .dout(n15619));
    jdff dff_A_dDbcnEjY4_0(.din(n15624), .dout(n15621));
    jdff dff_A_JIpFM2TJ9_0(.din(n15627), .dout(n15624));
    jdff dff_A_UivY7Xvx2_0(.din(n15630), .dout(n15627));
    jdff dff_A_66jSKIFW0_0(.din(n15633), .dout(n15630));
    jdff dff_A_c7SNGAbI1_0(.din(n15636), .dout(n15633));
    jdff dff_A_Qn1WG3OA6_0(.din(n15639), .dout(n15636));
    jdff dff_A_UX79hV7d6_0(.din(n15642), .dout(n15639));
    jdff dff_A_3QMeQRYx4_0(.din(n15645), .dout(n15642));
    jdff dff_A_AkiNZV2m3_0(.din(n15648), .dout(n15645));
    jdff dff_A_4GLBo9I30_0(.din(n15651), .dout(n15648));
    jdff dff_A_C6znERXG9_0(.din(n15654), .dout(n15651));
    jdff dff_A_OTrDjAso9_0(.din(n15657), .dout(n15654));
    jdff dff_A_M9TN7u1o8_0(.din(n15660), .dout(n15657));
    jdff dff_A_SpNUAerN7_0(.din(n15663), .dout(n15660));
    jdff dff_A_Li1BxMt35_0(.din(n15666), .dout(n15663));
    jdff dff_A_hVARLdF90_0(.din(n15669), .dout(n15666));
    jdff dff_A_KOyFnJ6P3_0(.din(n15672), .dout(n15669));
    jdff dff_A_heyaKFTt6_0(.din(n15675), .dout(n15672));
    jdff dff_A_IfoL8a475_0(.din(n15678), .dout(n15675));
    jdff dff_A_qzKxelDI9_0(.din(n15681), .dout(n15678));
    jdff dff_A_wrjPjiGi8_0(.din(n15684), .dout(n15681));
    jdff dff_A_U06rrlK61_0(.din(n15687), .dout(n15684));
    jdff dff_A_F7GGot049_0(.din(n1113), .dout(n15687));
    jdff dff_A_H5a6kMnc7_0(.din(n1312), .dout(n15690));
    jdff dff_B_YN9xniCe7_1(.din(n1120), .dout(n15694));
    jdff dff_A_B3WQpwTl4_0(.din(n15699), .dout(n15696));
    jdff dff_A_0YemFUP72_0(.din(n15702), .dout(n15699));
    jdff dff_A_KRiL7IEK0_0(.din(n15705), .dout(n15702));
    jdff dff_A_GBy94EUE8_0(.din(n15708), .dout(n15705));
    jdff dff_A_zaQIbnIG7_0(.din(n15711), .dout(n15708));
    jdff dff_A_TRKK8lrZ0_0(.din(n15714), .dout(n15711));
    jdff dff_A_fHLYcBzl5_0(.din(n15717), .dout(n15714));
    jdff dff_A_jeGCbEct3_0(.din(n15720), .dout(n15717));
    jdff dff_A_xwjJ8Hl73_0(.din(n15723), .dout(n15720));
    jdff dff_A_l0S9gEMM7_0(.din(n15726), .dout(n15723));
    jdff dff_A_4eGXOV3D3_0(.din(n15729), .dout(n15726));
    jdff dff_A_A5zXeENM3_0(.din(n15732), .dout(n15729));
    jdff dff_A_pH1V3gBq1_0(.din(n15735), .dout(n15732));
    jdff dff_A_O5YybVCM4_0(.din(n15738), .dout(n15735));
    jdff dff_A_AYkCkQii3_0(.din(n15741), .dout(n15738));
    jdff dff_A_E8GAXqDH7_0(.din(n15744), .dout(n15741));
    jdff dff_A_6XWz6aFm8_0(.din(n15747), .dout(n15744));
    jdff dff_A_cC0z3G040_0(.din(n15750), .dout(n15747));
    jdff dff_A_5pWPVmoE9_0(.din(n15753), .dout(n15750));
    jdff dff_A_bWWMFQmV5_0(.din(n893), .dout(n15753));
    jdff dff_A_vOuZa3lL8_0(.din(n1068), .dout(n15756));
    jdff dff_B_t7zGmDAA3_1(.din(n900), .dout(n15760));
    jdff dff_A_2UkcZ4Vf5_0(.din(n15765), .dout(n15762));
    jdff dff_A_3tkynaLc6_0(.din(n15768), .dout(n15765));
    jdff dff_A_Bn60p0gt6_0(.din(n15771), .dout(n15768));
    jdff dff_A_LBSeKYrW7_0(.din(n15774), .dout(n15771));
    jdff dff_A_ktP54q1O9_0(.din(n15777), .dout(n15774));
    jdff dff_A_oKlHnjZ98_0(.din(n15780), .dout(n15777));
    jdff dff_A_5fnwKwEV0_0(.din(n15783), .dout(n15780));
    jdff dff_A_28cwp9BN3_0(.din(n15786), .dout(n15783));
    jdff dff_A_TZyYsELy1_0(.din(n15789), .dout(n15786));
    jdff dff_A_PdIZnOZs0_0(.din(n15792), .dout(n15789));
    jdff dff_A_qu5JsAQ68_0(.din(n15795), .dout(n15792));
    jdff dff_A_iIdUagJN7_0(.din(n15798), .dout(n15795));
    jdff dff_A_7DmEP9vG1_0(.din(n15801), .dout(n15798));
    jdff dff_A_QHMsashP2_0(.din(n15804), .dout(n15801));
    jdff dff_A_Z335YrJW3_0(.din(n15807), .dout(n15804));
    jdff dff_A_YzF7m0cY7_0(.din(n15810), .dout(n15807));
    jdff dff_A_Q4WRj3c35_0(.din(n700), .dout(n15810));
    jdff dff_A_AoFzQpzy8_0(.din(n848), .dout(n15813));
    jdff dff_B_0Uuq0fZ45_1(.din(n707), .dout(n15817));
    jdff dff_A_2QI3qJVS2_0(.din(n15822), .dout(n15819));
    jdff dff_A_4TwJTyUU2_0(.din(n15825), .dout(n15822));
    jdff dff_A_zxDsxLGi9_0(.din(n15828), .dout(n15825));
    jdff dff_A_lCKEQrTs5_0(.din(n15831), .dout(n15828));
    jdff dff_A_D7FM4cfR4_0(.din(n15834), .dout(n15831));
    jdff dff_A_bh17kYxA5_0(.din(n15837), .dout(n15834));
    jdff dff_A_Y0CCq4A94_0(.din(n15840), .dout(n15837));
    jdff dff_A_NK5EfVlx2_0(.din(n15843), .dout(n15840));
    jdff dff_A_dLqodMmE1_0(.din(n15846), .dout(n15843));
    jdff dff_A_sagg0vuS4_0(.din(n15849), .dout(n15846));
    jdff dff_A_0LFcPuXD3_0(.din(n15852), .dout(n15849));
    jdff dff_A_cKBBEiH61_0(.din(n15855), .dout(n15852));
    jdff dff_A_NB7t1PsP8_0(.din(n15858), .dout(n15855));
    jdff dff_A_E3uuICfZ1_0(.din(n537), .dout(n15858));
    jdff dff_A_AGyhUYPC7_0(.din(n655), .dout(n15861));
    jdff dff_B_5lD7qqqs3_1(.din(n544), .dout(n15865));
    jdff dff_A_AeuZPtDG8_0(.din(n15870), .dout(n15867));
    jdff dff_A_vrALIgrq6_0(.din(n15873), .dout(n15870));
    jdff dff_A_qH8KSHAO7_0(.din(n15876), .dout(n15873));
    jdff dff_A_ilmxlb7E5_0(.din(n15879), .dout(n15876));
    jdff dff_A_ke8BPedF2_0(.din(n15882), .dout(n15879));
    jdff dff_A_inHWBLTv5_0(.din(n15885), .dout(n15882));
    jdff dff_A_pccu4gh62_0(.din(n15888), .dout(n15885));
    jdff dff_A_IbKovbYn7_0(.din(n15891), .dout(n15888));
    jdff dff_A_fu6aqHvG5_0(.din(n15894), .dout(n15891));
    jdff dff_A_0EY2T5k61_0(.din(n15897), .dout(n15894));
    jdff dff_A_VWcmwtMh6_0(.din(n393), .dout(n15897));
    jdff dff_A_m59HVWWN7_0(.din(n492), .dout(n15900));
    jdff dff_B_Mhfr6fth5_1(.din(n400), .dout(n15904));
    jdff dff_A_hyLvjgaq0_0(.din(n15909), .dout(n15906));
    jdff dff_A_fBk1XXtD8_0(.din(n15912), .dout(n15909));
    jdff dff_A_zOV19tar9_0(.din(n15915), .dout(n15912));
    jdff dff_A_cxfpP6D50_0(.din(n15918), .dout(n15915));
    jdff dff_A_e9mREQgc5_0(.din(n15921), .dout(n15918));
    jdff dff_A_dDUC5QbX1_0(.din(n15924), .dout(n15921));
    jdff dff_A_HeV4VCqy0_0(.din(n15927), .dout(n15924));
    jdff dff_A_lF7GCaFH7_0(.din(n261), .dout(n15927));
    jdff dff_A_SZD2cvwN7_0(.din(n348), .dout(n15930));
    jdff dff_A_ykQi1sID8_0(.din(n216), .dout(n15933));
    jdff dff_A_bcA037ij8_0(.din(n144), .dout(n15936));
    jdff dff_A_3cslWXqh6_1(.din(n133), .dout(n15939));
    jdff dff_A_FWT5Eskw0_0(.din(n15945), .dout(n15942));
    jdff dff_A_100ztZiO3_0(.din(n15948), .dout(n15945));
    jdff dff_A_rKcGLXn78_0(.din(n15951), .dout(n15948));
    jdff dff_A_zmkCMecj4_0(.din(n15954), .dout(n15951));
    jdff dff_A_K0SsOrCV3_0(.din(n178), .dout(n15954));
    jdff dff_A_dpwNAxEi6_0(.din(n15960), .dout(n15957));
    jdff dff_A_QvvnFDEe2_0(.din(n212), .dout(n15960));
    jdff dff_B_GTzGY71r8_1(.din(n189), .dout(n15964));
    jdff dff_A_JJnjh7cr5_1(.din(n133), .dout(n15966));
    jdff dff_A_O3sEcoDA0_2(.din(n15972), .dout(n15969));
    jdff dff_A_129vUXF14_2(.din(n133), .dout(n15972));
    jdff dff_A_58oNjSm74_0(.din(n15979), .dout(n15975));
    jdff dff_B_Xfkd7YaU7_2(.din(n4206), .dout(n15979));
    jdff dff_B_XYCnbEGk1_2(.din(n3798), .dout(n15982));
    jdff dff_B_ALEJVILM3_2(.din(n15982), .dout(n15985));
    jdff dff_B_hfXJN78t0_2(.din(n15985), .dout(n15988));
    jdff dff_B_IzVQw3Tg1_2(.din(n15988), .dout(n15991));
    jdff dff_B_86eJopzj1_2(.din(n15991), .dout(n15994));
    jdff dff_B_z0CKpGcV5_2(.din(n15994), .dout(n15997));
    jdff dff_B_VQGFMzn25_2(.din(n15997), .dout(n16000));
    jdff dff_B_pMLI55rQ1_2(.din(n16000), .dout(n16003));
    jdff dff_B_W07sIFpL5_2(.din(n16003), .dout(n16006));
    jdff dff_B_b4GITiFx9_2(.din(n16006), .dout(n16009));
    jdff dff_B_7vqDzFke6_2(.din(n16009), .dout(n16012));
    jdff dff_B_AFOV77Yp9_2(.din(n16012), .dout(n16015));
    jdff dff_B_LLMZEDco8_2(.din(n16015), .dout(n16018));
    jdff dff_B_IHcIAwtU1_2(.din(n16018), .dout(n16021));
    jdff dff_B_SX5AH0VY9_2(.din(n16021), .dout(n16024));
    jdff dff_B_skJe9Cz49_2(.din(n16024), .dout(n16027));
    jdff dff_B_GJkn4qjp1_2(.din(n16027), .dout(n16030));
    jdff dff_B_klc7ieDe0_2(.din(n16030), .dout(n16033));
    jdff dff_B_wwrrlaah7_2(.din(n16033), .dout(n16036));
    jdff dff_B_8JFqXxNQ4_2(.din(n16036), .dout(n16039));
    jdff dff_B_GXl8i9xh2_2(.din(n16039), .dout(n16042));
    jdff dff_B_1XnU7mGy5_2(.din(n16042), .dout(n16045));
    jdff dff_B_7yYzIjPa6_2(.din(n16045), .dout(n16048));
    jdff dff_B_E2v58dEj9_2(.din(n16048), .dout(n16051));
    jdff dff_B_GGvRfait7_2(.din(n16051), .dout(n16054));
    jdff dff_B_8421x3Dt3_2(.din(n16054), .dout(n16057));
    jdff dff_B_rIQAlWVs4_2(.din(n16057), .dout(n16060));
    jdff dff_B_FV3ApBIe9_2(.din(n16060), .dout(n16063));
    jdff dff_B_9QeiNDJJ8_2(.din(n16063), .dout(n16066));
    jdff dff_B_3Jm3eYIe2_2(.din(n16066), .dout(n16069));
    jdff dff_B_JaCMRJUa7_2(.din(n16069), .dout(n16072));
    jdff dff_B_7gh0oi4N6_2(.din(n16072), .dout(n16075));
    jdff dff_B_YrVzFK9A7_2(.din(n16075), .dout(n16078));
    jdff dff_B_LseRDJ8k7_2(.din(n16078), .dout(n16081));
    jdff dff_B_aYL9nx0e2_2(.din(n16081), .dout(n16084));
    jdff dff_B_77BJru3w1_2(.din(n16084), .dout(n16087));
    jdff dff_B_210xLPz89_2(.din(n16087), .dout(n16090));
    jdff dff_B_ai8Za3sR0_2(.din(n16090), .dout(n16093));
    jdff dff_B_7stG2Ylw7_2(.din(n16093), .dout(n16096));
    jdff dff_B_rD4XypI92_2(.din(n16096), .dout(n16099));
    jdff dff_B_9k8wHymZ8_2(.din(n16099), .dout(n16102));
    jdff dff_B_si7ZQzf03_2(.din(n16102), .dout(n16105));
    jdff dff_B_4MuhyZz56_2(.din(n16105), .dout(n16108));
    jdff dff_B_A3hoYYku9_2(.din(n16108), .dout(n16111));
    jdff dff_A_0WP8bNhx8_0(.din(n3813), .dout(n16113));
    jdff dff_B_ixj7yUiC0_1(.din(n3805), .dout(n16117));
    jdff dff_B_RdEFjcEE0_2(.din(n3411), .dout(n16120));
    jdff dff_B_MV4bqQJz9_2(.din(n16120), .dout(n16123));
    jdff dff_B_ClRaOHsw9_2(.din(n16123), .dout(n16126));
    jdff dff_B_UHV0fyxY3_2(.din(n16126), .dout(n16129));
    jdff dff_B_dygcDZ8r6_2(.din(n16129), .dout(n16132));
    jdff dff_B_6TgLpY779_2(.din(n16132), .dout(n16135));
    jdff dff_B_ir36mJq39_2(.din(n16135), .dout(n16138));
    jdff dff_B_8JZxrxqd7_2(.din(n16138), .dout(n16141));
    jdff dff_B_qmho1tvv5_2(.din(n16141), .dout(n16144));
    jdff dff_B_eA36qhs15_2(.din(n16144), .dout(n16147));
    jdff dff_B_vKHAUT8B3_2(.din(n16147), .dout(n16150));
    jdff dff_B_NHDgziGL8_2(.din(n16150), .dout(n16153));
    jdff dff_B_U12dkmG22_2(.din(n16153), .dout(n16156));
    jdff dff_B_qYCAoU1x6_2(.din(n16156), .dout(n16159));
    jdff dff_B_P1FziXA14_2(.din(n16159), .dout(n16162));
    jdff dff_B_KtVatRyz5_2(.din(n16162), .dout(n16165));
    jdff dff_B_manjh1NZ5_2(.din(n16165), .dout(n16168));
    jdff dff_B_QTwQ1JIM6_2(.din(n16168), .dout(n16171));
    jdff dff_B_9F3Cheqa6_2(.din(n16171), .dout(n16174));
    jdff dff_B_wYumgaWL6_2(.din(n16174), .dout(n16177));
    jdff dff_B_pCSDMmHc2_2(.din(n16177), .dout(n16180));
    jdff dff_B_WLlRa5yB2_2(.din(n16180), .dout(n16183));
    jdff dff_B_RlF98wIe1_2(.din(n16183), .dout(n16186));
    jdff dff_B_gSOEA2j56_2(.din(n16186), .dout(n16189));
    jdff dff_B_VXDqMmki5_2(.din(n16189), .dout(n16192));
    jdff dff_B_n8gUi5QA1_2(.din(n16192), .dout(n16195));
    jdff dff_B_PX2sR0uv3_2(.din(n16195), .dout(n16198));
    jdff dff_B_ZQyEPytw4_2(.din(n16198), .dout(n16201));
    jdff dff_B_9bhBoudj2_2(.din(n16201), .dout(n16204));
    jdff dff_B_CEJjXlkA2_2(.din(n16204), .dout(n16207));
    jdff dff_B_irtCtgqt4_2(.din(n16207), .dout(n16210));
    jdff dff_B_NtCTb9NO3_2(.din(n16210), .dout(n16213));
    jdff dff_B_QAMRhUhQ1_2(.din(n16213), .dout(n16216));
    jdff dff_B_L3KJJBar3_2(.din(n16216), .dout(n16219));
    jdff dff_B_X3hmDc9U0_2(.din(n16219), .dout(n16222));
    jdff dff_B_t8a7mpJc1_2(.din(n16222), .dout(n16225));
    jdff dff_B_eakJ78K88_2(.din(n16225), .dout(n16228));
    jdff dff_B_7Stnel8r1_2(.din(n16228), .dout(n16231));
    jdff dff_B_qFncmWYE3_2(.din(n16231), .dout(n16234));
    jdff dff_B_NK1cGy002_2(.din(n16234), .dout(n16237));
    jdff dff_B_0RTT3rWU7_2(.din(n16237), .dout(n16240));
    jdff dff_A_LiLLaKQ70_1(.din(n3751), .dout(n16242));
    jdff dff_A_JVFZYS5k2_0(.din(n16248), .dout(n16245));
    jdff dff_A_ThE4032i7_0(.din(n16251), .dout(n16248));
    jdff dff_A_b8dyL3Gc7_0(.din(n16254), .dout(n16251));
    jdff dff_A_MFmMa0Sk5_0(.din(n16257), .dout(n16254));
    jdff dff_A_hNVLQOt59_0(.din(n16260), .dout(n16257));
    jdff dff_A_aNJzPPnh5_0(.din(n16263), .dout(n16260));
    jdff dff_A_sTza9uYR8_0(.din(n16266), .dout(n16263));
    jdff dff_A_ucZrvFil5_0(.din(n16269), .dout(n16266));
    jdff dff_A_rujyZHXO7_0(.din(n16272), .dout(n16269));
    jdff dff_A_BTuUOtKP4_0(.din(n16275), .dout(n16272));
    jdff dff_A_oicvysoX1_0(.din(n16278), .dout(n16275));
    jdff dff_A_tmZXjUZJ1_0(.din(n16281), .dout(n16278));
    jdff dff_A_OP2JCiGM7_0(.din(n16284), .dout(n16281));
    jdff dff_A_X51ycMFW3_0(.din(n16287), .dout(n16284));
    jdff dff_A_ulWJkAd52_0(.din(n16290), .dout(n16287));
    jdff dff_A_wBkthbbs3_0(.din(n16293), .dout(n16290));
    jdff dff_A_efQbvt229_0(.din(n16296), .dout(n16293));
    jdff dff_A_QeXAeT9f6_0(.din(n16299), .dout(n16296));
    jdff dff_A_s7D7sebC2_0(.din(n16302), .dout(n16299));
    jdff dff_A_x885c7Ue6_0(.din(n16305), .dout(n16302));
    jdff dff_A_wiavjYbC8_0(.din(n16308), .dout(n16305));
    jdff dff_A_qLhJBFLE0_0(.din(n16311), .dout(n16308));
    jdff dff_A_1kIhnF6k7_0(.din(n16314), .dout(n16311));
    jdff dff_A_Z84DsC3x1_0(.din(n16317), .dout(n16314));
    jdff dff_A_O8e5PD9S4_0(.din(n16320), .dout(n16317));
    jdff dff_A_mxB2yEn90_0(.din(n16323), .dout(n16320));
    jdff dff_A_VLDufczS1_0(.din(n16326), .dout(n16323));
    jdff dff_A_tyScGpDV5_0(.din(n16329), .dout(n16326));
    jdff dff_A_CrJ0yvYZ5_0(.din(n16332), .dout(n16329));
    jdff dff_A_RrkunfDu4_0(.din(n16335), .dout(n16332));
    jdff dff_A_BZnmWBMG8_0(.din(n16338), .dout(n16335));
    jdff dff_A_JpAY9JLX4_0(.din(n16341), .dout(n16338));
    jdff dff_A_NN1WPiiH7_0(.din(n16344), .dout(n16341));
    jdff dff_A_ElRliAgJ8_0(.din(n16347), .dout(n16344));
    jdff dff_A_DqnCeYFm4_0(.din(n16350), .dout(n16347));
    jdff dff_A_Zrw86vAk2_0(.din(n16353), .dout(n16350));
    jdff dff_A_dfoK9Vu36_0(.din(n16356), .dout(n16353));
    jdff dff_A_PXYu4tFF2_0(.din(n3017), .dout(n16356));
    jdff dff_A_rNhfqppf1_1(.din(n3349), .dout(n16359));
    jdff dff_A_ERUtKZw50_2(.din(n3349), .dout(n16362));
    jdff dff_B_pFzgrlqQ6_1(.din(n3024), .dout(n16366));
    jdff dff_B_aqLqSVbb5_2(.din(n2641), .dout(n16369));
    jdff dff_B_8TtlUCFZ6_2(.din(n16369), .dout(n16372));
    jdff dff_B_fGoWAijM3_2(.din(n16372), .dout(n16375));
    jdff dff_B_LX6g5d3q0_2(.din(n16375), .dout(n16378));
    jdff dff_B_OxgyoqTX1_2(.din(n16378), .dout(n16381));
    jdff dff_B_ePUgQZSz9_2(.din(n16381), .dout(n16384));
    jdff dff_B_855WPIpP8_2(.din(n16384), .dout(n16387));
    jdff dff_B_1SLzG1sJ8_2(.din(n16387), .dout(n16390));
    jdff dff_B_ZONFmFUc2_2(.din(n16390), .dout(n16393));
    jdff dff_B_zgrMX4vu2_2(.din(n16393), .dout(n16396));
    jdff dff_B_CWoryAm58_2(.din(n16396), .dout(n16399));
    jdff dff_B_8PI4HxTW1_2(.din(n16399), .dout(n16402));
    jdff dff_B_W565hlja3_2(.din(n16402), .dout(n16405));
    jdff dff_B_goC2GtdM8_2(.din(n16405), .dout(n16408));
    jdff dff_B_zglewjTh2_2(.din(n16408), .dout(n16411));
    jdff dff_B_NCfsaHxY3_2(.din(n16411), .dout(n16414));
    jdff dff_B_izzFwD9P7_2(.din(n16414), .dout(n16417));
    jdff dff_B_jcVvnAzP3_2(.din(n16417), .dout(n16420));
    jdff dff_B_V8ljW9QM2_2(.din(n16420), .dout(n16423));
    jdff dff_B_RiDZEjDY7_2(.din(n16423), .dout(n16426));
    jdff dff_B_PiUefMaQ9_2(.din(n16426), .dout(n16429));
    jdff dff_B_l17r3wle0_2(.din(n16429), .dout(n16432));
    jdff dff_B_pjpfPEhq9_2(.din(n16432), .dout(n16435));
    jdff dff_B_DVx2s3wq5_2(.din(n16435), .dout(n16438));
    jdff dff_B_73GQfmpV4_2(.din(n16438), .dout(n16441));
    jdff dff_B_iiZJ8oQK7_2(.din(n16441), .dout(n16444));
    jdff dff_B_ETLGqHFC0_2(.din(n16444), .dout(n16447));
    jdff dff_B_wuc06J5x0_2(.din(n16447), .dout(n16450));
    jdff dff_B_2mWbSJ3u6_2(.din(n16450), .dout(n16453));
    jdff dff_B_UVLb67d54_2(.din(n16453), .dout(n16456));
    jdff dff_B_dXYrXhlm3_2(.din(n16456), .dout(n16459));
    jdff dff_B_sNZ6qBcz6_2(.din(n16459), .dout(n16462));
    jdff dff_B_GSt3l0oj2_2(.din(n16462), .dout(n16465));
    jdff dff_B_CGzaqclw9_2(.din(n16465), .dout(n16468));
    jdff dff_B_lsaBQh7J8_2(.din(n2944), .dout(n16471));
    jdff dff_B_YFGLmNff5_1(.din(n2645), .dout(n16474));
    jdff dff_B_qjeV4zON2_2(.din(n2286), .dout(n16477));
    jdff dff_B_8R7Ti3qY2_2(.din(n16477), .dout(n16480));
    jdff dff_B_84YqnIUj2_2(.din(n16480), .dout(n16483));
    jdff dff_B_IJnCaoWh3_2(.din(n16483), .dout(n16486));
    jdff dff_B_0OEM80xx5_2(.din(n16486), .dout(n16489));
    jdff dff_B_uV6ZS0iu8_2(.din(n16489), .dout(n16492));
    jdff dff_B_6Y0S37xe5_2(.din(n16492), .dout(n16495));
    jdff dff_B_lHV9p9xl7_2(.din(n16495), .dout(n16498));
    jdff dff_B_8REZEnvQ1_2(.din(n16498), .dout(n16501));
    jdff dff_B_VqROLeH34_2(.din(n16501), .dout(n16504));
    jdff dff_B_ogbzXqZ74_2(.din(n16504), .dout(n16507));
    jdff dff_B_t8uPvq429_2(.din(n16507), .dout(n16510));
    jdff dff_B_JaALiz3y5_2(.din(n16510), .dout(n16513));
    jdff dff_B_nRCTL3CB6_2(.din(n16513), .dout(n16516));
    jdff dff_B_rZWLath03_2(.din(n16516), .dout(n16519));
    jdff dff_B_8235HZRe8_2(.din(n16519), .dout(n16522));
    jdff dff_B_vj6GeHQl1_2(.din(n16522), .dout(n16525));
    jdff dff_B_wWrx1rJ38_2(.din(n16525), .dout(n16528));
    jdff dff_B_fYft93dk1_2(.din(n16528), .dout(n16531));
    jdff dff_B_3JYrxhaL4_2(.din(n16531), .dout(n16534));
    jdff dff_B_wNm6FKIX1_2(.din(n16534), .dout(n16537));
    jdff dff_B_2itOObFF4_2(.din(n16537), .dout(n16540));
    jdff dff_B_Rzkg6iNm6_2(.din(n16540), .dout(n16543));
    jdff dff_B_MkZbSH8v5_2(.din(n16543), .dout(n16546));
    jdff dff_B_LwCJR8VV8_2(.din(n16546), .dout(n16549));
    jdff dff_B_oPY21CCQ4_2(.din(n16549), .dout(n16552));
    jdff dff_B_vMqCSAr18_2(.din(n16552), .dout(n16555));
    jdff dff_B_vkit0yNc5_2(.din(n16555), .dout(n16558));
    jdff dff_B_LoFVokDw9_2(.din(n16558), .dout(n16561));
    jdff dff_B_JaDhI1AO8_2(.din(n16561), .dout(n16564));
    jdff dff_B_ZYWG448Y6_2(.din(n16564), .dout(n16567));
    jdff dff_B_XMyO4VcL9_2(.din(n2562), .dout(n16570));
    jdff dff_B_p7A5tY8K4_1(.din(n2290), .dout(n16573));
    jdff dff_B_SWE7pXwo9_2(.din(n1958), .dout(n16576));
    jdff dff_B_lOav3PfN0_2(.din(n16576), .dout(n16579));
    jdff dff_B_wFYf2lav8_2(.din(n16579), .dout(n16582));
    jdff dff_B_HZIKFsvb9_2(.din(n16582), .dout(n16585));
    jdff dff_B_R488Rsjb9_2(.din(n16585), .dout(n16588));
    jdff dff_B_098UAozT5_2(.din(n16588), .dout(n16591));
    jdff dff_B_iFUaAVA13_2(.din(n16591), .dout(n16594));
    jdff dff_B_IWrhjz9Z0_2(.din(n16594), .dout(n16597));
    jdff dff_B_4J5QOlcx4_2(.din(n16597), .dout(n16600));
    jdff dff_B_xfOBvoTR5_2(.din(n16600), .dout(n16603));
    jdff dff_B_03J3pO6K2_2(.din(n16603), .dout(n16606));
    jdff dff_B_aZn31KFm0_2(.din(n16606), .dout(n16609));
    jdff dff_B_226Xofee5_2(.din(n16609), .dout(n16612));
    jdff dff_B_lhKvZDVA2_2(.din(n16612), .dout(n16615));
    jdff dff_B_itQyYcEO2_2(.din(n16615), .dout(n16618));
    jdff dff_B_v2OoYA8f8_2(.din(n16618), .dout(n16621));
    jdff dff_B_w06hzSZz7_2(.din(n16621), .dout(n16624));
    jdff dff_B_TVmd71Bt5_2(.din(n16624), .dout(n16627));
    jdff dff_B_gAUP2gyM6_2(.din(n16627), .dout(n16630));
    jdff dff_B_pGZDE7MI4_2(.din(n16630), .dout(n16633));
    jdff dff_B_FF3Y9FHH8_2(.din(n16633), .dout(n16636));
    jdff dff_B_TlxNAIKP7_2(.din(n16636), .dout(n16639));
    jdff dff_B_uSV59Dl34_2(.din(n16639), .dout(n16642));
    jdff dff_B_r445SAU90_2(.din(n16642), .dout(n16645));
    jdff dff_B_pWXeHk9R5_2(.din(n16645), .dout(n16648));
    jdff dff_B_sVujVXx70_2(.din(n16648), .dout(n16651));
    jdff dff_B_IvwcZuZ52_2(.din(n16651), .dout(n16654));
    jdff dff_B_IqjvnNs23_2(.din(n16654), .dout(n16657));
    jdff dff_B_A0EP2u038_2(.din(n2207), .dout(n16660));
    jdff dff_B_LdbHXJz70_1(.din(n1962), .dout(n16663));
    jdff dff_B_remLdU3W7_2(.din(n1657), .dout(n16666));
    jdff dff_B_nSCTjnSp5_2(.din(n16666), .dout(n16669));
    jdff dff_B_EmZUjoei5_2(.din(n16669), .dout(n16672));
    jdff dff_B_kzvdLuxQ4_2(.din(n16672), .dout(n16675));
    jdff dff_B_j0nqz0qI3_2(.din(n16675), .dout(n16678));
    jdff dff_B_UF4stipx1_2(.din(n16678), .dout(n16681));
    jdff dff_B_Ong0mR9n3_2(.din(n16681), .dout(n16684));
    jdff dff_B_BoG9dJsj3_2(.din(n16684), .dout(n16687));
    jdff dff_B_4l8CMNvt4_2(.din(n16687), .dout(n16690));
    jdff dff_B_0AtmG2Cn7_2(.din(n16690), .dout(n16693));
    jdff dff_B_vaaTdudL8_2(.din(n16693), .dout(n16696));
    jdff dff_B_fJqk2wzJ0_2(.din(n16696), .dout(n16699));
    jdff dff_B_FPlSDfho2_2(.din(n16699), .dout(n16702));
    jdff dff_B_FukND1Vq8_2(.din(n16702), .dout(n16705));
    jdff dff_B_g0Om3uaU4_2(.din(n16705), .dout(n16708));
    jdff dff_B_Pj0dZwwN3_2(.din(n16708), .dout(n16711));
    jdff dff_B_Bh7jb3Mx6_2(.din(n16711), .dout(n16714));
    jdff dff_B_ffTQWIFS5_2(.din(n16714), .dout(n16717));
    jdff dff_B_wLMNGDU23_2(.din(n16717), .dout(n16720));
    jdff dff_B_A3BrkMmV3_2(.din(n16720), .dout(n16723));
    jdff dff_B_gSujsVYH1_2(.din(n16723), .dout(n16726));
    jdff dff_B_qErqbt8q0_2(.din(n16726), .dout(n16729));
    jdff dff_B_fOtmj0Vl2_2(.din(n16729), .dout(n16732));
    jdff dff_B_G3PK9Dmz9_2(.din(n16732), .dout(n16735));
    jdff dff_B_YZsqRtp03_2(.din(n16735), .dout(n16738));
    jdff dff_B_ahnDQaUE2_2(.din(n1879), .dout(n16741));
    jdff dff_B_VdB4vGKp5_1(.din(n1661), .dout(n16744));
    jdff dff_B_2VwStOel9_2(.din(n1383), .dout(n16747));
    jdff dff_B_kLxdcguU7_2(.din(n16747), .dout(n16750));
    jdff dff_B_7jOyGxjd9_2(.din(n16750), .dout(n16753));
    jdff dff_B_iAYneITv0_2(.din(n16753), .dout(n16756));
    jdff dff_B_7W1gMF8E6_2(.din(n16756), .dout(n16759));
    jdff dff_B_4heQCxFT6_2(.din(n16759), .dout(n16762));
    jdff dff_B_BmKSXrJd4_2(.din(n16762), .dout(n16765));
    jdff dff_B_YIhP0J3W2_2(.din(n16765), .dout(n16768));
    jdff dff_B_DxH8y57k0_2(.din(n16768), .dout(n16771));
    jdff dff_B_DxkGXL4K2_2(.din(n16771), .dout(n16774));
    jdff dff_B_LG1DRUM75_2(.din(n16774), .dout(n16777));
    jdff dff_B_gwkAKuOX3_2(.din(n16777), .dout(n16780));
    jdff dff_B_HZIXzl9R1_2(.din(n16780), .dout(n16783));
    jdff dff_B_t0YiUaOj3_2(.din(n16783), .dout(n16786));
    jdff dff_B_XaEkSQOJ5_2(.din(n16786), .dout(n16789));
    jdff dff_B_Ieuytx2k1_2(.din(n16789), .dout(n16792));
    jdff dff_B_rVH2xRnM3_2(.din(n16792), .dout(n16795));
    jdff dff_B_MNSiRIMK9_2(.din(n16795), .dout(n16798));
    jdff dff_B_gIFGXc919_2(.din(n16798), .dout(n16801));
    jdff dff_B_CrCxR1cm2_2(.din(n16801), .dout(n16804));
    jdff dff_B_gQ6syMS02_2(.din(n16804), .dout(n16807));
    jdff dff_B_B1MHIwkE4_2(.din(n16807), .dout(n16810));
    jdff dff_B_oai99Er00_2(.din(n1578), .dout(n16813));
    jdff dff_B_Ha01Stdo7_1(.din(n1387), .dout(n16816));
    jdff dff_B_kPzXdT731_2(.din(n1139), .dout(n16819));
    jdff dff_B_rtyGdkVm1_2(.din(n16819), .dout(n16822));
    jdff dff_B_vhAZV4Tc4_2(.din(n16822), .dout(n16825));
    jdff dff_B_gWd43pn36_2(.din(n16825), .dout(n16828));
    jdff dff_B_ZdFhonGr4_2(.din(n16828), .dout(n16831));
    jdff dff_B_Rtwqnh0h5_2(.din(n16831), .dout(n16834));
    jdff dff_B_HNe5PlZm0_2(.din(n16834), .dout(n16837));
    jdff dff_B_3SxQLx4g3_2(.din(n16837), .dout(n16840));
    jdff dff_B_okHSrSDq9_2(.din(n16840), .dout(n16843));
    jdff dff_B_3B9sHaTO1_2(.din(n16843), .dout(n16846));
    jdff dff_B_jpsQrg4H5_2(.din(n16846), .dout(n16849));
    jdff dff_B_DsHnBPqt4_2(.din(n16849), .dout(n16852));
    jdff dff_B_jZdjHIib2_2(.din(n16852), .dout(n16855));
    jdff dff_B_DBAuNXme7_2(.din(n16855), .dout(n16858));
    jdff dff_B_Z1xPljwx3_2(.din(n16858), .dout(n16861));
    jdff dff_B_a779KKf65_2(.din(n16861), .dout(n16864));
    jdff dff_B_t1I5GBDE3_2(.din(n16864), .dout(n16867));
    jdff dff_B_pLjYX2P31_2(.din(n16867), .dout(n16870));
    jdff dff_B_Jv3A2qaZ9_2(.din(n16870), .dout(n16873));
    jdff dff_B_rbZL3TVO2_2(.din(n1304), .dout(n16876));
    jdff dff_B_QhBkAYhP6_1(.din(n1143), .dout(n16879));
    jdff dff_B_3yKfvuf39_2(.din(n919), .dout(n16882));
    jdff dff_B_QAyCvtyq7_2(.din(n16882), .dout(n16885));
    jdff dff_B_Ob3yL81s1_2(.din(n16885), .dout(n16888));
    jdff dff_B_SW0GfjWC1_2(.din(n16888), .dout(n16891));
    jdff dff_B_pdfeUBWc5_2(.din(n16891), .dout(n16894));
    jdff dff_B_bzFlRNgb6_2(.din(n16894), .dout(n16897));
    jdff dff_B_reD8dfdd1_2(.din(n16897), .dout(n16900));
    jdff dff_B_HlnvGXCL2_2(.din(n16900), .dout(n16903));
    jdff dff_B_9R9D6Qrj3_2(.din(n16903), .dout(n16906));
    jdff dff_B_685BWqiP9_2(.din(n16906), .dout(n16909));
    jdff dff_B_OjdGeNKJ3_2(.din(n16909), .dout(n16912));
    jdff dff_B_ryEQoQyp0_2(.din(n16912), .dout(n16915));
    jdff dff_B_snitgZz50_2(.din(n16915), .dout(n16918));
    jdff dff_B_2EI7hVaw4_2(.din(n16918), .dout(n16921));
    jdff dff_B_1Huhmroh3_2(.din(n16921), .dout(n16924));
    jdff dff_B_OnVhSGaU0_2(.din(n16924), .dout(n16927));
    jdff dff_B_Flxa6Eko8_2(.din(n1060), .dout(n16930));
    jdff dff_B_6Fhf9Eju8_1(.din(n923), .dout(n16933));
    jdff dff_B_7OpAxnXt7_2(.din(n726), .dout(n16936));
    jdff dff_B_j0cy7ffD7_2(.din(n16936), .dout(n16939));
    jdff dff_B_Peeqc6VE0_2(.din(n16939), .dout(n16942));
    jdff dff_B_3ekBNrqu2_2(.din(n16942), .dout(n16945));
    jdff dff_B_Tvh1sZvk8_2(.din(n16945), .dout(n16948));
    jdff dff_B_iKrspdTh0_2(.din(n16948), .dout(n16951));
    jdff dff_B_NT2WauMy1_2(.din(n16951), .dout(n16954));
    jdff dff_B_OW93GX1A8_2(.din(n16954), .dout(n16957));
    jdff dff_B_wPlQyK8K5_2(.din(n16957), .dout(n16960));
    jdff dff_B_3gwdVvUv7_2(.din(n16960), .dout(n16963));
    jdff dff_B_QcrKqKi74_2(.din(n16963), .dout(n16966));
    jdff dff_B_7XhZKsfy9_2(.din(n16966), .dout(n16969));
    jdff dff_B_7t7VuDNg2_2(.din(n16969), .dout(n16972));
    jdff dff_B_5WzUuFtq7_2(.din(n840), .dout(n16975));
    jdff dff_B_ncfFgBcp6_1(.din(n730), .dout(n16978));
    jdff dff_B_1SQv2chZ3_2(.din(n563), .dout(n16981));
    jdff dff_B_kaNBOWuF6_2(.din(n16981), .dout(n16984));
    jdff dff_B_pMy8k2Y10_2(.din(n16984), .dout(n16987));
    jdff dff_B_CPnvODoO8_2(.din(n16987), .dout(n16990));
    jdff dff_B_BsS1fQvf8_2(.din(n16990), .dout(n16993));
    jdff dff_B_4KO8A3aG2_2(.din(n16993), .dout(n16996));
    jdff dff_B_WoJonN7K9_2(.din(n16996), .dout(n16999));
    jdff dff_B_cFRAFIlK7_2(.din(n16999), .dout(n17002));
    jdff dff_B_sE7s3cCi0_2(.din(n17002), .dout(n17005));
    jdff dff_B_2BHgDr6f3_2(.din(n17005), .dout(n17008));
    jdff dff_B_Hwp7sJGy6_2(.din(n647), .dout(n17011));
    jdff dff_B_Rn758qRw2_1(.din(n567), .dout(n17014));
    jdff dff_B_245dB2Vj1_2(.din(n419), .dout(n17017));
    jdff dff_B_GxmnUU2i9_2(.din(n17017), .dout(n17020));
    jdff dff_B_qMjk9fbg4_2(.din(n17020), .dout(n17023));
    jdff dff_B_HfWphmhP3_2(.din(n17023), .dout(n17026));
    jdff dff_B_QZE1CIaw1_2(.din(n17026), .dout(n17029));
    jdff dff_B_ht3rygSr0_2(.din(n17029), .dout(n17032));
    jdff dff_B_E9bULjDw7_2(.din(n17032), .dout(n17035));
    jdff dff_B_U2AtfufT8_2(.din(n484), .dout(n17038));
    jdff dff_B_6BySlTG00_1(.din(n430), .dout(n17041));
    jdff dff_B_jyMdLAoA5_1(.din(n17041), .dout(n17044));
    jdff dff_B_55AhhSfT5_2(.din(n306), .dout(n17047));
    jdff dff_B_AR0OBn1x1_2(.din(n17047), .dout(n17050));
    jdff dff_B_SKN6sspX6_2(.din(n17050), .dout(n17053));
    jdff dff_B_uXlhIgzZ4_2(.din(n17053), .dout(n17056));
    jdff dff_A_bcg8oVQH4_1(.din(n314), .dout(n17058));
    jdff dff_A_1G0AuNFk3_0(.din(n204), .dout(n17061));
    jdff dff_A_avonoj9j1_0(.din(n201), .dout(n17064));
    jdff dff_A_ixNCcfTv9_1(.din(n201), .dout(n17067));
    jdff dff_A_ir0jkoTy5_2(.din(n17073), .dout(n17070));
    jdff dff_A_srC73IwU0_2(.din(n201), .dout(n17073));
    jdff dff_B_iWR1jGX20_0(.din(n4889), .dout(n17077));
    jdff dff_A_vNJLJ28L9_1(.din(n17082), .dout(n17079));
    jdff dff_A_nsNq7sN28_1(.din(n4875), .dout(n17082));
    jdff dff_B_YGmA32BL2_1(.din(n4566), .dout(n17086));
    jdff dff_B_Xe2jUCZn7_1(.din(n17086), .dout(n17089));
    jdff dff_B_VrfINGLF2_2(.din(n4210), .dout(n17092));
    jdff dff_B_XRfA1XNS1_2(.din(n17092), .dout(n17095));
    jdff dff_B_OcDoaZCJ1_2(.din(n17095), .dout(n17098));
    jdff dff_B_TgjGHPTz1_2(.din(n17098), .dout(n17101));
    jdff dff_B_uirphLHQ6_2(.din(n17101), .dout(n17104));
    jdff dff_B_pXrGjQ6a9_2(.din(n17104), .dout(n17107));
    jdff dff_B_z75aXurF5_2(.din(n17107), .dout(n17110));
    jdff dff_B_gMdAcu1U7_2(.din(n17110), .dout(n17113));
    jdff dff_B_SAinsTPC1_2(.din(n17113), .dout(n17116));
    jdff dff_B_Vz6fifrE0_2(.din(n17116), .dout(n17119));
    jdff dff_B_G7rr8G725_2(.din(n17119), .dout(n17122));
    jdff dff_B_I2mQM6LX9_2(.din(n17122), .dout(n17125));
    jdff dff_B_QUJcTRdT2_2(.din(n17125), .dout(n17128));
    jdff dff_B_2BGDN8B65_2(.din(n17128), .dout(n17131));
    jdff dff_B_hBQWltrx1_2(.din(n17131), .dout(n17134));
    jdff dff_B_TdXrTcUA7_2(.din(n17134), .dout(n17137));
    jdff dff_B_IpKsEiml0_2(.din(n17137), .dout(n17140));
    jdff dff_B_VgYxqRs84_2(.din(n17140), .dout(n17143));
    jdff dff_B_Jr4pzSBm6_2(.din(n17143), .dout(n17146));
    jdff dff_B_9v4AewAA1_2(.din(n17146), .dout(n17149));
    jdff dff_B_sUyJAQLP2_2(.din(n17149), .dout(n17152));
    jdff dff_B_iIaN59k97_2(.din(n17152), .dout(n17155));
    jdff dff_B_7STjTvPY6_2(.din(n17155), .dout(n17158));
    jdff dff_B_SrNRAmR12_2(.din(n17158), .dout(n17161));
    jdff dff_B_O8jpz1An2_2(.din(n17161), .dout(n17164));
    jdff dff_B_7T1mB0cm9_2(.din(n17164), .dout(n17167));
    jdff dff_B_DmaFqNAH0_2(.din(n17167), .dout(n17170));
    jdff dff_B_WobrmUQu2_2(.din(n17170), .dout(n17173));
    jdff dff_B_D2JmnkdL1_2(.din(n17173), .dout(n17176));
    jdff dff_B_tpgvJ9CA8_2(.din(n17176), .dout(n17179));
    jdff dff_B_BSOTueR98_2(.din(n17179), .dout(n17182));
    jdff dff_B_VQH5x6mD1_2(.din(n17182), .dout(n17185));
    jdff dff_B_EbjNuSer1_2(.din(n17185), .dout(n17188));
    jdff dff_B_ka8jStj19_2(.din(n17188), .dout(n17191));
    jdff dff_B_kNTlWiqX7_2(.din(n17191), .dout(n17194));
    jdff dff_B_afMCcITk5_2(.din(n17194), .dout(n17197));
    jdff dff_B_bpOdG4iR4_2(.din(n17197), .dout(n17200));
    jdff dff_B_EH4SD5so8_2(.din(n17200), .dout(n17203));
    jdff dff_B_ebJun9CI7_2(.din(n17203), .dout(n17206));
    jdff dff_B_Rk1dtwek0_2(.din(n17206), .dout(n17209));
    jdff dff_B_71HUwSnK0_2(.din(n17209), .dout(n17212));
    jdff dff_B_dZZyLqHf4_2(.din(n17212), .dout(n17215));
    jdff dff_B_QSRCM4is5_2(.din(n17215), .dout(n17218));
    jdff dff_B_yiuIGVGX8_2(.din(n17218), .dout(n17221));
    jdff dff_B_fZaMNZMF5_2(.din(n17221), .dout(n17224));
    jdff dff_B_la2T5edW5_2(.din(n17224), .dout(n17227));
    jdff dff_B_GIJup5jm6_2(.din(n4525), .dout(n17230));
    jdff dff_B_KiUGehzL6_1(.din(n4217), .dout(n17233));
    jdff dff_B_rewq4jsN8_2(.din(n3817), .dout(n17236));
    jdff dff_B_FsJAHL7T8_2(.din(n17236), .dout(n17239));
    jdff dff_B_DxbEk9Do7_2(.din(n17239), .dout(n17242));
    jdff dff_B_qk9p5GUp6_2(.din(n17242), .dout(n17245));
    jdff dff_B_HZN6197g9_2(.din(n17245), .dout(n17248));
    jdff dff_B_ItHsGKyE2_2(.din(n17248), .dout(n17251));
    jdff dff_B_hRMkurKu0_2(.din(n17251), .dout(n17254));
    jdff dff_B_10g616Fd4_2(.din(n17254), .dout(n17257));
    jdff dff_B_AjD8ZvoK2_2(.din(n17257), .dout(n17260));
    jdff dff_B_EsPpHUED9_2(.din(n17260), .dout(n17263));
    jdff dff_B_z4QvrVIP4_2(.din(n17263), .dout(n17266));
    jdff dff_B_EdUwjeuf8_2(.din(n17266), .dout(n17269));
    jdff dff_B_nYnp5rFQ8_2(.din(n17269), .dout(n17272));
    jdff dff_B_aRSQi7JQ7_2(.din(n17272), .dout(n17275));
    jdff dff_B_5C1Bkj3z8_2(.din(n17275), .dout(n17278));
    jdff dff_B_FNBeGY117_2(.din(n17278), .dout(n17281));
    jdff dff_B_TQGFwaNc2_2(.din(n17281), .dout(n17284));
    jdff dff_B_nMaRYxcD2_2(.din(n17284), .dout(n17287));
    jdff dff_B_EqTgjE9Q8_2(.din(n17287), .dout(n17290));
    jdff dff_B_wSvHJhfE2_2(.din(n17290), .dout(n17293));
    jdff dff_B_Cm294iTF6_2(.din(n17293), .dout(n17296));
    jdff dff_B_xmhdO6RH9_2(.din(n17296), .dout(n17299));
    jdff dff_B_xtH2xk4b5_2(.din(n17299), .dout(n17302));
    jdff dff_B_9c9MD8zi2_2(.din(n17302), .dout(n17305));
    jdff dff_B_yRBYk8Oe2_2(.din(n17305), .dout(n17308));
    jdff dff_B_MGHYPV087_2(.din(n17308), .dout(n17311));
    jdff dff_B_yE4eQ1Uh3_2(.din(n17311), .dout(n17314));
    jdff dff_B_TqRH4DC72_2(.din(n17314), .dout(n17317));
    jdff dff_B_QTy9EYpY8_2(.din(n17317), .dout(n17320));
    jdff dff_B_LR2IAJHR2_2(.din(n17320), .dout(n17323));
    jdff dff_B_u2lXHmpz3_2(.din(n17323), .dout(n17326));
    jdff dff_B_9sNQnnWr0_2(.din(n17326), .dout(n17329));
    jdff dff_B_JvxBIJkd5_2(.din(n17329), .dout(n17332));
    jdff dff_B_bdNK3aFA1_2(.din(n17332), .dout(n17335));
    jdff dff_B_OXb66QLL0_2(.din(n17335), .dout(n17338));
    jdff dff_B_ui7AadZK3_2(.din(n17338), .dout(n17341));
    jdff dff_B_acAocIjr2_2(.din(n17341), .dout(n17344));
    jdff dff_B_uObjiOEf1_2(.din(n17344), .dout(n17347));
    jdff dff_B_RP3MClyb5_2(.din(n17347), .dout(n17350));
    jdff dff_B_6ZcaJYfa8_2(.din(n17350), .dout(n17353));
    jdff dff_B_hSsYxRe46_2(.din(n17353), .dout(n17356));
    jdff dff_B_LLAZKhDn3_2(.din(n17356), .dout(n17359));
    jdff dff_B_4OqqlQj08_2(.din(n4146), .dout(n17362));
    jdff dff_B_877gKBVH1_1(.din(n3821), .dout(n17365));
    jdff dff_B_5jft2Vwy6_2(.din(n3440), .dout(n17368));
    jdff dff_B_ZN8TJwuQ8_2(.din(n17368), .dout(n17371));
    jdff dff_B_zTZjp51P1_2(.din(n17371), .dout(n17374));
    jdff dff_B_hUvwZgQR1_2(.din(n17374), .dout(n17377));
    jdff dff_B_FVNmkt943_2(.din(n17377), .dout(n17380));
    jdff dff_B_sXLylmgx7_2(.din(n17380), .dout(n17383));
    jdff dff_B_WANgA7vs3_2(.din(n17383), .dout(n17386));
    jdff dff_B_fCC3zs2y6_2(.din(n17386), .dout(n17389));
    jdff dff_B_x2qKhbFB6_2(.din(n17389), .dout(n17392));
    jdff dff_B_GUNSKsCY0_2(.din(n17392), .dout(n17395));
    jdff dff_B_iQmc28Lc0_2(.din(n17395), .dout(n17398));
    jdff dff_B_uY4a52hs4_2(.din(n17398), .dout(n17401));
    jdff dff_B_3iCrlnnm9_2(.din(n17401), .dout(n17404));
    jdff dff_B_LJLGwmyK7_2(.din(n17404), .dout(n17407));
    jdff dff_B_NV4ochvg1_2(.din(n17407), .dout(n17410));
    jdff dff_B_cTAZdZuN9_2(.din(n17410), .dout(n17413));
    jdff dff_B_PrHX0WOD4_2(.din(n17413), .dout(n17416));
    jdff dff_B_rxkKwHsc1_2(.din(n17416), .dout(n17419));
    jdff dff_B_8rmTXVCC1_2(.din(n17419), .dout(n17422));
    jdff dff_B_6nCHpHQ83_2(.din(n17422), .dout(n17425));
    jdff dff_B_v9bxAY7j3_2(.din(n17425), .dout(n17428));
    jdff dff_B_dkFlagy72_2(.din(n17428), .dout(n17431));
    jdff dff_B_aXPHQdB68_2(.din(n17431), .dout(n17434));
    jdff dff_B_dnoxVV8M8_2(.din(n17434), .dout(n17437));
    jdff dff_B_siVuMN1S1_2(.din(n17437), .dout(n17440));
    jdff dff_B_OvKBIR2v5_2(.din(n17440), .dout(n17443));
    jdff dff_B_VGwR5a5V8_2(.din(n17443), .dout(n17446));
    jdff dff_B_PfZATf5Z7_2(.din(n17446), .dout(n17449));
    jdff dff_B_JO5e3owO8_2(.din(n17449), .dout(n17452));
    jdff dff_B_QOIGMBCv0_2(.din(n17452), .dout(n17455));
    jdff dff_B_cOEeJdOO5_2(.din(n17455), .dout(n17458));
    jdff dff_B_bLVjfL3e5_2(.din(n17458), .dout(n17461));
    jdff dff_B_RaWgKTIy8_2(.din(n17461), .dout(n17464));
    jdff dff_B_l22DOOKi2_2(.din(n17464), .dout(n17467));
    jdff dff_B_0GbXCiTa4_2(.din(n17467), .dout(n17470));
    jdff dff_B_ET3KHaJ89_2(.din(n17470), .dout(n17473));
    jdff dff_B_zFBisT5P4_2(.din(n17473), .dout(n17476));
    jdff dff_B_lwCdysTz7_2(.din(n3743), .dout(n17479));
    jdff dff_B_vxmO1t5E1_1(.din(n3444), .dout(n17482));
    jdff dff_B_KgNEIDdg7_2(.din(n3039), .dout(n17485));
    jdff dff_B_DyOciAqY6_2(.din(n17485), .dout(n17488));
    jdff dff_B_AO610JJm0_2(.din(n17488), .dout(n17491));
    jdff dff_B_4Bx7eUcR0_2(.din(n17491), .dout(n17494));
    jdff dff_B_Dce8WUZR6_2(.din(n17494), .dout(n17497));
    jdff dff_B_NTm7gPf28_2(.din(n17497), .dout(n17500));
    jdff dff_B_fU6SomYh0_2(.din(n17500), .dout(n17503));
    jdff dff_B_OdaSii8Z4_2(.din(n17503), .dout(n17506));
    jdff dff_B_1niVhtcy2_2(.din(n17506), .dout(n17509));
    jdff dff_B_GstPYLjk1_2(.din(n17509), .dout(n17512));
    jdff dff_B_T8Spe6jd9_2(.din(n17512), .dout(n17515));
    jdff dff_B_lPRBVp1C3_2(.din(n17515), .dout(n17518));
    jdff dff_B_pwA5AzaO2_2(.din(n17518), .dout(n17521));
    jdff dff_B_BI5zecxF9_2(.din(n17521), .dout(n17524));
    jdff dff_B_Rf3UPpIJ2_2(.din(n17524), .dout(n17527));
    jdff dff_B_NJz4azqW1_2(.din(n17527), .dout(n17530));
    jdff dff_B_NfQ241217_2(.din(n17530), .dout(n17533));
    jdff dff_B_awfMdEK42_2(.din(n17533), .dout(n17536));
    jdff dff_B_0PeRm2hj5_2(.din(n17536), .dout(n17539));
    jdff dff_B_Qmg3mdtc5_2(.din(n17539), .dout(n17542));
    jdff dff_B_wG7tUDtG6_2(.din(n17542), .dout(n17545));
    jdff dff_B_oB2hDlLM6_2(.din(n17545), .dout(n17548));
    jdff dff_B_P7fByLw52_2(.din(n17548), .dout(n17551));
    jdff dff_B_4lr70A8b7_2(.din(n17551), .dout(n17554));
    jdff dff_B_dhwmhWxF1_2(.din(n17554), .dout(n17557));
    jdff dff_B_jl7oPzYT6_2(.din(n17557), .dout(n17560));
    jdff dff_B_2extvQgJ6_2(.din(n17560), .dout(n17563));
    jdff dff_B_AuJWx6rf1_2(.din(n17563), .dout(n17566));
    jdff dff_B_tLaxWX5T1_2(.din(n17566), .dout(n17569));
    jdff dff_B_bBV8Rk6E4_2(.din(n17569), .dout(n17572));
    jdff dff_B_HpW7zvZH0_2(.din(n17572), .dout(n17575));
    jdff dff_B_EipvCePu1_2(.din(n17575), .dout(n17578));
    jdff dff_B_l7FlFbyc1_2(.din(n17578), .dout(n17581));
    jdff dff_B_X2kT5Udq3_2(.din(n17581), .dout(n17584));
    jdff dff_B_6Gtr6lbk5_2(.din(n3341), .dout(n17587));
    jdff dff_B_pkXP9ILj6_1(.din(n3043), .dout(n17590));
    jdff dff_B_7T2LisQI8_2(.din(n2660), .dout(n17593));
    jdff dff_B_83iD7Qxu4_2(.din(n17593), .dout(n17596));
    jdff dff_B_4jDij4Gy4_2(.din(n17596), .dout(n17599));
    jdff dff_B_7JujXeVW3_2(.din(n17599), .dout(n17602));
    jdff dff_B_Y591g1cA7_2(.din(n17602), .dout(n17605));
    jdff dff_B_OPsknhG53_2(.din(n17605), .dout(n17608));
    jdff dff_B_Oet3mOMN6_2(.din(n17608), .dout(n17611));
    jdff dff_B_dzqTfCik5_2(.din(n17611), .dout(n17614));
    jdff dff_B_5eDO5SmG6_2(.din(n17614), .dout(n17617));
    jdff dff_B_jPoroVdG8_2(.din(n17617), .dout(n17620));
    jdff dff_B_iIynPmaY5_2(.din(n17620), .dout(n17623));
    jdff dff_B_4aihdRmi2_2(.din(n17623), .dout(n17626));
    jdff dff_B_O3vtcIue1_2(.din(n17626), .dout(n17629));
    jdff dff_B_GinTlZ4E5_2(.din(n17629), .dout(n17632));
    jdff dff_B_8hOLKX822_2(.din(n17632), .dout(n17635));
    jdff dff_B_D4wy2Okt0_2(.din(n17635), .dout(n17638));
    jdff dff_B_zogtRBeB2_2(.din(n17638), .dout(n17641));
    jdff dff_B_kcYT7JJE9_2(.din(n17641), .dout(n17644));
    jdff dff_B_h74PmwWU9_2(.din(n17644), .dout(n17647));
    jdff dff_B_fxamom8A5_2(.din(n17647), .dout(n17650));
    jdff dff_B_7plIDstX4_2(.din(n17650), .dout(n17653));
    jdff dff_B_zwt3KlqH6_2(.din(n17653), .dout(n17656));
    jdff dff_B_F0e8ypID5_2(.din(n17656), .dout(n17659));
    jdff dff_B_INyCAKn87_2(.din(n17659), .dout(n17662));
    jdff dff_B_bG8EAJce6_2(.din(n17662), .dout(n17665));
    jdff dff_B_zqeQsN1F0_2(.din(n17665), .dout(n17668));
    jdff dff_B_vGlcpdYO4_2(.din(n17668), .dout(n17671));
    jdff dff_B_EGrDx8bY8_2(.din(n17671), .dout(n17674));
    jdff dff_B_M3k35jO77_2(.din(n17674), .dout(n17677));
    jdff dff_B_V8sBfmYO8_2(.din(n17677), .dout(n17680));
    jdff dff_B_HMm1T04d9_2(.din(n17680), .dout(n17683));
    jdff dff_B_pf4x7cqt6_2(.din(n2936), .dout(n17686));
    jdff dff_B_BJRhwV3R5_1(.din(n2664), .dout(n17689));
    jdff dff_B_BQnm9l3F7_2(.din(n2305), .dout(n17692));
    jdff dff_B_0fs6jalb2_2(.din(n17692), .dout(n17695));
    jdff dff_B_tWegmQyn5_2(.din(n17695), .dout(n17698));
    jdff dff_B_c8BeTa936_2(.din(n17698), .dout(n17701));
    jdff dff_B_UT333E6g5_2(.din(n17701), .dout(n17704));
    jdff dff_B_7aK2YLmc4_2(.din(n17704), .dout(n17707));
    jdff dff_B_YSRAgxvZ2_2(.din(n17707), .dout(n17710));
    jdff dff_B_hZO859T94_2(.din(n17710), .dout(n17713));
    jdff dff_B_Rjud5mMf3_2(.din(n17713), .dout(n17716));
    jdff dff_B_jKvJFixD2_2(.din(n17716), .dout(n17719));
    jdff dff_B_o2SywZtH9_2(.din(n17719), .dout(n17722));
    jdff dff_B_3K0e5WII4_2(.din(n17722), .dout(n17725));
    jdff dff_B_FM3HVfhi8_2(.din(n17725), .dout(n17728));
    jdff dff_B_zWDUI0Me3_2(.din(n17728), .dout(n17731));
    jdff dff_B_avZ27p1p6_2(.din(n17731), .dout(n17734));
    jdff dff_B_NEm5x4Wc3_2(.din(n17734), .dout(n17737));
    jdff dff_B_C5PNdhBg2_2(.din(n17737), .dout(n17740));
    jdff dff_B_VKCtOqN43_2(.din(n17740), .dout(n17743));
    jdff dff_B_lUwmlAeX7_2(.din(n17743), .dout(n17746));
    jdff dff_B_Fbiezlze8_2(.din(n17746), .dout(n17749));
    jdff dff_B_nufP5pcR3_2(.din(n17749), .dout(n17752));
    jdff dff_B_uakW9DrU9_2(.din(n17752), .dout(n17755));
    jdff dff_B_p9UZvedm1_2(.din(n17755), .dout(n17758));
    jdff dff_B_eucCY8Co8_2(.din(n17758), .dout(n17761));
    jdff dff_B_HTzDBLQN1_2(.din(n17761), .dout(n17764));
    jdff dff_B_LJb31AHq0_2(.din(n17764), .dout(n17767));
    jdff dff_B_DzISyPcN3_2(.din(n17767), .dout(n17770));
    jdff dff_B_ovFfKiA53_2(.din(n17770), .dout(n17773));
    jdff dff_B_LjFoFNip1_2(.din(n2554), .dout(n17776));
    jdff dff_B_yk77LfyS1_1(.din(n2309), .dout(n17779));
    jdff dff_B_vX247xk67_2(.din(n1977), .dout(n17782));
    jdff dff_B_sokSTcOG0_2(.din(n17782), .dout(n17785));
    jdff dff_B_Au02DbKr4_2(.din(n17785), .dout(n17788));
    jdff dff_B_xAKdDGgk1_2(.din(n17788), .dout(n17791));
    jdff dff_B_CKOuBb2H3_2(.din(n17791), .dout(n17794));
    jdff dff_B_J4gbxKKz7_2(.din(n17794), .dout(n17797));
    jdff dff_B_HmJft7fe1_2(.din(n17797), .dout(n17800));
    jdff dff_B_0o4AMnh69_2(.din(n17800), .dout(n17803));
    jdff dff_B_uotRdzng1_2(.din(n17803), .dout(n17806));
    jdff dff_B_7k9pINyR9_2(.din(n17806), .dout(n17809));
    jdff dff_B_yzGc4yFe4_2(.din(n17809), .dout(n17812));
    jdff dff_B_nNtGhztX6_2(.din(n17812), .dout(n17815));
    jdff dff_B_C3pVjf5o5_2(.din(n17815), .dout(n17818));
    jdff dff_B_SiadrbWM7_2(.din(n17818), .dout(n17821));
    jdff dff_B_VByJf3059_2(.din(n17821), .dout(n17824));
    jdff dff_B_yH2hGQCi7_2(.din(n17824), .dout(n17827));
    jdff dff_B_PHYtLVdL3_2(.din(n17827), .dout(n17830));
    jdff dff_B_aWFLV4zV8_2(.din(n17830), .dout(n17833));
    jdff dff_B_VreCK2Zn9_2(.din(n17833), .dout(n17836));
    jdff dff_B_vhbocJP33_2(.din(n17836), .dout(n17839));
    jdff dff_B_b36eqfI50_2(.din(n17839), .dout(n17842));
    jdff dff_B_tsznxY1O7_2(.din(n17842), .dout(n17845));
    jdff dff_B_cqMgiee46_2(.din(n17845), .dout(n17848));
    jdff dff_B_euIm4nAl6_2(.din(n17848), .dout(n17851));
    jdff dff_B_tVGUx8Nc5_2(.din(n17851), .dout(n17854));
    jdff dff_B_KPzLWWr84_2(.din(n2199), .dout(n17857));
    jdff dff_B_sfAyzdid9_1(.din(n1981), .dout(n17860));
    jdff dff_B_tBziSE9s9_2(.din(n1676), .dout(n17863));
    jdff dff_B_E3WiGHgg3_2(.din(n17863), .dout(n17866));
    jdff dff_B_3odx0bRh1_2(.din(n17866), .dout(n17869));
    jdff dff_B_5xvwF1AJ0_2(.din(n17869), .dout(n17872));
    jdff dff_B_PXwsmNAp1_2(.din(n17872), .dout(n17875));
    jdff dff_B_EPR7Gnig5_2(.din(n17875), .dout(n17878));
    jdff dff_B_BdDlnazm5_2(.din(n17878), .dout(n17881));
    jdff dff_B_MNrxvM1N4_2(.din(n17881), .dout(n17884));
    jdff dff_B_FktG2pVH6_2(.din(n17884), .dout(n17887));
    jdff dff_B_QO1tV3ur3_2(.din(n17887), .dout(n17890));
    jdff dff_B_cHrW7Fv70_2(.din(n17890), .dout(n17893));
    jdff dff_B_WpCoG4pw2_2(.din(n17893), .dout(n17896));
    jdff dff_B_hRKP4OTP6_2(.din(n17896), .dout(n17899));
    jdff dff_B_aMKpDt5s2_2(.din(n17899), .dout(n17902));
    jdff dff_B_SBAQuFqy8_2(.din(n17902), .dout(n17905));
    jdff dff_B_KfWZey4c7_2(.din(n17905), .dout(n17908));
    jdff dff_B_1sSUDwjL5_2(.din(n17908), .dout(n17911));
    jdff dff_B_kRM71OWs1_2(.din(n17911), .dout(n17914));
    jdff dff_B_L7Re6p556_2(.din(n17914), .dout(n17917));
    jdff dff_B_RLZ1sl8P5_2(.din(n17917), .dout(n17920));
    jdff dff_B_j7Hhtgq99_2(.din(n17920), .dout(n17923));
    jdff dff_B_fS3wTcsS6_2(.din(n17923), .dout(n17926));
    jdff dff_B_SXqyNsLN2_2(.din(n1871), .dout(n17929));
    jdff dff_B_P8KsRJix4_1(.din(n1680), .dout(n17932));
    jdff dff_B_ivtSATeg6_2(.din(n1402), .dout(n17935));
    jdff dff_B_bSck8pg16_2(.din(n17935), .dout(n17938));
    jdff dff_B_PPlnoxLt1_2(.din(n17938), .dout(n17941));
    jdff dff_B_gVRRjAkj5_2(.din(n17941), .dout(n17944));
    jdff dff_B_yXvRq2zm9_2(.din(n17944), .dout(n17947));
    jdff dff_B_udWu3Xpw1_2(.din(n17947), .dout(n17950));
    jdff dff_B_HPD2iSFG7_2(.din(n17950), .dout(n17953));
    jdff dff_B_3wR3YO3U4_2(.din(n17953), .dout(n17956));
    jdff dff_B_tjZYPU2Z4_2(.din(n17956), .dout(n17959));
    jdff dff_B_WQXKZcJ65_2(.din(n17959), .dout(n17962));
    jdff dff_B_cbevVVP57_2(.din(n17962), .dout(n17965));
    jdff dff_B_q1NKHPOc8_2(.din(n17965), .dout(n17968));
    jdff dff_B_DAKdFrKw1_2(.din(n17968), .dout(n17971));
    jdff dff_B_kSqrz5ax3_2(.din(n17971), .dout(n17974));
    jdff dff_B_jT95uDpE4_2(.din(n17974), .dout(n17977));
    jdff dff_B_tWTx0CE57_2(.din(n17977), .dout(n17980));
    jdff dff_B_OTXhif4F3_2(.din(n17980), .dout(n17983));
    jdff dff_B_2CSl2zK59_2(.din(n17983), .dout(n17986));
    jdff dff_B_OMGyWvRk1_2(.din(n17986), .dout(n17989));
    jdff dff_B_oiv1Ej0a7_2(.din(n1570), .dout(n17992));
    jdff dff_B_dq2zZtCe8_1(.din(n1406), .dout(n17995));
    jdff dff_B_xM74ADJ29_2(.din(n1158), .dout(n17998));
    jdff dff_B_3eiP6WyV9_2(.din(n17998), .dout(n18001));
    jdff dff_B_wwcWKxWg0_2(.din(n18001), .dout(n18004));
    jdff dff_B_6JXvXZL78_2(.din(n18004), .dout(n18007));
    jdff dff_B_nhQwA36v6_2(.din(n18007), .dout(n18010));
    jdff dff_B_tKbfhqnV1_2(.din(n18010), .dout(n18013));
    jdff dff_B_u3mx4Fm42_2(.din(n18013), .dout(n18016));
    jdff dff_B_AHTXeoLm0_2(.din(n18016), .dout(n18019));
    jdff dff_B_AC2GPz4U2_2(.din(n18019), .dout(n18022));
    jdff dff_B_1m42DFdN0_2(.din(n18022), .dout(n18025));
    jdff dff_B_M8rU20jP3_2(.din(n18025), .dout(n18028));
    jdff dff_B_D2qZE4Ho3_2(.din(n18028), .dout(n18031));
    jdff dff_B_0hHmznac2_2(.din(n18031), .dout(n18034));
    jdff dff_B_qIOTDY6n4_2(.din(n18034), .dout(n18037));
    jdff dff_B_EBfLEmbc8_2(.din(n18037), .dout(n18040));
    jdff dff_B_VzlPzLz94_2(.din(n18040), .dout(n18043));
    jdff dff_B_eVcoFSmM5_2(.din(n1296), .dout(n18046));
    jdff dff_B_YZOkLI4o6_1(.din(n1162), .dout(n18049));
    jdff dff_B_xuWjU0ax0_2(.din(n938), .dout(n18052));
    jdff dff_B_udVe7QZu4_2(.din(n18052), .dout(n18055));
    jdff dff_B_Klc1olYN9_2(.din(n18055), .dout(n18058));
    jdff dff_B_7yt3SJo93_2(.din(n18058), .dout(n18061));
    jdff dff_B_X0RUb1Vg3_2(.din(n18061), .dout(n18064));
    jdff dff_B_khSBdDmA2_2(.din(n18064), .dout(n18067));
    jdff dff_B_gmVkOzqQ9_2(.din(n18067), .dout(n18070));
    jdff dff_B_PJFu1ViR8_2(.din(n18070), .dout(n18073));
    jdff dff_B_HwKhKumH7_2(.din(n18073), .dout(n18076));
    jdff dff_B_OVKJk7MB5_2(.din(n18076), .dout(n18079));
    jdff dff_B_kFgG7cQJ0_2(.din(n18079), .dout(n18082));
    jdff dff_B_CgvGs1og2_2(.din(n18082), .dout(n18085));
    jdff dff_B_ZT1o73KG3_2(.din(n18085), .dout(n18088));
    jdff dff_B_Pwl0RWjL6_2(.din(n1052), .dout(n18091));
    jdff dff_B_emUlAaqO8_1(.din(n942), .dout(n18094));
    jdff dff_B_VhQFQa4L7_2(.din(n745), .dout(n18097));
    jdff dff_B_mI8afoDC6_2(.din(n18097), .dout(n18100));
    jdff dff_B_lD2EsLUg4_2(.din(n18100), .dout(n18103));
    jdff dff_B_hAofEnzJ7_2(.din(n18103), .dout(n18106));
    jdff dff_B_2jUyhUpQ3_2(.din(n18106), .dout(n18109));
    jdff dff_B_mEOz2IDu0_2(.din(n18109), .dout(n18112));
    jdff dff_B_21cavMbj0_2(.din(n18112), .dout(n18115));
    jdff dff_B_tOik5Oue3_2(.din(n18115), .dout(n18118));
    jdff dff_B_lfRjL2Zh3_2(.din(n18118), .dout(n18121));
    jdff dff_B_Eevn5yIO0_2(.din(n18121), .dout(n18124));
    jdff dff_B_HK1uxouA2_2(.din(n832), .dout(n18127));
    jdff dff_B_CzRkLVTi9_1(.din(n749), .dout(n18130));
    jdff dff_B_7w8WipcE5_2(.din(n582), .dout(n18133));
    jdff dff_B_dyrzvjCK6_2(.din(n18133), .dout(n18136));
    jdff dff_B_c4k9w88Y8_2(.din(n18136), .dout(n18139));
    jdff dff_B_KUDyAe7b5_2(.din(n18139), .dout(n18142));
    jdff dff_B_edYnSJi39_2(.din(n18142), .dout(n18145));
    jdff dff_B_Z1h68yYY9_2(.din(n18145), .dout(n18148));
    jdff dff_B_1YazrMbv9_2(.din(n18148), .dout(n18151));
    jdff dff_B_eHQGTVDo8_2(.din(n639), .dout(n18154));
    jdff dff_B_7gwb7JRl2_1(.din(n585), .dout(n18157));
    jdff dff_B_CraBrRg64_0(.din(n476), .dout(n18160));
    jdff dff_B_BzYavjYu2_2(.din(n445), .dout(n18163));
    jdff dff_B_uynEtcs31_2(.din(n18163), .dout(n18166));
    jdff dff_B_VjiOsel71_2(.din(n18166), .dout(n18169));
    jdff dff_B_LYuZZ2cD3_2(.din(n18169), .dout(n18172));
    jdff dff_B_owZoKCNi7_1(.din(n453), .dout(n18175));
    jdff dff_A_HULXV26v8_0(.din(n18180), .dout(n18177));
    jdff dff_A_g6UKxOzF8_0(.din(n322), .dout(n18180));
    jdff dff_A_5rzIXust7_1(.din(n322), .dout(n18183));
    jdff dff_B_xI4KtHss7_1(.din(n4911), .dout(n18187));
    jdff dff_B_UZHohOxC7_2(.din(n4578), .dout(n18190));
    jdff dff_B_TPMAldQH1_2(.din(n18190), .dout(n18193));
    jdff dff_B_5umnd9nw4_2(.din(n18193), .dout(n18196));
    jdff dff_B_0BLSgGkg2_2(.din(n18196), .dout(n18199));
    jdff dff_B_OXUIaxMq9_2(.din(n18199), .dout(n18202));
    jdff dff_B_S9W9NEpu2_2(.din(n18202), .dout(n18205));
    jdff dff_B_5LMjWyT50_2(.din(n18205), .dout(n18208));
    jdff dff_B_UEMTtNBy1_2(.din(n18208), .dout(n18211));
    jdff dff_B_eD72nMjZ9_2(.din(n18211), .dout(n18214));
    jdff dff_B_oNjwemyX7_2(.din(n18214), .dout(n18217));
    jdff dff_B_Bd2jz3141_2(.din(n18217), .dout(n18220));
    jdff dff_B_h9VDgHHg6_2(.din(n18220), .dout(n18223));
    jdff dff_B_hunrCV1g8_2(.din(n18223), .dout(n18226));
    jdff dff_B_Oip8vEve4_2(.din(n18226), .dout(n18229));
    jdff dff_B_CGb7fR6C3_2(.din(n18229), .dout(n18232));
    jdff dff_B_lhU3fi1G5_2(.din(n18232), .dout(n18235));
    jdff dff_B_LMRqX8TV9_2(.din(n18235), .dout(n18238));
    jdff dff_B_gbUfhRb91_2(.din(n18238), .dout(n18241));
    jdff dff_B_gTW28RTb5_2(.din(n18241), .dout(n18244));
    jdff dff_B_JzFV2ONK0_2(.din(n18244), .dout(n18247));
    jdff dff_B_wZ2WsLoG4_2(.din(n18247), .dout(n18250));
    jdff dff_B_32evhavQ6_2(.din(n18250), .dout(n18253));
    jdff dff_B_zRNwHgyq7_2(.din(n18253), .dout(n18256));
    jdff dff_B_CSIE9nZD5_2(.din(n18256), .dout(n18259));
    jdff dff_B_Hw8v52VP5_2(.din(n18259), .dout(n18262));
    jdff dff_B_Z0XSY5sY1_2(.din(n18262), .dout(n18265));
    jdff dff_B_hr8K6DLV8_2(.din(n18265), .dout(n18268));
    jdff dff_B_CpslQAyj1_2(.din(n18268), .dout(n18271));
    jdff dff_B_RY8Tk1dv4_2(.din(n18271), .dout(n18274));
    jdff dff_B_GBUU6KTQ5_2(.din(n18274), .dout(n18277));
    jdff dff_B_DjKzZ8ih2_2(.din(n18277), .dout(n18280));
    jdff dff_B_Novj0s5f8_2(.din(n18280), .dout(n18283));
    jdff dff_B_xk6Kvhft1_2(.din(n18283), .dout(n18286));
    jdff dff_B_OAoSmCH78_2(.din(n18286), .dout(n18289));
    jdff dff_B_apBZy1Lr3_2(.din(n18289), .dout(n18292));
    jdff dff_B_6vvQA9U62_2(.din(n18292), .dout(n18295));
    jdff dff_B_MZft0Rpa3_2(.din(n18295), .dout(n18298));
    jdff dff_B_Mlm0szhn8_2(.din(n18298), .dout(n18301));
    jdff dff_B_WmvtQHks0_2(.din(n18301), .dout(n18304));
    jdff dff_B_Hyy1Rhgv9_2(.din(n18304), .dout(n18307));
    jdff dff_B_vRqrLQ890_2(.din(n18307), .dout(n18310));
    jdff dff_B_4nmjdSV93_2(.din(n18310), .dout(n18313));
    jdff dff_B_GfL5xMsK7_2(.din(n18313), .dout(n18316));
    jdff dff_B_ZCZqkJND0_2(.din(n18316), .dout(n18319));
    jdff dff_B_aULq1Jt46_2(.din(n18319), .dout(n18322));
    jdff dff_B_RhxBNb8P7_0(.din(n4907), .dout(n18325));
    jdff dff_A_LfO3RIHK7_1(.din(n4864), .dout(n18327));
    jdff dff_B_JQvbpp403_1(.din(n4582), .dout(n18331));
    jdff dff_B_U90uMvAa1_2(.din(n4232), .dout(n18334));
    jdff dff_B_NoiBQRiJ2_2(.din(n18334), .dout(n18337));
    jdff dff_B_tL1mZXxV9_2(.din(n18337), .dout(n18340));
    jdff dff_B_enHzjiiw8_2(.din(n18340), .dout(n18343));
    jdff dff_B_rZPNWW4h8_2(.din(n18343), .dout(n18346));
    jdff dff_B_5d4oZ88T3_2(.din(n18346), .dout(n18349));
    jdff dff_B_LF8NBnL16_2(.din(n18349), .dout(n18352));
    jdff dff_B_aZ6ugA3w1_2(.din(n18352), .dout(n18355));
    jdff dff_B_6tSuWOSC7_2(.din(n18355), .dout(n18358));
    jdff dff_B_7VPh3tWa7_2(.din(n18358), .dout(n18361));
    jdff dff_B_IYxYnHIB6_2(.din(n18361), .dout(n18364));
    jdff dff_B_ZfUC2LkC6_2(.din(n18364), .dout(n18367));
    jdff dff_B_bJUgQ1XH8_2(.din(n18367), .dout(n18370));
    jdff dff_B_1nfqEaHb5_2(.din(n18370), .dout(n18373));
    jdff dff_B_HHn9aFlQ1_2(.din(n18373), .dout(n18376));
    jdff dff_B_GGXcCVo58_2(.din(n18376), .dout(n18379));
    jdff dff_B_Uuexpj197_2(.din(n18379), .dout(n18382));
    jdff dff_B_qmZSuspL3_2(.din(n18382), .dout(n18385));
    jdff dff_B_ujEsUb5c8_2(.din(n18385), .dout(n18388));
    jdff dff_B_WaY0OldU3_2(.din(n18388), .dout(n18391));
    jdff dff_B_8gIcdXQJ8_2(.din(n18391), .dout(n18394));
    jdff dff_B_XAq5HCEW5_2(.din(n18394), .dout(n18397));
    jdff dff_B_b152A6lN0_2(.din(n18397), .dout(n18400));
    jdff dff_B_k5sYsebK4_2(.din(n18400), .dout(n18403));
    jdff dff_B_p5e0Aezl2_2(.din(n18403), .dout(n18406));
    jdff dff_B_mIXScm0Q0_2(.din(n18406), .dout(n18409));
    jdff dff_B_pkiogah55_2(.din(n18409), .dout(n18412));
    jdff dff_B_y6dWHmgG4_2(.din(n18412), .dout(n18415));
    jdff dff_B_m9hCgzYF4_2(.din(n18415), .dout(n18418));
    jdff dff_B_QPQHOcDJ8_2(.din(n18418), .dout(n18421));
    jdff dff_B_Dm8NMg9V0_2(.din(n18421), .dout(n18424));
    jdff dff_B_5NYVmpA13_2(.din(n18424), .dout(n18427));
    jdff dff_B_QteqSDU96_2(.din(n18427), .dout(n18430));
    jdff dff_B_t2oKy07e8_2(.din(n18430), .dout(n18433));
    jdff dff_B_2a6sqRoH9_2(.din(n18433), .dout(n18436));
    jdff dff_B_AFtX9sIe1_2(.din(n18436), .dout(n18439));
    jdff dff_B_mv30Dwhi6_2(.din(n18439), .dout(n18442));
    jdff dff_B_YQa0O84W7_2(.din(n18442), .dout(n18445));
    jdff dff_B_Ot77QrI62_2(.din(n18445), .dout(n18448));
    jdff dff_B_Iuv5wbIc7_2(.din(n18448), .dout(n18451));
    jdff dff_B_O1NHPjoB7_2(.din(n4514), .dout(n18454));
    jdff dff_B_lOSBJ7tE3_1(.din(n4236), .dout(n18457));
    jdff dff_B_9RJNcfrF2_2(.din(n3836), .dout(n18460));
    jdff dff_B_aEoizBxe3_2(.din(n18460), .dout(n18463));
    jdff dff_B_HUhjX3n13_2(.din(n18463), .dout(n18466));
    jdff dff_B_FAnE5Wis5_2(.din(n18466), .dout(n18469));
    jdff dff_B_inS0zxTF9_2(.din(n18469), .dout(n18472));
    jdff dff_B_ocxw3Y8Y4_2(.din(n18472), .dout(n18475));
    jdff dff_B_jKQ9Slxc5_2(.din(n18475), .dout(n18478));
    jdff dff_B_K6n4O5zN0_2(.din(n18478), .dout(n18481));
    jdff dff_B_qOSioDeL5_2(.din(n18481), .dout(n18484));
    jdff dff_B_sqONaICq0_2(.din(n18484), .dout(n18487));
    jdff dff_B_Sn6e1hcZ3_2(.din(n18487), .dout(n18490));
    jdff dff_B_SeW8fSQC5_2(.din(n18490), .dout(n18493));
    jdff dff_B_HBLe2pbK5_2(.din(n18493), .dout(n18496));
    jdff dff_B_LW4q84Ob7_2(.din(n18496), .dout(n18499));
    jdff dff_B_SZByWkeP9_2(.din(n18499), .dout(n18502));
    jdff dff_B_efFwplAt5_2(.din(n18502), .dout(n18505));
    jdff dff_B_b34dtNXc7_2(.din(n18505), .dout(n18508));
    jdff dff_B_hUPtkb717_2(.din(n18508), .dout(n18511));
    jdff dff_B_iagk97iy3_2(.din(n18511), .dout(n18514));
    jdff dff_B_eEyigFEQ2_2(.din(n18514), .dout(n18517));
    jdff dff_B_Y2XLB0bw4_2(.din(n18517), .dout(n18520));
    jdff dff_B_upcuLzjl5_2(.din(n18520), .dout(n18523));
    jdff dff_B_Es71zjQl3_2(.din(n18523), .dout(n18526));
    jdff dff_B_CDVgHeAy7_2(.din(n18526), .dout(n18529));
    jdff dff_B_duaNfMR90_2(.din(n18529), .dout(n18532));
    jdff dff_B_PK063A7o8_2(.din(n18532), .dout(n18535));
    jdff dff_B_cavtLJ0J7_2(.din(n18535), .dout(n18538));
    jdff dff_B_Ta4lBXkR2_2(.din(n18538), .dout(n18541));
    jdff dff_B_nys8lKOj7_2(.din(n18541), .dout(n18544));
    jdff dff_B_K8vOuI1A7_2(.din(n18544), .dout(n18547));
    jdff dff_B_kcgKCWXT9_2(.din(n18547), .dout(n18550));
    jdff dff_B_w3iLftcQ4_2(.din(n18550), .dout(n18553));
    jdff dff_B_wyRUFoPh9_2(.din(n18553), .dout(n18556));
    jdff dff_B_XNdGnwWX0_2(.din(n18556), .dout(n18559));
    jdff dff_B_skBhd1sh3_2(.din(n18559), .dout(n18562));
    jdff dff_B_3azMdPCw2_2(.din(n18562), .dout(n18565));
    jdff dff_B_SzYlsXIl7_2(.din(n18565), .dout(n18568));
    jdff dff_B_dQDJWevx9_2(.din(n4138), .dout(n18571));
    jdff dff_B_eCtGb53e0_1(.din(n3840), .dout(n18574));
    jdff dff_B_TJ0XPJ058_2(.din(n3459), .dout(n18577));
    jdff dff_B_LFISirk68_2(.din(n18577), .dout(n18580));
    jdff dff_B_jKk0oP377_2(.din(n18580), .dout(n18583));
    jdff dff_B_42TnxQTR1_2(.din(n18583), .dout(n18586));
    jdff dff_B_eBVbqtvU6_2(.din(n18586), .dout(n18589));
    jdff dff_B_fmejP46P8_2(.din(n18589), .dout(n18592));
    jdff dff_B_P5Q0hKUW1_2(.din(n18592), .dout(n18595));
    jdff dff_B_tFj8JxWy3_2(.din(n18595), .dout(n18598));
    jdff dff_B_8kmoOYdH1_2(.din(n18598), .dout(n18601));
    jdff dff_B_xpmmf9ZZ5_2(.din(n18601), .dout(n18604));
    jdff dff_B_vVzBuWer4_2(.din(n18604), .dout(n18607));
    jdff dff_B_ia0jNExX5_2(.din(n18607), .dout(n18610));
    jdff dff_B_OxSmDrYf1_2(.din(n18610), .dout(n18613));
    jdff dff_B_yjNFD4bk2_2(.din(n18613), .dout(n18616));
    jdff dff_B_iN8QNmSG1_2(.din(n18616), .dout(n18619));
    jdff dff_B_DuOCbTw32_2(.din(n18619), .dout(n18622));
    jdff dff_B_v2omJpgm9_2(.din(n18622), .dout(n18625));
    jdff dff_B_9sJXtV8b3_2(.din(n18625), .dout(n18628));
    jdff dff_B_HyIdw98L7_2(.din(n18628), .dout(n18631));
    jdff dff_B_EmupylG62_2(.din(n18631), .dout(n18634));
    jdff dff_B_QFbOzZc40_2(.din(n18634), .dout(n18637));
    jdff dff_B_ECWOHVdg0_2(.din(n18637), .dout(n18640));
    jdff dff_B_Rw1BSHKQ9_2(.din(n18640), .dout(n18643));
    jdff dff_B_O5WmV9b73_2(.din(n18643), .dout(n18646));
    jdff dff_B_GxUPNd4x8_2(.din(n18646), .dout(n18649));
    jdff dff_B_vtbgzxZ13_2(.din(n18649), .dout(n18652));
    jdff dff_B_zpW5bKD34_2(.din(n18652), .dout(n18655));
    jdff dff_B_IJr7b9Kn5_2(.din(n18655), .dout(n18658));
    jdff dff_B_jpvW04FO2_2(.din(n18658), .dout(n18661));
    jdff dff_B_zcdynVVv1_2(.din(n18661), .dout(n18664));
    jdff dff_B_SOxiC8ch5_2(.din(n18664), .dout(n18667));
    jdff dff_B_yfTvDbjC5_2(.din(n18667), .dout(n18670));
    jdff dff_B_r9psN4dq6_2(.din(n18670), .dout(n18673));
    jdff dff_B_vZdHmVoe7_2(.din(n18673), .dout(n18676));
    jdff dff_B_pV0mhRZL3_2(.din(n3735), .dout(n18679));
    jdff dff_B_Rb5srVo57_1(.din(n3463), .dout(n18682));
    jdff dff_B_lZn9UF0Q4_2(.din(n3058), .dout(n18685));
    jdff dff_B_15z3pBvV7_2(.din(n18685), .dout(n18688));
    jdff dff_B_v8TT3key1_2(.din(n18688), .dout(n18691));
    jdff dff_B_3WxeF3as2_2(.din(n18691), .dout(n18694));
    jdff dff_B_cW4lRg5Y5_2(.din(n18694), .dout(n18697));
    jdff dff_B_on5C6lik6_2(.din(n18697), .dout(n18700));
    jdff dff_B_poWIt2H63_2(.din(n18700), .dout(n18703));
    jdff dff_B_keKaoNRj2_2(.din(n18703), .dout(n18706));
    jdff dff_B_YPAGzvB34_2(.din(n18706), .dout(n18709));
    jdff dff_B_sKfDDsa15_2(.din(n18709), .dout(n18712));
    jdff dff_B_145WmUMG5_2(.din(n18712), .dout(n18715));
    jdff dff_B_IDhYC0Mq0_2(.din(n18715), .dout(n18718));
    jdff dff_B_ltG2fnaH3_2(.din(n18718), .dout(n18721));
    jdff dff_B_fcwqtJuG0_2(.din(n18721), .dout(n18724));
    jdff dff_B_3iixEj0N7_2(.din(n18724), .dout(n18727));
    jdff dff_B_WrM8pzZb8_2(.din(n18727), .dout(n18730));
    jdff dff_B_4tTfQJlb0_2(.din(n18730), .dout(n18733));
    jdff dff_B_olsGP0uP6_2(.din(n18733), .dout(n18736));
    jdff dff_B_HoZJEgBU2_2(.din(n18736), .dout(n18739));
    jdff dff_B_26PZ9btN9_2(.din(n18739), .dout(n18742));
    jdff dff_B_wn9pbkMV8_2(.din(n18742), .dout(n18745));
    jdff dff_B_IKMYJJjS8_2(.din(n18745), .dout(n18748));
    jdff dff_B_0d4yX2xg0_2(.din(n18748), .dout(n18751));
    jdff dff_B_3XdOFMFu8_2(.din(n18751), .dout(n18754));
    jdff dff_B_WPiWKbN28_2(.din(n18754), .dout(n18757));
    jdff dff_B_3L6vqFYl4_2(.din(n18757), .dout(n18760));
    jdff dff_B_OtpxpA1G4_2(.din(n18760), .dout(n18763));
    jdff dff_B_5o0b8ZpA8_2(.din(n18763), .dout(n18766));
    jdff dff_B_pyChaReD3_2(.din(n18766), .dout(n18769));
    jdff dff_B_djIcuisx9_2(.din(n18769), .dout(n18772));
    jdff dff_B_E2Lm7Htj4_2(.din(n18772), .dout(n18775));
    jdff dff_B_eZBfBava6_2(.din(n3333), .dout(n18778));
    jdff dff_B_fWUgkO5b0_1(.din(n3062), .dout(n18781));
    jdff dff_B_6iUBDZHj4_2(.din(n2679), .dout(n18784));
    jdff dff_B_Fd0MyKka5_2(.din(n18784), .dout(n18787));
    jdff dff_B_ND8OBbwC0_2(.din(n18787), .dout(n18790));
    jdff dff_B_nErpmHl18_2(.din(n18790), .dout(n18793));
    jdff dff_B_2tEclMAK1_2(.din(n18793), .dout(n18796));
    jdff dff_B_lA9v8wsM5_2(.din(n18796), .dout(n18799));
    jdff dff_B_KnaG4l6K5_2(.din(n18799), .dout(n18802));
    jdff dff_B_m0I4GfXp4_2(.din(n18802), .dout(n18805));
    jdff dff_B_dwd3x7Ia6_2(.din(n18805), .dout(n18808));
    jdff dff_B_klRcr3bk7_2(.din(n18808), .dout(n18811));
    jdff dff_B_rl1m2nHq1_2(.din(n18811), .dout(n18814));
    jdff dff_B_gO1gN7Ik5_2(.din(n18814), .dout(n18817));
    jdff dff_B_GHym1I754_2(.din(n18817), .dout(n18820));
    jdff dff_B_jl9Ge0LM5_2(.din(n18820), .dout(n18823));
    jdff dff_B_x0QUaPVo7_2(.din(n18823), .dout(n18826));
    jdff dff_B_4qNuKCMZ4_2(.din(n18826), .dout(n18829));
    jdff dff_B_wWjawONr7_2(.din(n18829), .dout(n18832));
    jdff dff_B_YrfYcJyl0_2(.din(n18832), .dout(n18835));
    jdff dff_B_ALQWyxbg3_2(.din(n18835), .dout(n18838));
    jdff dff_B_VxcZ4zR37_2(.din(n18838), .dout(n18841));
    jdff dff_B_3SSxB3xy1_2(.din(n18841), .dout(n18844));
    jdff dff_B_r00RNczI8_2(.din(n18844), .dout(n18847));
    jdff dff_B_6TmPeOpD3_2(.din(n18847), .dout(n18850));
    jdff dff_B_QQGQvHcR2_2(.din(n18850), .dout(n18853));
    jdff dff_B_uwyEBFDM8_2(.din(n18853), .dout(n18856));
    jdff dff_B_PWGYKLKY5_2(.din(n18856), .dout(n18859));
    jdff dff_B_e6K5chWS2_2(.din(n18859), .dout(n18862));
    jdff dff_B_fj8Vgs8k0_2(.din(n18862), .dout(n18865));
    jdff dff_B_c0w64E9o7_2(.din(n2928), .dout(n18868));
    jdff dff_B_mxcrFEy75_1(.din(n2683), .dout(n18871));
    jdff dff_B_4OMtVokv1_2(.din(n2324), .dout(n18874));
    jdff dff_B_acoRmwt28_2(.din(n18874), .dout(n18877));
    jdff dff_B_9KkUNVVI6_2(.din(n18877), .dout(n18880));
    jdff dff_B_G1Bo0LPI7_2(.din(n18880), .dout(n18883));
    jdff dff_B_JICtEKpQ8_2(.din(n18883), .dout(n18886));
    jdff dff_B_pEUGoxrz8_2(.din(n18886), .dout(n18889));
    jdff dff_B_N306hy2O3_2(.din(n18889), .dout(n18892));
    jdff dff_B_lceEbzHj3_2(.din(n18892), .dout(n18895));
    jdff dff_B_gFD0s3mq0_2(.din(n18895), .dout(n18898));
    jdff dff_B_2lffssTC4_2(.din(n18898), .dout(n18901));
    jdff dff_B_Yxr7O1Uj6_2(.din(n18901), .dout(n18904));
    jdff dff_B_5YMx5so30_2(.din(n18904), .dout(n18907));
    jdff dff_B_oexpnFcj0_2(.din(n18907), .dout(n18910));
    jdff dff_B_AQJqsCTT4_2(.din(n18910), .dout(n18913));
    jdff dff_B_4psAA1UQ1_2(.din(n18913), .dout(n18916));
    jdff dff_B_0eo6v2GS3_2(.din(n18916), .dout(n18919));
    jdff dff_B_297USJ0g9_2(.din(n18919), .dout(n18922));
    jdff dff_B_mAYcP06y0_2(.din(n18922), .dout(n18925));
    jdff dff_B_NGHXSi535_2(.din(n18925), .dout(n18928));
    jdff dff_B_lU1WgcM25_2(.din(n18928), .dout(n18931));
    jdff dff_B_phJ4JOgn2_2(.din(n18931), .dout(n18934));
    jdff dff_B_6Lz8YEo09_2(.din(n18934), .dout(n18937));
    jdff dff_B_q7GzRp9T7_2(.din(n18937), .dout(n18940));
    jdff dff_B_43Y1xxIr5_2(.din(n18940), .dout(n18943));
    jdff dff_B_UDGVpLg17_2(.din(n18943), .dout(n18946));
    jdff dff_B_ycB40T2b3_2(.din(n2546), .dout(n18949));
    jdff dff_B_ygjs60Th7_1(.din(n2328), .dout(n18952));
    jdff dff_B_Z0Duo9dV0_2(.din(n1996), .dout(n18955));
    jdff dff_B_VRnX6mHH9_2(.din(n18955), .dout(n18958));
    jdff dff_B_hXfiWR3P6_2(.din(n18958), .dout(n18961));
    jdff dff_B_3jIfXF6T0_2(.din(n18961), .dout(n18964));
    jdff dff_B_vdyx2JQE5_2(.din(n18964), .dout(n18967));
    jdff dff_B_lOPKwDuT8_2(.din(n18967), .dout(n18970));
    jdff dff_B_l3MrveyU8_2(.din(n18970), .dout(n18973));
    jdff dff_B_4NWA4bwp0_2(.din(n18973), .dout(n18976));
    jdff dff_B_eOjGzMjl3_2(.din(n18976), .dout(n18979));
    jdff dff_B_x5te0b223_2(.din(n18979), .dout(n18982));
    jdff dff_B_ynbAoZOU9_2(.din(n18982), .dout(n18985));
    jdff dff_B_oaA6cAh42_2(.din(n18985), .dout(n18988));
    jdff dff_B_yBxAq33v3_2(.din(n18988), .dout(n18991));
    jdff dff_B_5faZdRXQ3_2(.din(n18991), .dout(n18994));
    jdff dff_B_DyBzSxvy7_2(.din(n18994), .dout(n18997));
    jdff dff_B_b2UQyiTc7_2(.din(n18997), .dout(n19000));
    jdff dff_B_EjFXhMjI9_2(.din(n19000), .dout(n19003));
    jdff dff_B_O4ZLzo7Q7_2(.din(n19003), .dout(n19006));
    jdff dff_B_OEPcdrkb7_2(.din(n19006), .dout(n19009));
    jdff dff_B_arWQVsp99_2(.din(n19009), .dout(n19012));
    jdff dff_B_xctT5K701_2(.din(n19012), .dout(n19015));
    jdff dff_B_DGBVxjsn9_2(.din(n19015), .dout(n19018));
    jdff dff_B_vZ6KDoV16_2(.din(n2191), .dout(n19021));
    jdff dff_B_WMEeveX70_1(.din(n2000), .dout(n19024));
    jdff dff_B_8xYkexNR0_2(.din(n1695), .dout(n19027));
    jdff dff_B_XchKCJZz6_2(.din(n19027), .dout(n19030));
    jdff dff_B_BcqWLi289_2(.din(n19030), .dout(n19033));
    jdff dff_B_7Ixca6yZ6_2(.din(n19033), .dout(n19036));
    jdff dff_B_GfjppUmw8_2(.din(n19036), .dout(n19039));
    jdff dff_B_TL87T78e5_2(.din(n19039), .dout(n19042));
    jdff dff_B_c6ACRB5u9_2(.din(n19042), .dout(n19045));
    jdff dff_B_7NIqPGV22_2(.din(n19045), .dout(n19048));
    jdff dff_B_648NKTum2_2(.din(n19048), .dout(n19051));
    jdff dff_B_uf0MxER77_2(.din(n19051), .dout(n19054));
    jdff dff_B_zrLxTw9F9_2(.din(n19054), .dout(n19057));
    jdff dff_B_8H5kqOg08_2(.din(n19057), .dout(n19060));
    jdff dff_B_lCivCT015_2(.din(n19060), .dout(n19063));
    jdff dff_B_qMyG07dM2_2(.din(n19063), .dout(n19066));
    jdff dff_B_TGb8nIso0_2(.din(n19066), .dout(n19069));
    jdff dff_B_HDWsRIIj2_2(.din(n19069), .dout(n19072));
    jdff dff_B_DsXCdJIH8_2(.din(n19072), .dout(n19075));
    jdff dff_B_sKSNMA531_2(.din(n19075), .dout(n19078));
    jdff dff_B_A3MxRWOn7_2(.din(n19078), .dout(n19081));
    jdff dff_B_DFyyoA0N0_2(.din(n1863), .dout(n19084));
    jdff dff_B_VvhQZ0NB6_1(.din(n1699), .dout(n19087));
    jdff dff_B_pgbrNAnr1_2(.din(n1421), .dout(n19090));
    jdff dff_B_bEdYUBvI7_2(.din(n19090), .dout(n19093));
    jdff dff_B_zugL85Ye3_2(.din(n19093), .dout(n19096));
    jdff dff_B_i48PGo582_2(.din(n19096), .dout(n19099));
    jdff dff_B_te4HLu1p9_2(.din(n19099), .dout(n19102));
    jdff dff_B_hwMFpPo93_2(.din(n19102), .dout(n19105));
    jdff dff_B_A60vuWWt2_2(.din(n19105), .dout(n19108));
    jdff dff_B_EQBRvvYW5_2(.din(n19108), .dout(n19111));
    jdff dff_B_QIrZ9R2b6_2(.din(n19111), .dout(n19114));
    jdff dff_B_aDMKBFu62_2(.din(n19114), .dout(n19117));
    jdff dff_B_HTRPVf4C5_2(.din(n19117), .dout(n19120));
    jdff dff_B_ziCjGJz67_2(.din(n19120), .dout(n19123));
    jdff dff_B_eIRFFKhB0_2(.din(n19123), .dout(n19126));
    jdff dff_B_txtJm3rF6_2(.din(n19126), .dout(n19129));
    jdff dff_B_k4XIAjuc1_2(.din(n19129), .dout(n19132));
    jdff dff_B_RNkWNosq9_2(.din(n19132), .dout(n19135));
    jdff dff_B_J6QBkd1c4_2(.din(n1562), .dout(n19138));
    jdff dff_B_UaNQnCtd9_1(.din(n1425), .dout(n19141));
    jdff dff_B_dighet794_2(.din(n1177), .dout(n19144));
    jdff dff_B_XMXdOW4Z5_2(.din(n19144), .dout(n19147));
    jdff dff_B_vKmnixM04_2(.din(n19147), .dout(n19150));
    jdff dff_B_MoWautym2_2(.din(n19150), .dout(n19153));
    jdff dff_B_758aSQuj9_2(.din(n19153), .dout(n19156));
    jdff dff_B_dFY0FqmX0_2(.din(n19156), .dout(n19159));
    jdff dff_B_ht9z6Nlz5_2(.din(n19159), .dout(n19162));
    jdff dff_B_6LLvWaqw6_2(.din(n19162), .dout(n19165));
    jdff dff_B_neqTqmG74_2(.din(n19165), .dout(n19168));
    jdff dff_B_NsYz8Tbc1_2(.din(n19168), .dout(n19171));
    jdff dff_B_0bhSfjpg3_2(.din(n19171), .dout(n19174));
    jdff dff_B_WSbE96bQ3_2(.din(n19174), .dout(n19177));
    jdff dff_B_TCa8Nxe60_2(.din(n19177), .dout(n19180));
    jdff dff_B_nnVOysn11_2(.din(n1288), .dout(n19183));
    jdff dff_B_ztAH3VDi4_1(.din(n1181), .dout(n19186));
    jdff dff_B_mwJc1BeS3_2(.din(n957), .dout(n19189));
    jdff dff_B_3sxCiYtf9_2(.din(n19189), .dout(n19192));
    jdff dff_B_RLpQhle37_2(.din(n19192), .dout(n19195));
    jdff dff_B_b01OVPTv4_2(.din(n19195), .dout(n19198));
    jdff dff_B_YVIsgybR5_2(.din(n19198), .dout(n19201));
    jdff dff_B_B7qquJtX8_2(.din(n19201), .dout(n19204));
    jdff dff_B_Ea8Tq7lI1_2(.din(n19204), .dout(n19207));
    jdff dff_B_qcWevvG74_2(.din(n19207), .dout(n19210));
    jdff dff_B_5s5oyIZD3_2(.din(n19210), .dout(n19213));
    jdff dff_B_BMfrFhAf7_2(.din(n19213), .dout(n19216));
    jdff dff_B_cFedhM6m6_2(.din(n1044), .dout(n19219));
    jdff dff_B_lIUTpAE80_1(.din(n961), .dout(n19222));
    jdff dff_B_uL5pjgHx5_2(.din(n764), .dout(n19225));
    jdff dff_B_tHoIgdej0_2(.din(n19225), .dout(n19228));
    jdff dff_B_VQfOBjtP3_2(.din(n19228), .dout(n19231));
    jdff dff_B_xiJINwsA5_2(.din(n19231), .dout(n19234));
    jdff dff_B_3ZyEqvnH6_2(.din(n19234), .dout(n19237));
    jdff dff_B_BG0lSzJ73_2(.din(n19237), .dout(n19240));
    jdff dff_B_9cmf9K3G9_2(.din(n19240), .dout(n19243));
    jdff dff_B_nalj3afZ5_2(.din(n824), .dout(n19246));
    jdff dff_B_BmR3h8NF0_1(.din(n767), .dout(n19249));
    jdff dff_B_fEsB0Ljq9_0(.din(n631), .dout(n19252));
    jdff dff_B_Su4WFigI8_2(.din(n600), .dout(n19255));
    jdff dff_B_jnLnM26k1_2(.din(n19255), .dout(n19258));
    jdff dff_B_nHW52yND5_2(.din(n19258), .dout(n19261));
    jdff dff_B_psp5KmyI1_2(.din(n19261), .dout(n19264));
    jdff dff_B_74u3CizV5_1(.din(n608), .dout(n19267));
    jdff dff_A_lY35Gf6q5_0(.din(n616), .dout(n19269));
    jdff dff_A_4KBjmpb35_0(.din(n19275), .dout(n19272));
    jdff dff_A_g6U8xrxE7_0(.din(n461), .dout(n19275));
    jdff dff_A_IX8YLItY8_1(.din(n461), .dout(n19278));
    jdff dff_B_5P4pp9zh5_2(.din(n5237), .dout(n19282));
    jdff dff_B_2YkkQ9rd3_1(.din(n5229), .dout(n19285));
    jdff dff_B_JuqYWJY15_2(.din(n4923), .dout(n19288));
    jdff dff_B_MFOTu59Z4_2(.din(n19288), .dout(n19291));
    jdff dff_B_pUrciEDZ6_2(.din(n19291), .dout(n19294));
    jdff dff_B_ae0rn1Vl9_2(.din(n19294), .dout(n19297));
    jdff dff_B_QQMrrVrk5_2(.din(n19297), .dout(n19300));
    jdff dff_B_4kSfgJ1w5_2(.din(n19300), .dout(n19303));
    jdff dff_B_lm8Xe7PB3_2(.din(n19303), .dout(n19306));
    jdff dff_B_oohCaw863_2(.din(n19306), .dout(n19309));
    jdff dff_B_ZKqaoZ7F4_2(.din(n19309), .dout(n19312));
    jdff dff_B_9n80JxzK0_2(.din(n19312), .dout(n19315));
    jdff dff_B_9GOdYVMe1_2(.din(n19315), .dout(n19318));
    jdff dff_B_W0HuBbm93_2(.din(n19318), .dout(n19321));
    jdff dff_B_2WXWACs30_2(.din(n19321), .dout(n19324));
    jdff dff_B_ItzjVcsw5_2(.din(n19324), .dout(n19327));
    jdff dff_B_jSscDheQ5_2(.din(n19327), .dout(n19330));
    jdff dff_B_IFADsWC58_2(.din(n19330), .dout(n19333));
    jdff dff_B_X2amMj6X1_2(.din(n19333), .dout(n19336));
    jdff dff_B_hz0cZMFW7_2(.din(n19336), .dout(n19339));
    jdff dff_B_R3E6d6yl4_2(.din(n19339), .dout(n19342));
    jdff dff_B_Jtl4fyGM1_2(.din(n19342), .dout(n19345));
    jdff dff_B_0iPHElpd8_2(.din(n19345), .dout(n19348));
    jdff dff_B_sCXxBtso0_2(.din(n19348), .dout(n19351));
    jdff dff_B_hgajkR5L3_2(.din(n19351), .dout(n19354));
    jdff dff_B_MflVSr1N3_2(.din(n19354), .dout(n19357));
    jdff dff_B_uFbs19s49_2(.din(n19357), .dout(n19360));
    jdff dff_B_JdRzqbq86_2(.din(n19360), .dout(n19363));
    jdff dff_B_uEbBayz01_2(.din(n19363), .dout(n19366));
    jdff dff_B_966hOrhk2_2(.din(n19366), .dout(n19369));
    jdff dff_B_TG4B0ySn7_2(.din(n19369), .dout(n19372));
    jdff dff_B_vUJgjzdo4_2(.din(n19372), .dout(n19375));
    jdff dff_B_1Zqukoio1_2(.din(n19375), .dout(n19378));
    jdff dff_B_QgioRiTJ3_2(.din(n19378), .dout(n19381));
    jdff dff_B_m8IPSO2E5_2(.din(n19381), .dout(n19384));
    jdff dff_B_z0uyovCq3_2(.din(n19384), .dout(n19387));
    jdff dff_B_6P9Ru5e75_2(.din(n19387), .dout(n19390));
    jdff dff_B_Mf8FdXk30_2(.din(n19390), .dout(n19393));
    jdff dff_B_2vxJTD2u6_2(.din(n19393), .dout(n19396));
    jdff dff_B_zKVWfg8V0_2(.din(n19396), .dout(n19399));
    jdff dff_B_tzpUw0ad2_2(.din(n19399), .dout(n19402));
    jdff dff_B_SicE7c7A6_2(.din(n19402), .dout(n19405));
    jdff dff_B_uumtACLN2_2(.din(n19405), .dout(n19408));
    jdff dff_B_FZ6IXBKU5_2(.din(n19408), .dout(n19411));
    jdff dff_B_cSvpNLU87_2(.din(n19411), .dout(n19414));
    jdff dff_B_GjTXKUHD5_2(.din(n19414), .dout(n19417));
    jdff dff_B_mJ9wVZH48_2(.din(n19417), .dout(n19420));
    jdff dff_B_Y7cEae5U1_1(.din(n4927), .dout(n19423));
    jdff dff_B_R0URrd2P3_2(.din(n4597), .dout(n19426));
    jdff dff_B_hwqMBUsx1_2(.din(n19426), .dout(n19429));
    jdff dff_B_YErTvJtL1_2(.din(n19429), .dout(n19432));
    jdff dff_B_zut8PZZn6_2(.din(n19432), .dout(n19435));
    jdff dff_B_UbOtM6RN0_2(.din(n19435), .dout(n19438));
    jdff dff_B_wieL0KOK9_2(.din(n19438), .dout(n19441));
    jdff dff_B_pej1ijAG6_2(.din(n19441), .dout(n19444));
    jdff dff_B_8IfK4BbJ0_2(.din(n19444), .dout(n19447));
    jdff dff_B_wzqxTmUW5_2(.din(n19447), .dout(n19450));
    jdff dff_B_3zUfbgfe6_2(.din(n19450), .dout(n19453));
    jdff dff_B_9u2PPMPm8_2(.din(n19453), .dout(n19456));
    jdff dff_B_somNHLV52_2(.din(n19456), .dout(n19459));
    jdff dff_B_wL41hHxW5_2(.din(n19459), .dout(n19462));
    jdff dff_B_j9GT010h3_2(.din(n19462), .dout(n19465));
    jdff dff_B_cX1W1JIx9_2(.din(n19465), .dout(n19468));
    jdff dff_B_8jhoHevL2_2(.din(n19468), .dout(n19471));
    jdff dff_B_uC7tnTzC1_2(.din(n19471), .dout(n19474));
    jdff dff_B_EbtojuWS9_2(.din(n19474), .dout(n19477));
    jdff dff_B_ev9XnmBM8_2(.din(n19477), .dout(n19480));
    jdff dff_B_wOC6kAbp3_2(.din(n19480), .dout(n19483));
    jdff dff_B_rgSopqSd3_2(.din(n19483), .dout(n19486));
    jdff dff_B_4LkbpIWS1_2(.din(n19486), .dout(n19489));
    jdff dff_B_Cd3jsIgJ2_2(.din(n19489), .dout(n19492));
    jdff dff_B_Jzi6yvEP6_2(.din(n19492), .dout(n19495));
    jdff dff_B_fF6d4owR2_2(.din(n19495), .dout(n19498));
    jdff dff_B_CBEP8Hgy4_2(.din(n19498), .dout(n19501));
    jdff dff_B_eEsFpIIl4_2(.din(n19501), .dout(n19504));
    jdff dff_B_b2m5Bg1A5_2(.din(n19504), .dout(n19507));
    jdff dff_B_h6bXhJra1_2(.din(n19507), .dout(n19510));
    jdff dff_B_PAMu7WGB0_2(.din(n19510), .dout(n19513));
    jdff dff_B_2Bnc9tCI2_2(.din(n19513), .dout(n19516));
    jdff dff_B_NyIK2i0x2_2(.din(n19516), .dout(n19519));
    jdff dff_B_KJkA6zte2_2(.din(n19519), .dout(n19522));
    jdff dff_B_DCwdtyls8_2(.din(n19522), .dout(n19525));
    jdff dff_B_nYNWCZCP3_2(.din(n19525), .dout(n19528));
    jdff dff_B_3jzPG3fB9_2(.din(n19528), .dout(n19531));
    jdff dff_B_fzmUEzNP9_2(.din(n19531), .dout(n19534));
    jdff dff_B_Krivrsg29_2(.din(n19534), .dout(n19537));
    jdff dff_B_MIEuH8hx6_2(.din(n19537), .dout(n19540));
    jdff dff_B_zS3qZF2g9_2(.din(n19540), .dout(n19543));
    jdff dff_B_veZHBUJv1_1(.din(n4601), .dout(n19546));
    jdff dff_B_lLeaJOqU6_2(.din(n4251), .dout(n19549));
    jdff dff_B_Gpc8TddJ5_2(.din(n19549), .dout(n19552));
    jdff dff_B_3dtFcCsZ5_2(.din(n19552), .dout(n19555));
    jdff dff_B_NgCwOr0u0_2(.din(n19555), .dout(n19558));
    jdff dff_B_4oDTmw7D5_2(.din(n19558), .dout(n19561));
    jdff dff_B_HJtdDzz43_2(.din(n19561), .dout(n19564));
    jdff dff_B_VEuFlud65_2(.din(n19564), .dout(n19567));
    jdff dff_B_JW6v6wyL5_2(.din(n19567), .dout(n19570));
    jdff dff_B_r83ELxry2_2(.din(n19570), .dout(n19573));
    jdff dff_B_LOIXOIv78_2(.din(n19573), .dout(n19576));
    jdff dff_B_F6yoJNjV6_2(.din(n19576), .dout(n19579));
    jdff dff_B_zLLd9rv06_2(.din(n19579), .dout(n19582));
    jdff dff_B_2BhHRQih1_2(.din(n19582), .dout(n19585));
    jdff dff_B_JB3k6geG3_2(.din(n19585), .dout(n19588));
    jdff dff_B_5q3NxEkH7_2(.din(n19588), .dout(n19591));
    jdff dff_B_eSBQStM02_2(.din(n19591), .dout(n19594));
    jdff dff_B_Y8TEAzYS5_2(.din(n19594), .dout(n19597));
    jdff dff_B_p9w5r6di2_2(.din(n19597), .dout(n19600));
    jdff dff_B_o7hHWP8Z2_2(.din(n19600), .dout(n19603));
    jdff dff_B_Nn3vFM4n8_2(.din(n19603), .dout(n19606));
    jdff dff_B_tSw5WrnD2_2(.din(n19606), .dout(n19609));
    jdff dff_B_61w3WLDm2_2(.din(n19609), .dout(n19612));
    jdff dff_B_P17ohZkU7_2(.din(n19612), .dout(n19615));
    jdff dff_B_RjHV7ITZ0_2(.din(n19615), .dout(n19618));
    jdff dff_B_9Tz4lley7_2(.din(n19618), .dout(n19621));
    jdff dff_B_QkGmoXMf7_2(.din(n19621), .dout(n19624));
    jdff dff_B_6sVUDqCe5_2(.din(n19624), .dout(n19627));
    jdff dff_B_VwWx60VY1_2(.din(n19627), .dout(n19630));
    jdff dff_B_czw2cOJi9_2(.din(n19630), .dout(n19633));
    jdff dff_B_NZD7xLZ20_2(.din(n19633), .dout(n19636));
    jdff dff_B_bXjCGVl78_2(.din(n19636), .dout(n19639));
    jdff dff_B_ViKNaZDL6_2(.din(n19639), .dout(n19642));
    jdff dff_B_xm6oSMuN9_2(.din(n19642), .dout(n19645));
    jdff dff_B_w1Q7IhUT5_2(.din(n19645), .dout(n19648));
    jdff dff_B_g0wfKieS7_2(.din(n19648), .dout(n19651));
    jdff dff_B_yb8ttNkF6_2(.din(n19651), .dout(n19654));
    jdff dff_B_WFUfie7T9_2(.din(n19654), .dout(n19657));
    jdff dff_B_uOEOZObL3_1(.din(n4255), .dout(n19660));
    jdff dff_B_1ojTqbuu5_2(.din(n3855), .dout(n19663));
    jdff dff_B_Mu1h62B41_2(.din(n19663), .dout(n19666));
    jdff dff_B_h48RORwK8_2(.din(n19666), .dout(n19669));
    jdff dff_B_M8KCaOh65_2(.din(n19669), .dout(n19672));
    jdff dff_B_id2XqKqF6_2(.din(n19672), .dout(n19675));
    jdff dff_B_477vbMIP6_2(.din(n19675), .dout(n19678));
    jdff dff_B_YARh4HJy9_2(.din(n19678), .dout(n19681));
    jdff dff_B_iaZlrNcx3_2(.din(n19681), .dout(n19684));
    jdff dff_B_cXwSHk198_2(.din(n19684), .dout(n19687));
    jdff dff_B_RUWyyqcD6_2(.din(n19687), .dout(n19690));
    jdff dff_B_Z0uOcxay9_2(.din(n19690), .dout(n19693));
    jdff dff_B_iYnFwR0M6_2(.din(n19693), .dout(n19696));
    jdff dff_B_kyLjDg9w9_2(.din(n19696), .dout(n19699));
    jdff dff_B_pVeZ9JKP0_2(.din(n19699), .dout(n19702));
    jdff dff_B_LMlpdPGc4_2(.din(n19702), .dout(n19705));
    jdff dff_B_0pEm2brJ7_2(.din(n19705), .dout(n19708));
    jdff dff_B_caSTd6PM9_2(.din(n19708), .dout(n19711));
    jdff dff_B_PePFdTAP5_2(.din(n19711), .dout(n19714));
    jdff dff_B_jsD4HgHt8_2(.din(n19714), .dout(n19717));
    jdff dff_B_Sg1wUg0H2_2(.din(n19717), .dout(n19720));
    jdff dff_B_yF28aubg9_2(.din(n19720), .dout(n19723));
    jdff dff_B_tvAuubX99_2(.din(n19723), .dout(n19726));
    jdff dff_B_4BqsZZHS4_2(.din(n19726), .dout(n19729));
    jdff dff_B_A81Y95J23_2(.din(n19729), .dout(n19732));
    jdff dff_B_kPfcUBLB3_2(.din(n19732), .dout(n19735));
    jdff dff_B_g2enGmPe7_2(.din(n19735), .dout(n19738));
    jdff dff_B_fZHCOcL76_2(.din(n19738), .dout(n19741));
    jdff dff_B_53SXnkVu4_2(.din(n19741), .dout(n19744));
    jdff dff_B_kCbt8Nyg5_2(.din(n19744), .dout(n19747));
    jdff dff_B_fJoq84PA2_2(.din(n19747), .dout(n19750));
    jdff dff_B_cRtX1KIi2_2(.din(n19750), .dout(n19753));
    jdff dff_B_TMcWbaYf7_2(.din(n19753), .dout(n19756));
    jdff dff_B_GOyUKeLb9_2(.din(n19756), .dout(n19759));
    jdff dff_B_4P83CbSp6_2(.din(n19759), .dout(n19762));
    jdff dff_B_UhIogdie1_1(.din(n3859), .dout(n19765));
    jdff dff_B_ar28uOhU3_2(.din(n3478), .dout(n19768));
    jdff dff_B_Mbxc45If8_2(.din(n19768), .dout(n19771));
    jdff dff_B_IRIz1hRJ5_2(.din(n19771), .dout(n19774));
    jdff dff_B_sAwZzgXI3_2(.din(n19774), .dout(n19777));
    jdff dff_B_Su7aprlm6_2(.din(n19777), .dout(n19780));
    jdff dff_B_0uBCu5Mm2_2(.din(n19780), .dout(n19783));
    jdff dff_B_zevdaLSW5_2(.din(n19783), .dout(n19786));
    jdff dff_B_Q7unzoo97_2(.din(n19786), .dout(n19789));
    jdff dff_B_mjsYeI5S9_2(.din(n19789), .dout(n19792));
    jdff dff_B_3un0WgMB5_2(.din(n19792), .dout(n19795));
    jdff dff_B_J0Da3LgN1_2(.din(n19795), .dout(n19798));
    jdff dff_B_u054pjDB7_2(.din(n19798), .dout(n19801));
    jdff dff_B_k3aJothM2_2(.din(n19801), .dout(n19804));
    jdff dff_B_C2ncuhDq0_2(.din(n19804), .dout(n19807));
    jdff dff_B_U3SgzjHC2_2(.din(n19807), .dout(n19810));
    jdff dff_B_Fuqn5Uxb5_2(.din(n19810), .dout(n19813));
    jdff dff_B_4jyMa10R5_2(.din(n19813), .dout(n19816));
    jdff dff_B_coKJHB6e8_2(.din(n19816), .dout(n19819));
    jdff dff_B_rmaE43Yd5_2(.din(n19819), .dout(n19822));
    jdff dff_B_j4sQzHwf7_2(.din(n19822), .dout(n19825));
    jdff dff_B_dN0cZSOu0_2(.din(n19825), .dout(n19828));
    jdff dff_B_UaO0raDX3_2(.din(n19828), .dout(n19831));
    jdff dff_B_zAux4gZk5_2(.din(n19831), .dout(n19834));
    jdff dff_B_lKn1YUqf5_2(.din(n19834), .dout(n19837));
    jdff dff_B_386CQtn60_2(.din(n19837), .dout(n19840));
    jdff dff_B_rpCfMSGh8_2(.din(n19840), .dout(n19843));
    jdff dff_B_Sivw5WCI8_2(.din(n19843), .dout(n19846));
    jdff dff_B_h1mTn8qL8_2(.din(n19846), .dout(n19849));
    jdff dff_B_zQTzwlJ39_2(.din(n19849), .dout(n19852));
    jdff dff_B_wHbRWiRb4_2(.din(n19852), .dout(n19855));
    jdff dff_B_eSqY2FEm1_2(.din(n19855), .dout(n19858));
    jdff dff_B_Ty6trjOr3_1(.din(n3482), .dout(n19861));
    jdff dff_B_zyptDpkY2_2(.din(n3077), .dout(n19864));
    jdff dff_B_y4Ube5an2_2(.din(n19864), .dout(n19867));
    jdff dff_B_I4zNbDoI3_2(.din(n19867), .dout(n19870));
    jdff dff_B_iC6EmDSr4_2(.din(n19870), .dout(n19873));
    jdff dff_B_MrZ7h7iX8_2(.din(n19873), .dout(n19876));
    jdff dff_B_9C48Tz4M7_2(.din(n19876), .dout(n19879));
    jdff dff_B_eY43w6qp7_2(.din(n19879), .dout(n19882));
    jdff dff_B_94bRS6Zc3_2(.din(n19882), .dout(n19885));
    jdff dff_B_MnxwYbbG6_2(.din(n19885), .dout(n19888));
    jdff dff_B_FcPa4WaH5_2(.din(n19888), .dout(n19891));
    jdff dff_B_yTvnrMGf7_2(.din(n19891), .dout(n19894));
    jdff dff_B_tmnxWpXx3_2(.din(n19894), .dout(n19897));
    jdff dff_B_mP67yWkI7_2(.din(n19897), .dout(n19900));
    jdff dff_B_ZVEW2Wgg7_2(.din(n19900), .dout(n19903));
    jdff dff_B_jEqc3vX75_2(.din(n19903), .dout(n19906));
    jdff dff_B_meSBabrK2_2(.din(n19906), .dout(n19909));
    jdff dff_B_js3dBYcS8_2(.din(n19909), .dout(n19912));
    jdff dff_B_BNKNvkt61_2(.din(n19912), .dout(n19915));
    jdff dff_B_0xtg43hz4_2(.din(n19915), .dout(n19918));
    jdff dff_B_lgd5mQvA2_2(.din(n19918), .dout(n19921));
    jdff dff_B_sCW2FjgQ1_2(.din(n19921), .dout(n19924));
    jdff dff_B_hMKtJyxY7_2(.din(n19924), .dout(n19927));
    jdff dff_B_SgOIII2a1_2(.din(n19927), .dout(n19930));
    jdff dff_B_LwYy6BIU8_2(.din(n19930), .dout(n19933));
    jdff dff_B_NdHpaAPw4_2(.din(n19933), .dout(n19936));
    jdff dff_B_na7o3CWK8_2(.din(n19936), .dout(n19939));
    jdff dff_B_o4fmtzml8_2(.din(n19939), .dout(n19942));
    jdff dff_B_j1yGSPFY8_2(.din(n19942), .dout(n19945));
    jdff dff_B_aOKnKsbI5_1(.din(n3081), .dout(n19948));
    jdff dff_B_t8WFISp08_2(.din(n2698), .dout(n19951));
    jdff dff_B_44nP9i2V4_2(.din(n19951), .dout(n19954));
    jdff dff_B_5bAK6Yg66_2(.din(n19954), .dout(n19957));
    jdff dff_B_wihg9dZv6_2(.din(n19957), .dout(n19960));
    jdff dff_B_y7sptAQY7_2(.din(n19960), .dout(n19963));
    jdff dff_B_r347IwI28_2(.din(n19963), .dout(n19966));
    jdff dff_B_OyhCjVUy9_2(.din(n19966), .dout(n19969));
    jdff dff_B_Ab5EYeQs5_2(.din(n19969), .dout(n19972));
    jdff dff_B_5E4cWV1U8_2(.din(n19972), .dout(n19975));
    jdff dff_B_usSTADm85_2(.din(n19975), .dout(n19978));
    jdff dff_B_C9OMeGqX5_2(.din(n19978), .dout(n19981));
    jdff dff_B_EVQJ2NAe5_2(.din(n19981), .dout(n19984));
    jdff dff_B_zaFgKXCb5_2(.din(n19984), .dout(n19987));
    jdff dff_B_B9iZeQ1Q6_2(.din(n19987), .dout(n19990));
    jdff dff_B_76jpFiPs1_2(.din(n19990), .dout(n19993));
    jdff dff_B_GMAX2RNd1_2(.din(n19993), .dout(n19996));
    jdff dff_B_oYUp9omq1_2(.din(n19996), .dout(n19999));
    jdff dff_B_qFhHMkon7_2(.din(n19999), .dout(n20002));
    jdff dff_B_o3ablrzL1_2(.din(n20002), .dout(n20005));
    jdff dff_B_UQv29VuB1_2(.din(n20005), .dout(n20008));
    jdff dff_B_M7jLzGgz1_2(.din(n20008), .dout(n20011));
    jdff dff_B_PwLVjtrM8_2(.din(n20011), .dout(n20014));
    jdff dff_B_KYXnVwUT0_2(.din(n20014), .dout(n20017));
    jdff dff_B_kmKD18UZ3_2(.din(n20017), .dout(n20020));
    jdff dff_B_zR9qlZKD4_2(.din(n20020), .dout(n20023));
    jdff dff_B_F4vP9F4i6_1(.din(n2702), .dout(n20026));
    jdff dff_B_1p18hD567_2(.din(n2343), .dout(n20029));
    jdff dff_B_MLapcce12_2(.din(n20029), .dout(n20032));
    jdff dff_B_EBSLFvWC5_2(.din(n20032), .dout(n20035));
    jdff dff_B_APz24RGh2_2(.din(n20035), .dout(n20038));
    jdff dff_B_6mYl2Ci25_2(.din(n20038), .dout(n20041));
    jdff dff_B_AKhJBG480_2(.din(n20041), .dout(n20044));
    jdff dff_B_5i0imjQS0_2(.din(n20044), .dout(n20047));
    jdff dff_B_NUXUo0vc7_2(.din(n20047), .dout(n20050));
    jdff dff_B_spQShVNE1_2(.din(n20050), .dout(n20053));
    jdff dff_B_EQeg9lbJ2_2(.din(n20053), .dout(n20056));
    jdff dff_B_tLQFADPr9_2(.din(n20056), .dout(n20059));
    jdff dff_B_EP7XPJMF7_2(.din(n20059), .dout(n20062));
    jdff dff_B_l5VjWV6J7_2(.din(n20062), .dout(n20065));
    jdff dff_B_EhiQJxor2_2(.din(n20065), .dout(n20068));
    jdff dff_B_HoUupqzo8_2(.din(n20068), .dout(n20071));
    jdff dff_B_8xTQIdKM1_2(.din(n20071), .dout(n20074));
    jdff dff_B_eXlfqz2o1_2(.din(n20074), .dout(n20077));
    jdff dff_B_FRfXUKr84_2(.din(n20077), .dout(n20080));
    jdff dff_B_9KiotzSZ4_2(.din(n20080), .dout(n20083));
    jdff dff_B_W62zzIzD4_2(.din(n20083), .dout(n20086));
    jdff dff_B_3KK4QQkq5_2(.din(n20086), .dout(n20089));
    jdff dff_B_QpjVlIc90_2(.din(n20089), .dout(n20092));
    jdff dff_B_9M5pmyQ40_1(.din(n2347), .dout(n20095));
    jdff dff_B_3Oy4zAc83_2(.din(n2015), .dout(n20098));
    jdff dff_B_RbVCnQe98_2(.din(n20098), .dout(n20101));
    jdff dff_B_1pczOuZR7_2(.din(n20101), .dout(n20104));
    jdff dff_B_6yB0xafJ0_2(.din(n20104), .dout(n20107));
    jdff dff_B_SuSjQcXD1_2(.din(n20107), .dout(n20110));
    jdff dff_B_DxiDnaAc5_2(.din(n20110), .dout(n20113));
    jdff dff_B_qiywJnVB2_2(.din(n20113), .dout(n20116));
    jdff dff_B_WVtFyks58_2(.din(n20116), .dout(n20119));
    jdff dff_B_16hPDcOk3_2(.din(n20119), .dout(n20122));
    jdff dff_B_GIDQdYSE8_2(.din(n20122), .dout(n20125));
    jdff dff_B_hjY8zbRe0_2(.din(n20125), .dout(n20128));
    jdff dff_B_flV9nWky7_2(.din(n20128), .dout(n20131));
    jdff dff_B_f6MA30B28_2(.din(n20131), .dout(n20134));
    jdff dff_B_rtRNaiLF9_2(.din(n20134), .dout(n20137));
    jdff dff_B_Weew9LTl7_2(.din(n20137), .dout(n20140));
    jdff dff_B_sPbCZpbO2_2(.din(n20140), .dout(n20143));
    jdff dff_B_UX0a4oAJ7_2(.din(n20143), .dout(n20146));
    jdff dff_B_ifbYKzyJ1_2(.din(n20146), .dout(n20149));
    jdff dff_B_qqduDE2g4_2(.din(n20149), .dout(n20152));
    jdff dff_B_s9Cd84hT8_1(.din(n2019), .dout(n20155));
    jdff dff_B_ZSz19q7P4_2(.din(n1714), .dout(n20158));
    jdff dff_B_Lq2hAwIk1_2(.din(n20158), .dout(n20161));
    jdff dff_B_R58AkyAS8_2(.din(n20161), .dout(n20164));
    jdff dff_B_2bS28fJ98_2(.din(n20164), .dout(n20167));
    jdff dff_B_X2Svo9sr2_2(.din(n20167), .dout(n20170));
    jdff dff_B_JEo17NHy5_2(.din(n20170), .dout(n20173));
    jdff dff_B_SgkybFcA6_2(.din(n20173), .dout(n20176));
    jdff dff_B_LY8odb8R5_2(.din(n20176), .dout(n20179));
    jdff dff_B_rVpjdAN79_2(.din(n20179), .dout(n20182));
    jdff dff_B_lyJmV2WD3_2(.din(n20182), .dout(n20185));
    jdff dff_B_yUNS7d8j9_2(.din(n20185), .dout(n20188));
    jdff dff_B_So8gVGsf1_2(.din(n20188), .dout(n20191));
    jdff dff_B_E31YnTJc1_2(.din(n20191), .dout(n20194));
    jdff dff_B_SeWOF00b6_2(.din(n20194), .dout(n20197));
    jdff dff_B_1g9pyNQd0_2(.din(n20197), .dout(n20200));
    jdff dff_B_1WJwsVqu8_2(.din(n20200), .dout(n20203));
    jdff dff_B_qAkQqxEW1_1(.din(n1718), .dout(n20206));
    jdff dff_B_DRRdmiDW3_2(.din(n1440), .dout(n20209));
    jdff dff_B_urIvva7L5_2(.din(n20209), .dout(n20212));
    jdff dff_B_MuWDCOfI2_2(.din(n20212), .dout(n20215));
    jdff dff_B_IKxz5faF8_2(.din(n20215), .dout(n20218));
    jdff dff_B_MUQ3CgdL6_2(.din(n20218), .dout(n20221));
    jdff dff_B_atjKpGNi7_2(.din(n20221), .dout(n20224));
    jdff dff_B_OXNf1yG70_2(.din(n20224), .dout(n20227));
    jdff dff_B_1UWUrrwO9_2(.din(n20227), .dout(n20230));
    jdff dff_B_qce8hfQB1_2(.din(n20230), .dout(n20233));
    jdff dff_B_mGHPOroW1_2(.din(n20233), .dout(n20236));
    jdff dff_B_mHDzVxhK5_2(.din(n20236), .dout(n20239));
    jdff dff_B_Vu6i6Fll3_2(.din(n20239), .dout(n20242));
    jdff dff_B_WVEh5NPZ2_2(.din(n20242), .dout(n20245));
    jdff dff_B_BnZj7UBm8_1(.din(n1444), .dout(n20248));
    jdff dff_B_4QyvSVSR8_2(.din(n1196), .dout(n20251));
    jdff dff_B_IIx56gXe0_2(.din(n20251), .dout(n20254));
    jdff dff_B_6wZH7Ok81_2(.din(n20254), .dout(n20257));
    jdff dff_B_gkNvJvQH7_2(.din(n20257), .dout(n20260));
    jdff dff_B_PUvLPEbX8_2(.din(n20260), .dout(n20263));
    jdff dff_B_613AM2O79_2(.din(n20263), .dout(n20266));
    jdff dff_B_xrCZWvcG0_2(.din(n20266), .dout(n20269));
    jdff dff_B_ly6g3P1U1_2(.din(n20269), .dout(n20272));
    jdff dff_B_QaJT2DOY0_2(.din(n20272), .dout(n20275));
    jdff dff_B_wVO3rB1a0_2(.din(n20275), .dout(n20278));
    jdff dff_B_OOIwGHPY4_2(.din(n1280), .dout(n20281));
    jdff dff_B_TK43nvRb3_1(.din(n1200), .dout(n20284));
    jdff dff_B_L7G2pKg59_2(.din(n976), .dout(n20287));
    jdff dff_B_0KwACUyX9_2(.din(n20287), .dout(n20290));
    jdff dff_B_kIK5WVBH9_2(.din(n20290), .dout(n20293));
    jdff dff_B_8YKbz1RU8_2(.din(n20293), .dout(n20296));
    jdff dff_B_F5ySW75Y5_2(.din(n20296), .dout(n20299));
    jdff dff_B_ffnSJ3H53_2(.din(n20299), .dout(n20302));
    jdff dff_B_JqLKAmu29_2(.din(n20302), .dout(n20305));
    jdff dff_B_NxEO5AfJ9_2(.din(n1036), .dout(n20308));
    jdff dff_B_p983pDwu3_1(.din(n979), .dout(n20311));
    jdff dff_B_Lj5YMUYh5_2(.din(n782), .dout(n20314));
    jdff dff_B_xBmmamQh7_2(.din(n20314), .dout(n20317));
    jdff dff_B_JlmFxbUl8_2(.din(n20317), .dout(n20320));
    jdff dff_B_Cjc6iVEW9_2(.din(n20320), .dout(n20323));
    jdff dff_B_9IuVKnvE7_1(.din(n790), .dout(n20326));
    jdff dff_A_pnxRAwe47_1(.din(n616), .dout(n20328));
    jdff dff_A_bReyMFdL4_2(.din(n20334), .dout(n20331));
    jdff dff_A_MHJ6KRGP1_2(.din(n616), .dout(n20334));
    jdff dff_B_1PbYWcAW4_2(.din(n5528), .dout(n20338));
    jdff dff_B_RRuD0sth9_1(.din(n5520), .dout(n20341));
    jdff dff_B_phbo0j6D0_2(.din(n5241), .dout(n20344));
    jdff dff_B_8YVilGzq5_2(.din(n20344), .dout(n20347));
    jdff dff_B_BmzU59om7_2(.din(n20347), .dout(n20350));
    jdff dff_B_YVIktdGg6_2(.din(n20350), .dout(n20353));
    jdff dff_B_8ydDYcP81_2(.din(n20353), .dout(n20356));
    jdff dff_B_OQgfeYhR3_2(.din(n20356), .dout(n20359));
    jdff dff_B_G11Lskv29_2(.din(n20359), .dout(n20362));
    jdff dff_B_CQCWSLBS8_2(.din(n20362), .dout(n20365));
    jdff dff_B_sUEr4TXq0_2(.din(n20365), .dout(n20368));
    jdff dff_B_7MbSH3721_2(.din(n20368), .dout(n20371));
    jdff dff_B_SePz8io24_2(.din(n20371), .dout(n20374));
    jdff dff_B_NGQ8Tdl15_2(.din(n20374), .dout(n20377));
    jdff dff_B_lt75ed062_2(.din(n20377), .dout(n20380));
    jdff dff_B_VWqlhZly4_2(.din(n20380), .dout(n20383));
    jdff dff_B_ntIG5aVD8_2(.din(n20383), .dout(n20386));
    jdff dff_B_W8LSHsh81_2(.din(n20386), .dout(n20389));
    jdff dff_B_tSTUgfPQ8_2(.din(n20389), .dout(n20392));
    jdff dff_B_upkqrRwu6_2(.din(n20392), .dout(n20395));
    jdff dff_B_jy1WydnB1_2(.din(n20395), .dout(n20398));
    jdff dff_B_ohhgsH8T8_2(.din(n20398), .dout(n20401));
    jdff dff_B_stsMYuIm9_2(.din(n20401), .dout(n20404));
    jdff dff_B_U1tVEron5_2(.din(n20404), .dout(n20407));
    jdff dff_B_ZiUT98Jd3_2(.din(n20407), .dout(n20410));
    jdff dff_B_LaBPyo2r3_2(.din(n20410), .dout(n20413));
    jdff dff_B_GkAN6Om21_2(.din(n20413), .dout(n20416));
    jdff dff_B_tejtAvzC6_2(.din(n20416), .dout(n20419));
    jdff dff_B_cVencumn7_2(.din(n20419), .dout(n20422));
    jdff dff_B_IpnrKMFN1_2(.din(n20422), .dout(n20425));
    jdff dff_B_LjnXAPnO4_2(.din(n20425), .dout(n20428));
    jdff dff_B_INSiJQO72_2(.din(n20428), .dout(n20431));
    jdff dff_B_hKsAMLUP0_2(.din(n20431), .dout(n20434));
    jdff dff_B_oEVqmzXk3_2(.din(n20434), .dout(n20437));
    jdff dff_B_684SEqpv1_2(.din(n20437), .dout(n20440));
    jdff dff_B_SZaKRMyP0_2(.din(n20440), .dout(n20443));
    jdff dff_B_b7TOsfdU2_2(.din(n20443), .dout(n20446));
    jdff dff_B_GRC7YGEg7_2(.din(n20446), .dout(n20449));
    jdff dff_B_wBGrFOu90_2(.din(n20449), .dout(n20452));
    jdff dff_B_2ld1AzU40_2(.din(n20452), .dout(n20455));
    jdff dff_B_inHNCpSI0_2(.din(n20455), .dout(n20458));
    jdff dff_B_Q5QfrRvA9_2(.din(n20458), .dout(n20461));
    jdff dff_B_4HYX0Wkp9_2(.din(n20461), .dout(n20464));
    jdff dff_B_Z7CtsIPD6_2(.din(n20464), .dout(n20467));
    jdff dff_B_VF1cx7eZ3_2(.din(n20467), .dout(n20470));
    jdff dff_B_fExNCCvN4_2(.din(n20470), .dout(n20473));
    jdff dff_B_QRalWrY44_2(.din(n20473), .dout(n20476));
    jdff dff_B_wthlQ4w61_2(.din(n20476), .dout(n20479));
    jdff dff_B_sIuJ0ldn2_1(.din(n5245), .dout(n20482));
    jdff dff_B_6KJiEFqY2_2(.din(n4942), .dout(n20485));
    jdff dff_B_mw3p6vg57_2(.din(n20485), .dout(n20488));
    jdff dff_B_g5ipnwXZ8_2(.din(n20488), .dout(n20491));
    jdff dff_B_B7gmGxNR2_2(.din(n20491), .dout(n20494));
    jdff dff_B_Ti3DIU192_2(.din(n20494), .dout(n20497));
    jdff dff_B_lXKsN52i6_2(.din(n20497), .dout(n20500));
    jdff dff_B_1W4sHzwi9_2(.din(n20500), .dout(n20503));
    jdff dff_B_RAn4t7HL8_2(.din(n20503), .dout(n20506));
    jdff dff_B_ELJ6mODA6_2(.din(n20506), .dout(n20509));
    jdff dff_B_dwQbV2VH6_2(.din(n20509), .dout(n20512));
    jdff dff_B_O7zE7Wi63_2(.din(n20512), .dout(n20515));
    jdff dff_B_FtPLZGxp7_2(.din(n20515), .dout(n20518));
    jdff dff_B_649zuP3T6_2(.din(n20518), .dout(n20521));
    jdff dff_B_cFneH57W6_2(.din(n20521), .dout(n20524));
    jdff dff_B_DqeffqpD8_2(.din(n20524), .dout(n20527));
    jdff dff_B_bvBe0FNz4_2(.din(n20527), .dout(n20530));
    jdff dff_B_tywvN8aH2_2(.din(n20530), .dout(n20533));
    jdff dff_B_gLWEqJuP2_2(.din(n20533), .dout(n20536));
    jdff dff_B_6gYaM4J94_2(.din(n20536), .dout(n20539));
    jdff dff_B_RT9Hkvei7_2(.din(n20539), .dout(n20542));
    jdff dff_B_Zxgv8LjW3_2(.din(n20542), .dout(n20545));
    jdff dff_B_ZFv2T1Bh8_2(.din(n20545), .dout(n20548));
    jdff dff_B_DeWHq8RW5_2(.din(n20548), .dout(n20551));
    jdff dff_B_Fn2Kytrg2_2(.din(n20551), .dout(n20554));
    jdff dff_B_fOcOOTkF3_2(.din(n20554), .dout(n20557));
    jdff dff_B_wqZknIfA0_2(.din(n20557), .dout(n20560));
    jdff dff_B_XqwC3bhT1_2(.din(n20560), .dout(n20563));
    jdff dff_B_jiJk4psO8_2(.din(n20563), .dout(n20566));
    jdff dff_B_i43SwWRs6_2(.din(n20566), .dout(n20569));
    jdff dff_B_dXh13j5K4_2(.din(n20569), .dout(n20572));
    jdff dff_B_Kc0wYyDf7_2(.din(n20572), .dout(n20575));
    jdff dff_B_EvRJKgDR7_2(.din(n20575), .dout(n20578));
    jdff dff_B_NjoHizA18_2(.din(n20578), .dout(n20581));
    jdff dff_B_lotqe8Oh9_2(.din(n20581), .dout(n20584));
    jdff dff_B_AXmoDAIb4_2(.din(n20584), .dout(n20587));
    jdff dff_B_eLZ0OLec7_2(.din(n20587), .dout(n20590));
    jdff dff_B_wAglXE6F0_2(.din(n20590), .dout(n20593));
    jdff dff_B_UrBfy7n78_2(.din(n20593), .dout(n20596));
    jdff dff_B_odXcaD7i8_2(.din(n20596), .dout(n20599));
    jdff dff_B_M0LYrLI80_2(.din(n20599), .dout(n20602));
    jdff dff_B_Cg2CwX5J4_2(.din(n20602), .dout(n20605));
    jdff dff_B_1csLnxFv0_1(.din(n4946), .dout(n20608));
    jdff dff_B_b4kl91Zv3_2(.din(n4616), .dout(n20611));
    jdff dff_B_QsZYzkpk1_2(.din(n20611), .dout(n20614));
    jdff dff_B_tNrblsGQ5_2(.din(n20614), .dout(n20617));
    jdff dff_B_XxOCstFK5_2(.din(n20617), .dout(n20620));
    jdff dff_B_5ws6GyMH6_2(.din(n20620), .dout(n20623));
    jdff dff_B_XiBkvPrz0_2(.din(n20623), .dout(n20626));
    jdff dff_B_ANZU9JIL9_2(.din(n20626), .dout(n20629));
    jdff dff_B_S7iFtZF05_2(.din(n20629), .dout(n20632));
    jdff dff_B_G8OgqTJ99_2(.din(n20632), .dout(n20635));
    jdff dff_B_nNTVIRhW9_2(.din(n20635), .dout(n20638));
    jdff dff_B_Fq3mlY0W3_2(.din(n20638), .dout(n20641));
    jdff dff_B_42xAzjpx3_2(.din(n20641), .dout(n20644));
    jdff dff_B_PBaV0l5S1_2(.din(n20644), .dout(n20647));
    jdff dff_B_uNJs50bg3_2(.din(n20647), .dout(n20650));
    jdff dff_B_nJdHJFwc2_2(.din(n20650), .dout(n20653));
    jdff dff_B_UTjvwtPY6_2(.din(n20653), .dout(n20656));
    jdff dff_B_IjWk86Bp9_2(.din(n20656), .dout(n20659));
    jdff dff_B_pnuPGRxD0_2(.din(n20659), .dout(n20662));
    jdff dff_B_x8cpswUn2_2(.din(n20662), .dout(n20665));
    jdff dff_B_fGzF0AhU7_2(.din(n20665), .dout(n20668));
    jdff dff_B_bFI6WgSD4_2(.din(n20668), .dout(n20671));
    jdff dff_B_095JIYNe4_2(.din(n20671), .dout(n20674));
    jdff dff_B_EiJlTDHF4_2(.din(n20674), .dout(n20677));
    jdff dff_B_bQNSlO170_2(.din(n20677), .dout(n20680));
    jdff dff_B_NB2NLA2v6_2(.din(n20680), .dout(n20683));
    jdff dff_B_MGxVDMPn2_2(.din(n20683), .dout(n20686));
    jdff dff_B_ZXh3Z5mH3_2(.din(n20686), .dout(n20689));
    jdff dff_B_lqvgRkIg5_2(.din(n20689), .dout(n20692));
    jdff dff_B_Ec17dfrk4_2(.din(n20692), .dout(n20695));
    jdff dff_B_ASikrecF2_2(.din(n20695), .dout(n20698));
    jdff dff_B_oUB0YSab3_2(.din(n20698), .dout(n20701));
    jdff dff_B_rR8EqmPP1_2(.din(n20701), .dout(n20704));
    jdff dff_B_zjR6gQcK8_2(.din(n20704), .dout(n20707));
    jdff dff_B_OwcYP0uH8_2(.din(n20707), .dout(n20710));
    jdff dff_B_3d7wCdrG2_2(.din(n20710), .dout(n20713));
    jdff dff_B_mahCikNx5_2(.din(n20713), .dout(n20716));
    jdff dff_B_si4xxSjr1_2(.din(n20716), .dout(n20719));
    jdff dff_B_qyzV3BIc3_2(.din(n20719), .dout(n20722));
    jdff dff_B_9SfuAkYY9_1(.din(n4620), .dout(n20725));
    jdff dff_B_FsMcM0tO7_2(.din(n4270), .dout(n20728));
    jdff dff_B_2ED1pqdD9_2(.din(n20728), .dout(n20731));
    jdff dff_B_jzNsQ8RR5_2(.din(n20731), .dout(n20734));
    jdff dff_B_PRx9EmQN4_2(.din(n20734), .dout(n20737));
    jdff dff_B_GtqUXrql6_2(.din(n20737), .dout(n20740));
    jdff dff_B_JnZ8EYwP5_2(.din(n20740), .dout(n20743));
    jdff dff_B_5tNGFGjg9_2(.din(n20743), .dout(n20746));
    jdff dff_B_ddYVAcUU7_2(.din(n20746), .dout(n20749));
    jdff dff_B_5YFqgaWt4_2(.din(n20749), .dout(n20752));
    jdff dff_B_oUbmb7iS9_2(.din(n20752), .dout(n20755));
    jdff dff_B_Kqs9sEQy3_2(.din(n20755), .dout(n20758));
    jdff dff_B_o7EUY3su9_2(.din(n20758), .dout(n20761));
    jdff dff_B_mFHopx8k7_2(.din(n20761), .dout(n20764));
    jdff dff_B_vPeapwCx7_2(.din(n20764), .dout(n20767));
    jdff dff_B_LntdU5Z96_2(.din(n20767), .dout(n20770));
    jdff dff_B_LlkzF4AE4_2(.din(n20770), .dout(n20773));
    jdff dff_B_UoDF4jVm3_2(.din(n20773), .dout(n20776));
    jdff dff_B_mlborhS82_2(.din(n20776), .dout(n20779));
    jdff dff_B_kv6fnce34_2(.din(n20779), .dout(n20782));
    jdff dff_B_F5EZnrfI6_2(.din(n20782), .dout(n20785));
    jdff dff_B_hg5VPneE7_2(.din(n20785), .dout(n20788));
    jdff dff_B_Zc12SvIE2_2(.din(n20788), .dout(n20791));
    jdff dff_B_9JW8665k2_2(.din(n20791), .dout(n20794));
    jdff dff_B_GC3jK5Dl2_2(.din(n20794), .dout(n20797));
    jdff dff_B_g7K8x2lD0_2(.din(n20797), .dout(n20800));
    jdff dff_B_9zfFNM3v5_2(.din(n20800), .dout(n20803));
    jdff dff_B_vfkppYBB0_2(.din(n20803), .dout(n20806));
    jdff dff_B_JWG6VLI99_2(.din(n20806), .dout(n20809));
    jdff dff_B_xwEi4aM58_2(.din(n20809), .dout(n20812));
    jdff dff_B_m2V0cs3H6_2(.din(n20812), .dout(n20815));
    jdff dff_B_uhzNH2U43_2(.din(n20815), .dout(n20818));
    jdff dff_B_y8yadeKv2_2(.din(n20818), .dout(n20821));
    jdff dff_B_J8TzKbhy6_2(.din(n20821), .dout(n20824));
    jdff dff_B_v8I2cg8R8_2(.din(n20824), .dout(n20827));
    jdff dff_B_22AifnwD9_2(.din(n20827), .dout(n20830));
    jdff dff_B_Ow6XnM5z2_1(.din(n4274), .dout(n20833));
    jdff dff_B_fXdVR7Yh4_2(.din(n3874), .dout(n20836));
    jdff dff_B_P4h4V8Nh2_2(.din(n20836), .dout(n20839));
    jdff dff_B_HxI3PnX11_2(.din(n20839), .dout(n20842));
    jdff dff_B_KWBjY2yn2_2(.din(n20842), .dout(n20845));
    jdff dff_B_mKkk714A4_2(.din(n20845), .dout(n20848));
    jdff dff_B_qJJthC0G1_2(.din(n20848), .dout(n20851));
    jdff dff_B_mxh4hOpr8_2(.din(n20851), .dout(n20854));
    jdff dff_B_M77jESMV4_2(.din(n20854), .dout(n20857));
    jdff dff_B_mW368jgu3_2(.din(n20857), .dout(n20860));
    jdff dff_B_3CodNuHe9_2(.din(n20860), .dout(n20863));
    jdff dff_B_qmSuJsmC7_2(.din(n20863), .dout(n20866));
    jdff dff_B_cOYrjpoi4_2(.din(n20866), .dout(n20869));
    jdff dff_B_Z18h3vrZ8_2(.din(n20869), .dout(n20872));
    jdff dff_B_lYFzWjRi4_2(.din(n20872), .dout(n20875));
    jdff dff_B_qvJ3F9DW2_2(.din(n20875), .dout(n20878));
    jdff dff_B_Hf6gstuf4_2(.din(n20878), .dout(n20881));
    jdff dff_B_C5NwgdrA5_2(.din(n20881), .dout(n20884));
    jdff dff_B_YvHI9ZI63_2(.din(n20884), .dout(n20887));
    jdff dff_B_P5xYgdSi5_2(.din(n20887), .dout(n20890));
    jdff dff_B_W5nzsXYb7_2(.din(n20890), .dout(n20893));
    jdff dff_B_vlnoy0995_2(.din(n20893), .dout(n20896));
    jdff dff_B_D3JC63K48_2(.din(n20896), .dout(n20899));
    jdff dff_B_PaiYz4uk8_2(.din(n20899), .dout(n20902));
    jdff dff_B_4dNax5Ww0_2(.din(n20902), .dout(n20905));
    jdff dff_B_QXnmCyxB3_2(.din(n20905), .dout(n20908));
    jdff dff_B_1OwSHxWC7_2(.din(n20908), .dout(n20911));
    jdff dff_B_K27QHcQL5_2(.din(n20911), .dout(n20914));
    jdff dff_B_dAPh4Opn0_2(.din(n20914), .dout(n20917));
    jdff dff_B_dAL4aXgJ4_2(.din(n20917), .dout(n20920));
    jdff dff_B_N9dgmGfc2_2(.din(n20920), .dout(n20923));
    jdff dff_B_ZWAQwnOr9_2(.din(n20923), .dout(n20926));
    jdff dff_B_PMFJBWlE4_2(.din(n20926), .dout(n20929));
    jdff dff_B_Z0oss8sb3_1(.din(n3878), .dout(n20932));
    jdff dff_B_Mwi8CdeB6_2(.din(n3497), .dout(n20935));
    jdff dff_B_z5EpUGAC6_2(.din(n20935), .dout(n20938));
    jdff dff_B_XH4IWRzp9_2(.din(n20938), .dout(n20941));
    jdff dff_B_K2wgqb1J8_2(.din(n20941), .dout(n20944));
    jdff dff_B_hbks4zt12_2(.din(n20944), .dout(n20947));
    jdff dff_B_qyTI3Nyt3_2(.din(n20947), .dout(n20950));
    jdff dff_B_Dyoe2unM8_2(.din(n20950), .dout(n20953));
    jdff dff_B_pBRBWnLh8_2(.din(n20953), .dout(n20956));
    jdff dff_B_QcXGHQf89_2(.din(n20956), .dout(n20959));
    jdff dff_B_Fw28KfIW4_2(.din(n20959), .dout(n20962));
    jdff dff_B_PIOMStCF6_2(.din(n20962), .dout(n20965));
    jdff dff_B_gShgcL5Z6_2(.din(n20965), .dout(n20968));
    jdff dff_B_rie49QFk7_2(.din(n20968), .dout(n20971));
    jdff dff_B_SuTYyFwc0_2(.din(n20971), .dout(n20974));
    jdff dff_B_3z9HK80M4_2(.din(n20974), .dout(n20977));
    jdff dff_B_riCzz8px7_2(.din(n20977), .dout(n20980));
    jdff dff_B_rWRAWtER1_2(.din(n20980), .dout(n20983));
    jdff dff_B_wxI1J3450_2(.din(n20983), .dout(n20986));
    jdff dff_B_3LSC9JC04_2(.din(n20986), .dout(n20989));
    jdff dff_B_H4NMfe866_2(.din(n20989), .dout(n20992));
    jdff dff_B_Be4zUztE7_2(.din(n20992), .dout(n20995));
    jdff dff_B_fnUFx6UZ3_2(.din(n20995), .dout(n20998));
    jdff dff_B_durrI5fz2_2(.din(n20998), .dout(n21001));
    jdff dff_B_AGj8QWtJ3_2(.din(n21001), .dout(n21004));
    jdff dff_B_70vRGkCI2_2(.din(n21004), .dout(n21007));
    jdff dff_B_RgH76awt7_2(.din(n21007), .dout(n21010));
    jdff dff_B_xFU6vod69_2(.din(n21010), .dout(n21013));
    jdff dff_B_SadRMwjg6_2(.din(n21013), .dout(n21016));
    jdff dff_B_vTxBxvLn4_2(.din(n21016), .dout(n21019));
    jdff dff_B_rM9QpD1R3_1(.din(n3501), .dout(n21022));
    jdff dff_B_5dAVkk415_2(.din(n3096), .dout(n21025));
    jdff dff_B_aEObCI7S3_2(.din(n21025), .dout(n21028));
    jdff dff_B_q4kr5DnY3_2(.din(n21028), .dout(n21031));
    jdff dff_B_TsoL5NO09_2(.din(n21031), .dout(n21034));
    jdff dff_B_w0g1rqsj8_2(.din(n21034), .dout(n21037));
    jdff dff_B_uz6FBTgE1_2(.din(n21037), .dout(n21040));
    jdff dff_B_ifSb8xnW1_2(.din(n21040), .dout(n21043));
    jdff dff_B_twNRafDj6_2(.din(n21043), .dout(n21046));
    jdff dff_B_RWbUv56y6_2(.din(n21046), .dout(n21049));
    jdff dff_B_wJEGs35L2_2(.din(n21049), .dout(n21052));
    jdff dff_B_wrFkDeYM7_2(.din(n21052), .dout(n21055));
    jdff dff_B_IDmoxZk77_2(.din(n21055), .dout(n21058));
    jdff dff_B_K1cx9ejt3_2(.din(n21058), .dout(n21061));
    jdff dff_B_Xz83PU8N3_2(.din(n21061), .dout(n21064));
    jdff dff_B_9MEZUAb25_2(.din(n21064), .dout(n21067));
    jdff dff_B_VJnHLuVn6_2(.din(n21067), .dout(n21070));
    jdff dff_B_u5l4rsjr6_2(.din(n21070), .dout(n21073));
    jdff dff_B_QLfIW2Nn0_2(.din(n21073), .dout(n21076));
    jdff dff_B_Tn4eHpk71_2(.din(n21076), .dout(n21079));
    jdff dff_B_pLlPYgku6_2(.din(n21079), .dout(n21082));
    jdff dff_B_1D5k8vXx1_2(.din(n21082), .dout(n21085));
    jdff dff_B_EkusFtkZ6_2(.din(n21085), .dout(n21088));
    jdff dff_B_7mTBadUp4_2(.din(n21088), .dout(n21091));
    jdff dff_B_gPHTXJU91_2(.din(n21091), .dout(n21094));
    jdff dff_B_eWwKaM8K4_2(.din(n21094), .dout(n21097));
    jdff dff_B_Bg6ghQej4_2(.din(n21097), .dout(n21100));
    jdff dff_B_QYADrKf36_1(.din(n3100), .dout(n21103));
    jdff dff_B_iqYUAous7_2(.din(n2717), .dout(n21106));
    jdff dff_B_IEgBySH99_2(.din(n21106), .dout(n21109));
    jdff dff_B_nmKsp4GW7_2(.din(n21109), .dout(n21112));
    jdff dff_B_sSrGumgj2_2(.din(n21112), .dout(n21115));
    jdff dff_B_2xqrFsFT3_2(.din(n21115), .dout(n21118));
    jdff dff_B_PeuKAcu55_2(.din(n21118), .dout(n21121));
    jdff dff_B_O6TyCTLV1_2(.din(n21121), .dout(n21124));
    jdff dff_B_V4O8t3vE8_2(.din(n21124), .dout(n21127));
    jdff dff_B_nh2rqO655_2(.din(n21127), .dout(n21130));
    jdff dff_B_tkHSC4hs7_2(.din(n21130), .dout(n21133));
    jdff dff_B_WVMS96HE7_2(.din(n21133), .dout(n21136));
    jdff dff_B_SklZIgxa3_2(.din(n21136), .dout(n21139));
    jdff dff_B_DqNHx9xf9_2(.din(n21139), .dout(n21142));
    jdff dff_B_Lc8xv4eH8_2(.din(n21142), .dout(n21145));
    jdff dff_B_0C8Y6kl37_2(.din(n21145), .dout(n21148));
    jdff dff_B_MusmQAan0_2(.din(n21148), .dout(n21151));
    jdff dff_B_2jQ2rd5G9_2(.din(n21151), .dout(n21154));
    jdff dff_B_bbKFYL1K1_2(.din(n21154), .dout(n21157));
    jdff dff_B_dGWY89kj9_2(.din(n21157), .dout(n21160));
    jdff dff_B_aUznYYAe2_2(.din(n21160), .dout(n21163));
    jdff dff_B_rGFNe1vY4_2(.din(n21163), .dout(n21166));
    jdff dff_B_mIlvcbW99_2(.din(n21166), .dout(n21169));
    jdff dff_B_GrOGSWfp7_2(.din(n21169), .dout(n21172));
    jdff dff_B_j9Ffr4DS0_1(.din(n2721), .dout(n21175));
    jdff dff_B_S7TvtqRR6_2(.din(n2362), .dout(n21178));
    jdff dff_B_wU3lPNwg6_2(.din(n21178), .dout(n21181));
    jdff dff_B_KvYMa5gq0_2(.din(n21181), .dout(n21184));
    jdff dff_B_JcfDtML31_2(.din(n21184), .dout(n21187));
    jdff dff_B_F6mLJgiV3_2(.din(n21187), .dout(n21190));
    jdff dff_B_HiaFSaBM4_2(.din(n21190), .dout(n21193));
    jdff dff_B_S2wL8ocN7_2(.din(n21193), .dout(n21196));
    jdff dff_B_6L2vsn9P1_2(.din(n21196), .dout(n21199));
    jdff dff_B_EXuGGKSs2_2(.din(n21199), .dout(n21202));
    jdff dff_B_j8iIcsy09_2(.din(n21202), .dout(n21205));
    jdff dff_B_8OE73jPJ3_2(.din(n21205), .dout(n21208));
    jdff dff_B_LPNmaUta7_2(.din(n21208), .dout(n21211));
    jdff dff_B_0gKLIgS97_2(.din(n21211), .dout(n21214));
    jdff dff_B_zJhJNn6o8_2(.din(n21214), .dout(n21217));
    jdff dff_B_f8npws4O8_2(.din(n21217), .dout(n21220));
    jdff dff_B_NJOTFBwo4_2(.din(n21220), .dout(n21223));
    jdff dff_B_PQd7iCdk7_2(.din(n21223), .dout(n21226));
    jdff dff_B_dgvqKwQl5_2(.din(n21226), .dout(n21229));
    jdff dff_B_9uQXoqq93_2(.din(n21229), .dout(n21232));
    jdff dff_B_BUOFNaTh0_2(.din(n21232), .dout(n21235));
    jdff dff_B_mW1TSD8L4_1(.din(n2366), .dout(n21238));
    jdff dff_B_WKBOTvv13_2(.din(n2034), .dout(n21241));
    jdff dff_B_sqn5zKLR6_2(.din(n21241), .dout(n21244));
    jdff dff_B_JV4GuYjx5_2(.din(n21244), .dout(n21247));
    jdff dff_B_69kkkViF9_2(.din(n21247), .dout(n21250));
    jdff dff_B_M0pxyStW1_2(.din(n21250), .dout(n21253));
    jdff dff_B_Es4cV7i55_2(.din(n21253), .dout(n21256));
    jdff dff_B_zMfhwVej3_2(.din(n21256), .dout(n21259));
    jdff dff_B_CtmUTiVC0_2(.din(n21259), .dout(n21262));
    jdff dff_B_zCyAhcLj0_2(.din(n21262), .dout(n21265));
    jdff dff_B_iKz7KXCa2_2(.din(n21265), .dout(n21268));
    jdff dff_B_a8n0zfU29_2(.din(n21268), .dout(n21271));
    jdff dff_B_PhDtRwzW1_2(.din(n21271), .dout(n21274));
    jdff dff_B_Dz0DTGEy6_2(.din(n21274), .dout(n21277));
    jdff dff_B_QU4yYePb4_2(.din(n21277), .dout(n21280));
    jdff dff_B_CS5SZ2Kk7_2(.din(n21280), .dout(n21283));
    jdff dff_B_ACczwGNs0_2(.din(n21283), .dout(n21286));
    jdff dff_B_8w35Olta4_2(.din(n21286), .dout(n21289));
    jdff dff_B_1jkOuCTe1_1(.din(n2038), .dout(n21292));
    jdff dff_B_UU0niQwW9_2(.din(n1733), .dout(n21295));
    jdff dff_B_KeVEyKMb1_2(.din(n21295), .dout(n21298));
    jdff dff_B_IfGQKgo49_2(.din(n21298), .dout(n21301));
    jdff dff_B_v8NkCyuF8_2(.din(n21301), .dout(n21304));
    jdff dff_B_DmBSNOsi5_2(.din(n21304), .dout(n21307));
    jdff dff_B_Bx2gnNGo9_2(.din(n21307), .dout(n21310));
    jdff dff_B_B5o8vsOp5_2(.din(n21310), .dout(n21313));
    jdff dff_B_8WFP1M3O3_2(.din(n21313), .dout(n21316));
    jdff dff_B_EtJZypqQ0_2(.din(n21316), .dout(n21319));
    jdff dff_B_2hTid2xz7_2(.din(n21319), .dout(n21322));
    jdff dff_B_wIPEjqCa4_2(.din(n21322), .dout(n21325));
    jdff dff_B_t2VXvQob3_2(.din(n21325), .dout(n21328));
    jdff dff_B_ugtxxaRF8_2(.din(n21328), .dout(n21331));
    jdff dff_B_4A2pXL0w9_2(.din(n21331), .dout(n21334));
    jdff dff_B_o1AElAy04_1(.din(n1737), .dout(n21337));
    jdff dff_B_yaTJdMX62_2(.din(n1459), .dout(n21340));
    jdff dff_B_0xzqZkN16_2(.din(n21340), .dout(n21343));
    jdff dff_B_x4Y8O32m2_2(.din(n21343), .dout(n21346));
    jdff dff_B_bjdxf3zh8_2(.din(n21346), .dout(n21349));
    jdff dff_B_QQPzpzg94_2(.din(n21349), .dout(n21352));
    jdff dff_B_Ygl76m6v6_2(.din(n21352), .dout(n21355));
    jdff dff_B_F1A8SqEE5_2(.din(n21355), .dout(n21358));
    jdff dff_B_9Ppv3XtM6_2(.din(n21358), .dout(n21361));
    jdff dff_B_csYC4KPe7_2(.din(n21361), .dout(n21364));
    jdff dff_B_REcqCrEE4_2(.din(n21364), .dout(n21367));
    jdff dff_B_t22o2eFd8_2(.din(n21367), .dout(n21370));
    jdff dff_B_1TPbLWoN5_2(.din(n1471), .dout(n21373));
    jdff dff_B_OO1D15tP2_1(.din(n1463), .dout(n21376));
    jdff dff_B_9zEPRubG3_2(.din(n1215), .dout(n21379));
    jdff dff_B_sqaADirs6_2(.din(n21379), .dout(n21382));
    jdff dff_B_fWKoUnXJ9_2(.din(n21382), .dout(n21385));
    jdff dff_B_QunNc8Us6_2(.din(n21385), .dout(n21388));
    jdff dff_B_feEC5aAb8_2(.din(n21388), .dout(n21391));
    jdff dff_B_ShoRSDqQ1_2(.din(n21391), .dout(n21394));
    jdff dff_B_xUKku5GK7_2(.din(n21394), .dout(n21397));
    jdff dff_B_03fXdbCs7_1(.din(n1218), .dout(n21400));
    jdff dff_B_wUHlHhtp4_2(.din(n994), .dout(n21403));
    jdff dff_B_YPvNkcuG0_2(.din(n21403), .dout(n21406));
    jdff dff_B_gIDleT7U8_2(.din(n21406), .dout(n21409));
    jdff dff_B_InSP26yk6_2(.din(n21409), .dout(n21412));
    jdff dff_B_pBKm8eeb1_1(.din(n1002), .dout(n21415));
    jdff dff_A_ND5nyXI76_0(.din(n798), .dout(n21417));
    jdff dff_A_Sleh7iQV6_1(.din(n21423), .dout(n21420));
    jdff dff_A_oB75lPv25_1(.din(n798), .dout(n21423));
    jdff dff_B_dscEN8CP3_1(.din(n5784), .dout(n21427));
    jdff dff_B_gZs9LaEz2_2(.din(n5532), .dout(n21430));
    jdff dff_B_PGEfNWI99_2(.din(n21430), .dout(n21433));
    jdff dff_B_W1Ek9dO77_2(.din(n21433), .dout(n21436));
    jdff dff_B_DDxqsWXw0_2(.din(n21436), .dout(n21439));
    jdff dff_B_OIYPBMRb4_2(.din(n21439), .dout(n21442));
    jdff dff_B_3syitiH25_2(.din(n21442), .dout(n21445));
    jdff dff_B_X0r7ewxt6_2(.din(n21445), .dout(n21448));
    jdff dff_B_YVKeeVHG7_2(.din(n21448), .dout(n21451));
    jdff dff_B_0KiXGFQ22_2(.din(n21451), .dout(n21454));
    jdff dff_B_OrxITFSE4_2(.din(n21454), .dout(n21457));
    jdff dff_B_p5XSaOeV3_2(.din(n21457), .dout(n21460));
    jdff dff_B_gX0PHthV9_2(.din(n21460), .dout(n21463));
    jdff dff_B_tSmN1HZK4_2(.din(n21463), .dout(n21466));
    jdff dff_B_bCg1fvIv9_2(.din(n21466), .dout(n21469));
    jdff dff_B_4rhMCbdM3_2(.din(n21469), .dout(n21472));
    jdff dff_B_zKAIuavT5_2(.din(n21472), .dout(n21475));
    jdff dff_B_WcE5HeEP9_2(.din(n21475), .dout(n21478));
    jdff dff_B_3v0Yo8XO9_2(.din(n21478), .dout(n21481));
    jdff dff_B_qz1XyZz10_2(.din(n21481), .dout(n21484));
    jdff dff_B_up5Fvazq8_2(.din(n21484), .dout(n21487));
    jdff dff_B_v26EmyiN3_2(.din(n21487), .dout(n21490));
    jdff dff_B_ybA0UQjG3_2(.din(n21490), .dout(n21493));
    jdff dff_B_gF3nxzH06_2(.din(n21493), .dout(n21496));
    jdff dff_B_iAAMCwx31_2(.din(n21496), .dout(n21499));
    jdff dff_B_3MjKph8N1_2(.din(n21499), .dout(n21502));
    jdff dff_B_5RdFssbW6_2(.din(n21502), .dout(n21505));
    jdff dff_B_uJfkE8X17_2(.din(n21505), .dout(n21508));
    jdff dff_B_w5zmZzTC5_2(.din(n21508), .dout(n21511));
    jdff dff_B_1goNVmJf8_2(.din(n21511), .dout(n21514));
    jdff dff_B_RwHDKR2h5_2(.din(n21514), .dout(n21517));
    jdff dff_B_SsVQtzwa4_2(.din(n21517), .dout(n21520));
    jdff dff_B_TzmBMLPI6_2(.din(n21520), .dout(n21523));
    jdff dff_B_H094nLHV7_2(.din(n21523), .dout(n21526));
    jdff dff_B_YWili5MT2_2(.din(n21526), .dout(n21529));
    jdff dff_B_NXZJJkEl4_2(.din(n21529), .dout(n21532));
    jdff dff_B_eODnW7n96_2(.din(n21532), .dout(n21535));
    jdff dff_B_VVeJMVTu0_2(.din(n21535), .dout(n21538));
    jdff dff_B_AFw9awkp9_2(.din(n21538), .dout(n21541));
    jdff dff_B_F4SSRS5d3_2(.din(n21541), .dout(n21544));
    jdff dff_B_unPgbOLe3_2(.din(n21544), .dout(n21547));
    jdff dff_B_xC7olaV15_2(.din(n21547), .dout(n21550));
    jdff dff_B_oWqxCd2C4_2(.din(n21550), .dout(n21553));
    jdff dff_B_XnMTc3tc5_2(.din(n21553), .dout(n21556));
    jdff dff_B_0UDdrsng6_2(.din(n21556), .dout(n21559));
    jdff dff_B_OdFVZsp64_2(.din(n21559), .dout(n21562));
    jdff dff_B_CeQ2fuut0_2(.din(n21562), .dout(n21565));
    jdff dff_B_ePm4FQ1L1_2(.din(n21565), .dout(n21568));
    jdff dff_B_xVbS7BIv1_0(.din(n5780), .dout(n21571));
    jdff dff_A_NoaSoI4S5_1(.din(n5737), .dout(n21573));
    jdff dff_B_lQf6csxZ2_1(.din(n5536), .dout(n21577));
    jdff dff_B_K8kUTWgq2_2(.din(n5260), .dout(n21580));
    jdff dff_B_CedpvwHs7_2(.din(n21580), .dout(n21583));
    jdff dff_B_7r2aTGij9_2(.din(n21583), .dout(n21586));
    jdff dff_B_dLvlGtDV0_2(.din(n21586), .dout(n21589));
    jdff dff_B_CMj8XDe25_2(.din(n21589), .dout(n21592));
    jdff dff_B_Y5UX4S5g2_2(.din(n21592), .dout(n21595));
    jdff dff_B_fGnOEmCY6_2(.din(n21595), .dout(n21598));
    jdff dff_B_dFvKUDWG2_2(.din(n21598), .dout(n21601));
    jdff dff_B_LZLEP57y7_2(.din(n21601), .dout(n21604));
    jdff dff_B_mL2VAuwq7_2(.din(n21604), .dout(n21607));
    jdff dff_B_QiyUvBsP5_2(.din(n21607), .dout(n21610));
    jdff dff_B_8zxexqDf3_2(.din(n21610), .dout(n21613));
    jdff dff_B_6oIlwFf77_2(.din(n21613), .dout(n21616));
    jdff dff_B_QIeW735N2_2(.din(n21616), .dout(n21619));
    jdff dff_B_t8xIgAYJ0_2(.din(n21619), .dout(n21622));
    jdff dff_B_WjDxrsoN8_2(.din(n21622), .dout(n21625));
    jdff dff_B_RJ1DzOCD2_2(.din(n21625), .dout(n21628));
    jdff dff_B_dPpnypC14_2(.din(n21628), .dout(n21631));
    jdff dff_B_YtEO3TLT3_2(.din(n21631), .dout(n21634));
    jdff dff_B_UarUl7fZ6_2(.din(n21634), .dout(n21637));
    jdff dff_B_Sj5WLCgo6_2(.din(n21637), .dout(n21640));
    jdff dff_B_s5q85r9E2_2(.din(n21640), .dout(n21643));
    jdff dff_B_ALefSdLr9_2(.din(n21643), .dout(n21646));
    jdff dff_B_24P93rEn5_2(.din(n21646), .dout(n21649));
    jdff dff_B_DouM5BnR5_2(.din(n21649), .dout(n21652));
    jdff dff_B_XicY1ay78_2(.din(n21652), .dout(n21655));
    jdff dff_B_MpMpxdGa3_2(.din(n21655), .dout(n21658));
    jdff dff_B_8XS9pli16_2(.din(n21658), .dout(n21661));
    jdff dff_B_dfwLvLV80_2(.din(n21661), .dout(n21664));
    jdff dff_B_eMQrLM579_2(.din(n21664), .dout(n21667));
    jdff dff_B_0g7HKPQi8_2(.din(n21667), .dout(n21670));
    jdff dff_B_gmFrnxSi7_2(.din(n21670), .dout(n21673));
    jdff dff_B_LHpRKbC69_2(.din(n21673), .dout(n21676));
    jdff dff_B_W5N0RPnN5_2(.din(n21676), .dout(n21679));
    jdff dff_B_RUCj2EVl5_2(.din(n21679), .dout(n21682));
    jdff dff_B_lfATVw4Z2_2(.din(n21682), .dout(n21685));
    jdff dff_B_9OaOwsta5_2(.din(n21685), .dout(n21688));
    jdff dff_B_5TU4Zch19_2(.din(n21688), .dout(n21691));
    jdff dff_B_mNTGIM3g0_2(.din(n21691), .dout(n21694));
    jdff dff_B_BNmq484u1_2(.din(n21694), .dout(n21697));
    jdff dff_B_ld4nXSo43_2(.din(n21697), .dout(n21700));
    jdff dff_B_hnjWvXPB6_2(.din(n21700), .dout(n21703));
    jdff dff_B_yDwue3896_2(.din(n5465), .dout(n21706));
    jdff dff_B_GNK67qew6_1(.din(n5264), .dout(n21709));
    jdff dff_B_mjwuSWFV6_2(.din(n4961), .dout(n21712));
    jdff dff_B_U9B1suxo8_2(.din(n21712), .dout(n21715));
    jdff dff_B_gb66n7Gz7_2(.din(n21715), .dout(n21718));
    jdff dff_B_M8ox9jiE1_2(.din(n21718), .dout(n21721));
    jdff dff_B_N6QIAid07_2(.din(n21721), .dout(n21724));
    jdff dff_B_Lx054sw25_2(.din(n21724), .dout(n21727));
    jdff dff_B_FCemGsSY4_2(.din(n21727), .dout(n21730));
    jdff dff_B_KJFQD4d71_2(.din(n21730), .dout(n21733));
    jdff dff_B_2u4iloU37_2(.din(n21733), .dout(n21736));
    jdff dff_B_nOkojfNl0_2(.din(n21736), .dout(n21739));
    jdff dff_B_23B6pC2S5_2(.din(n21739), .dout(n21742));
    jdff dff_B_MLegzzsA6_2(.din(n21742), .dout(n21745));
    jdff dff_B_qfg5kSDx2_2(.din(n21745), .dout(n21748));
    jdff dff_B_1abGkJLL3_2(.din(n21748), .dout(n21751));
    jdff dff_B_kRKuTYsx8_2(.din(n21751), .dout(n21754));
    jdff dff_B_Ku8lmRN92_2(.din(n21754), .dout(n21757));
    jdff dff_B_063y1oDD3_2(.din(n21757), .dout(n21760));
    jdff dff_B_4dR0k1Pe3_2(.din(n21760), .dout(n21763));
    jdff dff_B_uI4duSeb9_2(.din(n21763), .dout(n21766));
    jdff dff_B_ekNn9Kd60_2(.din(n21766), .dout(n21769));
    jdff dff_B_eNOnXkzs7_2(.din(n21769), .dout(n21772));
    jdff dff_B_pQ9JVMvA4_2(.din(n21772), .dout(n21775));
    jdff dff_B_91m689Lr0_2(.din(n21775), .dout(n21778));
    jdff dff_B_FXH8UVvw0_2(.din(n21778), .dout(n21781));
    jdff dff_B_7C8x3nza3_2(.din(n21781), .dout(n21784));
    jdff dff_B_sW6OVQP58_2(.din(n21784), .dout(n21787));
    jdff dff_B_k6h6274F0_2(.din(n21787), .dout(n21790));
    jdff dff_B_eQ2z22vz5_2(.din(n21790), .dout(n21793));
    jdff dff_B_qwQc6bcR9_2(.din(n21793), .dout(n21796));
    jdff dff_B_Pl7K4qeE4_2(.din(n21796), .dout(n21799));
    jdff dff_B_kjwtRpYF9_2(.din(n21799), .dout(n21802));
    jdff dff_B_3rpmHdA50_2(.din(n21802), .dout(n21805));
    jdff dff_B_lmYWVv327_2(.din(n21805), .dout(n21808));
    jdff dff_B_ymBku5oQ0_2(.din(n21808), .dout(n21811));
    jdff dff_B_JAcND1yG6_2(.din(n21811), .dout(n21814));
    jdff dff_B_dGRTS4v79_2(.din(n21814), .dout(n21817));
    jdff dff_B_c8zPlz7S7_2(.din(n21817), .dout(n21820));
    jdff dff_B_WBr45EPs8_2(.din(n21820), .dout(n21823));
    jdff dff_B_6NUDczgV1_2(.din(n21823), .dout(n21826));
    jdff dff_B_9ek3H3DE0_2(.din(n5166), .dout(n21829));
    jdff dff_B_faBXe0Lc1_1(.din(n4965), .dout(n21832));
    jdff dff_B_Zy0EmF5c8_2(.din(n4635), .dout(n21835));
    jdff dff_B_wxkXcXhe5_2(.din(n21835), .dout(n21838));
    jdff dff_B_6UXazMBB8_2(.din(n21838), .dout(n21841));
    jdff dff_B_0OQ4zjqZ5_2(.din(n21841), .dout(n21844));
    jdff dff_B_M37svjXN3_2(.din(n21844), .dout(n21847));
    jdff dff_B_48SDdk871_2(.din(n21847), .dout(n21850));
    jdff dff_B_tDVM4FSx0_2(.din(n21850), .dout(n21853));
    jdff dff_B_RnRX0C9p1_2(.din(n21853), .dout(n21856));
    jdff dff_B_jKbWh6lA2_2(.din(n21856), .dout(n21859));
    jdff dff_B_z1aBQxpj9_2(.din(n21859), .dout(n21862));
    jdff dff_B_zyFaztIQ2_2(.din(n21862), .dout(n21865));
    jdff dff_B_cX9Q2pET6_2(.din(n21865), .dout(n21868));
    jdff dff_B_kHfSLF8B6_2(.din(n21868), .dout(n21871));
    jdff dff_B_D5kFYsyw9_2(.din(n21871), .dout(n21874));
    jdff dff_B_rDwStpPN5_2(.din(n21874), .dout(n21877));
    jdff dff_B_vF3hEizx7_2(.din(n21877), .dout(n21880));
    jdff dff_B_AI8jw5il9_2(.din(n21880), .dout(n21883));
    jdff dff_B_lIeYby8V8_2(.din(n21883), .dout(n21886));
    jdff dff_B_nw4ESBAx9_2(.din(n21886), .dout(n21889));
    jdff dff_B_6qvCuHvB9_2(.din(n21889), .dout(n21892));
    jdff dff_B_bTUEaydP0_2(.din(n21892), .dout(n21895));
    jdff dff_B_9TVk05s40_2(.din(n21895), .dout(n21898));
    jdff dff_B_IMPzkTTk6_2(.din(n21898), .dout(n21901));
    jdff dff_B_IciobQ9S3_2(.din(n21901), .dout(n21904));
    jdff dff_B_olRmnmKX5_2(.din(n21904), .dout(n21907));
    jdff dff_B_D0Fo8iyw5_2(.din(n21907), .dout(n21910));
    jdff dff_B_XZfn5ScZ8_2(.din(n21910), .dout(n21913));
    jdff dff_B_xGr38sAj9_2(.din(n21913), .dout(n21916));
    jdff dff_B_iRazComT1_2(.din(n21916), .dout(n21919));
    jdff dff_B_6LfYAUrp2_2(.din(n21919), .dout(n21922));
    jdff dff_B_tMTFfhlg1_2(.din(n21922), .dout(n21925));
    jdff dff_B_KIPhj9SK0_2(.din(n21925), .dout(n21928));
    jdff dff_B_B4Ub5xnK4_2(.din(n21928), .dout(n21931));
    jdff dff_B_hVnXmHOG6_2(.din(n21931), .dout(n21934));
    jdff dff_B_Szd2QzRz4_2(.din(n21934), .dout(n21937));
    jdff dff_B_wK63IE4k2_2(.din(n21937), .dout(n21940));
    jdff dff_B_cN1DcKVD7_2(.din(n4840), .dout(n21943));
    jdff dff_B_ImpNrGtm4_1(.din(n4639), .dout(n21946));
    jdff dff_B_tupij4Nv5_2(.din(n4289), .dout(n21949));
    jdff dff_B_sHKsTPx80_2(.din(n21949), .dout(n21952));
    jdff dff_B_6vke0d8c0_2(.din(n21952), .dout(n21955));
    jdff dff_B_VLIgPtqg2_2(.din(n21955), .dout(n21958));
    jdff dff_B_yISFIlMI7_2(.din(n21958), .dout(n21961));
    jdff dff_B_vCX7vl4r7_2(.din(n21961), .dout(n21964));
    jdff dff_B_ROeHYyK89_2(.din(n21964), .dout(n21967));
    jdff dff_B_j8JRjkZw1_2(.din(n21967), .dout(n21970));
    jdff dff_B_OWIr4lcW8_2(.din(n21970), .dout(n21973));
    jdff dff_B_ihePhkrq9_2(.din(n21973), .dout(n21976));
    jdff dff_B_GVr11g0U7_2(.din(n21976), .dout(n21979));
    jdff dff_B_TvSbY1429_2(.din(n21979), .dout(n21982));
    jdff dff_B_KPrejBD39_2(.din(n21982), .dout(n21985));
    jdff dff_B_wBdZKpMH2_2(.din(n21985), .dout(n21988));
    jdff dff_B_AvTnVext5_2(.din(n21988), .dout(n21991));
    jdff dff_B_P9gTtpwK6_2(.din(n21991), .dout(n21994));
    jdff dff_B_ov0xG9pm8_2(.din(n21994), .dout(n21997));
    jdff dff_B_VGXCQCUd0_2(.din(n21997), .dout(n22000));
    jdff dff_B_kXYsHOV08_2(.din(n22000), .dout(n22003));
    jdff dff_B_1MMKTMfP2_2(.din(n22003), .dout(n22006));
    jdff dff_B_Of4YOxQd3_2(.din(n22006), .dout(n22009));
    jdff dff_B_4A2sPORL6_2(.din(n22009), .dout(n22012));
    jdff dff_B_fIhypljW9_2(.din(n22012), .dout(n22015));
    jdff dff_B_jWP9SUZ06_2(.din(n22015), .dout(n22018));
    jdff dff_B_D5aerA2U8_2(.din(n22018), .dout(n22021));
    jdff dff_B_CLOCFoYJ4_2(.din(n22021), .dout(n22024));
    jdff dff_B_9hCzTUK42_2(.din(n22024), .dout(n22027));
    jdff dff_B_fFiVH1kG4_2(.din(n22027), .dout(n22030));
    jdff dff_B_FKVraEVe9_2(.din(n22030), .dout(n22033));
    jdff dff_B_r3FGNd2r9_2(.din(n22033), .dout(n22036));
    jdff dff_B_2Xm7Rslv6_2(.din(n22036), .dout(n22039));
    jdff dff_B_HT9VLYAA6_2(.din(n22039), .dout(n22042));
    jdff dff_B_iArFbLF42_2(.din(n22042), .dout(n22045));
    jdff dff_B_X8PXlsSu2_2(.din(n4490), .dout(n22048));
    jdff dff_B_0sSPHn4O8_1(.din(n4293), .dout(n22051));
    jdff dff_B_c3Vd6GrN3_2(.din(n3893), .dout(n22054));
    jdff dff_B_lf3zomKh8_2(.din(n22054), .dout(n22057));
    jdff dff_B_FqoalI5p1_2(.din(n22057), .dout(n22060));
    jdff dff_B_BUS2HOza9_2(.din(n22060), .dout(n22063));
    jdff dff_B_NqlTAb3O0_2(.din(n22063), .dout(n22066));
    jdff dff_B_aJA2haG50_2(.din(n22066), .dout(n22069));
    jdff dff_B_MXv2KJ0H9_2(.din(n22069), .dout(n22072));
    jdff dff_B_5dIt3qRJ9_2(.din(n22072), .dout(n22075));
    jdff dff_B_tzWFpcnl3_2(.din(n22075), .dout(n22078));
    jdff dff_B_UE1XYbw51_2(.din(n22078), .dout(n22081));
    jdff dff_B_M4LX79iD3_2(.din(n22081), .dout(n22084));
    jdff dff_B_pMOogKxM1_2(.din(n22084), .dout(n22087));
    jdff dff_B_jQLXLeSi6_2(.din(n22087), .dout(n22090));
    jdff dff_B_m0zmUcfS8_2(.din(n22090), .dout(n22093));
    jdff dff_B_Umklu2qo4_2(.din(n22093), .dout(n22096));
    jdff dff_B_iIqrvonK1_2(.din(n22096), .dout(n22099));
    jdff dff_B_pRCVsK5J0_2(.din(n22099), .dout(n22102));
    jdff dff_B_FNJztTfC8_2(.din(n22102), .dout(n22105));
    jdff dff_B_prQxtbgJ4_2(.din(n22105), .dout(n22108));
    jdff dff_B_EyfdXWdF9_2(.din(n22108), .dout(n22111));
    jdff dff_B_MLxzRiDT8_2(.din(n22111), .dout(n22114));
    jdff dff_B_Scpb4JCl2_2(.din(n22114), .dout(n22117));
    jdff dff_B_al9HdKIK0_2(.din(n22117), .dout(n22120));
    jdff dff_B_JbQX7Hbj0_2(.din(n22120), .dout(n22123));
    jdff dff_B_BhDPqHiN3_2(.din(n22123), .dout(n22126));
    jdff dff_B_KCug5COe5_2(.din(n22126), .dout(n22129));
    jdff dff_B_vf3dco6h5_2(.din(n22129), .dout(n22132));
    jdff dff_B_MlpgTR5Q3_2(.din(n22132), .dout(n22135));
    jdff dff_B_MjcPfnJp5_2(.din(n22135), .dout(n22138));
    jdff dff_B_tE3GPyAT6_2(.din(n22138), .dout(n22141));
    jdff dff_B_Ey1mCoSe0_2(.din(n4114), .dout(n22144));
    jdff dff_B_EU9fSBA64_1(.din(n3897), .dout(n22147));
    jdff dff_B_msWHd3oh5_2(.din(n3516), .dout(n22150));
    jdff dff_B_Neyv2mKd0_2(.din(n22150), .dout(n22153));
    jdff dff_B_R6CN6o1L5_2(.din(n22153), .dout(n22156));
    jdff dff_B_qzQiVGiQ8_2(.din(n22156), .dout(n22159));
    jdff dff_B_EKLGHIcV9_2(.din(n22159), .dout(n22162));
    jdff dff_B_plfNoSIO3_2(.din(n22162), .dout(n22165));
    jdff dff_B_1twOcQB14_2(.din(n22165), .dout(n22168));
    jdff dff_B_DOMXe3GP5_2(.din(n22168), .dout(n22171));
    jdff dff_B_BPq00AG38_2(.din(n22171), .dout(n22174));
    jdff dff_B_OwlEvNCk5_2(.din(n22174), .dout(n22177));
    jdff dff_B_9691XIaT6_2(.din(n22177), .dout(n22180));
    jdff dff_B_Evd8MDCF3_2(.din(n22180), .dout(n22183));
    jdff dff_B_EWB6sXBG3_2(.din(n22183), .dout(n22186));
    jdff dff_B_7kx7y9Xv3_2(.din(n22186), .dout(n22189));
    jdff dff_B_7YH5rV9f4_2(.din(n22189), .dout(n22192));
    jdff dff_B_ol5XeFAm4_2(.din(n22192), .dout(n22195));
    jdff dff_B_nxNUkvJm1_2(.din(n22195), .dout(n22198));
    jdff dff_B_HHso2Rpj0_2(.din(n22198), .dout(n22201));
    jdff dff_B_W0w5z7bF8_2(.din(n22201), .dout(n22204));
    jdff dff_B_jTzzGAYl7_2(.din(n22204), .dout(n22207));
    jdff dff_B_Xuak1bne9_2(.din(n22207), .dout(n22210));
    jdff dff_B_Y4K0I4uD3_2(.din(n22210), .dout(n22213));
    jdff dff_B_vYRFEYbL2_2(.din(n22213), .dout(n22216));
    jdff dff_B_IpURNv8y7_2(.din(n22216), .dout(n22219));
    jdff dff_B_P3FSdtuF0_2(.din(n22219), .dout(n22222));
    jdff dff_B_6GbxEZyg9_2(.din(n22222), .dout(n22225));
    jdff dff_B_9B0pqAp15_2(.din(n22225), .dout(n22228));
    jdff dff_B_odIEMLG73_2(.din(n3711), .dout(n22231));
    jdff dff_B_P00V99xF6_1(.din(n3520), .dout(n22234));
    jdff dff_B_WJAPKH9r4_2(.din(n3115), .dout(n22237));
    jdff dff_B_Be2y1eLw1_2(.din(n22237), .dout(n22240));
    jdff dff_B_PP4BbTAx4_2(.din(n22240), .dout(n22243));
    jdff dff_B_knzvl6E08_2(.din(n22243), .dout(n22246));
    jdff dff_B_4SrQ0URV1_2(.din(n22246), .dout(n22249));
    jdff dff_B_yAIpMIn73_2(.din(n22249), .dout(n22252));
    jdff dff_B_UfsHC1C33_2(.din(n22252), .dout(n22255));
    jdff dff_B_5deEPxUu2_2(.din(n22255), .dout(n22258));
    jdff dff_B_ZQlbNdte0_2(.din(n22258), .dout(n22261));
    jdff dff_B_8ganj8Pt3_2(.din(n22261), .dout(n22264));
    jdff dff_B_wLDMP53B3_2(.din(n22264), .dout(n22267));
    jdff dff_B_QC9oHw9t2_2(.din(n22267), .dout(n22270));
    jdff dff_B_tkkr1hc26_2(.din(n22270), .dout(n22273));
    jdff dff_B_PBbUxTOK4_2(.din(n22273), .dout(n22276));
    jdff dff_B_GheVLLBZ8_2(.din(n22276), .dout(n22279));
    jdff dff_B_ygMLiikt8_2(.din(n22279), .dout(n22282));
    jdff dff_B_q5NYwUsE9_2(.din(n22282), .dout(n22285));
    jdff dff_B_3uzTq3Az3_2(.din(n22285), .dout(n22288));
    jdff dff_B_Rjet8Wn75_2(.din(n22288), .dout(n22291));
    jdff dff_B_J1iPLDCX0_2(.din(n22291), .dout(n22294));
    jdff dff_B_eF9Tk66p4_2(.din(n22294), .dout(n22297));
    jdff dff_B_47ZRFloy8_2(.din(n22297), .dout(n22300));
    jdff dff_B_H2RfDcbU6_2(.din(n22300), .dout(n22303));
    jdff dff_B_W4fjIvWG8_2(.din(n22303), .dout(n22306));
    jdff dff_B_SqSzmfJI2_2(.din(n3309), .dout(n22309));
    jdff dff_B_FwUjwLpg3_1(.din(n3119), .dout(n22312));
    jdff dff_B_sbiRgiuq9_2(.din(n2736), .dout(n22315));
    jdff dff_B_2qFNidnc3_2(.din(n22315), .dout(n22318));
    jdff dff_B_s8IYWgUJ6_2(.din(n22318), .dout(n22321));
    jdff dff_B_bfVDU8DR9_2(.din(n22321), .dout(n22324));
    jdff dff_B_Zsg35E7T0_2(.din(n22324), .dout(n22327));
    jdff dff_B_NIuS8Gao2_2(.din(n22327), .dout(n22330));
    jdff dff_B_2R3SzqrG6_2(.din(n22330), .dout(n22333));
    jdff dff_B_RnlveGLs4_2(.din(n22333), .dout(n22336));
    jdff dff_B_yKvtNNbC3_2(.din(n22336), .dout(n22339));
    jdff dff_B_nJLfIOD81_2(.din(n22339), .dout(n22342));
    jdff dff_B_XJEfy2eA2_2(.din(n22342), .dout(n22345));
    jdff dff_B_MjUiPWYF1_2(.din(n22345), .dout(n22348));
    jdff dff_B_2xI6hlF41_2(.din(n22348), .dout(n22351));
    jdff dff_B_rSF8CSo16_2(.din(n22351), .dout(n22354));
    jdff dff_B_W0mRZfbF5_2(.din(n22354), .dout(n22357));
    jdff dff_B_B6eRyLYW2_2(.din(n22357), .dout(n22360));
    jdff dff_B_kEoxd8r45_2(.din(n22360), .dout(n22363));
    jdff dff_B_DNoRZaMs0_2(.din(n22363), .dout(n22366));
    jdff dff_B_amQhJ1rp8_2(.din(n22366), .dout(n22369));
    jdff dff_B_hfBLVgxm8_2(.din(n22369), .dout(n22372));
    jdff dff_B_NJq9Mwmv8_2(.din(n22372), .dout(n22375));
    jdff dff_B_9rJcZFO74_2(.din(n2904), .dout(n22378));
    jdff dff_B_aLCONApw9_1(.din(n2740), .dout(n22381));
    jdff dff_B_eTKLcG3n9_2(.din(n2381), .dout(n22384));
    jdff dff_B_R6UHHqcU8_2(.din(n22384), .dout(n22387));
    jdff dff_B_hXhFr7N95_2(.din(n22387), .dout(n22390));
    jdff dff_B_NRLcLJR19_2(.din(n22390), .dout(n22393));
    jdff dff_B_dUEnkPYr7_2(.din(n22393), .dout(n22396));
    jdff dff_B_XLvcjCws7_2(.din(n22396), .dout(n22399));
    jdff dff_B_icyC7InA1_2(.din(n22399), .dout(n22402));
    jdff dff_B_Uqk8bYov4_2(.din(n22402), .dout(n22405));
    jdff dff_B_MpLiHoPy2_2(.din(n22405), .dout(n22408));
    jdff dff_B_F2gVclQR0_2(.din(n22408), .dout(n22411));
    jdff dff_B_DQ9DLNxE3_2(.din(n22411), .dout(n22414));
    jdff dff_B_F6QBbcuy4_2(.din(n22414), .dout(n22417));
    jdff dff_B_QjgN8iEH3_2(.din(n22417), .dout(n22420));
    jdff dff_B_7TsXYrYs6_2(.din(n22420), .dout(n22423));
    jdff dff_B_azhVPQdI9_2(.din(n22423), .dout(n22426));
    jdff dff_B_hbH2dvgo3_2(.din(n22426), .dout(n22429));
    jdff dff_B_9lYNUB6v6_2(.din(n22429), .dout(n22432));
    jdff dff_B_sWjd90256_2(.din(n22432), .dout(n22435));
    jdff dff_B_RHR0rDDN0_2(.din(n2522), .dout(n22438));
    jdff dff_B_myZc1rch3_1(.din(n2385), .dout(n22441));
    jdff dff_B_Wk0729rd9_2(.din(n2053), .dout(n22444));
    jdff dff_B_9j2TjyNq2_2(.din(n22444), .dout(n22447));
    jdff dff_B_0zH9w3kZ5_2(.din(n22447), .dout(n22450));
    jdff dff_B_hzUDXxsE8_2(.din(n22450), .dout(n22453));
    jdff dff_B_fDnBT49Y9_2(.din(n22453), .dout(n22456));
    jdff dff_B_AVfeqjyG7_2(.din(n22456), .dout(n22459));
    jdff dff_B_4BuUGYnX4_2(.din(n22459), .dout(n22462));
    jdff dff_B_mtqPUI0T1_2(.din(n22462), .dout(n22465));
    jdff dff_B_Mpp5fT8p6_2(.din(n22465), .dout(n22468));
    jdff dff_B_TViT5sPd4_2(.din(n22468), .dout(n22471));
    jdff dff_B_eQU8pXQN6_2(.din(n22471), .dout(n22474));
    jdff dff_B_hB9y8UTf7_2(.din(n22474), .dout(n22477));
    jdff dff_B_8lRcB4fm6_2(.din(n22477), .dout(n22480));
    jdff dff_B_aXuJiYt90_2(.din(n22480), .dout(n22483));
    jdff dff_B_N4qhkeI07_2(.din(n22483), .dout(n22486));
    jdff dff_B_rldC3BJ47_2(.din(n2167), .dout(n22489));
    jdff dff_B_JXDGhtOe4_1(.din(n2057), .dout(n22492));
    jdff dff_B_2RydlANO8_2(.din(n1752), .dout(n22495));
    jdff dff_B_CIScbIBQ6_2(.din(n22495), .dout(n22498));
    jdff dff_B_zH8a4xVO4_2(.din(n22498), .dout(n22501));
    jdff dff_B_sDahNV6J7_2(.din(n22501), .dout(n22504));
    jdff dff_B_94Su4Wyr7_2(.din(n22504), .dout(n22507));
    jdff dff_B_RRUJDn0M0_2(.din(n22507), .dout(n22510));
    jdff dff_B_PC0IDieh3_2(.din(n22510), .dout(n22513));
    jdff dff_B_Hd6Dvm0S6_2(.din(n22513), .dout(n22516));
    jdff dff_B_vnDs6X5n0_2(.din(n22516), .dout(n22519));
    jdff dff_B_SpKWs8qL6_2(.din(n22519), .dout(n22522));
    jdff dff_B_deIYh7Pd5_2(.din(n22522), .dout(n22525));
    jdff dff_B_StDSFw8h8_2(.din(n22525), .dout(n22528));
    jdff dff_B_CVnLg0kR4_2(.din(n1839), .dout(n22531));
    jdff dff_B_fr234X5Q7_1(.din(n1756), .dout(n22534));
    jdff dff_B_6tT9T7Su6_2(.din(n1478), .dout(n22537));
    jdff dff_B_Wqu20p4v5_2(.din(n22537), .dout(n22540));
    jdff dff_B_A8a4HFKX5_2(.din(n22540), .dout(n22543));
    jdff dff_B_nnvA88J42_2(.din(n22543), .dout(n22546));
    jdff dff_B_48uXmbWc9_2(.din(n22546), .dout(n22549));
    jdff dff_B_8H9EKZis3_2(.din(n22549), .dout(n22552));
    jdff dff_B_hIDVNv4n8_2(.din(n22552), .dout(n22555));
    jdff dff_B_wmccnfO15_2(.din(n22555), .dout(n22558));
    jdff dff_B_j23U0sOR6_2(.din(n22558), .dout(n22561));
    jdff dff_B_DENUeDNg6_2(.din(n1538), .dout(n22564));
    jdff dff_B_ugK7QYqi7_2(.din(n22564), .dout(n22567));
    jdff dff_B_MYapCTdd2_1(.din(n1481), .dout(n22570));
    jdff dff_B_xgmph9Mx5_1(.din(n22570), .dout(n22573));
    jdff dff_B_9kdLMMw17_1(.din(n22573), .dout(n22576));
    jdff dff_B_ou4UUd8m9_1(.din(n22576), .dout(n22579));
    jdff dff_B_Eg0G2rQK4_1(.din(n22579), .dout(n22582));
    jdff dff_B_zin7EFie7_1(.din(n22582), .dout(n22585));
    jdff dff_B_ayM6OZZT9_0(.din(n1264), .dout(n22588));
    jdff dff_B_L41QrBO30_0(.din(n22588), .dout(n22591));
    jdff dff_A_TmYr42cC0_0(.din(n22596), .dout(n22593));
    jdff dff_A_v2T2r6Bw5_0(.din(n22599), .dout(n22596));
    jdff dff_A_CFnGIAnQ4_0(.din(n1260), .dout(n22599));
    jdff dff_B_AuDEaiwK0_1(.din(n1238), .dout(n22603));
    jdff dff_A_CWv4PehF4_0(.din(n1010), .dout(n22605));
    jdff dff_A_PldyxTtr0_1(.din(n22611), .dout(n22608));
    jdff dff_A_IQZnHAAl3_1(.din(n1010), .dout(n22611));
    jdff dff_A_jlCOkuN10_1(.din(n22617), .dout(n22614));
    jdff dff_A_Vzuu0Vkz3_1(.din(n22620), .dout(n22617));
    jdff dff_A_5iOY39rK3_1(.din(n22623), .dout(n22620));
    jdff dff_A_fYxLTpdA0_1(.din(n22626), .dout(n22623));
    jdff dff_A_vkF2PkVD2_1(.din(n22629), .dout(n22626));
    jdff dff_A_AlngDwTI8_1(.din(n1230), .dout(n22629));
    jdff dff_B_tmATA0839_2(.din(n6029), .dout(n22633));
    jdff dff_B_qO9LQxKl1_2(.din(n22633), .dout(n22636));
    jdff dff_B_mP2VrqKQ6_1(.din(n6021), .dout(n22639));
    jdff dff_B_plqLQFNf4_2(.din(n5796), .dout(n22642));
    jdff dff_B_FSU4Fl4o1_2(.din(n22642), .dout(n22645));
    jdff dff_B_YCffW1NN1_2(.din(n22645), .dout(n22648));
    jdff dff_B_tnMY8Ikd0_2(.din(n22648), .dout(n22651));
    jdff dff_B_aRbZ0vuq7_2(.din(n22651), .dout(n22654));
    jdff dff_B_XjtbQkA16_2(.din(n22654), .dout(n22657));
    jdff dff_B_SZmuMXNF5_2(.din(n22657), .dout(n22660));
    jdff dff_B_8NpBifyg5_2(.din(n22660), .dout(n22663));
    jdff dff_B_EmYtTHYT5_2(.din(n22663), .dout(n22666));
    jdff dff_B_QWZjE07A5_2(.din(n22666), .dout(n22669));
    jdff dff_B_48xUDhoj6_2(.din(n22669), .dout(n22672));
    jdff dff_B_Yh5tGfSY6_2(.din(n22672), .dout(n22675));
    jdff dff_B_z2ELHyry4_2(.din(n22675), .dout(n22678));
    jdff dff_B_qW6Bg2YV3_2(.din(n22678), .dout(n22681));
    jdff dff_B_t36SaB8O2_2(.din(n22681), .dout(n22684));
    jdff dff_B_RKhaZqiF6_2(.din(n22684), .dout(n22687));
    jdff dff_B_knm0k8Xg4_2(.din(n22687), .dout(n22690));
    jdff dff_B_yEHtgwAw9_2(.din(n22690), .dout(n22693));
    jdff dff_B_CBPGj1Xr9_2(.din(n22693), .dout(n22696));
    jdff dff_B_wfNlrhA39_2(.din(n22696), .dout(n22699));
    jdff dff_B_XZWc1MA07_2(.din(n22699), .dout(n22702));
    jdff dff_B_tjYOlqZm1_2(.din(n22702), .dout(n22705));
    jdff dff_B_hELfrm557_2(.din(n22705), .dout(n22708));
    jdff dff_B_EeHt7nf20_2(.din(n22708), .dout(n22711));
    jdff dff_B_PUVktDH65_2(.din(n22711), .dout(n22714));
    jdff dff_B_e8tfmy4u5_2(.din(n22714), .dout(n22717));
    jdff dff_B_DE1T8EcF2_2(.din(n22717), .dout(n22720));
    jdff dff_B_DbnIVGSV5_2(.din(n22720), .dout(n22723));
    jdff dff_B_Semw6xyf3_2(.din(n22723), .dout(n22726));
    jdff dff_B_6HL6TPZi0_2(.din(n22726), .dout(n22729));
    jdff dff_B_dKWFuJb32_2(.din(n22729), .dout(n22732));
    jdff dff_B_tQwvjZBp2_2(.din(n22732), .dout(n22735));
    jdff dff_B_O3rmj7Hd0_2(.din(n22735), .dout(n22738));
    jdff dff_B_bSnaak8k2_2(.din(n22738), .dout(n22741));
    jdff dff_B_C3SRLnC69_2(.din(n22741), .dout(n22744));
    jdff dff_B_70Xy8b0j3_2(.din(n22744), .dout(n22747));
    jdff dff_B_zmavL6419_2(.din(n22747), .dout(n22750));
    jdff dff_B_0wlAA0ud1_2(.din(n22750), .dout(n22753));
    jdff dff_B_ow3Kdl3O0_2(.din(n22753), .dout(n22756));
    jdff dff_B_IXcVz9od3_2(.din(n22756), .dout(n22759));
    jdff dff_B_UIupoNSA5_2(.din(n22759), .dout(n22762));
    jdff dff_B_IxFvomfa6_2(.din(n22762), .dout(n22765));
    jdff dff_B_uivDMDmA9_2(.din(n22765), .dout(n22768));
    jdff dff_B_vJbzwzhe9_2(.din(n22768), .dout(n22771));
    jdff dff_B_y9QMcpst5_2(.din(n22771), .dout(n22774));
    jdff dff_B_KEC61UbN7_2(.din(n22774), .dout(n22777));
    jdff dff_B_4gjy0nN20_2(.din(n22777), .dout(n22780));
    jdff dff_B_ewia6aDz7_1(.din(n5800), .dout(n22783));
    jdff dff_B_SPXqW2dm1_2(.din(n5551), .dout(n22786));
    jdff dff_B_kTykYwNQ1_2(.din(n22786), .dout(n22789));
    jdff dff_B_OC4OnPtO3_2(.din(n22789), .dout(n22792));
    jdff dff_B_H1ekknui1_2(.din(n22792), .dout(n22795));
    jdff dff_B_ey9eU7cV7_2(.din(n22795), .dout(n22798));
    jdff dff_B_n7EoCFBQ3_2(.din(n22798), .dout(n22801));
    jdff dff_B_msYtl1oB4_2(.din(n22801), .dout(n22804));
    jdff dff_B_DhnOhXgm6_2(.din(n22804), .dout(n22807));
    jdff dff_B_hPp4pb6m3_2(.din(n22807), .dout(n22810));
    jdff dff_B_NcOOZW1C0_2(.din(n22810), .dout(n22813));
    jdff dff_B_H9TtCYDc6_2(.din(n22813), .dout(n22816));
    jdff dff_B_04DJ5N5p2_2(.din(n22816), .dout(n22819));
    jdff dff_B_1VzuVgi55_2(.din(n22819), .dout(n22822));
    jdff dff_B_jI0d8bc10_2(.din(n22822), .dout(n22825));
    jdff dff_B_W0I0efQf8_2(.din(n22825), .dout(n22828));
    jdff dff_B_w8oH05OQ2_2(.din(n22828), .dout(n22831));
    jdff dff_B_DCvcBuH23_2(.din(n22831), .dout(n22834));
    jdff dff_B_PQ9kNBfv0_2(.din(n22834), .dout(n22837));
    jdff dff_B_02MewigC3_2(.din(n22837), .dout(n22840));
    jdff dff_B_567YfJb48_2(.din(n22840), .dout(n22843));
    jdff dff_B_mv94IPBP5_2(.din(n22843), .dout(n22846));
    jdff dff_B_Rvyk1bc65_2(.din(n22846), .dout(n22849));
    jdff dff_B_u2ZuBt3E8_2(.din(n22849), .dout(n22852));
    jdff dff_B_4WU0sOu84_2(.din(n22852), .dout(n22855));
    jdff dff_B_nltW59Ju1_2(.din(n22855), .dout(n22858));
    jdff dff_B_1ZNXYIwD0_2(.din(n22858), .dout(n22861));
    jdff dff_B_o7z3vP909_2(.din(n22861), .dout(n22864));
    jdff dff_B_pZPftn4o4_2(.din(n22864), .dout(n22867));
    jdff dff_B_nROt5SIt4_2(.din(n22867), .dout(n22870));
    jdff dff_B_ivCzFx8c8_2(.din(n22870), .dout(n22873));
    jdff dff_B_D8shVlpO4_2(.din(n22873), .dout(n22876));
    jdff dff_B_HAGUHgsz6_2(.din(n22876), .dout(n22879));
    jdff dff_B_ASSS5cmR7_2(.din(n22879), .dout(n22882));
    jdff dff_B_B8QSHjaK1_2(.din(n22882), .dout(n22885));
    jdff dff_B_pBJ2Dndp1_2(.din(n22885), .dout(n22888));
    jdff dff_B_TnpgL7Sz4_2(.din(n22888), .dout(n22891));
    jdff dff_B_ZFryTQeT9_2(.din(n22891), .dout(n22894));
    jdff dff_B_vpmIoObM3_2(.din(n22894), .dout(n22897));
    jdff dff_B_7lS39wSh8_2(.din(n22897), .dout(n22900));
    jdff dff_B_t4TYKUIV5_2(.din(n22900), .dout(n22903));
    jdff dff_B_rG0GDWV04_2(.din(n22903), .dout(n22906));
    jdff dff_B_2Dc2Cqqv3_2(.din(n22906), .dout(n22909));
    jdff dff_B_DhnMH88a8_2(.din(n5729), .dout(n22912));
    jdff dff_B_t36JFZHW4_1(.din(n5555), .dout(n22915));
    jdff dff_B_W2D9LgdN6_2(.din(n5279), .dout(n22918));
    jdff dff_B_0WMAt5ZJ9_2(.din(n22918), .dout(n22921));
    jdff dff_B_27gtSKIT6_2(.din(n22921), .dout(n22924));
    jdff dff_B_2yeudNdz7_2(.din(n22924), .dout(n22927));
    jdff dff_B_mH2dwj8j0_2(.din(n22927), .dout(n22930));
    jdff dff_B_4ykKdkSo1_2(.din(n22930), .dout(n22933));
    jdff dff_B_YQPuyVSy9_2(.din(n22933), .dout(n22936));
    jdff dff_B_vRmFT9vW7_2(.din(n22936), .dout(n22939));
    jdff dff_B_AQ32ZqUO8_2(.din(n22939), .dout(n22942));
    jdff dff_B_NAzTCZhW0_2(.din(n22942), .dout(n22945));
    jdff dff_B_Xw5Zjdo61_2(.din(n22945), .dout(n22948));
    jdff dff_B_aHC6WF8t9_2(.din(n22948), .dout(n22951));
    jdff dff_B_hsBo7oyx7_2(.din(n22951), .dout(n22954));
    jdff dff_B_vl4HxP8H4_2(.din(n22954), .dout(n22957));
    jdff dff_B_AZ8Uq0Je9_2(.din(n22957), .dout(n22960));
    jdff dff_B_c77SKypD8_2(.din(n22960), .dout(n22963));
    jdff dff_B_4J9yUMTh4_2(.din(n22963), .dout(n22966));
    jdff dff_B_Kc4qZdze1_2(.din(n22966), .dout(n22969));
    jdff dff_B_FUUV2IFK0_2(.din(n22969), .dout(n22972));
    jdff dff_B_4IaHg2y39_2(.din(n22972), .dout(n22975));
    jdff dff_B_tSxKbDZx9_2(.din(n22975), .dout(n22978));
    jdff dff_B_XsHjt4T17_2(.din(n22978), .dout(n22981));
    jdff dff_B_zgWTXqDe3_2(.din(n22981), .dout(n22984));
    jdff dff_B_aQLIWByr2_2(.din(n22984), .dout(n22987));
    jdff dff_B_vjhBhKZL7_2(.din(n22987), .dout(n22990));
    jdff dff_B_15SdAugp4_2(.din(n22990), .dout(n22993));
    jdff dff_B_eZaSc35B2_2(.din(n22993), .dout(n22996));
    jdff dff_B_s0s7SrLJ2_2(.din(n22996), .dout(n22999));
    jdff dff_B_Pf8NYs0X7_2(.din(n22999), .dout(n23002));
    jdff dff_B_JS6VDofc4_2(.din(n23002), .dout(n23005));
    jdff dff_B_MxlpbtEz8_2(.din(n23005), .dout(n23008));
    jdff dff_B_ryAZhdJc6_2(.din(n23008), .dout(n23011));
    jdff dff_B_T8fmoYTS6_2(.din(n23011), .dout(n23014));
    jdff dff_B_XVlVHmCQ4_2(.din(n23014), .dout(n23017));
    jdff dff_B_RNOVQFcl9_2(.din(n23017), .dout(n23020));
    jdff dff_B_dgOO3eT99_2(.din(n23020), .dout(n23023));
    jdff dff_B_cHGSWxIC0_2(.din(n23023), .dout(n23026));
    jdff dff_B_p9L3JcAh3_2(.din(n23026), .dout(n23029));
    jdff dff_B_Gzmv50DE8_2(.din(n23029), .dout(n23032));
    jdff dff_B_A3R2VAa63_2(.din(n5457), .dout(n23035));
    jdff dff_B_NTWXxtiL6_1(.din(n5283), .dout(n23038));
    jdff dff_B_RNJJNCz87_2(.din(n4980), .dout(n23041));
    jdff dff_B_Ao0pvMLT7_2(.din(n23041), .dout(n23044));
    jdff dff_B_m5IhTBR80_2(.din(n23044), .dout(n23047));
    jdff dff_B_Fv0nOfa90_2(.din(n23047), .dout(n23050));
    jdff dff_B_rkybG2kM7_2(.din(n23050), .dout(n23053));
    jdff dff_B_l6mnBk3Z3_2(.din(n23053), .dout(n23056));
    jdff dff_B_WTfkTDFu1_2(.din(n23056), .dout(n23059));
    jdff dff_B_8PNFX68G2_2(.din(n23059), .dout(n23062));
    jdff dff_B_237ECkMK0_2(.din(n23062), .dout(n23065));
    jdff dff_B_iMGYnLzT3_2(.din(n23065), .dout(n23068));
    jdff dff_B_WUTQDFVG2_2(.din(n23068), .dout(n23071));
    jdff dff_B_ZjXT7OBx5_2(.din(n23071), .dout(n23074));
    jdff dff_B_kAhla4n08_2(.din(n23074), .dout(n23077));
    jdff dff_B_tomTPd9y1_2(.din(n23077), .dout(n23080));
    jdff dff_B_CfCdbbvS2_2(.din(n23080), .dout(n23083));
    jdff dff_B_3OUYU2I74_2(.din(n23083), .dout(n23086));
    jdff dff_B_pbxAkWNd0_2(.din(n23086), .dout(n23089));
    jdff dff_B_R5nBeBZ59_2(.din(n23089), .dout(n23092));
    jdff dff_B_QNOqrJ0A8_2(.din(n23092), .dout(n23095));
    jdff dff_B_MoKvDhTo5_2(.din(n23095), .dout(n23098));
    jdff dff_B_J7i9nfDu3_2(.din(n23098), .dout(n23101));
    jdff dff_B_TobCk7kL6_2(.din(n23101), .dout(n23104));
    jdff dff_B_xcs9joq36_2(.din(n23104), .dout(n23107));
    jdff dff_B_ZVqcZxM41_2(.din(n23107), .dout(n23110));
    jdff dff_B_P4niPtod4_2(.din(n23110), .dout(n23113));
    jdff dff_B_v92yHpEa5_2(.din(n23113), .dout(n23116));
    jdff dff_B_kfOIsyGW9_2(.din(n23116), .dout(n23119));
    jdff dff_B_1LofYttv4_2(.din(n23119), .dout(n23122));
    jdff dff_B_qrJBSzC89_2(.din(n23122), .dout(n23125));
    jdff dff_B_PB6FJwQ53_2(.din(n23125), .dout(n23128));
    jdff dff_B_MwzE1mE58_2(.din(n23128), .dout(n23131));
    jdff dff_B_7BAifTpZ3_2(.din(n23131), .dout(n23134));
    jdff dff_B_eRUPqLDn5_2(.din(n23134), .dout(n23137));
    jdff dff_B_gEpaOo1z1_2(.din(n23137), .dout(n23140));
    jdff dff_B_vJylCD1i2_2(.din(n23140), .dout(n23143));
    jdff dff_B_aVwQOu5d0_2(.din(n23143), .dout(n23146));
    jdff dff_B_1ibA4IKY8_2(.din(n5158), .dout(n23149));
    jdff dff_B_sP4Ejq843_1(.din(n4984), .dout(n23152));
    jdff dff_B_UPfBcQpT9_2(.din(n4654), .dout(n23155));
    jdff dff_B_Z5Iv1g5Q9_2(.din(n23155), .dout(n23158));
    jdff dff_B_jdLlyNxj6_2(.din(n23158), .dout(n23161));
    jdff dff_B_G4MVYnug1_2(.din(n23161), .dout(n23164));
    jdff dff_B_J4zpvQO48_2(.din(n23164), .dout(n23167));
    jdff dff_B_iXrriSKA5_2(.din(n23167), .dout(n23170));
    jdff dff_B_IML1f4pw4_2(.din(n23170), .dout(n23173));
    jdff dff_B_RCo6VYIV9_2(.din(n23173), .dout(n23176));
    jdff dff_B_Y0hH1vEO4_2(.din(n23176), .dout(n23179));
    jdff dff_B_nzvBuzoc2_2(.din(n23179), .dout(n23182));
    jdff dff_B_YeruEgU76_2(.din(n23182), .dout(n23185));
    jdff dff_B_LeEsOAyE2_2(.din(n23185), .dout(n23188));
    jdff dff_B_64IjW4vJ1_2(.din(n23188), .dout(n23191));
    jdff dff_B_sAwzFx3z9_2(.din(n23191), .dout(n23194));
    jdff dff_B_eP4KJ1Ce8_2(.din(n23194), .dout(n23197));
    jdff dff_B_cycacQty7_2(.din(n23197), .dout(n23200));
    jdff dff_B_C3SbwQnh2_2(.din(n23200), .dout(n23203));
    jdff dff_B_Eyqr2xo32_2(.din(n23203), .dout(n23206));
    jdff dff_B_HLctiEbA8_2(.din(n23206), .dout(n23209));
    jdff dff_B_EEFVhxNg0_2(.din(n23209), .dout(n23212));
    jdff dff_B_LOoSonQp4_2(.din(n23212), .dout(n23215));
    jdff dff_B_djsuKSzd7_2(.din(n23215), .dout(n23218));
    jdff dff_B_ZOROOSvj7_2(.din(n23218), .dout(n23221));
    jdff dff_B_95KqB4Id8_2(.din(n23221), .dout(n23224));
    jdff dff_B_KVdZoxK02_2(.din(n23224), .dout(n23227));
    jdff dff_B_LcUsYLLa3_2(.din(n23227), .dout(n23230));
    jdff dff_B_dFmMhxME2_2(.din(n23230), .dout(n23233));
    jdff dff_B_G4v4cB765_2(.din(n23233), .dout(n23236));
    jdff dff_B_txscnVFt6_2(.din(n23236), .dout(n23239));
    jdff dff_B_b0KI3EAq2_2(.din(n23239), .dout(n23242));
    jdff dff_B_5ndnb7647_2(.din(n23242), .dout(n23245));
    jdff dff_B_xTxfJX3d8_2(.din(n23245), .dout(n23248));
    jdff dff_B_7R0lN1O60_2(.din(n23248), .dout(n23251));
    jdff dff_B_gBIJsM8w9_2(.din(n4832), .dout(n23254));
    jdff dff_B_OV7ggkl04_1(.din(n4658), .dout(n23257));
    jdff dff_B_q7OUFDbZ9_2(.din(n4308), .dout(n23260));
    jdff dff_B_EdsKtupo0_2(.din(n23260), .dout(n23263));
    jdff dff_B_bbHw0lxs0_2(.din(n23263), .dout(n23266));
    jdff dff_B_Nj5M3Epq0_2(.din(n23266), .dout(n23269));
    jdff dff_B_oaFW9q362_2(.din(n23269), .dout(n23272));
    jdff dff_B_Gp1rMAbZ4_2(.din(n23272), .dout(n23275));
    jdff dff_B_tOq3sVn01_2(.din(n23275), .dout(n23278));
    jdff dff_B_o67CCh235_2(.din(n23278), .dout(n23281));
    jdff dff_B_MzV4yTXU7_2(.din(n23281), .dout(n23284));
    jdff dff_B_74rA2ppH0_2(.din(n23284), .dout(n23287));
    jdff dff_B_Aovb1Zli7_2(.din(n23287), .dout(n23290));
    jdff dff_B_T6WNXiWJ1_2(.din(n23290), .dout(n23293));
    jdff dff_B_RscgG0iQ7_2(.din(n23293), .dout(n23296));
    jdff dff_B_JnOtgfc76_2(.din(n23296), .dout(n23299));
    jdff dff_B_IxwqDl0d7_2(.din(n23299), .dout(n23302));
    jdff dff_B_8hqdvpSS9_2(.din(n23302), .dout(n23305));
    jdff dff_B_PeXW10J35_2(.din(n23305), .dout(n23308));
    jdff dff_B_9dZ3Len40_2(.din(n23308), .dout(n23311));
    jdff dff_B_5xM2FZkd0_2(.din(n23311), .dout(n23314));
    jdff dff_B_E1Fw6C7v8_2(.din(n23314), .dout(n23317));
    jdff dff_B_7Q8qCMYt1_2(.din(n23317), .dout(n23320));
    jdff dff_B_p90lf7R15_2(.din(n23320), .dout(n23323));
    jdff dff_B_zHe1xKuS3_2(.din(n23323), .dout(n23326));
    jdff dff_B_8ojM9xyx8_2(.din(n23326), .dout(n23329));
    jdff dff_B_rjS4bj6V0_2(.din(n23329), .dout(n23332));
    jdff dff_B_aruJWUHh6_2(.din(n23332), .dout(n23335));
    jdff dff_B_Y0cRz4VG2_2(.din(n23335), .dout(n23338));
    jdff dff_B_MhuYKNBv9_2(.din(n23338), .dout(n23341));
    jdff dff_B_EhXr46m92_2(.din(n23341), .dout(n23344));
    jdff dff_B_WTHNYiGv2_2(.din(n23344), .dout(n23347));
    jdff dff_B_lnYCOwVq2_2(.din(n4482), .dout(n23350));
    jdff dff_B_uzd3W8qA3_1(.din(n4312), .dout(n23353));
    jdff dff_B_xjj871zb0_2(.din(n3912), .dout(n23356));
    jdff dff_B_BZQu8nka9_2(.din(n23356), .dout(n23359));
    jdff dff_B_c8yZwTfn0_2(.din(n23359), .dout(n23362));
    jdff dff_B_yv4d6TTA5_2(.din(n23362), .dout(n23365));
    jdff dff_B_WDPk0vP99_2(.din(n23365), .dout(n23368));
    jdff dff_B_BtEugkbS4_2(.din(n23368), .dout(n23371));
    jdff dff_B_8CIlX0JD2_2(.din(n23371), .dout(n23374));
    jdff dff_B_vDtilpDP2_2(.din(n23374), .dout(n23377));
    jdff dff_B_b2SqLpvp0_2(.din(n23377), .dout(n23380));
    jdff dff_B_icSYXwrt0_2(.din(n23380), .dout(n23383));
    jdff dff_B_GTN6xiao0_2(.din(n23383), .dout(n23386));
    jdff dff_B_IkiyTq7T5_2(.din(n23386), .dout(n23389));
    jdff dff_B_sBy8yfAK0_2(.din(n23389), .dout(n23392));
    jdff dff_B_ayjmuoYy3_2(.din(n23392), .dout(n23395));
    jdff dff_B_c4HkXHup8_2(.din(n23395), .dout(n23398));
    jdff dff_B_ewLgdc4O5_2(.din(n23398), .dout(n23401));
    jdff dff_B_0rz40acQ1_2(.din(n23401), .dout(n23404));
    jdff dff_B_pDr0YIfu4_2(.din(n23404), .dout(n23407));
    jdff dff_B_ArYQ0XeZ8_2(.din(n23407), .dout(n23410));
    jdff dff_B_M7tjpi6J9_2(.din(n23410), .dout(n23413));
    jdff dff_B_K1ETa2s77_2(.din(n23413), .dout(n23416));
    jdff dff_B_dUA6h99e5_2(.din(n23416), .dout(n23419));
    jdff dff_B_YoWvCeLF3_2(.din(n23419), .dout(n23422));
    jdff dff_B_I2RdSUql2_2(.din(n23422), .dout(n23425));
    jdff dff_B_mGmdX3Wl9_2(.din(n23425), .dout(n23428));
    jdff dff_B_Aq25DpYO1_2(.din(n23428), .dout(n23431));
    jdff dff_B_0zxA06rf9_2(.din(n23431), .dout(n23434));
    jdff dff_B_xeE0Cf714_2(.din(n4106), .dout(n23437));
    jdff dff_B_Xewy7ynQ2_1(.din(n3916), .dout(n23440));
    jdff dff_B_ILqYK7GA6_2(.din(n3535), .dout(n23443));
    jdff dff_B_KefUfuQX2_2(.din(n23443), .dout(n23446));
    jdff dff_B_vbYQ3d9e6_2(.din(n23446), .dout(n23449));
    jdff dff_B_FxTI3rpf0_2(.din(n23449), .dout(n23452));
    jdff dff_B_eaz4wfXi4_2(.din(n23452), .dout(n23455));
    jdff dff_B_jHkGQAW51_2(.din(n23455), .dout(n23458));
    jdff dff_B_OsQFIn089_2(.din(n23458), .dout(n23461));
    jdff dff_B_yMkFgDtb4_2(.din(n23461), .dout(n23464));
    jdff dff_B_oxnhuztm1_2(.din(n23464), .dout(n23467));
    jdff dff_B_soxTaaV85_2(.din(n23467), .dout(n23470));
    jdff dff_B_PLudMCF56_2(.din(n23470), .dout(n23473));
    jdff dff_B_G3qFdKgE6_2(.din(n23473), .dout(n23476));
    jdff dff_B_ShZ6kQEh3_2(.din(n23476), .dout(n23479));
    jdff dff_B_ynNPUrKu4_2(.din(n23479), .dout(n23482));
    jdff dff_B_PPTnP7aQ2_2(.din(n23482), .dout(n23485));
    jdff dff_B_HmDCQnBm7_2(.din(n23485), .dout(n23488));
    jdff dff_B_snohWNGp8_2(.din(n23488), .dout(n23491));
    jdff dff_B_9o4564HU1_2(.din(n23491), .dout(n23494));
    jdff dff_B_fV8OAf4n9_2(.din(n23494), .dout(n23497));
    jdff dff_B_xzvpndms1_2(.din(n23497), .dout(n23500));
    jdff dff_B_cAiJ0cTE5_2(.din(n23500), .dout(n23503));
    jdff dff_B_LglNHTVx1_2(.din(n23503), .dout(n23506));
    jdff dff_B_AguJD1uK1_2(.din(n23506), .dout(n23509));
    jdff dff_B_jwFo8Crr7_2(.din(n23509), .dout(n23512));
    jdff dff_B_srM51NvW5_2(.din(n3703), .dout(n23515));
    jdff dff_B_KizjIKLD4_1(.din(n3539), .dout(n23518));
    jdff dff_B_kJbx6HmA4_2(.din(n3134), .dout(n23521));
    jdff dff_B_B2LcDPZV8_2(.din(n23521), .dout(n23524));
    jdff dff_B_VVtjfoL76_2(.din(n23524), .dout(n23527));
    jdff dff_B_D6V39gPe4_2(.din(n23527), .dout(n23530));
    jdff dff_B_I7fehIHE4_2(.din(n23530), .dout(n23533));
    jdff dff_B_Xv1jmA005_2(.din(n23533), .dout(n23536));
    jdff dff_B_AzezYvDp3_2(.din(n23536), .dout(n23539));
    jdff dff_B_Lfu3r4Qc2_2(.din(n23539), .dout(n23542));
    jdff dff_B_Vxrn0VrF8_2(.din(n23542), .dout(n23545));
    jdff dff_B_joRcfVxS5_2(.din(n23545), .dout(n23548));
    jdff dff_B_GIy6Ni797_2(.din(n23548), .dout(n23551));
    jdff dff_B_tEBNFMUf8_2(.din(n23551), .dout(n23554));
    jdff dff_B_aQAknhHc8_2(.din(n23554), .dout(n23557));
    jdff dff_B_C3FlaVdQ2_2(.din(n23557), .dout(n23560));
    jdff dff_B_4rN7hxPq4_2(.din(n23560), .dout(n23563));
    jdff dff_B_oStUWTwr1_2(.din(n23563), .dout(n23566));
    jdff dff_B_1FcR4dni7_2(.din(n23566), .dout(n23569));
    jdff dff_B_whimdm246_2(.din(n23569), .dout(n23572));
    jdff dff_B_kwEysLM92_2(.din(n23572), .dout(n23575));
    jdff dff_B_5f3kWY4S0_2(.din(n23575), .dout(n23578));
    jdff dff_B_kYkqdPMr6_2(.din(n23578), .dout(n23581));
    jdff dff_B_JcBbMAdb9_2(.din(n3301), .dout(n23584));
    jdff dff_B_c8K0u9p28_1(.din(n3138), .dout(n23587));
    jdff dff_B_HqPS48kr8_2(.din(n2755), .dout(n23590));
    jdff dff_B_JBOVN3QN0_2(.din(n23590), .dout(n23593));
    jdff dff_B_7TY5rIS07_2(.din(n23593), .dout(n23596));
    jdff dff_B_nP7lwz5r2_2(.din(n23596), .dout(n23599));
    jdff dff_B_e4hR2Ggt0_2(.din(n23599), .dout(n23602));
    jdff dff_B_wfs4P79U9_2(.din(n23602), .dout(n23605));
    jdff dff_B_AnLpgX643_2(.din(n23605), .dout(n23608));
    jdff dff_B_EPu3zuoE4_2(.din(n23608), .dout(n23611));
    jdff dff_B_jk0muqlY7_2(.din(n23611), .dout(n23614));
    jdff dff_B_Dbv7Pg6n5_2(.din(n23614), .dout(n23617));
    jdff dff_B_EM1pjMts4_2(.din(n23617), .dout(n23620));
    jdff dff_B_32uSxC0p3_2(.din(n23620), .dout(n23623));
    jdff dff_B_CRrFrIAr8_2(.din(n23623), .dout(n23626));
    jdff dff_B_T16sNmeR3_2(.din(n23626), .dout(n23629));
    jdff dff_B_j2u7iEnl2_2(.din(n23629), .dout(n23632));
    jdff dff_B_qVFpwbDJ5_2(.din(n23632), .dout(n23635));
    jdff dff_B_vIE5lVX17_2(.din(n23635), .dout(n23638));
    jdff dff_B_BcXpF4rI7_2(.din(n23638), .dout(n23641));
    jdff dff_B_FgF8KqwX0_2(.din(n2896), .dout(n23644));
    jdff dff_B_gkIHDYrP0_1(.din(n2759), .dout(n23647));
    jdff dff_B_KPE4BNW90_2(.din(n2400), .dout(n23650));
    jdff dff_B_IxD6OlcQ7_2(.din(n23650), .dout(n23653));
    jdff dff_B_Q6TigjFH5_2(.din(n23653), .dout(n23656));
    jdff dff_B_ORohxeBL6_2(.din(n23656), .dout(n23659));
    jdff dff_B_xfRwrgGu7_2(.din(n23659), .dout(n23662));
    jdff dff_B_JRz79APs0_2(.din(n23662), .dout(n23665));
    jdff dff_B_vI6OPqDp0_2(.din(n23665), .dout(n23668));
    jdff dff_B_VQPOLqxI8_2(.din(n23668), .dout(n23671));
    jdff dff_B_n3VJb7os0_2(.din(n23671), .dout(n23674));
    jdff dff_B_PXpKiGS69_2(.din(n23674), .dout(n23677));
    jdff dff_B_0NrkS6646_2(.din(n23677), .dout(n23680));
    jdff dff_B_JAffA4Ep7_2(.din(n23680), .dout(n23683));
    jdff dff_B_qZizcAE34_2(.din(n23683), .dout(n23686));
    jdff dff_B_Pec7xNWs6_2(.din(n23686), .dout(n23689));
    jdff dff_B_TGg6KFiC7_2(.din(n23689), .dout(n23692));
    jdff dff_B_4fGVicy57_2(.din(n2514), .dout(n23695));
    jdff dff_B_6qB0P92B1_1(.din(n2404), .dout(n23698));
    jdff dff_B_7blUpne13_2(.din(n2072), .dout(n23701));
    jdff dff_B_C4QfKUdZ7_2(.din(n23701), .dout(n23704));
    jdff dff_B_ekc50hko6_2(.din(n23704), .dout(n23707));
    jdff dff_B_LJBvSjCD6_2(.din(n23707), .dout(n23710));
    jdff dff_B_aK4zCiUF0_2(.din(n23710), .dout(n23713));
    jdff dff_B_4L345AdN8_2(.din(n23713), .dout(n23716));
    jdff dff_B_ieqWtctJ7_2(.din(n23716), .dout(n23719));
    jdff dff_B_jBAJX7Gd4_2(.din(n23719), .dout(n23722));
    jdff dff_B_27o1vert5_2(.din(n23722), .dout(n23725));
    jdff dff_B_emLOxp1V6_2(.din(n23725), .dout(n23728));
    jdff dff_B_FXgapH284_2(.din(n23728), .dout(n23731));
    jdff dff_B_DbqvFnC43_2(.din(n23731), .dout(n23734));
    jdff dff_B_oy8umolf6_2(.din(n2159), .dout(n23737));
    jdff dff_B_rAYAdfFl2_1(.din(n2076), .dout(n23740));
    jdff dff_B_ja1CMELV8_2(.din(n1771), .dout(n23743));
    jdff dff_B_5qSuCpD44_2(.din(n23743), .dout(n23746));
    jdff dff_B_f8f72HM14_2(.din(n23746), .dout(n23749));
    jdff dff_B_L2PET60S9_2(.din(n23749), .dout(n23752));
    jdff dff_B_4bgFc24M3_2(.din(n23752), .dout(n23755));
    jdff dff_B_dSKmSjOY5_2(.din(n23755), .dout(n23758));
    jdff dff_B_yx21GZjs0_2(.din(n23758), .dout(n23761));
    jdff dff_B_NnjONBx14_2(.din(n23761), .dout(n23764));
    jdff dff_B_aWyavlEF5_2(.din(n23764), .dout(n23767));
    jdff dff_B_CmShW5m65_2(.din(n1831), .dout(n23770));
    jdff dff_B_QiWXyrP18_2(.din(n23770), .dout(n23773));
    jdff dff_B_okGvTIfp4_1(.din(n1774), .dout(n23776));
    jdff dff_B_Ovga210J9_1(.din(n23776), .dout(n23779));
    jdff dff_B_cfkcpT9w5_1(.din(n23779), .dout(n23782));
    jdff dff_B_DNOyaLVM2_1(.din(n23782), .dout(n23785));
    jdff dff_B_N1MTUlbu6_1(.din(n23785), .dout(n23788));
    jdff dff_B_Oo0S0JvP8_1(.din(n23788), .dout(n23791));
    jdff dff_B_2LjfKZ2q1_0(.din(n1530), .dout(n23794));
    jdff dff_B_fzZDPGCA0_0(.din(n23794), .dout(n23797));
    jdff dff_A_uHGO6zZS9_0(.din(n23802), .dout(n23799));
    jdff dff_A_qXO6zwHi7_0(.din(n23805), .dout(n23802));
    jdff dff_A_PzvLBQM62_0(.din(n1526), .dout(n23805));
    jdff dff_B_kfrBW14e5_1(.din(n1504), .dout(n23809));
    jdff dff_A_OqaIikFK2_0(.din(n1246), .dout(n23811));
    jdff dff_A_OSxUYutW3_1(.din(n23817), .dout(n23814));
    jdff dff_A_RVoeUevc7_1(.din(n1246), .dout(n23817));
    jdff dff_A_teBB2hqj4_1(.din(n23823), .dout(n23820));
    jdff dff_A_tV7cHCuR6_1(.din(n23826), .dout(n23823));
    jdff dff_A_MwvqcJvR8_1(.din(n23829), .dout(n23826));
    jdff dff_A_i0ZkdQHk1_1(.din(n23832), .dout(n23829));
    jdff dff_A_WrFDIzY00_1(.din(n23835), .dout(n23832));
    jdff dff_A_mAPv3Wu33_1(.din(n1496), .dout(n23835));
    jdff dff_B_3RnJicDM9_2(.din(n6239), .dout(n23839));
    jdff dff_B_VVOCdBKQ9_1(.din(n6231), .dout(n23842));
    jdff dff_B_rQGk3lVe3_2(.din(n6033), .dout(n23845));
    jdff dff_B_H1sxGiWm9_2(.din(n23845), .dout(n23848));
    jdff dff_B_SJ3sHZQ76_2(.din(n23848), .dout(n23851));
    jdff dff_B_vdXYDhFr4_2(.din(n23851), .dout(n23854));
    jdff dff_B_gwD71AgJ4_2(.din(n23854), .dout(n23857));
    jdff dff_B_FLBhM1gE1_2(.din(n23857), .dout(n23860));
    jdff dff_B_k97zJxyz8_2(.din(n23860), .dout(n23863));
    jdff dff_B_TIjQOkkX5_2(.din(n23863), .dout(n23866));
    jdff dff_B_C9K4kJzr3_2(.din(n23866), .dout(n23869));
    jdff dff_B_N4ORJPVi3_2(.din(n23869), .dout(n23872));
    jdff dff_B_Z0giA0840_2(.din(n23872), .dout(n23875));
    jdff dff_B_MFFiOSBY4_2(.din(n23875), .dout(n23878));
    jdff dff_B_MANj7Cr24_2(.din(n23878), .dout(n23881));
    jdff dff_B_K50yHLw83_2(.din(n23881), .dout(n23884));
    jdff dff_B_04MGH8kK4_2(.din(n23884), .dout(n23887));
    jdff dff_B_yKcc2K6C6_2(.din(n23887), .dout(n23890));
    jdff dff_B_oUwf0fKg8_2(.din(n23890), .dout(n23893));
    jdff dff_B_BboUODOo8_2(.din(n23893), .dout(n23896));
    jdff dff_B_SHciex9f9_2(.din(n23896), .dout(n23899));
    jdff dff_B_OoS0rA8j2_2(.din(n23899), .dout(n23902));
    jdff dff_B_4lqdVSLO9_2(.din(n23902), .dout(n23905));
    jdff dff_B_46iNrCSM2_2(.din(n23905), .dout(n23908));
    jdff dff_B_SyTGHSIE7_2(.din(n23908), .dout(n23911));
    jdff dff_B_JsB3ySxS8_2(.din(n23911), .dout(n23914));
    jdff dff_B_t0h8V9m91_2(.din(n23914), .dout(n23917));
    jdff dff_B_jZQQWcrI5_2(.din(n23917), .dout(n23920));
    jdff dff_B_HGM76Mk49_2(.din(n23920), .dout(n23923));
    jdff dff_B_DjSDpkoM1_2(.din(n23923), .dout(n23926));
    jdff dff_B_dc9NxKfl2_2(.din(n23926), .dout(n23929));
    jdff dff_B_WnYEq7mm6_2(.din(n23929), .dout(n23932));
    jdff dff_B_6E6uATDr7_2(.din(n23932), .dout(n23935));
    jdff dff_B_nB2Qk6472_2(.din(n23935), .dout(n23938));
    jdff dff_B_eBpkP9O22_2(.din(n23938), .dout(n23941));
    jdff dff_B_RtIma7D91_2(.din(n23941), .dout(n23944));
    jdff dff_B_GGChZvOx8_2(.din(n23944), .dout(n23947));
    jdff dff_B_yeOGpDpF3_2(.din(n23947), .dout(n23950));
    jdff dff_B_zGTN5gvK3_2(.din(n23950), .dout(n23953));
    jdff dff_B_MxzjAqhn0_2(.din(n23953), .dout(n23956));
    jdff dff_B_bigACyS58_2(.din(n23956), .dout(n23959));
    jdff dff_B_cOGu1qVi3_2(.din(n23959), .dout(n23962));
    jdff dff_B_dLX3NpNs7_2(.din(n23962), .dout(n23965));
    jdff dff_B_z1i7qGpa8_2(.din(n23965), .dout(n23968));
    jdff dff_B_vFbDe1Cc7_2(.din(n23968), .dout(n23971));
    jdff dff_B_L0r0AVv03_2(.din(n23971), .dout(n23974));
    jdff dff_B_iJxvJt2Q7_2(.din(n23974), .dout(n23977));
    jdff dff_B_Hxpq3uqt4_2(.din(n23977), .dout(n23980));
    jdff dff_B_DRCkAmS47_2(.din(n23980), .dout(n23983));
    jdff dff_B_oshq8HRc1_2(.din(n23983), .dout(n23986));
    jdff dff_B_8udX8bne1_2(.din(n23986), .dout(n23989));
    jdff dff_B_rqcdsL8S1_1(.din(n6224), .dout(n23992));
    jdff dff_A_4JJX4vbh2_1(.din(n6045), .dout(n23994));
    jdff dff_B_caV1Uciq4_1(.din(n6037), .dout(n23998));
    jdff dff_B_00vZXMjC9_2(.din(n5815), .dout(n24001));
    jdff dff_B_OMYvfEqK5_2(.din(n24001), .dout(n24004));
    jdff dff_B_DsR74SI38_2(.din(n24004), .dout(n24007));
    jdff dff_B_2Knia5NI5_2(.din(n24007), .dout(n24010));
    jdff dff_B_T6O79sgf8_2(.din(n24010), .dout(n24013));
    jdff dff_B_z9TPqOtJ6_2(.din(n24013), .dout(n24016));
    jdff dff_B_6Fef7Z8Z2_2(.din(n24016), .dout(n24019));
    jdff dff_B_TRGcbW495_2(.din(n24019), .dout(n24022));
    jdff dff_B_Ue3RsntW9_2(.din(n24022), .dout(n24025));
    jdff dff_B_474AUWGh0_2(.din(n24025), .dout(n24028));
    jdff dff_B_ajBr2uW02_2(.din(n24028), .dout(n24031));
    jdff dff_B_fRCweLPu0_2(.din(n24031), .dout(n24034));
    jdff dff_B_I7lrImhF5_2(.din(n24034), .dout(n24037));
    jdff dff_B_2XBlZWlG4_2(.din(n24037), .dout(n24040));
    jdff dff_B_tKsrIPLH9_2(.din(n24040), .dout(n24043));
    jdff dff_B_ICsQXzqu8_2(.din(n24043), .dout(n24046));
    jdff dff_B_6QXffW1I2_2(.din(n24046), .dout(n24049));
    jdff dff_B_5Av5Qla75_2(.din(n24049), .dout(n24052));
    jdff dff_B_SGU9ONIy9_2(.din(n24052), .dout(n24055));
    jdff dff_B_AScHc9bz7_2(.din(n24055), .dout(n24058));
    jdff dff_B_rIh4aMwv5_2(.din(n24058), .dout(n24061));
    jdff dff_B_78i17mhF0_2(.din(n24061), .dout(n24064));
    jdff dff_B_ptYBTz6k8_2(.din(n24064), .dout(n24067));
    jdff dff_B_lIpR6Luf5_2(.din(n24067), .dout(n24070));
    jdff dff_B_sa5nhSK93_2(.din(n24070), .dout(n24073));
    jdff dff_B_9vYERfv13_2(.din(n24073), .dout(n24076));
    jdff dff_B_AmwdL0Gj9_2(.din(n24076), .dout(n24079));
    jdff dff_B_XJk98zk63_2(.din(n24079), .dout(n24082));
    jdff dff_B_mc0IQvLR4_2(.din(n24082), .dout(n24085));
    jdff dff_B_t9UkyfRx6_2(.din(n24085), .dout(n24088));
    jdff dff_B_rxn0rczN1_2(.din(n24088), .dout(n24091));
    jdff dff_B_HQz4GrLV4_2(.din(n24091), .dout(n24094));
    jdff dff_B_P6z2MrgN2_2(.din(n24094), .dout(n24097));
    jdff dff_B_Q3l6Dwu72_2(.din(n24097), .dout(n24100));
    jdff dff_B_TQORNAjw3_2(.din(n24100), .dout(n24103));
    jdff dff_B_Ni5NJVNp1_2(.din(n24103), .dout(n24106));
    jdff dff_B_oLOv9SCj5_2(.din(n24106), .dout(n24109));
    jdff dff_B_ue0jFElA2_2(.din(n24109), .dout(n24112));
    jdff dff_B_4Jvsh2GY7_2(.din(n24112), .dout(n24115));
    jdff dff_B_lo3ZEi1K0_2(.din(n24115), .dout(n24118));
    jdff dff_B_lc7UO8933_2(.din(n24118), .dout(n24121));
    jdff dff_B_svI6uF3k7_2(.din(n24121), .dout(n24124));
    jdff dff_B_zYjooRPh7_2(.din(n24124), .dout(n24127));
    jdff dff_B_rKUlpOpo5_2(.din(n5827), .dout(n24130));
    jdff dff_B_OVFaeoJQ4_1(.din(n5819), .dout(n24133));
    jdff dff_B_dxyA2MqL0_2(.din(n5570), .dout(n24136));
    jdff dff_B_F0NMUvbu7_2(.din(n24136), .dout(n24139));
    jdff dff_B_jMvfmP3p5_2(.din(n24139), .dout(n24142));
    jdff dff_B_q5vBtwrN5_2(.din(n24142), .dout(n24145));
    jdff dff_B_AwtR4eou3_2(.din(n24145), .dout(n24148));
    jdff dff_B_q1W5I5cG8_2(.din(n24148), .dout(n24151));
    jdff dff_B_8DqNIZRW2_2(.din(n24151), .dout(n24154));
    jdff dff_B_dtoVpleY8_2(.din(n24154), .dout(n24157));
    jdff dff_B_KpsN6g3A3_2(.din(n24157), .dout(n24160));
    jdff dff_B_UUpkqryu9_2(.din(n24160), .dout(n24163));
    jdff dff_B_Z0mBabTw8_2(.din(n24163), .dout(n24166));
    jdff dff_B_70Vadccr9_2(.din(n24166), .dout(n24169));
    jdff dff_B_BkAydNWi0_2(.din(n24169), .dout(n24172));
    jdff dff_B_Kc7AVJjm8_2(.din(n24172), .dout(n24175));
    jdff dff_B_QoXqCVU15_2(.din(n24175), .dout(n24178));
    jdff dff_B_RkQ1Wc8J6_2(.din(n24178), .dout(n24181));
    jdff dff_B_KsuwzJpz1_2(.din(n24181), .dout(n24184));
    jdff dff_B_aEWQcq2K0_2(.din(n24184), .dout(n24187));
    jdff dff_B_TdSHs97D6_2(.din(n24187), .dout(n24190));
    jdff dff_B_ojYdJ6xP7_2(.din(n24190), .dout(n24193));
    jdff dff_B_2aqGnBmB3_2(.din(n24193), .dout(n24196));
    jdff dff_B_BY9jdHMx3_2(.din(n24196), .dout(n24199));
    jdff dff_B_G75FPiZ94_2(.din(n24199), .dout(n24202));
    jdff dff_B_KH1bkfDM3_2(.din(n24202), .dout(n24205));
    jdff dff_B_ZCw7RZE63_2(.din(n24205), .dout(n24208));
    jdff dff_B_O5R55zZc6_2(.din(n24208), .dout(n24211));
    jdff dff_B_CltihA214_2(.din(n24211), .dout(n24214));
    jdff dff_B_NFs8nu665_2(.din(n24214), .dout(n24217));
    jdff dff_B_dA59S4zW5_2(.din(n24217), .dout(n24220));
    jdff dff_B_wZS7RfwH9_2(.din(n24220), .dout(n24223));
    jdff dff_B_ekZVA6Pp4_2(.din(n24223), .dout(n24226));
    jdff dff_B_qDnt8Nwe4_2(.din(n24226), .dout(n24229));
    jdff dff_B_5gyJeHCz5_2(.din(n24229), .dout(n24232));
    jdff dff_B_7IOPICYw1_2(.din(n24232), .dout(n24235));
    jdff dff_B_3b8WpZfL0_2(.din(n24235), .dout(n24238));
    jdff dff_B_YnabyG0G3_2(.din(n24238), .dout(n24241));
    jdff dff_B_n77vf1nt9_2(.din(n24241), .dout(n24244));
    jdff dff_B_Vm42VOx80_2(.din(n24244), .dout(n24247));
    jdff dff_B_m0eMMI8i3_2(.din(n24247), .dout(n24250));
    jdff dff_B_ep9J85lm5_1(.din(n5574), .dout(n24253));
    jdff dff_B_NITjvwZO1_2(.din(n5298), .dout(n24256));
    jdff dff_B_pp1IcoEZ3_2(.din(n24256), .dout(n24259));
    jdff dff_B_yCg6xIBm2_2(.din(n24259), .dout(n24262));
    jdff dff_B_AXH3ceeX4_2(.din(n24262), .dout(n24265));
    jdff dff_B_hBxhxHyA9_2(.din(n24265), .dout(n24268));
    jdff dff_B_2VNxjfxP7_2(.din(n24268), .dout(n24271));
    jdff dff_B_jUKy0EVc6_2(.din(n24271), .dout(n24274));
    jdff dff_B_pVmGhPvx3_2(.din(n24274), .dout(n24277));
    jdff dff_B_uKayVfot0_2(.din(n24277), .dout(n24280));
    jdff dff_B_vvfc7eE66_2(.din(n24280), .dout(n24283));
    jdff dff_B_5hX1zHPV4_2(.din(n24283), .dout(n24286));
    jdff dff_B_dcXSkwkr4_2(.din(n24286), .dout(n24289));
    jdff dff_B_wirYtMQL7_2(.din(n24289), .dout(n24292));
    jdff dff_B_o6umcOOP8_2(.din(n24292), .dout(n24295));
    jdff dff_B_d9CUyejE7_2(.din(n24295), .dout(n24298));
    jdff dff_B_L8ISDlfd1_2(.din(n24298), .dout(n24301));
    jdff dff_B_j1J6srgp4_2(.din(n24301), .dout(n24304));
    jdff dff_B_VQnKRV0Y2_2(.din(n24304), .dout(n24307));
    jdff dff_B_rhduM2fl6_2(.din(n24307), .dout(n24310));
    jdff dff_B_lG6L7IyP0_2(.din(n24310), .dout(n24313));
    jdff dff_B_I4ezPKmf1_2(.din(n24313), .dout(n24316));
    jdff dff_B_I5Mn5VT17_2(.din(n24316), .dout(n24319));
    jdff dff_B_63fQgczl7_2(.din(n24319), .dout(n24322));
    jdff dff_B_stByCNqY7_2(.din(n24322), .dout(n24325));
    jdff dff_B_PQDJDI380_2(.din(n24325), .dout(n24328));
    jdff dff_B_zFRQ0nHT0_2(.din(n24328), .dout(n24331));
    jdff dff_B_ErKhzT9D7_2(.din(n24331), .dout(n24334));
    jdff dff_B_yXmbOzmP5_2(.din(n24334), .dout(n24337));
    jdff dff_B_T5upasdN9_2(.din(n24337), .dout(n24340));
    jdff dff_B_JtUGBNnw2_2(.din(n24340), .dout(n24343));
    jdff dff_B_hI6yFXJz7_2(.din(n24343), .dout(n24346));
    jdff dff_B_PNQIdWr74_2(.din(n24346), .dout(n24349));
    jdff dff_B_wjpq9D6j9_2(.din(n24349), .dout(n24352));
    jdff dff_B_vRvr2wr26_2(.din(n24352), .dout(n24355));
    jdff dff_B_Nk3AB6I91_2(.din(n24355), .dout(n24358));
    jdff dff_B_2ywxSxKj8_2(.din(n24358), .dout(n24361));
    jdff dff_B_HISQ8N1N8_2(.din(n5449), .dout(n24364));
    jdff dff_B_bc8EOeQJ5_1(.din(n5302), .dout(n24367));
    jdff dff_B_9dobeQkJ7_2(.din(n4999), .dout(n24370));
    jdff dff_B_jyVHoDC70_2(.din(n24370), .dout(n24373));
    jdff dff_B_m7F28Hkb4_2(.din(n24373), .dout(n24376));
    jdff dff_B_eMQ3XJKt9_2(.din(n24376), .dout(n24379));
    jdff dff_B_fTpM45iT8_2(.din(n24379), .dout(n24382));
    jdff dff_B_hhwn8Kaf2_2(.din(n24382), .dout(n24385));
    jdff dff_B_1gBks4D78_2(.din(n24385), .dout(n24388));
    jdff dff_B_EUu8PYPN4_2(.din(n24388), .dout(n24391));
    jdff dff_B_dRIsLWDc5_2(.din(n24391), .dout(n24394));
    jdff dff_B_okH6juCc3_2(.din(n24394), .dout(n24397));
    jdff dff_B_HZpdYgyn7_2(.din(n24397), .dout(n24400));
    jdff dff_B_Pj4hLcsP1_2(.din(n24400), .dout(n24403));
    jdff dff_B_NYENvobe8_2(.din(n24403), .dout(n24406));
    jdff dff_B_wzcWJJa17_2(.din(n24406), .dout(n24409));
    jdff dff_B_Y17Tzvel4_2(.din(n24409), .dout(n24412));
    jdff dff_B_OAL4d9VV7_2(.din(n24412), .dout(n24415));
    jdff dff_B_uFMc3xi21_2(.din(n24415), .dout(n24418));
    jdff dff_B_1CWtZyUO2_2(.din(n24418), .dout(n24421));
    jdff dff_B_6sOJFOLV6_2(.din(n24421), .dout(n24424));
    jdff dff_B_PLWr5jKS6_2(.din(n24424), .dout(n24427));
    jdff dff_B_74DTXMSh3_2(.din(n24427), .dout(n24430));
    jdff dff_B_ajl8NgPG4_2(.din(n24430), .dout(n24433));
    jdff dff_B_fMU1GJRk7_2(.din(n24433), .dout(n24436));
    jdff dff_B_hoNMd5JW0_2(.din(n24436), .dout(n24439));
    jdff dff_B_Yn3XMZPW3_2(.din(n24439), .dout(n24442));
    jdff dff_B_muVvpKeL8_2(.din(n24442), .dout(n24445));
    jdff dff_B_ownsU5WY6_2(.din(n24445), .dout(n24448));
    jdff dff_B_KaOcZpno8_2(.din(n24448), .dout(n24451));
    jdff dff_B_X3GzVAcQ1_2(.din(n24451), .dout(n24454));
    jdff dff_B_0u3Qh3XZ2_2(.din(n24454), .dout(n24457));
    jdff dff_B_5S0Pu4gx2_2(.din(n24457), .dout(n24460));
    jdff dff_B_gtqgsyJ29_2(.din(n24460), .dout(n24463));
    jdff dff_B_ytPP6zC89_2(.din(n24463), .dout(n24466));
    jdff dff_B_1JzL5Mq57_2(.din(n5150), .dout(n24469));
    jdff dff_B_WVn4gxIs4_1(.din(n5003), .dout(n24472));
    jdff dff_B_ip10Dipr1_2(.din(n4673), .dout(n24475));
    jdff dff_B_F6lJWV9g8_2(.din(n24475), .dout(n24478));
    jdff dff_B_ZeC5lp6w7_2(.din(n24478), .dout(n24481));
    jdff dff_B_Fe3noJUt0_2(.din(n24481), .dout(n24484));
    jdff dff_B_6rMTpEze6_2(.din(n24484), .dout(n24487));
    jdff dff_B_iHGDDPCs5_2(.din(n24487), .dout(n24490));
    jdff dff_B_qAzHfZTW8_2(.din(n24490), .dout(n24493));
    jdff dff_B_toU4PPUN8_2(.din(n24493), .dout(n24496));
    jdff dff_B_ncnBoFdE2_2(.din(n24496), .dout(n24499));
    jdff dff_B_skqtymb74_2(.din(n24499), .dout(n24502));
    jdff dff_B_0VPZXGuf9_2(.din(n24502), .dout(n24505));
    jdff dff_B_YBZzA1aF4_2(.din(n24505), .dout(n24508));
    jdff dff_B_apHUwt5q6_2(.din(n24508), .dout(n24511));
    jdff dff_B_9iGDo3O46_2(.din(n24511), .dout(n24514));
    jdff dff_B_iAabzOLN2_2(.din(n24514), .dout(n24517));
    jdff dff_B_64YivDpv3_2(.din(n24517), .dout(n24520));
    jdff dff_B_GIcp11qT1_2(.din(n24520), .dout(n24523));
    jdff dff_B_Rr24kxsg3_2(.din(n24523), .dout(n24526));
    jdff dff_B_oxBHb8iV9_2(.din(n24526), .dout(n24529));
    jdff dff_B_BEKKcG2v0_2(.din(n24529), .dout(n24532));
    jdff dff_B_uM1nMhGN2_2(.din(n24532), .dout(n24535));
    jdff dff_B_Z3txKOzB0_2(.din(n24535), .dout(n24538));
    jdff dff_B_NsuF8KsE1_2(.din(n24538), .dout(n24541));
    jdff dff_B_SAvm11bq7_2(.din(n24541), .dout(n24544));
    jdff dff_B_L8G6ABRI2_2(.din(n24544), .dout(n24547));
    jdff dff_B_oFuVGFgH8_2(.din(n24547), .dout(n24550));
    jdff dff_B_eFMZsobE9_2(.din(n24550), .dout(n24553));
    jdff dff_B_2YLg9TQ78_2(.din(n24553), .dout(n24556));
    jdff dff_B_T1HO2Rd15_2(.din(n24556), .dout(n24559));
    jdff dff_B_7zpv10YT7_2(.din(n24559), .dout(n24562));
    jdff dff_B_mADqmqP18_2(.din(n4824), .dout(n24565));
    jdff dff_B_nwJXkFV64_1(.din(n4677), .dout(n24568));
    jdff dff_B_LiWGV6py7_2(.din(n4327), .dout(n24571));
    jdff dff_B_We4PU8jH9_2(.din(n24571), .dout(n24574));
    jdff dff_B_lcrIB0qU5_2(.din(n24574), .dout(n24577));
    jdff dff_B_cjjx011v3_2(.din(n24577), .dout(n24580));
    jdff dff_B_rrpxWGx76_2(.din(n24580), .dout(n24583));
    jdff dff_B_zWgXi6xT9_2(.din(n24583), .dout(n24586));
    jdff dff_B_eAkQYT9l8_2(.din(n24586), .dout(n24589));
    jdff dff_B_K8jmrcin0_2(.din(n24589), .dout(n24592));
    jdff dff_B_Uqjnyzse5_2(.din(n24592), .dout(n24595));
    jdff dff_B_2fxMLfWK8_2(.din(n24595), .dout(n24598));
    jdff dff_B_jAXTuAWY0_2(.din(n24598), .dout(n24601));
    jdff dff_B_WrljdxqX4_2(.din(n24601), .dout(n24604));
    jdff dff_B_G8Sh7LQa3_2(.din(n24604), .dout(n24607));
    jdff dff_B_VyJhSFsX7_2(.din(n24607), .dout(n24610));
    jdff dff_B_n4fjb4Hx4_2(.din(n24610), .dout(n24613));
    jdff dff_B_ctJpDmhB3_2(.din(n24613), .dout(n24616));
    jdff dff_B_dKvI9GS99_2(.din(n24616), .dout(n24619));
    jdff dff_B_kzUkZZI13_2(.din(n24619), .dout(n24622));
    jdff dff_B_7ZeqhotU4_2(.din(n24622), .dout(n24625));
    jdff dff_B_FgEaB1x25_2(.din(n24625), .dout(n24628));
    jdff dff_B_M6ZF9rCk4_2(.din(n24628), .dout(n24631));
    jdff dff_B_mRnJoWnI9_2(.din(n24631), .dout(n24634));
    jdff dff_B_uCuvAqPS5_2(.din(n24634), .dout(n24637));
    jdff dff_B_aZ27IuzA5_2(.din(n24637), .dout(n24640));
    jdff dff_B_x8ueRvEL4_2(.din(n24640), .dout(n24643));
    jdff dff_B_V7vgzhww6_2(.din(n24643), .dout(n24646));
    jdff dff_B_44hlovNk6_2(.din(n24646), .dout(n24649));
    jdff dff_B_MsvinaVe8_2(.din(n4474), .dout(n24652));
    jdff dff_B_k0AmojMX2_1(.din(n4331), .dout(n24655));
    jdff dff_B_dBxrUPST0_2(.din(n3931), .dout(n24658));
    jdff dff_B_6FQvDauU0_2(.din(n24658), .dout(n24661));
    jdff dff_B_On3kuz2s7_2(.din(n24661), .dout(n24664));
    jdff dff_B_i4PD0MDB5_2(.din(n24664), .dout(n24667));
    jdff dff_B_ZAyC6yzB2_2(.din(n24667), .dout(n24670));
    jdff dff_B_ACqCUdJK3_2(.din(n24670), .dout(n24673));
    jdff dff_B_7wAoJzCG3_2(.din(n24673), .dout(n24676));
    jdff dff_B_5imdgR868_2(.din(n24676), .dout(n24679));
    jdff dff_B_ezW95HMd0_2(.din(n24679), .dout(n24682));
    jdff dff_B_2hjVwVmF8_2(.din(n24682), .dout(n24685));
    jdff dff_B_QBlXEqT10_2(.din(n24685), .dout(n24688));
    jdff dff_B_uAyDHpfw6_2(.din(n24688), .dout(n24691));
    jdff dff_B_zMbHL9B32_2(.din(n24691), .dout(n24694));
    jdff dff_B_598SblUx5_2(.din(n24694), .dout(n24697));
    jdff dff_B_FFHcRYqL3_2(.din(n24697), .dout(n24700));
    jdff dff_B_xkdNef0i0_2(.din(n24700), .dout(n24703));
    jdff dff_B_mKinpzrY2_2(.din(n24703), .dout(n24706));
    jdff dff_B_sVlZZoUM2_2(.din(n24706), .dout(n24709));
    jdff dff_B_wizdV6E65_2(.din(n24709), .dout(n24712));
    jdff dff_B_WmzQRrq68_2(.din(n24712), .dout(n24715));
    jdff dff_B_RfEcLeU20_2(.din(n24715), .dout(n24718));
    jdff dff_B_hpnRPkPl8_2(.din(n24718), .dout(n24721));
    jdff dff_B_BOHMR4jD0_2(.din(n24721), .dout(n24724));
    jdff dff_B_zmFlblHR9_2(.din(n24724), .dout(n24727));
    jdff dff_B_ArKrp9Jo9_2(.din(n4098), .dout(n24730));
    jdff dff_B_IHPr1Lw29_1(.din(n3935), .dout(n24733));
    jdff dff_B_tXrxXVHm9_2(.din(n3554), .dout(n24736));
    jdff dff_B_MrHLKQ150_2(.din(n24736), .dout(n24739));
    jdff dff_B_ibuG9Ba73_2(.din(n24739), .dout(n24742));
    jdff dff_B_naOkVaFF0_2(.din(n24742), .dout(n24745));
    jdff dff_B_UTSv0xFq2_2(.din(n24745), .dout(n24748));
    jdff dff_B_H2a9u2ng7_2(.din(n24748), .dout(n24751));
    jdff dff_B_ERHndalF5_2(.din(n24751), .dout(n24754));
    jdff dff_B_q2HbTIzh3_2(.din(n24754), .dout(n24757));
    jdff dff_B_wrcCZKqo9_2(.din(n24757), .dout(n24760));
    jdff dff_B_ZDwDkWAI9_2(.din(n24760), .dout(n24763));
    jdff dff_B_HWroxUo33_2(.din(n24763), .dout(n24766));
    jdff dff_B_g1Lf0It04_2(.din(n24766), .dout(n24769));
    jdff dff_B_e6WgFQ6R8_2(.din(n24769), .dout(n24772));
    jdff dff_B_kpoUAvar0_2(.din(n24772), .dout(n24775));
    jdff dff_B_5xcht1sV5_2(.din(n24775), .dout(n24778));
    jdff dff_B_LIuaEXWL2_2(.din(n24778), .dout(n24781));
    jdff dff_B_JpvsrTgi6_2(.din(n24781), .dout(n24784));
    jdff dff_B_j5B9MQpc4_2(.din(n24784), .dout(n24787));
    jdff dff_B_0d3qYfrT5_2(.din(n24787), .dout(n24790));
    jdff dff_B_NlFy0QL04_2(.din(n24790), .dout(n24793));
    jdff dff_B_AU6jyrFE3_2(.din(n24793), .dout(n24796));
    jdff dff_B_hOikBsCD4_2(.din(n3695), .dout(n24799));
    jdff dff_B_xA5TsFm41_1(.din(n3558), .dout(n24802));
    jdff dff_B_5Xu7gypW2_2(.din(n3153), .dout(n24805));
    jdff dff_B_VbfjyOeY5_2(.din(n24805), .dout(n24808));
    jdff dff_B_rPfXnYEv0_2(.din(n24808), .dout(n24811));
    jdff dff_B_Whxa2VIo9_2(.din(n24811), .dout(n24814));
    jdff dff_B_JbtUBMFH5_2(.din(n24814), .dout(n24817));
    jdff dff_B_eCibOGKe4_2(.din(n24817), .dout(n24820));
    jdff dff_B_SofNfQdv7_2(.din(n24820), .dout(n24823));
    jdff dff_B_DxpG3HVZ7_2(.din(n24823), .dout(n24826));
    jdff dff_B_UMPJEe397_2(.din(n24826), .dout(n24829));
    jdff dff_B_DEN1JuF13_2(.din(n24829), .dout(n24832));
    jdff dff_B_SvVeqdPa7_2(.din(n24832), .dout(n24835));
    jdff dff_B_jwUptlux1_2(.din(n24835), .dout(n24838));
    jdff dff_B_WFlrYD1e1_2(.din(n24838), .dout(n24841));
    jdff dff_B_jiy5FE7l9_2(.din(n24841), .dout(n24844));
    jdff dff_B_BeVZ6VZy0_2(.din(n24844), .dout(n24847));
    jdff dff_B_hipvSVQU7_2(.din(n24847), .dout(n24850));
    jdff dff_B_LkHXZCBK7_2(.din(n24850), .dout(n24853));
    jdff dff_B_pfabGU1z4_2(.din(n24853), .dout(n24856));
    jdff dff_B_n9EISm401_2(.din(n3293), .dout(n24859));
    jdff dff_B_HJQyML745_1(.din(n3157), .dout(n24862));
    jdff dff_B_wQfdFuV10_2(.din(n2774), .dout(n24865));
    jdff dff_B_o73wuKI98_2(.din(n24865), .dout(n24868));
    jdff dff_B_wmM4FHRy8_2(.din(n24868), .dout(n24871));
    jdff dff_B_3FrgMzfP3_2(.din(n24871), .dout(n24874));
    jdff dff_B_zzCFyGPl5_2(.din(n24874), .dout(n24877));
    jdff dff_B_CTrWC2XS6_2(.din(n24877), .dout(n24880));
    jdff dff_B_7bFV2QGw0_2(.din(n24880), .dout(n24883));
    jdff dff_B_NeFY834T1_2(.din(n24883), .dout(n24886));
    jdff dff_B_7VkI8jLT7_2(.din(n24886), .dout(n24889));
    jdff dff_B_i1IxUYqg2_2(.din(n24889), .dout(n24892));
    jdff dff_B_knIISLSD0_2(.din(n24892), .dout(n24895));
    jdff dff_B_lARREP0g7_2(.din(n24895), .dout(n24898));
    jdff dff_B_g7j7Yk6r6_2(.din(n24898), .dout(n24901));
    jdff dff_B_XkKe7h4n6_2(.din(n24901), .dout(n24904));
    jdff dff_B_dOQjWle73_2(.din(n24904), .dout(n24907));
    jdff dff_B_yEpiPgRN8_2(.din(n2888), .dout(n24910));
    jdff dff_B_bSQO3Iix9_1(.din(n2778), .dout(n24913));
    jdff dff_B_KbwQes492_2(.din(n2419), .dout(n24916));
    jdff dff_B_IXmf1d398_2(.din(n24916), .dout(n24919));
    jdff dff_B_ix1OoRRr9_2(.din(n24919), .dout(n24922));
    jdff dff_B_uCJoVFSw0_2(.din(n24922), .dout(n24925));
    jdff dff_B_5xjfZ3Wp0_2(.din(n24925), .dout(n24928));
    jdff dff_B_X1viEgLQ7_2(.din(n24928), .dout(n24931));
    jdff dff_B_YuiNqHBZ8_2(.din(n24931), .dout(n24934));
    jdff dff_B_YOyAP99l4_2(.din(n24934), .dout(n24937));
    jdff dff_B_Uk4p2vjt6_2(.din(n24937), .dout(n24940));
    jdff dff_B_oQsncDie8_2(.din(n24940), .dout(n24943));
    jdff dff_B_PqihfLAO8_2(.din(n24943), .dout(n24946));
    jdff dff_B_7W6IBFpX8_2(.din(n24946), .dout(n24949));
    jdff dff_B_Q5STwsBo3_2(.din(n2506), .dout(n24952));
    jdff dff_B_vavzs6245_1(.din(n2423), .dout(n24955));
    jdff dff_B_uFybdbnK0_2(.din(n2091), .dout(n24958));
    jdff dff_B_0LVi9f7f4_2(.din(n24958), .dout(n24961));
    jdff dff_B_ZR15t9k95_2(.din(n24961), .dout(n24964));
    jdff dff_B_uoKljbTd4_2(.din(n24964), .dout(n24967));
    jdff dff_B_GalnD0kl1_2(.din(n24967), .dout(n24970));
    jdff dff_B_ykNEyVAn8_2(.din(n24970), .dout(n24973));
    jdff dff_B_WjD1AETW3_2(.din(n24973), .dout(n24976));
    jdff dff_B_bsuqZ2859_2(.din(n24976), .dout(n24979));
    jdff dff_B_jZe4YHWU3_2(.din(n24979), .dout(n24982));
    jdff dff_B_OhS1WdKY6_2(.din(n2151), .dout(n24985));
    jdff dff_B_Y11zjUIr9_2(.din(n24985), .dout(n24988));
    jdff dff_B_2NBhPVEo0_1(.din(n2094), .dout(n24991));
    jdff dff_B_yhRwLhSl0_1(.din(n24991), .dout(n24994));
    jdff dff_B_h5csbh3Q4_1(.din(n24994), .dout(n24997));
    jdff dff_B_A6id4RZi6_1(.din(n24997), .dout(n25000));
    jdff dff_B_tz6VrQ7D8_1(.din(n25000), .dout(n25003));
    jdff dff_B_CbMh0etk8_1(.din(n25003), .dout(n25006));
    jdff dff_B_clarPqnr6_0(.din(n1823), .dout(n25009));
    jdff dff_B_5EYqdB1x0_0(.din(n25009), .dout(n25012));
    jdff dff_A_yizNcz2A1_0(.din(n25017), .dout(n25014));
    jdff dff_A_sFCCDAuD8_0(.din(n25020), .dout(n25017));
    jdff dff_A_BnbUiBaX3_0(.din(n1819), .dout(n25020));
    jdff dff_B_pIrr73m08_1(.din(n1797), .dout(n25024));
    jdff dff_A_VEjDMFPq4_0(.din(n1512), .dout(n25026));
    jdff dff_A_SAfrAM5U4_1(.din(n25032), .dout(n25029));
    jdff dff_A_DzAcwloZ4_1(.din(n1512), .dout(n25032));
    jdff dff_A_ajZXznoi4_1(.din(n25038), .dout(n25035));
    jdff dff_A_2oHCCgGu6_1(.din(n25041), .dout(n25038));
    jdff dff_A_BK8X57VK0_1(.din(n25044), .dout(n25041));
    jdff dff_A_PbKr4Kqu4_1(.din(n25047), .dout(n25044));
    jdff dff_A_0GWR2Htb6_1(.din(n25050), .dout(n25047));
    jdff dff_A_6STtgGwI6_1(.din(n1789), .dout(n25050));
    jdff dff_B_TCewL5c97_1(.din(n6539), .dout(n25054));
    jdff dff_A_gs11IcZb5_1(.din(n6416), .dout(n25056));
    jdff dff_B_ZNA61zx23_1(.din(n6408), .dout(n25060));
    jdff dff_B_TkY1yLGK6_2(.din(n6246), .dout(n25063));
    jdff dff_B_diW2C7mX8_2(.din(n25063), .dout(n25066));
    jdff dff_B_rE5T2yVe7_2(.din(n25066), .dout(n25069));
    jdff dff_B_CS8zggMj5_2(.din(n25069), .dout(n25072));
    jdff dff_B_b2mo3lKz6_2(.din(n25072), .dout(n25075));
    jdff dff_B_KLT5Lpxt9_2(.din(n25075), .dout(n25078));
    jdff dff_B_b3FesVu59_2(.din(n25078), .dout(n25081));
    jdff dff_B_Ph3YzaFY7_2(.din(n25081), .dout(n25084));
    jdff dff_B_ANayHqti9_2(.din(n25084), .dout(n25087));
    jdff dff_B_4JXILDJZ6_2(.din(n25087), .dout(n25090));
    jdff dff_B_CfMFsKap0_2(.din(n25090), .dout(n25093));
    jdff dff_B_RWGSRGPx5_2(.din(n25093), .dout(n25096));
    jdff dff_B_9K3JBp0j7_2(.din(n25096), .dout(n25099));
    jdff dff_B_zJqTLJr99_2(.din(n25099), .dout(n25102));
    jdff dff_B_99CbURTR4_2(.din(n25102), .dout(n25105));
    jdff dff_B_GI3UMVU34_2(.din(n25105), .dout(n25108));
    jdff dff_B_5KSbgHdb9_2(.din(n25108), .dout(n25111));
    jdff dff_B_eGCNUpTC8_2(.din(n25111), .dout(n25114));
    jdff dff_B_bu3eTSlq2_2(.din(n25114), .dout(n25117));
    jdff dff_B_9otfr0AT1_2(.din(n25117), .dout(n25120));
    jdff dff_B_eh42FrmY0_2(.din(n25120), .dout(n25123));
    jdff dff_B_rawarsQ76_2(.din(n25123), .dout(n25126));
    jdff dff_B_FgThDuMj4_2(.din(n25126), .dout(n25129));
    jdff dff_B_vGmS6IKl5_2(.din(n25129), .dout(n25132));
    jdff dff_B_0C2ytVHC6_2(.din(n25132), .dout(n25135));
    jdff dff_B_Jq9SG4xc0_2(.din(n25135), .dout(n25138));
    jdff dff_B_fmhu7x7C5_2(.din(n25138), .dout(n25141));
    jdff dff_B_rWFzzuz68_2(.din(n25141), .dout(n25144));
    jdff dff_B_F5bXzkmW5_2(.din(n25144), .dout(n25147));
    jdff dff_B_n9uHyAWm4_2(.din(n25147), .dout(n25150));
    jdff dff_B_UWOLfndn8_2(.din(n25150), .dout(n25153));
    jdff dff_B_oXm7oNef5_2(.din(n25153), .dout(n25156));
    jdff dff_B_CBNzjB7B2_2(.din(n25156), .dout(n25159));
    jdff dff_B_Syiaelsg1_2(.din(n25159), .dout(n25162));
    jdff dff_B_3zQJlg3H0_2(.din(n25162), .dout(n25165));
    jdff dff_B_JI51UZ669_2(.din(n25165), .dout(n25168));
    jdff dff_B_vzn2Bcph8_2(.din(n25168), .dout(n25171));
    jdff dff_B_ppiBzVLm1_2(.din(n25171), .dout(n25174));
    jdff dff_B_Mftj1Eta7_2(.din(n25174), .dout(n25177));
    jdff dff_B_O4UpiI2e8_2(.din(n25177), .dout(n25180));
    jdff dff_B_eRtSiULM4_2(.din(n25180), .dout(n25183));
    jdff dff_B_aspaOuBq0_2(.din(n25183), .dout(n25186));
    jdff dff_B_9a1SXeoi0_2(.din(n25186), .dout(n25189));
    jdff dff_B_lWuhQ7km8_2(.din(n25189), .dout(n25192));
    jdff dff_B_yP0Jf2nB5_2(.din(n25192), .dout(n25195));
    jdff dff_B_JNbSNTFf9_2(.din(n25195), .dout(n25198));
    jdff dff_B_mAJPjSWK4_2(.din(n25198), .dout(n25201));
    jdff dff_B_tcULOzcr5_2(.din(n25201), .dout(n25204));
    jdff dff_B_1pDKIZ093_2(.din(n25204), .dout(n25207));
    jdff dff_B_N2jdzGk90_2(.din(n6258), .dout(n25210));
    jdff dff_B_OD8zsOFz3_1(.din(n6250), .dout(n25213));
    jdff dff_B_Le2aNLXW1_2(.din(n6052), .dout(n25216));
    jdff dff_B_X940kKQk4_2(.din(n25216), .dout(n25219));
    jdff dff_B_WQWOCGvC2_2(.din(n25219), .dout(n25222));
    jdff dff_B_KKy3QRSz1_2(.din(n25222), .dout(n25225));
    jdff dff_B_Dbr6G2PZ9_2(.din(n25225), .dout(n25228));
    jdff dff_B_G0ADHMuC9_2(.din(n25228), .dout(n25231));
    jdff dff_B_oEcDhbXk8_2(.din(n25231), .dout(n25234));
    jdff dff_B_l0jqOEwI9_2(.din(n25234), .dout(n25237));
    jdff dff_B_NZYnER997_2(.din(n25237), .dout(n25240));
    jdff dff_B_9eFXj9rZ8_2(.din(n25240), .dout(n25243));
    jdff dff_B_lATkhR9x2_2(.din(n25243), .dout(n25246));
    jdff dff_B_fjW11Uiw8_2(.din(n25246), .dout(n25249));
    jdff dff_B_AWWjL4iO7_2(.din(n25249), .dout(n25252));
    jdff dff_B_9zkz70Iy8_2(.din(n25252), .dout(n25255));
    jdff dff_B_4JdnowO17_2(.din(n25255), .dout(n25258));
    jdff dff_B_PFUZM9UN2_2(.din(n25258), .dout(n25261));
    jdff dff_B_eNZAHqET7_2(.din(n25261), .dout(n25264));
    jdff dff_B_23GPd94w8_2(.din(n25264), .dout(n25267));
    jdff dff_B_U06PEwPw6_2(.din(n25267), .dout(n25270));
    jdff dff_B_svnKd5Hb2_2(.din(n25270), .dout(n25273));
    jdff dff_B_WolfQb4C1_2(.din(n25273), .dout(n25276));
    jdff dff_B_8sef5ni97_2(.din(n25276), .dout(n25279));
    jdff dff_B_COQEwRTS3_2(.din(n25279), .dout(n25282));
    jdff dff_B_eNKHHtb45_2(.din(n25282), .dout(n25285));
    jdff dff_B_vZM6LUyC7_2(.din(n25285), .dout(n25288));
    jdff dff_B_O9ovA19C0_2(.din(n25288), .dout(n25291));
    jdff dff_B_0ayl8ijC5_2(.din(n25291), .dout(n25294));
    jdff dff_B_B3NPte5y2_2(.din(n25294), .dout(n25297));
    jdff dff_B_pkTmhiov8_2(.din(n25297), .dout(n25300));
    jdff dff_B_bU4njUtF6_2(.din(n25300), .dout(n25303));
    jdff dff_B_h9EIukWF0_2(.din(n25303), .dout(n25306));
    jdff dff_B_Qh8KRF7c1_2(.din(n25306), .dout(n25309));
    jdff dff_B_MdxlzSYs3_2(.din(n25309), .dout(n25312));
    jdff dff_B_5ocVLUiB6_2(.din(n25312), .dout(n25315));
    jdff dff_B_qwmLDYlS5_2(.din(n25315), .dout(n25318));
    jdff dff_B_K8LkMMUf4_2(.din(n25318), .dout(n25321));
    jdff dff_B_3QpEcBYS5_2(.din(n25321), .dout(n25324));
    jdff dff_B_B68IbSmN4_2(.din(n25324), .dout(n25327));
    jdff dff_B_q2UG8rry9_2(.din(n25327), .dout(n25330));
    jdff dff_B_GWmTiUBi7_2(.din(n25330), .dout(n25333));
    jdff dff_B_6czhGHEI7_2(.din(n25333), .dout(n25336));
    jdff dff_B_0dWJxbfB1_2(.din(n25336), .dout(n25339));
    jdff dff_B_Wiglwtz19_2(.din(n25339), .dout(n25342));
    jdff dff_B_e4hHRO710_2(.din(n25342), .dout(n25345));
    jdff dff_B_t7NTSo022_2(.din(n25345), .dout(n25348));
    jdff dff_B_gEWZXbi90_2(.din(n6064), .dout(n25351));
    jdff dff_B_4DM503qx1_1(.din(n6056), .dout(n25354));
    jdff dff_B_XSj0W33P0_2(.din(n5834), .dout(n25357));
    jdff dff_B_mF69VJTT3_2(.din(n25357), .dout(n25360));
    jdff dff_B_ucASIHuc0_2(.din(n25360), .dout(n25363));
    jdff dff_B_Qftq9QV42_2(.din(n25363), .dout(n25366));
    jdff dff_B_et16hyLE3_2(.din(n25366), .dout(n25369));
    jdff dff_B_9Nd1Zc0o6_2(.din(n25369), .dout(n25372));
    jdff dff_B_QzZVqoBh7_2(.din(n25372), .dout(n25375));
    jdff dff_B_IkSMX9aT1_2(.din(n25375), .dout(n25378));
    jdff dff_B_vQHBgyYe9_2(.din(n25378), .dout(n25381));
    jdff dff_B_vvAv7Okf5_2(.din(n25381), .dout(n25384));
    jdff dff_B_5e5HsEMC4_2(.din(n25384), .dout(n25387));
    jdff dff_B_pEBgNAwd1_2(.din(n25387), .dout(n25390));
    jdff dff_B_Vuefmv1m0_2(.din(n25390), .dout(n25393));
    jdff dff_B_COoAiAtz7_2(.din(n25393), .dout(n25396));
    jdff dff_B_DnnAyAKx2_2(.din(n25396), .dout(n25399));
    jdff dff_B_muPSitCL1_2(.din(n25399), .dout(n25402));
    jdff dff_B_muLNuAq94_2(.din(n25402), .dout(n25405));
    jdff dff_B_CAX2kDuR4_2(.din(n25405), .dout(n25408));
    jdff dff_B_TWbd1d8b4_2(.din(n25408), .dout(n25411));
    jdff dff_B_JI8RnBij7_2(.din(n25411), .dout(n25414));
    jdff dff_B_p95ohL3o8_2(.din(n25414), .dout(n25417));
    jdff dff_B_TxH64Jd20_2(.din(n25417), .dout(n25420));
    jdff dff_B_vlsk8rsp8_2(.din(n25420), .dout(n25423));
    jdff dff_B_HWi3T1sR2_2(.din(n25423), .dout(n25426));
    jdff dff_B_syxz5Bew5_2(.din(n25426), .dout(n25429));
    jdff dff_B_ViomdNKI7_2(.din(n25429), .dout(n25432));
    jdff dff_B_B2IHkcjU0_2(.din(n25432), .dout(n25435));
    jdff dff_B_JFXiRL2v5_2(.din(n25435), .dout(n25438));
    jdff dff_B_qnOSOI3J0_2(.din(n25438), .dout(n25441));
    jdff dff_B_o0aGfLs23_2(.din(n25441), .dout(n25444));
    jdff dff_B_2ZGwtNOI0_2(.din(n25444), .dout(n25447));
    jdff dff_B_oYfWgQwj4_2(.din(n25447), .dout(n25450));
    jdff dff_B_vrHRwwY64_2(.din(n25450), .dout(n25453));
    jdff dff_B_w6MhnlCF4_2(.din(n25453), .dout(n25456));
    jdff dff_B_dLFBpsyn4_2(.din(n25456), .dout(n25459));
    jdff dff_B_lOrcylcN4_2(.din(n25459), .dout(n25462));
    jdff dff_B_NTf9Cb4h1_2(.din(n25462), .dout(n25465));
    jdff dff_B_1xK1Vb336_2(.din(n25465), .dout(n25468));
    jdff dff_B_k00PbxRh3_2(.din(n25468), .dout(n25471));
    jdff dff_B_shqddaeU0_2(.din(n25471), .dout(n25474));
    jdff dff_B_PlW01fJO6_2(.din(n25474), .dout(n25477));
    jdff dff_B_k6Z3dM301_2(.din(n5846), .dout(n25480));
    jdff dff_B_KWsj1w4I1_1(.din(n5838), .dout(n25483));
    jdff dff_B_fnADqmUn2_2(.din(n5589), .dout(n25486));
    jdff dff_B_HtyjzvXR0_2(.din(n25486), .dout(n25489));
    jdff dff_B_niEEAyfw3_2(.din(n25489), .dout(n25492));
    jdff dff_B_nkqB8I3H3_2(.din(n25492), .dout(n25495));
    jdff dff_B_MBEf3onO7_2(.din(n25495), .dout(n25498));
    jdff dff_B_xExIR2Qf8_2(.din(n25498), .dout(n25501));
    jdff dff_B_ZZj8lqqf6_2(.din(n25501), .dout(n25504));
    jdff dff_B_wDnhVLNH7_2(.din(n25504), .dout(n25507));
    jdff dff_B_N5r9Gnzo9_2(.din(n25507), .dout(n25510));
    jdff dff_B_dFgESHhn5_2(.din(n25510), .dout(n25513));
    jdff dff_B_I5XpsT1x0_2(.din(n25513), .dout(n25516));
    jdff dff_B_qxrLQuA97_2(.din(n25516), .dout(n25519));
    jdff dff_B_TwS7Su2d1_2(.din(n25519), .dout(n25522));
    jdff dff_B_TI4D2na19_2(.din(n25522), .dout(n25525));
    jdff dff_B_wdtrvRXi8_2(.din(n25525), .dout(n25528));
    jdff dff_B_GE6M4kkh9_2(.din(n25528), .dout(n25531));
    jdff dff_B_1v9xkd8r2_2(.din(n25531), .dout(n25534));
    jdff dff_B_c8p1SSMr9_2(.din(n25534), .dout(n25537));
    jdff dff_B_rG8uYtic6_2(.din(n25537), .dout(n25540));
    jdff dff_B_G2qFkAGH0_2(.din(n25540), .dout(n25543));
    jdff dff_B_BmlNWpeI1_2(.din(n25543), .dout(n25546));
    jdff dff_B_8s4SRJPV3_2(.din(n25546), .dout(n25549));
    jdff dff_B_hxYpHBWI4_2(.din(n25549), .dout(n25552));
    jdff dff_B_iqOqpiti7_2(.din(n25552), .dout(n25555));
    jdff dff_B_1ap5ySk98_2(.din(n25555), .dout(n25558));
    jdff dff_B_ThBV1DCF0_2(.din(n25558), .dout(n25561));
    jdff dff_B_7iAodSeq2_2(.din(n25561), .dout(n25564));
    jdff dff_B_wopjOCEN2_2(.din(n25564), .dout(n25567));
    jdff dff_B_1WI3EKo63_2(.din(n25567), .dout(n25570));
    jdff dff_B_NR4hBKQh4_2(.din(n25570), .dout(n25573));
    jdff dff_B_G5gHnXfc5_2(.din(n25573), .dout(n25576));
    jdff dff_B_QN5lWEbu1_2(.din(n25576), .dout(n25579));
    jdff dff_B_hL6rvXJP4_2(.din(n25579), .dout(n25582));
    jdff dff_B_Xcz8bQt79_2(.din(n25582), .dout(n25585));
    jdff dff_B_lrITYiHD2_2(.din(n25585), .dout(n25588));
    jdff dff_B_BHbMM9XM6_2(.din(n25588), .dout(n25591));
    jdff dff_B_2q0oM0jv1_2(.din(n25591), .dout(n25594));
    jdff dff_B_f4y5ryhm3_2(.din(n5601), .dout(n25597));
    jdff dff_B_QlXDA0Gs6_1(.din(n5593), .dout(n25600));
    jdff dff_B_HFuURorS5_2(.din(n5317), .dout(n25603));
    jdff dff_B_HYtwev9K1_2(.din(n25603), .dout(n25606));
    jdff dff_B_jsr3QjnB4_2(.din(n25606), .dout(n25609));
    jdff dff_B_KLGBzTgE6_2(.din(n25609), .dout(n25612));
    jdff dff_B_6ChZadHj3_2(.din(n25612), .dout(n25615));
    jdff dff_B_UbqCyEjC9_2(.din(n25615), .dout(n25618));
    jdff dff_B_Hhwahzwe4_2(.din(n25618), .dout(n25621));
    jdff dff_B_2iJvjgP80_2(.din(n25621), .dout(n25624));
    jdff dff_B_0rAaLXo55_2(.din(n25624), .dout(n25627));
    jdff dff_B_WKRz6zFz4_2(.din(n25627), .dout(n25630));
    jdff dff_B_mYj8hEJG2_2(.din(n25630), .dout(n25633));
    jdff dff_B_2tDofd421_2(.din(n25633), .dout(n25636));
    jdff dff_B_BrDCQca44_2(.din(n25636), .dout(n25639));
    jdff dff_B_ovWFeDIW3_2(.din(n25639), .dout(n25642));
    jdff dff_B_UFvFRXVG7_2(.din(n25642), .dout(n25645));
    jdff dff_B_dWjQTx6d2_2(.din(n25645), .dout(n25648));
    jdff dff_B_Z1pQawyx2_2(.din(n25648), .dout(n25651));
    jdff dff_B_2Mws1gYY1_2(.din(n25651), .dout(n25654));
    jdff dff_B_tviATJVO9_2(.din(n25654), .dout(n25657));
    jdff dff_B_GTeB3NYr8_2(.din(n25657), .dout(n25660));
    jdff dff_B_Y6j6lNRV8_2(.din(n25660), .dout(n25663));
    jdff dff_B_unFGG66d8_2(.din(n25663), .dout(n25666));
    jdff dff_B_7aIpXPD49_2(.din(n25666), .dout(n25669));
    jdff dff_B_V2ISwFEN5_2(.din(n25669), .dout(n25672));
    jdff dff_B_LJw5olb82_2(.din(n25672), .dout(n25675));
    jdff dff_B_Fx76HhxW5_2(.din(n25675), .dout(n25678));
    jdff dff_B_0u5xo9Bq9_2(.din(n25678), .dout(n25681));
    jdff dff_B_GmD0ky7j3_2(.din(n25681), .dout(n25684));
    jdff dff_B_n9K19JA90_2(.din(n25684), .dout(n25687));
    jdff dff_B_fMOdFGYu5_2(.din(n25687), .dout(n25690));
    jdff dff_B_y2k1Dz5Y5_2(.din(n25690), .dout(n25693));
    jdff dff_B_ogX3M0e88_2(.din(n25693), .dout(n25696));
    jdff dff_B_NIiP5MnK3_2(.din(n25696), .dout(n25699));
    jdff dff_B_0Ke26RMA9_1(.din(n5321), .dout(n25702));
    jdff dff_B_zdur0rHx6_2(.din(n5018), .dout(n25705));
    jdff dff_B_NHoRZHjM0_2(.din(n25705), .dout(n25708));
    jdff dff_B_8SYQqcns8_2(.din(n25708), .dout(n25711));
    jdff dff_B_YBcxg5414_2(.din(n25711), .dout(n25714));
    jdff dff_B_erQ4fIHP6_2(.din(n25714), .dout(n25717));
    jdff dff_B_4PuvGxbi5_2(.din(n25717), .dout(n25720));
    jdff dff_B_HMFb1ltr6_2(.din(n25720), .dout(n25723));
    jdff dff_B_Ife0iku81_2(.din(n25723), .dout(n25726));
    jdff dff_B_f8cjXL9Z2_2(.din(n25726), .dout(n25729));
    jdff dff_B_UiOIbgrz5_2(.din(n25729), .dout(n25732));
    jdff dff_B_7jUvcbn46_2(.din(n25732), .dout(n25735));
    jdff dff_B_EVeQGmWW3_2(.din(n25735), .dout(n25738));
    jdff dff_B_H9Ffuray3_2(.din(n25738), .dout(n25741));
    jdff dff_B_3akg4uhZ2_2(.din(n25741), .dout(n25744));
    jdff dff_B_qlAL7DbF5_2(.din(n25744), .dout(n25747));
    jdff dff_B_rcyTbpPx5_2(.din(n25747), .dout(n25750));
    jdff dff_B_Egp1LORW2_2(.din(n25750), .dout(n25753));
    jdff dff_B_W59M4nOI8_2(.din(n25753), .dout(n25756));
    jdff dff_B_bxryLyCT7_2(.din(n25756), .dout(n25759));
    jdff dff_B_7WUGfm5W9_2(.din(n25759), .dout(n25762));
    jdff dff_B_4Lb1V7ce6_2(.din(n25762), .dout(n25765));
    jdff dff_B_VoDIUlxA7_2(.din(n25765), .dout(n25768));
    jdff dff_B_XTgZh5318_2(.din(n25768), .dout(n25771));
    jdff dff_B_CL2iF2yL3_2(.din(n25771), .dout(n25774));
    jdff dff_B_k9owATDD3_2(.din(n25774), .dout(n25777));
    jdff dff_B_iyU4cppo5_2(.din(n25777), .dout(n25780));
    jdff dff_B_MsQzurds4_2(.din(n25780), .dout(n25783));
    jdff dff_B_TTTi2UUd8_2(.din(n25783), .dout(n25786));
    jdff dff_B_WJEV09jc6_2(.din(n25786), .dout(n25789));
    jdff dff_B_iqpIQTzU2_2(.din(n25789), .dout(n25792));
    jdff dff_B_2gb9Bxer1_2(.din(n5142), .dout(n25795));
    jdff dff_B_jkB5FMPY5_1(.din(n5022), .dout(n25798));
    jdff dff_B_EHNiVPGa5_2(.din(n4692), .dout(n25801));
    jdff dff_B_R53KKUYP0_2(.din(n25801), .dout(n25804));
    jdff dff_B_cZjVBzQE5_2(.din(n25804), .dout(n25807));
    jdff dff_B_4j4JNBkS9_2(.din(n25807), .dout(n25810));
    jdff dff_B_qudDM4mX8_2(.din(n25810), .dout(n25813));
    jdff dff_B_I2hQy2mV6_2(.din(n25813), .dout(n25816));
    jdff dff_B_GUVxetKd4_2(.din(n25816), .dout(n25819));
    jdff dff_B_WlH3N3xI3_2(.din(n25819), .dout(n25822));
    jdff dff_B_qaD0liny8_2(.din(n25822), .dout(n25825));
    jdff dff_B_pskPLXQP5_2(.din(n25825), .dout(n25828));
    jdff dff_B_RY5mHMTT7_2(.din(n25828), .dout(n25831));
    jdff dff_B_w31ARI7p5_2(.din(n25831), .dout(n25834));
    jdff dff_B_q0iaNeqA5_2(.din(n25834), .dout(n25837));
    jdff dff_B_Ktf7kmeC2_2(.din(n25837), .dout(n25840));
    jdff dff_B_DQnPTe6U1_2(.din(n25840), .dout(n25843));
    jdff dff_B_s3baH0L16_2(.din(n25843), .dout(n25846));
    jdff dff_B_smTXGo765_2(.din(n25846), .dout(n25849));
    jdff dff_B_wqyk9ScC3_2(.din(n25849), .dout(n25852));
    jdff dff_B_MOC4qZHb7_2(.din(n25852), .dout(n25855));
    jdff dff_B_ypz8S9Q79_2(.din(n25855), .dout(n25858));
    jdff dff_B_NMepsmpw3_2(.din(n25858), .dout(n25861));
    jdff dff_B_mbJAJiPN0_2(.din(n25861), .dout(n25864));
    jdff dff_B_yLgDWa1g2_2(.din(n25864), .dout(n25867));
    jdff dff_B_DO6sKrzx2_2(.din(n25867), .dout(n25870));
    jdff dff_B_SnAK9J960_2(.din(n25870), .dout(n25873));
    jdff dff_B_EeLLnJ7g4_2(.din(n25873), .dout(n25876));
    jdff dff_B_1Klk0tMV1_2(.din(n25876), .dout(n25879));
    jdff dff_B_OyczPD237_2(.din(n4816), .dout(n25882));
    jdff dff_B_IZsyeWf28_1(.din(n4696), .dout(n25885));
    jdff dff_B_L1gaHzF19_2(.din(n4346), .dout(n25888));
    jdff dff_B_cihPYqz81_2(.din(n25888), .dout(n25891));
    jdff dff_B_GbGbOR9e9_2(.din(n25891), .dout(n25894));
    jdff dff_B_zOOFACYH8_2(.din(n25894), .dout(n25897));
    jdff dff_B_NrA7s80c8_2(.din(n25897), .dout(n25900));
    jdff dff_B_HsfuJafL4_2(.din(n25900), .dout(n25903));
    jdff dff_B_z8Spxi6f9_2(.din(n25903), .dout(n25906));
    jdff dff_B_TMGb5HZq1_2(.din(n25906), .dout(n25909));
    jdff dff_B_icSf5HTl1_2(.din(n25909), .dout(n25912));
    jdff dff_B_EAbTJmvu8_2(.din(n25912), .dout(n25915));
    jdff dff_B_MqnxQ0SH0_2(.din(n25915), .dout(n25918));
    jdff dff_B_TTRDu9L52_2(.din(n25918), .dout(n25921));
    jdff dff_B_UTsSfrOG5_2(.din(n25921), .dout(n25924));
    jdff dff_B_YY5hh0fQ9_2(.din(n25924), .dout(n25927));
    jdff dff_B_DhV318ib4_2(.din(n25927), .dout(n25930));
    jdff dff_B_Lf99Nr2G0_2(.din(n25930), .dout(n25933));
    jdff dff_B_GMR7TjrY2_2(.din(n25933), .dout(n25936));
    jdff dff_B_JLZtvhgW5_2(.din(n25936), .dout(n25939));
    jdff dff_B_ih9TGE8T8_2(.din(n25939), .dout(n25942));
    jdff dff_B_2WOqcq8D2_2(.din(n25942), .dout(n25945));
    jdff dff_B_NxtaKpLL8_2(.din(n25945), .dout(n25948));
    jdff dff_B_2FGWKC1H9_2(.din(n25948), .dout(n25951));
    jdff dff_B_uomZ3BfG8_2(.din(n25951), .dout(n25954));
    jdff dff_B_vuesWQg10_2(.din(n25954), .dout(n25957));
    jdff dff_B_0ln7i3yv3_2(.din(n4466), .dout(n25960));
    jdff dff_B_teh9vl1E7_1(.din(n4350), .dout(n25963));
    jdff dff_B_52OESfC01_2(.din(n3950), .dout(n25966));
    jdff dff_B_nySWuDaB3_2(.din(n25966), .dout(n25969));
    jdff dff_B_0j5IJlxb1_2(.din(n25969), .dout(n25972));
    jdff dff_B_xUnWSZUa1_2(.din(n25972), .dout(n25975));
    jdff dff_B_q6Jh4Fqk1_2(.din(n25975), .dout(n25978));
    jdff dff_B_VqFUs14A8_2(.din(n25978), .dout(n25981));
    jdff dff_B_PEclydIw9_2(.din(n25981), .dout(n25984));
    jdff dff_B_dwJuQe8d3_2(.din(n25984), .dout(n25987));
    jdff dff_B_bEUvZqBd9_2(.din(n25987), .dout(n25990));
    jdff dff_B_kn7fbtFZ0_2(.din(n25990), .dout(n25993));
    jdff dff_B_LARXZbmT2_2(.din(n25993), .dout(n25996));
    jdff dff_B_6HOxNdgJ9_2(.din(n25996), .dout(n25999));
    jdff dff_B_aX6E68Rs5_2(.din(n25999), .dout(n26002));
    jdff dff_B_IfY7yqZW1_2(.din(n26002), .dout(n26005));
    jdff dff_B_qxKB7DB39_2(.din(n26005), .dout(n26008));
    jdff dff_B_KBa7162e0_2(.din(n26008), .dout(n26011));
    jdff dff_B_KHTrgNUI6_2(.din(n26011), .dout(n26014));
    jdff dff_B_iNU01zlk3_2(.din(n26014), .dout(n26017));
    jdff dff_B_Y66iCzaW2_2(.din(n26017), .dout(n26020));
    jdff dff_B_FIAq9V0Q4_2(.din(n26020), .dout(n26023));
    jdff dff_B_F7lIEWSj0_2(.din(n26023), .dout(n26026));
    jdff dff_B_HKVoNoEe3_2(.din(n4090), .dout(n26029));
    jdff dff_B_g9P1r5ym0_1(.din(n3954), .dout(n26032));
    jdff dff_B_xiWu0dwT2_2(.din(n3573), .dout(n26035));
    jdff dff_B_YHrjbzBw9_2(.din(n26035), .dout(n26038));
    jdff dff_B_LEWog6le3_2(.din(n26038), .dout(n26041));
    jdff dff_B_gx8vGpJf7_2(.din(n26041), .dout(n26044));
    jdff dff_B_iXjk25ko9_2(.din(n26044), .dout(n26047));
    jdff dff_B_QmnEWcnm7_2(.din(n26047), .dout(n26050));
    jdff dff_B_Tk30aquB3_2(.din(n26050), .dout(n26053));
    jdff dff_B_XUzeh79p2_2(.din(n26053), .dout(n26056));
    jdff dff_B_9RsS1pdi9_2(.din(n26056), .dout(n26059));
    jdff dff_B_PvucHwYW2_2(.din(n26059), .dout(n26062));
    jdff dff_B_aHsH2MyB5_2(.din(n26062), .dout(n26065));
    jdff dff_B_dlJ8ddlK4_2(.din(n26065), .dout(n26068));
    jdff dff_B_xtYAbrtG5_2(.din(n26068), .dout(n26071));
    jdff dff_B_ic7GWx239_2(.din(n26071), .dout(n26074));
    jdff dff_B_ezXa3Q176_2(.din(n26074), .dout(n26077));
    jdff dff_B_M7KNXDcu3_2(.din(n26077), .dout(n26080));
    jdff dff_B_E60SA92c5_2(.din(n26080), .dout(n26083));
    jdff dff_B_A61RqbDr9_2(.din(n26083), .dout(n26086));
    jdff dff_B_RcsfpYi26_2(.din(n3687), .dout(n26089));
    jdff dff_B_nYni0s4q4_1(.din(n3577), .dout(n26092));
    jdff dff_B_16wA4Tok1_2(.din(n3172), .dout(n26095));
    jdff dff_B_HcoFhwj94_2(.din(n26095), .dout(n26098));
    jdff dff_B_ssb5h6nL8_2(.din(n26098), .dout(n26101));
    jdff dff_B_WhAQoRf68_2(.din(n26101), .dout(n26104));
    jdff dff_B_1W6cgkrg1_2(.din(n26104), .dout(n26107));
    jdff dff_B_qcw6OwS11_2(.din(n26107), .dout(n26110));
    jdff dff_B_eBYhpD1m0_2(.din(n26110), .dout(n26113));
    jdff dff_B_5Y0gQePj7_2(.din(n26113), .dout(n26116));
    jdff dff_B_gqcx2evk1_2(.din(n26116), .dout(n26119));
    jdff dff_B_rmOU3GDN6_2(.din(n26119), .dout(n26122));
    jdff dff_B_z7giTpya6_2(.din(n26122), .dout(n26125));
    jdff dff_B_Z3acxj7O5_2(.din(n26125), .dout(n26128));
    jdff dff_B_SG9yeJir4_2(.din(n26128), .dout(n26131));
    jdff dff_B_f9xz1iH55_2(.din(n26131), .dout(n26134));
    jdff dff_B_JmAnH8nQ3_2(.din(n26134), .dout(n26137));
    jdff dff_B_Lcdxw4Xr7_2(.din(n3285), .dout(n26140));
    jdff dff_B_6TftSVYF7_1(.din(n3176), .dout(n26143));
    jdff dff_B_fOZFgnN18_2(.din(n2793), .dout(n26146));
    jdff dff_B_J6dWZeOp2_2(.din(n26146), .dout(n26149));
    jdff dff_B_NEtTj2Mq9_2(.din(n26149), .dout(n26152));
    jdff dff_B_S3EBGOoQ6_2(.din(n26152), .dout(n26155));
    jdff dff_B_y1VeWTxt8_2(.din(n26155), .dout(n26158));
    jdff dff_B_jOoHe2UU8_2(.din(n26158), .dout(n26161));
    jdff dff_B_gsI5fYDQ3_2(.din(n26161), .dout(n26164));
    jdff dff_B_NBf5rh7b4_2(.din(n26164), .dout(n26167));
    jdff dff_B_OydbojVv2_2(.din(n26167), .dout(n26170));
    jdff dff_B_XepdfhXy6_2(.din(n26170), .dout(n26173));
    jdff dff_B_r2F1US2v5_2(.din(n26173), .dout(n26176));
    jdff dff_B_Fx7TQE1T8_2(.din(n26176), .dout(n26179));
    jdff dff_B_tWtJj8lm3_2(.din(n2880), .dout(n26182));
    jdff dff_B_R12el6iH1_1(.din(n2797), .dout(n26185));
    jdff dff_B_tdkRVyET1_2(.din(n2438), .dout(n26188));
    jdff dff_B_Dw7Hi8SV3_2(.din(n26188), .dout(n26191));
    jdff dff_B_frbER5xA9_2(.din(n26191), .dout(n26194));
    jdff dff_B_rmnmQTaV7_2(.din(n26194), .dout(n26197));
    jdff dff_B_qIGRpHMu2_2(.din(n26197), .dout(n26200));
    jdff dff_B_3QBsWR8H1_2(.din(n26200), .dout(n26203));
    jdff dff_B_zqHIAowd4_2(.din(n26203), .dout(n26206));
    jdff dff_B_y05Obsgc0_2(.din(n26206), .dout(n26209));
    jdff dff_B_PumEGzma6_2(.din(n26209), .dout(n26212));
    jdff dff_B_yd2VpjQb7_2(.din(n2498), .dout(n26215));
    jdff dff_B_GTmP2KeA8_2(.din(n26215), .dout(n26218));
    jdff dff_B_Y7u0ICTY3_1(.din(n2441), .dout(n26221));
    jdff dff_B_vMOoao6P2_1(.din(n26221), .dout(n26224));
    jdff dff_B_6wM3bMd49_1(.din(n26224), .dout(n26227));
    jdff dff_B_GKLQP4Ta8_1(.din(n26227), .dout(n26230));
    jdff dff_B_pEl37SFF6_1(.din(n26230), .dout(n26233));
    jdff dff_B_w4rI4dlB8_1(.din(n26233), .dout(n26236));
    jdff dff_B_uvHwSihO4_0(.din(n2143), .dout(n26239));
    jdff dff_B_yeWItqQb4_0(.din(n26239), .dout(n26242));
    jdff dff_A_sMSki8O07_0(.din(n26247), .dout(n26244));
    jdff dff_A_mV1ETtr76_0(.din(n26250), .dout(n26247));
    jdff dff_A_DwgwG6gr1_0(.din(n2139), .dout(n26250));
    jdff dff_B_wtlWOni45_1(.din(n2117), .dout(n26254));
    jdff dff_A_8UhmKZc75_0(.din(n1805), .dout(n26256));
    jdff dff_A_TaYnXwFq7_1(.din(n26262), .dout(n26259));
    jdff dff_A_NfLo46A38_1(.din(n1805), .dout(n26262));
    jdff dff_A_lD78zEp75_1(.din(n26268), .dout(n26265));
    jdff dff_A_iRN75Ff71_1(.din(n26271), .dout(n26268));
    jdff dff_A_U1GsVckW9_1(.din(n26274), .dout(n26271));
    jdff dff_A_kf5tlb256_1(.din(n26277), .dout(n26274));
    jdff dff_A_9RwiuLbM9_1(.din(n26280), .dout(n26277));
    jdff dff_A_7lPIcV558_1(.din(n2109), .dout(n26280));
    jdff dff_B_swAYl7xU4_1(.din(n6665), .dout(n26284));
    jdff dff_A_WItlfLpC4_1(.din(n6569), .dout(n26286));
    jdff dff_B_LzPbpWEu3_1(.din(n6561), .dout(n26290));
    jdff dff_B_H6mtBv1K6_2(.din(n6423), .dout(n26293));
    jdff dff_B_9XvtSTpv6_2(.din(n26293), .dout(n26296));
    jdff dff_B_yb1kLai44_2(.din(n26296), .dout(n26299));
    jdff dff_B_9JzcRiYJ3_2(.din(n26299), .dout(n26302));
    jdff dff_B_kdxV89qc4_2(.din(n26302), .dout(n26305));
    jdff dff_B_1nr48IKx1_2(.din(n26305), .dout(n26308));
    jdff dff_B_anXGj3Lk6_2(.din(n26308), .dout(n26311));
    jdff dff_B_gP6AfZ4R5_2(.din(n26311), .dout(n26314));
    jdff dff_B_l7rqyiSV9_2(.din(n26314), .dout(n26317));
    jdff dff_B_ShfQ0cvR2_2(.din(n26317), .dout(n26320));
    jdff dff_B_svNpG9i57_2(.din(n26320), .dout(n26323));
    jdff dff_B_xp2N5JwY0_2(.din(n26323), .dout(n26326));
    jdff dff_B_jlivo5LI9_2(.din(n26326), .dout(n26329));
    jdff dff_B_ej2HIOCH3_2(.din(n26329), .dout(n26332));
    jdff dff_B_6jU6beEu7_2(.din(n26332), .dout(n26335));
    jdff dff_B_aEVKyXID7_2(.din(n26335), .dout(n26338));
    jdff dff_B_ZU662TJJ7_2(.din(n26338), .dout(n26341));
    jdff dff_B_4qnuRD3s8_2(.din(n26341), .dout(n26344));
    jdff dff_B_9Gx5wGeG1_2(.din(n26344), .dout(n26347));
    jdff dff_B_Yo0Vf7SH7_2(.din(n26347), .dout(n26350));
    jdff dff_B_LbMODvhb2_2(.din(n26350), .dout(n26353));
    jdff dff_B_wrDSOEST9_2(.din(n26353), .dout(n26356));
    jdff dff_B_EIvnxcR78_2(.din(n26356), .dout(n26359));
    jdff dff_B_5v8GyuaA4_2(.din(n26359), .dout(n26362));
    jdff dff_B_Yhoexs5x1_2(.din(n26362), .dout(n26365));
    jdff dff_B_OrtWqyKA3_2(.din(n26365), .dout(n26368));
    jdff dff_B_tgn7m4K28_2(.din(n26368), .dout(n26371));
    jdff dff_B_yJcC1C7Q1_2(.din(n26371), .dout(n26374));
    jdff dff_B_UPcYNmSS2_2(.din(n26374), .dout(n26377));
    jdff dff_B_RIwApUQW6_2(.din(n26377), .dout(n26380));
    jdff dff_B_bQfhKYo91_2(.din(n26380), .dout(n26383));
    jdff dff_B_fMkyXAsr2_2(.din(n26383), .dout(n26386));
    jdff dff_B_zsGQLSGN9_2(.din(n26386), .dout(n26389));
    jdff dff_B_9FlxtoOI5_2(.din(n26389), .dout(n26392));
    jdff dff_B_IQdKcivU4_2(.din(n26392), .dout(n26395));
    jdff dff_B_CUKrA4Cw9_2(.din(n26395), .dout(n26398));
    jdff dff_B_Y9PhFo438_2(.din(n26398), .dout(n26401));
    jdff dff_B_LzbBETMS3_2(.din(n26401), .dout(n26404));
    jdff dff_B_957WxHNJ7_2(.din(n26404), .dout(n26407));
    jdff dff_B_rqZ2L9jc4_2(.din(n26407), .dout(n26410));
    jdff dff_B_tdgePMaP4_2(.din(n26410), .dout(n26413));
    jdff dff_B_gUyDHGLI0_2(.din(n26413), .dout(n26416));
    jdff dff_B_9MgmbgsI1_2(.din(n26416), .dout(n26419));
    jdff dff_B_syFGDCgS1_2(.din(n26419), .dout(n26422));
    jdff dff_B_utdgoEAV1_2(.din(n26422), .dout(n26425));
    jdff dff_B_YSxTucuZ5_2(.din(n26425), .dout(n26428));
    jdff dff_B_j7cEDYbT1_2(.din(n26428), .dout(n26431));
    jdff dff_B_wcq1zbGT0_2(.din(n26431), .dout(n26434));
    jdff dff_B_umlEhmbA0_2(.din(n26434), .dout(n26437));
    jdff dff_B_8T0UyFxb2_2(.din(n26437), .dout(n26440));
    jdff dff_B_xe0e7oJ50_2(.din(n26440), .dout(n26443));
    jdff dff_B_bUQI7BuH1_2(.din(n6435), .dout(n26446));
    jdff dff_B_cbqqkSOt3_1(.din(n6427), .dout(n26449));
    jdff dff_B_4WuJtOWd5_2(.din(n6265), .dout(n26452));
    jdff dff_B_YOyTYtVv5_2(.din(n26452), .dout(n26455));
    jdff dff_B_d9tLDOwU8_2(.din(n26455), .dout(n26458));
    jdff dff_B_BqLPgxoY5_2(.din(n26458), .dout(n26461));
    jdff dff_B_a0WegON35_2(.din(n26461), .dout(n26464));
    jdff dff_B_0Z9Q4Un26_2(.din(n26464), .dout(n26467));
    jdff dff_B_N1F4fEdb1_2(.din(n26467), .dout(n26470));
    jdff dff_B_eTMkIJLa1_2(.din(n26470), .dout(n26473));
    jdff dff_B_djqRUxpN1_2(.din(n26473), .dout(n26476));
    jdff dff_B_o3iJ7W9p2_2(.din(n26476), .dout(n26479));
    jdff dff_B_QkBUDKmJ9_2(.din(n26479), .dout(n26482));
    jdff dff_B_HMeZxEat8_2(.din(n26482), .dout(n26485));
    jdff dff_B_VgB0xkrC5_2(.din(n26485), .dout(n26488));
    jdff dff_B_edFqKEm53_2(.din(n26488), .dout(n26491));
    jdff dff_B_fH4Oxttf8_2(.din(n26491), .dout(n26494));
    jdff dff_B_NOTK3CBt7_2(.din(n26494), .dout(n26497));
    jdff dff_B_dPVSB4Nc7_2(.din(n26497), .dout(n26500));
    jdff dff_B_aFdUhKba3_2(.din(n26500), .dout(n26503));
    jdff dff_B_qMp8mdia4_2(.din(n26503), .dout(n26506));
    jdff dff_B_RoXPRaTS4_2(.din(n26506), .dout(n26509));
    jdff dff_B_bJhY5KSt2_2(.din(n26509), .dout(n26512));
    jdff dff_B_EZ6E0mIH9_2(.din(n26512), .dout(n26515));
    jdff dff_B_LiOHpp0s8_2(.din(n26515), .dout(n26518));
    jdff dff_B_UvNqbsXi3_2(.din(n26518), .dout(n26521));
    jdff dff_B_ZYkrU6122_2(.din(n26521), .dout(n26524));
    jdff dff_B_kyw1KR4g9_2(.din(n26524), .dout(n26527));
    jdff dff_B_P62hqi5Z4_2(.din(n26527), .dout(n26530));
    jdff dff_B_txPKKbPr8_2(.din(n26530), .dout(n26533));
    jdff dff_B_41AylPxe4_2(.din(n26533), .dout(n26536));
    jdff dff_B_mOKvSalK5_2(.din(n26536), .dout(n26539));
    jdff dff_B_z47xiuzn1_2(.din(n26539), .dout(n26542));
    jdff dff_B_K2Habuhe4_2(.din(n26542), .dout(n26545));
    jdff dff_B_KRwvONfS6_2(.din(n26545), .dout(n26548));
    jdff dff_B_3NSyxBTa3_2(.din(n26548), .dout(n26551));
    jdff dff_B_ExW8D8dv7_2(.din(n26551), .dout(n26554));
    jdff dff_B_GnmsHfMT3_2(.din(n26554), .dout(n26557));
    jdff dff_B_GJ6aRfhb6_2(.din(n26557), .dout(n26560));
    jdff dff_B_yQM7XMqw2_2(.din(n26560), .dout(n26563));
    jdff dff_B_vBvVXIyN1_2(.din(n26563), .dout(n26566));
    jdff dff_B_EN9LNgMC8_2(.din(n26566), .dout(n26569));
    jdff dff_B_sg1tNUUs7_2(.din(n26569), .dout(n26572));
    jdff dff_B_FcxZ8jjA7_2(.din(n26572), .dout(n26575));
    jdff dff_B_Z0iUD3KS2_2(.din(n26575), .dout(n26578));
    jdff dff_B_GnLQSwgO7_2(.din(n26578), .dout(n26581));
    jdff dff_B_mYHW4hAb0_2(.din(n26581), .dout(n26584));
    jdff dff_B_5F8Eq4700_2(.din(n26584), .dout(n26587));
    jdff dff_B_nj4zgaFg1_2(.din(n26587), .dout(n26590));
    jdff dff_B_jVVl5q6J8_2(.din(n6277), .dout(n26593));
    jdff dff_B_YNu2zp3w3_1(.din(n6269), .dout(n26596));
    jdff dff_B_TUQ9DmFl3_2(.din(n6071), .dout(n26599));
    jdff dff_B_2OdILCNc6_2(.din(n26599), .dout(n26602));
    jdff dff_B_OjvU5On85_2(.din(n26602), .dout(n26605));
    jdff dff_B_mLQhD9fW2_2(.din(n26605), .dout(n26608));
    jdff dff_B_oWwDZk5Y7_2(.din(n26608), .dout(n26611));
    jdff dff_B_GoOhqLBZ2_2(.din(n26611), .dout(n26614));
    jdff dff_B_eizSrCK38_2(.din(n26614), .dout(n26617));
    jdff dff_B_bcoynlxS0_2(.din(n26617), .dout(n26620));
    jdff dff_B_3A4MX6ls7_2(.din(n26620), .dout(n26623));
    jdff dff_B_tWhHESrw8_2(.din(n26623), .dout(n26626));
    jdff dff_B_VIfc0kX26_2(.din(n26626), .dout(n26629));
    jdff dff_B_zEMQBD2f6_2(.din(n26629), .dout(n26632));
    jdff dff_B_BKvZJwyW9_2(.din(n26632), .dout(n26635));
    jdff dff_B_yNQHINSw0_2(.din(n26635), .dout(n26638));
    jdff dff_B_qfR2ewqZ8_2(.din(n26638), .dout(n26641));
    jdff dff_B_K5ZmDyLb1_2(.din(n26641), .dout(n26644));
    jdff dff_B_0YAJk6Uj1_2(.din(n26644), .dout(n26647));
    jdff dff_B_z8BhNc4j2_2(.din(n26647), .dout(n26650));
    jdff dff_B_Y3ZIg1M75_2(.din(n26650), .dout(n26653));
    jdff dff_B_YSqnfV811_2(.din(n26653), .dout(n26656));
    jdff dff_B_ai8j6rzt5_2(.din(n26656), .dout(n26659));
    jdff dff_B_a98vFQd63_2(.din(n26659), .dout(n26662));
    jdff dff_B_CsJ1R2Tr4_2(.din(n26662), .dout(n26665));
    jdff dff_B_aDMptzkZ5_2(.din(n26665), .dout(n26668));
    jdff dff_B_ZLN7o7mO9_2(.din(n26668), .dout(n26671));
    jdff dff_B_W97JhkRO2_2(.din(n26671), .dout(n26674));
    jdff dff_B_GUzZIFy88_2(.din(n26674), .dout(n26677));
    jdff dff_B_5vcJ02eG7_2(.din(n26677), .dout(n26680));
    jdff dff_B_LgymVEUt2_2(.din(n26680), .dout(n26683));
    jdff dff_B_SrU3J8Tn8_2(.din(n26683), .dout(n26686));
    jdff dff_B_90hJe6is0_2(.din(n26686), .dout(n26689));
    jdff dff_B_An0iTvcV8_2(.din(n26689), .dout(n26692));
    jdff dff_B_CV5w5Dn94_2(.din(n26692), .dout(n26695));
    jdff dff_B_TMIYBPzl7_2(.din(n26695), .dout(n26698));
    jdff dff_B_GfeaITEK3_2(.din(n26698), .dout(n26701));
    jdff dff_B_o6gHOwCh1_2(.din(n26701), .dout(n26704));
    jdff dff_B_N1nDXXcd8_2(.din(n26704), .dout(n26707));
    jdff dff_B_X9SB6rxh9_2(.din(n26707), .dout(n26710));
    jdff dff_B_AvYioCkM2_2(.din(n26710), .dout(n26713));
    jdff dff_B_9ONkPx6P2_2(.din(n26713), .dout(n26716));
    jdff dff_B_sS0vzrBr8_2(.din(n26716), .dout(n26719));
    jdff dff_B_hSEr7CFm3_2(.din(n26719), .dout(n26722));
    jdff dff_B_gg96ixUT7_2(.din(n26722), .dout(n26725));
    jdff dff_B_RlKTCuxy7_2(.din(n6083), .dout(n26728));
    jdff dff_B_jPDNsV4f5_1(.din(n6075), .dout(n26731));
    jdff dff_B_FWhxwsyp1_2(.din(n5853), .dout(n26734));
    jdff dff_B_hN6NoHL09_2(.din(n26734), .dout(n26737));
    jdff dff_B_LmcKsD8k2_2(.din(n26737), .dout(n26740));
    jdff dff_B_HEZbZo4H0_2(.din(n26740), .dout(n26743));
    jdff dff_B_a5JieUma1_2(.din(n26743), .dout(n26746));
    jdff dff_B_SZllBtwh5_2(.din(n26746), .dout(n26749));
    jdff dff_B_CWE7WaOw3_2(.din(n26749), .dout(n26752));
    jdff dff_B_T5ucWDJP3_2(.din(n26752), .dout(n26755));
    jdff dff_B_vUhUwuC36_2(.din(n26755), .dout(n26758));
    jdff dff_B_qWV9Z5bT0_2(.din(n26758), .dout(n26761));
    jdff dff_B_S8Pv2Su02_2(.din(n26761), .dout(n26764));
    jdff dff_B_vTyWXmq13_2(.din(n26764), .dout(n26767));
    jdff dff_B_bPFVtFv45_2(.din(n26767), .dout(n26770));
    jdff dff_B_N6U4zmN03_2(.din(n26770), .dout(n26773));
    jdff dff_B_SSUob3hE8_2(.din(n26773), .dout(n26776));
    jdff dff_B_NT6MnoK61_2(.din(n26776), .dout(n26779));
    jdff dff_B_5oPMN6Tr6_2(.din(n26779), .dout(n26782));
    jdff dff_B_fIFqLAVR8_2(.din(n26782), .dout(n26785));
    jdff dff_B_A35TbZZY1_2(.din(n26785), .dout(n26788));
    jdff dff_B_TuHtGioY2_2(.din(n26788), .dout(n26791));
    jdff dff_B_EenB9Ik38_2(.din(n26791), .dout(n26794));
    jdff dff_B_zcY1HmAm6_2(.din(n26794), .dout(n26797));
    jdff dff_B_9DLkRjS03_2(.din(n26797), .dout(n26800));
    jdff dff_B_vGgx5UOl8_2(.din(n26800), .dout(n26803));
    jdff dff_B_0ss9W9jf0_2(.din(n26803), .dout(n26806));
    jdff dff_B_sQzvEDJH0_2(.din(n26806), .dout(n26809));
    jdff dff_B_Hj9Y9dzq5_2(.din(n26809), .dout(n26812));
    jdff dff_B_RE2q9mKr2_2(.din(n26812), .dout(n26815));
    jdff dff_B_cgkKqhsh2_2(.din(n26815), .dout(n26818));
    jdff dff_B_IllvyTv35_2(.din(n26818), .dout(n26821));
    jdff dff_B_OzYlfES70_2(.din(n26821), .dout(n26824));
    jdff dff_B_CupDJq5Y7_2(.din(n26824), .dout(n26827));
    jdff dff_B_V3vfjcVw0_2(.din(n26827), .dout(n26830));
    jdff dff_B_Cfb4vqSe7_2(.din(n26830), .dout(n26833));
    jdff dff_B_4C0WKNQH4_2(.din(n26833), .dout(n26836));
    jdff dff_B_i96nFEU98_2(.din(n26836), .dout(n26839));
    jdff dff_B_ypZ51DHP7_2(.din(n26839), .dout(n26842));
    jdff dff_B_zk0hrgOT6_2(.din(n26842), .dout(n26845));
    jdff dff_B_fmCt4rpQ0_2(.din(n26845), .dout(n26848));
    jdff dff_B_Us3zuZTo6_2(.din(n5865), .dout(n26851));
    jdff dff_B_8o2FsipG4_1(.din(n5857), .dout(n26854));
    jdff dff_B_yvHiPnQw7_2(.din(n5608), .dout(n26857));
    jdff dff_B_jUVPFEwC2_2(.din(n26857), .dout(n26860));
    jdff dff_B_GJuLF0m44_2(.din(n26860), .dout(n26863));
    jdff dff_B_b12wuBNb6_2(.din(n26863), .dout(n26866));
    jdff dff_B_qay5OBGx1_2(.din(n26866), .dout(n26869));
    jdff dff_B_lP0gwImO0_2(.din(n26869), .dout(n26872));
    jdff dff_B_k7XucLjP3_2(.din(n26872), .dout(n26875));
    jdff dff_B_NqDDxPS28_2(.din(n26875), .dout(n26878));
    jdff dff_B_0JQlx2xx9_2(.din(n26878), .dout(n26881));
    jdff dff_B_dDyXOI5Y6_2(.din(n26881), .dout(n26884));
    jdff dff_B_3T4EUipr5_2(.din(n26884), .dout(n26887));
    jdff dff_B_EmAbx1th6_2(.din(n26887), .dout(n26890));
    jdff dff_B_zDFDPh4S8_2(.din(n26890), .dout(n26893));
    jdff dff_B_MmorXoxh8_2(.din(n26893), .dout(n26896));
    jdff dff_B_7aMezkkc7_2(.din(n26896), .dout(n26899));
    jdff dff_B_PZUNlUiX7_2(.din(n26899), .dout(n26902));
    jdff dff_B_C1bhB9y15_2(.din(n26902), .dout(n26905));
    jdff dff_B_wL0SRZO77_2(.din(n26905), .dout(n26908));
    jdff dff_B_PQmflSPZ8_2(.din(n26908), .dout(n26911));
    jdff dff_B_2bVdqd6s8_2(.din(n26911), .dout(n26914));
    jdff dff_B_DQ6r8t1B7_2(.din(n26914), .dout(n26917));
    jdff dff_B_cIbBd5qZ7_2(.din(n26917), .dout(n26920));
    jdff dff_B_RacqNaBe5_2(.din(n26920), .dout(n26923));
    jdff dff_B_nD6vQqlA2_2(.din(n26923), .dout(n26926));
    jdff dff_B_uNVs8MvF4_2(.din(n26926), .dout(n26929));
    jdff dff_B_JQlG46sZ5_2(.din(n26929), .dout(n26932));
    jdff dff_B_VGko9RUY8_2(.din(n26932), .dout(n26935));
    jdff dff_B_HTldysDF6_2(.din(n26935), .dout(n26938));
    jdff dff_B_JzVxaj0z2_2(.din(n26938), .dout(n26941));
    jdff dff_B_NyAFTD8h7_2(.din(n26941), .dout(n26944));
    jdff dff_B_H3rhAmjQ4_2(.din(n26944), .dout(n26947));
    jdff dff_B_SUOXQVS70_2(.din(n26947), .dout(n26950));
    jdff dff_B_9UqHuJWk3_2(.din(n26950), .dout(n26953));
    jdff dff_B_5af9HRqt5_2(.din(n26953), .dout(n26956));
    jdff dff_B_68ngA5Vo5_2(.din(n26956), .dout(n26959));
    jdff dff_B_OMES7jqo9_2(.din(n5620), .dout(n26962));
    jdff dff_B_u5IVoq2a4_1(.din(n5612), .dout(n26965));
    jdff dff_B_YcFCBFPO3_2(.din(n5336), .dout(n26968));
    jdff dff_B_w4zDWyvm6_2(.din(n26968), .dout(n26971));
    jdff dff_B_2JWSzrzO0_2(.din(n26971), .dout(n26974));
    jdff dff_B_oTIs4USt9_2(.din(n26974), .dout(n26977));
    jdff dff_B_3zipsOJY5_2(.din(n26977), .dout(n26980));
    jdff dff_B_YIFSJtrs0_2(.din(n26980), .dout(n26983));
    jdff dff_B_N4acTxeA6_2(.din(n26983), .dout(n26986));
    jdff dff_B_eXEd1Tmq8_2(.din(n26986), .dout(n26989));
    jdff dff_B_21cSfqmk9_2(.din(n26989), .dout(n26992));
    jdff dff_B_OydAEvk49_2(.din(n26992), .dout(n26995));
    jdff dff_B_zLqu2rxX3_2(.din(n26995), .dout(n26998));
    jdff dff_B_zXzp0jIM8_2(.din(n26998), .dout(n27001));
    jdff dff_B_anhUD9a27_2(.din(n27001), .dout(n27004));
    jdff dff_B_eE1Wg2bl5_2(.din(n27004), .dout(n27007));
    jdff dff_B_MDKR1x8E2_2(.din(n27007), .dout(n27010));
    jdff dff_B_2O9MIAMb3_2(.din(n27010), .dout(n27013));
    jdff dff_B_iNFgzxZ08_2(.din(n27013), .dout(n27016));
    jdff dff_B_U8aDgk9d7_2(.din(n27016), .dout(n27019));
    jdff dff_B_ufLv9hl44_2(.din(n27019), .dout(n27022));
    jdff dff_B_8vwtoFUA6_2(.din(n27022), .dout(n27025));
    jdff dff_B_n7xiUSD47_2(.din(n27025), .dout(n27028));
    jdff dff_B_kciiJgb55_2(.din(n27028), .dout(n27031));
    jdff dff_B_zEkxCo4z3_2(.din(n27031), .dout(n27034));
    jdff dff_B_pgNjoc4F8_2(.din(n27034), .dout(n27037));
    jdff dff_B_u9kmetFt3_2(.din(n27037), .dout(n27040));
    jdff dff_B_ltVj1MsD6_2(.din(n27040), .dout(n27043));
    jdff dff_B_W2YPltbM3_2(.din(n27043), .dout(n27046));
    jdff dff_B_2oCdhB3n3_2(.din(n27046), .dout(n27049));
    jdff dff_B_ajPvAAUC4_2(.din(n27049), .dout(n27052));
    jdff dff_B_jYZV3R8I4_2(.din(n27052), .dout(n27055));
    jdff dff_B_jjedWkFG1_2(.din(n27055), .dout(n27058));
    jdff dff_B_njPQvG9e8_2(.din(n5348), .dout(n27061));
    jdff dff_B_DeIbx7lP9_1(.din(n5340), .dout(n27064));
    jdff dff_B_8e4NqzHw4_2(.din(n5037), .dout(n27067));
    jdff dff_B_9Vh8Bn5K4_2(.din(n27067), .dout(n27070));
    jdff dff_B_yRa6JZ6l7_2(.din(n27070), .dout(n27073));
    jdff dff_B_zdwx9JsP5_2(.din(n27073), .dout(n27076));
    jdff dff_B_3RknptOY1_2(.din(n27076), .dout(n27079));
    jdff dff_B_AOVLuSwa7_2(.din(n27079), .dout(n27082));
    jdff dff_B_wrNpn0Rv4_2(.din(n27082), .dout(n27085));
    jdff dff_B_SuxR5NWe6_2(.din(n27085), .dout(n27088));
    jdff dff_B_9Vxltf1N5_2(.din(n27088), .dout(n27091));
    jdff dff_B_oSCyB8iY8_2(.din(n27091), .dout(n27094));
    jdff dff_B_yrycadkq0_2(.din(n27094), .dout(n27097));
    jdff dff_B_vIIsJsSq8_2(.din(n27097), .dout(n27100));
    jdff dff_B_TgSk8gGZ1_2(.din(n27100), .dout(n27103));
    jdff dff_B_TFTtsks27_2(.din(n27103), .dout(n27106));
    jdff dff_B_RvZnRIGG5_2(.din(n27106), .dout(n27109));
    jdff dff_B_QD4U42DU1_2(.din(n27109), .dout(n27112));
    jdff dff_B_0sF7O7788_2(.din(n27112), .dout(n27115));
    jdff dff_B_VaE4exiy4_2(.din(n27115), .dout(n27118));
    jdff dff_B_xy9r5xCJ6_2(.din(n27118), .dout(n27121));
    jdff dff_B_rrP0XZrv6_2(.din(n27121), .dout(n27124));
    jdff dff_B_EjHAvBwx7_2(.din(n27124), .dout(n27127));
    jdff dff_B_dbN2Nquh8_2(.din(n27127), .dout(n27130));
    jdff dff_B_e34QdL9G8_2(.din(n27130), .dout(n27133));
    jdff dff_B_8cxraynF3_2(.din(n27133), .dout(n27136));
    jdff dff_B_QbmdQVPc6_2(.din(n27136), .dout(n27139));
    jdff dff_B_ouMsuwRl7_2(.din(n27139), .dout(n27142));
    jdff dff_B_kHJAgOSm2_2(.din(n27142), .dout(n27145));
    jdff dff_B_g4zIW2PC4_1(.din(n5041), .dout(n27148));
    jdff dff_B_AYwQZKXF4_2(.din(n4711), .dout(n27151));
    jdff dff_B_xaBHkDI30_2(.din(n27151), .dout(n27154));
    jdff dff_B_jeOGttWN8_2(.din(n27154), .dout(n27157));
    jdff dff_B_dHIOjesb1_2(.din(n27157), .dout(n27160));
    jdff dff_B_ygGQLR5W8_2(.din(n27160), .dout(n27163));
    jdff dff_B_WynmUHo74_2(.din(n27163), .dout(n27166));
    jdff dff_B_7KpYrw5Z4_2(.din(n27166), .dout(n27169));
    jdff dff_B_UVypv7lh7_2(.din(n27169), .dout(n27172));
    jdff dff_B_Ol5CSGFC4_2(.din(n27172), .dout(n27175));
    jdff dff_B_LUr1MXYX4_2(.din(n27175), .dout(n27178));
    jdff dff_B_URSG0eUG4_2(.din(n27178), .dout(n27181));
    jdff dff_B_7Jq3Nyio3_2(.din(n27181), .dout(n27184));
    jdff dff_B_k5Q1N5zD2_2(.din(n27184), .dout(n27187));
    jdff dff_B_OYPcVGBD1_2(.din(n27187), .dout(n27190));
    jdff dff_B_qXnGpUXg3_2(.din(n27190), .dout(n27193));
    jdff dff_B_IPPbY5Lz0_2(.din(n27193), .dout(n27196));
    jdff dff_B_1rwHte9Y5_2(.din(n27196), .dout(n27199));
    jdff dff_B_Np6mHN2u7_2(.din(n27199), .dout(n27202));
    jdff dff_B_jslJltsU6_2(.din(n27202), .dout(n27205));
    jdff dff_B_prf6axQ95_2(.din(n27205), .dout(n27208));
    jdff dff_B_AoafReTF8_2(.din(n27208), .dout(n27211));
    jdff dff_B_ikuXHfzF8_2(.din(n27211), .dout(n27214));
    jdff dff_B_5rfyVuhh2_2(.din(n27214), .dout(n27217));
    jdff dff_B_bpkdk6rt2_2(.din(n27217), .dout(n27220));
    jdff dff_B_JJRZtfhZ9_2(.din(n4808), .dout(n27223));
    jdff dff_B_uZ7dF0Vi0_1(.din(n4715), .dout(n27226));
    jdff dff_B_NOQlrnEz4_2(.din(n4365), .dout(n27229));
    jdff dff_B_ivEGhaFx0_2(.din(n27229), .dout(n27232));
    jdff dff_B_GRbcs1Zq0_2(.din(n27232), .dout(n27235));
    jdff dff_B_COEcUgMw3_2(.din(n27235), .dout(n27238));
    jdff dff_B_gJR63a2E9_2(.din(n27238), .dout(n27241));
    jdff dff_B_GG8SLyLe1_2(.din(n27241), .dout(n27244));
    jdff dff_B_q7RnC2cO8_2(.din(n27244), .dout(n27247));
    jdff dff_B_qG4cZdZk7_2(.din(n27247), .dout(n27250));
    jdff dff_B_9R7Dz9iL9_2(.din(n27250), .dout(n27253));
    jdff dff_B_vYsibJJa3_2(.din(n27253), .dout(n27256));
    jdff dff_B_eu0eYM0b0_2(.din(n27256), .dout(n27259));
    jdff dff_B_8myywXnU8_2(.din(n27259), .dout(n27262));
    jdff dff_B_mOsJWtyd9_2(.din(n27262), .dout(n27265));
    jdff dff_B_bH83fHp69_2(.din(n27265), .dout(n27268));
    jdff dff_B_Fzu3Vkti7_2(.din(n27268), .dout(n27271));
    jdff dff_B_zByCkGqu9_2(.din(n27271), .dout(n27274));
    jdff dff_B_Tcx4Y4gi5_2(.din(n27274), .dout(n27277));
    jdff dff_B_JkexPaGh0_2(.din(n27277), .dout(n27280));
    jdff dff_B_o4Lc9StX7_2(.din(n27280), .dout(n27283));
    jdff dff_B_n4cbJXyH0_2(.din(n27283), .dout(n27286));
    jdff dff_B_eXoYxCfj8_2(.din(n27286), .dout(n27289));
    jdff dff_B_cMtgVFzy1_2(.din(n4458), .dout(n27292));
    jdff dff_B_kK2ESgpI4_1(.din(n4369), .dout(n27295));
    jdff dff_B_mHn6A1TG5_2(.din(n3969), .dout(n27298));
    jdff dff_B_1vwQrPGr6_2(.din(n27298), .dout(n27301));
    jdff dff_B_qlumm9ey3_2(.din(n27301), .dout(n27304));
    jdff dff_B_buLk5kNv1_2(.din(n27304), .dout(n27307));
    jdff dff_B_brqUSC524_2(.din(n27307), .dout(n27310));
    jdff dff_B_hmKDX2123_2(.din(n27310), .dout(n27313));
    jdff dff_B_7a6b6YKa7_2(.din(n27313), .dout(n27316));
    jdff dff_B_KfiuQHT62_2(.din(n27316), .dout(n27319));
    jdff dff_B_UX5K9AA02_2(.din(n27319), .dout(n27322));
    jdff dff_B_5xw0O59C9_2(.din(n27322), .dout(n27325));
    jdff dff_B_XaBd5fvY9_2(.din(n27325), .dout(n27328));
    jdff dff_B_4Ajmh4Hz1_2(.din(n27328), .dout(n27331));
    jdff dff_B_GeeD8kzF0_2(.din(n27331), .dout(n27334));
    jdff dff_B_nEMqyReq9_2(.din(n27334), .dout(n27337));
    jdff dff_B_jiPdFc5v4_2(.din(n27337), .dout(n27340));
    jdff dff_B_7nqQFFA68_2(.din(n27340), .dout(n27343));
    jdff dff_B_KYByy9QX1_2(.din(n27343), .dout(n27346));
    jdff dff_B_9eFiQyfl7_2(.din(n27346), .dout(n27349));
    jdff dff_B_hZ2lehh50_2(.din(n4082), .dout(n27352));
    jdff dff_B_yk5YtVJ65_1(.din(n3973), .dout(n27355));
    jdff dff_B_iFI0Jw5b8_2(.din(n3592), .dout(n27358));
    jdff dff_B_Kv4pRacZ1_2(.din(n27358), .dout(n27361));
    jdff dff_B_bLaoZtQK9_2(.din(n27361), .dout(n27364));
    jdff dff_B_Tk3tCumm3_2(.din(n27364), .dout(n27367));
    jdff dff_B_RIbb9lo81_2(.din(n27367), .dout(n27370));
    jdff dff_B_fNkKkKfD6_2(.din(n27370), .dout(n27373));
    jdff dff_B_zRxHkNoV3_2(.din(n27373), .dout(n27376));
    jdff dff_B_FNNAJWGs8_2(.din(n27376), .dout(n27379));
    jdff dff_B_uVu1qw1Q7_2(.din(n27379), .dout(n27382));
    jdff dff_B_4lKUbKg04_2(.din(n27382), .dout(n27385));
    jdff dff_B_Tmmw64Qi2_2(.din(n27385), .dout(n27388));
    jdff dff_B_paeWwoNP1_2(.din(n27388), .dout(n27391));
    jdff dff_B_vV0WF0t53_2(.din(n27391), .dout(n27394));
    jdff dff_B_blbVkEUT9_2(.din(n27394), .dout(n27397));
    jdff dff_B_bflIGW7s7_2(.din(n27397), .dout(n27400));
    jdff dff_B_i5sM6kEZ8_2(.din(n3679), .dout(n27403));
    jdff dff_B_SB7dlvBc6_1(.din(n3596), .dout(n27406));
    jdff dff_B_Sklpz0k90_2(.din(n3191), .dout(n27409));
    jdff dff_B_W4v6kaYt6_2(.din(n27409), .dout(n27412));
    jdff dff_B_E09KK3E12_2(.din(n27412), .dout(n27415));
    jdff dff_B_lPn8Wxfn7_2(.din(n27415), .dout(n27418));
    jdff dff_B_jxOpEzbY9_2(.din(n27418), .dout(n27421));
    jdff dff_B_aE7bPIxk7_2(.din(n27421), .dout(n27424));
    jdff dff_B_kEUTOeIR7_2(.din(n27424), .dout(n27427));
    jdff dff_B_v4S3pv8l4_2(.din(n27427), .dout(n27430));
    jdff dff_B_EhWVhiBI6_2(.din(n27430), .dout(n27433));
    jdff dff_B_LIaiFfNQ6_2(.din(n27433), .dout(n27436));
    jdff dff_B_uKetQiRC1_2(.din(n27436), .dout(n27439));
    jdff dff_B_yAr04H9W1_2(.din(n27439), .dout(n27442));
    jdff dff_B_QPpQGM361_2(.din(n3277), .dout(n27445));
    jdff dff_B_UNbWXrTi5_1(.din(n3195), .dout(n27448));
    jdff dff_B_C5q94eMr1_2(.din(n2812), .dout(n27451));
    jdff dff_B_irBegRFQ8_2(.din(n27451), .dout(n27454));
    jdff dff_B_qwRekFJZ8_2(.din(n27454), .dout(n27457));
    jdff dff_B_eb8W9Ta22_2(.din(n27457), .dout(n27460));
    jdff dff_B_l2EDcrU55_2(.din(n27460), .dout(n27463));
    jdff dff_B_85hhOQCy4_2(.din(n27463), .dout(n27466));
    jdff dff_B_qsBeduna3_2(.din(n27466), .dout(n27469));
    jdff dff_B_XGOvkdA66_2(.din(n27469), .dout(n27472));
    jdff dff_B_4LFn6EgN7_2(.din(n27472), .dout(n27475));
    jdff dff_B_6JFRe99A8_2(.din(n2872), .dout(n27478));
    jdff dff_B_nzwKRckY6_2(.din(n27478), .dout(n27481));
    jdff dff_B_F6KKqp0I8_1(.din(n2815), .dout(n27484));
    jdff dff_B_208H61nz4_1(.din(n27484), .dout(n27487));
    jdff dff_B_nfh0Anse2_1(.din(n27487), .dout(n27490));
    jdff dff_B_aGehSRJq9_1(.din(n27490), .dout(n27493));
    jdff dff_B_pK6cNqnY1_1(.din(n27493), .dout(n27496));
    jdff dff_B_ycQziHRj5_1(.din(n27496), .dout(n27499));
    jdff dff_B_ghKvLSbr0_0(.din(n2490), .dout(n27502));
    jdff dff_B_PYhFfXDa8_0(.din(n27502), .dout(n27505));
    jdff dff_A_Iuo8bC7C8_0(.din(n27510), .dout(n27507));
    jdff dff_A_UmkstwiT2_0(.din(n27513), .dout(n27510));
    jdff dff_A_LRlOYx2p2_0(.din(n2486), .dout(n27513));
    jdff dff_B_j6eUikvB2_1(.din(n2464), .dout(n27517));
    jdff dff_A_Ai6ny8Yz9_0(.din(n2125), .dout(n27519));
    jdff dff_A_sWnJlBNP2_1(.din(n27525), .dout(n27522));
    jdff dff_A_MUWNUiji3_1(.din(n2125), .dout(n27525));
    jdff dff_A_DKGW4iE87_1(.din(n27531), .dout(n27528));
    jdff dff_A_ZtDRweVm1_1(.din(n27534), .dout(n27531));
    jdff dff_A_3Pzw6UTd0_1(.din(n27537), .dout(n27534));
    jdff dff_A_1d6TTFCT0_1(.din(n27540), .dout(n27537));
    jdff dff_A_Ophfcl6M1_1(.din(n27543), .dout(n27540));
    jdff dff_A_bBP3iweD3_1(.din(n2456), .dout(n27543));
    jdff dff_B_NiRQ0XUX0_1(.din(n6764), .dout(n27547));
    jdff dff_A_yvPCCEoS2_1(.din(n6695), .dout(n27549));
    jdff dff_B_CTe4bPiS3_1(.din(n6687), .dout(n27553));
    jdff dff_B_4nIVDGd25_2(.din(n6576), .dout(n27556));
    jdff dff_B_QUfPRJAv6_2(.din(n27556), .dout(n27559));
    jdff dff_B_quiluQjn1_2(.din(n27559), .dout(n27562));
    jdff dff_B_Lwpwq0Rs1_2(.din(n27562), .dout(n27565));
    jdff dff_B_go08VVGf3_2(.din(n27565), .dout(n27568));
    jdff dff_B_r02VsDN50_2(.din(n27568), .dout(n27571));
    jdff dff_B_AD3YtUdT3_2(.din(n27571), .dout(n27574));
    jdff dff_B_YidBgOfN1_2(.din(n27574), .dout(n27577));
    jdff dff_B_Eh6HP9FU7_2(.din(n27577), .dout(n27580));
    jdff dff_B_aCqiNgN90_2(.din(n27580), .dout(n27583));
    jdff dff_B_O7uZei4a2_2(.din(n27583), .dout(n27586));
    jdff dff_B_KlPistLC0_2(.din(n27586), .dout(n27589));
    jdff dff_B_5Uci0xnl4_2(.din(n27589), .dout(n27592));
    jdff dff_B_tsTNUwdT8_2(.din(n27592), .dout(n27595));
    jdff dff_B_IhEt0xlD8_2(.din(n27595), .dout(n27598));
    jdff dff_B_R5eYr6q44_2(.din(n27598), .dout(n27601));
    jdff dff_B_HF8XaDwQ5_2(.din(n27601), .dout(n27604));
    jdff dff_B_eCZCoMfL5_2(.din(n27604), .dout(n27607));
    jdff dff_B_65c9tFPw6_2(.din(n27607), .dout(n27610));
    jdff dff_B_c7nY5kDD2_2(.din(n27610), .dout(n27613));
    jdff dff_B_aUv76SM82_2(.din(n27613), .dout(n27616));
    jdff dff_B_NjvE3s542_2(.din(n27616), .dout(n27619));
    jdff dff_B_BeEC1Zg71_2(.din(n27619), .dout(n27622));
    jdff dff_B_8o94F5ir9_2(.din(n27622), .dout(n27625));
    jdff dff_B_6jffrsIL3_2(.din(n27625), .dout(n27628));
    jdff dff_B_obcOtCP87_2(.din(n27628), .dout(n27631));
    jdff dff_B_hwvu0FLI9_2(.din(n27631), .dout(n27634));
    jdff dff_B_pbZRBvRS6_2(.din(n27634), .dout(n27637));
    jdff dff_B_SPRwxoXi1_2(.din(n27637), .dout(n27640));
    jdff dff_B_W5tD9vhU1_2(.din(n27640), .dout(n27643));
    jdff dff_B_gKsJZiiL0_2(.din(n27643), .dout(n27646));
    jdff dff_B_kiKmBUMo3_2(.din(n27646), .dout(n27649));
    jdff dff_B_tROCr7Qy1_2(.din(n27649), .dout(n27652));
    jdff dff_B_9DKHQsVB6_2(.din(n27652), .dout(n27655));
    jdff dff_B_lvIOlS5B8_2(.din(n27655), .dout(n27658));
    jdff dff_B_aULnmtzK4_2(.din(n27658), .dout(n27661));
    jdff dff_B_gICv0iZF9_2(.din(n27661), .dout(n27664));
    jdff dff_B_qNV9so0P2_2(.din(n27664), .dout(n27667));
    jdff dff_B_ymtchohA0_2(.din(n27667), .dout(n27670));
    jdff dff_B_hzjYATWG7_2(.din(n27670), .dout(n27673));
    jdff dff_B_mX3K5PLX2_2(.din(n27673), .dout(n27676));
    jdff dff_B_CxOv5dCV8_2(.din(n27676), .dout(n27679));
    jdff dff_B_N9peuzqX8_2(.din(n27679), .dout(n27682));
    jdff dff_B_ia8C6Jxo2_2(.din(n27682), .dout(n27685));
    jdff dff_B_4h1mvUyI5_2(.din(n27685), .dout(n27688));
    jdff dff_B_dFVoXNyH6_2(.din(n27688), .dout(n27691));
    jdff dff_B_R2Uyxj707_2(.din(n27691), .dout(n27694));
    jdff dff_B_t6OTknWa2_2(.din(n27694), .dout(n27697));
    jdff dff_B_KJSXHFsq9_2(.din(n27697), .dout(n27700));
    jdff dff_B_ZaTVUDFY8_2(.din(n27700), .dout(n27703));
    jdff dff_B_NrKguckG2_2(.din(n27703), .dout(n27706));
    jdff dff_B_slftNcig9_2(.din(n27706), .dout(n27709));
    jdff dff_B_Yzc9RcZh4_2(.din(n27709), .dout(n27712));
    jdff dff_B_2XG2nvNA2_2(.din(n6588), .dout(n27715));
    jdff dff_B_b90Z7vXn8_1(.din(n6580), .dout(n27718));
    jdff dff_B_KXCtdLDY9_2(.din(n6442), .dout(n27721));
    jdff dff_B_ZPMbSx675_2(.din(n27721), .dout(n27724));
    jdff dff_B_oabqylBl9_2(.din(n27724), .dout(n27727));
    jdff dff_B_A0AcWmW61_2(.din(n27727), .dout(n27730));
    jdff dff_B_3pAKkzOx4_2(.din(n27730), .dout(n27733));
    jdff dff_B_qUoeQIKv6_2(.din(n27733), .dout(n27736));
    jdff dff_B_s4PK1PJk0_2(.din(n27736), .dout(n27739));
    jdff dff_B_5qVeG1Dk9_2(.din(n27739), .dout(n27742));
    jdff dff_B_ZdHKM6qD3_2(.din(n27742), .dout(n27745));
    jdff dff_B_i9an8hkh6_2(.din(n27745), .dout(n27748));
    jdff dff_B_5sjCzV3N6_2(.din(n27748), .dout(n27751));
    jdff dff_B_gPof9vDJ0_2(.din(n27751), .dout(n27754));
    jdff dff_B_Aq0lgHlt0_2(.din(n27754), .dout(n27757));
    jdff dff_B_Tres6fIH3_2(.din(n27757), .dout(n27760));
    jdff dff_B_b7EvgEKd2_2(.din(n27760), .dout(n27763));
    jdff dff_B_9vI8bOzX1_2(.din(n27763), .dout(n27766));
    jdff dff_B_2RDqrGKY7_2(.din(n27766), .dout(n27769));
    jdff dff_B_5TwqCLW80_2(.din(n27769), .dout(n27772));
    jdff dff_B_woQAuOM94_2(.din(n27772), .dout(n27775));
    jdff dff_B_f2G8Qthw2_2(.din(n27775), .dout(n27778));
    jdff dff_B_PG6hOt2x3_2(.din(n27778), .dout(n27781));
    jdff dff_B_m0ipGKvO8_2(.din(n27781), .dout(n27784));
    jdff dff_B_lUtFYRnr3_2(.din(n27784), .dout(n27787));
    jdff dff_B_KebbMlSm5_2(.din(n27787), .dout(n27790));
    jdff dff_B_oNxnqqyu5_2(.din(n27790), .dout(n27793));
    jdff dff_B_1l8dkLAa2_2(.din(n27793), .dout(n27796));
    jdff dff_B_nCz172J18_2(.din(n27796), .dout(n27799));
    jdff dff_B_AxL68lvD9_2(.din(n27799), .dout(n27802));
    jdff dff_B_f5mxh1ET3_2(.din(n27802), .dout(n27805));
    jdff dff_B_o20zr0du2_2(.din(n27805), .dout(n27808));
    jdff dff_B_ZeIq7Lxt3_2(.din(n27808), .dout(n27811));
    jdff dff_B_3OKcia3V4_2(.din(n27811), .dout(n27814));
    jdff dff_B_x1Y6veYi8_2(.din(n27814), .dout(n27817));
    jdff dff_B_mrBya4Ue2_2(.din(n27817), .dout(n27820));
    jdff dff_B_1rR9e1Ob7_2(.din(n27820), .dout(n27823));
    jdff dff_B_VgSSCo7L6_2(.din(n27823), .dout(n27826));
    jdff dff_B_4Inb6VYI6_2(.din(n27826), .dout(n27829));
    jdff dff_B_iFlcSjGb2_2(.din(n27829), .dout(n27832));
    jdff dff_B_Uc3LKQd95_2(.din(n27832), .dout(n27835));
    jdff dff_B_7uSCX6Ej2_2(.din(n27835), .dout(n27838));
    jdff dff_B_VTXlkmTV2_2(.din(n27838), .dout(n27841));
    jdff dff_B_ta4tm3Ee2_2(.din(n27841), .dout(n27844));
    jdff dff_B_ETpWHW4o5_2(.din(n27844), .dout(n27847));
    jdff dff_B_2PiFW1EC3_2(.din(n27847), .dout(n27850));
    jdff dff_B_hXelHWkr4_2(.din(n27850), .dout(n27853));
    jdff dff_B_1YHFoZHD0_2(.din(n27853), .dout(n27856));
    jdff dff_B_xCbISSsD1_2(.din(n27856), .dout(n27859));
    jdff dff_B_MIp6UnZx6_2(.din(n27859), .dout(n27862));
    jdff dff_B_09FlSBNU8_2(.din(n27862), .dout(n27865));
    jdff dff_B_Hto6pA017_2(.din(n6454), .dout(n27868));
    jdff dff_B_GBFhlqJt1_1(.din(n6446), .dout(n27871));
    jdff dff_B_4UDLIoq55_2(.din(n6284), .dout(n27874));
    jdff dff_B_6W6ZzYxM6_2(.din(n27874), .dout(n27877));
    jdff dff_B_XH1xguaG7_2(.din(n27877), .dout(n27880));
    jdff dff_B_wEzATMU09_2(.din(n27880), .dout(n27883));
    jdff dff_B_nndZOcyO3_2(.din(n27883), .dout(n27886));
    jdff dff_B_DFfnGP5J9_2(.din(n27886), .dout(n27889));
    jdff dff_B_BLdlEHzf0_2(.din(n27889), .dout(n27892));
    jdff dff_B_mh1EG16L9_2(.din(n27892), .dout(n27895));
    jdff dff_B_k5sQI2H94_2(.din(n27895), .dout(n27898));
    jdff dff_B_gIS3kEDz2_2(.din(n27898), .dout(n27901));
    jdff dff_B_WuTXHVMW8_2(.din(n27901), .dout(n27904));
    jdff dff_B_tVhIJKlQ7_2(.din(n27904), .dout(n27907));
    jdff dff_B_cWNrJTbM5_2(.din(n27907), .dout(n27910));
    jdff dff_B_kbAsr9uR3_2(.din(n27910), .dout(n27913));
    jdff dff_B_NipPy7uN2_2(.din(n27913), .dout(n27916));
    jdff dff_B_eiXdaOvx5_2(.din(n27916), .dout(n27919));
    jdff dff_B_vLi2tK112_2(.din(n27919), .dout(n27922));
    jdff dff_B_ksl1FEt55_2(.din(n27922), .dout(n27925));
    jdff dff_B_9juIz4GK3_2(.din(n27925), .dout(n27928));
    jdff dff_B_87lSFLpn4_2(.din(n27928), .dout(n27931));
    jdff dff_B_uX0s9TIR7_2(.din(n27931), .dout(n27934));
    jdff dff_B_K6W7jNUc1_2(.din(n27934), .dout(n27937));
    jdff dff_B_xBMYqHLV8_2(.din(n27937), .dout(n27940));
    jdff dff_B_D1VcgLeh7_2(.din(n27940), .dout(n27943));
    jdff dff_B_Kc3U1Dgf5_2(.din(n27943), .dout(n27946));
    jdff dff_B_fS7xFAsa4_2(.din(n27946), .dout(n27949));
    jdff dff_B_hJgONq219_2(.din(n27949), .dout(n27952));
    jdff dff_B_7HZ5Uspp5_2(.din(n27952), .dout(n27955));
    jdff dff_B_lRMMQxUd3_2(.din(n27955), .dout(n27958));
    jdff dff_B_NUYPluOB9_2(.din(n27958), .dout(n27961));
    jdff dff_B_M4hO2AI63_2(.din(n27961), .dout(n27964));
    jdff dff_B_E38pZlid0_2(.din(n27964), .dout(n27967));
    jdff dff_B_v3RGeEgj5_2(.din(n27967), .dout(n27970));
    jdff dff_B_0IskqFG09_2(.din(n27970), .dout(n27973));
    jdff dff_B_s5JImO5R6_2(.din(n27973), .dout(n27976));
    jdff dff_B_IFDitTZ19_2(.din(n27976), .dout(n27979));
    jdff dff_B_zqvwS3iM5_2(.din(n27979), .dout(n27982));
    jdff dff_B_i1aIOw928_2(.din(n27982), .dout(n27985));
    jdff dff_B_Gdc5TsG35_2(.din(n27985), .dout(n27988));
    jdff dff_B_CqHiyiZY7_2(.din(n27988), .dout(n27991));
    jdff dff_B_LfEiPaCA7_2(.din(n27991), .dout(n27994));
    jdff dff_B_Gpze2ohh9_2(.din(n27994), .dout(n27997));
    jdff dff_B_4OrxLSvx8_2(.din(n27997), .dout(n28000));
    jdff dff_B_lb9kz3zq0_2(.din(n28000), .dout(n28003));
    jdff dff_B_icbpygs14_2(.din(n28003), .dout(n28006));
    jdff dff_B_CWjW9Ljq8_2(.din(n6296), .dout(n28009));
    jdff dff_B_IVGV1hWr7_1(.din(n6288), .dout(n28012));
    jdff dff_B_273ZWcL18_2(.din(n6090), .dout(n28015));
    jdff dff_B_gLWEgUOH6_2(.din(n28015), .dout(n28018));
    jdff dff_B_oco2Xphf9_2(.din(n28018), .dout(n28021));
    jdff dff_B_xZiyinH49_2(.din(n28021), .dout(n28024));
    jdff dff_B_QtSkH6op7_2(.din(n28024), .dout(n28027));
    jdff dff_B_n6Yh4seq7_2(.din(n28027), .dout(n28030));
    jdff dff_B_7MxdhzbH0_2(.din(n28030), .dout(n28033));
    jdff dff_B_g5a79xU07_2(.din(n28033), .dout(n28036));
    jdff dff_B_W0GnBM7v9_2(.din(n28036), .dout(n28039));
    jdff dff_B_ApJ9mZ5m1_2(.din(n28039), .dout(n28042));
    jdff dff_B_BeobT1ZP5_2(.din(n28042), .dout(n28045));
    jdff dff_B_vW33an8Q9_2(.din(n28045), .dout(n28048));
    jdff dff_B_QOIXrkTW8_2(.din(n28048), .dout(n28051));
    jdff dff_B_NtK0a0m25_2(.din(n28051), .dout(n28054));
    jdff dff_B_VCgPFZcq9_2(.din(n28054), .dout(n28057));
    jdff dff_B_g26D1fnS9_2(.din(n28057), .dout(n28060));
    jdff dff_B_cUQTFXfz3_2(.din(n28060), .dout(n28063));
    jdff dff_B_fc7bjt8A9_2(.din(n28063), .dout(n28066));
    jdff dff_B_QTttfCQz4_2(.din(n28066), .dout(n28069));
    jdff dff_B_dN2AR35P0_2(.din(n28069), .dout(n28072));
    jdff dff_B_TOHUYWdZ1_2(.din(n28072), .dout(n28075));
    jdff dff_B_q6qrVm9B0_2(.din(n28075), .dout(n28078));
    jdff dff_B_OihMuvS32_2(.din(n28078), .dout(n28081));
    jdff dff_B_ndJRK4Ir6_2(.din(n28081), .dout(n28084));
    jdff dff_B_if7qqmyu3_2(.din(n28084), .dout(n28087));
    jdff dff_B_pksl8QHj3_2(.din(n28087), .dout(n28090));
    jdff dff_B_i6IMqcDR0_2(.din(n28090), .dout(n28093));
    jdff dff_B_k2vqLwNI5_2(.din(n28093), .dout(n28096));
    jdff dff_B_JnDYOcxb6_2(.din(n28096), .dout(n28099));
    jdff dff_B_u2SVdbn26_2(.din(n28099), .dout(n28102));
    jdff dff_B_uyYZNR952_2(.din(n28102), .dout(n28105));
    jdff dff_B_CaS43xin0_2(.din(n28105), .dout(n28108));
    jdff dff_B_iTqTfpYg1_2(.din(n28108), .dout(n28111));
    jdff dff_B_JzbMjfsx6_2(.din(n28111), .dout(n28114));
    jdff dff_B_Qe7aWXeH0_2(.din(n28114), .dout(n28117));
    jdff dff_B_045T1oLg8_2(.din(n28117), .dout(n28120));
    jdff dff_B_URcjHMWH7_2(.din(n28120), .dout(n28123));
    jdff dff_B_hyrv6va34_2(.din(n28123), .dout(n28126));
    jdff dff_B_dnZ792338_2(.din(n28126), .dout(n28129));
    jdff dff_B_mFUXl2Vr0_2(.din(n28129), .dout(n28132));
    jdff dff_B_49g8mCix4_2(.din(n28132), .dout(n28135));
    jdff dff_B_D0oz23es3_2(.din(n6102), .dout(n28138));
    jdff dff_B_BceJ9HAg2_1(.din(n6094), .dout(n28141));
    jdff dff_B_XU1ib5pi4_2(.din(n5872), .dout(n28144));
    jdff dff_B_4Hf9CiEg8_2(.din(n28144), .dout(n28147));
    jdff dff_B_PQbTCk5t0_2(.din(n28147), .dout(n28150));
    jdff dff_B_JwZJKHav3_2(.din(n28150), .dout(n28153));
    jdff dff_B_IU07JJ6l8_2(.din(n28153), .dout(n28156));
    jdff dff_B_iQyohNPb5_2(.din(n28156), .dout(n28159));
    jdff dff_B_2syLQrTk8_2(.din(n28159), .dout(n28162));
    jdff dff_B_c6BjeoqK3_2(.din(n28162), .dout(n28165));
    jdff dff_B_5CWHnyk14_2(.din(n28165), .dout(n28168));
    jdff dff_B_1ev366XH7_2(.din(n28168), .dout(n28171));
    jdff dff_B_kAPCeusT6_2(.din(n28171), .dout(n28174));
    jdff dff_B_Ui9tzaJe3_2(.din(n28174), .dout(n28177));
    jdff dff_B_8hseRavn4_2(.din(n28177), .dout(n28180));
    jdff dff_B_1hIBzhWY4_2(.din(n28180), .dout(n28183));
    jdff dff_B_yPUbsZcR6_2(.din(n28183), .dout(n28186));
    jdff dff_B_0Yx81Hka1_2(.din(n28186), .dout(n28189));
    jdff dff_B_0iY5WYrK6_2(.din(n28189), .dout(n28192));
    jdff dff_B_vIluE7Hi3_2(.din(n28192), .dout(n28195));
    jdff dff_B_jO7epaEW3_2(.din(n28195), .dout(n28198));
    jdff dff_B_Qwxy4cgT8_2(.din(n28198), .dout(n28201));
    jdff dff_B_6P7mbnmE0_2(.din(n28201), .dout(n28204));
    jdff dff_B_T9lmb8lD4_2(.din(n28204), .dout(n28207));
    jdff dff_B_uBmoyWnJ8_2(.din(n28207), .dout(n28210));
    jdff dff_B_aXfjF8iJ7_2(.din(n28210), .dout(n28213));
    jdff dff_B_L5RnNB3u8_2(.din(n28213), .dout(n28216));
    jdff dff_B_F3I74PE33_2(.din(n28216), .dout(n28219));
    jdff dff_B_OSC9w5fH6_2(.din(n28219), .dout(n28222));
    jdff dff_B_7aV4A1kK0_2(.din(n28222), .dout(n28225));
    jdff dff_B_Vqb8uKpm7_2(.din(n28225), .dout(n28228));
    jdff dff_B_VZEGaTD22_2(.din(n28228), .dout(n28231));
    jdff dff_B_e2dWQ5mI9_2(.din(n28231), .dout(n28234));
    jdff dff_B_eWJ0iAyU8_2(.din(n28234), .dout(n28237));
    jdff dff_B_yTiDZGKA7_2(.din(n28237), .dout(n28240));
    jdff dff_B_BB7c8lP05_2(.din(n28240), .dout(n28243));
    jdff dff_B_9VhKkMOn9_2(.din(n28243), .dout(n28246));
    jdff dff_B_gBhgOVnT1_2(.din(n28246), .dout(n28249));
    jdff dff_B_89y1K2Xs8_2(.din(n28249), .dout(n28252));
    jdff dff_B_mk4QHZQS7_2(.din(n5884), .dout(n28255));
    jdff dff_B_SAOoRhsC9_1(.din(n5876), .dout(n28258));
    jdff dff_B_XjefX4721_2(.din(n5627), .dout(n28261));
    jdff dff_B_NolhAyI60_2(.din(n28261), .dout(n28264));
    jdff dff_B_5Ux9wGwm5_2(.din(n28264), .dout(n28267));
    jdff dff_B_LD6nPV3L0_2(.din(n28267), .dout(n28270));
    jdff dff_B_qi2cPUYf2_2(.din(n28270), .dout(n28273));
    jdff dff_B_EnY0yLLv9_2(.din(n28273), .dout(n28276));
    jdff dff_B_aKQqJcDg9_2(.din(n28276), .dout(n28279));
    jdff dff_B_ZClTf7qy1_2(.din(n28279), .dout(n28282));
    jdff dff_B_IpAfcqwl0_2(.din(n28282), .dout(n28285));
    jdff dff_B_mrKCDw2q9_2(.din(n28285), .dout(n28288));
    jdff dff_B_U08s84Q54_2(.din(n28288), .dout(n28291));
    jdff dff_B_YVAuNIrv0_2(.din(n28291), .dout(n28294));
    jdff dff_B_0LxnTeCw2_2(.din(n28294), .dout(n28297));
    jdff dff_B_9xHkYdKc0_2(.din(n28297), .dout(n28300));
    jdff dff_B_l4Mnnc7U8_2(.din(n28300), .dout(n28303));
    jdff dff_B_W0QLLP3E9_2(.din(n28303), .dout(n28306));
    jdff dff_B_kJ4UVvww1_2(.din(n28306), .dout(n28309));
    jdff dff_B_iYxINs7f7_2(.din(n28309), .dout(n28312));
    jdff dff_B_IS2dR1B27_2(.din(n28312), .dout(n28315));
    jdff dff_B_7k2RvW6g1_2(.din(n28315), .dout(n28318));
    jdff dff_B_v75OYDqx0_2(.din(n28318), .dout(n28321));
    jdff dff_B_f3JmymHX2_2(.din(n28321), .dout(n28324));
    jdff dff_B_xnqkOxxm0_2(.din(n28324), .dout(n28327));
    jdff dff_B_s6uW2cIn2_2(.din(n28327), .dout(n28330));
    jdff dff_B_XRBAfsxD8_2(.din(n28330), .dout(n28333));
    jdff dff_B_YwwbrA3T6_2(.din(n28333), .dout(n28336));
    jdff dff_B_ndj0dHNJ8_2(.din(n28336), .dout(n28339));
    jdff dff_B_6bjCgydK2_2(.din(n28339), .dout(n28342));
    jdff dff_B_vpcUPsY24_2(.din(n28342), .dout(n28345));
    jdff dff_B_3eIUFEBL4_2(.din(n28345), .dout(n28348));
    jdff dff_B_yz6ItiD02_2(.din(n28348), .dout(n28351));
    jdff dff_B_OYI5TTQ27_2(.din(n28351), .dout(n28354));
    jdff dff_B_sEVUrz8g0_2(.din(n28354), .dout(n28357));
    jdff dff_B_4P5mUltv6_2(.din(n5639), .dout(n28360));
    jdff dff_B_TCdl79rD8_1(.din(n5631), .dout(n28363));
    jdff dff_B_edWN1NhW4_2(.din(n5355), .dout(n28366));
    jdff dff_B_HHx47qXL1_2(.din(n28366), .dout(n28369));
    jdff dff_B_rc7qgt0a3_2(.din(n28369), .dout(n28372));
    jdff dff_B_dIWe51b91_2(.din(n28372), .dout(n28375));
    jdff dff_B_HHe1uSsr2_2(.din(n28375), .dout(n28378));
    jdff dff_B_UUMlViDm1_2(.din(n28378), .dout(n28381));
    jdff dff_B_FACeCpGh4_2(.din(n28381), .dout(n28384));
    jdff dff_B_FRwGckXt5_2(.din(n28384), .dout(n28387));
    jdff dff_B_1DapE0cs9_2(.din(n28387), .dout(n28390));
    jdff dff_B_JVZC70tZ0_2(.din(n28390), .dout(n28393));
    jdff dff_B_ljxaKdkG0_2(.din(n28393), .dout(n28396));
    jdff dff_B_VOthYxX98_2(.din(n28396), .dout(n28399));
    jdff dff_B_fdfOxRjd5_2(.din(n28399), .dout(n28402));
    jdff dff_B_XKiqIZ5r4_2(.din(n28402), .dout(n28405));
    jdff dff_B_NeSmKgSE2_2(.din(n28405), .dout(n28408));
    jdff dff_B_F3SclU8R3_2(.din(n28408), .dout(n28411));
    jdff dff_B_XSyHIbcY0_2(.din(n28411), .dout(n28414));
    jdff dff_B_4LHxSwYK3_2(.din(n28414), .dout(n28417));
    jdff dff_B_P187kyDT4_2(.din(n28417), .dout(n28420));
    jdff dff_B_v0lmHB5I7_2(.din(n28420), .dout(n28423));
    jdff dff_B_wVKtpP5L9_2(.din(n28423), .dout(n28426));
    jdff dff_B_vYdEo0Fz2_2(.din(n28426), .dout(n28429));
    jdff dff_B_hz8Uspyn5_2(.din(n28429), .dout(n28432));
    jdff dff_B_zRU4CEaB0_2(.din(n28432), .dout(n28435));
    jdff dff_B_5zbn9sFc5_2(.din(n28435), .dout(n28438));
    jdff dff_B_7ubZMhHE7_2(.din(n28438), .dout(n28441));
    jdff dff_B_7EEoPkXK2_2(.din(n28441), .dout(n28444));
    jdff dff_B_VsStI1L86_2(.din(n28444), .dout(n28447));
    jdff dff_B_hT9Ev7Vt9_2(.din(n28447), .dout(n28450));
    jdff dff_B_qdYNCKvA2_2(.din(n5367), .dout(n28453));
    jdff dff_B_QsPz98oR1_1(.din(n5359), .dout(n28456));
    jdff dff_B_GrRxEaNu6_2(.din(n5056), .dout(n28459));
    jdff dff_B_rEGRSoG71_2(.din(n28459), .dout(n28462));
    jdff dff_B_tGa8r5Lc4_2(.din(n28462), .dout(n28465));
    jdff dff_B_ejkEqu0H3_2(.din(n28465), .dout(n28468));
    jdff dff_B_2NN5B2kf0_2(.din(n28468), .dout(n28471));
    jdff dff_B_RHDjHqwB8_2(.din(n28471), .dout(n28474));
    jdff dff_B_QEiEL3mN7_2(.din(n28474), .dout(n28477));
    jdff dff_B_JJKIdqw52_2(.din(n28477), .dout(n28480));
    jdff dff_B_OUNeJMVY8_2(.din(n28480), .dout(n28483));
    jdff dff_B_xkoXLOF85_2(.din(n28483), .dout(n28486));
    jdff dff_B_Jed5Tjm11_2(.din(n28486), .dout(n28489));
    jdff dff_B_mp4F1oZH8_2(.din(n28489), .dout(n28492));
    jdff dff_B_eEJfo6TG8_2(.din(n28492), .dout(n28495));
    jdff dff_B_RO0EvG131_2(.din(n28495), .dout(n28498));
    jdff dff_B_0hbscURz9_2(.din(n28498), .dout(n28501));
    jdff dff_B_uErcEyIz3_2(.din(n28501), .dout(n28504));
    jdff dff_B_8wOoISR05_2(.din(n28504), .dout(n28507));
    jdff dff_B_fKU9188e7_2(.din(n28507), .dout(n28510));
    jdff dff_B_ZbKGSvYT9_2(.din(n28510), .dout(n28513));
    jdff dff_B_MqbE7NgF3_2(.din(n28513), .dout(n28516));
    jdff dff_B_OoAHvFgV5_2(.din(n28516), .dout(n28519));
    jdff dff_B_qf2DMypr4_2(.din(n28519), .dout(n28522));
    jdff dff_B_pMKCDJvG9_2(.din(n28522), .dout(n28525));
    jdff dff_B_VrZdiStE9_2(.din(n28525), .dout(n28528));
    jdff dff_B_7bdxXkSP7_2(.din(n28528), .dout(n28531));
    jdff dff_B_c1BRs3pm3_2(.din(n5068), .dout(n28534));
    jdff dff_B_f3NceXEh7_1(.din(n5060), .dout(n28537));
    jdff dff_B_lCx35bWy3_2(.din(n4730), .dout(n28540));
    jdff dff_B_AztIEZv59_2(.din(n28540), .dout(n28543));
    jdff dff_B_d7TUXjew0_2(.din(n28543), .dout(n28546));
    jdff dff_B_k9Jg1eEh3_2(.din(n28546), .dout(n28549));
    jdff dff_B_124TKauY1_2(.din(n28549), .dout(n28552));
    jdff dff_B_mOF0fu9Y5_2(.din(n28552), .dout(n28555));
    jdff dff_B_Kl3R1ejy5_2(.din(n28555), .dout(n28558));
    jdff dff_B_qfbSuO2U5_2(.din(n28558), .dout(n28561));
    jdff dff_B_iPLNtMfH4_2(.din(n28561), .dout(n28564));
    jdff dff_B_LFvrOSLM2_2(.din(n28564), .dout(n28567));
    jdff dff_B_y5xnIrsl7_2(.din(n28567), .dout(n28570));
    jdff dff_B_KiJengFT6_2(.din(n28570), .dout(n28573));
    jdff dff_B_Ha11kADe9_2(.din(n28573), .dout(n28576));
    jdff dff_B_UrtMm4fC2_2(.din(n28576), .dout(n28579));
    jdff dff_B_n98Zh5Uc4_2(.din(n28579), .dout(n28582));
    jdff dff_B_6BtnarNa7_2(.din(n28582), .dout(n28585));
    jdff dff_B_WIL0cb5J4_2(.din(n28585), .dout(n28588));
    jdff dff_B_NqJgbb3l5_2(.din(n28588), .dout(n28591));
    jdff dff_B_bPKMX1LZ2_2(.din(n28591), .dout(n28594));
    jdff dff_B_gOxNeTZb8_2(.din(n28594), .dout(n28597));
    jdff dff_B_3XfacPBE0_2(.din(n28597), .dout(n28600));
    jdff dff_B_Za8DoiXy7_1(.din(n4734), .dout(n28603));
    jdff dff_B_r5fzfAxf9_2(.din(n4384), .dout(n28606));
    jdff dff_B_ePE49Jzy5_2(.din(n28606), .dout(n28609));
    jdff dff_B_Ve2RcBtt0_2(.din(n28609), .dout(n28612));
    jdff dff_B_Mz06rtE93_2(.din(n28612), .dout(n28615));
    jdff dff_B_9CMdKNfD5_2(.din(n28615), .dout(n28618));
    jdff dff_B_b8GLL0Nk3_2(.din(n28618), .dout(n28621));
    jdff dff_B_h7pYsV878_2(.din(n28621), .dout(n28624));
    jdff dff_B_lE00m7Z73_2(.din(n28624), .dout(n28627));
    jdff dff_B_eRPL2gmp0_2(.din(n28627), .dout(n28630));
    jdff dff_B_a6kvGCiD9_2(.din(n28630), .dout(n28633));
    jdff dff_B_L9TnrSUB8_2(.din(n28633), .dout(n28636));
    jdff dff_B_baOIVWVp9_2(.din(n28636), .dout(n28639));
    jdff dff_B_R8slybch4_2(.din(n28639), .dout(n28642));
    jdff dff_B_6hbSk1TN9_2(.din(n28642), .dout(n28645));
    jdff dff_B_ddo9L6QE0_2(.din(n28645), .dout(n28648));
    jdff dff_B_MczcRKuC2_2(.din(n28648), .dout(n28651));
    jdff dff_B_nvfTUSFu6_2(.din(n28651), .dout(n28654));
    jdff dff_B_Xiu0xkK29_2(.din(n28654), .dout(n28657));
    jdff dff_B_msSltTL19_2(.din(n4450), .dout(n28660));
    jdff dff_B_af6URBAC0_1(.din(n4388), .dout(n28663));
    jdff dff_B_oYP1l3rM5_2(.din(n3988), .dout(n28666));
    jdff dff_B_gRf78oQM8_2(.din(n28666), .dout(n28669));
    jdff dff_B_tgN7iGGJ7_2(.din(n28669), .dout(n28672));
    jdff dff_B_l7CesZvX9_2(.din(n28672), .dout(n28675));
    jdff dff_B_ezaZEJrp5_2(.din(n28675), .dout(n28678));
    jdff dff_B_RfHQRe791_2(.din(n28678), .dout(n28681));
    jdff dff_B_dsUBNTIy8_2(.din(n28681), .dout(n28684));
    jdff dff_B_nWAzqlwX2_2(.din(n28684), .dout(n28687));
    jdff dff_B_RaF2pSzQ5_2(.din(n28687), .dout(n28690));
    jdff dff_B_VZxdJc120_2(.din(n28690), .dout(n28693));
    jdff dff_B_L5Z5gPi44_2(.din(n28693), .dout(n28696));
    jdff dff_B_Px5rwGni0_2(.din(n28696), .dout(n28699));
    jdff dff_B_sbDZY1tI2_2(.din(n28699), .dout(n28702));
    jdff dff_B_WtGIh4183_2(.din(n28702), .dout(n28705));
    jdff dff_B_9P0YEedD2_2(.din(n28705), .dout(n28708));
    jdff dff_B_RSnN9Bqc6_2(.din(n4074), .dout(n28711));
    jdff dff_B_GbnFbinF7_2(.din(n28711), .dout(n28714));
    jdff dff_B_JdMX0b1g2_1(.din(n3992), .dout(n28717));
    jdff dff_B_eeCbMqGg7_2(.din(n3611), .dout(n28720));
    jdff dff_B_z1LRiTOE0_2(.din(n28720), .dout(n28723));
    jdff dff_B_gv3NYn6P6_2(.din(n28723), .dout(n28726));
    jdff dff_B_1ENQgEHy7_2(.din(n28726), .dout(n28729));
    jdff dff_B_vijbYQq07_2(.din(n28729), .dout(n28732));
    jdff dff_B_BhQpaSSH3_2(.din(n28732), .dout(n28735));
    jdff dff_B_CBo7bbq76_2(.din(n28735), .dout(n28738));
    jdff dff_B_JYBkCv3n7_2(.din(n28738), .dout(n28741));
    jdff dff_B_edUcnAT04_2(.din(n28741), .dout(n28744));
    jdff dff_B_yHYHauRk5_2(.din(n28744), .dout(n28747));
    jdff dff_B_eCVnUcVL2_2(.din(n28747), .dout(n28750));
    jdff dff_B_RN7mN8hd4_2(.din(n28750), .dout(n28753));
    jdff dff_B_DOAQMQjL2_2(.din(n3671), .dout(n28756));
    jdff dff_B_QkUk3v3e1_2(.din(n28756), .dout(n28759));
    jdff dff_B_PJf0cWwu9_1(.din(n3615), .dout(n28762));
    jdff dff_B_h9kLTsBE7_2(.din(n3210), .dout(n28765));
    jdff dff_B_3IuYWM1f7_2(.din(n28765), .dout(n28768));
    jdff dff_B_ZSeLQX9n7_2(.din(n28768), .dout(n28771));
    jdff dff_B_nGXJ12E88_2(.din(n28771), .dout(n28774));
    jdff dff_B_HdZ7ZILy2_2(.din(n28774), .dout(n28777));
    jdff dff_B_xWtGqVjE0_2(.din(n28777), .dout(n28780));
    jdff dff_B_aTqj50vP2_2(.din(n28780), .dout(n28783));
    jdff dff_B_FKjZDHFt8_2(.din(n28783), .dout(n28786));
    jdff dff_B_PJROlhI89_2(.din(n28786), .dout(n28789));
    jdff dff_B_WNF3HEs58_2(.din(n3269), .dout(n28792));
    jdff dff_B_6IN4EJlK2_2(.din(n28792), .dout(n28795));
    jdff dff_B_sYNSHnuN6_2(.din(n28795), .dout(n28798));
    jdff dff_B_yTJ3of4o1_1(.din(n3213), .dout(n28801));
    jdff dff_B_7Qv96jdo5_1(.din(n28801), .dout(n28804));
    jdff dff_B_qojY8BTd6_1(.din(n28804), .dout(n28807));
    jdff dff_B_3WH9b8qn6_1(.din(n28807), .dout(n28810));
    jdff dff_B_l0OJj6WW6_1(.din(n28810), .dout(n28813));
    jdff dff_B_Q36U5tAt1_1(.din(n28813), .dout(n28816));
    jdff dff_B_UmxfwUrb4_0(.din(n2864), .dout(n28819));
    jdff dff_B_l1FIUshX7_0(.din(n28819), .dout(n28822));
    jdff dff_A_IZ0xkOZa6_0(.din(n28827), .dout(n28824));
    jdff dff_A_Vp1im4IS8_0(.din(n28830), .dout(n28827));
    jdff dff_A_xxdJDKKt3_0(.din(n2860), .dout(n28830));
    jdff dff_B_fexZ1vyZ4_1(.din(n2838), .dout(n28834));
    jdff dff_A_PWnxLbLl4_0(.din(n2472), .dout(n28836));
    jdff dff_A_sW6BxUtj5_1(.din(n28842), .dout(n28839));
    jdff dff_A_j2EXnS4j2_1(.din(n2472), .dout(n28842));
    jdff dff_A_Bng07JI51_1(.din(n28848), .dout(n28845));
    jdff dff_A_DMRk3z007_1(.din(n28851), .dout(n28848));
    jdff dff_A_FPrhdtpG5_1(.din(n28854), .dout(n28851));
    jdff dff_A_kH63j8y58_1(.din(n28857), .dout(n28854));
    jdff dff_A_N3X0YXy17_1(.din(n28860), .dout(n28857));
    jdff dff_A_YFE1FYKA7_1(.din(n2830), .dout(n28860));
    jdff dff_B_G1Be0w1L8_1(.din(n6856), .dout(n28864));
    jdff dff_B_BJk9Dbvo7_1(.din(n6806), .dout(n28867));
    jdff dff_B_AxN3HC4J1_1(.din(n28867), .dout(n28870));
    jdff dff_B_9vMD6hbD0_2(.din(n6802), .dout(n28873));
    jdff dff_B_iR3Wwocn7_2(.din(n28873), .dout(n28876));
    jdff dff_B_y2CLNKJg3_2(.din(n28876), .dout(n28879));
    jdff dff_B_thMdE1km3_2(.din(n28879), .dout(n28882));
    jdff dff_B_gqRyL4kK8_2(.din(n28882), .dout(n28885));
    jdff dff_B_2A6sBGJO0_2(.din(n28885), .dout(n28888));
    jdff dff_B_1FX43Tc53_2(.din(n28888), .dout(n28891));
    jdff dff_B_6x2Ex84T7_2(.din(n28891), .dout(n28894));
    jdff dff_B_LYPyE8tY2_2(.din(n28894), .dout(n28897));
    jdff dff_B_zVhitRX36_2(.din(n28897), .dout(n28900));
    jdff dff_B_mtiAUmNd6_2(.din(n28900), .dout(n28903));
    jdff dff_B_7SoSryC90_2(.din(n28903), .dout(n28906));
    jdff dff_B_fP3eqyak0_2(.din(n28906), .dout(n28909));
    jdff dff_B_njOaAzGI0_2(.din(n28909), .dout(n28912));
    jdff dff_B_7tPl8Cjy8_2(.din(n28912), .dout(n28915));
    jdff dff_B_v8BIbjAg8_2(.din(n28915), .dout(n28918));
    jdff dff_B_StLRGRLP9_2(.din(n28918), .dout(n28921));
    jdff dff_B_QfVDqDwH8_2(.din(n28921), .dout(n28924));
    jdff dff_B_B3KWInmO7_2(.din(n28924), .dout(n28927));
    jdff dff_B_M7DCY9k03_2(.din(n28927), .dout(n28930));
    jdff dff_B_rAUwfWYI2_2(.din(n28930), .dout(n28933));
    jdff dff_B_52iviQen5_2(.din(n28933), .dout(n28936));
    jdff dff_B_nYhK47Pe4_2(.din(n28936), .dout(n28939));
    jdff dff_B_ETSoEChk3_2(.din(n28939), .dout(n28942));
    jdff dff_B_wJZ6jOMz5_2(.din(n28942), .dout(n28945));
    jdff dff_B_MnNlc0Ou7_2(.din(n28945), .dout(n28948));
    jdff dff_B_tEmivrTT0_2(.din(n28948), .dout(n28951));
    jdff dff_B_cE7dGaTG7_2(.din(n28951), .dout(n28954));
    jdff dff_B_eBmY3vh63_2(.din(n28954), .dout(n28957));
    jdff dff_B_UqrvQW5a4_2(.din(n28957), .dout(n28960));
    jdff dff_B_9S1WPhc23_2(.din(n28960), .dout(n28963));
    jdff dff_B_sgCui1Oh6_2(.din(n28963), .dout(n28966));
    jdff dff_B_dFFw3xfX4_2(.din(n28966), .dout(n28969));
    jdff dff_B_KykwPUDp1_2(.din(n28969), .dout(n28972));
    jdff dff_B_6nFXMZBp9_2(.din(n28972), .dout(n28975));
    jdff dff_B_Q4CBMmkC9_2(.din(n28975), .dout(n28978));
    jdff dff_B_UC5kuJaV0_2(.din(n28978), .dout(n28981));
    jdff dff_B_1fdUktiK4_2(.din(n28981), .dout(n28984));
    jdff dff_B_Pmflzgv54_2(.din(n28984), .dout(n28987));
    jdff dff_B_zhUTe2rp2_2(.din(n28987), .dout(n28990));
    jdff dff_B_D2PBaTFe8_2(.din(n28990), .dout(n28993));
    jdff dff_B_sH9z1PyZ3_2(.din(n28993), .dout(n28996));
    jdff dff_B_MvYL5r789_2(.din(n28996), .dout(n28999));
    jdff dff_B_5BFebvs10_2(.din(n28999), .dout(n29002));
    jdff dff_B_PULcOqeB0_2(.din(n29002), .dout(n29005));
    jdff dff_B_gXqmDAeT8_2(.din(n29005), .dout(n29008));
    jdff dff_B_xgFFtDeH6_2(.din(n29008), .dout(n29011));
    jdff dff_B_3H1iyCRn6_2(.din(n29011), .dout(n29014));
    jdff dff_B_06s29llU5_2(.din(n29014), .dout(n29017));
    jdff dff_B_NCg4KGXy8_2(.din(n29017), .dout(n29020));
    jdff dff_B_aDtcJ0ba2_2(.din(n29020), .dout(n29023));
    jdff dff_B_DBu9MS8x8_2(.din(n29023), .dout(n29026));
    jdff dff_B_WqK2XOQa0_2(.din(n29026), .dout(n29029));
    jdff dff_B_K12XMtUH4_2(.din(n29029), .dout(n29032));
    jdff dff_B_NX47Qo9X3_2(.din(n29032), .dout(n29035));
    jdff dff_B_1EHsxoj72_2(.din(n29035), .dout(n29038));
    jdff dff_B_XFzugYOA1_2(.din(n6798), .dout(n29041));
    jdff dff_B_T28lCIe81_2(.din(n29041), .dout(n29044));
    jdff dff_B_wkflulbq7_2(.din(n29044), .dout(n29047));
    jdff dff_B_U5frjtpA6_2(.din(n29047), .dout(n29050));
    jdff dff_B_O6i7BYTM1_2(.din(n29050), .dout(n29053));
    jdff dff_B_rwByXSln1_2(.din(n29053), .dout(n29056));
    jdff dff_B_rtwrQ7Tv5_2(.din(n29056), .dout(n29059));
    jdff dff_B_HDbnImm39_2(.din(n29059), .dout(n29062));
    jdff dff_B_AaMS8tfn6_2(.din(n29062), .dout(n29065));
    jdff dff_B_pVk1HtIl5_2(.din(n29065), .dout(n29068));
    jdff dff_B_FAc6RLLw4_2(.din(n29068), .dout(n29071));
    jdff dff_B_1TFpC6D21_2(.din(n29071), .dout(n29074));
    jdff dff_B_PfAeb9oB3_2(.din(n29074), .dout(n29077));
    jdff dff_B_MVQii1Gd8_2(.din(n29077), .dout(n29080));
    jdff dff_B_Djsn6kpn7_2(.din(n29080), .dout(n29083));
    jdff dff_B_xexikIMK3_2(.din(n29083), .dout(n29086));
    jdff dff_B_ggMbpQ1Y0_2(.din(n29086), .dout(n29089));
    jdff dff_B_vCgWseQY3_2(.din(n29089), .dout(n29092));
    jdff dff_B_JdEPa84d2_2(.din(n29092), .dout(n29095));
    jdff dff_B_4BkPHsBH0_2(.din(n29095), .dout(n29098));
    jdff dff_B_vHAFnp5x2_2(.din(n29098), .dout(n29101));
    jdff dff_B_nBcdnM9J5_2(.din(n29101), .dout(n29104));
    jdff dff_B_mqHpdWmB4_2(.din(n29104), .dout(n29107));
    jdff dff_B_XxhIOBW03_2(.din(n29107), .dout(n29110));
    jdff dff_B_YerTaQ5M3_2(.din(n29110), .dout(n29113));
    jdff dff_B_5qeh0qTg4_2(.din(n29113), .dout(n29116));
    jdff dff_B_N5mK56Ne9_2(.din(n29116), .dout(n29119));
    jdff dff_B_YvHSALV81_2(.din(n29119), .dout(n29122));
    jdff dff_B_SVjep5Kl0_2(.din(n29122), .dout(n29125));
    jdff dff_B_i2mWbpK86_2(.din(n29125), .dout(n29128));
    jdff dff_B_FxwMyqUs3_2(.din(n29128), .dout(n29131));
    jdff dff_B_cxmOkPJ61_2(.din(n29131), .dout(n29134));
    jdff dff_B_dyIoaoXw8_2(.din(n29134), .dout(n29137));
    jdff dff_B_SflPcyWR9_2(.din(n29137), .dout(n29140));
    jdff dff_B_jrItXETU6_2(.din(n29140), .dout(n29143));
    jdff dff_B_WK2EgIWG3_2(.din(n29143), .dout(n29146));
    jdff dff_B_xFAOHMdw9_2(.din(n29146), .dout(n29149));
    jdff dff_B_dhnAj0hT9_2(.din(n29149), .dout(n29152));
    jdff dff_B_QTDhhjWn0_2(.din(n29152), .dout(n29155));
    jdff dff_B_lN3EfoVL0_2(.din(n29155), .dout(n29158));
    jdff dff_B_8s5o3v5U4_2(.din(n29158), .dout(n29161));
    jdff dff_B_qde6tAky2_2(.din(n29161), .dout(n29164));
    jdff dff_B_In3gVkjm5_2(.din(n29164), .dout(n29167));
    jdff dff_B_STu83squ6_2(.din(n29167), .dout(n29170));
    jdff dff_B_gfdF8Odu5_2(.din(n29170), .dout(n29173));
    jdff dff_B_oyiBnt7S7_2(.din(n29173), .dout(n29176));
    jdff dff_B_ix5DV3Pj9_2(.din(n29176), .dout(n29179));
    jdff dff_B_DQziWUWh7_2(.din(n29179), .dout(n29182));
    jdff dff_B_tKKdVf3h6_2(.din(n29182), .dout(n29185));
    jdff dff_B_ZnvyxNqF0_2(.din(n29185), .dout(n29188));
    jdff dff_B_bVUR7K3M1_2(.din(n29188), .dout(n29191));
    jdff dff_B_NfQ7qjpF1_2(.din(n29191), .dout(n29194));
    jdff dff_B_KvjGBq3E4_2(.din(n29194), .dout(n29197));
    jdff dff_B_PFWPYXhD6_2(.din(n29197), .dout(n29200));
    jdff dff_B_JwSfpbBe7_2(.din(n29200), .dout(n29203));
    jdff dff_B_JRF5aHui3_2(.din(n29203), .dout(n29206));
    jdff dff_B_n6ngT6Yo2_2(.din(n29206), .dout(n29209));
    jdff dff_B_eP2sF8fc1_2(.din(n29209), .dout(n29212));
    jdff dff_A_Gl0YM9RQ1_1(.din(n6794), .dout(n29214));
    jdff dff_B_mgjKK9GJ3_1(.din(n6786), .dout(n29218));
    jdff dff_B_SCL5FPKf3_2(.din(n6702), .dout(n29221));
    jdff dff_B_rzXmh0BJ1_2(.din(n29221), .dout(n29224));
    jdff dff_B_qeZt0Tgx5_2(.din(n29224), .dout(n29227));
    jdff dff_B_f3WvnnPU4_2(.din(n29227), .dout(n29230));
    jdff dff_B_NyTNzeqe7_2(.din(n29230), .dout(n29233));
    jdff dff_B_bu82JbmM1_2(.din(n29233), .dout(n29236));
    jdff dff_B_PtMZMIJq2_2(.din(n29236), .dout(n29239));
    jdff dff_B_iAqmL0DB6_2(.din(n29239), .dout(n29242));
    jdff dff_B_ljIttL9l9_2(.din(n29242), .dout(n29245));
    jdff dff_B_nxCSWGlt7_2(.din(n29245), .dout(n29248));
    jdff dff_B_qwNFtUbC2_2(.din(n29248), .dout(n29251));
    jdff dff_B_eX9ZyAfw3_2(.din(n29251), .dout(n29254));
    jdff dff_B_d40C5jOH5_2(.din(n29254), .dout(n29257));
    jdff dff_B_QYCke47w0_2(.din(n29257), .dout(n29260));
    jdff dff_B_O7ZtqB7H8_2(.din(n29260), .dout(n29263));
    jdff dff_B_buJwVWIL1_2(.din(n29263), .dout(n29266));
    jdff dff_B_4wdRDvXP7_2(.din(n29266), .dout(n29269));
    jdff dff_B_M027ArTJ2_2(.din(n29269), .dout(n29272));
    jdff dff_B_IgbOy04R6_2(.din(n29272), .dout(n29275));
    jdff dff_B_JKKOcUY14_2(.din(n29275), .dout(n29278));
    jdff dff_B_uOyyPRu64_2(.din(n29278), .dout(n29281));
    jdff dff_B_Qq5pQ5Py1_2(.din(n29281), .dout(n29284));
    jdff dff_B_RNL4Jt5w8_2(.din(n29284), .dout(n29287));
    jdff dff_B_mDVG1MSg6_2(.din(n29287), .dout(n29290));
    jdff dff_B_qPSvWAOh0_2(.din(n29290), .dout(n29293));
    jdff dff_B_0OTCxfDP5_2(.din(n29293), .dout(n29296));
    jdff dff_B_e3nTQoLs9_2(.din(n29296), .dout(n29299));
    jdff dff_B_tpHaKlcI8_2(.din(n29299), .dout(n29302));
    jdff dff_B_2ux7tTVC2_2(.din(n29302), .dout(n29305));
    jdff dff_B_pVz0MthM3_2(.din(n29305), .dout(n29308));
    jdff dff_B_xpITjV6J8_2(.din(n29308), .dout(n29311));
    jdff dff_B_zCFukkEW2_2(.din(n29311), .dout(n29314));
    jdff dff_B_6GVByEGo9_2(.din(n29314), .dout(n29317));
    jdff dff_B_PzF4wiI91_2(.din(n29317), .dout(n29320));
    jdff dff_B_PZRbMNPF1_2(.din(n29320), .dout(n29323));
    jdff dff_B_wE8M9pSE6_2(.din(n29323), .dout(n29326));
    jdff dff_B_sxF7Nnto4_2(.din(n29326), .dout(n29329));
    jdff dff_B_0s4hG60m4_2(.din(n29329), .dout(n29332));
    jdff dff_B_5h7NepSj5_2(.din(n29332), .dout(n29335));
    jdff dff_B_pop4QW1h9_2(.din(n29335), .dout(n29338));
    jdff dff_B_upAQuHGD9_2(.din(n29338), .dout(n29341));
    jdff dff_B_vnGnmv5D6_2(.din(n29341), .dout(n29344));
    jdff dff_B_WsEJNZR41_2(.din(n29344), .dout(n29347));
    jdff dff_B_t8NUpRFL8_2(.din(n29347), .dout(n29350));
    jdff dff_B_n4UBlc7K0_2(.din(n29350), .dout(n29353));
    jdff dff_B_9QpmV5qC5_2(.din(n29353), .dout(n29356));
    jdff dff_B_LTNHYBTm5_2(.din(n29356), .dout(n29359));
    jdff dff_B_yZxKMZrc0_2(.din(n29359), .dout(n29362));
    jdff dff_B_t5UhvOzR9_2(.din(n29362), .dout(n29365));
    jdff dff_B_u4xfTwzc5_2(.din(n29365), .dout(n29368));
    jdff dff_B_f5WMARNu2_2(.din(n29368), .dout(n29371));
    jdff dff_B_kqOINCaK6_2(.din(n29371), .dout(n29374));
    jdff dff_B_pZhfJMe73_2(.din(n29374), .dout(n29377));
    jdff dff_B_DDLXVTVi5_2(.din(n29377), .dout(n29380));
    jdff dff_B_iy3NUKPE5_2(.din(n29380), .dout(n29383));
    jdff dff_B_C5PFZR9b4_1(.din(n6726), .dout(n29386));
    jdff dff_B_HF7UIH5v7_1(.din(n29386), .dout(n29389));
    jdff dff_B_wHsykZ4H0_2(.din(n6722), .dout(n29392));
    jdff dff_B_zhuPOkfj8_2(.din(n29392), .dout(n29395));
    jdff dff_B_0XaTQvYi4_2(.din(n29395), .dout(n29398));
    jdff dff_B_yDLhR7300_2(.din(n29398), .dout(n29401));
    jdff dff_B_Eex5LyVM5_2(.din(n29401), .dout(n29404));
    jdff dff_B_6ZvvSzvv7_2(.din(n29404), .dout(n29407));
    jdff dff_B_U9JaiPV90_2(.din(n29407), .dout(n29410));
    jdff dff_B_3HEWHJvJ7_2(.din(n29410), .dout(n29413));
    jdff dff_B_5tC6oTRG6_2(.din(n29413), .dout(n29416));
    jdff dff_B_kaXIRbLv3_2(.din(n29416), .dout(n29419));
    jdff dff_B_CP6JXgNu9_2(.din(n29419), .dout(n29422));
    jdff dff_B_gzs4q0lq2_2(.din(n29422), .dout(n29425));
    jdff dff_B_3esntLel3_2(.din(n29425), .dout(n29428));
    jdff dff_B_V4mb45DA0_2(.din(n29428), .dout(n29431));
    jdff dff_B_BelUqyhy5_2(.din(n29431), .dout(n29434));
    jdff dff_B_6H5KFKj60_2(.din(n29434), .dout(n29437));
    jdff dff_B_s8QpbDgg2_2(.din(n29437), .dout(n29440));
    jdff dff_B_U7g7E0915_2(.din(n29440), .dout(n29443));
    jdff dff_B_HQwyle1y5_2(.din(n29443), .dout(n29446));
    jdff dff_B_0TwLzO5A5_2(.din(n29446), .dout(n29449));
    jdff dff_B_jmKALU6T0_2(.din(n29449), .dout(n29452));
    jdff dff_B_eBUFuLKM9_2(.din(n29452), .dout(n29455));
    jdff dff_B_33O9jhYA3_2(.din(n29455), .dout(n29458));
    jdff dff_B_YJDYGVz93_2(.din(n29458), .dout(n29461));
    jdff dff_B_pG3Im42M8_2(.din(n29461), .dout(n29464));
    jdff dff_B_IST5TWf49_2(.din(n29464), .dout(n29467));
    jdff dff_B_Tl1UPHVz1_2(.din(n29467), .dout(n29470));
    jdff dff_B_oNE4NWWT9_2(.din(n29470), .dout(n29473));
    jdff dff_B_lyFbzixm0_2(.din(n29473), .dout(n29476));
    jdff dff_B_TocHg3WY7_2(.din(n29476), .dout(n29479));
    jdff dff_B_3cBaZWW75_2(.din(n29479), .dout(n29482));
    jdff dff_B_SDyoQ5iT4_2(.din(n29482), .dout(n29485));
    jdff dff_B_64TKNjo47_2(.din(n29485), .dout(n29488));
    jdff dff_B_uyHq7NzC1_2(.din(n29488), .dout(n29491));
    jdff dff_B_ZoiUq8a02_2(.din(n29491), .dout(n29494));
    jdff dff_B_Ba850tM69_2(.din(n29494), .dout(n29497));
    jdff dff_B_mnXNmXzB8_2(.din(n29497), .dout(n29500));
    jdff dff_B_4gS6xnRA7_2(.din(n29500), .dout(n29503));
    jdff dff_B_EbhUxANj2_2(.din(n29503), .dout(n29506));
    jdff dff_B_vuE5VV8D4_2(.din(n29506), .dout(n29509));
    jdff dff_B_eT333xhz5_2(.din(n29509), .dout(n29512));
    jdff dff_B_467KL0ma9_2(.din(n29512), .dout(n29515));
    jdff dff_B_0qy5Wpy23_2(.din(n29515), .dout(n29518));
    jdff dff_B_eFqEJzwg6_2(.din(n29518), .dout(n29521));
    jdff dff_B_a8QS7p6D1_2(.din(n29521), .dout(n29524));
    jdff dff_B_QPsg3qiV0_2(.din(n29524), .dout(n29527));
    jdff dff_B_VjQUnkm02_2(.din(n29527), .dout(n29530));
    jdff dff_B_Xv7fqjh14_2(.din(n29530), .dout(n29533));
    jdff dff_B_KY5ozMdg9_2(.din(n29533), .dout(n29536));
    jdff dff_B_fD031rCq7_2(.din(n29536), .dout(n29539));
    jdff dff_B_E57eyS4L2_2(.din(n29539), .dout(n29542));
    jdff dff_B_qDLH0N856_2(.din(n29542), .dout(n29545));
    jdff dff_B_2fPJuVhx8_2(.din(n6718), .dout(n29548));
    jdff dff_B_7dzdvXTd5_2(.din(n29548), .dout(n29551));
    jdff dff_B_0VyNcSpR3_2(.din(n29551), .dout(n29554));
    jdff dff_B_1P0ZU3AO1_2(.din(n29554), .dout(n29557));
    jdff dff_B_9eR9o1238_2(.din(n29557), .dout(n29560));
    jdff dff_B_Lt9yd9Dk1_2(.din(n29560), .dout(n29563));
    jdff dff_B_UuhZQnPW4_2(.din(n29563), .dout(n29566));
    jdff dff_B_bYhuYC8K5_2(.din(n29566), .dout(n29569));
    jdff dff_B_tCOv0GtU3_2(.din(n29569), .dout(n29572));
    jdff dff_B_LkK62bDd0_2(.din(n29572), .dout(n29575));
    jdff dff_B_FdqfFCXn2_2(.din(n29575), .dout(n29578));
    jdff dff_B_hxVovnc37_2(.din(n29578), .dout(n29581));
    jdff dff_B_tFMXEZ056_2(.din(n29581), .dout(n29584));
    jdff dff_B_YG1uLtQO4_2(.din(n29584), .dout(n29587));
    jdff dff_B_NIhudi1f7_2(.din(n29587), .dout(n29590));
    jdff dff_B_FBxUjoSz5_2(.din(n29590), .dout(n29593));
    jdff dff_B_c7fpcYcG8_2(.din(n29593), .dout(n29596));
    jdff dff_B_5NAKAHfi0_2(.din(n29596), .dout(n29599));
    jdff dff_B_P6j1z3zi3_2(.din(n29599), .dout(n29602));
    jdff dff_B_eaU1Od7X3_2(.din(n29602), .dout(n29605));
    jdff dff_B_luTLKIV70_2(.din(n29605), .dout(n29608));
    jdff dff_B_czYanEhE8_2(.din(n29608), .dout(n29611));
    jdff dff_B_X6ighRgX3_2(.din(n29611), .dout(n29614));
    jdff dff_B_asnk09Ta4_2(.din(n29614), .dout(n29617));
    jdff dff_B_ijlB5QAU4_2(.din(n29617), .dout(n29620));
    jdff dff_B_hmkodBnU9_2(.din(n29620), .dout(n29623));
    jdff dff_B_9m5MlGyv0_2(.din(n29623), .dout(n29626));
    jdff dff_B_oEHLFViE1_2(.din(n29626), .dout(n29629));
    jdff dff_B_7IopQFbk8_2(.din(n29629), .dout(n29632));
    jdff dff_B_FJXngTPx4_2(.din(n29632), .dout(n29635));
    jdff dff_B_CcvmYj4K1_2(.din(n29635), .dout(n29638));
    jdff dff_B_IcljosVj9_2(.din(n29638), .dout(n29641));
    jdff dff_B_D3OS0tOl8_2(.din(n29641), .dout(n29644));
    jdff dff_B_vLq7xXXe6_2(.din(n29644), .dout(n29647));
    jdff dff_B_Cxlbn2YH1_2(.din(n29647), .dout(n29650));
    jdff dff_B_bYDkw8ey7_2(.din(n29650), .dout(n29653));
    jdff dff_B_YsVtuTww3_2(.din(n29653), .dout(n29656));
    jdff dff_B_zeQHvMfS1_2(.din(n29656), .dout(n29659));
    jdff dff_B_xh3h0ZTH5_2(.din(n29659), .dout(n29662));
    jdff dff_B_Bxbj5GNR9_2(.din(n29662), .dout(n29665));
    jdff dff_B_DDQoObtD0_2(.din(n29665), .dout(n29668));
    jdff dff_B_WPWPEX9p4_2(.din(n29668), .dout(n29671));
    jdff dff_B_qe5l42G07_2(.din(n29671), .dout(n29674));
    jdff dff_B_5NwC0zyT1_2(.din(n29674), .dout(n29677));
    jdff dff_B_XMJKtRfu1_2(.din(n29677), .dout(n29680));
    jdff dff_B_gPYNN6We1_2(.din(n29680), .dout(n29683));
    jdff dff_B_4X61qpGa9_2(.din(n29683), .dout(n29686));
    jdff dff_B_g88UkIkL3_2(.din(n29686), .dout(n29689));
    jdff dff_B_xm3ajwH93_2(.din(n29689), .dout(n29692));
    jdff dff_B_LgYseWrf1_2(.din(n29692), .dout(n29695));
    jdff dff_B_fwwxPM7b0_2(.din(n29695), .dout(n29698));
    jdff dff_B_oawvuwEe3_2(.din(n29698), .dout(n29701));
    jdff dff_B_smj7f7QK1_2(.din(n29701), .dout(n29704));
    jdff dff_B_eAyBbxsi5_2(.din(n29704), .dout(n29707));
    jdff dff_B_qwcLaNmX5_2(.din(n6714), .dout(n29710));
    jdff dff_B_DCVTibQ27_1(.din(n6706), .dout(n29713));
    jdff dff_B_mBr9zinK6_2(.din(n6595), .dout(n29716));
    jdff dff_B_LULJaJzn4_2(.din(n29716), .dout(n29719));
    jdff dff_B_sUAEr5C76_2(.din(n29719), .dout(n29722));
    jdff dff_B_7O0dQzBl7_2(.din(n29722), .dout(n29725));
    jdff dff_B_2bRqSR7K4_2(.din(n29725), .dout(n29728));
    jdff dff_B_9oiuXmBM5_2(.din(n29728), .dout(n29731));
    jdff dff_B_CWyPJmsp1_2(.din(n29731), .dout(n29734));
    jdff dff_B_JQClPjCb6_2(.din(n29734), .dout(n29737));
    jdff dff_B_vmLGuPmO0_2(.din(n29737), .dout(n29740));
    jdff dff_B_M3aP8gb95_2(.din(n29740), .dout(n29743));
    jdff dff_B_wV5zPB190_2(.din(n29743), .dout(n29746));
    jdff dff_B_sjcZzzYF5_2(.din(n29746), .dout(n29749));
    jdff dff_B_430T1Hu07_2(.din(n29749), .dout(n29752));
    jdff dff_B_W97Gox2J2_2(.din(n29752), .dout(n29755));
    jdff dff_B_y0f3K5dY3_2(.din(n29755), .dout(n29758));
    jdff dff_B_6msuEzT60_2(.din(n29758), .dout(n29761));
    jdff dff_B_b4ApuG0W5_2(.din(n29761), .dout(n29764));
    jdff dff_B_f0i7id6f0_2(.din(n29764), .dout(n29767));
    jdff dff_B_fy0ZoZUL7_2(.din(n29767), .dout(n29770));
    jdff dff_B_DjY4juBD1_2(.din(n29770), .dout(n29773));
    jdff dff_B_NP1GV6ld1_2(.din(n29773), .dout(n29776));
    jdff dff_B_paD3DpxO7_2(.din(n29776), .dout(n29779));
    jdff dff_B_sDHHtcpz7_2(.din(n29779), .dout(n29782));
    jdff dff_B_wjppf0Bc1_2(.din(n29782), .dout(n29785));
    jdff dff_B_lbLrs8LF4_2(.din(n29785), .dout(n29788));
    jdff dff_B_L0DmwOYo7_2(.din(n29788), .dout(n29791));
    jdff dff_B_Ft5TVyL50_2(.din(n29791), .dout(n29794));
    jdff dff_B_9aue72Ua0_2(.din(n29794), .dout(n29797));
    jdff dff_B_cIwxU3zM3_2(.din(n29797), .dout(n29800));
    jdff dff_B_RHqIKApR7_2(.din(n29800), .dout(n29803));
    jdff dff_B_ujN89r0g6_2(.din(n29803), .dout(n29806));
    jdff dff_B_wvxQYmri1_2(.din(n29806), .dout(n29809));
    jdff dff_B_ePiEQjG64_2(.din(n29809), .dout(n29812));
    jdff dff_B_GrU9M4Jm8_2(.din(n29812), .dout(n29815));
    jdff dff_B_6f4JRWgK8_2(.din(n29815), .dout(n29818));
    jdff dff_B_D5mwCWO32_2(.din(n29818), .dout(n29821));
    jdff dff_B_xl4p3TSt5_2(.din(n29821), .dout(n29824));
    jdff dff_B_9GkEsjpZ8_2(.din(n29824), .dout(n29827));
    jdff dff_B_lAUcFlBh4_2(.din(n29827), .dout(n29830));
    jdff dff_B_DOaNXmBB7_2(.din(n29830), .dout(n29833));
    jdff dff_B_2MlMu2sh8_2(.din(n29833), .dout(n29836));
    jdff dff_B_74oQAdo70_2(.din(n29836), .dout(n29839));
    jdff dff_B_3wHcWuwi0_2(.din(n29839), .dout(n29842));
    jdff dff_B_R67BSxLW1_2(.din(n29842), .dout(n29845));
    jdff dff_B_Vw8N4D9R7_2(.din(n29845), .dout(n29848));
    jdff dff_B_00ZDp0qO0_2(.din(n29848), .dout(n29851));
    jdff dff_B_52nWTJBW9_2(.din(n29851), .dout(n29854));
    jdff dff_B_gh6p9pkQ1_2(.din(n29854), .dout(n29857));
    jdff dff_B_ov1qn2jK9_2(.din(n29857), .dout(n29860));
    jdff dff_B_gKuxhXwY3_2(.din(n29860), .dout(n29863));
    jdff dff_B_KRSHZt2L9_2(.din(n29863), .dout(n29866));
    jdff dff_B_1pa574RV7_1(.din(n6619), .dout(n29869));
    jdff dff_B_ab685Q2h6_1(.din(n29869), .dout(n29872));
    jdff dff_B_ZTQGXS6I4_2(.din(n6615), .dout(n29875));
    jdff dff_B_Lx3mjdSi3_2(.din(n29875), .dout(n29878));
    jdff dff_B_2yMd3pmf8_2(.din(n29878), .dout(n29881));
    jdff dff_B_GvLXw1Dy4_2(.din(n29881), .dout(n29884));
    jdff dff_B_Y34VWZRz1_2(.din(n29884), .dout(n29887));
    jdff dff_B_ASvUhJ8E6_2(.din(n29887), .dout(n29890));
    jdff dff_B_0DR97vdd7_2(.din(n29890), .dout(n29893));
    jdff dff_B_mhEG4gnA9_2(.din(n29893), .dout(n29896));
    jdff dff_B_NiVKBVR14_2(.din(n29896), .dout(n29899));
    jdff dff_B_zg14c5Ki7_2(.din(n29899), .dout(n29902));
    jdff dff_B_KW35wHnr4_2(.din(n29902), .dout(n29905));
    jdff dff_B_Lr2extkt9_2(.din(n29905), .dout(n29908));
    jdff dff_B_dTuSMScV1_2(.din(n29908), .dout(n29911));
    jdff dff_B_HUyS1SZJ5_2(.din(n29911), .dout(n29914));
    jdff dff_B_wi4EoFSo0_2(.din(n29914), .dout(n29917));
    jdff dff_B_JBWjeKvm9_2(.din(n29917), .dout(n29920));
    jdff dff_B_nPHj5vVo7_2(.din(n29920), .dout(n29923));
    jdff dff_B_zboqbU9m7_2(.din(n29923), .dout(n29926));
    jdff dff_B_Dpr5pW0F1_2(.din(n29926), .dout(n29929));
    jdff dff_B_4Rt9FTG91_2(.din(n29929), .dout(n29932));
    jdff dff_B_poSUiAYG0_2(.din(n29932), .dout(n29935));
    jdff dff_B_kIyNPvVA4_2(.din(n29935), .dout(n29938));
    jdff dff_B_jTSwfXPJ8_2(.din(n29938), .dout(n29941));
    jdff dff_B_nOxYfUo26_2(.din(n29941), .dout(n29944));
    jdff dff_B_h8cPlX6y5_2(.din(n29944), .dout(n29947));
    jdff dff_B_WPqMUme29_2(.din(n29947), .dout(n29950));
    jdff dff_B_MI5UAQtl8_2(.din(n29950), .dout(n29953));
    jdff dff_B_WRtTMCzU1_2(.din(n29953), .dout(n29956));
    jdff dff_B_5n4V0OA64_2(.din(n29956), .dout(n29959));
    jdff dff_B_O4WLllGz5_2(.din(n29959), .dout(n29962));
    jdff dff_B_qP2Freca0_2(.din(n29962), .dout(n29965));
    jdff dff_B_aYAGfY9R4_2(.din(n29965), .dout(n29968));
    jdff dff_B_HQbZyGRz8_2(.din(n29968), .dout(n29971));
    jdff dff_B_6XQUihbW8_2(.din(n29971), .dout(n29974));
    jdff dff_B_Hn32oo9u0_2(.din(n29974), .dout(n29977));
    jdff dff_B_aYmWKJlS1_2(.din(n29977), .dout(n29980));
    jdff dff_B_RddqjjSj7_2(.din(n29980), .dout(n29983));
    jdff dff_B_KzTHHdTZ9_2(.din(n29983), .dout(n29986));
    jdff dff_B_LQMIU07m6_2(.din(n29986), .dout(n29989));
    jdff dff_B_ANxyz6Kb5_2(.din(n29989), .dout(n29992));
    jdff dff_B_NCvwvwDQ1_2(.din(n29992), .dout(n29995));
    jdff dff_B_8ZyEKesh8_2(.din(n29995), .dout(n29998));
    jdff dff_B_12TJV3oR1_2(.din(n29998), .dout(n30001));
    jdff dff_B_6pviUdXw0_2(.din(n30001), .dout(n30004));
    jdff dff_B_Lgp6UKpm6_2(.din(n30004), .dout(n30007));
    jdff dff_B_vPpUmE0L7_2(.din(n30007), .dout(n30010));
    jdff dff_B_JTOL4DZN6_2(.din(n30010), .dout(n30013));
    jdff dff_B_T0DnmlcE6_2(.din(n30013), .dout(n30016));
    jdff dff_B_UTRszQtn2_2(.din(n6611), .dout(n30019));
    jdff dff_B_Cr8357xq0_2(.din(n30019), .dout(n30022));
    jdff dff_B_QZf6fSZk6_2(.din(n30022), .dout(n30025));
    jdff dff_B_KPhStNhc8_2(.din(n30025), .dout(n30028));
    jdff dff_B_vWPu9wjV8_2(.din(n30028), .dout(n30031));
    jdff dff_B_YYYBmQsF7_2(.din(n30031), .dout(n30034));
    jdff dff_B_ePWIeJ7V6_2(.din(n30034), .dout(n30037));
    jdff dff_B_bzgpolVd7_2(.din(n30037), .dout(n30040));
    jdff dff_B_JbbDq3Bd9_2(.din(n30040), .dout(n30043));
    jdff dff_B_05NofmFR7_2(.din(n30043), .dout(n30046));
    jdff dff_B_grb6c2iX6_2(.din(n30046), .dout(n30049));
    jdff dff_B_3T42BwSA4_2(.din(n30049), .dout(n30052));
    jdff dff_B_6MX5TUvy2_2(.din(n30052), .dout(n30055));
    jdff dff_B_vhJlguC05_2(.din(n30055), .dout(n30058));
    jdff dff_B_e7b6DkQD1_2(.din(n30058), .dout(n30061));
    jdff dff_B_Jlhw6XOj4_2(.din(n30061), .dout(n30064));
    jdff dff_B_BztSFJGT6_2(.din(n30064), .dout(n30067));
    jdff dff_B_WCvndrbo4_2(.din(n30067), .dout(n30070));
    jdff dff_B_O0eLY8gG7_2(.din(n30070), .dout(n30073));
    jdff dff_B_XRz4o72X2_2(.din(n30073), .dout(n30076));
    jdff dff_B_gdE9GhUH5_2(.din(n30076), .dout(n30079));
    jdff dff_B_owaIawDw8_2(.din(n30079), .dout(n30082));
    jdff dff_B_4DSfg6gF5_2(.din(n30082), .dout(n30085));
    jdff dff_B_2NbcAh0T1_2(.din(n30085), .dout(n30088));
    jdff dff_B_gdSaeRLj7_2(.din(n30088), .dout(n30091));
    jdff dff_B_9HrCLUZ11_2(.din(n30091), .dout(n30094));
    jdff dff_B_pm2HzBRZ3_2(.din(n30094), .dout(n30097));
    jdff dff_B_bGsG0aH45_2(.din(n30097), .dout(n30100));
    jdff dff_B_4EO0Me7n0_2(.din(n30100), .dout(n30103));
    jdff dff_B_xAwSMO3D1_2(.din(n30103), .dout(n30106));
    jdff dff_B_z2EjJ4dY6_2(.din(n30106), .dout(n30109));
    jdff dff_B_WsrsDtnA7_2(.din(n30109), .dout(n30112));
    jdff dff_B_Njbn7fqq4_2(.din(n30112), .dout(n30115));
    jdff dff_B_5El2Biyu2_2(.din(n30115), .dout(n30118));
    jdff dff_B_bYCIXVhK1_2(.din(n30118), .dout(n30121));
    jdff dff_B_Yq0xn5UJ7_2(.din(n30121), .dout(n30124));
    jdff dff_B_Sxnc3k794_2(.din(n30124), .dout(n30127));
    jdff dff_B_WM4jHbNO0_2(.din(n30127), .dout(n30130));
    jdff dff_B_8k2UQPcp3_2(.din(n30130), .dout(n30133));
    jdff dff_B_CQGVIHtp5_2(.din(n30133), .dout(n30136));
    jdff dff_B_WqHq0ZFJ8_2(.din(n30136), .dout(n30139));
    jdff dff_B_awSFrf515_2(.din(n30139), .dout(n30142));
    jdff dff_B_rlXqutju2_2(.din(n30142), .dout(n30145));
    jdff dff_B_inKx7PGA4_2(.din(n30145), .dout(n30148));
    jdff dff_B_RWuu1e251_2(.din(n30148), .dout(n30151));
    jdff dff_B_5rGmhKVO8_2(.din(n30151), .dout(n30154));
    jdff dff_B_dzzTHMoz6_2(.din(n30154), .dout(n30157));
    jdff dff_B_eIn0hFC26_2(.din(n30157), .dout(n30160));
    jdff dff_B_DigdRgnJ2_2(.din(n30160), .dout(n30163));
    jdff dff_B_qFmd4odf4_2(.din(n30163), .dout(n30166));
    jdff dff_B_agF8t62T8_2(.din(n6607), .dout(n30169));
    jdff dff_B_3hVnrSk46_1(.din(n6599), .dout(n30172));
    jdff dff_B_5T2MMC6t4_2(.din(n6461), .dout(n30175));
    jdff dff_B_jHJYw1tZ2_2(.din(n30175), .dout(n30178));
    jdff dff_B_ipwt0XsT6_2(.din(n30178), .dout(n30181));
    jdff dff_B_1eZUEalB9_2(.din(n30181), .dout(n30184));
    jdff dff_B_ZLREOlSh2_2(.din(n30184), .dout(n30187));
    jdff dff_B_3WHtvTS26_2(.din(n30187), .dout(n30190));
    jdff dff_B_r3UPrdIk0_2(.din(n30190), .dout(n30193));
    jdff dff_B_30ZujImX2_2(.din(n30193), .dout(n30196));
    jdff dff_B_LuAgpGXj1_2(.din(n30196), .dout(n30199));
    jdff dff_B_CueCAGRS1_2(.din(n30199), .dout(n30202));
    jdff dff_B_rR8nMODP8_2(.din(n30202), .dout(n30205));
    jdff dff_B_vlA4WHrT9_2(.din(n30205), .dout(n30208));
    jdff dff_B_hNPXYkr54_2(.din(n30208), .dout(n30211));
    jdff dff_B_CbJP7g9z3_2(.din(n30211), .dout(n30214));
    jdff dff_B_l7GiGpvr5_2(.din(n30214), .dout(n30217));
    jdff dff_B_TlmxsKRL8_2(.din(n30217), .dout(n30220));
    jdff dff_B_9TkOdnhg8_2(.din(n30220), .dout(n30223));
    jdff dff_B_o0H4G08Y3_2(.din(n30223), .dout(n30226));
    jdff dff_B_XlcvIfD08_2(.din(n30226), .dout(n30229));
    jdff dff_B_Rmq9Dlrt6_2(.din(n30229), .dout(n30232));
    jdff dff_B_fu5VFzlx7_2(.din(n30232), .dout(n30235));
    jdff dff_B_wIA6K3Ev7_2(.din(n30235), .dout(n30238));
    jdff dff_B_ub2kmoWX3_2(.din(n30238), .dout(n30241));
    jdff dff_B_U2zk2YV07_2(.din(n30241), .dout(n30244));
    jdff dff_B_aYTXs1Rt6_2(.din(n30244), .dout(n30247));
    jdff dff_B_4RGwT7B56_2(.din(n30247), .dout(n30250));
    jdff dff_B_opA2uA8u9_2(.din(n30250), .dout(n30253));
    jdff dff_B_znimIONV6_2(.din(n30253), .dout(n30256));
    jdff dff_B_0Is8eCHY6_2(.din(n30256), .dout(n30259));
    jdff dff_B_tqvDZqSD6_2(.din(n30259), .dout(n30262));
    jdff dff_B_fO3nrgpd7_2(.din(n30262), .dout(n30265));
    jdff dff_B_bVnvuLRV5_2(.din(n30265), .dout(n30268));
    jdff dff_B_peI1zMN58_2(.din(n30268), .dout(n30271));
    jdff dff_B_uVS5ZH7X4_2(.din(n30271), .dout(n30274));
    jdff dff_B_m8kkNvOa9_2(.din(n30274), .dout(n30277));
    jdff dff_B_zMTkOWJj4_2(.din(n30277), .dout(n30280));
    jdff dff_B_4VO5xxc52_2(.din(n30280), .dout(n30283));
    jdff dff_B_rsDZjJQp9_2(.din(n30283), .dout(n30286));
    jdff dff_B_Xx1zgopg7_2(.din(n30286), .dout(n30289));
    jdff dff_B_UJiMHZ1T7_2(.din(n30289), .dout(n30292));
    jdff dff_B_CqfMuxuq4_2(.din(n30292), .dout(n30295));
    jdff dff_B_fQriyvUs6_2(.din(n30295), .dout(n30298));
    jdff dff_B_rbfuiNGA4_2(.din(n30298), .dout(n30301));
    jdff dff_B_0L2gbH7y8_2(.din(n30301), .dout(n30304));
    jdff dff_B_IQenXnjK5_2(.din(n30304), .dout(n30307));
    jdff dff_B_gVBE3rh19_2(.din(n30307), .dout(n30310));
    jdff dff_B_DyB1IKPC5_2(.din(n30310), .dout(n30313));
    jdff dff_B_qT5sAETC5_1(.din(n6485), .dout(n30316));
    jdff dff_B_ITq5ODvv5_1(.din(n30316), .dout(n30319));
    jdff dff_B_sqPDmQhi6_2(.din(n6481), .dout(n30322));
    jdff dff_B_XHC47qVA8_2(.din(n30322), .dout(n30325));
    jdff dff_B_Lcsrw7ZW2_2(.din(n30325), .dout(n30328));
    jdff dff_B_AghjpGzh2_2(.din(n30328), .dout(n30331));
    jdff dff_B_AsT0YJje5_2(.din(n30331), .dout(n30334));
    jdff dff_B_jMrePLeH8_2(.din(n30334), .dout(n30337));
    jdff dff_B_Ra7XznvX7_2(.din(n30337), .dout(n30340));
    jdff dff_B_sPrRGCIl5_2(.din(n30340), .dout(n30343));
    jdff dff_B_9m5DIBku3_2(.din(n30343), .dout(n30346));
    jdff dff_B_wd47nu722_2(.din(n30346), .dout(n30349));
    jdff dff_B_kOheLc7A8_2(.din(n30349), .dout(n30352));
    jdff dff_B_UBxZJgp13_2(.din(n30352), .dout(n30355));
    jdff dff_B_W3z5arOG0_2(.din(n30355), .dout(n30358));
    jdff dff_B_nEPJvcAE5_2(.din(n30358), .dout(n30361));
    jdff dff_B_e9AZpvSL1_2(.din(n30361), .dout(n30364));
    jdff dff_B_34hCClRC5_2(.din(n30364), .dout(n30367));
    jdff dff_B_QtxlQDeo3_2(.din(n30367), .dout(n30370));
    jdff dff_B_A5G1GQsU1_2(.din(n30370), .dout(n30373));
    jdff dff_B_Z6WgYcih9_2(.din(n30373), .dout(n30376));
    jdff dff_B_Un0gvM0A3_2(.din(n30376), .dout(n30379));
    jdff dff_B_cEG43IBd2_2(.din(n30379), .dout(n30382));
    jdff dff_B_UmiKB51T9_2(.din(n30382), .dout(n30385));
    jdff dff_B_vmejwXTn7_2(.din(n30385), .dout(n30388));
    jdff dff_B_fBUGWA7r4_2(.din(n30388), .dout(n30391));
    jdff dff_B_RybLmypm7_2(.din(n30391), .dout(n30394));
    jdff dff_B_TrRCfxIc6_2(.din(n30394), .dout(n30397));
    jdff dff_B_NudGuLI28_2(.din(n30397), .dout(n30400));
    jdff dff_B_Udft1zug1_2(.din(n30400), .dout(n30403));
    jdff dff_B_bndFKDjV2_2(.din(n30403), .dout(n30406));
    jdff dff_B_tRLHHMq32_2(.din(n30406), .dout(n30409));
    jdff dff_B_6oO5qoZ88_2(.din(n30409), .dout(n30412));
    jdff dff_B_PPkq81yt1_2(.din(n30412), .dout(n30415));
    jdff dff_B_Up27UF968_2(.din(n30415), .dout(n30418));
    jdff dff_B_h8i0gn0l5_2(.din(n30418), .dout(n30421));
    jdff dff_B_pa97XfOY7_2(.din(n30421), .dout(n30424));
    jdff dff_B_9G0AjUt00_2(.din(n30424), .dout(n30427));
    jdff dff_B_hDkgm3b39_2(.din(n30427), .dout(n30430));
    jdff dff_B_gRhSfi7Y4_2(.din(n30430), .dout(n30433));
    jdff dff_B_kFbdzq0O6_2(.din(n30433), .dout(n30436));
    jdff dff_B_Vk0OT2gT7_2(.din(n30436), .dout(n30439));
    jdff dff_B_0NfvmgbE2_2(.din(n30439), .dout(n30442));
    jdff dff_B_IQFjwthz5_2(.din(n30442), .dout(n30445));
    jdff dff_B_MgjlpJUQ4_2(.din(n30445), .dout(n30448));
    jdff dff_B_XccXmWny7_2(.din(n30448), .dout(n30451));
    jdff dff_B_bIda4Wl94_2(.din(n6477), .dout(n30454));
    jdff dff_B_D2cKQdCD6_2(.din(n30454), .dout(n30457));
    jdff dff_B_WOviowce3_2(.din(n30457), .dout(n30460));
    jdff dff_B_RtvW9lIH1_2(.din(n30460), .dout(n30463));
    jdff dff_B_ngoc9Dr45_2(.din(n30463), .dout(n30466));
    jdff dff_B_yM6Mq15k2_2(.din(n30466), .dout(n30469));
    jdff dff_B_YYC0TVfN6_2(.din(n30469), .dout(n30472));
    jdff dff_B_LcvQ6Vel9_2(.din(n30472), .dout(n30475));
    jdff dff_B_Gj7zbwEj5_2(.din(n30475), .dout(n30478));
    jdff dff_B_NIhRWEWa3_2(.din(n30478), .dout(n30481));
    jdff dff_B_6RhbpRHq5_2(.din(n30481), .dout(n30484));
    jdff dff_B_xrjWXvYI5_2(.din(n30484), .dout(n30487));
    jdff dff_B_nOwczB7i9_2(.din(n30487), .dout(n30490));
    jdff dff_B_sw9dZln41_2(.din(n30490), .dout(n30493));
    jdff dff_B_zBpaf05x4_2(.din(n30493), .dout(n30496));
    jdff dff_B_HPBngvMO2_2(.din(n30496), .dout(n30499));
    jdff dff_B_V2xOTHGb5_2(.din(n30499), .dout(n30502));
    jdff dff_B_M9SZ4K9n7_2(.din(n30502), .dout(n30505));
    jdff dff_B_BVMznqHk9_2(.din(n30505), .dout(n30508));
    jdff dff_B_c1B8b2oY8_2(.din(n30508), .dout(n30511));
    jdff dff_B_idg30Hq10_2(.din(n30511), .dout(n30514));
    jdff dff_B_2RjKTG4C6_2(.din(n30514), .dout(n30517));
    jdff dff_B_ro5LUE5u7_2(.din(n30517), .dout(n30520));
    jdff dff_B_COgsj6Jh5_2(.din(n30520), .dout(n30523));
    jdff dff_B_IyAuwlPp5_2(.din(n30523), .dout(n30526));
    jdff dff_B_Iz5CJ1uM3_2(.din(n30526), .dout(n30529));
    jdff dff_B_HlG3ISFt2_2(.din(n30529), .dout(n30532));
    jdff dff_B_Rd4TqUI25_2(.din(n30532), .dout(n30535));
    jdff dff_B_cDI7qBXs5_2(.din(n30535), .dout(n30538));
    jdff dff_B_EqfTcMKK7_2(.din(n30538), .dout(n30541));
    jdff dff_B_dCEUnK2t6_2(.din(n30541), .dout(n30544));
    jdff dff_B_8Lpohban6_2(.din(n30544), .dout(n30547));
    jdff dff_B_3mIoPgG90_2(.din(n30547), .dout(n30550));
    jdff dff_B_0gNR8ukV1_2(.din(n30550), .dout(n30553));
    jdff dff_B_ZOUbpQuz2_2(.din(n30553), .dout(n30556));
    jdff dff_B_zi9iEQlJ1_2(.din(n30556), .dout(n30559));
    jdff dff_B_P4LaNWa51_2(.din(n30559), .dout(n30562));
    jdff dff_B_KWCFnulf0_2(.din(n30562), .dout(n30565));
    jdff dff_B_FqOHMpem9_2(.din(n30565), .dout(n30568));
    jdff dff_B_2Xg4DstL1_2(.din(n30568), .dout(n30571));
    jdff dff_B_1B3fioXq4_2(.din(n30571), .dout(n30574));
    jdff dff_B_SlOPBWUG4_2(.din(n30574), .dout(n30577));
    jdff dff_B_ZlrO80Xt4_2(.din(n30577), .dout(n30580));
    jdff dff_B_o2rqvsZX4_2(.din(n30580), .dout(n30583));
    jdff dff_B_DAygf4x11_2(.din(n30583), .dout(n30586));
    jdff dff_B_B7RNIbNT7_2(.din(n30586), .dout(n30589));
    jdff dff_B_0wdXCfdC9_2(.din(n6473), .dout(n30592));
    jdff dff_B_UFVwRiwo2_1(.din(n6465), .dout(n30595));
    jdff dff_B_4CbQx41F9_2(.din(n6303), .dout(n30598));
    jdff dff_B_tOzd0Gtu8_2(.din(n30598), .dout(n30601));
    jdff dff_B_3RK9jRb23_2(.din(n30601), .dout(n30604));
    jdff dff_B_aHLVSmPo4_2(.din(n30604), .dout(n30607));
    jdff dff_B_njx5V7RV3_2(.din(n30607), .dout(n30610));
    jdff dff_B_AWLuKZf47_2(.din(n30610), .dout(n30613));
    jdff dff_B_8yo0YQbD7_2(.din(n30613), .dout(n30616));
    jdff dff_B_R1JKiXfl3_2(.din(n30616), .dout(n30619));
    jdff dff_B_hPiNVPYx9_2(.din(n30619), .dout(n30622));
    jdff dff_B_xRtlWB7b4_2(.din(n30622), .dout(n30625));
    jdff dff_B_7g4ARltO2_2(.din(n30625), .dout(n30628));
    jdff dff_B_cl3vqZW91_2(.din(n30628), .dout(n30631));
    jdff dff_B_aifoDLxY3_2(.din(n30631), .dout(n30634));
    jdff dff_B_WZ7VcjL10_2(.din(n30634), .dout(n30637));
    jdff dff_B_6HbPTyBX3_2(.din(n30637), .dout(n30640));
    jdff dff_B_UlcXload6_2(.din(n30640), .dout(n30643));
    jdff dff_B_DWbaprGE6_2(.din(n30643), .dout(n30646));
    jdff dff_B_0v5qJSuu3_2(.din(n30646), .dout(n30649));
    jdff dff_B_rt0SGGiy8_2(.din(n30649), .dout(n30652));
    jdff dff_B_uYwP1HhH2_2(.din(n30652), .dout(n30655));
    jdff dff_B_8Gn5FTjb7_2(.din(n30655), .dout(n30658));
    jdff dff_B_thXTg66f1_2(.din(n30658), .dout(n30661));
    jdff dff_B_1C367qgX9_2(.din(n30661), .dout(n30664));
    jdff dff_B_d8ORhABr8_2(.din(n30664), .dout(n30667));
    jdff dff_B_5ixPI9vT5_2(.din(n30667), .dout(n30670));
    jdff dff_B_s2XpSyNf3_2(.din(n30670), .dout(n30673));
    jdff dff_B_FPkc7MQy5_2(.din(n30673), .dout(n30676));
    jdff dff_B_Lfo6DpxF6_2(.din(n30676), .dout(n30679));
    jdff dff_B_dgD72bWa6_2(.din(n30679), .dout(n30682));
    jdff dff_B_BY1kU5Ct4_2(.din(n30682), .dout(n30685));
    jdff dff_B_eFP3B0QO9_2(.din(n30685), .dout(n30688));
    jdff dff_B_HJR4GMn03_2(.din(n30688), .dout(n30691));
    jdff dff_B_pV2aBFeC8_2(.din(n30691), .dout(n30694));
    jdff dff_B_UM4RUzm44_2(.din(n30694), .dout(n30697));
    jdff dff_B_zr5HyVi01_2(.din(n30697), .dout(n30700));
    jdff dff_B_z2ACCUCN5_2(.din(n30700), .dout(n30703));
    jdff dff_B_szGS4o266_2(.din(n30703), .dout(n30706));
    jdff dff_B_gLEu3eWy3_2(.din(n30706), .dout(n30709));
    jdff dff_B_BMMSSA753_2(.din(n30709), .dout(n30712));
    jdff dff_B_BBLcp6S29_2(.din(n30712), .dout(n30715));
    jdff dff_B_9MIUmrvb4_2(.din(n30715), .dout(n30718));
    jdff dff_B_WvOsFQZ35_2(.din(n30718), .dout(n30721));
    jdff dff_B_YpBZ67h04_2(.din(n30721), .dout(n30724));
    jdff dff_B_YXZvJO2k0_1(.din(n6327), .dout(n30727));
    jdff dff_B_sl9LlNAT0_1(.din(n30727), .dout(n30730));
    jdff dff_B_a60FCBK10_2(.din(n6323), .dout(n30733));
    jdff dff_B_s1t0Ne6l1_2(.din(n30733), .dout(n30736));
    jdff dff_B_8txMS7B40_2(.din(n30736), .dout(n30739));
    jdff dff_B_DX4hwEel0_2(.din(n30739), .dout(n30742));
    jdff dff_B_UALV2Nvv2_2(.din(n30742), .dout(n30745));
    jdff dff_B_rbZtHZzC4_2(.din(n30745), .dout(n30748));
    jdff dff_B_Mckbp9AA5_2(.din(n30748), .dout(n30751));
    jdff dff_B_LqIoFn6Q8_2(.din(n30751), .dout(n30754));
    jdff dff_B_f3VAqxAh7_2(.din(n30754), .dout(n30757));
    jdff dff_B_CnYgRNZE5_2(.din(n30757), .dout(n30760));
    jdff dff_B_pVWbBQ752_2(.din(n30760), .dout(n30763));
    jdff dff_B_lQkJtgS43_2(.din(n30763), .dout(n30766));
    jdff dff_B_OoVrgO5r5_2(.din(n30766), .dout(n30769));
    jdff dff_B_01azvw9k8_2(.din(n30769), .dout(n30772));
    jdff dff_B_vvHpNv2c6_2(.din(n30772), .dout(n30775));
    jdff dff_B_0Nxn7GMb3_2(.din(n30775), .dout(n30778));
    jdff dff_B_oJBPUXTm8_2(.din(n30778), .dout(n30781));
    jdff dff_B_jtkDR4jN2_2(.din(n30781), .dout(n30784));
    jdff dff_B_0QZrmuTs4_2(.din(n30784), .dout(n30787));
    jdff dff_B_4ONyxXPC6_2(.din(n30787), .dout(n30790));
    jdff dff_B_9DXOjNco4_2(.din(n30790), .dout(n30793));
    jdff dff_B_plsApLue3_2(.din(n30793), .dout(n30796));
    jdff dff_B_iZ8OwxC19_2(.din(n30796), .dout(n30799));
    jdff dff_B_P7ODU0VS2_2(.din(n30799), .dout(n30802));
    jdff dff_B_7XkJH0Kl6_2(.din(n30802), .dout(n30805));
    jdff dff_B_J2CyJSVW3_2(.din(n30805), .dout(n30808));
    jdff dff_B_awG32zrH7_2(.din(n30808), .dout(n30811));
    jdff dff_B_G4phLsEV1_2(.din(n30811), .dout(n30814));
    jdff dff_B_1sSPCddY0_2(.din(n30814), .dout(n30817));
    jdff dff_B_1KItqeoN9_2(.din(n30817), .dout(n30820));
    jdff dff_B_bjkQGqVN7_2(.din(n30820), .dout(n30823));
    jdff dff_B_GnKywHke3_2(.din(n30823), .dout(n30826));
    jdff dff_B_hcg06UVb7_2(.din(n30826), .dout(n30829));
    jdff dff_B_KMgVGQSX8_2(.din(n30829), .dout(n30832));
    jdff dff_B_m8TLvjHr8_2(.din(n30832), .dout(n30835));
    jdff dff_B_lBGh094G6_2(.din(n30835), .dout(n30838));
    jdff dff_B_A9W44fyG5_2(.din(n30838), .dout(n30841));
    jdff dff_B_ITUO9W679_2(.din(n30841), .dout(n30844));
    jdff dff_B_jubSsqcg2_2(.din(n30844), .dout(n30847));
    jdff dff_B_ftAC1Tv30_2(.din(n30847), .dout(n30850));
    jdff dff_B_lQcMoh2d5_2(.din(n6319), .dout(n30853));
    jdff dff_B_RzhjSOY79_2(.din(n30853), .dout(n30856));
    jdff dff_B_IVtF71gj1_2(.din(n30856), .dout(n30859));
    jdff dff_B_ne5l9KOw5_2(.din(n30859), .dout(n30862));
    jdff dff_B_LZv7m9H48_2(.din(n30862), .dout(n30865));
    jdff dff_B_xLPZGdPs7_2(.din(n30865), .dout(n30868));
    jdff dff_B_WpcYmYiE8_2(.din(n30868), .dout(n30871));
    jdff dff_B_Xe29gkP29_2(.din(n30871), .dout(n30874));
    jdff dff_B_X8q39fkN9_2(.din(n30874), .dout(n30877));
    jdff dff_B_qEs4RS6u6_2(.din(n30877), .dout(n30880));
    jdff dff_B_wu1PItlE7_2(.din(n30880), .dout(n30883));
    jdff dff_B_b7iuyeou2_2(.din(n30883), .dout(n30886));
    jdff dff_B_VMXC3PbE2_2(.din(n30886), .dout(n30889));
    jdff dff_B_mHuU6GOr7_2(.din(n30889), .dout(n30892));
    jdff dff_B_7fl2GvwK8_2(.din(n30892), .dout(n30895));
    jdff dff_B_4YiJLsiw6_2(.din(n30895), .dout(n30898));
    jdff dff_B_eP5FJVGW1_2(.din(n30898), .dout(n30901));
    jdff dff_B_d4gPjic42_2(.din(n30901), .dout(n30904));
    jdff dff_B_JOLA9J4w9_2(.din(n30904), .dout(n30907));
    jdff dff_B_c2lYvNJ78_2(.din(n30907), .dout(n30910));
    jdff dff_B_hODBv9zx5_2(.din(n30910), .dout(n30913));
    jdff dff_B_zNY6mDat2_2(.din(n30913), .dout(n30916));
    jdff dff_B_x8AeANCb1_2(.din(n30916), .dout(n30919));
    jdff dff_B_gqMnlbSj4_2(.din(n30919), .dout(n30922));
    jdff dff_B_QR4AWM4t6_2(.din(n30922), .dout(n30925));
    jdff dff_B_eoTPu0120_2(.din(n30925), .dout(n30928));
    jdff dff_B_KRrr06ro0_2(.din(n30928), .dout(n30931));
    jdff dff_B_yPDbsUSp2_2(.din(n30931), .dout(n30934));
    jdff dff_B_4D4VzV5M7_2(.din(n30934), .dout(n30937));
    jdff dff_B_iAMWRmag3_2(.din(n30937), .dout(n30940));
    jdff dff_B_i7GRGFgO4_2(.din(n30940), .dout(n30943));
    jdff dff_B_QEukstIO4_2(.din(n30943), .dout(n30946));
    jdff dff_B_Q5QgZt8i7_2(.din(n30946), .dout(n30949));
    jdff dff_B_89Bz2bgh5_2(.din(n30949), .dout(n30952));
    jdff dff_B_X7fyyJgm1_2(.din(n30952), .dout(n30955));
    jdff dff_B_pvEecekj9_2(.din(n30955), .dout(n30958));
    jdff dff_B_epgzQZn99_2(.din(n30958), .dout(n30961));
    jdff dff_B_WbEVTkPs8_2(.din(n30961), .dout(n30964));
    jdff dff_B_QDa8gHla1_2(.din(n30964), .dout(n30967));
    jdff dff_B_mEwxybiH7_2(.din(n30967), .dout(n30970));
    jdff dff_B_7lJ4oeRx8_2(.din(n30970), .dout(n30973));
    jdff dff_B_kv4gH2Zd2_2(.din(n30973), .dout(n30976));
    jdff dff_B_hrir7I2z8_2(.din(n6315), .dout(n30979));
    jdff dff_B_LD9XSOiS3_1(.din(n6307), .dout(n30982));
    jdff dff_B_IO8osC6D0_2(.din(n6109), .dout(n30985));
    jdff dff_B_5YZ5C6Kq6_2(.din(n30985), .dout(n30988));
    jdff dff_B_mt6k1Qos2_2(.din(n30988), .dout(n30991));
    jdff dff_B_jtmtyrZ36_2(.din(n30991), .dout(n30994));
    jdff dff_B_M5YPqomP5_2(.din(n30994), .dout(n30997));
    jdff dff_B_HgGLTEMa7_2(.din(n30997), .dout(n31000));
    jdff dff_B_2QcuSjtX7_2(.din(n31000), .dout(n31003));
    jdff dff_B_wmwHp6Js4_2(.din(n31003), .dout(n31006));
    jdff dff_B_zzYyRr8p3_2(.din(n31006), .dout(n31009));
    jdff dff_B_VO1JxMWh7_2(.din(n31009), .dout(n31012));
    jdff dff_B_AqsmNwUX4_2(.din(n31012), .dout(n31015));
    jdff dff_B_B9KIpRH98_2(.din(n31015), .dout(n31018));
    jdff dff_B_V2zO15AL1_2(.din(n31018), .dout(n31021));
    jdff dff_B_WGas6kLb8_2(.din(n31021), .dout(n31024));
    jdff dff_B_dxtI1b3L5_2(.din(n31024), .dout(n31027));
    jdff dff_B_BNkXoz4z2_2(.din(n31027), .dout(n31030));
    jdff dff_B_p6AAIeBf7_2(.din(n31030), .dout(n31033));
    jdff dff_B_loF9KRgF4_2(.din(n31033), .dout(n31036));
    jdff dff_B_55OKPuuj6_2(.din(n31036), .dout(n31039));
    jdff dff_B_D5tdWEfJ1_2(.din(n31039), .dout(n31042));
    jdff dff_B_uT3CuPGq1_2(.din(n31042), .dout(n31045));
    jdff dff_B_2YkQPLcm9_2(.din(n31045), .dout(n31048));
    jdff dff_B_7Ie72Y0Y4_2(.din(n31048), .dout(n31051));
    jdff dff_B_LQYwPaLL0_2(.din(n31051), .dout(n31054));
    jdff dff_B_LuE6FoXo9_2(.din(n31054), .dout(n31057));
    jdff dff_B_VeGAicis8_2(.din(n31057), .dout(n31060));
    jdff dff_B_OAZR1hcB0_2(.din(n31060), .dout(n31063));
    jdff dff_B_z6tL5lTR1_2(.din(n31063), .dout(n31066));
    jdff dff_B_3SOP35U57_2(.din(n31066), .dout(n31069));
    jdff dff_B_4ldaTvvg9_2(.din(n31069), .dout(n31072));
    jdff dff_B_E4V7pNm14_2(.din(n31072), .dout(n31075));
    jdff dff_B_GjkRbhM33_2(.din(n31075), .dout(n31078));
    jdff dff_B_8RUqxONn7_2(.din(n31078), .dout(n31081));
    jdff dff_B_rjemjsH95_2(.din(n31081), .dout(n31084));
    jdff dff_B_pXfP7u089_2(.din(n31084), .dout(n31087));
    jdff dff_B_6fugebGy4_2(.din(n31087), .dout(n31090));
    jdff dff_B_SuRv9RT48_2(.din(n31090), .dout(n31093));
    jdff dff_B_grxZZwjR0_2(.din(n31093), .dout(n31096));
    jdff dff_B_FH7jW32D5_2(.din(n31096), .dout(n31099));
    jdff dff_B_11h2mnBb6_1(.din(n6133), .dout(n31102));
    jdff dff_B_QnrhvDJ39_1(.din(n31102), .dout(n31105));
    jdff dff_B_OjtRWkz85_2(.din(n6129), .dout(n31108));
    jdff dff_B_H4sLWXAM1_2(.din(n31108), .dout(n31111));
    jdff dff_B_rhKgKYmg2_2(.din(n31111), .dout(n31114));
    jdff dff_B_PrcewLJg3_2(.din(n31114), .dout(n31117));
    jdff dff_B_ciMQANda1_2(.din(n31117), .dout(n31120));
    jdff dff_B_BsoIaXf27_2(.din(n31120), .dout(n31123));
    jdff dff_B_oQWgyVv40_2(.din(n31123), .dout(n31126));
    jdff dff_B_yB01E5nB4_2(.din(n31126), .dout(n31129));
    jdff dff_B_7FeFVmGh3_2(.din(n31129), .dout(n31132));
    jdff dff_B_Tmxh3YeH3_2(.din(n31132), .dout(n31135));
    jdff dff_B_yCsTGjWz8_2(.din(n31135), .dout(n31138));
    jdff dff_B_y9zwp4Az5_2(.din(n31138), .dout(n31141));
    jdff dff_B_YFiH6sbf2_2(.din(n31141), .dout(n31144));
    jdff dff_B_FnzaljUV9_2(.din(n31144), .dout(n31147));
    jdff dff_B_ix1L4zjC8_2(.din(n31147), .dout(n31150));
    jdff dff_B_VVQpPhB32_2(.din(n31150), .dout(n31153));
    jdff dff_B_sSgwnOrU2_2(.din(n31153), .dout(n31156));
    jdff dff_B_UJZ3Wht43_2(.din(n31156), .dout(n31159));
    jdff dff_B_S6OOM1Kq2_2(.din(n31159), .dout(n31162));
    jdff dff_B_dBV8XEuL1_2(.din(n31162), .dout(n31165));
    jdff dff_B_sxWOfH029_2(.din(n31165), .dout(n31168));
    jdff dff_B_uwtfZuaL3_2(.din(n31168), .dout(n31171));
    jdff dff_B_PRHyGlfj1_2(.din(n31171), .dout(n31174));
    jdff dff_B_NwBrKywE1_2(.din(n31174), .dout(n31177));
    jdff dff_B_mI0wTFno9_2(.din(n31177), .dout(n31180));
    jdff dff_B_hX6AAV445_2(.din(n31180), .dout(n31183));
    jdff dff_B_5CvxOZxv5_2(.din(n31183), .dout(n31186));
    jdff dff_B_7c00OjEb2_2(.din(n31186), .dout(n31189));
    jdff dff_B_MbRKR5KN5_2(.din(n31189), .dout(n31192));
    jdff dff_B_BkYHmE6V4_2(.din(n31192), .dout(n31195));
    jdff dff_B_YE2rx8cE6_2(.din(n31195), .dout(n31198));
    jdff dff_B_Q2Bm8MuR8_2(.din(n31198), .dout(n31201));
    jdff dff_B_5MqNYOMH4_2(.din(n31201), .dout(n31204));
    jdff dff_B_lnxo9GcD3_2(.din(n31204), .dout(n31207));
    jdff dff_B_dOovRSgX9_2(.din(n31207), .dout(n31210));
    jdff dff_B_gllUR0MF3_2(.din(n31210), .dout(n31213));
    jdff dff_B_XnR8pnxw7_2(.din(n6125), .dout(n31216));
    jdff dff_B_GR15E4pp6_2(.din(n31216), .dout(n31219));
    jdff dff_B_PCIhFuYQ6_2(.din(n31219), .dout(n31222));
    jdff dff_B_IKYZ6lqQ6_2(.din(n31222), .dout(n31225));
    jdff dff_B_E65ue60G1_2(.din(n31225), .dout(n31228));
    jdff dff_B_CuRHdUgE3_2(.din(n31228), .dout(n31231));
    jdff dff_B_vf1kuXxr8_2(.din(n31231), .dout(n31234));
    jdff dff_B_jnb87pNR1_2(.din(n31234), .dout(n31237));
    jdff dff_B_8X9VvcrN1_2(.din(n31237), .dout(n31240));
    jdff dff_B_nrCLN1p26_2(.din(n31240), .dout(n31243));
    jdff dff_B_yog6ln8E5_2(.din(n31243), .dout(n31246));
    jdff dff_B_pEmW8hLs0_2(.din(n31246), .dout(n31249));
    jdff dff_B_TkCdXKA67_2(.din(n31249), .dout(n31252));
    jdff dff_B_FW6cNoW11_2(.din(n31252), .dout(n31255));
    jdff dff_B_ehuOBwyZ0_2(.din(n31255), .dout(n31258));
    jdff dff_B_0ZrObZ2m1_2(.din(n31258), .dout(n31261));
    jdff dff_B_Eq7tGFbb8_2(.din(n31261), .dout(n31264));
    jdff dff_B_10mGnbdy4_2(.din(n31264), .dout(n31267));
    jdff dff_B_cJiyqwCu8_2(.din(n31267), .dout(n31270));
    jdff dff_B_CVoOe6WP7_2(.din(n31270), .dout(n31273));
    jdff dff_B_868FyOFP4_2(.din(n31273), .dout(n31276));
    jdff dff_B_Q08SRK5p4_2(.din(n31276), .dout(n31279));
    jdff dff_B_alGe5RtK7_2(.din(n31279), .dout(n31282));
    jdff dff_B_Zp6xdwHW2_2(.din(n31282), .dout(n31285));
    jdff dff_B_I8DUJgua2_2(.din(n31285), .dout(n31288));
    jdff dff_B_31Sj8Rt25_2(.din(n31288), .dout(n31291));
    jdff dff_B_JV0yl0MZ1_2(.din(n31291), .dout(n31294));
    jdff dff_B_j9x3Q7nm3_2(.din(n31294), .dout(n31297));
    jdff dff_B_GnXLaZHG8_2(.din(n31297), .dout(n31300));
    jdff dff_B_Z3pLEOEH0_2(.din(n31300), .dout(n31303));
    jdff dff_B_HbzwnA556_2(.din(n31303), .dout(n31306));
    jdff dff_B_dv1s7Ykx1_2(.din(n31306), .dout(n31309));
    jdff dff_B_ObRThRGk1_2(.din(n31309), .dout(n31312));
    jdff dff_B_XwJ5JWuj3_2(.din(n31312), .dout(n31315));
    jdff dff_B_2q4SW0fe1_2(.din(n31315), .dout(n31318));
    jdff dff_B_ocKxbxSA6_2(.din(n31318), .dout(n31321));
    jdff dff_B_9PAd5v7J8_2(.din(n31321), .dout(n31324));
    jdff dff_B_NufzxXYp2_2(.din(n31324), .dout(n31327));
    jdff dff_B_IGBSwx534_2(.din(n6121), .dout(n31330));
    jdff dff_B_PRIZboWh1_1(.din(n6113), .dout(n31333));
    jdff dff_B_NracL9LR4_2(.din(n5891), .dout(n31336));
    jdff dff_B_0NUeyTxa8_2(.din(n31336), .dout(n31339));
    jdff dff_B_zRK2UE0c0_2(.din(n31339), .dout(n31342));
    jdff dff_B_FN3IRPQl4_2(.din(n31342), .dout(n31345));
    jdff dff_B_jAv1NIka7_2(.din(n31345), .dout(n31348));
    jdff dff_B_teeeHzWr1_2(.din(n31348), .dout(n31351));
    jdff dff_B_6fvY58Yc2_2(.din(n31351), .dout(n31354));
    jdff dff_B_Qwudmptu0_2(.din(n31354), .dout(n31357));
    jdff dff_B_MCD9BKO21_2(.din(n31357), .dout(n31360));
    jdff dff_B_dgyQrOCl3_2(.din(n31360), .dout(n31363));
    jdff dff_B_caS2ihKx8_2(.din(n31363), .dout(n31366));
    jdff dff_B_sERGt8je2_2(.din(n31366), .dout(n31369));
    jdff dff_B_wse96MkP4_2(.din(n31369), .dout(n31372));
    jdff dff_B_YVoBk29T8_2(.din(n31372), .dout(n31375));
    jdff dff_B_rNnEPmTd7_2(.din(n31375), .dout(n31378));
    jdff dff_B_91DkQBZA9_2(.din(n31378), .dout(n31381));
    jdff dff_B_WzkmCQyW8_2(.din(n31381), .dout(n31384));
    jdff dff_B_2Mjyl81S8_2(.din(n31384), .dout(n31387));
    jdff dff_B_RQRhDMSc3_2(.din(n31387), .dout(n31390));
    jdff dff_B_xLWUme7f7_2(.din(n31390), .dout(n31393));
    jdff dff_B_M4pE5sV05_2(.din(n31393), .dout(n31396));
    jdff dff_B_FiRVVw5h1_2(.din(n31396), .dout(n31399));
    jdff dff_B_4mzbmJPp6_2(.din(n31399), .dout(n31402));
    jdff dff_B_AOlAwuXk7_2(.din(n31402), .dout(n31405));
    jdff dff_B_BTHarfsS1_2(.din(n31405), .dout(n31408));
    jdff dff_B_4UvEFnxN4_2(.din(n31408), .dout(n31411));
    jdff dff_B_TbSFipsC5_2(.din(n31411), .dout(n31414));
    jdff dff_B_qCxYuplw6_2(.din(n31414), .dout(n31417));
    jdff dff_B_02PCvWrG3_2(.din(n31417), .dout(n31420));
    jdff dff_B_TwB6wEks6_2(.din(n31420), .dout(n31423));
    jdff dff_B_FDz5upXD3_2(.din(n31423), .dout(n31426));
    jdff dff_B_SiabVybH4_2(.din(n31426), .dout(n31429));
    jdff dff_B_VraM9NXu3_2(.din(n31429), .dout(n31432));
    jdff dff_B_qJzGZ17T5_2(.din(n31432), .dout(n31435));
    jdff dff_B_poyiy4tx3_2(.din(n31435), .dout(n31438));
    jdff dff_B_o269yUIt0_1(.din(n5915), .dout(n31441));
    jdff dff_B_F8seNExg6_1(.din(n31441), .dout(n31444));
    jdff dff_B_CKhLp4CL1_2(.din(n5911), .dout(n31447));
    jdff dff_B_xRDHZbVN6_2(.din(n31447), .dout(n31450));
    jdff dff_B_oqi26wSG4_2(.din(n31450), .dout(n31453));
    jdff dff_B_9tYi3ZoF6_2(.din(n31453), .dout(n31456));
    jdff dff_B_wZVMEj6s0_2(.din(n31456), .dout(n31459));
    jdff dff_B_tJibNlXw0_2(.din(n31459), .dout(n31462));
    jdff dff_B_JbuW4FVZ4_2(.din(n31462), .dout(n31465));
    jdff dff_B_JMyUr2pa2_2(.din(n31465), .dout(n31468));
    jdff dff_B_spw74YZt9_2(.din(n31468), .dout(n31471));
    jdff dff_B_68BhCiDL5_2(.din(n31471), .dout(n31474));
    jdff dff_B_9pAHtDJY3_2(.din(n31474), .dout(n31477));
    jdff dff_B_tD8IOVpw4_2(.din(n31477), .dout(n31480));
    jdff dff_B_lFHHKp1E1_2(.din(n31480), .dout(n31483));
    jdff dff_B_sYNlZP2V8_2(.din(n31483), .dout(n31486));
    jdff dff_B_6fJPR5jL1_2(.din(n31486), .dout(n31489));
    jdff dff_B_Z1351Jwl1_2(.din(n31489), .dout(n31492));
    jdff dff_B_NAhqd4hB7_2(.din(n31492), .dout(n31495));
    jdff dff_B_uftwVYDF0_2(.din(n31495), .dout(n31498));
    jdff dff_B_YTM6FdhP4_2(.din(n31498), .dout(n31501));
    jdff dff_B_XT5l0IX35_2(.din(n31501), .dout(n31504));
    jdff dff_B_gfi2GPms9_2(.din(n31504), .dout(n31507));
    jdff dff_B_7LGXwjJU3_2(.din(n31507), .dout(n31510));
    jdff dff_B_9Bl4KFyY8_2(.din(n31510), .dout(n31513));
    jdff dff_B_P7fVqXY20_2(.din(n31513), .dout(n31516));
    jdff dff_B_bcNGexlG7_2(.din(n31516), .dout(n31519));
    jdff dff_B_qkyEtRzg8_2(.din(n31519), .dout(n31522));
    jdff dff_B_5zXY9Bby4_2(.din(n31522), .dout(n31525));
    jdff dff_B_I9nvUdiI9_2(.din(n31525), .dout(n31528));
    jdff dff_B_Wzt3jgkN5_2(.din(n31528), .dout(n31531));
    jdff dff_B_qa9CpgJ81_2(.din(n31531), .dout(n31534));
    jdff dff_B_4MP7TjJv7_2(.din(n31534), .dout(n31537));
    jdff dff_B_k33KKcJH0_2(.din(n31537), .dout(n31540));
    jdff dff_B_z5sIHDtl4_2(.din(n5907), .dout(n31543));
    jdff dff_B_ceOKQeDm3_2(.din(n31543), .dout(n31546));
    jdff dff_B_OIwOBmQ74_2(.din(n31546), .dout(n31549));
    jdff dff_B_3VDPHyRE7_2(.din(n31549), .dout(n31552));
    jdff dff_B_45xF50ic2_2(.din(n31552), .dout(n31555));
    jdff dff_B_OkN2jMdi2_2(.din(n31555), .dout(n31558));
    jdff dff_B_oH16Peh98_2(.din(n31558), .dout(n31561));
    jdff dff_B_LR98fBSb3_2(.din(n31561), .dout(n31564));
    jdff dff_B_m2VBFUQB9_2(.din(n31564), .dout(n31567));
    jdff dff_B_ofV171bt6_2(.din(n31567), .dout(n31570));
    jdff dff_B_y2q5XDX69_2(.din(n31570), .dout(n31573));
    jdff dff_B_XP0fBp7V2_2(.din(n31573), .dout(n31576));
    jdff dff_B_W8vqF5TY8_2(.din(n31576), .dout(n31579));
    jdff dff_B_ieeJvNcR6_2(.din(n31579), .dout(n31582));
    jdff dff_B_qfeuUqiQ7_2(.din(n31582), .dout(n31585));
    jdff dff_B_rCIUZCPg8_2(.din(n31585), .dout(n31588));
    jdff dff_B_RJ14PlcM2_2(.din(n31588), .dout(n31591));
    jdff dff_B_3ZsxmYPr5_2(.din(n31591), .dout(n31594));
    jdff dff_B_M8SpTF1E4_2(.din(n31594), .dout(n31597));
    jdff dff_B_cXHeC0i30_2(.din(n31597), .dout(n31600));
    jdff dff_B_3pZV89Ul7_2(.din(n31600), .dout(n31603));
    jdff dff_B_vKJCAfLp4_2(.din(n31603), .dout(n31606));
    jdff dff_B_YlPJwVTa2_2(.din(n31606), .dout(n31609));
    jdff dff_B_Ag52ToH48_2(.din(n31609), .dout(n31612));
    jdff dff_B_In1xradN7_2(.din(n31612), .dout(n31615));
    jdff dff_B_Ssv5yBim0_2(.din(n31615), .dout(n31618));
    jdff dff_B_eW05ITvY5_2(.din(n31618), .dout(n31621));
    jdff dff_B_VOxdsDCI2_2(.din(n31621), .dout(n31624));
    jdff dff_B_u4nTYRW40_2(.din(n31624), .dout(n31627));
    jdff dff_B_3WN5ZGwT8_2(.din(n31627), .dout(n31630));
    jdff dff_B_qENnCH9B0_2(.din(n31630), .dout(n31633));
    jdff dff_B_KU1oYdmK9_2(.din(n31633), .dout(n31636));
    jdff dff_B_PCSE2ZYu5_2(.din(n31636), .dout(n31639));
    jdff dff_B_Dk0tMq5b9_2(.din(n31639), .dout(n31642));
    jdff dff_B_896xBcra0_2(.din(n5903), .dout(n31645));
    jdff dff_B_McwKnVtr5_1(.din(n5895), .dout(n31648));
    jdff dff_B_bZ6WEBNu7_2(.din(n5646), .dout(n31651));
    jdff dff_B_xzEVptqB3_2(.din(n31651), .dout(n31654));
    jdff dff_B_ea4bv41s1_2(.din(n31654), .dout(n31657));
    jdff dff_B_EEK7yyOR7_2(.din(n31657), .dout(n31660));
    jdff dff_B_G5rB0ymr7_2(.din(n31660), .dout(n31663));
    jdff dff_B_GLf2xhsH2_2(.din(n31663), .dout(n31666));
    jdff dff_B_dXmZjGWX2_2(.din(n31666), .dout(n31669));
    jdff dff_B_3muGzQyA3_2(.din(n31669), .dout(n31672));
    jdff dff_B_2FDjoapF1_2(.din(n31672), .dout(n31675));
    jdff dff_B_KEI8AuKV3_2(.din(n31675), .dout(n31678));
    jdff dff_B_VDBAvZfu0_2(.din(n31678), .dout(n31681));
    jdff dff_B_NgLvRoqM9_2(.din(n31681), .dout(n31684));
    jdff dff_B_2ab4lZzW5_2(.din(n31684), .dout(n31687));
    jdff dff_B_BrQETskv6_2(.din(n31687), .dout(n31690));
    jdff dff_B_7Y5AYlhf9_2(.din(n31690), .dout(n31693));
    jdff dff_B_ewG0hSRH3_2(.din(n31693), .dout(n31696));
    jdff dff_B_WPS5zvIH6_2(.din(n31696), .dout(n31699));
    jdff dff_B_CBfMUNlC8_2(.din(n31699), .dout(n31702));
    jdff dff_B_Q7SK2WP14_2(.din(n31702), .dout(n31705));
    jdff dff_B_9RdwN7NJ2_2(.din(n31705), .dout(n31708));
    jdff dff_B_utU1DPPF8_2(.din(n31708), .dout(n31711));
    jdff dff_B_dCgsYsmP2_2(.din(n31711), .dout(n31714));
    jdff dff_B_MD0JMfIu9_2(.din(n31714), .dout(n31717));
    jdff dff_B_gBZwyyzt0_2(.din(n31717), .dout(n31720));
    jdff dff_B_AhXiICfe0_2(.din(n31720), .dout(n31723));
    jdff dff_B_v8yKt9CW2_2(.din(n31723), .dout(n31726));
    jdff dff_B_lMxW56rO1_2(.din(n31726), .dout(n31729));
    jdff dff_B_M4PoGaBP3_2(.din(n31729), .dout(n31732));
    jdff dff_B_XT0Pvyyn6_2(.din(n31732), .dout(n31735));
    jdff dff_B_ZOu315Ty6_2(.din(n31735), .dout(n31738));
    jdff dff_B_ugBGSNfa3_2(.din(n31738), .dout(n31741));
    jdff dff_B_qoDRJVxL7_1(.din(n5670), .dout(n31744));
    jdff dff_B_2ezTw40N3_1(.din(n31744), .dout(n31747));
    jdff dff_B_58UfveQP3_2(.din(n5666), .dout(n31750));
    jdff dff_B_ADp3j63K0_2(.din(n31750), .dout(n31753));
    jdff dff_B_i7itV8O29_2(.din(n31753), .dout(n31756));
    jdff dff_B_UAApKXy27_2(.din(n31756), .dout(n31759));
    jdff dff_B_ualVowA88_2(.din(n31759), .dout(n31762));
    jdff dff_B_QcDY9brj0_2(.din(n31762), .dout(n31765));
    jdff dff_B_GdyBCVIk3_2(.din(n31765), .dout(n31768));
    jdff dff_B_TiogwJfi9_2(.din(n31768), .dout(n31771));
    jdff dff_B_gPw2qPn51_2(.din(n31771), .dout(n31774));
    jdff dff_B_3lSYcOmN9_2(.din(n31774), .dout(n31777));
    jdff dff_B_RqrDtsIH9_2(.din(n31777), .dout(n31780));
    jdff dff_B_nqltyu9W7_2(.din(n31780), .dout(n31783));
    jdff dff_B_Llt5KdTM8_2(.din(n31783), .dout(n31786));
    jdff dff_B_Cbi5UaaD9_2(.din(n31786), .dout(n31789));
    jdff dff_B_Y1QeJM9E6_2(.din(n31789), .dout(n31792));
    jdff dff_B_dPpWhZ6g2_2(.din(n31792), .dout(n31795));
    jdff dff_B_qwjEigGV2_2(.din(n31795), .dout(n31798));
    jdff dff_B_8rUETevF1_2(.din(n31798), .dout(n31801));
    jdff dff_B_igXJoIem2_2(.din(n31801), .dout(n31804));
    jdff dff_B_uZnQPvYp7_2(.din(n31804), .dout(n31807));
    jdff dff_B_y8rwqxq31_2(.din(n31807), .dout(n31810));
    jdff dff_B_FKTrVXhZ8_2(.din(n31810), .dout(n31813));
    jdff dff_B_3nv21eCL6_2(.din(n31813), .dout(n31816));
    jdff dff_B_F19CCd8T2_2(.din(n31816), .dout(n31819));
    jdff dff_B_kFLHSc7L3_2(.din(n31819), .dout(n31822));
    jdff dff_B_VeEQDDQO3_2(.din(n31822), .dout(n31825));
    jdff dff_B_vzwqLw0d9_2(.din(n31825), .dout(n31828));
    jdff dff_B_7nodYucn0_2(.din(n31828), .dout(n31831));
    jdff dff_B_60a6Xq1l9_2(.din(n5662), .dout(n31834));
    jdff dff_B_hodZAB5S2_2(.din(n31834), .dout(n31837));
    jdff dff_B_KXkbuGap5_2(.din(n31837), .dout(n31840));
    jdff dff_B_q24DgdNX2_2(.din(n31840), .dout(n31843));
    jdff dff_B_lI9Asubr5_2(.din(n31843), .dout(n31846));
    jdff dff_B_C9nG3yxR4_2(.din(n31846), .dout(n31849));
    jdff dff_B_YcRguUlg1_2(.din(n31849), .dout(n31852));
    jdff dff_B_3vZBWnPc9_2(.din(n31852), .dout(n31855));
    jdff dff_B_pbwmV0Pd3_2(.din(n31855), .dout(n31858));
    jdff dff_B_N8ZhIHqc4_2(.din(n31858), .dout(n31861));
    jdff dff_B_f70K9my72_2(.din(n31861), .dout(n31864));
    jdff dff_B_irg1wuLv2_2(.din(n31864), .dout(n31867));
    jdff dff_B_z4IAjJXj2_2(.din(n31867), .dout(n31870));
    jdff dff_B_cbLsPkEf9_2(.din(n31870), .dout(n31873));
    jdff dff_B_BRob48bd0_2(.din(n31873), .dout(n31876));
    jdff dff_B_9uiwO0Nl7_2(.din(n31876), .dout(n31879));
    jdff dff_B_SLiuM5ML4_2(.din(n31879), .dout(n31882));
    jdff dff_B_KYcwbfYM0_2(.din(n31882), .dout(n31885));
    jdff dff_B_zRRdla247_2(.din(n31885), .dout(n31888));
    jdff dff_B_VYh0AFar9_2(.din(n31888), .dout(n31891));
    jdff dff_B_BvHwI7er9_2(.din(n31891), .dout(n31894));
    jdff dff_B_SSqH70Pr3_2(.din(n31894), .dout(n31897));
    jdff dff_B_s0avIIv43_2(.din(n31897), .dout(n31900));
    jdff dff_B_e6Yqgxd20_2(.din(n31900), .dout(n31903));
    jdff dff_B_C41PjQDs7_2(.din(n31903), .dout(n31906));
    jdff dff_B_voCVrfKC1_2(.din(n31906), .dout(n31909));
    jdff dff_B_Kf2JBVjW1_2(.din(n31909), .dout(n31912));
    jdff dff_B_oFa4G7VG1_2(.din(n31912), .dout(n31915));
    jdff dff_B_3CPhrYIH7_2(.din(n31915), .dout(n31918));
    jdff dff_B_8YzArT0w9_2(.din(n31918), .dout(n31921));
    jdff dff_B_jyCedYn23_2(.din(n5658), .dout(n31924));
    jdff dff_B_4ZGyLYI34_1(.din(n5650), .dout(n31927));
    jdff dff_B_qFNYwrEz8_2(.din(n5374), .dout(n31930));
    jdff dff_B_aPMWol1E1_2(.din(n31930), .dout(n31933));
    jdff dff_B_YHzQ0G6b9_2(.din(n31933), .dout(n31936));
    jdff dff_B_7x82HizO4_2(.din(n31936), .dout(n31939));
    jdff dff_B_trzPZ1DV9_2(.din(n31939), .dout(n31942));
    jdff dff_B_iTpLJomj2_2(.din(n31942), .dout(n31945));
    jdff dff_B_Noac6bpN9_2(.din(n31945), .dout(n31948));
    jdff dff_B_ziRsvjyZ2_2(.din(n31948), .dout(n31951));
    jdff dff_B_tY7iefEe6_2(.din(n31951), .dout(n31954));
    jdff dff_B_sTQAvUcs4_2(.din(n31954), .dout(n31957));
    jdff dff_B_mXctcUt55_2(.din(n31957), .dout(n31960));
    jdff dff_B_29Y4etSI2_2(.din(n31960), .dout(n31963));
    jdff dff_B_WuFtF8pK6_2(.din(n31963), .dout(n31966));
    jdff dff_B_zO4t1JEV1_2(.din(n31966), .dout(n31969));
    jdff dff_B_Hb4tDzjv1_2(.din(n31969), .dout(n31972));
    jdff dff_B_mnmD1hQL7_2(.din(n31972), .dout(n31975));
    jdff dff_B_mMfPWLG28_2(.din(n31975), .dout(n31978));
    jdff dff_B_F3GEOyI63_2(.din(n31978), .dout(n31981));
    jdff dff_B_QeSoVTIQ9_2(.din(n31981), .dout(n31984));
    jdff dff_B_PXKRWx8c6_2(.din(n31984), .dout(n31987));
    jdff dff_B_ofihC0d07_2(.din(n31987), .dout(n31990));
    jdff dff_B_c656eRfT1_2(.din(n31990), .dout(n31993));
    jdff dff_B_lOISoo5H7_2(.din(n31993), .dout(n31996));
    jdff dff_B_rPZS3WR15_2(.din(n31996), .dout(n31999));
    jdff dff_B_t3HreJNU1_2(.din(n31999), .dout(n32002));
    jdff dff_B_gN63ag3Z0_2(.din(n32002), .dout(n32005));
    jdff dff_B_FDLZUWT77_2(.din(n32005), .dout(n32008));
    jdff dff_B_VA2S6U9k3_1(.din(n5398), .dout(n32011));
    jdff dff_B_RSFFa2ch4_1(.din(n32011), .dout(n32014));
    jdff dff_B_qYTGGBHQ4_2(.din(n5394), .dout(n32017));
    jdff dff_B_DnQe1eps2_2(.din(n32017), .dout(n32020));
    jdff dff_B_wOc0NqTM3_2(.din(n32020), .dout(n32023));
    jdff dff_B_l2LCdCB09_2(.din(n32023), .dout(n32026));
    jdff dff_B_fMjO1sZz7_2(.din(n32026), .dout(n32029));
    jdff dff_B_D2krJ9sU8_2(.din(n32029), .dout(n32032));
    jdff dff_B_V3Tvob7D8_2(.din(n32032), .dout(n32035));
    jdff dff_B_aoBNOexl5_2(.din(n32035), .dout(n32038));
    jdff dff_B_Igy2xp7q7_2(.din(n32038), .dout(n32041));
    jdff dff_B_fPLs186h5_2(.din(n32041), .dout(n32044));
    jdff dff_B_ooSGm1Wu3_2(.din(n32044), .dout(n32047));
    jdff dff_B_EPIkemYa6_2(.din(n32047), .dout(n32050));
    jdff dff_B_0srqfk369_2(.din(n32050), .dout(n32053));
    jdff dff_B_mDjfZofs0_2(.din(n32053), .dout(n32056));
    jdff dff_B_ONRmRIjR0_2(.din(n32056), .dout(n32059));
    jdff dff_B_Fn0cynub1_2(.din(n32059), .dout(n32062));
    jdff dff_B_Cy1ke8qC5_2(.din(n32062), .dout(n32065));
    jdff dff_B_l3P9r0Z05_2(.din(n32065), .dout(n32068));
    jdff dff_B_tn8Bj7vT3_2(.din(n32068), .dout(n32071));
    jdff dff_B_ZZfgxB8n9_2(.din(n32071), .dout(n32074));
    jdff dff_B_inr8OxK96_2(.din(n32074), .dout(n32077));
    jdff dff_B_zqSBWBxZ4_2(.din(n32077), .dout(n32080));
    jdff dff_B_XdgUDHoV7_2(.din(n32080), .dout(n32083));
    jdff dff_B_qLO6wcXk4_2(.din(n32083), .dout(n32086));
    jdff dff_B_2GUUuvJi6_2(.din(n5390), .dout(n32089));
    jdff dff_B_BcUnDo3x0_2(.din(n32089), .dout(n32092));
    jdff dff_B_ZTUmweih7_2(.din(n32092), .dout(n32095));
    jdff dff_B_mnxWbeaS7_2(.din(n32095), .dout(n32098));
    jdff dff_B_mly1ZQ6m9_2(.din(n32098), .dout(n32101));
    jdff dff_B_DsxJIYWN8_2(.din(n32101), .dout(n32104));
    jdff dff_B_cSN5Cmro0_2(.din(n32104), .dout(n32107));
    jdff dff_B_CBPklAv78_2(.din(n32107), .dout(n32110));
    jdff dff_B_eYqCWvtK9_2(.din(n32110), .dout(n32113));
    jdff dff_B_JzIh3nX11_2(.din(n32113), .dout(n32116));
    jdff dff_B_R1tHNeA23_2(.din(n32116), .dout(n32119));
    jdff dff_B_y3sOlxXo1_2(.din(n32119), .dout(n32122));
    jdff dff_B_FQuTkHes5_2(.din(n32122), .dout(n32125));
    jdff dff_B_hF9g4pqb5_2(.din(n32125), .dout(n32128));
    jdff dff_B_hYx4OPiE9_2(.din(n32128), .dout(n32131));
    jdff dff_B_wqBGXGS29_2(.din(n32131), .dout(n32134));
    jdff dff_B_EVUWCY8u1_2(.din(n32134), .dout(n32137));
    jdff dff_B_AVD8uGbv5_2(.din(n32137), .dout(n32140));
    jdff dff_B_LZAS6Ncv7_2(.din(n32140), .dout(n32143));
    jdff dff_B_9Ezn80wH8_2(.din(n32143), .dout(n32146));
    jdff dff_B_drNNHBSY3_2(.din(n32146), .dout(n32149));
    jdff dff_B_40GxfDLh2_2(.din(n32149), .dout(n32152));
    jdff dff_B_hkNq5KuS4_2(.din(n32152), .dout(n32155));
    jdff dff_B_0jv3VXap9_2(.din(n32155), .dout(n32158));
    jdff dff_B_cx3cJiul8_2(.din(n32158), .dout(n32161));
    jdff dff_B_9HjdEJhl7_2(.din(n32161), .dout(n32164));
    jdff dff_B_jUVca4ae9_2(.din(n5386), .dout(n32167));
    jdff dff_B_QnmaqLHI3_1(.din(n5378), .dout(n32170));
    jdff dff_B_RTYpZfbk8_2(.din(n5075), .dout(n32173));
    jdff dff_B_1h5JXzJ86_2(.din(n32173), .dout(n32176));
    jdff dff_B_AcHC6nNx6_2(.din(n32176), .dout(n32179));
    jdff dff_B_ocXo9ELj4_2(.din(n32179), .dout(n32182));
    jdff dff_B_jKH6hJgT0_2(.din(n32182), .dout(n32185));
    jdff dff_B_ilvAowbK1_2(.din(n32185), .dout(n32188));
    jdff dff_B_VLPeSxyM5_2(.din(n32188), .dout(n32191));
    jdff dff_B_XU5Xcd4s4_2(.din(n32191), .dout(n32194));
    jdff dff_B_B89o1cIh6_2(.din(n32194), .dout(n32197));
    jdff dff_B_msrWJA2I1_2(.din(n32197), .dout(n32200));
    jdff dff_B_EzqXSzlB0_2(.din(n32200), .dout(n32203));
    jdff dff_B_GSA0RLq28_2(.din(n32203), .dout(n32206));
    jdff dff_B_yF99YuQj5_2(.din(n32206), .dout(n32209));
    jdff dff_B_myVQmF2v8_2(.din(n32209), .dout(n32212));
    jdff dff_B_H9CCqDaM9_2(.din(n32212), .dout(n32215));
    jdff dff_B_CITYv9zH7_2(.din(n32215), .dout(n32218));
    jdff dff_B_IqlDVPEu7_2(.din(n32218), .dout(n32221));
    jdff dff_B_k5spDBxP4_2(.din(n32221), .dout(n32224));
    jdff dff_B_hGmShCwr1_2(.din(n32224), .dout(n32227));
    jdff dff_B_9OR9JLkl7_2(.din(n32227), .dout(n32230));
    jdff dff_B_kehTNLxI5_2(.din(n32230), .dout(n32233));
    jdff dff_B_XzFRErpm5_2(.din(n32233), .dout(n32236));
    jdff dff_B_XOoBHcnR4_2(.din(n32236), .dout(n32239));
    jdff dff_B_5yASU09a7_1(.din(n5099), .dout(n32242));
    jdff dff_B_OLZWrOjp4_1(.din(n32242), .dout(n32245));
    jdff dff_B_olLFN9c87_2(.din(n5095), .dout(n32248));
    jdff dff_B_Oy1yACP37_2(.din(n32248), .dout(n32251));
    jdff dff_B_hILtbE4e4_2(.din(n32251), .dout(n32254));
    jdff dff_B_jAZ0UAPM5_2(.din(n32254), .dout(n32257));
    jdff dff_B_tD6kzMRP0_2(.din(n32257), .dout(n32260));
    jdff dff_B_9EfIgV226_2(.din(n32260), .dout(n32263));
    jdff dff_B_2sTwPaFB7_2(.din(n32263), .dout(n32266));
    jdff dff_B_LGlJ9LGR6_2(.din(n32266), .dout(n32269));
    jdff dff_B_Gy1z6sy28_2(.din(n32269), .dout(n32272));
    jdff dff_B_qil5CCJE2_2(.din(n32272), .dout(n32275));
    jdff dff_B_ugPp0WhU1_2(.din(n32275), .dout(n32278));
    jdff dff_B_fqUOMK534_2(.din(n32278), .dout(n32281));
    jdff dff_B_mhWh2Hty5_2(.din(n32281), .dout(n32284));
    jdff dff_B_v5OiShYa0_2(.din(n32284), .dout(n32287));
    jdff dff_B_wVN5XThm4_2(.din(n32287), .dout(n32290));
    jdff dff_B_XR9ue4V19_2(.din(n32290), .dout(n32293));
    jdff dff_B_bKVQjgk65_2(.din(n32293), .dout(n32296));
    jdff dff_B_P6lI9vI11_2(.din(n32296), .dout(n32299));
    jdff dff_B_zQGYo7ns2_2(.din(n32299), .dout(n32302));
    jdff dff_B_2TsNxkrJ7_2(.din(n32302), .dout(n32305));
    jdff dff_B_u4OSFqmP6_2(.din(n5091), .dout(n32308));
    jdff dff_B_nlfaaTG72_2(.din(n32308), .dout(n32311));
    jdff dff_B_VJVzxNCg7_2(.din(n32311), .dout(n32314));
    jdff dff_B_30SkPjq55_2(.din(n32314), .dout(n32317));
    jdff dff_B_uSQi8yFR7_2(.din(n32317), .dout(n32320));
    jdff dff_B_3Ahs3CHu0_2(.din(n32320), .dout(n32323));
    jdff dff_B_1jT8OPdh5_2(.din(n32323), .dout(n32326));
    jdff dff_B_5JuWZToz2_2(.din(n32326), .dout(n32329));
    jdff dff_B_VtPQUMxf3_2(.din(n32329), .dout(n32332));
    jdff dff_B_YH45DRSu7_2(.din(n32332), .dout(n32335));
    jdff dff_B_4APZnBpN8_2(.din(n32335), .dout(n32338));
    jdff dff_B_c0tyCitH7_2(.din(n32338), .dout(n32341));
    jdff dff_B_b4kjQ4vj9_2(.din(n32341), .dout(n32344));
    jdff dff_B_GtTC14yz3_2(.din(n32344), .dout(n32347));
    jdff dff_B_J9YPhhVi8_2(.din(n32347), .dout(n32350));
    jdff dff_B_ce6ZBtkp1_2(.din(n32350), .dout(n32353));
    jdff dff_B_EagJwI7z3_2(.din(n32353), .dout(n32356));
    jdff dff_B_x5wcMjqP2_2(.din(n32356), .dout(n32359));
    jdff dff_B_dz69GAil1_2(.din(n32359), .dout(n32362));
    jdff dff_B_USR9CEH27_2(.din(n32362), .dout(n32365));
    jdff dff_B_IVvOEBOt9_2(.din(n32365), .dout(n32368));
    jdff dff_B_IEOErc0A7_2(.din(n32368), .dout(n32371));
    jdff dff_B_fYYk5f3O9_2(.din(n5087), .dout(n32374));
    jdff dff_B_8PWg07E36_1(.din(n5079), .dout(n32377));
    jdff dff_B_OzHhAVOr8_2(.din(n4749), .dout(n32380));
    jdff dff_B_VKHez9Q05_2(.din(n32380), .dout(n32383));
    jdff dff_B_wSxZEkEG6_2(.din(n32383), .dout(n32386));
    jdff dff_B_bgpXZGrs1_2(.din(n32386), .dout(n32389));
    jdff dff_B_TQyk5DZu4_2(.din(n32389), .dout(n32392));
    jdff dff_B_iiZ26NXU0_2(.din(n32392), .dout(n32395));
    jdff dff_B_u3ZcPFKs5_2(.din(n32395), .dout(n32398));
    jdff dff_B_NH2bHgDY3_2(.din(n32398), .dout(n32401));
    jdff dff_B_KOPAkTZ98_2(.din(n32401), .dout(n32404));
    jdff dff_B_GJyHhEcH6_2(.din(n32404), .dout(n32407));
    jdff dff_B_H7y5d9bZ3_2(.din(n32407), .dout(n32410));
    jdff dff_B_tslGbXB79_2(.din(n32410), .dout(n32413));
    jdff dff_B_N1htLnBN3_2(.din(n32413), .dout(n32416));
    jdff dff_B_w00JVhEH6_2(.din(n32416), .dout(n32419));
    jdff dff_B_oZbSLAm03_2(.din(n32419), .dout(n32422));
    jdff dff_B_GFeb4tGH0_2(.din(n32422), .dout(n32425));
    jdff dff_B_2V2Ugc569_2(.din(n32425), .dout(n32428));
    jdff dff_B_VOrXH5oj5_2(.din(n32428), .dout(n32431));
    jdff dff_B_EGF4byLT4_2(.din(n32431), .dout(n32434));
    jdff dff_B_Qv0e2HCL2_1(.din(n4773), .dout(n32437));
    jdff dff_B_e2ET3Y1E7_1(.din(n32437), .dout(n32440));
    jdff dff_B_Y3Dj646E0_2(.din(n4769), .dout(n32443));
    jdff dff_B_7CvXI7ia0_2(.din(n32443), .dout(n32446));
    jdff dff_B_9xXQQOur9_2(.din(n32446), .dout(n32449));
    jdff dff_B_7HO27aZ45_2(.din(n32449), .dout(n32452));
    jdff dff_B_jJNuFAOp9_2(.din(n32452), .dout(n32455));
    jdff dff_B_cYqN30bH0_2(.din(n32455), .dout(n32458));
    jdff dff_B_DlhQfQlF8_2(.din(n32458), .dout(n32461));
    jdff dff_B_exE0wN6I5_2(.din(n32461), .dout(n32464));
    jdff dff_B_vuCazIXF0_2(.din(n32464), .dout(n32467));
    jdff dff_B_BKjuYlam2_2(.din(n32467), .dout(n32470));
    jdff dff_B_wD24toJc9_2(.din(n32470), .dout(n32473));
    jdff dff_B_MQpUhRpQ3_2(.din(n32473), .dout(n32476));
    jdff dff_B_ziTNQ1Cx2_2(.din(n32476), .dout(n32479));
    jdff dff_B_RkkV6wiZ3_2(.din(n32479), .dout(n32482));
    jdff dff_B_AxdOm1kF0_2(.din(n32482), .dout(n32485));
    jdff dff_B_7a6jpQSa0_2(.din(n32485), .dout(n32488));
    jdff dff_B_LFO4qeg28_2(.din(n4765), .dout(n32491));
    jdff dff_B_Mw2zSURz3_2(.din(n32491), .dout(n32494));
    jdff dff_B_BlHRHpQm6_2(.din(n32494), .dout(n32497));
endmodule

