/*

c6288:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jcb: 312
	jdff: 5474
	jand: 664

Summary:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jcb: 312
	jdff: 5474
	jand: 664
*/

module c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G1gat_1;
	wire [2:0] w_G1gat_2;
	wire [2:0] w_G1gat_3;
	wire [2:0] w_G1gat_4;
	wire [2:0] w_G1gat_5;
	wire [2:0] w_G1gat_6;
	wire [1:0] w_G1gat_7;
	wire [2:0] w_G18gat_0;
	wire [2:0] w_G18gat_1;
	wire [2:0] w_G18gat_2;
	wire [2:0] w_G18gat_3;
	wire [2:0] w_G18gat_4;
	wire [2:0] w_G18gat_5;
	wire [2:0] w_G18gat_6;
	wire [1:0] w_G18gat_7;
	wire [2:0] w_G35gat_0;
	wire [2:0] w_G35gat_1;
	wire [2:0] w_G35gat_2;
	wire [2:0] w_G35gat_3;
	wire [2:0] w_G35gat_4;
	wire [2:0] w_G35gat_5;
	wire [2:0] w_G35gat_6;
	wire [2:0] w_G35gat_7;
	wire [2:0] w_G52gat_0;
	wire [2:0] w_G52gat_1;
	wire [2:0] w_G52gat_2;
	wire [2:0] w_G52gat_3;
	wire [2:0] w_G52gat_4;
	wire [2:0] w_G52gat_5;
	wire [2:0] w_G52gat_6;
	wire [2:0] w_G52gat_7;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G69gat_1;
	wire [2:0] w_G69gat_2;
	wire [2:0] w_G69gat_3;
	wire [2:0] w_G69gat_4;
	wire [2:0] w_G69gat_5;
	wire [2:0] w_G69gat_6;
	wire [1:0] w_G69gat_7;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G86gat_1;
	wire [2:0] w_G86gat_2;
	wire [2:0] w_G86gat_3;
	wire [2:0] w_G86gat_4;
	wire [2:0] w_G86gat_5;
	wire [2:0] w_G86gat_6;
	wire [1:0] w_G86gat_7;
	wire [2:0] w_G103gat_0;
	wire [2:0] w_G103gat_1;
	wire [2:0] w_G103gat_2;
	wire [2:0] w_G103gat_3;
	wire [2:0] w_G103gat_4;
	wire [2:0] w_G103gat_5;
	wire [2:0] w_G103gat_6;
	wire [1:0] w_G103gat_7;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G120gat_1;
	wire [2:0] w_G120gat_2;
	wire [2:0] w_G120gat_3;
	wire [2:0] w_G120gat_4;
	wire [2:0] w_G120gat_5;
	wire [2:0] w_G120gat_6;
	wire [1:0] w_G120gat_7;
	wire [2:0] w_G137gat_0;
	wire [2:0] w_G137gat_1;
	wire [2:0] w_G137gat_2;
	wire [2:0] w_G137gat_3;
	wire [2:0] w_G137gat_4;
	wire [2:0] w_G137gat_5;
	wire [2:0] w_G137gat_6;
	wire [1:0] w_G137gat_7;
	wire [2:0] w_G154gat_0;
	wire [2:0] w_G154gat_1;
	wire [2:0] w_G154gat_2;
	wire [2:0] w_G154gat_3;
	wire [2:0] w_G154gat_4;
	wire [2:0] w_G154gat_5;
	wire [2:0] w_G154gat_6;
	wire [1:0] w_G154gat_7;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G171gat_2;
	wire [2:0] w_G171gat_3;
	wire [2:0] w_G171gat_4;
	wire [2:0] w_G171gat_5;
	wire [2:0] w_G171gat_6;
	wire [1:0] w_G171gat_7;
	wire [2:0] w_G188gat_0;
	wire [2:0] w_G188gat_1;
	wire [2:0] w_G188gat_2;
	wire [2:0] w_G188gat_3;
	wire [2:0] w_G188gat_4;
	wire [2:0] w_G188gat_5;
	wire [2:0] w_G188gat_6;
	wire [1:0] w_G188gat_7;
	wire [2:0] w_G205gat_0;
	wire [2:0] w_G205gat_1;
	wire [2:0] w_G205gat_2;
	wire [2:0] w_G205gat_3;
	wire [2:0] w_G205gat_4;
	wire [2:0] w_G205gat_5;
	wire [2:0] w_G205gat_6;
	wire [1:0] w_G205gat_7;
	wire [2:0] w_G222gat_0;
	wire [2:0] w_G222gat_1;
	wire [2:0] w_G222gat_2;
	wire [2:0] w_G222gat_3;
	wire [2:0] w_G222gat_4;
	wire [2:0] w_G222gat_5;
	wire [2:0] w_G222gat_6;
	wire [1:0] w_G222gat_7;
	wire [2:0] w_G239gat_0;
	wire [2:0] w_G239gat_1;
	wire [2:0] w_G239gat_2;
	wire [2:0] w_G239gat_3;
	wire [2:0] w_G239gat_4;
	wire [2:0] w_G239gat_5;
	wire [2:0] w_G239gat_6;
	wire [1:0] w_G239gat_7;
	wire [2:0] w_G256gat_0;
	wire [2:0] w_G256gat_1;
	wire [2:0] w_G256gat_2;
	wire [2:0] w_G256gat_3;
	wire [2:0] w_G256gat_4;
	wire [2:0] w_G256gat_5;
	wire [2:0] w_G256gat_6;
	wire [1:0] w_G256gat_7;
	wire [2:0] w_G273gat_0;
	wire [2:0] w_G273gat_1;
	wire [2:0] w_G273gat_2;
	wire [2:0] w_G273gat_3;
	wire [2:0] w_G273gat_4;
	wire [2:0] w_G273gat_5;
	wire [2:0] w_G273gat_6;
	wire [1:0] w_G273gat_7;
	wire [2:0] w_G290gat_0;
	wire [2:0] w_G290gat_1;
	wire [2:0] w_G290gat_2;
	wire [2:0] w_G290gat_3;
	wire [2:0] w_G290gat_4;
	wire [2:0] w_G290gat_5;
	wire [2:0] w_G290gat_6;
	wire [2:0] w_G290gat_7;
	wire [2:0] w_G307gat_0;
	wire [2:0] w_G307gat_1;
	wire [2:0] w_G307gat_2;
	wire [2:0] w_G307gat_3;
	wire [2:0] w_G307gat_4;
	wire [2:0] w_G307gat_5;
	wire [2:0] w_G307gat_6;
	wire [1:0] w_G307gat_7;
	wire [2:0] w_G324gat_0;
	wire [2:0] w_G324gat_1;
	wire [2:0] w_G324gat_2;
	wire [2:0] w_G324gat_3;
	wire [2:0] w_G324gat_4;
	wire [2:0] w_G324gat_5;
	wire [2:0] w_G324gat_6;
	wire [1:0] w_G324gat_7;
	wire [2:0] w_G341gat_0;
	wire [2:0] w_G341gat_1;
	wire [2:0] w_G341gat_2;
	wire [2:0] w_G341gat_3;
	wire [2:0] w_G341gat_4;
	wire [2:0] w_G341gat_5;
	wire [2:0] w_G341gat_6;
	wire [1:0] w_G341gat_7;
	wire [2:0] w_G358gat_0;
	wire [2:0] w_G358gat_1;
	wire [2:0] w_G358gat_2;
	wire [2:0] w_G358gat_3;
	wire [2:0] w_G358gat_4;
	wire [2:0] w_G358gat_5;
	wire [2:0] w_G358gat_6;
	wire [1:0] w_G358gat_7;
	wire [2:0] w_G375gat_0;
	wire [2:0] w_G375gat_1;
	wire [2:0] w_G375gat_2;
	wire [2:0] w_G375gat_3;
	wire [2:0] w_G375gat_4;
	wire [2:0] w_G375gat_5;
	wire [2:0] w_G375gat_6;
	wire [1:0] w_G375gat_7;
	wire [2:0] w_G392gat_0;
	wire [2:0] w_G392gat_1;
	wire [2:0] w_G392gat_2;
	wire [2:0] w_G392gat_3;
	wire [2:0] w_G392gat_4;
	wire [2:0] w_G392gat_5;
	wire [2:0] w_G392gat_6;
	wire [1:0] w_G392gat_7;
	wire [2:0] w_G409gat_0;
	wire [2:0] w_G409gat_1;
	wire [2:0] w_G409gat_2;
	wire [2:0] w_G409gat_3;
	wire [2:0] w_G409gat_4;
	wire [2:0] w_G409gat_5;
	wire [2:0] w_G409gat_6;
	wire [1:0] w_G409gat_7;
	wire [2:0] w_G426gat_0;
	wire [2:0] w_G426gat_1;
	wire [2:0] w_G426gat_2;
	wire [2:0] w_G426gat_3;
	wire [2:0] w_G426gat_4;
	wire [2:0] w_G426gat_5;
	wire [2:0] w_G426gat_6;
	wire [1:0] w_G426gat_7;
	wire [2:0] w_G443gat_0;
	wire [2:0] w_G443gat_1;
	wire [2:0] w_G443gat_2;
	wire [2:0] w_G443gat_3;
	wire [2:0] w_G443gat_4;
	wire [2:0] w_G443gat_5;
	wire [2:0] w_G443gat_6;
	wire [1:0] w_G443gat_7;
	wire [2:0] w_G460gat_0;
	wire [2:0] w_G460gat_1;
	wire [2:0] w_G460gat_2;
	wire [2:0] w_G460gat_3;
	wire [2:0] w_G460gat_4;
	wire [2:0] w_G460gat_5;
	wire [2:0] w_G460gat_6;
	wire [1:0] w_G460gat_7;
	wire [2:0] w_G477gat_0;
	wire [2:0] w_G477gat_1;
	wire [2:0] w_G477gat_2;
	wire [2:0] w_G477gat_3;
	wire [2:0] w_G477gat_4;
	wire [2:0] w_G477gat_5;
	wire [2:0] w_G477gat_6;
	wire [1:0] w_G477gat_7;
	wire [2:0] w_G494gat_0;
	wire [2:0] w_G494gat_1;
	wire [2:0] w_G494gat_2;
	wire [2:0] w_G494gat_3;
	wire [2:0] w_G494gat_4;
	wire [2:0] w_G494gat_5;
	wire [2:0] w_G494gat_6;
	wire [1:0] w_G494gat_7;
	wire [2:0] w_G511gat_0;
	wire [2:0] w_G511gat_1;
	wire [2:0] w_G511gat_2;
	wire [2:0] w_G511gat_3;
	wire [2:0] w_G511gat_4;
	wire [2:0] w_G511gat_5;
	wire [2:0] w_G511gat_6;
	wire [1:0] w_G511gat_7;
	wire [2:0] w_G528gat_0;
	wire [2:0] w_G528gat_1;
	wire [2:0] w_G528gat_2;
	wire [2:0] w_G528gat_3;
	wire [2:0] w_G528gat_4;
	wire [2:0] w_G528gat_5;
	wire [2:0] w_G528gat_6;
	wire [1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire [1:0] w_n65_0;
	wire [1:0] w_n66_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [2:0] w_n80_0;
	wire [1:0] w_n83_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [1:0] w_n90_0;
	wire [1:0] w_n91_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n99_0;
	wire [2:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n112_0;
	wire [2:0] w_n117_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n123_0;
	wire [1:0] w_n125_0;
	wire [1:0] w_n127_0;
	wire [1:0] w_n128_0;
	wire [1:0] w_n129_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n132_0;
	wire [1:0] w_n133_0;
	wire [1:0] w_n135_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n141_0;
	wire [2:0] w_n146_0;
	wire [1:0] w_n148_0;
	wire [1:0] w_n152_0;
	wire [1:0] w_n154_0;
	wire [1:0] w_n155_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n157_0;
	wire [1:0] w_n158_0;
	wire [1:0] w_n160_0;
	wire [1:0] w_n161_0;
	wire [1:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n165_0;
	wire [1:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n175_0;
	wire [1:0] w_n176_0;
	wire [2:0] w_n181_0;
	wire [1:0] w_n183_0;
	wire [1:0] w_n186_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n192_0;
	wire [1:0] w_n194_0;
	wire [1:0] w_n195_0;
	wire [2:0] w_n196_0;
	wire [1:0] w_n198_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n203_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n209_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n212_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n218_0;
	wire [2:0] w_n223_0;
	wire [1:0] w_n225_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n230_0;
	wire [1:0] w_n233_0;
	wire [1:0] w_n235_0;
	wire [1:0] w_n239_0;
	wire [1:0] w_n241_0;
	wire [1:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [1:0] w_n245_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n248_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n250_0;
	wire [1:0] w_n251_0;
	wire [1:0] w_n252_0;
	wire [1:0] w_n253_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n256_0;
	wire [1:0] w_n258_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n266_0;
	wire [1:0] w_n267_0;
	wire [2:0] w_n272_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n277_0;
	wire [1:0] w_n279_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n284_0;
	wire [1:0] w_n287_0;
	wire [1:0] w_n289_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n296_0;
	wire [2:0] w_n297_0;
	wire [1:0] w_n299_0;
	wire [1:0] w_n301_0;
	wire [1:0] w_n302_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n304_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n306_0;
	wire [1:0] w_n307_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n309_0;
	wire [1:0] w_n310_0;
	wire [1:0] w_n311_0;
	wire [1:0] w_n312_0;
	wire [1:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n317_0;
	wire [1:0] w_n322_0;
	wire [1:0] w_n323_0;
	wire [2:0] w_n328_0;
	wire [1:0] w_n330_0;
	wire [1:0] w_n333_0;
	wire [1:0] w_n335_0;
	wire [1:0] w_n338_0;
	wire [1:0] w_n340_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n345_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n354_0;
	wire [1:0] w_n356_0;
	wire [1:0] w_n357_0;
	wire [2:0] w_n358_0;
	wire [1:0] w_n360_0;
	wire [1:0] w_n362_0;
	wire [1:0] w_n363_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n365_0;
	wire [1:0] w_n366_0;
	wire [1:0] w_n367_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n369_0;
	wire [1:0] w_n370_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n375_0;
	wire [1:0] w_n377_0;
	wire [1:0] w_n378_0;
	wire [1:0] w_n380_0;
	wire [1:0] w_n385_0;
	wire [1:0] w_n386_0;
	wire [2:0] w_n391_0;
	wire [1:0] w_n393_0;
	wire [1:0] w_n396_0;
	wire [1:0] w_n398_0;
	wire [1:0] w_n401_0;
	wire [1:0] w_n403_0;
	wire [1:0] w_n406_0;
	wire [1:0] w_n408_0;
	wire [1:0] w_n411_0;
	wire [1:0] w_n413_0;
	wire [1:0] w_n416_0;
	wire [1:0] w_n418_0;
	wire [1:0] w_n423_0;
	wire [1:0] w_n425_0;
	wire [1:0] w_n426_0;
	wire [2:0] w_n427_0;
	wire [1:0] w_n429_0;
	wire [1:0] w_n431_0;
	wire [1:0] w_n432_0;
	wire [1:0] w_n433_0;
	wire [1:0] w_n434_0;
	wire [1:0] w_n435_0;
	wire [1:0] w_n436_0;
	wire [1:0] w_n437_0;
	wire [1:0] w_n438_0;
	wire [1:0] w_n439_0;
	wire [1:0] w_n440_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n442_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n444_0;
	wire [1:0] w_n445_0;
	wire [1:0] w_n446_0;
	wire [1:0] w_n448_0;
	wire [1:0] w_n449_0;
	wire [1:0] w_n451_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n464_0;
	wire [1:0] w_n467_0;
	wire [1:0] w_n469_0;
	wire [1:0] w_n472_0;
	wire [1:0] w_n474_0;
	wire [1:0] w_n477_0;
	wire [1:0] w_n479_0;
	wire [1:0] w_n482_0;
	wire [1:0] w_n484_0;
	wire [1:0] w_n487_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n492_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n499_0;
	wire [1:0] w_n501_0;
	wire [1:0] w_n502_0;
	wire [2:0] w_n503_0;
	wire [1:0] w_n505_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n508_0;
	wire [1:0] w_n509_0;
	wire [1:0] w_n510_0;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n513_0;
	wire [1:0] w_n514_0;
	wire [1:0] w_n515_0;
	wire [1:0] w_n516_0;
	wire [1:0] w_n517_0;
	wire [1:0] w_n518_0;
	wire [1:0] w_n519_0;
	wire [1:0] w_n520_0;
	wire [1:0] w_n521_0;
	wire [1:0] w_n522_0;
	wire [1:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n526_0;
	wire [1:0] w_n527_0;
	wire [1:0] w_n529_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n535_0;
	wire [2:0] w_n540_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n545_0;
	wire [1:0] w_n547_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n552_0;
	wire [1:0] w_n555_0;
	wire [1:0] w_n557_0;
	wire [1:0] w_n560_0;
	wire [1:0] w_n562_0;
	wire [1:0] w_n565_0;
	wire [1:0] w_n567_0;
	wire [1:0] w_n570_0;
	wire [1:0] w_n572_0;
	wire [1:0] w_n575_0;
	wire [1:0] w_n577_0;
	wire [1:0] w_n582_0;
	wire [1:0] w_n584_0;
	wire [1:0] w_n585_0;
	wire [2:0] w_n586_0;
	wire [1:0] w_n588_0;
	wire [1:0] w_n590_0;
	wire [1:0] w_n591_0;
	wire [1:0] w_n592_0;
	wire [1:0] w_n593_0;
	wire [1:0] w_n594_0;
	wire [1:0] w_n595_0;
	wire [1:0] w_n596_0;
	wire [1:0] w_n597_0;
	wire [1:0] w_n598_0;
	wire [1:0] w_n599_0;
	wire [1:0] w_n600_0;
	wire [1:0] w_n601_0;
	wire [1:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [1:0] w_n604_0;
	wire [1:0] w_n605_0;
	wire [1:0] w_n606_0;
	wire [1:0] w_n607_0;
	wire [1:0] w_n608_0;
	wire [1:0] w_n609_0;
	wire [1:0] w_n611_0;
	wire [1:0] w_n612_0;
	wire [1:0] w_n614_0;
	wire [1:0] w_n619_0;
	wire [1:0] w_n620_0;
	wire [2:0] w_n625_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n630_0;
	wire [1:0] w_n632_0;
	wire [1:0] w_n635_0;
	wire [1:0] w_n637_0;
	wire [1:0] w_n640_0;
	wire [1:0] w_n642_0;
	wire [1:0] w_n645_0;
	wire [1:0] w_n647_0;
	wire [1:0] w_n650_0;
	wire [1:0] w_n652_0;
	wire [1:0] w_n655_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n660_0;
	wire [1:0] w_n662_0;
	wire [1:0] w_n665_0;
	wire [1:0] w_n667_0;
	wire [1:0] w_n672_0;
	wire [1:0] w_n674_0;
	wire [1:0] w_n675_0;
	wire [2:0] w_n676_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n680_0;
	wire [1:0] w_n681_0;
	wire [1:0] w_n682_0;
	wire [1:0] w_n683_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n688_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n691_0;
	wire [1:0] w_n692_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n694_0;
	wire [1:0] w_n695_0;
	wire [1:0] w_n696_0;
	wire [1:0] w_n697_0;
	wire [1:0] w_n698_0;
	wire [1:0] w_n699_0;
	wire [1:0] w_n700_0;
	wire [1:0] w_n701_0;
	wire [1:0] w_n703_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n706_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n712_0;
	wire [2:0] w_n717_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n722_0;
	wire [1:0] w_n724_0;
	wire [1:0] w_n727_0;
	wire [1:0] w_n729_0;
	wire [1:0] w_n732_0;
	wire [1:0] w_n734_0;
	wire [1:0] w_n737_0;
	wire [1:0] w_n739_0;
	wire [1:0] w_n742_0;
	wire [1:0] w_n744_0;
	wire [1:0] w_n747_0;
	wire [1:0] w_n749_0;
	wire [1:0] w_n752_0;
	wire [1:0] w_n754_0;
	wire [1:0] w_n757_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n762_0;
	wire [1:0] w_n764_0;
	wire [1:0] w_n769_0;
	wire [1:0] w_n771_0;
	wire [1:0] w_n772_0;
	wire [1:0] w_n773_0;
	wire [1:0] w_n774_0;
	wire [1:0] w_n775_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n778_0;
	wire [1:0] w_n779_0;
	wire [1:0] w_n780_0;
	wire [1:0] w_n781_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n783_0;
	wire [1:0] w_n784_0;
	wire [1:0] w_n785_0;
	wire [1:0] w_n786_0;
	wire [1:0] w_n787_0;
	wire [1:0] w_n788_0;
	wire [1:0] w_n789_0;
	wire [1:0] w_n790_0;
	wire [1:0] w_n791_0;
	wire [1:0] w_n792_0;
	wire [1:0] w_n793_0;
	wire [1:0] w_n794_0;
	wire [1:0] w_n795_0;
	wire [1:0] w_n796_0;
	wire [1:0] w_n797_0;
	wire [1:0] w_n798_0;
	wire [1:0] w_n799_0;
	wire [1:0] w_n800_0;
	wire [1:0] w_n802_0;
	wire [1:0] w_n803_0;
	wire [1:0] w_n805_0;
	wire [1:0] w_n810_0;
	wire [1:0] w_n811_0;
	wire [1:0] w_n815_0;
	wire [1:0] w_n816_0;
	wire [2:0] w_n820_0;
	wire [1:0] w_n822_0;
	wire [1:0] w_n825_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n830_0;
	wire [1:0] w_n832_0;
	wire [1:0] w_n835_0;
	wire [1:0] w_n837_0;
	wire [1:0] w_n840_0;
	wire [1:0] w_n842_0;
	wire [1:0] w_n845_0;
	wire [1:0] w_n847_0;
	wire [1:0] w_n850_0;
	wire [1:0] w_n852_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n857_0;
	wire [1:0] w_n860_0;
	wire [1:0] w_n862_0;
	wire [1:0] w_n865_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n872_0;
	wire [1:0] w_n874_0;
	wire [1:0] w_n875_0;
	wire [1:0] w_n877_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n880_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n882_0;
	wire [1:0] w_n883_0;
	wire [1:0] w_n884_0;
	wire [1:0] w_n885_0;
	wire [1:0] w_n886_0;
	wire [1:0] w_n887_0;
	wire [1:0] w_n888_0;
	wire [1:0] w_n889_0;
	wire [1:0] w_n890_0;
	wire [1:0] w_n891_0;
	wire [1:0] w_n892_0;
	wire [1:0] w_n893_0;
	wire [1:0] w_n894_0;
	wire [1:0] w_n895_0;
	wire [1:0] w_n896_0;
	wire [1:0] w_n897_0;
	wire [1:0] w_n898_0;
	wire [1:0] w_n899_0;
	wire [2:0] w_n900_0;
	wire [1:0] w_n902_0;
	wire [1:0] w_n903_0;
	wire [1:0] w_n904_0;
	wire [1:0] w_n905_0;
	wire [1:0] w_n910_0;
	wire [1:0] w_n911_0;
	wire [2:0] w_n915_0;
	wire [1:0] w_n916_0;
	wire [1:0] w_n922_0;
	wire [1:0] w_n924_0;
	wire [1:0] w_n927_0;
	wire [1:0] w_n929_0;
	wire [1:0] w_n932_0;
	wire [1:0] w_n934_0;
	wire [1:0] w_n937_0;
	wire [1:0] w_n939_0;
	wire [1:0] w_n942_0;
	wire [1:0] w_n944_0;
	wire [1:0] w_n947_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n952_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n959_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n967_0;
	wire [1:0] w_n969_0;
	wire [1:0] w_n972_0;
	wire [1:0] w_n974_0;
	wire [1:0] w_n978_0;
	wire [1:0] w_n980_0;
	wire [1:0] w_n982_0;
	wire [1:0] w_n983_0;
	wire [1:0] w_n984_0;
	wire [1:0] w_n985_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n987_0;
	wire [1:0] w_n988_0;
	wire [1:0] w_n989_0;
	wire [1:0] w_n990_0;
	wire [1:0] w_n991_0;
	wire [1:0] w_n992_0;
	wire [1:0] w_n993_0;
	wire [1:0] w_n994_0;
	wire [1:0] w_n995_0;
	wire [1:0] w_n996_0;
	wire [1:0] w_n997_0;
	wire [1:0] w_n998_0;
	wire [1:0] w_n999_0;
	wire [1:0] w_n1000_0;
	wire [1:0] w_n1001_0;
	wire [1:0] w_n1002_0;
	wire [1:0] w_n1003_0;
	wire [1:0] w_n1004_0;
	wire [1:0] w_n1005_0;
	wire [1:0] w_n1006_0;
	wire [1:0] w_n1007_0;
	wire [1:0] w_n1008_0;
	wire [1:0] w_n1009_0;
	wire [1:0] w_n1011_0;
	wire [1:0] w_n1013_0;
	wire [1:0] w_n1017_0;
	wire [1:0] w_n1018_0;
	wire [1:0] w_n1022_0;
	wire [1:0] w_n1023_0;
	wire [1:0] w_n1026_0;
	wire [1:0] w_n1028_0;
	wire [1:0] w_n1031_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1036_0;
	wire [1:0] w_n1038_0;
	wire [1:0] w_n1041_0;
	wire [1:0] w_n1043_0;
	wire [1:0] w_n1046_0;
	wire [1:0] w_n1048_0;
	wire [1:0] w_n1051_0;
	wire [1:0] w_n1053_0;
	wire [1:0] w_n1056_0;
	wire [1:0] w_n1058_0;
	wire [1:0] w_n1061_0;
	wire [1:0] w_n1063_0;
	wire [1:0] w_n1066_0;
	wire [1:0] w_n1068_0;
	wire [1:0] w_n1071_0;
	wire [1:0] w_n1073_0;
	wire [1:0] w_n1076_0;
	wire [1:0] w_n1077_0;
	wire [1:0] w_n1078_0;
	wire [1:0] w_n1080_0;
	wire [1:0] w_n1082_0;
	wire [1:0] w_n1083_0;
	wire [1:0] w_n1084_0;
	wire [1:0] w_n1085_0;
	wire [1:0] w_n1086_0;
	wire [1:0] w_n1087_0;
	wire [1:0] w_n1088_0;
	wire [1:0] w_n1089_0;
	wire [1:0] w_n1090_0;
	wire [1:0] w_n1091_0;
	wire [1:0] w_n1092_0;
	wire [1:0] w_n1093_0;
	wire [1:0] w_n1094_0;
	wire [1:0] w_n1095_0;
	wire [1:0] w_n1096_0;
	wire [1:0] w_n1097_0;
	wire [1:0] w_n1098_0;
	wire [1:0] w_n1099_0;
	wire [1:0] w_n1100_0;
	wire [1:0] w_n1101_0;
	wire [1:0] w_n1102_0;
	wire [1:0] w_n1103_0;
	wire [1:0] w_n1105_0;
	wire [1:0] w_n1106_0;
	wire [1:0] w_n1107_0;
	wire [1:0] w_n1108_0;
	wire [1:0] w_n1109_0;
	wire [1:0] w_n1115_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1120_0;
	wire [1:0] w_n1124_0;
	wire [1:0] w_n1126_0;
	wire [1:0] w_n1129_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1134_0;
	wire [1:0] w_n1136_0;
	wire [1:0] w_n1139_0;
	wire [1:0] w_n1141_0;
	wire [1:0] w_n1144_0;
	wire [1:0] w_n1146_0;
	wire [1:0] w_n1149_0;
	wire [1:0] w_n1151_0;
	wire [1:0] w_n1154_0;
	wire [1:0] w_n1156_0;
	wire [1:0] w_n1159_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1166_0;
	wire [1:0] w_n1169_0;
	wire [1:0] w_n1171_0;
	wire [1:0] w_n1174_0;
	wire [1:0] w_n1175_0;
	wire [1:0] w_n1176_0;
	wire [1:0] w_n1179_0;
	wire [1:0] w_n1181_0;
	wire [1:0] w_n1182_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1184_0;
	wire [1:0] w_n1185_0;
	wire [1:0] w_n1186_0;
	wire [1:0] w_n1187_0;
	wire [1:0] w_n1188_0;
	wire [1:0] w_n1189_0;
	wire [1:0] w_n1190_0;
	wire [1:0] w_n1191_0;
	wire [1:0] w_n1192_0;
	wire [1:0] w_n1193_0;
	wire [1:0] w_n1194_0;
	wire [1:0] w_n1195_0;
	wire [1:0] w_n1196_0;
	wire [1:0] w_n1197_0;
	wire [1:0] w_n1198_0;
	wire [1:0] w_n1199_0;
	wire [1:0] w_n1200_0;
	wire [1:0] w_n1201_0;
	wire [1:0] w_n1203_0;
	wire [1:0] w_n1205_0;
	wire [1:0] w_n1206_0;
	wire [1:0] w_n1207_0;
	wire [1:0] w_n1213_0;
	wire [1:0] w_n1216_0;
	wire [1:0] w_n1217_0;
	wire [1:0] w_n1220_0;
	wire [1:0] w_n1222_0;
	wire [1:0] w_n1225_0;
	wire [1:0] w_n1227_0;
	wire [1:0] w_n1230_0;
	wire [1:0] w_n1232_0;
	wire [1:0] w_n1235_0;
	wire [1:0] w_n1237_0;
	wire [1:0] w_n1240_0;
	wire [1:0] w_n1242_0;
	wire [1:0] w_n1245_0;
	wire [1:0] w_n1247_0;
	wire [1:0] w_n1250_0;
	wire [1:0] w_n1252_0;
	wire [1:0] w_n1255_0;
	wire [1:0] w_n1257_0;
	wire [1:0] w_n1260_0;
	wire [1:0] w_n1262_0;
	wire [1:0] w_n1265_0;
	wire [1:0] w_n1266_0;
	wire [1:0] w_n1267_0;
	wire [1:0] w_n1270_0;
	wire [1:0] w_n1272_0;
	wire [1:0] w_n1273_0;
	wire [1:0] w_n1274_0;
	wire [1:0] w_n1275_0;
	wire [1:0] w_n1276_0;
	wire [1:0] w_n1277_0;
	wire [1:0] w_n1278_0;
	wire [1:0] w_n1279_0;
	wire [1:0] w_n1280_0;
	wire [1:0] w_n1281_0;
	wire [1:0] w_n1282_0;
	wire [1:0] w_n1283_0;
	wire [1:0] w_n1284_0;
	wire [1:0] w_n1285_0;
	wire [1:0] w_n1286_0;
	wire [1:0] w_n1287_0;
	wire [1:0] w_n1288_0;
	wire [1:0] w_n1289_0;
	wire [1:0] w_n1290_0;
	wire [1:0] w_n1291_0;
	wire [1:0] w_n1293_0;
	wire [1:0] w_n1294_0;
	wire [1:0] w_n1295_0;
	wire [1:0] w_n1301_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1307_0;
	wire [1:0] w_n1310_0;
	wire [1:0] w_n1312_0;
	wire [1:0] w_n1315_0;
	wire [1:0] w_n1317_0;
	wire [1:0] w_n1320_0;
	wire [1:0] w_n1322_0;
	wire [1:0] w_n1325_0;
	wire [1:0] w_n1327_0;
	wire [1:0] w_n1330_0;
	wire [1:0] w_n1332_0;
	wire [1:0] w_n1335_0;
	wire [1:0] w_n1337_0;
	wire [1:0] w_n1340_0;
	wire [1:0] w_n1342_0;
	wire [1:0] w_n1345_0;
	wire [1:0] w_n1347_0;
	wire [1:0] w_n1350_0;
	wire [1:0] w_n1351_0;
	wire [1:0] w_n1352_0;
	wire [1:0] w_n1355_0;
	wire [1:0] w_n1357_0;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1359_0;
	wire [1:0] w_n1360_0;
	wire [1:0] w_n1361_0;
	wire [1:0] w_n1362_0;
	wire [1:0] w_n1363_0;
	wire [1:0] w_n1364_0;
	wire [1:0] w_n1365_0;
	wire [1:0] w_n1366_0;
	wire [1:0] w_n1367_0;
	wire [1:0] w_n1368_0;
	wire [1:0] w_n1369_0;
	wire [1:0] w_n1370_0;
	wire [1:0] w_n1371_0;
	wire [1:0] w_n1372_0;
	wire [1:0] w_n1373_0;
	wire [1:0] w_n1374_0;
	wire [1:0] w_n1376_0;
	wire [1:0] w_n1378_0;
	wire [1:0] w_n1379_0;
	wire [1:0] w_n1384_0;
	wire [1:0] w_n1389_0;
	wire [1:0] w_n1390_0;
	wire [1:0] w_n1393_0;
	wire [1:0] w_n1395_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1400_0;
	wire [1:0] w_n1403_0;
	wire [1:0] w_n1405_0;
	wire [1:0] w_n1408_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1413_0;
	wire [1:0] w_n1415_0;
	wire [1:0] w_n1418_0;
	wire [1:0] w_n1420_0;
	wire [1:0] w_n1423_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1428_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1430_0;
	wire [1:0] w_n1433_0;
	wire [1:0] w_n1435_0;
	wire [1:0] w_n1436_0;
	wire [1:0] w_n1437_0;
	wire [1:0] w_n1438_0;
	wire [1:0] w_n1439_0;
	wire [1:0] w_n1440_0;
	wire [1:0] w_n1441_0;
	wire [1:0] w_n1442_0;
	wire [1:0] w_n1443_0;
	wire [1:0] w_n1444_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1448_0;
	wire [1:0] w_n1449_0;
	wire [1:0] w_n1450_0;
	wire [1:0] w_n1452_0;
	wire [1:0] w_n1454_0;
	wire [1:0] w_n1455_0;
	wire [1:0] w_n1460_0;
	wire [1:0] w_n1465_0;
	wire [1:0] w_n1466_0;
	wire [1:0] w_n1469_0;
	wire [1:0] w_n1471_0;
	wire [1:0] w_n1474_0;
	wire [1:0] w_n1476_0;
	wire [1:0] w_n1479_0;
	wire [1:0] w_n1481_0;
	wire [1:0] w_n1484_0;
	wire [1:0] w_n1486_0;
	wire [1:0] w_n1489_0;
	wire [1:0] w_n1491_0;
	wire [1:0] w_n1494_0;
	wire [1:0] w_n1496_0;
	wire [1:0] w_n1499_0;
	wire [1:0] w_n1500_0;
	wire [1:0] w_n1501_0;
	wire [1:0] w_n1504_0;
	wire [1:0] w_n1506_0;
	wire [1:0] w_n1507_0;
	wire [1:0] w_n1508_0;
	wire [1:0] w_n1509_0;
	wire [1:0] w_n1510_0;
	wire [1:0] w_n1511_0;
	wire [1:0] w_n1512_0;
	wire [1:0] w_n1513_0;
	wire [1:0] w_n1514_0;
	wire [1:0] w_n1515_0;
	wire [1:0] w_n1516_0;
	wire [1:0] w_n1517_0;
	wire [1:0] w_n1518_0;
	wire [1:0] w_n1519_0;
	wire [1:0] w_n1521_0;
	wire [1:0] w_n1523_0;
	wire [1:0] w_n1524_0;
	wire [1:0] w_n1529_0;
	wire [1:0] w_n1534_0;
	wire [1:0] w_n1535_0;
	wire [1:0] w_n1538_0;
	wire [1:0] w_n1540_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1548_0;
	wire [1:0] w_n1550_0;
	wire [1:0] w_n1553_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1558_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1563_0;
	wire [1:0] w_n1564_0;
	wire [1:0] w_n1565_0;
	wire [1:0] w_n1568_0;
	wire [1:0] w_n1570_0;
	wire [1:0] w_n1571_0;
	wire [1:0] w_n1572_0;
	wire [1:0] w_n1573_0;
	wire [1:0] w_n1574_0;
	wire [1:0] w_n1575_0;
	wire [1:0] w_n1576_0;
	wire [1:0] w_n1577_0;
	wire [1:0] w_n1578_0;
	wire [1:0] w_n1579_0;
	wire [1:0] w_n1580_0;
	wire [1:0] w_n1581_0;
	wire [1:0] w_n1583_0;
	wire [1:0] w_n1585_0;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1597_0;
	wire [1:0] w_n1600_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1607_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1612_0;
	wire [1:0] w_n1615_0;
	wire [1:0] w_n1617_0;
	wire [1:0] w_n1620_0;
	wire [1:0] w_n1621_0;
	wire [1:0] w_n1622_0;
	wire [1:0] w_n1625_0;
	wire [1:0] w_n1627_0;
	wire [1:0] w_n1628_0;
	wire [1:0] w_n1629_0;
	wire [1:0] w_n1630_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1632_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1634_0;
	wire [1:0] w_n1635_0;
	wire [1:0] w_n1636_0;
	wire [1:0] w_n1638_0;
	wire [1:0] w_n1640_0;
	wire [1:0] w_n1641_0;
	wire [1:0] w_n1646_0;
	wire [1:0] w_n1651_0;
	wire [1:0] w_n1653_0;
	wire [1:0] w_n1656_0;
	wire [1:0] w_n1658_0;
	wire [1:0] w_n1661_0;
	wire [1:0] w_n1663_0;
	wire [1:0] w_n1666_0;
	wire [1:0] w_n1668_0;
	wire [1:0] w_n1671_0;
	wire [1:0] w_n1672_0;
	wire [1:0] w_n1673_0;
	wire [1:0] w_n1676_0;
	wire [1:0] w_n1678_0;
	wire [1:0] w_n1679_0;
	wire [1:0] w_n1680_0;
	wire [1:0] w_n1681_0;
	wire [1:0] w_n1682_0;
	wire [1:0] w_n1683_0;
	wire [1:0] w_n1684_0;
	wire [1:0] w_n1685_0;
	wire [1:0] w_n1686_0;
	wire [1:0] w_n1688_0;
	wire [1:0] w_n1689_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1697_0;
	wire [1:0] w_n1699_0;
	wire [1:0] w_n1702_0;
	wire [1:0] w_n1704_0;
	wire [1:0] w_n1707_0;
	wire [1:0] w_n1709_0;
	wire [1:0] w_n1712_0;
	wire [1:0] w_n1713_0;
	wire [1:0] w_n1714_0;
	wire [1:0] w_n1717_0;
	wire [1:0] w_n1719_0;
	wire [1:0] w_n1720_0;
	wire [1:0] w_n1721_0;
	wire [1:0] w_n1722_0;
	wire [1:0] w_n1723_0;
	wire [1:0] w_n1724_0;
	wire [1:0] w_n1725_0;
	wire [1:0] w_n1726_0;
	wire [1:0] w_n1727_0;
	wire [1:0] w_n1734_0;
	wire [1:0] w_n1737_0;
	wire [1:0] w_n1739_0;
	wire [1:0] w_n1742_0;
	wire [1:0] w_n1744_0;
	wire [1:0] w_n1747_0;
	wire [1:0] w_n1748_0;
	wire [1:0] w_n1749_0;
	wire [1:0] w_n1752_0;
	wire [1:0] w_n1754_0;
	wire [1:0] w_n1755_0;
	wire [1:0] w_n1756_0;
	wire [1:0] w_n1757_0;
	wire [1:0] w_n1758_0;
	wire [1:0] w_n1759_0;
	wire [1:0] w_n1760_0;
	wire [1:0] w_n1767_0;
	wire [1:0] w_n1770_0;
	wire [1:0] w_n1772_0;
	wire [1:0] w_n1775_0;
	wire [1:0] w_n1776_0;
	wire [1:0] w_n1777_0;
	wire [1:0] w_n1780_0;
	wire [1:0] w_n1782_0;
	wire [1:0] w_n1783_0;
	wire [1:0] w_n1784_0;
	wire [1:0] w_n1785_0;
	wire [1:0] w_n1786_0;
	wire [1:0] w_n1793_0;
	wire [1:0] w_n1796_0;
	wire [1:0] w_n1797_0;
	wire [1:0] w_n1798_0;
	wire [1:0] w_n1801_0;
	wire [1:0] w_n1803_0;
	wire [1:0] w_n1804_0;
	wire [1:0] w_n1805_0;
	wire [1:0] w_n1807_0;
	wire [1:0] w_n1810_0;
	wire [1:0] w_n1817_0;
	wire [1:0] w_n1818_0;
	wire w_dff_B_6HCBISXv8_0;
	wire w_dff_B_44QAozby7_0;
	wire w_dff_B_P1ly3IOS3_1;
	wire w_dff_B_ffyvxpWQ4_1;
	wire w_dff_B_AC3vnYzm4_1;
	wire w_dff_B_ZHAJKBDS4_1;
	wire w_dff_B_APaSBmRP6_1;
	wire w_dff_B_JZA2Vr1t8_1;
	wire w_dff_B_2Fxuiwdr8_1;
	wire w_dff_B_3FPIijzO9_1;
	wire w_dff_B_AQulzuKa3_1;
	wire w_dff_B_oRWhJ7ji7_1;
	wire w_dff_B_M3ZkKUfG3_1;
	wire w_dff_B_RzOqDIa92_1;
	wire w_dff_B_GiElhWcy4_1;
	wire w_dff_B_6lI0U1M62_1;
	wire w_dff_B_ZXRMAWNp2_1;
	wire w_dff_B_2h8wkNxg6_1;
	wire w_dff_B_RGGz8Q9K9_1;
	wire w_dff_B_EhBSwQtR6_1;
	wire w_dff_B_Zs2CFwyA2_1;
	wire w_dff_B_osBIpEl50_1;
	wire w_dff_B_p1KD1ZgB9_1;
	wire w_dff_B_b5hrTdYE4_1;
	wire w_dff_B_SPQ4uKhJ9_1;
	wire w_dff_B_2NBSrRwF8_1;
	wire w_dff_B_9MUDVhOy3_1;
	wire w_dff_B_rY0cHKBA7_1;
	wire w_dff_B_zezWY9qf2_1;
	wire w_dff_B_r6ZX9DFu5_1;
	wire w_dff_B_QN7GF7U64_1;
	wire w_dff_B_9tLIY7T60_1;
	wire w_dff_B_47zio2a76_1;
	wire w_dff_B_5y1P21MO3_1;
	wire w_dff_B_UmJB9HqK5_1;
	wire w_dff_B_2gQWOTyL9_1;
	wire w_dff_B_WYZafbxU0_1;
	wire w_dff_B_KLFHqAdj5_1;
	wire w_dff_B_mlpGvvNC4_1;
	wire w_dff_B_WTsUlwhd5_1;
	wire w_dff_B_G3Hg9CTa0_1;
	wire w_dff_B_1rPq1ELK7_1;
	wire w_dff_B_bhhnoe417_1;
	wire w_dff_B_GsgtfQa27_1;
	wire w_dff_B_bOxjIvyv2_1;
	wire w_dff_B_zaENAgzd0_1;
	wire w_dff_B_ZKOk38e58_1;
	wire w_dff_B_ZRCXMTqp0_1;
	wire w_dff_B_K0iH9oca7_1;
	wire w_dff_B_Pn7KYAtS2_1;
	wire w_dff_B_GvS6AMBC3_1;
	wire w_dff_B_Fd6u6okS6_1;
	wire w_dff_B_dHxcuFZv5_1;
	wire w_dff_B_eXbxvIVK6_1;
	wire w_dff_B_73mwioK95_1;
	wire w_dff_B_gkZRwCpI8_1;
	wire w_dff_B_PfcsKGKn9_1;
	wire w_dff_B_wANkVgu04_1;
	wire w_dff_B_SICmrVRM4_1;
	wire w_dff_B_WZmPXDDu0_1;
	wire w_dff_B_weYljKq51_1;
	wire w_dff_B_R6wPNhWs6_1;
	wire w_dff_B_e17I3Z3T3_1;
	wire w_dff_B_OYyNmgz28_1;
	wire w_dff_B_wpT0izjM6_1;
	wire w_dff_B_NDCYA0pf8_1;
	wire w_dff_B_vBSXl2Xc4_1;
	wire w_dff_B_MoG9tggT5_1;
	wire w_dff_B_lER1JFTz8_1;
	wire w_dff_B_v8rZBzxZ9_1;
	wire w_dff_B_rA12eeMp6_1;
	wire w_dff_B_337ugziS5_1;
	wire w_dff_B_GI4gaQTH8_1;
	wire w_dff_B_EsH4uZ5d2_1;
	wire w_dff_B_ionqlwBo7_1;
	wire w_dff_B_1lfLFahR2_1;
	wire w_dff_B_fAbvQ5Lh1_1;
	wire w_dff_B_H1AJWwLO1_1;
	wire w_dff_B_f0bdwSEM7_1;
	wire w_dff_B_gcplfyCN8_1;
	wire w_dff_B_slpYj5Sz2_1;
	wire w_dff_B_WAgK0wi61_1;
	wire w_dff_B_E2fepEw78_1;
	wire w_dff_B_KAaoo34K5_1;
	wire w_dff_B_h0pK2ZN59_1;
	wire w_dff_B_Vq2eGezB9_1;
	wire w_dff_B_eJBhluQ05_1;
	wire w_dff_B_db6P1TxI9_1;
	wire w_dff_B_z7sfF18P0_1;
	wire w_dff_B_r2WbuOzk7_1;
	wire w_dff_B_Vw3ANMGR6_1;
	wire w_dff_B_zIVdlYjI4_1;
	wire w_dff_B_piUAakqS0_1;
	wire w_dff_B_eNk1BIck3_1;
	wire w_dff_B_kZVeK0vh5_1;
	wire w_dff_B_To86uOx91_1;
	wire w_dff_B_hikmQHZC1_1;
	wire w_dff_B_xN1NM4QN6_1;
	wire w_dff_B_4t2gradw0_1;
	wire w_dff_B_Mswpm0uw4_1;
	wire w_dff_B_eJhFKHUS2_1;
	wire w_dff_B_nwUufPEM4_1;
	wire w_dff_B_CwUH8hIa5_1;
	wire w_dff_B_XEwaOo484_1;
	wire w_dff_B_s2M3ZHh94_1;
	wire w_dff_B_fk9C74SQ8_1;
	wire w_dff_B_sGQo05QB3_1;
	wire w_dff_B_jQt9tUQQ3_1;
	wire w_dff_B_75UviKYP7_1;
	wire w_dff_B_fNAOjXgj7_1;
	wire w_dff_B_yOZ9FPuE0_1;
	wire w_dff_B_DcOGLGC31_1;
	wire w_dff_B_Kvv5XlAD3_1;
	wire w_dff_B_RqZ8sDuB7_1;
	wire w_dff_B_6dW1A9a36_1;
	wire w_dff_B_dtvNKsfH7_1;
	wire w_dff_B_fAThyMH45_1;
	wire w_dff_B_J1kGCNu40_1;
	wire w_dff_B_jsxvJsVY9_1;
	wire w_dff_B_2JFBsbtW8_1;
	wire w_dff_B_lUcAy4X63_1;
	wire w_dff_B_pNShPGpz0_1;
	wire w_dff_B_0uDtAaaq6_1;
	wire w_dff_B_1bVWCKcC6_1;
	wire w_dff_B_NJIlRyTE6_1;
	wire w_dff_B_jwipN2CY1_1;
	wire w_dff_B_2kZXeCC49_1;
	wire w_dff_B_Aw8akPT04_1;
	wire w_dff_B_u3x12r8n9_1;
	wire w_dff_B_gouTXm9C8_1;
	wire w_dff_B_LOadvB4t1_1;
	wire w_dff_B_kWE5Tpjh0_1;
	wire w_dff_B_XAOBa3Mx5_1;
	wire w_dff_B_c1zz1fwu5_1;
	wire w_dff_B_NxYGl2uN6_1;
	wire w_dff_B_1L2ItabO4_1;
	wire w_dff_B_BafcEK5p1_1;
	wire w_dff_B_5BPUIjys6_1;
	wire w_dff_B_E8SJa8mo6_1;
	wire w_dff_B_vrV1saZx8_1;
	wire w_dff_B_8G05LpYR8_1;
	wire w_dff_B_VI28tZaS1_1;
	wire w_dff_B_DXE4c9xI2_1;
	wire w_dff_B_3Xfoueyt3_1;
	wire w_dff_B_YYRw8vvW0_1;
	wire w_dff_B_JUwEIWLz9_1;
	wire w_dff_B_5ZjePXzK5_1;
	wire w_dff_B_RpRR36822_1;
	wire w_dff_B_kW615ZDf3_1;
	wire w_dff_B_25PnaRh24_1;
	wire w_dff_B_OhLTnKcC2_1;
	wire w_dff_B_MhejmIW43_1;
	wire w_dff_B_WpY32sTM7_1;
	wire w_dff_B_ywyILbZb1_1;
	wire w_dff_B_CjdLPUiM5_1;
	wire w_dff_B_fPk6YKlx7_1;
	wire w_dff_B_3lifHEZd4_1;
	wire w_dff_B_z7vHNlC37_1;
	wire w_dff_B_YCOEgNde7_1;
	wire w_dff_B_q31oRVu59_1;
	wire w_dff_B_54U1Ebai6_1;
	wire w_dff_B_WgNOPtbR7_1;
	wire w_dff_B_pwhXadAr9_1;
	wire w_dff_B_D1uHqIK13_1;
	wire w_dff_B_UQuUMfDF6_1;
	wire w_dff_B_VHudfPek1_1;
	wire w_dff_B_FA28I9X16_1;
	wire w_dff_B_lustcrdz8_1;
	wire w_dff_B_B1sULxai5_1;
	wire w_dff_B_9NSKS4iH7_1;
	wire w_dff_B_BTC1j4ci8_1;
	wire w_dff_B_T4f05lYe2_1;
	wire w_dff_B_J7vC8etz5_1;
	wire w_dff_B_yfadh71H6_1;
	wire w_dff_B_lCvek3820_1;
	wire w_dff_B_Cb2FTDkZ0_1;
	wire w_dff_B_XDpT0z4L9_1;
	wire w_dff_B_ZWq9mVjX5_1;
	wire w_dff_B_ojxTvVzN8_1;
	wire w_dff_B_2n9rX5NF0_1;
	wire w_dff_B_xtAfkHVQ0_1;
	wire w_dff_B_d1E1EsaN5_1;
	wire w_dff_B_2xbHyuk16_1;
	wire w_dff_B_MywtW5J48_1;
	wire w_dff_B_zjo25QH17_1;
	wire w_dff_B_vjtwDPqG8_1;
	wire w_dff_B_o941zw169_1;
	wire w_dff_B_kZkDyc0g2_1;
	wire w_dff_B_FkzRXiDH9_1;
	wire w_dff_B_enIigK9G1_1;
	wire w_dff_B_DN4nkYGH0_1;
	wire w_dff_B_daZPsIaI8_1;
	wire w_dff_B_tYYbO5dn3_1;
	wire w_dff_B_uMpWvmzj5_1;
	wire w_dff_B_Zp53MIf52_1;
	wire w_dff_B_97zjeKu91_1;
	wire w_dff_B_Ek2XAlay5_1;
	wire w_dff_B_qD161yEY9_1;
	wire w_dff_B_A3v1x0ib6_1;
	wire w_dff_B_tBFU9LYF6_1;
	wire w_dff_B_em7tHQAn7_1;
	wire w_dff_B_yiVf1GD43_1;
	wire w_dff_B_UVEjgrBr8_1;
	wire w_dff_B_aEMieyYt2_1;
	wire w_dff_B_jZFb2SLn7_1;
	wire w_dff_B_rGb6IK2a2_1;
	wire w_dff_B_L1IzeLEC7_1;
	wire w_dff_B_dz67p68o8_1;
	wire w_dff_B_PD8HBJ9E5_1;
	wire w_dff_B_CP34vhPg4_1;
	wire w_dff_B_hYMNgODB1_1;
	wire w_dff_B_OETIUeAI6_1;
	wire w_dff_B_odBswDdc9_1;
	wire w_dff_B_lCDIlywy8_1;
	wire w_dff_B_0uBAdJ4d8_1;
	wire w_dff_B_C9He6REg3_1;
	wire w_dff_B_jhNC7s6L3_1;
	wire w_dff_B_yP7pFhl94_1;
	wire w_dff_B_AnNMTJn20_1;
	wire w_dff_B_LVkMcXWe4_1;
	wire w_dff_B_hOB0AtOD9_1;
	wire w_dff_B_Tk7wV1x59_1;
	wire w_dff_B_utRrxLn92_1;
	wire w_dff_B_Y8sUVSjt0_1;
	wire w_dff_B_fdES0JQs8_1;
	wire w_dff_B_cEXRX9cm0_1;
	wire w_dff_B_fakX5dCT6_1;
	wire w_dff_B_gr5uCgK71_1;
	wire w_dff_B_p5swbb7p8_1;
	wire w_dff_B_mrSl81Yl6_1;
	wire w_dff_B_QXICfYFg5_1;
	wire w_dff_B_gptQrV040_1;
	wire w_dff_B_4jjwyFOG0_1;
	wire w_dff_B_zfzNnqCc6_1;
	wire w_dff_B_qWMQWpFq9_1;
	wire w_dff_B_44qIIvi99_1;
	wire w_dff_B_lo1K324g8_1;
	wire w_dff_B_gJv09Qok4_1;
	wire w_dff_B_S1aAAp0O6_1;
	wire w_dff_B_u62KfPAb1_1;
	wire w_dff_B_2N0GWwYC9_1;
	wire w_dff_B_vx5kiSt78_1;
	wire w_dff_B_gvNJmRDX9_1;
	wire w_dff_B_OueJZUUO7_1;
	wire w_dff_B_kBVGO1xB8_1;
	wire w_dff_B_I66AOxMl8_1;
	wire w_dff_B_2pKtVac62_1;
	wire w_dff_B_yVQkM1H66_1;
	wire w_dff_B_to30z33n7_1;
	wire w_dff_B_FPhJtWp79_1;
	wire w_dff_B_lN9gcYhF1_1;
	wire w_dff_B_y2yx8tk69_1;
	wire w_dff_B_1z8N5QVY8_1;
	wire w_dff_B_bKVskMcs8_1;
	wire w_dff_B_pI24JtGM4_0;
	wire w_dff_B_L0lJCq0a1_1;
	wire w_dff_B_90IjmZ2U2_1;
	wire w_dff_B_zjc0t6o19_1;
	wire w_dff_B_kZYiTLjE5_1;
	wire w_dff_B_hiB8ofTa5_1;
	wire w_dff_B_AIOufWfd4_1;
	wire w_dff_B_SYkn1LZE6_1;
	wire w_dff_B_IqTVostd0_0;
	wire w_dff_B_K2FZU5Ca1_0;
	wire w_dff_B_1PHCjzAR5_0;
	wire w_dff_B_jDBZ49te8_0;
	wire w_dff_B_Hud6zxaB7_0;
	wire w_dff_A_W0ePeiK66_0;
	wire w_dff_A_MFPSpaIB9_0;
	wire w_dff_A_OBoyWszB3_0;
	wire w_dff_A_goyEREVc2_0;
	wire w_dff_A_xBmmHKr30_0;
	wire w_dff_A_Xwkf2BHt1_0;
	wire w_dff_B_xx6l7qui3_1;
	wire w_dff_B_mn4rCjzz0_1;
	wire w_dff_B_lE7QRb345_2;
	wire w_dff_B_8pCulNH83_2;
	wire w_dff_B_Qf6y5UA72_2;
	wire w_dff_B_ObuV6XP09_2;
	wire w_dff_B_u7Woywot6_2;
	wire w_dff_B_88T758w23_2;
	wire w_dff_B_zNi7oP3q8_2;
	wire w_dff_B_iYnjBo3z1_2;
	wire w_dff_B_yl7rMzmQ8_2;
	wire w_dff_B_AirbCeqY3_2;
	wire w_dff_B_PX3Ryoyl5_2;
	wire w_dff_B_OlxbPXNB9_2;
	wire w_dff_B_eiOJyZqL6_2;
	wire w_dff_B_jVuwhZvT8_2;
	wire w_dff_B_GL3slo7Z1_2;
	wire w_dff_B_1fIBqJmy8_2;
	wire w_dff_B_ZSRgh43m4_2;
	wire w_dff_B_RnSgaOmr8_2;
	wire w_dff_B_wgHEkmyy6_2;
	wire w_dff_B_DGdKhsWa1_2;
	wire w_dff_B_EuGidYqY6_2;
	wire w_dff_B_FYFisWGb9_2;
	wire w_dff_B_Yujf99G73_2;
	wire w_dff_B_VQizus1p1_2;
	wire w_dff_B_qUkau1RW4_2;
	wire w_dff_B_SjNiWd1k0_2;
	wire w_dff_B_mSM1Xl9R5_2;
	wire w_dff_B_hM7KeAsn4_2;
	wire w_dff_B_M9VDviPH7_2;
	wire w_dff_B_waMO7DUW5_2;
	wire w_dff_B_IleYBp5n1_2;
	wire w_dff_B_1KgAOyTA0_2;
	wire w_dff_B_VIDOZ50d4_2;
	wire w_dff_B_X62xnjUP3_2;
	wire w_dff_B_LZkHANrP5_2;
	wire w_dff_B_rH9JTWna4_2;
	wire w_dff_B_NPqX5pqK9_2;
	wire w_dff_B_iLKLZ3HG3_2;
	wire w_dff_B_jGz6bc6R3_2;
	wire w_dff_B_FSxwYpwN8_2;
	wire w_dff_B_faF78IKG6_2;
	wire w_dff_B_ZJgFeNct6_2;
	wire w_dff_B_CaMxzjt13_2;
	wire w_dff_B_UaMFD9u46_1;
	wire w_dff_B_2kjpgPmk6_1;
	wire w_dff_B_5LWtGzuY8_1;
	wire w_dff_B_aJP7bq8n8_1;
	wire w_dff_B_LWJ4q85k1_1;
	wire w_dff_B_tZ589fHD3_0;
	wire w_dff_B_jkygkTSI3_0;
	wire w_dff_B_GKJ3ibl99_0;
	wire w_dff_B_S4ltgIP69_0;
	wire w_dff_A_xuiwnLhZ9_1;
	wire w_dff_A_kKEoqttp9_1;
	wire w_dff_A_rBeQwzzF2_1;
	wire w_dff_A_J7NxZJ3L7_1;
	wire w_dff_A_7HgF2Ebz3_1;
	wire w_dff_B_zeANGTQO9_1;
	wire w_dff_B_W2fm52nh9_1;
	wire w_dff_B_tjxn3Cha9_1;
	wire w_dff_B_xy2ZCBsW6_1;
	wire w_dff_B_SeIcI13K2_1;
	wire w_dff_B_Bg2e2mZh0_0;
	wire w_dff_B_9LfwhznL4_0;
	wire w_dff_B_HjZbioiq5_0;
	wire w_dff_B_UKeQvCg87_0;
	wire w_dff_A_UmyjqEiB3_1;
	wire w_dff_A_g2W2EC9J8_1;
	wire w_dff_A_7nZHykkt0_1;
	wire w_dff_A_iKTDXahH9_1;
	wire w_dff_A_dLavTA406_1;
	wire w_dff_B_opUNiU9e4_1;
	wire w_dff_B_FXWqG8P88_1;
	wire w_dff_B_aTNh3bMG2_1;
	wire w_dff_B_9K7NBD5C3_1;
	wire w_dff_B_LBz8FDdd7_1;
	wire w_dff_B_lxBwEA4n3_0;
	wire w_dff_B_65s5OWsu0_0;
	wire w_dff_B_rYAiRxjA9_0;
	wire w_dff_B_5ubhJ4Ul9_0;
	wire w_dff_A_f238AYfa5_1;
	wire w_dff_A_E5jJywQ17_1;
	wire w_dff_A_6DUvxiW19_1;
	wire w_dff_A_32ZOwtlv4_1;
	wire w_dff_A_wwb1llDO5_1;
	wire w_dff_B_QVKlm6nG3_1;
	wire w_dff_B_2aPVKMdH7_1;
	wire w_dff_B_3LlaYMpX1_1;
	wire w_dff_B_xgLbS7ef2_1;
	wire w_dff_B_v9bnab3R2_1;
	wire w_dff_B_dsWpZ4tF8_0;
	wire w_dff_B_sotNSENx5_0;
	wire w_dff_B_mxLQyMKv5_0;
	wire w_dff_B_lculz7TR9_0;
	wire w_dff_A_haUmetS19_1;
	wire w_dff_A_9g1Wf2nE0_1;
	wire w_dff_A_9HZ3DGBc6_1;
	wire w_dff_A_GQ9guesq5_1;
	wire w_dff_A_nw0zklZx2_1;
	wire w_dff_B_7l0Me6jS2_1;
	wire w_dff_B_0sDZLPxK5_1;
	wire w_dff_B_oYxPY6s27_1;
	wire w_dff_B_dgNyMpz47_1;
	wire w_dff_B_3YCoDQeY1_1;
	wire w_dff_B_rMHj3k131_0;
	wire w_dff_B_fqTUIr7f6_0;
	wire w_dff_B_dN7mMsn83_0;
	wire w_dff_A_HmaB0Zgm4_1;
	wire w_dff_A_Ml8at2Oa9_1;
	wire w_dff_A_zEYZS2gD6_1;
	wire w_dff_A_ixcFa8oL9_1;
	wire w_dff_B_GG62YzVH8_1;
	wire w_dff_B_rGI26zXL7_1;
	wire w_dff_B_vCwvBcrj8_1;
	wire w_dff_B_8QhDajyx7_1;
	wire w_dff_B_EJmoYI6o3_0;
	wire w_dff_B_f4Eih3xY4_0;
	wire w_dff_A_nLDtfdqs7_1;
	wire w_dff_A_KeQP5j814_1;
	wire w_dff_A_my0cukNQ9_1;
	wire w_dff_B_lLTCaoQP0_1;
	wire w_dff_B_m9I7jFRb9_1;
	wire w_dff_B_qI9DitWk4_1;
	wire w_dff_B_UekR6NNa3_1;
	wire w_dff_B_q6FgAOK44_0;
	wire w_dff_B_FwpMwxfk6_0;
	wire w_dff_A_GRKxZznQ3_1;
	wire w_dff_A_BxhsF5cW3_1;
	wire w_dff_A_2W8eSvNS9_1;
	wire w_dff_B_lojryFKB0_1;
	wire w_dff_B_aJt4jwp71_1;
	wire w_dff_B_ErnfkFhA3_1;
	wire w_dff_B_AIG6bJtq8_1;
	wire w_dff_B_t5NPkjVm4_0;
	wire w_dff_B_xA4A4SQ38_0;
	wire w_dff_A_MhEnWH1e4_1;
	wire w_dff_A_OjP6DQj17_1;
	wire w_dff_A_Q4KL71pY0_1;
	wire w_dff_B_JhwNLh4z5_1;
	wire w_dff_B_MNJcPB5i0_1;
	wire w_dff_B_GL8yvwSr3_1;
	wire w_dff_B_zEQtFjHc9_1;
	wire w_dff_B_L7vuoqVx1_0;
	wire w_dff_B_UJiY7Bnj3_0;
	wire w_dff_A_9zNi1lLP1_1;
	wire w_dff_A_AYMSnguH9_1;
	wire w_dff_A_1RrEBp7h4_1;
	wire w_dff_B_czyWzkBd8_1;
	wire w_dff_B_clKURfb93_1;
	wire w_dff_B_vE7MgVrH1_1;
	wire w_dff_B_NAMTOoqD0_1;
	wire w_dff_B_s2uwMy4s4_0;
	wire w_dff_B_w2l7Nkfj6_0;
	wire w_dff_A_6S9ZFhC44_1;
	wire w_dff_A_ddKYqWmG2_1;
	wire w_dff_A_cFG0Ia5Z3_1;
	wire w_dff_B_Hqoe6YU48_1;
	wire w_dff_B_WSwqW1o59_1;
	wire w_dff_B_n6bnUqnb4_1;
	wire w_dff_A_uVhFRkNE4_0;
	wire w_dff_A_SX75LK7v5_0;
	wire w_dff_B_NpeQjmGC5_1;
	wire w_dff_A_BPfeRMEG5_0;
	wire w_dff_B_8GXt3znx8_1;
	wire w_dff_A_eim6TkIP3_0;
	wire w_dff_B_YNvCsceP4_2;
	wire w_dff_B_Xia3DPRR8_1;
	wire w_dff_A_662e2IZt3_0;
	wire w_dff_A_nYbpCc9b3_0;
	wire w_dff_A_ThMdp57M7_0;
	wire w_dff_A_kgFBWi1H8_0;
	wire w_dff_A_J2FjpTxz8_0;
	wire w_dff_A_nJSXpeTJ9_0;
	wire w_dff_A_f2sPAGvk7_0;
	wire w_dff_A_7r92TQdh3_0;
	wire w_dff_A_efvqtBPX6_0;
	wire w_dff_A_NpHji1wM6_0;
	wire w_dff_A_jkyacbFs5_0;
	wire w_dff_A_4aYeIp7H0_0;
	wire w_dff_A_Q1nZT9NW0_0;
	wire w_dff_A_2LBktEPd4_0;
	wire w_dff_A_RbA0scCG7_0;
	wire w_dff_A_LP7iEK6k7_0;
	wire w_dff_A_KMsGdlAA4_0;
	wire w_dff_A_jwKx4BaT1_0;
	wire w_dff_A_NesHmd2r2_0;
	wire w_dff_A_eSRf35sg1_0;
	wire w_dff_A_mZA5N4Dx4_0;
	wire w_dff_A_FaVWmzpk7_0;
	wire w_dff_A_l2grCAkI0_0;
	wire w_dff_A_vWvCWpLx2_0;
	wire w_dff_A_9TQiNsuW5_0;
	wire w_dff_A_WzVtAAyB4_0;
	wire w_dff_A_xWLrdaQV6_0;
	wire w_dff_A_S3D6GCMz9_0;
	wire w_dff_A_KGuhiddx0_0;
	wire w_dff_A_NowR9RrP5_0;
	wire w_dff_A_yK1ep4SU1_0;
	wire w_dff_A_FlWyKGHC0_0;
	wire w_dff_A_g7twgXVv7_0;
	wire w_dff_A_SHL8gzUL6_0;
	wire w_dff_A_r2CxQq4M1_1;
	wire w_dff_A_LjvnUsz49_0;
	wire w_dff_A_79GnhfdT0_0;
	wire w_dff_A_pf89cse13_0;
	wire w_dff_A_apu5ctas8_0;
	wire w_dff_A_Y44ODO1F3_0;
	wire w_dff_A_lqfcvZwT1_0;
	wire w_dff_A_ap2fhwR85_0;
	wire w_dff_A_NCqsT08l4_0;
	wire w_dff_A_X7MAs05s4_0;
	wire w_dff_A_vAceU8wQ5_0;
	wire w_dff_A_FuBDexXD0_0;
	wire w_dff_A_f77i4ZKS3_0;
	wire w_dff_A_Vkb2O4x28_0;
	wire w_dff_A_DoHLIW5U8_0;
	wire w_dff_A_EOJQe4B41_0;
	wire w_dff_A_xDlzd7Rw4_0;
	wire w_dff_A_eb5Z8V4x8_0;
	wire w_dff_A_HSdjzxSB4_0;
	wire w_dff_A_jxda1fWA3_0;
	wire w_dff_A_9C5Jn2vo2_0;
	wire w_dff_A_qsUQrKts7_0;
	wire w_dff_A_gocJm6ip5_0;
	wire w_dff_A_0UDK4Hgn9_0;
	wire w_dff_A_rzs4JHKQ7_0;
	wire w_dff_A_zU3szE2g4_0;
	wire w_dff_A_r3dRZP5F8_0;
	wire w_dff_A_XvnQLgZ65_0;
	wire w_dff_A_BGabRieq2_0;
	wire w_dff_A_u7MVywNI6_0;
	wire w_dff_A_J7GUCHDN2_0;
	wire w_dff_A_WWGZUu9N7_0;
	wire w_dff_A_4rh7ihgJ1_0;
	wire w_dff_B_fl0c5mED1_1;
	wire w_dff_B_EroCWDUZ0_1;
	wire w_dff_B_BcNIiExZ7_1;
	wire w_dff_B_FPU74JMr8_1;
	wire w_dff_B_LK183Sg95_1;
	wire w_dff_B_ihwmrTxG4_1;
	wire w_dff_B_9XK5f75c4_1;
	wire w_dff_B_azC47Q5P6_1;
	wire w_dff_B_vbp8zN347_1;
	wire w_dff_B_jufl5Zgt6_1;
	wire w_dff_B_o3X9hQLN0_1;
	wire w_dff_B_dkYp4EWn9_1;
	wire w_dff_B_tOd8JLdK9_1;
	wire w_dff_B_hVvAXGU58_1;
	wire w_dff_B_tp0VQJV27_1;
	wire w_dff_B_9WzvPrhm1_1;
	wire w_dff_B_L91TH4AG9_1;
	wire w_dff_B_1M9VXOi20_1;
	wire w_dff_B_i9uMggk96_1;
	wire w_dff_B_WkFeOUrA0_1;
	wire w_dff_B_xhaK2JqE9_1;
	wire w_dff_B_n4TMqiaz9_1;
	wire w_dff_B_T3L0LJUr4_1;
	wire w_dff_B_Cjp3A2X53_1;
	wire w_dff_B_Ai2Lm1r26_1;
	wire w_dff_B_OAZclFQB9_1;
	wire w_dff_B_moMqFGDf9_1;
	wire w_dff_B_aHmtZ6tl5_1;
	wire w_dff_B_Xr8BrdpT9_1;
	wire w_dff_A_u0s3Zbqb3_0;
	wire w_dff_A_DhJPKj8z5_0;
	wire w_dff_A_0NuIA5fv0_0;
	wire w_dff_A_aP1WtKMP3_0;
	wire w_dff_A_TfCsFiU43_0;
	wire w_dff_A_lrgq5xpY5_0;
	wire w_dff_A_Fmmh8k6N9_0;
	wire w_dff_A_BIpxdEPV2_0;
	wire w_dff_A_pQMKzbRF3_0;
	wire w_dff_A_Aolfnmco6_0;
	wire w_dff_A_xVRQm6lv1_0;
	wire w_dff_A_f2ZIWKq99_0;
	wire w_dff_A_ITW5vLeN9_0;
	wire w_dff_A_WlwAB7hE0_0;
	wire w_dff_A_8NxqBm351_0;
	wire w_dff_A_eryoXjcz8_0;
	wire w_dff_A_Z9yh2W5N9_0;
	wire w_dff_A_lk1UE25t6_0;
	wire w_dff_A_AXCjBpp53_0;
	wire w_dff_A_U4z4fEaq7_0;
	wire w_dff_A_rtaGv1At5_0;
	wire w_dff_A_q5UBzoSI8_0;
	wire w_dff_A_74bJ42Px2_0;
	wire w_dff_A_cKe8MsmW7_0;
	wire w_dff_A_YiKKVe339_0;
	wire w_dff_A_YlLS9Huu6_0;
	wire w_dff_A_UdzPKHV37_0;
	wire w_dff_A_1j8JjMbh9_0;
	wire w_dff_A_6jxhMHGT2_0;
	wire w_dff_A_VEaKGW435_0;
	wire w_dff_A_RK6NV3yY4_0;
	wire w_dff_B_yyVOwNSn6_1;
	wire w_dff_B_kDYN1VUs6_1;
	wire w_dff_B_pj3Ag8u10_1;
	wire w_dff_B_kuKkryOB8_1;
	wire w_dff_B_wV6ZTMw41_1;
	wire w_dff_B_zAKn2UZ08_1;
	wire w_dff_B_njclK8zl3_1;
	wire w_dff_B_vPpFkMWL7_1;
	wire w_dff_B_dxTpz6Ld8_1;
	wire w_dff_B_1ZlObyMt6_1;
	wire w_dff_B_pq7aIwPR5_1;
	wire w_dff_B_sfZo5COr3_1;
	wire w_dff_B_tPDdOh0K9_1;
	wire w_dff_B_xOif8gcl1_1;
	wire w_dff_B_ubcRyYBL4_1;
	wire w_dff_B_dxrBSLmP4_1;
	wire w_dff_B_nxT1jgfo7_1;
	wire w_dff_B_neV8O9dC9_1;
	wire w_dff_B_7UaYYAbM1_1;
	wire w_dff_B_Qaf57BRl0_1;
	wire w_dff_B_18iTE7CW6_1;
	wire w_dff_B_w28BwwaZ8_1;
	wire w_dff_B_k6QZNmAk0_1;
	wire w_dff_B_rFT5RGUN6_1;
	wire w_dff_B_DBuZFplD7_1;
	wire w_dff_B_JTC0kpu73_1;
	wire w_dff_B_b2d0OJvg0_1;
	wire w_dff_A_wpS1r5Ve3_0;
	wire w_dff_A_YA8c7Vsj6_0;
	wire w_dff_A_6VICeRBW3_0;
	wire w_dff_A_Pzz4ffo91_0;
	wire w_dff_A_6LsxZDxU1_0;
	wire w_dff_A_mstkAnUV8_0;
	wire w_dff_A_dvUsAZYt7_0;
	wire w_dff_A_apH9xc515_0;
	wire w_dff_A_k5sUWt6F5_0;
	wire w_dff_A_ZLA3LvBy4_0;
	wire w_dff_A_LJdIBqOY4_0;
	wire w_dff_A_atpe8yZE1_0;
	wire w_dff_A_nJ1njDy75_0;
	wire w_dff_A_XInLPycQ7_0;
	wire w_dff_A_lt8uivqi3_0;
	wire w_dff_A_8Tm8oo6L4_0;
	wire w_dff_A_wRK892fu0_0;
	wire w_dff_A_rmczvSi92_0;
	wire w_dff_A_4byYXUiP1_0;
	wire w_dff_A_eX2ryzXN3_0;
	wire w_dff_A_MJsbTHvp5_0;
	wire w_dff_A_8nXUk5064_0;
	wire w_dff_A_WALeyVol8_0;
	wire w_dff_A_gUgtPafd3_0;
	wire w_dff_A_mxvlQutG6_0;
	wire w_dff_A_7230e3rg5_0;
	wire w_dff_A_44f0VQ760_0;
	wire w_dff_A_XvAdRIwp2_0;
	wire w_dff_A_heUPJXR54_0;
	wire w_dff_B_lwbqDVIQ6_1;
	wire w_dff_B_KFB0YdQh2_1;
	wire w_dff_B_25UWo6Kx6_1;
	wire w_dff_B_x6Xp0fhs8_1;
	wire w_dff_B_FwpSVmFo7_1;
	wire w_dff_B_swzC9u0u5_1;
	wire w_dff_B_UmpXJIOF1_1;
	wire w_dff_B_LE85dAEu0_1;
	wire w_dff_B_k8Wmwwen9_1;
	wire w_dff_B_8foNXss18_1;
	wire w_dff_B_5zma2OI19_1;
	wire w_dff_B_G3W7TjME8_1;
	wire w_dff_B_9gqH5NdN3_1;
	wire w_dff_B_J2ZNqNcs7_1;
	wire w_dff_B_PK1mKeB32_1;
	wire w_dff_B_OCowzZ429_1;
	wire w_dff_B_JtjJyPBd8_1;
	wire w_dff_B_17PlxHih2_1;
	wire w_dff_B_8Pc8qrVl3_1;
	wire w_dff_B_cUQbM1Lk9_1;
	wire w_dff_B_02DVclHt9_1;
	wire w_dff_B_efRyBIxh2_1;
	wire w_dff_B_8DI3KBPB1_1;
	wire w_dff_B_xosNsz7v5_1;
	wire w_dff_B_fSWVXiTU0_1;
	wire w_dff_A_XGY45YLI0_0;
	wire w_dff_A_En2GioGH4_0;
	wire w_dff_A_GwkOOmRj8_0;
	wire w_dff_A_ae0vzBCp7_0;
	wire w_dff_A_k3lXcdZK0_0;
	wire w_dff_A_lw0rnrfI6_0;
	wire w_dff_A_D5XXFsMe3_0;
	wire w_dff_A_YQ1GHwYF8_0;
	wire w_dff_A_F2M2hjAQ7_0;
	wire w_dff_A_0t9o09RF1_0;
	wire w_dff_A_cqfiSJAM6_0;
	wire w_dff_A_eJSQsWRa4_0;
	wire w_dff_A_c79lqtLe4_0;
	wire w_dff_A_pobWB3Xf6_0;
	wire w_dff_A_rjG6rSI43_0;
	wire w_dff_A_ZFU39aD09_0;
	wire w_dff_A_zLwuAHox7_0;
	wire w_dff_A_7o1RRmWI5_0;
	wire w_dff_A_5ncj4DcK0_0;
	wire w_dff_A_SosMuBux0_0;
	wire w_dff_A_BxPeyYXQ6_0;
	wire w_dff_A_daNuyowd4_0;
	wire w_dff_A_1AsRAIib1_0;
	wire w_dff_A_c8Fuw6xd7_0;
	wire w_dff_A_yzoKD03O9_0;
	wire w_dff_A_m9b5JjKC8_0;
	wire w_dff_A_oHHeRJzx3_0;
	wire w_dff_B_autOpJMY4_1;
	wire w_dff_B_iwAisoDV7_1;
	wire w_dff_B_1UHCkcWA5_1;
	wire w_dff_B_U8bbVaYg7_1;
	wire w_dff_B_5wIgPplJ8_1;
	wire w_dff_B_EgztDzRY5_1;
	wire w_dff_B_rLWf9Khn9_1;
	wire w_dff_B_bioYfxHb3_1;
	wire w_dff_B_Y8J8XSz76_1;
	wire w_dff_B_30qpmITL7_1;
	wire w_dff_B_4uRb8raq6_1;
	wire w_dff_B_pLGfKK440_1;
	wire w_dff_B_GiH5w1Fx3_1;
	wire w_dff_B_iMZeQKvo0_1;
	wire w_dff_B_oWPvb8HD3_1;
	wire w_dff_B_2eJzP2Ax9_1;
	wire w_dff_B_dcjT6elr3_1;
	wire w_dff_B_lsJY1KAu1_1;
	wire w_dff_B_L9tQ05x56_1;
	wire w_dff_B_eOqGNY3X9_1;
	wire w_dff_B_E986NeAS8_1;
	wire w_dff_B_hwTqp9gH6_1;
	wire w_dff_B_ertSK6Qe6_1;
	wire w_dff_A_u8VsDPPC5_0;
	wire w_dff_A_ZXw6WQGz4_0;
	wire w_dff_A_VOZr7sxY7_0;
	wire w_dff_A_HBU1kEVA5_0;
	wire w_dff_A_3bS3gjp98_0;
	wire w_dff_A_1OXc49AO6_0;
	wire w_dff_A_hoFuVvjh6_0;
	wire w_dff_A_DOmHUwHf4_0;
	wire w_dff_A_jw2VlL2N9_0;
	wire w_dff_A_Gb0DUAz90_0;
	wire w_dff_A_gSuGt7599_0;
	wire w_dff_A_dmdBv8N27_0;
	wire w_dff_A_f9nTi06l8_0;
	wire w_dff_A_YlYbNnYc0_0;
	wire w_dff_A_HLjgf71D3_0;
	wire w_dff_A_kUyvyLAY3_0;
	wire w_dff_A_omMqnCze0_0;
	wire w_dff_A_2djNMAqW6_0;
	wire w_dff_A_q111pifi0_0;
	wire w_dff_A_VEnxGjTL4_0;
	wire w_dff_A_62OX3wJD5_0;
	wire w_dff_A_d1ul7Iot6_0;
	wire w_dff_A_jzHLlFiT5_0;
	wire w_dff_A_S2BPgjId0_0;
	wire w_dff_A_eEk6Vttx5_0;
	wire w_dff_B_ZBaLs8Xt5_1;
	wire w_dff_B_5OhO8aqw2_1;
	wire w_dff_B_uKNdESmR9_1;
	wire w_dff_B_a2bjLhg20_1;
	wire w_dff_B_mUUNlJ0V1_1;
	wire w_dff_B_xWGuQY4H3_1;
	wire w_dff_B_eFuyN7178_1;
	wire w_dff_B_LzCfgZce0_1;
	wire w_dff_B_klKHjjHP8_1;
	wire w_dff_B_q5cT0LaK9_1;
	wire w_dff_B_jLIAHJEB4_1;
	wire w_dff_B_40Rni9Ms8_1;
	wire w_dff_B_7sjyTkwd0_1;
	wire w_dff_B_I9lAXt8m1_1;
	wire w_dff_B_tF5ARYye3_1;
	wire w_dff_B_cuCAjS7Y9_1;
	wire w_dff_B_TTquGkNp2_1;
	wire w_dff_B_XurUm3wt5_1;
	wire w_dff_B_BdRZzR443_1;
	wire w_dff_B_lcf8fmva2_1;
	wire w_dff_B_VJscNDj46_1;
	wire w_dff_A_UPGQO3ku6_0;
	wire w_dff_B_YcJUKzoX3_2;
	wire w_dff_B_BgOGxSfx7_2;
	wire w_dff_B_WvtuT2Pi5_2;
	wire w_dff_A_ODBUwlKM2_0;
	wire w_dff_A_kuRBZquW6_0;
	wire w_dff_A_RnAKYu0I5_0;
	wire w_dff_A_vQIWDP8O7_0;
	wire w_dff_A_88dQwK2C2_0;
	wire w_dff_A_O2Z6KUF80_0;
	wire w_dff_A_zSQSs7UD4_0;
	wire w_dff_A_X7woO4tv3_0;
	wire w_dff_A_H463M3154_0;
	wire w_dff_A_EvwQHDzA9_0;
	wire w_dff_A_oRhAsIip2_0;
	wire w_dff_A_zvqnwvqG4_0;
	wire w_dff_A_ZxMd2Zpg2_0;
	wire w_dff_A_IybbEaTi6_0;
	wire w_dff_A_2mo7jEbm9_0;
	wire w_dff_A_W3pAHDV28_0;
	wire w_dff_A_wYQWRqgR0_0;
	wire w_dff_A_Vf3Vxb8B9_0;
	wire w_dff_A_hreXLba73_0;
	wire w_dff_B_ppvBdmk69_1;
	wire w_dff_B_wGq0fBei3_1;
	wire w_dff_B_52mRj8BX4_1;
	wire w_dff_B_EyZmbKQn1_1;
	wire w_dff_B_Ty4v1lhC6_1;
	wire w_dff_B_X6UfdxlN6_1;
	wire w_dff_B_OPTo0SHl1_1;
	wire w_dff_B_nJElXwyf0_1;
	wire w_dff_B_oAtWTKTZ8_1;
	wire w_dff_B_fDUpqPth8_1;
	wire w_dff_B_PWiVRgRp6_1;
	wire w_dff_B_FfGhO3UM8_1;
	wire w_dff_B_Kx8lPyYI3_1;
	wire w_dff_B_BvgUhpIb0_1;
	wire w_dff_B_nRx4sBmY5_1;
	wire w_dff_B_J2iYhzFI2_1;
	wire w_dff_A_tA5PPiBy4_0;
	wire w_dff_A_unjFYYcQ8_0;
	wire w_dff_A_nVzotmll3_0;
	wire w_dff_A_SMECIaB48_0;
	wire w_dff_A_yOxCL8S28_0;
	wire w_dff_A_z3DnaPuo7_0;
	wire w_dff_A_2ipbUAOX1_0;
	wire w_dff_A_NyWKRBh69_0;
	wire w_dff_A_puRTLCSS5_0;
	wire w_dff_A_pvox5kaB9_0;
	wire w_dff_A_2WKantat9_0;
	wire w_dff_A_AnYNbJGs3_0;
	wire w_dff_A_01AAbO2o1_0;
	wire w_dff_A_N8kmsmrQ9_0;
	wire w_dff_A_taOp7IB92_0;
	wire w_dff_A_nkWJqKJO7_0;
	wire w_dff_A_xtxI1w8u9_0;
	wire w_dff_A_a0Q0MiLY4_0;
	wire w_dff_B_wZLPf5rD3_1;
	wire w_dff_B_VgA1fXqw7_1;
	wire w_dff_B_6NwTz5RD3_1;
	wire w_dff_B_R5ILRlRx9_1;
	wire w_dff_B_zyrAS5QZ4_1;
	wire w_dff_B_5RJaNZTX0_1;
	wire w_dff_B_bcV2UJjf4_1;
	wire w_dff_B_tLbFtjrV9_1;
	wire w_dff_B_Nncg7cwm4_1;
	wire w_dff_B_AdnQVUDQ9_1;
	wire w_dff_B_FJjUJS5k8_1;
	wire w_dff_B_LRnOdHqb5_1;
	wire w_dff_B_yMMzxuTT9_1;
	wire w_dff_B_hp4iNseb0_1;
	wire w_dff_A_GJdiBsWB7_0;
	wire w_dff_A_5EXzJLuH3_0;
	wire w_dff_A_22WQMr4n0_0;
	wire w_dff_A_JaudKe7w0_0;
	wire w_dff_A_Rp14fa114_0;
	wire w_dff_A_dizxUtmd9_0;
	wire w_dff_A_dxVUt8yw9_0;
	wire w_dff_A_vNmnKIdx4_0;
	wire w_dff_A_e40IayJq1_0;
	wire w_dff_A_70k8EJs98_0;
	wire w_dff_A_8QRVLjO96_0;
	wire w_dff_A_pPh0vQUz9_0;
	wire w_dff_A_i338GVR02_0;
	wire w_dff_A_69oAD4ky3_0;
	wire w_dff_A_ZZzzjOXd1_0;
	wire w_dff_A_EEibSwoO2_0;
	wire w_dff_B_ehgFbZM29_1;
	wire w_dff_B_CfPz1sW61_1;
	wire w_dff_B_HQwbsi2q9_1;
	wire w_dff_B_uGVUTUZu2_1;
	wire w_dff_B_I0bJqcBs1_1;
	wire w_dff_B_mhJJuICq2_1;
	wire w_dff_B_3fkMhPZL9_1;
	wire w_dff_B_sVqsQlWz2_1;
	wire w_dff_B_2qC9ernC1_1;
	wire w_dff_B_l4AxyD8e1_1;
	wire w_dff_B_qqGPhaID0_1;
	wire w_dff_B_hkBaqYUO0_1;
	wire w_dff_A_oI3U0KAt2_0;
	wire w_dff_A_CZbsdVEy4_0;
	wire w_dff_A_l2rWvW2k6_0;
	wire w_dff_A_F5f6imAi0_0;
	wire w_dff_A_s9IBI8gC0_0;
	wire w_dff_A_L7VoPall2_0;
	wire w_dff_A_FZpxkJq41_0;
	wire w_dff_A_nSH68aSX5_0;
	wire w_dff_A_LfmZrE2x6_0;
	wire w_dff_A_J8sXJTQj3_0;
	wire w_dff_A_K2WTmrKj2_0;
	wire w_dff_A_nK8oxufB2_0;
	wire w_dff_A_1YlUi9QA2_0;
	wire w_dff_A_a0PbLUTj5_0;
	wire w_dff_B_0KXIUTjI6_1;
	wire w_dff_B_VjEdy8BS3_1;
	wire w_dff_B_1QgWNgf25_1;
	wire w_dff_B_Lm04xTtY7_1;
	wire w_dff_B_MjDQSxLh6_1;
	wire w_dff_B_xGYmIRLX6_1;
	wire w_dff_B_hWmYXbn75_1;
	wire w_dff_B_U1JzXxtl2_1;
	wire w_dff_B_yGIUHPSr3_1;
	wire w_dff_B_IV2jBIFP1_1;
	wire w_dff_A_urhleK3H5_0;
	wire w_dff_A_copowyB36_0;
	wire w_dff_A_u06mY1GP6_0;
	wire w_dff_A_rzp7B8dk5_0;
	wire w_dff_A_881PFUpB7_0;
	wire w_dff_A_hZgS5Bne6_0;
	wire w_dff_A_I2LyFV8Y8_0;
	wire w_dff_A_ylvADaxH1_0;
	wire w_dff_A_eVvk4y9j7_0;
	wire w_dff_A_IkWXygCx2_0;
	wire w_dff_A_lVJYfrnY4_0;
	wire w_dff_A_gUdkwqQc8_0;
	wire w_dff_B_dMneHK9C0_1;
	wire w_dff_B_mzwvJ4S71_1;
	wire w_dff_B_KAqqqU1e9_1;
	wire w_dff_B_di436h908_1;
	wire w_dff_B_TGYqgnsR9_1;
	wire w_dff_B_Z1Tp3tO33_1;
	wire w_dff_B_RFWMJ7Pm1_1;
	wire w_dff_B_fQZLEDiW3_1;
	wire w_dff_A_mwVSDR3y2_0;
	wire w_dff_A_caceFrAU7_0;
	wire w_dff_A_MLhWjLzD1_0;
	wire w_dff_A_RVlWy1fW8_0;
	wire w_dff_A_Q0Bag0Gl3_0;
	wire w_dff_A_sNTl6OET2_0;
	wire w_dff_A_jRTJA5X13_0;
	wire w_dff_A_2TqyeKPW3_0;
	wire w_dff_A_wcpvyPjQ9_0;
	wire w_dff_A_AFqrBfsz6_0;
	wire w_dff_B_oW5xUkWv9_1;
	wire w_dff_B_9WApEw879_1;
	wire w_dff_B_IewJZG8Z2_1;
	wire w_dff_B_AUVscL8l3_1;
	wire w_dff_B_Fts5z9WF7_1;
	wire w_dff_B_q9owYeI12_1;
	wire w_dff_A_xbYlxVGw3_0;
	wire w_dff_B_BBdFlk5W7_2;
	wire w_dff_B_CIHAMHnt6_2;
	wire w_dff_B_z1dMPwYz1_1;
	wire w_dff_A_7w36pcmb3_0;
	wire w_dff_A_FYmzH7fy9_0;
	wire w_dff_A_u5BQHdau1_0;
	wire w_dff_A_OBTyKFJL9_0;
	wire w_dff_A_Ck4bOiEB2_0;
	wire w_dff_A_Bv8lsQaE1_1;
	wire w_dff_B_sc9KY8Fy9_1;
	wire w_dff_B_E7g2rWZE1_1;
	wire w_dff_B_g0p1OFM37_1;
	wire w_dff_A_BhjmWNl43_0;
	wire w_dff_A_VGcuZtuh7_0;
	wire w_dff_A_D8ZagyVs8_0;
	wire w_dff_A_KsYCjYWA6_1;
	wire w_dff_A_gqHF4DZl2_0;
	wire w_dff_A_mXBLWQWm6_1;
	wire w_dff_B_pUEoHEdA2_2;
	wire w_dff_B_VjDpVPtW5_2;
	wire w_dff_B_CDiezGLX1_2;
	wire w_dff_B_hrNtueNY6_2;
	wire w_dff_B_xzXMQ78K6_2;
	wire w_dff_B_KnVJIlNm9_2;
	wire w_dff_B_GwgI0yLp5_2;
	wire w_dff_B_Sj5HycJh8_2;
	wire w_dff_B_uiEOOmkb8_2;
	wire w_dff_B_pw2WIRZJ3_2;
	wire w_dff_B_Mrqkuyqf2_2;
	wire w_dff_B_Y9sEi3Sb2_2;
	wire w_dff_B_ejez8uTU3_2;
	wire w_dff_B_srZchfgQ1_2;
	wire w_dff_B_mmxntYNI2_2;
	wire w_dff_B_0xu7klg74_2;
	wire w_dff_B_8n6gF85X6_2;
	wire w_dff_B_M41J3GWs9_2;
	wire w_dff_B_1NQNQZI22_2;
	wire w_dff_B_UKevyvjR8_2;
	wire w_dff_B_hXTjTZ819_2;
	wire w_dff_B_ec8USU462_2;
	wire w_dff_B_XHM6P4fV4_2;
	wire w_dff_B_nmxeaKC10_2;
	wire w_dff_B_QUSUmLwB4_2;
	wire w_dff_B_eIfUjQ2X7_2;
	wire w_dff_B_c5kKzlAa5_2;
	wire w_dff_B_dN2IENDA3_2;
	wire w_dff_B_zWIz0fXl1_2;
	wire w_dff_B_Dx5Vtea18_2;
	wire w_dff_B_Zu75j4Lr1_2;
	wire w_dff_B_BCStcs3G3_2;
	wire w_dff_B_Hws5aiKZ5_2;
	wire w_dff_B_GLO8DITt9_2;
	wire w_dff_A_03eNmzSV3_1;
	wire w_dff_A_UvcgMejF3_2;
	wire w_dff_B_Pl34Mh8Q8_3;
	wire w_dff_B_Babty6GB4_2;
	wire w_dff_B_nYw7Cytt7_2;
	wire w_dff_B_lqMIemrn7_2;
	wire w_dff_B_ZV3VsDIL2_2;
	wire w_dff_B_2MIdKlGR5_2;
	wire w_dff_B_LgUTvbRa3_2;
	wire w_dff_B_pAzOzIkd7_2;
	wire w_dff_B_6MWRjY6G2_2;
	wire w_dff_B_O7kF07mM5_2;
	wire w_dff_B_doLjYIdy4_2;
	wire w_dff_B_ErzC8j3T4_2;
	wire w_dff_B_lrDU8tK61_2;
	wire w_dff_B_XhXMM1HG7_2;
	wire w_dff_B_fMDKbW5C9_2;
	wire w_dff_B_DX9eR9X29_2;
	wire w_dff_B_cYuBZ7xA6_2;
	wire w_dff_B_9bpfnbwm4_2;
	wire w_dff_B_TNWgqI0m0_2;
	wire w_dff_B_DcQtgnxc5_2;
	wire w_dff_B_HAjKsZxT4_2;
	wire w_dff_B_cPlr3C5O0_2;
	wire w_dff_B_bz5LR08S5_2;
	wire w_dff_B_3LKMzIiD1_2;
	wire w_dff_B_Ov38ClNX8_2;
	wire w_dff_B_yZeCImj18_2;
	wire w_dff_B_xHUV53na8_2;
	wire w_dff_B_nJwKoeBn6_2;
	wire w_dff_B_ddw9zLfN6_2;
	wire w_dff_B_lTD0oQA26_2;
	wire w_dff_B_p388mCI49_2;
	wire w_dff_B_USy1Trii9_2;
	wire w_dff_B_kqnKkiIb2_1;
	wire w_dff_B_Hu1BJ9Py4_1;
	wire w_dff_B_7x97j8du0_1;
	wire w_dff_B_sLCnAuXu5_1;
	wire w_dff_B_DDd5QNhG3_1;
	wire w_dff_B_25yuYMur2_1;
	wire w_dff_B_Aln5U4oX1_1;
	wire w_dff_B_uAnphWv57_1;
	wire w_dff_B_FzFs4l730_1;
	wire w_dff_B_36YYKauh5_1;
	wire w_dff_B_fu8sMLXT9_1;
	wire w_dff_B_1tIyPv249_1;
	wire w_dff_B_GZXxZIVQ1_1;
	wire w_dff_B_aj8gI9Eh7_1;
	wire w_dff_B_aMcPJ7eC0_1;
	wire w_dff_B_XkpuDmtV4_1;
	wire w_dff_B_H7x1NHHF5_1;
	wire w_dff_B_I7qfQnZh2_1;
	wire w_dff_B_HhvaNsXh1_1;
	wire w_dff_B_yUOZu5MH2_1;
	wire w_dff_B_BnPStVUf6_1;
	wire w_dff_B_Fjf7Xnb44_1;
	wire w_dff_B_PYyFesMV4_1;
	wire w_dff_B_aTbs3Z4Y8_1;
	wire w_dff_B_s9FXjr378_1;
	wire w_dff_B_GhgI8sMn9_1;
	wire w_dff_B_b3OvboPa2_1;
	wire w_dff_B_tapHX3J87_1;
	wire w_dff_A_DcHsrmTj0_0;
	wire w_dff_A_X9EcOps89_0;
	wire w_dff_A_tDpBYWhs0_0;
	wire w_dff_A_PIoYYLe65_0;
	wire w_dff_A_TyrVEJwB5_0;
	wire w_dff_A_tUmYli7r3_0;
	wire w_dff_A_B5SWPUFX6_0;
	wire w_dff_A_qUjQ0fw15_0;
	wire w_dff_A_byfQ5dol3_0;
	wire w_dff_A_ADxtSsGn7_0;
	wire w_dff_A_R9DfQBYp6_0;
	wire w_dff_A_F7KZfXTX4_0;
	wire w_dff_A_DctNQRuQ9_0;
	wire w_dff_A_XZzIT9oc9_0;
	wire w_dff_A_rGgClRSu2_0;
	wire w_dff_A_1ArKhLZG5_0;
	wire w_dff_A_nd0uN8eP6_0;
	wire w_dff_A_6JNmbeze2_0;
	wire w_dff_A_861fChDR6_0;
	wire w_dff_A_R20mrMac7_0;
	wire w_dff_A_A1IAdkBD1_0;
	wire w_dff_A_ir0Ooy688_0;
	wire w_dff_A_bnnfhVE25_0;
	wire w_dff_A_SiTqRunJ6_0;
	wire w_dff_A_nimgtCq04_0;
	wire w_dff_A_0Hzxoq856_0;
	wire w_dff_A_tUjyESBT0_0;
	wire w_dff_A_08opqNZx2_0;
	wire w_dff_A_KhOaql1O5_0;
	wire w_dff_A_bENhUFb61_0;
	wire w_dff_A_QQiW9jHY7_1;
	wire w_dff_A_UZCyLOk90_2;
	wire w_dff_A_tT4vusQK8_0;
	wire w_dff_A_FJ0hg7Qw3_0;
	wire w_dff_A_PObZri7O3_0;
	wire w_dff_A_8oqumgGL0_0;
	wire w_dff_A_0qPY32M88_0;
	wire w_dff_A_QW3D3Aaz4_0;
	wire w_dff_A_wK2JlDMM7_0;
	wire w_dff_A_e8FCEq2U7_0;
	wire w_dff_A_HrpWBUEL6_0;
	wire w_dff_A_PM6eaZ0h4_0;
	wire w_dff_A_4Lmm1Ver6_0;
	wire w_dff_A_ZSzMyIF78_0;
	wire w_dff_A_uxSz08EX3_0;
	wire w_dff_A_l6Lu9EAc0_0;
	wire w_dff_A_fodFrSok9_0;
	wire w_dff_A_d4BkEOxs1_0;
	wire w_dff_A_yzBKiAe29_0;
	wire w_dff_A_D77r10yO3_0;
	wire w_dff_A_Kwtkl8wZ9_0;
	wire w_dff_A_VuFm5zs82_0;
	wire w_dff_A_z4S8U2114_0;
	wire w_dff_A_E0zGS5465_0;
	wire w_dff_A_doKv2wNU0_0;
	wire w_dff_A_p1w6RrO36_0;
	wire w_dff_A_TSP6erdd4_0;
	wire w_dff_A_wBTF6tG97_0;
	wire w_dff_A_lbCS54R79_0;
	wire w_dff_A_cjuBMvDR1_1;
	wire w_dff_A_1CFFVbwM8_2;
	wire w_dff_A_Egp6zTmU2_0;
	wire w_dff_A_xLqVU8W88_0;
	wire w_dff_A_Gt6SSnBR8_0;
	wire w_dff_A_6VHD1qXu6_0;
	wire w_dff_A_AiHNnsgj0_0;
	wire w_dff_A_iQ16p6fm1_0;
	wire w_dff_A_KJhlpZXr4_0;
	wire w_dff_A_OUM44gny1_0;
	wire w_dff_A_ivOB8jzk1_0;
	wire w_dff_A_15ZPBWxq5_0;
	wire w_dff_A_IeSFViUk8_0;
	wire w_dff_A_W1jKxoDm3_0;
	wire w_dff_A_UwHW28Du2_0;
	wire w_dff_A_BlSkSZEg8_0;
	wire w_dff_A_5b7OK6dR3_0;
	wire w_dff_A_XZ7qrrG87_0;
	wire w_dff_A_uCOA7kCG7_0;
	wire w_dff_A_M4IutWMU0_0;
	wire w_dff_A_RadhUKnM2_0;
	wire w_dff_A_Fct10wJE9_0;
	wire w_dff_A_kpmSESC04_0;
	wire w_dff_A_2yu0lIUe7_0;
	wire w_dff_A_dx5QL2HK5_0;
	wire w_dff_A_ngALKgO94_0;
	wire w_dff_A_A06Hb1ms3_0;
	wire w_dff_A_ZQVdk6Lq8_1;
	wire w_dff_A_gfmfUuPd7_2;
	wire w_dff_A_e0kImvxC3_0;
	wire w_dff_A_eD7Ix6Wj8_0;
	wire w_dff_A_3uGzoZuT4_0;
	wire w_dff_A_4RP6p57e9_0;
	wire w_dff_A_QW03tm6Y2_0;
	wire w_dff_A_9j1eNQgB5_0;
	wire w_dff_A_UTmAqdE04_0;
	wire w_dff_A_jZk2AhTA9_0;
	wire w_dff_A_zVwnH6Ss4_0;
	wire w_dff_A_VN2IVTXW2_0;
	wire w_dff_A_49Yn0lRu4_0;
	wire w_dff_A_MFXnEAzf0_0;
	wire w_dff_A_Giydvbdx5_0;
	wire w_dff_A_a5G4Tqy92_0;
	wire w_dff_A_nwlR48mJ8_0;
	wire w_dff_A_uHe5KRiu0_0;
	wire w_dff_A_oYEBCFhb0_0;
	wire w_dff_A_dOlZllaD2_0;
	wire w_dff_A_PLYszZBE0_0;
	wire w_dff_A_vtt2ordJ5_0;
	wire w_dff_A_WaCa1zKv0_0;
	wire w_dff_A_Ub49KRTY6_0;
	wire w_dff_A_ILxVErOV7_0;
	wire w_dff_A_I5tXqzfD0_1;
	wire w_dff_A_QfR65i8R2_2;
	wire w_dff_A_OgKaEuyH0_0;
	wire w_dff_A_JNRIqG7Q1_0;
	wire w_dff_A_kGZrLCOB5_0;
	wire w_dff_A_52cI6y6R4_0;
	wire w_dff_A_b10JSLqZ0_0;
	wire w_dff_A_Y2wZLREn3_0;
	wire w_dff_A_1JcpxVic2_0;
	wire w_dff_A_9qq9DEtF6_0;
	wire w_dff_A_WjyFuhvk7_0;
	wire w_dff_A_6eDZJBO78_0;
	wire w_dff_A_G48Bm8im9_0;
	wire w_dff_A_BHNaKbSr7_0;
	wire w_dff_A_S3fzd61M0_0;
	wire w_dff_A_njWEN1843_0;
	wire w_dff_A_AqQn5PND0_0;
	wire w_dff_A_j67mQTt59_0;
	wire w_dff_A_V714H1cc5_0;
	wire w_dff_A_ivOfx6Ti0_0;
	wire w_dff_A_PIIyxv3e4_0;
	wire w_dff_A_2o2IXzwD8_0;
	wire w_dff_A_91CmjfIu8_0;
	wire w_dff_A_X4AjoJhn4_1;
	wire w_dff_A_uXsEZDhL1_2;
	wire w_dff_B_ZgcXkTFS6_3;
	wire w_dff_B_tvsvbyGX0_3;
	wire w_dff_B_c9r1jGgp4_3;
	wire w_dff_A_xvNLAp835_0;
	wire w_dff_A_S9s49NdZ4_0;
	wire w_dff_A_eZYOnNfg9_0;
	wire w_dff_A_eiSqoekV6_0;
	wire w_dff_A_B3r5OUTw8_0;
	wire w_dff_A_WKlKpjuE4_0;
	wire w_dff_A_TFp0WR8M6_0;
	wire w_dff_A_u3MyCNRN6_0;
	wire w_dff_A_GSyojAc74_0;
	wire w_dff_A_AQoChlQw6_0;
	wire w_dff_A_wVj7xcz45_0;
	wire w_dff_A_r6LCIgO77_0;
	wire w_dff_A_ygdhYGnG1_0;
	wire w_dff_A_XiDKXq3e1_0;
	wire w_dff_A_52wPN3b80_0;
	wire w_dff_A_YabRlF152_0;
	wire w_dff_A_0eoWrf1S3_1;
	wire w_dff_A_iwaBUwCU1_2;
	wire w_dff_A_FrOgE1JG7_0;
	wire w_dff_A_PTUCHwB83_0;
	wire w_dff_A_nx9yNsZn8_0;
	wire w_dff_A_cTdyOx3I2_0;
	wire w_dff_A_FbsFObmB8_0;
	wire w_dff_A_lkubc8Xa2_0;
	wire w_dff_A_eeg1YH272_0;
	wire w_dff_A_zOYXO5LO6_0;
	wire w_dff_A_ufOV3YgE1_0;
	wire w_dff_A_ISQhXHx75_0;
	wire w_dff_A_LN0XjWtg3_0;
	wire w_dff_A_oFhOgkps0_0;
	wire w_dff_A_9yLDPtv77_0;
	wire w_dff_A_LOYtCh2c3_0;
	wire w_dff_A_0tGESKVt5_1;
	wire w_dff_A_naHyJ4d17_2;
	wire w_dff_A_5inedgFM2_0;
	wire w_dff_A_veKJvRCX5_0;
	wire w_dff_A_vauHgFrb2_0;
	wire w_dff_A_ET1t7Bcr2_0;
	wire w_dff_A_9KEQbPbd1_0;
	wire w_dff_A_HE5ukqLq5_0;
	wire w_dff_A_VHbxBVlD0_0;
	wire w_dff_A_k7H8XMyl3_0;
	wire w_dff_A_NQr1QQHL0_0;
	wire w_dff_A_V9tykzU10_0;
	wire w_dff_A_MvUuq6fk7_0;
	wire w_dff_A_AMQHIN923_0;
	wire w_dff_A_0A3wwcWf1_1;
	wire w_dff_A_c04hZHBx0_2;
	wire w_dff_A_dAiBishI8_0;
	wire w_dff_A_Aor2FHKo2_0;
	wire w_dff_A_SWnGiDW03_0;
	wire w_dff_A_yMoETBab4_0;
	wire w_dff_A_8v3CManF2_0;
	wire w_dff_A_ZmnPzlZr2_0;
	wire w_dff_A_PcH7twzX5_0;
	wire w_dff_A_Qu9OlvZc4_0;
	wire w_dff_A_Dcbj3qnk0_0;
	wire w_dff_A_BpAHiX1R2_0;
	wire w_dff_A_oiF60WcB7_1;
	wire w_dff_A_Cvh7nZWc3_2;
	wire w_dff_A_oumENl7w4_0;
	wire w_dff_A_PqWvTibw6_0;
	wire w_dff_A_augNwgFE2_0;
	wire w_dff_A_x4cVkPpp2_0;
	wire w_dff_A_3nmj66fQ7_0;
	wire w_dff_A_HOaGsRze1_0;
	wire w_dff_A_Pr58Vjkp3_0;
	wire w_dff_A_EVTnbB3G6_0;
	wire w_dff_A_t9jJ0Ax06_1;
	wire w_dff_A_ZnVzuhX42_2;
	wire w_dff_A_vzDX4kE98_0;
	wire w_dff_A_DCn4SF351_0;
	wire w_dff_A_MTsb8jqH3_0;
	wire w_dff_A_VBtoZvs29_0;
	wire w_dff_A_FwDOSz354_0;
	wire w_dff_A_YElQJLx72_0;
	wire w_dff_A_rLbe5iWw9_1;
	wire w_dff_A_WU05vbqJ5_2;
	wire w_dff_B_SdvaenAL9_3;
	wire w_dff_B_qOlwIYSL5_3;
	wire w_dff_B_7XBAQlWe7_1;
	wire w_dff_A_uVcTUwdv7_0;
	wire w_dff_A_ScPbN5a19_0;
	wire w_dff_A_4He3wXXc8_0;
	wire w_dff_A_V7rxrfus7_0;
	wire w_dff_B_5qk6RfLR5_2;
	wire w_dff_B_AwpYgIu32_2;
	wire w_dff_B_rxyDG2M89_2;
	wire w_dff_B_7wknFk848_2;
	wire w_dff_B_9DYGw7Dh6_2;
	wire w_dff_B_e8hpzakL7_2;
	wire w_dff_B_amro8CZb0_2;
	wire w_dff_B_YyeAAAiz1_2;
	wire w_dff_B_W0peWllr3_2;
	wire w_dff_B_hqaT3nBH6_2;
	wire w_dff_B_m9SCfVrB9_2;
	wire w_dff_B_GeMbTlVP7_2;
	wire w_dff_B_KzQo3o3R9_2;
	wire w_dff_B_0cdUS7TV9_2;
	wire w_dff_B_5rywKQS15_2;
	wire w_dff_B_kylEJjic3_2;
	wire w_dff_B_TptfY84m1_2;
	wire w_dff_B_brYRrtJW9_2;
	wire w_dff_B_Pt76kV2A9_2;
	wire w_dff_B_Wi3KLufh9_2;
	wire w_dff_B_QTdE5kJz2_2;
	wire w_dff_B_AQg3C7z21_2;
	wire w_dff_B_3w4zosuD7_2;
	wire w_dff_B_kiWf3GJU6_2;
	wire w_dff_B_FuVVGGMD1_2;
	wire w_dff_B_IGRs6V3n6_2;
	wire w_dff_B_Dyi1YIAH2_2;
	wire w_dff_B_90dv32rF7_2;
	wire w_dff_B_utK3GTcc2_2;
	wire w_dff_B_w8W9LDhj2_2;
	wire w_dff_B_4wMmvEWk7_2;
	wire w_dff_B_83MZuWrc5_2;
	wire w_dff_B_cLBThaVd3_2;
	wire w_dff_B_L1jNxXFS8_2;
	wire w_dff_B_ZG439JIz6_2;
	wire w_dff_A_dJHV3D2E4_0;
	wire w_dff_B_fLWRSZbu3_1;
	wire w_dff_B_5Gg4QPp35_2;
	wire w_dff_B_yqiSydbO6_2;
	wire w_dff_B_uJP7Zt6o2_2;
	wire w_dff_B_JHMxpmCT3_2;
	wire w_dff_B_wBob4Vtm3_2;
	wire w_dff_B_aJymxLPy8_2;
	wire w_dff_B_m3FvqUI57_2;
	wire w_dff_B_JhXFxKV94_2;
	wire w_dff_B_l6Jk3JnJ3_2;
	wire w_dff_B_63EujrUG6_2;
	wire w_dff_B_AxiXIGmo8_2;
	wire w_dff_B_YK2EEB5H0_2;
	wire w_dff_B_58771CmY8_2;
	wire w_dff_B_8Piz0tfp2_2;
	wire w_dff_B_mceGSAbA7_2;
	wire w_dff_B_4oEiDqDh3_2;
	wire w_dff_B_K1sfVUCj5_2;
	wire w_dff_B_yvGS4cgp2_2;
	wire w_dff_B_jQjRYNtY3_2;
	wire w_dff_B_jZRzcMb97_2;
	wire w_dff_B_4QPYsdQu2_2;
	wire w_dff_B_1REA3eFh0_2;
	wire w_dff_B_igXWHAIW3_2;
	wire w_dff_B_VjwhGhiQ1_2;
	wire w_dff_B_ZfPwlrQh7_2;
	wire w_dff_B_baM5UuUj9_2;
	wire w_dff_B_C97EUB5o5_2;
	wire w_dff_B_ay4RHgkB9_2;
	wire w_dff_B_PrqImqy58_2;
	wire w_dff_B_NFctmz8z3_2;
	wire w_dff_B_UGGY7aL27_2;
	wire w_dff_B_aGAepYLi9_2;
	wire w_dff_A_ifldbHus3_1;
	wire w_dff_A_Lk7C61MK4_0;
	wire w_dff_A_XTeS7fHm4_0;
	wire w_dff_A_CG1Whsdx0_0;
	wire w_dff_A_cgePzAdx2_0;
	wire w_dff_A_rPrYnz3m8_0;
	wire w_dff_A_snzH7SAi8_0;
	wire w_dff_A_ueBQLTmq2_0;
	wire w_dff_A_6BaDtHaP1_0;
	wire w_dff_A_lkVvhpXu5_0;
	wire w_dff_A_YaOjGzi51_0;
	wire w_dff_A_mqFlHYbJ9_0;
	wire w_dff_A_EXlWsVTM2_0;
	wire w_dff_A_fIUAoLko8_0;
	wire w_dff_A_XaNoVa8a3_0;
	wire w_dff_A_P0gIU8ib9_0;
	wire w_dff_A_rVVKLcIm2_0;
	wire w_dff_A_o261iGzt7_0;
	wire w_dff_A_tjK8g2Eb0_0;
	wire w_dff_A_kEephMl80_0;
	wire w_dff_A_KysHcyIl8_0;
	wire w_dff_A_ywZU3uOo5_0;
	wire w_dff_A_sbbrMCKZ9_0;
	wire w_dff_A_R3bd3qsZ2_0;
	wire w_dff_A_8yZubp9V5_0;
	wire w_dff_A_PygO025X9_0;
	wire w_dff_A_ElAq0Bqn2_0;
	wire w_dff_A_nJEAJzXB1_0;
	wire w_dff_A_b45eTMbn1_0;
	wire w_dff_A_dbuy7M5F6_0;
	wire w_dff_A_XGAWw9VZ5_0;
	wire w_dff_A_x6b9m6GW6_0;
	wire w_dff_B_cMTiWGax5_1;
	wire w_dff_B_uF6v6l9F4_2;
	wire w_dff_B_UJbDZzLl8_2;
	wire w_dff_B_33pWAx9J0_2;
	wire w_dff_B_5fZfaQUm0_2;
	wire w_dff_B_q4jJURHC3_2;
	wire w_dff_B_FNQhTGUT2_2;
	wire w_dff_B_OzDQ8Unp0_2;
	wire w_dff_B_52RZW9OQ6_2;
	wire w_dff_B_PsxwXRH22_2;
	wire w_dff_B_xxGuBGhD5_2;
	wire w_dff_B_SZaXjwHU5_2;
	wire w_dff_B_KAEC14Dg6_2;
	wire w_dff_B_QU9MbDhP0_2;
	wire w_dff_B_ySKUMeI93_2;
	wire w_dff_B_9h6NlaLw6_2;
	wire w_dff_B_O16Gc5wT2_2;
	wire w_dff_B_5IcWhh5n7_2;
	wire w_dff_B_hjkZlS5N2_2;
	wire w_dff_B_14T0t1lH1_2;
	wire w_dff_B_0JAEdSmU9_2;
	wire w_dff_B_XTMiFsPL7_2;
	wire w_dff_B_wyNebLeA6_2;
	wire w_dff_B_MJSKrjHa7_2;
	wire w_dff_B_oMDPKNTq5_2;
	wire w_dff_B_sZXq265h8_2;
	wire w_dff_B_7jkSTk9B6_2;
	wire w_dff_B_VTnCxu1s2_1;
	wire w_dff_B_o38pbutf8_2;
	wire w_dff_B_mqHkqoQt4_2;
	wire w_dff_B_DvdHCQfH6_2;
	wire w_dff_B_jIPfL9T36_2;
	wire w_dff_B_X7U5MrB34_2;
	wire w_dff_B_5W15h3EU7_2;
	wire w_dff_B_gztwS6fZ1_2;
	wire w_dff_B_z4S3XMLE1_2;
	wire w_dff_B_RFLBCUDz3_2;
	wire w_dff_B_PauOrJSC1_2;
	wire w_dff_B_zATPdLnJ5_2;
	wire w_dff_B_5YYgbd1u8_2;
	wire w_dff_B_SN1BSypw1_2;
	wire w_dff_B_LgNK6NPy1_2;
	wire w_dff_B_mLM8j9FV1_2;
	wire w_dff_B_9GAvwy2G2_2;
	wire w_dff_B_8XIIRcp81_2;
	wire w_dff_B_bhEX6O7d6_2;
	wire w_dff_B_pwNRDr5u7_2;
	wire w_dff_B_HNJeLkKb6_2;
	wire w_dff_B_fyN3ZaDT0_2;
	wire w_dff_B_EIspindm2_2;
	wire w_dff_B_hWChproN0_2;
	wire w_dff_B_HJozdlbv8_2;
	wire w_dff_B_DGB6GK2U4_1;
	wire w_dff_B_z5Mrl2d49_2;
	wire w_dff_B_ji1O4XeW8_2;
	wire w_dff_B_OGC6xtUR8_2;
	wire w_dff_B_U6VqR7Tu6_2;
	wire w_dff_B_BAP7ZMkT0_2;
	wire w_dff_B_EnyMka5z8_2;
	wire w_dff_B_SLbRyJW77_2;
	wire w_dff_B_TiEfzTcg3_2;
	wire w_dff_B_xfIGiNse3_2;
	wire w_dff_B_ZmuQ96UD1_2;
	wire w_dff_B_x3eC20vg7_2;
	wire w_dff_B_AgPuE6J71_2;
	wire w_dff_B_TJfFCRQk3_2;
	wire w_dff_B_fcLC42gh6_2;
	wire w_dff_B_9prlxDHj9_2;
	wire w_dff_B_4xxIRRzl4_2;
	wire w_dff_B_RBwEnbfL7_2;
	wire w_dff_B_yCQscvb85_2;
	wire w_dff_B_OqccJEAx6_2;
	wire w_dff_B_eItrhepZ7_2;
	wire w_dff_B_XJ4UuzMf0_2;
	wire w_dff_B_CtXZPoD54_2;
	wire w_dff_B_AYEMt2pb5_1;
	wire w_dff_B_yiFikY6S0_2;
	wire w_dff_B_9GWHbyoQ9_2;
	wire w_dff_B_mDMsgMjl5_2;
	wire w_dff_B_nnbUSo3H8_2;
	wire w_dff_B_1w7uZ2C55_2;
	wire w_dff_B_hwRikIEi1_2;
	wire w_dff_B_0DFTMkaz9_2;
	wire w_dff_B_0VweNF2b0_2;
	wire w_dff_B_A3vMFwbm9_2;
	wire w_dff_B_EYYS5jdu4_2;
	wire w_dff_B_NCfSB1RD5_2;
	wire w_dff_B_ZsEOCC6H8_2;
	wire w_dff_B_6I6clgRr8_2;
	wire w_dff_B_2MaNKVGT2_2;
	wire w_dff_B_bpGrHt7i6_2;
	wire w_dff_B_VXpvDMr24_2;
	wire w_dff_B_4ZTR1YRD0_2;
	wire w_dff_B_SOxsZYhb7_2;
	wire w_dff_B_ztEKzG725_2;
	wire w_dff_B_48wM55a46_2;
	wire w_dff_B_JRaUOXWj3_1;
	wire w_dff_B_o3o5kmgZ9_2;
	wire w_dff_B_i0dHUurS3_2;
	wire w_dff_B_92YhrZOP6_2;
	wire w_dff_B_WUM9aKaa4_2;
	wire w_dff_B_n4bOWrrF5_2;
	wire w_dff_B_dNzqswh10_2;
	wire w_dff_B_InYXbte39_2;
	wire w_dff_B_C2hvYceW0_2;
	wire w_dff_B_Iak6MvXc4_2;
	wire w_dff_B_icPAnBW05_2;
	wire w_dff_B_lOru7j3E7_2;
	wire w_dff_B_hnmhJOxM1_2;
	wire w_dff_B_VaZbsnba9_2;
	wire w_dff_B_Oxu1mLrj6_2;
	wire w_dff_B_SUxmqice2_2;
	wire w_dff_B_Qbc2p17A7_2;
	wire w_dff_B_j48qRoWx6_2;
	wire w_dff_B_fgyzPuhR6_2;
	wire w_dff_B_qwUALIAQ9_2;
	wire w_dff_B_vWAWZdc59_2;
	wire w_dff_B_N4sh3q5e5_2;
	wire w_dff_B_P93Tff5z4_1;
	wire w_dff_B_7sBlSo2X7_2;
	wire w_dff_B_dD1y967m9_2;
	wire w_dff_B_AC9zETx47_2;
	wire w_dff_B_JvXKLkmO7_2;
	wire w_dff_B_WjND6SVT6_2;
	wire w_dff_B_Aga9P3Bs4_2;
	wire w_dff_B_o3xOySRJ2_2;
	wire w_dff_B_QLSsXnrH2_2;
	wire w_dff_B_vsFXu0EJ6_2;
	wire w_dff_B_iwAi1GUU6_2;
	wire w_dff_B_oxmRtnfM1_2;
	wire w_dff_B_VCudCSLW9_2;
	wire w_dff_B_XG3grkrj8_2;
	wire w_dff_B_a6aAry2s3_1;
	wire w_dff_B_6BgSjQ4p0_2;
	wire w_dff_B_wSwAlr9b4_2;
	wire w_dff_B_5xNQ7vcN1_2;
	wire w_dff_B_BMKZfG7x8_2;
	wire w_dff_B_dITPWEAj9_2;
	wire w_dff_B_goRfSAGP9_2;
	wire w_dff_B_7hBaRknf8_2;
	wire w_dff_B_uUbNrxhr0_2;
	wire w_dff_B_ePYffLUN5_2;
	wire w_dff_B_XL44WUPg4_2;
	wire w_dff_B_aOXfa8sz8_2;
	wire w_dff_B_179JyEBS4_1;
	wire w_dff_B_wgfFPKcQ8_2;
	wire w_dff_B_4Mkdh8L65_2;
	wire w_dff_B_uzE8JzXO6_2;
	wire w_dff_B_Cx86ky2u9_2;
	wire w_dff_B_JEhgz6Oy5_2;
	wire w_dff_B_wESYyZfT3_2;
	wire w_dff_B_6SAplVxm9_2;
	wire w_dff_B_tC5J9qza7_2;
	wire w_dff_B_KZLo3TkJ9_2;
	wire w_dff_B_EK6M9CMC1_1;
	wire w_dff_B_eVakjd8v3_2;
	wire w_dff_B_sABgkMfb1_2;
	wire w_dff_B_L8BxoCXC8_2;
	wire w_dff_B_nx4Jfh7d1_2;
	wire w_dff_B_MI2MR9K84_2;
	wire w_dff_B_YljsIb8x7_2;
	wire w_dff_B_a0xbI5MR9_2;
	wire w_dff_B_0mJuPkMW1_1;
	wire w_dff_B_pycAoolc5_2;
	wire w_dff_B_jtqD1miP2_2;
	wire w_dff_B_BB597h2Q4_2;
	wire w_dff_B_si6JPCcA0_2;
	wire w_dff_B_U9BSC4ub3_2;
	wire w_dff_B_JOEeLthO3_1;
	wire w_dff_B_bJ3a7PNT8_2;
	wire w_dff_B_7EgRI1TZ8_2;
	wire w_dff_B_AmgMx0zO2_2;
	wire w_dff_B_2e37WqoN8_0;
	wire w_dff_B_KG6L1ole9_0;
	wire w_dff_B_R0DWTPDp5_2;
	wire w_dff_B_XyxqOr217_2;
	wire w_dff_A_XyCh9jAo8_1;
	wire w_dff_B_j8tgBVSe0_1;
	wire w_dff_B_CryD6Cfq3_1;
	wire w_dff_B_oilcDNtd4_2;
	wire w_dff_B_15zZ8kM33_2;
	wire w_dff_B_UbL0sGHz7_2;
	wire w_dff_B_cdtzEnhi5_2;
	wire w_dff_B_PRJkIcra5_2;
	wire w_dff_B_FzXg4FmR2_2;
	wire w_dff_B_vTFCoGC55_2;
	wire w_dff_B_wqfXGH9U4_2;
	wire w_dff_B_MsFJ0Z9w4_2;
	wire w_dff_B_qMH7nCs17_2;
	wire w_dff_B_nVJfKJMQ2_2;
	wire w_dff_B_paKERQX20_2;
	wire w_dff_B_7vOWv20M4_2;
	wire w_dff_B_i9DAn7Wh3_2;
	wire w_dff_B_cBjAkNjJ5_2;
	wire w_dff_B_a54AEM1u5_2;
	wire w_dff_B_YYsTaknn6_2;
	wire w_dff_B_rRDNzS7j6_2;
	wire w_dff_B_TLRYqo0p6_2;
	wire w_dff_B_Wy9Y70nD2_2;
	wire w_dff_B_CxVTMGzw1_2;
	wire w_dff_B_OWZ2oYMB0_2;
	wire w_dff_B_aBIHBdYF2_2;
	wire w_dff_B_cWwPpj9i9_2;
	wire w_dff_B_3mRUBu190_2;
	wire w_dff_B_PzJR96K57_2;
	wire w_dff_B_ZLBt1Kri8_2;
	wire w_dff_B_FUIbMm6V1_2;
	wire w_dff_B_P66wPTx76_2;
	wire w_dff_B_kRAFBaob1_2;
	wire w_dff_B_FXSYPZiZ0_2;
	wire w_dff_B_W0Fm7O9J0_2;
	wire w_dff_B_gxhM8V879_2;
	wire w_dff_B_zVNRmedN4_2;
	wire w_dff_B_IcVXHOmB8_2;
	wire w_dff_B_z2eft3Hx1_2;
	wire w_dff_B_5hCCQ6uO8_2;
	wire w_dff_B_R6efCo3Q3_2;
	wire w_dff_B_HHg7LBou9_2;
	wire w_dff_B_OZPvsSCI9_2;
	wire w_dff_B_cOmbRTJQ6_2;
	wire w_dff_B_JE1vqca74_2;
	wire w_dff_B_BjBDuWrd8_2;
	wire w_dff_B_vs2VIFTH1_2;
	wire w_dff_B_1Uf69JuG7_2;
	wire w_dff_B_SnvcmMeL2_2;
	wire w_dff_B_Y9GmZhvq2_2;
	wire w_dff_B_JDytO8bX0_2;
	wire w_dff_B_9jhhSUmO9_2;
	wire w_dff_B_sBmjEpyi9_2;
	wire w_dff_B_rn2e8mvC2_2;
	wire w_dff_B_sGVMbOxG4_2;
	wire w_dff_B_pM8lxuAE9_2;
	wire w_dff_B_YtEAZOW73_2;
	wire w_dff_B_93O3wBcX7_2;
	wire w_dff_B_bWjjSqsC9_2;
	wire w_dff_B_sRdUSWLX1_2;
	wire w_dff_B_gB2azBy89_2;
	wire w_dff_B_RP9SRDAQ2_2;
	wire w_dff_B_I0ZgTe0E6_2;
	wire w_dff_B_dfF5PRfQ1_2;
	wire w_dff_B_yA2vWf9f0_2;
	wire w_dff_B_OLpM4IRT2_2;
	wire w_dff_B_8hVdvtN82_2;
	wire w_dff_B_rBlPwu5Q4_2;
	wire w_dff_B_pyJdQncl1_2;
	wire w_dff_B_WGkBMv0o2_2;
	wire w_dff_B_sNTjJaJO2_1;
	wire w_dff_B_lMtLiVv80_2;
	wire w_dff_B_Kny7VouC8_2;
	wire w_dff_B_dZSAP3R21_2;
	wire w_dff_B_OwvQ85aW2_2;
	wire w_dff_B_4uMYYScH7_2;
	wire w_dff_B_v762xUcz5_2;
	wire w_dff_B_OQC4Q1wz8_2;
	wire w_dff_B_Lm7qDqoX9_2;
	wire w_dff_B_XSrmnJyZ8_2;
	wire w_dff_B_qWy7PIuP2_2;
	wire w_dff_B_TaaW1kKq3_2;
	wire w_dff_B_E1vGASyh0_2;
	wire w_dff_B_dvRv323c1_2;
	wire w_dff_B_7IEjVGqe0_2;
	wire w_dff_B_deC93HoG7_2;
	wire w_dff_B_hwcygG2j6_2;
	wire w_dff_B_WxEsqBZd6_2;
	wire w_dff_B_PXrT6IEk6_2;
	wire w_dff_B_4PMjx43R2_2;
	wire w_dff_B_uErkJBpM7_2;
	wire w_dff_B_GovHtXWP9_2;
	wire w_dff_B_T65xFP7s6_2;
	wire w_dff_B_lzAbEm1k0_2;
	wire w_dff_B_ZP2hEZ8b5_2;
	wire w_dff_B_2k3mJCGL0_2;
	wire w_dff_B_3jQ5aiW55_2;
	wire w_dff_B_5rwIkS546_2;
	wire w_dff_B_8HzqBeLN7_2;
	wire w_dff_B_8XmM6ZQT5_1;
	wire w_dff_B_oSUCqHoB3_2;
	wire w_dff_B_my9IvFGK1_2;
	wire w_dff_B_YiQWaEqU1_2;
	wire w_dff_B_u7lwJHaZ3_2;
	wire w_dff_B_9t7pxeCg7_2;
	wire w_dff_B_eUo8E2kU9_2;
	wire w_dff_B_LhF1i4Iz2_2;
	wire w_dff_B_T8FOXlNM3_2;
	wire w_dff_B_FYlCwDAt3_2;
	wire w_dff_B_1ZOHWq8R5_2;
	wire w_dff_B_CwkQDiPc0_2;
	wire w_dff_B_sYHeRNCk2_2;
	wire w_dff_B_aGjVGPL39_2;
	wire w_dff_B_YOVeNT463_2;
	wire w_dff_B_lnXAyMkZ6_2;
	wire w_dff_B_i4E5udyy3_2;
	wire w_dff_B_7JvJSi6F0_2;
	wire w_dff_B_wY4HfYA84_2;
	wire w_dff_B_ZU3J9brb8_2;
	wire w_dff_B_kgDElL1k1_2;
	wire w_dff_B_beOPmkz14_2;
	wire w_dff_B_aUowkf4D8_2;
	wire w_dff_B_I3GgmAax8_2;
	wire w_dff_B_8rOpwDjW9_2;
	wire w_dff_B_jji0w7VI7_2;
	wire w_dff_B_h6QApWVR7_2;
	wire w_dff_B_WJTzbYWo0_1;
	wire w_dff_B_tBD6Qgke8_2;
	wire w_dff_B_U7EKFjLC5_2;
	wire w_dff_B_HSiI8sUR0_2;
	wire w_dff_B_RoZtcD7e1_2;
	wire w_dff_B_vuSO3C1n0_2;
	wire w_dff_B_0ik5aAyt4_2;
	wire w_dff_B_iew6PsxQ6_2;
	wire w_dff_B_BmsOrLXp2_2;
	wire w_dff_B_viRx4J9i1_2;
	wire w_dff_B_sbPfn3469_2;
	wire w_dff_B_pxMrcd2p7_2;
	wire w_dff_B_IaNmMKtE9_2;
	wire w_dff_B_XpB7DWee3_2;
	wire w_dff_B_EabPG5Cm7_2;
	wire w_dff_B_RXrPWNiU2_2;
	wire w_dff_B_TFV84nU96_2;
	wire w_dff_B_3Cg8V9mk8_2;
	wire w_dff_B_aYVoHewh1_2;
	wire w_dff_B_fHJr7jH17_2;
	wire w_dff_B_KjBqay244_2;
	wire w_dff_B_2rsRrtsE7_2;
	wire w_dff_B_AF7UR4pz2_2;
	wire w_dff_B_VW950xfM8_2;
	wire w_dff_B_RAjW8tPC7_2;
	wire w_dff_B_6nBwJ9zZ6_1;
	wire w_dff_B_TJoJ2Hpf9_2;
	wire w_dff_B_FOmVx54i5_2;
	wire w_dff_B_IJ8YVhio0_2;
	wire w_dff_B_PUBPL4wg6_2;
	wire w_dff_B_8IKTRe025_2;
	wire w_dff_B_ydpiG5zF6_2;
	wire w_dff_B_8UhFquDK7_2;
	wire w_dff_B_4LjAfNAM1_2;
	wire w_dff_B_8Q4aZSdX8_2;
	wire w_dff_B_WucYABgL9_2;
	wire w_dff_B_qSpmCzeu1_2;
	wire w_dff_B_LUNfMWw72_2;
	wire w_dff_B_B5LDE6At9_2;
	wire w_dff_B_VNOsjfTr9_2;
	wire w_dff_B_oJqZbqpz0_2;
	wire w_dff_B_ixdC6bzi3_2;
	wire w_dff_B_v4S9lgTS6_2;
	wire w_dff_B_l4KhkdhZ9_2;
	wire w_dff_B_YEvaUqN93_2;
	wire w_dff_B_hc8EAVp60_2;
	wire w_dff_B_hg8srLWe7_2;
	wire w_dff_B_GTVULd038_2;
	wire w_dff_B_mvT3gYh79_1;
	wire w_dff_B_RVUS5a2h9_2;
	wire w_dff_B_ggDE6zDg3_2;
	wire w_dff_B_l7bTxlJX5_2;
	wire w_dff_B_4SLqWwqp8_2;
	wire w_dff_B_Ovj3rpTv1_2;
	wire w_dff_B_xaXNsIvP0_2;
	wire w_dff_B_cbr649zh8_2;
	wire w_dff_B_IzZig3L51_2;
	wire w_dff_B_cLwDYBZt7_2;
	wire w_dff_B_aFHeId8D9_2;
	wire w_dff_B_k8gJGjYO9_2;
	wire w_dff_B_dFzZABtA2_2;
	wire w_dff_B_di7Gth1s0_2;
	wire w_dff_B_qHK1YvLl7_2;
	wire w_dff_B_t9gbcdDy4_2;
	wire w_dff_B_gVa2kFoR4_2;
	wire w_dff_B_Vzh9OvP67_2;
	wire w_dff_B_a9wQwVAx2_2;
	wire w_dff_B_5UxDSrDo0_2;
	wire w_dff_B_U7tVD6sA5_2;
	wire w_dff_B_v8QRd6LZ4_1;
	wire w_dff_B_8w2BWKKy4_2;
	wire w_dff_B_X7BbLtuU9_2;
	wire w_dff_B_x3q2Bcwx9_2;
	wire w_dff_B_XWG9cLbQ4_2;
	wire w_dff_B_2jqGrJnV1_2;
	wire w_dff_B_sz7LAJru1_2;
	wire w_dff_B_WFwaxirL5_2;
	wire w_dff_B_iS8NsnM98_2;
	wire w_dff_B_tbhI4mFC6_2;
	wire w_dff_B_YrDirVu17_2;
	wire w_dff_B_BBG1u3ts7_2;
	wire w_dff_B_Gd0BBvtD0_2;
	wire w_dff_B_f7h8Dusw2_2;
	wire w_dff_B_klHxXJKr7_2;
	wire w_dff_B_9XVQ6UH09_2;
	wire w_dff_B_XSJYdEVn0_2;
	wire w_dff_B_D0wlWiL92_2;
	wire w_dff_B_mMtDY7Ft3_2;
	wire w_dff_B_zBQXm9a34_1;
	wire w_dff_B_1vcisxuE7_2;
	wire w_dff_B_RVCFi1c31_2;
	wire w_dff_B_ExsH5ryU0_2;
	wire w_dff_B_XdZN0oQW5_2;
	wire w_dff_B_IQQ7YdGG9_2;
	wire w_dff_B_B36eK0DP3_2;
	wire w_dff_B_FMjixvov4_2;
	wire w_dff_B_6CP1r0ny1_2;
	wire w_dff_B_KnvoEbWM2_2;
	wire w_dff_B_GafvfmSv4_2;
	wire w_dff_B_MtNYffRt7_2;
	wire w_dff_B_fd4wgxW34_2;
	wire w_dff_B_PE2x74zx9_2;
	wire w_dff_B_4r0V9rLA0_2;
	wire w_dff_B_fHZXDJi48_2;
	wire w_dff_B_gd3sCwu39_2;
	wire w_dff_B_DwbZPHca6_2;
	wire w_dff_B_8LSZcutg8_2;
	wire w_dff_B_1aTwimwz5_2;
	wire w_dff_B_YDTgA7rp3_1;
	wire w_dff_B_y7DxDGZo8_2;
	wire w_dff_B_5mrxDeXX1_2;
	wire w_dff_B_Fl8KEnUB2_2;
	wire w_dff_B_KofwOBxw2_2;
	wire w_dff_B_Nv0tesUh2_2;
	wire w_dff_B_7p5YZYKu8_2;
	wire w_dff_B_rsFCvRc05_2;
	wire w_dff_B_E0bbs0sO1_2;
	wire w_dff_B_lcKFYHoU3_2;
	wire w_dff_B_FEx3ty9d0_2;
	wire w_dff_B_bnx2wppo4_2;
	wire w_dff_B_TjKIPwAU4_1;
	wire w_dff_B_FrDCNQQy6_2;
	wire w_dff_B_vyUOjMeo3_2;
	wire w_dff_B_KsKCkddE8_2;
	wire w_dff_B_CSVUpzss6_2;
	wire w_dff_B_FtQPF6pV8_2;
	wire w_dff_B_zBpkpyB48_2;
	wire w_dff_B_tMW2Z0Vc1_2;
	wire w_dff_B_jPvqwdoK4_2;
	wire w_dff_B_xv1nQ7vz8_2;
	wire w_dff_B_TMXlGXGE2_1;
	wire w_dff_B_48mobnWy5_2;
	wire w_dff_B_Q1H5wwwU9_2;
	wire w_dff_B_nGFwCgmu1_2;
	wire w_dff_B_DMvDq34q2_2;
	wire w_dff_B_LuqvSgt21_2;
	wire w_dff_B_BhTaxGEE2_2;
	wire w_dff_B_hzjeHgL23_2;
	wire w_dff_B_H8Nf2bxb9_1;
	wire w_dff_B_8BOK5r7f5_2;
	wire w_dff_B_CxMuwOBI4_2;
	wire w_dff_B_EqHqyi9Y4_2;
	wire w_dff_B_ma8H6lte4_2;
	wire w_dff_B_AxwWbGXe2_2;
	wire w_dff_B_SM2C5eTN2_2;
	wire w_dff_B_B23Uh0Jm4_2;
	wire w_dff_B_IQchRE107_2;
	wire w_dff_B_RtYdSlrb2_0;
	wire w_dff_B_7heOTNru1_0;
	wire w_dff_A_A02n2DW34_0;
	wire w_dff_A_kkCyMRDe5_0;
	wire w_dff_A_D6DhIAUh2_0;
	wire w_dff_A_o1vhWlM35_0;
	wire w_dff_B_pxiAqJRP4_2;
	wire w_dff_B_fmTukOSK5_1;
	wire w_dff_B_Ze2a0qMu3_2;
	wire w_dff_B_YNHysRsW8_2;
	wire w_dff_B_vhuHWw3O6_2;
	wire w_dff_B_jOEJPwI61_2;
	wire w_dff_B_KB4AWD940_2;
	wire w_dff_B_qf5Yo19P0_2;
	wire w_dff_B_INZgAJQT9_2;
	wire w_dff_B_2MB8g3V94_2;
	wire w_dff_B_KiemjYa75_2;
	wire w_dff_B_m531pyuN3_2;
	wire w_dff_B_Nmk57WAB8_2;
	wire w_dff_B_sBmusA4K8_2;
	wire w_dff_B_GA5KIA3m8_2;
	wire w_dff_B_xwOSLHyZ4_2;
	wire w_dff_B_hU9xqo8f2_2;
	wire w_dff_B_mGMsgOJa8_2;
	wire w_dff_B_O3gYNr327_2;
	wire w_dff_B_cNU9WGg78_2;
	wire w_dff_B_4pN8YaBQ7_2;
	wire w_dff_B_AuWUyTAJ2_2;
	wire w_dff_B_WFN8QgVC2_2;
	wire w_dff_B_siZdu26O8_2;
	wire w_dff_B_9GhRiICd4_2;
	wire w_dff_B_zobSXAoj9_2;
	wire w_dff_B_cDE7uDpV1_2;
	wire w_dff_B_en5LGY3f9_2;
	wire w_dff_B_urn32Fvt0_2;
	wire w_dff_B_HAHz5OiS7_2;
	wire w_dff_B_9WiIpf7b4_2;
	wire w_dff_B_N6wxh4pV5_2;
	wire w_dff_B_CnkhAJF62_2;
	wire w_dff_B_RPWS1Gxo0_2;
	wire w_dff_B_Hej4yq6j7_2;
	wire w_dff_B_ovoLQTwy0_2;
	wire w_dff_B_yr9X1Uji1_1;
	wire w_dff_B_6Ig0Wrib6_2;
	wire w_dff_B_sBbrPwaD0_2;
	wire w_dff_B_s9hlSRkh7_2;
	wire w_dff_B_yIeyAk5M5_2;
	wire w_dff_B_9WotExv62_2;
	wire w_dff_B_gMlNety95_2;
	wire w_dff_B_rxj5pdJ56_2;
	wire w_dff_B_ylUgR8Pk1_2;
	wire w_dff_B_Qtva6Esw2_2;
	wire w_dff_B_49h92b0f8_2;
	wire w_dff_B_sCzqxtOy2_2;
	wire w_dff_B_TgGzpvF81_2;
	wire w_dff_B_UKZKDgEx1_2;
	wire w_dff_B_RUCec0kw1_2;
	wire w_dff_B_XuJUKu6A2_2;
	wire w_dff_B_5heccAfs4_2;
	wire w_dff_B_HwNprvhk8_2;
	wire w_dff_B_kfq9iLjj8_2;
	wire w_dff_B_gHajJhX94_2;
	wire w_dff_B_uXsq1X8p9_2;
	wire w_dff_B_veHxe9MD8_2;
	wire w_dff_B_ExQjT2xe0_2;
	wire w_dff_B_KF8C1XD12_2;
	wire w_dff_B_CDI0nxj59_2;
	wire w_dff_B_KDikc2b82_2;
	wire w_dff_B_bTUYfIJx8_2;
	wire w_dff_B_NA27Ky2t1_2;
	wire w_dff_B_qu7Z9csu7_2;
	wire w_dff_B_2ruYm7nD8_2;
	wire w_dff_B_hFHKLx7N3_2;
	wire w_dff_B_fZLq7QUg3_1;
	wire w_dff_B_EJMh1QQl6_2;
	wire w_dff_B_BWgqeZbH8_2;
	wire w_dff_B_bieWKeHu9_2;
	wire w_dff_B_CkQURvXS1_2;
	wire w_dff_B_ePCTChUN6_2;
	wire w_dff_B_810kvt9M8_2;
	wire w_dff_B_1uf4QUqx2_2;
	wire w_dff_B_gGGvKriD3_2;
	wire w_dff_B_KN7D9rK21_2;
	wire w_dff_B_GctTT3680_2;
	wire w_dff_B_DZt5sDHW2_2;
	wire w_dff_B_SBdJTp2B6_2;
	wire w_dff_B_m2tIKxb96_2;
	wire w_dff_B_YIOpxhuX9_2;
	wire w_dff_B_MbeO3Ngk5_2;
	wire w_dff_B_muqdDLpo7_2;
	wire w_dff_B_N6rH1bXL3_2;
	wire w_dff_B_vCumNGsD2_2;
	wire w_dff_B_JidzGYRu2_2;
	wire w_dff_B_dwxKcmGg2_2;
	wire w_dff_B_ahuWJ8uT9_2;
	wire w_dff_B_WfFv4OxZ1_2;
	wire w_dff_B_R0Cp8kF14_2;
	wire w_dff_B_PrHpp7u75_2;
	wire w_dff_B_cMdFCd0j0_2;
	wire w_dff_B_xdppXo9f3_2;
	wire w_dff_B_jSQvbZOs1_2;
	wire w_dff_B_kvmSRX9U9_2;
	wire w_dff_B_Vxbm8uDo5_1;
	wire w_dff_B_p4ZB1WcP1_2;
	wire w_dff_B_DlRZdn8u4_2;
	wire w_dff_B_N1aHqhFc7_2;
	wire w_dff_B_JJ9pVtSQ3_2;
	wire w_dff_B_hfbEGqzB6_2;
	wire w_dff_B_zmdeI1RR2_2;
	wire w_dff_B_OJm5394n6_2;
	wire w_dff_B_rpcW0TBT6_2;
	wire w_dff_B_KJeVeG0Y7_2;
	wire w_dff_B_EVCM8vJY2_2;
	wire w_dff_B_LvW401D86_2;
	wire w_dff_B_nGLDQ6Bm0_2;
	wire w_dff_B_gTY9Q1OR2_2;
	wire w_dff_B_sVh1yYi77_2;
	wire w_dff_B_X7kFy1Ak6_2;
	wire w_dff_B_sTlOQjPh4_2;
	wire w_dff_B_s4HKLGQL7_2;
	wire w_dff_B_wP4T2oEx5_2;
	wire w_dff_B_FKrWEXpt5_2;
	wire w_dff_B_rB8BmRK09_2;
	wire w_dff_B_upOfiIN43_2;
	wire w_dff_B_X8IGTZ6y3_2;
	wire w_dff_B_IF5z1V8o8_2;
	wire w_dff_B_Q1hnPCL74_2;
	wire w_dff_B_Yd3ecm9v4_2;
	wire w_dff_B_vj0XLNQO7_2;
	wire w_dff_B_IgYLrSL78_1;
	wire w_dff_B_5z43T4jN0_2;
	wire w_dff_B_osFMsEJI5_2;
	wire w_dff_B_oaULlXjH1_2;
	wire w_dff_B_kUScHdvo7_2;
	wire w_dff_B_W4eOKzJo8_2;
	wire w_dff_B_0ynQCqX17_2;
	wire w_dff_B_ybum0CE36_2;
	wire w_dff_B_W0s8vepI0_2;
	wire w_dff_B_Jqq5HyYy1_2;
	wire w_dff_B_X6MYm6fk0_2;
	wire w_dff_B_HQn0aSlA1_2;
	wire w_dff_B_botQhHke8_2;
	wire w_dff_B_AJTH37Jc3_2;
	wire w_dff_B_M9ftNkC68_2;
	wire w_dff_B_DCeyKkLr8_2;
	wire w_dff_B_nChQowO27_2;
	wire w_dff_B_XVfgfJ087_2;
	wire w_dff_B_vatxhv1J4_2;
	wire w_dff_B_Mhx8t4Wy6_2;
	wire w_dff_B_GUTVttjz0_2;
	wire w_dff_B_cd3ljYx34_2;
	wire w_dff_B_Xw0xS6fW9_2;
	wire w_dff_B_ZSvXv55q1_2;
	wire w_dff_B_Ur8YsLTJ9_2;
	wire w_dff_B_iZxUeO794_1;
	wire w_dff_B_9cHXJ6xI4_2;
	wire w_dff_B_sHQsWBYe6_2;
	wire w_dff_B_9O5Fk8Eq5_2;
	wire w_dff_B_QM5ycwpm5_2;
	wire w_dff_B_yIE2lwhV0_2;
	wire w_dff_B_J3tXTG7J3_2;
	wire w_dff_B_Fbg5e6d12_2;
	wire w_dff_B_ewcdukZ63_2;
	wire w_dff_B_cCy0cV929_2;
	wire w_dff_B_C3praiYw1_2;
	wire w_dff_B_9DzhZU3b4_2;
	wire w_dff_B_Ay1k8pSE1_2;
	wire w_dff_B_sygk0zuw1_2;
	wire w_dff_B_CxEx6bgT6_2;
	wire w_dff_B_d3lIxQyf4_2;
	wire w_dff_B_4ZWSruHv7_2;
	wire w_dff_B_xO1b3bP35_2;
	wire w_dff_B_DdJNGzU95_2;
	wire w_dff_B_5AbjnurS8_2;
	wire w_dff_B_4y032KLj5_2;
	wire w_dff_B_02o7Fihr9_2;
	wire w_dff_B_0G4BkaBJ6_2;
	wire w_dff_B_kYgnMuZK0_1;
	wire w_dff_B_HBoshp425_2;
	wire w_dff_B_nkw0MnBp6_2;
	wire w_dff_B_fRh20S9b6_2;
	wire w_dff_B_vsnzFCqZ0_2;
	wire w_dff_B_qDvcuv0O4_2;
	wire w_dff_B_JK8jTcXB1_2;
	wire w_dff_B_gKb7bFUd0_2;
	wire w_dff_B_mMyExi168_2;
	wire w_dff_B_uc6FLzr96_2;
	wire w_dff_B_Cw5oPujT1_2;
	wire w_dff_B_zDvQVPR20_2;
	wire w_dff_B_NL9AJev91_2;
	wire w_dff_B_RKhk3fWy1_2;
	wire w_dff_B_3Uosf91N7_2;
	wire w_dff_B_cUKRWuIn6_2;
	wire w_dff_B_MfjPzDl48_2;
	wire w_dff_B_6yAjG21H0_2;
	wire w_dff_B_0qJcRvyU2_2;
	wire w_dff_B_F7WlKSiL1_2;
	wire w_dff_B_Ja40IbTs7_2;
	wire w_dff_B_EzN5P6Er8_1;
	wire w_dff_B_WXFOOucF5_2;
	wire w_dff_B_wavBGGTY4_2;
	wire w_dff_B_rBodl2Rl4_2;
	wire w_dff_B_yjVaAvJd5_2;
	wire w_dff_B_p7n8aCKs6_2;
	wire w_dff_B_FBVDvcvc4_2;
	wire w_dff_B_RigZRfyr4_2;
	wire w_dff_B_TcRFPIOC3_2;
	wire w_dff_B_AfJC8Fe28_2;
	wire w_dff_B_sqLUfVGh3_2;
	wire w_dff_B_szrtYhym2_2;
	wire w_dff_B_ZGLPVILf7_2;
	wire w_dff_B_Ic8f7Rbe8_2;
	wire w_dff_B_VJQ29aMe2_2;
	wire w_dff_B_yik2uola1_2;
	wire w_dff_B_sApg5KCq0_2;
	wire w_dff_B_wxNgrRG15_2;
	wire w_dff_B_dGoD1wjK8_2;
	wire w_dff_B_2Ytn0KlC5_1;
	wire w_dff_B_wQeodYbi4_2;
	wire w_dff_B_WTx0HzLt9_2;
	wire w_dff_B_OzfKQF338_2;
	wire w_dff_B_aSKDJZTm6_2;
	wire w_dff_B_YLyfWVB10_2;
	wire w_dff_B_IPgcPpcI5_2;
	wire w_dff_B_P6X41ltl8_2;
	wire w_dff_B_rzKKLRbA1_2;
	wire w_dff_B_wmkluPFv3_2;
	wire w_dff_B_zY3c43w38_2;
	wire w_dff_B_EyvNzULS8_2;
	wire w_dff_B_GeqNlMIE0_2;
	wire w_dff_B_R0ZR6iCs3_2;
	wire w_dff_B_ULEgfoCS9_2;
	wire w_dff_B_nAuwTMlj1_2;
	wire w_dff_B_r65m0gHm0_2;
	wire w_dff_B_tc797yZk2_1;
	wire w_dff_B_SLa7yIMe6_2;
	wire w_dff_B_MjdljAZ27_2;
	wire w_dff_B_T9xnokmU6_2;
	wire w_dff_B_RsNr5UGG1_2;
	wire w_dff_B_SaLhkhMA3_2;
	wire w_dff_B_kBQ8eeqa9_2;
	wire w_dff_B_H22V1JKQ9_2;
	wire w_dff_B_7eeRBTvC4_2;
	wire w_dff_B_FONr2Ja70_2;
	wire w_dff_B_PF6eVLh83_2;
	wire w_dff_B_WlMjQp025_2;
	wire w_dff_B_cJwP2DIY5_2;
	wire w_dff_B_L1DTu0oL3_2;
	wire w_dff_B_1MUQayca2_2;
	wire w_dff_B_ZtbhKuhs5_2;
	wire w_dff_B_ajzQoUT25_2;
	wire w_dff_B_M9Ywdoct1_2;
	wire w_dff_B_4ZkH0V4J4_1;
	wire w_dff_B_4wZV470f8_2;
	wire w_dff_B_93m99Vn68_2;
	wire w_dff_B_c70jGVwM6_2;
	wire w_dff_B_9bfqCtGY2_2;
	wire w_dff_B_XrNXuaAF4_2;
	wire w_dff_B_HTD27yKz0_2;
	wire w_dff_B_MkPgHLIU9_2;
	wire w_dff_B_SkejRnpn0_2;
	wire w_dff_B_4Dj13Jvy2_2;
	wire w_dff_B_OsDt93ur4_1;
	wire w_dff_B_8VvdAJ4d8_2;
	wire w_dff_B_JltM7ZGy5_2;
	wire w_dff_B_aJGVUg9q7_2;
	wire w_dff_B_3juZpKTG2_2;
	wire w_dff_B_qgUAGqRV7_2;
	wire w_dff_B_z7lCqZki2_2;
	wire w_dff_B_dbs0Nf4r4_2;
	wire w_dff_B_Z0Y6Bzw53_1;
	wire w_dff_B_TkU64rgP2_2;
	wire w_dff_B_jvU8bwhf6_2;
	wire w_dff_B_TQSGHHTO7_2;
	wire w_dff_B_Dv1DFU4c7_2;
	wire w_dff_B_2vHWrEiA8_2;
	wire w_dff_B_3i3vPdau4_2;
	wire w_dff_B_rjgJwLKB0_2;
	wire w_dff_B_cbd2tEGR6_2;
	wire w_dff_B_AJL1rbdl4_0;
	wire w_dff_B_wD40bFgi9_0;
	wire w_dff_A_820aAthH5_0;
	wire w_dff_A_VFk9IOOo6_0;
	wire w_dff_A_RJf1Y65M4_0;
	wire w_dff_A_lXNE1JWt6_0;
	wire w_dff_B_2s9dHElE5_2;
	wire w_dff_B_X5KheESI6_2;
	wire w_dff_B_pruoaOri4_1;
	wire w_dff_B_jfR6X47k4_2;
	wire w_dff_B_S6g40pB57_2;
	wire w_dff_B_egYGi1Od2_2;
	wire w_dff_B_j2jZ3IJz0_2;
	wire w_dff_B_pg1SXlAp3_2;
	wire w_dff_B_zZ3ICMPW7_2;
	wire w_dff_B_wNnTB0qN1_2;
	wire w_dff_B_YkCeicYp4_2;
	wire w_dff_B_nhXQ1pFN1_2;
	wire w_dff_B_FDa1bFrG2_2;
	wire w_dff_B_KerW6clm1_2;
	wire w_dff_B_HIzLqiIZ4_2;
	wire w_dff_B_47Yn0VEd5_2;
	wire w_dff_B_6WAwCxhE8_2;
	wire w_dff_B_yzTges2q8_2;
	wire w_dff_B_yLXEaxdp0_2;
	wire w_dff_B_0ZxJP1fF8_2;
	wire w_dff_B_jaGU8V821_2;
	wire w_dff_B_C7ykZp4v7_2;
	wire w_dff_B_N3dAI3l63_2;
	wire w_dff_B_oY7ajPEx9_2;
	wire w_dff_B_rfZ8eDUg8_2;
	wire w_dff_B_uNHoWAuO3_2;
	wire w_dff_B_JKbuB6Mc2_2;
	wire w_dff_B_MYCLVb5o7_2;
	wire w_dff_B_aWeAeoS14_2;
	wire w_dff_B_fEu038fv1_2;
	wire w_dff_B_2JtvUI9V8_2;
	wire w_dff_B_VIa1jW1B9_2;
	wire w_dff_B_cDG4JfW54_2;
	wire w_dff_B_qGzVz2qc0_2;
	wire w_dff_B_VAvZLqhF2_2;
	wire w_dff_B_pgCfMrz43_2;
	wire w_dff_B_khNyTxgR1_2;
	wire w_dff_B_v3VgPoVA6_1;
	wire w_dff_B_IhY0Ds3Z3_2;
	wire w_dff_B_LjXWS6AA4_2;
	wire w_dff_B_JBSmMM8z3_2;
	wire w_dff_B_iBL2XGxJ0_2;
	wire w_dff_B_JMwULktA3_2;
	wire w_dff_B_RbmOlHMq9_2;
	wire w_dff_B_3yGlt62V6_2;
	wire w_dff_B_WxdKZAMv8_2;
	wire w_dff_B_MGBRD87w4_2;
	wire w_dff_B_XHs01P0X9_2;
	wire w_dff_B_qOayNJGz0_2;
	wire w_dff_B_BYuex7We0_2;
	wire w_dff_B_DmutNhWQ5_2;
	wire w_dff_B_F6OMPAFq7_2;
	wire w_dff_B_1RU4xIcQ4_2;
	wire w_dff_B_Zw3rbi1D3_2;
	wire w_dff_B_N7wWm7Uv0_2;
	wire w_dff_B_SZxqN9x08_2;
	wire w_dff_B_gR8OEe0h9_2;
	wire w_dff_B_eptCr87L8_2;
	wire w_dff_B_ma5NMSMI8_2;
	wire w_dff_B_njf8lLwo7_2;
	wire w_dff_B_MwvA4mZl4_2;
	wire w_dff_B_T5KgOxh74_2;
	wire w_dff_B_JX8pf6I34_2;
	wire w_dff_B_NqqxYUqI2_2;
	wire w_dff_B_FcjemT152_2;
	wire w_dff_B_AyQ9YqEA4_2;
	wire w_dff_B_zE7LPmHe3_2;
	wire w_dff_B_9iVFdk5t0_2;
	wire w_dff_B_QxnkdtK96_1;
	wire w_dff_B_xu18Wgd63_2;
	wire w_dff_B_SHi9O1wl0_2;
	wire w_dff_B_dhZIFRH02_2;
	wire w_dff_B_zwdWLX4l7_2;
	wire w_dff_B_HZ6uSPBh5_2;
	wire w_dff_B_oyBnS3GN8_2;
	wire w_dff_B_EUfySKTj9_2;
	wire w_dff_B_QxWT93uW6_2;
	wire w_dff_B_BdxFdJig0_2;
	wire w_dff_B_BNMW6Qob3_2;
	wire w_dff_B_LMW1Qgr25_2;
	wire w_dff_B_8pAhwc8G5_2;
	wire w_dff_B_hwozoBNM7_2;
	wire w_dff_B_zjNoWVwV1_2;
	wire w_dff_B_1fZK6CUp9_2;
	wire w_dff_B_Xm3JAaOh8_2;
	wire w_dff_B_ELlgVvUu7_2;
	wire w_dff_B_VBEBz7i95_2;
	wire w_dff_B_QEwiVNKB8_2;
	wire w_dff_B_EWohVFEg1_2;
	wire w_dff_B_3cujJYnU6_2;
	wire w_dff_B_dPyV0SGM2_2;
	wire w_dff_B_bVblJ1rf2_2;
	wire w_dff_B_5zbpitpD2_2;
	wire w_dff_B_74hQK1698_2;
	wire w_dff_B_k8cmLbAc7_2;
	wire w_dff_B_SrPYwD194_2;
	wire w_dff_B_LE4azKlA7_2;
	wire w_dff_B_ygGrrKsO1_1;
	wire w_dff_B_PnsullEO7_2;
	wire w_dff_B_Afhpwo7d3_2;
	wire w_dff_B_EKWG8set4_2;
	wire w_dff_B_O0EhHbYA9_2;
	wire w_dff_B_3V7ZAs4h9_2;
	wire w_dff_B_gtNfPWEz4_2;
	wire w_dff_B_FajFmzDy5_2;
	wire w_dff_B_vaVMa4NS6_2;
	wire w_dff_B_0YTtw7uS3_2;
	wire w_dff_B_jSTZrvy77_2;
	wire w_dff_B_yXsl5EKu5_2;
	wire w_dff_B_Q38pz4Jj3_2;
	wire w_dff_B_k0C6hbO88_2;
	wire w_dff_B_94O8dSav2_2;
	wire w_dff_B_GIkOKykb1_2;
	wire w_dff_B_lUfXqXAW7_2;
	wire w_dff_B_g7poNg7U3_2;
	wire w_dff_B_D5Y9i9q60_2;
	wire w_dff_B_EAOmlf739_2;
	wire w_dff_B_WLAcfqAC3_2;
	wire w_dff_B_PQB1mG6v1_2;
	wire w_dff_B_1RyHKKb59_2;
	wire w_dff_B_yKyGVzaj1_2;
	wire w_dff_B_DO9CrTUn1_2;
	wire w_dff_B_F3mr18MV6_2;
	wire w_dff_B_FeoLRdE16_2;
	wire w_dff_B_ED789YdO5_1;
	wire w_dff_B_stRJSPrO4_2;
	wire w_dff_B_uPCsLQqt9_2;
	wire w_dff_B_L7yLjOHe3_2;
	wire w_dff_B_kORukNq40_2;
	wire w_dff_B_1aKtioxn2_2;
	wire w_dff_B_UQNsoet96_2;
	wire w_dff_B_FWI24CPp1_2;
	wire w_dff_B_73oC28Ih7_2;
	wire w_dff_B_lRSgbmKP0_2;
	wire w_dff_B_x7hLgs4Y7_2;
	wire w_dff_B_d0ejrO6m1_2;
	wire w_dff_B_n25tirG72_2;
	wire w_dff_B_3FwuhAIb7_2;
	wire w_dff_B_Y0w0qHtz0_2;
	wire w_dff_B_PLRcf1md5_2;
	wire w_dff_B_yZH4XOE43_2;
	wire w_dff_B_CPSSX6F10_2;
	wire w_dff_B_bLZpHZRw5_2;
	wire w_dff_B_B2LPLQhR1_2;
	wire w_dff_B_NPNT7YiW8_2;
	wire w_dff_B_UPX9w7Ht8_2;
	wire w_dff_B_sPsAxl123_2;
	wire w_dff_B_Ria118Gd0_2;
	wire w_dff_B_PBlOLn9W3_2;
	wire w_dff_B_FgdnHYwK2_1;
	wire w_dff_B_ekgEtoUO2_2;
	wire w_dff_B_sYKDkzLF9_2;
	wire w_dff_B_Tr3LEl8r5_2;
	wire w_dff_B_zEK7cFsf1_2;
	wire w_dff_B_GfRMrhS61_2;
	wire w_dff_B_2FZCjvbg1_2;
	wire w_dff_B_XlyqA1IH5_2;
	wire w_dff_B_xP8AtX5Z5_2;
	wire w_dff_B_2yvGR2Ek1_2;
	wire w_dff_B_b1V6jxak8_2;
	wire w_dff_B_gN3pGbps7_2;
	wire w_dff_B_4BxoFDyC1_2;
	wire w_dff_B_O3PoVkvw4_2;
	wire w_dff_B_TVGJSBX56_2;
	wire w_dff_B_xtK5Rbih5_2;
	wire w_dff_B_3nCiWTnS1_2;
	wire w_dff_B_0NtUjsPQ1_2;
	wire w_dff_B_gjnnWyRi4_2;
	wire w_dff_B_h3n7iEUg1_2;
	wire w_dff_B_pMhNgscN4_2;
	wire w_dff_B_e0HsKxQf0_2;
	wire w_dff_B_mWheOF5C7_2;
	wire w_dff_B_q1b7ahO29_1;
	wire w_dff_B_veTLb8Vs8_2;
	wire w_dff_B_0ahfb7oG5_2;
	wire w_dff_B_dGm8vyB83_2;
	wire w_dff_B_fjUzNIqj5_2;
	wire w_dff_B_EL1xu06P2_2;
	wire w_dff_B_aSOYuojn0_2;
	wire w_dff_B_CZEOpvFt0_2;
	wire w_dff_B_E8omsfOG9_2;
	wire w_dff_B_18ffRcbz4_2;
	wire w_dff_B_uDT9w2XC3_2;
	wire w_dff_B_2M3DeORd4_2;
	wire w_dff_B_a0dAQvqn7_2;
	wire w_dff_B_SCiFj1xc9_2;
	wire w_dff_B_C36nM2X15_2;
	wire w_dff_B_NBsocNKy7_2;
	wire w_dff_B_8xdLxR9I9_2;
	wire w_dff_B_iP887MlT9_2;
	wire w_dff_B_3500toN99_2;
	wire w_dff_B_4ShIlRBK3_2;
	wire w_dff_B_vZt4kRgy3_2;
	wire w_dff_B_LVoVRGms8_1;
	wire w_dff_B_ClMo1ysm3_2;
	wire w_dff_B_uwuJcj5Z0_2;
	wire w_dff_B_r6WN8Ujm1_2;
	wire w_dff_B_q8VNmquh5_2;
	wire w_dff_B_umMJzL4H4_2;
	wire w_dff_B_qycJlDXy4_2;
	wire w_dff_B_8PxiXb4f7_2;
	wire w_dff_B_XELB2PkE5_2;
	wire w_dff_B_1OP0kEfm1_2;
	wire w_dff_B_l2VlOEbG5_2;
	wire w_dff_B_JE0GkGB96_2;
	wire w_dff_B_DwyTfFK09_2;
	wire w_dff_B_pxSpR05y1_2;
	wire w_dff_B_IN0dtKW29_2;
	wire w_dff_B_dm9LOI3q5_2;
	wire w_dff_B_i7FjBT1X6_2;
	wire w_dff_B_ZNGfFnnu0_2;
	wire w_dff_B_KJsm2iQ82_2;
	wire w_dff_B_4XFcQDTb2_1;
	wire w_dff_B_akRh96m98_2;
	wire w_dff_B_o3Hb8qRl9_2;
	wire w_dff_B_MdL5x2Um9_2;
	wire w_dff_B_iIuAZHJe0_2;
	wire w_dff_B_8nc1XJGJ6_2;
	wire w_dff_B_PW6VcZAH8_2;
	wire w_dff_B_wXTODCum4_2;
	wire w_dff_B_lT0uklDO9_2;
	wire w_dff_B_aVXoJ7u48_2;
	wire w_dff_B_VFC9A23N0_2;
	wire w_dff_B_T7RaTU3C0_2;
	wire w_dff_B_t8m4j8xr8_2;
	wire w_dff_B_Z4wJxIY12_2;
	wire w_dff_B_rruH8tJ20_2;
	wire w_dff_B_3zrRElB43_2;
	wire w_dff_B_xLVoL2A89_2;
	wire w_dff_B_EeRAn82r9_1;
	wire w_dff_B_7AI4Njhh6_2;
	wire w_dff_B_CREJbewt6_2;
	wire w_dff_B_aDc2gZMo1_2;
	wire w_dff_B_XGxtZviB5_2;
	wire w_dff_B_YZDPIdx77_2;
	wire w_dff_B_qoXoW2Br7_2;
	wire w_dff_B_nbGLUgVs8_2;
	wire w_dff_B_dvJqJAoi4_2;
	wire w_dff_B_O9G2zr9x4_2;
	wire w_dff_B_QMQyzwLw5_2;
	wire w_dff_B_2VWYOpj38_2;
	wire w_dff_B_Z1cr4aXq6_2;
	wire w_dff_B_JJeV97Np3_2;
	wire w_dff_B_tm99xvrP5_2;
	wire w_dff_B_t8UKOF9J6_1;
	wire w_dff_B_vmfqcjdR1_2;
	wire w_dff_B_zuHONWuS5_2;
	wire w_dff_B_Y8Ptgm9C0_2;
	wire w_dff_B_7CQ2v9EO7_2;
	wire w_dff_B_NLty3pQN6_2;
	wire w_dff_B_D8wmpClN2_2;
	wire w_dff_B_qJWLIZBO5_2;
	wire w_dff_B_AuvRTLi49_2;
	wire w_dff_B_wKwhIiQR9_2;
	wire w_dff_B_6LQjZsdB1_2;
	wire w_dff_B_Kj84ly7A4_2;
	wire w_dff_B_n8pcLXAT9_2;
	wire w_dff_B_QovX8Hk43_2;
	wire w_dff_B_GqB6oQRN9_2;
	wire w_dff_B_yFFnSilg5_2;
	wire w_dff_B_FvN6rCQc2_1;
	wire w_dff_B_cJDKDu5i9_2;
	wire w_dff_B_N14UW4li6_2;
	wire w_dff_B_3tCyqfK11_2;
	wire w_dff_B_v594jcT89_2;
	wire w_dff_B_jqC0T3Ib6_2;
	wire w_dff_B_ESlMcoRT9_2;
	wire w_dff_B_teCrdQ8K5_2;
	wire w_dff_B_JkEj9UbZ8_1;
	wire w_dff_B_i9xW1p9e3_2;
	wire w_dff_B_ZU1jIcRx3_2;
	wire w_dff_B_Pxtf12Fd3_2;
	wire w_dff_B_9JcfT8IA9_2;
	wire w_dff_B_ZXoeUWOj6_2;
	wire w_dff_B_7uz8IcC05_1;
	wire w_dff_B_YGy5Ezsl9_2;
	wire w_dff_B_x7IpbgK77_2;
	wire w_dff_B_IBrwA5D33_2;
	wire w_dff_B_wZMqDuih9_0;
	wire w_dff_B_VTHvwSX19_0;
	wire w_dff_A_retMBguq4_0;
	wire w_dff_A_hY78nFfS1_0;
	wire w_dff_A_xMoJ7StT8_1;
	wire w_dff_A_TMMq93Z77_1;
	wire w_dff_B_hU1vr8NB2_2;
	wire w_dff_B_w0qqjdMw7_2;
	wire w_dff_B_GKM8K4XL9_1;
	wire w_dff_B_maUi0Lzd7_2;
	wire w_dff_B_CxSPndrc1_2;
	wire w_dff_B_MhLCBSzF3_2;
	wire w_dff_B_a3dxtBr67_2;
	wire w_dff_B_8iSvPxTB5_2;
	wire w_dff_B_Ke6b32sX7_2;
	wire w_dff_B_1ExOcTyq1_2;
	wire w_dff_B_lgF1Qhfv7_2;
	wire w_dff_B_CGgVJdRW9_2;
	wire w_dff_B_PC55rC5Q2_2;
	wire w_dff_B_laNg1s5u2_2;
	wire w_dff_B_ek8eaccx1_2;
	wire w_dff_B_0boWsVUu9_2;
	wire w_dff_B_ifydVLx50_2;
	wire w_dff_B_bn7Bp5YP4_2;
	wire w_dff_B_IXmGDbx54_2;
	wire w_dff_B_5xAWax9B8_2;
	wire w_dff_B_KYHpEjRR4_2;
	wire w_dff_B_v8rEyMCD7_2;
	wire w_dff_B_wZvVc4L84_2;
	wire w_dff_B_3p9SAWRY2_2;
	wire w_dff_B_44dBfwXj8_2;
	wire w_dff_B_eILm0Hdd1_2;
	wire w_dff_B_SRB1jn3r4_2;
	wire w_dff_B_aMk3RGb47_2;
	wire w_dff_B_XIZvnHZf6_2;
	wire w_dff_B_1Bf0ttZE9_2;
	wire w_dff_B_mMW3aN4X6_2;
	wire w_dff_B_X85fratI2_2;
	wire w_dff_B_cqtq7KrZ3_2;
	wire w_dff_B_qkPFyqNd2_2;
	wire w_dff_B_uFiUg5zk1_2;
	wire w_dff_B_qQayyI4N9_2;
	wire w_dff_B_aSVJu1OY1_2;
	wire w_dff_B_PX4TXQFr3_2;
	wire w_dff_B_wYs9wv6H6_1;
	wire w_dff_A_cnLtIaDT5_1;
	wire w_dff_B_7bDJzS977_1;
	wire w_dff_B_wA5Gw0z84_2;
	wire w_dff_B_tMRehM009_2;
	wire w_dff_B_QPVHrLSu8_2;
	wire w_dff_B_poLOfYC04_2;
	wire w_dff_B_0TgQrXSf8_2;
	wire w_dff_B_WSVDKpfw1_2;
	wire w_dff_B_pAB45IqW3_2;
	wire w_dff_B_DSXpFfIh4_2;
	wire w_dff_B_TcuTRza81_2;
	wire w_dff_B_8aLhlURf9_2;
	wire w_dff_B_D7hHXQoh1_2;
	wire w_dff_B_Xv3tLuEo5_2;
	wire w_dff_B_orABP4fh7_2;
	wire w_dff_B_c9uSD6N01_2;
	wire w_dff_B_sdaqmCrV9_2;
	wire w_dff_B_pCkqAd235_2;
	wire w_dff_B_yUGJ1ABx7_2;
	wire w_dff_B_fHjw4xR85_2;
	wire w_dff_B_G9DlWunn7_2;
	wire w_dff_B_8ENxcvDx1_2;
	wire w_dff_B_UCLLO6K79_2;
	wire w_dff_B_F7Dp79Zo8_2;
	wire w_dff_B_Mk1Rz2mV3_2;
	wire w_dff_B_4cB1IIUp4_2;
	wire w_dff_B_V0wGUUrE2_2;
	wire w_dff_B_1DWqglps3_2;
	wire w_dff_B_NBvfBKSV9_2;
	wire w_dff_B_Vl22xVyp0_2;
	wire w_dff_B_nE2JIBPd8_2;
	wire w_dff_B_Mmu3qViy6_2;
	wire w_dff_B_RaRq5BB64_1;
	wire w_dff_B_jKS1znAl9_2;
	wire w_dff_B_IEldEdry3_2;
	wire w_dff_B_Wj2RZUHn7_2;
	wire w_dff_B_QOutNQxk7_2;
	wire w_dff_B_qgEb6KPh5_2;
	wire w_dff_B_enKxK3UM9_2;
	wire w_dff_B_8shtw70R2_2;
	wire w_dff_B_7fEHJGDL2_2;
	wire w_dff_B_qL08NAw01_2;
	wire w_dff_B_lT2NR7956_2;
	wire w_dff_B_H7hFTxHI7_2;
	wire w_dff_B_3KgJDtrk7_2;
	wire w_dff_B_ei8Sv0aK9_2;
	wire w_dff_B_jLu3wO3D8_2;
	wire w_dff_B_88Jx1Ykp3_2;
	wire w_dff_B_wvY57nQ62_2;
	wire w_dff_B_f5sIsrsv0_2;
	wire w_dff_B_QWY6R8Vv9_2;
	wire w_dff_B_iWuvyW2L8_2;
	wire w_dff_B_NtXmSGFY4_2;
	wire w_dff_B_mqC9gCbc5_2;
	wire w_dff_B_AJzHeA9K2_2;
	wire w_dff_B_MsKbgqrm1_2;
	wire w_dff_B_kWsbnAtx5_2;
	wire w_dff_B_jOB8gM1P1_2;
	wire w_dff_B_t5TkYjdu0_2;
	wire w_dff_B_u2C2UcnT0_2;
	wire w_dff_B_aNHEh6ZZ6_2;
	wire w_dff_B_Bd7910S22_1;
	wire w_dff_B_rrQgZzuG4_2;
	wire w_dff_B_pNIrZEG52_2;
	wire w_dff_B_LmDPB5aO5_2;
	wire w_dff_B_l5cg6R4B3_2;
	wire w_dff_B_zEAcGAwa4_2;
	wire w_dff_B_EupCZzFA2_2;
	wire w_dff_B_bQA6PJ652_2;
	wire w_dff_B_szrSiuWW1_2;
	wire w_dff_B_CGZlUZlS5_2;
	wire w_dff_B_HWsTwFSJ4_2;
	wire w_dff_B_h4WKwM6k2_2;
	wire w_dff_B_QgBNUGeA0_2;
	wire w_dff_B_SFD9oYE37_2;
	wire w_dff_B_8Zvk0iYL0_2;
	wire w_dff_B_zfekEoYl2_2;
	wire w_dff_B_HVBRvyDV0_2;
	wire w_dff_B_XeOabcEj5_2;
	wire w_dff_B_xFfop47F0_2;
	wire w_dff_B_Pnt7yk0J9_2;
	wire w_dff_B_7IzkV9ix1_2;
	wire w_dff_B_7ClHIuDo8_2;
	wire w_dff_B_bEO3POAo6_2;
	wire w_dff_B_Y9AFkIhl3_2;
	wire w_dff_B_YaQADm9V9_2;
	wire w_dff_B_Ew6GQxoc6_2;
	wire w_dff_B_DuRkClK69_2;
	wire w_dff_B_Mufn57ny6_1;
	wire w_dff_B_Ahh1psqS6_2;
	wire w_dff_B_ut37sD9P3_2;
	wire w_dff_B_q1BTJUjT5_2;
	wire w_dff_B_KTOszVOS9_2;
	wire w_dff_B_31q72oRG8_2;
	wire w_dff_B_M6EiS9eb5_2;
	wire w_dff_B_Ym9cUVec8_2;
	wire w_dff_B_wrd8rwdu6_2;
	wire w_dff_B_UPwZxG364_2;
	wire w_dff_B_C1B0sqnh7_2;
	wire w_dff_B_VF1RJEtp6_2;
	wire w_dff_B_swQSk3Ee8_2;
	wire w_dff_B_9a7cZNhN7_2;
	wire w_dff_B_SpWeiUL30_2;
	wire w_dff_B_8Yk8pSXQ5_2;
	wire w_dff_B_pJbpBqgm0_2;
	wire w_dff_B_YG6VkVdh7_2;
	wire w_dff_B_6HM1VqsS9_2;
	wire w_dff_B_14u4atyu2_2;
	wire w_dff_B_N3EFo4EA1_2;
	wire w_dff_B_e4zhWBgy9_2;
	wire w_dff_B_AEMtq3kd1_2;
	wire w_dff_B_aILTKOZt6_2;
	wire w_dff_B_i0Ted2BP2_2;
	wire w_dff_B_f7L6yJwE3_1;
	wire w_dff_B_b4J6Jsjq1_2;
	wire w_dff_B_P9SHxo5I4_2;
	wire w_dff_B_xLzQOyvP1_2;
	wire w_dff_B_yQUxV8S49_2;
	wire w_dff_B_FufbPb9v3_2;
	wire w_dff_B_CE8s2ibK8_2;
	wire w_dff_B_pmOtB5Vt7_2;
	wire w_dff_B_YwrX7H9T5_2;
	wire w_dff_B_GBzN1GgS7_2;
	wire w_dff_B_oTD8YeAJ6_2;
	wire w_dff_B_X1DeDsWc9_2;
	wire w_dff_B_fK9SMo8Y2_2;
	wire w_dff_B_fdMk5D4N6_2;
	wire w_dff_B_ZPHrhZsx2_2;
	wire w_dff_B_tGvA40Y17_2;
	wire w_dff_B_6X0smcHS3_2;
	wire w_dff_B_6qx6EC9Z1_2;
	wire w_dff_B_fU6iMUOy2_2;
	wire w_dff_B_74MAd6Bm5_2;
	wire w_dff_B_jId4Xbgr3_2;
	wire w_dff_B_zSWeITEe6_2;
	wire w_dff_B_RV3WkNZc5_2;
	wire w_dff_B_UA07Ppi04_1;
	wire w_dff_B_mLuleuuW0_2;
	wire w_dff_B_3HVmoRH91_2;
	wire w_dff_B_v24TIdmq9_2;
	wire w_dff_B_UiqP8xR29_2;
	wire w_dff_B_qE3SrZhB1_2;
	wire w_dff_B_SeiPQxnU4_2;
	wire w_dff_B_ab8tWZ0k3_2;
	wire w_dff_B_TC7iGZl78_2;
	wire w_dff_B_Z4Mvbzdo8_2;
	wire w_dff_B_W2zLnZtg9_2;
	wire w_dff_B_Lm9SP8yb6_2;
	wire w_dff_B_Vx26dSJb3_2;
	wire w_dff_B_RfERzzQF0_2;
	wire w_dff_B_dSeTHEyi8_2;
	wire w_dff_B_OWVazIu22_2;
	wire w_dff_B_gqlFadwb0_2;
	wire w_dff_B_px9xqlZb8_2;
	wire w_dff_B_8il9FhlR3_2;
	wire w_dff_B_MHn3v5bm5_2;
	wire w_dff_B_46mVB41B0_2;
	wire w_dff_B_MJOCAlLn4_1;
	wire w_dff_B_YlTZMmhF9_2;
	wire w_dff_B_BQBdGkrS6_2;
	wire w_dff_B_kV6mGeTN8_2;
	wire w_dff_B_juG7tBaw2_2;
	wire w_dff_B_wSYNEC4s3_2;
	wire w_dff_B_pwQUszuN1_2;
	wire w_dff_B_vHuksEov3_2;
	wire w_dff_B_3RSOZf3m2_2;
	wire w_dff_B_d2Nh74uB8_2;
	wire w_dff_B_XiXhp0LZ6_2;
	wire w_dff_B_QmdtSoxt5_2;
	wire w_dff_B_q0LHuPxt9_2;
	wire w_dff_B_boZKUdGN0_2;
	wire w_dff_B_ZXwtNYIJ0_2;
	wire w_dff_B_LXUXNYAJ1_2;
	wire w_dff_B_DeZzbMYc2_2;
	wire w_dff_B_WdGtINt84_2;
	wire w_dff_B_FAqUrTuV1_2;
	wire w_dff_B_eQvYoeCl6_1;
	wire w_dff_B_LE9eh2jq5_2;
	wire w_dff_B_S9YSBhFz2_2;
	wire w_dff_B_rfL8FXnI9_2;
	wire w_dff_B_93mCKM6Z4_2;
	wire w_dff_B_WghgYMo79_2;
	wire w_dff_B_00wZDapF8_2;
	wire w_dff_B_6Wtocq1f8_2;
	wire w_dff_B_ZqZ3KqWL5_2;
	wire w_dff_B_dH851IKM2_2;
	wire w_dff_B_FdMleJGZ8_2;
	wire w_dff_B_e1yJGDxr3_2;
	wire w_dff_B_7JXVf2JF2_2;
	wire w_dff_B_AQ1RrBGH6_2;
	wire w_dff_B_gMhffUhg5_2;
	wire w_dff_B_sWMeyzD53_2;
	wire w_dff_B_nQgUO1Pw2_2;
	wire w_dff_B_1P0ORXtM0_1;
	wire w_dff_B_7Tyh0ggS9_2;
	wire w_dff_B_KFHZ1Yb21_2;
	wire w_dff_B_ir9JsQlc5_2;
	wire w_dff_B_h9KxhMIl9_2;
	wire w_dff_B_G7Yk4JN51_2;
	wire w_dff_B_80vnigy17_2;
	wire w_dff_B_82JXgsKz1_2;
	wire w_dff_B_r0Xe9xzX9_2;
	wire w_dff_B_WcjxHfu34_2;
	wire w_dff_B_vtc9D6FF4_2;
	wire w_dff_B_mbeeLv1B3_2;
	wire w_dff_B_CIkdsVH92_2;
	wire w_dff_B_YxTpVFRc4_2;
	wire w_dff_B_9aOUgWIu3_2;
	wire w_dff_B_Y3iWifio0_1;
	wire w_dff_B_tYY4aaKe3_2;
	wire w_dff_B_wnadlOra2_2;
	wire w_dff_B_c8nsEbdb6_2;
	wire w_dff_B_kR158B877_2;
	wire w_dff_B_fUrG5sDI8_2;
	wire w_dff_B_JP2hJyNA1_2;
	wire w_dff_B_ZHVSF9JX1_2;
	wire w_dff_B_XUi64OdK7_2;
	wire w_dff_B_inSMvfMl8_2;
	wire w_dff_B_s5ZoFUJN4_2;
	wire w_dff_B_I31Na36j0_2;
	wire w_dff_B_W0AeNeTW6_2;
	wire w_dff_B_0ttUigoW2_1;
	wire w_dff_B_tutDU4Of6_2;
	wire w_dff_B_62YYaDSn3_2;
	wire w_dff_B_YRIm5N3Z8_2;
	wire w_dff_B_GVrHlklT3_2;
	wire w_dff_B_ub2s6Tib8_2;
	wire w_dff_B_Hah5zG2R3_2;
	wire w_dff_B_th4CQD6f5_2;
	wire w_dff_B_nyjW9aRJ9_2;
	wire w_dff_B_txcvjfHr9_2;
	wire w_dff_B_VdCinP0T1_2;
	wire w_dff_B_2eyN18HJ6_2;
	wire w_dff_B_Kf2vFNnD5_2;
	wire w_dff_B_RodJbxBX1_2;
	wire w_dff_B_aklalK3q6_1;
	wire w_dff_B_b58sizGw8_2;
	wire w_dff_B_puJmDR174_2;
	wire w_dff_B_fD4v50RS7_2;
	wire w_dff_B_dKdNc2dK3_2;
	wire w_dff_B_xso4Npzq4_2;
	wire w_dff_B_ZYD8hTSh7_1;
	wire w_dff_B_SbNQ4RCr9_2;
	wire w_dff_B_lJQVzpmo9_2;
	wire w_dff_B_1jyfj3PW8_2;
	wire w_dff_B_Q2Fswjgg1_0;
	wire w_dff_B_DIG1ikH87_0;
	wire w_dff_A_ZDNfXdBN8_0;
	wire w_dff_A_D70Zf41k4_0;
	wire w_dff_A_fsvH5Wdk4_1;
	wire w_dff_A_8uBIIrPF3_1;
	wire w_dff_B_ECy4dX4h6_2;
	wire w_dff_B_WFe17quy4_2;
	wire w_dff_B_ZIvl7ino7_1;
	wire w_dff_B_BEz0cK1R0_2;
	wire w_dff_B_M7MyesCO6_2;
	wire w_dff_B_RwZlw2uP8_2;
	wire w_dff_B_ZFfcxAnt4_2;
	wire w_dff_B_5ipsmv8G1_2;
	wire w_dff_B_lsj78i6I6_2;
	wire w_dff_B_wTpE2uP61_2;
	wire w_dff_B_Hk8JWjcv9_2;
	wire w_dff_B_Ge34LjSF4_2;
	wire w_dff_B_kodSHwjr0_2;
	wire w_dff_B_MVIxVjYi0_2;
	wire w_dff_B_Bp60VGvQ3_2;
	wire w_dff_B_mdOdkvQp7_2;
	wire w_dff_B_VMlaPO3N0_2;
	wire w_dff_B_TbibVkUy8_2;
	wire w_dff_B_ULTt1x6m0_2;
	wire w_dff_B_AbNtEIjL5_2;
	wire w_dff_B_lvE1obt88_2;
	wire w_dff_B_iBUngahR0_2;
	wire w_dff_B_I9h71T3S9_2;
	wire w_dff_B_i8zJOOv59_2;
	wire w_dff_B_IV3hgyvv5_2;
	wire w_dff_B_8Vh7H1n24_2;
	wire w_dff_B_jIWbACyW1_2;
	wire w_dff_B_JDTFM5R30_2;
	wire w_dff_B_xrfzY9ts9_2;
	wire w_dff_B_rw8SYItt1_2;
	wire w_dff_B_EmR8Mzgg3_2;
	wire w_dff_B_jMujvKHS0_2;
	wire w_dff_B_pjdjxP1g7_2;
	wire w_dff_B_bYs6Ix2a4_2;
	wire w_dff_B_EKJJA52A3_2;
	wire w_dff_B_i14y3HXd4_2;
	wire w_dff_B_FnD7VnyZ3_2;
	wire w_dff_B_mBUFPWuq2_2;
	wire w_dff_B_3uOXTrKJ1_2;
	wire w_dff_B_T1uQ9chI8_1;
	wire w_dff_A_CXO8gbcQ6_1;
	wire w_dff_B_JxXpUVSx0_1;
	wire w_dff_B_uVZaACIL5_2;
	wire w_dff_B_bHSTeePt1_2;
	wire w_dff_B_htlcsEFH0_2;
	wire w_dff_B_lcj2qm6t2_2;
	wire w_dff_B_EtghrVxC9_2;
	wire w_dff_B_5liMHcCa9_2;
	wire w_dff_B_Y9BODGAs9_2;
	wire w_dff_B_B9fvqJFy0_2;
	wire w_dff_B_abzMz8sP6_2;
	wire w_dff_B_iOLw0N4M6_2;
	wire w_dff_B_VTnpXutI6_2;
	wire w_dff_B_6NU93XRJ6_2;
	wire w_dff_B_GdKwB8Lv4_2;
	wire w_dff_B_14jSVvej2_2;
	wire w_dff_B_zZ9gawPG5_2;
	wire w_dff_B_TBrCzMc67_2;
	wire w_dff_B_wAy2h7Xi6_2;
	wire w_dff_B_pjFifiQt1_2;
	wire w_dff_B_aQQlawh42_2;
	wire w_dff_B_7fZWpBWh8_2;
	wire w_dff_B_2RVGEWwl0_2;
	wire w_dff_B_Dw2SbVdT4_2;
	wire w_dff_B_ZmmyUifv6_2;
	wire w_dff_B_E6mFrMLs9_2;
	wire w_dff_B_9ONz9mZI6_2;
	wire w_dff_B_YpinjtRB9_2;
	wire w_dff_B_wfU26BUj4_2;
	wire w_dff_B_ccnFoE9b3_2;
	wire w_dff_B_iyeVOivS0_2;
	wire w_dff_B_ouB1yI5z7_2;
	wire w_dff_B_YozbgheA4_2;
	wire w_dff_B_teb3lBS75_2;
	wire w_dff_B_bBMX1SXG4_1;
	wire w_dff_B_3tYya2XY0_2;
	wire w_dff_B_v1RQoMpg7_2;
	wire w_dff_B_WQcnvxIS1_2;
	wire w_dff_B_rw1dArzp0_2;
	wire w_dff_B_0IfI2JDD8_2;
	wire w_dff_B_3E7Ld6Bs0_2;
	wire w_dff_B_X30TRNvY3_2;
	wire w_dff_B_aeo0v2Tf2_2;
	wire w_dff_B_IgGgScUL5_2;
	wire w_dff_B_g5uEQv1I1_2;
	wire w_dff_B_T6fOICOU1_2;
	wire w_dff_B_OFyTDMBY4_2;
	wire w_dff_B_tmKxvrc41_2;
	wire w_dff_B_bKKRr2714_2;
	wire w_dff_B_U5ervHxI2_2;
	wire w_dff_B_lOBdCHeu6_2;
	wire w_dff_B_gqgheVp73_2;
	wire w_dff_B_gtuRSp407_2;
	wire w_dff_B_hcyNNc3Z9_2;
	wire w_dff_B_8eh2Lelk7_2;
	wire w_dff_B_5ze0fl2n3_2;
	wire w_dff_B_48bVh6RE8_2;
	wire w_dff_B_ZRZU8uOx3_2;
	wire w_dff_B_YHapp4X36_2;
	wire w_dff_B_mLXa6sQJ9_2;
	wire w_dff_B_e85M0g4m3_2;
	wire w_dff_B_PQn5RWsp2_2;
	wire w_dff_B_NV8HOxjN1_2;
	wire w_dff_B_tZqSwIO23_1;
	wire w_dff_B_P4joCQYg5_2;
	wire w_dff_B_QmfJxSJy7_2;
	wire w_dff_B_LV407I1u0_2;
	wire w_dff_B_oJFCao3m1_2;
	wire w_dff_B_V368PBcs7_2;
	wire w_dff_B_row4fal99_2;
	wire w_dff_B_kZp2BKhT6_2;
	wire w_dff_B_Pl7SyZlU7_2;
	wire w_dff_B_Xt4tnPcO7_2;
	wire w_dff_B_lpmOVdQ54_2;
	wire w_dff_B_LsgDdFIg8_2;
	wire w_dff_B_qElhWWo46_2;
	wire w_dff_B_F0JHrGAW2_2;
	wire w_dff_B_Vu9BHf0p0_2;
	wire w_dff_B_0VP4dFnq5_2;
	wire w_dff_B_0umoayER2_2;
	wire w_dff_B_B6g4u4xj8_2;
	wire w_dff_B_x5D2HBSH9_2;
	wire w_dff_B_i4IWkU3F9_2;
	wire w_dff_B_XplDPMIh4_2;
	wire w_dff_B_iehERLSP1_2;
	wire w_dff_B_cg2rVmTo2_2;
	wire w_dff_B_q7tsYwk66_2;
	wire w_dff_B_pWZC72y62_2;
	wire w_dff_B_9dnTYMnJ8_2;
	wire w_dff_B_p41h6Qti7_2;
	wire w_dff_B_9QvM6iid7_1;
	wire w_dff_B_BkfCbZWX6_2;
	wire w_dff_B_kUUHDAXv5_2;
	wire w_dff_B_9EZKI3by1_2;
	wire w_dff_B_fiFWuJxT7_2;
	wire w_dff_B_zdWlGihM1_2;
	wire w_dff_B_p3773nxj0_2;
	wire w_dff_B_16hmqoeA9_2;
	wire w_dff_B_wwUoVEIr5_2;
	wire w_dff_B_ZOXR1ScA0_2;
	wire w_dff_B_7MfeQt6P9_2;
	wire w_dff_B_0Bgro4s80_2;
	wire w_dff_B_SDkt6Y1F9_2;
	wire w_dff_B_IWldop6H8_2;
	wire w_dff_B_C5LSL2EQ1_2;
	wire w_dff_B_sDq8JODP6_2;
	wire w_dff_B_XZh9nUX64_2;
	wire w_dff_B_SGlk6sFj3_2;
	wire w_dff_B_Pyo4Rq5w3_2;
	wire w_dff_B_gsKldul77_2;
	wire w_dff_B_CKCIkqQH0_2;
	wire w_dff_B_yhzC7Sh76_2;
	wire w_dff_B_YDp39mFV0_2;
	wire w_dff_B_4fkW6JxK3_2;
	wire w_dff_B_jgJwiJ2Q9_2;
	wire w_dff_B_PyIWdvaA6_1;
	wire w_dff_B_lbmaXOJY1_2;
	wire w_dff_B_mPa3lmCK3_2;
	wire w_dff_B_8Yr477c90_2;
	wire w_dff_B_sW1WAFPS0_2;
	wire w_dff_B_CqnvPrmL2_2;
	wire w_dff_B_D50kcWaK7_2;
	wire w_dff_B_zrgel2Dy4_2;
	wire w_dff_B_4vwQvhhj3_2;
	wire w_dff_B_YxucSGjf8_2;
	wire w_dff_B_qZMGiOAX5_2;
	wire w_dff_B_TBWixOTo6_2;
	wire w_dff_B_wDv85QkS5_2;
	wire w_dff_B_emq3D8w50_2;
	wire w_dff_B_syYZUY0t3_2;
	wire w_dff_B_jmb5iSCv1_2;
	wire w_dff_B_eBgt6N6R7_2;
	wire w_dff_B_iuYDfpUc6_2;
	wire w_dff_B_nEfFQ1Go9_2;
	wire w_dff_B_3Dsugy110_2;
	wire w_dff_B_hVQDOkSS3_2;
	wire w_dff_B_yxiWYFnD1_2;
	wire w_dff_B_vzjEJ0329_2;
	wire w_dff_B_MkDHctiK9_1;
	wire w_dff_B_n9jsUks89_2;
	wire w_dff_B_k7slm72j0_2;
	wire w_dff_B_9RyLp5TZ7_2;
	wire w_dff_B_M3tKHR808_2;
	wire w_dff_B_xMlmvkvB0_2;
	wire w_dff_B_Ue5FMrYX7_2;
	wire w_dff_B_HwXYzmyU7_2;
	wire w_dff_B_cqgbEvwX6_2;
	wire w_dff_B_xjRsQbBv0_2;
	wire w_dff_B_9ustTMDn8_2;
	wire w_dff_B_g6wcwBbm0_2;
	wire w_dff_B_MLbn53373_2;
	wire w_dff_B_EdpKmaZt9_2;
	wire w_dff_B_bR52msFv3_2;
	wire w_dff_B_JmZUqjjP3_2;
	wire w_dff_B_avDZQ1ym1_2;
	wire w_dff_B_vbwOjNoj6_2;
	wire w_dff_B_eXa8awt02_2;
	wire w_dff_B_iDvLRFo35_2;
	wire w_dff_B_M9eT0cLQ5_2;
	wire w_dff_B_N1mDFkm30_1;
	wire w_dff_B_SZFPGhcw5_2;
	wire w_dff_B_GLOgjmtE3_2;
	wire w_dff_B_mb2sjTnx7_2;
	wire w_dff_B_sBmDC3pi0_2;
	wire w_dff_B_5oJ2qCnK8_2;
	wire w_dff_B_f2vb1aiX9_2;
	wire w_dff_B_zzTTdMZO1_2;
	wire w_dff_B_xSClVX798_2;
	wire w_dff_B_VdZFHFro3_2;
	wire w_dff_B_7Ple399Z8_2;
	wire w_dff_B_M9iIYBxB7_2;
	wire w_dff_B_KFdhiOFG1_2;
	wire w_dff_B_c1vI4eX01_2;
	wire w_dff_B_kAfTQgna7_2;
	wire w_dff_B_fs7Orvfl1_2;
	wire w_dff_B_LGWKeNzZ6_2;
	wire w_dff_B_EX2uFdos1_2;
	wire w_dff_B_pHEqSSlV6_2;
	wire w_dff_B_ve9g9IJh7_1;
	wire w_dff_B_tdFI5j512_2;
	wire w_dff_B_ChzGEBgH6_2;
	wire w_dff_B_fFnX7s5g8_2;
	wire w_dff_B_rIV2zthO5_2;
	wire w_dff_B_HdPFFl2T7_2;
	wire w_dff_B_sspUpihD2_2;
	wire w_dff_B_BvoygqHS8_2;
	wire w_dff_B_xG4vfSU18_2;
	wire w_dff_B_VdNyaOtG2_2;
	wire w_dff_B_Y8SZASBv8_2;
	wire w_dff_B_inuMOoXO9_2;
	wire w_dff_B_5n7KzOh11_2;
	wire w_dff_B_Im5zIJB11_2;
	wire w_dff_B_QbO8q9Q09_2;
	wire w_dff_B_UM1nxNZv0_2;
	wire w_dff_B_ej1hnLyh5_2;
	wire w_dff_B_2a025RzN9_1;
	wire w_dff_B_zHOavq1r9_2;
	wire w_dff_B_7w0CKtHm8_2;
	wire w_dff_B_wZOorxwm3_2;
	wire w_dff_B_D3blI8sS7_2;
	wire w_dff_B_TdeFe2XB0_2;
	wire w_dff_B_hvpPu6Ru7_2;
	wire w_dff_B_UdRzhJVA8_2;
	wire w_dff_B_mF9M2XuR7_2;
	wire w_dff_B_dXdjQlLA2_2;
	wire w_dff_B_pSK8wpHS9_2;
	wire w_dff_B_i7HXVwUz8_2;
	wire w_dff_B_3wFakej16_2;
	wire w_dff_B_mRDtuQqn9_2;
	wire w_dff_B_jbGt7EVX8_2;
	wire w_dff_B_SqHIZXkK4_1;
	wire w_dff_B_3ejax37o8_2;
	wire w_dff_B_kQXBoYYd9_2;
	wire w_dff_B_DHpCnyVw3_2;
	wire w_dff_B_j1iZgJm40_2;
	wire w_dff_B_nrbmUWzl7_2;
	wire w_dff_B_jTnUMRra7_2;
	wire w_dff_B_cuQh6nq22_2;
	wire w_dff_B_RGnWy5n37_2;
	wire w_dff_B_d8n4TBcx5_2;
	wire w_dff_B_2oWBBBKG2_2;
	wire w_dff_B_AIUdJpQ50_2;
	wire w_dff_B_55nlJBQr7_2;
	wire w_dff_B_vx7Y6eO44_1;
	wire w_dff_B_6TFfjaJL1_2;
	wire w_dff_B_ArwKlyIB6_2;
	wire w_dff_B_ZFTwEkfj3_2;
	wire w_dff_B_MuwePaIo5_2;
	wire w_dff_B_I7DNNgbm7_2;
	wire w_dff_B_S7AZXOhM1_2;
	wire w_dff_B_sxVOcIA26_2;
	wire w_dff_B_VBDX5PDy4_2;
	wire w_dff_B_ng7WXPmM5_2;
	wire w_dff_B_axgwUMrn3_2;
	wire w_dff_B_i45uaWzw6_1;
	wire w_dff_B_wGhaQFtC5_2;
	wire w_dff_B_ZVhZyt6A6_2;
	wire w_dff_B_dUocCLtD0_2;
	wire w_dff_B_nEblCyuF6_2;
	wire w_dff_B_Tvwx1Hh83_2;
	wire w_dff_B_ydDJ2MsK4_2;
	wire w_dff_B_hkWByp8s3_2;
	wire w_dff_B_2l0AIDKB1_2;
	wire w_dff_B_d3jWtuDe0_2;
	wire w_dff_B_abVjiXtl9_2;
	wire w_dff_B_NqcXKRfB2_2;
	wire w_dff_B_dPym85Zo9_1;
	wire w_dff_B_9uF4WiNa0_1;
	wire w_dff_B_FriOFbtv9_1;
	wire w_dff_B_g1z8XKt61_2;
	wire w_dff_B_AmXH2p9Z4_2;
	wire w_dff_B_fhv5ubir5_2;
	wire w_dff_B_WnY7mpGK0_0;
	wire w_dff_B_YuU6LOnn8_0;
	wire w_dff_A_deehWp9L1_0;
	wire w_dff_A_i0usyGzS7_0;
	wire w_dff_A_3nZsfIXV0_1;
	wire w_dff_A_q2evcYDZ5_1;
	wire w_dff_B_vcEbTGsI3_2;
	wire w_dff_B_lFsWGR3P7_2;
	wire w_dff_B_4BsIzBMw6_1;
	wire w_dff_B_HxXebcxg5_2;
	wire w_dff_B_WP1rxRCJ5_2;
	wire w_dff_B_Yf1v076c4_2;
	wire w_dff_B_hUP16nCm6_2;
	wire w_dff_B_Vj41LMhi1_2;
	wire w_dff_B_dTTekMdM3_2;
	wire w_dff_B_yyrGMbKm5_2;
	wire w_dff_B_3qqGqiIU2_2;
	wire w_dff_B_Thp5r74E6_2;
	wire w_dff_B_Mby9w92n0_2;
	wire w_dff_B_MFuCVV3z0_2;
	wire w_dff_B_mGugFnAj8_2;
	wire w_dff_B_GVrmcoad6_2;
	wire w_dff_B_XZuJnthB2_2;
	wire w_dff_B_ThixVkvE8_2;
	wire w_dff_B_UNNmP23o0_2;
	wire w_dff_B_vaXIHUKE7_2;
	wire w_dff_B_Qo6fIxKZ0_2;
	wire w_dff_B_2L78vnbn8_2;
	wire w_dff_B_YtP7SnK81_2;
	wire w_dff_B_xNPo3ieC2_2;
	wire w_dff_B_Ui3D5MDp5_2;
	wire w_dff_B_4je9YzJo3_2;
	wire w_dff_B_efMuE7CX6_2;
	wire w_dff_B_ecrc3ieh1_2;
	wire w_dff_B_wpLvLIuC4_2;
	wire w_dff_B_pKdxKnsb3_2;
	wire w_dff_B_ihlCNmq73_2;
	wire w_dff_B_kqhi5uqQ2_2;
	wire w_dff_B_OIOSvCgg7_2;
	wire w_dff_B_ORssjp738_2;
	wire w_dff_B_roNJYT814_2;
	wire w_dff_B_2E8EtbSU8_2;
	wire w_dff_B_XLsmYfGI7_2;
	wire w_dff_B_9VQXBh5r1_2;
	wire w_dff_B_CAQSRdEd6_2;
	wire w_dff_B_9XTlHHFv3_2;
	wire w_dff_B_vDgUCxtX0_1;
	wire w_dff_A_v4JB5FpV2_1;
	wire w_dff_B_liHWSXZD3_1;
	wire w_dff_B_bIGjJxxb3_2;
	wire w_dff_B_rXwZGBD63_2;
	wire w_dff_B_WgiHGz0s8_2;
	wire w_dff_B_rQdvQecD2_2;
	wire w_dff_B_UPUZWbIe6_2;
	wire w_dff_B_U0GE3S6W1_2;
	wire w_dff_B_KPzSsgjv0_2;
	wire w_dff_B_2rlnimY87_2;
	wire w_dff_B_3e3Cxr9A0_2;
	wire w_dff_B_0yrACB2p8_2;
	wire w_dff_B_eRvYyFQ85_2;
	wire w_dff_B_DBcj978o6_2;
	wire w_dff_B_FM96viRs2_2;
	wire w_dff_B_oMKWUdUF9_2;
	wire w_dff_B_dZprClE56_2;
	wire w_dff_B_jz1lDOW31_2;
	wire w_dff_B_HzEPq7uv5_2;
	wire w_dff_B_0POMQpTl9_2;
	wire w_dff_B_ZgMhr7PX9_2;
	wire w_dff_B_4t2MH9Fy3_2;
	wire w_dff_B_5g1oNCoa5_2;
	wire w_dff_B_WYoIOJ5w0_2;
	wire w_dff_B_AUnmZvQP7_2;
	wire w_dff_B_BCUUKeE94_2;
	wire w_dff_B_NCWoOmXz5_2;
	wire w_dff_B_tcSpubjx4_2;
	wire w_dff_B_ahk9aaSS2_2;
	wire w_dff_B_Cfb46NbZ0_2;
	wire w_dff_B_3jrur08M2_2;
	wire w_dff_B_guWsENKn1_2;
	wire w_dff_B_svpNUMGJ3_2;
	wire w_dff_B_vNogexnc8_2;
	wire w_dff_B_dmovVPEO7_2;
	wire w_dff_B_vbv4jbug2_1;
	wire w_dff_B_knh65Mub3_2;
	wire w_dff_B_rtbfUa4N3_2;
	wire w_dff_B_yZfi7oZz8_2;
	wire w_dff_B_pHTBo1wK1_2;
	wire w_dff_B_FKJmDMMY6_2;
	wire w_dff_B_wO0lpCBD3_2;
	wire w_dff_B_ACzMNpoF2_2;
	wire w_dff_B_dXGolllw6_2;
	wire w_dff_B_4GtaH4zl4_2;
	wire w_dff_B_6KZDl10G0_2;
	wire w_dff_B_Zeq3fLLW5_2;
	wire w_dff_B_Vt5KTL0r0_2;
	wire w_dff_B_pUeBZUWe6_2;
	wire w_dff_B_jUJvx4VH5_2;
	wire w_dff_B_nhokQXfo1_2;
	wire w_dff_B_QCeetsf33_2;
	wire w_dff_B_zNTkDR803_2;
	wire w_dff_B_v8vEdzaX0_2;
	wire w_dff_B_nYgwjDA91_2;
	wire w_dff_B_P00oN6iR2_2;
	wire w_dff_B_9XN3JhzY1_2;
	wire w_dff_B_RCRf1bmH3_2;
	wire w_dff_B_ljr7OGIX8_2;
	wire w_dff_B_0eOHq9LC7_2;
	wire w_dff_B_XPhQYgMY8_2;
	wire w_dff_B_nrTVaabD0_2;
	wire w_dff_B_tc8xiSLQ0_2;
	wire w_dff_B_eJQXBWSO6_2;
	wire w_dff_B_zVqLTIM78_2;
	wire w_dff_B_ISmDjF5k2_2;
	wire w_dff_B_tnlqCwf56_1;
	wire w_dff_B_Qj94JnIk7_2;
	wire w_dff_B_9VoRz78x1_2;
	wire w_dff_B_gBKYXQ4D7_2;
	wire w_dff_B_kG10tY4k1_2;
	wire w_dff_B_30qgJ2EH2_2;
	wire w_dff_B_M4Z8Hivs2_2;
	wire w_dff_B_F4KsOBJO1_2;
	wire w_dff_B_QQnBUEyp3_2;
	wire w_dff_B_7ZfPdFRY5_2;
	wire w_dff_B_J8dcXqrp4_2;
	wire w_dff_B_R6o0VXny5_2;
	wire w_dff_B_tafc9iqI9_2;
	wire w_dff_B_IzPDP5jB8_2;
	wire w_dff_B_Pu03p8sT7_2;
	wire w_dff_B_Y16q20xC2_2;
	wire w_dff_B_38saKqEP7_2;
	wire w_dff_B_TPlCHBjx9_2;
	wire w_dff_B_lYFNPIfF0_2;
	wire w_dff_B_O6js9CB48_2;
	wire w_dff_B_Qp7ehhEF1_2;
	wire w_dff_B_KKss5IRV7_2;
	wire w_dff_B_Ah2DniCw0_2;
	wire w_dff_B_HnjCamSK3_2;
	wire w_dff_B_igQdNCZt8_2;
	wire w_dff_B_pTLzZ28K6_2;
	wire w_dff_B_8I3X7dEL7_2;
	wire w_dff_B_32Ixfw7Z1_1;
	wire w_dff_B_05gSVpdw3_2;
	wire w_dff_B_yIJGvAp85_2;
	wire w_dff_B_4sCuC4yF3_2;
	wire w_dff_B_ZkSQfUkp6_2;
	wire w_dff_B_WkxIbYJK8_2;
	wire w_dff_B_1anvwL6R7_2;
	wire w_dff_B_nKqflDpN1_2;
	wire w_dff_B_jai23uj43_2;
	wire w_dff_B_Y8NEOlcL3_2;
	wire w_dff_B_TWFxZrgN2_2;
	wire w_dff_B_KpoPiNBM4_2;
	wire w_dff_B_jPO5Zibc1_2;
	wire w_dff_B_H3RETrgb0_2;
	wire w_dff_B_nBP5DtAl5_2;
	wire w_dff_B_AdWUsOxP8_2;
	wire w_dff_B_ufbezDiC3_2;
	wire w_dff_B_1hqYdLjg5_2;
	wire w_dff_B_QS1HdsCf1_2;
	wire w_dff_B_6qWUsFaA0_2;
	wire w_dff_B_kGukgcjl9_2;
	wire w_dff_B_mxkdFD5P6_2;
	wire w_dff_B_6n67HBBO9_2;
	wire w_dff_B_3CjuWQ8Z6_2;
	wire w_dff_B_NAXPIAqq6_2;
	wire w_dff_B_Q4Onb2760_1;
	wire w_dff_B_J1TpgkZa1_2;
	wire w_dff_B_t54vy7cw7_2;
	wire w_dff_B_DLSclZDo4_2;
	wire w_dff_B_7I7Xx8TQ5_2;
	wire w_dff_B_U4z9WrT53_2;
	wire w_dff_B_cPaktSpE2_2;
	wire w_dff_B_ckRVo5Xu4_2;
	wire w_dff_B_GBGJH0nS2_2;
	wire w_dff_B_RnMAILM42_2;
	wire w_dff_B_cUtcAg0O3_2;
	wire w_dff_B_D5LXQRvh7_2;
	wire w_dff_B_U0q6GnRr9_2;
	wire w_dff_B_gtCuGuHR7_2;
	wire w_dff_B_tcemRyZ50_2;
	wire w_dff_B_Xxend09L6_2;
	wire w_dff_B_ths3gjrN0_2;
	wire w_dff_B_5C92nWMz1_2;
	wire w_dff_B_Vk1ekSo52_2;
	wire w_dff_B_UHr93JyK7_2;
	wire w_dff_B_5vi4CxmF0_2;
	wire w_dff_B_5QJ5XjO55_2;
	wire w_dff_B_tZNJFONl2_2;
	wire w_dff_B_byEMZ9rd5_1;
	wire w_dff_B_5FYseBB29_2;
	wire w_dff_B_LiV73i203_2;
	wire w_dff_B_1XOHmA2o5_2;
	wire w_dff_B_DNfBUdyz0_2;
	wire w_dff_B_4i3vdge22_2;
	wire w_dff_B_JNGCyc2R0_2;
	wire w_dff_B_psIUSbKE4_2;
	wire w_dff_B_LJJNhOXG3_2;
	wire w_dff_B_RPOP7lpy4_2;
	wire w_dff_B_Dw1Yxqoj4_2;
	wire w_dff_B_BEa72CjN0_2;
	wire w_dff_B_VIr7JqWL2_2;
	wire w_dff_B_6L9BxnXQ0_2;
	wire w_dff_B_VJd2gfhQ2_2;
	wire w_dff_B_e6b5PeZB6_2;
	wire w_dff_B_Mi3PdvAa4_2;
	wire w_dff_B_VLVyVtTV6_2;
	wire w_dff_B_s82yRrnj0_2;
	wire w_dff_B_4Q9KcXTf9_2;
	wire w_dff_B_H8LlxpHs5_2;
	wire w_dff_B_XRr1dIOp7_1;
	wire w_dff_B_3o5rqsgq2_2;
	wire w_dff_B_4YMOUERR2_2;
	wire w_dff_B_U5JA5O9V8_2;
	wire w_dff_B_Rzrb5ZfJ1_2;
	wire w_dff_B_Ny8n0kyf1_2;
	wire w_dff_B_zF8eUwa44_2;
	wire w_dff_B_MoXylkxK3_2;
	wire w_dff_B_wSanp7K27_2;
	wire w_dff_B_0C9iyqU23_2;
	wire w_dff_B_08PxsBWl0_2;
	wire w_dff_B_QD6AugsZ3_2;
	wire w_dff_B_a3LTYmG01_2;
	wire w_dff_B_aHkiFuol9_2;
	wire w_dff_B_vVJLfvtI6_2;
	wire w_dff_B_TJjKZfoF1_2;
	wire w_dff_B_wl9s6AQB5_2;
	wire w_dff_B_ORs8uBqX0_2;
	wire w_dff_B_HZ2Qo92N7_2;
	wire w_dff_B_qeTXLU0b4_1;
	wire w_dff_B_MV4g2QNt1_2;
	wire w_dff_B_0eHZLoD04_2;
	wire w_dff_B_W7AdgweC5_2;
	wire w_dff_B_LS6ZICUD4_2;
	wire w_dff_B_PkFdBYLG5_2;
	wire w_dff_B_Fb2tyx6g7_2;
	wire w_dff_B_rJT8Zncn9_2;
	wire w_dff_B_j2p7VuyT1_2;
	wire w_dff_B_DC6MZPiF0_2;
	wire w_dff_B_gDN95RFl9_2;
	wire w_dff_B_M7hA9fv73_2;
	wire w_dff_B_DbPxRwwp4_2;
	wire w_dff_B_aAxi0Nzn0_2;
	wire w_dff_B_hBOGrQ0T1_2;
	wire w_dff_B_NHJGJXl27_2;
	wire w_dff_B_G3u1fkFI6_2;
	wire w_dff_B_pv43riop8_1;
	wire w_dff_B_wzwUUzUm6_2;
	wire w_dff_B_sGWruZf97_2;
	wire w_dff_B_H4z0HhCZ5_2;
	wire w_dff_B_ZJToBRjJ9_2;
	wire w_dff_B_VOnpvlJC5_2;
	wire w_dff_B_Z27iRV4o5_2;
	wire w_dff_B_ILFoDVZr5_2;
	wire w_dff_B_RHfHr3450_2;
	wire w_dff_B_ONCMmMQe1_2;
	wire w_dff_B_SM3xvBQ74_2;
	wire w_dff_B_sGBLMMv97_2;
	wire w_dff_B_85GcJfkc8_2;
	wire w_dff_B_EQkdYyZx9_2;
	wire w_dff_B_8lzSH3qA1_2;
	wire w_dff_B_yHDS6tVh6_1;
	wire w_dff_B_46lKdd870_2;
	wire w_dff_B_lbO1yTzX7_2;
	wire w_dff_B_E2FFnZge7_2;
	wire w_dff_B_FVVSrVpF4_2;
	wire w_dff_B_ni1JN2Xc0_2;
	wire w_dff_B_secEvfco7_2;
	wire w_dff_B_QSOhLVTd7_2;
	wire w_dff_B_dD4Wqlsh4_2;
	wire w_dff_B_PraNFw2U9_2;
	wire w_dff_B_Rb50kEvB0_2;
	wire w_dff_B_JXa4nZxj1_2;
	wire w_dff_B_nJrMpPDH9_2;
	wire w_dff_B_pqEVTRr14_1;
	wire w_dff_B_vZ7Tk3AX0_2;
	wire w_dff_B_FvkMsqtZ1_2;
	wire w_dff_B_a74mIRXI9_2;
	wire w_dff_B_xAWvAewH2_2;
	wire w_dff_B_ZjSdn17E9_2;
	wire w_dff_B_aLhjPEKB1_2;
	wire w_dff_B_DdgUgEna3_2;
	wire w_dff_B_tEaF8pVO8_2;
	wire w_dff_B_NBUfx7Fj6_2;
	wire w_dff_B_v8dDabgb2_2;
	wire w_dff_B_hJD0JWYq0_1;
	wire w_dff_B_VFwt9rHg2_2;
	wire w_dff_B_T9pbeyQO9_2;
	wire w_dff_B_6OL5UTYf6_2;
	wire w_dff_B_TPERxyw56_2;
	wire w_dff_B_A8gqdoZC5_2;
	wire w_dff_B_x5HBSNPC4_2;
	wire w_dff_B_Q4cWheUz4_2;
	wire w_dff_B_R9xRJ5ll5_2;
	wire w_dff_B_tMloJh7K6_2;
	wire w_dff_B_CFjS2mkS2_2;
	wire w_dff_B_UcTBY1zo6_2;
	wire w_dff_B_0Nzhwj1O0_1;
	wire w_dff_B_H81iEytJ1_1;
	wire w_dff_B_nZmWx5Sh4_1;
	wire w_dff_B_qE3ues0G9_2;
	wire w_dff_B_66EUHV0c6_2;
	wire w_dff_B_tL739E4x0_2;
	wire w_dff_B_UeAzmlqM4_0;
	wire w_dff_B_xsOacfNt7_0;
	wire w_dff_A_8d0lntMq6_0;
	wire w_dff_A_BwRsfu1h5_0;
	wire w_dff_A_Dof8RIBx2_1;
	wire w_dff_A_JeJnM9zr2_1;
	wire w_dff_B_xnQZKn1e6_2;
	wire w_dff_B_mkSi4f4V7_1;
	wire w_dff_B_VBW0ogTI6_2;
	wire w_dff_B_v1rfo64M4_2;
	wire w_dff_B_5uEtOVsX1_2;
	wire w_dff_B_vA7Gn5HE4_2;
	wire w_dff_B_cKb7ezjL7_2;
	wire w_dff_B_FyPHq40p4_2;
	wire w_dff_B_S3wNH8I13_2;
	wire w_dff_B_bYp6fC688_2;
	wire w_dff_B_XjrGQonB5_2;
	wire w_dff_B_PUetbgfh8_2;
	wire w_dff_B_IR4AG0en0_2;
	wire w_dff_B_iYvU3GlE3_2;
	wire w_dff_B_I1MDHbGc8_2;
	wire w_dff_B_l3Uq8J3R3_2;
	wire w_dff_B_fuC5iLKZ6_2;
	wire w_dff_B_dSrZ6e8f8_2;
	wire w_dff_B_giSfxoBs5_2;
	wire w_dff_B_YcJC36jV9_2;
	wire w_dff_B_UkU0bqgI9_2;
	wire w_dff_B_pbWx9hp86_2;
	wire w_dff_B_f535UBey5_2;
	wire w_dff_B_drC7sw329_2;
	wire w_dff_B_biQrQ1sy3_2;
	wire w_dff_B_PvuNGnTA0_2;
	wire w_dff_B_qEhnOnfS6_2;
	wire w_dff_B_UVALDTH68_2;
	wire w_dff_B_wb9MDVlw4_2;
	wire w_dff_B_kxeHh8gX1_2;
	wire w_dff_B_yQSN8lAV2_2;
	wire w_dff_B_59J1qeTa2_2;
	wire w_dff_B_Ni8wF5Du1_2;
	wire w_dff_B_V2TkmjJu0_2;
	wire w_dff_B_5cGNZfKr3_2;
	wire w_dff_B_ISv9F1e59_2;
	wire w_dff_B_RbBpgmtv8_2;
	wire w_dff_B_2jGGkJn77_2;
	wire w_dff_B_wqI2kAQe6_2;
	wire w_dff_B_TtcXziLy1_2;
	wire w_dff_B_e2z1JxOl1_1;
	wire w_dff_A_6pYNKldV8_1;
	wire w_dff_B_TSNOL1hx3_1;
	wire w_dff_B_mrDJFLs04_2;
	wire w_dff_B_W8cHUeGZ6_2;
	wire w_dff_B_1PnuUv3N0_2;
	wire w_dff_B_C9r2fK6t9_2;
	wire w_dff_B_zk2KIBey5_2;
	wire w_dff_B_I1Wo4Yuv6_2;
	wire w_dff_B_HPViOFY71_2;
	wire w_dff_B_Cv0Y47s56_2;
	wire w_dff_B_9RQSnSrE4_2;
	wire w_dff_B_QDUvAwlg1_2;
	wire w_dff_B_uy26qrPp3_2;
	wire w_dff_B_2FAmawaL9_2;
	wire w_dff_B_bblRoeif6_2;
	wire w_dff_B_NmDeHrv92_2;
	wire w_dff_B_iag5fKQv0_2;
	wire w_dff_B_UqmFmJSE5_2;
	wire w_dff_B_NUfuTtUN9_2;
	wire w_dff_B_KPj8zJaL3_2;
	wire w_dff_B_54Lssekp8_2;
	wire w_dff_B_MPCYk8OS1_2;
	wire w_dff_B_v9Qg1kqt6_2;
	wire w_dff_B_KPqy328H8_2;
	wire w_dff_B_h5sjxDfW7_2;
	wire w_dff_B_3B3PTyVI2_2;
	wire w_dff_B_1W9eD1rp9_2;
	wire w_dff_B_G9apCEHq0_2;
	wire w_dff_B_DebhzyCI5_2;
	wire w_dff_B_EeJqWmaU2_2;
	wire w_dff_B_mXaempWy3_2;
	wire w_dff_B_YOdfcH9A2_2;
	wire w_dff_B_KmXp3FyI1_2;
	wire w_dff_B_fkTswcPr6_2;
	wire w_dff_B_x51BuWjL3_2;
	wire w_dff_B_O0h7KmFr2_2;
	wire w_dff_B_u31k2Nk20_1;
	wire w_dff_B_H2OXBbe60_2;
	wire w_dff_B_bGnWXqi60_2;
	wire w_dff_B_P8ofvFfx7_2;
	wire w_dff_B_e1svo0Zp3_2;
	wire w_dff_B_jcTSoOaC6_2;
	wire w_dff_B_VCwa01U53_2;
	wire w_dff_B_3cFxOmPa2_2;
	wire w_dff_B_QKCVJ6FN0_2;
	wire w_dff_B_pmQdjvRI5_2;
	wire w_dff_B_zf69GMFj3_2;
	wire w_dff_B_KsRGGLFJ3_2;
	wire w_dff_B_moAuZaV85_2;
	wire w_dff_B_wFmrwfXv7_2;
	wire w_dff_B_TEwjkeF74_2;
	wire w_dff_B_7WNqZ5P39_2;
	wire w_dff_B_YP0FbpPG0_2;
	wire w_dff_B_YY09gFww6_2;
	wire w_dff_B_lwF4kr7x7_2;
	wire w_dff_B_jBAMjf907_2;
	wire w_dff_B_yq7oWzje7_2;
	wire w_dff_B_mRCykEN71_2;
	wire w_dff_B_0WDdaiKY2_2;
	wire w_dff_B_QT5TQdAh1_2;
	wire w_dff_B_3TdHUadp2_2;
	wire w_dff_B_d4Jc6hM94_2;
	wire w_dff_B_mi6L5EPP3_2;
	wire w_dff_B_Jle96uyH5_2;
	wire w_dff_B_b5EcWls47_2;
	wire w_dff_B_37bKEhBh2_2;
	wire w_dff_B_MDqnxK5G5_2;
	wire w_dff_B_zyA9jFjr4_2;
	wire w_dff_B_2vYE8m0s1_1;
	wire w_dff_B_Lp7qrQX68_2;
	wire w_dff_B_GOI2Y9Hg3_2;
	wire w_dff_B_cXlxZi112_2;
	wire w_dff_B_PLcetyJE8_2;
	wire w_dff_B_jZYNkq4D0_2;
	wire w_dff_B_tWsxuWkU3_2;
	wire w_dff_B_LSXcQq172_2;
	wire w_dff_B_PEIXlRVK9_2;
	wire w_dff_B_6wzu7IFF4_2;
	wire w_dff_B_ZmVlozeC0_2;
	wire w_dff_B_abLewnl91_2;
	wire w_dff_B_8Tzx9gzi2_2;
	wire w_dff_B_xEo1Kzkw9_2;
	wire w_dff_B_oyhSLhkL7_2;
	wire w_dff_B_V7ksLEFL8_2;
	wire w_dff_B_uhbOoM2d0_2;
	wire w_dff_B_UyWvtaUl7_2;
	wire w_dff_B_kbO544K39_2;
	wire w_dff_B_1cA5keYn5_2;
	wire w_dff_B_EfpL2XTI4_2;
	wire w_dff_B_sWd6KsID9_2;
	wire w_dff_B_QLWdYeyX0_2;
	wire w_dff_B_ybNKA7OT0_2;
	wire w_dff_B_h025lGvm0_2;
	wire w_dff_B_I81kX4pU9_2;
	wire w_dff_B_a0zie5520_2;
	wire w_dff_B_epbHyQ9n1_2;
	wire w_dff_B_LfDwkVxA7_2;
	wire w_dff_B_iLDdWkPX6_1;
	wire w_dff_B_LHZ4VKIQ4_2;
	wire w_dff_B_KezderHx2_2;
	wire w_dff_B_zZOMMQSe4_2;
	wire w_dff_B_8j2kBVfM4_2;
	wire w_dff_B_dCYtdT4w2_2;
	wire w_dff_B_EVyvL9BR6_2;
	wire w_dff_B_B6KoHIF87_2;
	wire w_dff_B_ZMqyKINg0_2;
	wire w_dff_B_CkXqgppJ3_2;
	wire w_dff_B_CyJj60EX0_2;
	wire w_dff_B_SeFTTevc0_2;
	wire w_dff_B_9IZW18Hb4_2;
	wire w_dff_B_7vaySFdw6_2;
	wire w_dff_B_jYSe9qsF4_2;
	wire w_dff_B_gyu3aPvi6_2;
	wire w_dff_B_GOicqNIt5_2;
	wire w_dff_B_awE6hmV85_2;
	wire w_dff_B_jslbRFA42_2;
	wire w_dff_B_Q4O5XPDp2_2;
	wire w_dff_B_ZAZKT3xQ9_2;
	wire w_dff_B_gxTUHhmZ6_2;
	wire w_dff_B_pCx6GYyo0_2;
	wire w_dff_B_qrtJTwc08_2;
	wire w_dff_B_RmbCiMPF6_2;
	wire w_dff_B_u4aSQSdF1_1;
	wire w_dff_B_Cx6My3pg9_2;
	wire w_dff_B_QXcIqmq80_2;
	wire w_dff_B_kkAoFUco2_2;
	wire w_dff_B_P73OyyiO4_2;
	wire w_dff_B_CZLw1cXT6_2;
	wire w_dff_B_HwFPJ4EA4_2;
	wire w_dff_B_NrFrBWx25_2;
	wire w_dff_B_mywMtiu13_2;
	wire w_dff_B_bB7dcx8R3_2;
	wire w_dff_B_uQPBbs0O3_2;
	wire w_dff_B_xN7pEiYJ9_2;
	wire w_dff_B_fM7Yq2WQ8_2;
	wire w_dff_B_aLxOuJhY3_2;
	wire w_dff_B_3Q4pkfNi1_2;
	wire w_dff_B_yYhd4daa7_2;
	wire w_dff_B_ZlA9nWD81_2;
	wire w_dff_B_QQcGgiGy7_2;
	wire w_dff_B_Lyn5RP2y2_2;
	wire w_dff_B_t0tqAlfT0_2;
	wire w_dff_B_SOP43ZMk1_2;
	wire w_dff_B_vRSC99dJ8_2;
	wire w_dff_B_pzaxuUlC1_2;
	wire w_dff_B_7NXe1aam5_1;
	wire w_dff_B_Je0dIbIX7_2;
	wire w_dff_B_szC91N574_2;
	wire w_dff_B_LXmzBUpG3_2;
	wire w_dff_B_Ey5AIvti9_2;
	wire w_dff_B_kyz0yeSz2_2;
	wire w_dff_B_JgHuZNH30_2;
	wire w_dff_B_kLGMyrwD4_2;
	wire w_dff_B_5M5P6f7G8_2;
	wire w_dff_B_NRndCDC24_2;
	wire w_dff_B_xEyC5FTv0_2;
	wire w_dff_B_SmXU5iOp1_2;
	wire w_dff_B_39Wr9A6V8_2;
	wire w_dff_B_u9R9wBej9_2;
	wire w_dff_B_WpCQmerQ5_2;
	wire w_dff_B_9czaz7Yk1_2;
	wire w_dff_B_W8Jkh4iC0_2;
	wire w_dff_B_i2HOhHua3_2;
	wire w_dff_B_rYLJkBLd3_2;
	wire w_dff_B_eZElVmW97_2;
	wire w_dff_B_Sr08VwJO8_2;
	wire w_dff_B_qXyM7Qwc6_1;
	wire w_dff_B_0TvzjfHU0_2;
	wire w_dff_B_ypmmE3C39_2;
	wire w_dff_B_K1R5TRh27_2;
	wire w_dff_B_3n3PnFyB1_2;
	wire w_dff_B_Sig101506_2;
	wire w_dff_B_bolEqkLW1_2;
	wire w_dff_B_fLhQkqRH7_2;
	wire w_dff_B_LHj4UaqR2_2;
	wire w_dff_B_iDje99eB5_2;
	wire w_dff_B_MskXIIxs6_2;
	wire w_dff_B_Od0FDlA80_2;
	wire w_dff_B_SkRX7Q4g9_2;
	wire w_dff_B_Z3rNbKFV1_2;
	wire w_dff_B_EBMd0cWs6_2;
	wire w_dff_B_WOqC9OdB8_2;
	wire w_dff_B_6vGPQelS1_2;
	wire w_dff_B_KWjXixrE8_2;
	wire w_dff_B_SU75RpGS3_2;
	wire w_dff_B_VVYYVHft7_1;
	wire w_dff_B_BfT0IfDy2_2;
	wire w_dff_B_OXIeXVOr8_2;
	wire w_dff_B_BSdDzozM3_2;
	wire w_dff_B_iNE26wtK5_2;
	wire w_dff_B_UNbIj7qn2_2;
	wire w_dff_B_R1mUILyP9_2;
	wire w_dff_B_i22bJWZf3_2;
	wire w_dff_B_XOmWZpx17_2;
	wire w_dff_B_Clb3lzXg2_2;
	wire w_dff_B_Y5DmB6y44_2;
	wire w_dff_B_l1NKi4vi9_2;
	wire w_dff_B_4wDrXFRU9_2;
	wire w_dff_B_KuIwdfcf8_2;
	wire w_dff_B_s7sd3LNW0_2;
	wire w_dff_B_qcPQIcQb7_2;
	wire w_dff_B_7EOlVDn41_2;
	wire w_dff_B_QeeoHfcw0_1;
	wire w_dff_B_r1S7Xluw5_2;
	wire w_dff_B_6zsibY9X8_2;
	wire w_dff_B_emK3KRQX6_2;
	wire w_dff_B_TIZwAch08_2;
	wire w_dff_B_B73Ro9kn2_2;
	wire w_dff_B_LlOJyFvd9_2;
	wire w_dff_B_rTAbZuoW4_2;
	wire w_dff_B_Tt00uwKb7_2;
	wire w_dff_B_0GwSHv5V9_2;
	wire w_dff_B_lm4pPCWv7_2;
	wire w_dff_B_fQTOUhIF3_2;
	wire w_dff_B_wIS1m3YM7_2;
	wire w_dff_B_S7K19t8L1_2;
	wire w_dff_B_44BG7z7r0_2;
	wire w_dff_B_KBFvPjWb1_1;
	wire w_dff_B_D2sIU5y97_2;
	wire w_dff_B_EVx0lc9W5_2;
	wire w_dff_B_2nkXRlqF9_2;
	wire w_dff_B_bAttG5yd2_2;
	wire w_dff_B_76T5mV5z6_2;
	wire w_dff_B_Z2P859FC9_2;
	wire w_dff_B_3bHjqqJB5_2;
	wire w_dff_B_j9H94ud07_2;
	wire w_dff_B_0xnVnBxE4_2;
	wire w_dff_B_H5M5tGWS7_2;
	wire w_dff_B_IAEuopXa7_2;
	wire w_dff_B_sglmE4pR1_2;
	wire w_dff_B_rotSg5d82_1;
	wire w_dff_B_XxAVYfDU5_2;
	wire w_dff_B_S2EemTn48_2;
	wire w_dff_B_cygVIqK89_2;
	wire w_dff_B_sFRzDL4a8_2;
	wire w_dff_B_jV1cZg2Q9_2;
	wire w_dff_B_VNar4xOi1_2;
	wire w_dff_B_z6V0r9oE0_2;
	wire w_dff_B_O7dbEXDU5_2;
	wire w_dff_B_oVoN5YBR6_2;
	wire w_dff_B_z6gQ9hNy3_2;
	wire w_dff_B_WREzFNmg8_1;
	wire w_dff_B_K1M8SoWB3_2;
	wire w_dff_B_wx5N0beU2_2;
	wire w_dff_B_Z8JK565X9_2;
	wire w_dff_B_nZiFLd5J9_2;
	wire w_dff_B_P4GtX4Xi9_2;
	wire w_dff_B_Z1Kc7rXZ8_2;
	wire w_dff_B_RmGjfVPt2_2;
	wire w_dff_B_1NLc7XxL1_2;
	wire w_dff_B_i8R0CmxG1_2;
	wire w_dff_B_7Rufg3Uj7_2;
	wire w_dff_B_N5Yqmrr39_2;
	wire w_dff_B_NUrjUkee4_1;
	wire w_dff_B_l32r1WdK3_1;
	wire w_dff_B_VFNjns4h3_1;
	wire w_dff_B_SdMVL1by0_2;
	wire w_dff_B_dM63tieg8_2;
	wire w_dff_B_tds3ch0X2_2;
	wire w_dff_B_RsaZpdi96_0;
	wire w_dff_B_fr6mKTAI4_0;
	wire w_dff_A_3Gg0Z0b75_0;
	wire w_dff_A_MVF4fcjn7_0;
	wire w_dff_A_VINnGMiS2_1;
	wire w_dff_A_BMAwMXjb2_1;
	wire w_dff_B_PE4m5ZCu8_1;
	wire w_dff_A_csoi6cFm2_1;
	wire w_dff_B_32RUcBr69_1;
	wire w_dff_B_QFG62Yqq9_2;
	wire w_dff_B_Ilcs4dY33_2;
	wire w_dff_B_QxHhpsNM5_2;
	wire w_dff_B_v44tIc602_2;
	wire w_dff_B_Flk4j5qc4_2;
	wire w_dff_B_kXpcI2eY9_2;
	wire w_dff_B_4BQSOL2l2_2;
	wire w_dff_B_aTFLY3PB2_2;
	wire w_dff_B_VLvrWuPZ5_2;
	wire w_dff_B_61sxVVWt4_2;
	wire w_dff_B_5QzWkgxD5_2;
	wire w_dff_B_qHmSAEz46_2;
	wire w_dff_B_s9zqOVEC5_2;
	wire w_dff_B_XO13hPQY3_2;
	wire w_dff_B_cSGCRgcZ1_2;
	wire w_dff_B_7pBR1iIP9_2;
	wire w_dff_B_e7xPARvF0_2;
	wire w_dff_B_WRyTq3sK4_2;
	wire w_dff_B_KE67mPxR4_2;
	wire w_dff_B_PLxFEBDJ1_2;
	wire w_dff_B_k4wOFEZD3_2;
	wire w_dff_B_mklHn2su3_2;
	wire w_dff_B_ip3aEDJF2_2;
	wire w_dff_B_rPDyahFY4_2;
	wire w_dff_B_Mf5Wy88i1_2;
	wire w_dff_B_joXVuqhp2_2;
	wire w_dff_B_FECT2AFU8_2;
	wire w_dff_B_vRZxbveO2_2;
	wire w_dff_B_EYgmD8Ne1_2;
	wire w_dff_B_Ezudp3L23_2;
	wire w_dff_B_BwBQcOWF6_2;
	wire w_dff_B_5ZcHfyEw7_2;
	wire w_dff_B_kHEsQ9Ld2_2;
	wire w_dff_B_mdSCRtuO2_2;
	wire w_dff_B_j3rHZW2q5_2;
	wire w_dff_B_62HyjOUL2_2;
	wire w_dff_B_9b7f8n6n3_2;
	wire w_dff_B_ezdYGMnN4_2;
	wire w_dff_B_QOTySqd87_1;
	wire w_dff_B_snGtzBvx5_2;
	wire w_dff_B_NBysoQ4p3_2;
	wire w_dff_B_gDaZSkVr3_2;
	wire w_dff_B_TEbkZlle4_2;
	wire w_dff_B_bHn8kcXD5_2;
	wire w_dff_B_LBRinYkX5_2;
	wire w_dff_B_4prf02q09_2;
	wire w_dff_B_M3dqth1M4_2;
	wire w_dff_B_gRGnvf8h5_2;
	wire w_dff_B_rpwoirJ62_2;
	wire w_dff_B_I7PBHofI5_2;
	wire w_dff_B_oViZ8m8C6_2;
	wire w_dff_B_55RINX5E8_2;
	wire w_dff_B_mvEzyRlR7_2;
	wire w_dff_B_zefmrKuf7_2;
	wire w_dff_B_3QkWOUJC9_2;
	wire w_dff_B_x8JYUs909_2;
	wire w_dff_B_eAFvx1Xe2_2;
	wire w_dff_B_pxEy49Oz7_2;
	wire w_dff_B_uqD9fGBQ8_2;
	wire w_dff_B_Y5uPpjE31_2;
	wire w_dff_B_1mgMYVK02_2;
	wire w_dff_B_S2zN05ch2_2;
	wire w_dff_B_1RI0rbVI0_2;
	wire w_dff_B_FWbA67yj3_2;
	wire w_dff_B_xHyk3nty9_2;
	wire w_dff_B_SFSMzVUo6_2;
	wire w_dff_B_HDWKiVzy6_2;
	wire w_dff_B_jlh42iic2_2;
	wire w_dff_B_mIy2pGjT3_2;
	wire w_dff_B_0ztbaOph2_2;
	wire w_dff_B_0FNj0ARD4_2;
	wire w_dff_B_2iv5EmEG0_2;
	wire w_dff_B_wbcx4oOg9_2;
	wire w_dff_B_Jm07S3Nn1_2;
	wire w_dff_B_m01alN119_1;
	wire w_dff_B_ermCbF732_2;
	wire w_dff_B_ZBX9aFZ51_2;
	wire w_dff_B_YFzwZPHy3_2;
	wire w_dff_B_mImqg4pu8_2;
	wire w_dff_B_FO0qQGWH9_2;
	wire w_dff_B_2EoKPnfP0_2;
	wire w_dff_B_eecEN4h19_2;
	wire w_dff_B_8ZCZzsU97_2;
	wire w_dff_B_gZpl0MII6_2;
	wire w_dff_B_5h4jZKRI8_2;
	wire w_dff_B_xXzivMBD0_2;
	wire w_dff_B_mPOjsurX1_2;
	wire w_dff_B_XcVyYVsk9_2;
	wire w_dff_B_BqVaqLSy3_2;
	wire w_dff_B_lz6MFlZF6_2;
	wire w_dff_B_cmQc13Iz5_2;
	wire w_dff_B_YrCD7PYW2_2;
	wire w_dff_B_vCbtqf1q7_2;
	wire w_dff_B_pp9o9R0J7_2;
	wire w_dff_B_Rk3wQcSV7_2;
	wire w_dff_B_uphxZ8yQ8_2;
	wire w_dff_B_LQgzsqpU9_2;
	wire w_dff_B_jBGzCqon4_2;
	wire w_dff_B_vVDunm8L6_2;
	wire w_dff_B_NTVXSH8x3_2;
	wire w_dff_B_0KlK6uy33_2;
	wire w_dff_B_gRXbMaD91_2;
	wire w_dff_B_Y2I6Z5fF7_2;
	wire w_dff_B_NkJEGTb19_2;
	wire w_dff_B_GbV6ToqS5_2;
	wire w_dff_B_bx6MHFYJ5_2;
	wire w_dff_B_5R5a4ZnB0_2;
	wire w_dff_B_3kuIQJaL6_1;
	wire w_dff_B_Nx6prODT8_2;
	wire w_dff_B_MmvvBlnb3_2;
	wire w_dff_B_L1ubTD0n1_2;
	wire w_dff_B_vxl184fQ4_2;
	wire w_dff_B_DXTahOtP4_2;
	wire w_dff_B_F5VknJy19_2;
	wire w_dff_B_g2fWq3F15_2;
	wire w_dff_B_mFRTmooO7_2;
	wire w_dff_B_Latnbfx71_2;
	wire w_dff_B_Erg1BIIt3_2;
	wire w_dff_B_uu3iam9e8_2;
	wire w_dff_B_owth1e5B6_2;
	wire w_dff_B_GaxctY0k4_2;
	wire w_dff_B_HEKkRr1X2_2;
	wire w_dff_B_AmlPPiku1_2;
	wire w_dff_B_natso62S0_2;
	wire w_dff_B_pK1nzeUa4_2;
	wire w_dff_B_cmARzKOa5_2;
	wire w_dff_B_ocWjzMWV2_2;
	wire w_dff_B_aD68uE3Q9_2;
	wire w_dff_B_n4EjIrH36_2;
	wire w_dff_B_8fwdlhds5_2;
	wire w_dff_B_olnEJeUQ0_2;
	wire w_dff_B_1Aunm1g73_2;
	wire w_dff_B_8zQr2RJb9_2;
	wire w_dff_B_AABk88Ph4_2;
	wire w_dff_B_0G3pVopU8_2;
	wire w_dff_B_meCKv3YC1_2;
	wire w_dff_B_yYSeLr7z7_2;
	wire w_dff_B_RIrmifht4_1;
	wire w_dff_B_7kgFtJlb4_2;
	wire w_dff_B_5PzBCSYi1_2;
	wire w_dff_B_O4CBBEIG3_2;
	wire w_dff_B_7Et7zRrX0_2;
	wire w_dff_B_N8nFr6Ah9_2;
	wire w_dff_B_qS3xw9qH4_2;
	wire w_dff_B_F0P9hycQ6_2;
	wire w_dff_B_EckjCATr2_2;
	wire w_dff_B_hfhgTPjF1_2;
	wire w_dff_B_dk3gJiMF1_2;
	wire w_dff_B_VQJ4USoi2_2;
	wire w_dff_B_sbq09ePv9_2;
	wire w_dff_B_8ET0SBc69_2;
	wire w_dff_B_8MgNKCBv6_2;
	wire w_dff_B_K0KcBQaj9_2;
	wire w_dff_B_A8WpoR518_2;
	wire w_dff_B_S3MWRViv5_2;
	wire w_dff_B_6woJ4yq17_2;
	wire w_dff_B_gWBK3IYt8_2;
	wire w_dff_B_EW08QSUF0_2;
	wire w_dff_B_HA4Rymwa9_2;
	wire w_dff_B_mYgJh4cX7_2;
	wire w_dff_B_LNvUpIxx0_2;
	wire w_dff_B_WJPC9az53_2;
	wire w_dff_B_EbO6FDzF9_2;
	wire w_dff_B_ArqXoQLF0_2;
	wire w_dff_B_TLtisFvc9_1;
	wire w_dff_B_4DWvxcdV9_2;
	wire w_dff_B_QDUfMgsb6_2;
	wire w_dff_B_I3cKe1RS8_2;
	wire w_dff_B_38Gw2lzi9_2;
	wire w_dff_B_iJMeS2Cm0_2;
	wire w_dff_B_iakj3AJ72_2;
	wire w_dff_B_2MWgvuZD9_2;
	wire w_dff_B_wsEJmLXr6_2;
	wire w_dff_B_qThltIpz6_2;
	wire w_dff_B_3CfE73JL3_2;
	wire w_dff_B_prXifrhR7_2;
	wire w_dff_B_TDt9EeZK8_2;
	wire w_dff_B_mt1TfKB29_2;
	wire w_dff_B_zD6LTIp08_2;
	wire w_dff_B_iDgjAlzy6_2;
	wire w_dff_B_EyqPd3UR0_2;
	wire w_dff_B_B8BD1BdN8_2;
	wire w_dff_B_IMsAsla93_2;
	wire w_dff_B_MDHoOfON6_2;
	wire w_dff_B_4N6NNVcz9_2;
	wire w_dff_B_OsPByg8L9_2;
	wire w_dff_B_x2InN0J80_2;
	wire w_dff_B_SblAxLOd8_1;
	wire w_dff_B_OJ4JnQJB2_2;
	wire w_dff_B_wCXotfUE3_2;
	wire w_dff_B_Ra8iuUCc6_2;
	wire w_dff_B_yeuLYKfg3_2;
	wire w_dff_B_Rq33UQ3B7_2;
	wire w_dff_B_uSeNHYCW1_2;
	wire w_dff_B_w3PZDCol5_2;
	wire w_dff_B_5kWWp7NJ8_2;
	wire w_dff_B_UwMDgdMW3_2;
	wire w_dff_B_qnTPUbn78_2;
	wire w_dff_B_6zyzZOQC8_2;
	wire w_dff_B_PgSGs52k4_2;
	wire w_dff_B_eHskGCaK9_2;
	wire w_dff_B_go5r6peb2_2;
	wire w_dff_B_OVpk8ql00_2;
	wire w_dff_B_me1KJaCE9_2;
	wire w_dff_B_kJkRFspF4_2;
	wire w_dff_B_fs2yL4LS9_2;
	wire w_dff_B_9CMwoNsU4_2;
	wire w_dff_B_xdbSe9VM5_2;
	wire w_dff_B_Q47A3wZg4_1;
	wire w_dff_B_sUti06fg7_2;
	wire w_dff_B_ZX0Jhod58_2;
	wire w_dff_B_DqVoTc2B6_2;
	wire w_dff_B_dLuNtJd85_2;
	wire w_dff_B_rlsgxYi46_2;
	wire w_dff_B_KUgsDlTU6_2;
	wire w_dff_B_RMENxy5T9_2;
	wire w_dff_B_EOoiShaq7_2;
	wire w_dff_B_hLGC8ap34_2;
	wire w_dff_B_B3K2sMmk2_2;
	wire w_dff_B_4LOcEv8e6_2;
	wire w_dff_B_RLG0ZDh45_2;
	wire w_dff_B_SWs2x6MT2_2;
	wire w_dff_B_BscJFiJj4_2;
	wire w_dff_B_69Bbgfkw4_2;
	wire w_dff_B_SkcNSFnk3_2;
	wire w_dff_B_5n1qQk7e4_2;
	wire w_dff_B_aPtSe8m90_2;
	wire w_dff_B_QsGqq5Sx7_1;
	wire w_dff_B_LA0y961X7_2;
	wire w_dff_B_inGyD92K1_2;
	wire w_dff_B_Gis1xd6E8_2;
	wire w_dff_B_GepeqIs48_2;
	wire w_dff_B_IkVdo9Kj0_2;
	wire w_dff_B_bRMPDL0D9_2;
	wire w_dff_B_e6JN9olU6_2;
	wire w_dff_B_ejxohMYf3_2;
	wire w_dff_B_5eMe5wWo5_2;
	wire w_dff_B_nHBUiJmd1_2;
	wire w_dff_B_tDydL1PX0_2;
	wire w_dff_B_eliUbxDp7_2;
	wire w_dff_B_AZZw5Ixz4_2;
	wire w_dff_B_198TQkrY6_2;
	wire w_dff_B_ukWplGiy0_2;
	wire w_dff_B_ZFYsJInP3_2;
	wire w_dff_B_DrhxwjcS0_1;
	wire w_dff_B_xwJhvg0Q4_2;
	wire w_dff_B_YRwg5mzY8_2;
	wire w_dff_B_epcv4njW1_2;
	wire w_dff_B_UeM2oomk1_2;
	wire w_dff_B_0AoTfTuT7_2;
	wire w_dff_B_19FKgTfh7_2;
	wire w_dff_B_fOUEpAxL8_2;
	wire w_dff_B_otOH1XqV2_2;
	wire w_dff_B_3lFqYNwn7_2;
	wire w_dff_B_QxsNpPkw7_2;
	wire w_dff_B_RAyjpQdF9_2;
	wire w_dff_B_92SXSXjX8_2;
	wire w_dff_B_cito59mb9_2;
	wire w_dff_B_EVtxD5999_2;
	wire w_dff_B_bYy1OwRT1_1;
	wire w_dff_B_kUHza9uG2_2;
	wire w_dff_B_bhwEK5bt2_2;
	wire w_dff_B_xEUE7uo23_2;
	wire w_dff_B_tSU0Z8BE5_2;
	wire w_dff_B_ts9UJt7J1_2;
	wire w_dff_B_FFpo0OqE6_2;
	wire w_dff_B_898eVje57_2;
	wire w_dff_B_wCegv5yY3_2;
	wire w_dff_B_s3clsBNy0_2;
	wire w_dff_B_P1tqOhQ32_2;
	wire w_dff_B_R4lCshcJ5_2;
	wire w_dff_B_Jii61y7X1_2;
	wire w_dff_B_0ZsMoynN4_1;
	wire w_dff_B_J08wHF7i5_2;
	wire w_dff_B_wTmm9n9Z9_2;
	wire w_dff_B_fUYcGxKE9_2;
	wire w_dff_B_cjdPkUFn9_2;
	wire w_dff_B_2EEc9zb23_2;
	wire w_dff_B_r0OWAUOU4_2;
	wire w_dff_B_yG45ZPEJ0_2;
	wire w_dff_B_mU0vltQ72_2;
	wire w_dff_B_NbvEfiLT5_2;
	wire w_dff_B_QriFem3S1_2;
	wire w_dff_B_cgMAQ9Lj0_1;
	wire w_dff_B_IihquM6n1_2;
	wire w_dff_B_r08S5zql6_2;
	wire w_dff_B_AOOHxe6x2_2;
	wire w_dff_B_jbniQ65W6_2;
	wire w_dff_B_6bcp0QCv6_2;
	wire w_dff_B_HMIz3pOd5_2;
	wire w_dff_B_nNQVii0L1_2;
	wire w_dff_B_pfmOU5sT4_2;
	wire w_dff_B_pJf4QxHE3_2;
	wire w_dff_B_rAK4d0JX2_2;
	wire w_dff_B_YIhjSKK65_2;
	wire w_dff_B_rwjqd2Fm2_1;
	wire w_dff_B_5cMpneYK2_1;
	wire w_dff_B_Rh8AN04i2_1;
	wire w_dff_B_jkdrcr0D2_2;
	wire w_dff_B_xi23xvLP7_2;
	wire w_dff_B_tLuPYHai7_2;
	wire w_dff_B_2FbvjWma8_0;
	wire w_dff_B_Xk0MFmbp8_0;
	wire w_dff_A_T2KRF8Fd3_0;
	wire w_dff_A_rrIgy5qa0_0;
	wire w_dff_A_SeewxzKt8_1;
	wire w_dff_A_DK2WnL0g7_1;
	wire w_dff_B_s9URHH6X8_1;
	wire w_dff_A_3cdlYTgW1_1;
	wire w_dff_B_zn1GqKHr3_1;
	wire w_dff_B_JQvsXwFq0_2;
	wire w_dff_B_URcEVwNy0_2;
	wire w_dff_B_OgpRmJbk3_2;
	wire w_dff_B_ziyCwVRs9_2;
	wire w_dff_B_wJ6XdJH00_2;
	wire w_dff_B_S57zhDqo1_2;
	wire w_dff_B_hYEZKbac0_2;
	wire w_dff_B_jy0fDjNG8_2;
	wire w_dff_B_lLQpOBoG7_2;
	wire w_dff_B_SQdAL7z73_2;
	wire w_dff_B_9rilH1Ps7_2;
	wire w_dff_B_ZiIHuY8R6_2;
	wire w_dff_B_m4H2Zib90_2;
	wire w_dff_B_1Of8N5Iu2_2;
	wire w_dff_B_REQtgeSP1_2;
	wire w_dff_B_LdXGDG7H5_2;
	wire w_dff_B_gFRCuXn28_2;
	wire w_dff_B_CMUmo4SJ6_2;
	wire w_dff_B_te1iNZRa8_2;
	wire w_dff_B_WU3W2Kx24_2;
	wire w_dff_B_LOHVeOO25_2;
	wire w_dff_B_BPSUXMde2_2;
	wire w_dff_B_v4hfpko45_2;
	wire w_dff_B_jsJhMGRl9_2;
	wire w_dff_B_pziGGJK40_2;
	wire w_dff_B_QFckyIIg6_2;
	wire w_dff_B_kvjlVmal4_2;
	wire w_dff_B_RWGR07XR3_2;
	wire w_dff_B_ouzKxJNe2_2;
	wire w_dff_B_MC8JN1nJ8_2;
	wire w_dff_B_4MJdl2Ka2_2;
	wire w_dff_B_nR8Mq71c3_2;
	wire w_dff_B_txStUAdM9_2;
	wire w_dff_B_lecib16x5_2;
	wire w_dff_B_6s6jQdzQ4_2;
	wire w_dff_B_lOrHr0yL6_2;
	wire w_dff_B_albXu4Yb6_2;
	wire w_dff_B_rpETgB5D8_2;
	wire w_dff_B_8F3sj5hl8_2;
	wire w_dff_B_bWhd0JRq4_1;
	wire w_dff_B_NceV2XFZ2_2;
	wire w_dff_B_78kZyxZz5_2;
	wire w_dff_B_eeeQodBV5_2;
	wire w_dff_B_WckFnbQ17_2;
	wire w_dff_B_Y60aYXNH9_2;
	wire w_dff_B_F7flt7i61_2;
	wire w_dff_B_aPHQpUby1_2;
	wire w_dff_B_5VgjWmd19_2;
	wire w_dff_B_UT0ULpdG5_2;
	wire w_dff_B_kdmJv8NN6_2;
	wire w_dff_B_y4ilG7I21_2;
	wire w_dff_B_6IOdWjSI4_2;
	wire w_dff_B_XYk7SIV42_2;
	wire w_dff_B_19xxkGM35_2;
	wire w_dff_B_qrrEeIxw5_2;
	wire w_dff_B_CgIY4SJD4_2;
	wire w_dff_B_fGn2kFiJ4_2;
	wire w_dff_B_PaB9nUod8_2;
	wire w_dff_B_NeTfnmOb4_2;
	wire w_dff_B_X4so6oJu2_2;
	wire w_dff_B_TqlBYD1S1_2;
	wire w_dff_B_oyyBpjv97_2;
	wire w_dff_B_tus45UP17_2;
	wire w_dff_B_MWNGRxcD5_2;
	wire w_dff_B_gKDuqa6h5_2;
	wire w_dff_B_KECTLfSI4_2;
	wire w_dff_B_M3YeJXZi2_2;
	wire w_dff_B_lVdRQTMn1_2;
	wire w_dff_B_N59cVE4J0_2;
	wire w_dff_B_cFjkWjwF7_2;
	wire w_dff_B_jyqf18H51_2;
	wire w_dff_B_Enhwv3RE0_2;
	wire w_dff_B_25s2XIJY6_2;
	wire w_dff_B_WDj3OuCc4_2;
	wire w_dff_B_dAEQBR6J5_2;
	wire w_dff_B_b59aqmGd7_2;
	wire w_dff_B_8YAqrqWn5_1;
	wire w_dff_B_z1FuxEoZ7_2;
	wire w_dff_B_2G83fqto0_2;
	wire w_dff_B_Emp1WiSE6_2;
	wire w_dff_B_DUiRXHXm0_2;
	wire w_dff_B_rx6JoiWH9_2;
	wire w_dff_B_3P1mNYXI8_2;
	wire w_dff_B_0bmjbqKn5_2;
	wire w_dff_B_MPcX7RhJ4_2;
	wire w_dff_B_dH1tXWpx3_2;
	wire w_dff_B_QlCD84lh4_2;
	wire w_dff_B_vSI0pBcb5_2;
	wire w_dff_B_0rBU27UG1_2;
	wire w_dff_B_WFE0MOd79_2;
	wire w_dff_B_YU2GDSQG5_2;
	wire w_dff_B_COLJEkRH1_2;
	wire w_dff_B_5H22GFfO1_2;
	wire w_dff_B_VRca994D1_2;
	wire w_dff_B_iBgBXIzs3_2;
	wire w_dff_B_tQpIQ05D8_2;
	wire w_dff_B_7Lc2N3YZ2_2;
	wire w_dff_B_dw78O9DL3_2;
	wire w_dff_B_zBLW9VIb7_2;
	wire w_dff_B_tpwqCFhn0_2;
	wire w_dff_B_cbEmSlcb6_2;
	wire w_dff_B_qerQYLyU5_2;
	wire w_dff_B_TxbnbpcG1_2;
	wire w_dff_B_aAouONU28_2;
	wire w_dff_B_ednQk6cC7_2;
	wire w_dff_B_wGC2Ykda3_2;
	wire w_dff_B_f3tfPW3Y8_2;
	wire w_dff_B_51TE2xvk5_2;
	wire w_dff_B_KzaSQKeX0_2;
	wire w_dff_B_6C8Bv70R4_2;
	wire w_dff_B_QUxCrnrP2_1;
	wire w_dff_B_rP1iXW1r8_2;
	wire w_dff_B_QnD1NCIy0_2;
	wire w_dff_B_lXZJx7kw6_2;
	wire w_dff_B_aegVVx8D7_2;
	wire w_dff_B_v86uZsZu2_2;
	wire w_dff_B_vjD5kRak6_2;
	wire w_dff_B_YAw1nIPB6_2;
	wire w_dff_B_toWiDd1w3_2;
	wire w_dff_B_WLL8pHkl4_2;
	wire w_dff_B_7mfRIqEx2_2;
	wire w_dff_B_fzD1B09G6_2;
	wire w_dff_B_sbxtOkAn9_2;
	wire w_dff_B_Z3WGGPwF1_2;
	wire w_dff_B_1lJUoyFi6_2;
	wire w_dff_B_LjAPldJH8_2;
	wire w_dff_B_zuBMIn6I7_2;
	wire w_dff_B_UliP24vG6_2;
	wire w_dff_B_38hELelm5_2;
	wire w_dff_B_UaT7octZ7_2;
	wire w_dff_B_v7YKJnwO5_2;
	wire w_dff_B_SqqV5f6z4_2;
	wire w_dff_B_yBm3HFis9_2;
	wire w_dff_B_qmTAj92z3_2;
	wire w_dff_B_g7DhUzlX9_2;
	wire w_dff_B_S3nUjeZH4_2;
	wire w_dff_B_m13h5eZ28_2;
	wire w_dff_B_gWym8VVz4_2;
	wire w_dff_B_el1QXwkV8_2;
	wire w_dff_B_00rP6kOR2_2;
	wire w_dff_B_moEMgU2N6_2;
	wire w_dff_B_xwntQN6w4_1;
	wire w_dff_B_uYcsPNOh4_2;
	wire w_dff_B_Lbb88Srh4_2;
	wire w_dff_B_GVcNLxHD1_2;
	wire w_dff_B_jOR1uSfS4_2;
	wire w_dff_B_z6asLAyO3_2;
	wire w_dff_B_ZSgPdKQo3_2;
	wire w_dff_B_FMGVvcrv2_2;
	wire w_dff_B_YyaB3ivC3_2;
	wire w_dff_B_Codtp45X7_2;
	wire w_dff_B_yCii9u252_2;
	wire w_dff_B_c0SJOclp1_2;
	wire w_dff_B_vP2xJAAq5_2;
	wire w_dff_B_Qt7bbinK7_2;
	wire w_dff_B_3HKBN7d94_2;
	wire w_dff_B_wHT9FuGU0_2;
	wire w_dff_B_SBpJVwLh4_2;
	wire w_dff_B_apWkk9hK8_2;
	wire w_dff_B_wIsP63or6_2;
	wire w_dff_B_lrvnhKSp0_2;
	wire w_dff_B_q9RLqorR2_2;
	wire w_dff_B_CGmpFAkC5_2;
	wire w_dff_B_Oqd0DyLu0_2;
	wire w_dff_B_SpR4f3xO2_2;
	wire w_dff_B_Szq79zXu1_2;
	wire w_dff_B_37DtKQN75_2;
	wire w_dff_B_4I6PdJS70_2;
	wire w_dff_B_9jxM2aiy2_2;
	wire w_dff_B_SqZb0rTo9_1;
	wire w_dff_B_DdI2bIv10_2;
	wire w_dff_B_meL1Vto37_2;
	wire w_dff_B_WKBfIGE80_2;
	wire w_dff_B_25LFaOna2_2;
	wire w_dff_B_YZYDP54h6_2;
	wire w_dff_B_oQq1cGES4_2;
	wire w_dff_B_ASgo0ttN3_2;
	wire w_dff_B_LlRcpt7T4_2;
	wire w_dff_B_drSK7fSF8_2;
	wire w_dff_B_67RF45jC1_2;
	wire w_dff_B_KFlzZAQE5_2;
	wire w_dff_B_72El23Cr9_2;
	wire w_dff_B_1u62Iwdf3_2;
	wire w_dff_B_67EWWzgp9_2;
	wire w_dff_B_ZYYnI4144_2;
	wire w_dff_B_idU947px2_2;
	wire w_dff_B_3ur6dyIE7_2;
	wire w_dff_B_FjvmHdvz1_2;
	wire w_dff_B_uhiHv0kY0_2;
	wire w_dff_B_hBp5jCZZ7_2;
	wire w_dff_B_VKUptWK73_2;
	wire w_dff_B_Of9tL9Os1_2;
	wire w_dff_B_DBt030OO6_2;
	wire w_dff_B_LU4nYTi48_2;
	wire w_dff_B_gUK6quCH9_1;
	wire w_dff_B_QpY56Rx47_2;
	wire w_dff_B_PNGYvlUO5_2;
	wire w_dff_B_mdO820bf6_2;
	wire w_dff_B_5vTE0yNV6_2;
	wire w_dff_B_MsaBUsDF1_2;
	wire w_dff_B_l1Tc5iua5_2;
	wire w_dff_B_9rgY2KeU3_2;
	wire w_dff_B_LHsCU7050_2;
	wire w_dff_B_YELg5juV5_2;
	wire w_dff_B_wnag1YGW5_2;
	wire w_dff_B_RGDX354s5_2;
	wire w_dff_B_IYpsZfBh1_2;
	wire w_dff_B_EoQkHSsE8_2;
	wire w_dff_B_eHSpO7N86_2;
	wire w_dff_B_5RmBExgl9_2;
	wire w_dff_B_nXdZS2gZ6_2;
	wire w_dff_B_uYsqBSRN2_2;
	wire w_dff_B_3wxf5Zom0_2;
	wire w_dff_B_qZ5SdUoN1_2;
	wire w_dff_B_TeMjtAcZ2_2;
	wire w_dff_B_jbWyQ2f59_1;
	wire w_dff_B_0ba8OZ1J0_2;
	wire w_dff_B_x1vg9g3C0_2;
	wire w_dff_B_G5DtcGGA6_2;
	wire w_dff_B_VkhB4F7C5_2;
	wire w_dff_B_x04ISGZH3_2;
	wire w_dff_B_mcBgZVSX6_2;
	wire w_dff_B_lsNpgKT07_2;
	wire w_dff_B_9bQ0KpVh3_2;
	wire w_dff_B_5xfSQFPC8_2;
	wire w_dff_B_JPwgvdJI1_2;
	wire w_dff_B_d7EkmAa06_2;
	wire w_dff_B_NbpgrCmA4_2;
	wire w_dff_B_95BlcFnV7_2;
	wire w_dff_B_XUVcPYcI5_2;
	wire w_dff_B_ukNE9JBI9_2;
	wire w_dff_B_LYKAZrm17_2;
	wire w_dff_B_TiTJtm369_2;
	wire w_dff_B_wmuiS3qd6_2;
	wire w_dff_B_AvhsdWwx0_1;
	wire w_dff_B_Oh1zq6Mh6_2;
	wire w_dff_B_oHnryv4o5_2;
	wire w_dff_B_yC4jijt47_2;
	wire w_dff_B_XfYe9kqy7_2;
	wire w_dff_B_iLeXhq9f2_2;
	wire w_dff_B_OL9yJHgO8_2;
	wire w_dff_B_J7aiNuZL2_2;
	wire w_dff_B_k3gITvSR1_2;
	wire w_dff_B_YeRToyGb0_2;
	wire w_dff_B_zBJ5tJdi9_2;
	wire w_dff_B_tMeUQAr51_2;
	wire w_dff_B_vyLppwd93_2;
	wire w_dff_B_guJvyLC42_2;
	wire w_dff_B_U0qPwURo8_2;
	wire w_dff_B_7XPxFGYO7_2;
	wire w_dff_B_SbRg2T466_2;
	wire w_dff_B_jDExplnb2_1;
	wire w_dff_B_hWqmaJz68_2;
	wire w_dff_B_Au2MqRS42_2;
	wire w_dff_B_K0rMzYeN2_2;
	wire w_dff_B_dOtyYH094_2;
	wire w_dff_B_FWho8mwh2_2;
	wire w_dff_B_cFjIApdh3_2;
	wire w_dff_B_Q8cwLoy62_2;
	wire w_dff_B_dnR4MMU02_2;
	wire w_dff_B_NZ6F6M5D1_2;
	wire w_dff_B_qty4MBao8_2;
	wire w_dff_B_zJ69d5Q91_2;
	wire w_dff_B_QonhRK344_2;
	wire w_dff_B_NbIEAUxQ8_2;
	wire w_dff_B_0BghZfKE4_2;
	wire w_dff_B_ZbX2H2M93_1;
	wire w_dff_B_byeQr5fB7_2;
	wire w_dff_B_Dj2olG4I4_2;
	wire w_dff_B_kfBuFU4K3_2;
	wire w_dff_B_ZY8BgPa79_2;
	wire w_dff_B_aKEU5xNU8_2;
	wire w_dff_B_wVQ1QvgF0_2;
	wire w_dff_B_Qu8sGOb56_2;
	wire w_dff_B_GWKSrfmK5_2;
	wire w_dff_B_YleM33fm8_2;
	wire w_dff_B_WqdSsM3X2_2;
	wire w_dff_B_BvutzHhp9_2;
	wire w_dff_B_5pO8copD6_2;
	wire w_dff_B_MZbWiYZP4_1;
	wire w_dff_B_SKbly1jy3_2;
	wire w_dff_B_xuApQhmg9_2;
	wire w_dff_B_hJVRdHFJ2_2;
	wire w_dff_B_HV9xsRd55_2;
	wire w_dff_B_iHUvig0Q5_2;
	wire w_dff_B_rTbsJc0U3_2;
	wire w_dff_B_hYKJftjW7_2;
	wire w_dff_B_IcvyUOpV9_2;
	wire w_dff_B_ZX1ox3bo8_2;
	wire w_dff_B_9QT1Zgay3_2;
	wire w_dff_B_4XuRTRbF5_1;
	wire w_dff_B_Yo4caIpC5_2;
	wire w_dff_B_so2WwinY5_2;
	wire w_dff_B_dPnlfqXA4_2;
	wire w_dff_B_PtlK4VvW2_2;
	wire w_dff_B_qpBA0bLC0_2;
	wire w_dff_B_TrqQCWBP1_2;
	wire w_dff_B_p8jGFLgk1_2;
	wire w_dff_B_jSQRXVU61_2;
	wire w_dff_B_kiu8i9rh1_2;
	wire w_dff_B_2iAqGD1d5_2;
	wire w_dff_B_CWBZljMi1_2;
	wire w_dff_B_tz9i5LDL6_1;
	wire w_dff_B_0RbaoSE57_1;
	wire w_dff_B_n1Y9jby81_1;
	wire w_dff_B_KH11dAwP7_2;
	wire w_dff_B_VYk08moP0_2;
	wire w_dff_B_WlqYnXpZ5_2;
	wire w_dff_B_7RAsqCfJ4_0;
	wire w_dff_B_wbmtKYiJ5_0;
	wire w_dff_A_gMUQkBHE4_0;
	wire w_dff_A_QsWz4K3z1_0;
	wire w_dff_A_boBTgFYQ0_1;
	wire w_dff_A_5I1E6S8T8_1;
	wire w_dff_B_wMZixJ0t3_1;
	wire w_dff_A_KNttCfjm4_1;
	wire w_dff_B_B1fTr3EQ0_1;
	wire w_dff_B_IKesATjm2_2;
	wire w_dff_B_Rai0w08W8_2;
	wire w_dff_B_BHpDV6SL2_2;
	wire w_dff_B_Ic9OiRAe4_2;
	wire w_dff_B_UeY8FAKR6_2;
	wire w_dff_B_dLcPpB2E1_2;
	wire w_dff_B_i1H8cDHp2_2;
	wire w_dff_B_PGXolDR15_2;
	wire w_dff_B_4fuqVPcN6_2;
	wire w_dff_B_1fTpE24b6_2;
	wire w_dff_B_BIO2Jqv37_2;
	wire w_dff_B_z0aytx1A7_2;
	wire w_dff_B_5KqVGXXJ5_2;
	wire w_dff_B_lkRuobfB7_2;
	wire w_dff_B_pBjD1pgZ8_2;
	wire w_dff_B_KnHscsVw9_2;
	wire w_dff_B_r6oHtWmn8_2;
	wire w_dff_B_9I2K4W1T5_2;
	wire w_dff_B_EpZG7LPc1_2;
	wire w_dff_B_ezVLhejA8_2;
	wire w_dff_B_IVpYyiNX3_2;
	wire w_dff_B_gJuf6WMv4_2;
	wire w_dff_B_AyvtIffD3_2;
	wire w_dff_B_i72cYq3q2_2;
	wire w_dff_B_E2NdmMMM5_2;
	wire w_dff_B_kqNXt3mr9_2;
	wire w_dff_B_m0lY1gc95_2;
	wire w_dff_B_zWGfcJdG2_2;
	wire w_dff_B_kDVPxAXA1_2;
	wire w_dff_B_7rArwP4H7_2;
	wire w_dff_B_fF0xbfAr5_2;
	wire w_dff_B_WP6hLDlV0_2;
	wire w_dff_B_bjdS5EFx7_2;
	wire w_dff_B_WsFgGShv2_2;
	wire w_dff_B_CwW7ib2w6_2;
	wire w_dff_B_Qjjt0w3S1_2;
	wire w_dff_B_n7DXsGIr8_2;
	wire w_dff_B_6pjK2m7T6_2;
	wire w_dff_B_Nsr8LsGd2_2;
	wire w_dff_B_9jwiKTXR0_2;
	wire w_dff_B_Ds0vKPck1_1;
	wire w_dff_B_de1NgIVY0_2;
	wire w_dff_B_b5W6mgeO0_2;
	wire w_dff_B_vijT05ax8_2;
	wire w_dff_B_06ECoTsA1_2;
	wire w_dff_B_4Opjvcgd9_2;
	wire w_dff_B_e4cTjmbp1_2;
	wire w_dff_B_MxMPcwTN8_2;
	wire w_dff_B_RlxPCt5t7_2;
	wire w_dff_B_Ov1Z5Iql3_2;
	wire w_dff_B_5sW30sEJ3_2;
	wire w_dff_B_IbpwfenH7_2;
	wire w_dff_B_Hp3WxBEw7_2;
	wire w_dff_B_W7J7j9fu3_2;
	wire w_dff_B_F9xq26UU0_2;
	wire w_dff_B_uss7Niaf0_2;
	wire w_dff_B_kHcqLz9C8_2;
	wire w_dff_B_kb6HjZos8_2;
	wire w_dff_B_6AtXfxs03_2;
	wire w_dff_B_vm4lwmeR7_2;
	wire w_dff_B_kwb45Ov56_2;
	wire w_dff_B_bfdsRwPH6_2;
	wire w_dff_B_fta1R7qd2_2;
	wire w_dff_B_qKCwzhgO0_2;
	wire w_dff_B_3e0gmAiY9_2;
	wire w_dff_B_D0jj3TBw8_2;
	wire w_dff_B_3DM79s4j6_2;
	wire w_dff_B_WDkaVjEG4_2;
	wire w_dff_B_mE720zBR7_2;
	wire w_dff_B_nnSDFqqO5_2;
	wire w_dff_B_FDLpQtwo4_2;
	wire w_dff_B_IFUkFm247_2;
	wire w_dff_B_IkRLZFXu5_2;
	wire w_dff_B_htxzZT5S3_2;
	wire w_dff_B_plmIA1TV1_2;
	wire w_dff_B_gkmta5bM2_2;
	wire w_dff_B_0kbzAFr32_2;
	wire w_dff_B_jnITGK5r1_2;
	wire w_dff_B_Q2VG2qeG7_1;
	wire w_dff_B_nEq5dsI15_2;
	wire w_dff_B_bt0OS5xJ5_2;
	wire w_dff_B_u6oKuM3D1_2;
	wire w_dff_B_imPLhoGZ6_2;
	wire w_dff_B_ZBchDq5z7_2;
	wire w_dff_B_lM5YyZWH9_2;
	wire w_dff_B_2tb0n7h61_2;
	wire w_dff_B_Oqer9GfB0_2;
	wire w_dff_B_yrnLnOZL7_2;
	wire w_dff_B_OhAdsSST3_2;
	wire w_dff_B_LL7oUxp97_2;
	wire w_dff_B_CEhMRDyD3_2;
	wire w_dff_B_3GH4dFwd9_2;
	wire w_dff_B_zun5r30O1_2;
	wire w_dff_B_su6K61sy8_2;
	wire w_dff_B_YVclku7K5_2;
	wire w_dff_B_wGYrY7Cg5_2;
	wire w_dff_B_UQ2rPhQl3_2;
	wire w_dff_B_TDkYhL5f6_2;
	wire w_dff_B_cA0IyRao7_2;
	wire w_dff_B_f0MxiaFR9_2;
	wire w_dff_B_8I4XB39R3_2;
	wire w_dff_B_wq7CeCXu6_2;
	wire w_dff_B_opQ4cZJN1_2;
	wire w_dff_B_fg2oMBcn2_2;
	wire w_dff_B_0S6KNmK59_2;
	wire w_dff_B_Yut8iCD26_2;
	wire w_dff_B_Jgtdt7or8_2;
	wire w_dff_B_FEzIH7wK5_2;
	wire w_dff_B_uzfU4WN12_2;
	wire w_dff_B_ILFyqgTb3_2;
	wire w_dff_B_qEikJNAa5_2;
	wire w_dff_B_dT6I9ojo5_2;
	wire w_dff_B_SwtKcqr72_2;
	wire w_dff_B_nxmiywbP2_1;
	wire w_dff_B_8AFNGO8B9_2;
	wire w_dff_B_k8dAsls96_2;
	wire w_dff_B_vOnenEBR8_2;
	wire w_dff_B_5oqkgYQU8_2;
	wire w_dff_B_MHA9LkyP6_2;
	wire w_dff_B_uYd7uQAA2_2;
	wire w_dff_B_obDSMITW2_2;
	wire w_dff_B_FcUHe5sT9_2;
	wire w_dff_B_OfmaWxW15_2;
	wire w_dff_B_3wc7Qi0x9_2;
	wire w_dff_B_SDpKUlTa3_2;
	wire w_dff_B_NMan6Nod9_2;
	wire w_dff_B_4z1umnXB9_2;
	wire w_dff_B_iSTT3HPX3_2;
	wire w_dff_B_7M8AIg5X6_2;
	wire w_dff_B_LrYpCf1R7_2;
	wire w_dff_B_YxLPl3QV6_2;
	wire w_dff_B_8Z78ucoJ0_2;
	wire w_dff_B_xnmuVipT2_2;
	wire w_dff_B_bRI5mEBV4_2;
	wire w_dff_B_besHd5Am9_2;
	wire w_dff_B_4kyFvT3S1_2;
	wire w_dff_B_v1DaeGCN4_2;
	wire w_dff_B_BgMvkOkL8_2;
	wire w_dff_B_4X0pw1Rd1_2;
	wire w_dff_B_ULUn1tQD4_2;
	wire w_dff_B_DOpKtcWe7_2;
	wire w_dff_B_fKbJoKPM1_2;
	wire w_dff_B_6bFjw2Xa8_2;
	wire w_dff_B_2HGFSGuf0_2;
	wire w_dff_B_SGwdY6Qc1_2;
	wire w_dff_B_xWWDbt2V5_1;
	wire w_dff_B_Zp9VLfbf2_2;
	wire w_dff_B_EFB1uhlB4_2;
	wire w_dff_B_KkAXeElX0_2;
	wire w_dff_B_pBU7uFsR5_2;
	wire w_dff_B_xrXG658n7_2;
	wire w_dff_B_QQus0tLD1_2;
	wire w_dff_B_i890ZlbO2_2;
	wire w_dff_B_1ei6fAKW2_2;
	wire w_dff_B_lPb9NTqD9_2;
	wire w_dff_B_r3JIv25B6_2;
	wire w_dff_B_MI18Tut26_2;
	wire w_dff_B_vTAunJB51_2;
	wire w_dff_B_Nh55hMhd8_2;
	wire w_dff_B_gMfX8drS2_2;
	wire w_dff_B_Sgw1XGVD3_2;
	wire w_dff_B_zjpAOmYz5_2;
	wire w_dff_B_zKk2AQBO1_2;
	wire w_dff_B_cl1IGK2H5_2;
	wire w_dff_B_rFyzzYzX9_2;
	wire w_dff_B_QEKXQ2at1_2;
	wire w_dff_B_ihq9HTqP9_2;
	wire w_dff_B_6dK7vAi15_2;
	wire w_dff_B_pTUQEWkH4_2;
	wire w_dff_B_JZ6jfiZk7_2;
	wire w_dff_B_p474wezT6_2;
	wire w_dff_B_nJTIuJgD8_2;
	wire w_dff_B_jJSpxOIK5_2;
	wire w_dff_B_CDoZxnYN5_2;
	wire w_dff_B_KSa9u7fX3_1;
	wire w_dff_B_O8ThttuR1_2;
	wire w_dff_B_8XbVtm7M3_2;
	wire w_dff_B_bz3kgK1s9_2;
	wire w_dff_B_g3m4722u4_2;
	wire w_dff_B_C6JHwCTn4_2;
	wire w_dff_B_zQknoiDg3_2;
	wire w_dff_B_cjrwAAy16_2;
	wire w_dff_B_ZT48QORD5_2;
	wire w_dff_B_9TRrKChU2_2;
	wire w_dff_B_rF5I3jvX1_2;
	wire w_dff_B_6fjpsBzQ9_2;
	wire w_dff_B_pF2QIoLs7_2;
	wire w_dff_B_hkB3C7qP2_2;
	wire w_dff_B_srW537b57_2;
	wire w_dff_B_THWA969h0_2;
	wire w_dff_B_eUIPKQ0i5_2;
	wire w_dff_B_ZOnrIuSA9_2;
	wire w_dff_B_s2c5LKeV8_2;
	wire w_dff_B_MVLQcRJq6_2;
	wire w_dff_B_0fmovR7g5_2;
	wire w_dff_B_rQgWs4YS9_2;
	wire w_dff_B_M5ubFsHp0_2;
	wire w_dff_B_QTETNQ1u7_2;
	wire w_dff_B_7bG69QOm0_2;
	wire w_dff_B_E7UOXUYz1_2;
	wire w_dff_B_ilQTpZAI4_1;
	wire w_dff_B_J3V8lbAN1_2;
	wire w_dff_B_Z2z1x4vr0_2;
	wire w_dff_B_i5fCaT5J1_2;
	wire w_dff_B_537e7v9Z6_2;
	wire w_dff_B_RVQwdxHp4_2;
	wire w_dff_B_kknwGhY53_2;
	wire w_dff_B_3UdbeDpG4_2;
	wire w_dff_B_0RqoV7tA2_2;
	wire w_dff_B_wRyfyGmV4_2;
	wire w_dff_B_MnPY1HCi9_2;
	wire w_dff_B_ZK6VhDlA9_2;
	wire w_dff_B_8Seups0i3_2;
	wire w_dff_B_biwGiqmq8_2;
	wire w_dff_B_UqoCI8AX2_2;
	wire w_dff_B_7PIRpC1j4_2;
	wire w_dff_B_GOkLcsT80_2;
	wire w_dff_B_UMCmhLl18_2;
	wire w_dff_B_yXv9mCPT4_2;
	wire w_dff_B_zBUICERP7_2;
	wire w_dff_B_Jue8yMXR6_2;
	wire w_dff_B_0BpSd3x59_2;
	wire w_dff_B_3ylLCC6d3_2;
	wire w_dff_B_TabAGmhm9_1;
	wire w_dff_B_tgXSQCd49_2;
	wire w_dff_B_OGGaluAV7_2;
	wire w_dff_B_cQaYg52C4_2;
	wire w_dff_B_08lXtpOw3_2;
	wire w_dff_B_lYuarRKj4_2;
	wire w_dff_B_snQFI0HS7_2;
	wire w_dff_B_EJGpQEYm5_2;
	wire w_dff_B_22UR10zD0_2;
	wire w_dff_B_uq4tktCi1_2;
	wire w_dff_B_5KA9qhZd1_2;
	wire w_dff_B_GyAEtiNK3_2;
	wire w_dff_B_v8zYFRii9_2;
	wire w_dff_B_vc9RdmFB7_2;
	wire w_dff_B_4L7LbXtC4_2;
	wire w_dff_B_w3VKHJfC4_2;
	wire w_dff_B_OfHnQNTx9_2;
	wire w_dff_B_ONsQwoUF5_2;
	wire w_dff_B_ICXqUIyS3_2;
	wire w_dff_B_13lUOBpt4_1;
	wire w_dff_B_XE8Zla7A7_2;
	wire w_dff_B_GBagAQh26_2;
	wire w_dff_B_W7beV2HV7_2;
	wire w_dff_B_3O8S6Rkd9_2;
	wire w_dff_B_RjHMUA5g0_2;
	wire w_dff_B_hkkAbBA62_2;
	wire w_dff_B_ds5nAQBH6_2;
	wire w_dff_B_osjiGzTg8_2;
	wire w_dff_B_AjtwBvk20_2;
	wire w_dff_B_LgQc05j61_2;
	wire w_dff_B_K5V3l6oe5_2;
	wire w_dff_B_jUhFgxou5_2;
	wire w_dff_B_HPAt1UAq8_2;
	wire w_dff_B_jWGxNwRn9_2;
	wire w_dff_B_IhcHGSeE9_2;
	wire w_dff_B_cUJKJhQb6_2;
	wire w_dff_B_le5ggeC59_2;
	wire w_dff_B_rX2mSMAu1_1;
	wire w_dff_B_OBXm2lG17_2;
	wire w_dff_B_1y6ZNWQn9_2;
	wire w_dff_B_TvRm66R32_2;
	wire w_dff_B_ZPw5bUAJ7_2;
	wire w_dff_B_SwwY8paL8_2;
	wire w_dff_B_MvsfIHOT3_2;
	wire w_dff_B_HnuoiPBJ9_2;
	wire w_dff_B_LqlLr0Gf2_2;
	wire w_dff_B_7uAjTiH48_2;
	wire w_dff_B_Asfhe3Xj1_2;
	wire w_dff_B_iYfvHzZn4_2;
	wire w_dff_B_8xwOzDuu7_2;
	wire w_dff_B_S75SklB48_2;
	wire w_dff_B_SVEDSDEi2_2;
	wire w_dff_B_B4HWDCRE2_2;
	wire w_dff_B_GZxrntJy9_1;
	wire w_dff_B_Nt7NuWTH8_2;
	wire w_dff_B_2cQPzvWm4_2;
	wire w_dff_B_2wTKKPzC0_2;
	wire w_dff_B_9catRUxp6_2;
	wire w_dff_B_pVensoYy4_2;
	wire w_dff_B_xRkTMFIC1_2;
	wire w_dff_B_wY2vCz325_2;
	wire w_dff_B_lJDYlO5t0_2;
	wire w_dff_B_JXXs8xIx6_2;
	wire w_dff_B_Ims85ujk8_2;
	wire w_dff_B_RK6kbfCp8_2;
	wire w_dff_B_pMPuw8w75_2;
	wire w_dff_B_YzE7vhIp1_2;
	wire w_dff_B_fBGJNpeL5_1;
	wire w_dff_B_e2Java6M1_2;
	wire w_dff_B_Yk9pl2oQ3_2;
	wire w_dff_B_k3JCi18x8_2;
	wire w_dff_B_qozo7iat7_2;
	wire w_dff_B_jEzkYGKY5_2;
	wire w_dff_B_FNNG2QIv1_2;
	wire w_dff_B_twRhjcnr3_2;
	wire w_dff_B_KphbzRRW0_2;
	wire w_dff_B_OZt0q0Bx8_2;
	wire w_dff_B_uWR791Wt7_2;
	wire w_dff_B_biMF5xiY2_2;
	wire w_dff_B_Qy0Xl20H1_1;
	wire w_dff_B_IprDgkyj1_2;
	wire w_dff_B_6R4J12MB3_2;
	wire w_dff_B_orbJmY5M4_2;
	wire w_dff_B_VRh20Rzh3_2;
	wire w_dff_B_RLopCCLL3_2;
	wire w_dff_B_Ne3ft27P3_2;
	wire w_dff_B_p49DaM4y5_2;
	wire w_dff_B_rnVyKTkM6_2;
	wire w_dff_B_xOc774nP5_2;
	wire w_dff_B_qpgK7ctZ7_2;
	wire w_dff_B_D84DGjHM1_2;
	wire w_dff_B_LAz1Hdqf1_2;
	wire w_dff_B_N0vnEraq2_1;
	wire w_dff_B_nZWTWXa57_1;
	wire w_dff_B_7msUnWsI5_1;
	wire w_dff_B_n8ACra2z8_2;
	wire w_dff_B_UGgeFQ3J6_2;
	wire w_dff_B_M7dKjfdi0_2;
	wire w_dff_B_KltZ9xIm0_0;
	wire w_dff_B_xvpOpkG77_0;
	wire w_dff_A_hsF3NyvZ2_0;
	wire w_dff_A_uEHtC4hr1_0;
	wire w_dff_A_kP1gabiN5_1;
	wire w_dff_A_7ZLP7fsA9_1;
	wire w_dff_B_uCql4FRT2_1;
	wire w_dff_B_rl9vlxdI6_1;
	wire w_dff_B_CF2m4dVa4_1;
	wire w_dff_B_nEFS87Ai0_2;
	wire w_dff_B_QIbqq9Zi8_2;
	wire w_dff_B_Anu3fJEK1_2;
	wire w_dff_B_Ivpi194A6_2;
	wire w_dff_B_wSeg0Sqm7_2;
	wire w_dff_B_q9zeoEoj4_2;
	wire w_dff_B_NM9Z7tEL3_2;
	wire w_dff_B_21PDXfCs1_2;
	wire w_dff_B_MS6ma5TJ0_2;
	wire w_dff_B_cWTYRXaf0_2;
	wire w_dff_B_edylnqdb4_2;
	wire w_dff_B_LONx44nf7_2;
	wire w_dff_B_RoR94wHC6_2;
	wire w_dff_B_RIHJWEMA6_2;
	wire w_dff_B_p6Z4JQWe1_2;
	wire w_dff_B_OuVLpQXI4_2;
	wire w_dff_B_gRbTJOSu6_2;
	wire w_dff_B_QQT2rHBu8_2;
	wire w_dff_B_G8L7C8to9_2;
	wire w_dff_B_X5lOdO0j9_2;
	wire w_dff_B_U2tAw60L8_2;
	wire w_dff_B_S3SZhNI05_2;
	wire w_dff_B_rCREUAou5_2;
	wire w_dff_B_YVSm7Ifz7_2;
	wire w_dff_B_oeVRQQCS1_2;
	wire w_dff_B_ZBBpgqqu1_2;
	wire w_dff_B_qqdARr595_2;
	wire w_dff_B_GQTXw5KC8_2;
	wire w_dff_B_TKBP6cBN4_2;
	wire w_dff_B_mwAC1SRx8_2;
	wire w_dff_B_8CR8RnnO8_2;
	wire w_dff_B_ulpok7JF8_2;
	wire w_dff_B_IqacMjtd3_2;
	wire w_dff_B_beenyYfC7_2;
	wire w_dff_B_piiYpN3z0_2;
	wire w_dff_B_3TSunjsR5_2;
	wire w_dff_B_PApem8KO0_2;
	wire w_dff_B_w8i6ZHGt6_2;
	wire w_dff_B_4rmOztLO7_2;
	wire w_dff_B_yB2mG7uE0_2;
	wire w_dff_B_x2k9ZlQs4_2;
	wire w_dff_B_vRibU5070_2;
	wire w_dff_B_l5NVgHt94_2;
	wire w_dff_B_LK7DGMTD3_2;
	wire w_dff_B_Ov1t8lOk6_2;
	wire w_dff_B_STCDMDJq9_2;
	wire w_dff_B_4yY9eZkn0_2;
	wire w_dff_B_3JoAIAof2_2;
	wire w_dff_B_Z22TOUEK3_2;
	wire w_dff_B_TYu2qYXa0_2;
	wire w_dff_B_otr8tp1c2_2;
	wire w_dff_B_ntKPQsXT6_2;
	wire w_dff_B_KpG2wTF57_2;
	wire w_dff_B_ouQnik5Y5_2;
	wire w_dff_B_67PgEyvu6_2;
	wire w_dff_B_G0W8jHBL3_2;
	wire w_dff_B_Z3cLKKX17_2;
	wire w_dff_B_gH85watT4_2;
	wire w_dff_B_y36MB31H5_2;
	wire w_dff_B_bPibAl636_2;
	wire w_dff_B_d0fz6zrI7_2;
	wire w_dff_B_zAaED1tm9_2;
	wire w_dff_B_RPMo3dtl2_2;
	wire w_dff_B_IJpghNJq6_2;
	wire w_dff_B_qFQ5aVNJ0_2;
	wire w_dff_B_kYQP5fqt3_2;
	wire w_dff_B_wRIcmDHZ4_2;
	wire w_dff_B_rlMoE8j13_2;
	wire w_dff_B_4QJhEaaP6_2;
	wire w_dff_B_gJzLfDV48_2;
	wire w_dff_B_3GpmEY7x0_2;
	wire w_dff_B_fyRqKogp5_2;
	wire w_dff_B_fIuVZdE61_2;
	wire w_dff_B_n0RBurjJ1_2;
	wire w_dff_B_630N5O5X1_2;
	wire w_dff_B_9f3XXe5K5_2;
	wire w_dff_B_vGdWOhNZ3_2;
	wire w_dff_B_htZaDNGr6_2;
	wire w_dff_B_RkC5OAzX7_2;
	wire w_dff_B_1c0MTidD8_2;
	wire w_dff_B_JOhg4HcK6_2;
	wire w_dff_B_MVv0CSar4_2;
	wire w_dff_A_KzNFY41T9_1;
	wire w_dff_B_Ve2vwywr3_1;
	wire w_dff_B_qHbWoxwg0_2;
	wire w_dff_B_f5l68lMe1_2;
	wire w_dff_B_gx3AzOuo8_2;
	wire w_dff_B_ZPxaJen13_2;
	wire w_dff_B_aczEN2C29_2;
	wire w_dff_B_pPJprndS1_2;
	wire w_dff_B_rZ9Xi93j3_2;
	wire w_dff_B_rvuYyjHg8_2;
	wire w_dff_B_0SIpv0ki1_2;
	wire w_dff_B_KXh5epmY6_2;
	wire w_dff_B_yK5G8RGe3_2;
	wire w_dff_B_xA6472Qr1_2;
	wire w_dff_B_sRlq7t2J1_2;
	wire w_dff_B_Csq2y3z53_2;
	wire w_dff_B_DOFbZy0i6_2;
	wire w_dff_B_rtN0sDRD3_2;
	wire w_dff_B_WDkQAfWS6_2;
	wire w_dff_B_qRM52eFs1_2;
	wire w_dff_B_fyAgyzEO8_2;
	wire w_dff_B_XrFIZvxS1_2;
	wire w_dff_B_FuAHmZEw7_2;
	wire w_dff_B_KcuMKJBl7_2;
	wire w_dff_B_ctYcNkls5_2;
	wire w_dff_B_yj77zrbg3_2;
	wire w_dff_B_xe8dbRAp8_2;
	wire w_dff_B_pR0pMSR62_2;
	wire w_dff_B_xk5RLVF85_2;
	wire w_dff_B_doxSpFA06_2;
	wire w_dff_B_4xesHF4G0_2;
	wire w_dff_B_oSmfh4520_2;
	wire w_dff_B_aeVapTJW4_2;
	wire w_dff_B_uFbkJfIW6_2;
	wire w_dff_B_JlqX9ns16_2;
	wire w_dff_B_8Skiq7x46_2;
	wire w_dff_B_3fns5Lo26_2;
	wire w_dff_B_waS7hUIH8_2;
	wire w_dff_B_le8oUxGK1_2;
	wire w_dff_B_YBxTBeR39_2;
	wire w_dff_B_ZRLwk30u8_2;
	wire w_dff_B_Dj7xdSpz2_2;
	wire w_dff_B_3auqZdgw9_1;
	wire w_dff_B_zYTpJKxQ4_1;
	wire w_dff_B_sg2mavvN5_2;
	wire w_dff_B_pS9fdlhH7_2;
	wire w_dff_B_9WDbVEhb6_2;
	wire w_dff_B_LJyNPkMQ0_2;
	wire w_dff_B_az27IJQC9_2;
	wire w_dff_B_1tDdINop6_2;
	wire w_dff_B_tRMX78DR5_2;
	wire w_dff_B_gE9WwGEE1_2;
	wire w_dff_B_Qw11cTgW3_2;
	wire w_dff_B_AbhvIrOf0_2;
	wire w_dff_B_i6TYpp8K0_2;
	wire w_dff_B_pFrzBEDu3_2;
	wire w_dff_B_aFwl7LdJ1_2;
	wire w_dff_B_0s1wmtCy3_2;
	wire w_dff_B_dWLZ40NO8_2;
	wire w_dff_B_qsU24Evg2_2;
	wire w_dff_B_VDvOjBsC3_2;
	wire w_dff_B_76rPRpns2_2;
	wire w_dff_B_NKPJvvii0_2;
	wire w_dff_B_wrnUSibZ5_2;
	wire w_dff_B_shyQeqna7_2;
	wire w_dff_B_fLAw8DzZ7_2;
	wire w_dff_B_0ovuIvrH5_2;
	wire w_dff_B_KDWTfekR0_2;
	wire w_dff_B_u834emlC2_2;
	wire w_dff_B_zNgEH4H47_2;
	wire w_dff_B_GnDBeocX5_2;
	wire w_dff_B_0WHItFsX6_2;
	wire w_dff_B_g2jzKlfp2_2;
	wire w_dff_B_3UH7pmWz8_2;
	wire w_dff_B_1yogI9wc9_2;
	wire w_dff_B_i3akOtyD8_2;
	wire w_dff_B_mr21e1yZ7_2;
	wire w_dff_B_R1t0GcMK1_2;
	wire w_dff_B_g2WeaEwB7_2;
	wire w_dff_B_3qezBYm26_2;
	wire w_dff_B_NcT0JcZ80_2;
	wire w_dff_B_8mc1lKV28_2;
	wire w_dff_B_GqPxBzMg0_2;
	wire w_dff_B_cr1DQ78h8_2;
	wire w_dff_B_ejgrpTFk1_2;
	wire w_dff_B_KqKqP7oH3_2;
	wire w_dff_B_uEsFci2l2_2;
	wire w_dff_B_5Tf6ZIM33_2;
	wire w_dff_B_smSF9p9H3_2;
	wire w_dff_B_gHaagsHU1_2;
	wire w_dff_B_6NzrWgCe6_2;
	wire w_dff_B_bWlLog5T2_2;
	wire w_dff_B_D1lVgHXe2_2;
	wire w_dff_B_Z40MKTgI9_2;
	wire w_dff_B_NDIuvHeO9_2;
	wire w_dff_B_ukxLGKj71_2;
	wire w_dff_B_lOpKA3VI3_2;
	wire w_dff_B_iTRW5P7E6_2;
	wire w_dff_B_qmBRteou8_2;
	wire w_dff_B_nRGPhBnc5_2;
	wire w_dff_B_4DovabGS0_2;
	wire w_dff_B_OVLMxxRT3_2;
	wire w_dff_B_IC4EYiKF8_2;
	wire w_dff_B_qzb9UkMo0_2;
	wire w_dff_B_eC85rIfO7_2;
	wire w_dff_B_ROHnfLMl0_2;
	wire w_dff_B_5SCm5VnK6_2;
	wire w_dff_B_K5y9wFPd3_2;
	wire w_dff_B_ptXQ1yug0_2;
	wire w_dff_B_4szw6T7j3_2;
	wire w_dff_B_Nm2Dtv0K2_2;
	wire w_dff_B_k9cqx16A9_2;
	wire w_dff_B_dEjuMNy99_2;
	wire w_dff_B_CAAMQcNK6_2;
	wire w_dff_B_tBM7LcQZ8_2;
	wire w_dff_B_h5pPy9Gq6_2;
	wire w_dff_B_U4BB5Ajd1_2;
	wire w_dff_B_Eh7djlWD7_2;
	wire w_dff_B_dh6cliBu6_2;
	wire w_dff_B_N7U1sZEN0_2;
	wire w_dff_B_QmpOAylZ8_2;
	wire w_dff_B_OVlA1riG1_1;
	wire w_dff_B_PudRumwI7_2;
	wire w_dff_B_G7WhFNlR7_2;
	wire w_dff_B_nHiYpvdv8_2;
	wire w_dff_B_dMAIWCWd5_2;
	wire w_dff_B_TV2lb9Qr7_2;
	wire w_dff_B_VfEjBzbS8_2;
	wire w_dff_B_EoPzviLr0_2;
	wire w_dff_B_HIUk1tbM9_2;
	wire w_dff_B_ID0UXKTq4_2;
	wire w_dff_B_5HarhjlT8_2;
	wire w_dff_B_WWeK4A9S3_2;
	wire w_dff_B_PWt0oHi46_2;
	wire w_dff_B_c5udqjXK0_2;
	wire w_dff_B_Y8UO8W862_2;
	wire w_dff_B_R83J7hPy8_2;
	wire w_dff_B_vYn5Rclj8_2;
	wire w_dff_B_q4gNGTDk7_2;
	wire w_dff_B_UAqestjT4_2;
	wire w_dff_B_4pQ4nEZ16_2;
	wire w_dff_B_CpkOYcdb4_2;
	wire w_dff_B_KRDvAaAB4_2;
	wire w_dff_B_YgcIZrnC6_2;
	wire w_dff_B_HGXYVM893_2;
	wire w_dff_B_rBz5WxrJ7_2;
	wire w_dff_B_Ss2BhEF81_2;
	wire w_dff_B_97g0Y8sw0_2;
	wire w_dff_B_MCCsQti76_2;
	wire w_dff_B_QJUaVTYR3_2;
	wire w_dff_B_3Vz9W5ri0_2;
	wire w_dff_B_FSODxsAg3_2;
	wire w_dff_B_yxrmKJhF4_2;
	wire w_dff_B_WqiElvCE5_2;
	wire w_dff_B_zaSjiBXE9_2;
	wire w_dff_B_IeF7Vl8X5_2;
	wire w_dff_B_ljm25N4D4_2;
	wire w_dff_B_5PF1bY5k4_2;
	wire w_dff_B_esALD8hJ7_2;
	wire w_dff_B_4ekOZUDN9_1;
	wire w_dff_B_C8UvJwn70_1;
	wire w_dff_B_VL9gpHbR8_2;
	wire w_dff_B_bvMksMx30_2;
	wire w_dff_B_lGOzT4o96_2;
	wire w_dff_B_eOwLewQw7_2;
	wire w_dff_B_2vA37C663_2;
	wire w_dff_B_DHJz70dY1_2;
	wire w_dff_B_5s2bCycI7_2;
	wire w_dff_B_a9twzAqb3_2;
	wire w_dff_B_JX562nkH3_2;
	wire w_dff_B_TydahiC79_2;
	wire w_dff_B_mUI8mGD98_2;
	wire w_dff_B_Aow0IKm28_2;
	wire w_dff_B_T10lSKPT1_2;
	wire w_dff_B_smu5n5i33_2;
	wire w_dff_B_5TYoeds34_2;
	wire w_dff_B_vMzbbPHs7_2;
	wire w_dff_B_LQS0kSTl9_2;
	wire w_dff_B_fnOuQwx36_2;
	wire w_dff_B_Z7k21gL23_2;
	wire w_dff_B_pPR7WpkX7_2;
	wire w_dff_B_9ORiV7NU0_2;
	wire w_dff_B_HZwUXxkj2_2;
	wire w_dff_B_29q95w5m4_2;
	wire w_dff_B_MGAjrWON1_2;
	wire w_dff_B_kGciZmGr4_2;
	wire w_dff_B_iKgUAloo5_2;
	wire w_dff_B_BaJPbYQH2_2;
	wire w_dff_B_1DBghht21_2;
	wire w_dff_B_Qu9kvEKb1_2;
	wire w_dff_B_1lmnw1El5_2;
	wire w_dff_B_6sUrJhUZ5_2;
	wire w_dff_B_NpxVmRyW3_2;
	wire w_dff_B_Pri80Zi09_2;
	wire w_dff_B_yP0NFXiX9_2;
	wire w_dff_B_Woql476Z1_2;
	wire w_dff_B_A2JzMxBB2_2;
	wire w_dff_B_r20sFKo12_2;
	wire w_dff_B_oleP03xa7_2;
	wire w_dff_B_21qc8pcD9_2;
	wire w_dff_B_UuZnL1N34_2;
	wire w_dff_B_ymgo2JbN4_2;
	wire w_dff_B_HjrqiORL1_2;
	wire w_dff_B_TSQbmhJl4_2;
	wire w_dff_B_9LJN5TX37_2;
	wire w_dff_B_8I0wKCJG3_2;
	wire w_dff_B_j0dfOK7A1_2;
	wire w_dff_B_f5KTIVCu3_2;
	wire w_dff_B_83Vm3xNJ7_2;
	wire w_dff_B_hPb3wsOR0_2;
	wire w_dff_B_9etpv8vD6_2;
	wire w_dff_B_UemEuhga8_2;
	wire w_dff_B_F44TWHRK4_2;
	wire w_dff_B_ZQKdpPTj7_2;
	wire w_dff_B_pKHb5SW60_2;
	wire w_dff_B_JVTya3gm1_2;
	wire w_dff_B_rF4N1plO2_2;
	wire w_dff_B_Zz8qDjjB5_2;
	wire w_dff_B_NT0WVFNs6_2;
	wire w_dff_B_Qy6zbgpi8_2;
	wire w_dff_B_3nhjBr1H5_2;
	wire w_dff_B_FTJWA3Wb0_2;
	wire w_dff_B_xsiyaY1M4_2;
	wire w_dff_B_LRvlqsUy2_2;
	wire w_dff_B_VyxlMqUh6_2;
	wire w_dff_B_pCqbXJPl6_2;
	wire w_dff_B_frj9NEkF7_2;
	wire w_dff_B_jZ2hx3oF8_2;
	wire w_dff_B_yqHE6R9N4_2;
	wire w_dff_B_dQZqkU7Z0_2;
	wire w_dff_B_ooyi4Dhj8_2;
	wire w_dff_B_uKa30N7n8_2;
	wire w_dff_B_KAPZZ2M51_1;
	wire w_dff_B_8KQSmLxP1_2;
	wire w_dff_B_cnm4pNU53_2;
	wire w_dff_B_NFKLhRmT6_2;
	wire w_dff_B_1PDCU8Ch8_2;
	wire w_dff_B_EFICxePJ5_2;
	wire w_dff_B_Rnrr9CHp0_2;
	wire w_dff_B_insuvd4Z9_2;
	wire w_dff_B_9nTySo4Z6_2;
	wire w_dff_B_xMufBLpJ6_2;
	wire w_dff_B_QbNkok730_2;
	wire w_dff_B_uqRpqt195_2;
	wire w_dff_B_Tia6Esri0_2;
	wire w_dff_B_XtenYsO29_2;
	wire w_dff_B_2uom0cBa3_2;
	wire w_dff_B_b25gftLS0_2;
	wire w_dff_B_R5PNm0si2_2;
	wire w_dff_B_0PFFGdyc2_2;
	wire w_dff_B_dsgKG87Q3_2;
	wire w_dff_B_seZZcPUD7_2;
	wire w_dff_B_UbrrY6Uw3_2;
	wire w_dff_B_PkNCOy2u6_2;
	wire w_dff_B_yWPTjqYi3_2;
	wire w_dff_B_XTqvdSER0_2;
	wire w_dff_B_blvJ59RF3_2;
	wire w_dff_B_3eWlahs43_2;
	wire w_dff_B_kqu4Jbls1_2;
	wire w_dff_B_YYwiy0Yh6_2;
	wire w_dff_B_xl5dLPUD7_2;
	wire w_dff_B_qvUOXcKk3_2;
	wire w_dff_B_k0Ka6w7K9_2;
	wire w_dff_B_WQwh4vy97_2;
	wire w_dff_B_R44vQg6Q5_2;
	wire w_dff_B_DhdwAVrR1_2;
	wire w_dff_B_ng7MdjRo8_2;
	wire w_dff_B_CFkAHw0j4_1;
	wire w_dff_B_wQmsM3qk1_1;
	wire w_dff_B_2HXbBIk07_2;
	wire w_dff_B_HBJaj7QS8_2;
	wire w_dff_B_AHSOSasA8_2;
	wire w_dff_B_kDCWsug17_2;
	wire w_dff_B_EaZG6X1D3_2;
	wire w_dff_B_YvPlzF8T3_2;
	wire w_dff_B_lVGBjZCS0_2;
	wire w_dff_B_ZmA2cTQN0_2;
	wire w_dff_B_C6pjOZAS9_2;
	wire w_dff_B_GOdzJMOV5_2;
	wire w_dff_B_HBgPADSC2_2;
	wire w_dff_B_Nbebmnft4_2;
	wire w_dff_B_xLOns4jM0_2;
	wire w_dff_B_6lmMNMfw7_2;
	wire w_dff_B_PgY44oFz5_2;
	wire w_dff_B_N1XXNetg8_2;
	wire w_dff_B_aSey69M92_2;
	wire w_dff_B_opsKTvnQ6_2;
	wire w_dff_B_Q5gwx0sm8_2;
	wire w_dff_B_5CLvqqWM2_2;
	wire w_dff_B_48RxOUUx8_2;
	wire w_dff_B_Cz1MBfmd8_2;
	wire w_dff_B_trv2bQy57_2;
	wire w_dff_B_DRpjh5Yl3_2;
	wire w_dff_B_qe0x86h46_2;
	wire w_dff_B_iCjHO4bM6_2;
	wire w_dff_B_rPKcuSzv0_2;
	wire w_dff_B_q1QBB7zv9_2;
	wire w_dff_B_SrxSrW0G3_2;
	wire w_dff_B_wNjID34g5_2;
	wire w_dff_B_J7N8fnvp0_2;
	wire w_dff_B_nFvh7y3i3_2;
	wire w_dff_B_i0Yvv1N56_2;
	wire w_dff_B_IQO3mTKG1_2;
	wire w_dff_B_3v0ADI9U9_2;
	wire w_dff_B_SBtpTMJZ5_2;
	wire w_dff_B_CNvUG9B36_2;
	wire w_dff_B_XKkhD4X06_2;
	wire w_dff_B_U0yjbSxp9_2;
	wire w_dff_B_MJHupzjb4_2;
	wire w_dff_B_dNBU1pdN0_2;
	wire w_dff_B_WyXfI5dU9_2;
	wire w_dff_B_qyILnLYn9_2;
	wire w_dff_B_DEw2b6Ni3_2;
	wire w_dff_B_CcSxBsZl0_2;
	wire w_dff_B_mfXXv0Vv0_2;
	wire w_dff_B_Ze9ugTDp0_2;
	wire w_dff_B_fpkHUbGs2_2;
	wire w_dff_B_DLqJCdGJ9_2;
	wire w_dff_B_eysHXuh48_2;
	wire w_dff_B_NrQ5MYUw1_2;
	wire w_dff_B_DKVkEJvC0_2;
	wire w_dff_B_LCT4YpCV1_2;
	wire w_dff_B_VHjWto203_2;
	wire w_dff_B_C9jrjA3o5_2;
	wire w_dff_B_26Q163G92_2;
	wire w_dff_B_uuzQMzJQ0_2;
	wire w_dff_B_Io0IbmwZ1_2;
	wire w_dff_B_aBRr0VjG5_2;
	wire w_dff_B_xgmijSJq7_2;
	wire w_dff_B_z7L8DSGO5_2;
	wire w_dff_B_11QQPtNf5_2;
	wire w_dff_B_D8krU0Ys7_2;
	wire w_dff_B_5MEgAAAv1_2;
	wire w_dff_B_FwikrSQf0_2;
	wire w_dff_B_sTlKSnnr0_1;
	wire w_dff_B_UWIdUfXK9_2;
	wire w_dff_B_qWDmvnZ22_2;
	wire w_dff_B_KxwnxxyK8_2;
	wire w_dff_B_ctu5O80e3_2;
	wire w_dff_B_ybng71f38_2;
	wire w_dff_B_aVfBNds87_2;
	wire w_dff_B_T3Kn75uS2_2;
	wire w_dff_B_JIrNpzIs4_2;
	wire w_dff_B_q1fXV2007_2;
	wire w_dff_B_lfstOxSI8_2;
	wire w_dff_B_Yw8iH4jl4_2;
	wire w_dff_B_6i0tAEd47_2;
	wire w_dff_B_Rl8xE0iy2_2;
	wire w_dff_B_PE1WyJXc6_2;
	wire w_dff_B_fwnWuWeg8_2;
	wire w_dff_B_RwL3Twf68_2;
	wire w_dff_B_NQRY5bSM3_2;
	wire w_dff_B_oD7Naomz3_2;
	wire w_dff_B_CqULvryu6_2;
	wire w_dff_B_OPL3znrp7_2;
	wire w_dff_B_JLRnP7sD5_2;
	wire w_dff_B_uZBsouB98_2;
	wire w_dff_B_Zg290EZQ2_2;
	wire w_dff_B_PixasGwK6_2;
	wire w_dff_B_DyJhSiRb9_2;
	wire w_dff_B_KcHzvtVe1_2;
	wire w_dff_B_wBXmdGKi8_2;
	wire w_dff_B_j8eaVuxS5_2;
	wire w_dff_B_wa4oXp9q4_2;
	wire w_dff_B_zxwx0PPF5_2;
	wire w_dff_B_hapB8zjH4_2;
	wire w_dff_B_CwM0rPiB5_1;
	wire w_dff_B_OLhctYmw4_1;
	wire w_dff_B_aKCpI4W40_2;
	wire w_dff_B_vg6D0js49_2;
	wire w_dff_B_fKiiRoqR3_2;
	wire w_dff_B_6IGJbsmP9_2;
	wire w_dff_B_NbgeeVgi4_2;
	wire w_dff_B_f3PwT8SZ4_2;
	wire w_dff_B_g0Si6Fu99_2;
	wire w_dff_B_f53rVkJu8_2;
	wire w_dff_B_0115tIk78_2;
	wire w_dff_B_637iVEJW7_2;
	wire w_dff_B_MuNNHNug7_2;
	wire w_dff_B_FoGxD9Oo3_2;
	wire w_dff_B_zm6CwYB79_2;
	wire w_dff_B_wN5lUYCb0_2;
	wire w_dff_B_scVsnS9Q6_2;
	wire w_dff_B_8aYoBSwx4_2;
	wire w_dff_B_Zi1D8kvU1_2;
	wire w_dff_B_7WdZfxw69_2;
	wire w_dff_B_wXT84iJF5_2;
	wire w_dff_B_lyGKtdyx4_2;
	wire w_dff_B_NfaMFL8B7_2;
	wire w_dff_B_G8oGNQ6C3_2;
	wire w_dff_B_CsFmnnYz9_2;
	wire w_dff_B_fJvYJ8zi7_2;
	wire w_dff_B_LmyQWHIX7_2;
	wire w_dff_B_UmN3Dyph0_2;
	wire w_dff_B_uTsoFDaG1_2;
	wire w_dff_B_FpLZbDWC4_2;
	wire w_dff_B_6dtxSjAr8_2;
	wire w_dff_B_EuWd9ZeP3_2;
	wire w_dff_B_qOayzeZa8_2;
	wire w_dff_B_oXfcGFna4_2;
	wire w_dff_B_f2F0H5Y09_2;
	wire w_dff_B_BPBtebEC6_2;
	wire w_dff_B_OUoVzMya5_2;
	wire w_dff_B_t4mGRhEk9_2;
	wire w_dff_B_AmJDgoIR5_2;
	wire w_dff_B_lxgtwjMq4_2;
	wire w_dff_B_xSR5WsxF3_2;
	wire w_dff_B_oAXnSN2Q4_2;
	wire w_dff_B_YBJjziKd2_2;
	wire w_dff_B_IUtx9uST3_2;
	wire w_dff_B_ynu59tw81_2;
	wire w_dff_B_CXdOWRCV6_2;
	wire w_dff_B_PAc7A3W79_2;
	wire w_dff_B_1oRHhMWH2_2;
	wire w_dff_B_ratrjSTf6_2;
	wire w_dff_B_tOKyTNL04_2;
	wire w_dff_B_OucVIWuq3_2;
	wire w_dff_B_898IZUov7_2;
	wire w_dff_B_9m1alUI77_2;
	wire w_dff_B_Nx1ICzwB2_2;
	wire w_dff_B_oYuSsp4l1_2;
	wire w_dff_B_dsxpN8f92_2;
	wire w_dff_B_3EZMwyX26_2;
	wire w_dff_B_ns77EYFo5_2;
	wire w_dff_B_YqiDvoCs3_2;
	wire w_dff_B_oOKqRdP05_2;
	wire w_dff_B_r3huhRxb0_2;
	wire w_dff_B_axwawoWk7_1;
	wire w_dff_B_pP1zO1dr1_2;
	wire w_dff_B_1jCzbY4i8_2;
	wire w_dff_B_zSpTN13E8_2;
	wire w_dff_B_BCucj8Jg2_2;
	wire w_dff_B_x9OfUCI92_2;
	wire w_dff_B_zn8hKTYi2_2;
	wire w_dff_B_WbuKOWZA5_2;
	wire w_dff_B_x5OgFASA0_2;
	wire w_dff_B_OqcEM6ry9_2;
	wire w_dff_B_VLBYan4f1_2;
	wire w_dff_B_CVeCeV9d8_2;
	wire w_dff_B_AYgZOObA1_2;
	wire w_dff_B_SWGQD5jE1_2;
	wire w_dff_B_8VMFlyWQ0_2;
	wire w_dff_B_Wt2wet0t6_2;
	wire w_dff_B_DMmIc6Li5_2;
	wire w_dff_B_17kVzHi07_2;
	wire w_dff_B_FWHTRLI31_2;
	wire w_dff_B_22KYK1pL5_2;
	wire w_dff_B_ClQDiSsc0_2;
	wire w_dff_B_yld00TSB7_2;
	wire w_dff_B_3sWcS0aT0_2;
	wire w_dff_B_32dytsvL2_2;
	wire w_dff_B_sRhPOV9Q7_2;
	wire w_dff_B_563zx3iX4_2;
	wire w_dff_B_o1oX2fjh2_2;
	wire w_dff_B_GG2ipBND6_2;
	wire w_dff_B_NpD8YZJA9_2;
	wire w_dff_B_KKo5uyzD1_1;
	wire w_dff_B_fUp5carD2_1;
	wire w_dff_B_iuKMDIcm1_2;
	wire w_dff_B_kjd9Dbyd1_2;
	wire w_dff_B_LDfN8eSa4_2;
	wire w_dff_B_nb5uT2GN5_2;
	wire w_dff_B_MLiRERpH6_2;
	wire w_dff_B_CduGgfau2_2;
	wire w_dff_B_NOSdq8cy0_2;
	wire w_dff_B_psunIQm47_2;
	wire w_dff_B_g2p7kXZc7_2;
	wire w_dff_B_B9lEuDsJ1_2;
	wire w_dff_B_y8oDhhuJ9_2;
	wire w_dff_B_xoodPjTG1_2;
	wire w_dff_B_0Mxu5Yft5_2;
	wire w_dff_B_Iwdzmfmy4_2;
	wire w_dff_B_99z39qjD3_2;
	wire w_dff_B_5FhJnfHY4_2;
	wire w_dff_B_X2idDRtj5_2;
	wire w_dff_B_XmqUqcaC9_2;
	wire w_dff_B_2fHsdkNh4_2;
	wire w_dff_B_qjpn0hwI8_2;
	wire w_dff_B_qObceB4j2_2;
	wire w_dff_B_jKouMlbX3_2;
	wire w_dff_B_SN1cEEHf9_2;
	wire w_dff_B_6h0sUWPv7_2;
	wire w_dff_B_gw1iOXXp7_2;
	wire w_dff_B_PiVM0ds34_2;
	wire w_dff_B_AeGB050M3_2;
	wire w_dff_B_6fe1ZZT72_2;
	wire w_dff_B_rbQzXhv49_2;
	wire w_dff_B_vpNtrClQ6_2;
	wire w_dff_B_zvCYuRT76_2;
	wire w_dff_B_6Wx6rueF9_2;
	wire w_dff_B_KywE32Fx1_2;
	wire w_dff_B_1leBmKF44_2;
	wire w_dff_B_2CqPL4yi0_2;
	wire w_dff_B_bMIAaMpA3_2;
	wire w_dff_B_QnRjZRUk0_2;
	wire w_dff_B_JEyLHMLm2_2;
	wire w_dff_B_4cANnGjV0_2;
	wire w_dff_B_BEziTMNN8_2;
	wire w_dff_B_HVJ59YLJ0_2;
	wire w_dff_B_4wvzxoic9_2;
	wire w_dff_B_BXTrh1J06_2;
	wire w_dff_B_xPlDu62I3_2;
	wire w_dff_B_Uva3JQDW0_2;
	wire w_dff_B_MluYXu587_2;
	wire w_dff_B_izJ6VbzU4_2;
	wire w_dff_B_gvN8qU1Z6_2;
	wire w_dff_B_YJrWGonY4_2;
	wire w_dff_B_IKiF4pOz3_2;
	wire w_dff_B_h1fyl2iW6_2;
	wire w_dff_B_1PFggV3Q2_2;
	wire w_dff_B_dfw6ZqK21_2;
	wire w_dff_B_MNUGWboP9_1;
	wire w_dff_B_0FQo1S0N8_2;
	wire w_dff_B_0Nobq94l0_2;
	wire w_dff_B_zSUR7HNA1_2;
	wire w_dff_B_xKJKMDGg2_2;
	wire w_dff_B_E41MIQhv0_2;
	wire w_dff_B_kQUQvBjL9_2;
	wire w_dff_B_HSEdLmDn3_2;
	wire w_dff_B_kfrP14b15_2;
	wire w_dff_B_O4Z4dzXu5_2;
	wire w_dff_B_oXCel9BL5_2;
	wire w_dff_B_Wn3kuzJG9_2;
	wire w_dff_B_23vHAYbw4_2;
	wire w_dff_B_KGTKr7ge0_2;
	wire w_dff_B_BGuARwc99_2;
	wire w_dff_B_tfGD2nFJ5_2;
	wire w_dff_B_ueNhaTmM7_2;
	wire w_dff_B_mtdXUTWK2_2;
	wire w_dff_B_5i8l131f1_2;
	wire w_dff_B_YXIQprDs0_2;
	wire w_dff_B_jhqLoEnP6_2;
	wire w_dff_B_Hk8ERIAI0_2;
	wire w_dff_B_j1tesltt5_2;
	wire w_dff_B_D39jm4sr1_2;
	wire w_dff_B_73KkxonX6_2;
	wire w_dff_B_3is5bFk90_2;
	wire w_dff_B_7mXJf0NA4_1;
	wire w_dff_B_rttLFnrN8_1;
	wire w_dff_B_20s5XONc9_2;
	wire w_dff_B_qHSG2b0c2_2;
	wire w_dff_B_ozevfPr46_2;
	wire w_dff_B_tkztgueh7_2;
	wire w_dff_B_uIfNoRPO2_2;
	wire w_dff_B_kRscPPRT2_2;
	wire w_dff_B_KhBHrXpY8_2;
	wire w_dff_B_6xGnlLq75_2;
	wire w_dff_B_dY5jxuO90_2;
	wire w_dff_B_D9bl3EcE9_2;
	wire w_dff_B_XYcQzRBz0_2;
	wire w_dff_B_URmY6v2R1_2;
	wire w_dff_B_sRD6j7Au3_2;
	wire w_dff_B_qvKa0wlw2_2;
	wire w_dff_B_iVO4tvig4_2;
	wire w_dff_B_IndCUCZF0_2;
	wire w_dff_B_TUXIBF0o1_2;
	wire w_dff_B_cTJkwEs64_2;
	wire w_dff_B_tHwxoFyi4_2;
	wire w_dff_B_UMOLD7XV5_2;
	wire w_dff_B_LxCUjF5H4_2;
	wire w_dff_B_eNP0hdtM1_2;
	wire w_dff_B_At0fZjz30_2;
	wire w_dff_B_A8uaYMKH2_2;
	wire w_dff_B_9gSPDxPc3_2;
	wire w_dff_B_djnkdzhD1_2;
	wire w_dff_B_RZ6YHp8E5_2;
	wire w_dff_B_MrqTEaHc6_2;
	wire w_dff_B_ev7Cdmy02_2;
	wire w_dff_B_COY2pKfh3_2;
	wire w_dff_B_QxQ2Sil13_2;
	wire w_dff_B_aiUSp1hR8_2;
	wire w_dff_B_QHXE6YZV1_2;
	wire w_dff_B_9wZfYbvL5_2;
	wire w_dff_B_uyhzLsEX9_2;
	wire w_dff_B_sgHepmNT8_2;
	wire w_dff_B_NKZjq98n6_2;
	wire w_dff_B_eoCahL8F1_2;
	wire w_dff_B_nTkXefiU5_2;
	wire w_dff_B_MIMdLjjW5_2;
	wire w_dff_B_lqViAUl30_2;
	wire w_dff_B_BZLKrAKe3_2;
	wire w_dff_B_Vh0D3MO12_2;
	wire w_dff_B_4hr0prvr4_2;
	wire w_dff_B_XSo3QIbe5_2;
	wire w_dff_B_SMT7j2uL7_2;
	wire w_dff_B_Tq1QvZat2_2;
	wire w_dff_B_UvPqCIej8_1;
	wire w_dff_B_W4KPgvEX4_2;
	wire w_dff_B_Uj9cySuM9_2;
	wire w_dff_B_CUMaRmay7_2;
	wire w_dff_B_pT4qGwsF0_2;
	wire w_dff_B_TvVosUeW1_2;
	wire w_dff_B_eA7Hi7LT6_2;
	wire w_dff_B_ngp5YqPy1_2;
	wire w_dff_B_F1D5UxXN3_2;
	wire w_dff_B_JyZ1M5lM7_2;
	wire w_dff_B_D0oT6NFZ3_2;
	wire w_dff_B_96Iv5nAP6_2;
	wire w_dff_B_iiEZY4z92_2;
	wire w_dff_B_74D5P7Ff4_2;
	wire w_dff_B_l8YfPTvn9_2;
	wire w_dff_B_4li1DH5p5_2;
	wire w_dff_B_fvkDwzAC3_2;
	wire w_dff_B_qyBezgsw6_2;
	wire w_dff_B_NijD4bqu9_2;
	wire w_dff_B_pIolcipT8_2;
	wire w_dff_B_VJZIoWdv9_2;
	wire w_dff_B_XNvcYRId0_2;
	wire w_dff_B_srWxmUGH1_2;
	wire w_dff_B_ckPjZXWm5_1;
	wire w_dff_B_H9FA1TvV4_1;
	wire w_dff_B_tXZbOlXK6_2;
	wire w_dff_B_Jwe3YR9W9_2;
	wire w_dff_B_uPHo45gm7_2;
	wire w_dff_B_kY3p7xUl8_2;
	wire w_dff_B_nsmmMEq34_2;
	wire w_dff_B_V35ZtRIk6_2;
	wire w_dff_B_l54mtnv53_2;
	wire w_dff_B_VWcvLOD40_2;
	wire w_dff_B_jAqZAYch5_2;
	wire w_dff_B_eLy6O99I6_2;
	wire w_dff_B_WG0M3gtT3_2;
	wire w_dff_B_znoe0lDQ7_2;
	wire w_dff_B_zGe1Xepb8_2;
	wire w_dff_B_SFrvPMuE3_2;
	wire w_dff_B_zY0wbfHt5_2;
	wire w_dff_B_bJHjr5z51_2;
	wire w_dff_B_j7mYsTgd0_2;
	wire w_dff_B_mA9KAMsF1_2;
	wire w_dff_B_iQjh87NT6_2;
	wire w_dff_B_jvcr6p3n7_2;
	wire w_dff_B_xNRjuCEd0_2;
	wire w_dff_B_VgK0fkjq6_2;
	wire w_dff_B_aVSHeBJJ3_2;
	wire w_dff_B_SZCVgi9k8_2;
	wire w_dff_B_HSgFmTUo9_2;
	wire w_dff_B_aCQJyS167_2;
	wire w_dff_B_EEAkD4rO9_2;
	wire w_dff_B_FPsrj22g8_2;
	wire w_dff_B_Yvglu0PZ3_2;
	wire w_dff_B_vEj4vuNa3_2;
	wire w_dff_B_2ck013Mi6_2;
	wire w_dff_B_g1lbKyY67_2;
	wire w_dff_B_h71LZwRD9_2;
	wire w_dff_B_jfWebrkp7_2;
	wire w_dff_B_RB8ktwhb8_2;
	wire w_dff_B_wvrPjaGA6_2;
	wire w_dff_B_dOxhdNAd2_2;
	wire w_dff_B_gC1xw0672_2;
	wire w_dff_B_ucxniJKP3_2;
	wire w_dff_B_GvYE6x427_2;
	wire w_dff_B_BdadzOvs7_2;
	wire w_dff_B_UAj1SjrY2_1;
	wire w_dff_B_ZURcfvPQ0_2;
	wire w_dff_B_WkGbWWub4_2;
	wire w_dff_B_eCMV28ii0_2;
	wire w_dff_B_YJh8Mtet8_2;
	wire w_dff_B_1GAI9xrm6_2;
	wire w_dff_B_vAw4yNn23_2;
	wire w_dff_B_Zz6DcGaK2_2;
	wire w_dff_B_fqzJZH849_2;
	wire w_dff_B_kwB6LRBl7_2;
	wire w_dff_B_GQsCX0NR3_2;
	wire w_dff_B_TipRNKVT4_2;
	wire w_dff_B_2gtpBNs35_2;
	wire w_dff_B_Flb76xP35_2;
	wire w_dff_B_d1ssITac7_2;
	wire w_dff_B_SlYxEG5Y8_2;
	wire w_dff_B_FIf92ijf8_2;
	wire w_dff_B_S3uJgSCE1_2;
	wire w_dff_B_zUWqdC8v8_2;
	wire w_dff_B_m2NcjGE91_2;
	wire w_dff_B_oNuiEidf0_1;
	wire w_dff_B_vUihC5lP1_1;
	wire w_dff_B_6ZZjHziA1_2;
	wire w_dff_B_G0LAQaai6_2;
	wire w_dff_B_MHj26KEy0_2;
	wire w_dff_B_PfTNKA7O1_2;
	wire w_dff_B_6n8B0bJc6_2;
	wire w_dff_B_u7Hog3wX1_2;
	wire w_dff_B_KpBUQ8wl7_2;
	wire w_dff_B_46KAuIWD5_2;
	wire w_dff_B_rHoMFQgi8_2;
	wire w_dff_B_2fW30ZPh7_2;
	wire w_dff_B_z83qEetY7_2;
	wire w_dff_B_vZjcRGP98_2;
	wire w_dff_B_9XesZivJ2_2;
	wire w_dff_B_NMAcy3rD7_2;
	wire w_dff_B_qFFFDnug7_2;
	wire w_dff_B_UX6p194Y7_2;
	wire w_dff_B_k6kywRH35_2;
	wire w_dff_B_D0jKwcVk4_2;
	wire w_dff_B_wzsN9kEW7_2;
	wire w_dff_B_8acDGkWu4_2;
	wire w_dff_B_z7WPkZ804_2;
	wire w_dff_B_2ZlohMTO4_2;
	wire w_dff_B_JqcmM7KS0_2;
	wire w_dff_B_vyg3BJSh4_2;
	wire w_dff_B_T23OO0co1_2;
	wire w_dff_B_1Ehd7qne6_2;
	wire w_dff_B_wqOXyipe2_2;
	wire w_dff_B_g2MKs5hz6_2;
	wire w_dff_B_YQ2qn2jF6_2;
	wire w_dff_B_sQN5eiBb7_2;
	wire w_dff_B_ZFtk1Kng5_2;
	wire w_dff_B_fPYMB1gx9_2;
	wire w_dff_B_YkNbzws61_2;
	wire w_dff_B_NZ65v4E38_2;
	wire w_dff_B_KiPv2Y083_2;
	wire w_dff_B_JOlWKl9O1_1;
	wire w_dff_B_XfLYnpdF6_2;
	wire w_dff_B_hcghk9XZ7_2;
	wire w_dff_B_NsWxy5j11_2;
	wire w_dff_B_6f6rUad83_2;
	wire w_dff_B_ZicVVwmB4_2;
	wire w_dff_B_GQ6zQRTI9_2;
	wire w_dff_B_iOcbgWV56_2;
	wire w_dff_B_sSVQtGts7_2;
	wire w_dff_B_sy4tdcVL2_2;
	wire w_dff_B_UeJXBPEt6_2;
	wire w_dff_B_GS14vH2t8_2;
	wire w_dff_B_xNa5kF7g2_2;
	wire w_dff_B_wKKe9xNQ8_2;
	wire w_dff_B_hfWUd8FK7_2;
	wire w_dff_B_3fmDMV6q8_2;
	wire w_dff_B_QZg7MbcJ4_2;
	wire w_dff_B_Fhdnx1eb8_1;
	wire w_dff_B_64BkNosx3_1;
	wire w_dff_B_AFSW1rJM9_2;
	wire w_dff_B_Lt57vjEl0_2;
	wire w_dff_B_snHSZHEI1_2;
	wire w_dff_B_dSD9j1M32_2;
	wire w_dff_B_wVcQnGcO0_2;
	wire w_dff_B_puNNTyc77_2;
	wire w_dff_B_yWjKXj6o8_2;
	wire w_dff_B_KDSMyLue3_2;
	wire w_dff_B_CgYGKt9D4_2;
	wire w_dff_B_zcbSCr4D8_2;
	wire w_dff_B_uJt3UDUC2_2;
	wire w_dff_B_l0mW5TPC9_2;
	wire w_dff_B_WYj5ns8X9_2;
	wire w_dff_B_wvtTIw738_2;
	wire w_dff_B_C1YSRQ7g6_2;
	wire w_dff_B_dHRuiRfN8_2;
	wire w_dff_B_gyIJUMMZ3_2;
	wire w_dff_B_g80eCCPX6_2;
	wire w_dff_B_qG9XMwlv3_2;
	wire w_dff_B_y2pTILfZ0_2;
	wire w_dff_B_3lPSPYKv0_2;
	wire w_dff_B_n7AMVRDS9_2;
	wire w_dff_B_dC3ZPlEE3_2;
	wire w_dff_B_efvfk0rc2_2;
	wire w_dff_B_yAhbeUEa0_2;
	wire w_dff_B_dcLt4VgG0_2;
	wire w_dff_B_A9qn4Qed0_2;
	wire w_dff_B_RapIJeDF9_2;
	wire w_dff_B_P6NmMIMJ3_2;
	wire w_dff_B_DXXp7Pxl5_1;
	wire w_dff_B_nRvwjuUq6_2;
	wire w_dff_B_Y3IwIJ952_2;
	wire w_dff_B_g56VptH23_2;
	wire w_dff_B_F4Zcur6t1_2;
	wire w_dff_B_QpK5AMUf8_2;
	wire w_dff_B_gCNhqQai0_2;
	wire w_dff_B_E5GXKQ5y1_2;
	wire w_dff_B_D4EnDcGT4_2;
	wire w_dff_B_u8dIuvGZ8_2;
	wire w_dff_B_sP4f4yKz7_2;
	wire w_dff_B_SZvkzbvI6_2;
	wire w_dff_B_40f00axQ4_2;
	wire w_dff_B_p0tOgi460_2;
	wire w_dff_B_4yk26g6X3_1;
	wire w_dff_B_J2DV1nKB9_1;
	wire w_dff_B_82hRT4OB5_2;
	wire w_dff_B_23VDLF7L9_2;
	wire w_dff_B_bNQIYJje6_2;
	wire w_dff_B_fO3eHuoT5_2;
	wire w_dff_B_joOBfP5k2_2;
	wire w_dff_B_wexHMndp0_2;
	wire w_dff_B_c4S10mQb8_2;
	wire w_dff_B_QUjYMaiX1_2;
	wire w_dff_B_U4AZ5aEj3_2;
	wire w_dff_B_rVQEiO3x4_2;
	wire w_dff_B_7CGIm1Xs9_2;
	wire w_dff_B_rWU2nklD9_2;
	wire w_dff_B_5hTvil179_2;
	wire w_dff_B_ER393EM95_2;
	wire w_dff_B_4WCWY19K4_2;
	wire w_dff_B_9pndhanH1_2;
	wire w_dff_B_PCUxEJIg2_2;
	wire w_dff_B_LrnxgylS7_2;
	wire w_dff_B_s6zl5eHJ9_2;
	wire w_dff_B_awqix9DE7_2;
	wire w_dff_B_RrL3WYwu1_2;
	wire w_dff_B_HO6FzM4K1_2;
	wire w_dff_B_9nPMHveG8_1;
	wire w_dff_B_XdtLQB7X6_2;
	wire w_dff_B_hwKN7OCW4_2;
	wire w_dff_B_6wYcFkxl1_2;
	wire w_dff_B_eaKJy4xE4_2;
	wire w_dff_B_0fGhoOSl2_2;
	wire w_dff_B_HOwsr0M04_2;
	wire w_dff_B_5KbKsbZn8_2;
	wire w_dff_B_J9IEz1r19_2;
	wire w_dff_B_ADuKv0yc5_2;
	wire w_dff_B_LKBWQccQ1_2;
	wire w_dff_B_3LF1fFik5_2;
	wire w_dff_B_KpCmnpil7_2;
	wire w_dff_B_0koEPZvE1_1;
	wire w_dff_B_mW7jJoG59_1;
	wire w_dff_B_bPZJas5R4_2;
	wire w_dff_B_4fhzi4Bd0_2;
	wire w_dff_B_97e0JX4Y1_2;
	wire w_dff_B_5CtKi17v4_2;
	wire w_dff_B_RHiQYOYh5_2;
	wire w_dff_B_s7rXv6oG9_2;
	wire w_dff_B_1YbWHAfd8_2;
	wire w_dff_B_XpA3bmsu4_2;
	wire w_dff_B_Un1YDpde2_2;
	wire w_dff_B_BXuAESMg7_2;
	wire w_dff_B_IFJ7U6Uv5_2;
	wire w_dff_B_VLnNGJHJ5_2;
	wire w_dff_B_1P3xHSq93_2;
	wire w_dff_B_fp6zLPHS6_2;
	wire w_dff_B_5t0S9Tc66_2;
	wire w_dff_B_ec9y6jOn3_2;
	wire w_dff_B_LvUd9uLj8_1;
	wire w_dff_B_kmHm9Wpt5_2;
	wire w_dff_B_X5V6kJyn2_2;
	wire w_dff_B_i8NYvCSz4_2;
	wire w_dff_B_gZBN4ew09_2;
	wire w_dff_B_sGm4xLkU6_2;
	wire w_dff_B_tYzdjnY44_2;
	wire w_dff_B_DTtGETrj7_2;
	wire w_dff_B_XrMHkfLs9_2;
	wire w_dff_B_1Wo4CiF30_2;
	wire w_dff_B_S5tqoVU85_2;
	wire w_dff_B_5RHH1Fax3_2;
	wire w_dff_B_Br8rk8lT2_2;
	wire w_dff_B_0t79R8j42_2;
	wire w_dff_B_O2P6ExlF7_2;
	wire w_dff_B_SSM5SvsX8_2;
	wire w_dff_B_fdbm5c8k8_2;
	wire w_dff_B_BjhJC7Mp1_2;
	wire w_dff_B_DL47iGsn1_2;
	wire w_dff_B_w74yMYTa7_2;
	wire w_dff_B_h0WeFLoh1_2;
	wire w_dff_B_HQl7EJU00_2;
	wire w_dff_B_cv0a7YUk9_1;
	wire w_dff_B_Gz9mkbZW3_2;
	wire w_dff_B_3j5auCwl7_2;
	wire w_dff_B_pOROb8Pk7_2;
	wire w_dff_B_3R0Sen8r1_2;
	wire w_dff_B_UfCzOdpd3_2;
	wire w_dff_B_ChYkX4iW9_2;
	wire w_dff_B_wCp8FuyK2_2;
	wire w_dff_B_TyAkCYbZ4_2;
	wire w_dff_B_ZorCzA459_2;
	wire w_dff_B_drOzPVID4_2;
	wire w_dff_B_0GefHd6l8_2;
	wire w_dff_B_6JgC3XOe7_2;
	wire w_dff_B_PNRnO2Eg7_2;
	wire w_dff_A_2dt4Jpqk0_0;
	wire w_dff_A_5ImTVvdP6_0;
	wire w_dff_B_cde1KABN0_2;
	wire w_dff_A_9MgiCG545_0;
	wire w_dff_A_jqTD4e0F0_0;
	wire w_dff_A_d5Hs080Z2_0;
	wire w_dff_B_NlKQY1ue6_2;
	wire w_dff_A_G9SnM9lB2_0;
	wire w_dff_A_64J3g8NG2_0;
	wire w_dff_B_ZBbanpTL9_2;
	wire w_dff_B_xjGe0H5j2_2;
	jand g0000(.dina(w_G273gat_7[1]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G290gat_7[2]),.dinb(w_G18gat_7[1]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_n65_0[1]),.dinb(w_G545gat_0),.dout(n66),.clk(gclk));
	jnot g0003(.din(w_n66_0[1]),.dout(n67),.clk(gclk));
	jnot g0004(.din(w_G18gat_7[0]),.dout(n68),.clk(gclk));
	jnot g0005(.din(w_G273gat_7[0]),.dout(n69),.clk(gclk));
	jcb g0006(.dina(w_n69_0[1]),.dinb(n68),.dout(n70));
	jnot g0007(.din(w_n70_0[1]),.dout(n71),.clk(gclk));
	jand g0008(.dina(w_G290gat_7[1]),.dinb(w_G1gat_7[0]),.dout(n72),.clk(gclk));
	jcb g0009(.dina(w_dff_B_44QAozby7_0),.dinb(n71),.dout(n73));
	jand g0010(.dina(w_dff_B_6HCBISXv8_0),.dinb(w_n67_0[1]),.dout(G1581gat),.clk(gclk));
	jand g0011(.dina(w_G307gat_7[1]),.dinb(w_G1gat_6[2]),.dout(n75),.clk(gclk));
	jnot g0012(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G290gat_7[0]),.dout(n78),.clk(gclk));
	jcb g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79));
	jcb g0016(.dina(n79),.dinb(w_n70_0[0]),.dout(n80));
	jand g0017(.dina(w_G273gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jcb g0018(.dina(n81),.dinb(w_n65_0[0]),.dout(n82));
	jand g0019(.dina(n82),.dinb(w_n80_0[2]),.dout(n83),.clk(gclk));
	jxor g0020(.dina(w_n83_0[1]),.dinb(w_n67_0[0]),.dout(n84),.clk(gclk));
	jxor g0021(.dina(w_n84_0[1]),.dinb(w_dff_B_ffyvxpWQ4_1),.dout(G1901gat),.clk(gclk));
	jand g0022(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n86),.clk(gclk));
	jnot g0023(.din(w_n86_0[1]),.dout(n87),.clk(gclk));
	jcb g0024(.dina(w_n83_0[0]),.dinb(w_n66_0[0]),.dout(n88));
	jcb g0025(.dina(w_n84_0[0]),.dinb(w_n75_0[0]),.dout(n89));
	jand g0026(.dina(n89),.dinb(w_dff_B_g0p1OFM37_1),.dout(n90),.clk(gclk));
	jand g0027(.dina(w_G307gat_7[0]),.dinb(w_G18gat_6[2]),.dout(n91),.clk(gclk));
	jnot g0028(.din(w_n91_0[1]),.dout(n92),.clk(gclk));
	jnot g0029(.din(w_n80_0[1]),.dout(n93),.clk(gclk));
	jcb g0030(.dina(w_n69_0[0]),.dinb(w_n77_0[0]),.dout(n94));
	jnot g0031(.din(w_G52gat_7[2]),.dout(n95),.clk(gclk));
	jcb g0032(.dina(w_n78_0[0]),.dinb(n95),.dout(n96));
	jcb g0033(.dina(n96),.dinb(n94),.dout(n97));
	jand g0034(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G273gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jcb g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100));
	jand g0037(.dina(n100),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g0038(.dina(w_n101_0[2]),.dinb(w_n93_0[1]),.dout(n102),.clk(gclk));
	jxor g0039(.dina(n102),.dinb(w_dff_B_sc9KY8Fy9_1),.dout(n103),.clk(gclk));
	jxor g0040(.dina(w_n103_0[1]),.dinb(w_n90_0[1]),.dout(n104),.clk(gclk));
	jxor g0041(.dina(w_n104_0[1]),.dinb(w_dff_B_JZA2Vr1t8_1),.dout(G2223gat),.clk(gclk));
	jand g0042(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n106),.clk(gclk));
	jnot g0043(.din(w_n106_0[1]),.dout(n107),.clk(gclk));
	jnot g0044(.din(w_n103_0[0]),.dout(n108),.clk(gclk));
	jcb g0045(.dina(n108),.dinb(w_n90_0[0]),.dout(n109));
	jcb g0046(.dina(w_n104_0[0]),.dinb(w_n86_0[0]),.dout(n110));
	jand g0047(.dina(n110),.dinb(w_dff_B_z1dMPwYz1_1),.dout(n111),.clk(gclk));
	jand g0048(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n112),.clk(gclk));
	jnot g0049(.din(w_n112_0[1]),.dout(n113),.clk(gclk));
	jcb g0050(.dina(w_n101_0[1]),.dinb(w_n93_0[0]),.dout(n114));
	jxor g0051(.dina(w_n101_0[0]),.dinb(w_n80_0[0]),.dout(n115),.clk(gclk));
	jcb g0052(.dina(n115),.dinb(w_n91_0[0]),.dout(n116));
	jand g0053(.dina(n116),.dinb(w_dff_B_7XBAQlWe7_1),.dout(n117),.clk(gclk));
	jand g0054(.dina(w_G307gat_6[2]),.dinb(w_G35gat_6[2]),.dout(n118),.clk(gclk));
	jnot g0055(.din(n118),.dout(n119),.clk(gclk));
	jnot g0056(.din(w_n97_0[0]),.dout(n120),.clk(gclk));
	jand g0057(.dina(w_G290gat_6[1]),.dinb(w_G69gat_7[1]),.dout(n121),.clk(gclk));
	jand g0058(.dina(w_n121_0[1]),.dinb(w_n99_0[0]),.dout(n122),.clk(gclk));
	jnot g0059(.din(w_n122_0[1]),.dout(n123),.clk(gclk));
	jand g0060(.dina(w_G290gat_6[0]),.dinb(w_G52gat_7[0]),.dout(n124),.clk(gclk));
	jand g0061(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n125),.clk(gclk));
	jcb g0062(.dina(w_n125_0[1]),.dinb(n124),.dout(n126));
	jand g0063(.dina(w_dff_B_KG6L1ole9_0),.dinb(w_n123_0[1]),.dout(n127),.clk(gclk));
	jxor g0064(.dina(w_n127_0[1]),.dinb(w_n120_0[1]),.dout(n128),.clk(gclk));
	jxor g0065(.dina(w_n128_0[1]),.dinb(w_n119_0[1]),.dout(n129),.clk(gclk));
	jnot g0066(.din(w_n129_0[1]),.dout(n130),.clk(gclk));
	jxor g0067(.dina(w_n130_0[1]),.dinb(w_n117_0[2]),.dout(n131),.clk(gclk));
	jxor g0068(.dina(n131),.dinb(w_dff_B_q9owYeI12_1),.dout(n132),.clk(gclk));
	jxor g0069(.dina(w_n132_0[1]),.dinb(w_n111_0[1]),.dout(n133),.clk(gclk));
	jxor g0070(.dina(w_n133_0[1]),.dinb(w_dff_B_6lI0U1M62_1),.dout(G2548gat),.clk(gclk));
	jand g0071(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n135),.clk(gclk));
	jnot g0072(.din(w_n135_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(w_n132_0[0]),.dout(n137),.clk(gclk));
	jcb g0074(.dina(n137),.dinb(w_n111_0[0]),.dout(n138));
	jcb g0075(.dina(w_n133_0[0]),.dinb(w_n106_0[0]),.dout(n139));
	jand g0076(.dina(n139),.dinb(n138),.dout(n140),.clk(gclk));
	jand g0077(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n141),.clk(gclk));
	jnot g0078(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jcb g0079(.dina(w_n130_0[0]),.dinb(w_n117_0[1]),.dout(n143));
	jxor g0080(.dina(w_n129_0[0]),.dinb(w_n117_0[0]),.dout(n144),.clk(gclk));
	jcb g0081(.dina(n144),.dinb(w_n112_0[0]),.dout(n145));
	jand g0082(.dina(n145),.dinb(n143),.dout(n146),.clk(gclk));
	jand g0083(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n147),.clk(gclk));
	jnot g0084(.din(n147),.dout(n148),.clk(gclk));
	jcb g0085(.dina(w_n127_0[0]),.dinb(w_n120_0[0]),.dout(n149));
	jnot g0086(.din(n149),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_n128_0[0]),.dinb(w_n119_0[0]),.dout(n151),.clk(gclk));
	jcb g0088(.dina(n151),.dinb(w_dff_B_JOEeLthO3_1),.dout(n152));
	jand g0089(.dina(w_G307gat_6[1]),.dinb(w_G52gat_6[2]),.dout(n153),.clk(gclk));
	jnot g0090(.din(n153),.dout(n154),.clk(gclk));
	jand g0091(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n155),.clk(gclk));
	jand g0092(.dina(w_n155_0[1]),.dinb(w_n125_0[0]),.dout(n156),.clk(gclk));
	jnot g0093(.din(w_n156_0[1]),.dout(n157),.clk(gclk));
	jand g0094(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n158),.clk(gclk));
	jcb g0095(.dina(w_n158_0[1]),.dinb(w_n121_0[0]),.dout(n159));
	jand g0096(.dina(w_dff_B_7heOTNru1_0),.dinb(w_n157_0[1]),.dout(n160),.clk(gclk));
	jxor g0097(.dina(w_n160_0[1]),.dinb(w_n122_0[0]),.dout(n161),.clk(gclk));
	jxor g0098(.dina(w_n161_0[1]),.dinb(w_n154_0[1]),.dout(n162),.clk(gclk));
	jxor g0099(.dina(w_n162_0[1]),.dinb(w_n152_0[1]),.dout(n163),.clk(gclk));
	jxor g0100(.dina(w_n163_0[1]),.dinb(w_n148_0[1]),.dout(n164),.clk(gclk));
	jnot g0101(.din(w_n164_0[1]),.dout(n165),.clk(gclk));
	jxor g0102(.dina(w_n165_0[1]),.dinb(w_n146_0[2]),.dout(n166),.clk(gclk));
	jxor g0103(.dina(n166),.dinb(w_dff_B_fQZLEDiW3_1),.dout(n167),.clk(gclk));
	jxor g0104(.dina(w_n167_0[1]),.dinb(w_n140_0[1]),.dout(n168),.clk(gclk));
	jxor g0105(.dina(w_n168_0[1]),.dinb(w_dff_B_2NBSrRwF8_1),.dout(G2877gat),.clk(gclk));
	jand g0106(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n170),.clk(gclk));
	jnot g0107(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jnot g0108(.din(w_n167_0[0]),.dout(n172),.clk(gclk));
	jcb g0109(.dina(n172),.dinb(w_n140_0[0]),.dout(n173));
	jcb g0110(.dina(w_n168_0[0]),.dinb(w_n135_0[0]),.dout(n174));
	jand g0111(.dina(n174),.dinb(n173),.dout(n175),.clk(gclk));
	jand g0112(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n176),.clk(gclk));
	jnot g0113(.din(w_n176_0[1]),.dout(n177),.clk(gclk));
	jcb g0114(.dina(w_n165_0[0]),.dinb(w_n146_0[1]),.dout(n178));
	jxor g0115(.dina(w_n164_0[0]),.dinb(w_n146_0[0]),.dout(n179),.clk(gclk));
	jcb g0116(.dina(n179),.dinb(w_n141_0[0]),.dout(n180));
	jand g0117(.dina(n180),.dinb(n178),.dout(n181),.clk(gclk));
	jand g0118(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n182),.clk(gclk));
	jnot g0119(.din(n182),.dout(n183),.clk(gclk));
	jand g0120(.dina(w_n162_0[0]),.dinb(w_n152_0[0]),.dout(n184),.clk(gclk));
	jand g0121(.dina(w_n163_0[0]),.dinb(w_n148_0[0]),.dout(n185),.clk(gclk));
	jcb g0122(.dina(n185),.dinb(w_dff_B_0mJuPkMW1_1),.dout(n186));
	jand g0123(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n187),.clk(gclk));
	jnot g0124(.din(n187),.dout(n188),.clk(gclk));
	jnot g0125(.din(w_n160_0[0]),.dout(n189),.clk(gclk));
	jand g0126(.dina(n189),.dinb(w_n123_0[0]),.dout(n190),.clk(gclk));
	jand g0127(.dina(w_n161_0[0]),.dinb(w_n154_0[0]),.dout(n191),.clk(gclk));
	jcb g0128(.dina(n191),.dinb(n190),.dout(n192));
	jand g0129(.dina(w_G307gat_6[0]),.dinb(w_G69gat_6[2]),.dout(n193),.clk(gclk));
	jnot g0130(.din(n193),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n195),.clk(gclk));
	jand g0132(.dina(w_n195_0[1]),.dinb(w_n158_0[0]),.dout(n196),.clk(gclk));
	jnot g0133(.din(w_n196_0[2]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n198),.clk(gclk));
	jcb g0135(.dina(w_n198_0[1]),.dinb(w_n155_0[0]),.dout(n199));
	jand g0136(.dina(w_dff_B_wD40bFgi9_0),.dinb(n197),.dout(n200),.clk(gclk));
	jxor g0137(.dina(w_n200_0[1]),.dinb(w_n156_0[0]),.dout(n201),.clk(gclk));
	jxor g0138(.dina(w_n201_0[1]),.dinb(w_n194_0[1]),.dout(n202),.clk(gclk));
	jxor g0139(.dina(w_n202_0[1]),.dinb(w_n192_0[1]),.dout(n203),.clk(gclk));
	jxor g0140(.dina(w_n203_0[1]),.dinb(w_n188_0[1]),.dout(n204),.clk(gclk));
	jxor g0141(.dina(w_n204_0[1]),.dinb(w_n186_0[1]),.dout(n205),.clk(gclk));
	jxor g0142(.dina(w_n205_0[1]),.dinb(w_n183_0[1]),.dout(n206),.clk(gclk));
	jnot g0143(.din(w_n206_0[1]),.dout(n207),.clk(gclk));
	jxor g0144(.dina(w_n207_0[1]),.dinb(w_n181_0[2]),.dout(n208),.clk(gclk));
	jxor g0145(.dina(n208),.dinb(w_dff_B_IV2jBIFP1_1),.dout(n209),.clk(gclk));
	jxor g0146(.dina(w_n209_0[1]),.dinb(w_n175_0[1]),.dout(n210),.clk(gclk));
	jxor g0147(.dina(w_n210_0[1]),.dinb(w_dff_B_KLFHqAdj5_1),.dout(G3211gat),.clk(gclk));
	jand g0148(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n212),.clk(gclk));
	jnot g0149(.din(w_n212_0[1]),.dout(n213),.clk(gclk));
	jnot g0150(.din(w_n209_0[0]),.dout(n214),.clk(gclk));
	jcb g0151(.dina(n214),.dinb(w_n175_0[0]),.dout(n215));
	jcb g0152(.dina(w_n210_0[0]),.dinb(w_n170_0[0]),.dout(n216));
	jand g0153(.dina(n216),.dinb(n215),.dout(n217),.clk(gclk));
	jand g0154(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n218),.clk(gclk));
	jnot g0155(.din(w_n218_0[1]),.dout(n219),.clk(gclk));
	jcb g0156(.dina(w_n207_0[0]),.dinb(w_n181_0[1]),.dout(n220));
	jxor g0157(.dina(w_n206_0[0]),.dinb(w_n181_0[0]),.dout(n221),.clk(gclk));
	jcb g0158(.dina(n221),.dinb(w_n176_0[0]),.dout(n222));
	jand g0159(.dina(n222),.dinb(n220),.dout(n223),.clk(gclk));
	jand g0160(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n224),.clk(gclk));
	jnot g0161(.din(n224),.dout(n225),.clk(gclk));
	jand g0162(.dina(w_n204_0[0]),.dinb(w_n186_0[0]),.dout(n226),.clk(gclk));
	jand g0163(.dina(w_n205_0[0]),.dinb(w_n183_0[0]),.dout(n227),.clk(gclk));
	jcb g0164(.dina(n227),.dinb(w_dff_B_EK6M9CMC1_1),.dout(n228));
	jand g0165(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n229),.clk(gclk));
	jnot g0166(.din(n229),.dout(n230),.clk(gclk));
	jand g0167(.dina(w_n202_0[0]),.dinb(w_n192_0[0]),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_n203_0[0]),.dinb(w_n188_0[0]),.dout(n232),.clk(gclk));
	jcb g0169(.dina(n232),.dinb(w_dff_B_H8Nf2bxb9_1),.dout(n233));
	jand g0170(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n234),.clk(gclk));
	jnot g0171(.din(n234),.dout(n235),.clk(gclk));
	jnot g0172(.din(w_n200_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_n157_0[0]),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_n201_0[0]),.dinb(w_n194_0[0]),.dout(n238),.clk(gclk));
	jcb g0175(.dina(n238),.dinb(n237),.dout(n239));
	jand g0176(.dina(w_G307gat_5[2]),.dinb(w_G86gat_6[2]),.dout(n240),.clk(gclk));
	jnot g0177(.din(n240),.dout(n241),.clk(gclk));
	jand g0178(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_n242_0[1]),.dinb(w_n198_0[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(w_n243_0[2]),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n245),.clk(gclk));
	jcb g0182(.dina(w_n245_0[1]),.dinb(w_n195_0[0]),.dout(n246));
	jand g0183(.dina(w_dff_B_VTHvwSX19_0),.dinb(n244),.dout(n247),.clk(gclk));
	jxor g0184(.dina(w_n247_0[1]),.dinb(w_n196_0[1]),.dout(n248),.clk(gclk));
	jxor g0185(.dina(w_n248_0[1]),.dinb(w_n241_0[1]),.dout(n249),.clk(gclk));
	jxor g0186(.dina(w_n249_0[1]),.dinb(w_n239_0[1]),.dout(n250),.clk(gclk));
	jxor g0187(.dina(w_n250_0[1]),.dinb(w_n235_0[1]),.dout(n251),.clk(gclk));
	jxor g0188(.dina(w_n251_0[1]),.dinb(w_n233_0[1]),.dout(n252),.clk(gclk));
	jxor g0189(.dina(w_n252_0[1]),.dinb(w_n230_0[1]),.dout(n253),.clk(gclk));
	jxor g0190(.dina(w_n253_0[1]),.dinb(w_n228_0[1]),.dout(n254),.clk(gclk));
	jxor g0191(.dina(w_n254_0[1]),.dinb(w_n225_0[1]),.dout(n255),.clk(gclk));
	jnot g0192(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jxor g0193(.dina(w_n256_0[1]),.dinb(w_n223_0[2]),.dout(n257),.clk(gclk));
	jxor g0194(.dina(n257),.dinb(w_dff_B_hkBaqYUO0_1),.dout(n258),.clk(gclk));
	jxor g0195(.dina(w_n258_0[1]),.dinb(w_n217_0[1]),.dout(n259),.clk(gclk));
	jxor g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_Fd6u6okS6_1),.dout(G3552gat),.clk(gclk));
	jand g0197(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n261),.clk(gclk));
	jnot g0198(.din(w_n261_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(w_n258_0[0]),.dout(n263),.clk(gclk));
	jcb g0200(.dina(n263),.dinb(w_n217_0[0]),.dout(n264));
	jcb g0201(.dina(w_n259_0[0]),.dinb(w_n212_0[0]),.dout(n265));
	jand g0202(.dina(n265),.dinb(n264),.dout(n266),.clk(gclk));
	jand g0203(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n267),.clk(gclk));
	jnot g0204(.din(w_n267_0[1]),.dout(n268),.clk(gclk));
	jcb g0205(.dina(w_n256_0[0]),.dinb(w_n223_0[1]),.dout(n269));
	jxor g0206(.dina(w_n255_0[0]),.dinb(w_n223_0[0]),.dout(n270),.clk(gclk));
	jcb g0207(.dina(n270),.dinb(w_n218_0[0]),.dout(n271));
	jand g0208(.dina(n271),.dinb(n269),.dout(n272),.clk(gclk));
	jand g0209(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n273),.clk(gclk));
	jnot g0210(.din(n273),.dout(n274),.clk(gclk));
	jand g0211(.dina(w_n253_0[0]),.dinb(w_n228_0[0]),.dout(n275),.clk(gclk));
	jand g0212(.dina(w_n254_0[0]),.dinb(w_n225_0[0]),.dout(n276),.clk(gclk));
	jcb g0213(.dina(n276),.dinb(w_dff_B_179JyEBS4_1),.dout(n277));
	jand g0214(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n278),.clk(gclk));
	jnot g0215(.din(n278),.dout(n279),.clk(gclk));
	jand g0216(.dina(w_n251_0[0]),.dinb(w_n233_0[0]),.dout(n280),.clk(gclk));
	jand g0217(.dina(w_n252_0[0]),.dinb(w_n230_0[0]),.dout(n281),.clk(gclk));
	jcb g0218(.dina(n281),.dinb(w_dff_B_TMXlGXGE2_1),.dout(n282));
	jand g0219(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(n283),.dout(n284),.clk(gclk));
	jand g0221(.dina(w_n249_0[0]),.dinb(w_n239_0[0]),.dout(n285),.clk(gclk));
	jand g0222(.dina(w_n250_0[0]),.dinb(w_n235_0[0]),.dout(n286),.clk(gclk));
	jcb g0223(.dina(n286),.dinb(w_dff_B_Z0Y6Bzw53_1),.dout(n287));
	jand g0224(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n288),.clk(gclk));
	jnot g0225(.din(n288),.dout(n289),.clk(gclk));
	jcb g0226(.dina(w_n247_0[0]),.dinb(w_n196_0[0]),.dout(n290));
	jnot g0227(.din(n290),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n248_0[0]),.dinb(w_n241_0[0]),.dout(n292),.clk(gclk));
	jcb g0229(.dina(n292),.dinb(w_dff_B_7uz8IcC05_1),.dout(n293));
	jand g0230(.dina(w_G307gat_5[1]),.dinb(w_G103gat_6[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n296_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g0234(.din(w_n297_0[2]),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n299),.clk(gclk));
	jcb g0236(.dina(w_n299_0[1]),.dinb(w_n242_0[0]),.dout(n300));
	jand g0237(.dina(w_dff_B_DIG1ikH87_0),.dinb(n298),.dout(n301),.clk(gclk));
	jxor g0238(.dina(w_n301_0[1]),.dinb(w_n243_0[1]),.dout(n302),.clk(gclk));
	jxor g0239(.dina(w_n302_0[1]),.dinb(w_n295_0[1]),.dout(n303),.clk(gclk));
	jxor g0240(.dina(w_n303_0[1]),.dinb(w_n293_0[1]),.dout(n304),.clk(gclk));
	jxor g0241(.dina(w_n304_0[1]),.dinb(w_n289_0[1]),.dout(n305),.clk(gclk));
	jxor g0242(.dina(w_n305_0[1]),.dinb(w_n287_0[1]),.dout(n306),.clk(gclk));
	jxor g0243(.dina(w_n306_0[1]),.dinb(w_n284_0[1]),.dout(n307),.clk(gclk));
	jxor g0244(.dina(w_n307_0[1]),.dinb(w_n282_0[1]),.dout(n308),.clk(gclk));
	jxor g0245(.dina(w_n308_0[1]),.dinb(w_n279_0[1]),.dout(n309),.clk(gclk));
	jxor g0246(.dina(w_n309_0[1]),.dinb(w_n277_0[1]),.dout(n310),.clk(gclk));
	jxor g0247(.dina(w_n310_0[1]),.dinb(w_n274_0[1]),.dout(n311),.clk(gclk));
	jnot g0248(.din(w_n311_0[1]),.dout(n312),.clk(gclk));
	jxor g0249(.dina(w_n312_0[1]),.dinb(w_n272_0[2]),.dout(n313),.clk(gclk));
	jxor g0250(.dina(n313),.dinb(w_dff_B_hp4iNseb0_1),.dout(n314),.clk(gclk));
	jxor g0251(.dina(w_n314_0[1]),.dinb(w_n266_0[1]),.dout(n315),.clk(gclk));
	jxor g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_MoG9tggT5_1),.dout(G3895gat),.clk(gclk));
	jand g0253(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n317),.clk(gclk));
	jnot g0254(.din(w_n317_0[1]),.dout(n318),.clk(gclk));
	jnot g0255(.din(w_n314_0[0]),.dout(n319),.clk(gclk));
	jcb g0256(.dina(n319),.dinb(w_n266_0[0]),.dout(n320));
	jcb g0257(.dina(w_n315_0[0]),.dinb(w_n261_0[0]),.dout(n321));
	jand g0258(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jand g0259(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n323),.clk(gclk));
	jnot g0260(.din(w_n323_0[1]),.dout(n324),.clk(gclk));
	jcb g0261(.dina(w_n312_0[0]),.dinb(w_n272_0[1]),.dout(n325));
	jxor g0262(.dina(w_n311_0[0]),.dinb(w_n272_0[0]),.dout(n326),.clk(gclk));
	jcb g0263(.dina(n326),.dinb(w_n267_0[0]),.dout(n327));
	jand g0264(.dina(n327),.dinb(n325),.dout(n328),.clk(gclk));
	jand g0265(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n329),.clk(gclk));
	jnot g0266(.din(n329),.dout(n330),.clk(gclk));
	jand g0267(.dina(w_n309_0[0]),.dinb(w_n277_0[0]),.dout(n331),.clk(gclk));
	jand g0268(.dina(w_n310_0[0]),.dinb(w_n274_0[0]),.dout(n332),.clk(gclk));
	jcb g0269(.dina(n332),.dinb(w_dff_B_a6aAry2s3_1),.dout(n333));
	jand g0270(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n334),.clk(gclk));
	jnot g0271(.din(n334),.dout(n335),.clk(gclk));
	jand g0272(.dina(w_n307_0[0]),.dinb(w_n282_0[0]),.dout(n336),.clk(gclk));
	jand g0273(.dina(w_n308_0[0]),.dinb(w_n279_0[0]),.dout(n337),.clk(gclk));
	jcb g0274(.dina(n337),.dinb(w_dff_B_TjKIPwAU4_1),.dout(n338));
	jand g0275(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n339),.clk(gclk));
	jnot g0276(.din(n339),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_n305_0[0]),.dinb(w_n287_0[0]),.dout(n341),.clk(gclk));
	jand g0278(.dina(w_n306_0[0]),.dinb(w_n284_0[0]),.dout(n342),.clk(gclk));
	jcb g0279(.dina(n342),.dinb(w_dff_B_OsDt93ur4_1),.dout(n343));
	jand g0280(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n344),.clk(gclk));
	jnot g0281(.din(n344),.dout(n345),.clk(gclk));
	jand g0282(.dina(w_n303_0[0]),.dinb(w_n293_0[0]),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_n304_0[0]),.dinb(w_n289_0[0]),.dout(n347),.clk(gclk));
	jcb g0284(.dina(n347),.dinb(w_dff_B_JkEj9UbZ8_1),.dout(n348));
	jand g0285(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n349),.clk(gclk));
	jnot g0286(.din(n349),.dout(n350),.clk(gclk));
	jcb g0287(.dina(w_n301_0[0]),.dinb(w_n243_0[0]),.dout(n351));
	jnot g0288(.din(n351),.dout(n352),.clk(gclk));
	jand g0289(.dina(w_n302_0[0]),.dinb(w_n295_0[0]),.dout(n353),.clk(gclk));
	jcb g0290(.dina(n353),.dinb(w_dff_B_ZYD8hTSh7_1),.dout(n354));
	jand g0291(.dina(w_G307gat_5[0]),.dinb(w_G120gat_6[2]),.dout(n355),.clk(gclk));
	jnot g0292(.din(n355),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n357),.clk(gclk));
	jand g0294(.dina(w_n357_0[1]),.dinb(w_n299_0[0]),.dout(n358),.clk(gclk));
	jnot g0295(.din(w_n358_0[2]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n360),.clk(gclk));
	jcb g0297(.dina(w_n360_0[1]),.dinb(w_n296_0[0]),.dout(n361));
	jand g0298(.dina(w_dff_B_YuU6LOnn8_0),.dinb(n359),.dout(n362),.clk(gclk));
	jxor g0299(.dina(w_n362_0[1]),.dinb(w_n297_0[1]),.dout(n363),.clk(gclk));
	jxor g0300(.dina(w_n363_0[1]),.dinb(w_n356_0[1]),.dout(n364),.clk(gclk));
	jxor g0301(.dina(w_n364_0[1]),.dinb(w_n354_0[1]),.dout(n365),.clk(gclk));
	jxor g0302(.dina(w_n365_0[1]),.dinb(w_n350_0[1]),.dout(n366),.clk(gclk));
	jxor g0303(.dina(w_n366_0[1]),.dinb(w_n348_0[1]),.dout(n367),.clk(gclk));
	jxor g0304(.dina(w_n367_0[1]),.dinb(w_n345_0[1]),.dout(n368),.clk(gclk));
	jxor g0305(.dina(w_n368_0[1]),.dinb(w_n343_0[1]),.dout(n369),.clk(gclk));
	jxor g0306(.dina(w_n369_0[1]),.dinb(w_n340_0[1]),.dout(n370),.clk(gclk));
	jxor g0307(.dina(w_n370_0[1]),.dinb(w_n338_0[1]),.dout(n371),.clk(gclk));
	jxor g0308(.dina(w_n371_0[1]),.dinb(w_n335_0[1]),.dout(n372),.clk(gclk));
	jxor g0309(.dina(w_n372_0[1]),.dinb(w_n333_0[1]),.dout(n373),.clk(gclk));
	jxor g0310(.dina(w_n373_0[1]),.dinb(w_n330_0[1]),.dout(n374),.clk(gclk));
	jnot g0311(.din(w_n374_0[1]),.dout(n375),.clk(gclk));
	jxor g0312(.dina(w_n375_0[1]),.dinb(w_n328_0[2]),.dout(n376),.clk(gclk));
	jxor g0313(.dina(n376),.dinb(w_dff_B_J2iYhzFI2_1),.dout(n377),.clk(gclk));
	jxor g0314(.dina(w_n377_0[1]),.dinb(w_n322_0[1]),.dout(n378),.clk(gclk));
	jxor g0315(.dina(w_n378_0[1]),.dinb(w_dff_B_Vq2eGezB9_1),.dout(G4241gat),.clk(gclk));
	jand g0316(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n380),.clk(gclk));
	jnot g0317(.din(w_n380_0[1]),.dout(n381),.clk(gclk));
	jnot g0318(.din(w_n377_0[0]),.dout(n382),.clk(gclk));
	jcb g0319(.dina(n382),.dinb(w_n322_0[0]),.dout(n383));
	jcb g0320(.dina(w_n378_0[0]),.dinb(w_n317_0[0]),.dout(n384));
	jand g0321(.dina(n384),.dinb(n383),.dout(n385),.clk(gclk));
	jand g0322(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n386),.clk(gclk));
	jnot g0323(.din(w_n386_0[1]),.dout(n387),.clk(gclk));
	jcb g0324(.dina(w_n375_0[0]),.dinb(w_n328_0[1]),.dout(n388));
	jxor g0325(.dina(w_n374_0[0]),.dinb(w_n328_0[0]),.dout(n389),.clk(gclk));
	jcb g0326(.dina(n389),.dinb(w_n323_0[0]),.dout(n390));
	jand g0327(.dina(n390),.dinb(n388),.dout(n391),.clk(gclk));
	jand g0328(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n392),.clk(gclk));
	jnot g0329(.din(n392),.dout(n393),.clk(gclk));
	jand g0330(.dina(w_n372_0[0]),.dinb(w_n333_0[0]),.dout(n394),.clk(gclk));
	jand g0331(.dina(w_n373_0[0]),.dinb(w_n330_0[0]),.dout(n395),.clk(gclk));
	jcb g0332(.dina(n395),.dinb(w_dff_B_P93Tff5z4_1),.dout(n396));
	jand g0333(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n397),.clk(gclk));
	jnot g0334(.din(n397),.dout(n398),.clk(gclk));
	jand g0335(.dina(w_n370_0[0]),.dinb(w_n338_0[0]),.dout(n399),.clk(gclk));
	jand g0336(.dina(w_n371_0[0]),.dinb(w_n335_0[0]),.dout(n400),.clk(gclk));
	jcb g0337(.dina(n400),.dinb(w_dff_B_YDTgA7rp3_1),.dout(n401));
	jand g0338(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n402),.clk(gclk));
	jnot g0339(.din(n402),.dout(n403),.clk(gclk));
	jand g0340(.dina(w_n368_0[0]),.dinb(w_n343_0[0]),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_n369_0[0]),.dinb(w_n340_0[0]),.dout(n405),.clk(gclk));
	jcb g0342(.dina(n405),.dinb(w_dff_B_4ZkH0V4J4_1),.dout(n406));
	jand g0343(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n407),.clk(gclk));
	jnot g0344(.din(n407),.dout(n408),.clk(gclk));
	jand g0345(.dina(w_n366_0[0]),.dinb(w_n348_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(w_n367_0[0]),.dinb(w_n345_0[0]),.dout(n410),.clk(gclk));
	jcb g0347(.dina(n410),.dinb(w_dff_B_FvN6rCQc2_1),.dout(n411));
	jand g0348(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n412),.clk(gclk));
	jnot g0349(.din(n412),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n364_0[0]),.dinb(w_n354_0[0]),.dout(n414),.clk(gclk));
	jand g0351(.dina(w_n365_0[0]),.dinb(w_n350_0[0]),.dout(n415),.clk(gclk));
	jcb g0352(.dina(n415),.dinb(w_dff_B_aklalK3q6_1),.dout(n416));
	jand g0353(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n417),.clk(gclk));
	jnot g0354(.din(n417),.dout(n418),.clk(gclk));
	jcb g0355(.dina(w_n362_0[0]),.dinb(w_n297_0[0]),.dout(n419));
	jand g0356(.dina(w_n363_0[0]),.dinb(w_n356_0[0]),.dout(n420),.clk(gclk));
	jnot g0357(.din(n420),.dout(n421),.clk(gclk));
	jand g0358(.dina(n421),.dinb(w_dff_B_FriOFbtv9_1),.dout(n422),.clk(gclk));
	jnot g0359(.din(n422),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_G307gat_4[2]),.dinb(w_G137gat_6[2]),.dout(n424),.clk(gclk));
	jnot g0361(.din(n424),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n426),.clk(gclk));
	jand g0363(.dina(w_n426_0[1]),.dinb(w_n360_0[0]),.dout(n427),.clk(gclk));
	jnot g0364(.din(w_n427_0[2]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n429),.clk(gclk));
	jcb g0366(.dina(w_n429_0[1]),.dinb(w_n357_0[0]),.dout(n430));
	jand g0367(.dina(w_dff_B_xsOacfNt7_0),.dinb(n428),.dout(n431),.clk(gclk));
	jxor g0368(.dina(w_n431_0[1]),.dinb(w_n358_0[1]),.dout(n432),.clk(gclk));
	jxor g0369(.dina(w_n432_0[1]),.dinb(w_n425_0[1]),.dout(n433),.clk(gclk));
	jxor g0370(.dina(w_n433_0[1]),.dinb(w_n423_0[1]),.dout(n434),.clk(gclk));
	jxor g0371(.dina(w_n434_0[1]),.dinb(w_n418_0[1]),.dout(n435),.clk(gclk));
	jxor g0372(.dina(w_n435_0[1]),.dinb(w_n416_0[1]),.dout(n436),.clk(gclk));
	jxor g0373(.dina(w_n436_0[1]),.dinb(w_n413_0[1]),.dout(n437),.clk(gclk));
	jxor g0374(.dina(w_n437_0[1]),.dinb(w_n411_0[1]),.dout(n438),.clk(gclk));
	jxor g0375(.dina(w_n438_0[1]),.dinb(w_n408_0[1]),.dout(n439),.clk(gclk));
	jxor g0376(.dina(w_n439_0[1]),.dinb(w_n406_0[1]),.dout(n440),.clk(gclk));
	jxor g0377(.dina(w_n440_0[1]),.dinb(w_n403_0[1]),.dout(n441),.clk(gclk));
	jxor g0378(.dina(w_n441_0[1]),.dinb(w_n401_0[1]),.dout(n442),.clk(gclk));
	jxor g0379(.dina(w_n442_0[1]),.dinb(w_n398_0[1]),.dout(n443),.clk(gclk));
	jxor g0380(.dina(w_n443_0[1]),.dinb(w_n396_0[1]),.dout(n444),.clk(gclk));
	jxor g0381(.dina(w_n444_0[1]),.dinb(w_n393_0[1]),.dout(n445),.clk(gclk));
	jnot g0382(.din(w_n445_0[1]),.dout(n446),.clk(gclk));
	jxor g0383(.dina(w_n446_0[1]),.dinb(w_n391_0[2]),.dout(n447),.clk(gclk));
	jxor g0384(.dina(n447),.dinb(w_dff_B_VJscNDj46_1),.dout(n448),.clk(gclk));
	jxor g0385(.dina(w_n448_0[1]),.dinb(w_n385_0[1]),.dout(n449),.clk(gclk));
	jxor g0386(.dina(w_n449_0[1]),.dinb(w_dff_B_75UviKYP7_1),.dout(G4591gat),.clk(gclk));
	jand g0387(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n451),.clk(gclk));
	jnot g0388(.din(w_n451_0[1]),.dout(n452),.clk(gclk));
	jnot g0389(.din(w_n448_0[0]),.dout(n453),.clk(gclk));
	jcb g0390(.dina(n453),.dinb(w_n385_0[0]),.dout(n454));
	jcb g0391(.dina(w_n449_0[0]),.dinb(w_n380_0[0]),.dout(n455));
	jand g0392(.dina(n455),.dinb(n454),.dout(n456),.clk(gclk));
	jand g0393(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n457),.clk(gclk));
	jnot g0394(.din(w_n457_0[1]),.dout(n458),.clk(gclk));
	jcb g0395(.dina(w_n446_0[0]),.dinb(w_n391_0[1]),.dout(n459));
	jxor g0396(.dina(w_n445_0[0]),.dinb(w_n391_0[0]),.dout(n460),.clk(gclk));
	jcb g0397(.dina(n460),.dinb(w_n386_0[0]),.dout(n461));
	jand g0398(.dina(n461),.dinb(n459),.dout(n462),.clk(gclk));
	jand g0399(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n463),.clk(gclk));
	jnot g0400(.din(n463),.dout(n464),.clk(gclk));
	jand g0401(.dina(w_n443_0[0]),.dinb(w_n396_0[0]),.dout(n465),.clk(gclk));
	jand g0402(.dina(w_n444_0[0]),.dinb(w_n393_0[0]),.dout(n466),.clk(gclk));
	jcb g0403(.dina(n466),.dinb(w_dff_B_JRaUOXWj3_1),.dout(n467));
	jand g0404(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n468),.clk(gclk));
	jnot g0405(.din(n468),.dout(n469),.clk(gclk));
	jand g0406(.dina(w_n441_0[0]),.dinb(w_n401_0[0]),.dout(n470),.clk(gclk));
	jand g0407(.dina(w_n442_0[0]),.dinb(w_n398_0[0]),.dout(n471),.clk(gclk));
	jcb g0408(.dina(n471),.dinb(w_dff_B_zBQXm9a34_1),.dout(n472));
	jand g0409(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n473),.clk(gclk));
	jnot g0410(.din(n473),.dout(n474),.clk(gclk));
	jand g0411(.dina(w_n439_0[0]),.dinb(w_n406_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(w_n440_0[0]),.dinb(w_n403_0[0]),.dout(n476),.clk(gclk));
	jcb g0413(.dina(n476),.dinb(w_dff_B_tc797yZk2_1),.dout(n477));
	jand g0414(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n478),.clk(gclk));
	jnot g0415(.din(n478),.dout(n479),.clk(gclk));
	jand g0416(.dina(w_n437_0[0]),.dinb(w_n411_0[0]),.dout(n480),.clk(gclk));
	jand g0417(.dina(w_n438_0[0]),.dinb(w_n408_0[0]),.dout(n481),.clk(gclk));
	jcb g0418(.dina(n481),.dinb(w_dff_B_t8UKOF9J6_1),.dout(n482));
	jand g0419(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n435_0[0]),.dinb(w_n416_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n436_0[0]),.dinb(w_n413_0[0]),.dout(n486),.clk(gclk));
	jcb g0423(.dina(n486),.dinb(w_dff_B_0ttUigoW2_1),.dout(n487));
	jand g0424(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n433_0[0]),.dinb(w_n423_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n434_0[0]),.dinb(w_n418_0[0]),.dout(n491),.clk(gclk));
	jcb g0428(.dina(n491),.dinb(w_dff_B_i45uaWzw6_1),.dout(n492));
	jand g0429(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jcb g0431(.dina(w_n431_0[0]),.dinb(w_n358_0[0]),.dout(n495));
	jand g0432(.dina(w_n432_0[0]),.dinb(w_n425_0[0]),.dout(n496),.clk(gclk));
	jnot g0433(.din(n496),.dout(n497),.clk(gclk));
	jand g0434(.dina(n497),.dinb(w_dff_B_nZmWx5Sh4_1),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_G307gat_4[1]),.dinb(w_G154gat_6[2]),.dout(n500),.clk(gclk));
	jnot g0437(.din(n500),.dout(n501),.clk(gclk));
	jand g0438(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_n502_0[1]),.dinb(w_n429_0[0]),.dout(n503),.clk(gclk));
	jnot g0440(.din(w_n503_0[2]),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n505),.clk(gclk));
	jcb g0442(.dina(w_n505_0[1]),.dinb(w_n426_0[0]),.dout(n506));
	jand g0443(.dina(w_dff_B_fr6mKTAI4_0),.dinb(n504),.dout(n507),.clk(gclk));
	jxor g0444(.dina(w_n507_0[1]),.dinb(w_n427_0[1]),.dout(n508),.clk(gclk));
	jxor g0445(.dina(w_n508_0[1]),.dinb(w_n501_0[1]),.dout(n509),.clk(gclk));
	jxor g0446(.dina(w_n509_0[1]),.dinb(w_n499_0[1]),.dout(n510),.clk(gclk));
	jxor g0447(.dina(w_n510_0[1]),.dinb(w_n494_0[1]),.dout(n511),.clk(gclk));
	jxor g0448(.dina(w_n511_0[1]),.dinb(w_n492_0[1]),.dout(n512),.clk(gclk));
	jxor g0449(.dina(w_n512_0[1]),.dinb(w_n489_0[1]),.dout(n513),.clk(gclk));
	jxor g0450(.dina(w_n513_0[1]),.dinb(w_n487_0[1]),.dout(n514),.clk(gclk));
	jxor g0451(.dina(w_n514_0[1]),.dinb(w_n484_0[1]),.dout(n515),.clk(gclk));
	jxor g0452(.dina(w_n515_0[1]),.dinb(w_n482_0[1]),.dout(n516),.clk(gclk));
	jxor g0453(.dina(w_n516_0[1]),.dinb(w_n479_0[1]),.dout(n517),.clk(gclk));
	jxor g0454(.dina(w_n517_0[1]),.dinb(w_n477_0[1]),.dout(n518),.clk(gclk));
	jxor g0455(.dina(w_n518_0[1]),.dinb(w_n474_0[1]),.dout(n519),.clk(gclk));
	jxor g0456(.dina(w_n519_0[1]),.dinb(w_n472_0[1]),.dout(n520),.clk(gclk));
	jxor g0457(.dina(w_n520_0[1]),.dinb(w_n469_0[1]),.dout(n521),.clk(gclk));
	jxor g0458(.dina(w_n521_0[1]),.dinb(w_n467_0[1]),.dout(n522),.clk(gclk));
	jxor g0459(.dina(w_n522_0[1]),.dinb(w_n464_0[1]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[1]),.dout(n524),.clk(gclk));
	jxor g0461(.dina(w_n524_0[1]),.dinb(w_n462_0[2]),.dout(n525),.clk(gclk));
	jxor g0462(.dina(n525),.dinb(w_dff_B_ertSK6Qe6_1),.dout(n526),.clk(gclk));
	jxor g0463(.dina(w_n526_0[1]),.dinb(w_n456_0[1]),.dout(n527),.clk(gclk));
	jxor g0464(.dina(w_n527_0[1]),.dinb(w_dff_B_c1zz1fwu5_1),.dout(G4946gat),.clk(gclk));
	jand g0465(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n529),.clk(gclk));
	jnot g0466(.din(w_n529_0[1]),.dout(n530),.clk(gclk));
	jnot g0467(.din(w_n526_0[0]),.dout(n531),.clk(gclk));
	jcb g0468(.dina(n531),.dinb(w_n456_0[0]),.dout(n532));
	jcb g0469(.dina(w_n527_0[0]),.dinb(w_n451_0[0]),.dout(n533));
	jand g0470(.dina(n533),.dinb(n532),.dout(n534),.clk(gclk));
	jand g0471(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n535),.clk(gclk));
	jnot g0472(.din(w_n535_0[1]),.dout(n536),.clk(gclk));
	jcb g0473(.dina(w_n524_0[0]),.dinb(w_n462_0[1]),.dout(n537));
	jxor g0474(.dina(w_n523_0[0]),.dinb(w_n462_0[0]),.dout(n538),.clk(gclk));
	jcb g0475(.dina(n538),.dinb(w_n457_0[0]),.dout(n539));
	jand g0476(.dina(n539),.dinb(n537),.dout(n540),.clk(gclk));
	jand g0477(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n541),.clk(gclk));
	jnot g0478(.din(n541),.dout(n542),.clk(gclk));
	jand g0479(.dina(w_n521_0[0]),.dinb(w_n467_0[0]),.dout(n543),.clk(gclk));
	jand g0480(.dina(w_n522_0[0]),.dinb(w_n464_0[0]),.dout(n544),.clk(gclk));
	jcb g0481(.dina(n544),.dinb(w_dff_B_AYEMt2pb5_1),.dout(n545));
	jand g0482(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n546),.clk(gclk));
	jnot g0483(.din(n546),.dout(n547),.clk(gclk));
	jand g0484(.dina(w_n519_0[0]),.dinb(w_n472_0[0]),.dout(n548),.clk(gclk));
	jand g0485(.dina(w_n520_0[0]),.dinb(w_n469_0[0]),.dout(n549),.clk(gclk));
	jcb g0486(.dina(n549),.dinb(w_dff_B_v8QRd6LZ4_1),.dout(n550));
	jand g0487(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n551),.clk(gclk));
	jnot g0488(.din(n551),.dout(n552),.clk(gclk));
	jand g0489(.dina(w_n517_0[0]),.dinb(w_n477_0[0]),.dout(n553),.clk(gclk));
	jand g0490(.dina(w_n518_0[0]),.dinb(w_n474_0[0]),.dout(n554),.clk(gclk));
	jcb g0491(.dina(n554),.dinb(w_dff_B_2Ytn0KlC5_1),.dout(n555));
	jand g0492(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n556),.clk(gclk));
	jnot g0493(.din(n556),.dout(n557),.clk(gclk));
	jand g0494(.dina(w_n515_0[0]),.dinb(w_n482_0[0]),.dout(n558),.clk(gclk));
	jand g0495(.dina(w_n516_0[0]),.dinb(w_n479_0[0]),.dout(n559),.clk(gclk));
	jcb g0496(.dina(n559),.dinb(w_dff_B_EeRAn82r9_1),.dout(n560));
	jand g0497(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n561),.clk(gclk));
	jnot g0498(.din(n561),.dout(n562),.clk(gclk));
	jand g0499(.dina(w_n513_0[0]),.dinb(w_n487_0[0]),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n514_0[0]),.dinb(w_n484_0[0]),.dout(n564),.clk(gclk));
	jcb g0501(.dina(n564),.dinb(w_dff_B_Y3iWifio0_1),.dout(n565));
	jand g0502(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n566),.clk(gclk));
	jnot g0503(.din(n566),.dout(n567),.clk(gclk));
	jand g0504(.dina(w_n511_0[0]),.dinb(w_n492_0[0]),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n512_0[0]),.dinb(w_n489_0[0]),.dout(n569),.clk(gclk));
	jcb g0506(.dina(n569),.dinb(w_dff_B_vx7Y6eO44_1),.dout(n570));
	jand g0507(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n571),.clk(gclk));
	jnot g0508(.din(n571),.dout(n572),.clk(gclk));
	jand g0509(.dina(w_n509_0[0]),.dinb(w_n499_0[0]),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n510_0[0]),.dinb(w_n494_0[0]),.dout(n574),.clk(gclk));
	jcb g0511(.dina(n574),.dinb(w_dff_B_hJD0JWYq0_1),.dout(n575));
	jand g0512(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n576),.clk(gclk));
	jnot g0513(.din(n576),.dout(n577),.clk(gclk));
	jcb g0514(.dina(w_n507_0[0]),.dinb(w_n427_0[0]),.dout(n578));
	jand g0515(.dina(w_n508_0[0]),.dinb(w_n501_0[0]),.dout(n579),.clk(gclk));
	jnot g0516(.din(n579),.dout(n580),.clk(gclk));
	jand g0517(.dina(n580),.dinb(w_dff_B_VFNjns4h3_1),.dout(n581),.clk(gclk));
	jnot g0518(.din(n581),.dout(n582),.clk(gclk));
	jand g0519(.dina(w_G307gat_4[0]),.dinb(w_G171gat_6[2]),.dout(n583),.clk(gclk));
	jnot g0520(.din(n583),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n585),.clk(gclk));
	jand g0522(.dina(w_n585_0[1]),.dinb(w_n505_0[0]),.dout(n586),.clk(gclk));
	jnot g0523(.din(w_n586_0[2]),.dout(n587),.clk(gclk));
	jand g0524(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n588),.clk(gclk));
	jcb g0525(.dina(w_n588_0[1]),.dinb(w_n502_0[0]),.dout(n589));
	jand g0526(.dina(w_dff_B_Xk0MFmbp8_0),.dinb(n587),.dout(n590),.clk(gclk));
	jxor g0527(.dina(w_n590_0[1]),.dinb(w_n503_0[1]),.dout(n591),.clk(gclk));
	jxor g0528(.dina(w_n591_0[1]),.dinb(w_n584_0[1]),.dout(n592),.clk(gclk));
	jxor g0529(.dina(w_n592_0[1]),.dinb(w_n582_0[1]),.dout(n593),.clk(gclk));
	jxor g0530(.dina(w_n593_0[1]),.dinb(w_n577_0[1]),.dout(n594),.clk(gclk));
	jxor g0531(.dina(w_n594_0[1]),.dinb(w_n575_0[1]),.dout(n595),.clk(gclk));
	jxor g0532(.dina(w_n595_0[1]),.dinb(w_n572_0[1]),.dout(n596),.clk(gclk));
	jxor g0533(.dina(w_n596_0[1]),.dinb(w_n570_0[1]),.dout(n597),.clk(gclk));
	jxor g0534(.dina(w_n597_0[1]),.dinb(w_n567_0[1]),.dout(n598),.clk(gclk));
	jxor g0535(.dina(w_n598_0[1]),.dinb(w_n565_0[1]),.dout(n599),.clk(gclk));
	jxor g0536(.dina(w_n599_0[1]),.dinb(w_n562_0[1]),.dout(n600),.clk(gclk));
	jxor g0537(.dina(w_n600_0[1]),.dinb(w_n560_0[1]),.dout(n601),.clk(gclk));
	jxor g0538(.dina(w_n601_0[1]),.dinb(w_n557_0[1]),.dout(n602),.clk(gclk));
	jxor g0539(.dina(w_n602_0[1]),.dinb(w_n555_0[1]),.dout(n603),.clk(gclk));
	jxor g0540(.dina(w_n603_0[1]),.dinb(w_n552_0[1]),.dout(n604),.clk(gclk));
	jxor g0541(.dina(w_n604_0[1]),.dinb(w_n550_0[1]),.dout(n605),.clk(gclk));
	jxor g0542(.dina(w_n605_0[1]),.dinb(w_n547_0[1]),.dout(n606),.clk(gclk));
	jxor g0543(.dina(w_n606_0[1]),.dinb(w_n545_0[1]),.dout(n607),.clk(gclk));
	jxor g0544(.dina(w_n607_0[1]),.dinb(w_n542_0[1]),.dout(n608),.clk(gclk));
	jnot g0545(.din(w_n608_0[1]),.dout(n609),.clk(gclk));
	jxor g0546(.dina(w_n609_0[1]),.dinb(w_n540_0[2]),.dout(n610),.clk(gclk));
	jxor g0547(.dina(n610),.dinb(w_dff_B_fSWVXiTU0_1),.dout(n611),.clk(gclk));
	jxor g0548(.dina(w_n611_0[1]),.dinb(w_n534_0[1]),.dout(n612),.clk(gclk));
	jxor g0549(.dina(w_n612_0[1]),.dinb(w_dff_B_54U1Ebai6_1),.dout(G5308gat),.clk(gclk));
	jand g0550(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n614),.clk(gclk));
	jnot g0551(.din(w_n614_0[1]),.dout(n615),.clk(gclk));
	jnot g0552(.din(w_n611_0[0]),.dout(n616),.clk(gclk));
	jcb g0553(.dina(n616),.dinb(w_n534_0[0]),.dout(n617));
	jcb g0554(.dina(w_n612_0[0]),.dinb(w_n529_0[0]),.dout(n618));
	jand g0555(.dina(n618),.dinb(n617),.dout(n619),.clk(gclk));
	jand g0556(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n620),.clk(gclk));
	jnot g0557(.din(w_n620_0[1]),.dout(n621),.clk(gclk));
	jcb g0558(.dina(w_n609_0[0]),.dinb(w_n540_0[1]),.dout(n622));
	jxor g0559(.dina(w_n608_0[0]),.dinb(w_n540_0[0]),.dout(n623),.clk(gclk));
	jcb g0560(.dina(n623),.dinb(w_n535_0[0]),.dout(n624));
	jand g0561(.dina(n624),.dinb(n622),.dout(n625),.clk(gclk));
	jand g0562(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n626),.clk(gclk));
	jnot g0563(.din(n626),.dout(n627),.clk(gclk));
	jand g0564(.dina(w_n606_0[0]),.dinb(w_n545_0[0]),.dout(n628),.clk(gclk));
	jand g0565(.dina(w_n607_0[0]),.dinb(w_n542_0[0]),.dout(n629),.clk(gclk));
	jcb g0566(.dina(n629),.dinb(w_dff_B_DGB6GK2U4_1),.dout(n630));
	jand g0567(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n631),.clk(gclk));
	jnot g0568(.din(n631),.dout(n632),.clk(gclk));
	jand g0569(.dina(w_n604_0[0]),.dinb(w_n550_0[0]),.dout(n633),.clk(gclk));
	jand g0570(.dina(w_n605_0[0]),.dinb(w_n547_0[0]),.dout(n634),.clk(gclk));
	jcb g0571(.dina(n634),.dinb(w_dff_B_mvT3gYh79_1),.dout(n635));
	jand g0572(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n636),.clk(gclk));
	jnot g0573(.din(n636),.dout(n637),.clk(gclk));
	jand g0574(.dina(w_n602_0[0]),.dinb(w_n555_0[0]),.dout(n638),.clk(gclk));
	jand g0575(.dina(w_n603_0[0]),.dinb(w_n552_0[0]),.dout(n639),.clk(gclk));
	jcb g0576(.dina(n639),.dinb(w_dff_B_EzN5P6Er8_1),.dout(n640));
	jand g0577(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n641),.clk(gclk));
	jnot g0578(.din(n641),.dout(n642),.clk(gclk));
	jand g0579(.dina(w_n600_0[0]),.dinb(w_n560_0[0]),.dout(n643),.clk(gclk));
	jand g0580(.dina(w_n601_0[0]),.dinb(w_n557_0[0]),.dout(n644),.clk(gclk));
	jcb g0581(.dina(n644),.dinb(w_dff_B_4XFcQDTb2_1),.dout(n645));
	jand g0582(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n646),.clk(gclk));
	jnot g0583(.din(n646),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_n598_0[0]),.dinb(w_n565_0[0]),.dout(n648),.clk(gclk));
	jand g0585(.dina(w_n599_0[0]),.dinb(w_n562_0[0]),.dout(n649),.clk(gclk));
	jcb g0586(.dina(n649),.dinb(w_dff_B_1P0ORXtM0_1),.dout(n650));
	jand g0587(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n651),.clk(gclk));
	jnot g0588(.din(n651),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_n596_0[0]),.dinb(w_n570_0[0]),.dout(n653),.clk(gclk));
	jand g0590(.dina(w_n597_0[0]),.dinb(w_n567_0[0]),.dout(n654),.clk(gclk));
	jcb g0591(.dina(n654),.dinb(w_dff_B_SqHIZXkK4_1),.dout(n655));
	jand g0592(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n656),.clk(gclk));
	jnot g0593(.din(n656),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_n594_0[0]),.dinb(w_n575_0[0]),.dout(n658),.clk(gclk));
	jand g0595(.dina(w_n595_0[0]),.dinb(w_n572_0[0]),.dout(n659),.clk(gclk));
	jcb g0596(.dina(n659),.dinb(w_dff_B_pqEVTRr14_1),.dout(n660));
	jand g0597(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n661),.clk(gclk));
	jnot g0598(.din(n661),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_n592_0[0]),.dinb(w_n582_0[0]),.dout(n663),.clk(gclk));
	jand g0600(.dina(w_n593_0[0]),.dinb(w_n577_0[0]),.dout(n664),.clk(gclk));
	jcb g0601(.dina(n664),.dinb(w_dff_B_WREzFNmg8_1),.dout(n665));
	jand g0602(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n666),.clk(gclk));
	jnot g0603(.din(n666),.dout(n667),.clk(gclk));
	jcb g0604(.dina(w_n590_0[0]),.dinb(w_n503_0[0]),.dout(n668));
	jand g0605(.dina(w_n591_0[0]),.dinb(w_n584_0[0]),.dout(n669),.clk(gclk));
	jnot g0606(.din(n669),.dout(n670),.clk(gclk));
	jand g0607(.dina(n670),.dinb(w_dff_B_Rh8AN04i2_1),.dout(n671),.clk(gclk));
	jnot g0608(.din(n671),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G307gat_3[2]),.dinb(w_G188gat_6[2]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n675_0[1]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jnot g0613(.din(w_n676_0[2]),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n678),.clk(gclk));
	jcb g0615(.dina(w_n678_0[1]),.dinb(w_n585_0[0]),.dout(n679));
	jand g0616(.dina(w_dff_B_wbmtKYiJ5_0),.dinb(n677),.dout(n680),.clk(gclk));
	jxor g0617(.dina(w_n680_0[1]),.dinb(w_n586_0[1]),.dout(n681),.clk(gclk));
	jxor g0618(.dina(w_n681_0[1]),.dinb(w_n674_0[1]),.dout(n682),.clk(gclk));
	jxor g0619(.dina(w_n682_0[1]),.dinb(w_n672_0[1]),.dout(n683),.clk(gclk));
	jxor g0620(.dina(w_n683_0[1]),.dinb(w_n667_0[1]),.dout(n684),.clk(gclk));
	jxor g0621(.dina(w_n684_0[1]),.dinb(w_n665_0[1]),.dout(n685),.clk(gclk));
	jxor g0622(.dina(w_n685_0[1]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jxor g0623(.dina(w_n686_0[1]),.dinb(w_n660_0[1]),.dout(n687),.clk(gclk));
	jxor g0624(.dina(w_n687_0[1]),.dinb(w_n657_0[1]),.dout(n688),.clk(gclk));
	jxor g0625(.dina(w_n688_0[1]),.dinb(w_n655_0[1]),.dout(n689),.clk(gclk));
	jxor g0626(.dina(w_n689_0[1]),.dinb(w_n652_0[1]),.dout(n690),.clk(gclk));
	jxor g0627(.dina(w_n690_0[1]),.dinb(w_n650_0[1]),.dout(n691),.clk(gclk));
	jxor g0628(.dina(w_n691_0[1]),.dinb(w_n647_0[1]),.dout(n692),.clk(gclk));
	jxor g0629(.dina(w_n692_0[1]),.dinb(w_n645_0[1]),.dout(n693),.clk(gclk));
	jxor g0630(.dina(w_n693_0[1]),.dinb(w_n642_0[1]),.dout(n694),.clk(gclk));
	jxor g0631(.dina(w_n694_0[1]),.dinb(w_n640_0[1]),.dout(n695),.clk(gclk));
	jxor g0632(.dina(w_n695_0[1]),.dinb(w_n637_0[1]),.dout(n696),.clk(gclk));
	jxor g0633(.dina(w_n696_0[1]),.dinb(w_n635_0[1]),.dout(n697),.clk(gclk));
	jxor g0634(.dina(w_n697_0[1]),.dinb(w_n632_0[1]),.dout(n698),.clk(gclk));
	jxor g0635(.dina(w_n698_0[1]),.dinb(w_n630_0[1]),.dout(n699),.clk(gclk));
	jxor g0636(.dina(w_n699_0[1]),.dinb(w_n627_0[1]),.dout(n700),.clk(gclk));
	jnot g0637(.din(w_n700_0[1]),.dout(n701),.clk(gclk));
	jxor g0638(.dina(w_n701_0[1]),.dinb(w_n625_0[2]),.dout(n702),.clk(gclk));
	jxor g0639(.dina(n702),.dinb(w_dff_B_b2d0OJvg0_1),.dout(n703),.clk(gclk));
	jxor g0640(.dina(w_n703_0[1]),.dinb(w_n619_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_dff_B_enIigK9G1_1),.dout(G5672gat),.clk(gclk));
	jand g0642(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n706),.clk(gclk));
	jnot g0643(.din(w_n706_0[1]),.dout(n707),.clk(gclk));
	jnot g0644(.din(w_n703_0[0]),.dout(n708),.clk(gclk));
	jcb g0645(.dina(n708),.dinb(w_n619_0[0]),.dout(n709));
	jcb g0646(.dina(w_n704_0[0]),.dinb(w_n614_0[0]),.dout(n710));
	jand g0647(.dina(n710),.dinb(n709),.dout(n711),.clk(gclk));
	jand g0648(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n712),.clk(gclk));
	jnot g0649(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jcb g0650(.dina(w_n701_0[0]),.dinb(w_n625_0[1]),.dout(n714));
	jxor g0651(.dina(w_n700_0[0]),.dinb(w_n625_0[0]),.dout(n715),.clk(gclk));
	jcb g0652(.dina(n715),.dinb(w_n620_0[0]),.dout(n716));
	jand g0653(.dina(n716),.dinb(n714),.dout(n717),.clk(gclk));
	jand g0654(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n718),.clk(gclk));
	jnot g0655(.din(n718),.dout(n719),.clk(gclk));
	jand g0656(.dina(w_n698_0[0]),.dinb(w_n630_0[0]),.dout(n720),.clk(gclk));
	jand g0657(.dina(w_n699_0[0]),.dinb(w_n627_0[0]),.dout(n721),.clk(gclk));
	jcb g0658(.dina(n721),.dinb(w_dff_B_VTnCxu1s2_1),.dout(n722));
	jand g0659(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n723),.clk(gclk));
	jnot g0660(.din(n723),.dout(n724),.clk(gclk));
	jand g0661(.dina(w_n696_0[0]),.dinb(w_n635_0[0]),.dout(n725),.clk(gclk));
	jand g0662(.dina(w_n697_0[0]),.dinb(w_n632_0[0]),.dout(n726),.clk(gclk));
	jcb g0663(.dina(n726),.dinb(w_dff_B_6nBwJ9zZ6_1),.dout(n727));
	jand g0664(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n728),.clk(gclk));
	jnot g0665(.din(n728),.dout(n729),.clk(gclk));
	jand g0666(.dina(w_n694_0[0]),.dinb(w_n640_0[0]),.dout(n730),.clk(gclk));
	jand g0667(.dina(w_n695_0[0]),.dinb(w_n637_0[0]),.dout(n731),.clk(gclk));
	jcb g0668(.dina(n731),.dinb(w_dff_B_kYgnMuZK0_1),.dout(n732));
	jand g0669(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n733),.clk(gclk));
	jnot g0670(.din(n733),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_n692_0[0]),.dinb(w_n645_0[0]),.dout(n735),.clk(gclk));
	jand g0672(.dina(w_n693_0[0]),.dinb(w_n642_0[0]),.dout(n736),.clk(gclk));
	jcb g0673(.dina(n736),.dinb(w_dff_B_LVoVRGms8_1),.dout(n737));
	jand g0674(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n738),.clk(gclk));
	jnot g0675(.din(n738),.dout(n739),.clk(gclk));
	jand g0676(.dina(w_n690_0[0]),.dinb(w_n650_0[0]),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_n691_0[0]),.dinb(w_n647_0[0]),.dout(n741),.clk(gclk));
	jcb g0678(.dina(n741),.dinb(w_dff_B_eQvYoeCl6_1),.dout(n742));
	jand g0679(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n743),.clk(gclk));
	jnot g0680(.din(n743),.dout(n744),.clk(gclk));
	jand g0681(.dina(w_n688_0[0]),.dinb(w_n655_0[0]),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_n689_0[0]),.dinb(w_n652_0[0]),.dout(n746),.clk(gclk));
	jcb g0683(.dina(n746),.dinb(w_dff_B_2a025RzN9_1),.dout(n747));
	jand g0684(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n748),.clk(gclk));
	jnot g0685(.din(n748),.dout(n749),.clk(gclk));
	jand g0686(.dina(w_n686_0[0]),.dinb(w_n660_0[0]),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_n687_0[0]),.dinb(w_n657_0[0]),.dout(n751),.clk(gclk));
	jcb g0688(.dina(n751),.dinb(w_dff_B_yHDS6tVh6_1),.dout(n752));
	jand g0689(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n753),.clk(gclk));
	jnot g0690(.din(n753),.dout(n754),.clk(gclk));
	jand g0691(.dina(w_n684_0[0]),.dinb(w_n665_0[0]),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_n685_0[0]),.dinb(w_n662_0[0]),.dout(n756),.clk(gclk));
	jcb g0693(.dina(n756),.dinb(w_dff_B_rotSg5d82_1),.dout(n757));
	jand g0694(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n758),.clk(gclk));
	jnot g0695(.din(n758),.dout(n759),.clk(gclk));
	jand g0696(.dina(w_n682_0[0]),.dinb(w_n672_0[0]),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_n683_0[0]),.dinb(w_n667_0[0]),.dout(n761),.clk(gclk));
	jcb g0698(.dina(n761),.dinb(w_dff_B_cgMAQ9Lj0_1),.dout(n762));
	jand g0699(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n763),.clk(gclk));
	jnot g0700(.din(n763),.dout(n764),.clk(gclk));
	jcb g0701(.dina(w_n680_0[0]),.dinb(w_n586_0[0]),.dout(n765));
	jand g0702(.dina(w_n681_0[0]),.dinb(w_n674_0[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(n767),.dinb(w_dff_B_n1Y9jby81_1),.dout(n768),.clk(gclk));
	jnot g0705(.din(n768),.dout(n769),.clk(gclk));
	jand g0706(.dina(w_G307gat_3[1]),.dinb(w_G205gat_6[2]),.dout(n770),.clk(gclk));
	jnot g0707(.din(n770),.dout(n771),.clk(gclk));
	jand g0708(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n772_0[1]),.dinb(w_n678_0[0]),.dout(n773),.clk(gclk));
	jnot g0710(.din(w_n773_0[1]),.dout(n774),.clk(gclk));
	jand g0711(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n775),.clk(gclk));
	jcb g0712(.dina(w_n775_0[1]),.dinb(w_n675_0[0]),.dout(n776));
	jand g0713(.dina(w_dff_B_xvpOpkG77_0),.dinb(w_n774_0[1]),.dout(n777),.clk(gclk));
	jxor g0714(.dina(w_n777_0[1]),.dinb(w_n676_0[1]),.dout(n778),.clk(gclk));
	jxor g0715(.dina(w_n778_0[1]),.dinb(w_n771_0[1]),.dout(n779),.clk(gclk));
	jxor g0716(.dina(w_n779_0[1]),.dinb(w_n769_0[1]),.dout(n780),.clk(gclk));
	jxor g0717(.dina(w_n780_0[1]),.dinb(w_n764_0[1]),.dout(n781),.clk(gclk));
	jxor g0718(.dina(w_n781_0[1]),.dinb(w_n762_0[1]),.dout(n782),.clk(gclk));
	jxor g0719(.dina(w_n782_0[1]),.dinb(w_n759_0[1]),.dout(n783),.clk(gclk));
	jxor g0720(.dina(w_n783_0[1]),.dinb(w_n757_0[1]),.dout(n784),.clk(gclk));
	jxor g0721(.dina(w_n784_0[1]),.dinb(w_n754_0[1]),.dout(n785),.clk(gclk));
	jxor g0722(.dina(w_n785_0[1]),.dinb(w_n752_0[1]),.dout(n786),.clk(gclk));
	jxor g0723(.dina(w_n786_0[1]),.dinb(w_n749_0[1]),.dout(n787),.clk(gclk));
	jxor g0724(.dina(w_n787_0[1]),.dinb(w_n747_0[1]),.dout(n788),.clk(gclk));
	jxor g0725(.dina(w_n788_0[1]),.dinb(w_n744_0[1]),.dout(n789),.clk(gclk));
	jxor g0726(.dina(w_n789_0[1]),.dinb(w_n742_0[1]),.dout(n790),.clk(gclk));
	jxor g0727(.dina(w_n790_0[1]),.dinb(w_n739_0[1]),.dout(n791),.clk(gclk));
	jxor g0728(.dina(w_n791_0[1]),.dinb(w_n737_0[1]),.dout(n792),.clk(gclk));
	jxor g0729(.dina(w_n792_0[1]),.dinb(w_n734_0[1]),.dout(n793),.clk(gclk));
	jxor g0730(.dina(w_n793_0[1]),.dinb(w_n732_0[1]),.dout(n794),.clk(gclk));
	jxor g0731(.dina(w_n794_0[1]),.dinb(w_n729_0[1]),.dout(n795),.clk(gclk));
	jxor g0732(.dina(w_n795_0[1]),.dinb(w_n727_0[1]),.dout(n796),.clk(gclk));
	jxor g0733(.dina(w_n796_0[1]),.dinb(w_n724_0[1]),.dout(n797),.clk(gclk));
	jxor g0734(.dina(w_n797_0[1]),.dinb(w_n722_0[1]),.dout(n798),.clk(gclk));
	jxor g0735(.dina(w_n798_0[1]),.dinb(w_n719_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(w_n799_0[1]),.dout(n800),.clk(gclk));
	jxor g0737(.dina(w_n800_0[1]),.dinb(w_n717_0[2]),.dout(n801),.clk(gclk));
	jxor g0738(.dina(n801),.dinb(w_dff_B_Xr8BrdpT9_1),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n711_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_dff_B_hOB0AtOD9_1),.dout(G5971gat),.clk(gclk));
	jand g0741(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n805),.clk(gclk));
	jnot g0742(.din(w_n805_0[1]),.dout(n806),.clk(gclk));
	jnot g0743(.din(w_n802_0[0]),.dout(n807),.clk(gclk));
	jcb g0744(.dina(n807),.dinb(w_n711_0[0]),.dout(n808));
	jcb g0745(.dina(w_n803_0[0]),.dinb(w_n706_0[0]),.dout(n809));
	jand g0746(.dina(n809),.dinb(n808),.dout(n810),.clk(gclk));
	jand g0747(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n811),.clk(gclk));
	jcb g0748(.dina(w_n800_0[0]),.dinb(w_n717_0[1]),.dout(n812));
	jxor g0749(.dina(w_n799_0[0]),.dinb(w_n717_0[0]),.dout(n813),.clk(gclk));
	jcb g0750(.dina(n813),.dinb(w_n712_0[0]),.dout(n814));
	jand g0751(.dina(n814),.dinb(n812),.dout(n815),.clk(gclk));
	jand g0752(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n816),.clk(gclk));
	jnot g0753(.din(w_n816_0[1]),.dout(n817),.clk(gclk));
	jand g0754(.dina(w_n797_0[0]),.dinb(w_n722_0[0]),.dout(n818),.clk(gclk));
	jand g0755(.dina(w_n798_0[0]),.dinb(w_n719_0[0]),.dout(n819),.clk(gclk));
	jcb g0756(.dina(n819),.dinb(w_dff_B_cMTiWGax5_1),.dout(n820));
	jand g0757(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n821),.clk(gclk));
	jnot g0758(.din(n821),.dout(n822),.clk(gclk));
	jand g0759(.dina(w_n795_0[0]),.dinb(w_n727_0[0]),.dout(n823),.clk(gclk));
	jand g0760(.dina(w_n796_0[0]),.dinb(w_n724_0[0]),.dout(n824),.clk(gclk));
	jcb g0761(.dina(n824),.dinb(w_dff_B_WJTzbYWo0_1),.dout(n825));
	jand g0762(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n826),.clk(gclk));
	jnot g0763(.din(n826),.dout(n827),.clk(gclk));
	jand g0764(.dina(w_n793_0[0]),.dinb(w_n732_0[0]),.dout(n828),.clk(gclk));
	jand g0765(.dina(w_n794_0[0]),.dinb(w_n729_0[0]),.dout(n829),.clk(gclk));
	jcb g0766(.dina(n829),.dinb(w_dff_B_iZxUeO794_1),.dout(n830));
	jand g0767(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n831),.clk(gclk));
	jnot g0768(.din(n831),.dout(n832),.clk(gclk));
	jand g0769(.dina(w_n791_0[0]),.dinb(w_n737_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(w_n792_0[0]),.dinb(w_n734_0[0]),.dout(n834),.clk(gclk));
	jcb g0771(.dina(n834),.dinb(w_dff_B_q1b7ahO29_1),.dout(n835));
	jand g0772(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n836),.clk(gclk));
	jnot g0773(.din(n836),.dout(n837),.clk(gclk));
	jand g0774(.dina(w_n789_0[0]),.dinb(w_n742_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(w_n790_0[0]),.dinb(w_n739_0[0]),.dout(n839),.clk(gclk));
	jcb g0776(.dina(n839),.dinb(w_dff_B_MJOCAlLn4_1),.dout(n840));
	jand g0777(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n841),.clk(gclk));
	jnot g0778(.din(n841),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n787_0[0]),.dinb(w_n747_0[0]),.dout(n843),.clk(gclk));
	jand g0780(.dina(w_n788_0[0]),.dinb(w_n744_0[0]),.dout(n844),.clk(gclk));
	jcb g0781(.dina(n844),.dinb(w_dff_B_ve9g9IJh7_1),.dout(n845));
	jand g0782(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n846),.clk(gclk));
	jnot g0783(.din(n846),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n785_0[0]),.dinb(w_n752_0[0]),.dout(n848),.clk(gclk));
	jand g0785(.dina(w_n786_0[0]),.dinb(w_n749_0[0]),.dout(n849),.clk(gclk));
	jcb g0786(.dina(n849),.dinb(w_dff_B_pv43riop8_1),.dout(n850));
	jand g0787(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n851),.clk(gclk));
	jnot g0788(.din(n851),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n783_0[0]),.dinb(w_n757_0[0]),.dout(n853),.clk(gclk));
	jand g0790(.dina(w_n784_0[0]),.dinb(w_n754_0[0]),.dout(n854),.clk(gclk));
	jcb g0791(.dina(n854),.dinb(w_dff_B_KBFvPjWb1_1),.dout(n855));
	jand g0792(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n856),.clk(gclk));
	jnot g0793(.din(n856),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n781_0[0]),.dinb(w_n762_0[0]),.dout(n858),.clk(gclk));
	jand g0795(.dina(w_n782_0[0]),.dinb(w_n759_0[0]),.dout(n859),.clk(gclk));
	jcb g0796(.dina(n859),.dinb(w_dff_B_0ZsMoynN4_1),.dout(n860));
	jand g0797(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n861),.clk(gclk));
	jnot g0798(.din(n861),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n779_0[0]),.dinb(w_n769_0[0]),.dout(n863),.clk(gclk));
	jand g0800(.dina(w_n780_0[0]),.dinb(w_n764_0[0]),.dout(n864),.clk(gclk));
	jcb g0801(.dina(n864),.dinb(w_dff_B_4XuRTRbF5_1),.dout(n865));
	jand g0802(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n866),.clk(gclk));
	jnot g0803(.din(n866),.dout(n867),.clk(gclk));
	jcb g0804(.dina(w_n777_0[0]),.dinb(w_n676_0[0]),.dout(n868));
	jand g0805(.dina(w_n778_0[0]),.dinb(w_n771_0[0]),.dout(n869),.clk(gclk));
	jnot g0806(.din(n869),.dout(n870),.clk(gclk));
	jand g0807(.dina(n870),.dinb(w_dff_B_7msUnWsI5_1),.dout(n871),.clk(gclk));
	jnot g0808(.din(n871),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_G307gat_3[0]),.dinb(w_G222gat_6[2]),.dout(n873),.clk(gclk));
	jnot g0810(.din(n873),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n875),.clk(gclk));
	jxor g0812(.dina(w_n875_0[1]),.dinb(w_n772_0[0]),.dout(n876),.clk(gclk));
	jcb g0813(.dina(n876),.dinb(w_n773_0[0]),.dout(n877));
	jcb g0814(.dina(w_n875_0[0]),.dinb(w_n774_0[0]),.dout(n878));
	jand g0815(.dina(n878),.dinb(w_n877_0[1]),.dout(n879),.clk(gclk));
	jxor g0816(.dina(w_n879_0[1]),.dinb(w_n874_0[1]),.dout(n880),.clk(gclk));
	jxor g0817(.dina(w_n880_0[1]),.dinb(w_n872_0[1]),.dout(n881),.clk(gclk));
	jxor g0818(.dina(w_n881_0[1]),.dinb(w_n867_0[1]),.dout(n882),.clk(gclk));
	jxor g0819(.dina(w_n882_0[1]),.dinb(w_n865_0[1]),.dout(n883),.clk(gclk));
	jxor g0820(.dina(w_n883_0[1]),.dinb(w_n862_0[1]),.dout(n884),.clk(gclk));
	jxor g0821(.dina(w_n884_0[1]),.dinb(w_n860_0[1]),.dout(n885),.clk(gclk));
	jxor g0822(.dina(w_n885_0[1]),.dinb(w_n857_0[1]),.dout(n886),.clk(gclk));
	jxor g0823(.dina(w_n886_0[1]),.dinb(w_n855_0[1]),.dout(n887),.clk(gclk));
	jxor g0824(.dina(w_n887_0[1]),.dinb(w_n852_0[1]),.dout(n888),.clk(gclk));
	jxor g0825(.dina(w_n888_0[1]),.dinb(w_n850_0[1]),.dout(n889),.clk(gclk));
	jxor g0826(.dina(w_n889_0[1]),.dinb(w_n847_0[1]),.dout(n890),.clk(gclk));
	jxor g0827(.dina(w_n890_0[1]),.dinb(w_n845_0[1]),.dout(n891),.clk(gclk));
	jxor g0828(.dina(w_n891_0[1]),.dinb(w_n842_0[1]),.dout(n892),.clk(gclk));
	jxor g0829(.dina(w_n892_0[1]),.dinb(w_n840_0[1]),.dout(n893),.clk(gclk));
	jxor g0830(.dina(w_n893_0[1]),.dinb(w_n837_0[1]),.dout(n894),.clk(gclk));
	jxor g0831(.dina(w_n894_0[1]),.dinb(w_n835_0[1]),.dout(n895),.clk(gclk));
	jxor g0832(.dina(w_n895_0[1]),.dinb(w_n832_0[1]),.dout(n896),.clk(gclk));
	jxor g0833(.dina(w_n896_0[1]),.dinb(w_n830_0[1]),.dout(n897),.clk(gclk));
	jxor g0834(.dina(w_n897_0[1]),.dinb(w_n827_0[1]),.dout(n898),.clk(gclk));
	jxor g0835(.dina(w_n898_0[1]),.dinb(w_n825_0[1]),.dout(n899),.clk(gclk));
	jxor g0836(.dina(w_n899_0[1]),.dinb(w_n822_0[1]),.dout(n900),.clk(gclk));
	jxor g0837(.dina(w_n900_0[2]),.dinb(w_n820_0[2]),.dout(n901),.clk(gclk));
	jxor g0838(.dina(n901),.dinb(w_dff_B_tapHX3J87_1),.dout(n902),.clk(gclk));
	jxor g0839(.dina(w_n902_0[1]),.dinb(w_n815_0[1]),.dout(n903),.clk(gclk));
	jxor g0840(.dina(w_n903_0[1]),.dinb(w_n811_0[1]),.dout(n904),.clk(gclk));
	jxor g0841(.dina(w_n904_0[1]),.dinb(w_n810_0[1]),.dout(n905),.clk(gclk));
	jxor g0842(.dina(w_n905_0[1]),.dinb(w_dff_B_bKVskMcs8_1),.dout(G6123gat),.clk(gclk));
	jnot g0843(.din(w_n904_0[0]),.dout(n907),.clk(gclk));
	jcb g0844(.dina(n907),.dinb(w_n810_0[0]),.dout(n908));
	jcb g0845(.dina(w_n905_0[0]),.dinb(w_n805_0[0]),.dout(n909));
	jand g0846(.dina(n909),.dinb(w_dff_B_Xia3DPRR8_1),.dout(n910),.clk(gclk));
	jand g0847(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n911),.clk(gclk));
	jnot g0848(.din(w_n902_0[0]),.dout(n912),.clk(gclk));
	jcb g0849(.dina(n912),.dinb(w_n815_0[0]),.dout(n913));
	jcb g0850(.dina(w_n903_0[0]),.dinb(w_n811_0[0]),.dout(n914));
	jand g0851(.dina(n914),.dinb(n913),.dout(n915),.clk(gclk));
	jand g0852(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n916),.clk(gclk));
	jand g0853(.dina(w_n900_0[1]),.dinb(w_n820_0[1]),.dout(n917),.clk(gclk));
	jnot g0854(.din(n917),.dout(n918),.clk(gclk));
	jnot g0855(.din(w_n900_0[0]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(n919),.dinb(w_n820_0[0]),.dout(n920),.clk(gclk));
	jcb g0857(.dina(n920),.dinb(w_n816_0[0]),.dout(n921));
	jand g0858(.dina(n921),.dinb(n918),.dout(n922),.clk(gclk));
	jand g0859(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n923),.clk(gclk));
	jnot g0860(.din(n923),.dout(n924),.clk(gclk));
	jand g0861(.dina(w_n898_0[0]),.dinb(w_n825_0[0]),.dout(n925),.clk(gclk));
	jand g0862(.dina(w_n899_0[0]),.dinb(w_n822_0[0]),.dout(n926),.clk(gclk));
	jcb g0863(.dina(n926),.dinb(w_dff_B_8XmM6ZQT5_1),.dout(n927));
	jand g0864(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n928),.clk(gclk));
	jnot g0865(.din(n928),.dout(n929),.clk(gclk));
	jand g0866(.dina(w_n896_0[0]),.dinb(w_n830_0[0]),.dout(n930),.clk(gclk));
	jand g0867(.dina(w_n897_0[0]),.dinb(w_n827_0[0]),.dout(n931),.clk(gclk));
	jcb g0868(.dina(n931),.dinb(w_dff_B_IgYLrSL78_1),.dout(n932));
	jand g0869(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n933),.clk(gclk));
	jnot g0870(.din(n933),.dout(n934),.clk(gclk));
	jand g0871(.dina(w_n894_0[0]),.dinb(w_n835_0[0]),.dout(n935),.clk(gclk));
	jand g0872(.dina(w_n895_0[0]),.dinb(w_n832_0[0]),.dout(n936),.clk(gclk));
	jcb g0873(.dina(n936),.dinb(w_dff_B_FgdnHYwK2_1),.dout(n937));
	jand g0874(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n938),.clk(gclk));
	jnot g0875(.din(n938),.dout(n939),.clk(gclk));
	jand g0876(.dina(w_n892_0[0]),.dinb(w_n840_0[0]),.dout(n940),.clk(gclk));
	jand g0877(.dina(w_n893_0[0]),.dinb(w_n837_0[0]),.dout(n941),.clk(gclk));
	jcb g0878(.dina(n941),.dinb(w_dff_B_UA07Ppi04_1),.dout(n942));
	jand g0879(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n943),.clk(gclk));
	jnot g0880(.din(n943),.dout(n944),.clk(gclk));
	jand g0881(.dina(w_n890_0[0]),.dinb(w_n845_0[0]),.dout(n945),.clk(gclk));
	jand g0882(.dina(w_n891_0[0]),.dinb(w_n842_0[0]),.dout(n946),.clk(gclk));
	jcb g0883(.dina(n946),.dinb(w_dff_B_N1mDFkm30_1),.dout(n947));
	jand g0884(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n948),.clk(gclk));
	jnot g0885(.din(n948),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_n888_0[0]),.dinb(w_n850_0[0]),.dout(n950),.clk(gclk));
	jand g0887(.dina(w_n889_0[0]),.dinb(w_n847_0[0]),.dout(n951),.clk(gclk));
	jcb g0888(.dina(n951),.dinb(w_dff_B_qeTXLU0b4_1),.dout(n952));
	jand g0889(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n953),.clk(gclk));
	jnot g0890(.din(n953),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_n886_0[0]),.dinb(w_n855_0[0]),.dout(n955),.clk(gclk));
	jand g0892(.dina(w_n887_0[0]),.dinb(w_n852_0[0]),.dout(n956),.clk(gclk));
	jcb g0893(.dina(n956),.dinb(w_dff_B_QeeoHfcw0_1),.dout(n957));
	jand g0894(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n958),.clk(gclk));
	jnot g0895(.din(n958),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_n884_0[0]),.dinb(w_n860_0[0]),.dout(n960),.clk(gclk));
	jand g0897(.dina(w_n885_0[0]),.dinb(w_n857_0[0]),.dout(n961),.clk(gclk));
	jcb g0898(.dina(n961),.dinb(w_dff_B_bYy1OwRT1_1),.dout(n962));
	jand g0899(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n963),.clk(gclk));
	jnot g0900(.din(n963),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_n882_0[0]),.dinb(w_n865_0[0]),.dout(n965),.clk(gclk));
	jand g0902(.dina(w_n883_0[0]),.dinb(w_n862_0[0]),.dout(n966),.clk(gclk));
	jcb g0903(.dina(n966),.dinb(w_dff_B_MZbWiYZP4_1),.dout(n967));
	jand g0904(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n968),.clk(gclk));
	jnot g0905(.din(n968),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_n880_0[0]),.dinb(w_n872_0[0]),.dout(n970),.clk(gclk));
	jand g0907(.dina(w_n881_0[0]),.dinb(w_n867_0[0]),.dout(n971),.clk(gclk));
	jcb g0908(.dina(n971),.dinb(w_dff_B_Qy0Xl20H1_1),.dout(n972));
	jand g0909(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n973),.clk(gclk));
	jnot g0910(.din(n973),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_n879_0[0]),.dinb(w_n874_0[0]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(n976),.dinb(w_n877_0[0]),.dout(n977),.clk(gclk));
	jnot g0914(.din(n977),.dout(n978),.clk(gclk));
	jnot g0915(.din(w_n775_0[0]),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n980),.clk(gclk));
	jand g0917(.dina(w_n980_0[1]),.dinb(n979),.dout(n981),.clk(gclk));
	jnot g0918(.din(n981),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_G307gat_2[2]),.dinb(w_G239gat_6[2]),.dout(n983),.clk(gclk));
	jxor g0920(.dina(w_n983_0[1]),.dinb(w_n982_0[1]),.dout(n984),.clk(gclk));
	jxor g0921(.dina(w_n984_0[1]),.dinb(w_n978_0[1]),.dout(n985),.clk(gclk));
	jxor g0922(.dina(w_n985_0[1]),.dinb(w_n974_0[1]),.dout(n986),.clk(gclk));
	jxor g0923(.dina(w_n986_0[1]),.dinb(w_n972_0[1]),.dout(n987),.clk(gclk));
	jxor g0924(.dina(w_n987_0[1]),.dinb(w_n969_0[1]),.dout(n988),.clk(gclk));
	jxor g0925(.dina(w_n988_0[1]),.dinb(w_n967_0[1]),.dout(n989),.clk(gclk));
	jxor g0926(.dina(w_n989_0[1]),.dinb(w_n964_0[1]),.dout(n990),.clk(gclk));
	jxor g0927(.dina(w_n990_0[1]),.dinb(w_n962_0[1]),.dout(n991),.clk(gclk));
	jxor g0928(.dina(w_n991_0[1]),.dinb(w_n959_0[1]),.dout(n992),.clk(gclk));
	jxor g0929(.dina(w_n992_0[1]),.dinb(w_n957_0[1]),.dout(n993),.clk(gclk));
	jxor g0930(.dina(w_n993_0[1]),.dinb(w_n954_0[1]),.dout(n994),.clk(gclk));
	jxor g0931(.dina(w_n994_0[1]),.dinb(w_n952_0[1]),.dout(n995),.clk(gclk));
	jxor g0932(.dina(w_n995_0[1]),.dinb(w_n949_0[1]),.dout(n996),.clk(gclk));
	jxor g0933(.dina(w_n996_0[1]),.dinb(w_n947_0[1]),.dout(n997),.clk(gclk));
	jxor g0934(.dina(w_n997_0[1]),.dinb(w_n944_0[1]),.dout(n998),.clk(gclk));
	jxor g0935(.dina(w_n998_0[1]),.dinb(w_n942_0[1]),.dout(n999),.clk(gclk));
	jxor g0936(.dina(w_n999_0[1]),.dinb(w_n939_0[1]),.dout(n1000),.clk(gclk));
	jxor g0937(.dina(w_n1000_0[1]),.dinb(w_n937_0[1]),.dout(n1001),.clk(gclk));
	jxor g0938(.dina(w_n1001_0[1]),.dinb(w_n934_0[1]),.dout(n1002),.clk(gclk));
	jxor g0939(.dina(w_n1002_0[1]),.dinb(w_n932_0[1]),.dout(n1003),.clk(gclk));
	jxor g0940(.dina(w_n1003_0[1]),.dinb(w_n929_0[1]),.dout(n1004),.clk(gclk));
	jxor g0941(.dina(w_n1004_0[1]),.dinb(w_n927_0[1]),.dout(n1005),.clk(gclk));
	jxor g0942(.dina(w_n1005_0[1]),.dinb(w_n924_0[1]),.dout(n1006),.clk(gclk));
	jxor g0943(.dina(w_n1006_0[1]),.dinb(w_n922_0[1]),.dout(n1007),.clk(gclk));
	jxor g0944(.dina(w_n1007_0[1]),.dinb(w_n916_0[1]),.dout(n1008),.clk(gclk));
	jnot g0945(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n915_0[2]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(n1010),.dinb(w_n911_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n910_0[1]),.dout(G6150gat),.clk(gclk));
	jand g0949(.dina(w_n1011_0[0]),.dinb(w_n910_0[0]),.dout(n1013),.clk(gclk));
	jcb g0950(.dina(w_n1009_0[0]),.dinb(w_n915_0[1]),.dout(n1014));
	jxor g0951(.dina(w_n1008_0[0]),.dinb(w_n915_0[0]),.dout(n1015),.clk(gclk));
	jcb g0952(.dina(n1015),.dinb(w_n911_0[0]),.dout(n1016));
	jand g0953(.dina(n1016),.dinb(n1014),.dout(n1017),.clk(gclk));
	jand g0954(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1018),.clk(gclk));
	jnot g0955(.din(w_n1006_0[0]),.dout(n1019),.clk(gclk));
	jcb g0956(.dina(n1019),.dinb(w_n922_0[0]),.dout(n1020));
	jcb g0957(.dina(w_n1007_0[0]),.dinb(w_n916_0[0]),.dout(n1021));
	jand g0958(.dina(n1021),.dinb(w_dff_B_fLWRSZbu3_1),.dout(n1022),.clk(gclk));
	jand g0959(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1023),.clk(gclk));
	jand g0960(.dina(w_n1004_0[0]),.dinb(w_n927_0[0]),.dout(n1024),.clk(gclk));
	jand g0961(.dina(w_n1005_0[0]),.dinb(w_n924_0[0]),.dout(n1025),.clk(gclk));
	jcb g0962(.dina(n1025),.dinb(w_dff_B_sNTjJaJO2_1),.dout(n1026));
	jand g0963(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1027),.clk(gclk));
	jnot g0964(.din(n1027),.dout(n1028),.clk(gclk));
	jand g0965(.dina(w_n1002_0[0]),.dinb(w_n932_0[0]),.dout(n1029),.clk(gclk));
	jand g0966(.dina(w_n1003_0[0]),.dinb(w_n929_0[0]),.dout(n1030),.clk(gclk));
	jcb g0967(.dina(n1030),.dinb(w_dff_B_Vxbm8uDo5_1),.dout(n1031));
	jand g0968(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1032),.clk(gclk));
	jnot g0969(.din(n1032),.dout(n1033),.clk(gclk));
	jand g0970(.dina(w_n1000_0[0]),.dinb(w_n937_0[0]),.dout(n1034),.clk(gclk));
	jand g0971(.dina(w_n1001_0[0]),.dinb(w_n934_0[0]),.dout(n1035),.clk(gclk));
	jcb g0972(.dina(n1035),.dinb(w_dff_B_ED789YdO5_1),.dout(n1036));
	jand g0973(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1037),.clk(gclk));
	jnot g0974(.din(n1037),.dout(n1038),.clk(gclk));
	jand g0975(.dina(w_n998_0[0]),.dinb(w_n942_0[0]),.dout(n1039),.clk(gclk));
	jand g0976(.dina(w_n999_0[0]),.dinb(w_n939_0[0]),.dout(n1040),.clk(gclk));
	jcb g0977(.dina(n1040),.dinb(w_dff_B_f7L6yJwE3_1),.dout(n1041));
	jand g0978(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1042),.clk(gclk));
	jnot g0979(.din(n1042),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_n996_0[0]),.dinb(w_n947_0[0]),.dout(n1044),.clk(gclk));
	jand g0981(.dina(w_n997_0[0]),.dinb(w_n944_0[0]),.dout(n1045),.clk(gclk));
	jcb g0982(.dina(n1045),.dinb(w_dff_B_MkDHctiK9_1),.dout(n1046));
	jand g0983(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1047),.clk(gclk));
	jnot g0984(.din(n1047),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_n994_0[0]),.dinb(w_n952_0[0]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n995_0[0]),.dinb(w_n949_0[0]),.dout(n1050),.clk(gclk));
	jcb g0987(.dina(n1050),.dinb(w_dff_B_XRr1dIOp7_1),.dout(n1051));
	jand g0988(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1052),.clk(gclk));
	jnot g0989(.din(n1052),.dout(n1053),.clk(gclk));
	jand g0990(.dina(w_n992_0[0]),.dinb(w_n957_0[0]),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n993_0[0]),.dinb(w_n954_0[0]),.dout(n1055),.clk(gclk));
	jcb g0992(.dina(n1055),.dinb(w_dff_B_VVYYVHft7_1),.dout(n1056));
	jand g0993(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1057),.clk(gclk));
	jnot g0994(.din(n1057),.dout(n1058),.clk(gclk));
	jand g0995(.dina(w_n990_0[0]),.dinb(w_n962_0[0]),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n991_0[0]),.dinb(w_n959_0[0]),.dout(n1060),.clk(gclk));
	jcb g0997(.dina(n1060),.dinb(w_dff_B_DrhxwjcS0_1),.dout(n1061));
	jand g0998(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1062),.clk(gclk));
	jnot g0999(.din(n1062),.dout(n1063),.clk(gclk));
	jand g1000(.dina(w_n988_0[0]),.dinb(w_n967_0[0]),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n989_0[0]),.dinb(w_n964_0[0]),.dout(n1065),.clk(gclk));
	jcb g1002(.dina(n1065),.dinb(w_dff_B_ZbX2H2M93_1),.dout(n1066));
	jand g1003(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1067),.clk(gclk));
	jnot g1004(.din(n1067),.dout(n1068),.clk(gclk));
	jand g1005(.dina(w_n986_0[0]),.dinb(w_n972_0[0]),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n987_0[0]),.dinb(w_n969_0[0]),.dout(n1070),.clk(gclk));
	jcb g1007(.dina(n1070),.dinb(w_dff_B_fBGJNpeL5_1),.dout(n1071));
	jand g1008(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1072),.clk(gclk));
	jnot g1009(.din(n1072),.dout(n1073),.clk(gclk));
	jand g1010(.dina(w_n984_0[0]),.dinb(w_n978_0[0]),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n985_0[0]),.dinb(w_n974_0[0]),.dout(n1075),.clk(gclk));
	jcb g1012(.dina(n1075),.dinb(w_dff_B_cv0a7YUk9_1),.dout(n1076));
	jand g1013(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G307gat_2[1]),.dinb(w_G256gat_6[2]),.dout(n1078),.clk(gclk));
	jcb g1015(.dina(w_n983_0[0]),.dinb(w_n982_0[0]),.dout(n1079));
	jand g1016(.dina(n1079),.dinb(w_n980_0[0]),.dout(n1080),.clk(gclk));
	jxor g1017(.dina(w_n1080_0[1]),.dinb(w_n1078_0[1]),.dout(n1081),.clk(gclk));
	jnot g1018(.din(n1081),.dout(n1082),.clk(gclk));
	jxor g1019(.dina(w_n1082_0[1]),.dinb(w_n1077_0[1]),.dout(n1083),.clk(gclk));
	jxor g1020(.dina(w_n1083_0[1]),.dinb(w_n1076_0[1]),.dout(n1084),.clk(gclk));
	jxor g1021(.dina(w_n1084_0[1]),.dinb(w_n1073_0[1]),.dout(n1085),.clk(gclk));
	jxor g1022(.dina(w_n1085_0[1]),.dinb(w_n1071_0[1]),.dout(n1086),.clk(gclk));
	jxor g1023(.dina(w_n1086_0[1]),.dinb(w_n1068_0[1]),.dout(n1087),.clk(gclk));
	jxor g1024(.dina(w_n1087_0[1]),.dinb(w_n1066_0[1]),.dout(n1088),.clk(gclk));
	jxor g1025(.dina(w_n1088_0[1]),.dinb(w_n1063_0[1]),.dout(n1089),.clk(gclk));
	jxor g1026(.dina(w_n1089_0[1]),.dinb(w_n1061_0[1]),.dout(n1090),.clk(gclk));
	jxor g1027(.dina(w_n1090_0[1]),.dinb(w_n1058_0[1]),.dout(n1091),.clk(gclk));
	jxor g1028(.dina(w_n1091_0[1]),.dinb(w_n1056_0[1]),.dout(n1092),.clk(gclk));
	jxor g1029(.dina(w_n1092_0[1]),.dinb(w_n1053_0[1]),.dout(n1093),.clk(gclk));
	jxor g1030(.dina(w_n1093_0[1]),.dinb(w_n1051_0[1]),.dout(n1094),.clk(gclk));
	jxor g1031(.dina(w_n1094_0[1]),.dinb(w_n1048_0[1]),.dout(n1095),.clk(gclk));
	jxor g1032(.dina(w_n1095_0[1]),.dinb(w_n1046_0[1]),.dout(n1096),.clk(gclk));
	jxor g1033(.dina(w_n1096_0[1]),.dinb(w_n1043_0[1]),.dout(n1097),.clk(gclk));
	jxor g1034(.dina(w_n1097_0[1]),.dinb(w_n1041_0[1]),.dout(n1098),.clk(gclk));
	jxor g1035(.dina(w_n1098_0[1]),.dinb(w_n1038_0[1]),.dout(n1099),.clk(gclk));
	jxor g1036(.dina(w_n1099_0[1]),.dinb(w_n1036_0[1]),.dout(n1100),.clk(gclk));
	jxor g1037(.dina(w_n1100_0[1]),.dinb(w_n1033_0[1]),.dout(n1101),.clk(gclk));
	jxor g1038(.dina(w_n1101_0[1]),.dinb(w_n1031_0[1]),.dout(n1102),.clk(gclk));
	jxor g1039(.dina(w_n1102_0[1]),.dinb(w_n1028_0[1]),.dout(n1103),.clk(gclk));
	jxor g1040(.dina(w_n1103_0[1]),.dinb(w_n1026_0[1]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(n1104),.dout(n1105),.clk(gclk));
	jxor g1042(.dina(w_n1105_0[1]),.dinb(w_n1023_0[1]),.dout(n1106),.clk(gclk));
	jxor g1043(.dina(w_n1106_0[1]),.dinb(w_n1022_0[1]),.dout(n1107),.clk(gclk));
	jxor g1044(.dina(w_n1107_0[1]),.dinb(w_n1018_0[1]),.dout(n1108),.clk(gclk));
	jxor g1045(.dina(w_n1108_0[1]),.dinb(w_n1017_0[1]),.dout(n1109),.clk(gclk));
	jnot g1046(.din(w_n1109_0[1]),.dout(n1110),.clk(gclk));
	jxor g1047(.dina(n1110),.dinb(w_n1013_0[1]),.dout(G6160gat),.clk(gclk));
	jnot g1048(.din(w_n1108_0[0]),.dout(n1112),.clk(gclk));
	jcb g1049(.dina(n1112),.dinb(w_n1017_0[0]),.dout(n1113));
	jcb g1050(.dina(w_n1109_0[0]),.dinb(w_n1013_0[0]),.dout(n1114));
	jand g1051(.dina(n1114),.dinb(w_dff_B_8GXt3znx8_1),.dout(n1115),.clk(gclk));
	jnot g1052(.din(w_n1106_0[0]),.dout(n1116),.clk(gclk));
	jcb g1053(.dina(n1116),.dinb(w_n1022_0[0]),.dout(n1117));
	jcb g1054(.dina(w_n1107_0[0]),.dinb(w_n1018_0[0]),.dout(n1118));
	jand g1055(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g1056(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1120),.clk(gclk));
	jand g1057(.dina(w_n1103_0[0]),.dinb(w_n1026_0[0]),.dout(n1121),.clk(gclk));
	jnot g1058(.din(n1121),.dout(n1122),.clk(gclk));
	jcb g1059(.dina(w_n1105_0[0]),.dinb(w_n1023_0[0]),.dout(n1123));
	jand g1060(.dina(n1123),.dinb(n1122),.dout(n1124),.clk(gclk));
	jand g1061(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1125),.clk(gclk));
	jnot g1062(.din(n1125),.dout(n1126),.clk(gclk));
	jand g1063(.dina(w_n1101_0[0]),.dinb(w_n1031_0[0]),.dout(n1127),.clk(gclk));
	jand g1064(.dina(w_n1102_0[0]),.dinb(w_n1028_0[0]),.dout(n1128),.clk(gclk));
	jcb g1065(.dina(n1128),.dinb(w_dff_B_fZLq7QUg3_1),.dout(n1129));
	jand g1066(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1130),.clk(gclk));
	jnot g1067(.din(n1130),.dout(n1131),.clk(gclk));
	jand g1068(.dina(w_n1099_0[0]),.dinb(w_n1036_0[0]),.dout(n1132),.clk(gclk));
	jand g1069(.dina(w_n1100_0[0]),.dinb(w_n1033_0[0]),.dout(n1133),.clk(gclk));
	jcb g1070(.dina(n1133),.dinb(w_dff_B_ygGrrKsO1_1),.dout(n1134));
	jand g1071(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1135),.clk(gclk));
	jnot g1072(.din(n1135),.dout(n1136),.clk(gclk));
	jand g1073(.dina(w_n1097_0[0]),.dinb(w_n1041_0[0]),.dout(n1137),.clk(gclk));
	jand g1074(.dina(w_n1098_0[0]),.dinb(w_n1038_0[0]),.dout(n1138),.clk(gclk));
	jcb g1075(.dina(n1138),.dinb(w_dff_B_Mufn57ny6_1),.dout(n1139));
	jand g1076(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1140),.clk(gclk));
	jnot g1077(.din(n1140),.dout(n1141),.clk(gclk));
	jand g1078(.dina(w_n1095_0[0]),.dinb(w_n1046_0[0]),.dout(n1142),.clk(gclk));
	jand g1079(.dina(w_n1096_0[0]),.dinb(w_n1043_0[0]),.dout(n1143),.clk(gclk));
	jcb g1080(.dina(n1143),.dinb(w_dff_B_PyIWdvaA6_1),.dout(n1144));
	jand g1081(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1145),.clk(gclk));
	jnot g1082(.din(n1145),.dout(n1146),.clk(gclk));
	jand g1083(.dina(w_n1093_0[0]),.dinb(w_n1051_0[0]),.dout(n1147),.clk(gclk));
	jand g1084(.dina(w_n1094_0[0]),.dinb(w_n1048_0[0]),.dout(n1148),.clk(gclk));
	jcb g1085(.dina(n1148),.dinb(w_dff_B_byEMZ9rd5_1),.dout(n1149));
	jand g1086(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1150),.clk(gclk));
	jnot g1087(.din(n1150),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_n1091_0[0]),.dinb(w_n1056_0[0]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1092_0[0]),.dinb(w_n1053_0[0]),.dout(n1153),.clk(gclk));
	jcb g1090(.dina(n1153),.dinb(w_dff_B_qXyM7Qwc6_1),.dout(n1154));
	jand g1091(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1155),.clk(gclk));
	jnot g1092(.din(n1155),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_n1089_0[0]),.dinb(w_n1061_0[0]),.dout(n1157),.clk(gclk));
	jand g1094(.dina(w_n1090_0[0]),.dinb(w_n1058_0[0]),.dout(n1158),.clk(gclk));
	jcb g1095(.dina(n1158),.dinb(w_dff_B_QsGqq5Sx7_1),.dout(n1159));
	jand g1096(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1160),.clk(gclk));
	jnot g1097(.din(n1160),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_n1087_0[0]),.dinb(w_n1066_0[0]),.dout(n1162),.clk(gclk));
	jand g1099(.dina(w_n1088_0[0]),.dinb(w_n1063_0[0]),.dout(n1163),.clk(gclk));
	jcb g1100(.dina(n1163),.dinb(w_dff_B_jDExplnb2_1),.dout(n1164));
	jand g1101(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1165),.clk(gclk));
	jnot g1102(.din(n1165),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_n1085_0[0]),.dinb(w_n1071_0[0]),.dout(n1167),.clk(gclk));
	jand g1104(.dina(w_n1086_0[0]),.dinb(w_n1068_0[0]),.dout(n1168),.clk(gclk));
	jcb g1105(.dina(n1168),.dinb(w_dff_B_GZxrntJy9_1),.dout(n1169));
	jand g1106(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1170),.clk(gclk));
	jnot g1107(.din(n1170),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_n1083_0[0]),.dinb(w_n1076_0[0]),.dout(n1172),.clk(gclk));
	jand g1109(.dina(w_n1084_0[0]),.dinb(w_n1073_0[0]),.dout(n1173),.clk(gclk));
	jcb g1110(.dina(n1173),.dinb(w_dff_B_LvUd9uLj8_1),.dout(n1174));
	jand g1111(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1175),.clk(gclk));
	jand g1112(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1176),.clk(gclk));
	jcb g1113(.dina(w_n1080_0[0]),.dinb(w_n1078_0[0]),.dout(n1177));
	jcb g1114(.dina(w_n1082_0[0]),.dinb(w_n1077_0[0]),.dout(n1178));
	jand g1115(.dina(n1178),.dinb(w_dff_B_mW7jJoG59_1),.dout(n1179),.clk(gclk));
	jxor g1116(.dina(w_n1179_0[1]),.dinb(w_n1176_0[1]),.dout(n1180),.clk(gclk));
	jnot g1117(.din(n1180),.dout(n1181),.clk(gclk));
	jxor g1118(.dina(w_n1181_0[1]),.dinb(w_n1175_0[1]),.dout(n1182),.clk(gclk));
	jxor g1119(.dina(w_n1182_0[1]),.dinb(w_n1174_0[1]),.dout(n1183),.clk(gclk));
	jxor g1120(.dina(w_n1183_0[1]),.dinb(w_n1171_0[1]),.dout(n1184),.clk(gclk));
	jxor g1121(.dina(w_n1184_0[1]),.dinb(w_n1169_0[1]),.dout(n1185),.clk(gclk));
	jxor g1122(.dina(w_n1185_0[1]),.dinb(w_n1166_0[1]),.dout(n1186),.clk(gclk));
	jxor g1123(.dina(w_n1186_0[1]),.dinb(w_n1164_0[1]),.dout(n1187),.clk(gclk));
	jxor g1124(.dina(w_n1187_0[1]),.dinb(w_n1161_0[1]),.dout(n1188),.clk(gclk));
	jxor g1125(.dina(w_n1188_0[1]),.dinb(w_n1159_0[1]),.dout(n1189),.clk(gclk));
	jxor g1126(.dina(w_n1189_0[1]),.dinb(w_n1156_0[1]),.dout(n1190),.clk(gclk));
	jxor g1127(.dina(w_n1190_0[1]),.dinb(w_n1154_0[1]),.dout(n1191),.clk(gclk));
	jxor g1128(.dina(w_n1191_0[1]),.dinb(w_n1151_0[1]),.dout(n1192),.clk(gclk));
	jxor g1129(.dina(w_n1192_0[1]),.dinb(w_n1149_0[1]),.dout(n1193),.clk(gclk));
	jxor g1130(.dina(w_n1193_0[1]),.dinb(w_n1146_0[1]),.dout(n1194),.clk(gclk));
	jxor g1131(.dina(w_n1194_0[1]),.dinb(w_n1144_0[1]),.dout(n1195),.clk(gclk));
	jxor g1132(.dina(w_n1195_0[1]),.dinb(w_n1141_0[1]),.dout(n1196),.clk(gclk));
	jxor g1133(.dina(w_n1196_0[1]),.dinb(w_n1139_0[1]),.dout(n1197),.clk(gclk));
	jxor g1134(.dina(w_n1197_0[1]),.dinb(w_n1136_0[1]),.dout(n1198),.clk(gclk));
	jxor g1135(.dina(w_n1198_0[1]),.dinb(w_n1134_0[1]),.dout(n1199),.clk(gclk));
	jxor g1136(.dina(w_n1199_0[1]),.dinb(w_n1131_0[1]),.dout(n1200),.clk(gclk));
	jxor g1137(.dina(w_n1200_0[1]),.dinb(w_n1129_0[1]),.dout(n1201),.clk(gclk));
	jxor g1138(.dina(w_n1201_0[1]),.dinb(w_n1126_0[1]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jxor g1140(.dina(w_n1203_0[1]),.dinb(w_n1124_0[1]),.dout(n1204),.clk(gclk));
	jnot g1141(.din(n1204),.dout(n1205),.clk(gclk));
	jxor g1142(.dina(w_n1205_0[1]),.dinb(w_n1120_0[1]),.dout(n1206),.clk(gclk));
	jxor g1143(.dina(w_n1206_0[1]),.dinb(w_n1119_0[1]),.dout(n1207),.clk(gclk));
	jnot g1144(.din(w_n1207_0[1]),.dout(n1208),.clk(gclk));
	jxor g1145(.dina(n1208),.dinb(w_n1115_0[1]),.dout(G6170gat),.clk(gclk));
	jnot g1146(.din(w_n1206_0[0]),.dout(n1210),.clk(gclk));
	jcb g1147(.dina(n1210),.dinb(w_n1119_0[0]),.dout(n1211));
	jcb g1148(.dina(w_n1207_0[0]),.dinb(w_n1115_0[0]),.dout(n1212));
	jand g1149(.dina(n1212),.dinb(w_dff_B_NpeQjmGC5_1),.dout(n1213),.clk(gclk));
	jcb g1150(.dina(w_n1203_0[0]),.dinb(w_n1124_0[0]),.dout(n1214));
	jcb g1151(.dina(w_n1205_0[0]),.dinb(w_n1120_0[0]),.dout(n1215));
	jand g1152(.dina(n1215),.dinb(w_dff_B_CryD6Cfq3_1),.dout(n1216),.clk(gclk));
	jand g1153(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1217),.clk(gclk));
	jand g1154(.dina(w_n1200_0[0]),.dinb(w_n1129_0[0]),.dout(n1218),.clk(gclk));
	jand g1155(.dina(w_n1201_0[0]),.dinb(w_n1126_0[0]),.dout(n1219),.clk(gclk));
	jcb g1156(.dina(n1219),.dinb(w_dff_B_yr9X1Uji1_1),.dout(n1220));
	jand g1157(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1221),.clk(gclk));
	jnot g1158(.din(n1221),.dout(n1222),.clk(gclk));
	jand g1159(.dina(w_n1198_0[0]),.dinb(w_n1134_0[0]),.dout(n1223),.clk(gclk));
	jand g1160(.dina(w_n1199_0[0]),.dinb(w_n1131_0[0]),.dout(n1224),.clk(gclk));
	jcb g1161(.dina(n1224),.dinb(w_dff_B_QxnkdtK96_1),.dout(n1225));
	jand g1162(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1226),.clk(gclk));
	jnot g1163(.din(n1226),.dout(n1227),.clk(gclk));
	jand g1164(.dina(w_n1196_0[0]),.dinb(w_n1139_0[0]),.dout(n1228),.clk(gclk));
	jand g1165(.dina(w_n1197_0[0]),.dinb(w_n1136_0[0]),.dout(n1229),.clk(gclk));
	jcb g1166(.dina(n1229),.dinb(w_dff_B_Bd7910S22_1),.dout(n1230));
	jand g1167(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1231),.clk(gclk));
	jnot g1168(.din(n1231),.dout(n1232),.clk(gclk));
	jand g1169(.dina(w_n1194_0[0]),.dinb(w_n1144_0[0]),.dout(n1233),.clk(gclk));
	jand g1170(.dina(w_n1195_0[0]),.dinb(w_n1141_0[0]),.dout(n1234),.clk(gclk));
	jcb g1171(.dina(n1234),.dinb(w_dff_B_9QvM6iid7_1),.dout(n1235));
	jand g1172(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1236),.clk(gclk));
	jnot g1173(.din(n1236),.dout(n1237),.clk(gclk));
	jand g1174(.dina(w_n1192_0[0]),.dinb(w_n1149_0[0]),.dout(n1238),.clk(gclk));
	jand g1175(.dina(w_n1193_0[0]),.dinb(w_n1146_0[0]),.dout(n1239),.clk(gclk));
	jcb g1176(.dina(n1239),.dinb(w_dff_B_Q4Onb2760_1),.dout(n1240));
	jand g1177(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1241),.clk(gclk));
	jnot g1178(.din(n1241),.dout(n1242),.clk(gclk));
	jand g1179(.dina(w_n1190_0[0]),.dinb(w_n1154_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(w_n1191_0[0]),.dinb(w_n1151_0[0]),.dout(n1244),.clk(gclk));
	jcb g1181(.dina(n1244),.dinb(w_dff_B_7NXe1aam5_1),.dout(n1245));
	jand g1182(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1246),.clk(gclk));
	jnot g1183(.din(n1246),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_n1188_0[0]),.dinb(w_n1159_0[0]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1189_0[0]),.dinb(w_n1156_0[0]),.dout(n1249),.clk(gclk));
	jcb g1186(.dina(n1249),.dinb(w_dff_B_Q47A3wZg4_1),.dout(n1250));
	jand g1187(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1251),.clk(gclk));
	jnot g1188(.din(n1251),.dout(n1252),.clk(gclk));
	jand g1189(.dina(w_n1186_0[0]),.dinb(w_n1164_0[0]),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1187_0[0]),.dinb(w_n1161_0[0]),.dout(n1254),.clk(gclk));
	jcb g1191(.dina(n1254),.dinb(w_dff_B_AvhsdWwx0_1),.dout(n1255));
	jand g1192(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1256),.clk(gclk));
	jnot g1193(.din(n1256),.dout(n1257),.clk(gclk));
	jand g1194(.dina(w_n1184_0[0]),.dinb(w_n1169_0[0]),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1185_0[0]),.dinb(w_n1166_0[0]),.dout(n1259),.clk(gclk));
	jcb g1196(.dina(n1259),.dinb(w_dff_B_rX2mSMAu1_1),.dout(n1260));
	jand g1197(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1261),.clk(gclk));
	jnot g1198(.din(n1261),.dout(n1262),.clk(gclk));
	jand g1199(.dina(w_n1182_0[0]),.dinb(w_n1174_0[0]),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1183_0[0]),.dinb(w_n1171_0[0]),.dout(n1264),.clk(gclk));
	jcb g1201(.dina(n1264),.dinb(w_dff_B_9nPMHveG8_1),.dout(n1265));
	jand g1202(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1267),.clk(gclk));
	jcb g1204(.dina(w_n1179_0[0]),.dinb(w_n1176_0[0]),.dout(n1268));
	jcb g1205(.dina(w_n1181_0[0]),.dinb(w_n1175_0[0]),.dout(n1269));
	jand g1206(.dina(n1269),.dinb(w_dff_B_J2DV1nKB9_1),.dout(n1270),.clk(gclk));
	jxor g1207(.dina(w_n1270_0[1]),.dinb(w_n1267_0[1]),.dout(n1271),.clk(gclk));
	jnot g1208(.din(n1271),.dout(n1272),.clk(gclk));
	jxor g1209(.dina(w_n1272_0[1]),.dinb(w_n1266_0[1]),.dout(n1273),.clk(gclk));
	jxor g1210(.dina(w_n1273_0[1]),.dinb(w_n1265_0[1]),.dout(n1274),.clk(gclk));
	jxor g1211(.dina(w_n1274_0[1]),.dinb(w_n1262_0[1]),.dout(n1275),.clk(gclk));
	jxor g1212(.dina(w_n1275_0[1]),.dinb(w_n1260_0[1]),.dout(n1276),.clk(gclk));
	jxor g1213(.dina(w_n1276_0[1]),.dinb(w_n1257_0[1]),.dout(n1277),.clk(gclk));
	jxor g1214(.dina(w_n1277_0[1]),.dinb(w_n1255_0[1]),.dout(n1278),.clk(gclk));
	jxor g1215(.dina(w_n1278_0[1]),.dinb(w_n1252_0[1]),.dout(n1279),.clk(gclk));
	jxor g1216(.dina(w_n1279_0[1]),.dinb(w_n1250_0[1]),.dout(n1280),.clk(gclk));
	jxor g1217(.dina(w_n1280_0[1]),.dinb(w_n1247_0[1]),.dout(n1281),.clk(gclk));
	jxor g1218(.dina(w_n1281_0[1]),.dinb(w_n1245_0[1]),.dout(n1282),.clk(gclk));
	jxor g1219(.dina(w_n1282_0[1]),.dinb(w_n1242_0[1]),.dout(n1283),.clk(gclk));
	jxor g1220(.dina(w_n1283_0[1]),.dinb(w_n1240_0[1]),.dout(n1284),.clk(gclk));
	jxor g1221(.dina(w_n1284_0[1]),.dinb(w_n1237_0[1]),.dout(n1285),.clk(gclk));
	jxor g1222(.dina(w_n1285_0[1]),.dinb(w_n1235_0[1]),.dout(n1286),.clk(gclk));
	jxor g1223(.dina(w_n1286_0[1]),.dinb(w_n1232_0[1]),.dout(n1287),.clk(gclk));
	jxor g1224(.dina(w_n1287_0[1]),.dinb(w_n1230_0[1]),.dout(n1288),.clk(gclk));
	jxor g1225(.dina(w_n1288_0[1]),.dinb(w_n1227_0[1]),.dout(n1289),.clk(gclk));
	jxor g1226(.dina(w_n1289_0[1]),.dinb(w_n1225_0[1]),.dout(n1290),.clk(gclk));
	jxor g1227(.dina(w_n1290_0[1]),.dinb(w_n1222_0[1]),.dout(n1291),.clk(gclk));
	jxor g1228(.dina(w_n1291_0[1]),.dinb(w_n1220_0[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jxor g1230(.dina(w_n1293_0[1]),.dinb(w_n1217_0[1]),.dout(n1294),.clk(gclk));
	jxor g1231(.dina(w_n1294_0[1]),.dinb(w_n1216_0[1]),.dout(n1295),.clk(gclk));
	jnot g1232(.din(w_n1295_0[1]),.dout(n1296),.clk(gclk));
	jxor g1233(.dina(w_dff_B_pI24JtGM4_0),.dinb(w_n1213_0[1]),.dout(G6180gat),.clk(gclk));
	jnot g1234(.din(w_n1294_0[0]),.dout(n1298),.clk(gclk));
	jcb g1235(.dina(n1298),.dinb(w_n1216_0[0]),.dout(n1299));
	jcb g1236(.dina(w_n1295_0[0]),.dinb(w_n1213_0[0]),.dout(n1300));
	jand g1237(.dina(n1300),.dinb(w_dff_B_n6bnUqnb4_1),.dout(n1301),.clk(gclk));
	jnot g1238(.din(w_n1220_0[0]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(w_n1291_0[0]),.dout(n1303),.clk(gclk));
	jcb g1240(.dina(n1303),.dinb(n1302),.dout(n1304));
	jcb g1241(.dina(w_n1293_0[0]),.dinb(w_n1217_0[0]),.dout(n1305));
	jand g1242(.dina(n1305),.dinb(w_dff_B_fmTukOSK5_1),.dout(n1306),.clk(gclk));
	jand g1243(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1307),.clk(gclk));
	jand g1244(.dina(w_n1289_0[0]),.dinb(w_n1225_0[0]),.dout(n1308),.clk(gclk));
	jand g1245(.dina(w_n1290_0[0]),.dinb(w_n1222_0[0]),.dout(n1309),.clk(gclk));
	jcb g1246(.dina(n1309),.dinb(w_dff_B_v3VgPoVA6_1),.dout(n1310));
	jand g1247(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1311),.clk(gclk));
	jnot g1248(.din(n1311),.dout(n1312),.clk(gclk));
	jand g1249(.dina(w_n1287_0[0]),.dinb(w_n1230_0[0]),.dout(n1313),.clk(gclk));
	jand g1250(.dina(w_n1288_0[0]),.dinb(w_n1227_0[0]),.dout(n1314),.clk(gclk));
	jcb g1251(.dina(n1314),.dinb(w_dff_B_RaRq5BB64_1),.dout(n1315));
	jand g1252(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1316),.clk(gclk));
	jnot g1253(.din(n1316),.dout(n1317),.clk(gclk));
	jand g1254(.dina(w_n1285_0[0]),.dinb(w_n1235_0[0]),.dout(n1318),.clk(gclk));
	jand g1255(.dina(w_n1286_0[0]),.dinb(w_n1232_0[0]),.dout(n1319),.clk(gclk));
	jcb g1256(.dina(n1319),.dinb(w_dff_B_tZqSwIO23_1),.dout(n1320));
	jand g1257(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1321),.clk(gclk));
	jnot g1258(.din(n1321),.dout(n1322),.clk(gclk));
	jand g1259(.dina(w_n1283_0[0]),.dinb(w_n1240_0[0]),.dout(n1323),.clk(gclk));
	jand g1260(.dina(w_n1284_0[0]),.dinb(w_n1237_0[0]),.dout(n1324),.clk(gclk));
	jcb g1261(.dina(n1324),.dinb(w_dff_B_32Ixfw7Z1_1),.dout(n1325));
	jand g1262(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(n1326),.dout(n1327),.clk(gclk));
	jand g1264(.dina(w_n1281_0[0]),.dinb(w_n1245_0[0]),.dout(n1328),.clk(gclk));
	jand g1265(.dina(w_n1282_0[0]),.dinb(w_n1242_0[0]),.dout(n1329),.clk(gclk));
	jcb g1266(.dina(n1329),.dinb(w_dff_B_u4aSQSdF1_1),.dout(n1330));
	jand g1267(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1331),.clk(gclk));
	jnot g1268(.din(n1331),.dout(n1332),.clk(gclk));
	jand g1269(.dina(w_n1279_0[0]),.dinb(w_n1250_0[0]),.dout(n1333),.clk(gclk));
	jand g1270(.dina(w_n1280_0[0]),.dinb(w_n1247_0[0]),.dout(n1334),.clk(gclk));
	jcb g1271(.dina(n1334),.dinb(w_dff_B_SblAxLOd8_1),.dout(n1335));
	jand g1272(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1336),.clk(gclk));
	jnot g1273(.din(n1336),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_n1277_0[0]),.dinb(w_n1255_0[0]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1278_0[0]),.dinb(w_n1252_0[0]),.dout(n1339),.clk(gclk));
	jcb g1276(.dina(n1339),.dinb(w_dff_B_jbWyQ2f59_1),.dout(n1340));
	jand g1277(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1341),.clk(gclk));
	jnot g1278(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1279(.dina(w_n1275_0[0]),.dinb(w_n1260_0[0]),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1276_0[0]),.dinb(w_n1257_0[0]),.dout(n1344),.clk(gclk));
	jcb g1281(.dina(n1344),.dinb(w_dff_B_13lUOBpt4_1),.dout(n1345));
	jand g1282(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1346),.clk(gclk));
	jnot g1283(.din(n1346),.dout(n1347),.clk(gclk));
	jand g1284(.dina(w_n1273_0[0]),.dinb(w_n1265_0[0]),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1274_0[0]),.dinb(w_n1262_0[0]),.dout(n1349),.clk(gclk));
	jcb g1286(.dina(n1349),.dinb(w_dff_B_DXXp7Pxl5_1),.dout(n1350));
	jand g1287(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1352),.clk(gclk));
	jcb g1289(.dina(w_n1270_0[0]),.dinb(w_n1267_0[0]),.dout(n1353));
	jcb g1290(.dina(w_n1272_0[0]),.dinb(w_n1266_0[0]),.dout(n1354));
	jand g1291(.dina(n1354),.dinb(w_dff_B_64BkNosx3_1),.dout(n1355),.clk(gclk));
	jxor g1292(.dina(w_n1355_0[1]),.dinb(w_n1352_0[1]),.dout(n1356),.clk(gclk));
	jnot g1293(.din(n1356),.dout(n1357),.clk(gclk));
	jxor g1294(.dina(w_n1357_0[1]),.dinb(w_n1351_0[1]),.dout(n1358),.clk(gclk));
	jxor g1295(.dina(w_n1358_0[1]),.dinb(w_n1350_0[1]),.dout(n1359),.clk(gclk));
	jxor g1296(.dina(w_n1359_0[1]),.dinb(w_n1347_0[1]),.dout(n1360),.clk(gclk));
	jxor g1297(.dina(w_n1360_0[1]),.dinb(w_n1345_0[1]),.dout(n1361),.clk(gclk));
	jxor g1298(.dina(w_n1361_0[1]),.dinb(w_n1342_0[1]),.dout(n1362),.clk(gclk));
	jxor g1299(.dina(w_n1362_0[1]),.dinb(w_n1340_0[1]),.dout(n1363),.clk(gclk));
	jxor g1300(.dina(w_n1363_0[1]),.dinb(w_n1337_0[1]),.dout(n1364),.clk(gclk));
	jxor g1301(.dina(w_n1364_0[1]),.dinb(w_n1335_0[1]),.dout(n1365),.clk(gclk));
	jxor g1302(.dina(w_n1365_0[1]),.dinb(w_n1332_0[1]),.dout(n1366),.clk(gclk));
	jxor g1303(.dina(w_n1366_0[1]),.dinb(w_n1330_0[1]),.dout(n1367),.clk(gclk));
	jxor g1304(.dina(w_n1367_0[1]),.dinb(w_n1327_0[1]),.dout(n1368),.clk(gclk));
	jxor g1305(.dina(w_n1368_0[1]),.dinb(w_n1325_0[1]),.dout(n1369),.clk(gclk));
	jxor g1306(.dina(w_n1369_0[1]),.dinb(w_n1322_0[1]),.dout(n1370),.clk(gclk));
	jxor g1307(.dina(w_n1370_0[1]),.dinb(w_n1320_0[1]),.dout(n1371),.clk(gclk));
	jxor g1308(.dina(w_n1371_0[1]),.dinb(w_n1317_0[1]),.dout(n1372),.clk(gclk));
	jxor g1309(.dina(w_n1372_0[1]),.dinb(w_n1315_0[1]),.dout(n1373),.clk(gclk));
	jxor g1310(.dina(w_n1373_0[1]),.dinb(w_n1312_0[1]),.dout(n1374),.clk(gclk));
	jxor g1311(.dina(w_n1374_0[1]),.dinb(w_n1310_0[1]),.dout(n1375),.clk(gclk));
	jnot g1312(.din(n1375),.dout(n1376),.clk(gclk));
	jxor g1313(.dina(w_n1376_0[1]),.dinb(w_n1307_0[1]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jxor g1315(.dina(w_n1378_0[1]),.dinb(w_n1306_0[1]),.dout(n1379),.clk(gclk));
	jxor g1316(.dina(w_n1379_0[1]),.dinb(w_n1301_0[1]),.dout(G6190gat),.clk(gclk));
	jcb g1317(.dina(w_n1378_0[0]),.dinb(w_n1306_0[0]),.dout(n1381));
	jnot g1318(.din(w_n1379_0[0]),.dout(n1382),.clk(gclk));
	jcb g1319(.dina(w_dff_B_w2l7Nkfj6_0),.dinb(w_n1301_0[0]),.dout(n1383));
	jand g1320(.dina(n1383),.dinb(w_dff_B_NAMTOoqD0_1),.dout(n1384),.clk(gclk));
	jnot g1321(.din(w_n1310_0[0]),.dout(n1385),.clk(gclk));
	jnot g1322(.din(w_n1374_0[0]),.dout(n1386),.clk(gclk));
	jcb g1323(.dina(n1386),.dinb(n1385),.dout(n1387));
	jcb g1324(.dina(w_n1376_0[0]),.dinb(w_n1307_0[0]),.dout(n1388));
	jand g1325(.dina(n1388),.dinb(w_dff_B_pruoaOri4_1),.dout(n1389),.clk(gclk));
	jand g1326(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1390),.clk(gclk));
	jand g1327(.dina(w_n1372_0[0]),.dinb(w_n1315_0[0]),.dout(n1391),.clk(gclk));
	jand g1328(.dina(w_n1373_0[0]),.dinb(w_n1312_0[0]),.dout(n1392),.clk(gclk));
	jcb g1329(.dina(n1392),.dinb(w_dff_B_7bDJzS977_1),.dout(n1393));
	jand g1330(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1394),.clk(gclk));
	jnot g1331(.din(n1394),.dout(n1395),.clk(gclk));
	jand g1332(.dina(w_n1370_0[0]),.dinb(w_n1320_0[0]),.dout(n1396),.clk(gclk));
	jand g1333(.dina(w_n1371_0[0]),.dinb(w_n1317_0[0]),.dout(n1397),.clk(gclk));
	jcb g1334(.dina(n1397),.dinb(w_dff_B_bBMX1SXG4_1),.dout(n1398));
	jand g1335(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1399),.clk(gclk));
	jnot g1336(.din(n1399),.dout(n1400),.clk(gclk));
	jand g1337(.dina(w_n1368_0[0]),.dinb(w_n1325_0[0]),.dout(n1401),.clk(gclk));
	jand g1338(.dina(w_n1369_0[0]),.dinb(w_n1322_0[0]),.dout(n1402),.clk(gclk));
	jcb g1339(.dina(n1402),.dinb(w_dff_B_tnlqCwf56_1),.dout(n1403));
	jand g1340(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1404),.clk(gclk));
	jnot g1341(.din(n1404),.dout(n1405),.clk(gclk));
	jand g1342(.dina(w_n1366_0[0]),.dinb(w_n1330_0[0]),.dout(n1406),.clk(gclk));
	jand g1343(.dina(w_n1367_0[0]),.dinb(w_n1327_0[0]),.dout(n1407),.clk(gclk));
	jcb g1344(.dina(n1407),.dinb(w_dff_B_iLDdWkPX6_1),.dout(n1408));
	jand g1345(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1409),.clk(gclk));
	jnot g1346(.din(n1409),.dout(n1410),.clk(gclk));
	jand g1347(.dina(w_n1364_0[0]),.dinb(w_n1335_0[0]),.dout(n1411),.clk(gclk));
	jand g1348(.dina(w_n1365_0[0]),.dinb(w_n1332_0[0]),.dout(n1412),.clk(gclk));
	jcb g1349(.dina(n1412),.dinb(w_dff_B_TLtisFvc9_1),.dout(n1413));
	jand g1350(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1414),.clk(gclk));
	jnot g1351(.din(n1414),.dout(n1415),.clk(gclk));
	jand g1352(.dina(w_n1362_0[0]),.dinb(w_n1340_0[0]),.dout(n1416),.clk(gclk));
	jand g1353(.dina(w_n1363_0[0]),.dinb(w_n1337_0[0]),.dout(n1417),.clk(gclk));
	jcb g1354(.dina(n1417),.dinb(w_dff_B_gUK6quCH9_1),.dout(n1418));
	jand g1355(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1419),.clk(gclk));
	jnot g1356(.din(n1419),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_n1360_0[0]),.dinb(w_n1345_0[0]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1361_0[0]),.dinb(w_n1342_0[0]),.dout(n1422),.clk(gclk));
	jcb g1359(.dina(n1422),.dinb(w_dff_B_TabAGmhm9_1),.dout(n1423));
	jand g1360(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1424),.clk(gclk));
	jnot g1361(.din(n1424),.dout(n1425),.clk(gclk));
	jand g1362(.dina(w_n1358_0[0]),.dinb(w_n1350_0[0]),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1359_0[0]),.dinb(w_n1347_0[0]),.dout(n1427),.clk(gclk));
	jcb g1364(.dina(n1427),.dinb(w_dff_B_JOlWKl9O1_1),.dout(n1428));
	jand g1365(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1430),.clk(gclk));
	jcb g1367(.dina(w_n1355_0[0]),.dinb(w_n1352_0[0]),.dout(n1431));
	jcb g1368(.dina(w_n1357_0[0]),.dinb(w_n1351_0[0]),.dout(n1432));
	jand g1369(.dina(n1432),.dinb(w_dff_B_vUihC5lP1_1),.dout(n1433),.clk(gclk));
	jxor g1370(.dina(w_n1433_0[1]),.dinb(w_n1430_0[1]),.dout(n1434),.clk(gclk));
	jnot g1371(.din(n1434),.dout(n1435),.clk(gclk));
	jxor g1372(.dina(w_n1435_0[1]),.dinb(w_n1429_0[1]),.dout(n1436),.clk(gclk));
	jxor g1373(.dina(w_n1436_0[1]),.dinb(w_n1428_0[1]),.dout(n1437),.clk(gclk));
	jxor g1374(.dina(w_n1437_0[1]),.dinb(w_n1425_0[1]),.dout(n1438),.clk(gclk));
	jxor g1375(.dina(w_n1438_0[1]),.dinb(w_n1423_0[1]),.dout(n1439),.clk(gclk));
	jxor g1376(.dina(w_n1439_0[1]),.dinb(w_n1420_0[1]),.dout(n1440),.clk(gclk));
	jxor g1377(.dina(w_n1440_0[1]),.dinb(w_n1418_0[1]),.dout(n1441),.clk(gclk));
	jxor g1378(.dina(w_n1441_0[1]),.dinb(w_n1415_0[1]),.dout(n1442),.clk(gclk));
	jxor g1379(.dina(w_n1442_0[1]),.dinb(w_n1413_0[1]),.dout(n1443),.clk(gclk));
	jxor g1380(.dina(w_n1443_0[1]),.dinb(w_n1410_0[1]),.dout(n1444),.clk(gclk));
	jxor g1381(.dina(w_n1444_0[1]),.dinb(w_n1408_0[1]),.dout(n1445),.clk(gclk));
	jxor g1382(.dina(w_n1445_0[1]),.dinb(w_n1405_0[1]),.dout(n1446),.clk(gclk));
	jxor g1383(.dina(w_n1446_0[1]),.dinb(w_n1403_0[1]),.dout(n1447),.clk(gclk));
	jxor g1384(.dina(w_n1447_0[1]),.dinb(w_n1400_0[1]),.dout(n1448),.clk(gclk));
	jxor g1385(.dina(w_n1448_0[1]),.dinb(w_n1398_0[1]),.dout(n1449),.clk(gclk));
	jxor g1386(.dina(w_n1449_0[1]),.dinb(w_n1395_0[1]),.dout(n1450),.clk(gclk));
	jxor g1387(.dina(w_n1450_0[1]),.dinb(w_n1393_0[1]),.dout(n1451),.clk(gclk));
	jnot g1388(.din(n1451),.dout(n1452),.clk(gclk));
	jxor g1389(.dina(w_n1452_0[1]),.dinb(w_n1390_0[1]),.dout(n1453),.clk(gclk));
	jnot g1390(.din(n1453),.dout(n1454),.clk(gclk));
	jxor g1391(.dina(w_n1454_0[1]),.dinb(w_n1389_0[1]),.dout(n1455),.clk(gclk));
	jxor g1392(.dina(w_n1455_0[1]),.dinb(w_n1384_0[1]),.dout(G6200gat),.clk(gclk));
	jcb g1393(.dina(w_n1454_0[0]),.dinb(w_n1389_0[0]),.dout(n1457));
	jnot g1394(.din(w_n1455_0[0]),.dout(n1458),.clk(gclk));
	jcb g1395(.dina(w_dff_B_UJiY7Bnj3_0),.dinb(w_n1384_0[0]),.dout(n1459));
	jand g1396(.dina(n1459),.dinb(w_dff_B_zEQtFjHc9_1),.dout(n1460),.clk(gclk));
	jnot g1397(.din(w_n1393_0[0]),.dout(n1461),.clk(gclk));
	jnot g1398(.din(w_n1450_0[0]),.dout(n1462),.clk(gclk));
	jcb g1399(.dina(n1462),.dinb(w_dff_B_wYs9wv6H6_1),.dout(n1463));
	jcb g1400(.dina(w_n1452_0[0]),.dinb(w_n1390_0[0]),.dout(n1464));
	jand g1401(.dina(n1464),.dinb(w_dff_B_GKM8K4XL9_1),.dout(n1465),.clk(gclk));
	jand g1402(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1466),.clk(gclk));
	jand g1403(.dina(w_n1448_0[0]),.dinb(w_n1398_0[0]),.dout(n1467),.clk(gclk));
	jand g1404(.dina(w_n1449_0[0]),.dinb(w_n1395_0[0]),.dout(n1468),.clk(gclk));
	jcb g1405(.dina(n1468),.dinb(w_dff_B_JxXpUVSx0_1),.dout(n1469));
	jand g1406(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1470),.clk(gclk));
	jnot g1407(.din(n1470),.dout(n1471),.clk(gclk));
	jand g1408(.dina(w_n1446_0[0]),.dinb(w_n1403_0[0]),.dout(n1472),.clk(gclk));
	jand g1409(.dina(w_n1447_0[0]),.dinb(w_n1400_0[0]),.dout(n1473),.clk(gclk));
	jcb g1410(.dina(n1473),.dinb(w_dff_B_vbv4jbug2_1),.dout(n1474));
	jand g1411(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1475),.clk(gclk));
	jnot g1412(.din(n1475),.dout(n1476),.clk(gclk));
	jand g1413(.dina(w_n1444_0[0]),.dinb(w_n1408_0[0]),.dout(n1477),.clk(gclk));
	jand g1414(.dina(w_n1445_0[0]),.dinb(w_n1405_0[0]),.dout(n1478),.clk(gclk));
	jcb g1415(.dina(n1478),.dinb(w_dff_B_2vYE8m0s1_1),.dout(n1479));
	jand g1416(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1480),.clk(gclk));
	jnot g1417(.din(n1480),.dout(n1481),.clk(gclk));
	jand g1418(.dina(w_n1442_0[0]),.dinb(w_n1413_0[0]),.dout(n1482),.clk(gclk));
	jand g1419(.dina(w_n1443_0[0]),.dinb(w_n1410_0[0]),.dout(n1483),.clk(gclk));
	jcb g1420(.dina(n1483),.dinb(w_dff_B_RIrmifht4_1),.dout(n1484));
	jand g1421(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1485),.clk(gclk));
	jnot g1422(.din(n1485),.dout(n1486),.clk(gclk));
	jand g1423(.dina(w_n1440_0[0]),.dinb(w_n1418_0[0]),.dout(n1487),.clk(gclk));
	jand g1424(.dina(w_n1441_0[0]),.dinb(w_n1415_0[0]),.dout(n1488),.clk(gclk));
	jcb g1425(.dina(n1488),.dinb(w_dff_B_SqZb0rTo9_1),.dout(n1489));
	jand g1426(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1490),.clk(gclk));
	jnot g1427(.din(n1490),.dout(n1491),.clk(gclk));
	jand g1428(.dina(w_n1438_0[0]),.dinb(w_n1423_0[0]),.dout(n1492),.clk(gclk));
	jand g1429(.dina(w_n1439_0[0]),.dinb(w_n1420_0[0]),.dout(n1493),.clk(gclk));
	jcb g1430(.dina(n1493),.dinb(w_dff_B_ilQTpZAI4_1),.dout(n1494));
	jand g1431(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1495),.clk(gclk));
	jnot g1432(.din(n1495),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_n1436_0[0]),.dinb(w_n1428_0[0]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1437_0[0]),.dinb(w_n1425_0[0]),.dout(n1498),.clk(gclk));
	jcb g1435(.dina(n1498),.dinb(w_dff_B_UAj1SjrY2_1),.dout(n1499));
	jand g1436(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1501),.clk(gclk));
	jcb g1438(.dina(w_n1433_0[0]),.dinb(w_n1430_0[0]),.dout(n1502));
	jcb g1439(.dina(w_n1435_0[0]),.dinb(w_n1429_0[0]),.dout(n1503));
	jand g1440(.dina(n1503),.dinb(w_dff_B_H9FA1TvV4_1),.dout(n1504),.clk(gclk));
	jxor g1441(.dina(w_n1504_0[1]),.dinb(w_n1501_0[1]),.dout(n1505),.clk(gclk));
	jnot g1442(.din(n1505),.dout(n1506),.clk(gclk));
	jxor g1443(.dina(w_n1506_0[1]),.dinb(w_n1500_0[1]),.dout(n1507),.clk(gclk));
	jxor g1444(.dina(w_n1507_0[1]),.dinb(w_n1499_0[1]),.dout(n1508),.clk(gclk));
	jxor g1445(.dina(w_n1508_0[1]),.dinb(w_n1496_0[1]),.dout(n1509),.clk(gclk));
	jxor g1446(.dina(w_n1509_0[1]),.dinb(w_n1494_0[1]),.dout(n1510),.clk(gclk));
	jxor g1447(.dina(w_n1510_0[1]),.dinb(w_n1491_0[1]),.dout(n1511),.clk(gclk));
	jxor g1448(.dina(w_n1511_0[1]),.dinb(w_n1489_0[1]),.dout(n1512),.clk(gclk));
	jxor g1449(.dina(w_n1512_0[1]),.dinb(w_n1486_0[1]),.dout(n1513),.clk(gclk));
	jxor g1450(.dina(w_n1513_0[1]),.dinb(w_n1484_0[1]),.dout(n1514),.clk(gclk));
	jxor g1451(.dina(w_n1514_0[1]),.dinb(w_n1481_0[1]),.dout(n1515),.clk(gclk));
	jxor g1452(.dina(w_n1515_0[1]),.dinb(w_n1479_0[1]),.dout(n1516),.clk(gclk));
	jxor g1453(.dina(w_n1516_0[1]),.dinb(w_n1476_0[1]),.dout(n1517),.clk(gclk));
	jxor g1454(.dina(w_n1517_0[1]),.dinb(w_n1474_0[1]),.dout(n1518),.clk(gclk));
	jxor g1455(.dina(w_n1518_0[1]),.dinb(w_n1471_0[1]),.dout(n1519),.clk(gclk));
	jxor g1456(.dina(w_n1519_0[1]),.dinb(w_n1469_0[1]),.dout(n1520),.clk(gclk));
	jnot g1457(.din(n1520),.dout(n1521),.clk(gclk));
	jxor g1458(.dina(w_n1521_0[1]),.dinb(w_n1466_0[1]),.dout(n1522),.clk(gclk));
	jnot g1459(.din(n1522),.dout(n1523),.clk(gclk));
	jxor g1460(.dina(w_n1523_0[1]),.dinb(w_n1465_0[1]),.dout(n1524),.clk(gclk));
	jxor g1461(.dina(w_n1524_0[1]),.dinb(w_n1460_0[1]),.dout(G6210gat),.clk(gclk));
	jcb g1462(.dina(w_n1523_0[0]),.dinb(w_n1465_0[0]),.dout(n1526));
	jnot g1463(.din(w_n1524_0[0]),.dout(n1527),.clk(gclk));
	jcb g1464(.dina(w_dff_B_xA4A4SQ38_0),.dinb(w_n1460_0[0]),.dout(n1528));
	jand g1465(.dina(n1528),.dinb(w_dff_B_AIG6bJtq8_1),.dout(n1529),.clk(gclk));
	jnot g1466(.din(w_n1469_0[0]),.dout(n1530),.clk(gclk));
	jnot g1467(.din(w_n1519_0[0]),.dout(n1531),.clk(gclk));
	jcb g1468(.dina(n1531),.dinb(w_dff_B_T1uQ9chI8_1),.dout(n1532));
	jcb g1469(.dina(w_n1521_0[0]),.dinb(w_n1466_0[0]),.dout(n1533));
	jand g1470(.dina(n1533),.dinb(w_dff_B_ZIvl7ino7_1),.dout(n1534),.clk(gclk));
	jand g1471(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1535),.clk(gclk));
	jand g1472(.dina(w_n1517_0[0]),.dinb(w_n1474_0[0]),.dout(n1536),.clk(gclk));
	jand g1473(.dina(w_n1518_0[0]),.dinb(w_n1471_0[0]),.dout(n1537),.clk(gclk));
	jcb g1474(.dina(n1537),.dinb(w_dff_B_liHWSXZD3_1),.dout(n1538));
	jand g1475(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1539),.clk(gclk));
	jnot g1476(.din(n1539),.dout(n1540),.clk(gclk));
	jand g1477(.dina(w_n1515_0[0]),.dinb(w_n1479_0[0]),.dout(n1541),.clk(gclk));
	jand g1478(.dina(w_n1516_0[0]),.dinb(w_n1476_0[0]),.dout(n1542),.clk(gclk));
	jcb g1479(.dina(n1542),.dinb(w_dff_B_u31k2Nk20_1),.dout(n1543));
	jand g1480(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1544),.clk(gclk));
	jnot g1481(.din(n1544),.dout(n1545),.clk(gclk));
	jand g1482(.dina(w_n1513_0[0]),.dinb(w_n1484_0[0]),.dout(n1546),.clk(gclk));
	jand g1483(.dina(w_n1514_0[0]),.dinb(w_n1481_0[0]),.dout(n1547),.clk(gclk));
	jcb g1484(.dina(n1547),.dinb(w_dff_B_3kuIQJaL6_1),.dout(n1548));
	jand g1485(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1549),.clk(gclk));
	jnot g1486(.din(n1549),.dout(n1550),.clk(gclk));
	jand g1487(.dina(w_n1511_0[0]),.dinb(w_n1489_0[0]),.dout(n1551),.clk(gclk));
	jand g1488(.dina(w_n1512_0[0]),.dinb(w_n1486_0[0]),.dout(n1552),.clk(gclk));
	jcb g1489(.dina(n1552),.dinb(w_dff_B_xwntQN6w4_1),.dout(n1553));
	jand g1490(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1554),.clk(gclk));
	jnot g1491(.din(n1554),.dout(n1555),.clk(gclk));
	jand g1492(.dina(w_n1509_0[0]),.dinb(w_n1494_0[0]),.dout(n1556),.clk(gclk));
	jand g1493(.dina(w_n1510_0[0]),.dinb(w_n1491_0[0]),.dout(n1557),.clk(gclk));
	jcb g1494(.dina(n1557),.dinb(w_dff_B_KSa9u7fX3_1),.dout(n1558));
	jand g1495(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1559),.clk(gclk));
	jnot g1496(.din(n1559),.dout(n1560),.clk(gclk));
	jand g1497(.dina(w_n1507_0[0]),.dinb(w_n1499_0[0]),.dout(n1561),.clk(gclk));
	jand g1498(.dina(w_n1508_0[0]),.dinb(w_n1496_0[0]),.dout(n1562),.clk(gclk));
	jcb g1499(.dina(n1562),.dinb(w_dff_B_UvPqCIej8_1),.dout(n1563));
	jand g1500(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1565),.clk(gclk));
	jcb g1502(.dina(w_n1504_0[0]),.dinb(w_n1501_0[0]),.dout(n1566));
	jcb g1503(.dina(w_n1506_0[0]),.dinb(w_n1500_0[0]),.dout(n1567));
	jand g1504(.dina(n1567),.dinb(w_dff_B_rttLFnrN8_1),.dout(n1568),.clk(gclk));
	jxor g1505(.dina(w_n1568_0[1]),.dinb(w_n1565_0[1]),.dout(n1569),.clk(gclk));
	jnot g1506(.din(n1569),.dout(n1570),.clk(gclk));
	jxor g1507(.dina(w_n1570_0[1]),.dinb(w_n1564_0[1]),.dout(n1571),.clk(gclk));
	jxor g1508(.dina(w_n1571_0[1]),.dinb(w_n1563_0[1]),.dout(n1572),.clk(gclk));
	jxor g1509(.dina(w_n1572_0[1]),.dinb(w_n1560_0[1]),.dout(n1573),.clk(gclk));
	jxor g1510(.dina(w_n1573_0[1]),.dinb(w_n1558_0[1]),.dout(n1574),.clk(gclk));
	jxor g1511(.dina(w_n1574_0[1]),.dinb(w_n1555_0[1]),.dout(n1575),.clk(gclk));
	jxor g1512(.dina(w_n1575_0[1]),.dinb(w_n1553_0[1]),.dout(n1576),.clk(gclk));
	jxor g1513(.dina(w_n1576_0[1]),.dinb(w_n1550_0[1]),.dout(n1577),.clk(gclk));
	jxor g1514(.dina(w_n1577_0[1]),.dinb(w_n1548_0[1]),.dout(n1578),.clk(gclk));
	jxor g1515(.dina(w_n1578_0[1]),.dinb(w_n1545_0[1]),.dout(n1579),.clk(gclk));
	jxor g1516(.dina(w_n1579_0[1]),.dinb(w_n1543_0[1]),.dout(n1580),.clk(gclk));
	jxor g1517(.dina(w_n1580_0[1]),.dinb(w_n1540_0[1]),.dout(n1581),.clk(gclk));
	jxor g1518(.dina(w_n1581_0[1]),.dinb(w_n1538_0[1]),.dout(n1582),.clk(gclk));
	jnot g1519(.din(n1582),.dout(n1583),.clk(gclk));
	jxor g1520(.dina(w_n1583_0[1]),.dinb(w_n1535_0[1]),.dout(n1584),.clk(gclk));
	jnot g1521(.din(n1584),.dout(n1585),.clk(gclk));
	jxor g1522(.dina(w_n1585_0[1]),.dinb(w_n1534_0[1]),.dout(n1586),.clk(gclk));
	jxor g1523(.dina(w_n1586_0[1]),.dinb(w_n1529_0[1]),.dout(G6220gat),.clk(gclk));
	jcb g1524(.dina(w_n1585_0[0]),.dinb(w_n1534_0[0]),.dout(n1588));
	jnot g1525(.din(w_n1586_0[0]),.dout(n1589),.clk(gclk));
	jcb g1526(.dina(w_dff_B_FwpMwxfk6_0),.dinb(w_n1529_0[0]),.dout(n1590));
	jand g1527(.dina(n1590),.dinb(w_dff_B_UekR6NNa3_1),.dout(n1591),.clk(gclk));
	jnot g1528(.din(w_n1538_0[0]),.dout(n1592),.clk(gclk));
	jnot g1529(.din(w_n1581_0[0]),.dout(n1593),.clk(gclk));
	jcb g1530(.dina(n1593),.dinb(w_dff_B_vDgUCxtX0_1),.dout(n1594));
	jcb g1531(.dina(w_n1583_0[0]),.dinb(w_n1535_0[0]),.dout(n1595));
	jand g1532(.dina(n1595),.dinb(w_dff_B_4BsIzBMw6_1),.dout(n1596),.clk(gclk));
	jand g1533(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1597),.clk(gclk));
	jand g1534(.dina(w_n1579_0[0]),.dinb(w_n1543_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(w_n1580_0[0]),.dinb(w_n1540_0[0]),.dout(n1599),.clk(gclk));
	jcb g1536(.dina(n1599),.dinb(w_dff_B_TSNOL1hx3_1),.dout(n1600));
	jand g1537(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1601),.clk(gclk));
	jnot g1538(.din(n1601),.dout(n1602),.clk(gclk));
	jand g1539(.dina(w_n1577_0[0]),.dinb(w_n1548_0[0]),.dout(n1603),.clk(gclk));
	jand g1540(.dina(w_n1578_0[0]),.dinb(w_n1545_0[0]),.dout(n1604),.clk(gclk));
	jcb g1541(.dina(n1604),.dinb(w_dff_B_m01alN119_1),.dout(n1605));
	jand g1542(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1606),.clk(gclk));
	jnot g1543(.din(n1606),.dout(n1607),.clk(gclk));
	jand g1544(.dina(w_n1575_0[0]),.dinb(w_n1553_0[0]),.dout(n1608),.clk(gclk));
	jand g1545(.dina(w_n1576_0[0]),.dinb(w_n1550_0[0]),.dout(n1609),.clk(gclk));
	jcb g1546(.dina(n1609),.dinb(w_dff_B_QUxCrnrP2_1),.dout(n1610));
	jand g1547(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1611),.clk(gclk));
	jnot g1548(.din(n1611),.dout(n1612),.clk(gclk));
	jand g1549(.dina(w_n1573_0[0]),.dinb(w_n1558_0[0]),.dout(n1613),.clk(gclk));
	jand g1550(.dina(w_n1574_0[0]),.dinb(w_n1555_0[0]),.dout(n1614),.clk(gclk));
	jcb g1551(.dina(n1614),.dinb(w_dff_B_xWWDbt2V5_1),.dout(n1615));
	jand g1552(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1616),.clk(gclk));
	jnot g1553(.din(n1616),.dout(n1617),.clk(gclk));
	jand g1554(.dina(w_n1571_0[0]),.dinb(w_n1563_0[0]),.dout(n1618),.clk(gclk));
	jand g1555(.dina(w_n1572_0[0]),.dinb(w_n1560_0[0]),.dout(n1619),.clk(gclk));
	jcb g1556(.dina(n1619),.dinb(w_dff_B_MNUGWboP9_1),.dout(n1620));
	jand g1557(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1622),.clk(gclk));
	jcb g1559(.dina(w_n1568_0[0]),.dinb(w_n1565_0[0]),.dout(n1623));
	jcb g1560(.dina(w_n1570_0[0]),.dinb(w_n1564_0[0]),.dout(n1624));
	jand g1561(.dina(n1624),.dinb(w_dff_B_fUp5carD2_1),.dout(n1625),.clk(gclk));
	jxor g1562(.dina(w_n1625_0[1]),.dinb(w_n1622_0[1]),.dout(n1626),.clk(gclk));
	jnot g1563(.din(n1626),.dout(n1627),.clk(gclk));
	jxor g1564(.dina(w_n1627_0[1]),.dinb(w_n1621_0[1]),.dout(n1628),.clk(gclk));
	jxor g1565(.dina(w_n1628_0[1]),.dinb(w_n1620_0[1]),.dout(n1629),.clk(gclk));
	jxor g1566(.dina(w_n1629_0[1]),.dinb(w_n1617_0[1]),.dout(n1630),.clk(gclk));
	jxor g1567(.dina(w_n1630_0[1]),.dinb(w_n1615_0[1]),.dout(n1631),.clk(gclk));
	jxor g1568(.dina(w_n1631_0[1]),.dinb(w_n1612_0[1]),.dout(n1632),.clk(gclk));
	jxor g1569(.dina(w_n1632_0[1]),.dinb(w_n1610_0[1]),.dout(n1633),.clk(gclk));
	jxor g1570(.dina(w_n1633_0[1]),.dinb(w_n1607_0[1]),.dout(n1634),.clk(gclk));
	jxor g1571(.dina(w_n1634_0[1]),.dinb(w_n1605_0[1]),.dout(n1635),.clk(gclk));
	jxor g1572(.dina(w_n1635_0[1]),.dinb(w_n1602_0[1]),.dout(n1636),.clk(gclk));
	jxor g1573(.dina(w_n1636_0[1]),.dinb(w_n1600_0[1]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jxor g1575(.dina(w_n1638_0[1]),.dinb(w_n1597_0[1]),.dout(n1639),.clk(gclk));
	jnot g1576(.din(n1639),.dout(n1640),.clk(gclk));
	jxor g1577(.dina(w_n1640_0[1]),.dinb(w_n1596_0[1]),.dout(n1641),.clk(gclk));
	jxor g1578(.dina(w_n1641_0[1]),.dinb(w_n1591_0[1]),.dout(G6230gat),.clk(gclk));
	jcb g1579(.dina(w_n1640_0[0]),.dinb(w_n1596_0[0]),.dout(n1643));
	jnot g1580(.din(w_n1641_0[0]),.dout(n1644),.clk(gclk));
	jcb g1581(.dina(w_dff_B_f4Eih3xY4_0),.dinb(w_n1591_0[0]),.dout(n1645));
	jand g1582(.dina(n1645),.dinb(w_dff_B_8QhDajyx7_1),.dout(n1646),.clk(gclk));
	jnot g1583(.din(w_n1600_0[0]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(w_n1636_0[0]),.dout(n1648),.clk(gclk));
	jcb g1585(.dina(n1648),.dinb(w_dff_B_e2z1JxOl1_1),.dout(n1649));
	jcb g1586(.dina(w_n1638_0[0]),.dinb(w_n1597_0[0]),.dout(n1650));
	jand g1587(.dina(n1650),.dinb(w_dff_B_mkSi4f4V7_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1652),.clk(gclk));
	jnot g1589(.din(n1652),.dout(n1653),.clk(gclk));
	jand g1590(.dina(w_n1634_0[0]),.dinb(w_n1605_0[0]),.dout(n1654),.clk(gclk));
	jand g1591(.dina(w_n1635_0[0]),.dinb(w_n1602_0[0]),.dout(n1655),.clk(gclk));
	jcb g1592(.dina(n1655),.dinb(w_dff_B_QOTySqd87_1),.dout(n1656));
	jand g1593(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jand g1595(.dina(w_n1632_0[0]),.dinb(w_n1610_0[0]),.dout(n1659),.clk(gclk));
	jand g1596(.dina(w_n1633_0[0]),.dinb(w_n1607_0[0]),.dout(n1660),.clk(gclk));
	jcb g1597(.dina(n1660),.dinb(w_dff_B_8YAqrqWn5_1),.dout(n1661));
	jand g1598(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1662),.clk(gclk));
	jnot g1599(.din(n1662),.dout(n1663),.clk(gclk));
	jand g1600(.dina(w_n1630_0[0]),.dinb(w_n1615_0[0]),.dout(n1664),.clk(gclk));
	jand g1601(.dina(w_n1631_0[0]),.dinb(w_n1612_0[0]),.dout(n1665),.clk(gclk));
	jcb g1602(.dina(n1665),.dinb(w_dff_B_nxmiywbP2_1),.dout(n1666));
	jand g1603(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1667),.clk(gclk));
	jnot g1604(.din(n1667),.dout(n1668),.clk(gclk));
	jand g1605(.dina(w_n1628_0[0]),.dinb(w_n1620_0[0]),.dout(n1669),.clk(gclk));
	jand g1606(.dina(w_n1629_0[0]),.dinb(w_n1617_0[0]),.dout(n1670),.clk(gclk));
	jcb g1607(.dina(n1670),.dinb(w_dff_B_axwawoWk7_1),.dout(n1671));
	jand g1608(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1672),.clk(gclk));
	jand g1609(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1673),.clk(gclk));
	jcb g1610(.dina(w_n1625_0[0]),.dinb(w_n1622_0[0]),.dout(n1674));
	jcb g1611(.dina(w_n1627_0[0]),.dinb(w_n1621_0[0]),.dout(n1675));
	jand g1612(.dina(n1675),.dinb(w_dff_B_OLhctYmw4_1),.dout(n1676),.clk(gclk));
	jxor g1613(.dina(w_n1676_0[1]),.dinb(w_n1673_0[1]),.dout(n1677),.clk(gclk));
	jnot g1614(.din(n1677),.dout(n1678),.clk(gclk));
	jxor g1615(.dina(w_n1678_0[1]),.dinb(w_n1672_0[1]),.dout(n1679),.clk(gclk));
	jxor g1616(.dina(w_n1679_0[1]),.dinb(w_n1671_0[1]),.dout(n1680),.clk(gclk));
	jxor g1617(.dina(w_n1680_0[1]),.dinb(w_n1668_0[1]),.dout(n1681),.clk(gclk));
	jxor g1618(.dina(w_n1681_0[1]),.dinb(w_n1666_0[1]),.dout(n1682),.clk(gclk));
	jxor g1619(.dina(w_n1682_0[1]),.dinb(w_n1663_0[1]),.dout(n1683),.clk(gclk));
	jxor g1620(.dina(w_n1683_0[1]),.dinb(w_n1661_0[1]),.dout(n1684),.clk(gclk));
	jxor g1621(.dina(w_n1684_0[1]),.dinb(w_n1658_0[1]),.dout(n1685),.clk(gclk));
	jxor g1622(.dina(w_n1685_0[1]),.dinb(w_n1656_0[1]),.dout(n1686),.clk(gclk));
	jxor g1623(.dina(w_n1686_0[1]),.dinb(w_n1653_0[1]),.dout(n1687),.clk(gclk));
	jnot g1624(.din(n1687),.dout(n1688),.clk(gclk));
	jxor g1625(.dina(w_n1688_0[1]),.dinb(w_n1651_0[1]),.dout(n1689),.clk(gclk));
	jxor g1626(.dina(w_n1689_0[1]),.dinb(w_n1646_0[1]),.dout(G6240gat),.clk(gclk));
	jcb g1627(.dina(w_n1688_0[0]),.dinb(w_n1651_0[0]),.dout(n1691));
	jnot g1628(.din(w_n1689_0[0]),.dout(n1692),.clk(gclk));
	jcb g1629(.dina(w_dff_B_dN7mMsn83_0),.dinb(w_n1646_0[0]),.dout(n1693));
	jand g1630(.dina(n1693),.dinb(w_dff_B_3YCoDQeY1_1),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1685_0[0]),.dinb(w_n1656_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1686_0[0]),.dinb(w_n1653_0[0]),.dout(n1696),.clk(gclk));
	jcb g1633(.dina(n1696),.dinb(w_dff_B_32RUcBr69_1),.dout(n1697));
	jand g1634(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1683_0[0]),.dinb(w_n1661_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1684_0[0]),.dinb(w_n1658_0[0]),.dout(n1701),.clk(gclk));
	jcb g1638(.dina(n1701),.dinb(w_dff_B_bWhd0JRq4_1),.dout(n1702));
	jand g1639(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1703),.clk(gclk));
	jnot g1640(.din(n1703),.dout(n1704),.clk(gclk));
	jand g1641(.dina(w_n1681_0[0]),.dinb(w_n1666_0[0]),.dout(n1705),.clk(gclk));
	jand g1642(.dina(w_n1682_0[0]),.dinb(w_n1663_0[0]),.dout(n1706),.clk(gclk));
	jcb g1643(.dina(n1706),.dinb(w_dff_B_Q2VG2qeG7_1),.dout(n1707));
	jand g1644(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jand g1646(.dina(w_n1679_0[0]),.dinb(w_n1671_0[0]),.dout(n1710),.clk(gclk));
	jand g1647(.dina(w_n1680_0[0]),.dinb(w_n1668_0[0]),.dout(n1711),.clk(gclk));
	jcb g1648(.dina(n1711),.dinb(w_dff_B_sTlKSnnr0_1),.dout(n1712));
	jand g1649(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1713),.clk(gclk));
	jand g1650(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1714),.clk(gclk));
	jcb g1651(.dina(w_n1676_0[0]),.dinb(w_n1673_0[0]),.dout(n1715));
	jcb g1652(.dina(w_n1678_0[0]),.dinb(w_n1672_0[0]),.dout(n1716));
	jand g1653(.dina(n1716),.dinb(w_dff_B_wQmsM3qk1_1),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1714_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1713_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1712_0[1]),.dout(n1721),.clk(gclk));
	jxor g1658(.dina(w_n1721_0[1]),.dinb(w_n1709_0[1]),.dout(n1722),.clk(gclk));
	jxor g1659(.dina(w_n1722_0[1]),.dinb(w_n1707_0[1]),.dout(n1723),.clk(gclk));
	jxor g1660(.dina(w_n1723_0[1]),.dinb(w_n1704_0[1]),.dout(n1724),.clk(gclk));
	jxor g1661(.dina(w_n1724_0[1]),.dinb(w_n1702_0[1]),.dout(n1725),.clk(gclk));
	jxor g1662(.dina(w_n1725_0[1]),.dinb(w_n1699_0[1]),.dout(n1726),.clk(gclk));
	jxor g1663(.dina(w_n1726_0[1]),.dinb(w_n1697_0[1]),.dout(n1727),.clk(gclk));
	jxor g1664(.dina(w_n1727_0[1]),.dinb(w_n1694_0[1]),.dout(G6250gat),.clk(gclk));
	jnot g1665(.din(w_n1697_0[0]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(w_n1726_0[0]),.dout(n1730),.clk(gclk));
	jcb g1667(.dina(n1730),.dinb(w_dff_B_PE4m5ZCu8_1),.dout(n1731));
	jnot g1668(.din(w_n1727_0[0]),.dout(n1732),.clk(gclk));
	jcb g1669(.dina(w_dff_B_lculz7TR9_0),.dinb(w_n1694_0[0]),.dout(n1733));
	jand g1670(.dina(n1733),.dinb(w_dff_B_v9bnab3R2_1),.dout(n1734),.clk(gclk));
	jand g1671(.dina(w_n1724_0[0]),.dinb(w_n1702_0[0]),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1725_0[0]),.dinb(w_n1699_0[0]),.dout(n1736),.clk(gclk));
	jcb g1673(.dina(n1736),.dinb(w_dff_B_zn1GqKHr3_1),.dout(n1737));
	jand g1674(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1738),.clk(gclk));
	jnot g1675(.din(n1738),.dout(n1739),.clk(gclk));
	jand g1676(.dina(w_n1722_0[0]),.dinb(w_n1707_0[0]),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1723_0[0]),.dinb(w_n1704_0[0]),.dout(n1741),.clk(gclk));
	jcb g1678(.dina(n1741),.dinb(w_dff_B_Ds0vKPck1_1),.dout(n1742));
	jand g1679(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1743),.clk(gclk));
	jnot g1680(.din(n1743),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_n1720_0[0]),.dinb(w_n1712_0[0]),.dout(n1745),.clk(gclk));
	jand g1682(.dina(w_n1721_0[0]),.dinb(w_n1709_0[0]),.dout(n1746),.clk(gclk));
	jcb g1683(.dina(n1746),.dinb(w_dff_B_KAPZZ2M51_1),.dout(n1747));
	jand g1684(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1748),.clk(gclk));
	jand g1685(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1749),.clk(gclk));
	jcb g1686(.dina(w_n1717_0[0]),.dinb(w_n1714_0[0]),.dout(n1750));
	jcb g1687(.dina(w_n1719_0[0]),.dinb(w_n1713_0[0]),.dout(n1751));
	jand g1688(.dina(n1751),.dinb(w_dff_B_C8UvJwn70_1),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1749_0[1]),.dout(n1753),.clk(gclk));
	jnot g1690(.din(n1753),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1748_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1747_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1744_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1742_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1739_0[1]),.dout(n1759),.clk(gclk));
	jxor g1696(.dina(w_n1759_0[1]),.dinb(w_n1737_0[1]),.dout(n1760),.clk(gclk));
	jxor g1697(.dina(w_n1760_0[1]),.dinb(w_n1734_0[1]),.dout(G6260gat),.clk(gclk));
	jnot g1698(.din(w_n1737_0[0]),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1759_0[0]),.dout(n1763),.clk(gclk));
	jcb g1700(.dina(n1763),.dinb(w_dff_B_s9URHH6X8_1),.dout(n1764));
	jnot g1701(.din(w_n1760_0[0]),.dout(n1765),.clk(gclk));
	jcb g1702(.dina(w_dff_B_5ubhJ4Ul9_0),.dinb(w_n1734_0[0]),.dout(n1766));
	jand g1703(.dina(n1766),.dinb(w_dff_B_LBz8FDdd7_1),.dout(n1767),.clk(gclk));
	jand g1704(.dina(w_n1757_0[0]),.dinb(w_n1742_0[0]),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_n1758_0[0]),.dinb(w_n1739_0[0]),.dout(n1769),.clk(gclk));
	jcb g1706(.dina(n1769),.dinb(w_dff_B_B1fTr3EQ0_1),.dout(n1770));
	jand g1707(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1771),.clk(gclk));
	jnot g1708(.din(n1771),.dout(n1772),.clk(gclk));
	jand g1709(.dina(w_n1755_0[0]),.dinb(w_n1747_0[0]),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_n1756_0[0]),.dinb(w_n1744_0[0]),.dout(n1774),.clk(gclk));
	jcb g1711(.dina(n1774),.dinb(w_dff_B_OVlA1riG1_1),.dout(n1775));
	jand g1712(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1777),.clk(gclk));
	jcb g1714(.dina(w_n1752_0[0]),.dinb(w_n1749_0[0]),.dout(n1778));
	jcb g1715(.dina(w_n1754_0[0]),.dinb(w_n1748_0[0]),.dout(n1779));
	jand g1716(.dina(n1779),.dinb(w_dff_B_zYTpJKxQ4_1),.dout(n1780),.clk(gclk));
	jxor g1717(.dina(w_n1780_0[1]),.dinb(w_n1777_0[1]),.dout(n1781),.clk(gclk));
	jnot g1718(.din(n1781),.dout(n1782),.clk(gclk));
	jxor g1719(.dina(w_n1782_0[1]),.dinb(w_n1776_0[1]),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1775_0[1]),.dout(n1784),.clk(gclk));
	jxor g1721(.dina(w_n1784_0[1]),.dinb(w_n1772_0[1]),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1770_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1767_0[1]),.dout(G6270gat),.clk(gclk));
	jnot g1724(.din(w_n1770_0[0]),.dout(n1788),.clk(gclk));
	jnot g1725(.din(w_n1785_0[0]),.dout(n1789),.clk(gclk));
	jcb g1726(.dina(n1789),.dinb(w_dff_B_wMZixJ0t3_1),.dout(n1790));
	jnot g1727(.din(w_n1786_0[0]),.dout(n1791),.clk(gclk));
	jcb g1728(.dina(w_dff_B_UKeQvCg87_0),.dinb(w_n1767_0[0]),.dout(n1792));
	jand g1729(.dina(n1792),.dinb(w_dff_B_SeIcI13K2_1),.dout(n1793),.clk(gclk));
	jand g1730(.dina(w_n1783_0[0]),.dinb(w_n1775_0[0]),.dout(n1794),.clk(gclk));
	jand g1731(.dina(w_n1784_0[0]),.dinb(w_n1772_0[0]),.dout(n1795),.clk(gclk));
	jcb g1732(.dina(n1795),.dinb(w_dff_B_Ve2vwywr3_1),.dout(n1796));
	jand g1733(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1798),.clk(gclk));
	jcb g1735(.dina(w_n1780_0[0]),.dinb(w_n1777_0[0]),.dout(n1799));
	jcb g1736(.dina(w_n1782_0[0]),.dinb(w_n1776_0[0]),.dout(n1800));
	jand g1737(.dina(n1800),.dinb(w_dff_B_CF2m4dVa4_1),.dout(n1801),.clk(gclk));
	jxor g1738(.dina(w_n1801_0[1]),.dinb(w_n1798_0[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jxor g1740(.dina(w_n1803_0[1]),.dinb(w_n1797_0[1]),.dout(n1804),.clk(gclk));
	jxor g1741(.dina(w_n1804_0[1]),.dinb(w_n1796_0[1]),.dout(n1805),.clk(gclk));
	jxor g1742(.dina(w_n1805_0[1]),.dinb(w_n1793_0[1]),.dout(G6280gat),.clk(gclk));
	jand g1743(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1807),.clk(gclk));
	jcb g1744(.dina(w_n1801_0[0]),.dinb(w_n1798_0[0]),.dout(n1808));
	jcb g1745(.dina(w_n1803_0[0]),.dinb(w_n1797_0[0]),.dout(n1809));
	jand g1746(.dina(n1809),.dinb(w_dff_B_mn4rCjzz0_1),.dout(n1810),.clk(gclk));
	jcb g1747(.dina(w_n1810_0[1]),.dinb(w_n1807_0[1]),.dout(n1811));
	jnot g1748(.din(w_n1796_0[0]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(w_n1804_0[0]),.dout(n1813),.clk(gclk));
	jcb g1750(.dina(n1813),.dinb(w_dff_B_uCql4FRT2_1),.dout(n1814));
	jnot g1751(.din(w_n1805_0[0]),.dout(n1815),.clk(gclk));
	jcb g1752(.dina(w_dff_B_S4ltgIP69_0),.dinb(w_n1793_0[0]),.dout(n1816));
	jand g1753(.dina(n1816),.dinb(w_dff_B_LWJ4q85k1_1),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1810_0[0]),.dinb(w_n1807_0[0]),.dout(n1818),.clk(gclk));
	jnot g1755(.din(w_n1818_0[1]),.dout(n1819),.clk(gclk));
	jcb g1756(.dina(w_dff_B_Hud6zxaB7_0),.dinb(w_n1817_0[1]),.dout(n1820));
	jand g1757(.dina(n1820),.dinb(w_dff_B_SYkn1LZE6_1),.dout(G6287gat),.clk(gclk));
	jxor g1758(.dina(w_n1818_0[0]),.dinb(w_n1817_0[0]),.dout(G6288gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl jspl_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl jspl_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_G307gat_2[1]),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl jspl_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(G545gat),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_n66_0[0]),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n75_0(.douta(w_dff_A_D8ZagyVs8_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n80_0(.douta(w_dff_A_4He3wXXc8_0),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_dff_A_KsYCjYWA6_1),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_Ck4bOiEB2_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_dff_A_ScPbN5a19_0),.doutb(w_n91_0[1]),.din(n91));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_Bv8lsQaE1_1),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_AFqrBfsz6_0),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n111_0(.douta(w_dff_A_xbYlxVGw3_0),.doutb(w_n111_0[1]),.din(w_dff_B_CIHAMHnt6_2));
	jspl jspl_w_n112_0(.douta(w_dff_A_YElQJLx72_0),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_rLbe5iWw9_1),.doutc(w_dff_A_WU05vbqJ5_2),.din(w_dff_B_qOlwIYSL5_3));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(w_dff_B_AmgMx0zO2_2));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(w_dff_B_XyxqOr217_2));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n122_0(.douta(w_dff_A_o1vhWlM35_0),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n123_0(.douta(w_dff_A_kkCyMRDe5_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.din(n133));
	jspl jspl_w_n135_0(.douta(w_dff_A_gUdkwqQc8_0),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n140_0(.douta(w_dff_A_mwVSDR3y2_0),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_EVTnbB3G6_0),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_t9jJ0Ax06_1),.doutc(w_dff_A_ZnVzuhX42_2),.din(n146));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(w_dff_B_U9BSC4ub3_2));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(w_dff_B_IQchRE107_2));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_dff_A_lXNE1JWt6_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_dff_A_VFk9IOOo6_0),.doutb(w_n157_0[1]),.din(n157));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl jspl_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl jspl_w_n170_0(.douta(w_dff_A_a0PbLUTj5_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n175_0(.douta(w_dff_A_urhleK3H5_0),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n176_0(.douta(w_dff_A_BpAHiX1R2_0),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_dff_A_oiF60WcB7_1),.doutc(w_dff_A_Cvh7nZWc3_2),.din(n181));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.din(w_dff_B_a0xbI5MR9_2));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(w_dff_B_AxwWbGXe2_2));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.din(w_dff_B_cbd2tEGR6_2));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_hY78nFfS1_0),.doutb(w_dff_A_TMMq93Z77_1),.doutc(w_n196_0[2]),.din(n196));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_dff_A_EEibSwoO2_0),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n217_0(.douta(w_dff_A_oI3U0KAt2_0),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_dff_A_AMQHIN923_0),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_dff_A_0A3wwcWf1_1),.doutc(w_dff_A_c04hZHBx0_2),.din(n223));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(w_dff_B_KZLo3TkJ9_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(w_dff_B_hzjeHgL23_2));
	jspl jspl_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.din(n233));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(w_dff_B_2vHWrEiA8_2));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(w_dff_B_IBrwA5D33_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_dff_A_D70Zf41k4_0),.doutb(w_dff_A_8uBIIrPF3_1),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(n251));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(n253));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_dff_A_a0Q0MiLY4_0),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n266_0(.douta(w_dff_A_GJdiBsWB7_0),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_dff_A_LOYtCh2c3_0),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n272_0(.douta(w_n272_0[0]),.doutb(w_dff_A_0tGESKVt5_1),.doutc(w_dff_A_naHyJ4d17_2),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_aOXfa8sz8_2));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_xv1nQ7vz8_2));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(w_dff_B_dbs0Nf4r4_2));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(w_dff_B_ZXoeUWOj6_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_1jyfj3PW8_2));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl3 jspl3_w_n297_0(.douta(w_dff_A_i0usyGzS7_0),.doutb(w_dff_A_q2evcYDZ5_1),.doutc(w_n297_0[2]),.din(n297));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.din(n306));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(n307));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_dff_A_hreXLba73_0),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n322_0(.douta(w_dff_A_tA5PPiBy4_0),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_dff_A_YabRlF152_0),.doutb(w_n323_0[1]),.din(n323));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_dff_A_0eoWrf1S3_1),.doutc(w_dff_A_iwaBUwCU1_2),.din(n328));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(w_dff_B_XG3grkrj8_2));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(w_dff_B_bnx2wppo4_2));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(w_dff_B_4Dj13Jvy2_2));
	jspl jspl_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(w_dff_B_teCrdQ8K5_2));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(w_dff_B_xso4Npzq4_2));
	jspl jspl_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.din(n354));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(w_dff_B_fhv5ubir5_2));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n358_0(.douta(w_dff_A_BwRsfu1h5_0),.doutb(w_dff_A_JeJnM9zr2_1),.doutc(w_n358_0[2]),.din(n358));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(n363));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl jspl_w_n380_0(.douta(w_dff_A_eEk6Vttx5_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n385_0(.douta(w_dff_A_UPGQO3ku6_0),.doutb(w_n385_0[1]),.din(w_dff_B_WvtuT2Pi5_2));
	jspl jspl_w_n386_0(.douta(w_dff_A_91CmjfIu8_0),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_dff_A_X4AjoJhn4_1),.doutc(w_dff_A_uXsEZDhL1_2),.din(w_dff_B_c9r1jGgp4_3));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(w_dff_B_fgyzPuhR6_2));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(w_dff_B_N4sh3q5e5_2));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(w_dff_B_gd3sCwu39_2));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(w_dff_B_1aTwimwz5_2));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(w_dff_B_1MUQayca2_2));
	jspl jspl_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.din(w_dff_B_M9Ywdoct1_2));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(w_dff_B_n8pcLXAT9_2));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(w_dff_B_yFFnSilg5_2));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(w_dff_B_VdCinP0T1_2));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(w_dff_B_RodJbxBX1_2));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(w_dff_B_2l0AIDKB1_2));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(w_dff_B_tL739E4x0_2));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_dff_A_MVF4fcjn7_0),.doutb(w_dff_A_BMAwMXjb2_1),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(n432));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(w_dff_B_NqcXKRfB2_2));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(n439));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl jspl_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.din(n449));
	jspl jspl_w_n451_0(.douta(w_dff_A_oHHeRJzx3_0),.doutb(w_n451_0[1]),.din(n451));
	jspl jspl_w_n456_0(.douta(w_dff_A_u8VsDPPC5_0),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_dff_A_ILxVErOV7_0),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_I5tXqzfD0_1),.doutc(w_dff_A_QfR65i8R2_2),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(w_dff_B_48wM55a46_2));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(w_dff_B_mMtDY7Ft3_2));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(w_dff_B_r65m0gHm0_2));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(w_dff_B_tm99xvrP5_2));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_W0AeNeTW6_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_axgwUMrn3_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_R9xRJ5ll5_2));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(w_dff_B_tds3ch0X2_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl3 jspl3_w_n503_0(.douta(w_dff_A_rrIgy5qa0_0),.doutb(w_dff_A_DK2WnL0g7_1),.doutc(w_n503_0[2]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_UcTBY1zo6_2));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.din(n515));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.din(n521));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl jspl_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n526_0(.douta(w_n526_0[0]),.doutb(w_n526_0[1]),.din(n526));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_dff_A_heUPJXR54_0),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n534_0(.douta(w_dff_A_XGY45YLI0_0),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_dff_A_A06Hb1ms3_0),.doutb(w_n535_0[1]),.din(n535));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_dff_A_ZQVdk6Lq8_1),.doutc(w_dff_A_gfmfUuPd7_2),.din(n540));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_CtXZPoD54_2));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(w_dff_B_U7tVD6sA5_2));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(w_dff_B_dGoD1wjK8_2));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(w_dff_B_xLVoL2A89_2));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(w_dff_B_9aOUgWIu3_2));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(w_dff_B_55nlJBQr7_2));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(w_dff_B_v8dDabgb2_2));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(w_dff_B_1NLc7XxL1_2));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(w_dff_B_tLuPYHai7_2));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n586_0(.douta(w_dff_A_QsWz4K3z1_0),.doutb(w_dff_A_5I1E6S8T8_1),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(w_dff_B_N5Yqmrr39_2));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.din(n594));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n611_0(.douta(w_n611_0[0]),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n614_0(.douta(w_dff_A_RK6NV3yY4_0),.doutb(w_n614_0[1]),.din(n614));
	jspl jspl_w_n619_0(.douta(w_dff_A_wpS1r5Ve3_0),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_dff_A_lbCS54R79_0),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_dff_A_cjuBMvDR1_1),.doutc(w_dff_A_1CFFVbwM8_2),.din(n625));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(w_dff_B_HJozdlbv8_2));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(w_dff_B_GTVULd038_2));
	jspl jspl_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(w_dff_B_Ja40IbTs7_2));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(w_dff_B_KJsm2iQ82_2));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(w_dff_B_nQgUO1Pw2_2));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_jbGt7EVX8_2));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(w_dff_B_nJrMpPDH9_2));
	jspl jspl_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.din(n660));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(w_dff_B_z6gQ9hNy3_2));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(w_dff_B_pfmOU5sT4_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_WlqYnXpZ5_2));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl3 jspl3_w_n676_0(.douta(w_dff_A_uEHtC4hr1_0),.doutb(w_dff_A_7ZLP7fsA9_1),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(w_dff_B_YIhjSKK65_2));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.din(n688));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(n694));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n706_0(.douta(w_dff_A_4rh7ihgJ1_0),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n711_0(.douta(w_dff_A_u0s3Zbqb3_0),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_dff_A_bENhUFb61_0),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_QQiW9jHY7_1),.doutc(w_dff_A_UZCyLOk90_2),.din(n717));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_7jkSTk9B6_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(w_dff_B_RAjW8tPC7_2));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(w_dff_B_0G4BkaBJ6_2));
	jspl jspl_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.din(n732));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(w_dff_B_vZt4kRgy3_2));
	jspl jspl_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.din(n737));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(w_dff_B_FAqUrTuV1_2));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.din(w_dff_B_ej1hnLyh5_2));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(w_dff_B_8lzSH3qA1_2));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(w_dff_B_sglmE4pR1_2));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(w_dff_B_QriFem3S1_2));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(w_dff_B_jSQRXVU61_2));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(w_dff_B_M7dKjfdi0_2));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(w_dff_B_CWBZljMi1_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(n781));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(n783));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(n787));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.din(n790));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.din(n794));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl jspl_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.din(n799));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n805_0(.douta(w_dff_A_SHL8gzUL6_0),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_USy1Trii9_2));
	jspl jspl_w_n815_0(.douta(w_dff_A_DcHsrmTj0_0),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_dff_A_XGAWw9VZ5_0),.doutb(w_n816_0[1]),.din(n816));
	jspl3 jspl3_w_n820_0(.douta(w_dff_A_x6b9m6GW6_0),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(w_dff_B_h6QApWVR7_2));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(w_dff_B_Ur8YsLTJ9_2));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(w_dff_B_mWheOF5C7_2));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(w_dff_B_46mVB41B0_2));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(w_dff_B_pHEqSSlV6_2));
	jspl jspl_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.din(n845));
	jspl jspl_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.din(w_dff_B_G3u1fkFI6_2));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(w_dff_B_44BG7z7r0_2));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(w_dff_B_Jii61y7X1_2));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(w_dff_B_9QT1Zgay3_2));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(w_dff_B_rnVyKTkM6_2));
	jspl jspl_w_n872_0(.douta(w_n872_0[0]),.doutb(w_n872_0[1]),.din(n872));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(w_dff_B_xjGe0H5j2_2));
	jspl jspl_w_n875_0(.douta(w_dff_A_64J3g8NG2_0),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n877_0(.douta(w_dff_A_d5Hs080Z2_0),.doutb(w_n877_0[1]),.din(w_dff_B_NlKQY1ue6_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(w_dff_B_LAz1Hdqf1_2));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(n882));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(n886));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.din(n888));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(n898));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.doutc(w_n900_0[2]),.din(n900));
	jspl jspl_w_n902_0(.douta(w_n902_0[0]),.doutb(w_n902_0[1]),.din(n902));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_dff_A_r2CxQq4M1_1),.din(n904));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(w_dff_B_YNvCsceP4_2));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_dff_A_mXBLWQWm6_1),.din(w_dff_B_GLO8DITt9_2));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_dff_A_03eNmzSV3_1),.doutc(w_dff_A_UvcgMejF3_2),.din(w_dff_B_Pl34Mh8Q8_3));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(w_dff_B_aGAepYLi9_2));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(w_dff_B_8HzqBeLN7_2));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(w_dff_B_vj0XLNQO7_2));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.din(w_dff_B_PBlOLn9W3_2));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(w_dff_B_RV3WkNZc5_2));
	jspl jspl_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.din(n942));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(w_dff_B_M9eT0cLQ5_2));
	jspl jspl_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.din(n947));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(w_dff_B_HZ2Qo92N7_2));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(w_dff_B_7EOlVDn41_2));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(w_dff_B_EVtxD5999_2));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(w_dff_B_5pO8copD6_2));
	jspl jspl_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.din(n967));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(w_dff_B_uWR791Wt7_2));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(w_dff_B_wCp8FuyK2_2));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n980_0(.douta(w_dff_A_5ImTVvdP6_0),.doutb(w_n980_0[1]),.din(w_dff_B_cde1KABN0_2));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(w_dff_B_PNRnO2Eg7_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(w_dff_B_drOzPVID4_2));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_biMF5xiY2_2));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(n988));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(n990));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(n996));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(n1004));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_ifldbHus3_1),.din(n1006));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1017_0(.douta(w_dff_A_gqHF4DZl2_0),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_ZG439JIz6_2));
	jspl jspl_w_n1022_0(.douta(w_dff_A_dJHV3D2E4_0),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(w_dff_B_WGkBMv0o2_2));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_kvmSRX9U9_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(w_dff_B_FeoLRdE16_2));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.din(w_dff_B_i0Ted2BP2_2));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(w_dff_B_vzjEJ0329_2));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(w_dff_B_H8LlxpHs5_2));
	jspl jspl_w_n1051_0(.douta(w_n1051_0[0]),.doutb(w_n1051_0[1]),.din(n1051));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(w_dff_B_SU75RpGS3_2));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.din(w_dff_B_ZFYsJInP3_2));
	jspl jspl_w_n1061_0(.douta(w_n1061_0[0]),.doutb(w_n1061_0[1]),.din(n1061));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(w_dff_B_0BghZfKE4_2));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(w_dff_B_pMPuw8w75_2));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(w_dff_B_1Wo4CiF30_2));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(w_dff_B_HQl7EJU00_2));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(w_dff_B_SSM5SvsX8_2));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(w_dff_B_5RHH1Fax3_2));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(w_dff_B_YzE7vhIp1_2));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(n1089));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(n1091));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(n1093));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(n1095));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1098_0(.douta(w_n1098_0[0]),.doutb(w_n1098_0[1]),.din(n1098));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.din(n1100));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(n1101));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(n1103));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.din(n1106));
	jspl jspl_w_n1107_0(.douta(w_n1107_0[0]),.doutb(w_n1107_0[1]),.din(n1107));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_n1108_0[1]),.din(n1108));
	jspl jspl_w_n1109_0(.douta(w_dff_A_eim6TkIP3_0),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1119_0(.douta(w_dff_A_V7rxrfus7_0),.doutb(w_n1119_0[1]),.din(w_dff_B_5qk6RfLR5_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(w_dff_B_IcVXHOmB8_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(w_dff_B_hFHKLx7N3_2));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(w_dff_B_LE4azKlA7_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.din(w_dff_B_DuRkClK69_2));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(w_dff_B_jgJwiJ2Q9_2));
	jspl jspl_w_n1144_0(.douta(w_n1144_0[0]),.doutb(w_n1144_0[1]),.din(n1144));
	jspl jspl_w_n1146_0(.douta(w_n1146_0[0]),.doutb(w_n1146_0[1]),.din(w_dff_B_tZNJFONl2_2));
	jspl jspl_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.din(n1149));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(w_dff_B_Sr08VwJO8_2));
	jspl jspl_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.din(n1154));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(w_dff_B_aPtSe8m90_2));
	jspl jspl_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(w_dff_B_SbRg2T466_2));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(w_dff_B_SVEDSDEi2_2));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(w_dff_B_3LF1fFik5_2));
	jspl jspl_w_n1174_0(.douta(w_n1174_0[0]),.doutb(w_n1174_0[1]),.din(n1174));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(w_dff_B_ec9y6jOn3_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(w_dff_B_1YbWHAfd8_2));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1182_0(.douta(w_n1182_0[0]),.doutb(w_n1182_0[1]),.din(w_dff_B_KpCmnpil7_2));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(w_dff_B_B4HWDCRE2_2));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.din(n1187));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(n1188));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(n1190));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(n1192));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl jspl_w_n1194_0(.douta(w_n1194_0[0]),.doutb(w_n1194_0[1]),.din(n1194));
	jspl jspl_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.din(n1195));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1199_0(.douta(w_n1199_0[0]),.doutb(w_n1199_0[1]),.din(n1199));
	jspl jspl_w_n1200_0(.douta(w_n1200_0[0]),.doutb(w_n1200_0[1]),.din(n1200));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(n1203));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1207_0(.douta(w_dff_A_BPfeRMEG5_0),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_ovoLQTwy0_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(w_dff_B_9iVFdk5t0_2));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(w_dff_B_aNHEh6ZZ6_2));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(w_dff_B_p41h6Qti7_2));
	jspl jspl_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.din(n1235));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(w_dff_B_NAXPIAqq6_2));
	jspl jspl_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.din(n1240));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(w_dff_B_pzaxuUlC1_2));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(w_dff_B_xdbSe9VM5_2));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(w_dff_B_wmuiS3qd6_2));
	jspl jspl_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.din(n1255));
	jspl jspl_w_n1257_0(.douta(w_n1257_0[0]),.doutb(w_n1257_0[1]),.din(w_dff_B_cUJKJhQb6_2));
	jspl jspl_w_n1260_0(.douta(w_n1260_0[0]),.doutb(w_n1260_0[1]),.din(n1260));
	jspl jspl_w_n1262_0(.douta(w_n1262_0[0]),.doutb(w_n1262_0[1]),.din(w_dff_B_p0tOgi460_2));
	jspl jspl_w_n1265_0(.douta(w_n1265_0[0]),.doutb(w_n1265_0[1]),.din(n1265));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(w_dff_B_HO6FzM4K1_2));
	jspl jspl_w_n1267_0(.douta(w_n1267_0[0]),.doutb(w_n1267_0[1]),.din(w_dff_B_rVQEiO3x4_2));
	jspl jspl_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.din(n1270));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(n1273));
	jspl jspl_w_n1274_0(.douta(w_n1274_0[0]),.doutb(w_n1274_0[1]),.din(n1274));
	jspl jspl_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.din(w_dff_B_le5ggeC59_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1277_0(.douta(w_n1277_0[0]),.doutb(w_n1277_0[1]),.din(n1277));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(n1279));
	jspl jspl_w_n1280_0(.douta(w_n1280_0[0]),.doutb(w_n1280_0[1]),.din(n1280));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(n1281));
	jspl jspl_w_n1282_0(.douta(w_n1282_0[0]),.doutb(w_n1282_0[1]),.din(n1282));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1284_0(.douta(w_n1284_0[0]),.doutb(w_n1284_0[1]),.din(n1284));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(n1285));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1287_0(.douta(w_n1287_0[0]),.doutb(w_n1287_0[1]),.din(n1287));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1289_0(.douta(w_n1289_0[0]),.doutb(w_n1289_0[1]),.din(n1289));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_dff_A_XyCh9jAo8_1),.din(n1294));
	jspl jspl_w_n1295_0(.douta(w_dff_A_SX75LK7v5_0),.doutb(w_n1295_0[1]),.din(n1295));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(w_dff_B_pxiAqJRP4_2));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(w_dff_B_khNyTxgR1_2));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_Mmu3qViy6_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(w_dff_B_NV8HOxjN1_2));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(w_dff_B_8I3X7dEL7_2));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1327_0(.douta(w_n1327_0[0]),.doutb(w_n1327_0[1]),.din(w_dff_B_RmbCiMPF6_2));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(w_dff_B_x2InN0J80_2));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(w_dff_B_TeMjtAcZ2_2));
	jspl jspl_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(w_dff_B_ICXqUIyS3_2));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.din(w_dff_B_QZg7MbcJ4_2));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(w_dff_B_P6NmMIMJ3_2));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(w_dff_B_RapIJeDF9_2));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(w_dff_B_WYj5ns8X9_2));
	jspl jspl_w_n1355_0(.douta(w_n1355_0[0]),.doutb(w_n1355_0[1]),.din(n1355));
	jspl jspl_w_n1357_0(.douta(w_n1357_0[0]),.doutb(w_n1357_0[1]),.din(n1357));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.din(n1360));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(n1362));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(n1364));
	jspl jspl_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.din(n1365));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(n1366));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(n1368));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_n1370_0[1]),.din(n1370));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.din(n1374));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_dff_A_cFG0Ia5Z3_1),.din(n1379));
	jspl jspl_w_n1384_0(.douta(w_n1384_0[0]),.doutb(w_n1384_0[1]),.din(n1384));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(w_dff_B_X5KheESI6_2));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(w_dff_B_PX4TXQFr3_2));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_dff_A_cnLtIaDT5_1),.din(n1393));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_YozbgheA4_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(w_dff_B_teb3lBS75_2));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(w_dff_B_zVqLTIM78_2));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(w_dff_B_ISmDjF5k2_2));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(w_dff_B_epbHyQ9n1_2));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(w_dff_B_LfDwkVxA7_2));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(w_dff_B_EbO6FDzF9_2));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(w_dff_B_ArqXoQLF0_2));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(w_dff_B_DBt030OO6_2));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(w_dff_B_LU4nYTi48_2));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_0BpSd3x59_2));
	jspl jspl_w_n1423_0(.douta(w_n1423_0[0]),.doutb(w_n1423_0[1]),.din(w_dff_B_3ylLCC6d3_2));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(w_dff_B_m2NcjGE91_2));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(w_dff_B_KiPv2Y083_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(w_dff_B_NZ65v4E38_2));
	jspl jspl_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.din(w_dff_B_UX6p194Y7_2));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.din(n1437));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.din(n1438));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(n1440));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.din(n1442));
	jspl jspl_w_n1443_0(.douta(w_n1443_0[0]),.doutb(w_n1443_0[1]),.din(n1443));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1448_0(.douta(w_n1448_0[0]),.doutb(w_n1448_0[1]),.din(n1448));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1450_0(.douta(w_n1450_0[0]),.doutb(w_n1450_0[1]),.din(n1450));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1455_0(.douta(w_n1455_0[0]),.doutb(w_dff_A_1RrEBp7h4_1),.din(n1455));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(w_dff_B_w0qqjdMw7_2));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(w_dff_B_3uOXTrKJ1_2));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_dff_A_CXO8gbcQ6_1),.din(n1469));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(w_dff_B_vNogexnc8_2));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(w_dff_B_dmovVPEO7_2));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(w_dff_B_MDqnxK5G5_2));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(w_dff_B_zyA9jFjr4_2));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(w_dff_B_meCKv3YC1_2));
	jspl jspl_w_n1484_0(.douta(w_n1484_0[0]),.doutb(w_n1484_0[1]),.din(w_dff_B_yYSeLr7z7_2));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(w_dff_B_4I6PdJS70_2));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(w_dff_B_9jxM2aiy2_2));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(w_dff_B_7bG69QOm0_2));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(w_dff_B_E7UOXUYz1_2));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_srWxmUGH1_2));
	jspl jspl_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.din(w_dff_B_BdadzOvs7_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(w_dff_B_GvYE6x427_2));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_n1501_0[1]),.din(w_dff_B_iQjh87NT6_2));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(n1513));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(n1515));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(n1517));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1519_0(.douta(w_n1519_0[0]),.doutb(w_n1519_0[1]),.din(n1519));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_dff_A_Q4KL71pY0_1),.din(n1524));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(w_dff_B_WFe17quy4_2));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(w_dff_B_9XTlHHFv3_2));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_dff_A_v4JB5FpV2_1),.din(n1538));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(w_dff_B_x51BuWjL3_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(w_dff_B_O0h7KmFr2_2));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(w_dff_B_bx6MHFYJ5_2));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(w_dff_B_5R5a4ZnB0_2));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(w_dff_B_00rP6kOR2_2));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_moEMgU2N6_2));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(w_dff_B_jJSpxOIK5_2));
	jspl jspl_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.din(w_dff_B_CDoZxnYN5_2));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(w_dff_B_3is5bFk90_2));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(w_dff_B_Tq1QvZat2_2));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(w_dff_B_SMT7j2uL7_2));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(w_dff_B_eNP0hdtM1_2));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.din(n1568));
	jspl jspl_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.din(n1570));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1572_0(.douta(w_n1572_0[0]),.doutb(w_n1572_0[1]),.din(n1572));
	jspl jspl_w_n1573_0(.douta(w_n1573_0[0]),.doutb(w_n1573_0[1]),.din(n1573));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(n1576));
	jspl jspl_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.din(n1577));
	jspl jspl_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.din(n1578));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(n1579));
	jspl jspl_w_n1580_0(.douta(w_n1580_0[0]),.doutb(w_n1580_0[1]),.din(n1580));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(n1581));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl jspl_w_n1585_0(.douta(w_n1585_0[0]),.doutb(w_n1585_0[1]),.din(n1585));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_dff_A_2W8eSvNS9_1),.din(n1586));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(w_dff_B_lFsWGR3P7_2));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(w_dff_B_TtcXziLy1_2));
	jspl jspl_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_dff_A_6pYNKldV8_1),.din(n1600));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(w_dff_B_wbcx4oOg9_2));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(w_dff_B_Jm07S3Nn1_2));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(w_dff_B_KzaSQKeX0_2));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(w_dff_B_6C8Bv70R4_2));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(w_dff_B_2HGFSGuf0_2));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(w_dff_B_SGwdY6Qc1_2));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_n1617_0[1]),.din(w_dff_B_NpD8YZJA9_2));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(w_dff_B_dfw6ZqK21_2));
	jspl jspl_w_n1621_0(.douta(w_n1621_0[0]),.doutb(w_n1621_0[1]),.din(w_dff_B_1PFggV3Q2_2));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(w_dff_B_gw1iOXXp7_2));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(n1628));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1630_0(.douta(w_n1630_0[0]),.doutb(w_n1630_0[1]),.din(n1630));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(n1636));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_dff_A_my0cukNQ9_1),.din(n1641));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_xnQZKn1e6_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_9b7f8n6n3_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(w_dff_B_ezdYGMnN4_2));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(w_dff_B_dAEQBR6J5_2));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(w_dff_B_b59aqmGd7_2));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(w_dff_B_dT6I9ojo5_2));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(w_dff_B_SwtKcqr72_2));
	jspl jspl_w_n1668_0(.douta(w_n1668_0[0]),.doutb(w_n1668_0[1]),.din(w_dff_B_hapB8zjH4_2));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(w_dff_B_r3huhRxb0_2));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(w_dff_B_oOKqRdP05_2));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(w_dff_B_FpLZbDWC4_2));
	jspl jspl_w_n1676_0(.douta(w_n1676_0[0]),.doutb(w_n1676_0[1]),.din(n1676));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.din(n1681));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl jspl_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.din(n1683));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1686_0(.douta(w_n1686_0[0]),.doutb(w_n1686_0[1]),.din(n1686));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_dff_A_ixcFa8oL9_1),.din(n1689));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_dff_A_csoi6cFm2_1),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_rpETgB5D8_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_8F3sj5hl8_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_0kbzAFr32_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(w_dff_B_jnITGK5r1_2));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(w_dff_B_ng7MdjRo8_2));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(w_dff_B_FwikrSQf0_2));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(w_dff_B_5MEgAAAv1_2));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(w_dff_B_J7N8fnvp0_2));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.din(n1721));
	jspl jspl_w_n1722_0(.douta(w_n1722_0[0]),.doutb(w_n1722_0[1]),.din(n1722));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_dff_A_nw0zklZx2_1),.din(n1727));
	jspl jspl_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.din(n1734));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_dff_A_3cdlYTgW1_1),.din(n1737));
	jspl jspl_w_n1739_0(.douta(w_n1739_0[0]),.doutb(w_n1739_0[1]),.din(w_dff_B_Nsr8LsGd2_2));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(w_dff_B_9jwiKTXR0_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_esALD8hJ7_2));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(w_dff_B_uKa30N7n8_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(w_dff_B_ooyi4Dhj8_2));
	jspl jspl_w_n1749_0(.douta(w_n1749_0[0]),.doutb(w_n1749_0[1]),.din(w_dff_B_yP0NFXiX9_2));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_dff_A_wwb1llDO5_1),.din(n1760));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_dff_A_KNttCfjm4_1),.din(n1770));
	jspl jspl_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.din(w_dff_B_Dj7xdSpz2_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_QmpOAylZ8_2));
	jspl jspl_w_n1776_0(.douta(w_n1776_0[0]),.doutb(w_n1776_0[1]),.din(w_dff_B_N7U1sZEN0_2));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(w_dff_B_NcT0JcZ80_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.din(n1782));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.din(n1784));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_dff_A_dLavTA406_1),.din(n1786));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_dff_A_KzNFY41T9_1),.din(n1796));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(w_dff_B_MVv0CSar4_2));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(w_dff_B_yB2mG7uE0_2));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_dff_A_7HgF2Ebz3_1),.din(n1805));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_CaMxzjt13_2));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1818_0(.douta(w_dff_A_Xwkf2BHt1_0),.doutb(w_n1818_0[1]),.din(n1818));
	jdff dff_B_6HCBISXv8_0(.din(n73),.dout(w_dff_B_6HCBISXv8_0),.clk(gclk));
	jdff dff_B_44QAozby7_0(.din(n72),.dout(w_dff_B_44QAozby7_0),.clk(gclk));
	jdff dff_B_P1ly3IOS3_1(.din(n76),.dout(w_dff_B_P1ly3IOS3_1),.clk(gclk));
	jdff dff_B_ffyvxpWQ4_1(.din(w_dff_B_P1ly3IOS3_1),.dout(w_dff_B_ffyvxpWQ4_1),.clk(gclk));
	jdff dff_B_AC3vnYzm4_1(.din(n87),.dout(w_dff_B_AC3vnYzm4_1),.clk(gclk));
	jdff dff_B_ZHAJKBDS4_1(.din(w_dff_B_AC3vnYzm4_1),.dout(w_dff_B_ZHAJKBDS4_1),.clk(gclk));
	jdff dff_B_APaSBmRP6_1(.din(w_dff_B_ZHAJKBDS4_1),.dout(w_dff_B_APaSBmRP6_1),.clk(gclk));
	jdff dff_B_JZA2Vr1t8_1(.din(w_dff_B_APaSBmRP6_1),.dout(w_dff_B_JZA2Vr1t8_1),.clk(gclk));
	jdff dff_B_2Fxuiwdr8_1(.din(n107),.dout(w_dff_B_2Fxuiwdr8_1),.clk(gclk));
	jdff dff_B_3FPIijzO9_1(.din(w_dff_B_2Fxuiwdr8_1),.dout(w_dff_B_3FPIijzO9_1),.clk(gclk));
	jdff dff_B_AQulzuKa3_1(.din(w_dff_B_3FPIijzO9_1),.dout(w_dff_B_AQulzuKa3_1),.clk(gclk));
	jdff dff_B_oRWhJ7ji7_1(.din(w_dff_B_AQulzuKa3_1),.dout(w_dff_B_oRWhJ7ji7_1),.clk(gclk));
	jdff dff_B_M3ZkKUfG3_1(.din(w_dff_B_oRWhJ7ji7_1),.dout(w_dff_B_M3ZkKUfG3_1),.clk(gclk));
	jdff dff_B_RzOqDIa92_1(.din(w_dff_B_M3ZkKUfG3_1),.dout(w_dff_B_RzOqDIa92_1),.clk(gclk));
	jdff dff_B_GiElhWcy4_1(.din(w_dff_B_RzOqDIa92_1),.dout(w_dff_B_GiElhWcy4_1),.clk(gclk));
	jdff dff_B_6lI0U1M62_1(.din(w_dff_B_GiElhWcy4_1),.dout(w_dff_B_6lI0U1M62_1),.clk(gclk));
	jdff dff_B_ZXRMAWNp2_1(.din(n136),.dout(w_dff_B_ZXRMAWNp2_1),.clk(gclk));
	jdff dff_B_2h8wkNxg6_1(.din(w_dff_B_ZXRMAWNp2_1),.dout(w_dff_B_2h8wkNxg6_1),.clk(gclk));
	jdff dff_B_RGGz8Q9K9_1(.din(w_dff_B_2h8wkNxg6_1),.dout(w_dff_B_RGGz8Q9K9_1),.clk(gclk));
	jdff dff_B_EhBSwQtR6_1(.din(w_dff_B_RGGz8Q9K9_1),.dout(w_dff_B_EhBSwQtR6_1),.clk(gclk));
	jdff dff_B_Zs2CFwyA2_1(.din(w_dff_B_EhBSwQtR6_1),.dout(w_dff_B_Zs2CFwyA2_1),.clk(gclk));
	jdff dff_B_osBIpEl50_1(.din(w_dff_B_Zs2CFwyA2_1),.dout(w_dff_B_osBIpEl50_1),.clk(gclk));
	jdff dff_B_p1KD1ZgB9_1(.din(w_dff_B_osBIpEl50_1),.dout(w_dff_B_p1KD1ZgB9_1),.clk(gclk));
	jdff dff_B_b5hrTdYE4_1(.din(w_dff_B_p1KD1ZgB9_1),.dout(w_dff_B_b5hrTdYE4_1),.clk(gclk));
	jdff dff_B_SPQ4uKhJ9_1(.din(w_dff_B_b5hrTdYE4_1),.dout(w_dff_B_SPQ4uKhJ9_1),.clk(gclk));
	jdff dff_B_2NBSrRwF8_1(.din(w_dff_B_SPQ4uKhJ9_1),.dout(w_dff_B_2NBSrRwF8_1),.clk(gclk));
	jdff dff_B_9MUDVhOy3_1(.din(n171),.dout(w_dff_B_9MUDVhOy3_1),.clk(gclk));
	jdff dff_B_rY0cHKBA7_1(.din(w_dff_B_9MUDVhOy3_1),.dout(w_dff_B_rY0cHKBA7_1),.clk(gclk));
	jdff dff_B_zezWY9qf2_1(.din(w_dff_B_rY0cHKBA7_1),.dout(w_dff_B_zezWY9qf2_1),.clk(gclk));
	jdff dff_B_r6ZX9DFu5_1(.din(w_dff_B_zezWY9qf2_1),.dout(w_dff_B_r6ZX9DFu5_1),.clk(gclk));
	jdff dff_B_QN7GF7U64_1(.din(w_dff_B_r6ZX9DFu5_1),.dout(w_dff_B_QN7GF7U64_1),.clk(gclk));
	jdff dff_B_9tLIY7T60_1(.din(w_dff_B_QN7GF7U64_1),.dout(w_dff_B_9tLIY7T60_1),.clk(gclk));
	jdff dff_B_47zio2a76_1(.din(w_dff_B_9tLIY7T60_1),.dout(w_dff_B_47zio2a76_1),.clk(gclk));
	jdff dff_B_5y1P21MO3_1(.din(w_dff_B_47zio2a76_1),.dout(w_dff_B_5y1P21MO3_1),.clk(gclk));
	jdff dff_B_UmJB9HqK5_1(.din(w_dff_B_5y1P21MO3_1),.dout(w_dff_B_UmJB9HqK5_1),.clk(gclk));
	jdff dff_B_2gQWOTyL9_1(.din(w_dff_B_UmJB9HqK5_1),.dout(w_dff_B_2gQWOTyL9_1),.clk(gclk));
	jdff dff_B_WYZafbxU0_1(.din(w_dff_B_2gQWOTyL9_1),.dout(w_dff_B_WYZafbxU0_1),.clk(gclk));
	jdff dff_B_KLFHqAdj5_1(.din(w_dff_B_WYZafbxU0_1),.dout(w_dff_B_KLFHqAdj5_1),.clk(gclk));
	jdff dff_B_mlpGvvNC4_1(.din(n213),.dout(w_dff_B_mlpGvvNC4_1),.clk(gclk));
	jdff dff_B_WTsUlwhd5_1(.din(w_dff_B_mlpGvvNC4_1),.dout(w_dff_B_WTsUlwhd5_1),.clk(gclk));
	jdff dff_B_G3Hg9CTa0_1(.din(w_dff_B_WTsUlwhd5_1),.dout(w_dff_B_G3Hg9CTa0_1),.clk(gclk));
	jdff dff_B_1rPq1ELK7_1(.din(w_dff_B_G3Hg9CTa0_1),.dout(w_dff_B_1rPq1ELK7_1),.clk(gclk));
	jdff dff_B_bhhnoe417_1(.din(w_dff_B_1rPq1ELK7_1),.dout(w_dff_B_bhhnoe417_1),.clk(gclk));
	jdff dff_B_GsgtfQa27_1(.din(w_dff_B_bhhnoe417_1),.dout(w_dff_B_GsgtfQa27_1),.clk(gclk));
	jdff dff_B_bOxjIvyv2_1(.din(w_dff_B_GsgtfQa27_1),.dout(w_dff_B_bOxjIvyv2_1),.clk(gclk));
	jdff dff_B_zaENAgzd0_1(.din(w_dff_B_bOxjIvyv2_1),.dout(w_dff_B_zaENAgzd0_1),.clk(gclk));
	jdff dff_B_ZKOk38e58_1(.din(w_dff_B_zaENAgzd0_1),.dout(w_dff_B_ZKOk38e58_1),.clk(gclk));
	jdff dff_B_ZRCXMTqp0_1(.din(w_dff_B_ZKOk38e58_1),.dout(w_dff_B_ZRCXMTqp0_1),.clk(gclk));
	jdff dff_B_K0iH9oca7_1(.din(w_dff_B_ZRCXMTqp0_1),.dout(w_dff_B_K0iH9oca7_1),.clk(gclk));
	jdff dff_B_Pn7KYAtS2_1(.din(w_dff_B_K0iH9oca7_1),.dout(w_dff_B_Pn7KYAtS2_1),.clk(gclk));
	jdff dff_B_GvS6AMBC3_1(.din(w_dff_B_Pn7KYAtS2_1),.dout(w_dff_B_GvS6AMBC3_1),.clk(gclk));
	jdff dff_B_Fd6u6okS6_1(.din(w_dff_B_GvS6AMBC3_1),.dout(w_dff_B_Fd6u6okS6_1),.clk(gclk));
	jdff dff_B_dHxcuFZv5_1(.din(n262),.dout(w_dff_B_dHxcuFZv5_1),.clk(gclk));
	jdff dff_B_eXbxvIVK6_1(.din(w_dff_B_dHxcuFZv5_1),.dout(w_dff_B_eXbxvIVK6_1),.clk(gclk));
	jdff dff_B_73mwioK95_1(.din(w_dff_B_eXbxvIVK6_1),.dout(w_dff_B_73mwioK95_1),.clk(gclk));
	jdff dff_B_gkZRwCpI8_1(.din(w_dff_B_73mwioK95_1),.dout(w_dff_B_gkZRwCpI8_1),.clk(gclk));
	jdff dff_B_PfcsKGKn9_1(.din(w_dff_B_gkZRwCpI8_1),.dout(w_dff_B_PfcsKGKn9_1),.clk(gclk));
	jdff dff_B_wANkVgu04_1(.din(w_dff_B_PfcsKGKn9_1),.dout(w_dff_B_wANkVgu04_1),.clk(gclk));
	jdff dff_B_SICmrVRM4_1(.din(w_dff_B_wANkVgu04_1),.dout(w_dff_B_SICmrVRM4_1),.clk(gclk));
	jdff dff_B_WZmPXDDu0_1(.din(w_dff_B_SICmrVRM4_1),.dout(w_dff_B_WZmPXDDu0_1),.clk(gclk));
	jdff dff_B_weYljKq51_1(.din(w_dff_B_WZmPXDDu0_1),.dout(w_dff_B_weYljKq51_1),.clk(gclk));
	jdff dff_B_R6wPNhWs6_1(.din(w_dff_B_weYljKq51_1),.dout(w_dff_B_R6wPNhWs6_1),.clk(gclk));
	jdff dff_B_e17I3Z3T3_1(.din(w_dff_B_R6wPNhWs6_1),.dout(w_dff_B_e17I3Z3T3_1),.clk(gclk));
	jdff dff_B_OYyNmgz28_1(.din(w_dff_B_e17I3Z3T3_1),.dout(w_dff_B_OYyNmgz28_1),.clk(gclk));
	jdff dff_B_wpT0izjM6_1(.din(w_dff_B_OYyNmgz28_1),.dout(w_dff_B_wpT0izjM6_1),.clk(gclk));
	jdff dff_B_NDCYA0pf8_1(.din(w_dff_B_wpT0izjM6_1),.dout(w_dff_B_NDCYA0pf8_1),.clk(gclk));
	jdff dff_B_vBSXl2Xc4_1(.din(w_dff_B_NDCYA0pf8_1),.dout(w_dff_B_vBSXl2Xc4_1),.clk(gclk));
	jdff dff_B_MoG9tggT5_1(.din(w_dff_B_vBSXl2Xc4_1),.dout(w_dff_B_MoG9tggT5_1),.clk(gclk));
	jdff dff_B_lER1JFTz8_1(.din(n318),.dout(w_dff_B_lER1JFTz8_1),.clk(gclk));
	jdff dff_B_v8rZBzxZ9_1(.din(w_dff_B_lER1JFTz8_1),.dout(w_dff_B_v8rZBzxZ9_1),.clk(gclk));
	jdff dff_B_rA12eeMp6_1(.din(w_dff_B_v8rZBzxZ9_1),.dout(w_dff_B_rA12eeMp6_1),.clk(gclk));
	jdff dff_B_337ugziS5_1(.din(w_dff_B_rA12eeMp6_1),.dout(w_dff_B_337ugziS5_1),.clk(gclk));
	jdff dff_B_GI4gaQTH8_1(.din(w_dff_B_337ugziS5_1),.dout(w_dff_B_GI4gaQTH8_1),.clk(gclk));
	jdff dff_B_EsH4uZ5d2_1(.din(w_dff_B_GI4gaQTH8_1),.dout(w_dff_B_EsH4uZ5d2_1),.clk(gclk));
	jdff dff_B_ionqlwBo7_1(.din(w_dff_B_EsH4uZ5d2_1),.dout(w_dff_B_ionqlwBo7_1),.clk(gclk));
	jdff dff_B_1lfLFahR2_1(.din(w_dff_B_ionqlwBo7_1),.dout(w_dff_B_1lfLFahR2_1),.clk(gclk));
	jdff dff_B_fAbvQ5Lh1_1(.din(w_dff_B_1lfLFahR2_1),.dout(w_dff_B_fAbvQ5Lh1_1),.clk(gclk));
	jdff dff_B_H1AJWwLO1_1(.din(w_dff_B_fAbvQ5Lh1_1),.dout(w_dff_B_H1AJWwLO1_1),.clk(gclk));
	jdff dff_B_f0bdwSEM7_1(.din(w_dff_B_H1AJWwLO1_1),.dout(w_dff_B_f0bdwSEM7_1),.clk(gclk));
	jdff dff_B_gcplfyCN8_1(.din(w_dff_B_f0bdwSEM7_1),.dout(w_dff_B_gcplfyCN8_1),.clk(gclk));
	jdff dff_B_slpYj5Sz2_1(.din(w_dff_B_gcplfyCN8_1),.dout(w_dff_B_slpYj5Sz2_1),.clk(gclk));
	jdff dff_B_WAgK0wi61_1(.din(w_dff_B_slpYj5Sz2_1),.dout(w_dff_B_WAgK0wi61_1),.clk(gclk));
	jdff dff_B_E2fepEw78_1(.din(w_dff_B_WAgK0wi61_1),.dout(w_dff_B_E2fepEw78_1),.clk(gclk));
	jdff dff_B_KAaoo34K5_1(.din(w_dff_B_E2fepEw78_1),.dout(w_dff_B_KAaoo34K5_1),.clk(gclk));
	jdff dff_B_h0pK2ZN59_1(.din(w_dff_B_KAaoo34K5_1),.dout(w_dff_B_h0pK2ZN59_1),.clk(gclk));
	jdff dff_B_Vq2eGezB9_1(.din(w_dff_B_h0pK2ZN59_1),.dout(w_dff_B_Vq2eGezB9_1),.clk(gclk));
	jdff dff_B_eJBhluQ05_1(.din(n381),.dout(w_dff_B_eJBhluQ05_1),.clk(gclk));
	jdff dff_B_db6P1TxI9_1(.din(w_dff_B_eJBhluQ05_1),.dout(w_dff_B_db6P1TxI9_1),.clk(gclk));
	jdff dff_B_z7sfF18P0_1(.din(w_dff_B_db6P1TxI9_1),.dout(w_dff_B_z7sfF18P0_1),.clk(gclk));
	jdff dff_B_r2WbuOzk7_1(.din(w_dff_B_z7sfF18P0_1),.dout(w_dff_B_r2WbuOzk7_1),.clk(gclk));
	jdff dff_B_Vw3ANMGR6_1(.din(w_dff_B_r2WbuOzk7_1),.dout(w_dff_B_Vw3ANMGR6_1),.clk(gclk));
	jdff dff_B_zIVdlYjI4_1(.din(w_dff_B_Vw3ANMGR6_1),.dout(w_dff_B_zIVdlYjI4_1),.clk(gclk));
	jdff dff_B_piUAakqS0_1(.din(w_dff_B_zIVdlYjI4_1),.dout(w_dff_B_piUAakqS0_1),.clk(gclk));
	jdff dff_B_eNk1BIck3_1(.din(w_dff_B_piUAakqS0_1),.dout(w_dff_B_eNk1BIck3_1),.clk(gclk));
	jdff dff_B_kZVeK0vh5_1(.din(w_dff_B_eNk1BIck3_1),.dout(w_dff_B_kZVeK0vh5_1),.clk(gclk));
	jdff dff_B_To86uOx91_1(.din(w_dff_B_kZVeK0vh5_1),.dout(w_dff_B_To86uOx91_1),.clk(gclk));
	jdff dff_B_hikmQHZC1_1(.din(w_dff_B_To86uOx91_1),.dout(w_dff_B_hikmQHZC1_1),.clk(gclk));
	jdff dff_B_xN1NM4QN6_1(.din(w_dff_B_hikmQHZC1_1),.dout(w_dff_B_xN1NM4QN6_1),.clk(gclk));
	jdff dff_B_4t2gradw0_1(.din(w_dff_B_xN1NM4QN6_1),.dout(w_dff_B_4t2gradw0_1),.clk(gclk));
	jdff dff_B_Mswpm0uw4_1(.din(w_dff_B_4t2gradw0_1),.dout(w_dff_B_Mswpm0uw4_1),.clk(gclk));
	jdff dff_B_eJhFKHUS2_1(.din(w_dff_B_Mswpm0uw4_1),.dout(w_dff_B_eJhFKHUS2_1),.clk(gclk));
	jdff dff_B_nwUufPEM4_1(.din(w_dff_B_eJhFKHUS2_1),.dout(w_dff_B_nwUufPEM4_1),.clk(gclk));
	jdff dff_B_CwUH8hIa5_1(.din(w_dff_B_nwUufPEM4_1),.dout(w_dff_B_CwUH8hIa5_1),.clk(gclk));
	jdff dff_B_XEwaOo484_1(.din(w_dff_B_CwUH8hIa5_1),.dout(w_dff_B_XEwaOo484_1),.clk(gclk));
	jdff dff_B_s2M3ZHh94_1(.din(w_dff_B_XEwaOo484_1),.dout(w_dff_B_s2M3ZHh94_1),.clk(gclk));
	jdff dff_B_fk9C74SQ8_1(.din(w_dff_B_s2M3ZHh94_1),.dout(w_dff_B_fk9C74SQ8_1),.clk(gclk));
	jdff dff_B_sGQo05QB3_1(.din(w_dff_B_fk9C74SQ8_1),.dout(w_dff_B_sGQo05QB3_1),.clk(gclk));
	jdff dff_B_jQt9tUQQ3_1(.din(w_dff_B_sGQo05QB3_1),.dout(w_dff_B_jQt9tUQQ3_1),.clk(gclk));
	jdff dff_B_75UviKYP7_1(.din(w_dff_B_jQt9tUQQ3_1),.dout(w_dff_B_75UviKYP7_1),.clk(gclk));
	jdff dff_B_fNAOjXgj7_1(.din(n452),.dout(w_dff_B_fNAOjXgj7_1),.clk(gclk));
	jdff dff_B_yOZ9FPuE0_1(.din(w_dff_B_fNAOjXgj7_1),.dout(w_dff_B_yOZ9FPuE0_1),.clk(gclk));
	jdff dff_B_DcOGLGC31_1(.din(w_dff_B_yOZ9FPuE0_1),.dout(w_dff_B_DcOGLGC31_1),.clk(gclk));
	jdff dff_B_Kvv5XlAD3_1(.din(w_dff_B_DcOGLGC31_1),.dout(w_dff_B_Kvv5XlAD3_1),.clk(gclk));
	jdff dff_B_RqZ8sDuB7_1(.din(w_dff_B_Kvv5XlAD3_1),.dout(w_dff_B_RqZ8sDuB7_1),.clk(gclk));
	jdff dff_B_6dW1A9a36_1(.din(w_dff_B_RqZ8sDuB7_1),.dout(w_dff_B_6dW1A9a36_1),.clk(gclk));
	jdff dff_B_dtvNKsfH7_1(.din(w_dff_B_6dW1A9a36_1),.dout(w_dff_B_dtvNKsfH7_1),.clk(gclk));
	jdff dff_B_fAThyMH45_1(.din(w_dff_B_dtvNKsfH7_1),.dout(w_dff_B_fAThyMH45_1),.clk(gclk));
	jdff dff_B_J1kGCNu40_1(.din(w_dff_B_fAThyMH45_1),.dout(w_dff_B_J1kGCNu40_1),.clk(gclk));
	jdff dff_B_jsxvJsVY9_1(.din(w_dff_B_J1kGCNu40_1),.dout(w_dff_B_jsxvJsVY9_1),.clk(gclk));
	jdff dff_B_2JFBsbtW8_1(.din(w_dff_B_jsxvJsVY9_1),.dout(w_dff_B_2JFBsbtW8_1),.clk(gclk));
	jdff dff_B_lUcAy4X63_1(.din(w_dff_B_2JFBsbtW8_1),.dout(w_dff_B_lUcAy4X63_1),.clk(gclk));
	jdff dff_B_pNShPGpz0_1(.din(w_dff_B_lUcAy4X63_1),.dout(w_dff_B_pNShPGpz0_1),.clk(gclk));
	jdff dff_B_0uDtAaaq6_1(.din(w_dff_B_pNShPGpz0_1),.dout(w_dff_B_0uDtAaaq6_1),.clk(gclk));
	jdff dff_B_1bVWCKcC6_1(.din(w_dff_B_0uDtAaaq6_1),.dout(w_dff_B_1bVWCKcC6_1),.clk(gclk));
	jdff dff_B_NJIlRyTE6_1(.din(w_dff_B_1bVWCKcC6_1),.dout(w_dff_B_NJIlRyTE6_1),.clk(gclk));
	jdff dff_B_jwipN2CY1_1(.din(w_dff_B_NJIlRyTE6_1),.dout(w_dff_B_jwipN2CY1_1),.clk(gclk));
	jdff dff_B_2kZXeCC49_1(.din(w_dff_B_jwipN2CY1_1),.dout(w_dff_B_2kZXeCC49_1),.clk(gclk));
	jdff dff_B_Aw8akPT04_1(.din(w_dff_B_2kZXeCC49_1),.dout(w_dff_B_Aw8akPT04_1),.clk(gclk));
	jdff dff_B_u3x12r8n9_1(.din(w_dff_B_Aw8akPT04_1),.dout(w_dff_B_u3x12r8n9_1),.clk(gclk));
	jdff dff_B_gouTXm9C8_1(.din(w_dff_B_u3x12r8n9_1),.dout(w_dff_B_gouTXm9C8_1),.clk(gclk));
	jdff dff_B_LOadvB4t1_1(.din(w_dff_B_gouTXm9C8_1),.dout(w_dff_B_LOadvB4t1_1),.clk(gclk));
	jdff dff_B_kWE5Tpjh0_1(.din(w_dff_B_LOadvB4t1_1),.dout(w_dff_B_kWE5Tpjh0_1),.clk(gclk));
	jdff dff_B_XAOBa3Mx5_1(.din(w_dff_B_kWE5Tpjh0_1),.dout(w_dff_B_XAOBa3Mx5_1),.clk(gclk));
	jdff dff_B_c1zz1fwu5_1(.din(w_dff_B_XAOBa3Mx5_1),.dout(w_dff_B_c1zz1fwu5_1),.clk(gclk));
	jdff dff_B_NxYGl2uN6_1(.din(n530),.dout(w_dff_B_NxYGl2uN6_1),.clk(gclk));
	jdff dff_B_1L2ItabO4_1(.din(w_dff_B_NxYGl2uN6_1),.dout(w_dff_B_1L2ItabO4_1),.clk(gclk));
	jdff dff_B_BafcEK5p1_1(.din(w_dff_B_1L2ItabO4_1),.dout(w_dff_B_BafcEK5p1_1),.clk(gclk));
	jdff dff_B_5BPUIjys6_1(.din(w_dff_B_BafcEK5p1_1),.dout(w_dff_B_5BPUIjys6_1),.clk(gclk));
	jdff dff_B_E8SJa8mo6_1(.din(w_dff_B_5BPUIjys6_1),.dout(w_dff_B_E8SJa8mo6_1),.clk(gclk));
	jdff dff_B_vrV1saZx8_1(.din(w_dff_B_E8SJa8mo6_1),.dout(w_dff_B_vrV1saZx8_1),.clk(gclk));
	jdff dff_B_8G05LpYR8_1(.din(w_dff_B_vrV1saZx8_1),.dout(w_dff_B_8G05LpYR8_1),.clk(gclk));
	jdff dff_B_VI28tZaS1_1(.din(w_dff_B_8G05LpYR8_1),.dout(w_dff_B_VI28tZaS1_1),.clk(gclk));
	jdff dff_B_DXE4c9xI2_1(.din(w_dff_B_VI28tZaS1_1),.dout(w_dff_B_DXE4c9xI2_1),.clk(gclk));
	jdff dff_B_3Xfoueyt3_1(.din(w_dff_B_DXE4c9xI2_1),.dout(w_dff_B_3Xfoueyt3_1),.clk(gclk));
	jdff dff_B_YYRw8vvW0_1(.din(w_dff_B_3Xfoueyt3_1),.dout(w_dff_B_YYRw8vvW0_1),.clk(gclk));
	jdff dff_B_JUwEIWLz9_1(.din(w_dff_B_YYRw8vvW0_1),.dout(w_dff_B_JUwEIWLz9_1),.clk(gclk));
	jdff dff_B_5ZjePXzK5_1(.din(w_dff_B_JUwEIWLz9_1),.dout(w_dff_B_5ZjePXzK5_1),.clk(gclk));
	jdff dff_B_RpRR36822_1(.din(w_dff_B_5ZjePXzK5_1),.dout(w_dff_B_RpRR36822_1),.clk(gclk));
	jdff dff_B_kW615ZDf3_1(.din(w_dff_B_RpRR36822_1),.dout(w_dff_B_kW615ZDf3_1),.clk(gclk));
	jdff dff_B_25PnaRh24_1(.din(w_dff_B_kW615ZDf3_1),.dout(w_dff_B_25PnaRh24_1),.clk(gclk));
	jdff dff_B_OhLTnKcC2_1(.din(w_dff_B_25PnaRh24_1),.dout(w_dff_B_OhLTnKcC2_1),.clk(gclk));
	jdff dff_B_MhejmIW43_1(.din(w_dff_B_OhLTnKcC2_1),.dout(w_dff_B_MhejmIW43_1),.clk(gclk));
	jdff dff_B_WpY32sTM7_1(.din(w_dff_B_MhejmIW43_1),.dout(w_dff_B_WpY32sTM7_1),.clk(gclk));
	jdff dff_B_ywyILbZb1_1(.din(w_dff_B_WpY32sTM7_1),.dout(w_dff_B_ywyILbZb1_1),.clk(gclk));
	jdff dff_B_CjdLPUiM5_1(.din(w_dff_B_ywyILbZb1_1),.dout(w_dff_B_CjdLPUiM5_1),.clk(gclk));
	jdff dff_B_fPk6YKlx7_1(.din(w_dff_B_CjdLPUiM5_1),.dout(w_dff_B_fPk6YKlx7_1),.clk(gclk));
	jdff dff_B_3lifHEZd4_1(.din(w_dff_B_fPk6YKlx7_1),.dout(w_dff_B_3lifHEZd4_1),.clk(gclk));
	jdff dff_B_z7vHNlC37_1(.din(w_dff_B_3lifHEZd4_1),.dout(w_dff_B_z7vHNlC37_1),.clk(gclk));
	jdff dff_B_YCOEgNde7_1(.din(w_dff_B_z7vHNlC37_1),.dout(w_dff_B_YCOEgNde7_1),.clk(gclk));
	jdff dff_B_q31oRVu59_1(.din(w_dff_B_YCOEgNde7_1),.dout(w_dff_B_q31oRVu59_1),.clk(gclk));
	jdff dff_B_54U1Ebai6_1(.din(w_dff_B_q31oRVu59_1),.dout(w_dff_B_54U1Ebai6_1),.clk(gclk));
	jdff dff_B_WgNOPtbR7_1(.din(n615),.dout(w_dff_B_WgNOPtbR7_1),.clk(gclk));
	jdff dff_B_pwhXadAr9_1(.din(w_dff_B_WgNOPtbR7_1),.dout(w_dff_B_pwhXadAr9_1),.clk(gclk));
	jdff dff_B_D1uHqIK13_1(.din(w_dff_B_pwhXadAr9_1),.dout(w_dff_B_D1uHqIK13_1),.clk(gclk));
	jdff dff_B_UQuUMfDF6_1(.din(w_dff_B_D1uHqIK13_1),.dout(w_dff_B_UQuUMfDF6_1),.clk(gclk));
	jdff dff_B_VHudfPek1_1(.din(w_dff_B_UQuUMfDF6_1),.dout(w_dff_B_VHudfPek1_1),.clk(gclk));
	jdff dff_B_FA28I9X16_1(.din(w_dff_B_VHudfPek1_1),.dout(w_dff_B_FA28I9X16_1),.clk(gclk));
	jdff dff_B_lustcrdz8_1(.din(w_dff_B_FA28I9X16_1),.dout(w_dff_B_lustcrdz8_1),.clk(gclk));
	jdff dff_B_B1sULxai5_1(.din(w_dff_B_lustcrdz8_1),.dout(w_dff_B_B1sULxai5_1),.clk(gclk));
	jdff dff_B_9NSKS4iH7_1(.din(w_dff_B_B1sULxai5_1),.dout(w_dff_B_9NSKS4iH7_1),.clk(gclk));
	jdff dff_B_BTC1j4ci8_1(.din(w_dff_B_9NSKS4iH7_1),.dout(w_dff_B_BTC1j4ci8_1),.clk(gclk));
	jdff dff_B_T4f05lYe2_1(.din(w_dff_B_BTC1j4ci8_1),.dout(w_dff_B_T4f05lYe2_1),.clk(gclk));
	jdff dff_B_J7vC8etz5_1(.din(w_dff_B_T4f05lYe2_1),.dout(w_dff_B_J7vC8etz5_1),.clk(gclk));
	jdff dff_B_yfadh71H6_1(.din(w_dff_B_J7vC8etz5_1),.dout(w_dff_B_yfadh71H6_1),.clk(gclk));
	jdff dff_B_lCvek3820_1(.din(w_dff_B_yfadh71H6_1),.dout(w_dff_B_lCvek3820_1),.clk(gclk));
	jdff dff_B_Cb2FTDkZ0_1(.din(w_dff_B_lCvek3820_1),.dout(w_dff_B_Cb2FTDkZ0_1),.clk(gclk));
	jdff dff_B_XDpT0z4L9_1(.din(w_dff_B_Cb2FTDkZ0_1),.dout(w_dff_B_XDpT0z4L9_1),.clk(gclk));
	jdff dff_B_ZWq9mVjX5_1(.din(w_dff_B_XDpT0z4L9_1),.dout(w_dff_B_ZWq9mVjX5_1),.clk(gclk));
	jdff dff_B_ojxTvVzN8_1(.din(w_dff_B_ZWq9mVjX5_1),.dout(w_dff_B_ojxTvVzN8_1),.clk(gclk));
	jdff dff_B_2n9rX5NF0_1(.din(w_dff_B_ojxTvVzN8_1),.dout(w_dff_B_2n9rX5NF0_1),.clk(gclk));
	jdff dff_B_xtAfkHVQ0_1(.din(w_dff_B_2n9rX5NF0_1),.dout(w_dff_B_xtAfkHVQ0_1),.clk(gclk));
	jdff dff_B_d1E1EsaN5_1(.din(w_dff_B_xtAfkHVQ0_1),.dout(w_dff_B_d1E1EsaN5_1),.clk(gclk));
	jdff dff_B_2xbHyuk16_1(.din(w_dff_B_d1E1EsaN5_1),.dout(w_dff_B_2xbHyuk16_1),.clk(gclk));
	jdff dff_B_MywtW5J48_1(.din(w_dff_B_2xbHyuk16_1),.dout(w_dff_B_MywtW5J48_1),.clk(gclk));
	jdff dff_B_zjo25QH17_1(.din(w_dff_B_MywtW5J48_1),.dout(w_dff_B_zjo25QH17_1),.clk(gclk));
	jdff dff_B_vjtwDPqG8_1(.din(w_dff_B_zjo25QH17_1),.dout(w_dff_B_vjtwDPqG8_1),.clk(gclk));
	jdff dff_B_o941zw169_1(.din(w_dff_B_vjtwDPqG8_1),.dout(w_dff_B_o941zw169_1),.clk(gclk));
	jdff dff_B_kZkDyc0g2_1(.din(w_dff_B_o941zw169_1),.dout(w_dff_B_kZkDyc0g2_1),.clk(gclk));
	jdff dff_B_FkzRXiDH9_1(.din(w_dff_B_kZkDyc0g2_1),.dout(w_dff_B_FkzRXiDH9_1),.clk(gclk));
	jdff dff_B_enIigK9G1_1(.din(w_dff_B_FkzRXiDH9_1),.dout(w_dff_B_enIigK9G1_1),.clk(gclk));
	jdff dff_B_DN4nkYGH0_1(.din(n707),.dout(w_dff_B_DN4nkYGH0_1),.clk(gclk));
	jdff dff_B_daZPsIaI8_1(.din(w_dff_B_DN4nkYGH0_1),.dout(w_dff_B_daZPsIaI8_1),.clk(gclk));
	jdff dff_B_tYYbO5dn3_1(.din(w_dff_B_daZPsIaI8_1),.dout(w_dff_B_tYYbO5dn3_1),.clk(gclk));
	jdff dff_B_uMpWvmzj5_1(.din(w_dff_B_tYYbO5dn3_1),.dout(w_dff_B_uMpWvmzj5_1),.clk(gclk));
	jdff dff_B_Zp53MIf52_1(.din(w_dff_B_uMpWvmzj5_1),.dout(w_dff_B_Zp53MIf52_1),.clk(gclk));
	jdff dff_B_97zjeKu91_1(.din(w_dff_B_Zp53MIf52_1),.dout(w_dff_B_97zjeKu91_1),.clk(gclk));
	jdff dff_B_Ek2XAlay5_1(.din(w_dff_B_97zjeKu91_1),.dout(w_dff_B_Ek2XAlay5_1),.clk(gclk));
	jdff dff_B_qD161yEY9_1(.din(w_dff_B_Ek2XAlay5_1),.dout(w_dff_B_qD161yEY9_1),.clk(gclk));
	jdff dff_B_A3v1x0ib6_1(.din(w_dff_B_qD161yEY9_1),.dout(w_dff_B_A3v1x0ib6_1),.clk(gclk));
	jdff dff_B_tBFU9LYF6_1(.din(w_dff_B_A3v1x0ib6_1),.dout(w_dff_B_tBFU9LYF6_1),.clk(gclk));
	jdff dff_B_em7tHQAn7_1(.din(w_dff_B_tBFU9LYF6_1),.dout(w_dff_B_em7tHQAn7_1),.clk(gclk));
	jdff dff_B_yiVf1GD43_1(.din(w_dff_B_em7tHQAn7_1),.dout(w_dff_B_yiVf1GD43_1),.clk(gclk));
	jdff dff_B_UVEjgrBr8_1(.din(w_dff_B_yiVf1GD43_1),.dout(w_dff_B_UVEjgrBr8_1),.clk(gclk));
	jdff dff_B_aEMieyYt2_1(.din(w_dff_B_UVEjgrBr8_1),.dout(w_dff_B_aEMieyYt2_1),.clk(gclk));
	jdff dff_B_jZFb2SLn7_1(.din(w_dff_B_aEMieyYt2_1),.dout(w_dff_B_jZFb2SLn7_1),.clk(gclk));
	jdff dff_B_rGb6IK2a2_1(.din(w_dff_B_jZFb2SLn7_1),.dout(w_dff_B_rGb6IK2a2_1),.clk(gclk));
	jdff dff_B_L1IzeLEC7_1(.din(w_dff_B_rGb6IK2a2_1),.dout(w_dff_B_L1IzeLEC7_1),.clk(gclk));
	jdff dff_B_dz67p68o8_1(.din(w_dff_B_L1IzeLEC7_1),.dout(w_dff_B_dz67p68o8_1),.clk(gclk));
	jdff dff_B_PD8HBJ9E5_1(.din(w_dff_B_dz67p68o8_1),.dout(w_dff_B_PD8HBJ9E5_1),.clk(gclk));
	jdff dff_B_CP34vhPg4_1(.din(w_dff_B_PD8HBJ9E5_1),.dout(w_dff_B_CP34vhPg4_1),.clk(gclk));
	jdff dff_B_hYMNgODB1_1(.din(w_dff_B_CP34vhPg4_1),.dout(w_dff_B_hYMNgODB1_1),.clk(gclk));
	jdff dff_B_OETIUeAI6_1(.din(w_dff_B_hYMNgODB1_1),.dout(w_dff_B_OETIUeAI6_1),.clk(gclk));
	jdff dff_B_odBswDdc9_1(.din(w_dff_B_OETIUeAI6_1),.dout(w_dff_B_odBswDdc9_1),.clk(gclk));
	jdff dff_B_lCDIlywy8_1(.din(w_dff_B_odBswDdc9_1),.dout(w_dff_B_lCDIlywy8_1),.clk(gclk));
	jdff dff_B_0uBAdJ4d8_1(.din(w_dff_B_lCDIlywy8_1),.dout(w_dff_B_0uBAdJ4d8_1),.clk(gclk));
	jdff dff_B_C9He6REg3_1(.din(w_dff_B_0uBAdJ4d8_1),.dout(w_dff_B_C9He6REg3_1),.clk(gclk));
	jdff dff_B_jhNC7s6L3_1(.din(w_dff_B_C9He6REg3_1),.dout(w_dff_B_jhNC7s6L3_1),.clk(gclk));
	jdff dff_B_yP7pFhl94_1(.din(w_dff_B_jhNC7s6L3_1),.dout(w_dff_B_yP7pFhl94_1),.clk(gclk));
	jdff dff_B_AnNMTJn20_1(.din(w_dff_B_yP7pFhl94_1),.dout(w_dff_B_AnNMTJn20_1),.clk(gclk));
	jdff dff_B_LVkMcXWe4_1(.din(w_dff_B_AnNMTJn20_1),.dout(w_dff_B_LVkMcXWe4_1),.clk(gclk));
	jdff dff_B_hOB0AtOD9_1(.din(w_dff_B_LVkMcXWe4_1),.dout(w_dff_B_hOB0AtOD9_1),.clk(gclk));
	jdff dff_B_Tk7wV1x59_1(.din(n806),.dout(w_dff_B_Tk7wV1x59_1),.clk(gclk));
	jdff dff_B_utRrxLn92_1(.din(w_dff_B_Tk7wV1x59_1),.dout(w_dff_B_utRrxLn92_1),.clk(gclk));
	jdff dff_B_Y8sUVSjt0_1(.din(w_dff_B_utRrxLn92_1),.dout(w_dff_B_Y8sUVSjt0_1),.clk(gclk));
	jdff dff_B_fdES0JQs8_1(.din(w_dff_B_Y8sUVSjt0_1),.dout(w_dff_B_fdES0JQs8_1),.clk(gclk));
	jdff dff_B_cEXRX9cm0_1(.din(w_dff_B_fdES0JQs8_1),.dout(w_dff_B_cEXRX9cm0_1),.clk(gclk));
	jdff dff_B_fakX5dCT6_1(.din(w_dff_B_cEXRX9cm0_1),.dout(w_dff_B_fakX5dCT6_1),.clk(gclk));
	jdff dff_B_gr5uCgK71_1(.din(w_dff_B_fakX5dCT6_1),.dout(w_dff_B_gr5uCgK71_1),.clk(gclk));
	jdff dff_B_p5swbb7p8_1(.din(w_dff_B_gr5uCgK71_1),.dout(w_dff_B_p5swbb7p8_1),.clk(gclk));
	jdff dff_B_mrSl81Yl6_1(.din(w_dff_B_p5swbb7p8_1),.dout(w_dff_B_mrSl81Yl6_1),.clk(gclk));
	jdff dff_B_QXICfYFg5_1(.din(w_dff_B_mrSl81Yl6_1),.dout(w_dff_B_QXICfYFg5_1),.clk(gclk));
	jdff dff_B_gptQrV040_1(.din(w_dff_B_QXICfYFg5_1),.dout(w_dff_B_gptQrV040_1),.clk(gclk));
	jdff dff_B_4jjwyFOG0_1(.din(w_dff_B_gptQrV040_1),.dout(w_dff_B_4jjwyFOG0_1),.clk(gclk));
	jdff dff_B_zfzNnqCc6_1(.din(w_dff_B_4jjwyFOG0_1),.dout(w_dff_B_zfzNnqCc6_1),.clk(gclk));
	jdff dff_B_qWMQWpFq9_1(.din(w_dff_B_zfzNnqCc6_1),.dout(w_dff_B_qWMQWpFq9_1),.clk(gclk));
	jdff dff_B_44qIIvi99_1(.din(w_dff_B_qWMQWpFq9_1),.dout(w_dff_B_44qIIvi99_1),.clk(gclk));
	jdff dff_B_lo1K324g8_1(.din(w_dff_B_44qIIvi99_1),.dout(w_dff_B_lo1K324g8_1),.clk(gclk));
	jdff dff_B_gJv09Qok4_1(.din(w_dff_B_lo1K324g8_1),.dout(w_dff_B_gJv09Qok4_1),.clk(gclk));
	jdff dff_B_S1aAAp0O6_1(.din(w_dff_B_gJv09Qok4_1),.dout(w_dff_B_S1aAAp0O6_1),.clk(gclk));
	jdff dff_B_u62KfPAb1_1(.din(w_dff_B_S1aAAp0O6_1),.dout(w_dff_B_u62KfPAb1_1),.clk(gclk));
	jdff dff_B_2N0GWwYC9_1(.din(w_dff_B_u62KfPAb1_1),.dout(w_dff_B_2N0GWwYC9_1),.clk(gclk));
	jdff dff_B_vx5kiSt78_1(.din(w_dff_B_2N0GWwYC9_1),.dout(w_dff_B_vx5kiSt78_1),.clk(gclk));
	jdff dff_B_gvNJmRDX9_1(.din(w_dff_B_vx5kiSt78_1),.dout(w_dff_B_gvNJmRDX9_1),.clk(gclk));
	jdff dff_B_OueJZUUO7_1(.din(w_dff_B_gvNJmRDX9_1),.dout(w_dff_B_OueJZUUO7_1),.clk(gclk));
	jdff dff_B_kBVGO1xB8_1(.din(w_dff_B_OueJZUUO7_1),.dout(w_dff_B_kBVGO1xB8_1),.clk(gclk));
	jdff dff_B_I66AOxMl8_1(.din(w_dff_B_kBVGO1xB8_1),.dout(w_dff_B_I66AOxMl8_1),.clk(gclk));
	jdff dff_B_2pKtVac62_1(.din(w_dff_B_I66AOxMl8_1),.dout(w_dff_B_2pKtVac62_1),.clk(gclk));
	jdff dff_B_yVQkM1H66_1(.din(w_dff_B_2pKtVac62_1),.dout(w_dff_B_yVQkM1H66_1),.clk(gclk));
	jdff dff_B_to30z33n7_1(.din(w_dff_B_yVQkM1H66_1),.dout(w_dff_B_to30z33n7_1),.clk(gclk));
	jdff dff_B_FPhJtWp79_1(.din(w_dff_B_to30z33n7_1),.dout(w_dff_B_FPhJtWp79_1),.clk(gclk));
	jdff dff_B_lN9gcYhF1_1(.din(w_dff_B_FPhJtWp79_1),.dout(w_dff_B_lN9gcYhF1_1),.clk(gclk));
	jdff dff_B_y2yx8tk69_1(.din(w_dff_B_lN9gcYhF1_1),.dout(w_dff_B_y2yx8tk69_1),.clk(gclk));
	jdff dff_B_1z8N5QVY8_1(.din(w_dff_B_y2yx8tk69_1),.dout(w_dff_B_1z8N5QVY8_1),.clk(gclk));
	jdff dff_B_bKVskMcs8_1(.din(w_dff_B_1z8N5QVY8_1),.dout(w_dff_B_bKVskMcs8_1),.clk(gclk));
	jdff dff_B_pI24JtGM4_0(.din(n1296),.dout(w_dff_B_pI24JtGM4_0),.clk(gclk));
	jdff dff_B_L0lJCq0a1_1(.din(n1811),.dout(w_dff_B_L0lJCq0a1_1),.clk(gclk));
	jdff dff_B_90IjmZ2U2_1(.din(w_dff_B_L0lJCq0a1_1),.dout(w_dff_B_90IjmZ2U2_1),.clk(gclk));
	jdff dff_B_zjc0t6o19_1(.din(w_dff_B_90IjmZ2U2_1),.dout(w_dff_B_zjc0t6o19_1),.clk(gclk));
	jdff dff_B_kZYiTLjE5_1(.din(w_dff_B_zjc0t6o19_1),.dout(w_dff_B_kZYiTLjE5_1),.clk(gclk));
	jdff dff_B_hiB8ofTa5_1(.din(w_dff_B_kZYiTLjE5_1),.dout(w_dff_B_hiB8ofTa5_1),.clk(gclk));
	jdff dff_B_AIOufWfd4_1(.din(w_dff_B_hiB8ofTa5_1),.dout(w_dff_B_AIOufWfd4_1),.clk(gclk));
	jdff dff_B_SYkn1LZE6_1(.din(w_dff_B_AIOufWfd4_1),.dout(w_dff_B_SYkn1LZE6_1),.clk(gclk));
	jdff dff_B_IqTVostd0_0(.din(n1819),.dout(w_dff_B_IqTVostd0_0),.clk(gclk));
	jdff dff_B_K2FZU5Ca1_0(.din(w_dff_B_IqTVostd0_0),.dout(w_dff_B_K2FZU5Ca1_0),.clk(gclk));
	jdff dff_B_1PHCjzAR5_0(.din(w_dff_B_K2FZU5Ca1_0),.dout(w_dff_B_1PHCjzAR5_0),.clk(gclk));
	jdff dff_B_jDBZ49te8_0(.din(w_dff_B_1PHCjzAR5_0),.dout(w_dff_B_jDBZ49te8_0),.clk(gclk));
	jdff dff_B_Hud6zxaB7_0(.din(w_dff_B_jDBZ49te8_0),.dout(w_dff_B_Hud6zxaB7_0),.clk(gclk));
	jdff dff_A_W0ePeiK66_0(.dout(w_n1818_0[0]),.din(w_dff_A_W0ePeiK66_0),.clk(gclk));
	jdff dff_A_MFPSpaIB9_0(.dout(w_dff_A_W0ePeiK66_0),.din(w_dff_A_MFPSpaIB9_0),.clk(gclk));
	jdff dff_A_OBoyWszB3_0(.dout(w_dff_A_MFPSpaIB9_0),.din(w_dff_A_OBoyWszB3_0),.clk(gclk));
	jdff dff_A_goyEREVc2_0(.dout(w_dff_A_OBoyWszB3_0),.din(w_dff_A_goyEREVc2_0),.clk(gclk));
	jdff dff_A_xBmmHKr30_0(.dout(w_dff_A_goyEREVc2_0),.din(w_dff_A_xBmmHKr30_0),.clk(gclk));
	jdff dff_A_Xwkf2BHt1_0(.dout(w_dff_A_xBmmHKr30_0),.din(w_dff_A_Xwkf2BHt1_0),.clk(gclk));
	jdff dff_B_xx6l7qui3_1(.din(n1808),.dout(w_dff_B_xx6l7qui3_1),.clk(gclk));
	jdff dff_B_mn4rCjzz0_1(.din(w_dff_B_xx6l7qui3_1),.dout(w_dff_B_mn4rCjzz0_1),.clk(gclk));
	jdff dff_B_lE7QRb345_2(.din(n1807),.dout(w_dff_B_lE7QRb345_2),.clk(gclk));
	jdff dff_B_8pCulNH83_2(.din(w_dff_B_lE7QRb345_2),.dout(w_dff_B_8pCulNH83_2),.clk(gclk));
	jdff dff_B_Qf6y5UA72_2(.din(w_dff_B_8pCulNH83_2),.dout(w_dff_B_Qf6y5UA72_2),.clk(gclk));
	jdff dff_B_ObuV6XP09_2(.din(w_dff_B_Qf6y5UA72_2),.dout(w_dff_B_ObuV6XP09_2),.clk(gclk));
	jdff dff_B_u7Woywot6_2(.din(w_dff_B_ObuV6XP09_2),.dout(w_dff_B_u7Woywot6_2),.clk(gclk));
	jdff dff_B_88T758w23_2(.din(w_dff_B_u7Woywot6_2),.dout(w_dff_B_88T758w23_2),.clk(gclk));
	jdff dff_B_zNi7oP3q8_2(.din(w_dff_B_88T758w23_2),.dout(w_dff_B_zNi7oP3q8_2),.clk(gclk));
	jdff dff_B_iYnjBo3z1_2(.din(w_dff_B_zNi7oP3q8_2),.dout(w_dff_B_iYnjBo3z1_2),.clk(gclk));
	jdff dff_B_yl7rMzmQ8_2(.din(w_dff_B_iYnjBo3z1_2),.dout(w_dff_B_yl7rMzmQ8_2),.clk(gclk));
	jdff dff_B_AirbCeqY3_2(.din(w_dff_B_yl7rMzmQ8_2),.dout(w_dff_B_AirbCeqY3_2),.clk(gclk));
	jdff dff_B_PX3Ryoyl5_2(.din(w_dff_B_AirbCeqY3_2),.dout(w_dff_B_PX3Ryoyl5_2),.clk(gclk));
	jdff dff_B_OlxbPXNB9_2(.din(w_dff_B_PX3Ryoyl5_2),.dout(w_dff_B_OlxbPXNB9_2),.clk(gclk));
	jdff dff_B_eiOJyZqL6_2(.din(w_dff_B_OlxbPXNB9_2),.dout(w_dff_B_eiOJyZqL6_2),.clk(gclk));
	jdff dff_B_jVuwhZvT8_2(.din(w_dff_B_eiOJyZqL6_2),.dout(w_dff_B_jVuwhZvT8_2),.clk(gclk));
	jdff dff_B_GL3slo7Z1_2(.din(w_dff_B_jVuwhZvT8_2),.dout(w_dff_B_GL3slo7Z1_2),.clk(gclk));
	jdff dff_B_1fIBqJmy8_2(.din(w_dff_B_GL3slo7Z1_2),.dout(w_dff_B_1fIBqJmy8_2),.clk(gclk));
	jdff dff_B_ZSRgh43m4_2(.din(w_dff_B_1fIBqJmy8_2),.dout(w_dff_B_ZSRgh43m4_2),.clk(gclk));
	jdff dff_B_RnSgaOmr8_2(.din(w_dff_B_ZSRgh43m4_2),.dout(w_dff_B_RnSgaOmr8_2),.clk(gclk));
	jdff dff_B_wgHEkmyy6_2(.din(w_dff_B_RnSgaOmr8_2),.dout(w_dff_B_wgHEkmyy6_2),.clk(gclk));
	jdff dff_B_DGdKhsWa1_2(.din(w_dff_B_wgHEkmyy6_2),.dout(w_dff_B_DGdKhsWa1_2),.clk(gclk));
	jdff dff_B_EuGidYqY6_2(.din(w_dff_B_DGdKhsWa1_2),.dout(w_dff_B_EuGidYqY6_2),.clk(gclk));
	jdff dff_B_FYFisWGb9_2(.din(w_dff_B_EuGidYqY6_2),.dout(w_dff_B_FYFisWGb9_2),.clk(gclk));
	jdff dff_B_Yujf99G73_2(.din(w_dff_B_FYFisWGb9_2),.dout(w_dff_B_Yujf99G73_2),.clk(gclk));
	jdff dff_B_VQizus1p1_2(.din(w_dff_B_Yujf99G73_2),.dout(w_dff_B_VQizus1p1_2),.clk(gclk));
	jdff dff_B_qUkau1RW4_2(.din(w_dff_B_VQizus1p1_2),.dout(w_dff_B_qUkau1RW4_2),.clk(gclk));
	jdff dff_B_SjNiWd1k0_2(.din(w_dff_B_qUkau1RW4_2),.dout(w_dff_B_SjNiWd1k0_2),.clk(gclk));
	jdff dff_B_mSM1Xl9R5_2(.din(w_dff_B_SjNiWd1k0_2),.dout(w_dff_B_mSM1Xl9R5_2),.clk(gclk));
	jdff dff_B_hM7KeAsn4_2(.din(w_dff_B_mSM1Xl9R5_2),.dout(w_dff_B_hM7KeAsn4_2),.clk(gclk));
	jdff dff_B_M9VDviPH7_2(.din(w_dff_B_hM7KeAsn4_2),.dout(w_dff_B_M9VDviPH7_2),.clk(gclk));
	jdff dff_B_waMO7DUW5_2(.din(w_dff_B_M9VDviPH7_2),.dout(w_dff_B_waMO7DUW5_2),.clk(gclk));
	jdff dff_B_IleYBp5n1_2(.din(w_dff_B_waMO7DUW5_2),.dout(w_dff_B_IleYBp5n1_2),.clk(gclk));
	jdff dff_B_1KgAOyTA0_2(.din(w_dff_B_IleYBp5n1_2),.dout(w_dff_B_1KgAOyTA0_2),.clk(gclk));
	jdff dff_B_VIDOZ50d4_2(.din(w_dff_B_1KgAOyTA0_2),.dout(w_dff_B_VIDOZ50d4_2),.clk(gclk));
	jdff dff_B_X62xnjUP3_2(.din(w_dff_B_VIDOZ50d4_2),.dout(w_dff_B_X62xnjUP3_2),.clk(gclk));
	jdff dff_B_LZkHANrP5_2(.din(w_dff_B_X62xnjUP3_2),.dout(w_dff_B_LZkHANrP5_2),.clk(gclk));
	jdff dff_B_rH9JTWna4_2(.din(w_dff_B_LZkHANrP5_2),.dout(w_dff_B_rH9JTWna4_2),.clk(gclk));
	jdff dff_B_NPqX5pqK9_2(.din(w_dff_B_rH9JTWna4_2),.dout(w_dff_B_NPqX5pqK9_2),.clk(gclk));
	jdff dff_B_iLKLZ3HG3_2(.din(w_dff_B_NPqX5pqK9_2),.dout(w_dff_B_iLKLZ3HG3_2),.clk(gclk));
	jdff dff_B_jGz6bc6R3_2(.din(w_dff_B_iLKLZ3HG3_2),.dout(w_dff_B_jGz6bc6R3_2),.clk(gclk));
	jdff dff_B_FSxwYpwN8_2(.din(w_dff_B_jGz6bc6R3_2),.dout(w_dff_B_FSxwYpwN8_2),.clk(gclk));
	jdff dff_B_faF78IKG6_2(.din(w_dff_B_FSxwYpwN8_2),.dout(w_dff_B_faF78IKG6_2),.clk(gclk));
	jdff dff_B_ZJgFeNct6_2(.din(w_dff_B_faF78IKG6_2),.dout(w_dff_B_ZJgFeNct6_2),.clk(gclk));
	jdff dff_B_CaMxzjt13_2(.din(w_dff_B_ZJgFeNct6_2),.dout(w_dff_B_CaMxzjt13_2),.clk(gclk));
	jdff dff_B_UaMFD9u46_1(.din(n1814),.dout(w_dff_B_UaMFD9u46_1),.clk(gclk));
	jdff dff_B_2kjpgPmk6_1(.din(w_dff_B_UaMFD9u46_1),.dout(w_dff_B_2kjpgPmk6_1),.clk(gclk));
	jdff dff_B_5LWtGzuY8_1(.din(w_dff_B_2kjpgPmk6_1),.dout(w_dff_B_5LWtGzuY8_1),.clk(gclk));
	jdff dff_B_aJP7bq8n8_1(.din(w_dff_B_5LWtGzuY8_1),.dout(w_dff_B_aJP7bq8n8_1),.clk(gclk));
	jdff dff_B_LWJ4q85k1_1(.din(w_dff_B_aJP7bq8n8_1),.dout(w_dff_B_LWJ4q85k1_1),.clk(gclk));
	jdff dff_B_tZ589fHD3_0(.din(n1815),.dout(w_dff_B_tZ589fHD3_0),.clk(gclk));
	jdff dff_B_jkygkTSI3_0(.din(w_dff_B_tZ589fHD3_0),.dout(w_dff_B_jkygkTSI3_0),.clk(gclk));
	jdff dff_B_GKJ3ibl99_0(.din(w_dff_B_jkygkTSI3_0),.dout(w_dff_B_GKJ3ibl99_0),.clk(gclk));
	jdff dff_B_S4ltgIP69_0(.din(w_dff_B_GKJ3ibl99_0),.dout(w_dff_B_S4ltgIP69_0),.clk(gclk));
	jdff dff_A_xuiwnLhZ9_1(.dout(w_n1805_0[1]),.din(w_dff_A_xuiwnLhZ9_1),.clk(gclk));
	jdff dff_A_kKEoqttp9_1(.dout(w_dff_A_xuiwnLhZ9_1),.din(w_dff_A_kKEoqttp9_1),.clk(gclk));
	jdff dff_A_rBeQwzzF2_1(.dout(w_dff_A_kKEoqttp9_1),.din(w_dff_A_rBeQwzzF2_1),.clk(gclk));
	jdff dff_A_J7NxZJ3L7_1(.dout(w_dff_A_rBeQwzzF2_1),.din(w_dff_A_J7NxZJ3L7_1),.clk(gclk));
	jdff dff_A_7HgF2Ebz3_1(.dout(w_dff_A_J7NxZJ3L7_1),.din(w_dff_A_7HgF2Ebz3_1),.clk(gclk));
	jdff dff_B_zeANGTQO9_1(.din(n1790),.dout(w_dff_B_zeANGTQO9_1),.clk(gclk));
	jdff dff_B_W2fm52nh9_1(.din(w_dff_B_zeANGTQO9_1),.dout(w_dff_B_W2fm52nh9_1),.clk(gclk));
	jdff dff_B_tjxn3Cha9_1(.din(w_dff_B_W2fm52nh9_1),.dout(w_dff_B_tjxn3Cha9_1),.clk(gclk));
	jdff dff_B_xy2ZCBsW6_1(.din(w_dff_B_tjxn3Cha9_1),.dout(w_dff_B_xy2ZCBsW6_1),.clk(gclk));
	jdff dff_B_SeIcI13K2_1(.din(w_dff_B_xy2ZCBsW6_1),.dout(w_dff_B_SeIcI13K2_1),.clk(gclk));
	jdff dff_B_Bg2e2mZh0_0(.din(n1791),.dout(w_dff_B_Bg2e2mZh0_0),.clk(gclk));
	jdff dff_B_9LfwhznL4_0(.din(w_dff_B_Bg2e2mZh0_0),.dout(w_dff_B_9LfwhznL4_0),.clk(gclk));
	jdff dff_B_HjZbioiq5_0(.din(w_dff_B_9LfwhznL4_0),.dout(w_dff_B_HjZbioiq5_0),.clk(gclk));
	jdff dff_B_UKeQvCg87_0(.din(w_dff_B_HjZbioiq5_0),.dout(w_dff_B_UKeQvCg87_0),.clk(gclk));
	jdff dff_A_UmyjqEiB3_1(.dout(w_n1786_0[1]),.din(w_dff_A_UmyjqEiB3_1),.clk(gclk));
	jdff dff_A_g2W2EC9J8_1(.dout(w_dff_A_UmyjqEiB3_1),.din(w_dff_A_g2W2EC9J8_1),.clk(gclk));
	jdff dff_A_7nZHykkt0_1(.dout(w_dff_A_g2W2EC9J8_1),.din(w_dff_A_7nZHykkt0_1),.clk(gclk));
	jdff dff_A_iKTDXahH9_1(.dout(w_dff_A_7nZHykkt0_1),.din(w_dff_A_iKTDXahH9_1),.clk(gclk));
	jdff dff_A_dLavTA406_1(.dout(w_dff_A_iKTDXahH9_1),.din(w_dff_A_dLavTA406_1),.clk(gclk));
	jdff dff_B_opUNiU9e4_1(.din(n1764),.dout(w_dff_B_opUNiU9e4_1),.clk(gclk));
	jdff dff_B_FXWqG8P88_1(.din(w_dff_B_opUNiU9e4_1),.dout(w_dff_B_FXWqG8P88_1),.clk(gclk));
	jdff dff_B_aTNh3bMG2_1(.din(w_dff_B_FXWqG8P88_1),.dout(w_dff_B_aTNh3bMG2_1),.clk(gclk));
	jdff dff_B_9K7NBD5C3_1(.din(w_dff_B_aTNh3bMG2_1),.dout(w_dff_B_9K7NBD5C3_1),.clk(gclk));
	jdff dff_B_LBz8FDdd7_1(.din(w_dff_B_9K7NBD5C3_1),.dout(w_dff_B_LBz8FDdd7_1),.clk(gclk));
	jdff dff_B_lxBwEA4n3_0(.din(n1765),.dout(w_dff_B_lxBwEA4n3_0),.clk(gclk));
	jdff dff_B_65s5OWsu0_0(.din(w_dff_B_lxBwEA4n3_0),.dout(w_dff_B_65s5OWsu0_0),.clk(gclk));
	jdff dff_B_rYAiRxjA9_0(.din(w_dff_B_65s5OWsu0_0),.dout(w_dff_B_rYAiRxjA9_0),.clk(gclk));
	jdff dff_B_5ubhJ4Ul9_0(.din(w_dff_B_rYAiRxjA9_0),.dout(w_dff_B_5ubhJ4Ul9_0),.clk(gclk));
	jdff dff_A_f238AYfa5_1(.dout(w_n1760_0[1]),.din(w_dff_A_f238AYfa5_1),.clk(gclk));
	jdff dff_A_E5jJywQ17_1(.dout(w_dff_A_f238AYfa5_1),.din(w_dff_A_E5jJywQ17_1),.clk(gclk));
	jdff dff_A_6DUvxiW19_1(.dout(w_dff_A_E5jJywQ17_1),.din(w_dff_A_6DUvxiW19_1),.clk(gclk));
	jdff dff_A_32ZOwtlv4_1(.dout(w_dff_A_6DUvxiW19_1),.din(w_dff_A_32ZOwtlv4_1),.clk(gclk));
	jdff dff_A_wwb1llDO5_1(.dout(w_dff_A_32ZOwtlv4_1),.din(w_dff_A_wwb1llDO5_1),.clk(gclk));
	jdff dff_B_QVKlm6nG3_1(.din(n1731),.dout(w_dff_B_QVKlm6nG3_1),.clk(gclk));
	jdff dff_B_2aPVKMdH7_1(.din(w_dff_B_QVKlm6nG3_1),.dout(w_dff_B_2aPVKMdH7_1),.clk(gclk));
	jdff dff_B_3LlaYMpX1_1(.din(w_dff_B_2aPVKMdH7_1),.dout(w_dff_B_3LlaYMpX1_1),.clk(gclk));
	jdff dff_B_xgLbS7ef2_1(.din(w_dff_B_3LlaYMpX1_1),.dout(w_dff_B_xgLbS7ef2_1),.clk(gclk));
	jdff dff_B_v9bnab3R2_1(.din(w_dff_B_xgLbS7ef2_1),.dout(w_dff_B_v9bnab3R2_1),.clk(gclk));
	jdff dff_B_dsWpZ4tF8_0(.din(n1732),.dout(w_dff_B_dsWpZ4tF8_0),.clk(gclk));
	jdff dff_B_sotNSENx5_0(.din(w_dff_B_dsWpZ4tF8_0),.dout(w_dff_B_sotNSENx5_0),.clk(gclk));
	jdff dff_B_mxLQyMKv5_0(.din(w_dff_B_sotNSENx5_0),.dout(w_dff_B_mxLQyMKv5_0),.clk(gclk));
	jdff dff_B_lculz7TR9_0(.din(w_dff_B_mxLQyMKv5_0),.dout(w_dff_B_lculz7TR9_0),.clk(gclk));
	jdff dff_A_haUmetS19_1(.dout(w_n1727_0[1]),.din(w_dff_A_haUmetS19_1),.clk(gclk));
	jdff dff_A_9g1Wf2nE0_1(.dout(w_dff_A_haUmetS19_1),.din(w_dff_A_9g1Wf2nE0_1),.clk(gclk));
	jdff dff_A_9HZ3DGBc6_1(.dout(w_dff_A_9g1Wf2nE0_1),.din(w_dff_A_9HZ3DGBc6_1),.clk(gclk));
	jdff dff_A_GQ9guesq5_1(.dout(w_dff_A_9HZ3DGBc6_1),.din(w_dff_A_GQ9guesq5_1),.clk(gclk));
	jdff dff_A_nw0zklZx2_1(.dout(w_dff_A_GQ9guesq5_1),.din(w_dff_A_nw0zklZx2_1),.clk(gclk));
	jdff dff_B_7l0Me6jS2_1(.din(n1691),.dout(w_dff_B_7l0Me6jS2_1),.clk(gclk));
	jdff dff_B_0sDZLPxK5_1(.din(w_dff_B_7l0Me6jS2_1),.dout(w_dff_B_0sDZLPxK5_1),.clk(gclk));
	jdff dff_B_oYxPY6s27_1(.din(w_dff_B_0sDZLPxK5_1),.dout(w_dff_B_oYxPY6s27_1),.clk(gclk));
	jdff dff_B_dgNyMpz47_1(.din(w_dff_B_oYxPY6s27_1),.dout(w_dff_B_dgNyMpz47_1),.clk(gclk));
	jdff dff_B_3YCoDQeY1_1(.din(w_dff_B_dgNyMpz47_1),.dout(w_dff_B_3YCoDQeY1_1),.clk(gclk));
	jdff dff_B_rMHj3k131_0(.din(n1692),.dout(w_dff_B_rMHj3k131_0),.clk(gclk));
	jdff dff_B_fqTUIr7f6_0(.din(w_dff_B_rMHj3k131_0),.dout(w_dff_B_fqTUIr7f6_0),.clk(gclk));
	jdff dff_B_dN7mMsn83_0(.din(w_dff_B_fqTUIr7f6_0),.dout(w_dff_B_dN7mMsn83_0),.clk(gclk));
	jdff dff_A_HmaB0Zgm4_1(.dout(w_n1689_0[1]),.din(w_dff_A_HmaB0Zgm4_1),.clk(gclk));
	jdff dff_A_Ml8at2Oa9_1(.dout(w_dff_A_HmaB0Zgm4_1),.din(w_dff_A_Ml8at2Oa9_1),.clk(gclk));
	jdff dff_A_zEYZS2gD6_1(.dout(w_dff_A_Ml8at2Oa9_1),.din(w_dff_A_zEYZS2gD6_1),.clk(gclk));
	jdff dff_A_ixcFa8oL9_1(.dout(w_dff_A_zEYZS2gD6_1),.din(w_dff_A_ixcFa8oL9_1),.clk(gclk));
	jdff dff_B_GG62YzVH8_1(.din(n1643),.dout(w_dff_B_GG62YzVH8_1),.clk(gclk));
	jdff dff_B_rGI26zXL7_1(.din(w_dff_B_GG62YzVH8_1),.dout(w_dff_B_rGI26zXL7_1),.clk(gclk));
	jdff dff_B_vCwvBcrj8_1(.din(w_dff_B_rGI26zXL7_1),.dout(w_dff_B_vCwvBcrj8_1),.clk(gclk));
	jdff dff_B_8QhDajyx7_1(.din(w_dff_B_vCwvBcrj8_1),.dout(w_dff_B_8QhDajyx7_1),.clk(gclk));
	jdff dff_B_EJmoYI6o3_0(.din(n1644),.dout(w_dff_B_EJmoYI6o3_0),.clk(gclk));
	jdff dff_B_f4Eih3xY4_0(.din(w_dff_B_EJmoYI6o3_0),.dout(w_dff_B_f4Eih3xY4_0),.clk(gclk));
	jdff dff_A_nLDtfdqs7_1(.dout(w_n1641_0[1]),.din(w_dff_A_nLDtfdqs7_1),.clk(gclk));
	jdff dff_A_KeQP5j814_1(.dout(w_dff_A_nLDtfdqs7_1),.din(w_dff_A_KeQP5j814_1),.clk(gclk));
	jdff dff_A_my0cukNQ9_1(.dout(w_dff_A_KeQP5j814_1),.din(w_dff_A_my0cukNQ9_1),.clk(gclk));
	jdff dff_B_lLTCaoQP0_1(.din(n1588),.dout(w_dff_B_lLTCaoQP0_1),.clk(gclk));
	jdff dff_B_m9I7jFRb9_1(.din(w_dff_B_lLTCaoQP0_1),.dout(w_dff_B_m9I7jFRb9_1),.clk(gclk));
	jdff dff_B_qI9DitWk4_1(.din(w_dff_B_m9I7jFRb9_1),.dout(w_dff_B_qI9DitWk4_1),.clk(gclk));
	jdff dff_B_UekR6NNa3_1(.din(w_dff_B_qI9DitWk4_1),.dout(w_dff_B_UekR6NNa3_1),.clk(gclk));
	jdff dff_B_q6FgAOK44_0(.din(n1589),.dout(w_dff_B_q6FgAOK44_0),.clk(gclk));
	jdff dff_B_FwpMwxfk6_0(.din(w_dff_B_q6FgAOK44_0),.dout(w_dff_B_FwpMwxfk6_0),.clk(gclk));
	jdff dff_A_GRKxZznQ3_1(.dout(w_n1586_0[1]),.din(w_dff_A_GRKxZznQ3_1),.clk(gclk));
	jdff dff_A_BxhsF5cW3_1(.dout(w_dff_A_GRKxZznQ3_1),.din(w_dff_A_BxhsF5cW3_1),.clk(gclk));
	jdff dff_A_2W8eSvNS9_1(.dout(w_dff_A_BxhsF5cW3_1),.din(w_dff_A_2W8eSvNS9_1),.clk(gclk));
	jdff dff_B_lojryFKB0_1(.din(n1526),.dout(w_dff_B_lojryFKB0_1),.clk(gclk));
	jdff dff_B_aJt4jwp71_1(.din(w_dff_B_lojryFKB0_1),.dout(w_dff_B_aJt4jwp71_1),.clk(gclk));
	jdff dff_B_ErnfkFhA3_1(.din(w_dff_B_aJt4jwp71_1),.dout(w_dff_B_ErnfkFhA3_1),.clk(gclk));
	jdff dff_B_AIG6bJtq8_1(.din(w_dff_B_ErnfkFhA3_1),.dout(w_dff_B_AIG6bJtq8_1),.clk(gclk));
	jdff dff_B_t5NPkjVm4_0(.din(n1527),.dout(w_dff_B_t5NPkjVm4_0),.clk(gclk));
	jdff dff_B_xA4A4SQ38_0(.din(w_dff_B_t5NPkjVm4_0),.dout(w_dff_B_xA4A4SQ38_0),.clk(gclk));
	jdff dff_A_MhEnWH1e4_1(.dout(w_n1524_0[1]),.din(w_dff_A_MhEnWH1e4_1),.clk(gclk));
	jdff dff_A_OjP6DQj17_1(.dout(w_dff_A_MhEnWH1e4_1),.din(w_dff_A_OjP6DQj17_1),.clk(gclk));
	jdff dff_A_Q4KL71pY0_1(.dout(w_dff_A_OjP6DQj17_1),.din(w_dff_A_Q4KL71pY0_1),.clk(gclk));
	jdff dff_B_JhwNLh4z5_1(.din(n1457),.dout(w_dff_B_JhwNLh4z5_1),.clk(gclk));
	jdff dff_B_MNJcPB5i0_1(.din(w_dff_B_JhwNLh4z5_1),.dout(w_dff_B_MNJcPB5i0_1),.clk(gclk));
	jdff dff_B_GL8yvwSr3_1(.din(w_dff_B_MNJcPB5i0_1),.dout(w_dff_B_GL8yvwSr3_1),.clk(gclk));
	jdff dff_B_zEQtFjHc9_1(.din(w_dff_B_GL8yvwSr3_1),.dout(w_dff_B_zEQtFjHc9_1),.clk(gclk));
	jdff dff_B_L7vuoqVx1_0(.din(n1458),.dout(w_dff_B_L7vuoqVx1_0),.clk(gclk));
	jdff dff_B_UJiY7Bnj3_0(.din(w_dff_B_L7vuoqVx1_0),.dout(w_dff_B_UJiY7Bnj3_0),.clk(gclk));
	jdff dff_A_9zNi1lLP1_1(.dout(w_n1455_0[1]),.din(w_dff_A_9zNi1lLP1_1),.clk(gclk));
	jdff dff_A_AYMSnguH9_1(.dout(w_dff_A_9zNi1lLP1_1),.din(w_dff_A_AYMSnguH9_1),.clk(gclk));
	jdff dff_A_1RrEBp7h4_1(.dout(w_dff_A_AYMSnguH9_1),.din(w_dff_A_1RrEBp7h4_1),.clk(gclk));
	jdff dff_B_czyWzkBd8_1(.din(n1381),.dout(w_dff_B_czyWzkBd8_1),.clk(gclk));
	jdff dff_B_clKURfb93_1(.din(w_dff_B_czyWzkBd8_1),.dout(w_dff_B_clKURfb93_1),.clk(gclk));
	jdff dff_B_vE7MgVrH1_1(.din(w_dff_B_clKURfb93_1),.dout(w_dff_B_vE7MgVrH1_1),.clk(gclk));
	jdff dff_B_NAMTOoqD0_1(.din(w_dff_B_vE7MgVrH1_1),.dout(w_dff_B_NAMTOoqD0_1),.clk(gclk));
	jdff dff_B_s2uwMy4s4_0(.din(n1382),.dout(w_dff_B_s2uwMy4s4_0),.clk(gclk));
	jdff dff_B_w2l7Nkfj6_0(.din(w_dff_B_s2uwMy4s4_0),.dout(w_dff_B_w2l7Nkfj6_0),.clk(gclk));
	jdff dff_A_6S9ZFhC44_1(.dout(w_n1379_0[1]),.din(w_dff_A_6S9ZFhC44_1),.clk(gclk));
	jdff dff_A_ddKYqWmG2_1(.dout(w_dff_A_6S9ZFhC44_1),.din(w_dff_A_ddKYqWmG2_1),.clk(gclk));
	jdff dff_A_cFG0Ia5Z3_1(.dout(w_dff_A_ddKYqWmG2_1),.din(w_dff_A_cFG0Ia5Z3_1),.clk(gclk));
	jdff dff_B_Hqoe6YU48_1(.din(n1299),.dout(w_dff_B_Hqoe6YU48_1),.clk(gclk));
	jdff dff_B_WSwqW1o59_1(.din(w_dff_B_Hqoe6YU48_1),.dout(w_dff_B_WSwqW1o59_1),.clk(gclk));
	jdff dff_B_n6bnUqnb4_1(.din(w_dff_B_WSwqW1o59_1),.dout(w_dff_B_n6bnUqnb4_1),.clk(gclk));
	jdff dff_A_uVhFRkNE4_0(.dout(w_n1295_0[0]),.din(w_dff_A_uVhFRkNE4_0),.clk(gclk));
	jdff dff_A_SX75LK7v5_0(.dout(w_dff_A_uVhFRkNE4_0),.din(w_dff_A_SX75LK7v5_0),.clk(gclk));
	jdff dff_B_NpeQjmGC5_1(.din(n1211),.dout(w_dff_B_NpeQjmGC5_1),.clk(gclk));
	jdff dff_A_BPfeRMEG5_0(.dout(w_n1207_0[0]),.din(w_dff_A_BPfeRMEG5_0),.clk(gclk));
	jdff dff_B_8GXt3znx8_1(.din(n1113),.dout(w_dff_B_8GXt3znx8_1),.clk(gclk));
	jdff dff_A_eim6TkIP3_0(.dout(w_n1109_0[0]),.din(w_dff_A_eim6TkIP3_0),.clk(gclk));
	jdff dff_B_YNvCsceP4_2(.din(n910),.dout(w_dff_B_YNvCsceP4_2),.clk(gclk));
	jdff dff_B_Xia3DPRR8_1(.din(n908),.dout(w_dff_B_Xia3DPRR8_1),.clk(gclk));
	jdff dff_A_662e2IZt3_0(.dout(w_n805_0[0]),.din(w_dff_A_662e2IZt3_0),.clk(gclk));
	jdff dff_A_nYbpCc9b3_0(.dout(w_dff_A_662e2IZt3_0),.din(w_dff_A_nYbpCc9b3_0),.clk(gclk));
	jdff dff_A_ThMdp57M7_0(.dout(w_dff_A_nYbpCc9b3_0),.din(w_dff_A_ThMdp57M7_0),.clk(gclk));
	jdff dff_A_kgFBWi1H8_0(.dout(w_dff_A_ThMdp57M7_0),.din(w_dff_A_kgFBWi1H8_0),.clk(gclk));
	jdff dff_A_J2FjpTxz8_0(.dout(w_dff_A_kgFBWi1H8_0),.din(w_dff_A_J2FjpTxz8_0),.clk(gclk));
	jdff dff_A_nJSXpeTJ9_0(.dout(w_dff_A_J2FjpTxz8_0),.din(w_dff_A_nJSXpeTJ9_0),.clk(gclk));
	jdff dff_A_f2sPAGvk7_0(.dout(w_dff_A_nJSXpeTJ9_0),.din(w_dff_A_f2sPAGvk7_0),.clk(gclk));
	jdff dff_A_7r92TQdh3_0(.dout(w_dff_A_f2sPAGvk7_0),.din(w_dff_A_7r92TQdh3_0),.clk(gclk));
	jdff dff_A_efvqtBPX6_0(.dout(w_dff_A_7r92TQdh3_0),.din(w_dff_A_efvqtBPX6_0),.clk(gclk));
	jdff dff_A_NpHji1wM6_0(.dout(w_dff_A_efvqtBPX6_0),.din(w_dff_A_NpHji1wM6_0),.clk(gclk));
	jdff dff_A_jkyacbFs5_0(.dout(w_dff_A_NpHji1wM6_0),.din(w_dff_A_jkyacbFs5_0),.clk(gclk));
	jdff dff_A_4aYeIp7H0_0(.dout(w_dff_A_jkyacbFs5_0),.din(w_dff_A_4aYeIp7H0_0),.clk(gclk));
	jdff dff_A_Q1nZT9NW0_0(.dout(w_dff_A_4aYeIp7H0_0),.din(w_dff_A_Q1nZT9NW0_0),.clk(gclk));
	jdff dff_A_2LBktEPd4_0(.dout(w_dff_A_Q1nZT9NW0_0),.din(w_dff_A_2LBktEPd4_0),.clk(gclk));
	jdff dff_A_RbA0scCG7_0(.dout(w_dff_A_2LBktEPd4_0),.din(w_dff_A_RbA0scCG7_0),.clk(gclk));
	jdff dff_A_LP7iEK6k7_0(.dout(w_dff_A_RbA0scCG7_0),.din(w_dff_A_LP7iEK6k7_0),.clk(gclk));
	jdff dff_A_KMsGdlAA4_0(.dout(w_dff_A_LP7iEK6k7_0),.din(w_dff_A_KMsGdlAA4_0),.clk(gclk));
	jdff dff_A_jwKx4BaT1_0(.dout(w_dff_A_KMsGdlAA4_0),.din(w_dff_A_jwKx4BaT1_0),.clk(gclk));
	jdff dff_A_NesHmd2r2_0(.dout(w_dff_A_jwKx4BaT1_0),.din(w_dff_A_NesHmd2r2_0),.clk(gclk));
	jdff dff_A_eSRf35sg1_0(.dout(w_dff_A_NesHmd2r2_0),.din(w_dff_A_eSRf35sg1_0),.clk(gclk));
	jdff dff_A_mZA5N4Dx4_0(.dout(w_dff_A_eSRf35sg1_0),.din(w_dff_A_mZA5N4Dx4_0),.clk(gclk));
	jdff dff_A_FaVWmzpk7_0(.dout(w_dff_A_mZA5N4Dx4_0),.din(w_dff_A_FaVWmzpk7_0),.clk(gclk));
	jdff dff_A_l2grCAkI0_0(.dout(w_dff_A_FaVWmzpk7_0),.din(w_dff_A_l2grCAkI0_0),.clk(gclk));
	jdff dff_A_vWvCWpLx2_0(.dout(w_dff_A_l2grCAkI0_0),.din(w_dff_A_vWvCWpLx2_0),.clk(gclk));
	jdff dff_A_9TQiNsuW5_0(.dout(w_dff_A_vWvCWpLx2_0),.din(w_dff_A_9TQiNsuW5_0),.clk(gclk));
	jdff dff_A_WzVtAAyB4_0(.dout(w_dff_A_9TQiNsuW5_0),.din(w_dff_A_WzVtAAyB4_0),.clk(gclk));
	jdff dff_A_xWLrdaQV6_0(.dout(w_dff_A_WzVtAAyB4_0),.din(w_dff_A_xWLrdaQV6_0),.clk(gclk));
	jdff dff_A_S3D6GCMz9_0(.dout(w_dff_A_xWLrdaQV6_0),.din(w_dff_A_S3D6GCMz9_0),.clk(gclk));
	jdff dff_A_KGuhiddx0_0(.dout(w_dff_A_S3D6GCMz9_0),.din(w_dff_A_KGuhiddx0_0),.clk(gclk));
	jdff dff_A_NowR9RrP5_0(.dout(w_dff_A_KGuhiddx0_0),.din(w_dff_A_NowR9RrP5_0),.clk(gclk));
	jdff dff_A_yK1ep4SU1_0(.dout(w_dff_A_NowR9RrP5_0),.din(w_dff_A_yK1ep4SU1_0),.clk(gclk));
	jdff dff_A_FlWyKGHC0_0(.dout(w_dff_A_yK1ep4SU1_0),.din(w_dff_A_FlWyKGHC0_0),.clk(gclk));
	jdff dff_A_g7twgXVv7_0(.dout(w_dff_A_FlWyKGHC0_0),.din(w_dff_A_g7twgXVv7_0),.clk(gclk));
	jdff dff_A_SHL8gzUL6_0(.dout(w_dff_A_g7twgXVv7_0),.din(w_dff_A_SHL8gzUL6_0),.clk(gclk));
	jdff dff_A_r2CxQq4M1_1(.dout(w_n904_0[1]),.din(w_dff_A_r2CxQq4M1_1),.clk(gclk));
	jdff dff_A_LjvnUsz49_0(.dout(w_n706_0[0]),.din(w_dff_A_LjvnUsz49_0),.clk(gclk));
	jdff dff_A_79GnhfdT0_0(.dout(w_dff_A_LjvnUsz49_0),.din(w_dff_A_79GnhfdT0_0),.clk(gclk));
	jdff dff_A_pf89cse13_0(.dout(w_dff_A_79GnhfdT0_0),.din(w_dff_A_pf89cse13_0),.clk(gclk));
	jdff dff_A_apu5ctas8_0(.dout(w_dff_A_pf89cse13_0),.din(w_dff_A_apu5ctas8_0),.clk(gclk));
	jdff dff_A_Y44ODO1F3_0(.dout(w_dff_A_apu5ctas8_0),.din(w_dff_A_Y44ODO1F3_0),.clk(gclk));
	jdff dff_A_lqfcvZwT1_0(.dout(w_dff_A_Y44ODO1F3_0),.din(w_dff_A_lqfcvZwT1_0),.clk(gclk));
	jdff dff_A_ap2fhwR85_0(.dout(w_dff_A_lqfcvZwT1_0),.din(w_dff_A_ap2fhwR85_0),.clk(gclk));
	jdff dff_A_NCqsT08l4_0(.dout(w_dff_A_ap2fhwR85_0),.din(w_dff_A_NCqsT08l4_0),.clk(gclk));
	jdff dff_A_X7MAs05s4_0(.dout(w_dff_A_NCqsT08l4_0),.din(w_dff_A_X7MAs05s4_0),.clk(gclk));
	jdff dff_A_vAceU8wQ5_0(.dout(w_dff_A_X7MAs05s4_0),.din(w_dff_A_vAceU8wQ5_0),.clk(gclk));
	jdff dff_A_FuBDexXD0_0(.dout(w_dff_A_vAceU8wQ5_0),.din(w_dff_A_FuBDexXD0_0),.clk(gclk));
	jdff dff_A_f77i4ZKS3_0(.dout(w_dff_A_FuBDexXD0_0),.din(w_dff_A_f77i4ZKS3_0),.clk(gclk));
	jdff dff_A_Vkb2O4x28_0(.dout(w_dff_A_f77i4ZKS3_0),.din(w_dff_A_Vkb2O4x28_0),.clk(gclk));
	jdff dff_A_DoHLIW5U8_0(.dout(w_dff_A_Vkb2O4x28_0),.din(w_dff_A_DoHLIW5U8_0),.clk(gclk));
	jdff dff_A_EOJQe4B41_0(.dout(w_dff_A_DoHLIW5U8_0),.din(w_dff_A_EOJQe4B41_0),.clk(gclk));
	jdff dff_A_xDlzd7Rw4_0(.dout(w_dff_A_EOJQe4B41_0),.din(w_dff_A_xDlzd7Rw4_0),.clk(gclk));
	jdff dff_A_eb5Z8V4x8_0(.dout(w_dff_A_xDlzd7Rw4_0),.din(w_dff_A_eb5Z8V4x8_0),.clk(gclk));
	jdff dff_A_HSdjzxSB4_0(.dout(w_dff_A_eb5Z8V4x8_0),.din(w_dff_A_HSdjzxSB4_0),.clk(gclk));
	jdff dff_A_jxda1fWA3_0(.dout(w_dff_A_HSdjzxSB4_0),.din(w_dff_A_jxda1fWA3_0),.clk(gclk));
	jdff dff_A_9C5Jn2vo2_0(.dout(w_dff_A_jxda1fWA3_0),.din(w_dff_A_9C5Jn2vo2_0),.clk(gclk));
	jdff dff_A_qsUQrKts7_0(.dout(w_dff_A_9C5Jn2vo2_0),.din(w_dff_A_qsUQrKts7_0),.clk(gclk));
	jdff dff_A_gocJm6ip5_0(.dout(w_dff_A_qsUQrKts7_0),.din(w_dff_A_gocJm6ip5_0),.clk(gclk));
	jdff dff_A_0UDK4Hgn9_0(.dout(w_dff_A_gocJm6ip5_0),.din(w_dff_A_0UDK4Hgn9_0),.clk(gclk));
	jdff dff_A_rzs4JHKQ7_0(.dout(w_dff_A_0UDK4Hgn9_0),.din(w_dff_A_rzs4JHKQ7_0),.clk(gclk));
	jdff dff_A_zU3szE2g4_0(.dout(w_dff_A_rzs4JHKQ7_0),.din(w_dff_A_zU3szE2g4_0),.clk(gclk));
	jdff dff_A_r3dRZP5F8_0(.dout(w_dff_A_zU3szE2g4_0),.din(w_dff_A_r3dRZP5F8_0),.clk(gclk));
	jdff dff_A_XvnQLgZ65_0(.dout(w_dff_A_r3dRZP5F8_0),.din(w_dff_A_XvnQLgZ65_0),.clk(gclk));
	jdff dff_A_BGabRieq2_0(.dout(w_dff_A_XvnQLgZ65_0),.din(w_dff_A_BGabRieq2_0),.clk(gclk));
	jdff dff_A_u7MVywNI6_0(.dout(w_dff_A_BGabRieq2_0),.din(w_dff_A_u7MVywNI6_0),.clk(gclk));
	jdff dff_A_J7GUCHDN2_0(.dout(w_dff_A_u7MVywNI6_0),.din(w_dff_A_J7GUCHDN2_0),.clk(gclk));
	jdff dff_A_WWGZUu9N7_0(.dout(w_dff_A_J7GUCHDN2_0),.din(w_dff_A_WWGZUu9N7_0),.clk(gclk));
	jdff dff_A_4rh7ihgJ1_0(.dout(w_dff_A_WWGZUu9N7_0),.din(w_dff_A_4rh7ihgJ1_0),.clk(gclk));
	jdff dff_B_fl0c5mED1_1(.din(n713),.dout(w_dff_B_fl0c5mED1_1),.clk(gclk));
	jdff dff_B_EroCWDUZ0_1(.din(w_dff_B_fl0c5mED1_1),.dout(w_dff_B_EroCWDUZ0_1),.clk(gclk));
	jdff dff_B_BcNIiExZ7_1(.din(w_dff_B_EroCWDUZ0_1),.dout(w_dff_B_BcNIiExZ7_1),.clk(gclk));
	jdff dff_B_FPU74JMr8_1(.din(w_dff_B_BcNIiExZ7_1),.dout(w_dff_B_FPU74JMr8_1),.clk(gclk));
	jdff dff_B_LK183Sg95_1(.din(w_dff_B_FPU74JMr8_1),.dout(w_dff_B_LK183Sg95_1),.clk(gclk));
	jdff dff_B_ihwmrTxG4_1(.din(w_dff_B_LK183Sg95_1),.dout(w_dff_B_ihwmrTxG4_1),.clk(gclk));
	jdff dff_B_9XK5f75c4_1(.din(w_dff_B_ihwmrTxG4_1),.dout(w_dff_B_9XK5f75c4_1),.clk(gclk));
	jdff dff_B_azC47Q5P6_1(.din(w_dff_B_9XK5f75c4_1),.dout(w_dff_B_azC47Q5P6_1),.clk(gclk));
	jdff dff_B_vbp8zN347_1(.din(w_dff_B_azC47Q5P6_1),.dout(w_dff_B_vbp8zN347_1),.clk(gclk));
	jdff dff_B_jufl5Zgt6_1(.din(w_dff_B_vbp8zN347_1),.dout(w_dff_B_jufl5Zgt6_1),.clk(gclk));
	jdff dff_B_o3X9hQLN0_1(.din(w_dff_B_jufl5Zgt6_1),.dout(w_dff_B_o3X9hQLN0_1),.clk(gclk));
	jdff dff_B_dkYp4EWn9_1(.din(w_dff_B_o3X9hQLN0_1),.dout(w_dff_B_dkYp4EWn9_1),.clk(gclk));
	jdff dff_B_tOd8JLdK9_1(.din(w_dff_B_dkYp4EWn9_1),.dout(w_dff_B_tOd8JLdK9_1),.clk(gclk));
	jdff dff_B_hVvAXGU58_1(.din(w_dff_B_tOd8JLdK9_1),.dout(w_dff_B_hVvAXGU58_1),.clk(gclk));
	jdff dff_B_tp0VQJV27_1(.din(w_dff_B_hVvAXGU58_1),.dout(w_dff_B_tp0VQJV27_1),.clk(gclk));
	jdff dff_B_9WzvPrhm1_1(.din(w_dff_B_tp0VQJV27_1),.dout(w_dff_B_9WzvPrhm1_1),.clk(gclk));
	jdff dff_B_L91TH4AG9_1(.din(w_dff_B_9WzvPrhm1_1),.dout(w_dff_B_L91TH4AG9_1),.clk(gclk));
	jdff dff_B_1M9VXOi20_1(.din(w_dff_B_L91TH4AG9_1),.dout(w_dff_B_1M9VXOi20_1),.clk(gclk));
	jdff dff_B_i9uMggk96_1(.din(w_dff_B_1M9VXOi20_1),.dout(w_dff_B_i9uMggk96_1),.clk(gclk));
	jdff dff_B_WkFeOUrA0_1(.din(w_dff_B_i9uMggk96_1),.dout(w_dff_B_WkFeOUrA0_1),.clk(gclk));
	jdff dff_B_xhaK2JqE9_1(.din(w_dff_B_WkFeOUrA0_1),.dout(w_dff_B_xhaK2JqE9_1),.clk(gclk));
	jdff dff_B_n4TMqiaz9_1(.din(w_dff_B_xhaK2JqE9_1),.dout(w_dff_B_n4TMqiaz9_1),.clk(gclk));
	jdff dff_B_T3L0LJUr4_1(.din(w_dff_B_n4TMqiaz9_1),.dout(w_dff_B_T3L0LJUr4_1),.clk(gclk));
	jdff dff_B_Cjp3A2X53_1(.din(w_dff_B_T3L0LJUr4_1),.dout(w_dff_B_Cjp3A2X53_1),.clk(gclk));
	jdff dff_B_Ai2Lm1r26_1(.din(w_dff_B_Cjp3A2X53_1),.dout(w_dff_B_Ai2Lm1r26_1),.clk(gclk));
	jdff dff_B_OAZclFQB9_1(.din(w_dff_B_Ai2Lm1r26_1),.dout(w_dff_B_OAZclFQB9_1),.clk(gclk));
	jdff dff_B_moMqFGDf9_1(.din(w_dff_B_OAZclFQB9_1),.dout(w_dff_B_moMqFGDf9_1),.clk(gclk));
	jdff dff_B_aHmtZ6tl5_1(.din(w_dff_B_moMqFGDf9_1),.dout(w_dff_B_aHmtZ6tl5_1),.clk(gclk));
	jdff dff_B_Xr8BrdpT9_1(.din(w_dff_B_aHmtZ6tl5_1),.dout(w_dff_B_Xr8BrdpT9_1),.clk(gclk));
	jdff dff_A_u0s3Zbqb3_0(.dout(w_n711_0[0]),.din(w_dff_A_u0s3Zbqb3_0),.clk(gclk));
	jdff dff_A_DhJPKj8z5_0(.dout(w_n614_0[0]),.din(w_dff_A_DhJPKj8z5_0),.clk(gclk));
	jdff dff_A_0NuIA5fv0_0(.dout(w_dff_A_DhJPKj8z5_0),.din(w_dff_A_0NuIA5fv0_0),.clk(gclk));
	jdff dff_A_aP1WtKMP3_0(.dout(w_dff_A_0NuIA5fv0_0),.din(w_dff_A_aP1WtKMP3_0),.clk(gclk));
	jdff dff_A_TfCsFiU43_0(.dout(w_dff_A_aP1WtKMP3_0),.din(w_dff_A_TfCsFiU43_0),.clk(gclk));
	jdff dff_A_lrgq5xpY5_0(.dout(w_dff_A_TfCsFiU43_0),.din(w_dff_A_lrgq5xpY5_0),.clk(gclk));
	jdff dff_A_Fmmh8k6N9_0(.dout(w_dff_A_lrgq5xpY5_0),.din(w_dff_A_Fmmh8k6N9_0),.clk(gclk));
	jdff dff_A_BIpxdEPV2_0(.dout(w_dff_A_Fmmh8k6N9_0),.din(w_dff_A_BIpxdEPV2_0),.clk(gclk));
	jdff dff_A_pQMKzbRF3_0(.dout(w_dff_A_BIpxdEPV2_0),.din(w_dff_A_pQMKzbRF3_0),.clk(gclk));
	jdff dff_A_Aolfnmco6_0(.dout(w_dff_A_pQMKzbRF3_0),.din(w_dff_A_Aolfnmco6_0),.clk(gclk));
	jdff dff_A_xVRQm6lv1_0(.dout(w_dff_A_Aolfnmco6_0),.din(w_dff_A_xVRQm6lv1_0),.clk(gclk));
	jdff dff_A_f2ZIWKq99_0(.dout(w_dff_A_xVRQm6lv1_0),.din(w_dff_A_f2ZIWKq99_0),.clk(gclk));
	jdff dff_A_ITW5vLeN9_0(.dout(w_dff_A_f2ZIWKq99_0),.din(w_dff_A_ITW5vLeN9_0),.clk(gclk));
	jdff dff_A_WlwAB7hE0_0(.dout(w_dff_A_ITW5vLeN9_0),.din(w_dff_A_WlwAB7hE0_0),.clk(gclk));
	jdff dff_A_8NxqBm351_0(.dout(w_dff_A_WlwAB7hE0_0),.din(w_dff_A_8NxqBm351_0),.clk(gclk));
	jdff dff_A_eryoXjcz8_0(.dout(w_dff_A_8NxqBm351_0),.din(w_dff_A_eryoXjcz8_0),.clk(gclk));
	jdff dff_A_Z9yh2W5N9_0(.dout(w_dff_A_eryoXjcz8_0),.din(w_dff_A_Z9yh2W5N9_0),.clk(gclk));
	jdff dff_A_lk1UE25t6_0(.dout(w_dff_A_Z9yh2W5N9_0),.din(w_dff_A_lk1UE25t6_0),.clk(gclk));
	jdff dff_A_AXCjBpp53_0(.dout(w_dff_A_lk1UE25t6_0),.din(w_dff_A_AXCjBpp53_0),.clk(gclk));
	jdff dff_A_U4z4fEaq7_0(.dout(w_dff_A_AXCjBpp53_0),.din(w_dff_A_U4z4fEaq7_0),.clk(gclk));
	jdff dff_A_rtaGv1At5_0(.dout(w_dff_A_U4z4fEaq7_0),.din(w_dff_A_rtaGv1At5_0),.clk(gclk));
	jdff dff_A_q5UBzoSI8_0(.dout(w_dff_A_rtaGv1At5_0),.din(w_dff_A_q5UBzoSI8_0),.clk(gclk));
	jdff dff_A_74bJ42Px2_0(.dout(w_dff_A_q5UBzoSI8_0),.din(w_dff_A_74bJ42Px2_0),.clk(gclk));
	jdff dff_A_cKe8MsmW7_0(.dout(w_dff_A_74bJ42Px2_0),.din(w_dff_A_cKe8MsmW7_0),.clk(gclk));
	jdff dff_A_YiKKVe339_0(.dout(w_dff_A_cKe8MsmW7_0),.din(w_dff_A_YiKKVe339_0),.clk(gclk));
	jdff dff_A_YlLS9Huu6_0(.dout(w_dff_A_YiKKVe339_0),.din(w_dff_A_YlLS9Huu6_0),.clk(gclk));
	jdff dff_A_UdzPKHV37_0(.dout(w_dff_A_YlLS9Huu6_0),.din(w_dff_A_UdzPKHV37_0),.clk(gclk));
	jdff dff_A_1j8JjMbh9_0(.dout(w_dff_A_UdzPKHV37_0),.din(w_dff_A_1j8JjMbh9_0),.clk(gclk));
	jdff dff_A_6jxhMHGT2_0(.dout(w_dff_A_1j8JjMbh9_0),.din(w_dff_A_6jxhMHGT2_0),.clk(gclk));
	jdff dff_A_VEaKGW435_0(.dout(w_dff_A_6jxhMHGT2_0),.din(w_dff_A_VEaKGW435_0),.clk(gclk));
	jdff dff_A_RK6NV3yY4_0(.dout(w_dff_A_VEaKGW435_0),.din(w_dff_A_RK6NV3yY4_0),.clk(gclk));
	jdff dff_B_yyVOwNSn6_1(.din(n621),.dout(w_dff_B_yyVOwNSn6_1),.clk(gclk));
	jdff dff_B_kDYN1VUs6_1(.din(w_dff_B_yyVOwNSn6_1),.dout(w_dff_B_kDYN1VUs6_1),.clk(gclk));
	jdff dff_B_pj3Ag8u10_1(.din(w_dff_B_kDYN1VUs6_1),.dout(w_dff_B_pj3Ag8u10_1),.clk(gclk));
	jdff dff_B_kuKkryOB8_1(.din(w_dff_B_pj3Ag8u10_1),.dout(w_dff_B_kuKkryOB8_1),.clk(gclk));
	jdff dff_B_wV6ZTMw41_1(.din(w_dff_B_kuKkryOB8_1),.dout(w_dff_B_wV6ZTMw41_1),.clk(gclk));
	jdff dff_B_zAKn2UZ08_1(.din(w_dff_B_wV6ZTMw41_1),.dout(w_dff_B_zAKn2UZ08_1),.clk(gclk));
	jdff dff_B_njclK8zl3_1(.din(w_dff_B_zAKn2UZ08_1),.dout(w_dff_B_njclK8zl3_1),.clk(gclk));
	jdff dff_B_vPpFkMWL7_1(.din(w_dff_B_njclK8zl3_1),.dout(w_dff_B_vPpFkMWL7_1),.clk(gclk));
	jdff dff_B_dxTpz6Ld8_1(.din(w_dff_B_vPpFkMWL7_1),.dout(w_dff_B_dxTpz6Ld8_1),.clk(gclk));
	jdff dff_B_1ZlObyMt6_1(.din(w_dff_B_dxTpz6Ld8_1),.dout(w_dff_B_1ZlObyMt6_1),.clk(gclk));
	jdff dff_B_pq7aIwPR5_1(.din(w_dff_B_1ZlObyMt6_1),.dout(w_dff_B_pq7aIwPR5_1),.clk(gclk));
	jdff dff_B_sfZo5COr3_1(.din(w_dff_B_pq7aIwPR5_1),.dout(w_dff_B_sfZo5COr3_1),.clk(gclk));
	jdff dff_B_tPDdOh0K9_1(.din(w_dff_B_sfZo5COr3_1),.dout(w_dff_B_tPDdOh0K9_1),.clk(gclk));
	jdff dff_B_xOif8gcl1_1(.din(w_dff_B_tPDdOh0K9_1),.dout(w_dff_B_xOif8gcl1_1),.clk(gclk));
	jdff dff_B_ubcRyYBL4_1(.din(w_dff_B_xOif8gcl1_1),.dout(w_dff_B_ubcRyYBL4_1),.clk(gclk));
	jdff dff_B_dxrBSLmP4_1(.din(w_dff_B_ubcRyYBL4_1),.dout(w_dff_B_dxrBSLmP4_1),.clk(gclk));
	jdff dff_B_nxT1jgfo7_1(.din(w_dff_B_dxrBSLmP4_1),.dout(w_dff_B_nxT1jgfo7_1),.clk(gclk));
	jdff dff_B_neV8O9dC9_1(.din(w_dff_B_nxT1jgfo7_1),.dout(w_dff_B_neV8O9dC9_1),.clk(gclk));
	jdff dff_B_7UaYYAbM1_1(.din(w_dff_B_neV8O9dC9_1),.dout(w_dff_B_7UaYYAbM1_1),.clk(gclk));
	jdff dff_B_Qaf57BRl0_1(.din(w_dff_B_7UaYYAbM1_1),.dout(w_dff_B_Qaf57BRl0_1),.clk(gclk));
	jdff dff_B_18iTE7CW6_1(.din(w_dff_B_Qaf57BRl0_1),.dout(w_dff_B_18iTE7CW6_1),.clk(gclk));
	jdff dff_B_w28BwwaZ8_1(.din(w_dff_B_18iTE7CW6_1),.dout(w_dff_B_w28BwwaZ8_1),.clk(gclk));
	jdff dff_B_k6QZNmAk0_1(.din(w_dff_B_w28BwwaZ8_1),.dout(w_dff_B_k6QZNmAk0_1),.clk(gclk));
	jdff dff_B_rFT5RGUN6_1(.din(w_dff_B_k6QZNmAk0_1),.dout(w_dff_B_rFT5RGUN6_1),.clk(gclk));
	jdff dff_B_DBuZFplD7_1(.din(w_dff_B_rFT5RGUN6_1),.dout(w_dff_B_DBuZFplD7_1),.clk(gclk));
	jdff dff_B_JTC0kpu73_1(.din(w_dff_B_DBuZFplD7_1),.dout(w_dff_B_JTC0kpu73_1),.clk(gclk));
	jdff dff_B_b2d0OJvg0_1(.din(w_dff_B_JTC0kpu73_1),.dout(w_dff_B_b2d0OJvg0_1),.clk(gclk));
	jdff dff_A_wpS1r5Ve3_0(.dout(w_n619_0[0]),.din(w_dff_A_wpS1r5Ve3_0),.clk(gclk));
	jdff dff_A_YA8c7Vsj6_0(.dout(w_n529_0[0]),.din(w_dff_A_YA8c7Vsj6_0),.clk(gclk));
	jdff dff_A_6VICeRBW3_0(.dout(w_dff_A_YA8c7Vsj6_0),.din(w_dff_A_6VICeRBW3_0),.clk(gclk));
	jdff dff_A_Pzz4ffo91_0(.dout(w_dff_A_6VICeRBW3_0),.din(w_dff_A_Pzz4ffo91_0),.clk(gclk));
	jdff dff_A_6LsxZDxU1_0(.dout(w_dff_A_Pzz4ffo91_0),.din(w_dff_A_6LsxZDxU1_0),.clk(gclk));
	jdff dff_A_mstkAnUV8_0(.dout(w_dff_A_6LsxZDxU1_0),.din(w_dff_A_mstkAnUV8_0),.clk(gclk));
	jdff dff_A_dvUsAZYt7_0(.dout(w_dff_A_mstkAnUV8_0),.din(w_dff_A_dvUsAZYt7_0),.clk(gclk));
	jdff dff_A_apH9xc515_0(.dout(w_dff_A_dvUsAZYt7_0),.din(w_dff_A_apH9xc515_0),.clk(gclk));
	jdff dff_A_k5sUWt6F5_0(.dout(w_dff_A_apH9xc515_0),.din(w_dff_A_k5sUWt6F5_0),.clk(gclk));
	jdff dff_A_ZLA3LvBy4_0(.dout(w_dff_A_k5sUWt6F5_0),.din(w_dff_A_ZLA3LvBy4_0),.clk(gclk));
	jdff dff_A_LJdIBqOY4_0(.dout(w_dff_A_ZLA3LvBy4_0),.din(w_dff_A_LJdIBqOY4_0),.clk(gclk));
	jdff dff_A_atpe8yZE1_0(.dout(w_dff_A_LJdIBqOY4_0),.din(w_dff_A_atpe8yZE1_0),.clk(gclk));
	jdff dff_A_nJ1njDy75_0(.dout(w_dff_A_atpe8yZE1_0),.din(w_dff_A_nJ1njDy75_0),.clk(gclk));
	jdff dff_A_XInLPycQ7_0(.dout(w_dff_A_nJ1njDy75_0),.din(w_dff_A_XInLPycQ7_0),.clk(gclk));
	jdff dff_A_lt8uivqi3_0(.dout(w_dff_A_XInLPycQ7_0),.din(w_dff_A_lt8uivqi3_0),.clk(gclk));
	jdff dff_A_8Tm8oo6L4_0(.dout(w_dff_A_lt8uivqi3_0),.din(w_dff_A_8Tm8oo6L4_0),.clk(gclk));
	jdff dff_A_wRK892fu0_0(.dout(w_dff_A_8Tm8oo6L4_0),.din(w_dff_A_wRK892fu0_0),.clk(gclk));
	jdff dff_A_rmczvSi92_0(.dout(w_dff_A_wRK892fu0_0),.din(w_dff_A_rmczvSi92_0),.clk(gclk));
	jdff dff_A_4byYXUiP1_0(.dout(w_dff_A_rmczvSi92_0),.din(w_dff_A_4byYXUiP1_0),.clk(gclk));
	jdff dff_A_eX2ryzXN3_0(.dout(w_dff_A_4byYXUiP1_0),.din(w_dff_A_eX2ryzXN3_0),.clk(gclk));
	jdff dff_A_MJsbTHvp5_0(.dout(w_dff_A_eX2ryzXN3_0),.din(w_dff_A_MJsbTHvp5_0),.clk(gclk));
	jdff dff_A_8nXUk5064_0(.dout(w_dff_A_MJsbTHvp5_0),.din(w_dff_A_8nXUk5064_0),.clk(gclk));
	jdff dff_A_WALeyVol8_0(.dout(w_dff_A_8nXUk5064_0),.din(w_dff_A_WALeyVol8_0),.clk(gclk));
	jdff dff_A_gUgtPafd3_0(.dout(w_dff_A_WALeyVol8_0),.din(w_dff_A_gUgtPafd3_0),.clk(gclk));
	jdff dff_A_mxvlQutG6_0(.dout(w_dff_A_gUgtPafd3_0),.din(w_dff_A_mxvlQutG6_0),.clk(gclk));
	jdff dff_A_7230e3rg5_0(.dout(w_dff_A_mxvlQutG6_0),.din(w_dff_A_7230e3rg5_0),.clk(gclk));
	jdff dff_A_44f0VQ760_0(.dout(w_dff_A_7230e3rg5_0),.din(w_dff_A_44f0VQ760_0),.clk(gclk));
	jdff dff_A_XvAdRIwp2_0(.dout(w_dff_A_44f0VQ760_0),.din(w_dff_A_XvAdRIwp2_0),.clk(gclk));
	jdff dff_A_heUPJXR54_0(.dout(w_dff_A_XvAdRIwp2_0),.din(w_dff_A_heUPJXR54_0),.clk(gclk));
	jdff dff_B_lwbqDVIQ6_1(.din(n536),.dout(w_dff_B_lwbqDVIQ6_1),.clk(gclk));
	jdff dff_B_KFB0YdQh2_1(.din(w_dff_B_lwbqDVIQ6_1),.dout(w_dff_B_KFB0YdQh2_1),.clk(gclk));
	jdff dff_B_25UWo6Kx6_1(.din(w_dff_B_KFB0YdQh2_1),.dout(w_dff_B_25UWo6Kx6_1),.clk(gclk));
	jdff dff_B_x6Xp0fhs8_1(.din(w_dff_B_25UWo6Kx6_1),.dout(w_dff_B_x6Xp0fhs8_1),.clk(gclk));
	jdff dff_B_FwpSVmFo7_1(.din(w_dff_B_x6Xp0fhs8_1),.dout(w_dff_B_FwpSVmFo7_1),.clk(gclk));
	jdff dff_B_swzC9u0u5_1(.din(w_dff_B_FwpSVmFo7_1),.dout(w_dff_B_swzC9u0u5_1),.clk(gclk));
	jdff dff_B_UmpXJIOF1_1(.din(w_dff_B_swzC9u0u5_1),.dout(w_dff_B_UmpXJIOF1_1),.clk(gclk));
	jdff dff_B_LE85dAEu0_1(.din(w_dff_B_UmpXJIOF1_1),.dout(w_dff_B_LE85dAEu0_1),.clk(gclk));
	jdff dff_B_k8Wmwwen9_1(.din(w_dff_B_LE85dAEu0_1),.dout(w_dff_B_k8Wmwwen9_1),.clk(gclk));
	jdff dff_B_8foNXss18_1(.din(w_dff_B_k8Wmwwen9_1),.dout(w_dff_B_8foNXss18_1),.clk(gclk));
	jdff dff_B_5zma2OI19_1(.din(w_dff_B_8foNXss18_1),.dout(w_dff_B_5zma2OI19_1),.clk(gclk));
	jdff dff_B_G3W7TjME8_1(.din(w_dff_B_5zma2OI19_1),.dout(w_dff_B_G3W7TjME8_1),.clk(gclk));
	jdff dff_B_9gqH5NdN3_1(.din(w_dff_B_G3W7TjME8_1),.dout(w_dff_B_9gqH5NdN3_1),.clk(gclk));
	jdff dff_B_J2ZNqNcs7_1(.din(w_dff_B_9gqH5NdN3_1),.dout(w_dff_B_J2ZNqNcs7_1),.clk(gclk));
	jdff dff_B_PK1mKeB32_1(.din(w_dff_B_J2ZNqNcs7_1),.dout(w_dff_B_PK1mKeB32_1),.clk(gclk));
	jdff dff_B_OCowzZ429_1(.din(w_dff_B_PK1mKeB32_1),.dout(w_dff_B_OCowzZ429_1),.clk(gclk));
	jdff dff_B_JtjJyPBd8_1(.din(w_dff_B_OCowzZ429_1),.dout(w_dff_B_JtjJyPBd8_1),.clk(gclk));
	jdff dff_B_17PlxHih2_1(.din(w_dff_B_JtjJyPBd8_1),.dout(w_dff_B_17PlxHih2_1),.clk(gclk));
	jdff dff_B_8Pc8qrVl3_1(.din(w_dff_B_17PlxHih2_1),.dout(w_dff_B_8Pc8qrVl3_1),.clk(gclk));
	jdff dff_B_cUQbM1Lk9_1(.din(w_dff_B_8Pc8qrVl3_1),.dout(w_dff_B_cUQbM1Lk9_1),.clk(gclk));
	jdff dff_B_02DVclHt9_1(.din(w_dff_B_cUQbM1Lk9_1),.dout(w_dff_B_02DVclHt9_1),.clk(gclk));
	jdff dff_B_efRyBIxh2_1(.din(w_dff_B_02DVclHt9_1),.dout(w_dff_B_efRyBIxh2_1),.clk(gclk));
	jdff dff_B_8DI3KBPB1_1(.din(w_dff_B_efRyBIxh2_1),.dout(w_dff_B_8DI3KBPB1_1),.clk(gclk));
	jdff dff_B_xosNsz7v5_1(.din(w_dff_B_8DI3KBPB1_1),.dout(w_dff_B_xosNsz7v5_1),.clk(gclk));
	jdff dff_B_fSWVXiTU0_1(.din(w_dff_B_xosNsz7v5_1),.dout(w_dff_B_fSWVXiTU0_1),.clk(gclk));
	jdff dff_A_XGY45YLI0_0(.dout(w_n534_0[0]),.din(w_dff_A_XGY45YLI0_0),.clk(gclk));
	jdff dff_A_En2GioGH4_0(.dout(w_n451_0[0]),.din(w_dff_A_En2GioGH4_0),.clk(gclk));
	jdff dff_A_GwkOOmRj8_0(.dout(w_dff_A_En2GioGH4_0),.din(w_dff_A_GwkOOmRj8_0),.clk(gclk));
	jdff dff_A_ae0vzBCp7_0(.dout(w_dff_A_GwkOOmRj8_0),.din(w_dff_A_ae0vzBCp7_0),.clk(gclk));
	jdff dff_A_k3lXcdZK0_0(.dout(w_dff_A_ae0vzBCp7_0),.din(w_dff_A_k3lXcdZK0_0),.clk(gclk));
	jdff dff_A_lw0rnrfI6_0(.dout(w_dff_A_k3lXcdZK0_0),.din(w_dff_A_lw0rnrfI6_0),.clk(gclk));
	jdff dff_A_D5XXFsMe3_0(.dout(w_dff_A_lw0rnrfI6_0),.din(w_dff_A_D5XXFsMe3_0),.clk(gclk));
	jdff dff_A_YQ1GHwYF8_0(.dout(w_dff_A_D5XXFsMe3_0),.din(w_dff_A_YQ1GHwYF8_0),.clk(gclk));
	jdff dff_A_F2M2hjAQ7_0(.dout(w_dff_A_YQ1GHwYF8_0),.din(w_dff_A_F2M2hjAQ7_0),.clk(gclk));
	jdff dff_A_0t9o09RF1_0(.dout(w_dff_A_F2M2hjAQ7_0),.din(w_dff_A_0t9o09RF1_0),.clk(gclk));
	jdff dff_A_cqfiSJAM6_0(.dout(w_dff_A_0t9o09RF1_0),.din(w_dff_A_cqfiSJAM6_0),.clk(gclk));
	jdff dff_A_eJSQsWRa4_0(.dout(w_dff_A_cqfiSJAM6_0),.din(w_dff_A_eJSQsWRa4_0),.clk(gclk));
	jdff dff_A_c79lqtLe4_0(.dout(w_dff_A_eJSQsWRa4_0),.din(w_dff_A_c79lqtLe4_0),.clk(gclk));
	jdff dff_A_pobWB3Xf6_0(.dout(w_dff_A_c79lqtLe4_0),.din(w_dff_A_pobWB3Xf6_0),.clk(gclk));
	jdff dff_A_rjG6rSI43_0(.dout(w_dff_A_pobWB3Xf6_0),.din(w_dff_A_rjG6rSI43_0),.clk(gclk));
	jdff dff_A_ZFU39aD09_0(.dout(w_dff_A_rjG6rSI43_0),.din(w_dff_A_ZFU39aD09_0),.clk(gclk));
	jdff dff_A_zLwuAHox7_0(.dout(w_dff_A_ZFU39aD09_0),.din(w_dff_A_zLwuAHox7_0),.clk(gclk));
	jdff dff_A_7o1RRmWI5_0(.dout(w_dff_A_zLwuAHox7_0),.din(w_dff_A_7o1RRmWI5_0),.clk(gclk));
	jdff dff_A_5ncj4DcK0_0(.dout(w_dff_A_7o1RRmWI5_0),.din(w_dff_A_5ncj4DcK0_0),.clk(gclk));
	jdff dff_A_SosMuBux0_0(.dout(w_dff_A_5ncj4DcK0_0),.din(w_dff_A_SosMuBux0_0),.clk(gclk));
	jdff dff_A_BxPeyYXQ6_0(.dout(w_dff_A_SosMuBux0_0),.din(w_dff_A_BxPeyYXQ6_0),.clk(gclk));
	jdff dff_A_daNuyowd4_0(.dout(w_dff_A_BxPeyYXQ6_0),.din(w_dff_A_daNuyowd4_0),.clk(gclk));
	jdff dff_A_1AsRAIib1_0(.dout(w_dff_A_daNuyowd4_0),.din(w_dff_A_1AsRAIib1_0),.clk(gclk));
	jdff dff_A_c8Fuw6xd7_0(.dout(w_dff_A_1AsRAIib1_0),.din(w_dff_A_c8Fuw6xd7_0),.clk(gclk));
	jdff dff_A_yzoKD03O9_0(.dout(w_dff_A_c8Fuw6xd7_0),.din(w_dff_A_yzoKD03O9_0),.clk(gclk));
	jdff dff_A_m9b5JjKC8_0(.dout(w_dff_A_yzoKD03O9_0),.din(w_dff_A_m9b5JjKC8_0),.clk(gclk));
	jdff dff_A_oHHeRJzx3_0(.dout(w_dff_A_m9b5JjKC8_0),.din(w_dff_A_oHHeRJzx3_0),.clk(gclk));
	jdff dff_B_autOpJMY4_1(.din(n458),.dout(w_dff_B_autOpJMY4_1),.clk(gclk));
	jdff dff_B_iwAisoDV7_1(.din(w_dff_B_autOpJMY4_1),.dout(w_dff_B_iwAisoDV7_1),.clk(gclk));
	jdff dff_B_1UHCkcWA5_1(.din(w_dff_B_iwAisoDV7_1),.dout(w_dff_B_1UHCkcWA5_1),.clk(gclk));
	jdff dff_B_U8bbVaYg7_1(.din(w_dff_B_1UHCkcWA5_1),.dout(w_dff_B_U8bbVaYg7_1),.clk(gclk));
	jdff dff_B_5wIgPplJ8_1(.din(w_dff_B_U8bbVaYg7_1),.dout(w_dff_B_5wIgPplJ8_1),.clk(gclk));
	jdff dff_B_EgztDzRY5_1(.din(w_dff_B_5wIgPplJ8_1),.dout(w_dff_B_EgztDzRY5_1),.clk(gclk));
	jdff dff_B_rLWf9Khn9_1(.din(w_dff_B_EgztDzRY5_1),.dout(w_dff_B_rLWf9Khn9_1),.clk(gclk));
	jdff dff_B_bioYfxHb3_1(.din(w_dff_B_rLWf9Khn9_1),.dout(w_dff_B_bioYfxHb3_1),.clk(gclk));
	jdff dff_B_Y8J8XSz76_1(.din(w_dff_B_bioYfxHb3_1),.dout(w_dff_B_Y8J8XSz76_1),.clk(gclk));
	jdff dff_B_30qpmITL7_1(.din(w_dff_B_Y8J8XSz76_1),.dout(w_dff_B_30qpmITL7_1),.clk(gclk));
	jdff dff_B_4uRb8raq6_1(.din(w_dff_B_30qpmITL7_1),.dout(w_dff_B_4uRb8raq6_1),.clk(gclk));
	jdff dff_B_pLGfKK440_1(.din(w_dff_B_4uRb8raq6_1),.dout(w_dff_B_pLGfKK440_1),.clk(gclk));
	jdff dff_B_GiH5w1Fx3_1(.din(w_dff_B_pLGfKK440_1),.dout(w_dff_B_GiH5w1Fx3_1),.clk(gclk));
	jdff dff_B_iMZeQKvo0_1(.din(w_dff_B_GiH5w1Fx3_1),.dout(w_dff_B_iMZeQKvo0_1),.clk(gclk));
	jdff dff_B_oWPvb8HD3_1(.din(w_dff_B_iMZeQKvo0_1),.dout(w_dff_B_oWPvb8HD3_1),.clk(gclk));
	jdff dff_B_2eJzP2Ax9_1(.din(w_dff_B_oWPvb8HD3_1),.dout(w_dff_B_2eJzP2Ax9_1),.clk(gclk));
	jdff dff_B_dcjT6elr3_1(.din(w_dff_B_2eJzP2Ax9_1),.dout(w_dff_B_dcjT6elr3_1),.clk(gclk));
	jdff dff_B_lsJY1KAu1_1(.din(w_dff_B_dcjT6elr3_1),.dout(w_dff_B_lsJY1KAu1_1),.clk(gclk));
	jdff dff_B_L9tQ05x56_1(.din(w_dff_B_lsJY1KAu1_1),.dout(w_dff_B_L9tQ05x56_1),.clk(gclk));
	jdff dff_B_eOqGNY3X9_1(.din(w_dff_B_L9tQ05x56_1),.dout(w_dff_B_eOqGNY3X9_1),.clk(gclk));
	jdff dff_B_E986NeAS8_1(.din(w_dff_B_eOqGNY3X9_1),.dout(w_dff_B_E986NeAS8_1),.clk(gclk));
	jdff dff_B_hwTqp9gH6_1(.din(w_dff_B_E986NeAS8_1),.dout(w_dff_B_hwTqp9gH6_1),.clk(gclk));
	jdff dff_B_ertSK6Qe6_1(.din(w_dff_B_hwTqp9gH6_1),.dout(w_dff_B_ertSK6Qe6_1),.clk(gclk));
	jdff dff_A_u8VsDPPC5_0(.dout(w_n456_0[0]),.din(w_dff_A_u8VsDPPC5_0),.clk(gclk));
	jdff dff_A_ZXw6WQGz4_0(.dout(w_n380_0[0]),.din(w_dff_A_ZXw6WQGz4_0),.clk(gclk));
	jdff dff_A_VOZr7sxY7_0(.dout(w_dff_A_ZXw6WQGz4_0),.din(w_dff_A_VOZr7sxY7_0),.clk(gclk));
	jdff dff_A_HBU1kEVA5_0(.dout(w_dff_A_VOZr7sxY7_0),.din(w_dff_A_HBU1kEVA5_0),.clk(gclk));
	jdff dff_A_3bS3gjp98_0(.dout(w_dff_A_HBU1kEVA5_0),.din(w_dff_A_3bS3gjp98_0),.clk(gclk));
	jdff dff_A_1OXc49AO6_0(.dout(w_dff_A_3bS3gjp98_0),.din(w_dff_A_1OXc49AO6_0),.clk(gclk));
	jdff dff_A_hoFuVvjh6_0(.dout(w_dff_A_1OXc49AO6_0),.din(w_dff_A_hoFuVvjh6_0),.clk(gclk));
	jdff dff_A_DOmHUwHf4_0(.dout(w_dff_A_hoFuVvjh6_0),.din(w_dff_A_DOmHUwHf4_0),.clk(gclk));
	jdff dff_A_jw2VlL2N9_0(.dout(w_dff_A_DOmHUwHf4_0),.din(w_dff_A_jw2VlL2N9_0),.clk(gclk));
	jdff dff_A_Gb0DUAz90_0(.dout(w_dff_A_jw2VlL2N9_0),.din(w_dff_A_Gb0DUAz90_0),.clk(gclk));
	jdff dff_A_gSuGt7599_0(.dout(w_dff_A_Gb0DUAz90_0),.din(w_dff_A_gSuGt7599_0),.clk(gclk));
	jdff dff_A_dmdBv8N27_0(.dout(w_dff_A_gSuGt7599_0),.din(w_dff_A_dmdBv8N27_0),.clk(gclk));
	jdff dff_A_f9nTi06l8_0(.dout(w_dff_A_dmdBv8N27_0),.din(w_dff_A_f9nTi06l8_0),.clk(gclk));
	jdff dff_A_YlYbNnYc0_0(.dout(w_dff_A_f9nTi06l8_0),.din(w_dff_A_YlYbNnYc0_0),.clk(gclk));
	jdff dff_A_HLjgf71D3_0(.dout(w_dff_A_YlYbNnYc0_0),.din(w_dff_A_HLjgf71D3_0),.clk(gclk));
	jdff dff_A_kUyvyLAY3_0(.dout(w_dff_A_HLjgf71D3_0),.din(w_dff_A_kUyvyLAY3_0),.clk(gclk));
	jdff dff_A_omMqnCze0_0(.dout(w_dff_A_kUyvyLAY3_0),.din(w_dff_A_omMqnCze0_0),.clk(gclk));
	jdff dff_A_2djNMAqW6_0(.dout(w_dff_A_omMqnCze0_0),.din(w_dff_A_2djNMAqW6_0),.clk(gclk));
	jdff dff_A_q111pifi0_0(.dout(w_dff_A_2djNMAqW6_0),.din(w_dff_A_q111pifi0_0),.clk(gclk));
	jdff dff_A_VEnxGjTL4_0(.dout(w_dff_A_q111pifi0_0),.din(w_dff_A_VEnxGjTL4_0),.clk(gclk));
	jdff dff_A_62OX3wJD5_0(.dout(w_dff_A_VEnxGjTL4_0),.din(w_dff_A_62OX3wJD5_0),.clk(gclk));
	jdff dff_A_d1ul7Iot6_0(.dout(w_dff_A_62OX3wJD5_0),.din(w_dff_A_d1ul7Iot6_0),.clk(gclk));
	jdff dff_A_jzHLlFiT5_0(.dout(w_dff_A_d1ul7Iot6_0),.din(w_dff_A_jzHLlFiT5_0),.clk(gclk));
	jdff dff_A_S2BPgjId0_0(.dout(w_dff_A_jzHLlFiT5_0),.din(w_dff_A_S2BPgjId0_0),.clk(gclk));
	jdff dff_A_eEk6Vttx5_0(.dout(w_dff_A_S2BPgjId0_0),.din(w_dff_A_eEk6Vttx5_0),.clk(gclk));
	jdff dff_B_ZBaLs8Xt5_1(.din(n387),.dout(w_dff_B_ZBaLs8Xt5_1),.clk(gclk));
	jdff dff_B_5OhO8aqw2_1(.din(w_dff_B_ZBaLs8Xt5_1),.dout(w_dff_B_5OhO8aqw2_1),.clk(gclk));
	jdff dff_B_uKNdESmR9_1(.din(w_dff_B_5OhO8aqw2_1),.dout(w_dff_B_uKNdESmR9_1),.clk(gclk));
	jdff dff_B_a2bjLhg20_1(.din(w_dff_B_uKNdESmR9_1),.dout(w_dff_B_a2bjLhg20_1),.clk(gclk));
	jdff dff_B_mUUNlJ0V1_1(.din(w_dff_B_a2bjLhg20_1),.dout(w_dff_B_mUUNlJ0V1_1),.clk(gclk));
	jdff dff_B_xWGuQY4H3_1(.din(w_dff_B_mUUNlJ0V1_1),.dout(w_dff_B_xWGuQY4H3_1),.clk(gclk));
	jdff dff_B_eFuyN7178_1(.din(w_dff_B_xWGuQY4H3_1),.dout(w_dff_B_eFuyN7178_1),.clk(gclk));
	jdff dff_B_LzCfgZce0_1(.din(w_dff_B_eFuyN7178_1),.dout(w_dff_B_LzCfgZce0_1),.clk(gclk));
	jdff dff_B_klKHjjHP8_1(.din(w_dff_B_LzCfgZce0_1),.dout(w_dff_B_klKHjjHP8_1),.clk(gclk));
	jdff dff_B_q5cT0LaK9_1(.din(w_dff_B_klKHjjHP8_1),.dout(w_dff_B_q5cT0LaK9_1),.clk(gclk));
	jdff dff_B_jLIAHJEB4_1(.din(w_dff_B_q5cT0LaK9_1),.dout(w_dff_B_jLIAHJEB4_1),.clk(gclk));
	jdff dff_B_40Rni9Ms8_1(.din(w_dff_B_jLIAHJEB4_1),.dout(w_dff_B_40Rni9Ms8_1),.clk(gclk));
	jdff dff_B_7sjyTkwd0_1(.din(w_dff_B_40Rni9Ms8_1),.dout(w_dff_B_7sjyTkwd0_1),.clk(gclk));
	jdff dff_B_I9lAXt8m1_1(.din(w_dff_B_7sjyTkwd0_1),.dout(w_dff_B_I9lAXt8m1_1),.clk(gclk));
	jdff dff_B_tF5ARYye3_1(.din(w_dff_B_I9lAXt8m1_1),.dout(w_dff_B_tF5ARYye3_1),.clk(gclk));
	jdff dff_B_cuCAjS7Y9_1(.din(w_dff_B_tF5ARYye3_1),.dout(w_dff_B_cuCAjS7Y9_1),.clk(gclk));
	jdff dff_B_TTquGkNp2_1(.din(w_dff_B_cuCAjS7Y9_1),.dout(w_dff_B_TTquGkNp2_1),.clk(gclk));
	jdff dff_B_XurUm3wt5_1(.din(w_dff_B_TTquGkNp2_1),.dout(w_dff_B_XurUm3wt5_1),.clk(gclk));
	jdff dff_B_BdRZzR443_1(.din(w_dff_B_XurUm3wt5_1),.dout(w_dff_B_BdRZzR443_1),.clk(gclk));
	jdff dff_B_lcf8fmva2_1(.din(w_dff_B_BdRZzR443_1),.dout(w_dff_B_lcf8fmva2_1),.clk(gclk));
	jdff dff_B_VJscNDj46_1(.din(w_dff_B_lcf8fmva2_1),.dout(w_dff_B_VJscNDj46_1),.clk(gclk));
	jdff dff_A_UPGQO3ku6_0(.dout(w_n385_0[0]),.din(w_dff_A_UPGQO3ku6_0),.clk(gclk));
	jdff dff_B_YcJUKzoX3_2(.din(n385),.dout(w_dff_B_YcJUKzoX3_2),.clk(gclk));
	jdff dff_B_BgOGxSfx7_2(.din(w_dff_B_YcJUKzoX3_2),.dout(w_dff_B_BgOGxSfx7_2),.clk(gclk));
	jdff dff_B_WvtuT2Pi5_2(.din(w_dff_B_BgOGxSfx7_2),.dout(w_dff_B_WvtuT2Pi5_2),.clk(gclk));
	jdff dff_A_ODBUwlKM2_0(.dout(w_n317_0[0]),.din(w_dff_A_ODBUwlKM2_0),.clk(gclk));
	jdff dff_A_kuRBZquW6_0(.dout(w_dff_A_ODBUwlKM2_0),.din(w_dff_A_kuRBZquW6_0),.clk(gclk));
	jdff dff_A_RnAKYu0I5_0(.dout(w_dff_A_kuRBZquW6_0),.din(w_dff_A_RnAKYu0I5_0),.clk(gclk));
	jdff dff_A_vQIWDP8O7_0(.dout(w_dff_A_RnAKYu0I5_0),.din(w_dff_A_vQIWDP8O7_0),.clk(gclk));
	jdff dff_A_88dQwK2C2_0(.dout(w_dff_A_vQIWDP8O7_0),.din(w_dff_A_88dQwK2C2_0),.clk(gclk));
	jdff dff_A_O2Z6KUF80_0(.dout(w_dff_A_88dQwK2C2_0),.din(w_dff_A_O2Z6KUF80_0),.clk(gclk));
	jdff dff_A_zSQSs7UD4_0(.dout(w_dff_A_O2Z6KUF80_0),.din(w_dff_A_zSQSs7UD4_0),.clk(gclk));
	jdff dff_A_X7woO4tv3_0(.dout(w_dff_A_zSQSs7UD4_0),.din(w_dff_A_X7woO4tv3_0),.clk(gclk));
	jdff dff_A_H463M3154_0(.dout(w_dff_A_X7woO4tv3_0),.din(w_dff_A_H463M3154_0),.clk(gclk));
	jdff dff_A_EvwQHDzA9_0(.dout(w_dff_A_H463M3154_0),.din(w_dff_A_EvwQHDzA9_0),.clk(gclk));
	jdff dff_A_oRhAsIip2_0(.dout(w_dff_A_EvwQHDzA9_0),.din(w_dff_A_oRhAsIip2_0),.clk(gclk));
	jdff dff_A_zvqnwvqG4_0(.dout(w_dff_A_oRhAsIip2_0),.din(w_dff_A_zvqnwvqG4_0),.clk(gclk));
	jdff dff_A_ZxMd2Zpg2_0(.dout(w_dff_A_zvqnwvqG4_0),.din(w_dff_A_ZxMd2Zpg2_0),.clk(gclk));
	jdff dff_A_IybbEaTi6_0(.dout(w_dff_A_ZxMd2Zpg2_0),.din(w_dff_A_IybbEaTi6_0),.clk(gclk));
	jdff dff_A_2mo7jEbm9_0(.dout(w_dff_A_IybbEaTi6_0),.din(w_dff_A_2mo7jEbm9_0),.clk(gclk));
	jdff dff_A_W3pAHDV28_0(.dout(w_dff_A_2mo7jEbm9_0),.din(w_dff_A_W3pAHDV28_0),.clk(gclk));
	jdff dff_A_wYQWRqgR0_0(.dout(w_dff_A_W3pAHDV28_0),.din(w_dff_A_wYQWRqgR0_0),.clk(gclk));
	jdff dff_A_Vf3Vxb8B9_0(.dout(w_dff_A_wYQWRqgR0_0),.din(w_dff_A_Vf3Vxb8B9_0),.clk(gclk));
	jdff dff_A_hreXLba73_0(.dout(w_dff_A_Vf3Vxb8B9_0),.din(w_dff_A_hreXLba73_0),.clk(gclk));
	jdff dff_B_ppvBdmk69_1(.din(n324),.dout(w_dff_B_ppvBdmk69_1),.clk(gclk));
	jdff dff_B_wGq0fBei3_1(.din(w_dff_B_ppvBdmk69_1),.dout(w_dff_B_wGq0fBei3_1),.clk(gclk));
	jdff dff_B_52mRj8BX4_1(.din(w_dff_B_wGq0fBei3_1),.dout(w_dff_B_52mRj8BX4_1),.clk(gclk));
	jdff dff_B_EyZmbKQn1_1(.din(w_dff_B_52mRj8BX4_1),.dout(w_dff_B_EyZmbKQn1_1),.clk(gclk));
	jdff dff_B_Ty4v1lhC6_1(.din(w_dff_B_EyZmbKQn1_1),.dout(w_dff_B_Ty4v1lhC6_1),.clk(gclk));
	jdff dff_B_X6UfdxlN6_1(.din(w_dff_B_Ty4v1lhC6_1),.dout(w_dff_B_X6UfdxlN6_1),.clk(gclk));
	jdff dff_B_OPTo0SHl1_1(.din(w_dff_B_X6UfdxlN6_1),.dout(w_dff_B_OPTo0SHl1_1),.clk(gclk));
	jdff dff_B_nJElXwyf0_1(.din(w_dff_B_OPTo0SHl1_1),.dout(w_dff_B_nJElXwyf0_1),.clk(gclk));
	jdff dff_B_oAtWTKTZ8_1(.din(w_dff_B_nJElXwyf0_1),.dout(w_dff_B_oAtWTKTZ8_1),.clk(gclk));
	jdff dff_B_fDUpqPth8_1(.din(w_dff_B_oAtWTKTZ8_1),.dout(w_dff_B_fDUpqPth8_1),.clk(gclk));
	jdff dff_B_PWiVRgRp6_1(.din(w_dff_B_fDUpqPth8_1),.dout(w_dff_B_PWiVRgRp6_1),.clk(gclk));
	jdff dff_B_FfGhO3UM8_1(.din(w_dff_B_PWiVRgRp6_1),.dout(w_dff_B_FfGhO3UM8_1),.clk(gclk));
	jdff dff_B_Kx8lPyYI3_1(.din(w_dff_B_FfGhO3UM8_1),.dout(w_dff_B_Kx8lPyYI3_1),.clk(gclk));
	jdff dff_B_BvgUhpIb0_1(.din(w_dff_B_Kx8lPyYI3_1),.dout(w_dff_B_BvgUhpIb0_1),.clk(gclk));
	jdff dff_B_nRx4sBmY5_1(.din(w_dff_B_BvgUhpIb0_1),.dout(w_dff_B_nRx4sBmY5_1),.clk(gclk));
	jdff dff_B_J2iYhzFI2_1(.din(w_dff_B_nRx4sBmY5_1),.dout(w_dff_B_J2iYhzFI2_1),.clk(gclk));
	jdff dff_A_tA5PPiBy4_0(.dout(w_n322_0[0]),.din(w_dff_A_tA5PPiBy4_0),.clk(gclk));
	jdff dff_A_unjFYYcQ8_0(.dout(w_n261_0[0]),.din(w_dff_A_unjFYYcQ8_0),.clk(gclk));
	jdff dff_A_nVzotmll3_0(.dout(w_dff_A_unjFYYcQ8_0),.din(w_dff_A_nVzotmll3_0),.clk(gclk));
	jdff dff_A_SMECIaB48_0(.dout(w_dff_A_nVzotmll3_0),.din(w_dff_A_SMECIaB48_0),.clk(gclk));
	jdff dff_A_yOxCL8S28_0(.dout(w_dff_A_SMECIaB48_0),.din(w_dff_A_yOxCL8S28_0),.clk(gclk));
	jdff dff_A_z3DnaPuo7_0(.dout(w_dff_A_yOxCL8S28_0),.din(w_dff_A_z3DnaPuo7_0),.clk(gclk));
	jdff dff_A_2ipbUAOX1_0(.dout(w_dff_A_z3DnaPuo7_0),.din(w_dff_A_2ipbUAOX1_0),.clk(gclk));
	jdff dff_A_NyWKRBh69_0(.dout(w_dff_A_2ipbUAOX1_0),.din(w_dff_A_NyWKRBh69_0),.clk(gclk));
	jdff dff_A_puRTLCSS5_0(.dout(w_dff_A_NyWKRBh69_0),.din(w_dff_A_puRTLCSS5_0),.clk(gclk));
	jdff dff_A_pvox5kaB9_0(.dout(w_dff_A_puRTLCSS5_0),.din(w_dff_A_pvox5kaB9_0),.clk(gclk));
	jdff dff_A_2WKantat9_0(.dout(w_dff_A_pvox5kaB9_0),.din(w_dff_A_2WKantat9_0),.clk(gclk));
	jdff dff_A_AnYNbJGs3_0(.dout(w_dff_A_2WKantat9_0),.din(w_dff_A_AnYNbJGs3_0),.clk(gclk));
	jdff dff_A_01AAbO2o1_0(.dout(w_dff_A_AnYNbJGs3_0),.din(w_dff_A_01AAbO2o1_0),.clk(gclk));
	jdff dff_A_N8kmsmrQ9_0(.dout(w_dff_A_01AAbO2o1_0),.din(w_dff_A_N8kmsmrQ9_0),.clk(gclk));
	jdff dff_A_taOp7IB92_0(.dout(w_dff_A_N8kmsmrQ9_0),.din(w_dff_A_taOp7IB92_0),.clk(gclk));
	jdff dff_A_nkWJqKJO7_0(.dout(w_dff_A_taOp7IB92_0),.din(w_dff_A_nkWJqKJO7_0),.clk(gclk));
	jdff dff_A_xtxI1w8u9_0(.dout(w_dff_A_nkWJqKJO7_0),.din(w_dff_A_xtxI1w8u9_0),.clk(gclk));
	jdff dff_A_a0Q0MiLY4_0(.dout(w_dff_A_xtxI1w8u9_0),.din(w_dff_A_a0Q0MiLY4_0),.clk(gclk));
	jdff dff_B_wZLPf5rD3_1(.din(n268),.dout(w_dff_B_wZLPf5rD3_1),.clk(gclk));
	jdff dff_B_VgA1fXqw7_1(.din(w_dff_B_wZLPf5rD3_1),.dout(w_dff_B_VgA1fXqw7_1),.clk(gclk));
	jdff dff_B_6NwTz5RD3_1(.din(w_dff_B_VgA1fXqw7_1),.dout(w_dff_B_6NwTz5RD3_1),.clk(gclk));
	jdff dff_B_R5ILRlRx9_1(.din(w_dff_B_6NwTz5RD3_1),.dout(w_dff_B_R5ILRlRx9_1),.clk(gclk));
	jdff dff_B_zyrAS5QZ4_1(.din(w_dff_B_R5ILRlRx9_1),.dout(w_dff_B_zyrAS5QZ4_1),.clk(gclk));
	jdff dff_B_5RJaNZTX0_1(.din(w_dff_B_zyrAS5QZ4_1),.dout(w_dff_B_5RJaNZTX0_1),.clk(gclk));
	jdff dff_B_bcV2UJjf4_1(.din(w_dff_B_5RJaNZTX0_1),.dout(w_dff_B_bcV2UJjf4_1),.clk(gclk));
	jdff dff_B_tLbFtjrV9_1(.din(w_dff_B_bcV2UJjf4_1),.dout(w_dff_B_tLbFtjrV9_1),.clk(gclk));
	jdff dff_B_Nncg7cwm4_1(.din(w_dff_B_tLbFtjrV9_1),.dout(w_dff_B_Nncg7cwm4_1),.clk(gclk));
	jdff dff_B_AdnQVUDQ9_1(.din(w_dff_B_Nncg7cwm4_1),.dout(w_dff_B_AdnQVUDQ9_1),.clk(gclk));
	jdff dff_B_FJjUJS5k8_1(.din(w_dff_B_AdnQVUDQ9_1),.dout(w_dff_B_FJjUJS5k8_1),.clk(gclk));
	jdff dff_B_LRnOdHqb5_1(.din(w_dff_B_FJjUJS5k8_1),.dout(w_dff_B_LRnOdHqb5_1),.clk(gclk));
	jdff dff_B_yMMzxuTT9_1(.din(w_dff_B_LRnOdHqb5_1),.dout(w_dff_B_yMMzxuTT9_1),.clk(gclk));
	jdff dff_B_hp4iNseb0_1(.din(w_dff_B_yMMzxuTT9_1),.dout(w_dff_B_hp4iNseb0_1),.clk(gclk));
	jdff dff_A_GJdiBsWB7_0(.dout(w_n266_0[0]),.din(w_dff_A_GJdiBsWB7_0),.clk(gclk));
	jdff dff_A_5EXzJLuH3_0(.dout(w_n212_0[0]),.din(w_dff_A_5EXzJLuH3_0),.clk(gclk));
	jdff dff_A_22WQMr4n0_0(.dout(w_dff_A_5EXzJLuH3_0),.din(w_dff_A_22WQMr4n0_0),.clk(gclk));
	jdff dff_A_JaudKe7w0_0(.dout(w_dff_A_22WQMr4n0_0),.din(w_dff_A_JaudKe7w0_0),.clk(gclk));
	jdff dff_A_Rp14fa114_0(.dout(w_dff_A_JaudKe7w0_0),.din(w_dff_A_Rp14fa114_0),.clk(gclk));
	jdff dff_A_dizxUtmd9_0(.dout(w_dff_A_Rp14fa114_0),.din(w_dff_A_dizxUtmd9_0),.clk(gclk));
	jdff dff_A_dxVUt8yw9_0(.dout(w_dff_A_dizxUtmd9_0),.din(w_dff_A_dxVUt8yw9_0),.clk(gclk));
	jdff dff_A_vNmnKIdx4_0(.dout(w_dff_A_dxVUt8yw9_0),.din(w_dff_A_vNmnKIdx4_0),.clk(gclk));
	jdff dff_A_e40IayJq1_0(.dout(w_dff_A_vNmnKIdx4_0),.din(w_dff_A_e40IayJq1_0),.clk(gclk));
	jdff dff_A_70k8EJs98_0(.dout(w_dff_A_e40IayJq1_0),.din(w_dff_A_70k8EJs98_0),.clk(gclk));
	jdff dff_A_8QRVLjO96_0(.dout(w_dff_A_70k8EJs98_0),.din(w_dff_A_8QRVLjO96_0),.clk(gclk));
	jdff dff_A_pPh0vQUz9_0(.dout(w_dff_A_8QRVLjO96_0),.din(w_dff_A_pPh0vQUz9_0),.clk(gclk));
	jdff dff_A_i338GVR02_0(.dout(w_dff_A_pPh0vQUz9_0),.din(w_dff_A_i338GVR02_0),.clk(gclk));
	jdff dff_A_69oAD4ky3_0(.dout(w_dff_A_i338GVR02_0),.din(w_dff_A_69oAD4ky3_0),.clk(gclk));
	jdff dff_A_ZZzzjOXd1_0(.dout(w_dff_A_69oAD4ky3_0),.din(w_dff_A_ZZzzjOXd1_0),.clk(gclk));
	jdff dff_A_EEibSwoO2_0(.dout(w_dff_A_ZZzzjOXd1_0),.din(w_dff_A_EEibSwoO2_0),.clk(gclk));
	jdff dff_B_ehgFbZM29_1(.din(n219),.dout(w_dff_B_ehgFbZM29_1),.clk(gclk));
	jdff dff_B_CfPz1sW61_1(.din(w_dff_B_ehgFbZM29_1),.dout(w_dff_B_CfPz1sW61_1),.clk(gclk));
	jdff dff_B_HQwbsi2q9_1(.din(w_dff_B_CfPz1sW61_1),.dout(w_dff_B_HQwbsi2q9_1),.clk(gclk));
	jdff dff_B_uGVUTUZu2_1(.din(w_dff_B_HQwbsi2q9_1),.dout(w_dff_B_uGVUTUZu2_1),.clk(gclk));
	jdff dff_B_I0bJqcBs1_1(.din(w_dff_B_uGVUTUZu2_1),.dout(w_dff_B_I0bJqcBs1_1),.clk(gclk));
	jdff dff_B_mhJJuICq2_1(.din(w_dff_B_I0bJqcBs1_1),.dout(w_dff_B_mhJJuICq2_1),.clk(gclk));
	jdff dff_B_3fkMhPZL9_1(.din(w_dff_B_mhJJuICq2_1),.dout(w_dff_B_3fkMhPZL9_1),.clk(gclk));
	jdff dff_B_sVqsQlWz2_1(.din(w_dff_B_3fkMhPZL9_1),.dout(w_dff_B_sVqsQlWz2_1),.clk(gclk));
	jdff dff_B_2qC9ernC1_1(.din(w_dff_B_sVqsQlWz2_1),.dout(w_dff_B_2qC9ernC1_1),.clk(gclk));
	jdff dff_B_l4AxyD8e1_1(.din(w_dff_B_2qC9ernC1_1),.dout(w_dff_B_l4AxyD8e1_1),.clk(gclk));
	jdff dff_B_qqGPhaID0_1(.din(w_dff_B_l4AxyD8e1_1),.dout(w_dff_B_qqGPhaID0_1),.clk(gclk));
	jdff dff_B_hkBaqYUO0_1(.din(w_dff_B_qqGPhaID0_1),.dout(w_dff_B_hkBaqYUO0_1),.clk(gclk));
	jdff dff_A_oI3U0KAt2_0(.dout(w_n217_0[0]),.din(w_dff_A_oI3U0KAt2_0),.clk(gclk));
	jdff dff_A_CZbsdVEy4_0(.dout(w_n170_0[0]),.din(w_dff_A_CZbsdVEy4_0),.clk(gclk));
	jdff dff_A_l2rWvW2k6_0(.dout(w_dff_A_CZbsdVEy4_0),.din(w_dff_A_l2rWvW2k6_0),.clk(gclk));
	jdff dff_A_F5f6imAi0_0(.dout(w_dff_A_l2rWvW2k6_0),.din(w_dff_A_F5f6imAi0_0),.clk(gclk));
	jdff dff_A_s9IBI8gC0_0(.dout(w_dff_A_F5f6imAi0_0),.din(w_dff_A_s9IBI8gC0_0),.clk(gclk));
	jdff dff_A_L7VoPall2_0(.dout(w_dff_A_s9IBI8gC0_0),.din(w_dff_A_L7VoPall2_0),.clk(gclk));
	jdff dff_A_FZpxkJq41_0(.dout(w_dff_A_L7VoPall2_0),.din(w_dff_A_FZpxkJq41_0),.clk(gclk));
	jdff dff_A_nSH68aSX5_0(.dout(w_dff_A_FZpxkJq41_0),.din(w_dff_A_nSH68aSX5_0),.clk(gclk));
	jdff dff_A_LfmZrE2x6_0(.dout(w_dff_A_nSH68aSX5_0),.din(w_dff_A_LfmZrE2x6_0),.clk(gclk));
	jdff dff_A_J8sXJTQj3_0(.dout(w_dff_A_LfmZrE2x6_0),.din(w_dff_A_J8sXJTQj3_0),.clk(gclk));
	jdff dff_A_K2WTmrKj2_0(.dout(w_dff_A_J8sXJTQj3_0),.din(w_dff_A_K2WTmrKj2_0),.clk(gclk));
	jdff dff_A_nK8oxufB2_0(.dout(w_dff_A_K2WTmrKj2_0),.din(w_dff_A_nK8oxufB2_0),.clk(gclk));
	jdff dff_A_1YlUi9QA2_0(.dout(w_dff_A_nK8oxufB2_0),.din(w_dff_A_1YlUi9QA2_0),.clk(gclk));
	jdff dff_A_a0PbLUTj5_0(.dout(w_dff_A_1YlUi9QA2_0),.din(w_dff_A_a0PbLUTj5_0),.clk(gclk));
	jdff dff_B_0KXIUTjI6_1(.din(n177),.dout(w_dff_B_0KXIUTjI6_1),.clk(gclk));
	jdff dff_B_VjEdy8BS3_1(.din(w_dff_B_0KXIUTjI6_1),.dout(w_dff_B_VjEdy8BS3_1),.clk(gclk));
	jdff dff_B_1QgWNgf25_1(.din(w_dff_B_VjEdy8BS3_1),.dout(w_dff_B_1QgWNgf25_1),.clk(gclk));
	jdff dff_B_Lm04xTtY7_1(.din(w_dff_B_1QgWNgf25_1),.dout(w_dff_B_Lm04xTtY7_1),.clk(gclk));
	jdff dff_B_MjDQSxLh6_1(.din(w_dff_B_Lm04xTtY7_1),.dout(w_dff_B_MjDQSxLh6_1),.clk(gclk));
	jdff dff_B_xGYmIRLX6_1(.din(w_dff_B_MjDQSxLh6_1),.dout(w_dff_B_xGYmIRLX6_1),.clk(gclk));
	jdff dff_B_hWmYXbn75_1(.din(w_dff_B_xGYmIRLX6_1),.dout(w_dff_B_hWmYXbn75_1),.clk(gclk));
	jdff dff_B_U1JzXxtl2_1(.din(w_dff_B_hWmYXbn75_1),.dout(w_dff_B_U1JzXxtl2_1),.clk(gclk));
	jdff dff_B_yGIUHPSr3_1(.din(w_dff_B_U1JzXxtl2_1),.dout(w_dff_B_yGIUHPSr3_1),.clk(gclk));
	jdff dff_B_IV2jBIFP1_1(.din(w_dff_B_yGIUHPSr3_1),.dout(w_dff_B_IV2jBIFP1_1),.clk(gclk));
	jdff dff_A_urhleK3H5_0(.dout(w_n175_0[0]),.din(w_dff_A_urhleK3H5_0),.clk(gclk));
	jdff dff_A_copowyB36_0(.dout(w_n135_0[0]),.din(w_dff_A_copowyB36_0),.clk(gclk));
	jdff dff_A_u06mY1GP6_0(.dout(w_dff_A_copowyB36_0),.din(w_dff_A_u06mY1GP6_0),.clk(gclk));
	jdff dff_A_rzp7B8dk5_0(.dout(w_dff_A_u06mY1GP6_0),.din(w_dff_A_rzp7B8dk5_0),.clk(gclk));
	jdff dff_A_881PFUpB7_0(.dout(w_dff_A_rzp7B8dk5_0),.din(w_dff_A_881PFUpB7_0),.clk(gclk));
	jdff dff_A_hZgS5Bne6_0(.dout(w_dff_A_881PFUpB7_0),.din(w_dff_A_hZgS5Bne6_0),.clk(gclk));
	jdff dff_A_I2LyFV8Y8_0(.dout(w_dff_A_hZgS5Bne6_0),.din(w_dff_A_I2LyFV8Y8_0),.clk(gclk));
	jdff dff_A_ylvADaxH1_0(.dout(w_dff_A_I2LyFV8Y8_0),.din(w_dff_A_ylvADaxH1_0),.clk(gclk));
	jdff dff_A_eVvk4y9j7_0(.dout(w_dff_A_ylvADaxH1_0),.din(w_dff_A_eVvk4y9j7_0),.clk(gclk));
	jdff dff_A_IkWXygCx2_0(.dout(w_dff_A_eVvk4y9j7_0),.din(w_dff_A_IkWXygCx2_0),.clk(gclk));
	jdff dff_A_lVJYfrnY4_0(.dout(w_dff_A_IkWXygCx2_0),.din(w_dff_A_lVJYfrnY4_0),.clk(gclk));
	jdff dff_A_gUdkwqQc8_0(.dout(w_dff_A_lVJYfrnY4_0),.din(w_dff_A_gUdkwqQc8_0),.clk(gclk));
	jdff dff_B_dMneHK9C0_1(.din(n142),.dout(w_dff_B_dMneHK9C0_1),.clk(gclk));
	jdff dff_B_mzwvJ4S71_1(.din(w_dff_B_dMneHK9C0_1),.dout(w_dff_B_mzwvJ4S71_1),.clk(gclk));
	jdff dff_B_KAqqqU1e9_1(.din(w_dff_B_mzwvJ4S71_1),.dout(w_dff_B_KAqqqU1e9_1),.clk(gclk));
	jdff dff_B_di436h908_1(.din(w_dff_B_KAqqqU1e9_1),.dout(w_dff_B_di436h908_1),.clk(gclk));
	jdff dff_B_TGYqgnsR9_1(.din(w_dff_B_di436h908_1),.dout(w_dff_B_TGYqgnsR9_1),.clk(gclk));
	jdff dff_B_Z1Tp3tO33_1(.din(w_dff_B_TGYqgnsR9_1),.dout(w_dff_B_Z1Tp3tO33_1),.clk(gclk));
	jdff dff_B_RFWMJ7Pm1_1(.din(w_dff_B_Z1Tp3tO33_1),.dout(w_dff_B_RFWMJ7Pm1_1),.clk(gclk));
	jdff dff_B_fQZLEDiW3_1(.din(w_dff_B_RFWMJ7Pm1_1),.dout(w_dff_B_fQZLEDiW3_1),.clk(gclk));
	jdff dff_A_mwVSDR3y2_0(.dout(w_n140_0[0]),.din(w_dff_A_mwVSDR3y2_0),.clk(gclk));
	jdff dff_A_caceFrAU7_0(.dout(w_n106_0[0]),.din(w_dff_A_caceFrAU7_0),.clk(gclk));
	jdff dff_A_MLhWjLzD1_0(.dout(w_dff_A_caceFrAU7_0),.din(w_dff_A_MLhWjLzD1_0),.clk(gclk));
	jdff dff_A_RVlWy1fW8_0(.dout(w_dff_A_MLhWjLzD1_0),.din(w_dff_A_RVlWy1fW8_0),.clk(gclk));
	jdff dff_A_Q0Bag0Gl3_0(.dout(w_dff_A_RVlWy1fW8_0),.din(w_dff_A_Q0Bag0Gl3_0),.clk(gclk));
	jdff dff_A_sNTl6OET2_0(.dout(w_dff_A_Q0Bag0Gl3_0),.din(w_dff_A_sNTl6OET2_0),.clk(gclk));
	jdff dff_A_jRTJA5X13_0(.dout(w_dff_A_sNTl6OET2_0),.din(w_dff_A_jRTJA5X13_0),.clk(gclk));
	jdff dff_A_2TqyeKPW3_0(.dout(w_dff_A_jRTJA5X13_0),.din(w_dff_A_2TqyeKPW3_0),.clk(gclk));
	jdff dff_A_wcpvyPjQ9_0(.dout(w_dff_A_2TqyeKPW3_0),.din(w_dff_A_wcpvyPjQ9_0),.clk(gclk));
	jdff dff_A_AFqrBfsz6_0(.dout(w_dff_A_wcpvyPjQ9_0),.din(w_dff_A_AFqrBfsz6_0),.clk(gclk));
	jdff dff_B_oW5xUkWv9_1(.din(n113),.dout(w_dff_B_oW5xUkWv9_1),.clk(gclk));
	jdff dff_B_9WApEw879_1(.din(w_dff_B_oW5xUkWv9_1),.dout(w_dff_B_9WApEw879_1),.clk(gclk));
	jdff dff_B_IewJZG8Z2_1(.din(w_dff_B_9WApEw879_1),.dout(w_dff_B_IewJZG8Z2_1),.clk(gclk));
	jdff dff_B_AUVscL8l3_1(.din(w_dff_B_IewJZG8Z2_1),.dout(w_dff_B_AUVscL8l3_1),.clk(gclk));
	jdff dff_B_Fts5z9WF7_1(.din(w_dff_B_AUVscL8l3_1),.dout(w_dff_B_Fts5z9WF7_1),.clk(gclk));
	jdff dff_B_q9owYeI12_1(.din(w_dff_B_Fts5z9WF7_1),.dout(w_dff_B_q9owYeI12_1),.clk(gclk));
	jdff dff_A_xbYlxVGw3_0(.dout(w_n111_0[0]),.din(w_dff_A_xbYlxVGw3_0),.clk(gclk));
	jdff dff_B_BBdFlk5W7_2(.din(n111),.dout(w_dff_B_BBdFlk5W7_2),.clk(gclk));
	jdff dff_B_CIHAMHnt6_2(.din(w_dff_B_BBdFlk5W7_2),.dout(w_dff_B_CIHAMHnt6_2),.clk(gclk));
	jdff dff_B_z1dMPwYz1_1(.din(n109),.dout(w_dff_B_z1dMPwYz1_1),.clk(gclk));
	jdff dff_A_7w36pcmb3_0(.dout(w_n86_0[0]),.din(w_dff_A_7w36pcmb3_0),.clk(gclk));
	jdff dff_A_FYmzH7fy9_0(.dout(w_dff_A_7w36pcmb3_0),.din(w_dff_A_FYmzH7fy9_0),.clk(gclk));
	jdff dff_A_u5BQHdau1_0(.dout(w_dff_A_FYmzH7fy9_0),.din(w_dff_A_u5BQHdau1_0),.clk(gclk));
	jdff dff_A_OBTyKFJL9_0(.dout(w_dff_A_u5BQHdau1_0),.din(w_dff_A_OBTyKFJL9_0),.clk(gclk));
	jdff dff_A_Ck4bOiEB2_0(.dout(w_dff_A_OBTyKFJL9_0),.din(w_dff_A_Ck4bOiEB2_0),.clk(gclk));
	jdff dff_A_Bv8lsQaE1_1(.dout(w_n103_0[1]),.din(w_dff_A_Bv8lsQaE1_1),.clk(gclk));
	jdff dff_B_sc9KY8Fy9_1(.din(n92),.dout(w_dff_B_sc9KY8Fy9_1),.clk(gclk));
	jdff dff_B_E7g2rWZE1_1(.din(n88),.dout(w_dff_B_E7g2rWZE1_1),.clk(gclk));
	jdff dff_B_g0p1OFM37_1(.din(w_dff_B_E7g2rWZE1_1),.dout(w_dff_B_g0p1OFM37_1),.clk(gclk));
	jdff dff_A_BhjmWNl43_0(.dout(w_n75_0[0]),.din(w_dff_A_BhjmWNl43_0),.clk(gclk));
	jdff dff_A_VGcuZtuh7_0(.dout(w_dff_A_BhjmWNl43_0),.din(w_dff_A_VGcuZtuh7_0),.clk(gclk));
	jdff dff_A_D8ZagyVs8_0(.dout(w_dff_A_VGcuZtuh7_0),.din(w_dff_A_D8ZagyVs8_0),.clk(gclk));
	jdff dff_A_KsYCjYWA6_1(.dout(w_n83_0[1]),.din(w_dff_A_KsYCjYWA6_1),.clk(gclk));
	jdff dff_A_gqHF4DZl2_0(.dout(w_n1017_0[0]),.din(w_dff_A_gqHF4DZl2_0),.clk(gclk));
	jdff dff_A_mXBLWQWm6_1(.dout(w_n911_0[1]),.din(w_dff_A_mXBLWQWm6_1),.clk(gclk));
	jdff dff_B_pUEoHEdA2_2(.din(n911),.dout(w_dff_B_pUEoHEdA2_2),.clk(gclk));
	jdff dff_B_VjDpVPtW5_2(.din(w_dff_B_pUEoHEdA2_2),.dout(w_dff_B_VjDpVPtW5_2),.clk(gclk));
	jdff dff_B_CDiezGLX1_2(.din(w_dff_B_VjDpVPtW5_2),.dout(w_dff_B_CDiezGLX1_2),.clk(gclk));
	jdff dff_B_hrNtueNY6_2(.din(w_dff_B_CDiezGLX1_2),.dout(w_dff_B_hrNtueNY6_2),.clk(gclk));
	jdff dff_B_xzXMQ78K6_2(.din(w_dff_B_hrNtueNY6_2),.dout(w_dff_B_xzXMQ78K6_2),.clk(gclk));
	jdff dff_B_KnVJIlNm9_2(.din(w_dff_B_xzXMQ78K6_2),.dout(w_dff_B_KnVJIlNm9_2),.clk(gclk));
	jdff dff_B_GwgI0yLp5_2(.din(w_dff_B_KnVJIlNm9_2),.dout(w_dff_B_GwgI0yLp5_2),.clk(gclk));
	jdff dff_B_Sj5HycJh8_2(.din(w_dff_B_GwgI0yLp5_2),.dout(w_dff_B_Sj5HycJh8_2),.clk(gclk));
	jdff dff_B_uiEOOmkb8_2(.din(w_dff_B_Sj5HycJh8_2),.dout(w_dff_B_uiEOOmkb8_2),.clk(gclk));
	jdff dff_B_pw2WIRZJ3_2(.din(w_dff_B_uiEOOmkb8_2),.dout(w_dff_B_pw2WIRZJ3_2),.clk(gclk));
	jdff dff_B_Mrqkuyqf2_2(.din(w_dff_B_pw2WIRZJ3_2),.dout(w_dff_B_Mrqkuyqf2_2),.clk(gclk));
	jdff dff_B_Y9sEi3Sb2_2(.din(w_dff_B_Mrqkuyqf2_2),.dout(w_dff_B_Y9sEi3Sb2_2),.clk(gclk));
	jdff dff_B_ejez8uTU3_2(.din(w_dff_B_Y9sEi3Sb2_2),.dout(w_dff_B_ejez8uTU3_2),.clk(gclk));
	jdff dff_B_srZchfgQ1_2(.din(w_dff_B_ejez8uTU3_2),.dout(w_dff_B_srZchfgQ1_2),.clk(gclk));
	jdff dff_B_mmxntYNI2_2(.din(w_dff_B_srZchfgQ1_2),.dout(w_dff_B_mmxntYNI2_2),.clk(gclk));
	jdff dff_B_0xu7klg74_2(.din(w_dff_B_mmxntYNI2_2),.dout(w_dff_B_0xu7klg74_2),.clk(gclk));
	jdff dff_B_8n6gF85X6_2(.din(w_dff_B_0xu7klg74_2),.dout(w_dff_B_8n6gF85X6_2),.clk(gclk));
	jdff dff_B_M41J3GWs9_2(.din(w_dff_B_8n6gF85X6_2),.dout(w_dff_B_M41J3GWs9_2),.clk(gclk));
	jdff dff_B_1NQNQZI22_2(.din(w_dff_B_M41J3GWs9_2),.dout(w_dff_B_1NQNQZI22_2),.clk(gclk));
	jdff dff_B_UKevyvjR8_2(.din(w_dff_B_1NQNQZI22_2),.dout(w_dff_B_UKevyvjR8_2),.clk(gclk));
	jdff dff_B_hXTjTZ819_2(.din(w_dff_B_UKevyvjR8_2),.dout(w_dff_B_hXTjTZ819_2),.clk(gclk));
	jdff dff_B_ec8USU462_2(.din(w_dff_B_hXTjTZ819_2),.dout(w_dff_B_ec8USU462_2),.clk(gclk));
	jdff dff_B_XHM6P4fV4_2(.din(w_dff_B_ec8USU462_2),.dout(w_dff_B_XHM6P4fV4_2),.clk(gclk));
	jdff dff_B_nmxeaKC10_2(.din(w_dff_B_XHM6P4fV4_2),.dout(w_dff_B_nmxeaKC10_2),.clk(gclk));
	jdff dff_B_QUSUmLwB4_2(.din(w_dff_B_nmxeaKC10_2),.dout(w_dff_B_QUSUmLwB4_2),.clk(gclk));
	jdff dff_B_eIfUjQ2X7_2(.din(w_dff_B_QUSUmLwB4_2),.dout(w_dff_B_eIfUjQ2X7_2),.clk(gclk));
	jdff dff_B_c5kKzlAa5_2(.din(w_dff_B_eIfUjQ2X7_2),.dout(w_dff_B_c5kKzlAa5_2),.clk(gclk));
	jdff dff_B_dN2IENDA3_2(.din(w_dff_B_c5kKzlAa5_2),.dout(w_dff_B_dN2IENDA3_2),.clk(gclk));
	jdff dff_B_zWIz0fXl1_2(.din(w_dff_B_dN2IENDA3_2),.dout(w_dff_B_zWIz0fXl1_2),.clk(gclk));
	jdff dff_B_Dx5Vtea18_2(.din(w_dff_B_zWIz0fXl1_2),.dout(w_dff_B_Dx5Vtea18_2),.clk(gclk));
	jdff dff_B_Zu75j4Lr1_2(.din(w_dff_B_Dx5Vtea18_2),.dout(w_dff_B_Zu75j4Lr1_2),.clk(gclk));
	jdff dff_B_BCStcs3G3_2(.din(w_dff_B_Zu75j4Lr1_2),.dout(w_dff_B_BCStcs3G3_2),.clk(gclk));
	jdff dff_B_Hws5aiKZ5_2(.din(w_dff_B_BCStcs3G3_2),.dout(w_dff_B_Hws5aiKZ5_2),.clk(gclk));
	jdff dff_B_GLO8DITt9_2(.din(w_dff_B_Hws5aiKZ5_2),.dout(w_dff_B_GLO8DITt9_2),.clk(gclk));
	jdff dff_A_03eNmzSV3_1(.dout(w_n915_0[1]),.din(w_dff_A_03eNmzSV3_1),.clk(gclk));
	jdff dff_A_UvcgMejF3_2(.dout(w_n915_0[2]),.din(w_dff_A_UvcgMejF3_2),.clk(gclk));
	jdff dff_B_Pl34Mh8Q8_3(.din(n915),.dout(w_dff_B_Pl34Mh8Q8_3),.clk(gclk));
	jdff dff_B_Babty6GB4_2(.din(n811),.dout(w_dff_B_Babty6GB4_2),.clk(gclk));
	jdff dff_B_nYw7Cytt7_2(.din(w_dff_B_Babty6GB4_2),.dout(w_dff_B_nYw7Cytt7_2),.clk(gclk));
	jdff dff_B_lqMIemrn7_2(.din(w_dff_B_nYw7Cytt7_2),.dout(w_dff_B_lqMIemrn7_2),.clk(gclk));
	jdff dff_B_ZV3VsDIL2_2(.din(w_dff_B_lqMIemrn7_2),.dout(w_dff_B_ZV3VsDIL2_2),.clk(gclk));
	jdff dff_B_2MIdKlGR5_2(.din(w_dff_B_ZV3VsDIL2_2),.dout(w_dff_B_2MIdKlGR5_2),.clk(gclk));
	jdff dff_B_LgUTvbRa3_2(.din(w_dff_B_2MIdKlGR5_2),.dout(w_dff_B_LgUTvbRa3_2),.clk(gclk));
	jdff dff_B_pAzOzIkd7_2(.din(w_dff_B_LgUTvbRa3_2),.dout(w_dff_B_pAzOzIkd7_2),.clk(gclk));
	jdff dff_B_6MWRjY6G2_2(.din(w_dff_B_pAzOzIkd7_2),.dout(w_dff_B_6MWRjY6G2_2),.clk(gclk));
	jdff dff_B_O7kF07mM5_2(.din(w_dff_B_6MWRjY6G2_2),.dout(w_dff_B_O7kF07mM5_2),.clk(gclk));
	jdff dff_B_doLjYIdy4_2(.din(w_dff_B_O7kF07mM5_2),.dout(w_dff_B_doLjYIdy4_2),.clk(gclk));
	jdff dff_B_ErzC8j3T4_2(.din(w_dff_B_doLjYIdy4_2),.dout(w_dff_B_ErzC8j3T4_2),.clk(gclk));
	jdff dff_B_lrDU8tK61_2(.din(w_dff_B_ErzC8j3T4_2),.dout(w_dff_B_lrDU8tK61_2),.clk(gclk));
	jdff dff_B_XhXMM1HG7_2(.din(w_dff_B_lrDU8tK61_2),.dout(w_dff_B_XhXMM1HG7_2),.clk(gclk));
	jdff dff_B_fMDKbW5C9_2(.din(w_dff_B_XhXMM1HG7_2),.dout(w_dff_B_fMDKbW5C9_2),.clk(gclk));
	jdff dff_B_DX9eR9X29_2(.din(w_dff_B_fMDKbW5C9_2),.dout(w_dff_B_DX9eR9X29_2),.clk(gclk));
	jdff dff_B_cYuBZ7xA6_2(.din(w_dff_B_DX9eR9X29_2),.dout(w_dff_B_cYuBZ7xA6_2),.clk(gclk));
	jdff dff_B_9bpfnbwm4_2(.din(w_dff_B_cYuBZ7xA6_2),.dout(w_dff_B_9bpfnbwm4_2),.clk(gclk));
	jdff dff_B_TNWgqI0m0_2(.din(w_dff_B_9bpfnbwm4_2),.dout(w_dff_B_TNWgqI0m0_2),.clk(gclk));
	jdff dff_B_DcQtgnxc5_2(.din(w_dff_B_TNWgqI0m0_2),.dout(w_dff_B_DcQtgnxc5_2),.clk(gclk));
	jdff dff_B_HAjKsZxT4_2(.din(w_dff_B_DcQtgnxc5_2),.dout(w_dff_B_HAjKsZxT4_2),.clk(gclk));
	jdff dff_B_cPlr3C5O0_2(.din(w_dff_B_HAjKsZxT4_2),.dout(w_dff_B_cPlr3C5O0_2),.clk(gclk));
	jdff dff_B_bz5LR08S5_2(.din(w_dff_B_cPlr3C5O0_2),.dout(w_dff_B_bz5LR08S5_2),.clk(gclk));
	jdff dff_B_3LKMzIiD1_2(.din(w_dff_B_bz5LR08S5_2),.dout(w_dff_B_3LKMzIiD1_2),.clk(gclk));
	jdff dff_B_Ov38ClNX8_2(.din(w_dff_B_3LKMzIiD1_2),.dout(w_dff_B_Ov38ClNX8_2),.clk(gclk));
	jdff dff_B_yZeCImj18_2(.din(w_dff_B_Ov38ClNX8_2),.dout(w_dff_B_yZeCImj18_2),.clk(gclk));
	jdff dff_B_xHUV53na8_2(.din(w_dff_B_yZeCImj18_2),.dout(w_dff_B_xHUV53na8_2),.clk(gclk));
	jdff dff_B_nJwKoeBn6_2(.din(w_dff_B_xHUV53na8_2),.dout(w_dff_B_nJwKoeBn6_2),.clk(gclk));
	jdff dff_B_ddw9zLfN6_2(.din(w_dff_B_nJwKoeBn6_2),.dout(w_dff_B_ddw9zLfN6_2),.clk(gclk));
	jdff dff_B_lTD0oQA26_2(.din(w_dff_B_ddw9zLfN6_2),.dout(w_dff_B_lTD0oQA26_2),.clk(gclk));
	jdff dff_B_p388mCI49_2(.din(w_dff_B_lTD0oQA26_2),.dout(w_dff_B_p388mCI49_2),.clk(gclk));
	jdff dff_B_USy1Trii9_2(.din(w_dff_B_p388mCI49_2),.dout(w_dff_B_USy1Trii9_2),.clk(gclk));
	jdff dff_B_kqnKkiIb2_1(.din(n817),.dout(w_dff_B_kqnKkiIb2_1),.clk(gclk));
	jdff dff_B_Hu1BJ9Py4_1(.din(w_dff_B_kqnKkiIb2_1),.dout(w_dff_B_Hu1BJ9Py4_1),.clk(gclk));
	jdff dff_B_7x97j8du0_1(.din(w_dff_B_Hu1BJ9Py4_1),.dout(w_dff_B_7x97j8du0_1),.clk(gclk));
	jdff dff_B_sLCnAuXu5_1(.din(w_dff_B_7x97j8du0_1),.dout(w_dff_B_sLCnAuXu5_1),.clk(gclk));
	jdff dff_B_DDd5QNhG3_1(.din(w_dff_B_sLCnAuXu5_1),.dout(w_dff_B_DDd5QNhG3_1),.clk(gclk));
	jdff dff_B_25yuYMur2_1(.din(w_dff_B_DDd5QNhG3_1),.dout(w_dff_B_25yuYMur2_1),.clk(gclk));
	jdff dff_B_Aln5U4oX1_1(.din(w_dff_B_25yuYMur2_1),.dout(w_dff_B_Aln5U4oX1_1),.clk(gclk));
	jdff dff_B_uAnphWv57_1(.din(w_dff_B_Aln5U4oX1_1),.dout(w_dff_B_uAnphWv57_1),.clk(gclk));
	jdff dff_B_FzFs4l730_1(.din(w_dff_B_uAnphWv57_1),.dout(w_dff_B_FzFs4l730_1),.clk(gclk));
	jdff dff_B_36YYKauh5_1(.din(w_dff_B_FzFs4l730_1),.dout(w_dff_B_36YYKauh5_1),.clk(gclk));
	jdff dff_B_fu8sMLXT9_1(.din(w_dff_B_36YYKauh5_1),.dout(w_dff_B_fu8sMLXT9_1),.clk(gclk));
	jdff dff_B_1tIyPv249_1(.din(w_dff_B_fu8sMLXT9_1),.dout(w_dff_B_1tIyPv249_1),.clk(gclk));
	jdff dff_B_GZXxZIVQ1_1(.din(w_dff_B_1tIyPv249_1),.dout(w_dff_B_GZXxZIVQ1_1),.clk(gclk));
	jdff dff_B_aj8gI9Eh7_1(.din(w_dff_B_GZXxZIVQ1_1),.dout(w_dff_B_aj8gI9Eh7_1),.clk(gclk));
	jdff dff_B_aMcPJ7eC0_1(.din(w_dff_B_aj8gI9Eh7_1),.dout(w_dff_B_aMcPJ7eC0_1),.clk(gclk));
	jdff dff_B_XkpuDmtV4_1(.din(w_dff_B_aMcPJ7eC0_1),.dout(w_dff_B_XkpuDmtV4_1),.clk(gclk));
	jdff dff_B_H7x1NHHF5_1(.din(w_dff_B_XkpuDmtV4_1),.dout(w_dff_B_H7x1NHHF5_1),.clk(gclk));
	jdff dff_B_I7qfQnZh2_1(.din(w_dff_B_H7x1NHHF5_1),.dout(w_dff_B_I7qfQnZh2_1),.clk(gclk));
	jdff dff_B_HhvaNsXh1_1(.din(w_dff_B_I7qfQnZh2_1),.dout(w_dff_B_HhvaNsXh1_1),.clk(gclk));
	jdff dff_B_yUOZu5MH2_1(.din(w_dff_B_HhvaNsXh1_1),.dout(w_dff_B_yUOZu5MH2_1),.clk(gclk));
	jdff dff_B_BnPStVUf6_1(.din(w_dff_B_yUOZu5MH2_1),.dout(w_dff_B_BnPStVUf6_1),.clk(gclk));
	jdff dff_B_Fjf7Xnb44_1(.din(w_dff_B_BnPStVUf6_1),.dout(w_dff_B_Fjf7Xnb44_1),.clk(gclk));
	jdff dff_B_PYyFesMV4_1(.din(w_dff_B_Fjf7Xnb44_1),.dout(w_dff_B_PYyFesMV4_1),.clk(gclk));
	jdff dff_B_aTbs3Z4Y8_1(.din(w_dff_B_PYyFesMV4_1),.dout(w_dff_B_aTbs3Z4Y8_1),.clk(gclk));
	jdff dff_B_s9FXjr378_1(.din(w_dff_B_aTbs3Z4Y8_1),.dout(w_dff_B_s9FXjr378_1),.clk(gclk));
	jdff dff_B_GhgI8sMn9_1(.din(w_dff_B_s9FXjr378_1),.dout(w_dff_B_GhgI8sMn9_1),.clk(gclk));
	jdff dff_B_b3OvboPa2_1(.din(w_dff_B_GhgI8sMn9_1),.dout(w_dff_B_b3OvboPa2_1),.clk(gclk));
	jdff dff_B_tapHX3J87_1(.din(w_dff_B_b3OvboPa2_1),.dout(w_dff_B_tapHX3J87_1),.clk(gclk));
	jdff dff_A_DcHsrmTj0_0(.dout(w_n815_0[0]),.din(w_dff_A_DcHsrmTj0_0),.clk(gclk));
	jdff dff_A_X9EcOps89_0(.dout(w_n712_0[0]),.din(w_dff_A_X9EcOps89_0),.clk(gclk));
	jdff dff_A_tDpBYWhs0_0(.dout(w_dff_A_X9EcOps89_0),.din(w_dff_A_tDpBYWhs0_0),.clk(gclk));
	jdff dff_A_PIoYYLe65_0(.dout(w_dff_A_tDpBYWhs0_0),.din(w_dff_A_PIoYYLe65_0),.clk(gclk));
	jdff dff_A_TyrVEJwB5_0(.dout(w_dff_A_PIoYYLe65_0),.din(w_dff_A_TyrVEJwB5_0),.clk(gclk));
	jdff dff_A_tUmYli7r3_0(.dout(w_dff_A_TyrVEJwB5_0),.din(w_dff_A_tUmYli7r3_0),.clk(gclk));
	jdff dff_A_B5SWPUFX6_0(.dout(w_dff_A_tUmYli7r3_0),.din(w_dff_A_B5SWPUFX6_0),.clk(gclk));
	jdff dff_A_qUjQ0fw15_0(.dout(w_dff_A_B5SWPUFX6_0),.din(w_dff_A_qUjQ0fw15_0),.clk(gclk));
	jdff dff_A_byfQ5dol3_0(.dout(w_dff_A_qUjQ0fw15_0),.din(w_dff_A_byfQ5dol3_0),.clk(gclk));
	jdff dff_A_ADxtSsGn7_0(.dout(w_dff_A_byfQ5dol3_0),.din(w_dff_A_ADxtSsGn7_0),.clk(gclk));
	jdff dff_A_R9DfQBYp6_0(.dout(w_dff_A_ADxtSsGn7_0),.din(w_dff_A_R9DfQBYp6_0),.clk(gclk));
	jdff dff_A_F7KZfXTX4_0(.dout(w_dff_A_R9DfQBYp6_0),.din(w_dff_A_F7KZfXTX4_0),.clk(gclk));
	jdff dff_A_DctNQRuQ9_0(.dout(w_dff_A_F7KZfXTX4_0),.din(w_dff_A_DctNQRuQ9_0),.clk(gclk));
	jdff dff_A_XZzIT9oc9_0(.dout(w_dff_A_DctNQRuQ9_0),.din(w_dff_A_XZzIT9oc9_0),.clk(gclk));
	jdff dff_A_rGgClRSu2_0(.dout(w_dff_A_XZzIT9oc9_0),.din(w_dff_A_rGgClRSu2_0),.clk(gclk));
	jdff dff_A_1ArKhLZG5_0(.dout(w_dff_A_rGgClRSu2_0),.din(w_dff_A_1ArKhLZG5_0),.clk(gclk));
	jdff dff_A_nd0uN8eP6_0(.dout(w_dff_A_1ArKhLZG5_0),.din(w_dff_A_nd0uN8eP6_0),.clk(gclk));
	jdff dff_A_6JNmbeze2_0(.dout(w_dff_A_nd0uN8eP6_0),.din(w_dff_A_6JNmbeze2_0),.clk(gclk));
	jdff dff_A_861fChDR6_0(.dout(w_dff_A_6JNmbeze2_0),.din(w_dff_A_861fChDR6_0),.clk(gclk));
	jdff dff_A_R20mrMac7_0(.dout(w_dff_A_861fChDR6_0),.din(w_dff_A_R20mrMac7_0),.clk(gclk));
	jdff dff_A_A1IAdkBD1_0(.dout(w_dff_A_R20mrMac7_0),.din(w_dff_A_A1IAdkBD1_0),.clk(gclk));
	jdff dff_A_ir0Ooy688_0(.dout(w_dff_A_A1IAdkBD1_0),.din(w_dff_A_ir0Ooy688_0),.clk(gclk));
	jdff dff_A_bnnfhVE25_0(.dout(w_dff_A_ir0Ooy688_0),.din(w_dff_A_bnnfhVE25_0),.clk(gclk));
	jdff dff_A_SiTqRunJ6_0(.dout(w_dff_A_bnnfhVE25_0),.din(w_dff_A_SiTqRunJ6_0),.clk(gclk));
	jdff dff_A_nimgtCq04_0(.dout(w_dff_A_SiTqRunJ6_0),.din(w_dff_A_nimgtCq04_0),.clk(gclk));
	jdff dff_A_0Hzxoq856_0(.dout(w_dff_A_nimgtCq04_0),.din(w_dff_A_0Hzxoq856_0),.clk(gclk));
	jdff dff_A_tUjyESBT0_0(.dout(w_dff_A_0Hzxoq856_0),.din(w_dff_A_tUjyESBT0_0),.clk(gclk));
	jdff dff_A_08opqNZx2_0(.dout(w_dff_A_tUjyESBT0_0),.din(w_dff_A_08opqNZx2_0),.clk(gclk));
	jdff dff_A_KhOaql1O5_0(.dout(w_dff_A_08opqNZx2_0),.din(w_dff_A_KhOaql1O5_0),.clk(gclk));
	jdff dff_A_bENhUFb61_0(.dout(w_dff_A_KhOaql1O5_0),.din(w_dff_A_bENhUFb61_0),.clk(gclk));
	jdff dff_A_QQiW9jHY7_1(.dout(w_n717_0[1]),.din(w_dff_A_QQiW9jHY7_1),.clk(gclk));
	jdff dff_A_UZCyLOk90_2(.dout(w_n717_0[2]),.din(w_dff_A_UZCyLOk90_2),.clk(gclk));
	jdff dff_A_tT4vusQK8_0(.dout(w_n620_0[0]),.din(w_dff_A_tT4vusQK8_0),.clk(gclk));
	jdff dff_A_FJ0hg7Qw3_0(.dout(w_dff_A_tT4vusQK8_0),.din(w_dff_A_FJ0hg7Qw3_0),.clk(gclk));
	jdff dff_A_PObZri7O3_0(.dout(w_dff_A_FJ0hg7Qw3_0),.din(w_dff_A_PObZri7O3_0),.clk(gclk));
	jdff dff_A_8oqumgGL0_0(.dout(w_dff_A_PObZri7O3_0),.din(w_dff_A_8oqumgGL0_0),.clk(gclk));
	jdff dff_A_0qPY32M88_0(.dout(w_dff_A_8oqumgGL0_0),.din(w_dff_A_0qPY32M88_0),.clk(gclk));
	jdff dff_A_QW3D3Aaz4_0(.dout(w_dff_A_0qPY32M88_0),.din(w_dff_A_QW3D3Aaz4_0),.clk(gclk));
	jdff dff_A_wK2JlDMM7_0(.dout(w_dff_A_QW3D3Aaz4_0),.din(w_dff_A_wK2JlDMM7_0),.clk(gclk));
	jdff dff_A_e8FCEq2U7_0(.dout(w_dff_A_wK2JlDMM7_0),.din(w_dff_A_e8FCEq2U7_0),.clk(gclk));
	jdff dff_A_HrpWBUEL6_0(.dout(w_dff_A_e8FCEq2U7_0),.din(w_dff_A_HrpWBUEL6_0),.clk(gclk));
	jdff dff_A_PM6eaZ0h4_0(.dout(w_dff_A_HrpWBUEL6_0),.din(w_dff_A_PM6eaZ0h4_0),.clk(gclk));
	jdff dff_A_4Lmm1Ver6_0(.dout(w_dff_A_PM6eaZ0h4_0),.din(w_dff_A_4Lmm1Ver6_0),.clk(gclk));
	jdff dff_A_ZSzMyIF78_0(.dout(w_dff_A_4Lmm1Ver6_0),.din(w_dff_A_ZSzMyIF78_0),.clk(gclk));
	jdff dff_A_uxSz08EX3_0(.dout(w_dff_A_ZSzMyIF78_0),.din(w_dff_A_uxSz08EX3_0),.clk(gclk));
	jdff dff_A_l6Lu9EAc0_0(.dout(w_dff_A_uxSz08EX3_0),.din(w_dff_A_l6Lu9EAc0_0),.clk(gclk));
	jdff dff_A_fodFrSok9_0(.dout(w_dff_A_l6Lu9EAc0_0),.din(w_dff_A_fodFrSok9_0),.clk(gclk));
	jdff dff_A_d4BkEOxs1_0(.dout(w_dff_A_fodFrSok9_0),.din(w_dff_A_d4BkEOxs1_0),.clk(gclk));
	jdff dff_A_yzBKiAe29_0(.dout(w_dff_A_d4BkEOxs1_0),.din(w_dff_A_yzBKiAe29_0),.clk(gclk));
	jdff dff_A_D77r10yO3_0(.dout(w_dff_A_yzBKiAe29_0),.din(w_dff_A_D77r10yO3_0),.clk(gclk));
	jdff dff_A_Kwtkl8wZ9_0(.dout(w_dff_A_D77r10yO3_0),.din(w_dff_A_Kwtkl8wZ9_0),.clk(gclk));
	jdff dff_A_VuFm5zs82_0(.dout(w_dff_A_Kwtkl8wZ9_0),.din(w_dff_A_VuFm5zs82_0),.clk(gclk));
	jdff dff_A_z4S8U2114_0(.dout(w_dff_A_VuFm5zs82_0),.din(w_dff_A_z4S8U2114_0),.clk(gclk));
	jdff dff_A_E0zGS5465_0(.dout(w_dff_A_z4S8U2114_0),.din(w_dff_A_E0zGS5465_0),.clk(gclk));
	jdff dff_A_doKv2wNU0_0(.dout(w_dff_A_E0zGS5465_0),.din(w_dff_A_doKv2wNU0_0),.clk(gclk));
	jdff dff_A_p1w6RrO36_0(.dout(w_dff_A_doKv2wNU0_0),.din(w_dff_A_p1w6RrO36_0),.clk(gclk));
	jdff dff_A_TSP6erdd4_0(.dout(w_dff_A_p1w6RrO36_0),.din(w_dff_A_TSP6erdd4_0),.clk(gclk));
	jdff dff_A_wBTF6tG97_0(.dout(w_dff_A_TSP6erdd4_0),.din(w_dff_A_wBTF6tG97_0),.clk(gclk));
	jdff dff_A_lbCS54R79_0(.dout(w_dff_A_wBTF6tG97_0),.din(w_dff_A_lbCS54R79_0),.clk(gclk));
	jdff dff_A_cjuBMvDR1_1(.dout(w_n625_0[1]),.din(w_dff_A_cjuBMvDR1_1),.clk(gclk));
	jdff dff_A_1CFFVbwM8_2(.dout(w_n625_0[2]),.din(w_dff_A_1CFFVbwM8_2),.clk(gclk));
	jdff dff_A_Egp6zTmU2_0(.dout(w_n535_0[0]),.din(w_dff_A_Egp6zTmU2_0),.clk(gclk));
	jdff dff_A_xLqVU8W88_0(.dout(w_dff_A_Egp6zTmU2_0),.din(w_dff_A_xLqVU8W88_0),.clk(gclk));
	jdff dff_A_Gt6SSnBR8_0(.dout(w_dff_A_xLqVU8W88_0),.din(w_dff_A_Gt6SSnBR8_0),.clk(gclk));
	jdff dff_A_6VHD1qXu6_0(.dout(w_dff_A_Gt6SSnBR8_0),.din(w_dff_A_6VHD1qXu6_0),.clk(gclk));
	jdff dff_A_AiHNnsgj0_0(.dout(w_dff_A_6VHD1qXu6_0),.din(w_dff_A_AiHNnsgj0_0),.clk(gclk));
	jdff dff_A_iQ16p6fm1_0(.dout(w_dff_A_AiHNnsgj0_0),.din(w_dff_A_iQ16p6fm1_0),.clk(gclk));
	jdff dff_A_KJhlpZXr4_0(.dout(w_dff_A_iQ16p6fm1_0),.din(w_dff_A_KJhlpZXr4_0),.clk(gclk));
	jdff dff_A_OUM44gny1_0(.dout(w_dff_A_KJhlpZXr4_0),.din(w_dff_A_OUM44gny1_0),.clk(gclk));
	jdff dff_A_ivOB8jzk1_0(.dout(w_dff_A_OUM44gny1_0),.din(w_dff_A_ivOB8jzk1_0),.clk(gclk));
	jdff dff_A_15ZPBWxq5_0(.dout(w_dff_A_ivOB8jzk1_0),.din(w_dff_A_15ZPBWxq5_0),.clk(gclk));
	jdff dff_A_IeSFViUk8_0(.dout(w_dff_A_15ZPBWxq5_0),.din(w_dff_A_IeSFViUk8_0),.clk(gclk));
	jdff dff_A_W1jKxoDm3_0(.dout(w_dff_A_IeSFViUk8_0),.din(w_dff_A_W1jKxoDm3_0),.clk(gclk));
	jdff dff_A_UwHW28Du2_0(.dout(w_dff_A_W1jKxoDm3_0),.din(w_dff_A_UwHW28Du2_0),.clk(gclk));
	jdff dff_A_BlSkSZEg8_0(.dout(w_dff_A_UwHW28Du2_0),.din(w_dff_A_BlSkSZEg8_0),.clk(gclk));
	jdff dff_A_5b7OK6dR3_0(.dout(w_dff_A_BlSkSZEg8_0),.din(w_dff_A_5b7OK6dR3_0),.clk(gclk));
	jdff dff_A_XZ7qrrG87_0(.dout(w_dff_A_5b7OK6dR3_0),.din(w_dff_A_XZ7qrrG87_0),.clk(gclk));
	jdff dff_A_uCOA7kCG7_0(.dout(w_dff_A_XZ7qrrG87_0),.din(w_dff_A_uCOA7kCG7_0),.clk(gclk));
	jdff dff_A_M4IutWMU0_0(.dout(w_dff_A_uCOA7kCG7_0),.din(w_dff_A_M4IutWMU0_0),.clk(gclk));
	jdff dff_A_RadhUKnM2_0(.dout(w_dff_A_M4IutWMU0_0),.din(w_dff_A_RadhUKnM2_0),.clk(gclk));
	jdff dff_A_Fct10wJE9_0(.dout(w_dff_A_RadhUKnM2_0),.din(w_dff_A_Fct10wJE9_0),.clk(gclk));
	jdff dff_A_kpmSESC04_0(.dout(w_dff_A_Fct10wJE9_0),.din(w_dff_A_kpmSESC04_0),.clk(gclk));
	jdff dff_A_2yu0lIUe7_0(.dout(w_dff_A_kpmSESC04_0),.din(w_dff_A_2yu0lIUe7_0),.clk(gclk));
	jdff dff_A_dx5QL2HK5_0(.dout(w_dff_A_2yu0lIUe7_0),.din(w_dff_A_dx5QL2HK5_0),.clk(gclk));
	jdff dff_A_ngALKgO94_0(.dout(w_dff_A_dx5QL2HK5_0),.din(w_dff_A_ngALKgO94_0),.clk(gclk));
	jdff dff_A_A06Hb1ms3_0(.dout(w_dff_A_ngALKgO94_0),.din(w_dff_A_A06Hb1ms3_0),.clk(gclk));
	jdff dff_A_ZQVdk6Lq8_1(.dout(w_n540_0[1]),.din(w_dff_A_ZQVdk6Lq8_1),.clk(gclk));
	jdff dff_A_gfmfUuPd7_2(.dout(w_n540_0[2]),.din(w_dff_A_gfmfUuPd7_2),.clk(gclk));
	jdff dff_A_e0kImvxC3_0(.dout(w_n457_0[0]),.din(w_dff_A_e0kImvxC3_0),.clk(gclk));
	jdff dff_A_eD7Ix6Wj8_0(.dout(w_dff_A_e0kImvxC3_0),.din(w_dff_A_eD7Ix6Wj8_0),.clk(gclk));
	jdff dff_A_3uGzoZuT4_0(.dout(w_dff_A_eD7Ix6Wj8_0),.din(w_dff_A_3uGzoZuT4_0),.clk(gclk));
	jdff dff_A_4RP6p57e9_0(.dout(w_dff_A_3uGzoZuT4_0),.din(w_dff_A_4RP6p57e9_0),.clk(gclk));
	jdff dff_A_QW03tm6Y2_0(.dout(w_dff_A_4RP6p57e9_0),.din(w_dff_A_QW03tm6Y2_0),.clk(gclk));
	jdff dff_A_9j1eNQgB5_0(.dout(w_dff_A_QW03tm6Y2_0),.din(w_dff_A_9j1eNQgB5_0),.clk(gclk));
	jdff dff_A_UTmAqdE04_0(.dout(w_dff_A_9j1eNQgB5_0),.din(w_dff_A_UTmAqdE04_0),.clk(gclk));
	jdff dff_A_jZk2AhTA9_0(.dout(w_dff_A_UTmAqdE04_0),.din(w_dff_A_jZk2AhTA9_0),.clk(gclk));
	jdff dff_A_zVwnH6Ss4_0(.dout(w_dff_A_jZk2AhTA9_0),.din(w_dff_A_zVwnH6Ss4_0),.clk(gclk));
	jdff dff_A_VN2IVTXW2_0(.dout(w_dff_A_zVwnH6Ss4_0),.din(w_dff_A_VN2IVTXW2_0),.clk(gclk));
	jdff dff_A_49Yn0lRu4_0(.dout(w_dff_A_VN2IVTXW2_0),.din(w_dff_A_49Yn0lRu4_0),.clk(gclk));
	jdff dff_A_MFXnEAzf0_0(.dout(w_dff_A_49Yn0lRu4_0),.din(w_dff_A_MFXnEAzf0_0),.clk(gclk));
	jdff dff_A_Giydvbdx5_0(.dout(w_dff_A_MFXnEAzf0_0),.din(w_dff_A_Giydvbdx5_0),.clk(gclk));
	jdff dff_A_a5G4Tqy92_0(.dout(w_dff_A_Giydvbdx5_0),.din(w_dff_A_a5G4Tqy92_0),.clk(gclk));
	jdff dff_A_nwlR48mJ8_0(.dout(w_dff_A_a5G4Tqy92_0),.din(w_dff_A_nwlR48mJ8_0),.clk(gclk));
	jdff dff_A_uHe5KRiu0_0(.dout(w_dff_A_nwlR48mJ8_0),.din(w_dff_A_uHe5KRiu0_0),.clk(gclk));
	jdff dff_A_oYEBCFhb0_0(.dout(w_dff_A_uHe5KRiu0_0),.din(w_dff_A_oYEBCFhb0_0),.clk(gclk));
	jdff dff_A_dOlZllaD2_0(.dout(w_dff_A_oYEBCFhb0_0),.din(w_dff_A_dOlZllaD2_0),.clk(gclk));
	jdff dff_A_PLYszZBE0_0(.dout(w_dff_A_dOlZllaD2_0),.din(w_dff_A_PLYszZBE0_0),.clk(gclk));
	jdff dff_A_vtt2ordJ5_0(.dout(w_dff_A_PLYszZBE0_0),.din(w_dff_A_vtt2ordJ5_0),.clk(gclk));
	jdff dff_A_WaCa1zKv0_0(.dout(w_dff_A_vtt2ordJ5_0),.din(w_dff_A_WaCa1zKv0_0),.clk(gclk));
	jdff dff_A_Ub49KRTY6_0(.dout(w_dff_A_WaCa1zKv0_0),.din(w_dff_A_Ub49KRTY6_0),.clk(gclk));
	jdff dff_A_ILxVErOV7_0(.dout(w_dff_A_Ub49KRTY6_0),.din(w_dff_A_ILxVErOV7_0),.clk(gclk));
	jdff dff_A_I5tXqzfD0_1(.dout(w_n462_0[1]),.din(w_dff_A_I5tXqzfD0_1),.clk(gclk));
	jdff dff_A_QfR65i8R2_2(.dout(w_n462_0[2]),.din(w_dff_A_QfR65i8R2_2),.clk(gclk));
	jdff dff_A_OgKaEuyH0_0(.dout(w_n386_0[0]),.din(w_dff_A_OgKaEuyH0_0),.clk(gclk));
	jdff dff_A_JNRIqG7Q1_0(.dout(w_dff_A_OgKaEuyH0_0),.din(w_dff_A_JNRIqG7Q1_0),.clk(gclk));
	jdff dff_A_kGZrLCOB5_0(.dout(w_dff_A_JNRIqG7Q1_0),.din(w_dff_A_kGZrLCOB5_0),.clk(gclk));
	jdff dff_A_52cI6y6R4_0(.dout(w_dff_A_kGZrLCOB5_0),.din(w_dff_A_52cI6y6R4_0),.clk(gclk));
	jdff dff_A_b10JSLqZ0_0(.dout(w_dff_A_52cI6y6R4_0),.din(w_dff_A_b10JSLqZ0_0),.clk(gclk));
	jdff dff_A_Y2wZLREn3_0(.dout(w_dff_A_b10JSLqZ0_0),.din(w_dff_A_Y2wZLREn3_0),.clk(gclk));
	jdff dff_A_1JcpxVic2_0(.dout(w_dff_A_Y2wZLREn3_0),.din(w_dff_A_1JcpxVic2_0),.clk(gclk));
	jdff dff_A_9qq9DEtF6_0(.dout(w_dff_A_1JcpxVic2_0),.din(w_dff_A_9qq9DEtF6_0),.clk(gclk));
	jdff dff_A_WjyFuhvk7_0(.dout(w_dff_A_9qq9DEtF6_0),.din(w_dff_A_WjyFuhvk7_0),.clk(gclk));
	jdff dff_A_6eDZJBO78_0(.dout(w_dff_A_WjyFuhvk7_0),.din(w_dff_A_6eDZJBO78_0),.clk(gclk));
	jdff dff_A_G48Bm8im9_0(.dout(w_dff_A_6eDZJBO78_0),.din(w_dff_A_G48Bm8im9_0),.clk(gclk));
	jdff dff_A_BHNaKbSr7_0(.dout(w_dff_A_G48Bm8im9_0),.din(w_dff_A_BHNaKbSr7_0),.clk(gclk));
	jdff dff_A_S3fzd61M0_0(.dout(w_dff_A_BHNaKbSr7_0),.din(w_dff_A_S3fzd61M0_0),.clk(gclk));
	jdff dff_A_njWEN1843_0(.dout(w_dff_A_S3fzd61M0_0),.din(w_dff_A_njWEN1843_0),.clk(gclk));
	jdff dff_A_AqQn5PND0_0(.dout(w_dff_A_njWEN1843_0),.din(w_dff_A_AqQn5PND0_0),.clk(gclk));
	jdff dff_A_j67mQTt59_0(.dout(w_dff_A_AqQn5PND0_0),.din(w_dff_A_j67mQTt59_0),.clk(gclk));
	jdff dff_A_V714H1cc5_0(.dout(w_dff_A_j67mQTt59_0),.din(w_dff_A_V714H1cc5_0),.clk(gclk));
	jdff dff_A_ivOfx6Ti0_0(.dout(w_dff_A_V714H1cc5_0),.din(w_dff_A_ivOfx6Ti0_0),.clk(gclk));
	jdff dff_A_PIIyxv3e4_0(.dout(w_dff_A_ivOfx6Ti0_0),.din(w_dff_A_PIIyxv3e4_0),.clk(gclk));
	jdff dff_A_2o2IXzwD8_0(.dout(w_dff_A_PIIyxv3e4_0),.din(w_dff_A_2o2IXzwD8_0),.clk(gclk));
	jdff dff_A_91CmjfIu8_0(.dout(w_dff_A_2o2IXzwD8_0),.din(w_dff_A_91CmjfIu8_0),.clk(gclk));
	jdff dff_A_X4AjoJhn4_1(.dout(w_n391_0[1]),.din(w_dff_A_X4AjoJhn4_1),.clk(gclk));
	jdff dff_A_uXsEZDhL1_2(.dout(w_n391_0[2]),.din(w_dff_A_uXsEZDhL1_2),.clk(gclk));
	jdff dff_B_ZgcXkTFS6_3(.din(n391),.dout(w_dff_B_ZgcXkTFS6_3),.clk(gclk));
	jdff dff_B_tvsvbyGX0_3(.din(w_dff_B_ZgcXkTFS6_3),.dout(w_dff_B_tvsvbyGX0_3),.clk(gclk));
	jdff dff_B_c9r1jGgp4_3(.din(w_dff_B_tvsvbyGX0_3),.dout(w_dff_B_c9r1jGgp4_3),.clk(gclk));
	jdff dff_A_xvNLAp835_0(.dout(w_n323_0[0]),.din(w_dff_A_xvNLAp835_0),.clk(gclk));
	jdff dff_A_S9s49NdZ4_0(.dout(w_dff_A_xvNLAp835_0),.din(w_dff_A_S9s49NdZ4_0),.clk(gclk));
	jdff dff_A_eZYOnNfg9_0(.dout(w_dff_A_S9s49NdZ4_0),.din(w_dff_A_eZYOnNfg9_0),.clk(gclk));
	jdff dff_A_eiSqoekV6_0(.dout(w_dff_A_eZYOnNfg9_0),.din(w_dff_A_eiSqoekV6_0),.clk(gclk));
	jdff dff_A_B3r5OUTw8_0(.dout(w_dff_A_eiSqoekV6_0),.din(w_dff_A_B3r5OUTw8_0),.clk(gclk));
	jdff dff_A_WKlKpjuE4_0(.dout(w_dff_A_B3r5OUTw8_0),.din(w_dff_A_WKlKpjuE4_0),.clk(gclk));
	jdff dff_A_TFp0WR8M6_0(.dout(w_dff_A_WKlKpjuE4_0),.din(w_dff_A_TFp0WR8M6_0),.clk(gclk));
	jdff dff_A_u3MyCNRN6_0(.dout(w_dff_A_TFp0WR8M6_0),.din(w_dff_A_u3MyCNRN6_0),.clk(gclk));
	jdff dff_A_GSyojAc74_0(.dout(w_dff_A_u3MyCNRN6_0),.din(w_dff_A_GSyojAc74_0),.clk(gclk));
	jdff dff_A_AQoChlQw6_0(.dout(w_dff_A_GSyojAc74_0),.din(w_dff_A_AQoChlQw6_0),.clk(gclk));
	jdff dff_A_wVj7xcz45_0(.dout(w_dff_A_AQoChlQw6_0),.din(w_dff_A_wVj7xcz45_0),.clk(gclk));
	jdff dff_A_r6LCIgO77_0(.dout(w_dff_A_wVj7xcz45_0),.din(w_dff_A_r6LCIgO77_0),.clk(gclk));
	jdff dff_A_ygdhYGnG1_0(.dout(w_dff_A_r6LCIgO77_0),.din(w_dff_A_ygdhYGnG1_0),.clk(gclk));
	jdff dff_A_XiDKXq3e1_0(.dout(w_dff_A_ygdhYGnG1_0),.din(w_dff_A_XiDKXq3e1_0),.clk(gclk));
	jdff dff_A_52wPN3b80_0(.dout(w_dff_A_XiDKXq3e1_0),.din(w_dff_A_52wPN3b80_0),.clk(gclk));
	jdff dff_A_YabRlF152_0(.dout(w_dff_A_52wPN3b80_0),.din(w_dff_A_YabRlF152_0),.clk(gclk));
	jdff dff_A_0eoWrf1S3_1(.dout(w_n328_0[1]),.din(w_dff_A_0eoWrf1S3_1),.clk(gclk));
	jdff dff_A_iwaBUwCU1_2(.dout(w_n328_0[2]),.din(w_dff_A_iwaBUwCU1_2),.clk(gclk));
	jdff dff_A_FrOgE1JG7_0(.dout(w_n267_0[0]),.din(w_dff_A_FrOgE1JG7_0),.clk(gclk));
	jdff dff_A_PTUCHwB83_0(.dout(w_dff_A_FrOgE1JG7_0),.din(w_dff_A_PTUCHwB83_0),.clk(gclk));
	jdff dff_A_nx9yNsZn8_0(.dout(w_dff_A_PTUCHwB83_0),.din(w_dff_A_nx9yNsZn8_0),.clk(gclk));
	jdff dff_A_cTdyOx3I2_0(.dout(w_dff_A_nx9yNsZn8_0),.din(w_dff_A_cTdyOx3I2_0),.clk(gclk));
	jdff dff_A_FbsFObmB8_0(.dout(w_dff_A_cTdyOx3I2_0),.din(w_dff_A_FbsFObmB8_0),.clk(gclk));
	jdff dff_A_lkubc8Xa2_0(.dout(w_dff_A_FbsFObmB8_0),.din(w_dff_A_lkubc8Xa2_0),.clk(gclk));
	jdff dff_A_eeg1YH272_0(.dout(w_dff_A_lkubc8Xa2_0),.din(w_dff_A_eeg1YH272_0),.clk(gclk));
	jdff dff_A_zOYXO5LO6_0(.dout(w_dff_A_eeg1YH272_0),.din(w_dff_A_zOYXO5LO6_0),.clk(gclk));
	jdff dff_A_ufOV3YgE1_0(.dout(w_dff_A_zOYXO5LO6_0),.din(w_dff_A_ufOV3YgE1_0),.clk(gclk));
	jdff dff_A_ISQhXHx75_0(.dout(w_dff_A_ufOV3YgE1_0),.din(w_dff_A_ISQhXHx75_0),.clk(gclk));
	jdff dff_A_LN0XjWtg3_0(.dout(w_dff_A_ISQhXHx75_0),.din(w_dff_A_LN0XjWtg3_0),.clk(gclk));
	jdff dff_A_oFhOgkps0_0(.dout(w_dff_A_LN0XjWtg3_0),.din(w_dff_A_oFhOgkps0_0),.clk(gclk));
	jdff dff_A_9yLDPtv77_0(.dout(w_dff_A_oFhOgkps0_0),.din(w_dff_A_9yLDPtv77_0),.clk(gclk));
	jdff dff_A_LOYtCh2c3_0(.dout(w_dff_A_9yLDPtv77_0),.din(w_dff_A_LOYtCh2c3_0),.clk(gclk));
	jdff dff_A_0tGESKVt5_1(.dout(w_n272_0[1]),.din(w_dff_A_0tGESKVt5_1),.clk(gclk));
	jdff dff_A_naHyJ4d17_2(.dout(w_n272_0[2]),.din(w_dff_A_naHyJ4d17_2),.clk(gclk));
	jdff dff_A_5inedgFM2_0(.dout(w_n218_0[0]),.din(w_dff_A_5inedgFM2_0),.clk(gclk));
	jdff dff_A_veKJvRCX5_0(.dout(w_dff_A_5inedgFM2_0),.din(w_dff_A_veKJvRCX5_0),.clk(gclk));
	jdff dff_A_vauHgFrb2_0(.dout(w_dff_A_veKJvRCX5_0),.din(w_dff_A_vauHgFrb2_0),.clk(gclk));
	jdff dff_A_ET1t7Bcr2_0(.dout(w_dff_A_vauHgFrb2_0),.din(w_dff_A_ET1t7Bcr2_0),.clk(gclk));
	jdff dff_A_9KEQbPbd1_0(.dout(w_dff_A_ET1t7Bcr2_0),.din(w_dff_A_9KEQbPbd1_0),.clk(gclk));
	jdff dff_A_HE5ukqLq5_0(.dout(w_dff_A_9KEQbPbd1_0),.din(w_dff_A_HE5ukqLq5_0),.clk(gclk));
	jdff dff_A_VHbxBVlD0_0(.dout(w_dff_A_HE5ukqLq5_0),.din(w_dff_A_VHbxBVlD0_0),.clk(gclk));
	jdff dff_A_k7H8XMyl3_0(.dout(w_dff_A_VHbxBVlD0_0),.din(w_dff_A_k7H8XMyl3_0),.clk(gclk));
	jdff dff_A_NQr1QQHL0_0(.dout(w_dff_A_k7H8XMyl3_0),.din(w_dff_A_NQr1QQHL0_0),.clk(gclk));
	jdff dff_A_V9tykzU10_0(.dout(w_dff_A_NQr1QQHL0_0),.din(w_dff_A_V9tykzU10_0),.clk(gclk));
	jdff dff_A_MvUuq6fk7_0(.dout(w_dff_A_V9tykzU10_0),.din(w_dff_A_MvUuq6fk7_0),.clk(gclk));
	jdff dff_A_AMQHIN923_0(.dout(w_dff_A_MvUuq6fk7_0),.din(w_dff_A_AMQHIN923_0),.clk(gclk));
	jdff dff_A_0A3wwcWf1_1(.dout(w_n223_0[1]),.din(w_dff_A_0A3wwcWf1_1),.clk(gclk));
	jdff dff_A_c04hZHBx0_2(.dout(w_n223_0[2]),.din(w_dff_A_c04hZHBx0_2),.clk(gclk));
	jdff dff_A_dAiBishI8_0(.dout(w_n176_0[0]),.din(w_dff_A_dAiBishI8_0),.clk(gclk));
	jdff dff_A_Aor2FHKo2_0(.dout(w_dff_A_dAiBishI8_0),.din(w_dff_A_Aor2FHKo2_0),.clk(gclk));
	jdff dff_A_SWnGiDW03_0(.dout(w_dff_A_Aor2FHKo2_0),.din(w_dff_A_SWnGiDW03_0),.clk(gclk));
	jdff dff_A_yMoETBab4_0(.dout(w_dff_A_SWnGiDW03_0),.din(w_dff_A_yMoETBab4_0),.clk(gclk));
	jdff dff_A_8v3CManF2_0(.dout(w_dff_A_yMoETBab4_0),.din(w_dff_A_8v3CManF2_0),.clk(gclk));
	jdff dff_A_ZmnPzlZr2_0(.dout(w_dff_A_8v3CManF2_0),.din(w_dff_A_ZmnPzlZr2_0),.clk(gclk));
	jdff dff_A_PcH7twzX5_0(.dout(w_dff_A_ZmnPzlZr2_0),.din(w_dff_A_PcH7twzX5_0),.clk(gclk));
	jdff dff_A_Qu9OlvZc4_0(.dout(w_dff_A_PcH7twzX5_0),.din(w_dff_A_Qu9OlvZc4_0),.clk(gclk));
	jdff dff_A_Dcbj3qnk0_0(.dout(w_dff_A_Qu9OlvZc4_0),.din(w_dff_A_Dcbj3qnk0_0),.clk(gclk));
	jdff dff_A_BpAHiX1R2_0(.dout(w_dff_A_Dcbj3qnk0_0),.din(w_dff_A_BpAHiX1R2_0),.clk(gclk));
	jdff dff_A_oiF60WcB7_1(.dout(w_n181_0[1]),.din(w_dff_A_oiF60WcB7_1),.clk(gclk));
	jdff dff_A_Cvh7nZWc3_2(.dout(w_n181_0[2]),.din(w_dff_A_Cvh7nZWc3_2),.clk(gclk));
	jdff dff_A_oumENl7w4_0(.dout(w_n141_0[0]),.din(w_dff_A_oumENl7w4_0),.clk(gclk));
	jdff dff_A_PqWvTibw6_0(.dout(w_dff_A_oumENl7w4_0),.din(w_dff_A_PqWvTibw6_0),.clk(gclk));
	jdff dff_A_augNwgFE2_0(.dout(w_dff_A_PqWvTibw6_0),.din(w_dff_A_augNwgFE2_0),.clk(gclk));
	jdff dff_A_x4cVkPpp2_0(.dout(w_dff_A_augNwgFE2_0),.din(w_dff_A_x4cVkPpp2_0),.clk(gclk));
	jdff dff_A_3nmj66fQ7_0(.dout(w_dff_A_x4cVkPpp2_0),.din(w_dff_A_3nmj66fQ7_0),.clk(gclk));
	jdff dff_A_HOaGsRze1_0(.dout(w_dff_A_3nmj66fQ7_0),.din(w_dff_A_HOaGsRze1_0),.clk(gclk));
	jdff dff_A_Pr58Vjkp3_0(.dout(w_dff_A_HOaGsRze1_0),.din(w_dff_A_Pr58Vjkp3_0),.clk(gclk));
	jdff dff_A_EVTnbB3G6_0(.dout(w_dff_A_Pr58Vjkp3_0),.din(w_dff_A_EVTnbB3G6_0),.clk(gclk));
	jdff dff_A_t9jJ0Ax06_1(.dout(w_n146_0[1]),.din(w_dff_A_t9jJ0Ax06_1),.clk(gclk));
	jdff dff_A_ZnVzuhX42_2(.dout(w_n146_0[2]),.din(w_dff_A_ZnVzuhX42_2),.clk(gclk));
	jdff dff_A_vzDX4kE98_0(.dout(w_n112_0[0]),.din(w_dff_A_vzDX4kE98_0),.clk(gclk));
	jdff dff_A_DCn4SF351_0(.dout(w_dff_A_vzDX4kE98_0),.din(w_dff_A_DCn4SF351_0),.clk(gclk));
	jdff dff_A_MTsb8jqH3_0(.dout(w_dff_A_DCn4SF351_0),.din(w_dff_A_MTsb8jqH3_0),.clk(gclk));
	jdff dff_A_VBtoZvs29_0(.dout(w_dff_A_MTsb8jqH3_0),.din(w_dff_A_VBtoZvs29_0),.clk(gclk));
	jdff dff_A_FwDOSz354_0(.dout(w_dff_A_VBtoZvs29_0),.din(w_dff_A_FwDOSz354_0),.clk(gclk));
	jdff dff_A_YElQJLx72_0(.dout(w_dff_A_FwDOSz354_0),.din(w_dff_A_YElQJLx72_0),.clk(gclk));
	jdff dff_A_rLbe5iWw9_1(.dout(w_n117_0[1]),.din(w_dff_A_rLbe5iWw9_1),.clk(gclk));
	jdff dff_A_WU05vbqJ5_2(.dout(w_n117_0[2]),.din(w_dff_A_WU05vbqJ5_2),.clk(gclk));
	jdff dff_B_SdvaenAL9_3(.din(n117),.dout(w_dff_B_SdvaenAL9_3),.clk(gclk));
	jdff dff_B_qOlwIYSL5_3(.din(w_dff_B_SdvaenAL9_3),.dout(w_dff_B_qOlwIYSL5_3),.clk(gclk));
	jdff dff_B_7XBAQlWe7_1(.din(n114),.dout(w_dff_B_7XBAQlWe7_1),.clk(gclk));
	jdff dff_A_uVcTUwdv7_0(.dout(w_n91_0[0]),.din(w_dff_A_uVcTUwdv7_0),.clk(gclk));
	jdff dff_A_ScPbN5a19_0(.dout(w_dff_A_uVcTUwdv7_0),.din(w_dff_A_ScPbN5a19_0),.clk(gclk));
	jdff dff_A_4He3wXXc8_0(.dout(w_n80_0[0]),.din(w_dff_A_4He3wXXc8_0),.clk(gclk));
	jdff dff_A_V7rxrfus7_0(.dout(w_n1119_0[0]),.din(w_dff_A_V7rxrfus7_0),.clk(gclk));
	jdff dff_B_5qk6RfLR5_2(.din(n1119),.dout(w_dff_B_5qk6RfLR5_2),.clk(gclk));
	jdff dff_B_AwpYgIu32_2(.din(n1018),.dout(w_dff_B_AwpYgIu32_2),.clk(gclk));
	jdff dff_B_rxyDG2M89_2(.din(w_dff_B_AwpYgIu32_2),.dout(w_dff_B_rxyDG2M89_2),.clk(gclk));
	jdff dff_B_7wknFk848_2(.din(w_dff_B_rxyDG2M89_2),.dout(w_dff_B_7wknFk848_2),.clk(gclk));
	jdff dff_B_9DYGw7Dh6_2(.din(w_dff_B_7wknFk848_2),.dout(w_dff_B_9DYGw7Dh6_2),.clk(gclk));
	jdff dff_B_e8hpzakL7_2(.din(w_dff_B_9DYGw7Dh6_2),.dout(w_dff_B_e8hpzakL7_2),.clk(gclk));
	jdff dff_B_amro8CZb0_2(.din(w_dff_B_e8hpzakL7_2),.dout(w_dff_B_amro8CZb0_2),.clk(gclk));
	jdff dff_B_YyeAAAiz1_2(.din(w_dff_B_amro8CZb0_2),.dout(w_dff_B_YyeAAAiz1_2),.clk(gclk));
	jdff dff_B_W0peWllr3_2(.din(w_dff_B_YyeAAAiz1_2),.dout(w_dff_B_W0peWllr3_2),.clk(gclk));
	jdff dff_B_hqaT3nBH6_2(.din(w_dff_B_W0peWllr3_2),.dout(w_dff_B_hqaT3nBH6_2),.clk(gclk));
	jdff dff_B_m9SCfVrB9_2(.din(w_dff_B_hqaT3nBH6_2),.dout(w_dff_B_m9SCfVrB9_2),.clk(gclk));
	jdff dff_B_GeMbTlVP7_2(.din(w_dff_B_m9SCfVrB9_2),.dout(w_dff_B_GeMbTlVP7_2),.clk(gclk));
	jdff dff_B_KzQo3o3R9_2(.din(w_dff_B_GeMbTlVP7_2),.dout(w_dff_B_KzQo3o3R9_2),.clk(gclk));
	jdff dff_B_0cdUS7TV9_2(.din(w_dff_B_KzQo3o3R9_2),.dout(w_dff_B_0cdUS7TV9_2),.clk(gclk));
	jdff dff_B_5rywKQS15_2(.din(w_dff_B_0cdUS7TV9_2),.dout(w_dff_B_5rywKQS15_2),.clk(gclk));
	jdff dff_B_kylEJjic3_2(.din(w_dff_B_5rywKQS15_2),.dout(w_dff_B_kylEJjic3_2),.clk(gclk));
	jdff dff_B_TptfY84m1_2(.din(w_dff_B_kylEJjic3_2),.dout(w_dff_B_TptfY84m1_2),.clk(gclk));
	jdff dff_B_brYRrtJW9_2(.din(w_dff_B_TptfY84m1_2),.dout(w_dff_B_brYRrtJW9_2),.clk(gclk));
	jdff dff_B_Pt76kV2A9_2(.din(w_dff_B_brYRrtJW9_2),.dout(w_dff_B_Pt76kV2A9_2),.clk(gclk));
	jdff dff_B_Wi3KLufh9_2(.din(w_dff_B_Pt76kV2A9_2),.dout(w_dff_B_Wi3KLufh9_2),.clk(gclk));
	jdff dff_B_QTdE5kJz2_2(.din(w_dff_B_Wi3KLufh9_2),.dout(w_dff_B_QTdE5kJz2_2),.clk(gclk));
	jdff dff_B_AQg3C7z21_2(.din(w_dff_B_QTdE5kJz2_2),.dout(w_dff_B_AQg3C7z21_2),.clk(gclk));
	jdff dff_B_3w4zosuD7_2(.din(w_dff_B_AQg3C7z21_2),.dout(w_dff_B_3w4zosuD7_2),.clk(gclk));
	jdff dff_B_kiWf3GJU6_2(.din(w_dff_B_3w4zosuD7_2),.dout(w_dff_B_kiWf3GJU6_2),.clk(gclk));
	jdff dff_B_FuVVGGMD1_2(.din(w_dff_B_kiWf3GJU6_2),.dout(w_dff_B_FuVVGGMD1_2),.clk(gclk));
	jdff dff_B_IGRs6V3n6_2(.din(w_dff_B_FuVVGGMD1_2),.dout(w_dff_B_IGRs6V3n6_2),.clk(gclk));
	jdff dff_B_Dyi1YIAH2_2(.din(w_dff_B_IGRs6V3n6_2),.dout(w_dff_B_Dyi1YIAH2_2),.clk(gclk));
	jdff dff_B_90dv32rF7_2(.din(w_dff_B_Dyi1YIAH2_2),.dout(w_dff_B_90dv32rF7_2),.clk(gclk));
	jdff dff_B_utK3GTcc2_2(.din(w_dff_B_90dv32rF7_2),.dout(w_dff_B_utK3GTcc2_2),.clk(gclk));
	jdff dff_B_w8W9LDhj2_2(.din(w_dff_B_utK3GTcc2_2),.dout(w_dff_B_w8W9LDhj2_2),.clk(gclk));
	jdff dff_B_4wMmvEWk7_2(.din(w_dff_B_w8W9LDhj2_2),.dout(w_dff_B_4wMmvEWk7_2),.clk(gclk));
	jdff dff_B_83MZuWrc5_2(.din(w_dff_B_4wMmvEWk7_2),.dout(w_dff_B_83MZuWrc5_2),.clk(gclk));
	jdff dff_B_cLBThaVd3_2(.din(w_dff_B_83MZuWrc5_2),.dout(w_dff_B_cLBThaVd3_2),.clk(gclk));
	jdff dff_B_L1jNxXFS8_2(.din(w_dff_B_cLBThaVd3_2),.dout(w_dff_B_L1jNxXFS8_2),.clk(gclk));
	jdff dff_B_ZG439JIz6_2(.din(w_dff_B_L1jNxXFS8_2),.dout(w_dff_B_ZG439JIz6_2),.clk(gclk));
	jdff dff_A_dJHV3D2E4_0(.dout(w_n1022_0[0]),.din(w_dff_A_dJHV3D2E4_0),.clk(gclk));
	jdff dff_B_fLWRSZbu3_1(.din(n1020),.dout(w_dff_B_fLWRSZbu3_1),.clk(gclk));
	jdff dff_B_5Gg4QPp35_2(.din(n916),.dout(w_dff_B_5Gg4QPp35_2),.clk(gclk));
	jdff dff_B_yqiSydbO6_2(.din(w_dff_B_5Gg4QPp35_2),.dout(w_dff_B_yqiSydbO6_2),.clk(gclk));
	jdff dff_B_uJP7Zt6o2_2(.din(w_dff_B_yqiSydbO6_2),.dout(w_dff_B_uJP7Zt6o2_2),.clk(gclk));
	jdff dff_B_JHMxpmCT3_2(.din(w_dff_B_uJP7Zt6o2_2),.dout(w_dff_B_JHMxpmCT3_2),.clk(gclk));
	jdff dff_B_wBob4Vtm3_2(.din(w_dff_B_JHMxpmCT3_2),.dout(w_dff_B_wBob4Vtm3_2),.clk(gclk));
	jdff dff_B_aJymxLPy8_2(.din(w_dff_B_wBob4Vtm3_2),.dout(w_dff_B_aJymxLPy8_2),.clk(gclk));
	jdff dff_B_m3FvqUI57_2(.din(w_dff_B_aJymxLPy8_2),.dout(w_dff_B_m3FvqUI57_2),.clk(gclk));
	jdff dff_B_JhXFxKV94_2(.din(w_dff_B_m3FvqUI57_2),.dout(w_dff_B_JhXFxKV94_2),.clk(gclk));
	jdff dff_B_l6Jk3JnJ3_2(.din(w_dff_B_JhXFxKV94_2),.dout(w_dff_B_l6Jk3JnJ3_2),.clk(gclk));
	jdff dff_B_63EujrUG6_2(.din(w_dff_B_l6Jk3JnJ3_2),.dout(w_dff_B_63EujrUG6_2),.clk(gclk));
	jdff dff_B_AxiXIGmo8_2(.din(w_dff_B_63EujrUG6_2),.dout(w_dff_B_AxiXIGmo8_2),.clk(gclk));
	jdff dff_B_YK2EEB5H0_2(.din(w_dff_B_AxiXIGmo8_2),.dout(w_dff_B_YK2EEB5H0_2),.clk(gclk));
	jdff dff_B_58771CmY8_2(.din(w_dff_B_YK2EEB5H0_2),.dout(w_dff_B_58771CmY8_2),.clk(gclk));
	jdff dff_B_8Piz0tfp2_2(.din(w_dff_B_58771CmY8_2),.dout(w_dff_B_8Piz0tfp2_2),.clk(gclk));
	jdff dff_B_mceGSAbA7_2(.din(w_dff_B_8Piz0tfp2_2),.dout(w_dff_B_mceGSAbA7_2),.clk(gclk));
	jdff dff_B_4oEiDqDh3_2(.din(w_dff_B_mceGSAbA7_2),.dout(w_dff_B_4oEiDqDh3_2),.clk(gclk));
	jdff dff_B_K1sfVUCj5_2(.din(w_dff_B_4oEiDqDh3_2),.dout(w_dff_B_K1sfVUCj5_2),.clk(gclk));
	jdff dff_B_yvGS4cgp2_2(.din(w_dff_B_K1sfVUCj5_2),.dout(w_dff_B_yvGS4cgp2_2),.clk(gclk));
	jdff dff_B_jQjRYNtY3_2(.din(w_dff_B_yvGS4cgp2_2),.dout(w_dff_B_jQjRYNtY3_2),.clk(gclk));
	jdff dff_B_jZRzcMb97_2(.din(w_dff_B_jQjRYNtY3_2),.dout(w_dff_B_jZRzcMb97_2),.clk(gclk));
	jdff dff_B_4QPYsdQu2_2(.din(w_dff_B_jZRzcMb97_2),.dout(w_dff_B_4QPYsdQu2_2),.clk(gclk));
	jdff dff_B_1REA3eFh0_2(.din(w_dff_B_4QPYsdQu2_2),.dout(w_dff_B_1REA3eFh0_2),.clk(gclk));
	jdff dff_B_igXWHAIW3_2(.din(w_dff_B_1REA3eFh0_2),.dout(w_dff_B_igXWHAIW3_2),.clk(gclk));
	jdff dff_B_VjwhGhiQ1_2(.din(w_dff_B_igXWHAIW3_2),.dout(w_dff_B_VjwhGhiQ1_2),.clk(gclk));
	jdff dff_B_ZfPwlrQh7_2(.din(w_dff_B_VjwhGhiQ1_2),.dout(w_dff_B_ZfPwlrQh7_2),.clk(gclk));
	jdff dff_B_baM5UuUj9_2(.din(w_dff_B_ZfPwlrQh7_2),.dout(w_dff_B_baM5UuUj9_2),.clk(gclk));
	jdff dff_B_C97EUB5o5_2(.din(w_dff_B_baM5UuUj9_2),.dout(w_dff_B_C97EUB5o5_2),.clk(gclk));
	jdff dff_B_ay4RHgkB9_2(.din(w_dff_B_C97EUB5o5_2),.dout(w_dff_B_ay4RHgkB9_2),.clk(gclk));
	jdff dff_B_PrqImqy58_2(.din(w_dff_B_ay4RHgkB9_2),.dout(w_dff_B_PrqImqy58_2),.clk(gclk));
	jdff dff_B_NFctmz8z3_2(.din(w_dff_B_PrqImqy58_2),.dout(w_dff_B_NFctmz8z3_2),.clk(gclk));
	jdff dff_B_UGGY7aL27_2(.din(w_dff_B_NFctmz8z3_2),.dout(w_dff_B_UGGY7aL27_2),.clk(gclk));
	jdff dff_B_aGAepYLi9_2(.din(w_dff_B_UGGY7aL27_2),.dout(w_dff_B_aGAepYLi9_2),.clk(gclk));
	jdff dff_A_ifldbHus3_1(.dout(w_n1006_0[1]),.din(w_dff_A_ifldbHus3_1),.clk(gclk));
	jdff dff_A_Lk7C61MK4_0(.dout(w_n816_0[0]),.din(w_dff_A_Lk7C61MK4_0),.clk(gclk));
	jdff dff_A_XTeS7fHm4_0(.dout(w_dff_A_Lk7C61MK4_0),.din(w_dff_A_XTeS7fHm4_0),.clk(gclk));
	jdff dff_A_CG1Whsdx0_0(.dout(w_dff_A_XTeS7fHm4_0),.din(w_dff_A_CG1Whsdx0_0),.clk(gclk));
	jdff dff_A_cgePzAdx2_0(.dout(w_dff_A_CG1Whsdx0_0),.din(w_dff_A_cgePzAdx2_0),.clk(gclk));
	jdff dff_A_rPrYnz3m8_0(.dout(w_dff_A_cgePzAdx2_0),.din(w_dff_A_rPrYnz3m8_0),.clk(gclk));
	jdff dff_A_snzH7SAi8_0(.dout(w_dff_A_rPrYnz3m8_0),.din(w_dff_A_snzH7SAi8_0),.clk(gclk));
	jdff dff_A_ueBQLTmq2_0(.dout(w_dff_A_snzH7SAi8_0),.din(w_dff_A_ueBQLTmq2_0),.clk(gclk));
	jdff dff_A_6BaDtHaP1_0(.dout(w_dff_A_ueBQLTmq2_0),.din(w_dff_A_6BaDtHaP1_0),.clk(gclk));
	jdff dff_A_lkVvhpXu5_0(.dout(w_dff_A_6BaDtHaP1_0),.din(w_dff_A_lkVvhpXu5_0),.clk(gclk));
	jdff dff_A_YaOjGzi51_0(.dout(w_dff_A_lkVvhpXu5_0),.din(w_dff_A_YaOjGzi51_0),.clk(gclk));
	jdff dff_A_mqFlHYbJ9_0(.dout(w_dff_A_YaOjGzi51_0),.din(w_dff_A_mqFlHYbJ9_0),.clk(gclk));
	jdff dff_A_EXlWsVTM2_0(.dout(w_dff_A_mqFlHYbJ9_0),.din(w_dff_A_EXlWsVTM2_0),.clk(gclk));
	jdff dff_A_fIUAoLko8_0(.dout(w_dff_A_EXlWsVTM2_0),.din(w_dff_A_fIUAoLko8_0),.clk(gclk));
	jdff dff_A_XaNoVa8a3_0(.dout(w_dff_A_fIUAoLko8_0),.din(w_dff_A_XaNoVa8a3_0),.clk(gclk));
	jdff dff_A_P0gIU8ib9_0(.dout(w_dff_A_XaNoVa8a3_0),.din(w_dff_A_P0gIU8ib9_0),.clk(gclk));
	jdff dff_A_rVVKLcIm2_0(.dout(w_dff_A_P0gIU8ib9_0),.din(w_dff_A_rVVKLcIm2_0),.clk(gclk));
	jdff dff_A_o261iGzt7_0(.dout(w_dff_A_rVVKLcIm2_0),.din(w_dff_A_o261iGzt7_0),.clk(gclk));
	jdff dff_A_tjK8g2Eb0_0(.dout(w_dff_A_o261iGzt7_0),.din(w_dff_A_tjK8g2Eb0_0),.clk(gclk));
	jdff dff_A_kEephMl80_0(.dout(w_dff_A_tjK8g2Eb0_0),.din(w_dff_A_kEephMl80_0),.clk(gclk));
	jdff dff_A_KysHcyIl8_0(.dout(w_dff_A_kEephMl80_0),.din(w_dff_A_KysHcyIl8_0),.clk(gclk));
	jdff dff_A_ywZU3uOo5_0(.dout(w_dff_A_KysHcyIl8_0),.din(w_dff_A_ywZU3uOo5_0),.clk(gclk));
	jdff dff_A_sbbrMCKZ9_0(.dout(w_dff_A_ywZU3uOo5_0),.din(w_dff_A_sbbrMCKZ9_0),.clk(gclk));
	jdff dff_A_R3bd3qsZ2_0(.dout(w_dff_A_sbbrMCKZ9_0),.din(w_dff_A_R3bd3qsZ2_0),.clk(gclk));
	jdff dff_A_8yZubp9V5_0(.dout(w_dff_A_R3bd3qsZ2_0),.din(w_dff_A_8yZubp9V5_0),.clk(gclk));
	jdff dff_A_PygO025X9_0(.dout(w_dff_A_8yZubp9V5_0),.din(w_dff_A_PygO025X9_0),.clk(gclk));
	jdff dff_A_ElAq0Bqn2_0(.dout(w_dff_A_PygO025X9_0),.din(w_dff_A_ElAq0Bqn2_0),.clk(gclk));
	jdff dff_A_nJEAJzXB1_0(.dout(w_dff_A_ElAq0Bqn2_0),.din(w_dff_A_nJEAJzXB1_0),.clk(gclk));
	jdff dff_A_b45eTMbn1_0(.dout(w_dff_A_nJEAJzXB1_0),.din(w_dff_A_b45eTMbn1_0),.clk(gclk));
	jdff dff_A_dbuy7M5F6_0(.dout(w_dff_A_b45eTMbn1_0),.din(w_dff_A_dbuy7M5F6_0),.clk(gclk));
	jdff dff_A_XGAWw9VZ5_0(.dout(w_dff_A_dbuy7M5F6_0),.din(w_dff_A_XGAWw9VZ5_0),.clk(gclk));
	jdff dff_A_x6b9m6GW6_0(.dout(w_n820_0[0]),.din(w_dff_A_x6b9m6GW6_0),.clk(gclk));
	jdff dff_B_cMTiWGax5_1(.din(n818),.dout(w_dff_B_cMTiWGax5_1),.clk(gclk));
	jdff dff_B_uF6v6l9F4_2(.din(n719),.dout(w_dff_B_uF6v6l9F4_2),.clk(gclk));
	jdff dff_B_UJbDZzLl8_2(.din(w_dff_B_uF6v6l9F4_2),.dout(w_dff_B_UJbDZzLl8_2),.clk(gclk));
	jdff dff_B_33pWAx9J0_2(.din(w_dff_B_UJbDZzLl8_2),.dout(w_dff_B_33pWAx9J0_2),.clk(gclk));
	jdff dff_B_5fZfaQUm0_2(.din(w_dff_B_33pWAx9J0_2),.dout(w_dff_B_5fZfaQUm0_2),.clk(gclk));
	jdff dff_B_q4jJURHC3_2(.din(w_dff_B_5fZfaQUm0_2),.dout(w_dff_B_q4jJURHC3_2),.clk(gclk));
	jdff dff_B_FNQhTGUT2_2(.din(w_dff_B_q4jJURHC3_2),.dout(w_dff_B_FNQhTGUT2_2),.clk(gclk));
	jdff dff_B_OzDQ8Unp0_2(.din(w_dff_B_FNQhTGUT2_2),.dout(w_dff_B_OzDQ8Unp0_2),.clk(gclk));
	jdff dff_B_52RZW9OQ6_2(.din(w_dff_B_OzDQ8Unp0_2),.dout(w_dff_B_52RZW9OQ6_2),.clk(gclk));
	jdff dff_B_PsxwXRH22_2(.din(w_dff_B_52RZW9OQ6_2),.dout(w_dff_B_PsxwXRH22_2),.clk(gclk));
	jdff dff_B_xxGuBGhD5_2(.din(w_dff_B_PsxwXRH22_2),.dout(w_dff_B_xxGuBGhD5_2),.clk(gclk));
	jdff dff_B_SZaXjwHU5_2(.din(w_dff_B_xxGuBGhD5_2),.dout(w_dff_B_SZaXjwHU5_2),.clk(gclk));
	jdff dff_B_KAEC14Dg6_2(.din(w_dff_B_SZaXjwHU5_2),.dout(w_dff_B_KAEC14Dg6_2),.clk(gclk));
	jdff dff_B_QU9MbDhP0_2(.din(w_dff_B_KAEC14Dg6_2),.dout(w_dff_B_QU9MbDhP0_2),.clk(gclk));
	jdff dff_B_ySKUMeI93_2(.din(w_dff_B_QU9MbDhP0_2),.dout(w_dff_B_ySKUMeI93_2),.clk(gclk));
	jdff dff_B_9h6NlaLw6_2(.din(w_dff_B_ySKUMeI93_2),.dout(w_dff_B_9h6NlaLw6_2),.clk(gclk));
	jdff dff_B_O16Gc5wT2_2(.din(w_dff_B_9h6NlaLw6_2),.dout(w_dff_B_O16Gc5wT2_2),.clk(gclk));
	jdff dff_B_5IcWhh5n7_2(.din(w_dff_B_O16Gc5wT2_2),.dout(w_dff_B_5IcWhh5n7_2),.clk(gclk));
	jdff dff_B_hjkZlS5N2_2(.din(w_dff_B_5IcWhh5n7_2),.dout(w_dff_B_hjkZlS5N2_2),.clk(gclk));
	jdff dff_B_14T0t1lH1_2(.din(w_dff_B_hjkZlS5N2_2),.dout(w_dff_B_14T0t1lH1_2),.clk(gclk));
	jdff dff_B_0JAEdSmU9_2(.din(w_dff_B_14T0t1lH1_2),.dout(w_dff_B_0JAEdSmU9_2),.clk(gclk));
	jdff dff_B_XTMiFsPL7_2(.din(w_dff_B_0JAEdSmU9_2),.dout(w_dff_B_XTMiFsPL7_2),.clk(gclk));
	jdff dff_B_wyNebLeA6_2(.din(w_dff_B_XTMiFsPL7_2),.dout(w_dff_B_wyNebLeA6_2),.clk(gclk));
	jdff dff_B_MJSKrjHa7_2(.din(w_dff_B_wyNebLeA6_2),.dout(w_dff_B_MJSKrjHa7_2),.clk(gclk));
	jdff dff_B_oMDPKNTq5_2(.din(w_dff_B_MJSKrjHa7_2),.dout(w_dff_B_oMDPKNTq5_2),.clk(gclk));
	jdff dff_B_sZXq265h8_2(.din(w_dff_B_oMDPKNTq5_2),.dout(w_dff_B_sZXq265h8_2),.clk(gclk));
	jdff dff_B_7jkSTk9B6_2(.din(w_dff_B_sZXq265h8_2),.dout(w_dff_B_7jkSTk9B6_2),.clk(gclk));
	jdff dff_B_VTnCxu1s2_1(.din(n720),.dout(w_dff_B_VTnCxu1s2_1),.clk(gclk));
	jdff dff_B_o38pbutf8_2(.din(n627),.dout(w_dff_B_o38pbutf8_2),.clk(gclk));
	jdff dff_B_mqHkqoQt4_2(.din(w_dff_B_o38pbutf8_2),.dout(w_dff_B_mqHkqoQt4_2),.clk(gclk));
	jdff dff_B_DvdHCQfH6_2(.din(w_dff_B_mqHkqoQt4_2),.dout(w_dff_B_DvdHCQfH6_2),.clk(gclk));
	jdff dff_B_jIPfL9T36_2(.din(w_dff_B_DvdHCQfH6_2),.dout(w_dff_B_jIPfL9T36_2),.clk(gclk));
	jdff dff_B_X7U5MrB34_2(.din(w_dff_B_jIPfL9T36_2),.dout(w_dff_B_X7U5MrB34_2),.clk(gclk));
	jdff dff_B_5W15h3EU7_2(.din(w_dff_B_X7U5MrB34_2),.dout(w_dff_B_5W15h3EU7_2),.clk(gclk));
	jdff dff_B_gztwS6fZ1_2(.din(w_dff_B_5W15h3EU7_2),.dout(w_dff_B_gztwS6fZ1_2),.clk(gclk));
	jdff dff_B_z4S3XMLE1_2(.din(w_dff_B_gztwS6fZ1_2),.dout(w_dff_B_z4S3XMLE1_2),.clk(gclk));
	jdff dff_B_RFLBCUDz3_2(.din(w_dff_B_z4S3XMLE1_2),.dout(w_dff_B_RFLBCUDz3_2),.clk(gclk));
	jdff dff_B_PauOrJSC1_2(.din(w_dff_B_RFLBCUDz3_2),.dout(w_dff_B_PauOrJSC1_2),.clk(gclk));
	jdff dff_B_zATPdLnJ5_2(.din(w_dff_B_PauOrJSC1_2),.dout(w_dff_B_zATPdLnJ5_2),.clk(gclk));
	jdff dff_B_5YYgbd1u8_2(.din(w_dff_B_zATPdLnJ5_2),.dout(w_dff_B_5YYgbd1u8_2),.clk(gclk));
	jdff dff_B_SN1BSypw1_2(.din(w_dff_B_5YYgbd1u8_2),.dout(w_dff_B_SN1BSypw1_2),.clk(gclk));
	jdff dff_B_LgNK6NPy1_2(.din(w_dff_B_SN1BSypw1_2),.dout(w_dff_B_LgNK6NPy1_2),.clk(gclk));
	jdff dff_B_mLM8j9FV1_2(.din(w_dff_B_LgNK6NPy1_2),.dout(w_dff_B_mLM8j9FV1_2),.clk(gclk));
	jdff dff_B_9GAvwy2G2_2(.din(w_dff_B_mLM8j9FV1_2),.dout(w_dff_B_9GAvwy2G2_2),.clk(gclk));
	jdff dff_B_8XIIRcp81_2(.din(w_dff_B_9GAvwy2G2_2),.dout(w_dff_B_8XIIRcp81_2),.clk(gclk));
	jdff dff_B_bhEX6O7d6_2(.din(w_dff_B_8XIIRcp81_2),.dout(w_dff_B_bhEX6O7d6_2),.clk(gclk));
	jdff dff_B_pwNRDr5u7_2(.din(w_dff_B_bhEX6O7d6_2),.dout(w_dff_B_pwNRDr5u7_2),.clk(gclk));
	jdff dff_B_HNJeLkKb6_2(.din(w_dff_B_pwNRDr5u7_2),.dout(w_dff_B_HNJeLkKb6_2),.clk(gclk));
	jdff dff_B_fyN3ZaDT0_2(.din(w_dff_B_HNJeLkKb6_2),.dout(w_dff_B_fyN3ZaDT0_2),.clk(gclk));
	jdff dff_B_EIspindm2_2(.din(w_dff_B_fyN3ZaDT0_2),.dout(w_dff_B_EIspindm2_2),.clk(gclk));
	jdff dff_B_hWChproN0_2(.din(w_dff_B_EIspindm2_2),.dout(w_dff_B_hWChproN0_2),.clk(gclk));
	jdff dff_B_HJozdlbv8_2(.din(w_dff_B_hWChproN0_2),.dout(w_dff_B_HJozdlbv8_2),.clk(gclk));
	jdff dff_B_DGB6GK2U4_1(.din(n628),.dout(w_dff_B_DGB6GK2U4_1),.clk(gclk));
	jdff dff_B_z5Mrl2d49_2(.din(n542),.dout(w_dff_B_z5Mrl2d49_2),.clk(gclk));
	jdff dff_B_ji1O4XeW8_2(.din(w_dff_B_z5Mrl2d49_2),.dout(w_dff_B_ji1O4XeW8_2),.clk(gclk));
	jdff dff_B_OGC6xtUR8_2(.din(w_dff_B_ji1O4XeW8_2),.dout(w_dff_B_OGC6xtUR8_2),.clk(gclk));
	jdff dff_B_U6VqR7Tu6_2(.din(w_dff_B_OGC6xtUR8_2),.dout(w_dff_B_U6VqR7Tu6_2),.clk(gclk));
	jdff dff_B_BAP7ZMkT0_2(.din(w_dff_B_U6VqR7Tu6_2),.dout(w_dff_B_BAP7ZMkT0_2),.clk(gclk));
	jdff dff_B_EnyMka5z8_2(.din(w_dff_B_BAP7ZMkT0_2),.dout(w_dff_B_EnyMka5z8_2),.clk(gclk));
	jdff dff_B_SLbRyJW77_2(.din(w_dff_B_EnyMka5z8_2),.dout(w_dff_B_SLbRyJW77_2),.clk(gclk));
	jdff dff_B_TiEfzTcg3_2(.din(w_dff_B_SLbRyJW77_2),.dout(w_dff_B_TiEfzTcg3_2),.clk(gclk));
	jdff dff_B_xfIGiNse3_2(.din(w_dff_B_TiEfzTcg3_2),.dout(w_dff_B_xfIGiNse3_2),.clk(gclk));
	jdff dff_B_ZmuQ96UD1_2(.din(w_dff_B_xfIGiNse3_2),.dout(w_dff_B_ZmuQ96UD1_2),.clk(gclk));
	jdff dff_B_x3eC20vg7_2(.din(w_dff_B_ZmuQ96UD1_2),.dout(w_dff_B_x3eC20vg7_2),.clk(gclk));
	jdff dff_B_AgPuE6J71_2(.din(w_dff_B_x3eC20vg7_2),.dout(w_dff_B_AgPuE6J71_2),.clk(gclk));
	jdff dff_B_TJfFCRQk3_2(.din(w_dff_B_AgPuE6J71_2),.dout(w_dff_B_TJfFCRQk3_2),.clk(gclk));
	jdff dff_B_fcLC42gh6_2(.din(w_dff_B_TJfFCRQk3_2),.dout(w_dff_B_fcLC42gh6_2),.clk(gclk));
	jdff dff_B_9prlxDHj9_2(.din(w_dff_B_fcLC42gh6_2),.dout(w_dff_B_9prlxDHj9_2),.clk(gclk));
	jdff dff_B_4xxIRRzl4_2(.din(w_dff_B_9prlxDHj9_2),.dout(w_dff_B_4xxIRRzl4_2),.clk(gclk));
	jdff dff_B_RBwEnbfL7_2(.din(w_dff_B_4xxIRRzl4_2),.dout(w_dff_B_RBwEnbfL7_2),.clk(gclk));
	jdff dff_B_yCQscvb85_2(.din(w_dff_B_RBwEnbfL7_2),.dout(w_dff_B_yCQscvb85_2),.clk(gclk));
	jdff dff_B_OqccJEAx6_2(.din(w_dff_B_yCQscvb85_2),.dout(w_dff_B_OqccJEAx6_2),.clk(gclk));
	jdff dff_B_eItrhepZ7_2(.din(w_dff_B_OqccJEAx6_2),.dout(w_dff_B_eItrhepZ7_2),.clk(gclk));
	jdff dff_B_XJ4UuzMf0_2(.din(w_dff_B_eItrhepZ7_2),.dout(w_dff_B_XJ4UuzMf0_2),.clk(gclk));
	jdff dff_B_CtXZPoD54_2(.din(w_dff_B_XJ4UuzMf0_2),.dout(w_dff_B_CtXZPoD54_2),.clk(gclk));
	jdff dff_B_AYEMt2pb5_1(.din(n543),.dout(w_dff_B_AYEMt2pb5_1),.clk(gclk));
	jdff dff_B_yiFikY6S0_2(.din(n464),.dout(w_dff_B_yiFikY6S0_2),.clk(gclk));
	jdff dff_B_9GWHbyoQ9_2(.din(w_dff_B_yiFikY6S0_2),.dout(w_dff_B_9GWHbyoQ9_2),.clk(gclk));
	jdff dff_B_mDMsgMjl5_2(.din(w_dff_B_9GWHbyoQ9_2),.dout(w_dff_B_mDMsgMjl5_2),.clk(gclk));
	jdff dff_B_nnbUSo3H8_2(.din(w_dff_B_mDMsgMjl5_2),.dout(w_dff_B_nnbUSo3H8_2),.clk(gclk));
	jdff dff_B_1w7uZ2C55_2(.din(w_dff_B_nnbUSo3H8_2),.dout(w_dff_B_1w7uZ2C55_2),.clk(gclk));
	jdff dff_B_hwRikIEi1_2(.din(w_dff_B_1w7uZ2C55_2),.dout(w_dff_B_hwRikIEi1_2),.clk(gclk));
	jdff dff_B_0DFTMkaz9_2(.din(w_dff_B_hwRikIEi1_2),.dout(w_dff_B_0DFTMkaz9_2),.clk(gclk));
	jdff dff_B_0VweNF2b0_2(.din(w_dff_B_0DFTMkaz9_2),.dout(w_dff_B_0VweNF2b0_2),.clk(gclk));
	jdff dff_B_A3vMFwbm9_2(.din(w_dff_B_0VweNF2b0_2),.dout(w_dff_B_A3vMFwbm9_2),.clk(gclk));
	jdff dff_B_EYYS5jdu4_2(.din(w_dff_B_A3vMFwbm9_2),.dout(w_dff_B_EYYS5jdu4_2),.clk(gclk));
	jdff dff_B_NCfSB1RD5_2(.din(w_dff_B_EYYS5jdu4_2),.dout(w_dff_B_NCfSB1RD5_2),.clk(gclk));
	jdff dff_B_ZsEOCC6H8_2(.din(w_dff_B_NCfSB1RD5_2),.dout(w_dff_B_ZsEOCC6H8_2),.clk(gclk));
	jdff dff_B_6I6clgRr8_2(.din(w_dff_B_ZsEOCC6H8_2),.dout(w_dff_B_6I6clgRr8_2),.clk(gclk));
	jdff dff_B_2MaNKVGT2_2(.din(w_dff_B_6I6clgRr8_2),.dout(w_dff_B_2MaNKVGT2_2),.clk(gclk));
	jdff dff_B_bpGrHt7i6_2(.din(w_dff_B_2MaNKVGT2_2),.dout(w_dff_B_bpGrHt7i6_2),.clk(gclk));
	jdff dff_B_VXpvDMr24_2(.din(w_dff_B_bpGrHt7i6_2),.dout(w_dff_B_VXpvDMr24_2),.clk(gclk));
	jdff dff_B_4ZTR1YRD0_2(.din(w_dff_B_VXpvDMr24_2),.dout(w_dff_B_4ZTR1YRD0_2),.clk(gclk));
	jdff dff_B_SOxsZYhb7_2(.din(w_dff_B_4ZTR1YRD0_2),.dout(w_dff_B_SOxsZYhb7_2),.clk(gclk));
	jdff dff_B_ztEKzG725_2(.din(w_dff_B_SOxsZYhb7_2),.dout(w_dff_B_ztEKzG725_2),.clk(gclk));
	jdff dff_B_48wM55a46_2(.din(w_dff_B_ztEKzG725_2),.dout(w_dff_B_48wM55a46_2),.clk(gclk));
	jdff dff_B_JRaUOXWj3_1(.din(n465),.dout(w_dff_B_JRaUOXWj3_1),.clk(gclk));
	jdff dff_B_o3o5kmgZ9_2(.din(n393),.dout(w_dff_B_o3o5kmgZ9_2),.clk(gclk));
	jdff dff_B_i0dHUurS3_2(.din(w_dff_B_o3o5kmgZ9_2),.dout(w_dff_B_i0dHUurS3_2),.clk(gclk));
	jdff dff_B_92YhrZOP6_2(.din(w_dff_B_i0dHUurS3_2),.dout(w_dff_B_92YhrZOP6_2),.clk(gclk));
	jdff dff_B_WUM9aKaa4_2(.din(w_dff_B_92YhrZOP6_2),.dout(w_dff_B_WUM9aKaa4_2),.clk(gclk));
	jdff dff_B_n4bOWrrF5_2(.din(w_dff_B_WUM9aKaa4_2),.dout(w_dff_B_n4bOWrrF5_2),.clk(gclk));
	jdff dff_B_dNzqswh10_2(.din(w_dff_B_n4bOWrrF5_2),.dout(w_dff_B_dNzqswh10_2),.clk(gclk));
	jdff dff_B_InYXbte39_2(.din(w_dff_B_dNzqswh10_2),.dout(w_dff_B_InYXbte39_2),.clk(gclk));
	jdff dff_B_C2hvYceW0_2(.din(w_dff_B_InYXbte39_2),.dout(w_dff_B_C2hvYceW0_2),.clk(gclk));
	jdff dff_B_Iak6MvXc4_2(.din(w_dff_B_C2hvYceW0_2),.dout(w_dff_B_Iak6MvXc4_2),.clk(gclk));
	jdff dff_B_icPAnBW05_2(.din(w_dff_B_Iak6MvXc4_2),.dout(w_dff_B_icPAnBW05_2),.clk(gclk));
	jdff dff_B_lOru7j3E7_2(.din(w_dff_B_icPAnBW05_2),.dout(w_dff_B_lOru7j3E7_2),.clk(gclk));
	jdff dff_B_hnmhJOxM1_2(.din(w_dff_B_lOru7j3E7_2),.dout(w_dff_B_hnmhJOxM1_2),.clk(gclk));
	jdff dff_B_VaZbsnba9_2(.din(w_dff_B_hnmhJOxM1_2),.dout(w_dff_B_VaZbsnba9_2),.clk(gclk));
	jdff dff_B_Oxu1mLrj6_2(.din(w_dff_B_VaZbsnba9_2),.dout(w_dff_B_Oxu1mLrj6_2),.clk(gclk));
	jdff dff_B_SUxmqice2_2(.din(w_dff_B_Oxu1mLrj6_2),.dout(w_dff_B_SUxmqice2_2),.clk(gclk));
	jdff dff_B_Qbc2p17A7_2(.din(w_dff_B_SUxmqice2_2),.dout(w_dff_B_Qbc2p17A7_2),.clk(gclk));
	jdff dff_B_j48qRoWx6_2(.din(w_dff_B_Qbc2p17A7_2),.dout(w_dff_B_j48qRoWx6_2),.clk(gclk));
	jdff dff_B_fgyzPuhR6_2(.din(w_dff_B_j48qRoWx6_2),.dout(w_dff_B_fgyzPuhR6_2),.clk(gclk));
	jdff dff_B_qwUALIAQ9_2(.din(n396),.dout(w_dff_B_qwUALIAQ9_2),.clk(gclk));
	jdff dff_B_vWAWZdc59_2(.din(w_dff_B_qwUALIAQ9_2),.dout(w_dff_B_vWAWZdc59_2),.clk(gclk));
	jdff dff_B_N4sh3q5e5_2(.din(w_dff_B_vWAWZdc59_2),.dout(w_dff_B_N4sh3q5e5_2),.clk(gclk));
	jdff dff_B_P93Tff5z4_1(.din(n394),.dout(w_dff_B_P93Tff5z4_1),.clk(gclk));
	jdff dff_B_7sBlSo2X7_2(.din(n330),.dout(w_dff_B_7sBlSo2X7_2),.clk(gclk));
	jdff dff_B_dD1y967m9_2(.din(w_dff_B_7sBlSo2X7_2),.dout(w_dff_B_dD1y967m9_2),.clk(gclk));
	jdff dff_B_AC9zETx47_2(.din(w_dff_B_dD1y967m9_2),.dout(w_dff_B_AC9zETx47_2),.clk(gclk));
	jdff dff_B_JvXKLkmO7_2(.din(w_dff_B_AC9zETx47_2),.dout(w_dff_B_JvXKLkmO7_2),.clk(gclk));
	jdff dff_B_WjND6SVT6_2(.din(w_dff_B_JvXKLkmO7_2),.dout(w_dff_B_WjND6SVT6_2),.clk(gclk));
	jdff dff_B_Aga9P3Bs4_2(.din(w_dff_B_WjND6SVT6_2),.dout(w_dff_B_Aga9P3Bs4_2),.clk(gclk));
	jdff dff_B_o3xOySRJ2_2(.din(w_dff_B_Aga9P3Bs4_2),.dout(w_dff_B_o3xOySRJ2_2),.clk(gclk));
	jdff dff_B_QLSsXnrH2_2(.din(w_dff_B_o3xOySRJ2_2),.dout(w_dff_B_QLSsXnrH2_2),.clk(gclk));
	jdff dff_B_vsFXu0EJ6_2(.din(w_dff_B_QLSsXnrH2_2),.dout(w_dff_B_vsFXu0EJ6_2),.clk(gclk));
	jdff dff_B_iwAi1GUU6_2(.din(w_dff_B_vsFXu0EJ6_2),.dout(w_dff_B_iwAi1GUU6_2),.clk(gclk));
	jdff dff_B_oxmRtnfM1_2(.din(w_dff_B_iwAi1GUU6_2),.dout(w_dff_B_oxmRtnfM1_2),.clk(gclk));
	jdff dff_B_VCudCSLW9_2(.din(w_dff_B_oxmRtnfM1_2),.dout(w_dff_B_VCudCSLW9_2),.clk(gclk));
	jdff dff_B_XG3grkrj8_2(.din(w_dff_B_VCudCSLW9_2),.dout(w_dff_B_XG3grkrj8_2),.clk(gclk));
	jdff dff_B_a6aAry2s3_1(.din(n331),.dout(w_dff_B_a6aAry2s3_1),.clk(gclk));
	jdff dff_B_6BgSjQ4p0_2(.din(n274),.dout(w_dff_B_6BgSjQ4p0_2),.clk(gclk));
	jdff dff_B_wSwAlr9b4_2(.din(w_dff_B_6BgSjQ4p0_2),.dout(w_dff_B_wSwAlr9b4_2),.clk(gclk));
	jdff dff_B_5xNQ7vcN1_2(.din(w_dff_B_wSwAlr9b4_2),.dout(w_dff_B_5xNQ7vcN1_2),.clk(gclk));
	jdff dff_B_BMKZfG7x8_2(.din(w_dff_B_5xNQ7vcN1_2),.dout(w_dff_B_BMKZfG7x8_2),.clk(gclk));
	jdff dff_B_dITPWEAj9_2(.din(w_dff_B_BMKZfG7x8_2),.dout(w_dff_B_dITPWEAj9_2),.clk(gclk));
	jdff dff_B_goRfSAGP9_2(.din(w_dff_B_dITPWEAj9_2),.dout(w_dff_B_goRfSAGP9_2),.clk(gclk));
	jdff dff_B_7hBaRknf8_2(.din(w_dff_B_goRfSAGP9_2),.dout(w_dff_B_7hBaRknf8_2),.clk(gclk));
	jdff dff_B_uUbNrxhr0_2(.din(w_dff_B_7hBaRknf8_2),.dout(w_dff_B_uUbNrxhr0_2),.clk(gclk));
	jdff dff_B_ePYffLUN5_2(.din(w_dff_B_uUbNrxhr0_2),.dout(w_dff_B_ePYffLUN5_2),.clk(gclk));
	jdff dff_B_XL44WUPg4_2(.din(w_dff_B_ePYffLUN5_2),.dout(w_dff_B_XL44WUPg4_2),.clk(gclk));
	jdff dff_B_aOXfa8sz8_2(.din(w_dff_B_XL44WUPg4_2),.dout(w_dff_B_aOXfa8sz8_2),.clk(gclk));
	jdff dff_B_179JyEBS4_1(.din(n275),.dout(w_dff_B_179JyEBS4_1),.clk(gclk));
	jdff dff_B_wgfFPKcQ8_2(.din(n225),.dout(w_dff_B_wgfFPKcQ8_2),.clk(gclk));
	jdff dff_B_4Mkdh8L65_2(.din(w_dff_B_wgfFPKcQ8_2),.dout(w_dff_B_4Mkdh8L65_2),.clk(gclk));
	jdff dff_B_uzE8JzXO6_2(.din(w_dff_B_4Mkdh8L65_2),.dout(w_dff_B_uzE8JzXO6_2),.clk(gclk));
	jdff dff_B_Cx86ky2u9_2(.din(w_dff_B_uzE8JzXO6_2),.dout(w_dff_B_Cx86ky2u9_2),.clk(gclk));
	jdff dff_B_JEhgz6Oy5_2(.din(w_dff_B_Cx86ky2u9_2),.dout(w_dff_B_JEhgz6Oy5_2),.clk(gclk));
	jdff dff_B_wESYyZfT3_2(.din(w_dff_B_JEhgz6Oy5_2),.dout(w_dff_B_wESYyZfT3_2),.clk(gclk));
	jdff dff_B_6SAplVxm9_2(.din(w_dff_B_wESYyZfT3_2),.dout(w_dff_B_6SAplVxm9_2),.clk(gclk));
	jdff dff_B_tC5J9qza7_2(.din(w_dff_B_6SAplVxm9_2),.dout(w_dff_B_tC5J9qza7_2),.clk(gclk));
	jdff dff_B_KZLo3TkJ9_2(.din(w_dff_B_tC5J9qza7_2),.dout(w_dff_B_KZLo3TkJ9_2),.clk(gclk));
	jdff dff_B_EK6M9CMC1_1(.din(n226),.dout(w_dff_B_EK6M9CMC1_1),.clk(gclk));
	jdff dff_B_eVakjd8v3_2(.din(n183),.dout(w_dff_B_eVakjd8v3_2),.clk(gclk));
	jdff dff_B_sABgkMfb1_2(.din(w_dff_B_eVakjd8v3_2),.dout(w_dff_B_sABgkMfb1_2),.clk(gclk));
	jdff dff_B_L8BxoCXC8_2(.din(w_dff_B_sABgkMfb1_2),.dout(w_dff_B_L8BxoCXC8_2),.clk(gclk));
	jdff dff_B_nx4Jfh7d1_2(.din(w_dff_B_L8BxoCXC8_2),.dout(w_dff_B_nx4Jfh7d1_2),.clk(gclk));
	jdff dff_B_MI2MR9K84_2(.din(w_dff_B_nx4Jfh7d1_2),.dout(w_dff_B_MI2MR9K84_2),.clk(gclk));
	jdff dff_B_YljsIb8x7_2(.din(w_dff_B_MI2MR9K84_2),.dout(w_dff_B_YljsIb8x7_2),.clk(gclk));
	jdff dff_B_a0xbI5MR9_2(.din(w_dff_B_YljsIb8x7_2),.dout(w_dff_B_a0xbI5MR9_2),.clk(gclk));
	jdff dff_B_0mJuPkMW1_1(.din(n184),.dout(w_dff_B_0mJuPkMW1_1),.clk(gclk));
	jdff dff_B_pycAoolc5_2(.din(n148),.dout(w_dff_B_pycAoolc5_2),.clk(gclk));
	jdff dff_B_jtqD1miP2_2(.din(w_dff_B_pycAoolc5_2),.dout(w_dff_B_jtqD1miP2_2),.clk(gclk));
	jdff dff_B_BB597h2Q4_2(.din(w_dff_B_jtqD1miP2_2),.dout(w_dff_B_BB597h2Q4_2),.clk(gclk));
	jdff dff_B_si6JPCcA0_2(.din(w_dff_B_BB597h2Q4_2),.dout(w_dff_B_si6JPCcA0_2),.clk(gclk));
	jdff dff_B_U9BSC4ub3_2(.din(w_dff_B_si6JPCcA0_2),.dout(w_dff_B_U9BSC4ub3_2),.clk(gclk));
	jdff dff_B_JOEeLthO3_1(.din(n150),.dout(w_dff_B_JOEeLthO3_1),.clk(gclk));
	jdff dff_B_bJ3a7PNT8_2(.din(n119),.dout(w_dff_B_bJ3a7PNT8_2),.clk(gclk));
	jdff dff_B_7EgRI1TZ8_2(.din(w_dff_B_bJ3a7PNT8_2),.dout(w_dff_B_7EgRI1TZ8_2),.clk(gclk));
	jdff dff_B_AmgMx0zO2_2(.din(w_dff_B_7EgRI1TZ8_2),.dout(w_dff_B_AmgMx0zO2_2),.clk(gclk));
	jdff dff_B_2e37WqoN8_0(.din(n126),.dout(w_dff_B_2e37WqoN8_0),.clk(gclk));
	jdff dff_B_KG6L1ole9_0(.din(w_dff_B_2e37WqoN8_0),.dout(w_dff_B_KG6L1ole9_0),.clk(gclk));
	jdff dff_B_R0DWTPDp5_2(.din(n120),.dout(w_dff_B_R0DWTPDp5_2),.clk(gclk));
	jdff dff_B_XyxqOr217_2(.din(w_dff_B_R0DWTPDp5_2),.dout(w_dff_B_XyxqOr217_2),.clk(gclk));
	jdff dff_A_XyCh9jAo8_1(.dout(w_n1294_0[1]),.din(w_dff_A_XyCh9jAo8_1),.clk(gclk));
	jdff dff_B_j8tgBVSe0_1(.din(n1214),.dout(w_dff_B_j8tgBVSe0_1),.clk(gclk));
	jdff dff_B_CryD6Cfq3_1(.din(w_dff_B_j8tgBVSe0_1),.dout(w_dff_B_CryD6Cfq3_1),.clk(gclk));
	jdff dff_B_oilcDNtd4_2(.din(n1120),.dout(w_dff_B_oilcDNtd4_2),.clk(gclk));
	jdff dff_B_15zZ8kM33_2(.din(w_dff_B_oilcDNtd4_2),.dout(w_dff_B_15zZ8kM33_2),.clk(gclk));
	jdff dff_B_UbL0sGHz7_2(.din(w_dff_B_15zZ8kM33_2),.dout(w_dff_B_UbL0sGHz7_2),.clk(gclk));
	jdff dff_B_cdtzEnhi5_2(.din(w_dff_B_UbL0sGHz7_2),.dout(w_dff_B_cdtzEnhi5_2),.clk(gclk));
	jdff dff_B_PRJkIcra5_2(.din(w_dff_B_cdtzEnhi5_2),.dout(w_dff_B_PRJkIcra5_2),.clk(gclk));
	jdff dff_B_FzXg4FmR2_2(.din(w_dff_B_PRJkIcra5_2),.dout(w_dff_B_FzXg4FmR2_2),.clk(gclk));
	jdff dff_B_vTFCoGC55_2(.din(w_dff_B_FzXg4FmR2_2),.dout(w_dff_B_vTFCoGC55_2),.clk(gclk));
	jdff dff_B_wqfXGH9U4_2(.din(w_dff_B_vTFCoGC55_2),.dout(w_dff_B_wqfXGH9U4_2),.clk(gclk));
	jdff dff_B_MsFJ0Z9w4_2(.din(w_dff_B_wqfXGH9U4_2),.dout(w_dff_B_MsFJ0Z9w4_2),.clk(gclk));
	jdff dff_B_qMH7nCs17_2(.din(w_dff_B_MsFJ0Z9w4_2),.dout(w_dff_B_qMH7nCs17_2),.clk(gclk));
	jdff dff_B_nVJfKJMQ2_2(.din(w_dff_B_qMH7nCs17_2),.dout(w_dff_B_nVJfKJMQ2_2),.clk(gclk));
	jdff dff_B_paKERQX20_2(.din(w_dff_B_nVJfKJMQ2_2),.dout(w_dff_B_paKERQX20_2),.clk(gclk));
	jdff dff_B_7vOWv20M4_2(.din(w_dff_B_paKERQX20_2),.dout(w_dff_B_7vOWv20M4_2),.clk(gclk));
	jdff dff_B_i9DAn7Wh3_2(.din(w_dff_B_7vOWv20M4_2),.dout(w_dff_B_i9DAn7Wh3_2),.clk(gclk));
	jdff dff_B_cBjAkNjJ5_2(.din(w_dff_B_i9DAn7Wh3_2),.dout(w_dff_B_cBjAkNjJ5_2),.clk(gclk));
	jdff dff_B_a54AEM1u5_2(.din(w_dff_B_cBjAkNjJ5_2),.dout(w_dff_B_a54AEM1u5_2),.clk(gclk));
	jdff dff_B_YYsTaknn6_2(.din(w_dff_B_a54AEM1u5_2),.dout(w_dff_B_YYsTaknn6_2),.clk(gclk));
	jdff dff_B_rRDNzS7j6_2(.din(w_dff_B_YYsTaknn6_2),.dout(w_dff_B_rRDNzS7j6_2),.clk(gclk));
	jdff dff_B_TLRYqo0p6_2(.din(w_dff_B_rRDNzS7j6_2),.dout(w_dff_B_TLRYqo0p6_2),.clk(gclk));
	jdff dff_B_Wy9Y70nD2_2(.din(w_dff_B_TLRYqo0p6_2),.dout(w_dff_B_Wy9Y70nD2_2),.clk(gclk));
	jdff dff_B_CxVTMGzw1_2(.din(w_dff_B_Wy9Y70nD2_2),.dout(w_dff_B_CxVTMGzw1_2),.clk(gclk));
	jdff dff_B_OWZ2oYMB0_2(.din(w_dff_B_CxVTMGzw1_2),.dout(w_dff_B_OWZ2oYMB0_2),.clk(gclk));
	jdff dff_B_aBIHBdYF2_2(.din(w_dff_B_OWZ2oYMB0_2),.dout(w_dff_B_aBIHBdYF2_2),.clk(gclk));
	jdff dff_B_cWwPpj9i9_2(.din(w_dff_B_aBIHBdYF2_2),.dout(w_dff_B_cWwPpj9i9_2),.clk(gclk));
	jdff dff_B_3mRUBu190_2(.din(w_dff_B_cWwPpj9i9_2),.dout(w_dff_B_3mRUBu190_2),.clk(gclk));
	jdff dff_B_PzJR96K57_2(.din(w_dff_B_3mRUBu190_2),.dout(w_dff_B_PzJR96K57_2),.clk(gclk));
	jdff dff_B_ZLBt1Kri8_2(.din(w_dff_B_PzJR96K57_2),.dout(w_dff_B_ZLBt1Kri8_2),.clk(gclk));
	jdff dff_B_FUIbMm6V1_2(.din(w_dff_B_ZLBt1Kri8_2),.dout(w_dff_B_FUIbMm6V1_2),.clk(gclk));
	jdff dff_B_P66wPTx76_2(.din(w_dff_B_FUIbMm6V1_2),.dout(w_dff_B_P66wPTx76_2),.clk(gclk));
	jdff dff_B_kRAFBaob1_2(.din(w_dff_B_P66wPTx76_2),.dout(w_dff_B_kRAFBaob1_2),.clk(gclk));
	jdff dff_B_FXSYPZiZ0_2(.din(w_dff_B_kRAFBaob1_2),.dout(w_dff_B_FXSYPZiZ0_2),.clk(gclk));
	jdff dff_B_W0Fm7O9J0_2(.din(w_dff_B_FXSYPZiZ0_2),.dout(w_dff_B_W0Fm7O9J0_2),.clk(gclk));
	jdff dff_B_gxhM8V879_2(.din(w_dff_B_W0Fm7O9J0_2),.dout(w_dff_B_gxhM8V879_2),.clk(gclk));
	jdff dff_B_zVNRmedN4_2(.din(w_dff_B_gxhM8V879_2),.dout(w_dff_B_zVNRmedN4_2),.clk(gclk));
	jdff dff_B_IcVXHOmB8_2(.din(w_dff_B_zVNRmedN4_2),.dout(w_dff_B_IcVXHOmB8_2),.clk(gclk));
	jdff dff_B_z2eft3Hx1_2(.din(n1023),.dout(w_dff_B_z2eft3Hx1_2),.clk(gclk));
	jdff dff_B_5hCCQ6uO8_2(.din(w_dff_B_z2eft3Hx1_2),.dout(w_dff_B_5hCCQ6uO8_2),.clk(gclk));
	jdff dff_B_R6efCo3Q3_2(.din(w_dff_B_5hCCQ6uO8_2),.dout(w_dff_B_R6efCo3Q3_2),.clk(gclk));
	jdff dff_B_HHg7LBou9_2(.din(w_dff_B_R6efCo3Q3_2),.dout(w_dff_B_HHg7LBou9_2),.clk(gclk));
	jdff dff_B_OZPvsSCI9_2(.din(w_dff_B_HHg7LBou9_2),.dout(w_dff_B_OZPvsSCI9_2),.clk(gclk));
	jdff dff_B_cOmbRTJQ6_2(.din(w_dff_B_OZPvsSCI9_2),.dout(w_dff_B_cOmbRTJQ6_2),.clk(gclk));
	jdff dff_B_JE1vqca74_2(.din(w_dff_B_cOmbRTJQ6_2),.dout(w_dff_B_JE1vqca74_2),.clk(gclk));
	jdff dff_B_BjBDuWrd8_2(.din(w_dff_B_JE1vqca74_2),.dout(w_dff_B_BjBDuWrd8_2),.clk(gclk));
	jdff dff_B_vs2VIFTH1_2(.din(w_dff_B_BjBDuWrd8_2),.dout(w_dff_B_vs2VIFTH1_2),.clk(gclk));
	jdff dff_B_1Uf69JuG7_2(.din(w_dff_B_vs2VIFTH1_2),.dout(w_dff_B_1Uf69JuG7_2),.clk(gclk));
	jdff dff_B_SnvcmMeL2_2(.din(w_dff_B_1Uf69JuG7_2),.dout(w_dff_B_SnvcmMeL2_2),.clk(gclk));
	jdff dff_B_Y9GmZhvq2_2(.din(w_dff_B_SnvcmMeL2_2),.dout(w_dff_B_Y9GmZhvq2_2),.clk(gclk));
	jdff dff_B_JDytO8bX0_2(.din(w_dff_B_Y9GmZhvq2_2),.dout(w_dff_B_JDytO8bX0_2),.clk(gclk));
	jdff dff_B_9jhhSUmO9_2(.din(w_dff_B_JDytO8bX0_2),.dout(w_dff_B_9jhhSUmO9_2),.clk(gclk));
	jdff dff_B_sBmjEpyi9_2(.din(w_dff_B_9jhhSUmO9_2),.dout(w_dff_B_sBmjEpyi9_2),.clk(gclk));
	jdff dff_B_rn2e8mvC2_2(.din(w_dff_B_sBmjEpyi9_2),.dout(w_dff_B_rn2e8mvC2_2),.clk(gclk));
	jdff dff_B_sGVMbOxG4_2(.din(w_dff_B_rn2e8mvC2_2),.dout(w_dff_B_sGVMbOxG4_2),.clk(gclk));
	jdff dff_B_pM8lxuAE9_2(.din(w_dff_B_sGVMbOxG4_2),.dout(w_dff_B_pM8lxuAE9_2),.clk(gclk));
	jdff dff_B_YtEAZOW73_2(.din(w_dff_B_pM8lxuAE9_2),.dout(w_dff_B_YtEAZOW73_2),.clk(gclk));
	jdff dff_B_93O3wBcX7_2(.din(w_dff_B_YtEAZOW73_2),.dout(w_dff_B_93O3wBcX7_2),.clk(gclk));
	jdff dff_B_bWjjSqsC9_2(.din(w_dff_B_93O3wBcX7_2),.dout(w_dff_B_bWjjSqsC9_2),.clk(gclk));
	jdff dff_B_sRdUSWLX1_2(.din(w_dff_B_bWjjSqsC9_2),.dout(w_dff_B_sRdUSWLX1_2),.clk(gclk));
	jdff dff_B_gB2azBy89_2(.din(w_dff_B_sRdUSWLX1_2),.dout(w_dff_B_gB2azBy89_2),.clk(gclk));
	jdff dff_B_RP9SRDAQ2_2(.din(w_dff_B_gB2azBy89_2),.dout(w_dff_B_RP9SRDAQ2_2),.clk(gclk));
	jdff dff_B_I0ZgTe0E6_2(.din(w_dff_B_RP9SRDAQ2_2),.dout(w_dff_B_I0ZgTe0E6_2),.clk(gclk));
	jdff dff_B_dfF5PRfQ1_2(.din(w_dff_B_I0ZgTe0E6_2),.dout(w_dff_B_dfF5PRfQ1_2),.clk(gclk));
	jdff dff_B_yA2vWf9f0_2(.din(w_dff_B_dfF5PRfQ1_2),.dout(w_dff_B_yA2vWf9f0_2),.clk(gclk));
	jdff dff_B_OLpM4IRT2_2(.din(w_dff_B_yA2vWf9f0_2),.dout(w_dff_B_OLpM4IRT2_2),.clk(gclk));
	jdff dff_B_8hVdvtN82_2(.din(w_dff_B_OLpM4IRT2_2),.dout(w_dff_B_8hVdvtN82_2),.clk(gclk));
	jdff dff_B_rBlPwu5Q4_2(.din(w_dff_B_8hVdvtN82_2),.dout(w_dff_B_rBlPwu5Q4_2),.clk(gclk));
	jdff dff_B_pyJdQncl1_2(.din(w_dff_B_rBlPwu5Q4_2),.dout(w_dff_B_pyJdQncl1_2),.clk(gclk));
	jdff dff_B_WGkBMv0o2_2(.din(w_dff_B_pyJdQncl1_2),.dout(w_dff_B_WGkBMv0o2_2),.clk(gclk));
	jdff dff_B_sNTjJaJO2_1(.din(n1024),.dout(w_dff_B_sNTjJaJO2_1),.clk(gclk));
	jdff dff_B_lMtLiVv80_2(.din(n924),.dout(w_dff_B_lMtLiVv80_2),.clk(gclk));
	jdff dff_B_Kny7VouC8_2(.din(w_dff_B_lMtLiVv80_2),.dout(w_dff_B_Kny7VouC8_2),.clk(gclk));
	jdff dff_B_dZSAP3R21_2(.din(w_dff_B_Kny7VouC8_2),.dout(w_dff_B_dZSAP3R21_2),.clk(gclk));
	jdff dff_B_OwvQ85aW2_2(.din(w_dff_B_dZSAP3R21_2),.dout(w_dff_B_OwvQ85aW2_2),.clk(gclk));
	jdff dff_B_4uMYYScH7_2(.din(w_dff_B_OwvQ85aW2_2),.dout(w_dff_B_4uMYYScH7_2),.clk(gclk));
	jdff dff_B_v762xUcz5_2(.din(w_dff_B_4uMYYScH7_2),.dout(w_dff_B_v762xUcz5_2),.clk(gclk));
	jdff dff_B_OQC4Q1wz8_2(.din(w_dff_B_v762xUcz5_2),.dout(w_dff_B_OQC4Q1wz8_2),.clk(gclk));
	jdff dff_B_Lm7qDqoX9_2(.din(w_dff_B_OQC4Q1wz8_2),.dout(w_dff_B_Lm7qDqoX9_2),.clk(gclk));
	jdff dff_B_XSrmnJyZ8_2(.din(w_dff_B_Lm7qDqoX9_2),.dout(w_dff_B_XSrmnJyZ8_2),.clk(gclk));
	jdff dff_B_qWy7PIuP2_2(.din(w_dff_B_XSrmnJyZ8_2),.dout(w_dff_B_qWy7PIuP2_2),.clk(gclk));
	jdff dff_B_TaaW1kKq3_2(.din(w_dff_B_qWy7PIuP2_2),.dout(w_dff_B_TaaW1kKq3_2),.clk(gclk));
	jdff dff_B_E1vGASyh0_2(.din(w_dff_B_TaaW1kKq3_2),.dout(w_dff_B_E1vGASyh0_2),.clk(gclk));
	jdff dff_B_dvRv323c1_2(.din(w_dff_B_E1vGASyh0_2),.dout(w_dff_B_dvRv323c1_2),.clk(gclk));
	jdff dff_B_7IEjVGqe0_2(.din(w_dff_B_dvRv323c1_2),.dout(w_dff_B_7IEjVGqe0_2),.clk(gclk));
	jdff dff_B_deC93HoG7_2(.din(w_dff_B_7IEjVGqe0_2),.dout(w_dff_B_deC93HoG7_2),.clk(gclk));
	jdff dff_B_hwcygG2j6_2(.din(w_dff_B_deC93HoG7_2),.dout(w_dff_B_hwcygG2j6_2),.clk(gclk));
	jdff dff_B_WxEsqBZd6_2(.din(w_dff_B_hwcygG2j6_2),.dout(w_dff_B_WxEsqBZd6_2),.clk(gclk));
	jdff dff_B_PXrT6IEk6_2(.din(w_dff_B_WxEsqBZd6_2),.dout(w_dff_B_PXrT6IEk6_2),.clk(gclk));
	jdff dff_B_4PMjx43R2_2(.din(w_dff_B_PXrT6IEk6_2),.dout(w_dff_B_4PMjx43R2_2),.clk(gclk));
	jdff dff_B_uErkJBpM7_2(.din(w_dff_B_4PMjx43R2_2),.dout(w_dff_B_uErkJBpM7_2),.clk(gclk));
	jdff dff_B_GovHtXWP9_2(.din(w_dff_B_uErkJBpM7_2),.dout(w_dff_B_GovHtXWP9_2),.clk(gclk));
	jdff dff_B_T65xFP7s6_2(.din(w_dff_B_GovHtXWP9_2),.dout(w_dff_B_T65xFP7s6_2),.clk(gclk));
	jdff dff_B_lzAbEm1k0_2(.din(w_dff_B_T65xFP7s6_2),.dout(w_dff_B_lzAbEm1k0_2),.clk(gclk));
	jdff dff_B_ZP2hEZ8b5_2(.din(w_dff_B_lzAbEm1k0_2),.dout(w_dff_B_ZP2hEZ8b5_2),.clk(gclk));
	jdff dff_B_2k3mJCGL0_2(.din(w_dff_B_ZP2hEZ8b5_2),.dout(w_dff_B_2k3mJCGL0_2),.clk(gclk));
	jdff dff_B_3jQ5aiW55_2(.din(w_dff_B_2k3mJCGL0_2),.dout(w_dff_B_3jQ5aiW55_2),.clk(gclk));
	jdff dff_B_5rwIkS546_2(.din(w_dff_B_3jQ5aiW55_2),.dout(w_dff_B_5rwIkS546_2),.clk(gclk));
	jdff dff_B_8HzqBeLN7_2(.din(w_dff_B_5rwIkS546_2),.dout(w_dff_B_8HzqBeLN7_2),.clk(gclk));
	jdff dff_B_8XmM6ZQT5_1(.din(n925),.dout(w_dff_B_8XmM6ZQT5_1),.clk(gclk));
	jdff dff_B_oSUCqHoB3_2(.din(n822),.dout(w_dff_B_oSUCqHoB3_2),.clk(gclk));
	jdff dff_B_my9IvFGK1_2(.din(w_dff_B_oSUCqHoB3_2),.dout(w_dff_B_my9IvFGK1_2),.clk(gclk));
	jdff dff_B_YiQWaEqU1_2(.din(w_dff_B_my9IvFGK1_2),.dout(w_dff_B_YiQWaEqU1_2),.clk(gclk));
	jdff dff_B_u7lwJHaZ3_2(.din(w_dff_B_YiQWaEqU1_2),.dout(w_dff_B_u7lwJHaZ3_2),.clk(gclk));
	jdff dff_B_9t7pxeCg7_2(.din(w_dff_B_u7lwJHaZ3_2),.dout(w_dff_B_9t7pxeCg7_2),.clk(gclk));
	jdff dff_B_eUo8E2kU9_2(.din(w_dff_B_9t7pxeCg7_2),.dout(w_dff_B_eUo8E2kU9_2),.clk(gclk));
	jdff dff_B_LhF1i4Iz2_2(.din(w_dff_B_eUo8E2kU9_2),.dout(w_dff_B_LhF1i4Iz2_2),.clk(gclk));
	jdff dff_B_T8FOXlNM3_2(.din(w_dff_B_LhF1i4Iz2_2),.dout(w_dff_B_T8FOXlNM3_2),.clk(gclk));
	jdff dff_B_FYlCwDAt3_2(.din(w_dff_B_T8FOXlNM3_2),.dout(w_dff_B_FYlCwDAt3_2),.clk(gclk));
	jdff dff_B_1ZOHWq8R5_2(.din(w_dff_B_FYlCwDAt3_2),.dout(w_dff_B_1ZOHWq8R5_2),.clk(gclk));
	jdff dff_B_CwkQDiPc0_2(.din(w_dff_B_1ZOHWq8R5_2),.dout(w_dff_B_CwkQDiPc0_2),.clk(gclk));
	jdff dff_B_sYHeRNCk2_2(.din(w_dff_B_CwkQDiPc0_2),.dout(w_dff_B_sYHeRNCk2_2),.clk(gclk));
	jdff dff_B_aGjVGPL39_2(.din(w_dff_B_sYHeRNCk2_2),.dout(w_dff_B_aGjVGPL39_2),.clk(gclk));
	jdff dff_B_YOVeNT463_2(.din(w_dff_B_aGjVGPL39_2),.dout(w_dff_B_YOVeNT463_2),.clk(gclk));
	jdff dff_B_lnXAyMkZ6_2(.din(w_dff_B_YOVeNT463_2),.dout(w_dff_B_lnXAyMkZ6_2),.clk(gclk));
	jdff dff_B_i4E5udyy3_2(.din(w_dff_B_lnXAyMkZ6_2),.dout(w_dff_B_i4E5udyy3_2),.clk(gclk));
	jdff dff_B_7JvJSi6F0_2(.din(w_dff_B_i4E5udyy3_2),.dout(w_dff_B_7JvJSi6F0_2),.clk(gclk));
	jdff dff_B_wY4HfYA84_2(.din(w_dff_B_7JvJSi6F0_2),.dout(w_dff_B_wY4HfYA84_2),.clk(gclk));
	jdff dff_B_ZU3J9brb8_2(.din(w_dff_B_wY4HfYA84_2),.dout(w_dff_B_ZU3J9brb8_2),.clk(gclk));
	jdff dff_B_kgDElL1k1_2(.din(w_dff_B_ZU3J9brb8_2),.dout(w_dff_B_kgDElL1k1_2),.clk(gclk));
	jdff dff_B_beOPmkz14_2(.din(w_dff_B_kgDElL1k1_2),.dout(w_dff_B_beOPmkz14_2),.clk(gclk));
	jdff dff_B_aUowkf4D8_2(.din(w_dff_B_beOPmkz14_2),.dout(w_dff_B_aUowkf4D8_2),.clk(gclk));
	jdff dff_B_I3GgmAax8_2(.din(w_dff_B_aUowkf4D8_2),.dout(w_dff_B_I3GgmAax8_2),.clk(gclk));
	jdff dff_B_8rOpwDjW9_2(.din(w_dff_B_I3GgmAax8_2),.dout(w_dff_B_8rOpwDjW9_2),.clk(gclk));
	jdff dff_B_jji0w7VI7_2(.din(w_dff_B_8rOpwDjW9_2),.dout(w_dff_B_jji0w7VI7_2),.clk(gclk));
	jdff dff_B_h6QApWVR7_2(.din(w_dff_B_jji0w7VI7_2),.dout(w_dff_B_h6QApWVR7_2),.clk(gclk));
	jdff dff_B_WJTzbYWo0_1(.din(n823),.dout(w_dff_B_WJTzbYWo0_1),.clk(gclk));
	jdff dff_B_tBD6Qgke8_2(.din(n724),.dout(w_dff_B_tBD6Qgke8_2),.clk(gclk));
	jdff dff_B_U7EKFjLC5_2(.din(w_dff_B_tBD6Qgke8_2),.dout(w_dff_B_U7EKFjLC5_2),.clk(gclk));
	jdff dff_B_HSiI8sUR0_2(.din(w_dff_B_U7EKFjLC5_2),.dout(w_dff_B_HSiI8sUR0_2),.clk(gclk));
	jdff dff_B_RoZtcD7e1_2(.din(w_dff_B_HSiI8sUR0_2),.dout(w_dff_B_RoZtcD7e1_2),.clk(gclk));
	jdff dff_B_vuSO3C1n0_2(.din(w_dff_B_RoZtcD7e1_2),.dout(w_dff_B_vuSO3C1n0_2),.clk(gclk));
	jdff dff_B_0ik5aAyt4_2(.din(w_dff_B_vuSO3C1n0_2),.dout(w_dff_B_0ik5aAyt4_2),.clk(gclk));
	jdff dff_B_iew6PsxQ6_2(.din(w_dff_B_0ik5aAyt4_2),.dout(w_dff_B_iew6PsxQ6_2),.clk(gclk));
	jdff dff_B_BmsOrLXp2_2(.din(w_dff_B_iew6PsxQ6_2),.dout(w_dff_B_BmsOrLXp2_2),.clk(gclk));
	jdff dff_B_viRx4J9i1_2(.din(w_dff_B_BmsOrLXp2_2),.dout(w_dff_B_viRx4J9i1_2),.clk(gclk));
	jdff dff_B_sbPfn3469_2(.din(w_dff_B_viRx4J9i1_2),.dout(w_dff_B_sbPfn3469_2),.clk(gclk));
	jdff dff_B_pxMrcd2p7_2(.din(w_dff_B_sbPfn3469_2),.dout(w_dff_B_pxMrcd2p7_2),.clk(gclk));
	jdff dff_B_IaNmMKtE9_2(.din(w_dff_B_pxMrcd2p7_2),.dout(w_dff_B_IaNmMKtE9_2),.clk(gclk));
	jdff dff_B_XpB7DWee3_2(.din(w_dff_B_IaNmMKtE9_2),.dout(w_dff_B_XpB7DWee3_2),.clk(gclk));
	jdff dff_B_EabPG5Cm7_2(.din(w_dff_B_XpB7DWee3_2),.dout(w_dff_B_EabPG5Cm7_2),.clk(gclk));
	jdff dff_B_RXrPWNiU2_2(.din(w_dff_B_EabPG5Cm7_2),.dout(w_dff_B_RXrPWNiU2_2),.clk(gclk));
	jdff dff_B_TFV84nU96_2(.din(w_dff_B_RXrPWNiU2_2),.dout(w_dff_B_TFV84nU96_2),.clk(gclk));
	jdff dff_B_3Cg8V9mk8_2(.din(w_dff_B_TFV84nU96_2),.dout(w_dff_B_3Cg8V9mk8_2),.clk(gclk));
	jdff dff_B_aYVoHewh1_2(.din(w_dff_B_3Cg8V9mk8_2),.dout(w_dff_B_aYVoHewh1_2),.clk(gclk));
	jdff dff_B_fHJr7jH17_2(.din(w_dff_B_aYVoHewh1_2),.dout(w_dff_B_fHJr7jH17_2),.clk(gclk));
	jdff dff_B_KjBqay244_2(.din(w_dff_B_fHJr7jH17_2),.dout(w_dff_B_KjBqay244_2),.clk(gclk));
	jdff dff_B_2rsRrtsE7_2(.din(w_dff_B_KjBqay244_2),.dout(w_dff_B_2rsRrtsE7_2),.clk(gclk));
	jdff dff_B_AF7UR4pz2_2(.din(w_dff_B_2rsRrtsE7_2),.dout(w_dff_B_AF7UR4pz2_2),.clk(gclk));
	jdff dff_B_VW950xfM8_2(.din(w_dff_B_AF7UR4pz2_2),.dout(w_dff_B_VW950xfM8_2),.clk(gclk));
	jdff dff_B_RAjW8tPC7_2(.din(w_dff_B_VW950xfM8_2),.dout(w_dff_B_RAjW8tPC7_2),.clk(gclk));
	jdff dff_B_6nBwJ9zZ6_1(.din(n725),.dout(w_dff_B_6nBwJ9zZ6_1),.clk(gclk));
	jdff dff_B_TJoJ2Hpf9_2(.din(n632),.dout(w_dff_B_TJoJ2Hpf9_2),.clk(gclk));
	jdff dff_B_FOmVx54i5_2(.din(w_dff_B_TJoJ2Hpf9_2),.dout(w_dff_B_FOmVx54i5_2),.clk(gclk));
	jdff dff_B_IJ8YVhio0_2(.din(w_dff_B_FOmVx54i5_2),.dout(w_dff_B_IJ8YVhio0_2),.clk(gclk));
	jdff dff_B_PUBPL4wg6_2(.din(w_dff_B_IJ8YVhio0_2),.dout(w_dff_B_PUBPL4wg6_2),.clk(gclk));
	jdff dff_B_8IKTRe025_2(.din(w_dff_B_PUBPL4wg6_2),.dout(w_dff_B_8IKTRe025_2),.clk(gclk));
	jdff dff_B_ydpiG5zF6_2(.din(w_dff_B_8IKTRe025_2),.dout(w_dff_B_ydpiG5zF6_2),.clk(gclk));
	jdff dff_B_8UhFquDK7_2(.din(w_dff_B_ydpiG5zF6_2),.dout(w_dff_B_8UhFquDK7_2),.clk(gclk));
	jdff dff_B_4LjAfNAM1_2(.din(w_dff_B_8UhFquDK7_2),.dout(w_dff_B_4LjAfNAM1_2),.clk(gclk));
	jdff dff_B_8Q4aZSdX8_2(.din(w_dff_B_4LjAfNAM1_2),.dout(w_dff_B_8Q4aZSdX8_2),.clk(gclk));
	jdff dff_B_WucYABgL9_2(.din(w_dff_B_8Q4aZSdX8_2),.dout(w_dff_B_WucYABgL9_2),.clk(gclk));
	jdff dff_B_qSpmCzeu1_2(.din(w_dff_B_WucYABgL9_2),.dout(w_dff_B_qSpmCzeu1_2),.clk(gclk));
	jdff dff_B_LUNfMWw72_2(.din(w_dff_B_qSpmCzeu1_2),.dout(w_dff_B_LUNfMWw72_2),.clk(gclk));
	jdff dff_B_B5LDE6At9_2(.din(w_dff_B_LUNfMWw72_2),.dout(w_dff_B_B5LDE6At9_2),.clk(gclk));
	jdff dff_B_VNOsjfTr9_2(.din(w_dff_B_B5LDE6At9_2),.dout(w_dff_B_VNOsjfTr9_2),.clk(gclk));
	jdff dff_B_oJqZbqpz0_2(.din(w_dff_B_VNOsjfTr9_2),.dout(w_dff_B_oJqZbqpz0_2),.clk(gclk));
	jdff dff_B_ixdC6bzi3_2(.din(w_dff_B_oJqZbqpz0_2),.dout(w_dff_B_ixdC6bzi3_2),.clk(gclk));
	jdff dff_B_v4S9lgTS6_2(.din(w_dff_B_ixdC6bzi3_2),.dout(w_dff_B_v4S9lgTS6_2),.clk(gclk));
	jdff dff_B_l4KhkdhZ9_2(.din(w_dff_B_v4S9lgTS6_2),.dout(w_dff_B_l4KhkdhZ9_2),.clk(gclk));
	jdff dff_B_YEvaUqN93_2(.din(w_dff_B_l4KhkdhZ9_2),.dout(w_dff_B_YEvaUqN93_2),.clk(gclk));
	jdff dff_B_hc8EAVp60_2(.din(w_dff_B_YEvaUqN93_2),.dout(w_dff_B_hc8EAVp60_2),.clk(gclk));
	jdff dff_B_hg8srLWe7_2(.din(w_dff_B_hc8EAVp60_2),.dout(w_dff_B_hg8srLWe7_2),.clk(gclk));
	jdff dff_B_GTVULd038_2(.din(w_dff_B_hg8srLWe7_2),.dout(w_dff_B_GTVULd038_2),.clk(gclk));
	jdff dff_B_mvT3gYh79_1(.din(n633),.dout(w_dff_B_mvT3gYh79_1),.clk(gclk));
	jdff dff_B_RVUS5a2h9_2(.din(n547),.dout(w_dff_B_RVUS5a2h9_2),.clk(gclk));
	jdff dff_B_ggDE6zDg3_2(.din(w_dff_B_RVUS5a2h9_2),.dout(w_dff_B_ggDE6zDg3_2),.clk(gclk));
	jdff dff_B_l7bTxlJX5_2(.din(w_dff_B_ggDE6zDg3_2),.dout(w_dff_B_l7bTxlJX5_2),.clk(gclk));
	jdff dff_B_4SLqWwqp8_2(.din(w_dff_B_l7bTxlJX5_2),.dout(w_dff_B_4SLqWwqp8_2),.clk(gclk));
	jdff dff_B_Ovj3rpTv1_2(.din(w_dff_B_4SLqWwqp8_2),.dout(w_dff_B_Ovj3rpTv1_2),.clk(gclk));
	jdff dff_B_xaXNsIvP0_2(.din(w_dff_B_Ovj3rpTv1_2),.dout(w_dff_B_xaXNsIvP0_2),.clk(gclk));
	jdff dff_B_cbr649zh8_2(.din(w_dff_B_xaXNsIvP0_2),.dout(w_dff_B_cbr649zh8_2),.clk(gclk));
	jdff dff_B_IzZig3L51_2(.din(w_dff_B_cbr649zh8_2),.dout(w_dff_B_IzZig3L51_2),.clk(gclk));
	jdff dff_B_cLwDYBZt7_2(.din(w_dff_B_IzZig3L51_2),.dout(w_dff_B_cLwDYBZt7_2),.clk(gclk));
	jdff dff_B_aFHeId8D9_2(.din(w_dff_B_cLwDYBZt7_2),.dout(w_dff_B_aFHeId8D9_2),.clk(gclk));
	jdff dff_B_k8gJGjYO9_2(.din(w_dff_B_aFHeId8D9_2),.dout(w_dff_B_k8gJGjYO9_2),.clk(gclk));
	jdff dff_B_dFzZABtA2_2(.din(w_dff_B_k8gJGjYO9_2),.dout(w_dff_B_dFzZABtA2_2),.clk(gclk));
	jdff dff_B_di7Gth1s0_2(.din(w_dff_B_dFzZABtA2_2),.dout(w_dff_B_di7Gth1s0_2),.clk(gclk));
	jdff dff_B_qHK1YvLl7_2(.din(w_dff_B_di7Gth1s0_2),.dout(w_dff_B_qHK1YvLl7_2),.clk(gclk));
	jdff dff_B_t9gbcdDy4_2(.din(w_dff_B_qHK1YvLl7_2),.dout(w_dff_B_t9gbcdDy4_2),.clk(gclk));
	jdff dff_B_gVa2kFoR4_2(.din(w_dff_B_t9gbcdDy4_2),.dout(w_dff_B_gVa2kFoR4_2),.clk(gclk));
	jdff dff_B_Vzh9OvP67_2(.din(w_dff_B_gVa2kFoR4_2),.dout(w_dff_B_Vzh9OvP67_2),.clk(gclk));
	jdff dff_B_a9wQwVAx2_2(.din(w_dff_B_Vzh9OvP67_2),.dout(w_dff_B_a9wQwVAx2_2),.clk(gclk));
	jdff dff_B_5UxDSrDo0_2(.din(w_dff_B_a9wQwVAx2_2),.dout(w_dff_B_5UxDSrDo0_2),.clk(gclk));
	jdff dff_B_U7tVD6sA5_2(.din(w_dff_B_5UxDSrDo0_2),.dout(w_dff_B_U7tVD6sA5_2),.clk(gclk));
	jdff dff_B_v8QRd6LZ4_1(.din(n548),.dout(w_dff_B_v8QRd6LZ4_1),.clk(gclk));
	jdff dff_B_8w2BWKKy4_2(.din(n469),.dout(w_dff_B_8w2BWKKy4_2),.clk(gclk));
	jdff dff_B_X7BbLtuU9_2(.din(w_dff_B_8w2BWKKy4_2),.dout(w_dff_B_X7BbLtuU9_2),.clk(gclk));
	jdff dff_B_x3q2Bcwx9_2(.din(w_dff_B_X7BbLtuU9_2),.dout(w_dff_B_x3q2Bcwx9_2),.clk(gclk));
	jdff dff_B_XWG9cLbQ4_2(.din(w_dff_B_x3q2Bcwx9_2),.dout(w_dff_B_XWG9cLbQ4_2),.clk(gclk));
	jdff dff_B_2jqGrJnV1_2(.din(w_dff_B_XWG9cLbQ4_2),.dout(w_dff_B_2jqGrJnV1_2),.clk(gclk));
	jdff dff_B_sz7LAJru1_2(.din(w_dff_B_2jqGrJnV1_2),.dout(w_dff_B_sz7LAJru1_2),.clk(gclk));
	jdff dff_B_WFwaxirL5_2(.din(w_dff_B_sz7LAJru1_2),.dout(w_dff_B_WFwaxirL5_2),.clk(gclk));
	jdff dff_B_iS8NsnM98_2(.din(w_dff_B_WFwaxirL5_2),.dout(w_dff_B_iS8NsnM98_2),.clk(gclk));
	jdff dff_B_tbhI4mFC6_2(.din(w_dff_B_iS8NsnM98_2),.dout(w_dff_B_tbhI4mFC6_2),.clk(gclk));
	jdff dff_B_YrDirVu17_2(.din(w_dff_B_tbhI4mFC6_2),.dout(w_dff_B_YrDirVu17_2),.clk(gclk));
	jdff dff_B_BBG1u3ts7_2(.din(w_dff_B_YrDirVu17_2),.dout(w_dff_B_BBG1u3ts7_2),.clk(gclk));
	jdff dff_B_Gd0BBvtD0_2(.din(w_dff_B_BBG1u3ts7_2),.dout(w_dff_B_Gd0BBvtD0_2),.clk(gclk));
	jdff dff_B_f7h8Dusw2_2(.din(w_dff_B_Gd0BBvtD0_2),.dout(w_dff_B_f7h8Dusw2_2),.clk(gclk));
	jdff dff_B_klHxXJKr7_2(.din(w_dff_B_f7h8Dusw2_2),.dout(w_dff_B_klHxXJKr7_2),.clk(gclk));
	jdff dff_B_9XVQ6UH09_2(.din(w_dff_B_klHxXJKr7_2),.dout(w_dff_B_9XVQ6UH09_2),.clk(gclk));
	jdff dff_B_XSJYdEVn0_2(.din(w_dff_B_9XVQ6UH09_2),.dout(w_dff_B_XSJYdEVn0_2),.clk(gclk));
	jdff dff_B_D0wlWiL92_2(.din(w_dff_B_XSJYdEVn0_2),.dout(w_dff_B_D0wlWiL92_2),.clk(gclk));
	jdff dff_B_mMtDY7Ft3_2(.din(w_dff_B_D0wlWiL92_2),.dout(w_dff_B_mMtDY7Ft3_2),.clk(gclk));
	jdff dff_B_zBQXm9a34_1(.din(n470),.dout(w_dff_B_zBQXm9a34_1),.clk(gclk));
	jdff dff_B_1vcisxuE7_2(.din(n398),.dout(w_dff_B_1vcisxuE7_2),.clk(gclk));
	jdff dff_B_RVCFi1c31_2(.din(w_dff_B_1vcisxuE7_2),.dout(w_dff_B_RVCFi1c31_2),.clk(gclk));
	jdff dff_B_ExsH5ryU0_2(.din(w_dff_B_RVCFi1c31_2),.dout(w_dff_B_ExsH5ryU0_2),.clk(gclk));
	jdff dff_B_XdZN0oQW5_2(.din(w_dff_B_ExsH5ryU0_2),.dout(w_dff_B_XdZN0oQW5_2),.clk(gclk));
	jdff dff_B_IQQ7YdGG9_2(.din(w_dff_B_XdZN0oQW5_2),.dout(w_dff_B_IQQ7YdGG9_2),.clk(gclk));
	jdff dff_B_B36eK0DP3_2(.din(w_dff_B_IQQ7YdGG9_2),.dout(w_dff_B_B36eK0DP3_2),.clk(gclk));
	jdff dff_B_FMjixvov4_2(.din(w_dff_B_B36eK0DP3_2),.dout(w_dff_B_FMjixvov4_2),.clk(gclk));
	jdff dff_B_6CP1r0ny1_2(.din(w_dff_B_FMjixvov4_2),.dout(w_dff_B_6CP1r0ny1_2),.clk(gclk));
	jdff dff_B_KnvoEbWM2_2(.din(w_dff_B_6CP1r0ny1_2),.dout(w_dff_B_KnvoEbWM2_2),.clk(gclk));
	jdff dff_B_GafvfmSv4_2(.din(w_dff_B_KnvoEbWM2_2),.dout(w_dff_B_GafvfmSv4_2),.clk(gclk));
	jdff dff_B_MtNYffRt7_2(.din(w_dff_B_GafvfmSv4_2),.dout(w_dff_B_MtNYffRt7_2),.clk(gclk));
	jdff dff_B_fd4wgxW34_2(.din(w_dff_B_MtNYffRt7_2),.dout(w_dff_B_fd4wgxW34_2),.clk(gclk));
	jdff dff_B_PE2x74zx9_2(.din(w_dff_B_fd4wgxW34_2),.dout(w_dff_B_PE2x74zx9_2),.clk(gclk));
	jdff dff_B_4r0V9rLA0_2(.din(w_dff_B_PE2x74zx9_2),.dout(w_dff_B_4r0V9rLA0_2),.clk(gclk));
	jdff dff_B_fHZXDJi48_2(.din(w_dff_B_4r0V9rLA0_2),.dout(w_dff_B_fHZXDJi48_2),.clk(gclk));
	jdff dff_B_gd3sCwu39_2(.din(w_dff_B_fHZXDJi48_2),.dout(w_dff_B_gd3sCwu39_2),.clk(gclk));
	jdff dff_B_DwbZPHca6_2(.din(n401),.dout(w_dff_B_DwbZPHca6_2),.clk(gclk));
	jdff dff_B_8LSZcutg8_2(.din(w_dff_B_DwbZPHca6_2),.dout(w_dff_B_8LSZcutg8_2),.clk(gclk));
	jdff dff_B_1aTwimwz5_2(.din(w_dff_B_8LSZcutg8_2),.dout(w_dff_B_1aTwimwz5_2),.clk(gclk));
	jdff dff_B_YDTgA7rp3_1(.din(n399),.dout(w_dff_B_YDTgA7rp3_1),.clk(gclk));
	jdff dff_B_y7DxDGZo8_2(.din(n335),.dout(w_dff_B_y7DxDGZo8_2),.clk(gclk));
	jdff dff_B_5mrxDeXX1_2(.din(w_dff_B_y7DxDGZo8_2),.dout(w_dff_B_5mrxDeXX1_2),.clk(gclk));
	jdff dff_B_Fl8KEnUB2_2(.din(w_dff_B_5mrxDeXX1_2),.dout(w_dff_B_Fl8KEnUB2_2),.clk(gclk));
	jdff dff_B_KofwOBxw2_2(.din(w_dff_B_Fl8KEnUB2_2),.dout(w_dff_B_KofwOBxw2_2),.clk(gclk));
	jdff dff_B_Nv0tesUh2_2(.din(w_dff_B_KofwOBxw2_2),.dout(w_dff_B_Nv0tesUh2_2),.clk(gclk));
	jdff dff_B_7p5YZYKu8_2(.din(w_dff_B_Nv0tesUh2_2),.dout(w_dff_B_7p5YZYKu8_2),.clk(gclk));
	jdff dff_B_rsFCvRc05_2(.din(w_dff_B_7p5YZYKu8_2),.dout(w_dff_B_rsFCvRc05_2),.clk(gclk));
	jdff dff_B_E0bbs0sO1_2(.din(w_dff_B_rsFCvRc05_2),.dout(w_dff_B_E0bbs0sO1_2),.clk(gclk));
	jdff dff_B_lcKFYHoU3_2(.din(w_dff_B_E0bbs0sO1_2),.dout(w_dff_B_lcKFYHoU3_2),.clk(gclk));
	jdff dff_B_FEx3ty9d0_2(.din(w_dff_B_lcKFYHoU3_2),.dout(w_dff_B_FEx3ty9d0_2),.clk(gclk));
	jdff dff_B_bnx2wppo4_2(.din(w_dff_B_FEx3ty9d0_2),.dout(w_dff_B_bnx2wppo4_2),.clk(gclk));
	jdff dff_B_TjKIPwAU4_1(.din(n336),.dout(w_dff_B_TjKIPwAU4_1),.clk(gclk));
	jdff dff_B_FrDCNQQy6_2(.din(n279),.dout(w_dff_B_FrDCNQQy6_2),.clk(gclk));
	jdff dff_B_vyUOjMeo3_2(.din(w_dff_B_FrDCNQQy6_2),.dout(w_dff_B_vyUOjMeo3_2),.clk(gclk));
	jdff dff_B_KsKCkddE8_2(.din(w_dff_B_vyUOjMeo3_2),.dout(w_dff_B_KsKCkddE8_2),.clk(gclk));
	jdff dff_B_CSVUpzss6_2(.din(w_dff_B_KsKCkddE8_2),.dout(w_dff_B_CSVUpzss6_2),.clk(gclk));
	jdff dff_B_FtQPF6pV8_2(.din(w_dff_B_CSVUpzss6_2),.dout(w_dff_B_FtQPF6pV8_2),.clk(gclk));
	jdff dff_B_zBpkpyB48_2(.din(w_dff_B_FtQPF6pV8_2),.dout(w_dff_B_zBpkpyB48_2),.clk(gclk));
	jdff dff_B_tMW2Z0Vc1_2(.din(w_dff_B_zBpkpyB48_2),.dout(w_dff_B_tMW2Z0Vc1_2),.clk(gclk));
	jdff dff_B_jPvqwdoK4_2(.din(w_dff_B_tMW2Z0Vc1_2),.dout(w_dff_B_jPvqwdoK4_2),.clk(gclk));
	jdff dff_B_xv1nQ7vz8_2(.din(w_dff_B_jPvqwdoK4_2),.dout(w_dff_B_xv1nQ7vz8_2),.clk(gclk));
	jdff dff_B_TMXlGXGE2_1(.din(n280),.dout(w_dff_B_TMXlGXGE2_1),.clk(gclk));
	jdff dff_B_48mobnWy5_2(.din(n230),.dout(w_dff_B_48mobnWy5_2),.clk(gclk));
	jdff dff_B_Q1H5wwwU9_2(.din(w_dff_B_48mobnWy5_2),.dout(w_dff_B_Q1H5wwwU9_2),.clk(gclk));
	jdff dff_B_nGFwCgmu1_2(.din(w_dff_B_Q1H5wwwU9_2),.dout(w_dff_B_nGFwCgmu1_2),.clk(gclk));
	jdff dff_B_DMvDq34q2_2(.din(w_dff_B_nGFwCgmu1_2),.dout(w_dff_B_DMvDq34q2_2),.clk(gclk));
	jdff dff_B_LuqvSgt21_2(.din(w_dff_B_DMvDq34q2_2),.dout(w_dff_B_LuqvSgt21_2),.clk(gclk));
	jdff dff_B_BhTaxGEE2_2(.din(w_dff_B_LuqvSgt21_2),.dout(w_dff_B_BhTaxGEE2_2),.clk(gclk));
	jdff dff_B_hzjeHgL23_2(.din(w_dff_B_BhTaxGEE2_2),.dout(w_dff_B_hzjeHgL23_2),.clk(gclk));
	jdff dff_B_H8Nf2bxb9_1(.din(n231),.dout(w_dff_B_H8Nf2bxb9_1),.clk(gclk));
	jdff dff_B_8BOK5r7f5_2(.din(n188),.dout(w_dff_B_8BOK5r7f5_2),.clk(gclk));
	jdff dff_B_CxMuwOBI4_2(.din(w_dff_B_8BOK5r7f5_2),.dout(w_dff_B_CxMuwOBI4_2),.clk(gclk));
	jdff dff_B_EqHqyi9Y4_2(.din(w_dff_B_CxMuwOBI4_2),.dout(w_dff_B_EqHqyi9Y4_2),.clk(gclk));
	jdff dff_B_ma8H6lte4_2(.din(w_dff_B_EqHqyi9Y4_2),.dout(w_dff_B_ma8H6lte4_2),.clk(gclk));
	jdff dff_B_AxwWbGXe2_2(.din(w_dff_B_ma8H6lte4_2),.dout(w_dff_B_AxwWbGXe2_2),.clk(gclk));
	jdff dff_B_SM2C5eTN2_2(.din(n154),.dout(w_dff_B_SM2C5eTN2_2),.clk(gclk));
	jdff dff_B_B23Uh0Jm4_2(.din(w_dff_B_SM2C5eTN2_2),.dout(w_dff_B_B23Uh0Jm4_2),.clk(gclk));
	jdff dff_B_IQchRE107_2(.din(w_dff_B_B23Uh0Jm4_2),.dout(w_dff_B_IQchRE107_2),.clk(gclk));
	jdff dff_B_RtYdSlrb2_0(.din(n159),.dout(w_dff_B_RtYdSlrb2_0),.clk(gclk));
	jdff dff_B_7heOTNru1_0(.din(w_dff_B_RtYdSlrb2_0),.dout(w_dff_B_7heOTNru1_0),.clk(gclk));
	jdff dff_A_A02n2DW34_0(.dout(w_n123_0[0]),.din(w_dff_A_A02n2DW34_0),.clk(gclk));
	jdff dff_A_kkCyMRDe5_0(.dout(w_dff_A_A02n2DW34_0),.din(w_dff_A_kkCyMRDe5_0),.clk(gclk));
	jdff dff_A_D6DhIAUh2_0(.dout(w_n122_0[0]),.din(w_dff_A_D6DhIAUh2_0),.clk(gclk));
	jdff dff_A_o1vhWlM35_0(.dout(w_dff_A_D6DhIAUh2_0),.din(w_dff_A_o1vhWlM35_0),.clk(gclk));
	jdff dff_B_pxiAqJRP4_2(.din(n1306),.dout(w_dff_B_pxiAqJRP4_2),.clk(gclk));
	jdff dff_B_fmTukOSK5_1(.din(n1304),.dout(w_dff_B_fmTukOSK5_1),.clk(gclk));
	jdff dff_B_Ze2a0qMu3_2(.din(n1217),.dout(w_dff_B_Ze2a0qMu3_2),.clk(gclk));
	jdff dff_B_YNHysRsW8_2(.din(w_dff_B_Ze2a0qMu3_2),.dout(w_dff_B_YNHysRsW8_2),.clk(gclk));
	jdff dff_B_vhuHWw3O6_2(.din(w_dff_B_YNHysRsW8_2),.dout(w_dff_B_vhuHWw3O6_2),.clk(gclk));
	jdff dff_B_jOEJPwI61_2(.din(w_dff_B_vhuHWw3O6_2),.dout(w_dff_B_jOEJPwI61_2),.clk(gclk));
	jdff dff_B_KB4AWD940_2(.din(w_dff_B_jOEJPwI61_2),.dout(w_dff_B_KB4AWD940_2),.clk(gclk));
	jdff dff_B_qf5Yo19P0_2(.din(w_dff_B_KB4AWD940_2),.dout(w_dff_B_qf5Yo19P0_2),.clk(gclk));
	jdff dff_B_INZgAJQT9_2(.din(w_dff_B_qf5Yo19P0_2),.dout(w_dff_B_INZgAJQT9_2),.clk(gclk));
	jdff dff_B_2MB8g3V94_2(.din(w_dff_B_INZgAJQT9_2),.dout(w_dff_B_2MB8g3V94_2),.clk(gclk));
	jdff dff_B_KiemjYa75_2(.din(w_dff_B_2MB8g3V94_2),.dout(w_dff_B_KiemjYa75_2),.clk(gclk));
	jdff dff_B_m531pyuN3_2(.din(w_dff_B_KiemjYa75_2),.dout(w_dff_B_m531pyuN3_2),.clk(gclk));
	jdff dff_B_Nmk57WAB8_2(.din(w_dff_B_m531pyuN3_2),.dout(w_dff_B_Nmk57WAB8_2),.clk(gclk));
	jdff dff_B_sBmusA4K8_2(.din(w_dff_B_Nmk57WAB8_2),.dout(w_dff_B_sBmusA4K8_2),.clk(gclk));
	jdff dff_B_GA5KIA3m8_2(.din(w_dff_B_sBmusA4K8_2),.dout(w_dff_B_GA5KIA3m8_2),.clk(gclk));
	jdff dff_B_xwOSLHyZ4_2(.din(w_dff_B_GA5KIA3m8_2),.dout(w_dff_B_xwOSLHyZ4_2),.clk(gclk));
	jdff dff_B_hU9xqo8f2_2(.din(w_dff_B_xwOSLHyZ4_2),.dout(w_dff_B_hU9xqo8f2_2),.clk(gclk));
	jdff dff_B_mGMsgOJa8_2(.din(w_dff_B_hU9xqo8f2_2),.dout(w_dff_B_mGMsgOJa8_2),.clk(gclk));
	jdff dff_B_O3gYNr327_2(.din(w_dff_B_mGMsgOJa8_2),.dout(w_dff_B_O3gYNr327_2),.clk(gclk));
	jdff dff_B_cNU9WGg78_2(.din(w_dff_B_O3gYNr327_2),.dout(w_dff_B_cNU9WGg78_2),.clk(gclk));
	jdff dff_B_4pN8YaBQ7_2(.din(w_dff_B_cNU9WGg78_2),.dout(w_dff_B_4pN8YaBQ7_2),.clk(gclk));
	jdff dff_B_AuWUyTAJ2_2(.din(w_dff_B_4pN8YaBQ7_2),.dout(w_dff_B_AuWUyTAJ2_2),.clk(gclk));
	jdff dff_B_WFN8QgVC2_2(.din(w_dff_B_AuWUyTAJ2_2),.dout(w_dff_B_WFN8QgVC2_2),.clk(gclk));
	jdff dff_B_siZdu26O8_2(.din(w_dff_B_WFN8QgVC2_2),.dout(w_dff_B_siZdu26O8_2),.clk(gclk));
	jdff dff_B_9GhRiICd4_2(.din(w_dff_B_siZdu26O8_2),.dout(w_dff_B_9GhRiICd4_2),.clk(gclk));
	jdff dff_B_zobSXAoj9_2(.din(w_dff_B_9GhRiICd4_2),.dout(w_dff_B_zobSXAoj9_2),.clk(gclk));
	jdff dff_B_cDE7uDpV1_2(.din(w_dff_B_zobSXAoj9_2),.dout(w_dff_B_cDE7uDpV1_2),.clk(gclk));
	jdff dff_B_en5LGY3f9_2(.din(w_dff_B_cDE7uDpV1_2),.dout(w_dff_B_en5LGY3f9_2),.clk(gclk));
	jdff dff_B_urn32Fvt0_2(.din(w_dff_B_en5LGY3f9_2),.dout(w_dff_B_urn32Fvt0_2),.clk(gclk));
	jdff dff_B_HAHz5OiS7_2(.din(w_dff_B_urn32Fvt0_2),.dout(w_dff_B_HAHz5OiS7_2),.clk(gclk));
	jdff dff_B_9WiIpf7b4_2(.din(w_dff_B_HAHz5OiS7_2),.dout(w_dff_B_9WiIpf7b4_2),.clk(gclk));
	jdff dff_B_N6wxh4pV5_2(.din(w_dff_B_9WiIpf7b4_2),.dout(w_dff_B_N6wxh4pV5_2),.clk(gclk));
	jdff dff_B_CnkhAJF62_2(.din(w_dff_B_N6wxh4pV5_2),.dout(w_dff_B_CnkhAJF62_2),.clk(gclk));
	jdff dff_B_RPWS1Gxo0_2(.din(w_dff_B_CnkhAJF62_2),.dout(w_dff_B_RPWS1Gxo0_2),.clk(gclk));
	jdff dff_B_Hej4yq6j7_2(.din(w_dff_B_RPWS1Gxo0_2),.dout(w_dff_B_Hej4yq6j7_2),.clk(gclk));
	jdff dff_B_ovoLQTwy0_2(.din(w_dff_B_Hej4yq6j7_2),.dout(w_dff_B_ovoLQTwy0_2),.clk(gclk));
	jdff dff_B_yr9X1Uji1_1(.din(n1218),.dout(w_dff_B_yr9X1Uji1_1),.clk(gclk));
	jdff dff_B_6Ig0Wrib6_2(.din(n1126),.dout(w_dff_B_6Ig0Wrib6_2),.clk(gclk));
	jdff dff_B_sBbrPwaD0_2(.din(w_dff_B_6Ig0Wrib6_2),.dout(w_dff_B_sBbrPwaD0_2),.clk(gclk));
	jdff dff_B_s9hlSRkh7_2(.din(w_dff_B_sBbrPwaD0_2),.dout(w_dff_B_s9hlSRkh7_2),.clk(gclk));
	jdff dff_B_yIeyAk5M5_2(.din(w_dff_B_s9hlSRkh7_2),.dout(w_dff_B_yIeyAk5M5_2),.clk(gclk));
	jdff dff_B_9WotExv62_2(.din(w_dff_B_yIeyAk5M5_2),.dout(w_dff_B_9WotExv62_2),.clk(gclk));
	jdff dff_B_gMlNety95_2(.din(w_dff_B_9WotExv62_2),.dout(w_dff_B_gMlNety95_2),.clk(gclk));
	jdff dff_B_rxj5pdJ56_2(.din(w_dff_B_gMlNety95_2),.dout(w_dff_B_rxj5pdJ56_2),.clk(gclk));
	jdff dff_B_ylUgR8Pk1_2(.din(w_dff_B_rxj5pdJ56_2),.dout(w_dff_B_ylUgR8Pk1_2),.clk(gclk));
	jdff dff_B_Qtva6Esw2_2(.din(w_dff_B_ylUgR8Pk1_2),.dout(w_dff_B_Qtva6Esw2_2),.clk(gclk));
	jdff dff_B_49h92b0f8_2(.din(w_dff_B_Qtva6Esw2_2),.dout(w_dff_B_49h92b0f8_2),.clk(gclk));
	jdff dff_B_sCzqxtOy2_2(.din(w_dff_B_49h92b0f8_2),.dout(w_dff_B_sCzqxtOy2_2),.clk(gclk));
	jdff dff_B_TgGzpvF81_2(.din(w_dff_B_sCzqxtOy2_2),.dout(w_dff_B_TgGzpvF81_2),.clk(gclk));
	jdff dff_B_UKZKDgEx1_2(.din(w_dff_B_TgGzpvF81_2),.dout(w_dff_B_UKZKDgEx1_2),.clk(gclk));
	jdff dff_B_RUCec0kw1_2(.din(w_dff_B_UKZKDgEx1_2),.dout(w_dff_B_RUCec0kw1_2),.clk(gclk));
	jdff dff_B_XuJUKu6A2_2(.din(w_dff_B_RUCec0kw1_2),.dout(w_dff_B_XuJUKu6A2_2),.clk(gclk));
	jdff dff_B_5heccAfs4_2(.din(w_dff_B_XuJUKu6A2_2),.dout(w_dff_B_5heccAfs4_2),.clk(gclk));
	jdff dff_B_HwNprvhk8_2(.din(w_dff_B_5heccAfs4_2),.dout(w_dff_B_HwNprvhk8_2),.clk(gclk));
	jdff dff_B_kfq9iLjj8_2(.din(w_dff_B_HwNprvhk8_2),.dout(w_dff_B_kfq9iLjj8_2),.clk(gclk));
	jdff dff_B_gHajJhX94_2(.din(w_dff_B_kfq9iLjj8_2),.dout(w_dff_B_gHajJhX94_2),.clk(gclk));
	jdff dff_B_uXsq1X8p9_2(.din(w_dff_B_gHajJhX94_2),.dout(w_dff_B_uXsq1X8p9_2),.clk(gclk));
	jdff dff_B_veHxe9MD8_2(.din(w_dff_B_uXsq1X8p9_2),.dout(w_dff_B_veHxe9MD8_2),.clk(gclk));
	jdff dff_B_ExQjT2xe0_2(.din(w_dff_B_veHxe9MD8_2),.dout(w_dff_B_ExQjT2xe0_2),.clk(gclk));
	jdff dff_B_KF8C1XD12_2(.din(w_dff_B_ExQjT2xe0_2),.dout(w_dff_B_KF8C1XD12_2),.clk(gclk));
	jdff dff_B_CDI0nxj59_2(.din(w_dff_B_KF8C1XD12_2),.dout(w_dff_B_CDI0nxj59_2),.clk(gclk));
	jdff dff_B_KDikc2b82_2(.din(w_dff_B_CDI0nxj59_2),.dout(w_dff_B_KDikc2b82_2),.clk(gclk));
	jdff dff_B_bTUYfIJx8_2(.din(w_dff_B_KDikc2b82_2),.dout(w_dff_B_bTUYfIJx8_2),.clk(gclk));
	jdff dff_B_NA27Ky2t1_2(.din(w_dff_B_bTUYfIJx8_2),.dout(w_dff_B_NA27Ky2t1_2),.clk(gclk));
	jdff dff_B_qu7Z9csu7_2(.din(w_dff_B_NA27Ky2t1_2),.dout(w_dff_B_qu7Z9csu7_2),.clk(gclk));
	jdff dff_B_2ruYm7nD8_2(.din(w_dff_B_qu7Z9csu7_2),.dout(w_dff_B_2ruYm7nD8_2),.clk(gclk));
	jdff dff_B_hFHKLx7N3_2(.din(w_dff_B_2ruYm7nD8_2),.dout(w_dff_B_hFHKLx7N3_2),.clk(gclk));
	jdff dff_B_fZLq7QUg3_1(.din(n1127),.dout(w_dff_B_fZLq7QUg3_1),.clk(gclk));
	jdff dff_B_EJMh1QQl6_2(.din(n1028),.dout(w_dff_B_EJMh1QQl6_2),.clk(gclk));
	jdff dff_B_BWgqeZbH8_2(.din(w_dff_B_EJMh1QQl6_2),.dout(w_dff_B_BWgqeZbH8_2),.clk(gclk));
	jdff dff_B_bieWKeHu9_2(.din(w_dff_B_BWgqeZbH8_2),.dout(w_dff_B_bieWKeHu9_2),.clk(gclk));
	jdff dff_B_CkQURvXS1_2(.din(w_dff_B_bieWKeHu9_2),.dout(w_dff_B_CkQURvXS1_2),.clk(gclk));
	jdff dff_B_ePCTChUN6_2(.din(w_dff_B_CkQURvXS1_2),.dout(w_dff_B_ePCTChUN6_2),.clk(gclk));
	jdff dff_B_810kvt9M8_2(.din(w_dff_B_ePCTChUN6_2),.dout(w_dff_B_810kvt9M8_2),.clk(gclk));
	jdff dff_B_1uf4QUqx2_2(.din(w_dff_B_810kvt9M8_2),.dout(w_dff_B_1uf4QUqx2_2),.clk(gclk));
	jdff dff_B_gGGvKriD3_2(.din(w_dff_B_1uf4QUqx2_2),.dout(w_dff_B_gGGvKriD3_2),.clk(gclk));
	jdff dff_B_KN7D9rK21_2(.din(w_dff_B_gGGvKriD3_2),.dout(w_dff_B_KN7D9rK21_2),.clk(gclk));
	jdff dff_B_GctTT3680_2(.din(w_dff_B_KN7D9rK21_2),.dout(w_dff_B_GctTT3680_2),.clk(gclk));
	jdff dff_B_DZt5sDHW2_2(.din(w_dff_B_GctTT3680_2),.dout(w_dff_B_DZt5sDHW2_2),.clk(gclk));
	jdff dff_B_SBdJTp2B6_2(.din(w_dff_B_DZt5sDHW2_2),.dout(w_dff_B_SBdJTp2B6_2),.clk(gclk));
	jdff dff_B_m2tIKxb96_2(.din(w_dff_B_SBdJTp2B6_2),.dout(w_dff_B_m2tIKxb96_2),.clk(gclk));
	jdff dff_B_YIOpxhuX9_2(.din(w_dff_B_m2tIKxb96_2),.dout(w_dff_B_YIOpxhuX9_2),.clk(gclk));
	jdff dff_B_MbeO3Ngk5_2(.din(w_dff_B_YIOpxhuX9_2),.dout(w_dff_B_MbeO3Ngk5_2),.clk(gclk));
	jdff dff_B_muqdDLpo7_2(.din(w_dff_B_MbeO3Ngk5_2),.dout(w_dff_B_muqdDLpo7_2),.clk(gclk));
	jdff dff_B_N6rH1bXL3_2(.din(w_dff_B_muqdDLpo7_2),.dout(w_dff_B_N6rH1bXL3_2),.clk(gclk));
	jdff dff_B_vCumNGsD2_2(.din(w_dff_B_N6rH1bXL3_2),.dout(w_dff_B_vCumNGsD2_2),.clk(gclk));
	jdff dff_B_JidzGYRu2_2(.din(w_dff_B_vCumNGsD2_2),.dout(w_dff_B_JidzGYRu2_2),.clk(gclk));
	jdff dff_B_dwxKcmGg2_2(.din(w_dff_B_JidzGYRu2_2),.dout(w_dff_B_dwxKcmGg2_2),.clk(gclk));
	jdff dff_B_ahuWJ8uT9_2(.din(w_dff_B_dwxKcmGg2_2),.dout(w_dff_B_ahuWJ8uT9_2),.clk(gclk));
	jdff dff_B_WfFv4OxZ1_2(.din(w_dff_B_ahuWJ8uT9_2),.dout(w_dff_B_WfFv4OxZ1_2),.clk(gclk));
	jdff dff_B_R0Cp8kF14_2(.din(w_dff_B_WfFv4OxZ1_2),.dout(w_dff_B_R0Cp8kF14_2),.clk(gclk));
	jdff dff_B_PrHpp7u75_2(.din(w_dff_B_R0Cp8kF14_2),.dout(w_dff_B_PrHpp7u75_2),.clk(gclk));
	jdff dff_B_cMdFCd0j0_2(.din(w_dff_B_PrHpp7u75_2),.dout(w_dff_B_cMdFCd0j0_2),.clk(gclk));
	jdff dff_B_xdppXo9f3_2(.din(w_dff_B_cMdFCd0j0_2),.dout(w_dff_B_xdppXo9f3_2),.clk(gclk));
	jdff dff_B_jSQvbZOs1_2(.din(w_dff_B_xdppXo9f3_2),.dout(w_dff_B_jSQvbZOs1_2),.clk(gclk));
	jdff dff_B_kvmSRX9U9_2(.din(w_dff_B_jSQvbZOs1_2),.dout(w_dff_B_kvmSRX9U9_2),.clk(gclk));
	jdff dff_B_Vxbm8uDo5_1(.din(n1029),.dout(w_dff_B_Vxbm8uDo5_1),.clk(gclk));
	jdff dff_B_p4ZB1WcP1_2(.din(n929),.dout(w_dff_B_p4ZB1WcP1_2),.clk(gclk));
	jdff dff_B_DlRZdn8u4_2(.din(w_dff_B_p4ZB1WcP1_2),.dout(w_dff_B_DlRZdn8u4_2),.clk(gclk));
	jdff dff_B_N1aHqhFc7_2(.din(w_dff_B_DlRZdn8u4_2),.dout(w_dff_B_N1aHqhFc7_2),.clk(gclk));
	jdff dff_B_JJ9pVtSQ3_2(.din(w_dff_B_N1aHqhFc7_2),.dout(w_dff_B_JJ9pVtSQ3_2),.clk(gclk));
	jdff dff_B_hfbEGqzB6_2(.din(w_dff_B_JJ9pVtSQ3_2),.dout(w_dff_B_hfbEGqzB6_2),.clk(gclk));
	jdff dff_B_zmdeI1RR2_2(.din(w_dff_B_hfbEGqzB6_2),.dout(w_dff_B_zmdeI1RR2_2),.clk(gclk));
	jdff dff_B_OJm5394n6_2(.din(w_dff_B_zmdeI1RR2_2),.dout(w_dff_B_OJm5394n6_2),.clk(gclk));
	jdff dff_B_rpcW0TBT6_2(.din(w_dff_B_OJm5394n6_2),.dout(w_dff_B_rpcW0TBT6_2),.clk(gclk));
	jdff dff_B_KJeVeG0Y7_2(.din(w_dff_B_rpcW0TBT6_2),.dout(w_dff_B_KJeVeG0Y7_2),.clk(gclk));
	jdff dff_B_EVCM8vJY2_2(.din(w_dff_B_KJeVeG0Y7_2),.dout(w_dff_B_EVCM8vJY2_2),.clk(gclk));
	jdff dff_B_LvW401D86_2(.din(w_dff_B_EVCM8vJY2_2),.dout(w_dff_B_LvW401D86_2),.clk(gclk));
	jdff dff_B_nGLDQ6Bm0_2(.din(w_dff_B_LvW401D86_2),.dout(w_dff_B_nGLDQ6Bm0_2),.clk(gclk));
	jdff dff_B_gTY9Q1OR2_2(.din(w_dff_B_nGLDQ6Bm0_2),.dout(w_dff_B_gTY9Q1OR2_2),.clk(gclk));
	jdff dff_B_sVh1yYi77_2(.din(w_dff_B_gTY9Q1OR2_2),.dout(w_dff_B_sVh1yYi77_2),.clk(gclk));
	jdff dff_B_X7kFy1Ak6_2(.din(w_dff_B_sVh1yYi77_2),.dout(w_dff_B_X7kFy1Ak6_2),.clk(gclk));
	jdff dff_B_sTlOQjPh4_2(.din(w_dff_B_X7kFy1Ak6_2),.dout(w_dff_B_sTlOQjPh4_2),.clk(gclk));
	jdff dff_B_s4HKLGQL7_2(.din(w_dff_B_sTlOQjPh4_2),.dout(w_dff_B_s4HKLGQL7_2),.clk(gclk));
	jdff dff_B_wP4T2oEx5_2(.din(w_dff_B_s4HKLGQL7_2),.dout(w_dff_B_wP4T2oEx5_2),.clk(gclk));
	jdff dff_B_FKrWEXpt5_2(.din(w_dff_B_wP4T2oEx5_2),.dout(w_dff_B_FKrWEXpt5_2),.clk(gclk));
	jdff dff_B_rB8BmRK09_2(.din(w_dff_B_FKrWEXpt5_2),.dout(w_dff_B_rB8BmRK09_2),.clk(gclk));
	jdff dff_B_upOfiIN43_2(.din(w_dff_B_rB8BmRK09_2),.dout(w_dff_B_upOfiIN43_2),.clk(gclk));
	jdff dff_B_X8IGTZ6y3_2(.din(w_dff_B_upOfiIN43_2),.dout(w_dff_B_X8IGTZ6y3_2),.clk(gclk));
	jdff dff_B_IF5z1V8o8_2(.din(w_dff_B_X8IGTZ6y3_2),.dout(w_dff_B_IF5z1V8o8_2),.clk(gclk));
	jdff dff_B_Q1hnPCL74_2(.din(w_dff_B_IF5z1V8o8_2),.dout(w_dff_B_Q1hnPCL74_2),.clk(gclk));
	jdff dff_B_Yd3ecm9v4_2(.din(w_dff_B_Q1hnPCL74_2),.dout(w_dff_B_Yd3ecm9v4_2),.clk(gclk));
	jdff dff_B_vj0XLNQO7_2(.din(w_dff_B_Yd3ecm9v4_2),.dout(w_dff_B_vj0XLNQO7_2),.clk(gclk));
	jdff dff_B_IgYLrSL78_1(.din(n930),.dout(w_dff_B_IgYLrSL78_1),.clk(gclk));
	jdff dff_B_5z43T4jN0_2(.din(n827),.dout(w_dff_B_5z43T4jN0_2),.clk(gclk));
	jdff dff_B_osFMsEJI5_2(.din(w_dff_B_5z43T4jN0_2),.dout(w_dff_B_osFMsEJI5_2),.clk(gclk));
	jdff dff_B_oaULlXjH1_2(.din(w_dff_B_osFMsEJI5_2),.dout(w_dff_B_oaULlXjH1_2),.clk(gclk));
	jdff dff_B_kUScHdvo7_2(.din(w_dff_B_oaULlXjH1_2),.dout(w_dff_B_kUScHdvo7_2),.clk(gclk));
	jdff dff_B_W4eOKzJo8_2(.din(w_dff_B_kUScHdvo7_2),.dout(w_dff_B_W4eOKzJo8_2),.clk(gclk));
	jdff dff_B_0ynQCqX17_2(.din(w_dff_B_W4eOKzJo8_2),.dout(w_dff_B_0ynQCqX17_2),.clk(gclk));
	jdff dff_B_ybum0CE36_2(.din(w_dff_B_0ynQCqX17_2),.dout(w_dff_B_ybum0CE36_2),.clk(gclk));
	jdff dff_B_W0s8vepI0_2(.din(w_dff_B_ybum0CE36_2),.dout(w_dff_B_W0s8vepI0_2),.clk(gclk));
	jdff dff_B_Jqq5HyYy1_2(.din(w_dff_B_W0s8vepI0_2),.dout(w_dff_B_Jqq5HyYy1_2),.clk(gclk));
	jdff dff_B_X6MYm6fk0_2(.din(w_dff_B_Jqq5HyYy1_2),.dout(w_dff_B_X6MYm6fk0_2),.clk(gclk));
	jdff dff_B_HQn0aSlA1_2(.din(w_dff_B_X6MYm6fk0_2),.dout(w_dff_B_HQn0aSlA1_2),.clk(gclk));
	jdff dff_B_botQhHke8_2(.din(w_dff_B_HQn0aSlA1_2),.dout(w_dff_B_botQhHke8_2),.clk(gclk));
	jdff dff_B_AJTH37Jc3_2(.din(w_dff_B_botQhHke8_2),.dout(w_dff_B_AJTH37Jc3_2),.clk(gclk));
	jdff dff_B_M9ftNkC68_2(.din(w_dff_B_AJTH37Jc3_2),.dout(w_dff_B_M9ftNkC68_2),.clk(gclk));
	jdff dff_B_DCeyKkLr8_2(.din(w_dff_B_M9ftNkC68_2),.dout(w_dff_B_DCeyKkLr8_2),.clk(gclk));
	jdff dff_B_nChQowO27_2(.din(w_dff_B_DCeyKkLr8_2),.dout(w_dff_B_nChQowO27_2),.clk(gclk));
	jdff dff_B_XVfgfJ087_2(.din(w_dff_B_nChQowO27_2),.dout(w_dff_B_XVfgfJ087_2),.clk(gclk));
	jdff dff_B_vatxhv1J4_2(.din(w_dff_B_XVfgfJ087_2),.dout(w_dff_B_vatxhv1J4_2),.clk(gclk));
	jdff dff_B_Mhx8t4Wy6_2(.din(w_dff_B_vatxhv1J4_2),.dout(w_dff_B_Mhx8t4Wy6_2),.clk(gclk));
	jdff dff_B_GUTVttjz0_2(.din(w_dff_B_Mhx8t4Wy6_2),.dout(w_dff_B_GUTVttjz0_2),.clk(gclk));
	jdff dff_B_cd3ljYx34_2(.din(w_dff_B_GUTVttjz0_2),.dout(w_dff_B_cd3ljYx34_2),.clk(gclk));
	jdff dff_B_Xw0xS6fW9_2(.din(w_dff_B_cd3ljYx34_2),.dout(w_dff_B_Xw0xS6fW9_2),.clk(gclk));
	jdff dff_B_ZSvXv55q1_2(.din(w_dff_B_Xw0xS6fW9_2),.dout(w_dff_B_ZSvXv55q1_2),.clk(gclk));
	jdff dff_B_Ur8YsLTJ9_2(.din(w_dff_B_ZSvXv55q1_2),.dout(w_dff_B_Ur8YsLTJ9_2),.clk(gclk));
	jdff dff_B_iZxUeO794_1(.din(n828),.dout(w_dff_B_iZxUeO794_1),.clk(gclk));
	jdff dff_B_9cHXJ6xI4_2(.din(n729),.dout(w_dff_B_9cHXJ6xI4_2),.clk(gclk));
	jdff dff_B_sHQsWBYe6_2(.din(w_dff_B_9cHXJ6xI4_2),.dout(w_dff_B_sHQsWBYe6_2),.clk(gclk));
	jdff dff_B_9O5Fk8Eq5_2(.din(w_dff_B_sHQsWBYe6_2),.dout(w_dff_B_9O5Fk8Eq5_2),.clk(gclk));
	jdff dff_B_QM5ycwpm5_2(.din(w_dff_B_9O5Fk8Eq5_2),.dout(w_dff_B_QM5ycwpm5_2),.clk(gclk));
	jdff dff_B_yIE2lwhV0_2(.din(w_dff_B_QM5ycwpm5_2),.dout(w_dff_B_yIE2lwhV0_2),.clk(gclk));
	jdff dff_B_J3tXTG7J3_2(.din(w_dff_B_yIE2lwhV0_2),.dout(w_dff_B_J3tXTG7J3_2),.clk(gclk));
	jdff dff_B_Fbg5e6d12_2(.din(w_dff_B_J3tXTG7J3_2),.dout(w_dff_B_Fbg5e6d12_2),.clk(gclk));
	jdff dff_B_ewcdukZ63_2(.din(w_dff_B_Fbg5e6d12_2),.dout(w_dff_B_ewcdukZ63_2),.clk(gclk));
	jdff dff_B_cCy0cV929_2(.din(w_dff_B_ewcdukZ63_2),.dout(w_dff_B_cCy0cV929_2),.clk(gclk));
	jdff dff_B_C3praiYw1_2(.din(w_dff_B_cCy0cV929_2),.dout(w_dff_B_C3praiYw1_2),.clk(gclk));
	jdff dff_B_9DzhZU3b4_2(.din(w_dff_B_C3praiYw1_2),.dout(w_dff_B_9DzhZU3b4_2),.clk(gclk));
	jdff dff_B_Ay1k8pSE1_2(.din(w_dff_B_9DzhZU3b4_2),.dout(w_dff_B_Ay1k8pSE1_2),.clk(gclk));
	jdff dff_B_sygk0zuw1_2(.din(w_dff_B_Ay1k8pSE1_2),.dout(w_dff_B_sygk0zuw1_2),.clk(gclk));
	jdff dff_B_CxEx6bgT6_2(.din(w_dff_B_sygk0zuw1_2),.dout(w_dff_B_CxEx6bgT6_2),.clk(gclk));
	jdff dff_B_d3lIxQyf4_2(.din(w_dff_B_CxEx6bgT6_2),.dout(w_dff_B_d3lIxQyf4_2),.clk(gclk));
	jdff dff_B_4ZWSruHv7_2(.din(w_dff_B_d3lIxQyf4_2),.dout(w_dff_B_4ZWSruHv7_2),.clk(gclk));
	jdff dff_B_xO1b3bP35_2(.din(w_dff_B_4ZWSruHv7_2),.dout(w_dff_B_xO1b3bP35_2),.clk(gclk));
	jdff dff_B_DdJNGzU95_2(.din(w_dff_B_xO1b3bP35_2),.dout(w_dff_B_DdJNGzU95_2),.clk(gclk));
	jdff dff_B_5AbjnurS8_2(.din(w_dff_B_DdJNGzU95_2),.dout(w_dff_B_5AbjnurS8_2),.clk(gclk));
	jdff dff_B_4y032KLj5_2(.din(w_dff_B_5AbjnurS8_2),.dout(w_dff_B_4y032KLj5_2),.clk(gclk));
	jdff dff_B_02o7Fihr9_2(.din(w_dff_B_4y032KLj5_2),.dout(w_dff_B_02o7Fihr9_2),.clk(gclk));
	jdff dff_B_0G4BkaBJ6_2(.din(w_dff_B_02o7Fihr9_2),.dout(w_dff_B_0G4BkaBJ6_2),.clk(gclk));
	jdff dff_B_kYgnMuZK0_1(.din(n730),.dout(w_dff_B_kYgnMuZK0_1),.clk(gclk));
	jdff dff_B_HBoshp425_2(.din(n637),.dout(w_dff_B_HBoshp425_2),.clk(gclk));
	jdff dff_B_nkw0MnBp6_2(.din(w_dff_B_HBoshp425_2),.dout(w_dff_B_nkw0MnBp6_2),.clk(gclk));
	jdff dff_B_fRh20S9b6_2(.din(w_dff_B_nkw0MnBp6_2),.dout(w_dff_B_fRh20S9b6_2),.clk(gclk));
	jdff dff_B_vsnzFCqZ0_2(.din(w_dff_B_fRh20S9b6_2),.dout(w_dff_B_vsnzFCqZ0_2),.clk(gclk));
	jdff dff_B_qDvcuv0O4_2(.din(w_dff_B_vsnzFCqZ0_2),.dout(w_dff_B_qDvcuv0O4_2),.clk(gclk));
	jdff dff_B_JK8jTcXB1_2(.din(w_dff_B_qDvcuv0O4_2),.dout(w_dff_B_JK8jTcXB1_2),.clk(gclk));
	jdff dff_B_gKb7bFUd0_2(.din(w_dff_B_JK8jTcXB1_2),.dout(w_dff_B_gKb7bFUd0_2),.clk(gclk));
	jdff dff_B_mMyExi168_2(.din(w_dff_B_gKb7bFUd0_2),.dout(w_dff_B_mMyExi168_2),.clk(gclk));
	jdff dff_B_uc6FLzr96_2(.din(w_dff_B_mMyExi168_2),.dout(w_dff_B_uc6FLzr96_2),.clk(gclk));
	jdff dff_B_Cw5oPujT1_2(.din(w_dff_B_uc6FLzr96_2),.dout(w_dff_B_Cw5oPujT1_2),.clk(gclk));
	jdff dff_B_zDvQVPR20_2(.din(w_dff_B_Cw5oPujT1_2),.dout(w_dff_B_zDvQVPR20_2),.clk(gclk));
	jdff dff_B_NL9AJev91_2(.din(w_dff_B_zDvQVPR20_2),.dout(w_dff_B_NL9AJev91_2),.clk(gclk));
	jdff dff_B_RKhk3fWy1_2(.din(w_dff_B_NL9AJev91_2),.dout(w_dff_B_RKhk3fWy1_2),.clk(gclk));
	jdff dff_B_3Uosf91N7_2(.din(w_dff_B_RKhk3fWy1_2),.dout(w_dff_B_3Uosf91N7_2),.clk(gclk));
	jdff dff_B_cUKRWuIn6_2(.din(w_dff_B_3Uosf91N7_2),.dout(w_dff_B_cUKRWuIn6_2),.clk(gclk));
	jdff dff_B_MfjPzDl48_2(.din(w_dff_B_cUKRWuIn6_2),.dout(w_dff_B_MfjPzDl48_2),.clk(gclk));
	jdff dff_B_6yAjG21H0_2(.din(w_dff_B_MfjPzDl48_2),.dout(w_dff_B_6yAjG21H0_2),.clk(gclk));
	jdff dff_B_0qJcRvyU2_2(.din(w_dff_B_6yAjG21H0_2),.dout(w_dff_B_0qJcRvyU2_2),.clk(gclk));
	jdff dff_B_F7WlKSiL1_2(.din(w_dff_B_0qJcRvyU2_2),.dout(w_dff_B_F7WlKSiL1_2),.clk(gclk));
	jdff dff_B_Ja40IbTs7_2(.din(w_dff_B_F7WlKSiL1_2),.dout(w_dff_B_Ja40IbTs7_2),.clk(gclk));
	jdff dff_B_EzN5P6Er8_1(.din(n638),.dout(w_dff_B_EzN5P6Er8_1),.clk(gclk));
	jdff dff_B_WXFOOucF5_2(.din(n552),.dout(w_dff_B_WXFOOucF5_2),.clk(gclk));
	jdff dff_B_wavBGGTY4_2(.din(w_dff_B_WXFOOucF5_2),.dout(w_dff_B_wavBGGTY4_2),.clk(gclk));
	jdff dff_B_rBodl2Rl4_2(.din(w_dff_B_wavBGGTY4_2),.dout(w_dff_B_rBodl2Rl4_2),.clk(gclk));
	jdff dff_B_yjVaAvJd5_2(.din(w_dff_B_rBodl2Rl4_2),.dout(w_dff_B_yjVaAvJd5_2),.clk(gclk));
	jdff dff_B_p7n8aCKs6_2(.din(w_dff_B_yjVaAvJd5_2),.dout(w_dff_B_p7n8aCKs6_2),.clk(gclk));
	jdff dff_B_FBVDvcvc4_2(.din(w_dff_B_p7n8aCKs6_2),.dout(w_dff_B_FBVDvcvc4_2),.clk(gclk));
	jdff dff_B_RigZRfyr4_2(.din(w_dff_B_FBVDvcvc4_2),.dout(w_dff_B_RigZRfyr4_2),.clk(gclk));
	jdff dff_B_TcRFPIOC3_2(.din(w_dff_B_RigZRfyr4_2),.dout(w_dff_B_TcRFPIOC3_2),.clk(gclk));
	jdff dff_B_AfJC8Fe28_2(.din(w_dff_B_TcRFPIOC3_2),.dout(w_dff_B_AfJC8Fe28_2),.clk(gclk));
	jdff dff_B_sqLUfVGh3_2(.din(w_dff_B_AfJC8Fe28_2),.dout(w_dff_B_sqLUfVGh3_2),.clk(gclk));
	jdff dff_B_szrtYhym2_2(.din(w_dff_B_sqLUfVGh3_2),.dout(w_dff_B_szrtYhym2_2),.clk(gclk));
	jdff dff_B_ZGLPVILf7_2(.din(w_dff_B_szrtYhym2_2),.dout(w_dff_B_ZGLPVILf7_2),.clk(gclk));
	jdff dff_B_Ic8f7Rbe8_2(.din(w_dff_B_ZGLPVILf7_2),.dout(w_dff_B_Ic8f7Rbe8_2),.clk(gclk));
	jdff dff_B_VJQ29aMe2_2(.din(w_dff_B_Ic8f7Rbe8_2),.dout(w_dff_B_VJQ29aMe2_2),.clk(gclk));
	jdff dff_B_yik2uola1_2(.din(w_dff_B_VJQ29aMe2_2),.dout(w_dff_B_yik2uola1_2),.clk(gclk));
	jdff dff_B_sApg5KCq0_2(.din(w_dff_B_yik2uola1_2),.dout(w_dff_B_sApg5KCq0_2),.clk(gclk));
	jdff dff_B_wxNgrRG15_2(.din(w_dff_B_sApg5KCq0_2),.dout(w_dff_B_wxNgrRG15_2),.clk(gclk));
	jdff dff_B_dGoD1wjK8_2(.din(w_dff_B_wxNgrRG15_2),.dout(w_dff_B_dGoD1wjK8_2),.clk(gclk));
	jdff dff_B_2Ytn0KlC5_1(.din(n553),.dout(w_dff_B_2Ytn0KlC5_1),.clk(gclk));
	jdff dff_B_wQeodYbi4_2(.din(n474),.dout(w_dff_B_wQeodYbi4_2),.clk(gclk));
	jdff dff_B_WTx0HzLt9_2(.din(w_dff_B_wQeodYbi4_2),.dout(w_dff_B_WTx0HzLt9_2),.clk(gclk));
	jdff dff_B_OzfKQF338_2(.din(w_dff_B_WTx0HzLt9_2),.dout(w_dff_B_OzfKQF338_2),.clk(gclk));
	jdff dff_B_aSKDJZTm6_2(.din(w_dff_B_OzfKQF338_2),.dout(w_dff_B_aSKDJZTm6_2),.clk(gclk));
	jdff dff_B_YLyfWVB10_2(.din(w_dff_B_aSKDJZTm6_2),.dout(w_dff_B_YLyfWVB10_2),.clk(gclk));
	jdff dff_B_IPgcPpcI5_2(.din(w_dff_B_YLyfWVB10_2),.dout(w_dff_B_IPgcPpcI5_2),.clk(gclk));
	jdff dff_B_P6X41ltl8_2(.din(w_dff_B_IPgcPpcI5_2),.dout(w_dff_B_P6X41ltl8_2),.clk(gclk));
	jdff dff_B_rzKKLRbA1_2(.din(w_dff_B_P6X41ltl8_2),.dout(w_dff_B_rzKKLRbA1_2),.clk(gclk));
	jdff dff_B_wmkluPFv3_2(.din(w_dff_B_rzKKLRbA1_2),.dout(w_dff_B_wmkluPFv3_2),.clk(gclk));
	jdff dff_B_zY3c43w38_2(.din(w_dff_B_wmkluPFv3_2),.dout(w_dff_B_zY3c43w38_2),.clk(gclk));
	jdff dff_B_EyvNzULS8_2(.din(w_dff_B_zY3c43w38_2),.dout(w_dff_B_EyvNzULS8_2),.clk(gclk));
	jdff dff_B_GeqNlMIE0_2(.din(w_dff_B_EyvNzULS8_2),.dout(w_dff_B_GeqNlMIE0_2),.clk(gclk));
	jdff dff_B_R0ZR6iCs3_2(.din(w_dff_B_GeqNlMIE0_2),.dout(w_dff_B_R0ZR6iCs3_2),.clk(gclk));
	jdff dff_B_ULEgfoCS9_2(.din(w_dff_B_R0ZR6iCs3_2),.dout(w_dff_B_ULEgfoCS9_2),.clk(gclk));
	jdff dff_B_nAuwTMlj1_2(.din(w_dff_B_ULEgfoCS9_2),.dout(w_dff_B_nAuwTMlj1_2),.clk(gclk));
	jdff dff_B_r65m0gHm0_2(.din(w_dff_B_nAuwTMlj1_2),.dout(w_dff_B_r65m0gHm0_2),.clk(gclk));
	jdff dff_B_tc797yZk2_1(.din(n475),.dout(w_dff_B_tc797yZk2_1),.clk(gclk));
	jdff dff_B_SLa7yIMe6_2(.din(n403),.dout(w_dff_B_SLa7yIMe6_2),.clk(gclk));
	jdff dff_B_MjdljAZ27_2(.din(w_dff_B_SLa7yIMe6_2),.dout(w_dff_B_MjdljAZ27_2),.clk(gclk));
	jdff dff_B_T9xnokmU6_2(.din(w_dff_B_MjdljAZ27_2),.dout(w_dff_B_T9xnokmU6_2),.clk(gclk));
	jdff dff_B_RsNr5UGG1_2(.din(w_dff_B_T9xnokmU6_2),.dout(w_dff_B_RsNr5UGG1_2),.clk(gclk));
	jdff dff_B_SaLhkhMA3_2(.din(w_dff_B_RsNr5UGG1_2),.dout(w_dff_B_SaLhkhMA3_2),.clk(gclk));
	jdff dff_B_kBQ8eeqa9_2(.din(w_dff_B_SaLhkhMA3_2),.dout(w_dff_B_kBQ8eeqa9_2),.clk(gclk));
	jdff dff_B_H22V1JKQ9_2(.din(w_dff_B_kBQ8eeqa9_2),.dout(w_dff_B_H22V1JKQ9_2),.clk(gclk));
	jdff dff_B_7eeRBTvC4_2(.din(w_dff_B_H22V1JKQ9_2),.dout(w_dff_B_7eeRBTvC4_2),.clk(gclk));
	jdff dff_B_FONr2Ja70_2(.din(w_dff_B_7eeRBTvC4_2),.dout(w_dff_B_FONr2Ja70_2),.clk(gclk));
	jdff dff_B_PF6eVLh83_2(.din(w_dff_B_FONr2Ja70_2),.dout(w_dff_B_PF6eVLh83_2),.clk(gclk));
	jdff dff_B_WlMjQp025_2(.din(w_dff_B_PF6eVLh83_2),.dout(w_dff_B_WlMjQp025_2),.clk(gclk));
	jdff dff_B_cJwP2DIY5_2(.din(w_dff_B_WlMjQp025_2),.dout(w_dff_B_cJwP2DIY5_2),.clk(gclk));
	jdff dff_B_L1DTu0oL3_2(.din(w_dff_B_cJwP2DIY5_2),.dout(w_dff_B_L1DTu0oL3_2),.clk(gclk));
	jdff dff_B_1MUQayca2_2(.din(w_dff_B_L1DTu0oL3_2),.dout(w_dff_B_1MUQayca2_2),.clk(gclk));
	jdff dff_B_ZtbhKuhs5_2(.din(n406),.dout(w_dff_B_ZtbhKuhs5_2),.clk(gclk));
	jdff dff_B_ajzQoUT25_2(.din(w_dff_B_ZtbhKuhs5_2),.dout(w_dff_B_ajzQoUT25_2),.clk(gclk));
	jdff dff_B_M9Ywdoct1_2(.din(w_dff_B_ajzQoUT25_2),.dout(w_dff_B_M9Ywdoct1_2),.clk(gclk));
	jdff dff_B_4ZkH0V4J4_1(.din(n404),.dout(w_dff_B_4ZkH0V4J4_1),.clk(gclk));
	jdff dff_B_4wZV470f8_2(.din(n340),.dout(w_dff_B_4wZV470f8_2),.clk(gclk));
	jdff dff_B_93m99Vn68_2(.din(w_dff_B_4wZV470f8_2),.dout(w_dff_B_93m99Vn68_2),.clk(gclk));
	jdff dff_B_c70jGVwM6_2(.din(w_dff_B_93m99Vn68_2),.dout(w_dff_B_c70jGVwM6_2),.clk(gclk));
	jdff dff_B_9bfqCtGY2_2(.din(w_dff_B_c70jGVwM6_2),.dout(w_dff_B_9bfqCtGY2_2),.clk(gclk));
	jdff dff_B_XrNXuaAF4_2(.din(w_dff_B_9bfqCtGY2_2),.dout(w_dff_B_XrNXuaAF4_2),.clk(gclk));
	jdff dff_B_HTD27yKz0_2(.din(w_dff_B_XrNXuaAF4_2),.dout(w_dff_B_HTD27yKz0_2),.clk(gclk));
	jdff dff_B_MkPgHLIU9_2(.din(w_dff_B_HTD27yKz0_2),.dout(w_dff_B_MkPgHLIU9_2),.clk(gclk));
	jdff dff_B_SkejRnpn0_2(.din(w_dff_B_MkPgHLIU9_2),.dout(w_dff_B_SkejRnpn0_2),.clk(gclk));
	jdff dff_B_4Dj13Jvy2_2(.din(w_dff_B_SkejRnpn0_2),.dout(w_dff_B_4Dj13Jvy2_2),.clk(gclk));
	jdff dff_B_OsDt93ur4_1(.din(n341),.dout(w_dff_B_OsDt93ur4_1),.clk(gclk));
	jdff dff_B_8VvdAJ4d8_2(.din(n284),.dout(w_dff_B_8VvdAJ4d8_2),.clk(gclk));
	jdff dff_B_JltM7ZGy5_2(.din(w_dff_B_8VvdAJ4d8_2),.dout(w_dff_B_JltM7ZGy5_2),.clk(gclk));
	jdff dff_B_aJGVUg9q7_2(.din(w_dff_B_JltM7ZGy5_2),.dout(w_dff_B_aJGVUg9q7_2),.clk(gclk));
	jdff dff_B_3juZpKTG2_2(.din(w_dff_B_aJGVUg9q7_2),.dout(w_dff_B_3juZpKTG2_2),.clk(gclk));
	jdff dff_B_qgUAGqRV7_2(.din(w_dff_B_3juZpKTG2_2),.dout(w_dff_B_qgUAGqRV7_2),.clk(gclk));
	jdff dff_B_z7lCqZki2_2(.din(w_dff_B_qgUAGqRV7_2),.dout(w_dff_B_z7lCqZki2_2),.clk(gclk));
	jdff dff_B_dbs0Nf4r4_2(.din(w_dff_B_z7lCqZki2_2),.dout(w_dff_B_dbs0Nf4r4_2),.clk(gclk));
	jdff dff_B_Z0Y6Bzw53_1(.din(n285),.dout(w_dff_B_Z0Y6Bzw53_1),.clk(gclk));
	jdff dff_B_TkU64rgP2_2(.din(n235),.dout(w_dff_B_TkU64rgP2_2),.clk(gclk));
	jdff dff_B_jvU8bwhf6_2(.din(w_dff_B_TkU64rgP2_2),.dout(w_dff_B_jvU8bwhf6_2),.clk(gclk));
	jdff dff_B_TQSGHHTO7_2(.din(w_dff_B_jvU8bwhf6_2),.dout(w_dff_B_TQSGHHTO7_2),.clk(gclk));
	jdff dff_B_Dv1DFU4c7_2(.din(w_dff_B_TQSGHHTO7_2),.dout(w_dff_B_Dv1DFU4c7_2),.clk(gclk));
	jdff dff_B_2vHWrEiA8_2(.din(w_dff_B_Dv1DFU4c7_2),.dout(w_dff_B_2vHWrEiA8_2),.clk(gclk));
	jdff dff_B_3i3vPdau4_2(.din(n194),.dout(w_dff_B_3i3vPdau4_2),.clk(gclk));
	jdff dff_B_rjgJwLKB0_2(.din(w_dff_B_3i3vPdau4_2),.dout(w_dff_B_rjgJwLKB0_2),.clk(gclk));
	jdff dff_B_cbd2tEGR6_2(.din(w_dff_B_rjgJwLKB0_2),.dout(w_dff_B_cbd2tEGR6_2),.clk(gclk));
	jdff dff_B_AJL1rbdl4_0(.din(n199),.dout(w_dff_B_AJL1rbdl4_0),.clk(gclk));
	jdff dff_B_wD40bFgi9_0(.din(w_dff_B_AJL1rbdl4_0),.dout(w_dff_B_wD40bFgi9_0),.clk(gclk));
	jdff dff_A_820aAthH5_0(.dout(w_n157_0[0]),.din(w_dff_A_820aAthH5_0),.clk(gclk));
	jdff dff_A_VFk9IOOo6_0(.dout(w_dff_A_820aAthH5_0),.din(w_dff_A_VFk9IOOo6_0),.clk(gclk));
	jdff dff_A_RJf1Y65M4_0(.dout(w_n156_0[0]),.din(w_dff_A_RJf1Y65M4_0),.clk(gclk));
	jdff dff_A_lXNE1JWt6_0(.dout(w_dff_A_RJf1Y65M4_0),.din(w_dff_A_lXNE1JWt6_0),.clk(gclk));
	jdff dff_B_2s9dHElE5_2(.din(n1389),.dout(w_dff_B_2s9dHElE5_2),.clk(gclk));
	jdff dff_B_X5KheESI6_2(.din(w_dff_B_2s9dHElE5_2),.dout(w_dff_B_X5KheESI6_2),.clk(gclk));
	jdff dff_B_pruoaOri4_1(.din(n1387),.dout(w_dff_B_pruoaOri4_1),.clk(gclk));
	jdff dff_B_jfR6X47k4_2(.din(n1307),.dout(w_dff_B_jfR6X47k4_2),.clk(gclk));
	jdff dff_B_S6g40pB57_2(.din(w_dff_B_jfR6X47k4_2),.dout(w_dff_B_S6g40pB57_2),.clk(gclk));
	jdff dff_B_egYGi1Od2_2(.din(w_dff_B_S6g40pB57_2),.dout(w_dff_B_egYGi1Od2_2),.clk(gclk));
	jdff dff_B_j2jZ3IJz0_2(.din(w_dff_B_egYGi1Od2_2),.dout(w_dff_B_j2jZ3IJz0_2),.clk(gclk));
	jdff dff_B_pg1SXlAp3_2(.din(w_dff_B_j2jZ3IJz0_2),.dout(w_dff_B_pg1SXlAp3_2),.clk(gclk));
	jdff dff_B_zZ3ICMPW7_2(.din(w_dff_B_pg1SXlAp3_2),.dout(w_dff_B_zZ3ICMPW7_2),.clk(gclk));
	jdff dff_B_wNnTB0qN1_2(.din(w_dff_B_zZ3ICMPW7_2),.dout(w_dff_B_wNnTB0qN1_2),.clk(gclk));
	jdff dff_B_YkCeicYp4_2(.din(w_dff_B_wNnTB0qN1_2),.dout(w_dff_B_YkCeicYp4_2),.clk(gclk));
	jdff dff_B_nhXQ1pFN1_2(.din(w_dff_B_YkCeicYp4_2),.dout(w_dff_B_nhXQ1pFN1_2),.clk(gclk));
	jdff dff_B_FDa1bFrG2_2(.din(w_dff_B_nhXQ1pFN1_2),.dout(w_dff_B_FDa1bFrG2_2),.clk(gclk));
	jdff dff_B_KerW6clm1_2(.din(w_dff_B_FDa1bFrG2_2),.dout(w_dff_B_KerW6clm1_2),.clk(gclk));
	jdff dff_B_HIzLqiIZ4_2(.din(w_dff_B_KerW6clm1_2),.dout(w_dff_B_HIzLqiIZ4_2),.clk(gclk));
	jdff dff_B_47Yn0VEd5_2(.din(w_dff_B_HIzLqiIZ4_2),.dout(w_dff_B_47Yn0VEd5_2),.clk(gclk));
	jdff dff_B_6WAwCxhE8_2(.din(w_dff_B_47Yn0VEd5_2),.dout(w_dff_B_6WAwCxhE8_2),.clk(gclk));
	jdff dff_B_yzTges2q8_2(.din(w_dff_B_6WAwCxhE8_2),.dout(w_dff_B_yzTges2q8_2),.clk(gclk));
	jdff dff_B_yLXEaxdp0_2(.din(w_dff_B_yzTges2q8_2),.dout(w_dff_B_yLXEaxdp0_2),.clk(gclk));
	jdff dff_B_0ZxJP1fF8_2(.din(w_dff_B_yLXEaxdp0_2),.dout(w_dff_B_0ZxJP1fF8_2),.clk(gclk));
	jdff dff_B_jaGU8V821_2(.din(w_dff_B_0ZxJP1fF8_2),.dout(w_dff_B_jaGU8V821_2),.clk(gclk));
	jdff dff_B_C7ykZp4v7_2(.din(w_dff_B_jaGU8V821_2),.dout(w_dff_B_C7ykZp4v7_2),.clk(gclk));
	jdff dff_B_N3dAI3l63_2(.din(w_dff_B_C7ykZp4v7_2),.dout(w_dff_B_N3dAI3l63_2),.clk(gclk));
	jdff dff_B_oY7ajPEx9_2(.din(w_dff_B_N3dAI3l63_2),.dout(w_dff_B_oY7ajPEx9_2),.clk(gclk));
	jdff dff_B_rfZ8eDUg8_2(.din(w_dff_B_oY7ajPEx9_2),.dout(w_dff_B_rfZ8eDUg8_2),.clk(gclk));
	jdff dff_B_uNHoWAuO3_2(.din(w_dff_B_rfZ8eDUg8_2),.dout(w_dff_B_uNHoWAuO3_2),.clk(gclk));
	jdff dff_B_JKbuB6Mc2_2(.din(w_dff_B_uNHoWAuO3_2),.dout(w_dff_B_JKbuB6Mc2_2),.clk(gclk));
	jdff dff_B_MYCLVb5o7_2(.din(w_dff_B_JKbuB6Mc2_2),.dout(w_dff_B_MYCLVb5o7_2),.clk(gclk));
	jdff dff_B_aWeAeoS14_2(.din(w_dff_B_MYCLVb5o7_2),.dout(w_dff_B_aWeAeoS14_2),.clk(gclk));
	jdff dff_B_fEu038fv1_2(.din(w_dff_B_aWeAeoS14_2),.dout(w_dff_B_fEu038fv1_2),.clk(gclk));
	jdff dff_B_2JtvUI9V8_2(.din(w_dff_B_fEu038fv1_2),.dout(w_dff_B_2JtvUI9V8_2),.clk(gclk));
	jdff dff_B_VIa1jW1B9_2(.din(w_dff_B_2JtvUI9V8_2),.dout(w_dff_B_VIa1jW1B9_2),.clk(gclk));
	jdff dff_B_cDG4JfW54_2(.din(w_dff_B_VIa1jW1B9_2),.dout(w_dff_B_cDG4JfW54_2),.clk(gclk));
	jdff dff_B_qGzVz2qc0_2(.din(w_dff_B_cDG4JfW54_2),.dout(w_dff_B_qGzVz2qc0_2),.clk(gclk));
	jdff dff_B_VAvZLqhF2_2(.din(w_dff_B_qGzVz2qc0_2),.dout(w_dff_B_VAvZLqhF2_2),.clk(gclk));
	jdff dff_B_pgCfMrz43_2(.din(w_dff_B_VAvZLqhF2_2),.dout(w_dff_B_pgCfMrz43_2),.clk(gclk));
	jdff dff_B_khNyTxgR1_2(.din(w_dff_B_pgCfMrz43_2),.dout(w_dff_B_khNyTxgR1_2),.clk(gclk));
	jdff dff_B_v3VgPoVA6_1(.din(n1308),.dout(w_dff_B_v3VgPoVA6_1),.clk(gclk));
	jdff dff_B_IhY0Ds3Z3_2(.din(n1222),.dout(w_dff_B_IhY0Ds3Z3_2),.clk(gclk));
	jdff dff_B_LjXWS6AA4_2(.din(w_dff_B_IhY0Ds3Z3_2),.dout(w_dff_B_LjXWS6AA4_2),.clk(gclk));
	jdff dff_B_JBSmMM8z3_2(.din(w_dff_B_LjXWS6AA4_2),.dout(w_dff_B_JBSmMM8z3_2),.clk(gclk));
	jdff dff_B_iBL2XGxJ0_2(.din(w_dff_B_JBSmMM8z3_2),.dout(w_dff_B_iBL2XGxJ0_2),.clk(gclk));
	jdff dff_B_JMwULktA3_2(.din(w_dff_B_iBL2XGxJ0_2),.dout(w_dff_B_JMwULktA3_2),.clk(gclk));
	jdff dff_B_RbmOlHMq9_2(.din(w_dff_B_JMwULktA3_2),.dout(w_dff_B_RbmOlHMq9_2),.clk(gclk));
	jdff dff_B_3yGlt62V6_2(.din(w_dff_B_RbmOlHMq9_2),.dout(w_dff_B_3yGlt62V6_2),.clk(gclk));
	jdff dff_B_WxdKZAMv8_2(.din(w_dff_B_3yGlt62V6_2),.dout(w_dff_B_WxdKZAMv8_2),.clk(gclk));
	jdff dff_B_MGBRD87w4_2(.din(w_dff_B_WxdKZAMv8_2),.dout(w_dff_B_MGBRD87w4_2),.clk(gclk));
	jdff dff_B_XHs01P0X9_2(.din(w_dff_B_MGBRD87w4_2),.dout(w_dff_B_XHs01P0X9_2),.clk(gclk));
	jdff dff_B_qOayNJGz0_2(.din(w_dff_B_XHs01P0X9_2),.dout(w_dff_B_qOayNJGz0_2),.clk(gclk));
	jdff dff_B_BYuex7We0_2(.din(w_dff_B_qOayNJGz0_2),.dout(w_dff_B_BYuex7We0_2),.clk(gclk));
	jdff dff_B_DmutNhWQ5_2(.din(w_dff_B_BYuex7We0_2),.dout(w_dff_B_DmutNhWQ5_2),.clk(gclk));
	jdff dff_B_F6OMPAFq7_2(.din(w_dff_B_DmutNhWQ5_2),.dout(w_dff_B_F6OMPAFq7_2),.clk(gclk));
	jdff dff_B_1RU4xIcQ4_2(.din(w_dff_B_F6OMPAFq7_2),.dout(w_dff_B_1RU4xIcQ4_2),.clk(gclk));
	jdff dff_B_Zw3rbi1D3_2(.din(w_dff_B_1RU4xIcQ4_2),.dout(w_dff_B_Zw3rbi1D3_2),.clk(gclk));
	jdff dff_B_N7wWm7Uv0_2(.din(w_dff_B_Zw3rbi1D3_2),.dout(w_dff_B_N7wWm7Uv0_2),.clk(gclk));
	jdff dff_B_SZxqN9x08_2(.din(w_dff_B_N7wWm7Uv0_2),.dout(w_dff_B_SZxqN9x08_2),.clk(gclk));
	jdff dff_B_gR8OEe0h9_2(.din(w_dff_B_SZxqN9x08_2),.dout(w_dff_B_gR8OEe0h9_2),.clk(gclk));
	jdff dff_B_eptCr87L8_2(.din(w_dff_B_gR8OEe0h9_2),.dout(w_dff_B_eptCr87L8_2),.clk(gclk));
	jdff dff_B_ma5NMSMI8_2(.din(w_dff_B_eptCr87L8_2),.dout(w_dff_B_ma5NMSMI8_2),.clk(gclk));
	jdff dff_B_njf8lLwo7_2(.din(w_dff_B_ma5NMSMI8_2),.dout(w_dff_B_njf8lLwo7_2),.clk(gclk));
	jdff dff_B_MwvA4mZl4_2(.din(w_dff_B_njf8lLwo7_2),.dout(w_dff_B_MwvA4mZl4_2),.clk(gclk));
	jdff dff_B_T5KgOxh74_2(.din(w_dff_B_MwvA4mZl4_2),.dout(w_dff_B_T5KgOxh74_2),.clk(gclk));
	jdff dff_B_JX8pf6I34_2(.din(w_dff_B_T5KgOxh74_2),.dout(w_dff_B_JX8pf6I34_2),.clk(gclk));
	jdff dff_B_NqqxYUqI2_2(.din(w_dff_B_JX8pf6I34_2),.dout(w_dff_B_NqqxYUqI2_2),.clk(gclk));
	jdff dff_B_FcjemT152_2(.din(w_dff_B_NqqxYUqI2_2),.dout(w_dff_B_FcjemT152_2),.clk(gclk));
	jdff dff_B_AyQ9YqEA4_2(.din(w_dff_B_FcjemT152_2),.dout(w_dff_B_AyQ9YqEA4_2),.clk(gclk));
	jdff dff_B_zE7LPmHe3_2(.din(w_dff_B_AyQ9YqEA4_2),.dout(w_dff_B_zE7LPmHe3_2),.clk(gclk));
	jdff dff_B_9iVFdk5t0_2(.din(w_dff_B_zE7LPmHe3_2),.dout(w_dff_B_9iVFdk5t0_2),.clk(gclk));
	jdff dff_B_QxnkdtK96_1(.din(n1223),.dout(w_dff_B_QxnkdtK96_1),.clk(gclk));
	jdff dff_B_xu18Wgd63_2(.din(n1131),.dout(w_dff_B_xu18Wgd63_2),.clk(gclk));
	jdff dff_B_SHi9O1wl0_2(.din(w_dff_B_xu18Wgd63_2),.dout(w_dff_B_SHi9O1wl0_2),.clk(gclk));
	jdff dff_B_dhZIFRH02_2(.din(w_dff_B_SHi9O1wl0_2),.dout(w_dff_B_dhZIFRH02_2),.clk(gclk));
	jdff dff_B_zwdWLX4l7_2(.din(w_dff_B_dhZIFRH02_2),.dout(w_dff_B_zwdWLX4l7_2),.clk(gclk));
	jdff dff_B_HZ6uSPBh5_2(.din(w_dff_B_zwdWLX4l7_2),.dout(w_dff_B_HZ6uSPBh5_2),.clk(gclk));
	jdff dff_B_oyBnS3GN8_2(.din(w_dff_B_HZ6uSPBh5_2),.dout(w_dff_B_oyBnS3GN8_2),.clk(gclk));
	jdff dff_B_EUfySKTj9_2(.din(w_dff_B_oyBnS3GN8_2),.dout(w_dff_B_EUfySKTj9_2),.clk(gclk));
	jdff dff_B_QxWT93uW6_2(.din(w_dff_B_EUfySKTj9_2),.dout(w_dff_B_QxWT93uW6_2),.clk(gclk));
	jdff dff_B_BdxFdJig0_2(.din(w_dff_B_QxWT93uW6_2),.dout(w_dff_B_BdxFdJig0_2),.clk(gclk));
	jdff dff_B_BNMW6Qob3_2(.din(w_dff_B_BdxFdJig0_2),.dout(w_dff_B_BNMW6Qob3_2),.clk(gclk));
	jdff dff_B_LMW1Qgr25_2(.din(w_dff_B_BNMW6Qob3_2),.dout(w_dff_B_LMW1Qgr25_2),.clk(gclk));
	jdff dff_B_8pAhwc8G5_2(.din(w_dff_B_LMW1Qgr25_2),.dout(w_dff_B_8pAhwc8G5_2),.clk(gclk));
	jdff dff_B_hwozoBNM7_2(.din(w_dff_B_8pAhwc8G5_2),.dout(w_dff_B_hwozoBNM7_2),.clk(gclk));
	jdff dff_B_zjNoWVwV1_2(.din(w_dff_B_hwozoBNM7_2),.dout(w_dff_B_zjNoWVwV1_2),.clk(gclk));
	jdff dff_B_1fZK6CUp9_2(.din(w_dff_B_zjNoWVwV1_2),.dout(w_dff_B_1fZK6CUp9_2),.clk(gclk));
	jdff dff_B_Xm3JAaOh8_2(.din(w_dff_B_1fZK6CUp9_2),.dout(w_dff_B_Xm3JAaOh8_2),.clk(gclk));
	jdff dff_B_ELlgVvUu7_2(.din(w_dff_B_Xm3JAaOh8_2),.dout(w_dff_B_ELlgVvUu7_2),.clk(gclk));
	jdff dff_B_VBEBz7i95_2(.din(w_dff_B_ELlgVvUu7_2),.dout(w_dff_B_VBEBz7i95_2),.clk(gclk));
	jdff dff_B_QEwiVNKB8_2(.din(w_dff_B_VBEBz7i95_2),.dout(w_dff_B_QEwiVNKB8_2),.clk(gclk));
	jdff dff_B_EWohVFEg1_2(.din(w_dff_B_QEwiVNKB8_2),.dout(w_dff_B_EWohVFEg1_2),.clk(gclk));
	jdff dff_B_3cujJYnU6_2(.din(w_dff_B_EWohVFEg1_2),.dout(w_dff_B_3cujJYnU6_2),.clk(gclk));
	jdff dff_B_dPyV0SGM2_2(.din(w_dff_B_3cujJYnU6_2),.dout(w_dff_B_dPyV0SGM2_2),.clk(gclk));
	jdff dff_B_bVblJ1rf2_2(.din(w_dff_B_dPyV0SGM2_2),.dout(w_dff_B_bVblJ1rf2_2),.clk(gclk));
	jdff dff_B_5zbpitpD2_2(.din(w_dff_B_bVblJ1rf2_2),.dout(w_dff_B_5zbpitpD2_2),.clk(gclk));
	jdff dff_B_74hQK1698_2(.din(w_dff_B_5zbpitpD2_2),.dout(w_dff_B_74hQK1698_2),.clk(gclk));
	jdff dff_B_k8cmLbAc7_2(.din(w_dff_B_74hQK1698_2),.dout(w_dff_B_k8cmLbAc7_2),.clk(gclk));
	jdff dff_B_SrPYwD194_2(.din(w_dff_B_k8cmLbAc7_2),.dout(w_dff_B_SrPYwD194_2),.clk(gclk));
	jdff dff_B_LE4azKlA7_2(.din(w_dff_B_SrPYwD194_2),.dout(w_dff_B_LE4azKlA7_2),.clk(gclk));
	jdff dff_B_ygGrrKsO1_1(.din(n1132),.dout(w_dff_B_ygGrrKsO1_1),.clk(gclk));
	jdff dff_B_PnsullEO7_2(.din(n1033),.dout(w_dff_B_PnsullEO7_2),.clk(gclk));
	jdff dff_B_Afhpwo7d3_2(.din(w_dff_B_PnsullEO7_2),.dout(w_dff_B_Afhpwo7d3_2),.clk(gclk));
	jdff dff_B_EKWG8set4_2(.din(w_dff_B_Afhpwo7d3_2),.dout(w_dff_B_EKWG8set4_2),.clk(gclk));
	jdff dff_B_O0EhHbYA9_2(.din(w_dff_B_EKWG8set4_2),.dout(w_dff_B_O0EhHbYA9_2),.clk(gclk));
	jdff dff_B_3V7ZAs4h9_2(.din(w_dff_B_O0EhHbYA9_2),.dout(w_dff_B_3V7ZAs4h9_2),.clk(gclk));
	jdff dff_B_gtNfPWEz4_2(.din(w_dff_B_3V7ZAs4h9_2),.dout(w_dff_B_gtNfPWEz4_2),.clk(gclk));
	jdff dff_B_FajFmzDy5_2(.din(w_dff_B_gtNfPWEz4_2),.dout(w_dff_B_FajFmzDy5_2),.clk(gclk));
	jdff dff_B_vaVMa4NS6_2(.din(w_dff_B_FajFmzDy5_2),.dout(w_dff_B_vaVMa4NS6_2),.clk(gclk));
	jdff dff_B_0YTtw7uS3_2(.din(w_dff_B_vaVMa4NS6_2),.dout(w_dff_B_0YTtw7uS3_2),.clk(gclk));
	jdff dff_B_jSTZrvy77_2(.din(w_dff_B_0YTtw7uS3_2),.dout(w_dff_B_jSTZrvy77_2),.clk(gclk));
	jdff dff_B_yXsl5EKu5_2(.din(w_dff_B_jSTZrvy77_2),.dout(w_dff_B_yXsl5EKu5_2),.clk(gclk));
	jdff dff_B_Q38pz4Jj3_2(.din(w_dff_B_yXsl5EKu5_2),.dout(w_dff_B_Q38pz4Jj3_2),.clk(gclk));
	jdff dff_B_k0C6hbO88_2(.din(w_dff_B_Q38pz4Jj3_2),.dout(w_dff_B_k0C6hbO88_2),.clk(gclk));
	jdff dff_B_94O8dSav2_2(.din(w_dff_B_k0C6hbO88_2),.dout(w_dff_B_94O8dSav2_2),.clk(gclk));
	jdff dff_B_GIkOKykb1_2(.din(w_dff_B_94O8dSav2_2),.dout(w_dff_B_GIkOKykb1_2),.clk(gclk));
	jdff dff_B_lUfXqXAW7_2(.din(w_dff_B_GIkOKykb1_2),.dout(w_dff_B_lUfXqXAW7_2),.clk(gclk));
	jdff dff_B_g7poNg7U3_2(.din(w_dff_B_lUfXqXAW7_2),.dout(w_dff_B_g7poNg7U3_2),.clk(gclk));
	jdff dff_B_D5Y9i9q60_2(.din(w_dff_B_g7poNg7U3_2),.dout(w_dff_B_D5Y9i9q60_2),.clk(gclk));
	jdff dff_B_EAOmlf739_2(.din(w_dff_B_D5Y9i9q60_2),.dout(w_dff_B_EAOmlf739_2),.clk(gclk));
	jdff dff_B_WLAcfqAC3_2(.din(w_dff_B_EAOmlf739_2),.dout(w_dff_B_WLAcfqAC3_2),.clk(gclk));
	jdff dff_B_PQB1mG6v1_2(.din(w_dff_B_WLAcfqAC3_2),.dout(w_dff_B_PQB1mG6v1_2),.clk(gclk));
	jdff dff_B_1RyHKKb59_2(.din(w_dff_B_PQB1mG6v1_2),.dout(w_dff_B_1RyHKKb59_2),.clk(gclk));
	jdff dff_B_yKyGVzaj1_2(.din(w_dff_B_1RyHKKb59_2),.dout(w_dff_B_yKyGVzaj1_2),.clk(gclk));
	jdff dff_B_DO9CrTUn1_2(.din(w_dff_B_yKyGVzaj1_2),.dout(w_dff_B_DO9CrTUn1_2),.clk(gclk));
	jdff dff_B_F3mr18MV6_2(.din(w_dff_B_DO9CrTUn1_2),.dout(w_dff_B_F3mr18MV6_2),.clk(gclk));
	jdff dff_B_FeoLRdE16_2(.din(w_dff_B_F3mr18MV6_2),.dout(w_dff_B_FeoLRdE16_2),.clk(gclk));
	jdff dff_B_ED789YdO5_1(.din(n1034),.dout(w_dff_B_ED789YdO5_1),.clk(gclk));
	jdff dff_B_stRJSPrO4_2(.din(n934),.dout(w_dff_B_stRJSPrO4_2),.clk(gclk));
	jdff dff_B_uPCsLQqt9_2(.din(w_dff_B_stRJSPrO4_2),.dout(w_dff_B_uPCsLQqt9_2),.clk(gclk));
	jdff dff_B_L7yLjOHe3_2(.din(w_dff_B_uPCsLQqt9_2),.dout(w_dff_B_L7yLjOHe3_2),.clk(gclk));
	jdff dff_B_kORukNq40_2(.din(w_dff_B_L7yLjOHe3_2),.dout(w_dff_B_kORukNq40_2),.clk(gclk));
	jdff dff_B_1aKtioxn2_2(.din(w_dff_B_kORukNq40_2),.dout(w_dff_B_1aKtioxn2_2),.clk(gclk));
	jdff dff_B_UQNsoet96_2(.din(w_dff_B_1aKtioxn2_2),.dout(w_dff_B_UQNsoet96_2),.clk(gclk));
	jdff dff_B_FWI24CPp1_2(.din(w_dff_B_UQNsoet96_2),.dout(w_dff_B_FWI24CPp1_2),.clk(gclk));
	jdff dff_B_73oC28Ih7_2(.din(w_dff_B_FWI24CPp1_2),.dout(w_dff_B_73oC28Ih7_2),.clk(gclk));
	jdff dff_B_lRSgbmKP0_2(.din(w_dff_B_73oC28Ih7_2),.dout(w_dff_B_lRSgbmKP0_2),.clk(gclk));
	jdff dff_B_x7hLgs4Y7_2(.din(w_dff_B_lRSgbmKP0_2),.dout(w_dff_B_x7hLgs4Y7_2),.clk(gclk));
	jdff dff_B_d0ejrO6m1_2(.din(w_dff_B_x7hLgs4Y7_2),.dout(w_dff_B_d0ejrO6m1_2),.clk(gclk));
	jdff dff_B_n25tirG72_2(.din(w_dff_B_d0ejrO6m1_2),.dout(w_dff_B_n25tirG72_2),.clk(gclk));
	jdff dff_B_3FwuhAIb7_2(.din(w_dff_B_n25tirG72_2),.dout(w_dff_B_3FwuhAIb7_2),.clk(gclk));
	jdff dff_B_Y0w0qHtz0_2(.din(w_dff_B_3FwuhAIb7_2),.dout(w_dff_B_Y0w0qHtz0_2),.clk(gclk));
	jdff dff_B_PLRcf1md5_2(.din(w_dff_B_Y0w0qHtz0_2),.dout(w_dff_B_PLRcf1md5_2),.clk(gclk));
	jdff dff_B_yZH4XOE43_2(.din(w_dff_B_PLRcf1md5_2),.dout(w_dff_B_yZH4XOE43_2),.clk(gclk));
	jdff dff_B_CPSSX6F10_2(.din(w_dff_B_yZH4XOE43_2),.dout(w_dff_B_CPSSX6F10_2),.clk(gclk));
	jdff dff_B_bLZpHZRw5_2(.din(w_dff_B_CPSSX6F10_2),.dout(w_dff_B_bLZpHZRw5_2),.clk(gclk));
	jdff dff_B_B2LPLQhR1_2(.din(w_dff_B_bLZpHZRw5_2),.dout(w_dff_B_B2LPLQhR1_2),.clk(gclk));
	jdff dff_B_NPNT7YiW8_2(.din(w_dff_B_B2LPLQhR1_2),.dout(w_dff_B_NPNT7YiW8_2),.clk(gclk));
	jdff dff_B_UPX9w7Ht8_2(.din(w_dff_B_NPNT7YiW8_2),.dout(w_dff_B_UPX9w7Ht8_2),.clk(gclk));
	jdff dff_B_sPsAxl123_2(.din(w_dff_B_UPX9w7Ht8_2),.dout(w_dff_B_sPsAxl123_2),.clk(gclk));
	jdff dff_B_Ria118Gd0_2(.din(w_dff_B_sPsAxl123_2),.dout(w_dff_B_Ria118Gd0_2),.clk(gclk));
	jdff dff_B_PBlOLn9W3_2(.din(w_dff_B_Ria118Gd0_2),.dout(w_dff_B_PBlOLn9W3_2),.clk(gclk));
	jdff dff_B_FgdnHYwK2_1(.din(n935),.dout(w_dff_B_FgdnHYwK2_1),.clk(gclk));
	jdff dff_B_ekgEtoUO2_2(.din(n832),.dout(w_dff_B_ekgEtoUO2_2),.clk(gclk));
	jdff dff_B_sYKDkzLF9_2(.din(w_dff_B_ekgEtoUO2_2),.dout(w_dff_B_sYKDkzLF9_2),.clk(gclk));
	jdff dff_B_Tr3LEl8r5_2(.din(w_dff_B_sYKDkzLF9_2),.dout(w_dff_B_Tr3LEl8r5_2),.clk(gclk));
	jdff dff_B_zEK7cFsf1_2(.din(w_dff_B_Tr3LEl8r5_2),.dout(w_dff_B_zEK7cFsf1_2),.clk(gclk));
	jdff dff_B_GfRMrhS61_2(.din(w_dff_B_zEK7cFsf1_2),.dout(w_dff_B_GfRMrhS61_2),.clk(gclk));
	jdff dff_B_2FZCjvbg1_2(.din(w_dff_B_GfRMrhS61_2),.dout(w_dff_B_2FZCjvbg1_2),.clk(gclk));
	jdff dff_B_XlyqA1IH5_2(.din(w_dff_B_2FZCjvbg1_2),.dout(w_dff_B_XlyqA1IH5_2),.clk(gclk));
	jdff dff_B_xP8AtX5Z5_2(.din(w_dff_B_XlyqA1IH5_2),.dout(w_dff_B_xP8AtX5Z5_2),.clk(gclk));
	jdff dff_B_2yvGR2Ek1_2(.din(w_dff_B_xP8AtX5Z5_2),.dout(w_dff_B_2yvGR2Ek1_2),.clk(gclk));
	jdff dff_B_b1V6jxak8_2(.din(w_dff_B_2yvGR2Ek1_2),.dout(w_dff_B_b1V6jxak8_2),.clk(gclk));
	jdff dff_B_gN3pGbps7_2(.din(w_dff_B_b1V6jxak8_2),.dout(w_dff_B_gN3pGbps7_2),.clk(gclk));
	jdff dff_B_4BxoFDyC1_2(.din(w_dff_B_gN3pGbps7_2),.dout(w_dff_B_4BxoFDyC1_2),.clk(gclk));
	jdff dff_B_O3PoVkvw4_2(.din(w_dff_B_4BxoFDyC1_2),.dout(w_dff_B_O3PoVkvw4_2),.clk(gclk));
	jdff dff_B_TVGJSBX56_2(.din(w_dff_B_O3PoVkvw4_2),.dout(w_dff_B_TVGJSBX56_2),.clk(gclk));
	jdff dff_B_xtK5Rbih5_2(.din(w_dff_B_TVGJSBX56_2),.dout(w_dff_B_xtK5Rbih5_2),.clk(gclk));
	jdff dff_B_3nCiWTnS1_2(.din(w_dff_B_xtK5Rbih5_2),.dout(w_dff_B_3nCiWTnS1_2),.clk(gclk));
	jdff dff_B_0NtUjsPQ1_2(.din(w_dff_B_3nCiWTnS1_2),.dout(w_dff_B_0NtUjsPQ1_2),.clk(gclk));
	jdff dff_B_gjnnWyRi4_2(.din(w_dff_B_0NtUjsPQ1_2),.dout(w_dff_B_gjnnWyRi4_2),.clk(gclk));
	jdff dff_B_h3n7iEUg1_2(.din(w_dff_B_gjnnWyRi4_2),.dout(w_dff_B_h3n7iEUg1_2),.clk(gclk));
	jdff dff_B_pMhNgscN4_2(.din(w_dff_B_h3n7iEUg1_2),.dout(w_dff_B_pMhNgscN4_2),.clk(gclk));
	jdff dff_B_e0HsKxQf0_2(.din(w_dff_B_pMhNgscN4_2),.dout(w_dff_B_e0HsKxQf0_2),.clk(gclk));
	jdff dff_B_mWheOF5C7_2(.din(w_dff_B_e0HsKxQf0_2),.dout(w_dff_B_mWheOF5C7_2),.clk(gclk));
	jdff dff_B_q1b7ahO29_1(.din(n833),.dout(w_dff_B_q1b7ahO29_1),.clk(gclk));
	jdff dff_B_veTLb8Vs8_2(.din(n734),.dout(w_dff_B_veTLb8Vs8_2),.clk(gclk));
	jdff dff_B_0ahfb7oG5_2(.din(w_dff_B_veTLb8Vs8_2),.dout(w_dff_B_0ahfb7oG5_2),.clk(gclk));
	jdff dff_B_dGm8vyB83_2(.din(w_dff_B_0ahfb7oG5_2),.dout(w_dff_B_dGm8vyB83_2),.clk(gclk));
	jdff dff_B_fjUzNIqj5_2(.din(w_dff_B_dGm8vyB83_2),.dout(w_dff_B_fjUzNIqj5_2),.clk(gclk));
	jdff dff_B_EL1xu06P2_2(.din(w_dff_B_fjUzNIqj5_2),.dout(w_dff_B_EL1xu06P2_2),.clk(gclk));
	jdff dff_B_aSOYuojn0_2(.din(w_dff_B_EL1xu06P2_2),.dout(w_dff_B_aSOYuojn0_2),.clk(gclk));
	jdff dff_B_CZEOpvFt0_2(.din(w_dff_B_aSOYuojn0_2),.dout(w_dff_B_CZEOpvFt0_2),.clk(gclk));
	jdff dff_B_E8omsfOG9_2(.din(w_dff_B_CZEOpvFt0_2),.dout(w_dff_B_E8omsfOG9_2),.clk(gclk));
	jdff dff_B_18ffRcbz4_2(.din(w_dff_B_E8omsfOG9_2),.dout(w_dff_B_18ffRcbz4_2),.clk(gclk));
	jdff dff_B_uDT9w2XC3_2(.din(w_dff_B_18ffRcbz4_2),.dout(w_dff_B_uDT9w2XC3_2),.clk(gclk));
	jdff dff_B_2M3DeORd4_2(.din(w_dff_B_uDT9w2XC3_2),.dout(w_dff_B_2M3DeORd4_2),.clk(gclk));
	jdff dff_B_a0dAQvqn7_2(.din(w_dff_B_2M3DeORd4_2),.dout(w_dff_B_a0dAQvqn7_2),.clk(gclk));
	jdff dff_B_SCiFj1xc9_2(.din(w_dff_B_a0dAQvqn7_2),.dout(w_dff_B_SCiFj1xc9_2),.clk(gclk));
	jdff dff_B_C36nM2X15_2(.din(w_dff_B_SCiFj1xc9_2),.dout(w_dff_B_C36nM2X15_2),.clk(gclk));
	jdff dff_B_NBsocNKy7_2(.din(w_dff_B_C36nM2X15_2),.dout(w_dff_B_NBsocNKy7_2),.clk(gclk));
	jdff dff_B_8xdLxR9I9_2(.din(w_dff_B_NBsocNKy7_2),.dout(w_dff_B_8xdLxR9I9_2),.clk(gclk));
	jdff dff_B_iP887MlT9_2(.din(w_dff_B_8xdLxR9I9_2),.dout(w_dff_B_iP887MlT9_2),.clk(gclk));
	jdff dff_B_3500toN99_2(.din(w_dff_B_iP887MlT9_2),.dout(w_dff_B_3500toN99_2),.clk(gclk));
	jdff dff_B_4ShIlRBK3_2(.din(w_dff_B_3500toN99_2),.dout(w_dff_B_4ShIlRBK3_2),.clk(gclk));
	jdff dff_B_vZt4kRgy3_2(.din(w_dff_B_4ShIlRBK3_2),.dout(w_dff_B_vZt4kRgy3_2),.clk(gclk));
	jdff dff_B_LVoVRGms8_1(.din(n735),.dout(w_dff_B_LVoVRGms8_1),.clk(gclk));
	jdff dff_B_ClMo1ysm3_2(.din(n642),.dout(w_dff_B_ClMo1ysm3_2),.clk(gclk));
	jdff dff_B_uwuJcj5Z0_2(.din(w_dff_B_ClMo1ysm3_2),.dout(w_dff_B_uwuJcj5Z0_2),.clk(gclk));
	jdff dff_B_r6WN8Ujm1_2(.din(w_dff_B_uwuJcj5Z0_2),.dout(w_dff_B_r6WN8Ujm1_2),.clk(gclk));
	jdff dff_B_q8VNmquh5_2(.din(w_dff_B_r6WN8Ujm1_2),.dout(w_dff_B_q8VNmquh5_2),.clk(gclk));
	jdff dff_B_umMJzL4H4_2(.din(w_dff_B_q8VNmquh5_2),.dout(w_dff_B_umMJzL4H4_2),.clk(gclk));
	jdff dff_B_qycJlDXy4_2(.din(w_dff_B_umMJzL4H4_2),.dout(w_dff_B_qycJlDXy4_2),.clk(gclk));
	jdff dff_B_8PxiXb4f7_2(.din(w_dff_B_qycJlDXy4_2),.dout(w_dff_B_8PxiXb4f7_2),.clk(gclk));
	jdff dff_B_XELB2PkE5_2(.din(w_dff_B_8PxiXb4f7_2),.dout(w_dff_B_XELB2PkE5_2),.clk(gclk));
	jdff dff_B_1OP0kEfm1_2(.din(w_dff_B_XELB2PkE5_2),.dout(w_dff_B_1OP0kEfm1_2),.clk(gclk));
	jdff dff_B_l2VlOEbG5_2(.din(w_dff_B_1OP0kEfm1_2),.dout(w_dff_B_l2VlOEbG5_2),.clk(gclk));
	jdff dff_B_JE0GkGB96_2(.din(w_dff_B_l2VlOEbG5_2),.dout(w_dff_B_JE0GkGB96_2),.clk(gclk));
	jdff dff_B_DwyTfFK09_2(.din(w_dff_B_JE0GkGB96_2),.dout(w_dff_B_DwyTfFK09_2),.clk(gclk));
	jdff dff_B_pxSpR05y1_2(.din(w_dff_B_DwyTfFK09_2),.dout(w_dff_B_pxSpR05y1_2),.clk(gclk));
	jdff dff_B_IN0dtKW29_2(.din(w_dff_B_pxSpR05y1_2),.dout(w_dff_B_IN0dtKW29_2),.clk(gclk));
	jdff dff_B_dm9LOI3q5_2(.din(w_dff_B_IN0dtKW29_2),.dout(w_dff_B_dm9LOI3q5_2),.clk(gclk));
	jdff dff_B_i7FjBT1X6_2(.din(w_dff_B_dm9LOI3q5_2),.dout(w_dff_B_i7FjBT1X6_2),.clk(gclk));
	jdff dff_B_ZNGfFnnu0_2(.din(w_dff_B_i7FjBT1X6_2),.dout(w_dff_B_ZNGfFnnu0_2),.clk(gclk));
	jdff dff_B_KJsm2iQ82_2(.din(w_dff_B_ZNGfFnnu0_2),.dout(w_dff_B_KJsm2iQ82_2),.clk(gclk));
	jdff dff_B_4XFcQDTb2_1(.din(n643),.dout(w_dff_B_4XFcQDTb2_1),.clk(gclk));
	jdff dff_B_akRh96m98_2(.din(n557),.dout(w_dff_B_akRh96m98_2),.clk(gclk));
	jdff dff_B_o3Hb8qRl9_2(.din(w_dff_B_akRh96m98_2),.dout(w_dff_B_o3Hb8qRl9_2),.clk(gclk));
	jdff dff_B_MdL5x2Um9_2(.din(w_dff_B_o3Hb8qRl9_2),.dout(w_dff_B_MdL5x2Um9_2),.clk(gclk));
	jdff dff_B_iIuAZHJe0_2(.din(w_dff_B_MdL5x2Um9_2),.dout(w_dff_B_iIuAZHJe0_2),.clk(gclk));
	jdff dff_B_8nc1XJGJ6_2(.din(w_dff_B_iIuAZHJe0_2),.dout(w_dff_B_8nc1XJGJ6_2),.clk(gclk));
	jdff dff_B_PW6VcZAH8_2(.din(w_dff_B_8nc1XJGJ6_2),.dout(w_dff_B_PW6VcZAH8_2),.clk(gclk));
	jdff dff_B_wXTODCum4_2(.din(w_dff_B_PW6VcZAH8_2),.dout(w_dff_B_wXTODCum4_2),.clk(gclk));
	jdff dff_B_lT0uklDO9_2(.din(w_dff_B_wXTODCum4_2),.dout(w_dff_B_lT0uklDO9_2),.clk(gclk));
	jdff dff_B_aVXoJ7u48_2(.din(w_dff_B_lT0uklDO9_2),.dout(w_dff_B_aVXoJ7u48_2),.clk(gclk));
	jdff dff_B_VFC9A23N0_2(.din(w_dff_B_aVXoJ7u48_2),.dout(w_dff_B_VFC9A23N0_2),.clk(gclk));
	jdff dff_B_T7RaTU3C0_2(.din(w_dff_B_VFC9A23N0_2),.dout(w_dff_B_T7RaTU3C0_2),.clk(gclk));
	jdff dff_B_t8m4j8xr8_2(.din(w_dff_B_T7RaTU3C0_2),.dout(w_dff_B_t8m4j8xr8_2),.clk(gclk));
	jdff dff_B_Z4wJxIY12_2(.din(w_dff_B_t8m4j8xr8_2),.dout(w_dff_B_Z4wJxIY12_2),.clk(gclk));
	jdff dff_B_rruH8tJ20_2(.din(w_dff_B_Z4wJxIY12_2),.dout(w_dff_B_rruH8tJ20_2),.clk(gclk));
	jdff dff_B_3zrRElB43_2(.din(w_dff_B_rruH8tJ20_2),.dout(w_dff_B_3zrRElB43_2),.clk(gclk));
	jdff dff_B_xLVoL2A89_2(.din(w_dff_B_3zrRElB43_2),.dout(w_dff_B_xLVoL2A89_2),.clk(gclk));
	jdff dff_B_EeRAn82r9_1(.din(n558),.dout(w_dff_B_EeRAn82r9_1),.clk(gclk));
	jdff dff_B_7AI4Njhh6_2(.din(n479),.dout(w_dff_B_7AI4Njhh6_2),.clk(gclk));
	jdff dff_B_CREJbewt6_2(.din(w_dff_B_7AI4Njhh6_2),.dout(w_dff_B_CREJbewt6_2),.clk(gclk));
	jdff dff_B_aDc2gZMo1_2(.din(w_dff_B_CREJbewt6_2),.dout(w_dff_B_aDc2gZMo1_2),.clk(gclk));
	jdff dff_B_XGxtZviB5_2(.din(w_dff_B_aDc2gZMo1_2),.dout(w_dff_B_XGxtZviB5_2),.clk(gclk));
	jdff dff_B_YZDPIdx77_2(.din(w_dff_B_XGxtZviB5_2),.dout(w_dff_B_YZDPIdx77_2),.clk(gclk));
	jdff dff_B_qoXoW2Br7_2(.din(w_dff_B_YZDPIdx77_2),.dout(w_dff_B_qoXoW2Br7_2),.clk(gclk));
	jdff dff_B_nbGLUgVs8_2(.din(w_dff_B_qoXoW2Br7_2),.dout(w_dff_B_nbGLUgVs8_2),.clk(gclk));
	jdff dff_B_dvJqJAoi4_2(.din(w_dff_B_nbGLUgVs8_2),.dout(w_dff_B_dvJqJAoi4_2),.clk(gclk));
	jdff dff_B_O9G2zr9x4_2(.din(w_dff_B_dvJqJAoi4_2),.dout(w_dff_B_O9G2zr9x4_2),.clk(gclk));
	jdff dff_B_QMQyzwLw5_2(.din(w_dff_B_O9G2zr9x4_2),.dout(w_dff_B_QMQyzwLw5_2),.clk(gclk));
	jdff dff_B_2VWYOpj38_2(.din(w_dff_B_QMQyzwLw5_2),.dout(w_dff_B_2VWYOpj38_2),.clk(gclk));
	jdff dff_B_Z1cr4aXq6_2(.din(w_dff_B_2VWYOpj38_2),.dout(w_dff_B_Z1cr4aXq6_2),.clk(gclk));
	jdff dff_B_JJeV97Np3_2(.din(w_dff_B_Z1cr4aXq6_2),.dout(w_dff_B_JJeV97Np3_2),.clk(gclk));
	jdff dff_B_tm99xvrP5_2(.din(w_dff_B_JJeV97Np3_2),.dout(w_dff_B_tm99xvrP5_2),.clk(gclk));
	jdff dff_B_t8UKOF9J6_1(.din(n480),.dout(w_dff_B_t8UKOF9J6_1),.clk(gclk));
	jdff dff_B_vmfqcjdR1_2(.din(n408),.dout(w_dff_B_vmfqcjdR1_2),.clk(gclk));
	jdff dff_B_zuHONWuS5_2(.din(w_dff_B_vmfqcjdR1_2),.dout(w_dff_B_zuHONWuS5_2),.clk(gclk));
	jdff dff_B_Y8Ptgm9C0_2(.din(w_dff_B_zuHONWuS5_2),.dout(w_dff_B_Y8Ptgm9C0_2),.clk(gclk));
	jdff dff_B_7CQ2v9EO7_2(.din(w_dff_B_Y8Ptgm9C0_2),.dout(w_dff_B_7CQ2v9EO7_2),.clk(gclk));
	jdff dff_B_NLty3pQN6_2(.din(w_dff_B_7CQ2v9EO7_2),.dout(w_dff_B_NLty3pQN6_2),.clk(gclk));
	jdff dff_B_D8wmpClN2_2(.din(w_dff_B_NLty3pQN6_2),.dout(w_dff_B_D8wmpClN2_2),.clk(gclk));
	jdff dff_B_qJWLIZBO5_2(.din(w_dff_B_D8wmpClN2_2),.dout(w_dff_B_qJWLIZBO5_2),.clk(gclk));
	jdff dff_B_AuvRTLi49_2(.din(w_dff_B_qJWLIZBO5_2),.dout(w_dff_B_AuvRTLi49_2),.clk(gclk));
	jdff dff_B_wKwhIiQR9_2(.din(w_dff_B_AuvRTLi49_2),.dout(w_dff_B_wKwhIiQR9_2),.clk(gclk));
	jdff dff_B_6LQjZsdB1_2(.din(w_dff_B_wKwhIiQR9_2),.dout(w_dff_B_6LQjZsdB1_2),.clk(gclk));
	jdff dff_B_Kj84ly7A4_2(.din(w_dff_B_6LQjZsdB1_2),.dout(w_dff_B_Kj84ly7A4_2),.clk(gclk));
	jdff dff_B_n8pcLXAT9_2(.din(w_dff_B_Kj84ly7A4_2),.dout(w_dff_B_n8pcLXAT9_2),.clk(gclk));
	jdff dff_B_QovX8Hk43_2(.din(n411),.dout(w_dff_B_QovX8Hk43_2),.clk(gclk));
	jdff dff_B_GqB6oQRN9_2(.din(w_dff_B_QovX8Hk43_2),.dout(w_dff_B_GqB6oQRN9_2),.clk(gclk));
	jdff dff_B_yFFnSilg5_2(.din(w_dff_B_GqB6oQRN9_2),.dout(w_dff_B_yFFnSilg5_2),.clk(gclk));
	jdff dff_B_FvN6rCQc2_1(.din(n409),.dout(w_dff_B_FvN6rCQc2_1),.clk(gclk));
	jdff dff_B_cJDKDu5i9_2(.din(n345),.dout(w_dff_B_cJDKDu5i9_2),.clk(gclk));
	jdff dff_B_N14UW4li6_2(.din(w_dff_B_cJDKDu5i9_2),.dout(w_dff_B_N14UW4li6_2),.clk(gclk));
	jdff dff_B_3tCyqfK11_2(.din(w_dff_B_N14UW4li6_2),.dout(w_dff_B_3tCyqfK11_2),.clk(gclk));
	jdff dff_B_v594jcT89_2(.din(w_dff_B_3tCyqfK11_2),.dout(w_dff_B_v594jcT89_2),.clk(gclk));
	jdff dff_B_jqC0T3Ib6_2(.din(w_dff_B_v594jcT89_2),.dout(w_dff_B_jqC0T3Ib6_2),.clk(gclk));
	jdff dff_B_ESlMcoRT9_2(.din(w_dff_B_jqC0T3Ib6_2),.dout(w_dff_B_ESlMcoRT9_2),.clk(gclk));
	jdff dff_B_teCrdQ8K5_2(.din(w_dff_B_ESlMcoRT9_2),.dout(w_dff_B_teCrdQ8K5_2),.clk(gclk));
	jdff dff_B_JkEj9UbZ8_1(.din(n346),.dout(w_dff_B_JkEj9UbZ8_1),.clk(gclk));
	jdff dff_B_i9xW1p9e3_2(.din(n289),.dout(w_dff_B_i9xW1p9e3_2),.clk(gclk));
	jdff dff_B_ZU1jIcRx3_2(.din(w_dff_B_i9xW1p9e3_2),.dout(w_dff_B_ZU1jIcRx3_2),.clk(gclk));
	jdff dff_B_Pxtf12Fd3_2(.din(w_dff_B_ZU1jIcRx3_2),.dout(w_dff_B_Pxtf12Fd3_2),.clk(gclk));
	jdff dff_B_9JcfT8IA9_2(.din(w_dff_B_Pxtf12Fd3_2),.dout(w_dff_B_9JcfT8IA9_2),.clk(gclk));
	jdff dff_B_ZXoeUWOj6_2(.din(w_dff_B_9JcfT8IA9_2),.dout(w_dff_B_ZXoeUWOj6_2),.clk(gclk));
	jdff dff_B_7uz8IcC05_1(.din(n291),.dout(w_dff_B_7uz8IcC05_1),.clk(gclk));
	jdff dff_B_YGy5Ezsl9_2(.din(n241),.dout(w_dff_B_YGy5Ezsl9_2),.clk(gclk));
	jdff dff_B_x7IpbgK77_2(.din(w_dff_B_YGy5Ezsl9_2),.dout(w_dff_B_x7IpbgK77_2),.clk(gclk));
	jdff dff_B_IBrwA5D33_2(.din(w_dff_B_x7IpbgK77_2),.dout(w_dff_B_IBrwA5D33_2),.clk(gclk));
	jdff dff_B_wZMqDuih9_0(.din(n246),.dout(w_dff_B_wZMqDuih9_0),.clk(gclk));
	jdff dff_B_VTHvwSX19_0(.din(w_dff_B_wZMqDuih9_0),.dout(w_dff_B_VTHvwSX19_0),.clk(gclk));
	jdff dff_A_retMBguq4_0(.dout(w_n196_0[0]),.din(w_dff_A_retMBguq4_0),.clk(gclk));
	jdff dff_A_hY78nFfS1_0(.dout(w_dff_A_retMBguq4_0),.din(w_dff_A_hY78nFfS1_0),.clk(gclk));
	jdff dff_A_xMoJ7StT8_1(.dout(w_n196_0[1]),.din(w_dff_A_xMoJ7StT8_1),.clk(gclk));
	jdff dff_A_TMMq93Z77_1(.dout(w_dff_A_xMoJ7StT8_1),.din(w_dff_A_TMMq93Z77_1),.clk(gclk));
	jdff dff_B_hU1vr8NB2_2(.din(n1465),.dout(w_dff_B_hU1vr8NB2_2),.clk(gclk));
	jdff dff_B_w0qqjdMw7_2(.din(w_dff_B_hU1vr8NB2_2),.dout(w_dff_B_w0qqjdMw7_2),.clk(gclk));
	jdff dff_B_GKM8K4XL9_1(.din(n1463),.dout(w_dff_B_GKM8K4XL9_1),.clk(gclk));
	jdff dff_B_maUi0Lzd7_2(.din(n1390),.dout(w_dff_B_maUi0Lzd7_2),.clk(gclk));
	jdff dff_B_CxSPndrc1_2(.din(w_dff_B_maUi0Lzd7_2),.dout(w_dff_B_CxSPndrc1_2),.clk(gclk));
	jdff dff_B_MhLCBSzF3_2(.din(w_dff_B_CxSPndrc1_2),.dout(w_dff_B_MhLCBSzF3_2),.clk(gclk));
	jdff dff_B_a3dxtBr67_2(.din(w_dff_B_MhLCBSzF3_2),.dout(w_dff_B_a3dxtBr67_2),.clk(gclk));
	jdff dff_B_8iSvPxTB5_2(.din(w_dff_B_a3dxtBr67_2),.dout(w_dff_B_8iSvPxTB5_2),.clk(gclk));
	jdff dff_B_Ke6b32sX7_2(.din(w_dff_B_8iSvPxTB5_2),.dout(w_dff_B_Ke6b32sX7_2),.clk(gclk));
	jdff dff_B_1ExOcTyq1_2(.din(w_dff_B_Ke6b32sX7_2),.dout(w_dff_B_1ExOcTyq1_2),.clk(gclk));
	jdff dff_B_lgF1Qhfv7_2(.din(w_dff_B_1ExOcTyq1_2),.dout(w_dff_B_lgF1Qhfv7_2),.clk(gclk));
	jdff dff_B_CGgVJdRW9_2(.din(w_dff_B_lgF1Qhfv7_2),.dout(w_dff_B_CGgVJdRW9_2),.clk(gclk));
	jdff dff_B_PC55rC5Q2_2(.din(w_dff_B_CGgVJdRW9_2),.dout(w_dff_B_PC55rC5Q2_2),.clk(gclk));
	jdff dff_B_laNg1s5u2_2(.din(w_dff_B_PC55rC5Q2_2),.dout(w_dff_B_laNg1s5u2_2),.clk(gclk));
	jdff dff_B_ek8eaccx1_2(.din(w_dff_B_laNg1s5u2_2),.dout(w_dff_B_ek8eaccx1_2),.clk(gclk));
	jdff dff_B_0boWsVUu9_2(.din(w_dff_B_ek8eaccx1_2),.dout(w_dff_B_0boWsVUu9_2),.clk(gclk));
	jdff dff_B_ifydVLx50_2(.din(w_dff_B_0boWsVUu9_2),.dout(w_dff_B_ifydVLx50_2),.clk(gclk));
	jdff dff_B_bn7Bp5YP4_2(.din(w_dff_B_ifydVLx50_2),.dout(w_dff_B_bn7Bp5YP4_2),.clk(gclk));
	jdff dff_B_IXmGDbx54_2(.din(w_dff_B_bn7Bp5YP4_2),.dout(w_dff_B_IXmGDbx54_2),.clk(gclk));
	jdff dff_B_5xAWax9B8_2(.din(w_dff_B_IXmGDbx54_2),.dout(w_dff_B_5xAWax9B8_2),.clk(gclk));
	jdff dff_B_KYHpEjRR4_2(.din(w_dff_B_5xAWax9B8_2),.dout(w_dff_B_KYHpEjRR4_2),.clk(gclk));
	jdff dff_B_v8rEyMCD7_2(.din(w_dff_B_KYHpEjRR4_2),.dout(w_dff_B_v8rEyMCD7_2),.clk(gclk));
	jdff dff_B_wZvVc4L84_2(.din(w_dff_B_v8rEyMCD7_2),.dout(w_dff_B_wZvVc4L84_2),.clk(gclk));
	jdff dff_B_3p9SAWRY2_2(.din(w_dff_B_wZvVc4L84_2),.dout(w_dff_B_3p9SAWRY2_2),.clk(gclk));
	jdff dff_B_44dBfwXj8_2(.din(w_dff_B_3p9SAWRY2_2),.dout(w_dff_B_44dBfwXj8_2),.clk(gclk));
	jdff dff_B_eILm0Hdd1_2(.din(w_dff_B_44dBfwXj8_2),.dout(w_dff_B_eILm0Hdd1_2),.clk(gclk));
	jdff dff_B_SRB1jn3r4_2(.din(w_dff_B_eILm0Hdd1_2),.dout(w_dff_B_SRB1jn3r4_2),.clk(gclk));
	jdff dff_B_aMk3RGb47_2(.din(w_dff_B_SRB1jn3r4_2),.dout(w_dff_B_aMk3RGb47_2),.clk(gclk));
	jdff dff_B_XIZvnHZf6_2(.din(w_dff_B_aMk3RGb47_2),.dout(w_dff_B_XIZvnHZf6_2),.clk(gclk));
	jdff dff_B_1Bf0ttZE9_2(.din(w_dff_B_XIZvnHZf6_2),.dout(w_dff_B_1Bf0ttZE9_2),.clk(gclk));
	jdff dff_B_mMW3aN4X6_2(.din(w_dff_B_1Bf0ttZE9_2),.dout(w_dff_B_mMW3aN4X6_2),.clk(gclk));
	jdff dff_B_X85fratI2_2(.din(w_dff_B_mMW3aN4X6_2),.dout(w_dff_B_X85fratI2_2),.clk(gclk));
	jdff dff_B_cqtq7KrZ3_2(.din(w_dff_B_X85fratI2_2),.dout(w_dff_B_cqtq7KrZ3_2),.clk(gclk));
	jdff dff_B_qkPFyqNd2_2(.din(w_dff_B_cqtq7KrZ3_2),.dout(w_dff_B_qkPFyqNd2_2),.clk(gclk));
	jdff dff_B_uFiUg5zk1_2(.din(w_dff_B_qkPFyqNd2_2),.dout(w_dff_B_uFiUg5zk1_2),.clk(gclk));
	jdff dff_B_qQayyI4N9_2(.din(w_dff_B_uFiUg5zk1_2),.dout(w_dff_B_qQayyI4N9_2),.clk(gclk));
	jdff dff_B_aSVJu1OY1_2(.din(w_dff_B_qQayyI4N9_2),.dout(w_dff_B_aSVJu1OY1_2),.clk(gclk));
	jdff dff_B_PX4TXQFr3_2(.din(w_dff_B_aSVJu1OY1_2),.dout(w_dff_B_PX4TXQFr3_2),.clk(gclk));
	jdff dff_B_wYs9wv6H6_1(.din(n1461),.dout(w_dff_B_wYs9wv6H6_1),.clk(gclk));
	jdff dff_A_cnLtIaDT5_1(.dout(w_n1393_0[1]),.din(w_dff_A_cnLtIaDT5_1),.clk(gclk));
	jdff dff_B_7bDJzS977_1(.din(n1391),.dout(w_dff_B_7bDJzS977_1),.clk(gclk));
	jdff dff_B_wA5Gw0z84_2(.din(n1312),.dout(w_dff_B_wA5Gw0z84_2),.clk(gclk));
	jdff dff_B_tMRehM009_2(.din(w_dff_B_wA5Gw0z84_2),.dout(w_dff_B_tMRehM009_2),.clk(gclk));
	jdff dff_B_QPVHrLSu8_2(.din(w_dff_B_tMRehM009_2),.dout(w_dff_B_QPVHrLSu8_2),.clk(gclk));
	jdff dff_B_poLOfYC04_2(.din(w_dff_B_QPVHrLSu8_2),.dout(w_dff_B_poLOfYC04_2),.clk(gclk));
	jdff dff_B_0TgQrXSf8_2(.din(w_dff_B_poLOfYC04_2),.dout(w_dff_B_0TgQrXSf8_2),.clk(gclk));
	jdff dff_B_WSVDKpfw1_2(.din(w_dff_B_0TgQrXSf8_2),.dout(w_dff_B_WSVDKpfw1_2),.clk(gclk));
	jdff dff_B_pAB45IqW3_2(.din(w_dff_B_WSVDKpfw1_2),.dout(w_dff_B_pAB45IqW3_2),.clk(gclk));
	jdff dff_B_DSXpFfIh4_2(.din(w_dff_B_pAB45IqW3_2),.dout(w_dff_B_DSXpFfIh4_2),.clk(gclk));
	jdff dff_B_TcuTRza81_2(.din(w_dff_B_DSXpFfIh4_2),.dout(w_dff_B_TcuTRza81_2),.clk(gclk));
	jdff dff_B_8aLhlURf9_2(.din(w_dff_B_TcuTRza81_2),.dout(w_dff_B_8aLhlURf9_2),.clk(gclk));
	jdff dff_B_D7hHXQoh1_2(.din(w_dff_B_8aLhlURf9_2),.dout(w_dff_B_D7hHXQoh1_2),.clk(gclk));
	jdff dff_B_Xv3tLuEo5_2(.din(w_dff_B_D7hHXQoh1_2),.dout(w_dff_B_Xv3tLuEo5_2),.clk(gclk));
	jdff dff_B_orABP4fh7_2(.din(w_dff_B_Xv3tLuEo5_2),.dout(w_dff_B_orABP4fh7_2),.clk(gclk));
	jdff dff_B_c9uSD6N01_2(.din(w_dff_B_orABP4fh7_2),.dout(w_dff_B_c9uSD6N01_2),.clk(gclk));
	jdff dff_B_sdaqmCrV9_2(.din(w_dff_B_c9uSD6N01_2),.dout(w_dff_B_sdaqmCrV9_2),.clk(gclk));
	jdff dff_B_pCkqAd235_2(.din(w_dff_B_sdaqmCrV9_2),.dout(w_dff_B_pCkqAd235_2),.clk(gclk));
	jdff dff_B_yUGJ1ABx7_2(.din(w_dff_B_pCkqAd235_2),.dout(w_dff_B_yUGJ1ABx7_2),.clk(gclk));
	jdff dff_B_fHjw4xR85_2(.din(w_dff_B_yUGJ1ABx7_2),.dout(w_dff_B_fHjw4xR85_2),.clk(gclk));
	jdff dff_B_G9DlWunn7_2(.din(w_dff_B_fHjw4xR85_2),.dout(w_dff_B_G9DlWunn7_2),.clk(gclk));
	jdff dff_B_8ENxcvDx1_2(.din(w_dff_B_G9DlWunn7_2),.dout(w_dff_B_8ENxcvDx1_2),.clk(gclk));
	jdff dff_B_UCLLO6K79_2(.din(w_dff_B_8ENxcvDx1_2),.dout(w_dff_B_UCLLO6K79_2),.clk(gclk));
	jdff dff_B_F7Dp79Zo8_2(.din(w_dff_B_UCLLO6K79_2),.dout(w_dff_B_F7Dp79Zo8_2),.clk(gclk));
	jdff dff_B_Mk1Rz2mV3_2(.din(w_dff_B_F7Dp79Zo8_2),.dout(w_dff_B_Mk1Rz2mV3_2),.clk(gclk));
	jdff dff_B_4cB1IIUp4_2(.din(w_dff_B_Mk1Rz2mV3_2),.dout(w_dff_B_4cB1IIUp4_2),.clk(gclk));
	jdff dff_B_V0wGUUrE2_2(.din(w_dff_B_4cB1IIUp4_2),.dout(w_dff_B_V0wGUUrE2_2),.clk(gclk));
	jdff dff_B_1DWqglps3_2(.din(w_dff_B_V0wGUUrE2_2),.dout(w_dff_B_1DWqglps3_2),.clk(gclk));
	jdff dff_B_NBvfBKSV9_2(.din(w_dff_B_1DWqglps3_2),.dout(w_dff_B_NBvfBKSV9_2),.clk(gclk));
	jdff dff_B_Vl22xVyp0_2(.din(w_dff_B_NBvfBKSV9_2),.dout(w_dff_B_Vl22xVyp0_2),.clk(gclk));
	jdff dff_B_nE2JIBPd8_2(.din(w_dff_B_Vl22xVyp0_2),.dout(w_dff_B_nE2JIBPd8_2),.clk(gclk));
	jdff dff_B_Mmu3qViy6_2(.din(w_dff_B_nE2JIBPd8_2),.dout(w_dff_B_Mmu3qViy6_2),.clk(gclk));
	jdff dff_B_RaRq5BB64_1(.din(n1313),.dout(w_dff_B_RaRq5BB64_1),.clk(gclk));
	jdff dff_B_jKS1znAl9_2(.din(n1227),.dout(w_dff_B_jKS1znAl9_2),.clk(gclk));
	jdff dff_B_IEldEdry3_2(.din(w_dff_B_jKS1znAl9_2),.dout(w_dff_B_IEldEdry3_2),.clk(gclk));
	jdff dff_B_Wj2RZUHn7_2(.din(w_dff_B_IEldEdry3_2),.dout(w_dff_B_Wj2RZUHn7_2),.clk(gclk));
	jdff dff_B_QOutNQxk7_2(.din(w_dff_B_Wj2RZUHn7_2),.dout(w_dff_B_QOutNQxk7_2),.clk(gclk));
	jdff dff_B_qgEb6KPh5_2(.din(w_dff_B_QOutNQxk7_2),.dout(w_dff_B_qgEb6KPh5_2),.clk(gclk));
	jdff dff_B_enKxK3UM9_2(.din(w_dff_B_qgEb6KPh5_2),.dout(w_dff_B_enKxK3UM9_2),.clk(gclk));
	jdff dff_B_8shtw70R2_2(.din(w_dff_B_enKxK3UM9_2),.dout(w_dff_B_8shtw70R2_2),.clk(gclk));
	jdff dff_B_7fEHJGDL2_2(.din(w_dff_B_8shtw70R2_2),.dout(w_dff_B_7fEHJGDL2_2),.clk(gclk));
	jdff dff_B_qL08NAw01_2(.din(w_dff_B_7fEHJGDL2_2),.dout(w_dff_B_qL08NAw01_2),.clk(gclk));
	jdff dff_B_lT2NR7956_2(.din(w_dff_B_qL08NAw01_2),.dout(w_dff_B_lT2NR7956_2),.clk(gclk));
	jdff dff_B_H7hFTxHI7_2(.din(w_dff_B_lT2NR7956_2),.dout(w_dff_B_H7hFTxHI7_2),.clk(gclk));
	jdff dff_B_3KgJDtrk7_2(.din(w_dff_B_H7hFTxHI7_2),.dout(w_dff_B_3KgJDtrk7_2),.clk(gclk));
	jdff dff_B_ei8Sv0aK9_2(.din(w_dff_B_3KgJDtrk7_2),.dout(w_dff_B_ei8Sv0aK9_2),.clk(gclk));
	jdff dff_B_jLu3wO3D8_2(.din(w_dff_B_ei8Sv0aK9_2),.dout(w_dff_B_jLu3wO3D8_2),.clk(gclk));
	jdff dff_B_88Jx1Ykp3_2(.din(w_dff_B_jLu3wO3D8_2),.dout(w_dff_B_88Jx1Ykp3_2),.clk(gclk));
	jdff dff_B_wvY57nQ62_2(.din(w_dff_B_88Jx1Ykp3_2),.dout(w_dff_B_wvY57nQ62_2),.clk(gclk));
	jdff dff_B_f5sIsrsv0_2(.din(w_dff_B_wvY57nQ62_2),.dout(w_dff_B_f5sIsrsv0_2),.clk(gclk));
	jdff dff_B_QWY6R8Vv9_2(.din(w_dff_B_f5sIsrsv0_2),.dout(w_dff_B_QWY6R8Vv9_2),.clk(gclk));
	jdff dff_B_iWuvyW2L8_2(.din(w_dff_B_QWY6R8Vv9_2),.dout(w_dff_B_iWuvyW2L8_2),.clk(gclk));
	jdff dff_B_NtXmSGFY4_2(.din(w_dff_B_iWuvyW2L8_2),.dout(w_dff_B_NtXmSGFY4_2),.clk(gclk));
	jdff dff_B_mqC9gCbc5_2(.din(w_dff_B_NtXmSGFY4_2),.dout(w_dff_B_mqC9gCbc5_2),.clk(gclk));
	jdff dff_B_AJzHeA9K2_2(.din(w_dff_B_mqC9gCbc5_2),.dout(w_dff_B_AJzHeA9K2_2),.clk(gclk));
	jdff dff_B_MsKbgqrm1_2(.din(w_dff_B_AJzHeA9K2_2),.dout(w_dff_B_MsKbgqrm1_2),.clk(gclk));
	jdff dff_B_kWsbnAtx5_2(.din(w_dff_B_MsKbgqrm1_2),.dout(w_dff_B_kWsbnAtx5_2),.clk(gclk));
	jdff dff_B_jOB8gM1P1_2(.din(w_dff_B_kWsbnAtx5_2),.dout(w_dff_B_jOB8gM1P1_2),.clk(gclk));
	jdff dff_B_t5TkYjdu0_2(.din(w_dff_B_jOB8gM1P1_2),.dout(w_dff_B_t5TkYjdu0_2),.clk(gclk));
	jdff dff_B_u2C2UcnT0_2(.din(w_dff_B_t5TkYjdu0_2),.dout(w_dff_B_u2C2UcnT0_2),.clk(gclk));
	jdff dff_B_aNHEh6ZZ6_2(.din(w_dff_B_u2C2UcnT0_2),.dout(w_dff_B_aNHEh6ZZ6_2),.clk(gclk));
	jdff dff_B_Bd7910S22_1(.din(n1228),.dout(w_dff_B_Bd7910S22_1),.clk(gclk));
	jdff dff_B_rrQgZzuG4_2(.din(n1136),.dout(w_dff_B_rrQgZzuG4_2),.clk(gclk));
	jdff dff_B_pNIrZEG52_2(.din(w_dff_B_rrQgZzuG4_2),.dout(w_dff_B_pNIrZEG52_2),.clk(gclk));
	jdff dff_B_LmDPB5aO5_2(.din(w_dff_B_pNIrZEG52_2),.dout(w_dff_B_LmDPB5aO5_2),.clk(gclk));
	jdff dff_B_l5cg6R4B3_2(.din(w_dff_B_LmDPB5aO5_2),.dout(w_dff_B_l5cg6R4B3_2),.clk(gclk));
	jdff dff_B_zEAcGAwa4_2(.din(w_dff_B_l5cg6R4B3_2),.dout(w_dff_B_zEAcGAwa4_2),.clk(gclk));
	jdff dff_B_EupCZzFA2_2(.din(w_dff_B_zEAcGAwa4_2),.dout(w_dff_B_EupCZzFA2_2),.clk(gclk));
	jdff dff_B_bQA6PJ652_2(.din(w_dff_B_EupCZzFA2_2),.dout(w_dff_B_bQA6PJ652_2),.clk(gclk));
	jdff dff_B_szrSiuWW1_2(.din(w_dff_B_bQA6PJ652_2),.dout(w_dff_B_szrSiuWW1_2),.clk(gclk));
	jdff dff_B_CGZlUZlS5_2(.din(w_dff_B_szrSiuWW1_2),.dout(w_dff_B_CGZlUZlS5_2),.clk(gclk));
	jdff dff_B_HWsTwFSJ4_2(.din(w_dff_B_CGZlUZlS5_2),.dout(w_dff_B_HWsTwFSJ4_2),.clk(gclk));
	jdff dff_B_h4WKwM6k2_2(.din(w_dff_B_HWsTwFSJ4_2),.dout(w_dff_B_h4WKwM6k2_2),.clk(gclk));
	jdff dff_B_QgBNUGeA0_2(.din(w_dff_B_h4WKwM6k2_2),.dout(w_dff_B_QgBNUGeA0_2),.clk(gclk));
	jdff dff_B_SFD9oYE37_2(.din(w_dff_B_QgBNUGeA0_2),.dout(w_dff_B_SFD9oYE37_2),.clk(gclk));
	jdff dff_B_8Zvk0iYL0_2(.din(w_dff_B_SFD9oYE37_2),.dout(w_dff_B_8Zvk0iYL0_2),.clk(gclk));
	jdff dff_B_zfekEoYl2_2(.din(w_dff_B_8Zvk0iYL0_2),.dout(w_dff_B_zfekEoYl2_2),.clk(gclk));
	jdff dff_B_HVBRvyDV0_2(.din(w_dff_B_zfekEoYl2_2),.dout(w_dff_B_HVBRvyDV0_2),.clk(gclk));
	jdff dff_B_XeOabcEj5_2(.din(w_dff_B_HVBRvyDV0_2),.dout(w_dff_B_XeOabcEj5_2),.clk(gclk));
	jdff dff_B_xFfop47F0_2(.din(w_dff_B_XeOabcEj5_2),.dout(w_dff_B_xFfop47F0_2),.clk(gclk));
	jdff dff_B_Pnt7yk0J9_2(.din(w_dff_B_xFfop47F0_2),.dout(w_dff_B_Pnt7yk0J9_2),.clk(gclk));
	jdff dff_B_7IzkV9ix1_2(.din(w_dff_B_Pnt7yk0J9_2),.dout(w_dff_B_7IzkV9ix1_2),.clk(gclk));
	jdff dff_B_7ClHIuDo8_2(.din(w_dff_B_7IzkV9ix1_2),.dout(w_dff_B_7ClHIuDo8_2),.clk(gclk));
	jdff dff_B_bEO3POAo6_2(.din(w_dff_B_7ClHIuDo8_2),.dout(w_dff_B_bEO3POAo6_2),.clk(gclk));
	jdff dff_B_Y9AFkIhl3_2(.din(w_dff_B_bEO3POAo6_2),.dout(w_dff_B_Y9AFkIhl3_2),.clk(gclk));
	jdff dff_B_YaQADm9V9_2(.din(w_dff_B_Y9AFkIhl3_2),.dout(w_dff_B_YaQADm9V9_2),.clk(gclk));
	jdff dff_B_Ew6GQxoc6_2(.din(w_dff_B_YaQADm9V9_2),.dout(w_dff_B_Ew6GQxoc6_2),.clk(gclk));
	jdff dff_B_DuRkClK69_2(.din(w_dff_B_Ew6GQxoc6_2),.dout(w_dff_B_DuRkClK69_2),.clk(gclk));
	jdff dff_B_Mufn57ny6_1(.din(n1137),.dout(w_dff_B_Mufn57ny6_1),.clk(gclk));
	jdff dff_B_Ahh1psqS6_2(.din(n1038),.dout(w_dff_B_Ahh1psqS6_2),.clk(gclk));
	jdff dff_B_ut37sD9P3_2(.din(w_dff_B_Ahh1psqS6_2),.dout(w_dff_B_ut37sD9P3_2),.clk(gclk));
	jdff dff_B_q1BTJUjT5_2(.din(w_dff_B_ut37sD9P3_2),.dout(w_dff_B_q1BTJUjT5_2),.clk(gclk));
	jdff dff_B_KTOszVOS9_2(.din(w_dff_B_q1BTJUjT5_2),.dout(w_dff_B_KTOszVOS9_2),.clk(gclk));
	jdff dff_B_31q72oRG8_2(.din(w_dff_B_KTOszVOS9_2),.dout(w_dff_B_31q72oRG8_2),.clk(gclk));
	jdff dff_B_M6EiS9eb5_2(.din(w_dff_B_31q72oRG8_2),.dout(w_dff_B_M6EiS9eb5_2),.clk(gclk));
	jdff dff_B_Ym9cUVec8_2(.din(w_dff_B_M6EiS9eb5_2),.dout(w_dff_B_Ym9cUVec8_2),.clk(gclk));
	jdff dff_B_wrd8rwdu6_2(.din(w_dff_B_Ym9cUVec8_2),.dout(w_dff_B_wrd8rwdu6_2),.clk(gclk));
	jdff dff_B_UPwZxG364_2(.din(w_dff_B_wrd8rwdu6_2),.dout(w_dff_B_UPwZxG364_2),.clk(gclk));
	jdff dff_B_C1B0sqnh7_2(.din(w_dff_B_UPwZxG364_2),.dout(w_dff_B_C1B0sqnh7_2),.clk(gclk));
	jdff dff_B_VF1RJEtp6_2(.din(w_dff_B_C1B0sqnh7_2),.dout(w_dff_B_VF1RJEtp6_2),.clk(gclk));
	jdff dff_B_swQSk3Ee8_2(.din(w_dff_B_VF1RJEtp6_2),.dout(w_dff_B_swQSk3Ee8_2),.clk(gclk));
	jdff dff_B_9a7cZNhN7_2(.din(w_dff_B_swQSk3Ee8_2),.dout(w_dff_B_9a7cZNhN7_2),.clk(gclk));
	jdff dff_B_SpWeiUL30_2(.din(w_dff_B_9a7cZNhN7_2),.dout(w_dff_B_SpWeiUL30_2),.clk(gclk));
	jdff dff_B_8Yk8pSXQ5_2(.din(w_dff_B_SpWeiUL30_2),.dout(w_dff_B_8Yk8pSXQ5_2),.clk(gclk));
	jdff dff_B_pJbpBqgm0_2(.din(w_dff_B_8Yk8pSXQ5_2),.dout(w_dff_B_pJbpBqgm0_2),.clk(gclk));
	jdff dff_B_YG6VkVdh7_2(.din(w_dff_B_pJbpBqgm0_2),.dout(w_dff_B_YG6VkVdh7_2),.clk(gclk));
	jdff dff_B_6HM1VqsS9_2(.din(w_dff_B_YG6VkVdh7_2),.dout(w_dff_B_6HM1VqsS9_2),.clk(gclk));
	jdff dff_B_14u4atyu2_2(.din(w_dff_B_6HM1VqsS9_2),.dout(w_dff_B_14u4atyu2_2),.clk(gclk));
	jdff dff_B_N3EFo4EA1_2(.din(w_dff_B_14u4atyu2_2),.dout(w_dff_B_N3EFo4EA1_2),.clk(gclk));
	jdff dff_B_e4zhWBgy9_2(.din(w_dff_B_N3EFo4EA1_2),.dout(w_dff_B_e4zhWBgy9_2),.clk(gclk));
	jdff dff_B_AEMtq3kd1_2(.din(w_dff_B_e4zhWBgy9_2),.dout(w_dff_B_AEMtq3kd1_2),.clk(gclk));
	jdff dff_B_aILTKOZt6_2(.din(w_dff_B_AEMtq3kd1_2),.dout(w_dff_B_aILTKOZt6_2),.clk(gclk));
	jdff dff_B_i0Ted2BP2_2(.din(w_dff_B_aILTKOZt6_2),.dout(w_dff_B_i0Ted2BP2_2),.clk(gclk));
	jdff dff_B_f7L6yJwE3_1(.din(n1039),.dout(w_dff_B_f7L6yJwE3_1),.clk(gclk));
	jdff dff_B_b4J6Jsjq1_2(.din(n939),.dout(w_dff_B_b4J6Jsjq1_2),.clk(gclk));
	jdff dff_B_P9SHxo5I4_2(.din(w_dff_B_b4J6Jsjq1_2),.dout(w_dff_B_P9SHxo5I4_2),.clk(gclk));
	jdff dff_B_xLzQOyvP1_2(.din(w_dff_B_P9SHxo5I4_2),.dout(w_dff_B_xLzQOyvP1_2),.clk(gclk));
	jdff dff_B_yQUxV8S49_2(.din(w_dff_B_xLzQOyvP1_2),.dout(w_dff_B_yQUxV8S49_2),.clk(gclk));
	jdff dff_B_FufbPb9v3_2(.din(w_dff_B_yQUxV8S49_2),.dout(w_dff_B_FufbPb9v3_2),.clk(gclk));
	jdff dff_B_CE8s2ibK8_2(.din(w_dff_B_FufbPb9v3_2),.dout(w_dff_B_CE8s2ibK8_2),.clk(gclk));
	jdff dff_B_pmOtB5Vt7_2(.din(w_dff_B_CE8s2ibK8_2),.dout(w_dff_B_pmOtB5Vt7_2),.clk(gclk));
	jdff dff_B_YwrX7H9T5_2(.din(w_dff_B_pmOtB5Vt7_2),.dout(w_dff_B_YwrX7H9T5_2),.clk(gclk));
	jdff dff_B_GBzN1GgS7_2(.din(w_dff_B_YwrX7H9T5_2),.dout(w_dff_B_GBzN1GgS7_2),.clk(gclk));
	jdff dff_B_oTD8YeAJ6_2(.din(w_dff_B_GBzN1GgS7_2),.dout(w_dff_B_oTD8YeAJ6_2),.clk(gclk));
	jdff dff_B_X1DeDsWc9_2(.din(w_dff_B_oTD8YeAJ6_2),.dout(w_dff_B_X1DeDsWc9_2),.clk(gclk));
	jdff dff_B_fK9SMo8Y2_2(.din(w_dff_B_X1DeDsWc9_2),.dout(w_dff_B_fK9SMo8Y2_2),.clk(gclk));
	jdff dff_B_fdMk5D4N6_2(.din(w_dff_B_fK9SMo8Y2_2),.dout(w_dff_B_fdMk5D4N6_2),.clk(gclk));
	jdff dff_B_ZPHrhZsx2_2(.din(w_dff_B_fdMk5D4N6_2),.dout(w_dff_B_ZPHrhZsx2_2),.clk(gclk));
	jdff dff_B_tGvA40Y17_2(.din(w_dff_B_ZPHrhZsx2_2),.dout(w_dff_B_tGvA40Y17_2),.clk(gclk));
	jdff dff_B_6X0smcHS3_2(.din(w_dff_B_tGvA40Y17_2),.dout(w_dff_B_6X0smcHS3_2),.clk(gclk));
	jdff dff_B_6qx6EC9Z1_2(.din(w_dff_B_6X0smcHS3_2),.dout(w_dff_B_6qx6EC9Z1_2),.clk(gclk));
	jdff dff_B_fU6iMUOy2_2(.din(w_dff_B_6qx6EC9Z1_2),.dout(w_dff_B_fU6iMUOy2_2),.clk(gclk));
	jdff dff_B_74MAd6Bm5_2(.din(w_dff_B_fU6iMUOy2_2),.dout(w_dff_B_74MAd6Bm5_2),.clk(gclk));
	jdff dff_B_jId4Xbgr3_2(.din(w_dff_B_74MAd6Bm5_2),.dout(w_dff_B_jId4Xbgr3_2),.clk(gclk));
	jdff dff_B_zSWeITEe6_2(.din(w_dff_B_jId4Xbgr3_2),.dout(w_dff_B_zSWeITEe6_2),.clk(gclk));
	jdff dff_B_RV3WkNZc5_2(.din(w_dff_B_zSWeITEe6_2),.dout(w_dff_B_RV3WkNZc5_2),.clk(gclk));
	jdff dff_B_UA07Ppi04_1(.din(n940),.dout(w_dff_B_UA07Ppi04_1),.clk(gclk));
	jdff dff_B_mLuleuuW0_2(.din(n837),.dout(w_dff_B_mLuleuuW0_2),.clk(gclk));
	jdff dff_B_3HVmoRH91_2(.din(w_dff_B_mLuleuuW0_2),.dout(w_dff_B_3HVmoRH91_2),.clk(gclk));
	jdff dff_B_v24TIdmq9_2(.din(w_dff_B_3HVmoRH91_2),.dout(w_dff_B_v24TIdmq9_2),.clk(gclk));
	jdff dff_B_UiqP8xR29_2(.din(w_dff_B_v24TIdmq9_2),.dout(w_dff_B_UiqP8xR29_2),.clk(gclk));
	jdff dff_B_qE3SrZhB1_2(.din(w_dff_B_UiqP8xR29_2),.dout(w_dff_B_qE3SrZhB1_2),.clk(gclk));
	jdff dff_B_SeiPQxnU4_2(.din(w_dff_B_qE3SrZhB1_2),.dout(w_dff_B_SeiPQxnU4_2),.clk(gclk));
	jdff dff_B_ab8tWZ0k3_2(.din(w_dff_B_SeiPQxnU4_2),.dout(w_dff_B_ab8tWZ0k3_2),.clk(gclk));
	jdff dff_B_TC7iGZl78_2(.din(w_dff_B_ab8tWZ0k3_2),.dout(w_dff_B_TC7iGZl78_2),.clk(gclk));
	jdff dff_B_Z4Mvbzdo8_2(.din(w_dff_B_TC7iGZl78_2),.dout(w_dff_B_Z4Mvbzdo8_2),.clk(gclk));
	jdff dff_B_W2zLnZtg9_2(.din(w_dff_B_Z4Mvbzdo8_2),.dout(w_dff_B_W2zLnZtg9_2),.clk(gclk));
	jdff dff_B_Lm9SP8yb6_2(.din(w_dff_B_W2zLnZtg9_2),.dout(w_dff_B_Lm9SP8yb6_2),.clk(gclk));
	jdff dff_B_Vx26dSJb3_2(.din(w_dff_B_Lm9SP8yb6_2),.dout(w_dff_B_Vx26dSJb3_2),.clk(gclk));
	jdff dff_B_RfERzzQF0_2(.din(w_dff_B_Vx26dSJb3_2),.dout(w_dff_B_RfERzzQF0_2),.clk(gclk));
	jdff dff_B_dSeTHEyi8_2(.din(w_dff_B_RfERzzQF0_2),.dout(w_dff_B_dSeTHEyi8_2),.clk(gclk));
	jdff dff_B_OWVazIu22_2(.din(w_dff_B_dSeTHEyi8_2),.dout(w_dff_B_OWVazIu22_2),.clk(gclk));
	jdff dff_B_gqlFadwb0_2(.din(w_dff_B_OWVazIu22_2),.dout(w_dff_B_gqlFadwb0_2),.clk(gclk));
	jdff dff_B_px9xqlZb8_2(.din(w_dff_B_gqlFadwb0_2),.dout(w_dff_B_px9xqlZb8_2),.clk(gclk));
	jdff dff_B_8il9FhlR3_2(.din(w_dff_B_px9xqlZb8_2),.dout(w_dff_B_8il9FhlR3_2),.clk(gclk));
	jdff dff_B_MHn3v5bm5_2(.din(w_dff_B_8il9FhlR3_2),.dout(w_dff_B_MHn3v5bm5_2),.clk(gclk));
	jdff dff_B_46mVB41B0_2(.din(w_dff_B_MHn3v5bm5_2),.dout(w_dff_B_46mVB41B0_2),.clk(gclk));
	jdff dff_B_MJOCAlLn4_1(.din(n838),.dout(w_dff_B_MJOCAlLn4_1),.clk(gclk));
	jdff dff_B_YlTZMmhF9_2(.din(n739),.dout(w_dff_B_YlTZMmhF9_2),.clk(gclk));
	jdff dff_B_BQBdGkrS6_2(.din(w_dff_B_YlTZMmhF9_2),.dout(w_dff_B_BQBdGkrS6_2),.clk(gclk));
	jdff dff_B_kV6mGeTN8_2(.din(w_dff_B_BQBdGkrS6_2),.dout(w_dff_B_kV6mGeTN8_2),.clk(gclk));
	jdff dff_B_juG7tBaw2_2(.din(w_dff_B_kV6mGeTN8_2),.dout(w_dff_B_juG7tBaw2_2),.clk(gclk));
	jdff dff_B_wSYNEC4s3_2(.din(w_dff_B_juG7tBaw2_2),.dout(w_dff_B_wSYNEC4s3_2),.clk(gclk));
	jdff dff_B_pwQUszuN1_2(.din(w_dff_B_wSYNEC4s3_2),.dout(w_dff_B_pwQUszuN1_2),.clk(gclk));
	jdff dff_B_vHuksEov3_2(.din(w_dff_B_pwQUszuN1_2),.dout(w_dff_B_vHuksEov3_2),.clk(gclk));
	jdff dff_B_3RSOZf3m2_2(.din(w_dff_B_vHuksEov3_2),.dout(w_dff_B_3RSOZf3m2_2),.clk(gclk));
	jdff dff_B_d2Nh74uB8_2(.din(w_dff_B_3RSOZf3m2_2),.dout(w_dff_B_d2Nh74uB8_2),.clk(gclk));
	jdff dff_B_XiXhp0LZ6_2(.din(w_dff_B_d2Nh74uB8_2),.dout(w_dff_B_XiXhp0LZ6_2),.clk(gclk));
	jdff dff_B_QmdtSoxt5_2(.din(w_dff_B_XiXhp0LZ6_2),.dout(w_dff_B_QmdtSoxt5_2),.clk(gclk));
	jdff dff_B_q0LHuPxt9_2(.din(w_dff_B_QmdtSoxt5_2),.dout(w_dff_B_q0LHuPxt9_2),.clk(gclk));
	jdff dff_B_boZKUdGN0_2(.din(w_dff_B_q0LHuPxt9_2),.dout(w_dff_B_boZKUdGN0_2),.clk(gclk));
	jdff dff_B_ZXwtNYIJ0_2(.din(w_dff_B_boZKUdGN0_2),.dout(w_dff_B_ZXwtNYIJ0_2),.clk(gclk));
	jdff dff_B_LXUXNYAJ1_2(.din(w_dff_B_ZXwtNYIJ0_2),.dout(w_dff_B_LXUXNYAJ1_2),.clk(gclk));
	jdff dff_B_DeZzbMYc2_2(.din(w_dff_B_LXUXNYAJ1_2),.dout(w_dff_B_DeZzbMYc2_2),.clk(gclk));
	jdff dff_B_WdGtINt84_2(.din(w_dff_B_DeZzbMYc2_2),.dout(w_dff_B_WdGtINt84_2),.clk(gclk));
	jdff dff_B_FAqUrTuV1_2(.din(w_dff_B_WdGtINt84_2),.dout(w_dff_B_FAqUrTuV1_2),.clk(gclk));
	jdff dff_B_eQvYoeCl6_1(.din(n740),.dout(w_dff_B_eQvYoeCl6_1),.clk(gclk));
	jdff dff_B_LE9eh2jq5_2(.din(n647),.dout(w_dff_B_LE9eh2jq5_2),.clk(gclk));
	jdff dff_B_S9YSBhFz2_2(.din(w_dff_B_LE9eh2jq5_2),.dout(w_dff_B_S9YSBhFz2_2),.clk(gclk));
	jdff dff_B_rfL8FXnI9_2(.din(w_dff_B_S9YSBhFz2_2),.dout(w_dff_B_rfL8FXnI9_2),.clk(gclk));
	jdff dff_B_93mCKM6Z4_2(.din(w_dff_B_rfL8FXnI9_2),.dout(w_dff_B_93mCKM6Z4_2),.clk(gclk));
	jdff dff_B_WghgYMo79_2(.din(w_dff_B_93mCKM6Z4_2),.dout(w_dff_B_WghgYMo79_2),.clk(gclk));
	jdff dff_B_00wZDapF8_2(.din(w_dff_B_WghgYMo79_2),.dout(w_dff_B_00wZDapF8_2),.clk(gclk));
	jdff dff_B_6Wtocq1f8_2(.din(w_dff_B_00wZDapF8_2),.dout(w_dff_B_6Wtocq1f8_2),.clk(gclk));
	jdff dff_B_ZqZ3KqWL5_2(.din(w_dff_B_6Wtocq1f8_2),.dout(w_dff_B_ZqZ3KqWL5_2),.clk(gclk));
	jdff dff_B_dH851IKM2_2(.din(w_dff_B_ZqZ3KqWL5_2),.dout(w_dff_B_dH851IKM2_2),.clk(gclk));
	jdff dff_B_FdMleJGZ8_2(.din(w_dff_B_dH851IKM2_2),.dout(w_dff_B_FdMleJGZ8_2),.clk(gclk));
	jdff dff_B_e1yJGDxr3_2(.din(w_dff_B_FdMleJGZ8_2),.dout(w_dff_B_e1yJGDxr3_2),.clk(gclk));
	jdff dff_B_7JXVf2JF2_2(.din(w_dff_B_e1yJGDxr3_2),.dout(w_dff_B_7JXVf2JF2_2),.clk(gclk));
	jdff dff_B_AQ1RrBGH6_2(.din(w_dff_B_7JXVf2JF2_2),.dout(w_dff_B_AQ1RrBGH6_2),.clk(gclk));
	jdff dff_B_gMhffUhg5_2(.din(w_dff_B_AQ1RrBGH6_2),.dout(w_dff_B_gMhffUhg5_2),.clk(gclk));
	jdff dff_B_sWMeyzD53_2(.din(w_dff_B_gMhffUhg5_2),.dout(w_dff_B_sWMeyzD53_2),.clk(gclk));
	jdff dff_B_nQgUO1Pw2_2(.din(w_dff_B_sWMeyzD53_2),.dout(w_dff_B_nQgUO1Pw2_2),.clk(gclk));
	jdff dff_B_1P0ORXtM0_1(.din(n648),.dout(w_dff_B_1P0ORXtM0_1),.clk(gclk));
	jdff dff_B_7Tyh0ggS9_2(.din(n562),.dout(w_dff_B_7Tyh0ggS9_2),.clk(gclk));
	jdff dff_B_KFHZ1Yb21_2(.din(w_dff_B_7Tyh0ggS9_2),.dout(w_dff_B_KFHZ1Yb21_2),.clk(gclk));
	jdff dff_B_ir9JsQlc5_2(.din(w_dff_B_KFHZ1Yb21_2),.dout(w_dff_B_ir9JsQlc5_2),.clk(gclk));
	jdff dff_B_h9KxhMIl9_2(.din(w_dff_B_ir9JsQlc5_2),.dout(w_dff_B_h9KxhMIl9_2),.clk(gclk));
	jdff dff_B_G7Yk4JN51_2(.din(w_dff_B_h9KxhMIl9_2),.dout(w_dff_B_G7Yk4JN51_2),.clk(gclk));
	jdff dff_B_80vnigy17_2(.din(w_dff_B_G7Yk4JN51_2),.dout(w_dff_B_80vnigy17_2),.clk(gclk));
	jdff dff_B_82JXgsKz1_2(.din(w_dff_B_80vnigy17_2),.dout(w_dff_B_82JXgsKz1_2),.clk(gclk));
	jdff dff_B_r0Xe9xzX9_2(.din(w_dff_B_82JXgsKz1_2),.dout(w_dff_B_r0Xe9xzX9_2),.clk(gclk));
	jdff dff_B_WcjxHfu34_2(.din(w_dff_B_r0Xe9xzX9_2),.dout(w_dff_B_WcjxHfu34_2),.clk(gclk));
	jdff dff_B_vtc9D6FF4_2(.din(w_dff_B_WcjxHfu34_2),.dout(w_dff_B_vtc9D6FF4_2),.clk(gclk));
	jdff dff_B_mbeeLv1B3_2(.din(w_dff_B_vtc9D6FF4_2),.dout(w_dff_B_mbeeLv1B3_2),.clk(gclk));
	jdff dff_B_CIkdsVH92_2(.din(w_dff_B_mbeeLv1B3_2),.dout(w_dff_B_CIkdsVH92_2),.clk(gclk));
	jdff dff_B_YxTpVFRc4_2(.din(w_dff_B_CIkdsVH92_2),.dout(w_dff_B_YxTpVFRc4_2),.clk(gclk));
	jdff dff_B_9aOUgWIu3_2(.din(w_dff_B_YxTpVFRc4_2),.dout(w_dff_B_9aOUgWIu3_2),.clk(gclk));
	jdff dff_B_Y3iWifio0_1(.din(n563),.dout(w_dff_B_Y3iWifio0_1),.clk(gclk));
	jdff dff_B_tYY4aaKe3_2(.din(n484),.dout(w_dff_B_tYY4aaKe3_2),.clk(gclk));
	jdff dff_B_wnadlOra2_2(.din(w_dff_B_tYY4aaKe3_2),.dout(w_dff_B_wnadlOra2_2),.clk(gclk));
	jdff dff_B_c8nsEbdb6_2(.din(w_dff_B_wnadlOra2_2),.dout(w_dff_B_c8nsEbdb6_2),.clk(gclk));
	jdff dff_B_kR158B877_2(.din(w_dff_B_c8nsEbdb6_2),.dout(w_dff_B_kR158B877_2),.clk(gclk));
	jdff dff_B_fUrG5sDI8_2(.din(w_dff_B_kR158B877_2),.dout(w_dff_B_fUrG5sDI8_2),.clk(gclk));
	jdff dff_B_JP2hJyNA1_2(.din(w_dff_B_fUrG5sDI8_2),.dout(w_dff_B_JP2hJyNA1_2),.clk(gclk));
	jdff dff_B_ZHVSF9JX1_2(.din(w_dff_B_JP2hJyNA1_2),.dout(w_dff_B_ZHVSF9JX1_2),.clk(gclk));
	jdff dff_B_XUi64OdK7_2(.din(w_dff_B_ZHVSF9JX1_2),.dout(w_dff_B_XUi64OdK7_2),.clk(gclk));
	jdff dff_B_inSMvfMl8_2(.din(w_dff_B_XUi64OdK7_2),.dout(w_dff_B_inSMvfMl8_2),.clk(gclk));
	jdff dff_B_s5ZoFUJN4_2(.din(w_dff_B_inSMvfMl8_2),.dout(w_dff_B_s5ZoFUJN4_2),.clk(gclk));
	jdff dff_B_I31Na36j0_2(.din(w_dff_B_s5ZoFUJN4_2),.dout(w_dff_B_I31Na36j0_2),.clk(gclk));
	jdff dff_B_W0AeNeTW6_2(.din(w_dff_B_I31Na36j0_2),.dout(w_dff_B_W0AeNeTW6_2),.clk(gclk));
	jdff dff_B_0ttUigoW2_1(.din(n485),.dout(w_dff_B_0ttUigoW2_1),.clk(gclk));
	jdff dff_B_tutDU4Of6_2(.din(n413),.dout(w_dff_B_tutDU4Of6_2),.clk(gclk));
	jdff dff_B_62YYaDSn3_2(.din(w_dff_B_tutDU4Of6_2),.dout(w_dff_B_62YYaDSn3_2),.clk(gclk));
	jdff dff_B_YRIm5N3Z8_2(.din(w_dff_B_62YYaDSn3_2),.dout(w_dff_B_YRIm5N3Z8_2),.clk(gclk));
	jdff dff_B_GVrHlklT3_2(.din(w_dff_B_YRIm5N3Z8_2),.dout(w_dff_B_GVrHlklT3_2),.clk(gclk));
	jdff dff_B_ub2s6Tib8_2(.din(w_dff_B_GVrHlklT3_2),.dout(w_dff_B_ub2s6Tib8_2),.clk(gclk));
	jdff dff_B_Hah5zG2R3_2(.din(w_dff_B_ub2s6Tib8_2),.dout(w_dff_B_Hah5zG2R3_2),.clk(gclk));
	jdff dff_B_th4CQD6f5_2(.din(w_dff_B_Hah5zG2R3_2),.dout(w_dff_B_th4CQD6f5_2),.clk(gclk));
	jdff dff_B_nyjW9aRJ9_2(.din(w_dff_B_th4CQD6f5_2),.dout(w_dff_B_nyjW9aRJ9_2),.clk(gclk));
	jdff dff_B_txcvjfHr9_2(.din(w_dff_B_nyjW9aRJ9_2),.dout(w_dff_B_txcvjfHr9_2),.clk(gclk));
	jdff dff_B_VdCinP0T1_2(.din(w_dff_B_txcvjfHr9_2),.dout(w_dff_B_VdCinP0T1_2),.clk(gclk));
	jdff dff_B_2eyN18HJ6_2(.din(n416),.dout(w_dff_B_2eyN18HJ6_2),.clk(gclk));
	jdff dff_B_Kf2vFNnD5_2(.din(w_dff_B_2eyN18HJ6_2),.dout(w_dff_B_Kf2vFNnD5_2),.clk(gclk));
	jdff dff_B_RodJbxBX1_2(.din(w_dff_B_Kf2vFNnD5_2),.dout(w_dff_B_RodJbxBX1_2),.clk(gclk));
	jdff dff_B_aklalK3q6_1(.din(n414),.dout(w_dff_B_aklalK3q6_1),.clk(gclk));
	jdff dff_B_b58sizGw8_2(.din(n350),.dout(w_dff_B_b58sizGw8_2),.clk(gclk));
	jdff dff_B_puJmDR174_2(.din(w_dff_B_b58sizGw8_2),.dout(w_dff_B_puJmDR174_2),.clk(gclk));
	jdff dff_B_fD4v50RS7_2(.din(w_dff_B_puJmDR174_2),.dout(w_dff_B_fD4v50RS7_2),.clk(gclk));
	jdff dff_B_dKdNc2dK3_2(.din(w_dff_B_fD4v50RS7_2),.dout(w_dff_B_dKdNc2dK3_2),.clk(gclk));
	jdff dff_B_xso4Npzq4_2(.din(w_dff_B_dKdNc2dK3_2),.dout(w_dff_B_xso4Npzq4_2),.clk(gclk));
	jdff dff_B_ZYD8hTSh7_1(.din(n352),.dout(w_dff_B_ZYD8hTSh7_1),.clk(gclk));
	jdff dff_B_SbNQ4RCr9_2(.din(n295),.dout(w_dff_B_SbNQ4RCr9_2),.clk(gclk));
	jdff dff_B_lJQVzpmo9_2(.din(w_dff_B_SbNQ4RCr9_2),.dout(w_dff_B_lJQVzpmo9_2),.clk(gclk));
	jdff dff_B_1jyfj3PW8_2(.din(w_dff_B_lJQVzpmo9_2),.dout(w_dff_B_1jyfj3PW8_2),.clk(gclk));
	jdff dff_B_Q2Fswjgg1_0(.din(n300),.dout(w_dff_B_Q2Fswjgg1_0),.clk(gclk));
	jdff dff_B_DIG1ikH87_0(.din(w_dff_B_Q2Fswjgg1_0),.dout(w_dff_B_DIG1ikH87_0),.clk(gclk));
	jdff dff_A_ZDNfXdBN8_0(.dout(w_n243_0[0]),.din(w_dff_A_ZDNfXdBN8_0),.clk(gclk));
	jdff dff_A_D70Zf41k4_0(.dout(w_dff_A_ZDNfXdBN8_0),.din(w_dff_A_D70Zf41k4_0),.clk(gclk));
	jdff dff_A_fsvH5Wdk4_1(.dout(w_n243_0[1]),.din(w_dff_A_fsvH5Wdk4_1),.clk(gclk));
	jdff dff_A_8uBIIrPF3_1(.dout(w_dff_A_fsvH5Wdk4_1),.din(w_dff_A_8uBIIrPF3_1),.clk(gclk));
	jdff dff_B_ECy4dX4h6_2(.din(n1534),.dout(w_dff_B_ECy4dX4h6_2),.clk(gclk));
	jdff dff_B_WFe17quy4_2(.din(w_dff_B_ECy4dX4h6_2),.dout(w_dff_B_WFe17quy4_2),.clk(gclk));
	jdff dff_B_ZIvl7ino7_1(.din(n1532),.dout(w_dff_B_ZIvl7ino7_1),.clk(gclk));
	jdff dff_B_BEz0cK1R0_2(.din(n1466),.dout(w_dff_B_BEz0cK1R0_2),.clk(gclk));
	jdff dff_B_M7MyesCO6_2(.din(w_dff_B_BEz0cK1R0_2),.dout(w_dff_B_M7MyesCO6_2),.clk(gclk));
	jdff dff_B_RwZlw2uP8_2(.din(w_dff_B_M7MyesCO6_2),.dout(w_dff_B_RwZlw2uP8_2),.clk(gclk));
	jdff dff_B_ZFfcxAnt4_2(.din(w_dff_B_RwZlw2uP8_2),.dout(w_dff_B_ZFfcxAnt4_2),.clk(gclk));
	jdff dff_B_5ipsmv8G1_2(.din(w_dff_B_ZFfcxAnt4_2),.dout(w_dff_B_5ipsmv8G1_2),.clk(gclk));
	jdff dff_B_lsj78i6I6_2(.din(w_dff_B_5ipsmv8G1_2),.dout(w_dff_B_lsj78i6I6_2),.clk(gclk));
	jdff dff_B_wTpE2uP61_2(.din(w_dff_B_lsj78i6I6_2),.dout(w_dff_B_wTpE2uP61_2),.clk(gclk));
	jdff dff_B_Hk8JWjcv9_2(.din(w_dff_B_wTpE2uP61_2),.dout(w_dff_B_Hk8JWjcv9_2),.clk(gclk));
	jdff dff_B_Ge34LjSF4_2(.din(w_dff_B_Hk8JWjcv9_2),.dout(w_dff_B_Ge34LjSF4_2),.clk(gclk));
	jdff dff_B_kodSHwjr0_2(.din(w_dff_B_Ge34LjSF4_2),.dout(w_dff_B_kodSHwjr0_2),.clk(gclk));
	jdff dff_B_MVIxVjYi0_2(.din(w_dff_B_kodSHwjr0_2),.dout(w_dff_B_MVIxVjYi0_2),.clk(gclk));
	jdff dff_B_Bp60VGvQ3_2(.din(w_dff_B_MVIxVjYi0_2),.dout(w_dff_B_Bp60VGvQ3_2),.clk(gclk));
	jdff dff_B_mdOdkvQp7_2(.din(w_dff_B_Bp60VGvQ3_2),.dout(w_dff_B_mdOdkvQp7_2),.clk(gclk));
	jdff dff_B_VMlaPO3N0_2(.din(w_dff_B_mdOdkvQp7_2),.dout(w_dff_B_VMlaPO3N0_2),.clk(gclk));
	jdff dff_B_TbibVkUy8_2(.din(w_dff_B_VMlaPO3N0_2),.dout(w_dff_B_TbibVkUy8_2),.clk(gclk));
	jdff dff_B_ULTt1x6m0_2(.din(w_dff_B_TbibVkUy8_2),.dout(w_dff_B_ULTt1x6m0_2),.clk(gclk));
	jdff dff_B_AbNtEIjL5_2(.din(w_dff_B_ULTt1x6m0_2),.dout(w_dff_B_AbNtEIjL5_2),.clk(gclk));
	jdff dff_B_lvE1obt88_2(.din(w_dff_B_AbNtEIjL5_2),.dout(w_dff_B_lvE1obt88_2),.clk(gclk));
	jdff dff_B_iBUngahR0_2(.din(w_dff_B_lvE1obt88_2),.dout(w_dff_B_iBUngahR0_2),.clk(gclk));
	jdff dff_B_I9h71T3S9_2(.din(w_dff_B_iBUngahR0_2),.dout(w_dff_B_I9h71T3S9_2),.clk(gclk));
	jdff dff_B_i8zJOOv59_2(.din(w_dff_B_I9h71T3S9_2),.dout(w_dff_B_i8zJOOv59_2),.clk(gclk));
	jdff dff_B_IV3hgyvv5_2(.din(w_dff_B_i8zJOOv59_2),.dout(w_dff_B_IV3hgyvv5_2),.clk(gclk));
	jdff dff_B_8Vh7H1n24_2(.din(w_dff_B_IV3hgyvv5_2),.dout(w_dff_B_8Vh7H1n24_2),.clk(gclk));
	jdff dff_B_jIWbACyW1_2(.din(w_dff_B_8Vh7H1n24_2),.dout(w_dff_B_jIWbACyW1_2),.clk(gclk));
	jdff dff_B_JDTFM5R30_2(.din(w_dff_B_jIWbACyW1_2),.dout(w_dff_B_JDTFM5R30_2),.clk(gclk));
	jdff dff_B_xrfzY9ts9_2(.din(w_dff_B_JDTFM5R30_2),.dout(w_dff_B_xrfzY9ts9_2),.clk(gclk));
	jdff dff_B_rw8SYItt1_2(.din(w_dff_B_xrfzY9ts9_2),.dout(w_dff_B_rw8SYItt1_2),.clk(gclk));
	jdff dff_B_EmR8Mzgg3_2(.din(w_dff_B_rw8SYItt1_2),.dout(w_dff_B_EmR8Mzgg3_2),.clk(gclk));
	jdff dff_B_jMujvKHS0_2(.din(w_dff_B_EmR8Mzgg3_2),.dout(w_dff_B_jMujvKHS0_2),.clk(gclk));
	jdff dff_B_pjdjxP1g7_2(.din(w_dff_B_jMujvKHS0_2),.dout(w_dff_B_pjdjxP1g7_2),.clk(gclk));
	jdff dff_B_bYs6Ix2a4_2(.din(w_dff_B_pjdjxP1g7_2),.dout(w_dff_B_bYs6Ix2a4_2),.clk(gclk));
	jdff dff_B_EKJJA52A3_2(.din(w_dff_B_bYs6Ix2a4_2),.dout(w_dff_B_EKJJA52A3_2),.clk(gclk));
	jdff dff_B_i14y3HXd4_2(.din(w_dff_B_EKJJA52A3_2),.dout(w_dff_B_i14y3HXd4_2),.clk(gclk));
	jdff dff_B_FnD7VnyZ3_2(.din(w_dff_B_i14y3HXd4_2),.dout(w_dff_B_FnD7VnyZ3_2),.clk(gclk));
	jdff dff_B_mBUFPWuq2_2(.din(w_dff_B_FnD7VnyZ3_2),.dout(w_dff_B_mBUFPWuq2_2),.clk(gclk));
	jdff dff_B_3uOXTrKJ1_2(.din(w_dff_B_mBUFPWuq2_2),.dout(w_dff_B_3uOXTrKJ1_2),.clk(gclk));
	jdff dff_B_T1uQ9chI8_1(.din(n1530),.dout(w_dff_B_T1uQ9chI8_1),.clk(gclk));
	jdff dff_A_CXO8gbcQ6_1(.dout(w_n1469_0[1]),.din(w_dff_A_CXO8gbcQ6_1),.clk(gclk));
	jdff dff_B_JxXpUVSx0_1(.din(n1467),.dout(w_dff_B_JxXpUVSx0_1),.clk(gclk));
	jdff dff_B_uVZaACIL5_2(.din(n1395),.dout(w_dff_B_uVZaACIL5_2),.clk(gclk));
	jdff dff_B_bHSTeePt1_2(.din(w_dff_B_uVZaACIL5_2),.dout(w_dff_B_bHSTeePt1_2),.clk(gclk));
	jdff dff_B_htlcsEFH0_2(.din(w_dff_B_bHSTeePt1_2),.dout(w_dff_B_htlcsEFH0_2),.clk(gclk));
	jdff dff_B_lcj2qm6t2_2(.din(w_dff_B_htlcsEFH0_2),.dout(w_dff_B_lcj2qm6t2_2),.clk(gclk));
	jdff dff_B_EtghrVxC9_2(.din(w_dff_B_lcj2qm6t2_2),.dout(w_dff_B_EtghrVxC9_2),.clk(gclk));
	jdff dff_B_5liMHcCa9_2(.din(w_dff_B_EtghrVxC9_2),.dout(w_dff_B_5liMHcCa9_2),.clk(gclk));
	jdff dff_B_Y9BODGAs9_2(.din(w_dff_B_5liMHcCa9_2),.dout(w_dff_B_Y9BODGAs9_2),.clk(gclk));
	jdff dff_B_B9fvqJFy0_2(.din(w_dff_B_Y9BODGAs9_2),.dout(w_dff_B_B9fvqJFy0_2),.clk(gclk));
	jdff dff_B_abzMz8sP6_2(.din(w_dff_B_B9fvqJFy0_2),.dout(w_dff_B_abzMz8sP6_2),.clk(gclk));
	jdff dff_B_iOLw0N4M6_2(.din(w_dff_B_abzMz8sP6_2),.dout(w_dff_B_iOLw0N4M6_2),.clk(gclk));
	jdff dff_B_VTnpXutI6_2(.din(w_dff_B_iOLw0N4M6_2),.dout(w_dff_B_VTnpXutI6_2),.clk(gclk));
	jdff dff_B_6NU93XRJ6_2(.din(w_dff_B_VTnpXutI6_2),.dout(w_dff_B_6NU93XRJ6_2),.clk(gclk));
	jdff dff_B_GdKwB8Lv4_2(.din(w_dff_B_6NU93XRJ6_2),.dout(w_dff_B_GdKwB8Lv4_2),.clk(gclk));
	jdff dff_B_14jSVvej2_2(.din(w_dff_B_GdKwB8Lv4_2),.dout(w_dff_B_14jSVvej2_2),.clk(gclk));
	jdff dff_B_zZ9gawPG5_2(.din(w_dff_B_14jSVvej2_2),.dout(w_dff_B_zZ9gawPG5_2),.clk(gclk));
	jdff dff_B_TBrCzMc67_2(.din(w_dff_B_zZ9gawPG5_2),.dout(w_dff_B_TBrCzMc67_2),.clk(gclk));
	jdff dff_B_wAy2h7Xi6_2(.din(w_dff_B_TBrCzMc67_2),.dout(w_dff_B_wAy2h7Xi6_2),.clk(gclk));
	jdff dff_B_pjFifiQt1_2(.din(w_dff_B_wAy2h7Xi6_2),.dout(w_dff_B_pjFifiQt1_2),.clk(gclk));
	jdff dff_B_aQQlawh42_2(.din(w_dff_B_pjFifiQt1_2),.dout(w_dff_B_aQQlawh42_2),.clk(gclk));
	jdff dff_B_7fZWpBWh8_2(.din(w_dff_B_aQQlawh42_2),.dout(w_dff_B_7fZWpBWh8_2),.clk(gclk));
	jdff dff_B_2RVGEWwl0_2(.din(w_dff_B_7fZWpBWh8_2),.dout(w_dff_B_2RVGEWwl0_2),.clk(gclk));
	jdff dff_B_Dw2SbVdT4_2(.din(w_dff_B_2RVGEWwl0_2),.dout(w_dff_B_Dw2SbVdT4_2),.clk(gclk));
	jdff dff_B_ZmmyUifv6_2(.din(w_dff_B_Dw2SbVdT4_2),.dout(w_dff_B_ZmmyUifv6_2),.clk(gclk));
	jdff dff_B_E6mFrMLs9_2(.din(w_dff_B_ZmmyUifv6_2),.dout(w_dff_B_E6mFrMLs9_2),.clk(gclk));
	jdff dff_B_9ONz9mZI6_2(.din(w_dff_B_E6mFrMLs9_2),.dout(w_dff_B_9ONz9mZI6_2),.clk(gclk));
	jdff dff_B_YpinjtRB9_2(.din(w_dff_B_9ONz9mZI6_2),.dout(w_dff_B_YpinjtRB9_2),.clk(gclk));
	jdff dff_B_wfU26BUj4_2(.din(w_dff_B_YpinjtRB9_2),.dout(w_dff_B_wfU26BUj4_2),.clk(gclk));
	jdff dff_B_ccnFoE9b3_2(.din(w_dff_B_wfU26BUj4_2),.dout(w_dff_B_ccnFoE9b3_2),.clk(gclk));
	jdff dff_B_iyeVOivS0_2(.din(w_dff_B_ccnFoE9b3_2),.dout(w_dff_B_iyeVOivS0_2),.clk(gclk));
	jdff dff_B_ouB1yI5z7_2(.din(w_dff_B_iyeVOivS0_2),.dout(w_dff_B_ouB1yI5z7_2),.clk(gclk));
	jdff dff_B_YozbgheA4_2(.din(w_dff_B_ouB1yI5z7_2),.dout(w_dff_B_YozbgheA4_2),.clk(gclk));
	jdff dff_B_teb3lBS75_2(.din(n1398),.dout(w_dff_B_teb3lBS75_2),.clk(gclk));
	jdff dff_B_bBMX1SXG4_1(.din(n1396),.dout(w_dff_B_bBMX1SXG4_1),.clk(gclk));
	jdff dff_B_3tYya2XY0_2(.din(n1317),.dout(w_dff_B_3tYya2XY0_2),.clk(gclk));
	jdff dff_B_v1RQoMpg7_2(.din(w_dff_B_3tYya2XY0_2),.dout(w_dff_B_v1RQoMpg7_2),.clk(gclk));
	jdff dff_B_WQcnvxIS1_2(.din(w_dff_B_v1RQoMpg7_2),.dout(w_dff_B_WQcnvxIS1_2),.clk(gclk));
	jdff dff_B_rw1dArzp0_2(.din(w_dff_B_WQcnvxIS1_2),.dout(w_dff_B_rw1dArzp0_2),.clk(gclk));
	jdff dff_B_0IfI2JDD8_2(.din(w_dff_B_rw1dArzp0_2),.dout(w_dff_B_0IfI2JDD8_2),.clk(gclk));
	jdff dff_B_3E7Ld6Bs0_2(.din(w_dff_B_0IfI2JDD8_2),.dout(w_dff_B_3E7Ld6Bs0_2),.clk(gclk));
	jdff dff_B_X30TRNvY3_2(.din(w_dff_B_3E7Ld6Bs0_2),.dout(w_dff_B_X30TRNvY3_2),.clk(gclk));
	jdff dff_B_aeo0v2Tf2_2(.din(w_dff_B_X30TRNvY3_2),.dout(w_dff_B_aeo0v2Tf2_2),.clk(gclk));
	jdff dff_B_IgGgScUL5_2(.din(w_dff_B_aeo0v2Tf2_2),.dout(w_dff_B_IgGgScUL5_2),.clk(gclk));
	jdff dff_B_g5uEQv1I1_2(.din(w_dff_B_IgGgScUL5_2),.dout(w_dff_B_g5uEQv1I1_2),.clk(gclk));
	jdff dff_B_T6fOICOU1_2(.din(w_dff_B_g5uEQv1I1_2),.dout(w_dff_B_T6fOICOU1_2),.clk(gclk));
	jdff dff_B_OFyTDMBY4_2(.din(w_dff_B_T6fOICOU1_2),.dout(w_dff_B_OFyTDMBY4_2),.clk(gclk));
	jdff dff_B_tmKxvrc41_2(.din(w_dff_B_OFyTDMBY4_2),.dout(w_dff_B_tmKxvrc41_2),.clk(gclk));
	jdff dff_B_bKKRr2714_2(.din(w_dff_B_tmKxvrc41_2),.dout(w_dff_B_bKKRr2714_2),.clk(gclk));
	jdff dff_B_U5ervHxI2_2(.din(w_dff_B_bKKRr2714_2),.dout(w_dff_B_U5ervHxI2_2),.clk(gclk));
	jdff dff_B_lOBdCHeu6_2(.din(w_dff_B_U5ervHxI2_2),.dout(w_dff_B_lOBdCHeu6_2),.clk(gclk));
	jdff dff_B_gqgheVp73_2(.din(w_dff_B_lOBdCHeu6_2),.dout(w_dff_B_gqgheVp73_2),.clk(gclk));
	jdff dff_B_gtuRSp407_2(.din(w_dff_B_gqgheVp73_2),.dout(w_dff_B_gtuRSp407_2),.clk(gclk));
	jdff dff_B_hcyNNc3Z9_2(.din(w_dff_B_gtuRSp407_2),.dout(w_dff_B_hcyNNc3Z9_2),.clk(gclk));
	jdff dff_B_8eh2Lelk7_2(.din(w_dff_B_hcyNNc3Z9_2),.dout(w_dff_B_8eh2Lelk7_2),.clk(gclk));
	jdff dff_B_5ze0fl2n3_2(.din(w_dff_B_8eh2Lelk7_2),.dout(w_dff_B_5ze0fl2n3_2),.clk(gclk));
	jdff dff_B_48bVh6RE8_2(.din(w_dff_B_5ze0fl2n3_2),.dout(w_dff_B_48bVh6RE8_2),.clk(gclk));
	jdff dff_B_ZRZU8uOx3_2(.din(w_dff_B_48bVh6RE8_2),.dout(w_dff_B_ZRZU8uOx3_2),.clk(gclk));
	jdff dff_B_YHapp4X36_2(.din(w_dff_B_ZRZU8uOx3_2),.dout(w_dff_B_YHapp4X36_2),.clk(gclk));
	jdff dff_B_mLXa6sQJ9_2(.din(w_dff_B_YHapp4X36_2),.dout(w_dff_B_mLXa6sQJ9_2),.clk(gclk));
	jdff dff_B_e85M0g4m3_2(.din(w_dff_B_mLXa6sQJ9_2),.dout(w_dff_B_e85M0g4m3_2),.clk(gclk));
	jdff dff_B_PQn5RWsp2_2(.din(w_dff_B_e85M0g4m3_2),.dout(w_dff_B_PQn5RWsp2_2),.clk(gclk));
	jdff dff_B_NV8HOxjN1_2(.din(w_dff_B_PQn5RWsp2_2),.dout(w_dff_B_NV8HOxjN1_2),.clk(gclk));
	jdff dff_B_tZqSwIO23_1(.din(n1318),.dout(w_dff_B_tZqSwIO23_1),.clk(gclk));
	jdff dff_B_P4joCQYg5_2(.din(n1232),.dout(w_dff_B_P4joCQYg5_2),.clk(gclk));
	jdff dff_B_QmfJxSJy7_2(.din(w_dff_B_P4joCQYg5_2),.dout(w_dff_B_QmfJxSJy7_2),.clk(gclk));
	jdff dff_B_LV407I1u0_2(.din(w_dff_B_QmfJxSJy7_2),.dout(w_dff_B_LV407I1u0_2),.clk(gclk));
	jdff dff_B_oJFCao3m1_2(.din(w_dff_B_LV407I1u0_2),.dout(w_dff_B_oJFCao3m1_2),.clk(gclk));
	jdff dff_B_V368PBcs7_2(.din(w_dff_B_oJFCao3m1_2),.dout(w_dff_B_V368PBcs7_2),.clk(gclk));
	jdff dff_B_row4fal99_2(.din(w_dff_B_V368PBcs7_2),.dout(w_dff_B_row4fal99_2),.clk(gclk));
	jdff dff_B_kZp2BKhT6_2(.din(w_dff_B_row4fal99_2),.dout(w_dff_B_kZp2BKhT6_2),.clk(gclk));
	jdff dff_B_Pl7SyZlU7_2(.din(w_dff_B_kZp2BKhT6_2),.dout(w_dff_B_Pl7SyZlU7_2),.clk(gclk));
	jdff dff_B_Xt4tnPcO7_2(.din(w_dff_B_Pl7SyZlU7_2),.dout(w_dff_B_Xt4tnPcO7_2),.clk(gclk));
	jdff dff_B_lpmOVdQ54_2(.din(w_dff_B_Xt4tnPcO7_2),.dout(w_dff_B_lpmOVdQ54_2),.clk(gclk));
	jdff dff_B_LsgDdFIg8_2(.din(w_dff_B_lpmOVdQ54_2),.dout(w_dff_B_LsgDdFIg8_2),.clk(gclk));
	jdff dff_B_qElhWWo46_2(.din(w_dff_B_LsgDdFIg8_2),.dout(w_dff_B_qElhWWo46_2),.clk(gclk));
	jdff dff_B_F0JHrGAW2_2(.din(w_dff_B_qElhWWo46_2),.dout(w_dff_B_F0JHrGAW2_2),.clk(gclk));
	jdff dff_B_Vu9BHf0p0_2(.din(w_dff_B_F0JHrGAW2_2),.dout(w_dff_B_Vu9BHf0p0_2),.clk(gclk));
	jdff dff_B_0VP4dFnq5_2(.din(w_dff_B_Vu9BHf0p0_2),.dout(w_dff_B_0VP4dFnq5_2),.clk(gclk));
	jdff dff_B_0umoayER2_2(.din(w_dff_B_0VP4dFnq5_2),.dout(w_dff_B_0umoayER2_2),.clk(gclk));
	jdff dff_B_B6g4u4xj8_2(.din(w_dff_B_0umoayER2_2),.dout(w_dff_B_B6g4u4xj8_2),.clk(gclk));
	jdff dff_B_x5D2HBSH9_2(.din(w_dff_B_B6g4u4xj8_2),.dout(w_dff_B_x5D2HBSH9_2),.clk(gclk));
	jdff dff_B_i4IWkU3F9_2(.din(w_dff_B_x5D2HBSH9_2),.dout(w_dff_B_i4IWkU3F9_2),.clk(gclk));
	jdff dff_B_XplDPMIh4_2(.din(w_dff_B_i4IWkU3F9_2),.dout(w_dff_B_XplDPMIh4_2),.clk(gclk));
	jdff dff_B_iehERLSP1_2(.din(w_dff_B_XplDPMIh4_2),.dout(w_dff_B_iehERLSP1_2),.clk(gclk));
	jdff dff_B_cg2rVmTo2_2(.din(w_dff_B_iehERLSP1_2),.dout(w_dff_B_cg2rVmTo2_2),.clk(gclk));
	jdff dff_B_q7tsYwk66_2(.din(w_dff_B_cg2rVmTo2_2),.dout(w_dff_B_q7tsYwk66_2),.clk(gclk));
	jdff dff_B_pWZC72y62_2(.din(w_dff_B_q7tsYwk66_2),.dout(w_dff_B_pWZC72y62_2),.clk(gclk));
	jdff dff_B_9dnTYMnJ8_2(.din(w_dff_B_pWZC72y62_2),.dout(w_dff_B_9dnTYMnJ8_2),.clk(gclk));
	jdff dff_B_p41h6Qti7_2(.din(w_dff_B_9dnTYMnJ8_2),.dout(w_dff_B_p41h6Qti7_2),.clk(gclk));
	jdff dff_B_9QvM6iid7_1(.din(n1233),.dout(w_dff_B_9QvM6iid7_1),.clk(gclk));
	jdff dff_B_BkfCbZWX6_2(.din(n1141),.dout(w_dff_B_BkfCbZWX6_2),.clk(gclk));
	jdff dff_B_kUUHDAXv5_2(.din(w_dff_B_BkfCbZWX6_2),.dout(w_dff_B_kUUHDAXv5_2),.clk(gclk));
	jdff dff_B_9EZKI3by1_2(.din(w_dff_B_kUUHDAXv5_2),.dout(w_dff_B_9EZKI3by1_2),.clk(gclk));
	jdff dff_B_fiFWuJxT7_2(.din(w_dff_B_9EZKI3by1_2),.dout(w_dff_B_fiFWuJxT7_2),.clk(gclk));
	jdff dff_B_zdWlGihM1_2(.din(w_dff_B_fiFWuJxT7_2),.dout(w_dff_B_zdWlGihM1_2),.clk(gclk));
	jdff dff_B_p3773nxj0_2(.din(w_dff_B_zdWlGihM1_2),.dout(w_dff_B_p3773nxj0_2),.clk(gclk));
	jdff dff_B_16hmqoeA9_2(.din(w_dff_B_p3773nxj0_2),.dout(w_dff_B_16hmqoeA9_2),.clk(gclk));
	jdff dff_B_wwUoVEIr5_2(.din(w_dff_B_16hmqoeA9_2),.dout(w_dff_B_wwUoVEIr5_2),.clk(gclk));
	jdff dff_B_ZOXR1ScA0_2(.din(w_dff_B_wwUoVEIr5_2),.dout(w_dff_B_ZOXR1ScA0_2),.clk(gclk));
	jdff dff_B_7MfeQt6P9_2(.din(w_dff_B_ZOXR1ScA0_2),.dout(w_dff_B_7MfeQt6P9_2),.clk(gclk));
	jdff dff_B_0Bgro4s80_2(.din(w_dff_B_7MfeQt6P9_2),.dout(w_dff_B_0Bgro4s80_2),.clk(gclk));
	jdff dff_B_SDkt6Y1F9_2(.din(w_dff_B_0Bgro4s80_2),.dout(w_dff_B_SDkt6Y1F9_2),.clk(gclk));
	jdff dff_B_IWldop6H8_2(.din(w_dff_B_SDkt6Y1F9_2),.dout(w_dff_B_IWldop6H8_2),.clk(gclk));
	jdff dff_B_C5LSL2EQ1_2(.din(w_dff_B_IWldop6H8_2),.dout(w_dff_B_C5LSL2EQ1_2),.clk(gclk));
	jdff dff_B_sDq8JODP6_2(.din(w_dff_B_C5LSL2EQ1_2),.dout(w_dff_B_sDq8JODP6_2),.clk(gclk));
	jdff dff_B_XZh9nUX64_2(.din(w_dff_B_sDq8JODP6_2),.dout(w_dff_B_XZh9nUX64_2),.clk(gclk));
	jdff dff_B_SGlk6sFj3_2(.din(w_dff_B_XZh9nUX64_2),.dout(w_dff_B_SGlk6sFj3_2),.clk(gclk));
	jdff dff_B_Pyo4Rq5w3_2(.din(w_dff_B_SGlk6sFj3_2),.dout(w_dff_B_Pyo4Rq5w3_2),.clk(gclk));
	jdff dff_B_gsKldul77_2(.din(w_dff_B_Pyo4Rq5w3_2),.dout(w_dff_B_gsKldul77_2),.clk(gclk));
	jdff dff_B_CKCIkqQH0_2(.din(w_dff_B_gsKldul77_2),.dout(w_dff_B_CKCIkqQH0_2),.clk(gclk));
	jdff dff_B_yhzC7Sh76_2(.din(w_dff_B_CKCIkqQH0_2),.dout(w_dff_B_yhzC7Sh76_2),.clk(gclk));
	jdff dff_B_YDp39mFV0_2(.din(w_dff_B_yhzC7Sh76_2),.dout(w_dff_B_YDp39mFV0_2),.clk(gclk));
	jdff dff_B_4fkW6JxK3_2(.din(w_dff_B_YDp39mFV0_2),.dout(w_dff_B_4fkW6JxK3_2),.clk(gclk));
	jdff dff_B_jgJwiJ2Q9_2(.din(w_dff_B_4fkW6JxK3_2),.dout(w_dff_B_jgJwiJ2Q9_2),.clk(gclk));
	jdff dff_B_PyIWdvaA6_1(.din(n1142),.dout(w_dff_B_PyIWdvaA6_1),.clk(gclk));
	jdff dff_B_lbmaXOJY1_2(.din(n1043),.dout(w_dff_B_lbmaXOJY1_2),.clk(gclk));
	jdff dff_B_mPa3lmCK3_2(.din(w_dff_B_lbmaXOJY1_2),.dout(w_dff_B_mPa3lmCK3_2),.clk(gclk));
	jdff dff_B_8Yr477c90_2(.din(w_dff_B_mPa3lmCK3_2),.dout(w_dff_B_8Yr477c90_2),.clk(gclk));
	jdff dff_B_sW1WAFPS0_2(.din(w_dff_B_8Yr477c90_2),.dout(w_dff_B_sW1WAFPS0_2),.clk(gclk));
	jdff dff_B_CqnvPrmL2_2(.din(w_dff_B_sW1WAFPS0_2),.dout(w_dff_B_CqnvPrmL2_2),.clk(gclk));
	jdff dff_B_D50kcWaK7_2(.din(w_dff_B_CqnvPrmL2_2),.dout(w_dff_B_D50kcWaK7_2),.clk(gclk));
	jdff dff_B_zrgel2Dy4_2(.din(w_dff_B_D50kcWaK7_2),.dout(w_dff_B_zrgel2Dy4_2),.clk(gclk));
	jdff dff_B_4vwQvhhj3_2(.din(w_dff_B_zrgel2Dy4_2),.dout(w_dff_B_4vwQvhhj3_2),.clk(gclk));
	jdff dff_B_YxucSGjf8_2(.din(w_dff_B_4vwQvhhj3_2),.dout(w_dff_B_YxucSGjf8_2),.clk(gclk));
	jdff dff_B_qZMGiOAX5_2(.din(w_dff_B_YxucSGjf8_2),.dout(w_dff_B_qZMGiOAX5_2),.clk(gclk));
	jdff dff_B_TBWixOTo6_2(.din(w_dff_B_qZMGiOAX5_2),.dout(w_dff_B_TBWixOTo6_2),.clk(gclk));
	jdff dff_B_wDv85QkS5_2(.din(w_dff_B_TBWixOTo6_2),.dout(w_dff_B_wDv85QkS5_2),.clk(gclk));
	jdff dff_B_emq3D8w50_2(.din(w_dff_B_wDv85QkS5_2),.dout(w_dff_B_emq3D8w50_2),.clk(gclk));
	jdff dff_B_syYZUY0t3_2(.din(w_dff_B_emq3D8w50_2),.dout(w_dff_B_syYZUY0t3_2),.clk(gclk));
	jdff dff_B_jmb5iSCv1_2(.din(w_dff_B_syYZUY0t3_2),.dout(w_dff_B_jmb5iSCv1_2),.clk(gclk));
	jdff dff_B_eBgt6N6R7_2(.din(w_dff_B_jmb5iSCv1_2),.dout(w_dff_B_eBgt6N6R7_2),.clk(gclk));
	jdff dff_B_iuYDfpUc6_2(.din(w_dff_B_eBgt6N6R7_2),.dout(w_dff_B_iuYDfpUc6_2),.clk(gclk));
	jdff dff_B_nEfFQ1Go9_2(.din(w_dff_B_iuYDfpUc6_2),.dout(w_dff_B_nEfFQ1Go9_2),.clk(gclk));
	jdff dff_B_3Dsugy110_2(.din(w_dff_B_nEfFQ1Go9_2),.dout(w_dff_B_3Dsugy110_2),.clk(gclk));
	jdff dff_B_hVQDOkSS3_2(.din(w_dff_B_3Dsugy110_2),.dout(w_dff_B_hVQDOkSS3_2),.clk(gclk));
	jdff dff_B_yxiWYFnD1_2(.din(w_dff_B_hVQDOkSS3_2),.dout(w_dff_B_yxiWYFnD1_2),.clk(gclk));
	jdff dff_B_vzjEJ0329_2(.din(w_dff_B_yxiWYFnD1_2),.dout(w_dff_B_vzjEJ0329_2),.clk(gclk));
	jdff dff_B_MkDHctiK9_1(.din(n1044),.dout(w_dff_B_MkDHctiK9_1),.clk(gclk));
	jdff dff_B_n9jsUks89_2(.din(n944),.dout(w_dff_B_n9jsUks89_2),.clk(gclk));
	jdff dff_B_k7slm72j0_2(.din(w_dff_B_n9jsUks89_2),.dout(w_dff_B_k7slm72j0_2),.clk(gclk));
	jdff dff_B_9RyLp5TZ7_2(.din(w_dff_B_k7slm72j0_2),.dout(w_dff_B_9RyLp5TZ7_2),.clk(gclk));
	jdff dff_B_M3tKHR808_2(.din(w_dff_B_9RyLp5TZ7_2),.dout(w_dff_B_M3tKHR808_2),.clk(gclk));
	jdff dff_B_xMlmvkvB0_2(.din(w_dff_B_M3tKHR808_2),.dout(w_dff_B_xMlmvkvB0_2),.clk(gclk));
	jdff dff_B_Ue5FMrYX7_2(.din(w_dff_B_xMlmvkvB0_2),.dout(w_dff_B_Ue5FMrYX7_2),.clk(gclk));
	jdff dff_B_HwXYzmyU7_2(.din(w_dff_B_Ue5FMrYX7_2),.dout(w_dff_B_HwXYzmyU7_2),.clk(gclk));
	jdff dff_B_cqgbEvwX6_2(.din(w_dff_B_HwXYzmyU7_2),.dout(w_dff_B_cqgbEvwX6_2),.clk(gclk));
	jdff dff_B_xjRsQbBv0_2(.din(w_dff_B_cqgbEvwX6_2),.dout(w_dff_B_xjRsQbBv0_2),.clk(gclk));
	jdff dff_B_9ustTMDn8_2(.din(w_dff_B_xjRsQbBv0_2),.dout(w_dff_B_9ustTMDn8_2),.clk(gclk));
	jdff dff_B_g6wcwBbm0_2(.din(w_dff_B_9ustTMDn8_2),.dout(w_dff_B_g6wcwBbm0_2),.clk(gclk));
	jdff dff_B_MLbn53373_2(.din(w_dff_B_g6wcwBbm0_2),.dout(w_dff_B_MLbn53373_2),.clk(gclk));
	jdff dff_B_EdpKmaZt9_2(.din(w_dff_B_MLbn53373_2),.dout(w_dff_B_EdpKmaZt9_2),.clk(gclk));
	jdff dff_B_bR52msFv3_2(.din(w_dff_B_EdpKmaZt9_2),.dout(w_dff_B_bR52msFv3_2),.clk(gclk));
	jdff dff_B_JmZUqjjP3_2(.din(w_dff_B_bR52msFv3_2),.dout(w_dff_B_JmZUqjjP3_2),.clk(gclk));
	jdff dff_B_avDZQ1ym1_2(.din(w_dff_B_JmZUqjjP3_2),.dout(w_dff_B_avDZQ1ym1_2),.clk(gclk));
	jdff dff_B_vbwOjNoj6_2(.din(w_dff_B_avDZQ1ym1_2),.dout(w_dff_B_vbwOjNoj6_2),.clk(gclk));
	jdff dff_B_eXa8awt02_2(.din(w_dff_B_vbwOjNoj6_2),.dout(w_dff_B_eXa8awt02_2),.clk(gclk));
	jdff dff_B_iDvLRFo35_2(.din(w_dff_B_eXa8awt02_2),.dout(w_dff_B_iDvLRFo35_2),.clk(gclk));
	jdff dff_B_M9eT0cLQ5_2(.din(w_dff_B_iDvLRFo35_2),.dout(w_dff_B_M9eT0cLQ5_2),.clk(gclk));
	jdff dff_B_N1mDFkm30_1(.din(n945),.dout(w_dff_B_N1mDFkm30_1),.clk(gclk));
	jdff dff_B_SZFPGhcw5_2(.din(n842),.dout(w_dff_B_SZFPGhcw5_2),.clk(gclk));
	jdff dff_B_GLOgjmtE3_2(.din(w_dff_B_SZFPGhcw5_2),.dout(w_dff_B_GLOgjmtE3_2),.clk(gclk));
	jdff dff_B_mb2sjTnx7_2(.din(w_dff_B_GLOgjmtE3_2),.dout(w_dff_B_mb2sjTnx7_2),.clk(gclk));
	jdff dff_B_sBmDC3pi0_2(.din(w_dff_B_mb2sjTnx7_2),.dout(w_dff_B_sBmDC3pi0_2),.clk(gclk));
	jdff dff_B_5oJ2qCnK8_2(.din(w_dff_B_sBmDC3pi0_2),.dout(w_dff_B_5oJ2qCnK8_2),.clk(gclk));
	jdff dff_B_f2vb1aiX9_2(.din(w_dff_B_5oJ2qCnK8_2),.dout(w_dff_B_f2vb1aiX9_2),.clk(gclk));
	jdff dff_B_zzTTdMZO1_2(.din(w_dff_B_f2vb1aiX9_2),.dout(w_dff_B_zzTTdMZO1_2),.clk(gclk));
	jdff dff_B_xSClVX798_2(.din(w_dff_B_zzTTdMZO1_2),.dout(w_dff_B_xSClVX798_2),.clk(gclk));
	jdff dff_B_VdZFHFro3_2(.din(w_dff_B_xSClVX798_2),.dout(w_dff_B_VdZFHFro3_2),.clk(gclk));
	jdff dff_B_7Ple399Z8_2(.din(w_dff_B_VdZFHFro3_2),.dout(w_dff_B_7Ple399Z8_2),.clk(gclk));
	jdff dff_B_M9iIYBxB7_2(.din(w_dff_B_7Ple399Z8_2),.dout(w_dff_B_M9iIYBxB7_2),.clk(gclk));
	jdff dff_B_KFdhiOFG1_2(.din(w_dff_B_M9iIYBxB7_2),.dout(w_dff_B_KFdhiOFG1_2),.clk(gclk));
	jdff dff_B_c1vI4eX01_2(.din(w_dff_B_KFdhiOFG1_2),.dout(w_dff_B_c1vI4eX01_2),.clk(gclk));
	jdff dff_B_kAfTQgna7_2(.din(w_dff_B_c1vI4eX01_2),.dout(w_dff_B_kAfTQgna7_2),.clk(gclk));
	jdff dff_B_fs7Orvfl1_2(.din(w_dff_B_kAfTQgna7_2),.dout(w_dff_B_fs7Orvfl1_2),.clk(gclk));
	jdff dff_B_LGWKeNzZ6_2(.din(w_dff_B_fs7Orvfl1_2),.dout(w_dff_B_LGWKeNzZ6_2),.clk(gclk));
	jdff dff_B_EX2uFdos1_2(.din(w_dff_B_LGWKeNzZ6_2),.dout(w_dff_B_EX2uFdos1_2),.clk(gclk));
	jdff dff_B_pHEqSSlV6_2(.din(w_dff_B_EX2uFdos1_2),.dout(w_dff_B_pHEqSSlV6_2),.clk(gclk));
	jdff dff_B_ve9g9IJh7_1(.din(n843),.dout(w_dff_B_ve9g9IJh7_1),.clk(gclk));
	jdff dff_B_tdFI5j512_2(.din(n744),.dout(w_dff_B_tdFI5j512_2),.clk(gclk));
	jdff dff_B_ChzGEBgH6_2(.din(w_dff_B_tdFI5j512_2),.dout(w_dff_B_ChzGEBgH6_2),.clk(gclk));
	jdff dff_B_fFnX7s5g8_2(.din(w_dff_B_ChzGEBgH6_2),.dout(w_dff_B_fFnX7s5g8_2),.clk(gclk));
	jdff dff_B_rIV2zthO5_2(.din(w_dff_B_fFnX7s5g8_2),.dout(w_dff_B_rIV2zthO5_2),.clk(gclk));
	jdff dff_B_HdPFFl2T7_2(.din(w_dff_B_rIV2zthO5_2),.dout(w_dff_B_HdPFFl2T7_2),.clk(gclk));
	jdff dff_B_sspUpihD2_2(.din(w_dff_B_HdPFFl2T7_2),.dout(w_dff_B_sspUpihD2_2),.clk(gclk));
	jdff dff_B_BvoygqHS8_2(.din(w_dff_B_sspUpihD2_2),.dout(w_dff_B_BvoygqHS8_2),.clk(gclk));
	jdff dff_B_xG4vfSU18_2(.din(w_dff_B_BvoygqHS8_2),.dout(w_dff_B_xG4vfSU18_2),.clk(gclk));
	jdff dff_B_VdNyaOtG2_2(.din(w_dff_B_xG4vfSU18_2),.dout(w_dff_B_VdNyaOtG2_2),.clk(gclk));
	jdff dff_B_Y8SZASBv8_2(.din(w_dff_B_VdNyaOtG2_2),.dout(w_dff_B_Y8SZASBv8_2),.clk(gclk));
	jdff dff_B_inuMOoXO9_2(.din(w_dff_B_Y8SZASBv8_2),.dout(w_dff_B_inuMOoXO9_2),.clk(gclk));
	jdff dff_B_5n7KzOh11_2(.din(w_dff_B_inuMOoXO9_2),.dout(w_dff_B_5n7KzOh11_2),.clk(gclk));
	jdff dff_B_Im5zIJB11_2(.din(w_dff_B_5n7KzOh11_2),.dout(w_dff_B_Im5zIJB11_2),.clk(gclk));
	jdff dff_B_QbO8q9Q09_2(.din(w_dff_B_Im5zIJB11_2),.dout(w_dff_B_QbO8q9Q09_2),.clk(gclk));
	jdff dff_B_UM1nxNZv0_2(.din(w_dff_B_QbO8q9Q09_2),.dout(w_dff_B_UM1nxNZv0_2),.clk(gclk));
	jdff dff_B_ej1hnLyh5_2(.din(w_dff_B_UM1nxNZv0_2),.dout(w_dff_B_ej1hnLyh5_2),.clk(gclk));
	jdff dff_B_2a025RzN9_1(.din(n745),.dout(w_dff_B_2a025RzN9_1),.clk(gclk));
	jdff dff_B_zHOavq1r9_2(.din(n652),.dout(w_dff_B_zHOavq1r9_2),.clk(gclk));
	jdff dff_B_7w0CKtHm8_2(.din(w_dff_B_zHOavq1r9_2),.dout(w_dff_B_7w0CKtHm8_2),.clk(gclk));
	jdff dff_B_wZOorxwm3_2(.din(w_dff_B_7w0CKtHm8_2),.dout(w_dff_B_wZOorxwm3_2),.clk(gclk));
	jdff dff_B_D3blI8sS7_2(.din(w_dff_B_wZOorxwm3_2),.dout(w_dff_B_D3blI8sS7_2),.clk(gclk));
	jdff dff_B_TdeFe2XB0_2(.din(w_dff_B_D3blI8sS7_2),.dout(w_dff_B_TdeFe2XB0_2),.clk(gclk));
	jdff dff_B_hvpPu6Ru7_2(.din(w_dff_B_TdeFe2XB0_2),.dout(w_dff_B_hvpPu6Ru7_2),.clk(gclk));
	jdff dff_B_UdRzhJVA8_2(.din(w_dff_B_hvpPu6Ru7_2),.dout(w_dff_B_UdRzhJVA8_2),.clk(gclk));
	jdff dff_B_mF9M2XuR7_2(.din(w_dff_B_UdRzhJVA8_2),.dout(w_dff_B_mF9M2XuR7_2),.clk(gclk));
	jdff dff_B_dXdjQlLA2_2(.din(w_dff_B_mF9M2XuR7_2),.dout(w_dff_B_dXdjQlLA2_2),.clk(gclk));
	jdff dff_B_pSK8wpHS9_2(.din(w_dff_B_dXdjQlLA2_2),.dout(w_dff_B_pSK8wpHS9_2),.clk(gclk));
	jdff dff_B_i7HXVwUz8_2(.din(w_dff_B_pSK8wpHS9_2),.dout(w_dff_B_i7HXVwUz8_2),.clk(gclk));
	jdff dff_B_3wFakej16_2(.din(w_dff_B_i7HXVwUz8_2),.dout(w_dff_B_3wFakej16_2),.clk(gclk));
	jdff dff_B_mRDtuQqn9_2(.din(w_dff_B_3wFakej16_2),.dout(w_dff_B_mRDtuQqn9_2),.clk(gclk));
	jdff dff_B_jbGt7EVX8_2(.din(w_dff_B_mRDtuQqn9_2),.dout(w_dff_B_jbGt7EVX8_2),.clk(gclk));
	jdff dff_B_SqHIZXkK4_1(.din(n653),.dout(w_dff_B_SqHIZXkK4_1),.clk(gclk));
	jdff dff_B_3ejax37o8_2(.din(n567),.dout(w_dff_B_3ejax37o8_2),.clk(gclk));
	jdff dff_B_kQXBoYYd9_2(.din(w_dff_B_3ejax37o8_2),.dout(w_dff_B_kQXBoYYd9_2),.clk(gclk));
	jdff dff_B_DHpCnyVw3_2(.din(w_dff_B_kQXBoYYd9_2),.dout(w_dff_B_DHpCnyVw3_2),.clk(gclk));
	jdff dff_B_j1iZgJm40_2(.din(w_dff_B_DHpCnyVw3_2),.dout(w_dff_B_j1iZgJm40_2),.clk(gclk));
	jdff dff_B_nrbmUWzl7_2(.din(w_dff_B_j1iZgJm40_2),.dout(w_dff_B_nrbmUWzl7_2),.clk(gclk));
	jdff dff_B_jTnUMRra7_2(.din(w_dff_B_nrbmUWzl7_2),.dout(w_dff_B_jTnUMRra7_2),.clk(gclk));
	jdff dff_B_cuQh6nq22_2(.din(w_dff_B_jTnUMRra7_2),.dout(w_dff_B_cuQh6nq22_2),.clk(gclk));
	jdff dff_B_RGnWy5n37_2(.din(w_dff_B_cuQh6nq22_2),.dout(w_dff_B_RGnWy5n37_2),.clk(gclk));
	jdff dff_B_d8n4TBcx5_2(.din(w_dff_B_RGnWy5n37_2),.dout(w_dff_B_d8n4TBcx5_2),.clk(gclk));
	jdff dff_B_2oWBBBKG2_2(.din(w_dff_B_d8n4TBcx5_2),.dout(w_dff_B_2oWBBBKG2_2),.clk(gclk));
	jdff dff_B_AIUdJpQ50_2(.din(w_dff_B_2oWBBBKG2_2),.dout(w_dff_B_AIUdJpQ50_2),.clk(gclk));
	jdff dff_B_55nlJBQr7_2(.din(w_dff_B_AIUdJpQ50_2),.dout(w_dff_B_55nlJBQr7_2),.clk(gclk));
	jdff dff_B_vx7Y6eO44_1(.din(n568),.dout(w_dff_B_vx7Y6eO44_1),.clk(gclk));
	jdff dff_B_6TFfjaJL1_2(.din(n489),.dout(w_dff_B_6TFfjaJL1_2),.clk(gclk));
	jdff dff_B_ArwKlyIB6_2(.din(w_dff_B_6TFfjaJL1_2),.dout(w_dff_B_ArwKlyIB6_2),.clk(gclk));
	jdff dff_B_ZFTwEkfj3_2(.din(w_dff_B_ArwKlyIB6_2),.dout(w_dff_B_ZFTwEkfj3_2),.clk(gclk));
	jdff dff_B_MuwePaIo5_2(.din(w_dff_B_ZFTwEkfj3_2),.dout(w_dff_B_MuwePaIo5_2),.clk(gclk));
	jdff dff_B_I7DNNgbm7_2(.din(w_dff_B_MuwePaIo5_2),.dout(w_dff_B_I7DNNgbm7_2),.clk(gclk));
	jdff dff_B_S7AZXOhM1_2(.din(w_dff_B_I7DNNgbm7_2),.dout(w_dff_B_S7AZXOhM1_2),.clk(gclk));
	jdff dff_B_sxVOcIA26_2(.din(w_dff_B_S7AZXOhM1_2),.dout(w_dff_B_sxVOcIA26_2),.clk(gclk));
	jdff dff_B_VBDX5PDy4_2(.din(w_dff_B_sxVOcIA26_2),.dout(w_dff_B_VBDX5PDy4_2),.clk(gclk));
	jdff dff_B_ng7WXPmM5_2(.din(w_dff_B_VBDX5PDy4_2),.dout(w_dff_B_ng7WXPmM5_2),.clk(gclk));
	jdff dff_B_axgwUMrn3_2(.din(w_dff_B_ng7WXPmM5_2),.dout(w_dff_B_axgwUMrn3_2),.clk(gclk));
	jdff dff_B_i45uaWzw6_1(.din(n490),.dout(w_dff_B_i45uaWzw6_1),.clk(gclk));
	jdff dff_B_wGhaQFtC5_2(.din(n418),.dout(w_dff_B_wGhaQFtC5_2),.clk(gclk));
	jdff dff_B_ZVhZyt6A6_2(.din(w_dff_B_wGhaQFtC5_2),.dout(w_dff_B_ZVhZyt6A6_2),.clk(gclk));
	jdff dff_B_dUocCLtD0_2(.din(w_dff_B_ZVhZyt6A6_2),.dout(w_dff_B_dUocCLtD0_2),.clk(gclk));
	jdff dff_B_nEblCyuF6_2(.din(w_dff_B_dUocCLtD0_2),.dout(w_dff_B_nEblCyuF6_2),.clk(gclk));
	jdff dff_B_Tvwx1Hh83_2(.din(w_dff_B_nEblCyuF6_2),.dout(w_dff_B_Tvwx1Hh83_2),.clk(gclk));
	jdff dff_B_ydDJ2MsK4_2(.din(w_dff_B_Tvwx1Hh83_2),.dout(w_dff_B_ydDJ2MsK4_2),.clk(gclk));
	jdff dff_B_hkWByp8s3_2(.din(w_dff_B_ydDJ2MsK4_2),.dout(w_dff_B_hkWByp8s3_2),.clk(gclk));
	jdff dff_B_2l0AIDKB1_2(.din(w_dff_B_hkWByp8s3_2),.dout(w_dff_B_2l0AIDKB1_2),.clk(gclk));
	jdff dff_B_d3jWtuDe0_2(.din(n433),.dout(w_dff_B_d3jWtuDe0_2),.clk(gclk));
	jdff dff_B_abVjiXtl9_2(.din(w_dff_B_d3jWtuDe0_2),.dout(w_dff_B_abVjiXtl9_2),.clk(gclk));
	jdff dff_B_NqcXKRfB2_2(.din(w_dff_B_abVjiXtl9_2),.dout(w_dff_B_NqcXKRfB2_2),.clk(gclk));
	jdff dff_B_dPym85Zo9_1(.din(n419),.dout(w_dff_B_dPym85Zo9_1),.clk(gclk));
	jdff dff_B_9uF4WiNa0_1(.din(w_dff_B_dPym85Zo9_1),.dout(w_dff_B_9uF4WiNa0_1),.clk(gclk));
	jdff dff_B_FriOFbtv9_1(.din(w_dff_B_9uF4WiNa0_1),.dout(w_dff_B_FriOFbtv9_1),.clk(gclk));
	jdff dff_B_g1z8XKt61_2(.din(n356),.dout(w_dff_B_g1z8XKt61_2),.clk(gclk));
	jdff dff_B_AmXH2p9Z4_2(.din(w_dff_B_g1z8XKt61_2),.dout(w_dff_B_AmXH2p9Z4_2),.clk(gclk));
	jdff dff_B_fhv5ubir5_2(.din(w_dff_B_AmXH2p9Z4_2),.dout(w_dff_B_fhv5ubir5_2),.clk(gclk));
	jdff dff_B_WnY7mpGK0_0(.din(n361),.dout(w_dff_B_WnY7mpGK0_0),.clk(gclk));
	jdff dff_B_YuU6LOnn8_0(.din(w_dff_B_WnY7mpGK0_0),.dout(w_dff_B_YuU6LOnn8_0),.clk(gclk));
	jdff dff_A_deehWp9L1_0(.dout(w_n297_0[0]),.din(w_dff_A_deehWp9L1_0),.clk(gclk));
	jdff dff_A_i0usyGzS7_0(.dout(w_dff_A_deehWp9L1_0),.din(w_dff_A_i0usyGzS7_0),.clk(gclk));
	jdff dff_A_3nZsfIXV0_1(.dout(w_n297_0[1]),.din(w_dff_A_3nZsfIXV0_1),.clk(gclk));
	jdff dff_A_q2evcYDZ5_1(.dout(w_dff_A_3nZsfIXV0_1),.din(w_dff_A_q2evcYDZ5_1),.clk(gclk));
	jdff dff_B_vcEbTGsI3_2(.din(n1596),.dout(w_dff_B_vcEbTGsI3_2),.clk(gclk));
	jdff dff_B_lFsWGR3P7_2(.din(w_dff_B_vcEbTGsI3_2),.dout(w_dff_B_lFsWGR3P7_2),.clk(gclk));
	jdff dff_B_4BsIzBMw6_1(.din(n1594),.dout(w_dff_B_4BsIzBMw6_1),.clk(gclk));
	jdff dff_B_HxXebcxg5_2(.din(n1535),.dout(w_dff_B_HxXebcxg5_2),.clk(gclk));
	jdff dff_B_WP1rxRCJ5_2(.din(w_dff_B_HxXebcxg5_2),.dout(w_dff_B_WP1rxRCJ5_2),.clk(gclk));
	jdff dff_B_Yf1v076c4_2(.din(w_dff_B_WP1rxRCJ5_2),.dout(w_dff_B_Yf1v076c4_2),.clk(gclk));
	jdff dff_B_hUP16nCm6_2(.din(w_dff_B_Yf1v076c4_2),.dout(w_dff_B_hUP16nCm6_2),.clk(gclk));
	jdff dff_B_Vj41LMhi1_2(.din(w_dff_B_hUP16nCm6_2),.dout(w_dff_B_Vj41LMhi1_2),.clk(gclk));
	jdff dff_B_dTTekMdM3_2(.din(w_dff_B_Vj41LMhi1_2),.dout(w_dff_B_dTTekMdM3_2),.clk(gclk));
	jdff dff_B_yyrGMbKm5_2(.din(w_dff_B_dTTekMdM3_2),.dout(w_dff_B_yyrGMbKm5_2),.clk(gclk));
	jdff dff_B_3qqGqiIU2_2(.din(w_dff_B_yyrGMbKm5_2),.dout(w_dff_B_3qqGqiIU2_2),.clk(gclk));
	jdff dff_B_Thp5r74E6_2(.din(w_dff_B_3qqGqiIU2_2),.dout(w_dff_B_Thp5r74E6_2),.clk(gclk));
	jdff dff_B_Mby9w92n0_2(.din(w_dff_B_Thp5r74E6_2),.dout(w_dff_B_Mby9w92n0_2),.clk(gclk));
	jdff dff_B_MFuCVV3z0_2(.din(w_dff_B_Mby9w92n0_2),.dout(w_dff_B_MFuCVV3z0_2),.clk(gclk));
	jdff dff_B_mGugFnAj8_2(.din(w_dff_B_MFuCVV3z0_2),.dout(w_dff_B_mGugFnAj8_2),.clk(gclk));
	jdff dff_B_GVrmcoad6_2(.din(w_dff_B_mGugFnAj8_2),.dout(w_dff_B_GVrmcoad6_2),.clk(gclk));
	jdff dff_B_XZuJnthB2_2(.din(w_dff_B_GVrmcoad6_2),.dout(w_dff_B_XZuJnthB2_2),.clk(gclk));
	jdff dff_B_ThixVkvE8_2(.din(w_dff_B_XZuJnthB2_2),.dout(w_dff_B_ThixVkvE8_2),.clk(gclk));
	jdff dff_B_UNNmP23o0_2(.din(w_dff_B_ThixVkvE8_2),.dout(w_dff_B_UNNmP23o0_2),.clk(gclk));
	jdff dff_B_vaXIHUKE7_2(.din(w_dff_B_UNNmP23o0_2),.dout(w_dff_B_vaXIHUKE7_2),.clk(gclk));
	jdff dff_B_Qo6fIxKZ0_2(.din(w_dff_B_vaXIHUKE7_2),.dout(w_dff_B_Qo6fIxKZ0_2),.clk(gclk));
	jdff dff_B_2L78vnbn8_2(.din(w_dff_B_Qo6fIxKZ0_2),.dout(w_dff_B_2L78vnbn8_2),.clk(gclk));
	jdff dff_B_YtP7SnK81_2(.din(w_dff_B_2L78vnbn8_2),.dout(w_dff_B_YtP7SnK81_2),.clk(gclk));
	jdff dff_B_xNPo3ieC2_2(.din(w_dff_B_YtP7SnK81_2),.dout(w_dff_B_xNPo3ieC2_2),.clk(gclk));
	jdff dff_B_Ui3D5MDp5_2(.din(w_dff_B_xNPo3ieC2_2),.dout(w_dff_B_Ui3D5MDp5_2),.clk(gclk));
	jdff dff_B_4je9YzJo3_2(.din(w_dff_B_Ui3D5MDp5_2),.dout(w_dff_B_4je9YzJo3_2),.clk(gclk));
	jdff dff_B_efMuE7CX6_2(.din(w_dff_B_4je9YzJo3_2),.dout(w_dff_B_efMuE7CX6_2),.clk(gclk));
	jdff dff_B_ecrc3ieh1_2(.din(w_dff_B_efMuE7CX6_2),.dout(w_dff_B_ecrc3ieh1_2),.clk(gclk));
	jdff dff_B_wpLvLIuC4_2(.din(w_dff_B_ecrc3ieh1_2),.dout(w_dff_B_wpLvLIuC4_2),.clk(gclk));
	jdff dff_B_pKdxKnsb3_2(.din(w_dff_B_wpLvLIuC4_2),.dout(w_dff_B_pKdxKnsb3_2),.clk(gclk));
	jdff dff_B_ihlCNmq73_2(.din(w_dff_B_pKdxKnsb3_2),.dout(w_dff_B_ihlCNmq73_2),.clk(gclk));
	jdff dff_B_kqhi5uqQ2_2(.din(w_dff_B_ihlCNmq73_2),.dout(w_dff_B_kqhi5uqQ2_2),.clk(gclk));
	jdff dff_B_OIOSvCgg7_2(.din(w_dff_B_kqhi5uqQ2_2),.dout(w_dff_B_OIOSvCgg7_2),.clk(gclk));
	jdff dff_B_ORssjp738_2(.din(w_dff_B_OIOSvCgg7_2),.dout(w_dff_B_ORssjp738_2),.clk(gclk));
	jdff dff_B_roNJYT814_2(.din(w_dff_B_ORssjp738_2),.dout(w_dff_B_roNJYT814_2),.clk(gclk));
	jdff dff_B_2E8EtbSU8_2(.din(w_dff_B_roNJYT814_2),.dout(w_dff_B_2E8EtbSU8_2),.clk(gclk));
	jdff dff_B_XLsmYfGI7_2(.din(w_dff_B_2E8EtbSU8_2),.dout(w_dff_B_XLsmYfGI7_2),.clk(gclk));
	jdff dff_B_9VQXBh5r1_2(.din(w_dff_B_XLsmYfGI7_2),.dout(w_dff_B_9VQXBh5r1_2),.clk(gclk));
	jdff dff_B_CAQSRdEd6_2(.din(w_dff_B_9VQXBh5r1_2),.dout(w_dff_B_CAQSRdEd6_2),.clk(gclk));
	jdff dff_B_9XTlHHFv3_2(.din(w_dff_B_CAQSRdEd6_2),.dout(w_dff_B_9XTlHHFv3_2),.clk(gclk));
	jdff dff_B_vDgUCxtX0_1(.din(n1592),.dout(w_dff_B_vDgUCxtX0_1),.clk(gclk));
	jdff dff_A_v4JB5FpV2_1(.dout(w_n1538_0[1]),.din(w_dff_A_v4JB5FpV2_1),.clk(gclk));
	jdff dff_B_liHWSXZD3_1(.din(n1536),.dout(w_dff_B_liHWSXZD3_1),.clk(gclk));
	jdff dff_B_bIGjJxxb3_2(.din(n1471),.dout(w_dff_B_bIGjJxxb3_2),.clk(gclk));
	jdff dff_B_rXwZGBD63_2(.din(w_dff_B_bIGjJxxb3_2),.dout(w_dff_B_rXwZGBD63_2),.clk(gclk));
	jdff dff_B_WgiHGz0s8_2(.din(w_dff_B_rXwZGBD63_2),.dout(w_dff_B_WgiHGz0s8_2),.clk(gclk));
	jdff dff_B_rQdvQecD2_2(.din(w_dff_B_WgiHGz0s8_2),.dout(w_dff_B_rQdvQecD2_2),.clk(gclk));
	jdff dff_B_UPUZWbIe6_2(.din(w_dff_B_rQdvQecD2_2),.dout(w_dff_B_UPUZWbIe6_2),.clk(gclk));
	jdff dff_B_U0GE3S6W1_2(.din(w_dff_B_UPUZWbIe6_2),.dout(w_dff_B_U0GE3S6W1_2),.clk(gclk));
	jdff dff_B_KPzSsgjv0_2(.din(w_dff_B_U0GE3S6W1_2),.dout(w_dff_B_KPzSsgjv0_2),.clk(gclk));
	jdff dff_B_2rlnimY87_2(.din(w_dff_B_KPzSsgjv0_2),.dout(w_dff_B_2rlnimY87_2),.clk(gclk));
	jdff dff_B_3e3Cxr9A0_2(.din(w_dff_B_2rlnimY87_2),.dout(w_dff_B_3e3Cxr9A0_2),.clk(gclk));
	jdff dff_B_0yrACB2p8_2(.din(w_dff_B_3e3Cxr9A0_2),.dout(w_dff_B_0yrACB2p8_2),.clk(gclk));
	jdff dff_B_eRvYyFQ85_2(.din(w_dff_B_0yrACB2p8_2),.dout(w_dff_B_eRvYyFQ85_2),.clk(gclk));
	jdff dff_B_DBcj978o6_2(.din(w_dff_B_eRvYyFQ85_2),.dout(w_dff_B_DBcj978o6_2),.clk(gclk));
	jdff dff_B_FM96viRs2_2(.din(w_dff_B_DBcj978o6_2),.dout(w_dff_B_FM96viRs2_2),.clk(gclk));
	jdff dff_B_oMKWUdUF9_2(.din(w_dff_B_FM96viRs2_2),.dout(w_dff_B_oMKWUdUF9_2),.clk(gclk));
	jdff dff_B_dZprClE56_2(.din(w_dff_B_oMKWUdUF9_2),.dout(w_dff_B_dZprClE56_2),.clk(gclk));
	jdff dff_B_jz1lDOW31_2(.din(w_dff_B_dZprClE56_2),.dout(w_dff_B_jz1lDOW31_2),.clk(gclk));
	jdff dff_B_HzEPq7uv5_2(.din(w_dff_B_jz1lDOW31_2),.dout(w_dff_B_HzEPq7uv5_2),.clk(gclk));
	jdff dff_B_0POMQpTl9_2(.din(w_dff_B_HzEPq7uv5_2),.dout(w_dff_B_0POMQpTl9_2),.clk(gclk));
	jdff dff_B_ZgMhr7PX9_2(.din(w_dff_B_0POMQpTl9_2),.dout(w_dff_B_ZgMhr7PX9_2),.clk(gclk));
	jdff dff_B_4t2MH9Fy3_2(.din(w_dff_B_ZgMhr7PX9_2),.dout(w_dff_B_4t2MH9Fy3_2),.clk(gclk));
	jdff dff_B_5g1oNCoa5_2(.din(w_dff_B_4t2MH9Fy3_2),.dout(w_dff_B_5g1oNCoa5_2),.clk(gclk));
	jdff dff_B_WYoIOJ5w0_2(.din(w_dff_B_5g1oNCoa5_2),.dout(w_dff_B_WYoIOJ5w0_2),.clk(gclk));
	jdff dff_B_AUnmZvQP7_2(.din(w_dff_B_WYoIOJ5w0_2),.dout(w_dff_B_AUnmZvQP7_2),.clk(gclk));
	jdff dff_B_BCUUKeE94_2(.din(w_dff_B_AUnmZvQP7_2),.dout(w_dff_B_BCUUKeE94_2),.clk(gclk));
	jdff dff_B_NCWoOmXz5_2(.din(w_dff_B_BCUUKeE94_2),.dout(w_dff_B_NCWoOmXz5_2),.clk(gclk));
	jdff dff_B_tcSpubjx4_2(.din(w_dff_B_NCWoOmXz5_2),.dout(w_dff_B_tcSpubjx4_2),.clk(gclk));
	jdff dff_B_ahk9aaSS2_2(.din(w_dff_B_tcSpubjx4_2),.dout(w_dff_B_ahk9aaSS2_2),.clk(gclk));
	jdff dff_B_Cfb46NbZ0_2(.din(w_dff_B_ahk9aaSS2_2),.dout(w_dff_B_Cfb46NbZ0_2),.clk(gclk));
	jdff dff_B_3jrur08M2_2(.din(w_dff_B_Cfb46NbZ0_2),.dout(w_dff_B_3jrur08M2_2),.clk(gclk));
	jdff dff_B_guWsENKn1_2(.din(w_dff_B_3jrur08M2_2),.dout(w_dff_B_guWsENKn1_2),.clk(gclk));
	jdff dff_B_svpNUMGJ3_2(.din(w_dff_B_guWsENKn1_2),.dout(w_dff_B_svpNUMGJ3_2),.clk(gclk));
	jdff dff_B_vNogexnc8_2(.din(w_dff_B_svpNUMGJ3_2),.dout(w_dff_B_vNogexnc8_2),.clk(gclk));
	jdff dff_B_dmovVPEO7_2(.din(n1474),.dout(w_dff_B_dmovVPEO7_2),.clk(gclk));
	jdff dff_B_vbv4jbug2_1(.din(n1472),.dout(w_dff_B_vbv4jbug2_1),.clk(gclk));
	jdff dff_B_knh65Mub3_2(.din(n1400),.dout(w_dff_B_knh65Mub3_2),.clk(gclk));
	jdff dff_B_rtbfUa4N3_2(.din(w_dff_B_knh65Mub3_2),.dout(w_dff_B_rtbfUa4N3_2),.clk(gclk));
	jdff dff_B_yZfi7oZz8_2(.din(w_dff_B_rtbfUa4N3_2),.dout(w_dff_B_yZfi7oZz8_2),.clk(gclk));
	jdff dff_B_pHTBo1wK1_2(.din(w_dff_B_yZfi7oZz8_2),.dout(w_dff_B_pHTBo1wK1_2),.clk(gclk));
	jdff dff_B_FKJmDMMY6_2(.din(w_dff_B_pHTBo1wK1_2),.dout(w_dff_B_FKJmDMMY6_2),.clk(gclk));
	jdff dff_B_wO0lpCBD3_2(.din(w_dff_B_FKJmDMMY6_2),.dout(w_dff_B_wO0lpCBD3_2),.clk(gclk));
	jdff dff_B_ACzMNpoF2_2(.din(w_dff_B_wO0lpCBD3_2),.dout(w_dff_B_ACzMNpoF2_2),.clk(gclk));
	jdff dff_B_dXGolllw6_2(.din(w_dff_B_ACzMNpoF2_2),.dout(w_dff_B_dXGolllw6_2),.clk(gclk));
	jdff dff_B_4GtaH4zl4_2(.din(w_dff_B_dXGolllw6_2),.dout(w_dff_B_4GtaH4zl4_2),.clk(gclk));
	jdff dff_B_6KZDl10G0_2(.din(w_dff_B_4GtaH4zl4_2),.dout(w_dff_B_6KZDl10G0_2),.clk(gclk));
	jdff dff_B_Zeq3fLLW5_2(.din(w_dff_B_6KZDl10G0_2),.dout(w_dff_B_Zeq3fLLW5_2),.clk(gclk));
	jdff dff_B_Vt5KTL0r0_2(.din(w_dff_B_Zeq3fLLW5_2),.dout(w_dff_B_Vt5KTL0r0_2),.clk(gclk));
	jdff dff_B_pUeBZUWe6_2(.din(w_dff_B_Vt5KTL0r0_2),.dout(w_dff_B_pUeBZUWe6_2),.clk(gclk));
	jdff dff_B_jUJvx4VH5_2(.din(w_dff_B_pUeBZUWe6_2),.dout(w_dff_B_jUJvx4VH5_2),.clk(gclk));
	jdff dff_B_nhokQXfo1_2(.din(w_dff_B_jUJvx4VH5_2),.dout(w_dff_B_nhokQXfo1_2),.clk(gclk));
	jdff dff_B_QCeetsf33_2(.din(w_dff_B_nhokQXfo1_2),.dout(w_dff_B_QCeetsf33_2),.clk(gclk));
	jdff dff_B_zNTkDR803_2(.din(w_dff_B_QCeetsf33_2),.dout(w_dff_B_zNTkDR803_2),.clk(gclk));
	jdff dff_B_v8vEdzaX0_2(.din(w_dff_B_zNTkDR803_2),.dout(w_dff_B_v8vEdzaX0_2),.clk(gclk));
	jdff dff_B_nYgwjDA91_2(.din(w_dff_B_v8vEdzaX0_2),.dout(w_dff_B_nYgwjDA91_2),.clk(gclk));
	jdff dff_B_P00oN6iR2_2(.din(w_dff_B_nYgwjDA91_2),.dout(w_dff_B_P00oN6iR2_2),.clk(gclk));
	jdff dff_B_9XN3JhzY1_2(.din(w_dff_B_P00oN6iR2_2),.dout(w_dff_B_9XN3JhzY1_2),.clk(gclk));
	jdff dff_B_RCRf1bmH3_2(.din(w_dff_B_9XN3JhzY1_2),.dout(w_dff_B_RCRf1bmH3_2),.clk(gclk));
	jdff dff_B_ljr7OGIX8_2(.din(w_dff_B_RCRf1bmH3_2),.dout(w_dff_B_ljr7OGIX8_2),.clk(gclk));
	jdff dff_B_0eOHq9LC7_2(.din(w_dff_B_ljr7OGIX8_2),.dout(w_dff_B_0eOHq9LC7_2),.clk(gclk));
	jdff dff_B_XPhQYgMY8_2(.din(w_dff_B_0eOHq9LC7_2),.dout(w_dff_B_XPhQYgMY8_2),.clk(gclk));
	jdff dff_B_nrTVaabD0_2(.din(w_dff_B_XPhQYgMY8_2),.dout(w_dff_B_nrTVaabD0_2),.clk(gclk));
	jdff dff_B_tc8xiSLQ0_2(.din(w_dff_B_nrTVaabD0_2),.dout(w_dff_B_tc8xiSLQ0_2),.clk(gclk));
	jdff dff_B_eJQXBWSO6_2(.din(w_dff_B_tc8xiSLQ0_2),.dout(w_dff_B_eJQXBWSO6_2),.clk(gclk));
	jdff dff_B_zVqLTIM78_2(.din(w_dff_B_eJQXBWSO6_2),.dout(w_dff_B_zVqLTIM78_2),.clk(gclk));
	jdff dff_B_ISmDjF5k2_2(.din(n1403),.dout(w_dff_B_ISmDjF5k2_2),.clk(gclk));
	jdff dff_B_tnlqCwf56_1(.din(n1401),.dout(w_dff_B_tnlqCwf56_1),.clk(gclk));
	jdff dff_B_Qj94JnIk7_2(.din(n1322),.dout(w_dff_B_Qj94JnIk7_2),.clk(gclk));
	jdff dff_B_9VoRz78x1_2(.din(w_dff_B_Qj94JnIk7_2),.dout(w_dff_B_9VoRz78x1_2),.clk(gclk));
	jdff dff_B_gBKYXQ4D7_2(.din(w_dff_B_9VoRz78x1_2),.dout(w_dff_B_gBKYXQ4D7_2),.clk(gclk));
	jdff dff_B_kG10tY4k1_2(.din(w_dff_B_gBKYXQ4D7_2),.dout(w_dff_B_kG10tY4k1_2),.clk(gclk));
	jdff dff_B_30qgJ2EH2_2(.din(w_dff_B_kG10tY4k1_2),.dout(w_dff_B_30qgJ2EH2_2),.clk(gclk));
	jdff dff_B_M4Z8Hivs2_2(.din(w_dff_B_30qgJ2EH2_2),.dout(w_dff_B_M4Z8Hivs2_2),.clk(gclk));
	jdff dff_B_F4KsOBJO1_2(.din(w_dff_B_M4Z8Hivs2_2),.dout(w_dff_B_F4KsOBJO1_2),.clk(gclk));
	jdff dff_B_QQnBUEyp3_2(.din(w_dff_B_F4KsOBJO1_2),.dout(w_dff_B_QQnBUEyp3_2),.clk(gclk));
	jdff dff_B_7ZfPdFRY5_2(.din(w_dff_B_QQnBUEyp3_2),.dout(w_dff_B_7ZfPdFRY5_2),.clk(gclk));
	jdff dff_B_J8dcXqrp4_2(.din(w_dff_B_7ZfPdFRY5_2),.dout(w_dff_B_J8dcXqrp4_2),.clk(gclk));
	jdff dff_B_R6o0VXny5_2(.din(w_dff_B_J8dcXqrp4_2),.dout(w_dff_B_R6o0VXny5_2),.clk(gclk));
	jdff dff_B_tafc9iqI9_2(.din(w_dff_B_R6o0VXny5_2),.dout(w_dff_B_tafc9iqI9_2),.clk(gclk));
	jdff dff_B_IzPDP5jB8_2(.din(w_dff_B_tafc9iqI9_2),.dout(w_dff_B_IzPDP5jB8_2),.clk(gclk));
	jdff dff_B_Pu03p8sT7_2(.din(w_dff_B_IzPDP5jB8_2),.dout(w_dff_B_Pu03p8sT7_2),.clk(gclk));
	jdff dff_B_Y16q20xC2_2(.din(w_dff_B_Pu03p8sT7_2),.dout(w_dff_B_Y16q20xC2_2),.clk(gclk));
	jdff dff_B_38saKqEP7_2(.din(w_dff_B_Y16q20xC2_2),.dout(w_dff_B_38saKqEP7_2),.clk(gclk));
	jdff dff_B_TPlCHBjx9_2(.din(w_dff_B_38saKqEP7_2),.dout(w_dff_B_TPlCHBjx9_2),.clk(gclk));
	jdff dff_B_lYFNPIfF0_2(.din(w_dff_B_TPlCHBjx9_2),.dout(w_dff_B_lYFNPIfF0_2),.clk(gclk));
	jdff dff_B_O6js9CB48_2(.din(w_dff_B_lYFNPIfF0_2),.dout(w_dff_B_O6js9CB48_2),.clk(gclk));
	jdff dff_B_Qp7ehhEF1_2(.din(w_dff_B_O6js9CB48_2),.dout(w_dff_B_Qp7ehhEF1_2),.clk(gclk));
	jdff dff_B_KKss5IRV7_2(.din(w_dff_B_Qp7ehhEF1_2),.dout(w_dff_B_KKss5IRV7_2),.clk(gclk));
	jdff dff_B_Ah2DniCw0_2(.din(w_dff_B_KKss5IRV7_2),.dout(w_dff_B_Ah2DniCw0_2),.clk(gclk));
	jdff dff_B_HnjCamSK3_2(.din(w_dff_B_Ah2DniCw0_2),.dout(w_dff_B_HnjCamSK3_2),.clk(gclk));
	jdff dff_B_igQdNCZt8_2(.din(w_dff_B_HnjCamSK3_2),.dout(w_dff_B_igQdNCZt8_2),.clk(gclk));
	jdff dff_B_pTLzZ28K6_2(.din(w_dff_B_igQdNCZt8_2),.dout(w_dff_B_pTLzZ28K6_2),.clk(gclk));
	jdff dff_B_8I3X7dEL7_2(.din(w_dff_B_pTLzZ28K6_2),.dout(w_dff_B_8I3X7dEL7_2),.clk(gclk));
	jdff dff_B_32Ixfw7Z1_1(.din(n1323),.dout(w_dff_B_32Ixfw7Z1_1),.clk(gclk));
	jdff dff_B_05gSVpdw3_2(.din(n1237),.dout(w_dff_B_05gSVpdw3_2),.clk(gclk));
	jdff dff_B_yIJGvAp85_2(.din(w_dff_B_05gSVpdw3_2),.dout(w_dff_B_yIJGvAp85_2),.clk(gclk));
	jdff dff_B_4sCuC4yF3_2(.din(w_dff_B_yIJGvAp85_2),.dout(w_dff_B_4sCuC4yF3_2),.clk(gclk));
	jdff dff_B_ZkSQfUkp6_2(.din(w_dff_B_4sCuC4yF3_2),.dout(w_dff_B_ZkSQfUkp6_2),.clk(gclk));
	jdff dff_B_WkxIbYJK8_2(.din(w_dff_B_ZkSQfUkp6_2),.dout(w_dff_B_WkxIbYJK8_2),.clk(gclk));
	jdff dff_B_1anvwL6R7_2(.din(w_dff_B_WkxIbYJK8_2),.dout(w_dff_B_1anvwL6R7_2),.clk(gclk));
	jdff dff_B_nKqflDpN1_2(.din(w_dff_B_1anvwL6R7_2),.dout(w_dff_B_nKqflDpN1_2),.clk(gclk));
	jdff dff_B_jai23uj43_2(.din(w_dff_B_nKqflDpN1_2),.dout(w_dff_B_jai23uj43_2),.clk(gclk));
	jdff dff_B_Y8NEOlcL3_2(.din(w_dff_B_jai23uj43_2),.dout(w_dff_B_Y8NEOlcL3_2),.clk(gclk));
	jdff dff_B_TWFxZrgN2_2(.din(w_dff_B_Y8NEOlcL3_2),.dout(w_dff_B_TWFxZrgN2_2),.clk(gclk));
	jdff dff_B_KpoPiNBM4_2(.din(w_dff_B_TWFxZrgN2_2),.dout(w_dff_B_KpoPiNBM4_2),.clk(gclk));
	jdff dff_B_jPO5Zibc1_2(.din(w_dff_B_KpoPiNBM4_2),.dout(w_dff_B_jPO5Zibc1_2),.clk(gclk));
	jdff dff_B_H3RETrgb0_2(.din(w_dff_B_jPO5Zibc1_2),.dout(w_dff_B_H3RETrgb0_2),.clk(gclk));
	jdff dff_B_nBP5DtAl5_2(.din(w_dff_B_H3RETrgb0_2),.dout(w_dff_B_nBP5DtAl5_2),.clk(gclk));
	jdff dff_B_AdWUsOxP8_2(.din(w_dff_B_nBP5DtAl5_2),.dout(w_dff_B_AdWUsOxP8_2),.clk(gclk));
	jdff dff_B_ufbezDiC3_2(.din(w_dff_B_AdWUsOxP8_2),.dout(w_dff_B_ufbezDiC3_2),.clk(gclk));
	jdff dff_B_1hqYdLjg5_2(.din(w_dff_B_ufbezDiC3_2),.dout(w_dff_B_1hqYdLjg5_2),.clk(gclk));
	jdff dff_B_QS1HdsCf1_2(.din(w_dff_B_1hqYdLjg5_2),.dout(w_dff_B_QS1HdsCf1_2),.clk(gclk));
	jdff dff_B_6qWUsFaA0_2(.din(w_dff_B_QS1HdsCf1_2),.dout(w_dff_B_6qWUsFaA0_2),.clk(gclk));
	jdff dff_B_kGukgcjl9_2(.din(w_dff_B_6qWUsFaA0_2),.dout(w_dff_B_kGukgcjl9_2),.clk(gclk));
	jdff dff_B_mxkdFD5P6_2(.din(w_dff_B_kGukgcjl9_2),.dout(w_dff_B_mxkdFD5P6_2),.clk(gclk));
	jdff dff_B_6n67HBBO9_2(.din(w_dff_B_mxkdFD5P6_2),.dout(w_dff_B_6n67HBBO9_2),.clk(gclk));
	jdff dff_B_3CjuWQ8Z6_2(.din(w_dff_B_6n67HBBO9_2),.dout(w_dff_B_3CjuWQ8Z6_2),.clk(gclk));
	jdff dff_B_NAXPIAqq6_2(.din(w_dff_B_3CjuWQ8Z6_2),.dout(w_dff_B_NAXPIAqq6_2),.clk(gclk));
	jdff dff_B_Q4Onb2760_1(.din(n1238),.dout(w_dff_B_Q4Onb2760_1),.clk(gclk));
	jdff dff_B_J1TpgkZa1_2(.din(n1146),.dout(w_dff_B_J1TpgkZa1_2),.clk(gclk));
	jdff dff_B_t54vy7cw7_2(.din(w_dff_B_J1TpgkZa1_2),.dout(w_dff_B_t54vy7cw7_2),.clk(gclk));
	jdff dff_B_DLSclZDo4_2(.din(w_dff_B_t54vy7cw7_2),.dout(w_dff_B_DLSclZDo4_2),.clk(gclk));
	jdff dff_B_7I7Xx8TQ5_2(.din(w_dff_B_DLSclZDo4_2),.dout(w_dff_B_7I7Xx8TQ5_2),.clk(gclk));
	jdff dff_B_U4z9WrT53_2(.din(w_dff_B_7I7Xx8TQ5_2),.dout(w_dff_B_U4z9WrT53_2),.clk(gclk));
	jdff dff_B_cPaktSpE2_2(.din(w_dff_B_U4z9WrT53_2),.dout(w_dff_B_cPaktSpE2_2),.clk(gclk));
	jdff dff_B_ckRVo5Xu4_2(.din(w_dff_B_cPaktSpE2_2),.dout(w_dff_B_ckRVo5Xu4_2),.clk(gclk));
	jdff dff_B_GBGJH0nS2_2(.din(w_dff_B_ckRVo5Xu4_2),.dout(w_dff_B_GBGJH0nS2_2),.clk(gclk));
	jdff dff_B_RnMAILM42_2(.din(w_dff_B_GBGJH0nS2_2),.dout(w_dff_B_RnMAILM42_2),.clk(gclk));
	jdff dff_B_cUtcAg0O3_2(.din(w_dff_B_RnMAILM42_2),.dout(w_dff_B_cUtcAg0O3_2),.clk(gclk));
	jdff dff_B_D5LXQRvh7_2(.din(w_dff_B_cUtcAg0O3_2),.dout(w_dff_B_D5LXQRvh7_2),.clk(gclk));
	jdff dff_B_U0q6GnRr9_2(.din(w_dff_B_D5LXQRvh7_2),.dout(w_dff_B_U0q6GnRr9_2),.clk(gclk));
	jdff dff_B_gtCuGuHR7_2(.din(w_dff_B_U0q6GnRr9_2),.dout(w_dff_B_gtCuGuHR7_2),.clk(gclk));
	jdff dff_B_tcemRyZ50_2(.din(w_dff_B_gtCuGuHR7_2),.dout(w_dff_B_tcemRyZ50_2),.clk(gclk));
	jdff dff_B_Xxend09L6_2(.din(w_dff_B_tcemRyZ50_2),.dout(w_dff_B_Xxend09L6_2),.clk(gclk));
	jdff dff_B_ths3gjrN0_2(.din(w_dff_B_Xxend09L6_2),.dout(w_dff_B_ths3gjrN0_2),.clk(gclk));
	jdff dff_B_5C92nWMz1_2(.din(w_dff_B_ths3gjrN0_2),.dout(w_dff_B_5C92nWMz1_2),.clk(gclk));
	jdff dff_B_Vk1ekSo52_2(.din(w_dff_B_5C92nWMz1_2),.dout(w_dff_B_Vk1ekSo52_2),.clk(gclk));
	jdff dff_B_UHr93JyK7_2(.din(w_dff_B_Vk1ekSo52_2),.dout(w_dff_B_UHr93JyK7_2),.clk(gclk));
	jdff dff_B_5vi4CxmF0_2(.din(w_dff_B_UHr93JyK7_2),.dout(w_dff_B_5vi4CxmF0_2),.clk(gclk));
	jdff dff_B_5QJ5XjO55_2(.din(w_dff_B_5vi4CxmF0_2),.dout(w_dff_B_5QJ5XjO55_2),.clk(gclk));
	jdff dff_B_tZNJFONl2_2(.din(w_dff_B_5QJ5XjO55_2),.dout(w_dff_B_tZNJFONl2_2),.clk(gclk));
	jdff dff_B_byEMZ9rd5_1(.din(n1147),.dout(w_dff_B_byEMZ9rd5_1),.clk(gclk));
	jdff dff_B_5FYseBB29_2(.din(n1048),.dout(w_dff_B_5FYseBB29_2),.clk(gclk));
	jdff dff_B_LiV73i203_2(.din(w_dff_B_5FYseBB29_2),.dout(w_dff_B_LiV73i203_2),.clk(gclk));
	jdff dff_B_1XOHmA2o5_2(.din(w_dff_B_LiV73i203_2),.dout(w_dff_B_1XOHmA2o5_2),.clk(gclk));
	jdff dff_B_DNfBUdyz0_2(.din(w_dff_B_1XOHmA2o5_2),.dout(w_dff_B_DNfBUdyz0_2),.clk(gclk));
	jdff dff_B_4i3vdge22_2(.din(w_dff_B_DNfBUdyz0_2),.dout(w_dff_B_4i3vdge22_2),.clk(gclk));
	jdff dff_B_JNGCyc2R0_2(.din(w_dff_B_4i3vdge22_2),.dout(w_dff_B_JNGCyc2R0_2),.clk(gclk));
	jdff dff_B_psIUSbKE4_2(.din(w_dff_B_JNGCyc2R0_2),.dout(w_dff_B_psIUSbKE4_2),.clk(gclk));
	jdff dff_B_LJJNhOXG3_2(.din(w_dff_B_psIUSbKE4_2),.dout(w_dff_B_LJJNhOXG3_2),.clk(gclk));
	jdff dff_B_RPOP7lpy4_2(.din(w_dff_B_LJJNhOXG3_2),.dout(w_dff_B_RPOP7lpy4_2),.clk(gclk));
	jdff dff_B_Dw1Yxqoj4_2(.din(w_dff_B_RPOP7lpy4_2),.dout(w_dff_B_Dw1Yxqoj4_2),.clk(gclk));
	jdff dff_B_BEa72CjN0_2(.din(w_dff_B_Dw1Yxqoj4_2),.dout(w_dff_B_BEa72CjN0_2),.clk(gclk));
	jdff dff_B_VIr7JqWL2_2(.din(w_dff_B_BEa72CjN0_2),.dout(w_dff_B_VIr7JqWL2_2),.clk(gclk));
	jdff dff_B_6L9BxnXQ0_2(.din(w_dff_B_VIr7JqWL2_2),.dout(w_dff_B_6L9BxnXQ0_2),.clk(gclk));
	jdff dff_B_VJd2gfhQ2_2(.din(w_dff_B_6L9BxnXQ0_2),.dout(w_dff_B_VJd2gfhQ2_2),.clk(gclk));
	jdff dff_B_e6b5PeZB6_2(.din(w_dff_B_VJd2gfhQ2_2),.dout(w_dff_B_e6b5PeZB6_2),.clk(gclk));
	jdff dff_B_Mi3PdvAa4_2(.din(w_dff_B_e6b5PeZB6_2),.dout(w_dff_B_Mi3PdvAa4_2),.clk(gclk));
	jdff dff_B_VLVyVtTV6_2(.din(w_dff_B_Mi3PdvAa4_2),.dout(w_dff_B_VLVyVtTV6_2),.clk(gclk));
	jdff dff_B_s82yRrnj0_2(.din(w_dff_B_VLVyVtTV6_2),.dout(w_dff_B_s82yRrnj0_2),.clk(gclk));
	jdff dff_B_4Q9KcXTf9_2(.din(w_dff_B_s82yRrnj0_2),.dout(w_dff_B_4Q9KcXTf9_2),.clk(gclk));
	jdff dff_B_H8LlxpHs5_2(.din(w_dff_B_4Q9KcXTf9_2),.dout(w_dff_B_H8LlxpHs5_2),.clk(gclk));
	jdff dff_B_XRr1dIOp7_1(.din(n1049),.dout(w_dff_B_XRr1dIOp7_1),.clk(gclk));
	jdff dff_B_3o5rqsgq2_2(.din(n949),.dout(w_dff_B_3o5rqsgq2_2),.clk(gclk));
	jdff dff_B_4YMOUERR2_2(.din(w_dff_B_3o5rqsgq2_2),.dout(w_dff_B_4YMOUERR2_2),.clk(gclk));
	jdff dff_B_U5JA5O9V8_2(.din(w_dff_B_4YMOUERR2_2),.dout(w_dff_B_U5JA5O9V8_2),.clk(gclk));
	jdff dff_B_Rzrb5ZfJ1_2(.din(w_dff_B_U5JA5O9V8_2),.dout(w_dff_B_Rzrb5ZfJ1_2),.clk(gclk));
	jdff dff_B_Ny8n0kyf1_2(.din(w_dff_B_Rzrb5ZfJ1_2),.dout(w_dff_B_Ny8n0kyf1_2),.clk(gclk));
	jdff dff_B_zF8eUwa44_2(.din(w_dff_B_Ny8n0kyf1_2),.dout(w_dff_B_zF8eUwa44_2),.clk(gclk));
	jdff dff_B_MoXylkxK3_2(.din(w_dff_B_zF8eUwa44_2),.dout(w_dff_B_MoXylkxK3_2),.clk(gclk));
	jdff dff_B_wSanp7K27_2(.din(w_dff_B_MoXylkxK3_2),.dout(w_dff_B_wSanp7K27_2),.clk(gclk));
	jdff dff_B_0C9iyqU23_2(.din(w_dff_B_wSanp7K27_2),.dout(w_dff_B_0C9iyqU23_2),.clk(gclk));
	jdff dff_B_08PxsBWl0_2(.din(w_dff_B_0C9iyqU23_2),.dout(w_dff_B_08PxsBWl0_2),.clk(gclk));
	jdff dff_B_QD6AugsZ3_2(.din(w_dff_B_08PxsBWl0_2),.dout(w_dff_B_QD6AugsZ3_2),.clk(gclk));
	jdff dff_B_a3LTYmG01_2(.din(w_dff_B_QD6AugsZ3_2),.dout(w_dff_B_a3LTYmG01_2),.clk(gclk));
	jdff dff_B_aHkiFuol9_2(.din(w_dff_B_a3LTYmG01_2),.dout(w_dff_B_aHkiFuol9_2),.clk(gclk));
	jdff dff_B_vVJLfvtI6_2(.din(w_dff_B_aHkiFuol9_2),.dout(w_dff_B_vVJLfvtI6_2),.clk(gclk));
	jdff dff_B_TJjKZfoF1_2(.din(w_dff_B_vVJLfvtI6_2),.dout(w_dff_B_TJjKZfoF1_2),.clk(gclk));
	jdff dff_B_wl9s6AQB5_2(.din(w_dff_B_TJjKZfoF1_2),.dout(w_dff_B_wl9s6AQB5_2),.clk(gclk));
	jdff dff_B_ORs8uBqX0_2(.din(w_dff_B_wl9s6AQB5_2),.dout(w_dff_B_ORs8uBqX0_2),.clk(gclk));
	jdff dff_B_HZ2Qo92N7_2(.din(w_dff_B_ORs8uBqX0_2),.dout(w_dff_B_HZ2Qo92N7_2),.clk(gclk));
	jdff dff_B_qeTXLU0b4_1(.din(n950),.dout(w_dff_B_qeTXLU0b4_1),.clk(gclk));
	jdff dff_B_MV4g2QNt1_2(.din(n847),.dout(w_dff_B_MV4g2QNt1_2),.clk(gclk));
	jdff dff_B_0eHZLoD04_2(.din(w_dff_B_MV4g2QNt1_2),.dout(w_dff_B_0eHZLoD04_2),.clk(gclk));
	jdff dff_B_W7AdgweC5_2(.din(w_dff_B_0eHZLoD04_2),.dout(w_dff_B_W7AdgweC5_2),.clk(gclk));
	jdff dff_B_LS6ZICUD4_2(.din(w_dff_B_W7AdgweC5_2),.dout(w_dff_B_LS6ZICUD4_2),.clk(gclk));
	jdff dff_B_PkFdBYLG5_2(.din(w_dff_B_LS6ZICUD4_2),.dout(w_dff_B_PkFdBYLG5_2),.clk(gclk));
	jdff dff_B_Fb2tyx6g7_2(.din(w_dff_B_PkFdBYLG5_2),.dout(w_dff_B_Fb2tyx6g7_2),.clk(gclk));
	jdff dff_B_rJT8Zncn9_2(.din(w_dff_B_Fb2tyx6g7_2),.dout(w_dff_B_rJT8Zncn9_2),.clk(gclk));
	jdff dff_B_j2p7VuyT1_2(.din(w_dff_B_rJT8Zncn9_2),.dout(w_dff_B_j2p7VuyT1_2),.clk(gclk));
	jdff dff_B_DC6MZPiF0_2(.din(w_dff_B_j2p7VuyT1_2),.dout(w_dff_B_DC6MZPiF0_2),.clk(gclk));
	jdff dff_B_gDN95RFl9_2(.din(w_dff_B_DC6MZPiF0_2),.dout(w_dff_B_gDN95RFl9_2),.clk(gclk));
	jdff dff_B_M7hA9fv73_2(.din(w_dff_B_gDN95RFl9_2),.dout(w_dff_B_M7hA9fv73_2),.clk(gclk));
	jdff dff_B_DbPxRwwp4_2(.din(w_dff_B_M7hA9fv73_2),.dout(w_dff_B_DbPxRwwp4_2),.clk(gclk));
	jdff dff_B_aAxi0Nzn0_2(.din(w_dff_B_DbPxRwwp4_2),.dout(w_dff_B_aAxi0Nzn0_2),.clk(gclk));
	jdff dff_B_hBOGrQ0T1_2(.din(w_dff_B_aAxi0Nzn0_2),.dout(w_dff_B_hBOGrQ0T1_2),.clk(gclk));
	jdff dff_B_NHJGJXl27_2(.din(w_dff_B_hBOGrQ0T1_2),.dout(w_dff_B_NHJGJXl27_2),.clk(gclk));
	jdff dff_B_G3u1fkFI6_2(.din(w_dff_B_NHJGJXl27_2),.dout(w_dff_B_G3u1fkFI6_2),.clk(gclk));
	jdff dff_B_pv43riop8_1(.din(n848),.dout(w_dff_B_pv43riop8_1),.clk(gclk));
	jdff dff_B_wzwUUzUm6_2(.din(n749),.dout(w_dff_B_wzwUUzUm6_2),.clk(gclk));
	jdff dff_B_sGWruZf97_2(.din(w_dff_B_wzwUUzUm6_2),.dout(w_dff_B_sGWruZf97_2),.clk(gclk));
	jdff dff_B_H4z0HhCZ5_2(.din(w_dff_B_sGWruZf97_2),.dout(w_dff_B_H4z0HhCZ5_2),.clk(gclk));
	jdff dff_B_ZJToBRjJ9_2(.din(w_dff_B_H4z0HhCZ5_2),.dout(w_dff_B_ZJToBRjJ9_2),.clk(gclk));
	jdff dff_B_VOnpvlJC5_2(.din(w_dff_B_ZJToBRjJ9_2),.dout(w_dff_B_VOnpvlJC5_2),.clk(gclk));
	jdff dff_B_Z27iRV4o5_2(.din(w_dff_B_VOnpvlJC5_2),.dout(w_dff_B_Z27iRV4o5_2),.clk(gclk));
	jdff dff_B_ILFoDVZr5_2(.din(w_dff_B_Z27iRV4o5_2),.dout(w_dff_B_ILFoDVZr5_2),.clk(gclk));
	jdff dff_B_RHfHr3450_2(.din(w_dff_B_ILFoDVZr5_2),.dout(w_dff_B_RHfHr3450_2),.clk(gclk));
	jdff dff_B_ONCMmMQe1_2(.din(w_dff_B_RHfHr3450_2),.dout(w_dff_B_ONCMmMQe1_2),.clk(gclk));
	jdff dff_B_SM3xvBQ74_2(.din(w_dff_B_ONCMmMQe1_2),.dout(w_dff_B_SM3xvBQ74_2),.clk(gclk));
	jdff dff_B_sGBLMMv97_2(.din(w_dff_B_SM3xvBQ74_2),.dout(w_dff_B_sGBLMMv97_2),.clk(gclk));
	jdff dff_B_85GcJfkc8_2(.din(w_dff_B_sGBLMMv97_2),.dout(w_dff_B_85GcJfkc8_2),.clk(gclk));
	jdff dff_B_EQkdYyZx9_2(.din(w_dff_B_85GcJfkc8_2),.dout(w_dff_B_EQkdYyZx9_2),.clk(gclk));
	jdff dff_B_8lzSH3qA1_2(.din(w_dff_B_EQkdYyZx9_2),.dout(w_dff_B_8lzSH3qA1_2),.clk(gclk));
	jdff dff_B_yHDS6tVh6_1(.din(n750),.dout(w_dff_B_yHDS6tVh6_1),.clk(gclk));
	jdff dff_B_46lKdd870_2(.din(n657),.dout(w_dff_B_46lKdd870_2),.clk(gclk));
	jdff dff_B_lbO1yTzX7_2(.din(w_dff_B_46lKdd870_2),.dout(w_dff_B_lbO1yTzX7_2),.clk(gclk));
	jdff dff_B_E2FFnZge7_2(.din(w_dff_B_lbO1yTzX7_2),.dout(w_dff_B_E2FFnZge7_2),.clk(gclk));
	jdff dff_B_FVVSrVpF4_2(.din(w_dff_B_E2FFnZge7_2),.dout(w_dff_B_FVVSrVpF4_2),.clk(gclk));
	jdff dff_B_ni1JN2Xc0_2(.din(w_dff_B_FVVSrVpF4_2),.dout(w_dff_B_ni1JN2Xc0_2),.clk(gclk));
	jdff dff_B_secEvfco7_2(.din(w_dff_B_ni1JN2Xc0_2),.dout(w_dff_B_secEvfco7_2),.clk(gclk));
	jdff dff_B_QSOhLVTd7_2(.din(w_dff_B_secEvfco7_2),.dout(w_dff_B_QSOhLVTd7_2),.clk(gclk));
	jdff dff_B_dD4Wqlsh4_2(.din(w_dff_B_QSOhLVTd7_2),.dout(w_dff_B_dD4Wqlsh4_2),.clk(gclk));
	jdff dff_B_PraNFw2U9_2(.din(w_dff_B_dD4Wqlsh4_2),.dout(w_dff_B_PraNFw2U9_2),.clk(gclk));
	jdff dff_B_Rb50kEvB0_2(.din(w_dff_B_PraNFw2U9_2),.dout(w_dff_B_Rb50kEvB0_2),.clk(gclk));
	jdff dff_B_JXa4nZxj1_2(.din(w_dff_B_Rb50kEvB0_2),.dout(w_dff_B_JXa4nZxj1_2),.clk(gclk));
	jdff dff_B_nJrMpPDH9_2(.din(w_dff_B_JXa4nZxj1_2),.dout(w_dff_B_nJrMpPDH9_2),.clk(gclk));
	jdff dff_B_pqEVTRr14_1(.din(n658),.dout(w_dff_B_pqEVTRr14_1),.clk(gclk));
	jdff dff_B_vZ7Tk3AX0_2(.din(n572),.dout(w_dff_B_vZ7Tk3AX0_2),.clk(gclk));
	jdff dff_B_FvkMsqtZ1_2(.din(w_dff_B_vZ7Tk3AX0_2),.dout(w_dff_B_FvkMsqtZ1_2),.clk(gclk));
	jdff dff_B_a74mIRXI9_2(.din(w_dff_B_FvkMsqtZ1_2),.dout(w_dff_B_a74mIRXI9_2),.clk(gclk));
	jdff dff_B_xAWvAewH2_2(.din(w_dff_B_a74mIRXI9_2),.dout(w_dff_B_xAWvAewH2_2),.clk(gclk));
	jdff dff_B_ZjSdn17E9_2(.din(w_dff_B_xAWvAewH2_2),.dout(w_dff_B_ZjSdn17E9_2),.clk(gclk));
	jdff dff_B_aLhjPEKB1_2(.din(w_dff_B_ZjSdn17E9_2),.dout(w_dff_B_aLhjPEKB1_2),.clk(gclk));
	jdff dff_B_DdgUgEna3_2(.din(w_dff_B_aLhjPEKB1_2),.dout(w_dff_B_DdgUgEna3_2),.clk(gclk));
	jdff dff_B_tEaF8pVO8_2(.din(w_dff_B_DdgUgEna3_2),.dout(w_dff_B_tEaF8pVO8_2),.clk(gclk));
	jdff dff_B_NBUfx7Fj6_2(.din(w_dff_B_tEaF8pVO8_2),.dout(w_dff_B_NBUfx7Fj6_2),.clk(gclk));
	jdff dff_B_v8dDabgb2_2(.din(w_dff_B_NBUfx7Fj6_2),.dout(w_dff_B_v8dDabgb2_2),.clk(gclk));
	jdff dff_B_hJD0JWYq0_1(.din(n573),.dout(w_dff_B_hJD0JWYq0_1),.clk(gclk));
	jdff dff_B_VFwt9rHg2_2(.din(n494),.dout(w_dff_B_VFwt9rHg2_2),.clk(gclk));
	jdff dff_B_T9pbeyQO9_2(.din(w_dff_B_VFwt9rHg2_2),.dout(w_dff_B_T9pbeyQO9_2),.clk(gclk));
	jdff dff_B_6OL5UTYf6_2(.din(w_dff_B_T9pbeyQO9_2),.dout(w_dff_B_6OL5UTYf6_2),.clk(gclk));
	jdff dff_B_TPERxyw56_2(.din(w_dff_B_6OL5UTYf6_2),.dout(w_dff_B_TPERxyw56_2),.clk(gclk));
	jdff dff_B_A8gqdoZC5_2(.din(w_dff_B_TPERxyw56_2),.dout(w_dff_B_A8gqdoZC5_2),.clk(gclk));
	jdff dff_B_x5HBSNPC4_2(.din(w_dff_B_A8gqdoZC5_2),.dout(w_dff_B_x5HBSNPC4_2),.clk(gclk));
	jdff dff_B_Q4cWheUz4_2(.din(w_dff_B_x5HBSNPC4_2),.dout(w_dff_B_Q4cWheUz4_2),.clk(gclk));
	jdff dff_B_R9xRJ5ll5_2(.din(w_dff_B_Q4cWheUz4_2),.dout(w_dff_B_R9xRJ5ll5_2),.clk(gclk));
	jdff dff_B_tMloJh7K6_2(.din(n509),.dout(w_dff_B_tMloJh7K6_2),.clk(gclk));
	jdff dff_B_CFjS2mkS2_2(.din(w_dff_B_tMloJh7K6_2),.dout(w_dff_B_CFjS2mkS2_2),.clk(gclk));
	jdff dff_B_UcTBY1zo6_2(.din(w_dff_B_CFjS2mkS2_2),.dout(w_dff_B_UcTBY1zo6_2),.clk(gclk));
	jdff dff_B_0Nzhwj1O0_1(.din(n495),.dout(w_dff_B_0Nzhwj1O0_1),.clk(gclk));
	jdff dff_B_H81iEytJ1_1(.din(w_dff_B_0Nzhwj1O0_1),.dout(w_dff_B_H81iEytJ1_1),.clk(gclk));
	jdff dff_B_nZmWx5Sh4_1(.din(w_dff_B_H81iEytJ1_1),.dout(w_dff_B_nZmWx5Sh4_1),.clk(gclk));
	jdff dff_B_qE3ues0G9_2(.din(n425),.dout(w_dff_B_qE3ues0G9_2),.clk(gclk));
	jdff dff_B_66EUHV0c6_2(.din(w_dff_B_qE3ues0G9_2),.dout(w_dff_B_66EUHV0c6_2),.clk(gclk));
	jdff dff_B_tL739E4x0_2(.din(w_dff_B_66EUHV0c6_2),.dout(w_dff_B_tL739E4x0_2),.clk(gclk));
	jdff dff_B_UeAzmlqM4_0(.din(n430),.dout(w_dff_B_UeAzmlqM4_0),.clk(gclk));
	jdff dff_B_xsOacfNt7_0(.din(w_dff_B_UeAzmlqM4_0),.dout(w_dff_B_xsOacfNt7_0),.clk(gclk));
	jdff dff_A_8d0lntMq6_0(.dout(w_n358_0[0]),.din(w_dff_A_8d0lntMq6_0),.clk(gclk));
	jdff dff_A_BwRsfu1h5_0(.dout(w_dff_A_8d0lntMq6_0),.din(w_dff_A_BwRsfu1h5_0),.clk(gclk));
	jdff dff_A_Dof8RIBx2_1(.dout(w_n358_0[1]),.din(w_dff_A_Dof8RIBx2_1),.clk(gclk));
	jdff dff_A_JeJnM9zr2_1(.dout(w_dff_A_Dof8RIBx2_1),.din(w_dff_A_JeJnM9zr2_1),.clk(gclk));
	jdff dff_B_xnQZKn1e6_2(.din(n1651),.dout(w_dff_B_xnQZKn1e6_2),.clk(gclk));
	jdff dff_B_mkSi4f4V7_1(.din(n1649),.dout(w_dff_B_mkSi4f4V7_1),.clk(gclk));
	jdff dff_B_VBW0ogTI6_2(.din(n1597),.dout(w_dff_B_VBW0ogTI6_2),.clk(gclk));
	jdff dff_B_v1rfo64M4_2(.din(w_dff_B_VBW0ogTI6_2),.dout(w_dff_B_v1rfo64M4_2),.clk(gclk));
	jdff dff_B_5uEtOVsX1_2(.din(w_dff_B_v1rfo64M4_2),.dout(w_dff_B_5uEtOVsX1_2),.clk(gclk));
	jdff dff_B_vA7Gn5HE4_2(.din(w_dff_B_5uEtOVsX1_2),.dout(w_dff_B_vA7Gn5HE4_2),.clk(gclk));
	jdff dff_B_cKb7ezjL7_2(.din(w_dff_B_vA7Gn5HE4_2),.dout(w_dff_B_cKb7ezjL7_2),.clk(gclk));
	jdff dff_B_FyPHq40p4_2(.din(w_dff_B_cKb7ezjL7_2),.dout(w_dff_B_FyPHq40p4_2),.clk(gclk));
	jdff dff_B_S3wNH8I13_2(.din(w_dff_B_FyPHq40p4_2),.dout(w_dff_B_S3wNH8I13_2),.clk(gclk));
	jdff dff_B_bYp6fC688_2(.din(w_dff_B_S3wNH8I13_2),.dout(w_dff_B_bYp6fC688_2),.clk(gclk));
	jdff dff_B_XjrGQonB5_2(.din(w_dff_B_bYp6fC688_2),.dout(w_dff_B_XjrGQonB5_2),.clk(gclk));
	jdff dff_B_PUetbgfh8_2(.din(w_dff_B_XjrGQonB5_2),.dout(w_dff_B_PUetbgfh8_2),.clk(gclk));
	jdff dff_B_IR4AG0en0_2(.din(w_dff_B_PUetbgfh8_2),.dout(w_dff_B_IR4AG0en0_2),.clk(gclk));
	jdff dff_B_iYvU3GlE3_2(.din(w_dff_B_IR4AG0en0_2),.dout(w_dff_B_iYvU3GlE3_2),.clk(gclk));
	jdff dff_B_I1MDHbGc8_2(.din(w_dff_B_iYvU3GlE3_2),.dout(w_dff_B_I1MDHbGc8_2),.clk(gclk));
	jdff dff_B_l3Uq8J3R3_2(.din(w_dff_B_I1MDHbGc8_2),.dout(w_dff_B_l3Uq8J3R3_2),.clk(gclk));
	jdff dff_B_fuC5iLKZ6_2(.din(w_dff_B_l3Uq8J3R3_2),.dout(w_dff_B_fuC5iLKZ6_2),.clk(gclk));
	jdff dff_B_dSrZ6e8f8_2(.din(w_dff_B_fuC5iLKZ6_2),.dout(w_dff_B_dSrZ6e8f8_2),.clk(gclk));
	jdff dff_B_giSfxoBs5_2(.din(w_dff_B_dSrZ6e8f8_2),.dout(w_dff_B_giSfxoBs5_2),.clk(gclk));
	jdff dff_B_YcJC36jV9_2(.din(w_dff_B_giSfxoBs5_2),.dout(w_dff_B_YcJC36jV9_2),.clk(gclk));
	jdff dff_B_UkU0bqgI9_2(.din(w_dff_B_YcJC36jV9_2),.dout(w_dff_B_UkU0bqgI9_2),.clk(gclk));
	jdff dff_B_pbWx9hp86_2(.din(w_dff_B_UkU0bqgI9_2),.dout(w_dff_B_pbWx9hp86_2),.clk(gclk));
	jdff dff_B_f535UBey5_2(.din(w_dff_B_pbWx9hp86_2),.dout(w_dff_B_f535UBey5_2),.clk(gclk));
	jdff dff_B_drC7sw329_2(.din(w_dff_B_f535UBey5_2),.dout(w_dff_B_drC7sw329_2),.clk(gclk));
	jdff dff_B_biQrQ1sy3_2(.din(w_dff_B_drC7sw329_2),.dout(w_dff_B_biQrQ1sy3_2),.clk(gclk));
	jdff dff_B_PvuNGnTA0_2(.din(w_dff_B_biQrQ1sy3_2),.dout(w_dff_B_PvuNGnTA0_2),.clk(gclk));
	jdff dff_B_qEhnOnfS6_2(.din(w_dff_B_PvuNGnTA0_2),.dout(w_dff_B_qEhnOnfS6_2),.clk(gclk));
	jdff dff_B_UVALDTH68_2(.din(w_dff_B_qEhnOnfS6_2),.dout(w_dff_B_UVALDTH68_2),.clk(gclk));
	jdff dff_B_wb9MDVlw4_2(.din(w_dff_B_UVALDTH68_2),.dout(w_dff_B_wb9MDVlw4_2),.clk(gclk));
	jdff dff_B_kxeHh8gX1_2(.din(w_dff_B_wb9MDVlw4_2),.dout(w_dff_B_kxeHh8gX1_2),.clk(gclk));
	jdff dff_B_yQSN8lAV2_2(.din(w_dff_B_kxeHh8gX1_2),.dout(w_dff_B_yQSN8lAV2_2),.clk(gclk));
	jdff dff_B_59J1qeTa2_2(.din(w_dff_B_yQSN8lAV2_2),.dout(w_dff_B_59J1qeTa2_2),.clk(gclk));
	jdff dff_B_Ni8wF5Du1_2(.din(w_dff_B_59J1qeTa2_2),.dout(w_dff_B_Ni8wF5Du1_2),.clk(gclk));
	jdff dff_B_V2TkmjJu0_2(.din(w_dff_B_Ni8wF5Du1_2),.dout(w_dff_B_V2TkmjJu0_2),.clk(gclk));
	jdff dff_B_5cGNZfKr3_2(.din(w_dff_B_V2TkmjJu0_2),.dout(w_dff_B_5cGNZfKr3_2),.clk(gclk));
	jdff dff_B_ISv9F1e59_2(.din(w_dff_B_5cGNZfKr3_2),.dout(w_dff_B_ISv9F1e59_2),.clk(gclk));
	jdff dff_B_RbBpgmtv8_2(.din(w_dff_B_ISv9F1e59_2),.dout(w_dff_B_RbBpgmtv8_2),.clk(gclk));
	jdff dff_B_2jGGkJn77_2(.din(w_dff_B_RbBpgmtv8_2),.dout(w_dff_B_2jGGkJn77_2),.clk(gclk));
	jdff dff_B_wqI2kAQe6_2(.din(w_dff_B_2jGGkJn77_2),.dout(w_dff_B_wqI2kAQe6_2),.clk(gclk));
	jdff dff_B_TtcXziLy1_2(.din(w_dff_B_wqI2kAQe6_2),.dout(w_dff_B_TtcXziLy1_2),.clk(gclk));
	jdff dff_B_e2z1JxOl1_1(.din(n1647),.dout(w_dff_B_e2z1JxOl1_1),.clk(gclk));
	jdff dff_A_6pYNKldV8_1(.dout(w_n1600_0[1]),.din(w_dff_A_6pYNKldV8_1),.clk(gclk));
	jdff dff_B_TSNOL1hx3_1(.din(n1598),.dout(w_dff_B_TSNOL1hx3_1),.clk(gclk));
	jdff dff_B_mrDJFLs04_2(.din(n1540),.dout(w_dff_B_mrDJFLs04_2),.clk(gclk));
	jdff dff_B_W8cHUeGZ6_2(.din(w_dff_B_mrDJFLs04_2),.dout(w_dff_B_W8cHUeGZ6_2),.clk(gclk));
	jdff dff_B_1PnuUv3N0_2(.din(w_dff_B_W8cHUeGZ6_2),.dout(w_dff_B_1PnuUv3N0_2),.clk(gclk));
	jdff dff_B_C9r2fK6t9_2(.din(w_dff_B_1PnuUv3N0_2),.dout(w_dff_B_C9r2fK6t9_2),.clk(gclk));
	jdff dff_B_zk2KIBey5_2(.din(w_dff_B_C9r2fK6t9_2),.dout(w_dff_B_zk2KIBey5_2),.clk(gclk));
	jdff dff_B_I1Wo4Yuv6_2(.din(w_dff_B_zk2KIBey5_2),.dout(w_dff_B_I1Wo4Yuv6_2),.clk(gclk));
	jdff dff_B_HPViOFY71_2(.din(w_dff_B_I1Wo4Yuv6_2),.dout(w_dff_B_HPViOFY71_2),.clk(gclk));
	jdff dff_B_Cv0Y47s56_2(.din(w_dff_B_HPViOFY71_2),.dout(w_dff_B_Cv0Y47s56_2),.clk(gclk));
	jdff dff_B_9RQSnSrE4_2(.din(w_dff_B_Cv0Y47s56_2),.dout(w_dff_B_9RQSnSrE4_2),.clk(gclk));
	jdff dff_B_QDUvAwlg1_2(.din(w_dff_B_9RQSnSrE4_2),.dout(w_dff_B_QDUvAwlg1_2),.clk(gclk));
	jdff dff_B_uy26qrPp3_2(.din(w_dff_B_QDUvAwlg1_2),.dout(w_dff_B_uy26qrPp3_2),.clk(gclk));
	jdff dff_B_2FAmawaL9_2(.din(w_dff_B_uy26qrPp3_2),.dout(w_dff_B_2FAmawaL9_2),.clk(gclk));
	jdff dff_B_bblRoeif6_2(.din(w_dff_B_2FAmawaL9_2),.dout(w_dff_B_bblRoeif6_2),.clk(gclk));
	jdff dff_B_NmDeHrv92_2(.din(w_dff_B_bblRoeif6_2),.dout(w_dff_B_NmDeHrv92_2),.clk(gclk));
	jdff dff_B_iag5fKQv0_2(.din(w_dff_B_NmDeHrv92_2),.dout(w_dff_B_iag5fKQv0_2),.clk(gclk));
	jdff dff_B_UqmFmJSE5_2(.din(w_dff_B_iag5fKQv0_2),.dout(w_dff_B_UqmFmJSE5_2),.clk(gclk));
	jdff dff_B_NUfuTtUN9_2(.din(w_dff_B_UqmFmJSE5_2),.dout(w_dff_B_NUfuTtUN9_2),.clk(gclk));
	jdff dff_B_KPj8zJaL3_2(.din(w_dff_B_NUfuTtUN9_2),.dout(w_dff_B_KPj8zJaL3_2),.clk(gclk));
	jdff dff_B_54Lssekp8_2(.din(w_dff_B_KPj8zJaL3_2),.dout(w_dff_B_54Lssekp8_2),.clk(gclk));
	jdff dff_B_MPCYk8OS1_2(.din(w_dff_B_54Lssekp8_2),.dout(w_dff_B_MPCYk8OS1_2),.clk(gclk));
	jdff dff_B_v9Qg1kqt6_2(.din(w_dff_B_MPCYk8OS1_2),.dout(w_dff_B_v9Qg1kqt6_2),.clk(gclk));
	jdff dff_B_KPqy328H8_2(.din(w_dff_B_v9Qg1kqt6_2),.dout(w_dff_B_KPqy328H8_2),.clk(gclk));
	jdff dff_B_h5sjxDfW7_2(.din(w_dff_B_KPqy328H8_2),.dout(w_dff_B_h5sjxDfW7_2),.clk(gclk));
	jdff dff_B_3B3PTyVI2_2(.din(w_dff_B_h5sjxDfW7_2),.dout(w_dff_B_3B3PTyVI2_2),.clk(gclk));
	jdff dff_B_1W9eD1rp9_2(.din(w_dff_B_3B3PTyVI2_2),.dout(w_dff_B_1W9eD1rp9_2),.clk(gclk));
	jdff dff_B_G9apCEHq0_2(.din(w_dff_B_1W9eD1rp9_2),.dout(w_dff_B_G9apCEHq0_2),.clk(gclk));
	jdff dff_B_DebhzyCI5_2(.din(w_dff_B_G9apCEHq0_2),.dout(w_dff_B_DebhzyCI5_2),.clk(gclk));
	jdff dff_B_EeJqWmaU2_2(.din(w_dff_B_DebhzyCI5_2),.dout(w_dff_B_EeJqWmaU2_2),.clk(gclk));
	jdff dff_B_mXaempWy3_2(.din(w_dff_B_EeJqWmaU2_2),.dout(w_dff_B_mXaempWy3_2),.clk(gclk));
	jdff dff_B_YOdfcH9A2_2(.din(w_dff_B_mXaempWy3_2),.dout(w_dff_B_YOdfcH9A2_2),.clk(gclk));
	jdff dff_B_KmXp3FyI1_2(.din(w_dff_B_YOdfcH9A2_2),.dout(w_dff_B_KmXp3FyI1_2),.clk(gclk));
	jdff dff_B_fkTswcPr6_2(.din(w_dff_B_KmXp3FyI1_2),.dout(w_dff_B_fkTswcPr6_2),.clk(gclk));
	jdff dff_B_x51BuWjL3_2(.din(w_dff_B_fkTswcPr6_2),.dout(w_dff_B_x51BuWjL3_2),.clk(gclk));
	jdff dff_B_O0h7KmFr2_2(.din(n1543),.dout(w_dff_B_O0h7KmFr2_2),.clk(gclk));
	jdff dff_B_u31k2Nk20_1(.din(n1541),.dout(w_dff_B_u31k2Nk20_1),.clk(gclk));
	jdff dff_B_H2OXBbe60_2(.din(n1476),.dout(w_dff_B_H2OXBbe60_2),.clk(gclk));
	jdff dff_B_bGnWXqi60_2(.din(w_dff_B_H2OXBbe60_2),.dout(w_dff_B_bGnWXqi60_2),.clk(gclk));
	jdff dff_B_P8ofvFfx7_2(.din(w_dff_B_bGnWXqi60_2),.dout(w_dff_B_P8ofvFfx7_2),.clk(gclk));
	jdff dff_B_e1svo0Zp3_2(.din(w_dff_B_P8ofvFfx7_2),.dout(w_dff_B_e1svo0Zp3_2),.clk(gclk));
	jdff dff_B_jcTSoOaC6_2(.din(w_dff_B_e1svo0Zp3_2),.dout(w_dff_B_jcTSoOaC6_2),.clk(gclk));
	jdff dff_B_VCwa01U53_2(.din(w_dff_B_jcTSoOaC6_2),.dout(w_dff_B_VCwa01U53_2),.clk(gclk));
	jdff dff_B_3cFxOmPa2_2(.din(w_dff_B_VCwa01U53_2),.dout(w_dff_B_3cFxOmPa2_2),.clk(gclk));
	jdff dff_B_QKCVJ6FN0_2(.din(w_dff_B_3cFxOmPa2_2),.dout(w_dff_B_QKCVJ6FN0_2),.clk(gclk));
	jdff dff_B_pmQdjvRI5_2(.din(w_dff_B_QKCVJ6FN0_2),.dout(w_dff_B_pmQdjvRI5_2),.clk(gclk));
	jdff dff_B_zf69GMFj3_2(.din(w_dff_B_pmQdjvRI5_2),.dout(w_dff_B_zf69GMFj3_2),.clk(gclk));
	jdff dff_B_KsRGGLFJ3_2(.din(w_dff_B_zf69GMFj3_2),.dout(w_dff_B_KsRGGLFJ3_2),.clk(gclk));
	jdff dff_B_moAuZaV85_2(.din(w_dff_B_KsRGGLFJ3_2),.dout(w_dff_B_moAuZaV85_2),.clk(gclk));
	jdff dff_B_wFmrwfXv7_2(.din(w_dff_B_moAuZaV85_2),.dout(w_dff_B_wFmrwfXv7_2),.clk(gclk));
	jdff dff_B_TEwjkeF74_2(.din(w_dff_B_wFmrwfXv7_2),.dout(w_dff_B_TEwjkeF74_2),.clk(gclk));
	jdff dff_B_7WNqZ5P39_2(.din(w_dff_B_TEwjkeF74_2),.dout(w_dff_B_7WNqZ5P39_2),.clk(gclk));
	jdff dff_B_YP0FbpPG0_2(.din(w_dff_B_7WNqZ5P39_2),.dout(w_dff_B_YP0FbpPG0_2),.clk(gclk));
	jdff dff_B_YY09gFww6_2(.din(w_dff_B_YP0FbpPG0_2),.dout(w_dff_B_YY09gFww6_2),.clk(gclk));
	jdff dff_B_lwF4kr7x7_2(.din(w_dff_B_YY09gFww6_2),.dout(w_dff_B_lwF4kr7x7_2),.clk(gclk));
	jdff dff_B_jBAMjf907_2(.din(w_dff_B_lwF4kr7x7_2),.dout(w_dff_B_jBAMjf907_2),.clk(gclk));
	jdff dff_B_yq7oWzje7_2(.din(w_dff_B_jBAMjf907_2),.dout(w_dff_B_yq7oWzje7_2),.clk(gclk));
	jdff dff_B_mRCykEN71_2(.din(w_dff_B_yq7oWzje7_2),.dout(w_dff_B_mRCykEN71_2),.clk(gclk));
	jdff dff_B_0WDdaiKY2_2(.din(w_dff_B_mRCykEN71_2),.dout(w_dff_B_0WDdaiKY2_2),.clk(gclk));
	jdff dff_B_QT5TQdAh1_2(.din(w_dff_B_0WDdaiKY2_2),.dout(w_dff_B_QT5TQdAh1_2),.clk(gclk));
	jdff dff_B_3TdHUadp2_2(.din(w_dff_B_QT5TQdAh1_2),.dout(w_dff_B_3TdHUadp2_2),.clk(gclk));
	jdff dff_B_d4Jc6hM94_2(.din(w_dff_B_3TdHUadp2_2),.dout(w_dff_B_d4Jc6hM94_2),.clk(gclk));
	jdff dff_B_mi6L5EPP3_2(.din(w_dff_B_d4Jc6hM94_2),.dout(w_dff_B_mi6L5EPP3_2),.clk(gclk));
	jdff dff_B_Jle96uyH5_2(.din(w_dff_B_mi6L5EPP3_2),.dout(w_dff_B_Jle96uyH5_2),.clk(gclk));
	jdff dff_B_b5EcWls47_2(.din(w_dff_B_Jle96uyH5_2),.dout(w_dff_B_b5EcWls47_2),.clk(gclk));
	jdff dff_B_37bKEhBh2_2(.din(w_dff_B_b5EcWls47_2),.dout(w_dff_B_37bKEhBh2_2),.clk(gclk));
	jdff dff_B_MDqnxK5G5_2(.din(w_dff_B_37bKEhBh2_2),.dout(w_dff_B_MDqnxK5G5_2),.clk(gclk));
	jdff dff_B_zyA9jFjr4_2(.din(n1479),.dout(w_dff_B_zyA9jFjr4_2),.clk(gclk));
	jdff dff_B_2vYE8m0s1_1(.din(n1477),.dout(w_dff_B_2vYE8m0s1_1),.clk(gclk));
	jdff dff_B_Lp7qrQX68_2(.din(n1405),.dout(w_dff_B_Lp7qrQX68_2),.clk(gclk));
	jdff dff_B_GOI2Y9Hg3_2(.din(w_dff_B_Lp7qrQX68_2),.dout(w_dff_B_GOI2Y9Hg3_2),.clk(gclk));
	jdff dff_B_cXlxZi112_2(.din(w_dff_B_GOI2Y9Hg3_2),.dout(w_dff_B_cXlxZi112_2),.clk(gclk));
	jdff dff_B_PLcetyJE8_2(.din(w_dff_B_cXlxZi112_2),.dout(w_dff_B_PLcetyJE8_2),.clk(gclk));
	jdff dff_B_jZYNkq4D0_2(.din(w_dff_B_PLcetyJE8_2),.dout(w_dff_B_jZYNkq4D0_2),.clk(gclk));
	jdff dff_B_tWsxuWkU3_2(.din(w_dff_B_jZYNkq4D0_2),.dout(w_dff_B_tWsxuWkU3_2),.clk(gclk));
	jdff dff_B_LSXcQq172_2(.din(w_dff_B_tWsxuWkU3_2),.dout(w_dff_B_LSXcQq172_2),.clk(gclk));
	jdff dff_B_PEIXlRVK9_2(.din(w_dff_B_LSXcQq172_2),.dout(w_dff_B_PEIXlRVK9_2),.clk(gclk));
	jdff dff_B_6wzu7IFF4_2(.din(w_dff_B_PEIXlRVK9_2),.dout(w_dff_B_6wzu7IFF4_2),.clk(gclk));
	jdff dff_B_ZmVlozeC0_2(.din(w_dff_B_6wzu7IFF4_2),.dout(w_dff_B_ZmVlozeC0_2),.clk(gclk));
	jdff dff_B_abLewnl91_2(.din(w_dff_B_ZmVlozeC0_2),.dout(w_dff_B_abLewnl91_2),.clk(gclk));
	jdff dff_B_8Tzx9gzi2_2(.din(w_dff_B_abLewnl91_2),.dout(w_dff_B_8Tzx9gzi2_2),.clk(gclk));
	jdff dff_B_xEo1Kzkw9_2(.din(w_dff_B_8Tzx9gzi2_2),.dout(w_dff_B_xEo1Kzkw9_2),.clk(gclk));
	jdff dff_B_oyhSLhkL7_2(.din(w_dff_B_xEo1Kzkw9_2),.dout(w_dff_B_oyhSLhkL7_2),.clk(gclk));
	jdff dff_B_V7ksLEFL8_2(.din(w_dff_B_oyhSLhkL7_2),.dout(w_dff_B_V7ksLEFL8_2),.clk(gclk));
	jdff dff_B_uhbOoM2d0_2(.din(w_dff_B_V7ksLEFL8_2),.dout(w_dff_B_uhbOoM2d0_2),.clk(gclk));
	jdff dff_B_UyWvtaUl7_2(.din(w_dff_B_uhbOoM2d0_2),.dout(w_dff_B_UyWvtaUl7_2),.clk(gclk));
	jdff dff_B_kbO544K39_2(.din(w_dff_B_UyWvtaUl7_2),.dout(w_dff_B_kbO544K39_2),.clk(gclk));
	jdff dff_B_1cA5keYn5_2(.din(w_dff_B_kbO544K39_2),.dout(w_dff_B_1cA5keYn5_2),.clk(gclk));
	jdff dff_B_EfpL2XTI4_2(.din(w_dff_B_1cA5keYn5_2),.dout(w_dff_B_EfpL2XTI4_2),.clk(gclk));
	jdff dff_B_sWd6KsID9_2(.din(w_dff_B_EfpL2XTI4_2),.dout(w_dff_B_sWd6KsID9_2),.clk(gclk));
	jdff dff_B_QLWdYeyX0_2(.din(w_dff_B_sWd6KsID9_2),.dout(w_dff_B_QLWdYeyX0_2),.clk(gclk));
	jdff dff_B_ybNKA7OT0_2(.din(w_dff_B_QLWdYeyX0_2),.dout(w_dff_B_ybNKA7OT0_2),.clk(gclk));
	jdff dff_B_h025lGvm0_2(.din(w_dff_B_ybNKA7OT0_2),.dout(w_dff_B_h025lGvm0_2),.clk(gclk));
	jdff dff_B_I81kX4pU9_2(.din(w_dff_B_h025lGvm0_2),.dout(w_dff_B_I81kX4pU9_2),.clk(gclk));
	jdff dff_B_a0zie5520_2(.din(w_dff_B_I81kX4pU9_2),.dout(w_dff_B_a0zie5520_2),.clk(gclk));
	jdff dff_B_epbHyQ9n1_2(.din(w_dff_B_a0zie5520_2),.dout(w_dff_B_epbHyQ9n1_2),.clk(gclk));
	jdff dff_B_LfDwkVxA7_2(.din(n1408),.dout(w_dff_B_LfDwkVxA7_2),.clk(gclk));
	jdff dff_B_iLDdWkPX6_1(.din(n1406),.dout(w_dff_B_iLDdWkPX6_1),.clk(gclk));
	jdff dff_B_LHZ4VKIQ4_2(.din(n1327),.dout(w_dff_B_LHZ4VKIQ4_2),.clk(gclk));
	jdff dff_B_KezderHx2_2(.din(w_dff_B_LHZ4VKIQ4_2),.dout(w_dff_B_KezderHx2_2),.clk(gclk));
	jdff dff_B_zZOMMQSe4_2(.din(w_dff_B_KezderHx2_2),.dout(w_dff_B_zZOMMQSe4_2),.clk(gclk));
	jdff dff_B_8j2kBVfM4_2(.din(w_dff_B_zZOMMQSe4_2),.dout(w_dff_B_8j2kBVfM4_2),.clk(gclk));
	jdff dff_B_dCYtdT4w2_2(.din(w_dff_B_8j2kBVfM4_2),.dout(w_dff_B_dCYtdT4w2_2),.clk(gclk));
	jdff dff_B_EVyvL9BR6_2(.din(w_dff_B_dCYtdT4w2_2),.dout(w_dff_B_EVyvL9BR6_2),.clk(gclk));
	jdff dff_B_B6KoHIF87_2(.din(w_dff_B_EVyvL9BR6_2),.dout(w_dff_B_B6KoHIF87_2),.clk(gclk));
	jdff dff_B_ZMqyKINg0_2(.din(w_dff_B_B6KoHIF87_2),.dout(w_dff_B_ZMqyKINg0_2),.clk(gclk));
	jdff dff_B_CkXqgppJ3_2(.din(w_dff_B_ZMqyKINg0_2),.dout(w_dff_B_CkXqgppJ3_2),.clk(gclk));
	jdff dff_B_CyJj60EX0_2(.din(w_dff_B_CkXqgppJ3_2),.dout(w_dff_B_CyJj60EX0_2),.clk(gclk));
	jdff dff_B_SeFTTevc0_2(.din(w_dff_B_CyJj60EX0_2),.dout(w_dff_B_SeFTTevc0_2),.clk(gclk));
	jdff dff_B_9IZW18Hb4_2(.din(w_dff_B_SeFTTevc0_2),.dout(w_dff_B_9IZW18Hb4_2),.clk(gclk));
	jdff dff_B_7vaySFdw6_2(.din(w_dff_B_9IZW18Hb4_2),.dout(w_dff_B_7vaySFdw6_2),.clk(gclk));
	jdff dff_B_jYSe9qsF4_2(.din(w_dff_B_7vaySFdw6_2),.dout(w_dff_B_jYSe9qsF4_2),.clk(gclk));
	jdff dff_B_gyu3aPvi6_2(.din(w_dff_B_jYSe9qsF4_2),.dout(w_dff_B_gyu3aPvi6_2),.clk(gclk));
	jdff dff_B_GOicqNIt5_2(.din(w_dff_B_gyu3aPvi6_2),.dout(w_dff_B_GOicqNIt5_2),.clk(gclk));
	jdff dff_B_awE6hmV85_2(.din(w_dff_B_GOicqNIt5_2),.dout(w_dff_B_awE6hmV85_2),.clk(gclk));
	jdff dff_B_jslbRFA42_2(.din(w_dff_B_awE6hmV85_2),.dout(w_dff_B_jslbRFA42_2),.clk(gclk));
	jdff dff_B_Q4O5XPDp2_2(.din(w_dff_B_jslbRFA42_2),.dout(w_dff_B_Q4O5XPDp2_2),.clk(gclk));
	jdff dff_B_ZAZKT3xQ9_2(.din(w_dff_B_Q4O5XPDp2_2),.dout(w_dff_B_ZAZKT3xQ9_2),.clk(gclk));
	jdff dff_B_gxTUHhmZ6_2(.din(w_dff_B_ZAZKT3xQ9_2),.dout(w_dff_B_gxTUHhmZ6_2),.clk(gclk));
	jdff dff_B_pCx6GYyo0_2(.din(w_dff_B_gxTUHhmZ6_2),.dout(w_dff_B_pCx6GYyo0_2),.clk(gclk));
	jdff dff_B_qrtJTwc08_2(.din(w_dff_B_pCx6GYyo0_2),.dout(w_dff_B_qrtJTwc08_2),.clk(gclk));
	jdff dff_B_RmbCiMPF6_2(.din(w_dff_B_qrtJTwc08_2),.dout(w_dff_B_RmbCiMPF6_2),.clk(gclk));
	jdff dff_B_u4aSQSdF1_1(.din(n1328),.dout(w_dff_B_u4aSQSdF1_1),.clk(gclk));
	jdff dff_B_Cx6My3pg9_2(.din(n1242),.dout(w_dff_B_Cx6My3pg9_2),.clk(gclk));
	jdff dff_B_QXcIqmq80_2(.din(w_dff_B_Cx6My3pg9_2),.dout(w_dff_B_QXcIqmq80_2),.clk(gclk));
	jdff dff_B_kkAoFUco2_2(.din(w_dff_B_QXcIqmq80_2),.dout(w_dff_B_kkAoFUco2_2),.clk(gclk));
	jdff dff_B_P73OyyiO4_2(.din(w_dff_B_kkAoFUco2_2),.dout(w_dff_B_P73OyyiO4_2),.clk(gclk));
	jdff dff_B_CZLw1cXT6_2(.din(w_dff_B_P73OyyiO4_2),.dout(w_dff_B_CZLw1cXT6_2),.clk(gclk));
	jdff dff_B_HwFPJ4EA4_2(.din(w_dff_B_CZLw1cXT6_2),.dout(w_dff_B_HwFPJ4EA4_2),.clk(gclk));
	jdff dff_B_NrFrBWx25_2(.din(w_dff_B_HwFPJ4EA4_2),.dout(w_dff_B_NrFrBWx25_2),.clk(gclk));
	jdff dff_B_mywMtiu13_2(.din(w_dff_B_NrFrBWx25_2),.dout(w_dff_B_mywMtiu13_2),.clk(gclk));
	jdff dff_B_bB7dcx8R3_2(.din(w_dff_B_mywMtiu13_2),.dout(w_dff_B_bB7dcx8R3_2),.clk(gclk));
	jdff dff_B_uQPBbs0O3_2(.din(w_dff_B_bB7dcx8R3_2),.dout(w_dff_B_uQPBbs0O3_2),.clk(gclk));
	jdff dff_B_xN7pEiYJ9_2(.din(w_dff_B_uQPBbs0O3_2),.dout(w_dff_B_xN7pEiYJ9_2),.clk(gclk));
	jdff dff_B_fM7Yq2WQ8_2(.din(w_dff_B_xN7pEiYJ9_2),.dout(w_dff_B_fM7Yq2WQ8_2),.clk(gclk));
	jdff dff_B_aLxOuJhY3_2(.din(w_dff_B_fM7Yq2WQ8_2),.dout(w_dff_B_aLxOuJhY3_2),.clk(gclk));
	jdff dff_B_3Q4pkfNi1_2(.din(w_dff_B_aLxOuJhY3_2),.dout(w_dff_B_3Q4pkfNi1_2),.clk(gclk));
	jdff dff_B_yYhd4daa7_2(.din(w_dff_B_3Q4pkfNi1_2),.dout(w_dff_B_yYhd4daa7_2),.clk(gclk));
	jdff dff_B_ZlA9nWD81_2(.din(w_dff_B_yYhd4daa7_2),.dout(w_dff_B_ZlA9nWD81_2),.clk(gclk));
	jdff dff_B_QQcGgiGy7_2(.din(w_dff_B_ZlA9nWD81_2),.dout(w_dff_B_QQcGgiGy7_2),.clk(gclk));
	jdff dff_B_Lyn5RP2y2_2(.din(w_dff_B_QQcGgiGy7_2),.dout(w_dff_B_Lyn5RP2y2_2),.clk(gclk));
	jdff dff_B_t0tqAlfT0_2(.din(w_dff_B_Lyn5RP2y2_2),.dout(w_dff_B_t0tqAlfT0_2),.clk(gclk));
	jdff dff_B_SOP43ZMk1_2(.din(w_dff_B_t0tqAlfT0_2),.dout(w_dff_B_SOP43ZMk1_2),.clk(gclk));
	jdff dff_B_vRSC99dJ8_2(.din(w_dff_B_SOP43ZMk1_2),.dout(w_dff_B_vRSC99dJ8_2),.clk(gclk));
	jdff dff_B_pzaxuUlC1_2(.din(w_dff_B_vRSC99dJ8_2),.dout(w_dff_B_pzaxuUlC1_2),.clk(gclk));
	jdff dff_B_7NXe1aam5_1(.din(n1243),.dout(w_dff_B_7NXe1aam5_1),.clk(gclk));
	jdff dff_B_Je0dIbIX7_2(.din(n1151),.dout(w_dff_B_Je0dIbIX7_2),.clk(gclk));
	jdff dff_B_szC91N574_2(.din(w_dff_B_Je0dIbIX7_2),.dout(w_dff_B_szC91N574_2),.clk(gclk));
	jdff dff_B_LXmzBUpG3_2(.din(w_dff_B_szC91N574_2),.dout(w_dff_B_LXmzBUpG3_2),.clk(gclk));
	jdff dff_B_Ey5AIvti9_2(.din(w_dff_B_LXmzBUpG3_2),.dout(w_dff_B_Ey5AIvti9_2),.clk(gclk));
	jdff dff_B_kyz0yeSz2_2(.din(w_dff_B_Ey5AIvti9_2),.dout(w_dff_B_kyz0yeSz2_2),.clk(gclk));
	jdff dff_B_JgHuZNH30_2(.din(w_dff_B_kyz0yeSz2_2),.dout(w_dff_B_JgHuZNH30_2),.clk(gclk));
	jdff dff_B_kLGMyrwD4_2(.din(w_dff_B_JgHuZNH30_2),.dout(w_dff_B_kLGMyrwD4_2),.clk(gclk));
	jdff dff_B_5M5P6f7G8_2(.din(w_dff_B_kLGMyrwD4_2),.dout(w_dff_B_5M5P6f7G8_2),.clk(gclk));
	jdff dff_B_NRndCDC24_2(.din(w_dff_B_5M5P6f7G8_2),.dout(w_dff_B_NRndCDC24_2),.clk(gclk));
	jdff dff_B_xEyC5FTv0_2(.din(w_dff_B_NRndCDC24_2),.dout(w_dff_B_xEyC5FTv0_2),.clk(gclk));
	jdff dff_B_SmXU5iOp1_2(.din(w_dff_B_xEyC5FTv0_2),.dout(w_dff_B_SmXU5iOp1_2),.clk(gclk));
	jdff dff_B_39Wr9A6V8_2(.din(w_dff_B_SmXU5iOp1_2),.dout(w_dff_B_39Wr9A6V8_2),.clk(gclk));
	jdff dff_B_u9R9wBej9_2(.din(w_dff_B_39Wr9A6V8_2),.dout(w_dff_B_u9R9wBej9_2),.clk(gclk));
	jdff dff_B_WpCQmerQ5_2(.din(w_dff_B_u9R9wBej9_2),.dout(w_dff_B_WpCQmerQ5_2),.clk(gclk));
	jdff dff_B_9czaz7Yk1_2(.din(w_dff_B_WpCQmerQ5_2),.dout(w_dff_B_9czaz7Yk1_2),.clk(gclk));
	jdff dff_B_W8Jkh4iC0_2(.din(w_dff_B_9czaz7Yk1_2),.dout(w_dff_B_W8Jkh4iC0_2),.clk(gclk));
	jdff dff_B_i2HOhHua3_2(.din(w_dff_B_W8Jkh4iC0_2),.dout(w_dff_B_i2HOhHua3_2),.clk(gclk));
	jdff dff_B_rYLJkBLd3_2(.din(w_dff_B_i2HOhHua3_2),.dout(w_dff_B_rYLJkBLd3_2),.clk(gclk));
	jdff dff_B_eZElVmW97_2(.din(w_dff_B_rYLJkBLd3_2),.dout(w_dff_B_eZElVmW97_2),.clk(gclk));
	jdff dff_B_Sr08VwJO8_2(.din(w_dff_B_eZElVmW97_2),.dout(w_dff_B_Sr08VwJO8_2),.clk(gclk));
	jdff dff_B_qXyM7Qwc6_1(.din(n1152),.dout(w_dff_B_qXyM7Qwc6_1),.clk(gclk));
	jdff dff_B_0TvzjfHU0_2(.din(n1053),.dout(w_dff_B_0TvzjfHU0_2),.clk(gclk));
	jdff dff_B_ypmmE3C39_2(.din(w_dff_B_0TvzjfHU0_2),.dout(w_dff_B_ypmmE3C39_2),.clk(gclk));
	jdff dff_B_K1R5TRh27_2(.din(w_dff_B_ypmmE3C39_2),.dout(w_dff_B_K1R5TRh27_2),.clk(gclk));
	jdff dff_B_3n3PnFyB1_2(.din(w_dff_B_K1R5TRh27_2),.dout(w_dff_B_3n3PnFyB1_2),.clk(gclk));
	jdff dff_B_Sig101506_2(.din(w_dff_B_3n3PnFyB1_2),.dout(w_dff_B_Sig101506_2),.clk(gclk));
	jdff dff_B_bolEqkLW1_2(.din(w_dff_B_Sig101506_2),.dout(w_dff_B_bolEqkLW1_2),.clk(gclk));
	jdff dff_B_fLhQkqRH7_2(.din(w_dff_B_bolEqkLW1_2),.dout(w_dff_B_fLhQkqRH7_2),.clk(gclk));
	jdff dff_B_LHj4UaqR2_2(.din(w_dff_B_fLhQkqRH7_2),.dout(w_dff_B_LHj4UaqR2_2),.clk(gclk));
	jdff dff_B_iDje99eB5_2(.din(w_dff_B_LHj4UaqR2_2),.dout(w_dff_B_iDje99eB5_2),.clk(gclk));
	jdff dff_B_MskXIIxs6_2(.din(w_dff_B_iDje99eB5_2),.dout(w_dff_B_MskXIIxs6_2),.clk(gclk));
	jdff dff_B_Od0FDlA80_2(.din(w_dff_B_MskXIIxs6_2),.dout(w_dff_B_Od0FDlA80_2),.clk(gclk));
	jdff dff_B_SkRX7Q4g9_2(.din(w_dff_B_Od0FDlA80_2),.dout(w_dff_B_SkRX7Q4g9_2),.clk(gclk));
	jdff dff_B_Z3rNbKFV1_2(.din(w_dff_B_SkRX7Q4g9_2),.dout(w_dff_B_Z3rNbKFV1_2),.clk(gclk));
	jdff dff_B_EBMd0cWs6_2(.din(w_dff_B_Z3rNbKFV1_2),.dout(w_dff_B_EBMd0cWs6_2),.clk(gclk));
	jdff dff_B_WOqC9OdB8_2(.din(w_dff_B_EBMd0cWs6_2),.dout(w_dff_B_WOqC9OdB8_2),.clk(gclk));
	jdff dff_B_6vGPQelS1_2(.din(w_dff_B_WOqC9OdB8_2),.dout(w_dff_B_6vGPQelS1_2),.clk(gclk));
	jdff dff_B_KWjXixrE8_2(.din(w_dff_B_6vGPQelS1_2),.dout(w_dff_B_KWjXixrE8_2),.clk(gclk));
	jdff dff_B_SU75RpGS3_2(.din(w_dff_B_KWjXixrE8_2),.dout(w_dff_B_SU75RpGS3_2),.clk(gclk));
	jdff dff_B_VVYYVHft7_1(.din(n1054),.dout(w_dff_B_VVYYVHft7_1),.clk(gclk));
	jdff dff_B_BfT0IfDy2_2(.din(n954),.dout(w_dff_B_BfT0IfDy2_2),.clk(gclk));
	jdff dff_B_OXIeXVOr8_2(.din(w_dff_B_BfT0IfDy2_2),.dout(w_dff_B_OXIeXVOr8_2),.clk(gclk));
	jdff dff_B_BSdDzozM3_2(.din(w_dff_B_OXIeXVOr8_2),.dout(w_dff_B_BSdDzozM3_2),.clk(gclk));
	jdff dff_B_iNE26wtK5_2(.din(w_dff_B_BSdDzozM3_2),.dout(w_dff_B_iNE26wtK5_2),.clk(gclk));
	jdff dff_B_UNbIj7qn2_2(.din(w_dff_B_iNE26wtK5_2),.dout(w_dff_B_UNbIj7qn2_2),.clk(gclk));
	jdff dff_B_R1mUILyP9_2(.din(w_dff_B_UNbIj7qn2_2),.dout(w_dff_B_R1mUILyP9_2),.clk(gclk));
	jdff dff_B_i22bJWZf3_2(.din(w_dff_B_R1mUILyP9_2),.dout(w_dff_B_i22bJWZf3_2),.clk(gclk));
	jdff dff_B_XOmWZpx17_2(.din(w_dff_B_i22bJWZf3_2),.dout(w_dff_B_XOmWZpx17_2),.clk(gclk));
	jdff dff_B_Clb3lzXg2_2(.din(w_dff_B_XOmWZpx17_2),.dout(w_dff_B_Clb3lzXg2_2),.clk(gclk));
	jdff dff_B_Y5DmB6y44_2(.din(w_dff_B_Clb3lzXg2_2),.dout(w_dff_B_Y5DmB6y44_2),.clk(gclk));
	jdff dff_B_l1NKi4vi9_2(.din(w_dff_B_Y5DmB6y44_2),.dout(w_dff_B_l1NKi4vi9_2),.clk(gclk));
	jdff dff_B_4wDrXFRU9_2(.din(w_dff_B_l1NKi4vi9_2),.dout(w_dff_B_4wDrXFRU9_2),.clk(gclk));
	jdff dff_B_KuIwdfcf8_2(.din(w_dff_B_4wDrXFRU9_2),.dout(w_dff_B_KuIwdfcf8_2),.clk(gclk));
	jdff dff_B_s7sd3LNW0_2(.din(w_dff_B_KuIwdfcf8_2),.dout(w_dff_B_s7sd3LNW0_2),.clk(gclk));
	jdff dff_B_qcPQIcQb7_2(.din(w_dff_B_s7sd3LNW0_2),.dout(w_dff_B_qcPQIcQb7_2),.clk(gclk));
	jdff dff_B_7EOlVDn41_2(.din(w_dff_B_qcPQIcQb7_2),.dout(w_dff_B_7EOlVDn41_2),.clk(gclk));
	jdff dff_B_QeeoHfcw0_1(.din(n955),.dout(w_dff_B_QeeoHfcw0_1),.clk(gclk));
	jdff dff_B_r1S7Xluw5_2(.din(n852),.dout(w_dff_B_r1S7Xluw5_2),.clk(gclk));
	jdff dff_B_6zsibY9X8_2(.din(w_dff_B_r1S7Xluw5_2),.dout(w_dff_B_6zsibY9X8_2),.clk(gclk));
	jdff dff_B_emK3KRQX6_2(.din(w_dff_B_6zsibY9X8_2),.dout(w_dff_B_emK3KRQX6_2),.clk(gclk));
	jdff dff_B_TIZwAch08_2(.din(w_dff_B_emK3KRQX6_2),.dout(w_dff_B_TIZwAch08_2),.clk(gclk));
	jdff dff_B_B73Ro9kn2_2(.din(w_dff_B_TIZwAch08_2),.dout(w_dff_B_B73Ro9kn2_2),.clk(gclk));
	jdff dff_B_LlOJyFvd9_2(.din(w_dff_B_B73Ro9kn2_2),.dout(w_dff_B_LlOJyFvd9_2),.clk(gclk));
	jdff dff_B_rTAbZuoW4_2(.din(w_dff_B_LlOJyFvd9_2),.dout(w_dff_B_rTAbZuoW4_2),.clk(gclk));
	jdff dff_B_Tt00uwKb7_2(.din(w_dff_B_rTAbZuoW4_2),.dout(w_dff_B_Tt00uwKb7_2),.clk(gclk));
	jdff dff_B_0GwSHv5V9_2(.din(w_dff_B_Tt00uwKb7_2),.dout(w_dff_B_0GwSHv5V9_2),.clk(gclk));
	jdff dff_B_lm4pPCWv7_2(.din(w_dff_B_0GwSHv5V9_2),.dout(w_dff_B_lm4pPCWv7_2),.clk(gclk));
	jdff dff_B_fQTOUhIF3_2(.din(w_dff_B_lm4pPCWv7_2),.dout(w_dff_B_fQTOUhIF3_2),.clk(gclk));
	jdff dff_B_wIS1m3YM7_2(.din(w_dff_B_fQTOUhIF3_2),.dout(w_dff_B_wIS1m3YM7_2),.clk(gclk));
	jdff dff_B_S7K19t8L1_2(.din(w_dff_B_wIS1m3YM7_2),.dout(w_dff_B_S7K19t8L1_2),.clk(gclk));
	jdff dff_B_44BG7z7r0_2(.din(w_dff_B_S7K19t8L1_2),.dout(w_dff_B_44BG7z7r0_2),.clk(gclk));
	jdff dff_B_KBFvPjWb1_1(.din(n853),.dout(w_dff_B_KBFvPjWb1_1),.clk(gclk));
	jdff dff_B_D2sIU5y97_2(.din(n754),.dout(w_dff_B_D2sIU5y97_2),.clk(gclk));
	jdff dff_B_EVx0lc9W5_2(.din(w_dff_B_D2sIU5y97_2),.dout(w_dff_B_EVx0lc9W5_2),.clk(gclk));
	jdff dff_B_2nkXRlqF9_2(.din(w_dff_B_EVx0lc9W5_2),.dout(w_dff_B_2nkXRlqF9_2),.clk(gclk));
	jdff dff_B_bAttG5yd2_2(.din(w_dff_B_2nkXRlqF9_2),.dout(w_dff_B_bAttG5yd2_2),.clk(gclk));
	jdff dff_B_76T5mV5z6_2(.din(w_dff_B_bAttG5yd2_2),.dout(w_dff_B_76T5mV5z6_2),.clk(gclk));
	jdff dff_B_Z2P859FC9_2(.din(w_dff_B_76T5mV5z6_2),.dout(w_dff_B_Z2P859FC9_2),.clk(gclk));
	jdff dff_B_3bHjqqJB5_2(.din(w_dff_B_Z2P859FC9_2),.dout(w_dff_B_3bHjqqJB5_2),.clk(gclk));
	jdff dff_B_j9H94ud07_2(.din(w_dff_B_3bHjqqJB5_2),.dout(w_dff_B_j9H94ud07_2),.clk(gclk));
	jdff dff_B_0xnVnBxE4_2(.din(w_dff_B_j9H94ud07_2),.dout(w_dff_B_0xnVnBxE4_2),.clk(gclk));
	jdff dff_B_H5M5tGWS7_2(.din(w_dff_B_0xnVnBxE4_2),.dout(w_dff_B_H5M5tGWS7_2),.clk(gclk));
	jdff dff_B_IAEuopXa7_2(.din(w_dff_B_H5M5tGWS7_2),.dout(w_dff_B_IAEuopXa7_2),.clk(gclk));
	jdff dff_B_sglmE4pR1_2(.din(w_dff_B_IAEuopXa7_2),.dout(w_dff_B_sglmE4pR1_2),.clk(gclk));
	jdff dff_B_rotSg5d82_1(.din(n755),.dout(w_dff_B_rotSg5d82_1),.clk(gclk));
	jdff dff_B_XxAVYfDU5_2(.din(n662),.dout(w_dff_B_XxAVYfDU5_2),.clk(gclk));
	jdff dff_B_S2EemTn48_2(.din(w_dff_B_XxAVYfDU5_2),.dout(w_dff_B_S2EemTn48_2),.clk(gclk));
	jdff dff_B_cygVIqK89_2(.din(w_dff_B_S2EemTn48_2),.dout(w_dff_B_cygVIqK89_2),.clk(gclk));
	jdff dff_B_sFRzDL4a8_2(.din(w_dff_B_cygVIqK89_2),.dout(w_dff_B_sFRzDL4a8_2),.clk(gclk));
	jdff dff_B_jV1cZg2Q9_2(.din(w_dff_B_sFRzDL4a8_2),.dout(w_dff_B_jV1cZg2Q9_2),.clk(gclk));
	jdff dff_B_VNar4xOi1_2(.din(w_dff_B_jV1cZg2Q9_2),.dout(w_dff_B_VNar4xOi1_2),.clk(gclk));
	jdff dff_B_z6V0r9oE0_2(.din(w_dff_B_VNar4xOi1_2),.dout(w_dff_B_z6V0r9oE0_2),.clk(gclk));
	jdff dff_B_O7dbEXDU5_2(.din(w_dff_B_z6V0r9oE0_2),.dout(w_dff_B_O7dbEXDU5_2),.clk(gclk));
	jdff dff_B_oVoN5YBR6_2(.din(w_dff_B_O7dbEXDU5_2),.dout(w_dff_B_oVoN5YBR6_2),.clk(gclk));
	jdff dff_B_z6gQ9hNy3_2(.din(w_dff_B_oVoN5YBR6_2),.dout(w_dff_B_z6gQ9hNy3_2),.clk(gclk));
	jdff dff_B_WREzFNmg8_1(.din(n663),.dout(w_dff_B_WREzFNmg8_1),.clk(gclk));
	jdff dff_B_K1M8SoWB3_2(.din(n577),.dout(w_dff_B_K1M8SoWB3_2),.clk(gclk));
	jdff dff_B_wx5N0beU2_2(.din(w_dff_B_K1M8SoWB3_2),.dout(w_dff_B_wx5N0beU2_2),.clk(gclk));
	jdff dff_B_Z8JK565X9_2(.din(w_dff_B_wx5N0beU2_2),.dout(w_dff_B_Z8JK565X9_2),.clk(gclk));
	jdff dff_B_nZiFLd5J9_2(.din(w_dff_B_Z8JK565X9_2),.dout(w_dff_B_nZiFLd5J9_2),.clk(gclk));
	jdff dff_B_P4GtX4Xi9_2(.din(w_dff_B_nZiFLd5J9_2),.dout(w_dff_B_P4GtX4Xi9_2),.clk(gclk));
	jdff dff_B_Z1Kc7rXZ8_2(.din(w_dff_B_P4GtX4Xi9_2),.dout(w_dff_B_Z1Kc7rXZ8_2),.clk(gclk));
	jdff dff_B_RmGjfVPt2_2(.din(w_dff_B_Z1Kc7rXZ8_2),.dout(w_dff_B_RmGjfVPt2_2),.clk(gclk));
	jdff dff_B_1NLc7XxL1_2(.din(w_dff_B_RmGjfVPt2_2),.dout(w_dff_B_1NLc7XxL1_2),.clk(gclk));
	jdff dff_B_i8R0CmxG1_2(.din(n592),.dout(w_dff_B_i8R0CmxG1_2),.clk(gclk));
	jdff dff_B_7Rufg3Uj7_2(.din(w_dff_B_i8R0CmxG1_2),.dout(w_dff_B_7Rufg3Uj7_2),.clk(gclk));
	jdff dff_B_N5Yqmrr39_2(.din(w_dff_B_7Rufg3Uj7_2),.dout(w_dff_B_N5Yqmrr39_2),.clk(gclk));
	jdff dff_B_NUrjUkee4_1(.din(n578),.dout(w_dff_B_NUrjUkee4_1),.clk(gclk));
	jdff dff_B_l32r1WdK3_1(.din(w_dff_B_NUrjUkee4_1),.dout(w_dff_B_l32r1WdK3_1),.clk(gclk));
	jdff dff_B_VFNjns4h3_1(.din(w_dff_B_l32r1WdK3_1),.dout(w_dff_B_VFNjns4h3_1),.clk(gclk));
	jdff dff_B_SdMVL1by0_2(.din(n501),.dout(w_dff_B_SdMVL1by0_2),.clk(gclk));
	jdff dff_B_dM63tieg8_2(.din(w_dff_B_SdMVL1by0_2),.dout(w_dff_B_dM63tieg8_2),.clk(gclk));
	jdff dff_B_tds3ch0X2_2(.din(w_dff_B_dM63tieg8_2),.dout(w_dff_B_tds3ch0X2_2),.clk(gclk));
	jdff dff_B_RsaZpdi96_0(.din(n506),.dout(w_dff_B_RsaZpdi96_0),.clk(gclk));
	jdff dff_B_fr6mKTAI4_0(.din(w_dff_B_RsaZpdi96_0),.dout(w_dff_B_fr6mKTAI4_0),.clk(gclk));
	jdff dff_A_3Gg0Z0b75_0(.dout(w_n427_0[0]),.din(w_dff_A_3Gg0Z0b75_0),.clk(gclk));
	jdff dff_A_MVF4fcjn7_0(.dout(w_dff_A_3Gg0Z0b75_0),.din(w_dff_A_MVF4fcjn7_0),.clk(gclk));
	jdff dff_A_VINnGMiS2_1(.dout(w_n427_0[1]),.din(w_dff_A_VINnGMiS2_1),.clk(gclk));
	jdff dff_A_BMAwMXjb2_1(.dout(w_dff_A_VINnGMiS2_1),.din(w_dff_A_BMAwMXjb2_1),.clk(gclk));
	jdff dff_B_PE4m5ZCu8_1(.din(n1729),.dout(w_dff_B_PE4m5ZCu8_1),.clk(gclk));
	jdff dff_A_csoi6cFm2_1(.dout(w_n1697_0[1]),.din(w_dff_A_csoi6cFm2_1),.clk(gclk));
	jdff dff_B_32RUcBr69_1(.din(n1695),.dout(w_dff_B_32RUcBr69_1),.clk(gclk));
	jdff dff_B_QFG62Yqq9_2(.din(n1653),.dout(w_dff_B_QFG62Yqq9_2),.clk(gclk));
	jdff dff_B_Ilcs4dY33_2(.din(w_dff_B_QFG62Yqq9_2),.dout(w_dff_B_Ilcs4dY33_2),.clk(gclk));
	jdff dff_B_QxHhpsNM5_2(.din(w_dff_B_Ilcs4dY33_2),.dout(w_dff_B_QxHhpsNM5_2),.clk(gclk));
	jdff dff_B_v44tIc602_2(.din(w_dff_B_QxHhpsNM5_2),.dout(w_dff_B_v44tIc602_2),.clk(gclk));
	jdff dff_B_Flk4j5qc4_2(.din(w_dff_B_v44tIc602_2),.dout(w_dff_B_Flk4j5qc4_2),.clk(gclk));
	jdff dff_B_kXpcI2eY9_2(.din(w_dff_B_Flk4j5qc4_2),.dout(w_dff_B_kXpcI2eY9_2),.clk(gclk));
	jdff dff_B_4BQSOL2l2_2(.din(w_dff_B_kXpcI2eY9_2),.dout(w_dff_B_4BQSOL2l2_2),.clk(gclk));
	jdff dff_B_aTFLY3PB2_2(.din(w_dff_B_4BQSOL2l2_2),.dout(w_dff_B_aTFLY3PB2_2),.clk(gclk));
	jdff dff_B_VLvrWuPZ5_2(.din(w_dff_B_aTFLY3PB2_2),.dout(w_dff_B_VLvrWuPZ5_2),.clk(gclk));
	jdff dff_B_61sxVVWt4_2(.din(w_dff_B_VLvrWuPZ5_2),.dout(w_dff_B_61sxVVWt4_2),.clk(gclk));
	jdff dff_B_5QzWkgxD5_2(.din(w_dff_B_61sxVVWt4_2),.dout(w_dff_B_5QzWkgxD5_2),.clk(gclk));
	jdff dff_B_qHmSAEz46_2(.din(w_dff_B_5QzWkgxD5_2),.dout(w_dff_B_qHmSAEz46_2),.clk(gclk));
	jdff dff_B_s9zqOVEC5_2(.din(w_dff_B_qHmSAEz46_2),.dout(w_dff_B_s9zqOVEC5_2),.clk(gclk));
	jdff dff_B_XO13hPQY3_2(.din(w_dff_B_s9zqOVEC5_2),.dout(w_dff_B_XO13hPQY3_2),.clk(gclk));
	jdff dff_B_cSGCRgcZ1_2(.din(w_dff_B_XO13hPQY3_2),.dout(w_dff_B_cSGCRgcZ1_2),.clk(gclk));
	jdff dff_B_7pBR1iIP9_2(.din(w_dff_B_cSGCRgcZ1_2),.dout(w_dff_B_7pBR1iIP9_2),.clk(gclk));
	jdff dff_B_e7xPARvF0_2(.din(w_dff_B_7pBR1iIP9_2),.dout(w_dff_B_e7xPARvF0_2),.clk(gclk));
	jdff dff_B_WRyTq3sK4_2(.din(w_dff_B_e7xPARvF0_2),.dout(w_dff_B_WRyTq3sK4_2),.clk(gclk));
	jdff dff_B_KE67mPxR4_2(.din(w_dff_B_WRyTq3sK4_2),.dout(w_dff_B_KE67mPxR4_2),.clk(gclk));
	jdff dff_B_PLxFEBDJ1_2(.din(w_dff_B_KE67mPxR4_2),.dout(w_dff_B_PLxFEBDJ1_2),.clk(gclk));
	jdff dff_B_k4wOFEZD3_2(.din(w_dff_B_PLxFEBDJ1_2),.dout(w_dff_B_k4wOFEZD3_2),.clk(gclk));
	jdff dff_B_mklHn2su3_2(.din(w_dff_B_k4wOFEZD3_2),.dout(w_dff_B_mklHn2su3_2),.clk(gclk));
	jdff dff_B_ip3aEDJF2_2(.din(w_dff_B_mklHn2su3_2),.dout(w_dff_B_ip3aEDJF2_2),.clk(gclk));
	jdff dff_B_rPDyahFY4_2(.din(w_dff_B_ip3aEDJF2_2),.dout(w_dff_B_rPDyahFY4_2),.clk(gclk));
	jdff dff_B_Mf5Wy88i1_2(.din(w_dff_B_rPDyahFY4_2),.dout(w_dff_B_Mf5Wy88i1_2),.clk(gclk));
	jdff dff_B_joXVuqhp2_2(.din(w_dff_B_Mf5Wy88i1_2),.dout(w_dff_B_joXVuqhp2_2),.clk(gclk));
	jdff dff_B_FECT2AFU8_2(.din(w_dff_B_joXVuqhp2_2),.dout(w_dff_B_FECT2AFU8_2),.clk(gclk));
	jdff dff_B_vRZxbveO2_2(.din(w_dff_B_FECT2AFU8_2),.dout(w_dff_B_vRZxbveO2_2),.clk(gclk));
	jdff dff_B_EYgmD8Ne1_2(.din(w_dff_B_vRZxbveO2_2),.dout(w_dff_B_EYgmD8Ne1_2),.clk(gclk));
	jdff dff_B_Ezudp3L23_2(.din(w_dff_B_EYgmD8Ne1_2),.dout(w_dff_B_Ezudp3L23_2),.clk(gclk));
	jdff dff_B_BwBQcOWF6_2(.din(w_dff_B_Ezudp3L23_2),.dout(w_dff_B_BwBQcOWF6_2),.clk(gclk));
	jdff dff_B_5ZcHfyEw7_2(.din(w_dff_B_BwBQcOWF6_2),.dout(w_dff_B_5ZcHfyEw7_2),.clk(gclk));
	jdff dff_B_kHEsQ9Ld2_2(.din(w_dff_B_5ZcHfyEw7_2),.dout(w_dff_B_kHEsQ9Ld2_2),.clk(gclk));
	jdff dff_B_mdSCRtuO2_2(.din(w_dff_B_kHEsQ9Ld2_2),.dout(w_dff_B_mdSCRtuO2_2),.clk(gclk));
	jdff dff_B_j3rHZW2q5_2(.din(w_dff_B_mdSCRtuO2_2),.dout(w_dff_B_j3rHZW2q5_2),.clk(gclk));
	jdff dff_B_62HyjOUL2_2(.din(w_dff_B_j3rHZW2q5_2),.dout(w_dff_B_62HyjOUL2_2),.clk(gclk));
	jdff dff_B_9b7f8n6n3_2(.din(w_dff_B_62HyjOUL2_2),.dout(w_dff_B_9b7f8n6n3_2),.clk(gclk));
	jdff dff_B_ezdYGMnN4_2(.din(n1656),.dout(w_dff_B_ezdYGMnN4_2),.clk(gclk));
	jdff dff_B_QOTySqd87_1(.din(n1654),.dout(w_dff_B_QOTySqd87_1),.clk(gclk));
	jdff dff_B_snGtzBvx5_2(.din(n1602),.dout(w_dff_B_snGtzBvx5_2),.clk(gclk));
	jdff dff_B_NBysoQ4p3_2(.din(w_dff_B_snGtzBvx5_2),.dout(w_dff_B_NBysoQ4p3_2),.clk(gclk));
	jdff dff_B_gDaZSkVr3_2(.din(w_dff_B_NBysoQ4p3_2),.dout(w_dff_B_gDaZSkVr3_2),.clk(gclk));
	jdff dff_B_TEbkZlle4_2(.din(w_dff_B_gDaZSkVr3_2),.dout(w_dff_B_TEbkZlle4_2),.clk(gclk));
	jdff dff_B_bHn8kcXD5_2(.din(w_dff_B_TEbkZlle4_2),.dout(w_dff_B_bHn8kcXD5_2),.clk(gclk));
	jdff dff_B_LBRinYkX5_2(.din(w_dff_B_bHn8kcXD5_2),.dout(w_dff_B_LBRinYkX5_2),.clk(gclk));
	jdff dff_B_4prf02q09_2(.din(w_dff_B_LBRinYkX5_2),.dout(w_dff_B_4prf02q09_2),.clk(gclk));
	jdff dff_B_M3dqth1M4_2(.din(w_dff_B_4prf02q09_2),.dout(w_dff_B_M3dqth1M4_2),.clk(gclk));
	jdff dff_B_gRGnvf8h5_2(.din(w_dff_B_M3dqth1M4_2),.dout(w_dff_B_gRGnvf8h5_2),.clk(gclk));
	jdff dff_B_rpwoirJ62_2(.din(w_dff_B_gRGnvf8h5_2),.dout(w_dff_B_rpwoirJ62_2),.clk(gclk));
	jdff dff_B_I7PBHofI5_2(.din(w_dff_B_rpwoirJ62_2),.dout(w_dff_B_I7PBHofI5_2),.clk(gclk));
	jdff dff_B_oViZ8m8C6_2(.din(w_dff_B_I7PBHofI5_2),.dout(w_dff_B_oViZ8m8C6_2),.clk(gclk));
	jdff dff_B_55RINX5E8_2(.din(w_dff_B_oViZ8m8C6_2),.dout(w_dff_B_55RINX5E8_2),.clk(gclk));
	jdff dff_B_mvEzyRlR7_2(.din(w_dff_B_55RINX5E8_2),.dout(w_dff_B_mvEzyRlR7_2),.clk(gclk));
	jdff dff_B_zefmrKuf7_2(.din(w_dff_B_mvEzyRlR7_2),.dout(w_dff_B_zefmrKuf7_2),.clk(gclk));
	jdff dff_B_3QkWOUJC9_2(.din(w_dff_B_zefmrKuf7_2),.dout(w_dff_B_3QkWOUJC9_2),.clk(gclk));
	jdff dff_B_x8JYUs909_2(.din(w_dff_B_3QkWOUJC9_2),.dout(w_dff_B_x8JYUs909_2),.clk(gclk));
	jdff dff_B_eAFvx1Xe2_2(.din(w_dff_B_x8JYUs909_2),.dout(w_dff_B_eAFvx1Xe2_2),.clk(gclk));
	jdff dff_B_pxEy49Oz7_2(.din(w_dff_B_eAFvx1Xe2_2),.dout(w_dff_B_pxEy49Oz7_2),.clk(gclk));
	jdff dff_B_uqD9fGBQ8_2(.din(w_dff_B_pxEy49Oz7_2),.dout(w_dff_B_uqD9fGBQ8_2),.clk(gclk));
	jdff dff_B_Y5uPpjE31_2(.din(w_dff_B_uqD9fGBQ8_2),.dout(w_dff_B_Y5uPpjE31_2),.clk(gclk));
	jdff dff_B_1mgMYVK02_2(.din(w_dff_B_Y5uPpjE31_2),.dout(w_dff_B_1mgMYVK02_2),.clk(gclk));
	jdff dff_B_S2zN05ch2_2(.din(w_dff_B_1mgMYVK02_2),.dout(w_dff_B_S2zN05ch2_2),.clk(gclk));
	jdff dff_B_1RI0rbVI0_2(.din(w_dff_B_S2zN05ch2_2),.dout(w_dff_B_1RI0rbVI0_2),.clk(gclk));
	jdff dff_B_FWbA67yj3_2(.din(w_dff_B_1RI0rbVI0_2),.dout(w_dff_B_FWbA67yj3_2),.clk(gclk));
	jdff dff_B_xHyk3nty9_2(.din(w_dff_B_FWbA67yj3_2),.dout(w_dff_B_xHyk3nty9_2),.clk(gclk));
	jdff dff_B_SFSMzVUo6_2(.din(w_dff_B_xHyk3nty9_2),.dout(w_dff_B_SFSMzVUo6_2),.clk(gclk));
	jdff dff_B_HDWKiVzy6_2(.din(w_dff_B_SFSMzVUo6_2),.dout(w_dff_B_HDWKiVzy6_2),.clk(gclk));
	jdff dff_B_jlh42iic2_2(.din(w_dff_B_HDWKiVzy6_2),.dout(w_dff_B_jlh42iic2_2),.clk(gclk));
	jdff dff_B_mIy2pGjT3_2(.din(w_dff_B_jlh42iic2_2),.dout(w_dff_B_mIy2pGjT3_2),.clk(gclk));
	jdff dff_B_0ztbaOph2_2(.din(w_dff_B_mIy2pGjT3_2),.dout(w_dff_B_0ztbaOph2_2),.clk(gclk));
	jdff dff_B_0FNj0ARD4_2(.din(w_dff_B_0ztbaOph2_2),.dout(w_dff_B_0FNj0ARD4_2),.clk(gclk));
	jdff dff_B_2iv5EmEG0_2(.din(w_dff_B_0FNj0ARD4_2),.dout(w_dff_B_2iv5EmEG0_2),.clk(gclk));
	jdff dff_B_wbcx4oOg9_2(.din(w_dff_B_2iv5EmEG0_2),.dout(w_dff_B_wbcx4oOg9_2),.clk(gclk));
	jdff dff_B_Jm07S3Nn1_2(.din(n1605),.dout(w_dff_B_Jm07S3Nn1_2),.clk(gclk));
	jdff dff_B_m01alN119_1(.din(n1603),.dout(w_dff_B_m01alN119_1),.clk(gclk));
	jdff dff_B_ermCbF732_2(.din(n1545),.dout(w_dff_B_ermCbF732_2),.clk(gclk));
	jdff dff_B_ZBX9aFZ51_2(.din(w_dff_B_ermCbF732_2),.dout(w_dff_B_ZBX9aFZ51_2),.clk(gclk));
	jdff dff_B_YFzwZPHy3_2(.din(w_dff_B_ZBX9aFZ51_2),.dout(w_dff_B_YFzwZPHy3_2),.clk(gclk));
	jdff dff_B_mImqg4pu8_2(.din(w_dff_B_YFzwZPHy3_2),.dout(w_dff_B_mImqg4pu8_2),.clk(gclk));
	jdff dff_B_FO0qQGWH9_2(.din(w_dff_B_mImqg4pu8_2),.dout(w_dff_B_FO0qQGWH9_2),.clk(gclk));
	jdff dff_B_2EoKPnfP0_2(.din(w_dff_B_FO0qQGWH9_2),.dout(w_dff_B_2EoKPnfP0_2),.clk(gclk));
	jdff dff_B_eecEN4h19_2(.din(w_dff_B_2EoKPnfP0_2),.dout(w_dff_B_eecEN4h19_2),.clk(gclk));
	jdff dff_B_8ZCZzsU97_2(.din(w_dff_B_eecEN4h19_2),.dout(w_dff_B_8ZCZzsU97_2),.clk(gclk));
	jdff dff_B_gZpl0MII6_2(.din(w_dff_B_8ZCZzsU97_2),.dout(w_dff_B_gZpl0MII6_2),.clk(gclk));
	jdff dff_B_5h4jZKRI8_2(.din(w_dff_B_gZpl0MII6_2),.dout(w_dff_B_5h4jZKRI8_2),.clk(gclk));
	jdff dff_B_xXzivMBD0_2(.din(w_dff_B_5h4jZKRI8_2),.dout(w_dff_B_xXzivMBD0_2),.clk(gclk));
	jdff dff_B_mPOjsurX1_2(.din(w_dff_B_xXzivMBD0_2),.dout(w_dff_B_mPOjsurX1_2),.clk(gclk));
	jdff dff_B_XcVyYVsk9_2(.din(w_dff_B_mPOjsurX1_2),.dout(w_dff_B_XcVyYVsk9_2),.clk(gclk));
	jdff dff_B_BqVaqLSy3_2(.din(w_dff_B_XcVyYVsk9_2),.dout(w_dff_B_BqVaqLSy3_2),.clk(gclk));
	jdff dff_B_lz6MFlZF6_2(.din(w_dff_B_BqVaqLSy3_2),.dout(w_dff_B_lz6MFlZF6_2),.clk(gclk));
	jdff dff_B_cmQc13Iz5_2(.din(w_dff_B_lz6MFlZF6_2),.dout(w_dff_B_cmQc13Iz5_2),.clk(gclk));
	jdff dff_B_YrCD7PYW2_2(.din(w_dff_B_cmQc13Iz5_2),.dout(w_dff_B_YrCD7PYW2_2),.clk(gclk));
	jdff dff_B_vCbtqf1q7_2(.din(w_dff_B_YrCD7PYW2_2),.dout(w_dff_B_vCbtqf1q7_2),.clk(gclk));
	jdff dff_B_pp9o9R0J7_2(.din(w_dff_B_vCbtqf1q7_2),.dout(w_dff_B_pp9o9R0J7_2),.clk(gclk));
	jdff dff_B_Rk3wQcSV7_2(.din(w_dff_B_pp9o9R0J7_2),.dout(w_dff_B_Rk3wQcSV7_2),.clk(gclk));
	jdff dff_B_uphxZ8yQ8_2(.din(w_dff_B_Rk3wQcSV7_2),.dout(w_dff_B_uphxZ8yQ8_2),.clk(gclk));
	jdff dff_B_LQgzsqpU9_2(.din(w_dff_B_uphxZ8yQ8_2),.dout(w_dff_B_LQgzsqpU9_2),.clk(gclk));
	jdff dff_B_jBGzCqon4_2(.din(w_dff_B_LQgzsqpU9_2),.dout(w_dff_B_jBGzCqon4_2),.clk(gclk));
	jdff dff_B_vVDunm8L6_2(.din(w_dff_B_jBGzCqon4_2),.dout(w_dff_B_vVDunm8L6_2),.clk(gclk));
	jdff dff_B_NTVXSH8x3_2(.din(w_dff_B_vVDunm8L6_2),.dout(w_dff_B_NTVXSH8x3_2),.clk(gclk));
	jdff dff_B_0KlK6uy33_2(.din(w_dff_B_NTVXSH8x3_2),.dout(w_dff_B_0KlK6uy33_2),.clk(gclk));
	jdff dff_B_gRXbMaD91_2(.din(w_dff_B_0KlK6uy33_2),.dout(w_dff_B_gRXbMaD91_2),.clk(gclk));
	jdff dff_B_Y2I6Z5fF7_2(.din(w_dff_B_gRXbMaD91_2),.dout(w_dff_B_Y2I6Z5fF7_2),.clk(gclk));
	jdff dff_B_NkJEGTb19_2(.din(w_dff_B_Y2I6Z5fF7_2),.dout(w_dff_B_NkJEGTb19_2),.clk(gclk));
	jdff dff_B_GbV6ToqS5_2(.din(w_dff_B_NkJEGTb19_2),.dout(w_dff_B_GbV6ToqS5_2),.clk(gclk));
	jdff dff_B_bx6MHFYJ5_2(.din(w_dff_B_GbV6ToqS5_2),.dout(w_dff_B_bx6MHFYJ5_2),.clk(gclk));
	jdff dff_B_5R5a4ZnB0_2(.din(n1548),.dout(w_dff_B_5R5a4ZnB0_2),.clk(gclk));
	jdff dff_B_3kuIQJaL6_1(.din(n1546),.dout(w_dff_B_3kuIQJaL6_1),.clk(gclk));
	jdff dff_B_Nx6prODT8_2(.din(n1481),.dout(w_dff_B_Nx6prODT8_2),.clk(gclk));
	jdff dff_B_MmvvBlnb3_2(.din(w_dff_B_Nx6prODT8_2),.dout(w_dff_B_MmvvBlnb3_2),.clk(gclk));
	jdff dff_B_L1ubTD0n1_2(.din(w_dff_B_MmvvBlnb3_2),.dout(w_dff_B_L1ubTD0n1_2),.clk(gclk));
	jdff dff_B_vxl184fQ4_2(.din(w_dff_B_L1ubTD0n1_2),.dout(w_dff_B_vxl184fQ4_2),.clk(gclk));
	jdff dff_B_DXTahOtP4_2(.din(w_dff_B_vxl184fQ4_2),.dout(w_dff_B_DXTahOtP4_2),.clk(gclk));
	jdff dff_B_F5VknJy19_2(.din(w_dff_B_DXTahOtP4_2),.dout(w_dff_B_F5VknJy19_2),.clk(gclk));
	jdff dff_B_g2fWq3F15_2(.din(w_dff_B_F5VknJy19_2),.dout(w_dff_B_g2fWq3F15_2),.clk(gclk));
	jdff dff_B_mFRTmooO7_2(.din(w_dff_B_g2fWq3F15_2),.dout(w_dff_B_mFRTmooO7_2),.clk(gclk));
	jdff dff_B_Latnbfx71_2(.din(w_dff_B_mFRTmooO7_2),.dout(w_dff_B_Latnbfx71_2),.clk(gclk));
	jdff dff_B_Erg1BIIt3_2(.din(w_dff_B_Latnbfx71_2),.dout(w_dff_B_Erg1BIIt3_2),.clk(gclk));
	jdff dff_B_uu3iam9e8_2(.din(w_dff_B_Erg1BIIt3_2),.dout(w_dff_B_uu3iam9e8_2),.clk(gclk));
	jdff dff_B_owth1e5B6_2(.din(w_dff_B_uu3iam9e8_2),.dout(w_dff_B_owth1e5B6_2),.clk(gclk));
	jdff dff_B_GaxctY0k4_2(.din(w_dff_B_owth1e5B6_2),.dout(w_dff_B_GaxctY0k4_2),.clk(gclk));
	jdff dff_B_HEKkRr1X2_2(.din(w_dff_B_GaxctY0k4_2),.dout(w_dff_B_HEKkRr1X2_2),.clk(gclk));
	jdff dff_B_AmlPPiku1_2(.din(w_dff_B_HEKkRr1X2_2),.dout(w_dff_B_AmlPPiku1_2),.clk(gclk));
	jdff dff_B_natso62S0_2(.din(w_dff_B_AmlPPiku1_2),.dout(w_dff_B_natso62S0_2),.clk(gclk));
	jdff dff_B_pK1nzeUa4_2(.din(w_dff_B_natso62S0_2),.dout(w_dff_B_pK1nzeUa4_2),.clk(gclk));
	jdff dff_B_cmARzKOa5_2(.din(w_dff_B_pK1nzeUa4_2),.dout(w_dff_B_cmARzKOa5_2),.clk(gclk));
	jdff dff_B_ocWjzMWV2_2(.din(w_dff_B_cmARzKOa5_2),.dout(w_dff_B_ocWjzMWV2_2),.clk(gclk));
	jdff dff_B_aD68uE3Q9_2(.din(w_dff_B_ocWjzMWV2_2),.dout(w_dff_B_aD68uE3Q9_2),.clk(gclk));
	jdff dff_B_n4EjIrH36_2(.din(w_dff_B_aD68uE3Q9_2),.dout(w_dff_B_n4EjIrH36_2),.clk(gclk));
	jdff dff_B_8fwdlhds5_2(.din(w_dff_B_n4EjIrH36_2),.dout(w_dff_B_8fwdlhds5_2),.clk(gclk));
	jdff dff_B_olnEJeUQ0_2(.din(w_dff_B_8fwdlhds5_2),.dout(w_dff_B_olnEJeUQ0_2),.clk(gclk));
	jdff dff_B_1Aunm1g73_2(.din(w_dff_B_olnEJeUQ0_2),.dout(w_dff_B_1Aunm1g73_2),.clk(gclk));
	jdff dff_B_8zQr2RJb9_2(.din(w_dff_B_1Aunm1g73_2),.dout(w_dff_B_8zQr2RJb9_2),.clk(gclk));
	jdff dff_B_AABk88Ph4_2(.din(w_dff_B_8zQr2RJb9_2),.dout(w_dff_B_AABk88Ph4_2),.clk(gclk));
	jdff dff_B_0G3pVopU8_2(.din(w_dff_B_AABk88Ph4_2),.dout(w_dff_B_0G3pVopU8_2),.clk(gclk));
	jdff dff_B_meCKv3YC1_2(.din(w_dff_B_0G3pVopU8_2),.dout(w_dff_B_meCKv3YC1_2),.clk(gclk));
	jdff dff_B_yYSeLr7z7_2(.din(n1484),.dout(w_dff_B_yYSeLr7z7_2),.clk(gclk));
	jdff dff_B_RIrmifht4_1(.din(n1482),.dout(w_dff_B_RIrmifht4_1),.clk(gclk));
	jdff dff_B_7kgFtJlb4_2(.din(n1410),.dout(w_dff_B_7kgFtJlb4_2),.clk(gclk));
	jdff dff_B_5PzBCSYi1_2(.din(w_dff_B_7kgFtJlb4_2),.dout(w_dff_B_5PzBCSYi1_2),.clk(gclk));
	jdff dff_B_O4CBBEIG3_2(.din(w_dff_B_5PzBCSYi1_2),.dout(w_dff_B_O4CBBEIG3_2),.clk(gclk));
	jdff dff_B_7Et7zRrX0_2(.din(w_dff_B_O4CBBEIG3_2),.dout(w_dff_B_7Et7zRrX0_2),.clk(gclk));
	jdff dff_B_N8nFr6Ah9_2(.din(w_dff_B_7Et7zRrX0_2),.dout(w_dff_B_N8nFr6Ah9_2),.clk(gclk));
	jdff dff_B_qS3xw9qH4_2(.din(w_dff_B_N8nFr6Ah9_2),.dout(w_dff_B_qS3xw9qH4_2),.clk(gclk));
	jdff dff_B_F0P9hycQ6_2(.din(w_dff_B_qS3xw9qH4_2),.dout(w_dff_B_F0P9hycQ6_2),.clk(gclk));
	jdff dff_B_EckjCATr2_2(.din(w_dff_B_F0P9hycQ6_2),.dout(w_dff_B_EckjCATr2_2),.clk(gclk));
	jdff dff_B_hfhgTPjF1_2(.din(w_dff_B_EckjCATr2_2),.dout(w_dff_B_hfhgTPjF1_2),.clk(gclk));
	jdff dff_B_dk3gJiMF1_2(.din(w_dff_B_hfhgTPjF1_2),.dout(w_dff_B_dk3gJiMF1_2),.clk(gclk));
	jdff dff_B_VQJ4USoi2_2(.din(w_dff_B_dk3gJiMF1_2),.dout(w_dff_B_VQJ4USoi2_2),.clk(gclk));
	jdff dff_B_sbq09ePv9_2(.din(w_dff_B_VQJ4USoi2_2),.dout(w_dff_B_sbq09ePv9_2),.clk(gclk));
	jdff dff_B_8ET0SBc69_2(.din(w_dff_B_sbq09ePv9_2),.dout(w_dff_B_8ET0SBc69_2),.clk(gclk));
	jdff dff_B_8MgNKCBv6_2(.din(w_dff_B_8ET0SBc69_2),.dout(w_dff_B_8MgNKCBv6_2),.clk(gclk));
	jdff dff_B_K0KcBQaj9_2(.din(w_dff_B_8MgNKCBv6_2),.dout(w_dff_B_K0KcBQaj9_2),.clk(gclk));
	jdff dff_B_A8WpoR518_2(.din(w_dff_B_K0KcBQaj9_2),.dout(w_dff_B_A8WpoR518_2),.clk(gclk));
	jdff dff_B_S3MWRViv5_2(.din(w_dff_B_A8WpoR518_2),.dout(w_dff_B_S3MWRViv5_2),.clk(gclk));
	jdff dff_B_6woJ4yq17_2(.din(w_dff_B_S3MWRViv5_2),.dout(w_dff_B_6woJ4yq17_2),.clk(gclk));
	jdff dff_B_gWBK3IYt8_2(.din(w_dff_B_6woJ4yq17_2),.dout(w_dff_B_gWBK3IYt8_2),.clk(gclk));
	jdff dff_B_EW08QSUF0_2(.din(w_dff_B_gWBK3IYt8_2),.dout(w_dff_B_EW08QSUF0_2),.clk(gclk));
	jdff dff_B_HA4Rymwa9_2(.din(w_dff_B_EW08QSUF0_2),.dout(w_dff_B_HA4Rymwa9_2),.clk(gclk));
	jdff dff_B_mYgJh4cX7_2(.din(w_dff_B_HA4Rymwa9_2),.dout(w_dff_B_mYgJh4cX7_2),.clk(gclk));
	jdff dff_B_LNvUpIxx0_2(.din(w_dff_B_mYgJh4cX7_2),.dout(w_dff_B_LNvUpIxx0_2),.clk(gclk));
	jdff dff_B_WJPC9az53_2(.din(w_dff_B_LNvUpIxx0_2),.dout(w_dff_B_WJPC9az53_2),.clk(gclk));
	jdff dff_B_EbO6FDzF9_2(.din(w_dff_B_WJPC9az53_2),.dout(w_dff_B_EbO6FDzF9_2),.clk(gclk));
	jdff dff_B_ArqXoQLF0_2(.din(n1413),.dout(w_dff_B_ArqXoQLF0_2),.clk(gclk));
	jdff dff_B_TLtisFvc9_1(.din(n1411),.dout(w_dff_B_TLtisFvc9_1),.clk(gclk));
	jdff dff_B_4DWvxcdV9_2(.din(n1332),.dout(w_dff_B_4DWvxcdV9_2),.clk(gclk));
	jdff dff_B_QDUfMgsb6_2(.din(w_dff_B_4DWvxcdV9_2),.dout(w_dff_B_QDUfMgsb6_2),.clk(gclk));
	jdff dff_B_I3cKe1RS8_2(.din(w_dff_B_QDUfMgsb6_2),.dout(w_dff_B_I3cKe1RS8_2),.clk(gclk));
	jdff dff_B_38Gw2lzi9_2(.din(w_dff_B_I3cKe1RS8_2),.dout(w_dff_B_38Gw2lzi9_2),.clk(gclk));
	jdff dff_B_iJMeS2Cm0_2(.din(w_dff_B_38Gw2lzi9_2),.dout(w_dff_B_iJMeS2Cm0_2),.clk(gclk));
	jdff dff_B_iakj3AJ72_2(.din(w_dff_B_iJMeS2Cm0_2),.dout(w_dff_B_iakj3AJ72_2),.clk(gclk));
	jdff dff_B_2MWgvuZD9_2(.din(w_dff_B_iakj3AJ72_2),.dout(w_dff_B_2MWgvuZD9_2),.clk(gclk));
	jdff dff_B_wsEJmLXr6_2(.din(w_dff_B_2MWgvuZD9_2),.dout(w_dff_B_wsEJmLXr6_2),.clk(gclk));
	jdff dff_B_qThltIpz6_2(.din(w_dff_B_wsEJmLXr6_2),.dout(w_dff_B_qThltIpz6_2),.clk(gclk));
	jdff dff_B_3CfE73JL3_2(.din(w_dff_B_qThltIpz6_2),.dout(w_dff_B_3CfE73JL3_2),.clk(gclk));
	jdff dff_B_prXifrhR7_2(.din(w_dff_B_3CfE73JL3_2),.dout(w_dff_B_prXifrhR7_2),.clk(gclk));
	jdff dff_B_TDt9EeZK8_2(.din(w_dff_B_prXifrhR7_2),.dout(w_dff_B_TDt9EeZK8_2),.clk(gclk));
	jdff dff_B_mt1TfKB29_2(.din(w_dff_B_TDt9EeZK8_2),.dout(w_dff_B_mt1TfKB29_2),.clk(gclk));
	jdff dff_B_zD6LTIp08_2(.din(w_dff_B_mt1TfKB29_2),.dout(w_dff_B_zD6LTIp08_2),.clk(gclk));
	jdff dff_B_iDgjAlzy6_2(.din(w_dff_B_zD6LTIp08_2),.dout(w_dff_B_iDgjAlzy6_2),.clk(gclk));
	jdff dff_B_EyqPd3UR0_2(.din(w_dff_B_iDgjAlzy6_2),.dout(w_dff_B_EyqPd3UR0_2),.clk(gclk));
	jdff dff_B_B8BD1BdN8_2(.din(w_dff_B_EyqPd3UR0_2),.dout(w_dff_B_B8BD1BdN8_2),.clk(gclk));
	jdff dff_B_IMsAsla93_2(.din(w_dff_B_B8BD1BdN8_2),.dout(w_dff_B_IMsAsla93_2),.clk(gclk));
	jdff dff_B_MDHoOfON6_2(.din(w_dff_B_IMsAsla93_2),.dout(w_dff_B_MDHoOfON6_2),.clk(gclk));
	jdff dff_B_4N6NNVcz9_2(.din(w_dff_B_MDHoOfON6_2),.dout(w_dff_B_4N6NNVcz9_2),.clk(gclk));
	jdff dff_B_OsPByg8L9_2(.din(w_dff_B_4N6NNVcz9_2),.dout(w_dff_B_OsPByg8L9_2),.clk(gclk));
	jdff dff_B_x2InN0J80_2(.din(w_dff_B_OsPByg8L9_2),.dout(w_dff_B_x2InN0J80_2),.clk(gclk));
	jdff dff_B_SblAxLOd8_1(.din(n1333),.dout(w_dff_B_SblAxLOd8_1),.clk(gclk));
	jdff dff_B_OJ4JnQJB2_2(.din(n1247),.dout(w_dff_B_OJ4JnQJB2_2),.clk(gclk));
	jdff dff_B_wCXotfUE3_2(.din(w_dff_B_OJ4JnQJB2_2),.dout(w_dff_B_wCXotfUE3_2),.clk(gclk));
	jdff dff_B_Ra8iuUCc6_2(.din(w_dff_B_wCXotfUE3_2),.dout(w_dff_B_Ra8iuUCc6_2),.clk(gclk));
	jdff dff_B_yeuLYKfg3_2(.din(w_dff_B_Ra8iuUCc6_2),.dout(w_dff_B_yeuLYKfg3_2),.clk(gclk));
	jdff dff_B_Rq33UQ3B7_2(.din(w_dff_B_yeuLYKfg3_2),.dout(w_dff_B_Rq33UQ3B7_2),.clk(gclk));
	jdff dff_B_uSeNHYCW1_2(.din(w_dff_B_Rq33UQ3B7_2),.dout(w_dff_B_uSeNHYCW1_2),.clk(gclk));
	jdff dff_B_w3PZDCol5_2(.din(w_dff_B_uSeNHYCW1_2),.dout(w_dff_B_w3PZDCol5_2),.clk(gclk));
	jdff dff_B_5kWWp7NJ8_2(.din(w_dff_B_w3PZDCol5_2),.dout(w_dff_B_5kWWp7NJ8_2),.clk(gclk));
	jdff dff_B_UwMDgdMW3_2(.din(w_dff_B_5kWWp7NJ8_2),.dout(w_dff_B_UwMDgdMW3_2),.clk(gclk));
	jdff dff_B_qnTPUbn78_2(.din(w_dff_B_UwMDgdMW3_2),.dout(w_dff_B_qnTPUbn78_2),.clk(gclk));
	jdff dff_B_6zyzZOQC8_2(.din(w_dff_B_qnTPUbn78_2),.dout(w_dff_B_6zyzZOQC8_2),.clk(gclk));
	jdff dff_B_PgSGs52k4_2(.din(w_dff_B_6zyzZOQC8_2),.dout(w_dff_B_PgSGs52k4_2),.clk(gclk));
	jdff dff_B_eHskGCaK9_2(.din(w_dff_B_PgSGs52k4_2),.dout(w_dff_B_eHskGCaK9_2),.clk(gclk));
	jdff dff_B_go5r6peb2_2(.din(w_dff_B_eHskGCaK9_2),.dout(w_dff_B_go5r6peb2_2),.clk(gclk));
	jdff dff_B_OVpk8ql00_2(.din(w_dff_B_go5r6peb2_2),.dout(w_dff_B_OVpk8ql00_2),.clk(gclk));
	jdff dff_B_me1KJaCE9_2(.din(w_dff_B_OVpk8ql00_2),.dout(w_dff_B_me1KJaCE9_2),.clk(gclk));
	jdff dff_B_kJkRFspF4_2(.din(w_dff_B_me1KJaCE9_2),.dout(w_dff_B_kJkRFspF4_2),.clk(gclk));
	jdff dff_B_fs2yL4LS9_2(.din(w_dff_B_kJkRFspF4_2),.dout(w_dff_B_fs2yL4LS9_2),.clk(gclk));
	jdff dff_B_9CMwoNsU4_2(.din(w_dff_B_fs2yL4LS9_2),.dout(w_dff_B_9CMwoNsU4_2),.clk(gclk));
	jdff dff_B_xdbSe9VM5_2(.din(w_dff_B_9CMwoNsU4_2),.dout(w_dff_B_xdbSe9VM5_2),.clk(gclk));
	jdff dff_B_Q47A3wZg4_1(.din(n1248),.dout(w_dff_B_Q47A3wZg4_1),.clk(gclk));
	jdff dff_B_sUti06fg7_2(.din(n1156),.dout(w_dff_B_sUti06fg7_2),.clk(gclk));
	jdff dff_B_ZX0Jhod58_2(.din(w_dff_B_sUti06fg7_2),.dout(w_dff_B_ZX0Jhod58_2),.clk(gclk));
	jdff dff_B_DqVoTc2B6_2(.din(w_dff_B_ZX0Jhod58_2),.dout(w_dff_B_DqVoTc2B6_2),.clk(gclk));
	jdff dff_B_dLuNtJd85_2(.din(w_dff_B_DqVoTc2B6_2),.dout(w_dff_B_dLuNtJd85_2),.clk(gclk));
	jdff dff_B_rlsgxYi46_2(.din(w_dff_B_dLuNtJd85_2),.dout(w_dff_B_rlsgxYi46_2),.clk(gclk));
	jdff dff_B_KUgsDlTU6_2(.din(w_dff_B_rlsgxYi46_2),.dout(w_dff_B_KUgsDlTU6_2),.clk(gclk));
	jdff dff_B_RMENxy5T9_2(.din(w_dff_B_KUgsDlTU6_2),.dout(w_dff_B_RMENxy5T9_2),.clk(gclk));
	jdff dff_B_EOoiShaq7_2(.din(w_dff_B_RMENxy5T9_2),.dout(w_dff_B_EOoiShaq7_2),.clk(gclk));
	jdff dff_B_hLGC8ap34_2(.din(w_dff_B_EOoiShaq7_2),.dout(w_dff_B_hLGC8ap34_2),.clk(gclk));
	jdff dff_B_B3K2sMmk2_2(.din(w_dff_B_hLGC8ap34_2),.dout(w_dff_B_B3K2sMmk2_2),.clk(gclk));
	jdff dff_B_4LOcEv8e6_2(.din(w_dff_B_B3K2sMmk2_2),.dout(w_dff_B_4LOcEv8e6_2),.clk(gclk));
	jdff dff_B_RLG0ZDh45_2(.din(w_dff_B_4LOcEv8e6_2),.dout(w_dff_B_RLG0ZDh45_2),.clk(gclk));
	jdff dff_B_SWs2x6MT2_2(.din(w_dff_B_RLG0ZDh45_2),.dout(w_dff_B_SWs2x6MT2_2),.clk(gclk));
	jdff dff_B_BscJFiJj4_2(.din(w_dff_B_SWs2x6MT2_2),.dout(w_dff_B_BscJFiJj4_2),.clk(gclk));
	jdff dff_B_69Bbgfkw4_2(.din(w_dff_B_BscJFiJj4_2),.dout(w_dff_B_69Bbgfkw4_2),.clk(gclk));
	jdff dff_B_SkcNSFnk3_2(.din(w_dff_B_69Bbgfkw4_2),.dout(w_dff_B_SkcNSFnk3_2),.clk(gclk));
	jdff dff_B_5n1qQk7e4_2(.din(w_dff_B_SkcNSFnk3_2),.dout(w_dff_B_5n1qQk7e4_2),.clk(gclk));
	jdff dff_B_aPtSe8m90_2(.din(w_dff_B_5n1qQk7e4_2),.dout(w_dff_B_aPtSe8m90_2),.clk(gclk));
	jdff dff_B_QsGqq5Sx7_1(.din(n1157),.dout(w_dff_B_QsGqq5Sx7_1),.clk(gclk));
	jdff dff_B_LA0y961X7_2(.din(n1058),.dout(w_dff_B_LA0y961X7_2),.clk(gclk));
	jdff dff_B_inGyD92K1_2(.din(w_dff_B_LA0y961X7_2),.dout(w_dff_B_inGyD92K1_2),.clk(gclk));
	jdff dff_B_Gis1xd6E8_2(.din(w_dff_B_inGyD92K1_2),.dout(w_dff_B_Gis1xd6E8_2),.clk(gclk));
	jdff dff_B_GepeqIs48_2(.din(w_dff_B_Gis1xd6E8_2),.dout(w_dff_B_GepeqIs48_2),.clk(gclk));
	jdff dff_B_IkVdo9Kj0_2(.din(w_dff_B_GepeqIs48_2),.dout(w_dff_B_IkVdo9Kj0_2),.clk(gclk));
	jdff dff_B_bRMPDL0D9_2(.din(w_dff_B_IkVdo9Kj0_2),.dout(w_dff_B_bRMPDL0D9_2),.clk(gclk));
	jdff dff_B_e6JN9olU6_2(.din(w_dff_B_bRMPDL0D9_2),.dout(w_dff_B_e6JN9olU6_2),.clk(gclk));
	jdff dff_B_ejxohMYf3_2(.din(w_dff_B_e6JN9olU6_2),.dout(w_dff_B_ejxohMYf3_2),.clk(gclk));
	jdff dff_B_5eMe5wWo5_2(.din(w_dff_B_ejxohMYf3_2),.dout(w_dff_B_5eMe5wWo5_2),.clk(gclk));
	jdff dff_B_nHBUiJmd1_2(.din(w_dff_B_5eMe5wWo5_2),.dout(w_dff_B_nHBUiJmd1_2),.clk(gclk));
	jdff dff_B_tDydL1PX0_2(.din(w_dff_B_nHBUiJmd1_2),.dout(w_dff_B_tDydL1PX0_2),.clk(gclk));
	jdff dff_B_eliUbxDp7_2(.din(w_dff_B_tDydL1PX0_2),.dout(w_dff_B_eliUbxDp7_2),.clk(gclk));
	jdff dff_B_AZZw5Ixz4_2(.din(w_dff_B_eliUbxDp7_2),.dout(w_dff_B_AZZw5Ixz4_2),.clk(gclk));
	jdff dff_B_198TQkrY6_2(.din(w_dff_B_AZZw5Ixz4_2),.dout(w_dff_B_198TQkrY6_2),.clk(gclk));
	jdff dff_B_ukWplGiy0_2(.din(w_dff_B_198TQkrY6_2),.dout(w_dff_B_ukWplGiy0_2),.clk(gclk));
	jdff dff_B_ZFYsJInP3_2(.din(w_dff_B_ukWplGiy0_2),.dout(w_dff_B_ZFYsJInP3_2),.clk(gclk));
	jdff dff_B_DrhxwjcS0_1(.din(n1059),.dout(w_dff_B_DrhxwjcS0_1),.clk(gclk));
	jdff dff_B_xwJhvg0Q4_2(.din(n959),.dout(w_dff_B_xwJhvg0Q4_2),.clk(gclk));
	jdff dff_B_YRwg5mzY8_2(.din(w_dff_B_xwJhvg0Q4_2),.dout(w_dff_B_YRwg5mzY8_2),.clk(gclk));
	jdff dff_B_epcv4njW1_2(.din(w_dff_B_YRwg5mzY8_2),.dout(w_dff_B_epcv4njW1_2),.clk(gclk));
	jdff dff_B_UeM2oomk1_2(.din(w_dff_B_epcv4njW1_2),.dout(w_dff_B_UeM2oomk1_2),.clk(gclk));
	jdff dff_B_0AoTfTuT7_2(.din(w_dff_B_UeM2oomk1_2),.dout(w_dff_B_0AoTfTuT7_2),.clk(gclk));
	jdff dff_B_19FKgTfh7_2(.din(w_dff_B_0AoTfTuT7_2),.dout(w_dff_B_19FKgTfh7_2),.clk(gclk));
	jdff dff_B_fOUEpAxL8_2(.din(w_dff_B_19FKgTfh7_2),.dout(w_dff_B_fOUEpAxL8_2),.clk(gclk));
	jdff dff_B_otOH1XqV2_2(.din(w_dff_B_fOUEpAxL8_2),.dout(w_dff_B_otOH1XqV2_2),.clk(gclk));
	jdff dff_B_3lFqYNwn7_2(.din(w_dff_B_otOH1XqV2_2),.dout(w_dff_B_3lFqYNwn7_2),.clk(gclk));
	jdff dff_B_QxsNpPkw7_2(.din(w_dff_B_3lFqYNwn7_2),.dout(w_dff_B_QxsNpPkw7_2),.clk(gclk));
	jdff dff_B_RAyjpQdF9_2(.din(w_dff_B_QxsNpPkw7_2),.dout(w_dff_B_RAyjpQdF9_2),.clk(gclk));
	jdff dff_B_92SXSXjX8_2(.din(w_dff_B_RAyjpQdF9_2),.dout(w_dff_B_92SXSXjX8_2),.clk(gclk));
	jdff dff_B_cito59mb9_2(.din(w_dff_B_92SXSXjX8_2),.dout(w_dff_B_cito59mb9_2),.clk(gclk));
	jdff dff_B_EVtxD5999_2(.din(w_dff_B_cito59mb9_2),.dout(w_dff_B_EVtxD5999_2),.clk(gclk));
	jdff dff_B_bYy1OwRT1_1(.din(n960),.dout(w_dff_B_bYy1OwRT1_1),.clk(gclk));
	jdff dff_B_kUHza9uG2_2(.din(n857),.dout(w_dff_B_kUHza9uG2_2),.clk(gclk));
	jdff dff_B_bhwEK5bt2_2(.din(w_dff_B_kUHza9uG2_2),.dout(w_dff_B_bhwEK5bt2_2),.clk(gclk));
	jdff dff_B_xEUE7uo23_2(.din(w_dff_B_bhwEK5bt2_2),.dout(w_dff_B_xEUE7uo23_2),.clk(gclk));
	jdff dff_B_tSU0Z8BE5_2(.din(w_dff_B_xEUE7uo23_2),.dout(w_dff_B_tSU0Z8BE5_2),.clk(gclk));
	jdff dff_B_ts9UJt7J1_2(.din(w_dff_B_tSU0Z8BE5_2),.dout(w_dff_B_ts9UJt7J1_2),.clk(gclk));
	jdff dff_B_FFpo0OqE6_2(.din(w_dff_B_ts9UJt7J1_2),.dout(w_dff_B_FFpo0OqE6_2),.clk(gclk));
	jdff dff_B_898eVje57_2(.din(w_dff_B_FFpo0OqE6_2),.dout(w_dff_B_898eVje57_2),.clk(gclk));
	jdff dff_B_wCegv5yY3_2(.din(w_dff_B_898eVje57_2),.dout(w_dff_B_wCegv5yY3_2),.clk(gclk));
	jdff dff_B_s3clsBNy0_2(.din(w_dff_B_wCegv5yY3_2),.dout(w_dff_B_s3clsBNy0_2),.clk(gclk));
	jdff dff_B_P1tqOhQ32_2(.din(w_dff_B_s3clsBNy0_2),.dout(w_dff_B_P1tqOhQ32_2),.clk(gclk));
	jdff dff_B_R4lCshcJ5_2(.din(w_dff_B_P1tqOhQ32_2),.dout(w_dff_B_R4lCshcJ5_2),.clk(gclk));
	jdff dff_B_Jii61y7X1_2(.din(w_dff_B_R4lCshcJ5_2),.dout(w_dff_B_Jii61y7X1_2),.clk(gclk));
	jdff dff_B_0ZsMoynN4_1(.din(n858),.dout(w_dff_B_0ZsMoynN4_1),.clk(gclk));
	jdff dff_B_J08wHF7i5_2(.din(n759),.dout(w_dff_B_J08wHF7i5_2),.clk(gclk));
	jdff dff_B_wTmm9n9Z9_2(.din(w_dff_B_J08wHF7i5_2),.dout(w_dff_B_wTmm9n9Z9_2),.clk(gclk));
	jdff dff_B_fUYcGxKE9_2(.din(w_dff_B_wTmm9n9Z9_2),.dout(w_dff_B_fUYcGxKE9_2),.clk(gclk));
	jdff dff_B_cjdPkUFn9_2(.din(w_dff_B_fUYcGxKE9_2),.dout(w_dff_B_cjdPkUFn9_2),.clk(gclk));
	jdff dff_B_2EEc9zb23_2(.din(w_dff_B_cjdPkUFn9_2),.dout(w_dff_B_2EEc9zb23_2),.clk(gclk));
	jdff dff_B_r0OWAUOU4_2(.din(w_dff_B_2EEc9zb23_2),.dout(w_dff_B_r0OWAUOU4_2),.clk(gclk));
	jdff dff_B_yG45ZPEJ0_2(.din(w_dff_B_r0OWAUOU4_2),.dout(w_dff_B_yG45ZPEJ0_2),.clk(gclk));
	jdff dff_B_mU0vltQ72_2(.din(w_dff_B_yG45ZPEJ0_2),.dout(w_dff_B_mU0vltQ72_2),.clk(gclk));
	jdff dff_B_NbvEfiLT5_2(.din(w_dff_B_mU0vltQ72_2),.dout(w_dff_B_NbvEfiLT5_2),.clk(gclk));
	jdff dff_B_QriFem3S1_2(.din(w_dff_B_NbvEfiLT5_2),.dout(w_dff_B_QriFem3S1_2),.clk(gclk));
	jdff dff_B_cgMAQ9Lj0_1(.din(n760),.dout(w_dff_B_cgMAQ9Lj0_1),.clk(gclk));
	jdff dff_B_IihquM6n1_2(.din(n667),.dout(w_dff_B_IihquM6n1_2),.clk(gclk));
	jdff dff_B_r08S5zql6_2(.din(w_dff_B_IihquM6n1_2),.dout(w_dff_B_r08S5zql6_2),.clk(gclk));
	jdff dff_B_AOOHxe6x2_2(.din(w_dff_B_r08S5zql6_2),.dout(w_dff_B_AOOHxe6x2_2),.clk(gclk));
	jdff dff_B_jbniQ65W6_2(.din(w_dff_B_AOOHxe6x2_2),.dout(w_dff_B_jbniQ65W6_2),.clk(gclk));
	jdff dff_B_6bcp0QCv6_2(.din(w_dff_B_jbniQ65W6_2),.dout(w_dff_B_6bcp0QCv6_2),.clk(gclk));
	jdff dff_B_HMIz3pOd5_2(.din(w_dff_B_6bcp0QCv6_2),.dout(w_dff_B_HMIz3pOd5_2),.clk(gclk));
	jdff dff_B_nNQVii0L1_2(.din(w_dff_B_HMIz3pOd5_2),.dout(w_dff_B_nNQVii0L1_2),.clk(gclk));
	jdff dff_B_pfmOU5sT4_2(.din(w_dff_B_nNQVii0L1_2),.dout(w_dff_B_pfmOU5sT4_2),.clk(gclk));
	jdff dff_B_pJf4QxHE3_2(.din(n682),.dout(w_dff_B_pJf4QxHE3_2),.clk(gclk));
	jdff dff_B_rAK4d0JX2_2(.din(w_dff_B_pJf4QxHE3_2),.dout(w_dff_B_rAK4d0JX2_2),.clk(gclk));
	jdff dff_B_YIhjSKK65_2(.din(w_dff_B_rAK4d0JX2_2),.dout(w_dff_B_YIhjSKK65_2),.clk(gclk));
	jdff dff_B_rwjqd2Fm2_1(.din(n668),.dout(w_dff_B_rwjqd2Fm2_1),.clk(gclk));
	jdff dff_B_5cMpneYK2_1(.din(w_dff_B_rwjqd2Fm2_1),.dout(w_dff_B_5cMpneYK2_1),.clk(gclk));
	jdff dff_B_Rh8AN04i2_1(.din(w_dff_B_5cMpneYK2_1),.dout(w_dff_B_Rh8AN04i2_1),.clk(gclk));
	jdff dff_B_jkdrcr0D2_2(.din(n584),.dout(w_dff_B_jkdrcr0D2_2),.clk(gclk));
	jdff dff_B_xi23xvLP7_2(.din(w_dff_B_jkdrcr0D2_2),.dout(w_dff_B_xi23xvLP7_2),.clk(gclk));
	jdff dff_B_tLuPYHai7_2(.din(w_dff_B_xi23xvLP7_2),.dout(w_dff_B_tLuPYHai7_2),.clk(gclk));
	jdff dff_B_2FbvjWma8_0(.din(n589),.dout(w_dff_B_2FbvjWma8_0),.clk(gclk));
	jdff dff_B_Xk0MFmbp8_0(.din(w_dff_B_2FbvjWma8_0),.dout(w_dff_B_Xk0MFmbp8_0),.clk(gclk));
	jdff dff_A_T2KRF8Fd3_0(.dout(w_n503_0[0]),.din(w_dff_A_T2KRF8Fd3_0),.clk(gclk));
	jdff dff_A_rrIgy5qa0_0(.dout(w_dff_A_T2KRF8Fd3_0),.din(w_dff_A_rrIgy5qa0_0),.clk(gclk));
	jdff dff_A_SeewxzKt8_1(.dout(w_n503_0[1]),.din(w_dff_A_SeewxzKt8_1),.clk(gclk));
	jdff dff_A_DK2WnL0g7_1(.dout(w_dff_A_SeewxzKt8_1),.din(w_dff_A_DK2WnL0g7_1),.clk(gclk));
	jdff dff_B_s9URHH6X8_1(.din(n1762),.dout(w_dff_B_s9URHH6X8_1),.clk(gclk));
	jdff dff_A_3cdlYTgW1_1(.dout(w_n1737_0[1]),.din(w_dff_A_3cdlYTgW1_1),.clk(gclk));
	jdff dff_B_zn1GqKHr3_1(.din(n1735),.dout(w_dff_B_zn1GqKHr3_1),.clk(gclk));
	jdff dff_B_JQvsXwFq0_2(.din(n1699),.dout(w_dff_B_JQvsXwFq0_2),.clk(gclk));
	jdff dff_B_URcEVwNy0_2(.din(w_dff_B_JQvsXwFq0_2),.dout(w_dff_B_URcEVwNy0_2),.clk(gclk));
	jdff dff_B_OgpRmJbk3_2(.din(w_dff_B_URcEVwNy0_2),.dout(w_dff_B_OgpRmJbk3_2),.clk(gclk));
	jdff dff_B_ziyCwVRs9_2(.din(w_dff_B_OgpRmJbk3_2),.dout(w_dff_B_ziyCwVRs9_2),.clk(gclk));
	jdff dff_B_wJ6XdJH00_2(.din(w_dff_B_ziyCwVRs9_2),.dout(w_dff_B_wJ6XdJH00_2),.clk(gclk));
	jdff dff_B_S57zhDqo1_2(.din(w_dff_B_wJ6XdJH00_2),.dout(w_dff_B_S57zhDqo1_2),.clk(gclk));
	jdff dff_B_hYEZKbac0_2(.din(w_dff_B_S57zhDqo1_2),.dout(w_dff_B_hYEZKbac0_2),.clk(gclk));
	jdff dff_B_jy0fDjNG8_2(.din(w_dff_B_hYEZKbac0_2),.dout(w_dff_B_jy0fDjNG8_2),.clk(gclk));
	jdff dff_B_lLQpOBoG7_2(.din(w_dff_B_jy0fDjNG8_2),.dout(w_dff_B_lLQpOBoG7_2),.clk(gclk));
	jdff dff_B_SQdAL7z73_2(.din(w_dff_B_lLQpOBoG7_2),.dout(w_dff_B_SQdAL7z73_2),.clk(gclk));
	jdff dff_B_9rilH1Ps7_2(.din(w_dff_B_SQdAL7z73_2),.dout(w_dff_B_9rilH1Ps7_2),.clk(gclk));
	jdff dff_B_ZiIHuY8R6_2(.din(w_dff_B_9rilH1Ps7_2),.dout(w_dff_B_ZiIHuY8R6_2),.clk(gclk));
	jdff dff_B_m4H2Zib90_2(.din(w_dff_B_ZiIHuY8R6_2),.dout(w_dff_B_m4H2Zib90_2),.clk(gclk));
	jdff dff_B_1Of8N5Iu2_2(.din(w_dff_B_m4H2Zib90_2),.dout(w_dff_B_1Of8N5Iu2_2),.clk(gclk));
	jdff dff_B_REQtgeSP1_2(.din(w_dff_B_1Of8N5Iu2_2),.dout(w_dff_B_REQtgeSP1_2),.clk(gclk));
	jdff dff_B_LdXGDG7H5_2(.din(w_dff_B_REQtgeSP1_2),.dout(w_dff_B_LdXGDG7H5_2),.clk(gclk));
	jdff dff_B_gFRCuXn28_2(.din(w_dff_B_LdXGDG7H5_2),.dout(w_dff_B_gFRCuXn28_2),.clk(gclk));
	jdff dff_B_CMUmo4SJ6_2(.din(w_dff_B_gFRCuXn28_2),.dout(w_dff_B_CMUmo4SJ6_2),.clk(gclk));
	jdff dff_B_te1iNZRa8_2(.din(w_dff_B_CMUmo4SJ6_2),.dout(w_dff_B_te1iNZRa8_2),.clk(gclk));
	jdff dff_B_WU3W2Kx24_2(.din(w_dff_B_te1iNZRa8_2),.dout(w_dff_B_WU3W2Kx24_2),.clk(gclk));
	jdff dff_B_LOHVeOO25_2(.din(w_dff_B_WU3W2Kx24_2),.dout(w_dff_B_LOHVeOO25_2),.clk(gclk));
	jdff dff_B_BPSUXMde2_2(.din(w_dff_B_LOHVeOO25_2),.dout(w_dff_B_BPSUXMde2_2),.clk(gclk));
	jdff dff_B_v4hfpko45_2(.din(w_dff_B_BPSUXMde2_2),.dout(w_dff_B_v4hfpko45_2),.clk(gclk));
	jdff dff_B_jsJhMGRl9_2(.din(w_dff_B_v4hfpko45_2),.dout(w_dff_B_jsJhMGRl9_2),.clk(gclk));
	jdff dff_B_pziGGJK40_2(.din(w_dff_B_jsJhMGRl9_2),.dout(w_dff_B_pziGGJK40_2),.clk(gclk));
	jdff dff_B_QFckyIIg6_2(.din(w_dff_B_pziGGJK40_2),.dout(w_dff_B_QFckyIIg6_2),.clk(gclk));
	jdff dff_B_kvjlVmal4_2(.din(w_dff_B_QFckyIIg6_2),.dout(w_dff_B_kvjlVmal4_2),.clk(gclk));
	jdff dff_B_RWGR07XR3_2(.din(w_dff_B_kvjlVmal4_2),.dout(w_dff_B_RWGR07XR3_2),.clk(gclk));
	jdff dff_B_ouzKxJNe2_2(.din(w_dff_B_RWGR07XR3_2),.dout(w_dff_B_ouzKxJNe2_2),.clk(gclk));
	jdff dff_B_MC8JN1nJ8_2(.din(w_dff_B_ouzKxJNe2_2),.dout(w_dff_B_MC8JN1nJ8_2),.clk(gclk));
	jdff dff_B_4MJdl2Ka2_2(.din(w_dff_B_MC8JN1nJ8_2),.dout(w_dff_B_4MJdl2Ka2_2),.clk(gclk));
	jdff dff_B_nR8Mq71c3_2(.din(w_dff_B_4MJdl2Ka2_2),.dout(w_dff_B_nR8Mq71c3_2),.clk(gclk));
	jdff dff_B_txStUAdM9_2(.din(w_dff_B_nR8Mq71c3_2),.dout(w_dff_B_txStUAdM9_2),.clk(gclk));
	jdff dff_B_lecib16x5_2(.din(w_dff_B_txStUAdM9_2),.dout(w_dff_B_lecib16x5_2),.clk(gclk));
	jdff dff_B_6s6jQdzQ4_2(.din(w_dff_B_lecib16x5_2),.dout(w_dff_B_6s6jQdzQ4_2),.clk(gclk));
	jdff dff_B_lOrHr0yL6_2(.din(w_dff_B_6s6jQdzQ4_2),.dout(w_dff_B_lOrHr0yL6_2),.clk(gclk));
	jdff dff_B_albXu4Yb6_2(.din(w_dff_B_lOrHr0yL6_2),.dout(w_dff_B_albXu4Yb6_2),.clk(gclk));
	jdff dff_B_rpETgB5D8_2(.din(w_dff_B_albXu4Yb6_2),.dout(w_dff_B_rpETgB5D8_2),.clk(gclk));
	jdff dff_B_8F3sj5hl8_2(.din(n1702),.dout(w_dff_B_8F3sj5hl8_2),.clk(gclk));
	jdff dff_B_bWhd0JRq4_1(.din(n1700),.dout(w_dff_B_bWhd0JRq4_1),.clk(gclk));
	jdff dff_B_NceV2XFZ2_2(.din(n1658),.dout(w_dff_B_NceV2XFZ2_2),.clk(gclk));
	jdff dff_B_78kZyxZz5_2(.din(w_dff_B_NceV2XFZ2_2),.dout(w_dff_B_78kZyxZz5_2),.clk(gclk));
	jdff dff_B_eeeQodBV5_2(.din(w_dff_B_78kZyxZz5_2),.dout(w_dff_B_eeeQodBV5_2),.clk(gclk));
	jdff dff_B_WckFnbQ17_2(.din(w_dff_B_eeeQodBV5_2),.dout(w_dff_B_WckFnbQ17_2),.clk(gclk));
	jdff dff_B_Y60aYXNH9_2(.din(w_dff_B_WckFnbQ17_2),.dout(w_dff_B_Y60aYXNH9_2),.clk(gclk));
	jdff dff_B_F7flt7i61_2(.din(w_dff_B_Y60aYXNH9_2),.dout(w_dff_B_F7flt7i61_2),.clk(gclk));
	jdff dff_B_aPHQpUby1_2(.din(w_dff_B_F7flt7i61_2),.dout(w_dff_B_aPHQpUby1_2),.clk(gclk));
	jdff dff_B_5VgjWmd19_2(.din(w_dff_B_aPHQpUby1_2),.dout(w_dff_B_5VgjWmd19_2),.clk(gclk));
	jdff dff_B_UT0ULpdG5_2(.din(w_dff_B_5VgjWmd19_2),.dout(w_dff_B_UT0ULpdG5_2),.clk(gclk));
	jdff dff_B_kdmJv8NN6_2(.din(w_dff_B_UT0ULpdG5_2),.dout(w_dff_B_kdmJv8NN6_2),.clk(gclk));
	jdff dff_B_y4ilG7I21_2(.din(w_dff_B_kdmJv8NN6_2),.dout(w_dff_B_y4ilG7I21_2),.clk(gclk));
	jdff dff_B_6IOdWjSI4_2(.din(w_dff_B_y4ilG7I21_2),.dout(w_dff_B_6IOdWjSI4_2),.clk(gclk));
	jdff dff_B_XYk7SIV42_2(.din(w_dff_B_6IOdWjSI4_2),.dout(w_dff_B_XYk7SIV42_2),.clk(gclk));
	jdff dff_B_19xxkGM35_2(.din(w_dff_B_XYk7SIV42_2),.dout(w_dff_B_19xxkGM35_2),.clk(gclk));
	jdff dff_B_qrrEeIxw5_2(.din(w_dff_B_19xxkGM35_2),.dout(w_dff_B_qrrEeIxw5_2),.clk(gclk));
	jdff dff_B_CgIY4SJD4_2(.din(w_dff_B_qrrEeIxw5_2),.dout(w_dff_B_CgIY4SJD4_2),.clk(gclk));
	jdff dff_B_fGn2kFiJ4_2(.din(w_dff_B_CgIY4SJD4_2),.dout(w_dff_B_fGn2kFiJ4_2),.clk(gclk));
	jdff dff_B_PaB9nUod8_2(.din(w_dff_B_fGn2kFiJ4_2),.dout(w_dff_B_PaB9nUod8_2),.clk(gclk));
	jdff dff_B_NeTfnmOb4_2(.din(w_dff_B_PaB9nUod8_2),.dout(w_dff_B_NeTfnmOb4_2),.clk(gclk));
	jdff dff_B_X4so6oJu2_2(.din(w_dff_B_NeTfnmOb4_2),.dout(w_dff_B_X4so6oJu2_2),.clk(gclk));
	jdff dff_B_TqlBYD1S1_2(.din(w_dff_B_X4so6oJu2_2),.dout(w_dff_B_TqlBYD1S1_2),.clk(gclk));
	jdff dff_B_oyyBpjv97_2(.din(w_dff_B_TqlBYD1S1_2),.dout(w_dff_B_oyyBpjv97_2),.clk(gclk));
	jdff dff_B_tus45UP17_2(.din(w_dff_B_oyyBpjv97_2),.dout(w_dff_B_tus45UP17_2),.clk(gclk));
	jdff dff_B_MWNGRxcD5_2(.din(w_dff_B_tus45UP17_2),.dout(w_dff_B_MWNGRxcD5_2),.clk(gclk));
	jdff dff_B_gKDuqa6h5_2(.din(w_dff_B_MWNGRxcD5_2),.dout(w_dff_B_gKDuqa6h5_2),.clk(gclk));
	jdff dff_B_KECTLfSI4_2(.din(w_dff_B_gKDuqa6h5_2),.dout(w_dff_B_KECTLfSI4_2),.clk(gclk));
	jdff dff_B_M3YeJXZi2_2(.din(w_dff_B_KECTLfSI4_2),.dout(w_dff_B_M3YeJXZi2_2),.clk(gclk));
	jdff dff_B_lVdRQTMn1_2(.din(w_dff_B_M3YeJXZi2_2),.dout(w_dff_B_lVdRQTMn1_2),.clk(gclk));
	jdff dff_B_N59cVE4J0_2(.din(w_dff_B_lVdRQTMn1_2),.dout(w_dff_B_N59cVE4J0_2),.clk(gclk));
	jdff dff_B_cFjkWjwF7_2(.din(w_dff_B_N59cVE4J0_2),.dout(w_dff_B_cFjkWjwF7_2),.clk(gclk));
	jdff dff_B_jyqf18H51_2(.din(w_dff_B_cFjkWjwF7_2),.dout(w_dff_B_jyqf18H51_2),.clk(gclk));
	jdff dff_B_Enhwv3RE0_2(.din(w_dff_B_jyqf18H51_2),.dout(w_dff_B_Enhwv3RE0_2),.clk(gclk));
	jdff dff_B_25s2XIJY6_2(.din(w_dff_B_Enhwv3RE0_2),.dout(w_dff_B_25s2XIJY6_2),.clk(gclk));
	jdff dff_B_WDj3OuCc4_2(.din(w_dff_B_25s2XIJY6_2),.dout(w_dff_B_WDj3OuCc4_2),.clk(gclk));
	jdff dff_B_dAEQBR6J5_2(.din(w_dff_B_WDj3OuCc4_2),.dout(w_dff_B_dAEQBR6J5_2),.clk(gclk));
	jdff dff_B_b59aqmGd7_2(.din(n1661),.dout(w_dff_B_b59aqmGd7_2),.clk(gclk));
	jdff dff_B_8YAqrqWn5_1(.din(n1659),.dout(w_dff_B_8YAqrqWn5_1),.clk(gclk));
	jdff dff_B_z1FuxEoZ7_2(.din(n1607),.dout(w_dff_B_z1FuxEoZ7_2),.clk(gclk));
	jdff dff_B_2G83fqto0_2(.din(w_dff_B_z1FuxEoZ7_2),.dout(w_dff_B_2G83fqto0_2),.clk(gclk));
	jdff dff_B_Emp1WiSE6_2(.din(w_dff_B_2G83fqto0_2),.dout(w_dff_B_Emp1WiSE6_2),.clk(gclk));
	jdff dff_B_DUiRXHXm0_2(.din(w_dff_B_Emp1WiSE6_2),.dout(w_dff_B_DUiRXHXm0_2),.clk(gclk));
	jdff dff_B_rx6JoiWH9_2(.din(w_dff_B_DUiRXHXm0_2),.dout(w_dff_B_rx6JoiWH9_2),.clk(gclk));
	jdff dff_B_3P1mNYXI8_2(.din(w_dff_B_rx6JoiWH9_2),.dout(w_dff_B_3P1mNYXI8_2),.clk(gclk));
	jdff dff_B_0bmjbqKn5_2(.din(w_dff_B_3P1mNYXI8_2),.dout(w_dff_B_0bmjbqKn5_2),.clk(gclk));
	jdff dff_B_MPcX7RhJ4_2(.din(w_dff_B_0bmjbqKn5_2),.dout(w_dff_B_MPcX7RhJ4_2),.clk(gclk));
	jdff dff_B_dH1tXWpx3_2(.din(w_dff_B_MPcX7RhJ4_2),.dout(w_dff_B_dH1tXWpx3_2),.clk(gclk));
	jdff dff_B_QlCD84lh4_2(.din(w_dff_B_dH1tXWpx3_2),.dout(w_dff_B_QlCD84lh4_2),.clk(gclk));
	jdff dff_B_vSI0pBcb5_2(.din(w_dff_B_QlCD84lh4_2),.dout(w_dff_B_vSI0pBcb5_2),.clk(gclk));
	jdff dff_B_0rBU27UG1_2(.din(w_dff_B_vSI0pBcb5_2),.dout(w_dff_B_0rBU27UG1_2),.clk(gclk));
	jdff dff_B_WFE0MOd79_2(.din(w_dff_B_0rBU27UG1_2),.dout(w_dff_B_WFE0MOd79_2),.clk(gclk));
	jdff dff_B_YU2GDSQG5_2(.din(w_dff_B_WFE0MOd79_2),.dout(w_dff_B_YU2GDSQG5_2),.clk(gclk));
	jdff dff_B_COLJEkRH1_2(.din(w_dff_B_YU2GDSQG5_2),.dout(w_dff_B_COLJEkRH1_2),.clk(gclk));
	jdff dff_B_5H22GFfO1_2(.din(w_dff_B_COLJEkRH1_2),.dout(w_dff_B_5H22GFfO1_2),.clk(gclk));
	jdff dff_B_VRca994D1_2(.din(w_dff_B_5H22GFfO1_2),.dout(w_dff_B_VRca994D1_2),.clk(gclk));
	jdff dff_B_iBgBXIzs3_2(.din(w_dff_B_VRca994D1_2),.dout(w_dff_B_iBgBXIzs3_2),.clk(gclk));
	jdff dff_B_tQpIQ05D8_2(.din(w_dff_B_iBgBXIzs3_2),.dout(w_dff_B_tQpIQ05D8_2),.clk(gclk));
	jdff dff_B_7Lc2N3YZ2_2(.din(w_dff_B_tQpIQ05D8_2),.dout(w_dff_B_7Lc2N3YZ2_2),.clk(gclk));
	jdff dff_B_dw78O9DL3_2(.din(w_dff_B_7Lc2N3YZ2_2),.dout(w_dff_B_dw78O9DL3_2),.clk(gclk));
	jdff dff_B_zBLW9VIb7_2(.din(w_dff_B_dw78O9DL3_2),.dout(w_dff_B_zBLW9VIb7_2),.clk(gclk));
	jdff dff_B_tpwqCFhn0_2(.din(w_dff_B_zBLW9VIb7_2),.dout(w_dff_B_tpwqCFhn0_2),.clk(gclk));
	jdff dff_B_cbEmSlcb6_2(.din(w_dff_B_tpwqCFhn0_2),.dout(w_dff_B_cbEmSlcb6_2),.clk(gclk));
	jdff dff_B_qerQYLyU5_2(.din(w_dff_B_cbEmSlcb6_2),.dout(w_dff_B_qerQYLyU5_2),.clk(gclk));
	jdff dff_B_TxbnbpcG1_2(.din(w_dff_B_qerQYLyU5_2),.dout(w_dff_B_TxbnbpcG1_2),.clk(gclk));
	jdff dff_B_aAouONU28_2(.din(w_dff_B_TxbnbpcG1_2),.dout(w_dff_B_aAouONU28_2),.clk(gclk));
	jdff dff_B_ednQk6cC7_2(.din(w_dff_B_aAouONU28_2),.dout(w_dff_B_ednQk6cC7_2),.clk(gclk));
	jdff dff_B_wGC2Ykda3_2(.din(w_dff_B_ednQk6cC7_2),.dout(w_dff_B_wGC2Ykda3_2),.clk(gclk));
	jdff dff_B_f3tfPW3Y8_2(.din(w_dff_B_wGC2Ykda3_2),.dout(w_dff_B_f3tfPW3Y8_2),.clk(gclk));
	jdff dff_B_51TE2xvk5_2(.din(w_dff_B_f3tfPW3Y8_2),.dout(w_dff_B_51TE2xvk5_2),.clk(gclk));
	jdff dff_B_KzaSQKeX0_2(.din(w_dff_B_51TE2xvk5_2),.dout(w_dff_B_KzaSQKeX0_2),.clk(gclk));
	jdff dff_B_6C8Bv70R4_2(.din(n1610),.dout(w_dff_B_6C8Bv70R4_2),.clk(gclk));
	jdff dff_B_QUxCrnrP2_1(.din(n1608),.dout(w_dff_B_QUxCrnrP2_1),.clk(gclk));
	jdff dff_B_rP1iXW1r8_2(.din(n1550),.dout(w_dff_B_rP1iXW1r8_2),.clk(gclk));
	jdff dff_B_QnD1NCIy0_2(.din(w_dff_B_rP1iXW1r8_2),.dout(w_dff_B_QnD1NCIy0_2),.clk(gclk));
	jdff dff_B_lXZJx7kw6_2(.din(w_dff_B_QnD1NCIy0_2),.dout(w_dff_B_lXZJx7kw6_2),.clk(gclk));
	jdff dff_B_aegVVx8D7_2(.din(w_dff_B_lXZJx7kw6_2),.dout(w_dff_B_aegVVx8D7_2),.clk(gclk));
	jdff dff_B_v86uZsZu2_2(.din(w_dff_B_aegVVx8D7_2),.dout(w_dff_B_v86uZsZu2_2),.clk(gclk));
	jdff dff_B_vjD5kRak6_2(.din(w_dff_B_v86uZsZu2_2),.dout(w_dff_B_vjD5kRak6_2),.clk(gclk));
	jdff dff_B_YAw1nIPB6_2(.din(w_dff_B_vjD5kRak6_2),.dout(w_dff_B_YAw1nIPB6_2),.clk(gclk));
	jdff dff_B_toWiDd1w3_2(.din(w_dff_B_YAw1nIPB6_2),.dout(w_dff_B_toWiDd1w3_2),.clk(gclk));
	jdff dff_B_WLL8pHkl4_2(.din(w_dff_B_toWiDd1w3_2),.dout(w_dff_B_WLL8pHkl4_2),.clk(gclk));
	jdff dff_B_7mfRIqEx2_2(.din(w_dff_B_WLL8pHkl4_2),.dout(w_dff_B_7mfRIqEx2_2),.clk(gclk));
	jdff dff_B_fzD1B09G6_2(.din(w_dff_B_7mfRIqEx2_2),.dout(w_dff_B_fzD1B09G6_2),.clk(gclk));
	jdff dff_B_sbxtOkAn9_2(.din(w_dff_B_fzD1B09G6_2),.dout(w_dff_B_sbxtOkAn9_2),.clk(gclk));
	jdff dff_B_Z3WGGPwF1_2(.din(w_dff_B_sbxtOkAn9_2),.dout(w_dff_B_Z3WGGPwF1_2),.clk(gclk));
	jdff dff_B_1lJUoyFi6_2(.din(w_dff_B_Z3WGGPwF1_2),.dout(w_dff_B_1lJUoyFi6_2),.clk(gclk));
	jdff dff_B_LjAPldJH8_2(.din(w_dff_B_1lJUoyFi6_2),.dout(w_dff_B_LjAPldJH8_2),.clk(gclk));
	jdff dff_B_zuBMIn6I7_2(.din(w_dff_B_LjAPldJH8_2),.dout(w_dff_B_zuBMIn6I7_2),.clk(gclk));
	jdff dff_B_UliP24vG6_2(.din(w_dff_B_zuBMIn6I7_2),.dout(w_dff_B_UliP24vG6_2),.clk(gclk));
	jdff dff_B_38hELelm5_2(.din(w_dff_B_UliP24vG6_2),.dout(w_dff_B_38hELelm5_2),.clk(gclk));
	jdff dff_B_UaT7octZ7_2(.din(w_dff_B_38hELelm5_2),.dout(w_dff_B_UaT7octZ7_2),.clk(gclk));
	jdff dff_B_v7YKJnwO5_2(.din(w_dff_B_UaT7octZ7_2),.dout(w_dff_B_v7YKJnwO5_2),.clk(gclk));
	jdff dff_B_SqqV5f6z4_2(.din(w_dff_B_v7YKJnwO5_2),.dout(w_dff_B_SqqV5f6z4_2),.clk(gclk));
	jdff dff_B_yBm3HFis9_2(.din(w_dff_B_SqqV5f6z4_2),.dout(w_dff_B_yBm3HFis9_2),.clk(gclk));
	jdff dff_B_qmTAj92z3_2(.din(w_dff_B_yBm3HFis9_2),.dout(w_dff_B_qmTAj92z3_2),.clk(gclk));
	jdff dff_B_g7DhUzlX9_2(.din(w_dff_B_qmTAj92z3_2),.dout(w_dff_B_g7DhUzlX9_2),.clk(gclk));
	jdff dff_B_S3nUjeZH4_2(.din(w_dff_B_g7DhUzlX9_2),.dout(w_dff_B_S3nUjeZH4_2),.clk(gclk));
	jdff dff_B_m13h5eZ28_2(.din(w_dff_B_S3nUjeZH4_2),.dout(w_dff_B_m13h5eZ28_2),.clk(gclk));
	jdff dff_B_gWym8VVz4_2(.din(w_dff_B_m13h5eZ28_2),.dout(w_dff_B_gWym8VVz4_2),.clk(gclk));
	jdff dff_B_el1QXwkV8_2(.din(w_dff_B_gWym8VVz4_2),.dout(w_dff_B_el1QXwkV8_2),.clk(gclk));
	jdff dff_B_00rP6kOR2_2(.din(w_dff_B_el1QXwkV8_2),.dout(w_dff_B_00rP6kOR2_2),.clk(gclk));
	jdff dff_B_moEMgU2N6_2(.din(n1553),.dout(w_dff_B_moEMgU2N6_2),.clk(gclk));
	jdff dff_B_xwntQN6w4_1(.din(n1551),.dout(w_dff_B_xwntQN6w4_1),.clk(gclk));
	jdff dff_B_uYcsPNOh4_2(.din(n1486),.dout(w_dff_B_uYcsPNOh4_2),.clk(gclk));
	jdff dff_B_Lbb88Srh4_2(.din(w_dff_B_uYcsPNOh4_2),.dout(w_dff_B_Lbb88Srh4_2),.clk(gclk));
	jdff dff_B_GVcNLxHD1_2(.din(w_dff_B_Lbb88Srh4_2),.dout(w_dff_B_GVcNLxHD1_2),.clk(gclk));
	jdff dff_B_jOR1uSfS4_2(.din(w_dff_B_GVcNLxHD1_2),.dout(w_dff_B_jOR1uSfS4_2),.clk(gclk));
	jdff dff_B_z6asLAyO3_2(.din(w_dff_B_jOR1uSfS4_2),.dout(w_dff_B_z6asLAyO3_2),.clk(gclk));
	jdff dff_B_ZSgPdKQo3_2(.din(w_dff_B_z6asLAyO3_2),.dout(w_dff_B_ZSgPdKQo3_2),.clk(gclk));
	jdff dff_B_FMGVvcrv2_2(.din(w_dff_B_ZSgPdKQo3_2),.dout(w_dff_B_FMGVvcrv2_2),.clk(gclk));
	jdff dff_B_YyaB3ivC3_2(.din(w_dff_B_FMGVvcrv2_2),.dout(w_dff_B_YyaB3ivC3_2),.clk(gclk));
	jdff dff_B_Codtp45X7_2(.din(w_dff_B_YyaB3ivC3_2),.dout(w_dff_B_Codtp45X7_2),.clk(gclk));
	jdff dff_B_yCii9u252_2(.din(w_dff_B_Codtp45X7_2),.dout(w_dff_B_yCii9u252_2),.clk(gclk));
	jdff dff_B_c0SJOclp1_2(.din(w_dff_B_yCii9u252_2),.dout(w_dff_B_c0SJOclp1_2),.clk(gclk));
	jdff dff_B_vP2xJAAq5_2(.din(w_dff_B_c0SJOclp1_2),.dout(w_dff_B_vP2xJAAq5_2),.clk(gclk));
	jdff dff_B_Qt7bbinK7_2(.din(w_dff_B_vP2xJAAq5_2),.dout(w_dff_B_Qt7bbinK7_2),.clk(gclk));
	jdff dff_B_3HKBN7d94_2(.din(w_dff_B_Qt7bbinK7_2),.dout(w_dff_B_3HKBN7d94_2),.clk(gclk));
	jdff dff_B_wHT9FuGU0_2(.din(w_dff_B_3HKBN7d94_2),.dout(w_dff_B_wHT9FuGU0_2),.clk(gclk));
	jdff dff_B_SBpJVwLh4_2(.din(w_dff_B_wHT9FuGU0_2),.dout(w_dff_B_SBpJVwLh4_2),.clk(gclk));
	jdff dff_B_apWkk9hK8_2(.din(w_dff_B_SBpJVwLh4_2),.dout(w_dff_B_apWkk9hK8_2),.clk(gclk));
	jdff dff_B_wIsP63or6_2(.din(w_dff_B_apWkk9hK8_2),.dout(w_dff_B_wIsP63or6_2),.clk(gclk));
	jdff dff_B_lrvnhKSp0_2(.din(w_dff_B_wIsP63or6_2),.dout(w_dff_B_lrvnhKSp0_2),.clk(gclk));
	jdff dff_B_q9RLqorR2_2(.din(w_dff_B_lrvnhKSp0_2),.dout(w_dff_B_q9RLqorR2_2),.clk(gclk));
	jdff dff_B_CGmpFAkC5_2(.din(w_dff_B_q9RLqorR2_2),.dout(w_dff_B_CGmpFAkC5_2),.clk(gclk));
	jdff dff_B_Oqd0DyLu0_2(.din(w_dff_B_CGmpFAkC5_2),.dout(w_dff_B_Oqd0DyLu0_2),.clk(gclk));
	jdff dff_B_SpR4f3xO2_2(.din(w_dff_B_Oqd0DyLu0_2),.dout(w_dff_B_SpR4f3xO2_2),.clk(gclk));
	jdff dff_B_Szq79zXu1_2(.din(w_dff_B_SpR4f3xO2_2),.dout(w_dff_B_Szq79zXu1_2),.clk(gclk));
	jdff dff_B_37DtKQN75_2(.din(w_dff_B_Szq79zXu1_2),.dout(w_dff_B_37DtKQN75_2),.clk(gclk));
	jdff dff_B_4I6PdJS70_2(.din(w_dff_B_37DtKQN75_2),.dout(w_dff_B_4I6PdJS70_2),.clk(gclk));
	jdff dff_B_9jxM2aiy2_2(.din(n1489),.dout(w_dff_B_9jxM2aiy2_2),.clk(gclk));
	jdff dff_B_SqZb0rTo9_1(.din(n1487),.dout(w_dff_B_SqZb0rTo9_1),.clk(gclk));
	jdff dff_B_DdI2bIv10_2(.din(n1415),.dout(w_dff_B_DdI2bIv10_2),.clk(gclk));
	jdff dff_B_meL1Vto37_2(.din(w_dff_B_DdI2bIv10_2),.dout(w_dff_B_meL1Vto37_2),.clk(gclk));
	jdff dff_B_WKBfIGE80_2(.din(w_dff_B_meL1Vto37_2),.dout(w_dff_B_WKBfIGE80_2),.clk(gclk));
	jdff dff_B_25LFaOna2_2(.din(w_dff_B_WKBfIGE80_2),.dout(w_dff_B_25LFaOna2_2),.clk(gclk));
	jdff dff_B_YZYDP54h6_2(.din(w_dff_B_25LFaOna2_2),.dout(w_dff_B_YZYDP54h6_2),.clk(gclk));
	jdff dff_B_oQq1cGES4_2(.din(w_dff_B_YZYDP54h6_2),.dout(w_dff_B_oQq1cGES4_2),.clk(gclk));
	jdff dff_B_ASgo0ttN3_2(.din(w_dff_B_oQq1cGES4_2),.dout(w_dff_B_ASgo0ttN3_2),.clk(gclk));
	jdff dff_B_LlRcpt7T4_2(.din(w_dff_B_ASgo0ttN3_2),.dout(w_dff_B_LlRcpt7T4_2),.clk(gclk));
	jdff dff_B_drSK7fSF8_2(.din(w_dff_B_LlRcpt7T4_2),.dout(w_dff_B_drSK7fSF8_2),.clk(gclk));
	jdff dff_B_67RF45jC1_2(.din(w_dff_B_drSK7fSF8_2),.dout(w_dff_B_67RF45jC1_2),.clk(gclk));
	jdff dff_B_KFlzZAQE5_2(.din(w_dff_B_67RF45jC1_2),.dout(w_dff_B_KFlzZAQE5_2),.clk(gclk));
	jdff dff_B_72El23Cr9_2(.din(w_dff_B_KFlzZAQE5_2),.dout(w_dff_B_72El23Cr9_2),.clk(gclk));
	jdff dff_B_1u62Iwdf3_2(.din(w_dff_B_72El23Cr9_2),.dout(w_dff_B_1u62Iwdf3_2),.clk(gclk));
	jdff dff_B_67EWWzgp9_2(.din(w_dff_B_1u62Iwdf3_2),.dout(w_dff_B_67EWWzgp9_2),.clk(gclk));
	jdff dff_B_ZYYnI4144_2(.din(w_dff_B_67EWWzgp9_2),.dout(w_dff_B_ZYYnI4144_2),.clk(gclk));
	jdff dff_B_idU947px2_2(.din(w_dff_B_ZYYnI4144_2),.dout(w_dff_B_idU947px2_2),.clk(gclk));
	jdff dff_B_3ur6dyIE7_2(.din(w_dff_B_idU947px2_2),.dout(w_dff_B_3ur6dyIE7_2),.clk(gclk));
	jdff dff_B_FjvmHdvz1_2(.din(w_dff_B_3ur6dyIE7_2),.dout(w_dff_B_FjvmHdvz1_2),.clk(gclk));
	jdff dff_B_uhiHv0kY0_2(.din(w_dff_B_FjvmHdvz1_2),.dout(w_dff_B_uhiHv0kY0_2),.clk(gclk));
	jdff dff_B_hBp5jCZZ7_2(.din(w_dff_B_uhiHv0kY0_2),.dout(w_dff_B_hBp5jCZZ7_2),.clk(gclk));
	jdff dff_B_VKUptWK73_2(.din(w_dff_B_hBp5jCZZ7_2),.dout(w_dff_B_VKUptWK73_2),.clk(gclk));
	jdff dff_B_Of9tL9Os1_2(.din(w_dff_B_VKUptWK73_2),.dout(w_dff_B_Of9tL9Os1_2),.clk(gclk));
	jdff dff_B_DBt030OO6_2(.din(w_dff_B_Of9tL9Os1_2),.dout(w_dff_B_DBt030OO6_2),.clk(gclk));
	jdff dff_B_LU4nYTi48_2(.din(n1418),.dout(w_dff_B_LU4nYTi48_2),.clk(gclk));
	jdff dff_B_gUK6quCH9_1(.din(n1416),.dout(w_dff_B_gUK6quCH9_1),.clk(gclk));
	jdff dff_B_QpY56Rx47_2(.din(n1337),.dout(w_dff_B_QpY56Rx47_2),.clk(gclk));
	jdff dff_B_PNGYvlUO5_2(.din(w_dff_B_QpY56Rx47_2),.dout(w_dff_B_PNGYvlUO5_2),.clk(gclk));
	jdff dff_B_mdO820bf6_2(.din(w_dff_B_PNGYvlUO5_2),.dout(w_dff_B_mdO820bf6_2),.clk(gclk));
	jdff dff_B_5vTE0yNV6_2(.din(w_dff_B_mdO820bf6_2),.dout(w_dff_B_5vTE0yNV6_2),.clk(gclk));
	jdff dff_B_MsaBUsDF1_2(.din(w_dff_B_5vTE0yNV6_2),.dout(w_dff_B_MsaBUsDF1_2),.clk(gclk));
	jdff dff_B_l1Tc5iua5_2(.din(w_dff_B_MsaBUsDF1_2),.dout(w_dff_B_l1Tc5iua5_2),.clk(gclk));
	jdff dff_B_9rgY2KeU3_2(.din(w_dff_B_l1Tc5iua5_2),.dout(w_dff_B_9rgY2KeU3_2),.clk(gclk));
	jdff dff_B_LHsCU7050_2(.din(w_dff_B_9rgY2KeU3_2),.dout(w_dff_B_LHsCU7050_2),.clk(gclk));
	jdff dff_B_YELg5juV5_2(.din(w_dff_B_LHsCU7050_2),.dout(w_dff_B_YELg5juV5_2),.clk(gclk));
	jdff dff_B_wnag1YGW5_2(.din(w_dff_B_YELg5juV5_2),.dout(w_dff_B_wnag1YGW5_2),.clk(gclk));
	jdff dff_B_RGDX354s5_2(.din(w_dff_B_wnag1YGW5_2),.dout(w_dff_B_RGDX354s5_2),.clk(gclk));
	jdff dff_B_IYpsZfBh1_2(.din(w_dff_B_RGDX354s5_2),.dout(w_dff_B_IYpsZfBh1_2),.clk(gclk));
	jdff dff_B_EoQkHSsE8_2(.din(w_dff_B_IYpsZfBh1_2),.dout(w_dff_B_EoQkHSsE8_2),.clk(gclk));
	jdff dff_B_eHSpO7N86_2(.din(w_dff_B_EoQkHSsE8_2),.dout(w_dff_B_eHSpO7N86_2),.clk(gclk));
	jdff dff_B_5RmBExgl9_2(.din(w_dff_B_eHSpO7N86_2),.dout(w_dff_B_5RmBExgl9_2),.clk(gclk));
	jdff dff_B_nXdZS2gZ6_2(.din(w_dff_B_5RmBExgl9_2),.dout(w_dff_B_nXdZS2gZ6_2),.clk(gclk));
	jdff dff_B_uYsqBSRN2_2(.din(w_dff_B_nXdZS2gZ6_2),.dout(w_dff_B_uYsqBSRN2_2),.clk(gclk));
	jdff dff_B_3wxf5Zom0_2(.din(w_dff_B_uYsqBSRN2_2),.dout(w_dff_B_3wxf5Zom0_2),.clk(gclk));
	jdff dff_B_qZ5SdUoN1_2(.din(w_dff_B_3wxf5Zom0_2),.dout(w_dff_B_qZ5SdUoN1_2),.clk(gclk));
	jdff dff_B_TeMjtAcZ2_2(.din(w_dff_B_qZ5SdUoN1_2),.dout(w_dff_B_TeMjtAcZ2_2),.clk(gclk));
	jdff dff_B_jbWyQ2f59_1(.din(n1338),.dout(w_dff_B_jbWyQ2f59_1),.clk(gclk));
	jdff dff_B_0ba8OZ1J0_2(.din(n1252),.dout(w_dff_B_0ba8OZ1J0_2),.clk(gclk));
	jdff dff_B_x1vg9g3C0_2(.din(w_dff_B_0ba8OZ1J0_2),.dout(w_dff_B_x1vg9g3C0_2),.clk(gclk));
	jdff dff_B_G5DtcGGA6_2(.din(w_dff_B_x1vg9g3C0_2),.dout(w_dff_B_G5DtcGGA6_2),.clk(gclk));
	jdff dff_B_VkhB4F7C5_2(.din(w_dff_B_G5DtcGGA6_2),.dout(w_dff_B_VkhB4F7C5_2),.clk(gclk));
	jdff dff_B_x04ISGZH3_2(.din(w_dff_B_VkhB4F7C5_2),.dout(w_dff_B_x04ISGZH3_2),.clk(gclk));
	jdff dff_B_mcBgZVSX6_2(.din(w_dff_B_x04ISGZH3_2),.dout(w_dff_B_mcBgZVSX6_2),.clk(gclk));
	jdff dff_B_lsNpgKT07_2(.din(w_dff_B_mcBgZVSX6_2),.dout(w_dff_B_lsNpgKT07_2),.clk(gclk));
	jdff dff_B_9bQ0KpVh3_2(.din(w_dff_B_lsNpgKT07_2),.dout(w_dff_B_9bQ0KpVh3_2),.clk(gclk));
	jdff dff_B_5xfSQFPC8_2(.din(w_dff_B_9bQ0KpVh3_2),.dout(w_dff_B_5xfSQFPC8_2),.clk(gclk));
	jdff dff_B_JPwgvdJI1_2(.din(w_dff_B_5xfSQFPC8_2),.dout(w_dff_B_JPwgvdJI1_2),.clk(gclk));
	jdff dff_B_d7EkmAa06_2(.din(w_dff_B_JPwgvdJI1_2),.dout(w_dff_B_d7EkmAa06_2),.clk(gclk));
	jdff dff_B_NbpgrCmA4_2(.din(w_dff_B_d7EkmAa06_2),.dout(w_dff_B_NbpgrCmA4_2),.clk(gclk));
	jdff dff_B_95BlcFnV7_2(.din(w_dff_B_NbpgrCmA4_2),.dout(w_dff_B_95BlcFnV7_2),.clk(gclk));
	jdff dff_B_XUVcPYcI5_2(.din(w_dff_B_95BlcFnV7_2),.dout(w_dff_B_XUVcPYcI5_2),.clk(gclk));
	jdff dff_B_ukNE9JBI9_2(.din(w_dff_B_XUVcPYcI5_2),.dout(w_dff_B_ukNE9JBI9_2),.clk(gclk));
	jdff dff_B_LYKAZrm17_2(.din(w_dff_B_ukNE9JBI9_2),.dout(w_dff_B_LYKAZrm17_2),.clk(gclk));
	jdff dff_B_TiTJtm369_2(.din(w_dff_B_LYKAZrm17_2),.dout(w_dff_B_TiTJtm369_2),.clk(gclk));
	jdff dff_B_wmuiS3qd6_2(.din(w_dff_B_TiTJtm369_2),.dout(w_dff_B_wmuiS3qd6_2),.clk(gclk));
	jdff dff_B_AvhsdWwx0_1(.din(n1253),.dout(w_dff_B_AvhsdWwx0_1),.clk(gclk));
	jdff dff_B_Oh1zq6Mh6_2(.din(n1161),.dout(w_dff_B_Oh1zq6Mh6_2),.clk(gclk));
	jdff dff_B_oHnryv4o5_2(.din(w_dff_B_Oh1zq6Mh6_2),.dout(w_dff_B_oHnryv4o5_2),.clk(gclk));
	jdff dff_B_yC4jijt47_2(.din(w_dff_B_oHnryv4o5_2),.dout(w_dff_B_yC4jijt47_2),.clk(gclk));
	jdff dff_B_XfYe9kqy7_2(.din(w_dff_B_yC4jijt47_2),.dout(w_dff_B_XfYe9kqy7_2),.clk(gclk));
	jdff dff_B_iLeXhq9f2_2(.din(w_dff_B_XfYe9kqy7_2),.dout(w_dff_B_iLeXhq9f2_2),.clk(gclk));
	jdff dff_B_OL9yJHgO8_2(.din(w_dff_B_iLeXhq9f2_2),.dout(w_dff_B_OL9yJHgO8_2),.clk(gclk));
	jdff dff_B_J7aiNuZL2_2(.din(w_dff_B_OL9yJHgO8_2),.dout(w_dff_B_J7aiNuZL2_2),.clk(gclk));
	jdff dff_B_k3gITvSR1_2(.din(w_dff_B_J7aiNuZL2_2),.dout(w_dff_B_k3gITvSR1_2),.clk(gclk));
	jdff dff_B_YeRToyGb0_2(.din(w_dff_B_k3gITvSR1_2),.dout(w_dff_B_YeRToyGb0_2),.clk(gclk));
	jdff dff_B_zBJ5tJdi9_2(.din(w_dff_B_YeRToyGb0_2),.dout(w_dff_B_zBJ5tJdi9_2),.clk(gclk));
	jdff dff_B_tMeUQAr51_2(.din(w_dff_B_zBJ5tJdi9_2),.dout(w_dff_B_tMeUQAr51_2),.clk(gclk));
	jdff dff_B_vyLppwd93_2(.din(w_dff_B_tMeUQAr51_2),.dout(w_dff_B_vyLppwd93_2),.clk(gclk));
	jdff dff_B_guJvyLC42_2(.din(w_dff_B_vyLppwd93_2),.dout(w_dff_B_guJvyLC42_2),.clk(gclk));
	jdff dff_B_U0qPwURo8_2(.din(w_dff_B_guJvyLC42_2),.dout(w_dff_B_U0qPwURo8_2),.clk(gclk));
	jdff dff_B_7XPxFGYO7_2(.din(w_dff_B_U0qPwURo8_2),.dout(w_dff_B_7XPxFGYO7_2),.clk(gclk));
	jdff dff_B_SbRg2T466_2(.din(w_dff_B_7XPxFGYO7_2),.dout(w_dff_B_SbRg2T466_2),.clk(gclk));
	jdff dff_B_jDExplnb2_1(.din(n1162),.dout(w_dff_B_jDExplnb2_1),.clk(gclk));
	jdff dff_B_hWqmaJz68_2(.din(n1063),.dout(w_dff_B_hWqmaJz68_2),.clk(gclk));
	jdff dff_B_Au2MqRS42_2(.din(w_dff_B_hWqmaJz68_2),.dout(w_dff_B_Au2MqRS42_2),.clk(gclk));
	jdff dff_B_K0rMzYeN2_2(.din(w_dff_B_Au2MqRS42_2),.dout(w_dff_B_K0rMzYeN2_2),.clk(gclk));
	jdff dff_B_dOtyYH094_2(.din(w_dff_B_K0rMzYeN2_2),.dout(w_dff_B_dOtyYH094_2),.clk(gclk));
	jdff dff_B_FWho8mwh2_2(.din(w_dff_B_dOtyYH094_2),.dout(w_dff_B_FWho8mwh2_2),.clk(gclk));
	jdff dff_B_cFjIApdh3_2(.din(w_dff_B_FWho8mwh2_2),.dout(w_dff_B_cFjIApdh3_2),.clk(gclk));
	jdff dff_B_Q8cwLoy62_2(.din(w_dff_B_cFjIApdh3_2),.dout(w_dff_B_Q8cwLoy62_2),.clk(gclk));
	jdff dff_B_dnR4MMU02_2(.din(w_dff_B_Q8cwLoy62_2),.dout(w_dff_B_dnR4MMU02_2),.clk(gclk));
	jdff dff_B_NZ6F6M5D1_2(.din(w_dff_B_dnR4MMU02_2),.dout(w_dff_B_NZ6F6M5D1_2),.clk(gclk));
	jdff dff_B_qty4MBao8_2(.din(w_dff_B_NZ6F6M5D1_2),.dout(w_dff_B_qty4MBao8_2),.clk(gclk));
	jdff dff_B_zJ69d5Q91_2(.din(w_dff_B_qty4MBao8_2),.dout(w_dff_B_zJ69d5Q91_2),.clk(gclk));
	jdff dff_B_QonhRK344_2(.din(w_dff_B_zJ69d5Q91_2),.dout(w_dff_B_QonhRK344_2),.clk(gclk));
	jdff dff_B_NbIEAUxQ8_2(.din(w_dff_B_QonhRK344_2),.dout(w_dff_B_NbIEAUxQ8_2),.clk(gclk));
	jdff dff_B_0BghZfKE4_2(.din(w_dff_B_NbIEAUxQ8_2),.dout(w_dff_B_0BghZfKE4_2),.clk(gclk));
	jdff dff_B_ZbX2H2M93_1(.din(n1064),.dout(w_dff_B_ZbX2H2M93_1),.clk(gclk));
	jdff dff_B_byeQr5fB7_2(.din(n964),.dout(w_dff_B_byeQr5fB7_2),.clk(gclk));
	jdff dff_B_Dj2olG4I4_2(.din(w_dff_B_byeQr5fB7_2),.dout(w_dff_B_Dj2olG4I4_2),.clk(gclk));
	jdff dff_B_kfBuFU4K3_2(.din(w_dff_B_Dj2olG4I4_2),.dout(w_dff_B_kfBuFU4K3_2),.clk(gclk));
	jdff dff_B_ZY8BgPa79_2(.din(w_dff_B_kfBuFU4K3_2),.dout(w_dff_B_ZY8BgPa79_2),.clk(gclk));
	jdff dff_B_aKEU5xNU8_2(.din(w_dff_B_ZY8BgPa79_2),.dout(w_dff_B_aKEU5xNU8_2),.clk(gclk));
	jdff dff_B_wVQ1QvgF0_2(.din(w_dff_B_aKEU5xNU8_2),.dout(w_dff_B_wVQ1QvgF0_2),.clk(gclk));
	jdff dff_B_Qu8sGOb56_2(.din(w_dff_B_wVQ1QvgF0_2),.dout(w_dff_B_Qu8sGOb56_2),.clk(gclk));
	jdff dff_B_GWKSrfmK5_2(.din(w_dff_B_Qu8sGOb56_2),.dout(w_dff_B_GWKSrfmK5_2),.clk(gclk));
	jdff dff_B_YleM33fm8_2(.din(w_dff_B_GWKSrfmK5_2),.dout(w_dff_B_YleM33fm8_2),.clk(gclk));
	jdff dff_B_WqdSsM3X2_2(.din(w_dff_B_YleM33fm8_2),.dout(w_dff_B_WqdSsM3X2_2),.clk(gclk));
	jdff dff_B_BvutzHhp9_2(.din(w_dff_B_WqdSsM3X2_2),.dout(w_dff_B_BvutzHhp9_2),.clk(gclk));
	jdff dff_B_5pO8copD6_2(.din(w_dff_B_BvutzHhp9_2),.dout(w_dff_B_5pO8copD6_2),.clk(gclk));
	jdff dff_B_MZbWiYZP4_1(.din(n965),.dout(w_dff_B_MZbWiYZP4_1),.clk(gclk));
	jdff dff_B_SKbly1jy3_2(.din(n862),.dout(w_dff_B_SKbly1jy3_2),.clk(gclk));
	jdff dff_B_xuApQhmg9_2(.din(w_dff_B_SKbly1jy3_2),.dout(w_dff_B_xuApQhmg9_2),.clk(gclk));
	jdff dff_B_hJVRdHFJ2_2(.din(w_dff_B_xuApQhmg9_2),.dout(w_dff_B_hJVRdHFJ2_2),.clk(gclk));
	jdff dff_B_HV9xsRd55_2(.din(w_dff_B_hJVRdHFJ2_2),.dout(w_dff_B_HV9xsRd55_2),.clk(gclk));
	jdff dff_B_iHUvig0Q5_2(.din(w_dff_B_HV9xsRd55_2),.dout(w_dff_B_iHUvig0Q5_2),.clk(gclk));
	jdff dff_B_rTbsJc0U3_2(.din(w_dff_B_iHUvig0Q5_2),.dout(w_dff_B_rTbsJc0U3_2),.clk(gclk));
	jdff dff_B_hYKJftjW7_2(.din(w_dff_B_rTbsJc0U3_2),.dout(w_dff_B_hYKJftjW7_2),.clk(gclk));
	jdff dff_B_IcvyUOpV9_2(.din(w_dff_B_hYKJftjW7_2),.dout(w_dff_B_IcvyUOpV9_2),.clk(gclk));
	jdff dff_B_ZX1ox3bo8_2(.din(w_dff_B_IcvyUOpV9_2),.dout(w_dff_B_ZX1ox3bo8_2),.clk(gclk));
	jdff dff_B_9QT1Zgay3_2(.din(w_dff_B_ZX1ox3bo8_2),.dout(w_dff_B_9QT1Zgay3_2),.clk(gclk));
	jdff dff_B_4XuRTRbF5_1(.din(n863),.dout(w_dff_B_4XuRTRbF5_1),.clk(gclk));
	jdff dff_B_Yo4caIpC5_2(.din(n764),.dout(w_dff_B_Yo4caIpC5_2),.clk(gclk));
	jdff dff_B_so2WwinY5_2(.din(w_dff_B_Yo4caIpC5_2),.dout(w_dff_B_so2WwinY5_2),.clk(gclk));
	jdff dff_B_dPnlfqXA4_2(.din(w_dff_B_so2WwinY5_2),.dout(w_dff_B_dPnlfqXA4_2),.clk(gclk));
	jdff dff_B_PtlK4VvW2_2(.din(w_dff_B_dPnlfqXA4_2),.dout(w_dff_B_PtlK4VvW2_2),.clk(gclk));
	jdff dff_B_qpBA0bLC0_2(.din(w_dff_B_PtlK4VvW2_2),.dout(w_dff_B_qpBA0bLC0_2),.clk(gclk));
	jdff dff_B_TrqQCWBP1_2(.din(w_dff_B_qpBA0bLC0_2),.dout(w_dff_B_TrqQCWBP1_2),.clk(gclk));
	jdff dff_B_p8jGFLgk1_2(.din(w_dff_B_TrqQCWBP1_2),.dout(w_dff_B_p8jGFLgk1_2),.clk(gclk));
	jdff dff_B_jSQRXVU61_2(.din(w_dff_B_p8jGFLgk1_2),.dout(w_dff_B_jSQRXVU61_2),.clk(gclk));
	jdff dff_B_kiu8i9rh1_2(.din(n779),.dout(w_dff_B_kiu8i9rh1_2),.clk(gclk));
	jdff dff_B_2iAqGD1d5_2(.din(w_dff_B_kiu8i9rh1_2),.dout(w_dff_B_2iAqGD1d5_2),.clk(gclk));
	jdff dff_B_CWBZljMi1_2(.din(w_dff_B_2iAqGD1d5_2),.dout(w_dff_B_CWBZljMi1_2),.clk(gclk));
	jdff dff_B_tz9i5LDL6_1(.din(n765),.dout(w_dff_B_tz9i5LDL6_1),.clk(gclk));
	jdff dff_B_0RbaoSE57_1(.din(w_dff_B_tz9i5LDL6_1),.dout(w_dff_B_0RbaoSE57_1),.clk(gclk));
	jdff dff_B_n1Y9jby81_1(.din(w_dff_B_0RbaoSE57_1),.dout(w_dff_B_n1Y9jby81_1),.clk(gclk));
	jdff dff_B_KH11dAwP7_2(.din(n674),.dout(w_dff_B_KH11dAwP7_2),.clk(gclk));
	jdff dff_B_VYk08moP0_2(.din(w_dff_B_KH11dAwP7_2),.dout(w_dff_B_VYk08moP0_2),.clk(gclk));
	jdff dff_B_WlqYnXpZ5_2(.din(w_dff_B_VYk08moP0_2),.dout(w_dff_B_WlqYnXpZ5_2),.clk(gclk));
	jdff dff_B_7RAsqCfJ4_0(.din(n679),.dout(w_dff_B_7RAsqCfJ4_0),.clk(gclk));
	jdff dff_B_wbmtKYiJ5_0(.din(w_dff_B_7RAsqCfJ4_0),.dout(w_dff_B_wbmtKYiJ5_0),.clk(gclk));
	jdff dff_A_gMUQkBHE4_0(.dout(w_n586_0[0]),.din(w_dff_A_gMUQkBHE4_0),.clk(gclk));
	jdff dff_A_QsWz4K3z1_0(.dout(w_dff_A_gMUQkBHE4_0),.din(w_dff_A_QsWz4K3z1_0),.clk(gclk));
	jdff dff_A_boBTgFYQ0_1(.dout(w_n586_0[1]),.din(w_dff_A_boBTgFYQ0_1),.clk(gclk));
	jdff dff_A_5I1E6S8T8_1(.dout(w_dff_A_boBTgFYQ0_1),.din(w_dff_A_5I1E6S8T8_1),.clk(gclk));
	jdff dff_B_wMZixJ0t3_1(.din(n1788),.dout(w_dff_B_wMZixJ0t3_1),.clk(gclk));
	jdff dff_A_KNttCfjm4_1(.dout(w_n1770_0[1]),.din(w_dff_A_KNttCfjm4_1),.clk(gclk));
	jdff dff_B_B1fTr3EQ0_1(.din(n1768),.dout(w_dff_B_B1fTr3EQ0_1),.clk(gclk));
	jdff dff_B_IKesATjm2_2(.din(n1739),.dout(w_dff_B_IKesATjm2_2),.clk(gclk));
	jdff dff_B_Rai0w08W8_2(.din(w_dff_B_IKesATjm2_2),.dout(w_dff_B_Rai0w08W8_2),.clk(gclk));
	jdff dff_B_BHpDV6SL2_2(.din(w_dff_B_Rai0w08W8_2),.dout(w_dff_B_BHpDV6SL2_2),.clk(gclk));
	jdff dff_B_Ic9OiRAe4_2(.din(w_dff_B_BHpDV6SL2_2),.dout(w_dff_B_Ic9OiRAe4_2),.clk(gclk));
	jdff dff_B_UeY8FAKR6_2(.din(w_dff_B_Ic9OiRAe4_2),.dout(w_dff_B_UeY8FAKR6_2),.clk(gclk));
	jdff dff_B_dLcPpB2E1_2(.din(w_dff_B_UeY8FAKR6_2),.dout(w_dff_B_dLcPpB2E1_2),.clk(gclk));
	jdff dff_B_i1H8cDHp2_2(.din(w_dff_B_dLcPpB2E1_2),.dout(w_dff_B_i1H8cDHp2_2),.clk(gclk));
	jdff dff_B_PGXolDR15_2(.din(w_dff_B_i1H8cDHp2_2),.dout(w_dff_B_PGXolDR15_2),.clk(gclk));
	jdff dff_B_4fuqVPcN6_2(.din(w_dff_B_PGXolDR15_2),.dout(w_dff_B_4fuqVPcN6_2),.clk(gclk));
	jdff dff_B_1fTpE24b6_2(.din(w_dff_B_4fuqVPcN6_2),.dout(w_dff_B_1fTpE24b6_2),.clk(gclk));
	jdff dff_B_BIO2Jqv37_2(.din(w_dff_B_1fTpE24b6_2),.dout(w_dff_B_BIO2Jqv37_2),.clk(gclk));
	jdff dff_B_z0aytx1A7_2(.din(w_dff_B_BIO2Jqv37_2),.dout(w_dff_B_z0aytx1A7_2),.clk(gclk));
	jdff dff_B_5KqVGXXJ5_2(.din(w_dff_B_z0aytx1A7_2),.dout(w_dff_B_5KqVGXXJ5_2),.clk(gclk));
	jdff dff_B_lkRuobfB7_2(.din(w_dff_B_5KqVGXXJ5_2),.dout(w_dff_B_lkRuobfB7_2),.clk(gclk));
	jdff dff_B_pBjD1pgZ8_2(.din(w_dff_B_lkRuobfB7_2),.dout(w_dff_B_pBjD1pgZ8_2),.clk(gclk));
	jdff dff_B_KnHscsVw9_2(.din(w_dff_B_pBjD1pgZ8_2),.dout(w_dff_B_KnHscsVw9_2),.clk(gclk));
	jdff dff_B_r6oHtWmn8_2(.din(w_dff_B_KnHscsVw9_2),.dout(w_dff_B_r6oHtWmn8_2),.clk(gclk));
	jdff dff_B_9I2K4W1T5_2(.din(w_dff_B_r6oHtWmn8_2),.dout(w_dff_B_9I2K4W1T5_2),.clk(gclk));
	jdff dff_B_EpZG7LPc1_2(.din(w_dff_B_9I2K4W1T5_2),.dout(w_dff_B_EpZG7LPc1_2),.clk(gclk));
	jdff dff_B_ezVLhejA8_2(.din(w_dff_B_EpZG7LPc1_2),.dout(w_dff_B_ezVLhejA8_2),.clk(gclk));
	jdff dff_B_IVpYyiNX3_2(.din(w_dff_B_ezVLhejA8_2),.dout(w_dff_B_IVpYyiNX3_2),.clk(gclk));
	jdff dff_B_gJuf6WMv4_2(.din(w_dff_B_IVpYyiNX3_2),.dout(w_dff_B_gJuf6WMv4_2),.clk(gclk));
	jdff dff_B_AyvtIffD3_2(.din(w_dff_B_gJuf6WMv4_2),.dout(w_dff_B_AyvtIffD3_2),.clk(gclk));
	jdff dff_B_i72cYq3q2_2(.din(w_dff_B_AyvtIffD3_2),.dout(w_dff_B_i72cYq3q2_2),.clk(gclk));
	jdff dff_B_E2NdmMMM5_2(.din(w_dff_B_i72cYq3q2_2),.dout(w_dff_B_E2NdmMMM5_2),.clk(gclk));
	jdff dff_B_kqNXt3mr9_2(.din(w_dff_B_E2NdmMMM5_2),.dout(w_dff_B_kqNXt3mr9_2),.clk(gclk));
	jdff dff_B_m0lY1gc95_2(.din(w_dff_B_kqNXt3mr9_2),.dout(w_dff_B_m0lY1gc95_2),.clk(gclk));
	jdff dff_B_zWGfcJdG2_2(.din(w_dff_B_m0lY1gc95_2),.dout(w_dff_B_zWGfcJdG2_2),.clk(gclk));
	jdff dff_B_kDVPxAXA1_2(.din(w_dff_B_zWGfcJdG2_2),.dout(w_dff_B_kDVPxAXA1_2),.clk(gclk));
	jdff dff_B_7rArwP4H7_2(.din(w_dff_B_kDVPxAXA1_2),.dout(w_dff_B_7rArwP4H7_2),.clk(gclk));
	jdff dff_B_fF0xbfAr5_2(.din(w_dff_B_7rArwP4H7_2),.dout(w_dff_B_fF0xbfAr5_2),.clk(gclk));
	jdff dff_B_WP6hLDlV0_2(.din(w_dff_B_fF0xbfAr5_2),.dout(w_dff_B_WP6hLDlV0_2),.clk(gclk));
	jdff dff_B_bjdS5EFx7_2(.din(w_dff_B_WP6hLDlV0_2),.dout(w_dff_B_bjdS5EFx7_2),.clk(gclk));
	jdff dff_B_WsFgGShv2_2(.din(w_dff_B_bjdS5EFx7_2),.dout(w_dff_B_WsFgGShv2_2),.clk(gclk));
	jdff dff_B_CwW7ib2w6_2(.din(w_dff_B_WsFgGShv2_2),.dout(w_dff_B_CwW7ib2w6_2),.clk(gclk));
	jdff dff_B_Qjjt0w3S1_2(.din(w_dff_B_CwW7ib2w6_2),.dout(w_dff_B_Qjjt0w3S1_2),.clk(gclk));
	jdff dff_B_n7DXsGIr8_2(.din(w_dff_B_Qjjt0w3S1_2),.dout(w_dff_B_n7DXsGIr8_2),.clk(gclk));
	jdff dff_B_6pjK2m7T6_2(.din(w_dff_B_n7DXsGIr8_2),.dout(w_dff_B_6pjK2m7T6_2),.clk(gclk));
	jdff dff_B_Nsr8LsGd2_2(.din(w_dff_B_6pjK2m7T6_2),.dout(w_dff_B_Nsr8LsGd2_2),.clk(gclk));
	jdff dff_B_9jwiKTXR0_2(.din(n1742),.dout(w_dff_B_9jwiKTXR0_2),.clk(gclk));
	jdff dff_B_Ds0vKPck1_1(.din(n1740),.dout(w_dff_B_Ds0vKPck1_1),.clk(gclk));
	jdff dff_B_de1NgIVY0_2(.din(n1704),.dout(w_dff_B_de1NgIVY0_2),.clk(gclk));
	jdff dff_B_b5W6mgeO0_2(.din(w_dff_B_de1NgIVY0_2),.dout(w_dff_B_b5W6mgeO0_2),.clk(gclk));
	jdff dff_B_vijT05ax8_2(.din(w_dff_B_b5W6mgeO0_2),.dout(w_dff_B_vijT05ax8_2),.clk(gclk));
	jdff dff_B_06ECoTsA1_2(.din(w_dff_B_vijT05ax8_2),.dout(w_dff_B_06ECoTsA1_2),.clk(gclk));
	jdff dff_B_4Opjvcgd9_2(.din(w_dff_B_06ECoTsA1_2),.dout(w_dff_B_4Opjvcgd9_2),.clk(gclk));
	jdff dff_B_e4cTjmbp1_2(.din(w_dff_B_4Opjvcgd9_2),.dout(w_dff_B_e4cTjmbp1_2),.clk(gclk));
	jdff dff_B_MxMPcwTN8_2(.din(w_dff_B_e4cTjmbp1_2),.dout(w_dff_B_MxMPcwTN8_2),.clk(gclk));
	jdff dff_B_RlxPCt5t7_2(.din(w_dff_B_MxMPcwTN8_2),.dout(w_dff_B_RlxPCt5t7_2),.clk(gclk));
	jdff dff_B_Ov1Z5Iql3_2(.din(w_dff_B_RlxPCt5t7_2),.dout(w_dff_B_Ov1Z5Iql3_2),.clk(gclk));
	jdff dff_B_5sW30sEJ3_2(.din(w_dff_B_Ov1Z5Iql3_2),.dout(w_dff_B_5sW30sEJ3_2),.clk(gclk));
	jdff dff_B_IbpwfenH7_2(.din(w_dff_B_5sW30sEJ3_2),.dout(w_dff_B_IbpwfenH7_2),.clk(gclk));
	jdff dff_B_Hp3WxBEw7_2(.din(w_dff_B_IbpwfenH7_2),.dout(w_dff_B_Hp3WxBEw7_2),.clk(gclk));
	jdff dff_B_W7J7j9fu3_2(.din(w_dff_B_Hp3WxBEw7_2),.dout(w_dff_B_W7J7j9fu3_2),.clk(gclk));
	jdff dff_B_F9xq26UU0_2(.din(w_dff_B_W7J7j9fu3_2),.dout(w_dff_B_F9xq26UU0_2),.clk(gclk));
	jdff dff_B_uss7Niaf0_2(.din(w_dff_B_F9xq26UU0_2),.dout(w_dff_B_uss7Niaf0_2),.clk(gclk));
	jdff dff_B_kHcqLz9C8_2(.din(w_dff_B_uss7Niaf0_2),.dout(w_dff_B_kHcqLz9C8_2),.clk(gclk));
	jdff dff_B_kb6HjZos8_2(.din(w_dff_B_kHcqLz9C8_2),.dout(w_dff_B_kb6HjZos8_2),.clk(gclk));
	jdff dff_B_6AtXfxs03_2(.din(w_dff_B_kb6HjZos8_2),.dout(w_dff_B_6AtXfxs03_2),.clk(gclk));
	jdff dff_B_vm4lwmeR7_2(.din(w_dff_B_6AtXfxs03_2),.dout(w_dff_B_vm4lwmeR7_2),.clk(gclk));
	jdff dff_B_kwb45Ov56_2(.din(w_dff_B_vm4lwmeR7_2),.dout(w_dff_B_kwb45Ov56_2),.clk(gclk));
	jdff dff_B_bfdsRwPH6_2(.din(w_dff_B_kwb45Ov56_2),.dout(w_dff_B_bfdsRwPH6_2),.clk(gclk));
	jdff dff_B_fta1R7qd2_2(.din(w_dff_B_bfdsRwPH6_2),.dout(w_dff_B_fta1R7qd2_2),.clk(gclk));
	jdff dff_B_qKCwzhgO0_2(.din(w_dff_B_fta1R7qd2_2),.dout(w_dff_B_qKCwzhgO0_2),.clk(gclk));
	jdff dff_B_3e0gmAiY9_2(.din(w_dff_B_qKCwzhgO0_2),.dout(w_dff_B_3e0gmAiY9_2),.clk(gclk));
	jdff dff_B_D0jj3TBw8_2(.din(w_dff_B_3e0gmAiY9_2),.dout(w_dff_B_D0jj3TBw8_2),.clk(gclk));
	jdff dff_B_3DM79s4j6_2(.din(w_dff_B_D0jj3TBw8_2),.dout(w_dff_B_3DM79s4j6_2),.clk(gclk));
	jdff dff_B_WDkaVjEG4_2(.din(w_dff_B_3DM79s4j6_2),.dout(w_dff_B_WDkaVjEG4_2),.clk(gclk));
	jdff dff_B_mE720zBR7_2(.din(w_dff_B_WDkaVjEG4_2),.dout(w_dff_B_mE720zBR7_2),.clk(gclk));
	jdff dff_B_nnSDFqqO5_2(.din(w_dff_B_mE720zBR7_2),.dout(w_dff_B_nnSDFqqO5_2),.clk(gclk));
	jdff dff_B_FDLpQtwo4_2(.din(w_dff_B_nnSDFqqO5_2),.dout(w_dff_B_FDLpQtwo4_2),.clk(gclk));
	jdff dff_B_IFUkFm247_2(.din(w_dff_B_FDLpQtwo4_2),.dout(w_dff_B_IFUkFm247_2),.clk(gclk));
	jdff dff_B_IkRLZFXu5_2(.din(w_dff_B_IFUkFm247_2),.dout(w_dff_B_IkRLZFXu5_2),.clk(gclk));
	jdff dff_B_htxzZT5S3_2(.din(w_dff_B_IkRLZFXu5_2),.dout(w_dff_B_htxzZT5S3_2),.clk(gclk));
	jdff dff_B_plmIA1TV1_2(.din(w_dff_B_htxzZT5S3_2),.dout(w_dff_B_plmIA1TV1_2),.clk(gclk));
	jdff dff_B_gkmta5bM2_2(.din(w_dff_B_plmIA1TV1_2),.dout(w_dff_B_gkmta5bM2_2),.clk(gclk));
	jdff dff_B_0kbzAFr32_2(.din(w_dff_B_gkmta5bM2_2),.dout(w_dff_B_0kbzAFr32_2),.clk(gclk));
	jdff dff_B_jnITGK5r1_2(.din(n1707),.dout(w_dff_B_jnITGK5r1_2),.clk(gclk));
	jdff dff_B_Q2VG2qeG7_1(.din(n1705),.dout(w_dff_B_Q2VG2qeG7_1),.clk(gclk));
	jdff dff_B_nEq5dsI15_2(.din(n1663),.dout(w_dff_B_nEq5dsI15_2),.clk(gclk));
	jdff dff_B_bt0OS5xJ5_2(.din(w_dff_B_nEq5dsI15_2),.dout(w_dff_B_bt0OS5xJ5_2),.clk(gclk));
	jdff dff_B_u6oKuM3D1_2(.din(w_dff_B_bt0OS5xJ5_2),.dout(w_dff_B_u6oKuM3D1_2),.clk(gclk));
	jdff dff_B_imPLhoGZ6_2(.din(w_dff_B_u6oKuM3D1_2),.dout(w_dff_B_imPLhoGZ6_2),.clk(gclk));
	jdff dff_B_ZBchDq5z7_2(.din(w_dff_B_imPLhoGZ6_2),.dout(w_dff_B_ZBchDq5z7_2),.clk(gclk));
	jdff dff_B_lM5YyZWH9_2(.din(w_dff_B_ZBchDq5z7_2),.dout(w_dff_B_lM5YyZWH9_2),.clk(gclk));
	jdff dff_B_2tb0n7h61_2(.din(w_dff_B_lM5YyZWH9_2),.dout(w_dff_B_2tb0n7h61_2),.clk(gclk));
	jdff dff_B_Oqer9GfB0_2(.din(w_dff_B_2tb0n7h61_2),.dout(w_dff_B_Oqer9GfB0_2),.clk(gclk));
	jdff dff_B_yrnLnOZL7_2(.din(w_dff_B_Oqer9GfB0_2),.dout(w_dff_B_yrnLnOZL7_2),.clk(gclk));
	jdff dff_B_OhAdsSST3_2(.din(w_dff_B_yrnLnOZL7_2),.dout(w_dff_B_OhAdsSST3_2),.clk(gclk));
	jdff dff_B_LL7oUxp97_2(.din(w_dff_B_OhAdsSST3_2),.dout(w_dff_B_LL7oUxp97_2),.clk(gclk));
	jdff dff_B_CEhMRDyD3_2(.din(w_dff_B_LL7oUxp97_2),.dout(w_dff_B_CEhMRDyD3_2),.clk(gclk));
	jdff dff_B_3GH4dFwd9_2(.din(w_dff_B_CEhMRDyD3_2),.dout(w_dff_B_3GH4dFwd9_2),.clk(gclk));
	jdff dff_B_zun5r30O1_2(.din(w_dff_B_3GH4dFwd9_2),.dout(w_dff_B_zun5r30O1_2),.clk(gclk));
	jdff dff_B_su6K61sy8_2(.din(w_dff_B_zun5r30O1_2),.dout(w_dff_B_su6K61sy8_2),.clk(gclk));
	jdff dff_B_YVclku7K5_2(.din(w_dff_B_su6K61sy8_2),.dout(w_dff_B_YVclku7K5_2),.clk(gclk));
	jdff dff_B_wGYrY7Cg5_2(.din(w_dff_B_YVclku7K5_2),.dout(w_dff_B_wGYrY7Cg5_2),.clk(gclk));
	jdff dff_B_UQ2rPhQl3_2(.din(w_dff_B_wGYrY7Cg5_2),.dout(w_dff_B_UQ2rPhQl3_2),.clk(gclk));
	jdff dff_B_TDkYhL5f6_2(.din(w_dff_B_UQ2rPhQl3_2),.dout(w_dff_B_TDkYhL5f6_2),.clk(gclk));
	jdff dff_B_cA0IyRao7_2(.din(w_dff_B_TDkYhL5f6_2),.dout(w_dff_B_cA0IyRao7_2),.clk(gclk));
	jdff dff_B_f0MxiaFR9_2(.din(w_dff_B_cA0IyRao7_2),.dout(w_dff_B_f0MxiaFR9_2),.clk(gclk));
	jdff dff_B_8I4XB39R3_2(.din(w_dff_B_f0MxiaFR9_2),.dout(w_dff_B_8I4XB39R3_2),.clk(gclk));
	jdff dff_B_wq7CeCXu6_2(.din(w_dff_B_8I4XB39R3_2),.dout(w_dff_B_wq7CeCXu6_2),.clk(gclk));
	jdff dff_B_opQ4cZJN1_2(.din(w_dff_B_wq7CeCXu6_2),.dout(w_dff_B_opQ4cZJN1_2),.clk(gclk));
	jdff dff_B_fg2oMBcn2_2(.din(w_dff_B_opQ4cZJN1_2),.dout(w_dff_B_fg2oMBcn2_2),.clk(gclk));
	jdff dff_B_0S6KNmK59_2(.din(w_dff_B_fg2oMBcn2_2),.dout(w_dff_B_0S6KNmK59_2),.clk(gclk));
	jdff dff_B_Yut8iCD26_2(.din(w_dff_B_0S6KNmK59_2),.dout(w_dff_B_Yut8iCD26_2),.clk(gclk));
	jdff dff_B_Jgtdt7or8_2(.din(w_dff_B_Yut8iCD26_2),.dout(w_dff_B_Jgtdt7or8_2),.clk(gclk));
	jdff dff_B_FEzIH7wK5_2(.din(w_dff_B_Jgtdt7or8_2),.dout(w_dff_B_FEzIH7wK5_2),.clk(gclk));
	jdff dff_B_uzfU4WN12_2(.din(w_dff_B_FEzIH7wK5_2),.dout(w_dff_B_uzfU4WN12_2),.clk(gclk));
	jdff dff_B_ILFyqgTb3_2(.din(w_dff_B_uzfU4WN12_2),.dout(w_dff_B_ILFyqgTb3_2),.clk(gclk));
	jdff dff_B_qEikJNAa5_2(.din(w_dff_B_ILFyqgTb3_2),.dout(w_dff_B_qEikJNAa5_2),.clk(gclk));
	jdff dff_B_dT6I9ojo5_2(.din(w_dff_B_qEikJNAa5_2),.dout(w_dff_B_dT6I9ojo5_2),.clk(gclk));
	jdff dff_B_SwtKcqr72_2(.din(n1666),.dout(w_dff_B_SwtKcqr72_2),.clk(gclk));
	jdff dff_B_nxmiywbP2_1(.din(n1664),.dout(w_dff_B_nxmiywbP2_1),.clk(gclk));
	jdff dff_B_8AFNGO8B9_2(.din(n1612),.dout(w_dff_B_8AFNGO8B9_2),.clk(gclk));
	jdff dff_B_k8dAsls96_2(.din(w_dff_B_8AFNGO8B9_2),.dout(w_dff_B_k8dAsls96_2),.clk(gclk));
	jdff dff_B_vOnenEBR8_2(.din(w_dff_B_k8dAsls96_2),.dout(w_dff_B_vOnenEBR8_2),.clk(gclk));
	jdff dff_B_5oqkgYQU8_2(.din(w_dff_B_vOnenEBR8_2),.dout(w_dff_B_5oqkgYQU8_2),.clk(gclk));
	jdff dff_B_MHA9LkyP6_2(.din(w_dff_B_5oqkgYQU8_2),.dout(w_dff_B_MHA9LkyP6_2),.clk(gclk));
	jdff dff_B_uYd7uQAA2_2(.din(w_dff_B_MHA9LkyP6_2),.dout(w_dff_B_uYd7uQAA2_2),.clk(gclk));
	jdff dff_B_obDSMITW2_2(.din(w_dff_B_uYd7uQAA2_2),.dout(w_dff_B_obDSMITW2_2),.clk(gclk));
	jdff dff_B_FcUHe5sT9_2(.din(w_dff_B_obDSMITW2_2),.dout(w_dff_B_FcUHe5sT9_2),.clk(gclk));
	jdff dff_B_OfmaWxW15_2(.din(w_dff_B_FcUHe5sT9_2),.dout(w_dff_B_OfmaWxW15_2),.clk(gclk));
	jdff dff_B_3wc7Qi0x9_2(.din(w_dff_B_OfmaWxW15_2),.dout(w_dff_B_3wc7Qi0x9_2),.clk(gclk));
	jdff dff_B_SDpKUlTa3_2(.din(w_dff_B_3wc7Qi0x9_2),.dout(w_dff_B_SDpKUlTa3_2),.clk(gclk));
	jdff dff_B_NMan6Nod9_2(.din(w_dff_B_SDpKUlTa3_2),.dout(w_dff_B_NMan6Nod9_2),.clk(gclk));
	jdff dff_B_4z1umnXB9_2(.din(w_dff_B_NMan6Nod9_2),.dout(w_dff_B_4z1umnXB9_2),.clk(gclk));
	jdff dff_B_iSTT3HPX3_2(.din(w_dff_B_4z1umnXB9_2),.dout(w_dff_B_iSTT3HPX3_2),.clk(gclk));
	jdff dff_B_7M8AIg5X6_2(.din(w_dff_B_iSTT3HPX3_2),.dout(w_dff_B_7M8AIg5X6_2),.clk(gclk));
	jdff dff_B_LrYpCf1R7_2(.din(w_dff_B_7M8AIg5X6_2),.dout(w_dff_B_LrYpCf1R7_2),.clk(gclk));
	jdff dff_B_YxLPl3QV6_2(.din(w_dff_B_LrYpCf1R7_2),.dout(w_dff_B_YxLPl3QV6_2),.clk(gclk));
	jdff dff_B_8Z78ucoJ0_2(.din(w_dff_B_YxLPl3QV6_2),.dout(w_dff_B_8Z78ucoJ0_2),.clk(gclk));
	jdff dff_B_xnmuVipT2_2(.din(w_dff_B_8Z78ucoJ0_2),.dout(w_dff_B_xnmuVipT2_2),.clk(gclk));
	jdff dff_B_bRI5mEBV4_2(.din(w_dff_B_xnmuVipT2_2),.dout(w_dff_B_bRI5mEBV4_2),.clk(gclk));
	jdff dff_B_besHd5Am9_2(.din(w_dff_B_bRI5mEBV4_2),.dout(w_dff_B_besHd5Am9_2),.clk(gclk));
	jdff dff_B_4kyFvT3S1_2(.din(w_dff_B_besHd5Am9_2),.dout(w_dff_B_4kyFvT3S1_2),.clk(gclk));
	jdff dff_B_v1DaeGCN4_2(.din(w_dff_B_4kyFvT3S1_2),.dout(w_dff_B_v1DaeGCN4_2),.clk(gclk));
	jdff dff_B_BgMvkOkL8_2(.din(w_dff_B_v1DaeGCN4_2),.dout(w_dff_B_BgMvkOkL8_2),.clk(gclk));
	jdff dff_B_4X0pw1Rd1_2(.din(w_dff_B_BgMvkOkL8_2),.dout(w_dff_B_4X0pw1Rd1_2),.clk(gclk));
	jdff dff_B_ULUn1tQD4_2(.din(w_dff_B_4X0pw1Rd1_2),.dout(w_dff_B_ULUn1tQD4_2),.clk(gclk));
	jdff dff_B_DOpKtcWe7_2(.din(w_dff_B_ULUn1tQD4_2),.dout(w_dff_B_DOpKtcWe7_2),.clk(gclk));
	jdff dff_B_fKbJoKPM1_2(.din(w_dff_B_DOpKtcWe7_2),.dout(w_dff_B_fKbJoKPM1_2),.clk(gclk));
	jdff dff_B_6bFjw2Xa8_2(.din(w_dff_B_fKbJoKPM1_2),.dout(w_dff_B_6bFjw2Xa8_2),.clk(gclk));
	jdff dff_B_2HGFSGuf0_2(.din(w_dff_B_6bFjw2Xa8_2),.dout(w_dff_B_2HGFSGuf0_2),.clk(gclk));
	jdff dff_B_SGwdY6Qc1_2(.din(n1615),.dout(w_dff_B_SGwdY6Qc1_2),.clk(gclk));
	jdff dff_B_xWWDbt2V5_1(.din(n1613),.dout(w_dff_B_xWWDbt2V5_1),.clk(gclk));
	jdff dff_B_Zp9VLfbf2_2(.din(n1555),.dout(w_dff_B_Zp9VLfbf2_2),.clk(gclk));
	jdff dff_B_EFB1uhlB4_2(.din(w_dff_B_Zp9VLfbf2_2),.dout(w_dff_B_EFB1uhlB4_2),.clk(gclk));
	jdff dff_B_KkAXeElX0_2(.din(w_dff_B_EFB1uhlB4_2),.dout(w_dff_B_KkAXeElX0_2),.clk(gclk));
	jdff dff_B_pBU7uFsR5_2(.din(w_dff_B_KkAXeElX0_2),.dout(w_dff_B_pBU7uFsR5_2),.clk(gclk));
	jdff dff_B_xrXG658n7_2(.din(w_dff_B_pBU7uFsR5_2),.dout(w_dff_B_xrXG658n7_2),.clk(gclk));
	jdff dff_B_QQus0tLD1_2(.din(w_dff_B_xrXG658n7_2),.dout(w_dff_B_QQus0tLD1_2),.clk(gclk));
	jdff dff_B_i890ZlbO2_2(.din(w_dff_B_QQus0tLD1_2),.dout(w_dff_B_i890ZlbO2_2),.clk(gclk));
	jdff dff_B_1ei6fAKW2_2(.din(w_dff_B_i890ZlbO2_2),.dout(w_dff_B_1ei6fAKW2_2),.clk(gclk));
	jdff dff_B_lPb9NTqD9_2(.din(w_dff_B_1ei6fAKW2_2),.dout(w_dff_B_lPb9NTqD9_2),.clk(gclk));
	jdff dff_B_r3JIv25B6_2(.din(w_dff_B_lPb9NTqD9_2),.dout(w_dff_B_r3JIv25B6_2),.clk(gclk));
	jdff dff_B_MI18Tut26_2(.din(w_dff_B_r3JIv25B6_2),.dout(w_dff_B_MI18Tut26_2),.clk(gclk));
	jdff dff_B_vTAunJB51_2(.din(w_dff_B_MI18Tut26_2),.dout(w_dff_B_vTAunJB51_2),.clk(gclk));
	jdff dff_B_Nh55hMhd8_2(.din(w_dff_B_vTAunJB51_2),.dout(w_dff_B_Nh55hMhd8_2),.clk(gclk));
	jdff dff_B_gMfX8drS2_2(.din(w_dff_B_Nh55hMhd8_2),.dout(w_dff_B_gMfX8drS2_2),.clk(gclk));
	jdff dff_B_Sgw1XGVD3_2(.din(w_dff_B_gMfX8drS2_2),.dout(w_dff_B_Sgw1XGVD3_2),.clk(gclk));
	jdff dff_B_zjpAOmYz5_2(.din(w_dff_B_Sgw1XGVD3_2),.dout(w_dff_B_zjpAOmYz5_2),.clk(gclk));
	jdff dff_B_zKk2AQBO1_2(.din(w_dff_B_zjpAOmYz5_2),.dout(w_dff_B_zKk2AQBO1_2),.clk(gclk));
	jdff dff_B_cl1IGK2H5_2(.din(w_dff_B_zKk2AQBO1_2),.dout(w_dff_B_cl1IGK2H5_2),.clk(gclk));
	jdff dff_B_rFyzzYzX9_2(.din(w_dff_B_cl1IGK2H5_2),.dout(w_dff_B_rFyzzYzX9_2),.clk(gclk));
	jdff dff_B_QEKXQ2at1_2(.din(w_dff_B_rFyzzYzX9_2),.dout(w_dff_B_QEKXQ2at1_2),.clk(gclk));
	jdff dff_B_ihq9HTqP9_2(.din(w_dff_B_QEKXQ2at1_2),.dout(w_dff_B_ihq9HTqP9_2),.clk(gclk));
	jdff dff_B_6dK7vAi15_2(.din(w_dff_B_ihq9HTqP9_2),.dout(w_dff_B_6dK7vAi15_2),.clk(gclk));
	jdff dff_B_pTUQEWkH4_2(.din(w_dff_B_6dK7vAi15_2),.dout(w_dff_B_pTUQEWkH4_2),.clk(gclk));
	jdff dff_B_JZ6jfiZk7_2(.din(w_dff_B_pTUQEWkH4_2),.dout(w_dff_B_JZ6jfiZk7_2),.clk(gclk));
	jdff dff_B_p474wezT6_2(.din(w_dff_B_JZ6jfiZk7_2),.dout(w_dff_B_p474wezT6_2),.clk(gclk));
	jdff dff_B_nJTIuJgD8_2(.din(w_dff_B_p474wezT6_2),.dout(w_dff_B_nJTIuJgD8_2),.clk(gclk));
	jdff dff_B_jJSpxOIK5_2(.din(w_dff_B_nJTIuJgD8_2),.dout(w_dff_B_jJSpxOIK5_2),.clk(gclk));
	jdff dff_B_CDoZxnYN5_2(.din(n1558),.dout(w_dff_B_CDoZxnYN5_2),.clk(gclk));
	jdff dff_B_KSa9u7fX3_1(.din(n1556),.dout(w_dff_B_KSa9u7fX3_1),.clk(gclk));
	jdff dff_B_O8ThttuR1_2(.din(n1491),.dout(w_dff_B_O8ThttuR1_2),.clk(gclk));
	jdff dff_B_8XbVtm7M3_2(.din(w_dff_B_O8ThttuR1_2),.dout(w_dff_B_8XbVtm7M3_2),.clk(gclk));
	jdff dff_B_bz3kgK1s9_2(.din(w_dff_B_8XbVtm7M3_2),.dout(w_dff_B_bz3kgK1s9_2),.clk(gclk));
	jdff dff_B_g3m4722u4_2(.din(w_dff_B_bz3kgK1s9_2),.dout(w_dff_B_g3m4722u4_2),.clk(gclk));
	jdff dff_B_C6JHwCTn4_2(.din(w_dff_B_g3m4722u4_2),.dout(w_dff_B_C6JHwCTn4_2),.clk(gclk));
	jdff dff_B_zQknoiDg3_2(.din(w_dff_B_C6JHwCTn4_2),.dout(w_dff_B_zQknoiDg3_2),.clk(gclk));
	jdff dff_B_cjrwAAy16_2(.din(w_dff_B_zQknoiDg3_2),.dout(w_dff_B_cjrwAAy16_2),.clk(gclk));
	jdff dff_B_ZT48QORD5_2(.din(w_dff_B_cjrwAAy16_2),.dout(w_dff_B_ZT48QORD5_2),.clk(gclk));
	jdff dff_B_9TRrKChU2_2(.din(w_dff_B_ZT48QORD5_2),.dout(w_dff_B_9TRrKChU2_2),.clk(gclk));
	jdff dff_B_rF5I3jvX1_2(.din(w_dff_B_9TRrKChU2_2),.dout(w_dff_B_rF5I3jvX1_2),.clk(gclk));
	jdff dff_B_6fjpsBzQ9_2(.din(w_dff_B_rF5I3jvX1_2),.dout(w_dff_B_6fjpsBzQ9_2),.clk(gclk));
	jdff dff_B_pF2QIoLs7_2(.din(w_dff_B_6fjpsBzQ9_2),.dout(w_dff_B_pF2QIoLs7_2),.clk(gclk));
	jdff dff_B_hkB3C7qP2_2(.din(w_dff_B_pF2QIoLs7_2),.dout(w_dff_B_hkB3C7qP2_2),.clk(gclk));
	jdff dff_B_srW537b57_2(.din(w_dff_B_hkB3C7qP2_2),.dout(w_dff_B_srW537b57_2),.clk(gclk));
	jdff dff_B_THWA969h0_2(.din(w_dff_B_srW537b57_2),.dout(w_dff_B_THWA969h0_2),.clk(gclk));
	jdff dff_B_eUIPKQ0i5_2(.din(w_dff_B_THWA969h0_2),.dout(w_dff_B_eUIPKQ0i5_2),.clk(gclk));
	jdff dff_B_ZOnrIuSA9_2(.din(w_dff_B_eUIPKQ0i5_2),.dout(w_dff_B_ZOnrIuSA9_2),.clk(gclk));
	jdff dff_B_s2c5LKeV8_2(.din(w_dff_B_ZOnrIuSA9_2),.dout(w_dff_B_s2c5LKeV8_2),.clk(gclk));
	jdff dff_B_MVLQcRJq6_2(.din(w_dff_B_s2c5LKeV8_2),.dout(w_dff_B_MVLQcRJq6_2),.clk(gclk));
	jdff dff_B_0fmovR7g5_2(.din(w_dff_B_MVLQcRJq6_2),.dout(w_dff_B_0fmovR7g5_2),.clk(gclk));
	jdff dff_B_rQgWs4YS9_2(.din(w_dff_B_0fmovR7g5_2),.dout(w_dff_B_rQgWs4YS9_2),.clk(gclk));
	jdff dff_B_M5ubFsHp0_2(.din(w_dff_B_rQgWs4YS9_2),.dout(w_dff_B_M5ubFsHp0_2),.clk(gclk));
	jdff dff_B_QTETNQ1u7_2(.din(w_dff_B_M5ubFsHp0_2),.dout(w_dff_B_QTETNQ1u7_2),.clk(gclk));
	jdff dff_B_7bG69QOm0_2(.din(w_dff_B_QTETNQ1u7_2),.dout(w_dff_B_7bG69QOm0_2),.clk(gclk));
	jdff dff_B_E7UOXUYz1_2(.din(n1494),.dout(w_dff_B_E7UOXUYz1_2),.clk(gclk));
	jdff dff_B_ilQTpZAI4_1(.din(n1492),.dout(w_dff_B_ilQTpZAI4_1),.clk(gclk));
	jdff dff_B_J3V8lbAN1_2(.din(n1420),.dout(w_dff_B_J3V8lbAN1_2),.clk(gclk));
	jdff dff_B_Z2z1x4vr0_2(.din(w_dff_B_J3V8lbAN1_2),.dout(w_dff_B_Z2z1x4vr0_2),.clk(gclk));
	jdff dff_B_i5fCaT5J1_2(.din(w_dff_B_Z2z1x4vr0_2),.dout(w_dff_B_i5fCaT5J1_2),.clk(gclk));
	jdff dff_B_537e7v9Z6_2(.din(w_dff_B_i5fCaT5J1_2),.dout(w_dff_B_537e7v9Z6_2),.clk(gclk));
	jdff dff_B_RVQwdxHp4_2(.din(w_dff_B_537e7v9Z6_2),.dout(w_dff_B_RVQwdxHp4_2),.clk(gclk));
	jdff dff_B_kknwGhY53_2(.din(w_dff_B_RVQwdxHp4_2),.dout(w_dff_B_kknwGhY53_2),.clk(gclk));
	jdff dff_B_3UdbeDpG4_2(.din(w_dff_B_kknwGhY53_2),.dout(w_dff_B_3UdbeDpG4_2),.clk(gclk));
	jdff dff_B_0RqoV7tA2_2(.din(w_dff_B_3UdbeDpG4_2),.dout(w_dff_B_0RqoV7tA2_2),.clk(gclk));
	jdff dff_B_wRyfyGmV4_2(.din(w_dff_B_0RqoV7tA2_2),.dout(w_dff_B_wRyfyGmV4_2),.clk(gclk));
	jdff dff_B_MnPY1HCi9_2(.din(w_dff_B_wRyfyGmV4_2),.dout(w_dff_B_MnPY1HCi9_2),.clk(gclk));
	jdff dff_B_ZK6VhDlA9_2(.din(w_dff_B_MnPY1HCi9_2),.dout(w_dff_B_ZK6VhDlA9_2),.clk(gclk));
	jdff dff_B_8Seups0i3_2(.din(w_dff_B_ZK6VhDlA9_2),.dout(w_dff_B_8Seups0i3_2),.clk(gclk));
	jdff dff_B_biwGiqmq8_2(.din(w_dff_B_8Seups0i3_2),.dout(w_dff_B_biwGiqmq8_2),.clk(gclk));
	jdff dff_B_UqoCI8AX2_2(.din(w_dff_B_biwGiqmq8_2),.dout(w_dff_B_UqoCI8AX2_2),.clk(gclk));
	jdff dff_B_7PIRpC1j4_2(.din(w_dff_B_UqoCI8AX2_2),.dout(w_dff_B_7PIRpC1j4_2),.clk(gclk));
	jdff dff_B_GOkLcsT80_2(.din(w_dff_B_7PIRpC1j4_2),.dout(w_dff_B_GOkLcsT80_2),.clk(gclk));
	jdff dff_B_UMCmhLl18_2(.din(w_dff_B_GOkLcsT80_2),.dout(w_dff_B_UMCmhLl18_2),.clk(gclk));
	jdff dff_B_yXv9mCPT4_2(.din(w_dff_B_UMCmhLl18_2),.dout(w_dff_B_yXv9mCPT4_2),.clk(gclk));
	jdff dff_B_zBUICERP7_2(.din(w_dff_B_yXv9mCPT4_2),.dout(w_dff_B_zBUICERP7_2),.clk(gclk));
	jdff dff_B_Jue8yMXR6_2(.din(w_dff_B_zBUICERP7_2),.dout(w_dff_B_Jue8yMXR6_2),.clk(gclk));
	jdff dff_B_0BpSd3x59_2(.din(w_dff_B_Jue8yMXR6_2),.dout(w_dff_B_0BpSd3x59_2),.clk(gclk));
	jdff dff_B_3ylLCC6d3_2(.din(n1423),.dout(w_dff_B_3ylLCC6d3_2),.clk(gclk));
	jdff dff_B_TabAGmhm9_1(.din(n1421),.dout(w_dff_B_TabAGmhm9_1),.clk(gclk));
	jdff dff_B_tgXSQCd49_2(.din(n1342),.dout(w_dff_B_tgXSQCd49_2),.clk(gclk));
	jdff dff_B_OGGaluAV7_2(.din(w_dff_B_tgXSQCd49_2),.dout(w_dff_B_OGGaluAV7_2),.clk(gclk));
	jdff dff_B_cQaYg52C4_2(.din(w_dff_B_OGGaluAV7_2),.dout(w_dff_B_cQaYg52C4_2),.clk(gclk));
	jdff dff_B_08lXtpOw3_2(.din(w_dff_B_cQaYg52C4_2),.dout(w_dff_B_08lXtpOw3_2),.clk(gclk));
	jdff dff_B_lYuarRKj4_2(.din(w_dff_B_08lXtpOw3_2),.dout(w_dff_B_lYuarRKj4_2),.clk(gclk));
	jdff dff_B_snQFI0HS7_2(.din(w_dff_B_lYuarRKj4_2),.dout(w_dff_B_snQFI0HS7_2),.clk(gclk));
	jdff dff_B_EJGpQEYm5_2(.din(w_dff_B_snQFI0HS7_2),.dout(w_dff_B_EJGpQEYm5_2),.clk(gclk));
	jdff dff_B_22UR10zD0_2(.din(w_dff_B_EJGpQEYm5_2),.dout(w_dff_B_22UR10zD0_2),.clk(gclk));
	jdff dff_B_uq4tktCi1_2(.din(w_dff_B_22UR10zD0_2),.dout(w_dff_B_uq4tktCi1_2),.clk(gclk));
	jdff dff_B_5KA9qhZd1_2(.din(w_dff_B_uq4tktCi1_2),.dout(w_dff_B_5KA9qhZd1_2),.clk(gclk));
	jdff dff_B_GyAEtiNK3_2(.din(w_dff_B_5KA9qhZd1_2),.dout(w_dff_B_GyAEtiNK3_2),.clk(gclk));
	jdff dff_B_v8zYFRii9_2(.din(w_dff_B_GyAEtiNK3_2),.dout(w_dff_B_v8zYFRii9_2),.clk(gclk));
	jdff dff_B_vc9RdmFB7_2(.din(w_dff_B_v8zYFRii9_2),.dout(w_dff_B_vc9RdmFB7_2),.clk(gclk));
	jdff dff_B_4L7LbXtC4_2(.din(w_dff_B_vc9RdmFB7_2),.dout(w_dff_B_4L7LbXtC4_2),.clk(gclk));
	jdff dff_B_w3VKHJfC4_2(.din(w_dff_B_4L7LbXtC4_2),.dout(w_dff_B_w3VKHJfC4_2),.clk(gclk));
	jdff dff_B_OfHnQNTx9_2(.din(w_dff_B_w3VKHJfC4_2),.dout(w_dff_B_OfHnQNTx9_2),.clk(gclk));
	jdff dff_B_ONsQwoUF5_2(.din(w_dff_B_OfHnQNTx9_2),.dout(w_dff_B_ONsQwoUF5_2),.clk(gclk));
	jdff dff_B_ICXqUIyS3_2(.din(w_dff_B_ONsQwoUF5_2),.dout(w_dff_B_ICXqUIyS3_2),.clk(gclk));
	jdff dff_B_13lUOBpt4_1(.din(n1343),.dout(w_dff_B_13lUOBpt4_1),.clk(gclk));
	jdff dff_B_XE8Zla7A7_2(.din(n1257),.dout(w_dff_B_XE8Zla7A7_2),.clk(gclk));
	jdff dff_B_GBagAQh26_2(.din(w_dff_B_XE8Zla7A7_2),.dout(w_dff_B_GBagAQh26_2),.clk(gclk));
	jdff dff_B_W7beV2HV7_2(.din(w_dff_B_GBagAQh26_2),.dout(w_dff_B_W7beV2HV7_2),.clk(gclk));
	jdff dff_B_3O8S6Rkd9_2(.din(w_dff_B_W7beV2HV7_2),.dout(w_dff_B_3O8S6Rkd9_2),.clk(gclk));
	jdff dff_B_RjHMUA5g0_2(.din(w_dff_B_3O8S6Rkd9_2),.dout(w_dff_B_RjHMUA5g0_2),.clk(gclk));
	jdff dff_B_hkkAbBA62_2(.din(w_dff_B_RjHMUA5g0_2),.dout(w_dff_B_hkkAbBA62_2),.clk(gclk));
	jdff dff_B_ds5nAQBH6_2(.din(w_dff_B_hkkAbBA62_2),.dout(w_dff_B_ds5nAQBH6_2),.clk(gclk));
	jdff dff_B_osjiGzTg8_2(.din(w_dff_B_ds5nAQBH6_2),.dout(w_dff_B_osjiGzTg8_2),.clk(gclk));
	jdff dff_B_AjtwBvk20_2(.din(w_dff_B_osjiGzTg8_2),.dout(w_dff_B_AjtwBvk20_2),.clk(gclk));
	jdff dff_B_LgQc05j61_2(.din(w_dff_B_AjtwBvk20_2),.dout(w_dff_B_LgQc05j61_2),.clk(gclk));
	jdff dff_B_K5V3l6oe5_2(.din(w_dff_B_LgQc05j61_2),.dout(w_dff_B_K5V3l6oe5_2),.clk(gclk));
	jdff dff_B_jUhFgxou5_2(.din(w_dff_B_K5V3l6oe5_2),.dout(w_dff_B_jUhFgxou5_2),.clk(gclk));
	jdff dff_B_HPAt1UAq8_2(.din(w_dff_B_jUhFgxou5_2),.dout(w_dff_B_HPAt1UAq8_2),.clk(gclk));
	jdff dff_B_jWGxNwRn9_2(.din(w_dff_B_HPAt1UAq8_2),.dout(w_dff_B_jWGxNwRn9_2),.clk(gclk));
	jdff dff_B_IhcHGSeE9_2(.din(w_dff_B_jWGxNwRn9_2),.dout(w_dff_B_IhcHGSeE9_2),.clk(gclk));
	jdff dff_B_cUJKJhQb6_2(.din(w_dff_B_IhcHGSeE9_2),.dout(w_dff_B_cUJKJhQb6_2),.clk(gclk));
	jdff dff_B_le5ggeC59_2(.din(n1275),.dout(w_dff_B_le5ggeC59_2),.clk(gclk));
	jdff dff_B_rX2mSMAu1_1(.din(n1258),.dout(w_dff_B_rX2mSMAu1_1),.clk(gclk));
	jdff dff_B_OBXm2lG17_2(.din(n1166),.dout(w_dff_B_OBXm2lG17_2),.clk(gclk));
	jdff dff_B_1y6ZNWQn9_2(.din(w_dff_B_OBXm2lG17_2),.dout(w_dff_B_1y6ZNWQn9_2),.clk(gclk));
	jdff dff_B_TvRm66R32_2(.din(w_dff_B_1y6ZNWQn9_2),.dout(w_dff_B_TvRm66R32_2),.clk(gclk));
	jdff dff_B_ZPw5bUAJ7_2(.din(w_dff_B_TvRm66R32_2),.dout(w_dff_B_ZPw5bUAJ7_2),.clk(gclk));
	jdff dff_B_SwwY8paL8_2(.din(w_dff_B_ZPw5bUAJ7_2),.dout(w_dff_B_SwwY8paL8_2),.clk(gclk));
	jdff dff_B_MvsfIHOT3_2(.din(w_dff_B_SwwY8paL8_2),.dout(w_dff_B_MvsfIHOT3_2),.clk(gclk));
	jdff dff_B_HnuoiPBJ9_2(.din(w_dff_B_MvsfIHOT3_2),.dout(w_dff_B_HnuoiPBJ9_2),.clk(gclk));
	jdff dff_B_LqlLr0Gf2_2(.din(w_dff_B_HnuoiPBJ9_2),.dout(w_dff_B_LqlLr0Gf2_2),.clk(gclk));
	jdff dff_B_7uAjTiH48_2(.din(w_dff_B_LqlLr0Gf2_2),.dout(w_dff_B_7uAjTiH48_2),.clk(gclk));
	jdff dff_B_Asfhe3Xj1_2(.din(w_dff_B_7uAjTiH48_2),.dout(w_dff_B_Asfhe3Xj1_2),.clk(gclk));
	jdff dff_B_iYfvHzZn4_2(.din(w_dff_B_Asfhe3Xj1_2),.dout(w_dff_B_iYfvHzZn4_2),.clk(gclk));
	jdff dff_B_8xwOzDuu7_2(.din(w_dff_B_iYfvHzZn4_2),.dout(w_dff_B_8xwOzDuu7_2),.clk(gclk));
	jdff dff_B_S75SklB48_2(.din(w_dff_B_8xwOzDuu7_2),.dout(w_dff_B_S75SklB48_2),.clk(gclk));
	jdff dff_B_SVEDSDEi2_2(.din(w_dff_B_S75SklB48_2),.dout(w_dff_B_SVEDSDEi2_2),.clk(gclk));
	jdff dff_B_B4HWDCRE2_2(.din(n1184),.dout(w_dff_B_B4HWDCRE2_2),.clk(gclk));
	jdff dff_B_GZxrntJy9_1(.din(n1167),.dout(w_dff_B_GZxrntJy9_1),.clk(gclk));
	jdff dff_B_Nt7NuWTH8_2(.din(n1068),.dout(w_dff_B_Nt7NuWTH8_2),.clk(gclk));
	jdff dff_B_2cQPzvWm4_2(.din(w_dff_B_Nt7NuWTH8_2),.dout(w_dff_B_2cQPzvWm4_2),.clk(gclk));
	jdff dff_B_2wTKKPzC0_2(.din(w_dff_B_2cQPzvWm4_2),.dout(w_dff_B_2wTKKPzC0_2),.clk(gclk));
	jdff dff_B_9catRUxp6_2(.din(w_dff_B_2wTKKPzC0_2),.dout(w_dff_B_9catRUxp6_2),.clk(gclk));
	jdff dff_B_pVensoYy4_2(.din(w_dff_B_9catRUxp6_2),.dout(w_dff_B_pVensoYy4_2),.clk(gclk));
	jdff dff_B_xRkTMFIC1_2(.din(w_dff_B_pVensoYy4_2),.dout(w_dff_B_xRkTMFIC1_2),.clk(gclk));
	jdff dff_B_wY2vCz325_2(.din(w_dff_B_xRkTMFIC1_2),.dout(w_dff_B_wY2vCz325_2),.clk(gclk));
	jdff dff_B_lJDYlO5t0_2(.din(w_dff_B_wY2vCz325_2),.dout(w_dff_B_lJDYlO5t0_2),.clk(gclk));
	jdff dff_B_JXXs8xIx6_2(.din(w_dff_B_lJDYlO5t0_2),.dout(w_dff_B_JXXs8xIx6_2),.clk(gclk));
	jdff dff_B_Ims85ujk8_2(.din(w_dff_B_JXXs8xIx6_2),.dout(w_dff_B_Ims85ujk8_2),.clk(gclk));
	jdff dff_B_RK6kbfCp8_2(.din(w_dff_B_Ims85ujk8_2),.dout(w_dff_B_RK6kbfCp8_2),.clk(gclk));
	jdff dff_B_pMPuw8w75_2(.din(w_dff_B_RK6kbfCp8_2),.dout(w_dff_B_pMPuw8w75_2),.clk(gclk));
	jdff dff_B_YzE7vhIp1_2(.din(n1085),.dout(w_dff_B_YzE7vhIp1_2),.clk(gclk));
	jdff dff_B_fBGJNpeL5_1(.din(n1069),.dout(w_dff_B_fBGJNpeL5_1),.clk(gclk));
	jdff dff_B_e2Java6M1_2(.din(n969),.dout(w_dff_B_e2Java6M1_2),.clk(gclk));
	jdff dff_B_Yk9pl2oQ3_2(.din(w_dff_B_e2Java6M1_2),.dout(w_dff_B_Yk9pl2oQ3_2),.clk(gclk));
	jdff dff_B_k3JCi18x8_2(.din(w_dff_B_Yk9pl2oQ3_2),.dout(w_dff_B_k3JCi18x8_2),.clk(gclk));
	jdff dff_B_qozo7iat7_2(.din(w_dff_B_k3JCi18x8_2),.dout(w_dff_B_qozo7iat7_2),.clk(gclk));
	jdff dff_B_jEzkYGKY5_2(.din(w_dff_B_qozo7iat7_2),.dout(w_dff_B_jEzkYGKY5_2),.clk(gclk));
	jdff dff_B_FNNG2QIv1_2(.din(w_dff_B_jEzkYGKY5_2),.dout(w_dff_B_FNNG2QIv1_2),.clk(gclk));
	jdff dff_B_twRhjcnr3_2(.din(w_dff_B_FNNG2QIv1_2),.dout(w_dff_B_twRhjcnr3_2),.clk(gclk));
	jdff dff_B_KphbzRRW0_2(.din(w_dff_B_twRhjcnr3_2),.dout(w_dff_B_KphbzRRW0_2),.clk(gclk));
	jdff dff_B_OZt0q0Bx8_2(.din(w_dff_B_KphbzRRW0_2),.dout(w_dff_B_OZt0q0Bx8_2),.clk(gclk));
	jdff dff_B_uWR791Wt7_2(.din(w_dff_B_OZt0q0Bx8_2),.dout(w_dff_B_uWR791Wt7_2),.clk(gclk));
	jdff dff_B_biMF5xiY2_2(.din(n986),.dout(w_dff_B_biMF5xiY2_2),.clk(gclk));
	jdff dff_B_Qy0Xl20H1_1(.din(n970),.dout(w_dff_B_Qy0Xl20H1_1),.clk(gclk));
	jdff dff_B_IprDgkyj1_2(.din(n867),.dout(w_dff_B_IprDgkyj1_2),.clk(gclk));
	jdff dff_B_6R4J12MB3_2(.din(w_dff_B_IprDgkyj1_2),.dout(w_dff_B_6R4J12MB3_2),.clk(gclk));
	jdff dff_B_orbJmY5M4_2(.din(w_dff_B_6R4J12MB3_2),.dout(w_dff_B_orbJmY5M4_2),.clk(gclk));
	jdff dff_B_VRh20Rzh3_2(.din(w_dff_B_orbJmY5M4_2),.dout(w_dff_B_VRh20Rzh3_2),.clk(gclk));
	jdff dff_B_RLopCCLL3_2(.din(w_dff_B_VRh20Rzh3_2),.dout(w_dff_B_RLopCCLL3_2),.clk(gclk));
	jdff dff_B_Ne3ft27P3_2(.din(w_dff_B_RLopCCLL3_2),.dout(w_dff_B_Ne3ft27P3_2),.clk(gclk));
	jdff dff_B_p49DaM4y5_2(.din(w_dff_B_Ne3ft27P3_2),.dout(w_dff_B_p49DaM4y5_2),.clk(gclk));
	jdff dff_B_rnVyKTkM6_2(.din(w_dff_B_p49DaM4y5_2),.dout(w_dff_B_rnVyKTkM6_2),.clk(gclk));
	jdff dff_B_xOc774nP5_2(.din(n880),.dout(w_dff_B_xOc774nP5_2),.clk(gclk));
	jdff dff_B_qpgK7ctZ7_2(.din(w_dff_B_xOc774nP5_2),.dout(w_dff_B_qpgK7ctZ7_2),.clk(gclk));
	jdff dff_B_D84DGjHM1_2(.din(w_dff_B_qpgK7ctZ7_2),.dout(w_dff_B_D84DGjHM1_2),.clk(gclk));
	jdff dff_B_LAz1Hdqf1_2(.din(w_dff_B_D84DGjHM1_2),.dout(w_dff_B_LAz1Hdqf1_2),.clk(gclk));
	jdff dff_B_N0vnEraq2_1(.din(n868),.dout(w_dff_B_N0vnEraq2_1),.clk(gclk));
	jdff dff_B_nZWTWXa57_1(.din(w_dff_B_N0vnEraq2_1),.dout(w_dff_B_nZWTWXa57_1),.clk(gclk));
	jdff dff_B_7msUnWsI5_1(.din(w_dff_B_nZWTWXa57_1),.dout(w_dff_B_7msUnWsI5_1),.clk(gclk));
	jdff dff_B_n8ACra2z8_2(.din(n771),.dout(w_dff_B_n8ACra2z8_2),.clk(gclk));
	jdff dff_B_UGgeFQ3J6_2(.din(w_dff_B_n8ACra2z8_2),.dout(w_dff_B_UGgeFQ3J6_2),.clk(gclk));
	jdff dff_B_M7dKjfdi0_2(.din(w_dff_B_UGgeFQ3J6_2),.dout(w_dff_B_M7dKjfdi0_2),.clk(gclk));
	jdff dff_B_KltZ9xIm0_0(.din(n776),.dout(w_dff_B_KltZ9xIm0_0),.clk(gclk));
	jdff dff_B_xvpOpkG77_0(.din(w_dff_B_KltZ9xIm0_0),.dout(w_dff_B_xvpOpkG77_0),.clk(gclk));
	jdff dff_A_hsF3NyvZ2_0(.dout(w_n676_0[0]),.din(w_dff_A_hsF3NyvZ2_0),.clk(gclk));
	jdff dff_A_uEHtC4hr1_0(.dout(w_dff_A_hsF3NyvZ2_0),.din(w_dff_A_uEHtC4hr1_0),.clk(gclk));
	jdff dff_A_kP1gabiN5_1(.dout(w_n676_0[1]),.din(w_dff_A_kP1gabiN5_1),.clk(gclk));
	jdff dff_A_7ZLP7fsA9_1(.dout(w_dff_A_kP1gabiN5_1),.din(w_dff_A_7ZLP7fsA9_1),.clk(gclk));
	jdff dff_B_uCql4FRT2_1(.din(n1812),.dout(w_dff_B_uCql4FRT2_1),.clk(gclk));
	jdff dff_B_rl9vlxdI6_1(.din(n1799),.dout(w_dff_B_rl9vlxdI6_1),.clk(gclk));
	jdff dff_B_CF2m4dVa4_1(.din(w_dff_B_rl9vlxdI6_1),.dout(w_dff_B_CF2m4dVa4_1),.clk(gclk));
	jdff dff_B_nEFS87Ai0_2(.din(n1798),.dout(w_dff_B_nEFS87Ai0_2),.clk(gclk));
	jdff dff_B_QIbqq9Zi8_2(.din(w_dff_B_nEFS87Ai0_2),.dout(w_dff_B_QIbqq9Zi8_2),.clk(gclk));
	jdff dff_B_Anu3fJEK1_2(.din(w_dff_B_QIbqq9Zi8_2),.dout(w_dff_B_Anu3fJEK1_2),.clk(gclk));
	jdff dff_B_Ivpi194A6_2(.din(w_dff_B_Anu3fJEK1_2),.dout(w_dff_B_Ivpi194A6_2),.clk(gclk));
	jdff dff_B_wSeg0Sqm7_2(.din(w_dff_B_Ivpi194A6_2),.dout(w_dff_B_wSeg0Sqm7_2),.clk(gclk));
	jdff dff_B_q9zeoEoj4_2(.din(w_dff_B_wSeg0Sqm7_2),.dout(w_dff_B_q9zeoEoj4_2),.clk(gclk));
	jdff dff_B_NM9Z7tEL3_2(.din(w_dff_B_q9zeoEoj4_2),.dout(w_dff_B_NM9Z7tEL3_2),.clk(gclk));
	jdff dff_B_21PDXfCs1_2(.din(w_dff_B_NM9Z7tEL3_2),.dout(w_dff_B_21PDXfCs1_2),.clk(gclk));
	jdff dff_B_MS6ma5TJ0_2(.din(w_dff_B_21PDXfCs1_2),.dout(w_dff_B_MS6ma5TJ0_2),.clk(gclk));
	jdff dff_B_cWTYRXaf0_2(.din(w_dff_B_MS6ma5TJ0_2),.dout(w_dff_B_cWTYRXaf0_2),.clk(gclk));
	jdff dff_B_edylnqdb4_2(.din(w_dff_B_cWTYRXaf0_2),.dout(w_dff_B_edylnqdb4_2),.clk(gclk));
	jdff dff_B_LONx44nf7_2(.din(w_dff_B_edylnqdb4_2),.dout(w_dff_B_LONx44nf7_2),.clk(gclk));
	jdff dff_B_RoR94wHC6_2(.din(w_dff_B_LONx44nf7_2),.dout(w_dff_B_RoR94wHC6_2),.clk(gclk));
	jdff dff_B_RIHJWEMA6_2(.din(w_dff_B_RoR94wHC6_2),.dout(w_dff_B_RIHJWEMA6_2),.clk(gclk));
	jdff dff_B_p6Z4JQWe1_2(.din(w_dff_B_RIHJWEMA6_2),.dout(w_dff_B_p6Z4JQWe1_2),.clk(gclk));
	jdff dff_B_OuVLpQXI4_2(.din(w_dff_B_p6Z4JQWe1_2),.dout(w_dff_B_OuVLpQXI4_2),.clk(gclk));
	jdff dff_B_gRbTJOSu6_2(.din(w_dff_B_OuVLpQXI4_2),.dout(w_dff_B_gRbTJOSu6_2),.clk(gclk));
	jdff dff_B_QQT2rHBu8_2(.din(w_dff_B_gRbTJOSu6_2),.dout(w_dff_B_QQT2rHBu8_2),.clk(gclk));
	jdff dff_B_G8L7C8to9_2(.din(w_dff_B_QQT2rHBu8_2),.dout(w_dff_B_G8L7C8to9_2),.clk(gclk));
	jdff dff_B_X5lOdO0j9_2(.din(w_dff_B_G8L7C8to9_2),.dout(w_dff_B_X5lOdO0j9_2),.clk(gclk));
	jdff dff_B_U2tAw60L8_2(.din(w_dff_B_X5lOdO0j9_2),.dout(w_dff_B_U2tAw60L8_2),.clk(gclk));
	jdff dff_B_S3SZhNI05_2(.din(w_dff_B_U2tAw60L8_2),.dout(w_dff_B_S3SZhNI05_2),.clk(gclk));
	jdff dff_B_rCREUAou5_2(.din(w_dff_B_S3SZhNI05_2),.dout(w_dff_B_rCREUAou5_2),.clk(gclk));
	jdff dff_B_YVSm7Ifz7_2(.din(w_dff_B_rCREUAou5_2),.dout(w_dff_B_YVSm7Ifz7_2),.clk(gclk));
	jdff dff_B_oeVRQQCS1_2(.din(w_dff_B_YVSm7Ifz7_2),.dout(w_dff_B_oeVRQQCS1_2),.clk(gclk));
	jdff dff_B_ZBBpgqqu1_2(.din(w_dff_B_oeVRQQCS1_2),.dout(w_dff_B_ZBBpgqqu1_2),.clk(gclk));
	jdff dff_B_qqdARr595_2(.din(w_dff_B_ZBBpgqqu1_2),.dout(w_dff_B_qqdARr595_2),.clk(gclk));
	jdff dff_B_GQTXw5KC8_2(.din(w_dff_B_qqdARr595_2),.dout(w_dff_B_GQTXw5KC8_2),.clk(gclk));
	jdff dff_B_TKBP6cBN4_2(.din(w_dff_B_GQTXw5KC8_2),.dout(w_dff_B_TKBP6cBN4_2),.clk(gclk));
	jdff dff_B_mwAC1SRx8_2(.din(w_dff_B_TKBP6cBN4_2),.dout(w_dff_B_mwAC1SRx8_2),.clk(gclk));
	jdff dff_B_8CR8RnnO8_2(.din(w_dff_B_mwAC1SRx8_2),.dout(w_dff_B_8CR8RnnO8_2),.clk(gclk));
	jdff dff_B_ulpok7JF8_2(.din(w_dff_B_8CR8RnnO8_2),.dout(w_dff_B_ulpok7JF8_2),.clk(gclk));
	jdff dff_B_IqacMjtd3_2(.din(w_dff_B_ulpok7JF8_2),.dout(w_dff_B_IqacMjtd3_2),.clk(gclk));
	jdff dff_B_beenyYfC7_2(.din(w_dff_B_IqacMjtd3_2),.dout(w_dff_B_beenyYfC7_2),.clk(gclk));
	jdff dff_B_piiYpN3z0_2(.din(w_dff_B_beenyYfC7_2),.dout(w_dff_B_piiYpN3z0_2),.clk(gclk));
	jdff dff_B_3TSunjsR5_2(.din(w_dff_B_piiYpN3z0_2),.dout(w_dff_B_3TSunjsR5_2),.clk(gclk));
	jdff dff_B_PApem8KO0_2(.din(w_dff_B_3TSunjsR5_2),.dout(w_dff_B_PApem8KO0_2),.clk(gclk));
	jdff dff_B_w8i6ZHGt6_2(.din(w_dff_B_PApem8KO0_2),.dout(w_dff_B_w8i6ZHGt6_2),.clk(gclk));
	jdff dff_B_4rmOztLO7_2(.din(w_dff_B_w8i6ZHGt6_2),.dout(w_dff_B_4rmOztLO7_2),.clk(gclk));
	jdff dff_B_yB2mG7uE0_2(.din(w_dff_B_4rmOztLO7_2),.dout(w_dff_B_yB2mG7uE0_2),.clk(gclk));
	jdff dff_B_x2k9ZlQs4_2(.din(n1797),.dout(w_dff_B_x2k9ZlQs4_2),.clk(gclk));
	jdff dff_B_vRibU5070_2(.din(w_dff_B_x2k9ZlQs4_2),.dout(w_dff_B_vRibU5070_2),.clk(gclk));
	jdff dff_B_l5NVgHt94_2(.din(w_dff_B_vRibU5070_2),.dout(w_dff_B_l5NVgHt94_2),.clk(gclk));
	jdff dff_B_LK7DGMTD3_2(.din(w_dff_B_l5NVgHt94_2),.dout(w_dff_B_LK7DGMTD3_2),.clk(gclk));
	jdff dff_B_Ov1t8lOk6_2(.din(w_dff_B_LK7DGMTD3_2),.dout(w_dff_B_Ov1t8lOk6_2),.clk(gclk));
	jdff dff_B_STCDMDJq9_2(.din(w_dff_B_Ov1t8lOk6_2),.dout(w_dff_B_STCDMDJq9_2),.clk(gclk));
	jdff dff_B_4yY9eZkn0_2(.din(w_dff_B_STCDMDJq9_2),.dout(w_dff_B_4yY9eZkn0_2),.clk(gclk));
	jdff dff_B_3JoAIAof2_2(.din(w_dff_B_4yY9eZkn0_2),.dout(w_dff_B_3JoAIAof2_2),.clk(gclk));
	jdff dff_B_Z22TOUEK3_2(.din(w_dff_B_3JoAIAof2_2),.dout(w_dff_B_Z22TOUEK3_2),.clk(gclk));
	jdff dff_B_TYu2qYXa0_2(.din(w_dff_B_Z22TOUEK3_2),.dout(w_dff_B_TYu2qYXa0_2),.clk(gclk));
	jdff dff_B_otr8tp1c2_2(.din(w_dff_B_TYu2qYXa0_2),.dout(w_dff_B_otr8tp1c2_2),.clk(gclk));
	jdff dff_B_ntKPQsXT6_2(.din(w_dff_B_otr8tp1c2_2),.dout(w_dff_B_ntKPQsXT6_2),.clk(gclk));
	jdff dff_B_KpG2wTF57_2(.din(w_dff_B_ntKPQsXT6_2),.dout(w_dff_B_KpG2wTF57_2),.clk(gclk));
	jdff dff_B_ouQnik5Y5_2(.din(w_dff_B_KpG2wTF57_2),.dout(w_dff_B_ouQnik5Y5_2),.clk(gclk));
	jdff dff_B_67PgEyvu6_2(.din(w_dff_B_ouQnik5Y5_2),.dout(w_dff_B_67PgEyvu6_2),.clk(gclk));
	jdff dff_B_G0W8jHBL3_2(.din(w_dff_B_67PgEyvu6_2),.dout(w_dff_B_G0W8jHBL3_2),.clk(gclk));
	jdff dff_B_Z3cLKKX17_2(.din(w_dff_B_G0W8jHBL3_2),.dout(w_dff_B_Z3cLKKX17_2),.clk(gclk));
	jdff dff_B_gH85watT4_2(.din(w_dff_B_Z3cLKKX17_2),.dout(w_dff_B_gH85watT4_2),.clk(gclk));
	jdff dff_B_y36MB31H5_2(.din(w_dff_B_gH85watT4_2),.dout(w_dff_B_y36MB31H5_2),.clk(gclk));
	jdff dff_B_bPibAl636_2(.din(w_dff_B_y36MB31H5_2),.dout(w_dff_B_bPibAl636_2),.clk(gclk));
	jdff dff_B_d0fz6zrI7_2(.din(w_dff_B_bPibAl636_2),.dout(w_dff_B_d0fz6zrI7_2),.clk(gclk));
	jdff dff_B_zAaED1tm9_2(.din(w_dff_B_d0fz6zrI7_2),.dout(w_dff_B_zAaED1tm9_2),.clk(gclk));
	jdff dff_B_RPMo3dtl2_2(.din(w_dff_B_zAaED1tm9_2),.dout(w_dff_B_RPMo3dtl2_2),.clk(gclk));
	jdff dff_B_IJpghNJq6_2(.din(w_dff_B_RPMo3dtl2_2),.dout(w_dff_B_IJpghNJq6_2),.clk(gclk));
	jdff dff_B_qFQ5aVNJ0_2(.din(w_dff_B_IJpghNJq6_2),.dout(w_dff_B_qFQ5aVNJ0_2),.clk(gclk));
	jdff dff_B_kYQP5fqt3_2(.din(w_dff_B_qFQ5aVNJ0_2),.dout(w_dff_B_kYQP5fqt3_2),.clk(gclk));
	jdff dff_B_wRIcmDHZ4_2(.din(w_dff_B_kYQP5fqt3_2),.dout(w_dff_B_wRIcmDHZ4_2),.clk(gclk));
	jdff dff_B_rlMoE8j13_2(.din(w_dff_B_wRIcmDHZ4_2),.dout(w_dff_B_rlMoE8j13_2),.clk(gclk));
	jdff dff_B_4QJhEaaP6_2(.din(w_dff_B_rlMoE8j13_2),.dout(w_dff_B_4QJhEaaP6_2),.clk(gclk));
	jdff dff_B_gJzLfDV48_2(.din(w_dff_B_4QJhEaaP6_2),.dout(w_dff_B_gJzLfDV48_2),.clk(gclk));
	jdff dff_B_3GpmEY7x0_2(.din(w_dff_B_gJzLfDV48_2),.dout(w_dff_B_3GpmEY7x0_2),.clk(gclk));
	jdff dff_B_fyRqKogp5_2(.din(w_dff_B_3GpmEY7x0_2),.dout(w_dff_B_fyRqKogp5_2),.clk(gclk));
	jdff dff_B_fIuVZdE61_2(.din(w_dff_B_fyRqKogp5_2),.dout(w_dff_B_fIuVZdE61_2),.clk(gclk));
	jdff dff_B_n0RBurjJ1_2(.din(w_dff_B_fIuVZdE61_2),.dout(w_dff_B_n0RBurjJ1_2),.clk(gclk));
	jdff dff_B_630N5O5X1_2(.din(w_dff_B_n0RBurjJ1_2),.dout(w_dff_B_630N5O5X1_2),.clk(gclk));
	jdff dff_B_9f3XXe5K5_2(.din(w_dff_B_630N5O5X1_2),.dout(w_dff_B_9f3XXe5K5_2),.clk(gclk));
	jdff dff_B_vGdWOhNZ3_2(.din(w_dff_B_9f3XXe5K5_2),.dout(w_dff_B_vGdWOhNZ3_2),.clk(gclk));
	jdff dff_B_htZaDNGr6_2(.din(w_dff_B_vGdWOhNZ3_2),.dout(w_dff_B_htZaDNGr6_2),.clk(gclk));
	jdff dff_B_RkC5OAzX7_2(.din(w_dff_B_htZaDNGr6_2),.dout(w_dff_B_RkC5OAzX7_2),.clk(gclk));
	jdff dff_B_1c0MTidD8_2(.din(w_dff_B_RkC5OAzX7_2),.dout(w_dff_B_1c0MTidD8_2),.clk(gclk));
	jdff dff_B_JOhg4HcK6_2(.din(w_dff_B_1c0MTidD8_2),.dout(w_dff_B_JOhg4HcK6_2),.clk(gclk));
	jdff dff_B_MVv0CSar4_2(.din(w_dff_B_JOhg4HcK6_2),.dout(w_dff_B_MVv0CSar4_2),.clk(gclk));
	jdff dff_A_KzNFY41T9_1(.dout(w_n1796_0[1]),.din(w_dff_A_KzNFY41T9_1),.clk(gclk));
	jdff dff_B_Ve2vwywr3_1(.din(n1794),.dout(w_dff_B_Ve2vwywr3_1),.clk(gclk));
	jdff dff_B_qHbWoxwg0_2(.din(n1772),.dout(w_dff_B_qHbWoxwg0_2),.clk(gclk));
	jdff dff_B_f5l68lMe1_2(.din(w_dff_B_qHbWoxwg0_2),.dout(w_dff_B_f5l68lMe1_2),.clk(gclk));
	jdff dff_B_gx3AzOuo8_2(.din(w_dff_B_f5l68lMe1_2),.dout(w_dff_B_gx3AzOuo8_2),.clk(gclk));
	jdff dff_B_ZPxaJen13_2(.din(w_dff_B_gx3AzOuo8_2),.dout(w_dff_B_ZPxaJen13_2),.clk(gclk));
	jdff dff_B_aczEN2C29_2(.din(w_dff_B_ZPxaJen13_2),.dout(w_dff_B_aczEN2C29_2),.clk(gclk));
	jdff dff_B_pPJprndS1_2(.din(w_dff_B_aczEN2C29_2),.dout(w_dff_B_pPJprndS1_2),.clk(gclk));
	jdff dff_B_rZ9Xi93j3_2(.din(w_dff_B_pPJprndS1_2),.dout(w_dff_B_rZ9Xi93j3_2),.clk(gclk));
	jdff dff_B_rvuYyjHg8_2(.din(w_dff_B_rZ9Xi93j3_2),.dout(w_dff_B_rvuYyjHg8_2),.clk(gclk));
	jdff dff_B_0SIpv0ki1_2(.din(w_dff_B_rvuYyjHg8_2),.dout(w_dff_B_0SIpv0ki1_2),.clk(gclk));
	jdff dff_B_KXh5epmY6_2(.din(w_dff_B_0SIpv0ki1_2),.dout(w_dff_B_KXh5epmY6_2),.clk(gclk));
	jdff dff_B_yK5G8RGe3_2(.din(w_dff_B_KXh5epmY6_2),.dout(w_dff_B_yK5G8RGe3_2),.clk(gclk));
	jdff dff_B_xA6472Qr1_2(.din(w_dff_B_yK5G8RGe3_2),.dout(w_dff_B_xA6472Qr1_2),.clk(gclk));
	jdff dff_B_sRlq7t2J1_2(.din(w_dff_B_xA6472Qr1_2),.dout(w_dff_B_sRlq7t2J1_2),.clk(gclk));
	jdff dff_B_Csq2y3z53_2(.din(w_dff_B_sRlq7t2J1_2),.dout(w_dff_B_Csq2y3z53_2),.clk(gclk));
	jdff dff_B_DOFbZy0i6_2(.din(w_dff_B_Csq2y3z53_2),.dout(w_dff_B_DOFbZy0i6_2),.clk(gclk));
	jdff dff_B_rtN0sDRD3_2(.din(w_dff_B_DOFbZy0i6_2),.dout(w_dff_B_rtN0sDRD3_2),.clk(gclk));
	jdff dff_B_WDkQAfWS6_2(.din(w_dff_B_rtN0sDRD3_2),.dout(w_dff_B_WDkQAfWS6_2),.clk(gclk));
	jdff dff_B_qRM52eFs1_2(.din(w_dff_B_WDkQAfWS6_2),.dout(w_dff_B_qRM52eFs1_2),.clk(gclk));
	jdff dff_B_fyAgyzEO8_2(.din(w_dff_B_qRM52eFs1_2),.dout(w_dff_B_fyAgyzEO8_2),.clk(gclk));
	jdff dff_B_XrFIZvxS1_2(.din(w_dff_B_fyAgyzEO8_2),.dout(w_dff_B_XrFIZvxS1_2),.clk(gclk));
	jdff dff_B_FuAHmZEw7_2(.din(w_dff_B_XrFIZvxS1_2),.dout(w_dff_B_FuAHmZEw7_2),.clk(gclk));
	jdff dff_B_KcuMKJBl7_2(.din(w_dff_B_FuAHmZEw7_2),.dout(w_dff_B_KcuMKJBl7_2),.clk(gclk));
	jdff dff_B_ctYcNkls5_2(.din(w_dff_B_KcuMKJBl7_2),.dout(w_dff_B_ctYcNkls5_2),.clk(gclk));
	jdff dff_B_yj77zrbg3_2(.din(w_dff_B_ctYcNkls5_2),.dout(w_dff_B_yj77zrbg3_2),.clk(gclk));
	jdff dff_B_xe8dbRAp8_2(.din(w_dff_B_yj77zrbg3_2),.dout(w_dff_B_xe8dbRAp8_2),.clk(gclk));
	jdff dff_B_pR0pMSR62_2(.din(w_dff_B_xe8dbRAp8_2),.dout(w_dff_B_pR0pMSR62_2),.clk(gclk));
	jdff dff_B_xk5RLVF85_2(.din(w_dff_B_pR0pMSR62_2),.dout(w_dff_B_xk5RLVF85_2),.clk(gclk));
	jdff dff_B_doxSpFA06_2(.din(w_dff_B_xk5RLVF85_2),.dout(w_dff_B_doxSpFA06_2),.clk(gclk));
	jdff dff_B_4xesHF4G0_2(.din(w_dff_B_doxSpFA06_2),.dout(w_dff_B_4xesHF4G0_2),.clk(gclk));
	jdff dff_B_oSmfh4520_2(.din(w_dff_B_4xesHF4G0_2),.dout(w_dff_B_oSmfh4520_2),.clk(gclk));
	jdff dff_B_aeVapTJW4_2(.din(w_dff_B_oSmfh4520_2),.dout(w_dff_B_aeVapTJW4_2),.clk(gclk));
	jdff dff_B_uFbkJfIW6_2(.din(w_dff_B_aeVapTJW4_2),.dout(w_dff_B_uFbkJfIW6_2),.clk(gclk));
	jdff dff_B_JlqX9ns16_2(.din(w_dff_B_uFbkJfIW6_2),.dout(w_dff_B_JlqX9ns16_2),.clk(gclk));
	jdff dff_B_8Skiq7x46_2(.din(w_dff_B_JlqX9ns16_2),.dout(w_dff_B_8Skiq7x46_2),.clk(gclk));
	jdff dff_B_3fns5Lo26_2(.din(w_dff_B_8Skiq7x46_2),.dout(w_dff_B_3fns5Lo26_2),.clk(gclk));
	jdff dff_B_waS7hUIH8_2(.din(w_dff_B_3fns5Lo26_2),.dout(w_dff_B_waS7hUIH8_2),.clk(gclk));
	jdff dff_B_le8oUxGK1_2(.din(w_dff_B_waS7hUIH8_2),.dout(w_dff_B_le8oUxGK1_2),.clk(gclk));
	jdff dff_B_YBxTBeR39_2(.din(w_dff_B_le8oUxGK1_2),.dout(w_dff_B_YBxTBeR39_2),.clk(gclk));
	jdff dff_B_ZRLwk30u8_2(.din(w_dff_B_YBxTBeR39_2),.dout(w_dff_B_ZRLwk30u8_2),.clk(gclk));
	jdff dff_B_Dj7xdSpz2_2(.din(w_dff_B_ZRLwk30u8_2),.dout(w_dff_B_Dj7xdSpz2_2),.clk(gclk));
	jdff dff_B_3auqZdgw9_1(.din(n1778),.dout(w_dff_B_3auqZdgw9_1),.clk(gclk));
	jdff dff_B_zYTpJKxQ4_1(.din(w_dff_B_3auqZdgw9_1),.dout(w_dff_B_zYTpJKxQ4_1),.clk(gclk));
	jdff dff_B_sg2mavvN5_2(.din(n1777),.dout(w_dff_B_sg2mavvN5_2),.clk(gclk));
	jdff dff_B_pS9fdlhH7_2(.din(w_dff_B_sg2mavvN5_2),.dout(w_dff_B_pS9fdlhH7_2),.clk(gclk));
	jdff dff_B_9WDbVEhb6_2(.din(w_dff_B_pS9fdlhH7_2),.dout(w_dff_B_9WDbVEhb6_2),.clk(gclk));
	jdff dff_B_LJyNPkMQ0_2(.din(w_dff_B_9WDbVEhb6_2),.dout(w_dff_B_LJyNPkMQ0_2),.clk(gclk));
	jdff dff_B_az27IJQC9_2(.din(w_dff_B_LJyNPkMQ0_2),.dout(w_dff_B_az27IJQC9_2),.clk(gclk));
	jdff dff_B_1tDdINop6_2(.din(w_dff_B_az27IJQC9_2),.dout(w_dff_B_1tDdINop6_2),.clk(gclk));
	jdff dff_B_tRMX78DR5_2(.din(w_dff_B_1tDdINop6_2),.dout(w_dff_B_tRMX78DR5_2),.clk(gclk));
	jdff dff_B_gE9WwGEE1_2(.din(w_dff_B_tRMX78DR5_2),.dout(w_dff_B_gE9WwGEE1_2),.clk(gclk));
	jdff dff_B_Qw11cTgW3_2(.din(w_dff_B_gE9WwGEE1_2),.dout(w_dff_B_Qw11cTgW3_2),.clk(gclk));
	jdff dff_B_AbhvIrOf0_2(.din(w_dff_B_Qw11cTgW3_2),.dout(w_dff_B_AbhvIrOf0_2),.clk(gclk));
	jdff dff_B_i6TYpp8K0_2(.din(w_dff_B_AbhvIrOf0_2),.dout(w_dff_B_i6TYpp8K0_2),.clk(gclk));
	jdff dff_B_pFrzBEDu3_2(.din(w_dff_B_i6TYpp8K0_2),.dout(w_dff_B_pFrzBEDu3_2),.clk(gclk));
	jdff dff_B_aFwl7LdJ1_2(.din(w_dff_B_pFrzBEDu3_2),.dout(w_dff_B_aFwl7LdJ1_2),.clk(gclk));
	jdff dff_B_0s1wmtCy3_2(.din(w_dff_B_aFwl7LdJ1_2),.dout(w_dff_B_0s1wmtCy3_2),.clk(gclk));
	jdff dff_B_dWLZ40NO8_2(.din(w_dff_B_0s1wmtCy3_2),.dout(w_dff_B_dWLZ40NO8_2),.clk(gclk));
	jdff dff_B_qsU24Evg2_2(.din(w_dff_B_dWLZ40NO8_2),.dout(w_dff_B_qsU24Evg2_2),.clk(gclk));
	jdff dff_B_VDvOjBsC3_2(.din(w_dff_B_qsU24Evg2_2),.dout(w_dff_B_VDvOjBsC3_2),.clk(gclk));
	jdff dff_B_76rPRpns2_2(.din(w_dff_B_VDvOjBsC3_2),.dout(w_dff_B_76rPRpns2_2),.clk(gclk));
	jdff dff_B_NKPJvvii0_2(.din(w_dff_B_76rPRpns2_2),.dout(w_dff_B_NKPJvvii0_2),.clk(gclk));
	jdff dff_B_wrnUSibZ5_2(.din(w_dff_B_NKPJvvii0_2),.dout(w_dff_B_wrnUSibZ5_2),.clk(gclk));
	jdff dff_B_shyQeqna7_2(.din(w_dff_B_wrnUSibZ5_2),.dout(w_dff_B_shyQeqna7_2),.clk(gclk));
	jdff dff_B_fLAw8DzZ7_2(.din(w_dff_B_shyQeqna7_2),.dout(w_dff_B_fLAw8DzZ7_2),.clk(gclk));
	jdff dff_B_0ovuIvrH5_2(.din(w_dff_B_fLAw8DzZ7_2),.dout(w_dff_B_0ovuIvrH5_2),.clk(gclk));
	jdff dff_B_KDWTfekR0_2(.din(w_dff_B_0ovuIvrH5_2),.dout(w_dff_B_KDWTfekR0_2),.clk(gclk));
	jdff dff_B_u834emlC2_2(.din(w_dff_B_KDWTfekR0_2),.dout(w_dff_B_u834emlC2_2),.clk(gclk));
	jdff dff_B_zNgEH4H47_2(.din(w_dff_B_u834emlC2_2),.dout(w_dff_B_zNgEH4H47_2),.clk(gclk));
	jdff dff_B_GnDBeocX5_2(.din(w_dff_B_zNgEH4H47_2),.dout(w_dff_B_GnDBeocX5_2),.clk(gclk));
	jdff dff_B_0WHItFsX6_2(.din(w_dff_B_GnDBeocX5_2),.dout(w_dff_B_0WHItFsX6_2),.clk(gclk));
	jdff dff_B_g2jzKlfp2_2(.din(w_dff_B_0WHItFsX6_2),.dout(w_dff_B_g2jzKlfp2_2),.clk(gclk));
	jdff dff_B_3UH7pmWz8_2(.din(w_dff_B_g2jzKlfp2_2),.dout(w_dff_B_3UH7pmWz8_2),.clk(gclk));
	jdff dff_B_1yogI9wc9_2(.din(w_dff_B_3UH7pmWz8_2),.dout(w_dff_B_1yogI9wc9_2),.clk(gclk));
	jdff dff_B_i3akOtyD8_2(.din(w_dff_B_1yogI9wc9_2),.dout(w_dff_B_i3akOtyD8_2),.clk(gclk));
	jdff dff_B_mr21e1yZ7_2(.din(w_dff_B_i3akOtyD8_2),.dout(w_dff_B_mr21e1yZ7_2),.clk(gclk));
	jdff dff_B_R1t0GcMK1_2(.din(w_dff_B_mr21e1yZ7_2),.dout(w_dff_B_R1t0GcMK1_2),.clk(gclk));
	jdff dff_B_g2WeaEwB7_2(.din(w_dff_B_R1t0GcMK1_2),.dout(w_dff_B_g2WeaEwB7_2),.clk(gclk));
	jdff dff_B_3qezBYm26_2(.din(w_dff_B_g2WeaEwB7_2),.dout(w_dff_B_3qezBYm26_2),.clk(gclk));
	jdff dff_B_NcT0JcZ80_2(.din(w_dff_B_3qezBYm26_2),.dout(w_dff_B_NcT0JcZ80_2),.clk(gclk));
	jdff dff_B_8mc1lKV28_2(.din(n1776),.dout(w_dff_B_8mc1lKV28_2),.clk(gclk));
	jdff dff_B_GqPxBzMg0_2(.din(w_dff_B_8mc1lKV28_2),.dout(w_dff_B_GqPxBzMg0_2),.clk(gclk));
	jdff dff_B_cr1DQ78h8_2(.din(w_dff_B_GqPxBzMg0_2),.dout(w_dff_B_cr1DQ78h8_2),.clk(gclk));
	jdff dff_B_ejgrpTFk1_2(.din(w_dff_B_cr1DQ78h8_2),.dout(w_dff_B_ejgrpTFk1_2),.clk(gclk));
	jdff dff_B_KqKqP7oH3_2(.din(w_dff_B_ejgrpTFk1_2),.dout(w_dff_B_KqKqP7oH3_2),.clk(gclk));
	jdff dff_B_uEsFci2l2_2(.din(w_dff_B_KqKqP7oH3_2),.dout(w_dff_B_uEsFci2l2_2),.clk(gclk));
	jdff dff_B_5Tf6ZIM33_2(.din(w_dff_B_uEsFci2l2_2),.dout(w_dff_B_5Tf6ZIM33_2),.clk(gclk));
	jdff dff_B_smSF9p9H3_2(.din(w_dff_B_5Tf6ZIM33_2),.dout(w_dff_B_smSF9p9H3_2),.clk(gclk));
	jdff dff_B_gHaagsHU1_2(.din(w_dff_B_smSF9p9H3_2),.dout(w_dff_B_gHaagsHU1_2),.clk(gclk));
	jdff dff_B_6NzrWgCe6_2(.din(w_dff_B_gHaagsHU1_2),.dout(w_dff_B_6NzrWgCe6_2),.clk(gclk));
	jdff dff_B_bWlLog5T2_2(.din(w_dff_B_6NzrWgCe6_2),.dout(w_dff_B_bWlLog5T2_2),.clk(gclk));
	jdff dff_B_D1lVgHXe2_2(.din(w_dff_B_bWlLog5T2_2),.dout(w_dff_B_D1lVgHXe2_2),.clk(gclk));
	jdff dff_B_Z40MKTgI9_2(.din(w_dff_B_D1lVgHXe2_2),.dout(w_dff_B_Z40MKTgI9_2),.clk(gclk));
	jdff dff_B_NDIuvHeO9_2(.din(w_dff_B_Z40MKTgI9_2),.dout(w_dff_B_NDIuvHeO9_2),.clk(gclk));
	jdff dff_B_ukxLGKj71_2(.din(w_dff_B_NDIuvHeO9_2),.dout(w_dff_B_ukxLGKj71_2),.clk(gclk));
	jdff dff_B_lOpKA3VI3_2(.din(w_dff_B_ukxLGKj71_2),.dout(w_dff_B_lOpKA3VI3_2),.clk(gclk));
	jdff dff_B_iTRW5P7E6_2(.din(w_dff_B_lOpKA3VI3_2),.dout(w_dff_B_iTRW5P7E6_2),.clk(gclk));
	jdff dff_B_qmBRteou8_2(.din(w_dff_B_iTRW5P7E6_2),.dout(w_dff_B_qmBRteou8_2),.clk(gclk));
	jdff dff_B_nRGPhBnc5_2(.din(w_dff_B_qmBRteou8_2),.dout(w_dff_B_nRGPhBnc5_2),.clk(gclk));
	jdff dff_B_4DovabGS0_2(.din(w_dff_B_nRGPhBnc5_2),.dout(w_dff_B_4DovabGS0_2),.clk(gclk));
	jdff dff_B_OVLMxxRT3_2(.din(w_dff_B_4DovabGS0_2),.dout(w_dff_B_OVLMxxRT3_2),.clk(gclk));
	jdff dff_B_IC4EYiKF8_2(.din(w_dff_B_OVLMxxRT3_2),.dout(w_dff_B_IC4EYiKF8_2),.clk(gclk));
	jdff dff_B_qzb9UkMo0_2(.din(w_dff_B_IC4EYiKF8_2),.dout(w_dff_B_qzb9UkMo0_2),.clk(gclk));
	jdff dff_B_eC85rIfO7_2(.din(w_dff_B_qzb9UkMo0_2),.dout(w_dff_B_eC85rIfO7_2),.clk(gclk));
	jdff dff_B_ROHnfLMl0_2(.din(w_dff_B_eC85rIfO7_2),.dout(w_dff_B_ROHnfLMl0_2),.clk(gclk));
	jdff dff_B_5SCm5VnK6_2(.din(w_dff_B_ROHnfLMl0_2),.dout(w_dff_B_5SCm5VnK6_2),.clk(gclk));
	jdff dff_B_K5y9wFPd3_2(.din(w_dff_B_5SCm5VnK6_2),.dout(w_dff_B_K5y9wFPd3_2),.clk(gclk));
	jdff dff_B_ptXQ1yug0_2(.din(w_dff_B_K5y9wFPd3_2),.dout(w_dff_B_ptXQ1yug0_2),.clk(gclk));
	jdff dff_B_4szw6T7j3_2(.din(w_dff_B_ptXQ1yug0_2),.dout(w_dff_B_4szw6T7j3_2),.clk(gclk));
	jdff dff_B_Nm2Dtv0K2_2(.din(w_dff_B_4szw6T7j3_2),.dout(w_dff_B_Nm2Dtv0K2_2),.clk(gclk));
	jdff dff_B_k9cqx16A9_2(.din(w_dff_B_Nm2Dtv0K2_2),.dout(w_dff_B_k9cqx16A9_2),.clk(gclk));
	jdff dff_B_dEjuMNy99_2(.din(w_dff_B_k9cqx16A9_2),.dout(w_dff_B_dEjuMNy99_2),.clk(gclk));
	jdff dff_B_CAAMQcNK6_2(.din(w_dff_B_dEjuMNy99_2),.dout(w_dff_B_CAAMQcNK6_2),.clk(gclk));
	jdff dff_B_tBM7LcQZ8_2(.din(w_dff_B_CAAMQcNK6_2),.dout(w_dff_B_tBM7LcQZ8_2),.clk(gclk));
	jdff dff_B_h5pPy9Gq6_2(.din(w_dff_B_tBM7LcQZ8_2),.dout(w_dff_B_h5pPy9Gq6_2),.clk(gclk));
	jdff dff_B_U4BB5Ajd1_2(.din(w_dff_B_h5pPy9Gq6_2),.dout(w_dff_B_U4BB5Ajd1_2),.clk(gclk));
	jdff dff_B_Eh7djlWD7_2(.din(w_dff_B_U4BB5Ajd1_2),.dout(w_dff_B_Eh7djlWD7_2),.clk(gclk));
	jdff dff_B_dh6cliBu6_2(.din(w_dff_B_Eh7djlWD7_2),.dout(w_dff_B_dh6cliBu6_2),.clk(gclk));
	jdff dff_B_N7U1sZEN0_2(.din(w_dff_B_dh6cliBu6_2),.dout(w_dff_B_N7U1sZEN0_2),.clk(gclk));
	jdff dff_B_QmpOAylZ8_2(.din(n1775),.dout(w_dff_B_QmpOAylZ8_2),.clk(gclk));
	jdff dff_B_OVlA1riG1_1(.din(n1773),.dout(w_dff_B_OVlA1riG1_1),.clk(gclk));
	jdff dff_B_PudRumwI7_2(.din(n1744),.dout(w_dff_B_PudRumwI7_2),.clk(gclk));
	jdff dff_B_G7WhFNlR7_2(.din(w_dff_B_PudRumwI7_2),.dout(w_dff_B_G7WhFNlR7_2),.clk(gclk));
	jdff dff_B_nHiYpvdv8_2(.din(w_dff_B_G7WhFNlR7_2),.dout(w_dff_B_nHiYpvdv8_2),.clk(gclk));
	jdff dff_B_dMAIWCWd5_2(.din(w_dff_B_nHiYpvdv8_2),.dout(w_dff_B_dMAIWCWd5_2),.clk(gclk));
	jdff dff_B_TV2lb9Qr7_2(.din(w_dff_B_dMAIWCWd5_2),.dout(w_dff_B_TV2lb9Qr7_2),.clk(gclk));
	jdff dff_B_VfEjBzbS8_2(.din(w_dff_B_TV2lb9Qr7_2),.dout(w_dff_B_VfEjBzbS8_2),.clk(gclk));
	jdff dff_B_EoPzviLr0_2(.din(w_dff_B_VfEjBzbS8_2),.dout(w_dff_B_EoPzviLr0_2),.clk(gclk));
	jdff dff_B_HIUk1tbM9_2(.din(w_dff_B_EoPzviLr0_2),.dout(w_dff_B_HIUk1tbM9_2),.clk(gclk));
	jdff dff_B_ID0UXKTq4_2(.din(w_dff_B_HIUk1tbM9_2),.dout(w_dff_B_ID0UXKTq4_2),.clk(gclk));
	jdff dff_B_5HarhjlT8_2(.din(w_dff_B_ID0UXKTq4_2),.dout(w_dff_B_5HarhjlT8_2),.clk(gclk));
	jdff dff_B_WWeK4A9S3_2(.din(w_dff_B_5HarhjlT8_2),.dout(w_dff_B_WWeK4A9S3_2),.clk(gclk));
	jdff dff_B_PWt0oHi46_2(.din(w_dff_B_WWeK4A9S3_2),.dout(w_dff_B_PWt0oHi46_2),.clk(gclk));
	jdff dff_B_c5udqjXK0_2(.din(w_dff_B_PWt0oHi46_2),.dout(w_dff_B_c5udqjXK0_2),.clk(gclk));
	jdff dff_B_Y8UO8W862_2(.din(w_dff_B_c5udqjXK0_2),.dout(w_dff_B_Y8UO8W862_2),.clk(gclk));
	jdff dff_B_R83J7hPy8_2(.din(w_dff_B_Y8UO8W862_2),.dout(w_dff_B_R83J7hPy8_2),.clk(gclk));
	jdff dff_B_vYn5Rclj8_2(.din(w_dff_B_R83J7hPy8_2),.dout(w_dff_B_vYn5Rclj8_2),.clk(gclk));
	jdff dff_B_q4gNGTDk7_2(.din(w_dff_B_vYn5Rclj8_2),.dout(w_dff_B_q4gNGTDk7_2),.clk(gclk));
	jdff dff_B_UAqestjT4_2(.din(w_dff_B_q4gNGTDk7_2),.dout(w_dff_B_UAqestjT4_2),.clk(gclk));
	jdff dff_B_4pQ4nEZ16_2(.din(w_dff_B_UAqestjT4_2),.dout(w_dff_B_4pQ4nEZ16_2),.clk(gclk));
	jdff dff_B_CpkOYcdb4_2(.din(w_dff_B_4pQ4nEZ16_2),.dout(w_dff_B_CpkOYcdb4_2),.clk(gclk));
	jdff dff_B_KRDvAaAB4_2(.din(w_dff_B_CpkOYcdb4_2),.dout(w_dff_B_KRDvAaAB4_2),.clk(gclk));
	jdff dff_B_YgcIZrnC6_2(.din(w_dff_B_KRDvAaAB4_2),.dout(w_dff_B_YgcIZrnC6_2),.clk(gclk));
	jdff dff_B_HGXYVM893_2(.din(w_dff_B_YgcIZrnC6_2),.dout(w_dff_B_HGXYVM893_2),.clk(gclk));
	jdff dff_B_rBz5WxrJ7_2(.din(w_dff_B_HGXYVM893_2),.dout(w_dff_B_rBz5WxrJ7_2),.clk(gclk));
	jdff dff_B_Ss2BhEF81_2(.din(w_dff_B_rBz5WxrJ7_2),.dout(w_dff_B_Ss2BhEF81_2),.clk(gclk));
	jdff dff_B_97g0Y8sw0_2(.din(w_dff_B_Ss2BhEF81_2),.dout(w_dff_B_97g0Y8sw0_2),.clk(gclk));
	jdff dff_B_MCCsQti76_2(.din(w_dff_B_97g0Y8sw0_2),.dout(w_dff_B_MCCsQti76_2),.clk(gclk));
	jdff dff_B_QJUaVTYR3_2(.din(w_dff_B_MCCsQti76_2),.dout(w_dff_B_QJUaVTYR3_2),.clk(gclk));
	jdff dff_B_3Vz9W5ri0_2(.din(w_dff_B_QJUaVTYR3_2),.dout(w_dff_B_3Vz9W5ri0_2),.clk(gclk));
	jdff dff_B_FSODxsAg3_2(.din(w_dff_B_3Vz9W5ri0_2),.dout(w_dff_B_FSODxsAg3_2),.clk(gclk));
	jdff dff_B_yxrmKJhF4_2(.din(w_dff_B_FSODxsAg3_2),.dout(w_dff_B_yxrmKJhF4_2),.clk(gclk));
	jdff dff_B_WqiElvCE5_2(.din(w_dff_B_yxrmKJhF4_2),.dout(w_dff_B_WqiElvCE5_2),.clk(gclk));
	jdff dff_B_zaSjiBXE9_2(.din(w_dff_B_WqiElvCE5_2),.dout(w_dff_B_zaSjiBXE9_2),.clk(gclk));
	jdff dff_B_IeF7Vl8X5_2(.din(w_dff_B_zaSjiBXE9_2),.dout(w_dff_B_IeF7Vl8X5_2),.clk(gclk));
	jdff dff_B_ljm25N4D4_2(.din(w_dff_B_IeF7Vl8X5_2),.dout(w_dff_B_ljm25N4D4_2),.clk(gclk));
	jdff dff_B_5PF1bY5k4_2(.din(w_dff_B_ljm25N4D4_2),.dout(w_dff_B_5PF1bY5k4_2),.clk(gclk));
	jdff dff_B_esALD8hJ7_2(.din(w_dff_B_5PF1bY5k4_2),.dout(w_dff_B_esALD8hJ7_2),.clk(gclk));
	jdff dff_B_4ekOZUDN9_1(.din(n1750),.dout(w_dff_B_4ekOZUDN9_1),.clk(gclk));
	jdff dff_B_C8UvJwn70_1(.din(w_dff_B_4ekOZUDN9_1),.dout(w_dff_B_C8UvJwn70_1),.clk(gclk));
	jdff dff_B_VL9gpHbR8_2(.din(n1749),.dout(w_dff_B_VL9gpHbR8_2),.clk(gclk));
	jdff dff_B_bvMksMx30_2(.din(w_dff_B_VL9gpHbR8_2),.dout(w_dff_B_bvMksMx30_2),.clk(gclk));
	jdff dff_B_lGOzT4o96_2(.din(w_dff_B_bvMksMx30_2),.dout(w_dff_B_lGOzT4o96_2),.clk(gclk));
	jdff dff_B_eOwLewQw7_2(.din(w_dff_B_lGOzT4o96_2),.dout(w_dff_B_eOwLewQw7_2),.clk(gclk));
	jdff dff_B_2vA37C663_2(.din(w_dff_B_eOwLewQw7_2),.dout(w_dff_B_2vA37C663_2),.clk(gclk));
	jdff dff_B_DHJz70dY1_2(.din(w_dff_B_2vA37C663_2),.dout(w_dff_B_DHJz70dY1_2),.clk(gclk));
	jdff dff_B_5s2bCycI7_2(.din(w_dff_B_DHJz70dY1_2),.dout(w_dff_B_5s2bCycI7_2),.clk(gclk));
	jdff dff_B_a9twzAqb3_2(.din(w_dff_B_5s2bCycI7_2),.dout(w_dff_B_a9twzAqb3_2),.clk(gclk));
	jdff dff_B_JX562nkH3_2(.din(w_dff_B_a9twzAqb3_2),.dout(w_dff_B_JX562nkH3_2),.clk(gclk));
	jdff dff_B_TydahiC79_2(.din(w_dff_B_JX562nkH3_2),.dout(w_dff_B_TydahiC79_2),.clk(gclk));
	jdff dff_B_mUI8mGD98_2(.din(w_dff_B_TydahiC79_2),.dout(w_dff_B_mUI8mGD98_2),.clk(gclk));
	jdff dff_B_Aow0IKm28_2(.din(w_dff_B_mUI8mGD98_2),.dout(w_dff_B_Aow0IKm28_2),.clk(gclk));
	jdff dff_B_T10lSKPT1_2(.din(w_dff_B_Aow0IKm28_2),.dout(w_dff_B_T10lSKPT1_2),.clk(gclk));
	jdff dff_B_smu5n5i33_2(.din(w_dff_B_T10lSKPT1_2),.dout(w_dff_B_smu5n5i33_2),.clk(gclk));
	jdff dff_B_5TYoeds34_2(.din(w_dff_B_smu5n5i33_2),.dout(w_dff_B_5TYoeds34_2),.clk(gclk));
	jdff dff_B_vMzbbPHs7_2(.din(w_dff_B_5TYoeds34_2),.dout(w_dff_B_vMzbbPHs7_2),.clk(gclk));
	jdff dff_B_LQS0kSTl9_2(.din(w_dff_B_vMzbbPHs7_2),.dout(w_dff_B_LQS0kSTl9_2),.clk(gclk));
	jdff dff_B_fnOuQwx36_2(.din(w_dff_B_LQS0kSTl9_2),.dout(w_dff_B_fnOuQwx36_2),.clk(gclk));
	jdff dff_B_Z7k21gL23_2(.din(w_dff_B_fnOuQwx36_2),.dout(w_dff_B_Z7k21gL23_2),.clk(gclk));
	jdff dff_B_pPR7WpkX7_2(.din(w_dff_B_Z7k21gL23_2),.dout(w_dff_B_pPR7WpkX7_2),.clk(gclk));
	jdff dff_B_9ORiV7NU0_2(.din(w_dff_B_pPR7WpkX7_2),.dout(w_dff_B_9ORiV7NU0_2),.clk(gclk));
	jdff dff_B_HZwUXxkj2_2(.din(w_dff_B_9ORiV7NU0_2),.dout(w_dff_B_HZwUXxkj2_2),.clk(gclk));
	jdff dff_B_29q95w5m4_2(.din(w_dff_B_HZwUXxkj2_2),.dout(w_dff_B_29q95w5m4_2),.clk(gclk));
	jdff dff_B_MGAjrWON1_2(.din(w_dff_B_29q95w5m4_2),.dout(w_dff_B_MGAjrWON1_2),.clk(gclk));
	jdff dff_B_kGciZmGr4_2(.din(w_dff_B_MGAjrWON1_2),.dout(w_dff_B_kGciZmGr4_2),.clk(gclk));
	jdff dff_B_iKgUAloo5_2(.din(w_dff_B_kGciZmGr4_2),.dout(w_dff_B_iKgUAloo5_2),.clk(gclk));
	jdff dff_B_BaJPbYQH2_2(.din(w_dff_B_iKgUAloo5_2),.dout(w_dff_B_BaJPbYQH2_2),.clk(gclk));
	jdff dff_B_1DBghht21_2(.din(w_dff_B_BaJPbYQH2_2),.dout(w_dff_B_1DBghht21_2),.clk(gclk));
	jdff dff_B_Qu9kvEKb1_2(.din(w_dff_B_1DBghht21_2),.dout(w_dff_B_Qu9kvEKb1_2),.clk(gclk));
	jdff dff_B_1lmnw1El5_2(.din(w_dff_B_Qu9kvEKb1_2),.dout(w_dff_B_1lmnw1El5_2),.clk(gclk));
	jdff dff_B_6sUrJhUZ5_2(.din(w_dff_B_1lmnw1El5_2),.dout(w_dff_B_6sUrJhUZ5_2),.clk(gclk));
	jdff dff_B_NpxVmRyW3_2(.din(w_dff_B_6sUrJhUZ5_2),.dout(w_dff_B_NpxVmRyW3_2),.clk(gclk));
	jdff dff_B_Pri80Zi09_2(.din(w_dff_B_NpxVmRyW3_2),.dout(w_dff_B_Pri80Zi09_2),.clk(gclk));
	jdff dff_B_yP0NFXiX9_2(.din(w_dff_B_Pri80Zi09_2),.dout(w_dff_B_yP0NFXiX9_2),.clk(gclk));
	jdff dff_B_Woql476Z1_2(.din(n1748),.dout(w_dff_B_Woql476Z1_2),.clk(gclk));
	jdff dff_B_A2JzMxBB2_2(.din(w_dff_B_Woql476Z1_2),.dout(w_dff_B_A2JzMxBB2_2),.clk(gclk));
	jdff dff_B_r20sFKo12_2(.din(w_dff_B_A2JzMxBB2_2),.dout(w_dff_B_r20sFKo12_2),.clk(gclk));
	jdff dff_B_oleP03xa7_2(.din(w_dff_B_r20sFKo12_2),.dout(w_dff_B_oleP03xa7_2),.clk(gclk));
	jdff dff_B_21qc8pcD9_2(.din(w_dff_B_oleP03xa7_2),.dout(w_dff_B_21qc8pcD9_2),.clk(gclk));
	jdff dff_B_UuZnL1N34_2(.din(w_dff_B_21qc8pcD9_2),.dout(w_dff_B_UuZnL1N34_2),.clk(gclk));
	jdff dff_B_ymgo2JbN4_2(.din(w_dff_B_UuZnL1N34_2),.dout(w_dff_B_ymgo2JbN4_2),.clk(gclk));
	jdff dff_B_HjrqiORL1_2(.din(w_dff_B_ymgo2JbN4_2),.dout(w_dff_B_HjrqiORL1_2),.clk(gclk));
	jdff dff_B_TSQbmhJl4_2(.din(w_dff_B_HjrqiORL1_2),.dout(w_dff_B_TSQbmhJl4_2),.clk(gclk));
	jdff dff_B_9LJN5TX37_2(.din(w_dff_B_TSQbmhJl4_2),.dout(w_dff_B_9LJN5TX37_2),.clk(gclk));
	jdff dff_B_8I0wKCJG3_2(.din(w_dff_B_9LJN5TX37_2),.dout(w_dff_B_8I0wKCJG3_2),.clk(gclk));
	jdff dff_B_j0dfOK7A1_2(.din(w_dff_B_8I0wKCJG3_2),.dout(w_dff_B_j0dfOK7A1_2),.clk(gclk));
	jdff dff_B_f5KTIVCu3_2(.din(w_dff_B_j0dfOK7A1_2),.dout(w_dff_B_f5KTIVCu3_2),.clk(gclk));
	jdff dff_B_83Vm3xNJ7_2(.din(w_dff_B_f5KTIVCu3_2),.dout(w_dff_B_83Vm3xNJ7_2),.clk(gclk));
	jdff dff_B_hPb3wsOR0_2(.din(w_dff_B_83Vm3xNJ7_2),.dout(w_dff_B_hPb3wsOR0_2),.clk(gclk));
	jdff dff_B_9etpv8vD6_2(.din(w_dff_B_hPb3wsOR0_2),.dout(w_dff_B_9etpv8vD6_2),.clk(gclk));
	jdff dff_B_UemEuhga8_2(.din(w_dff_B_9etpv8vD6_2),.dout(w_dff_B_UemEuhga8_2),.clk(gclk));
	jdff dff_B_F44TWHRK4_2(.din(w_dff_B_UemEuhga8_2),.dout(w_dff_B_F44TWHRK4_2),.clk(gclk));
	jdff dff_B_ZQKdpPTj7_2(.din(w_dff_B_F44TWHRK4_2),.dout(w_dff_B_ZQKdpPTj7_2),.clk(gclk));
	jdff dff_B_pKHb5SW60_2(.din(w_dff_B_ZQKdpPTj7_2),.dout(w_dff_B_pKHb5SW60_2),.clk(gclk));
	jdff dff_B_JVTya3gm1_2(.din(w_dff_B_pKHb5SW60_2),.dout(w_dff_B_JVTya3gm1_2),.clk(gclk));
	jdff dff_B_rF4N1plO2_2(.din(w_dff_B_JVTya3gm1_2),.dout(w_dff_B_rF4N1plO2_2),.clk(gclk));
	jdff dff_B_Zz8qDjjB5_2(.din(w_dff_B_rF4N1plO2_2),.dout(w_dff_B_Zz8qDjjB5_2),.clk(gclk));
	jdff dff_B_NT0WVFNs6_2(.din(w_dff_B_Zz8qDjjB5_2),.dout(w_dff_B_NT0WVFNs6_2),.clk(gclk));
	jdff dff_B_Qy6zbgpi8_2(.din(w_dff_B_NT0WVFNs6_2),.dout(w_dff_B_Qy6zbgpi8_2),.clk(gclk));
	jdff dff_B_3nhjBr1H5_2(.din(w_dff_B_Qy6zbgpi8_2),.dout(w_dff_B_3nhjBr1H5_2),.clk(gclk));
	jdff dff_B_FTJWA3Wb0_2(.din(w_dff_B_3nhjBr1H5_2),.dout(w_dff_B_FTJWA3Wb0_2),.clk(gclk));
	jdff dff_B_xsiyaY1M4_2(.din(w_dff_B_FTJWA3Wb0_2),.dout(w_dff_B_xsiyaY1M4_2),.clk(gclk));
	jdff dff_B_LRvlqsUy2_2(.din(w_dff_B_xsiyaY1M4_2),.dout(w_dff_B_LRvlqsUy2_2),.clk(gclk));
	jdff dff_B_VyxlMqUh6_2(.din(w_dff_B_LRvlqsUy2_2),.dout(w_dff_B_VyxlMqUh6_2),.clk(gclk));
	jdff dff_B_pCqbXJPl6_2(.din(w_dff_B_VyxlMqUh6_2),.dout(w_dff_B_pCqbXJPl6_2),.clk(gclk));
	jdff dff_B_frj9NEkF7_2(.din(w_dff_B_pCqbXJPl6_2),.dout(w_dff_B_frj9NEkF7_2),.clk(gclk));
	jdff dff_B_jZ2hx3oF8_2(.din(w_dff_B_frj9NEkF7_2),.dout(w_dff_B_jZ2hx3oF8_2),.clk(gclk));
	jdff dff_B_yqHE6R9N4_2(.din(w_dff_B_jZ2hx3oF8_2),.dout(w_dff_B_yqHE6R9N4_2),.clk(gclk));
	jdff dff_B_dQZqkU7Z0_2(.din(w_dff_B_yqHE6R9N4_2),.dout(w_dff_B_dQZqkU7Z0_2),.clk(gclk));
	jdff dff_B_ooyi4Dhj8_2(.din(w_dff_B_dQZqkU7Z0_2),.dout(w_dff_B_ooyi4Dhj8_2),.clk(gclk));
	jdff dff_B_uKa30N7n8_2(.din(n1747),.dout(w_dff_B_uKa30N7n8_2),.clk(gclk));
	jdff dff_B_KAPZZ2M51_1(.din(n1745),.dout(w_dff_B_KAPZZ2M51_1),.clk(gclk));
	jdff dff_B_8KQSmLxP1_2(.din(n1709),.dout(w_dff_B_8KQSmLxP1_2),.clk(gclk));
	jdff dff_B_cnm4pNU53_2(.din(w_dff_B_8KQSmLxP1_2),.dout(w_dff_B_cnm4pNU53_2),.clk(gclk));
	jdff dff_B_NFKLhRmT6_2(.din(w_dff_B_cnm4pNU53_2),.dout(w_dff_B_NFKLhRmT6_2),.clk(gclk));
	jdff dff_B_1PDCU8Ch8_2(.din(w_dff_B_NFKLhRmT6_2),.dout(w_dff_B_1PDCU8Ch8_2),.clk(gclk));
	jdff dff_B_EFICxePJ5_2(.din(w_dff_B_1PDCU8Ch8_2),.dout(w_dff_B_EFICxePJ5_2),.clk(gclk));
	jdff dff_B_Rnrr9CHp0_2(.din(w_dff_B_EFICxePJ5_2),.dout(w_dff_B_Rnrr9CHp0_2),.clk(gclk));
	jdff dff_B_insuvd4Z9_2(.din(w_dff_B_Rnrr9CHp0_2),.dout(w_dff_B_insuvd4Z9_2),.clk(gclk));
	jdff dff_B_9nTySo4Z6_2(.din(w_dff_B_insuvd4Z9_2),.dout(w_dff_B_9nTySo4Z6_2),.clk(gclk));
	jdff dff_B_xMufBLpJ6_2(.din(w_dff_B_9nTySo4Z6_2),.dout(w_dff_B_xMufBLpJ6_2),.clk(gclk));
	jdff dff_B_QbNkok730_2(.din(w_dff_B_xMufBLpJ6_2),.dout(w_dff_B_QbNkok730_2),.clk(gclk));
	jdff dff_B_uqRpqt195_2(.din(w_dff_B_QbNkok730_2),.dout(w_dff_B_uqRpqt195_2),.clk(gclk));
	jdff dff_B_Tia6Esri0_2(.din(w_dff_B_uqRpqt195_2),.dout(w_dff_B_Tia6Esri0_2),.clk(gclk));
	jdff dff_B_XtenYsO29_2(.din(w_dff_B_Tia6Esri0_2),.dout(w_dff_B_XtenYsO29_2),.clk(gclk));
	jdff dff_B_2uom0cBa3_2(.din(w_dff_B_XtenYsO29_2),.dout(w_dff_B_2uom0cBa3_2),.clk(gclk));
	jdff dff_B_b25gftLS0_2(.din(w_dff_B_2uom0cBa3_2),.dout(w_dff_B_b25gftLS0_2),.clk(gclk));
	jdff dff_B_R5PNm0si2_2(.din(w_dff_B_b25gftLS0_2),.dout(w_dff_B_R5PNm0si2_2),.clk(gclk));
	jdff dff_B_0PFFGdyc2_2(.din(w_dff_B_R5PNm0si2_2),.dout(w_dff_B_0PFFGdyc2_2),.clk(gclk));
	jdff dff_B_dsgKG87Q3_2(.din(w_dff_B_0PFFGdyc2_2),.dout(w_dff_B_dsgKG87Q3_2),.clk(gclk));
	jdff dff_B_seZZcPUD7_2(.din(w_dff_B_dsgKG87Q3_2),.dout(w_dff_B_seZZcPUD7_2),.clk(gclk));
	jdff dff_B_UbrrY6Uw3_2(.din(w_dff_B_seZZcPUD7_2),.dout(w_dff_B_UbrrY6Uw3_2),.clk(gclk));
	jdff dff_B_PkNCOy2u6_2(.din(w_dff_B_UbrrY6Uw3_2),.dout(w_dff_B_PkNCOy2u6_2),.clk(gclk));
	jdff dff_B_yWPTjqYi3_2(.din(w_dff_B_PkNCOy2u6_2),.dout(w_dff_B_yWPTjqYi3_2),.clk(gclk));
	jdff dff_B_XTqvdSER0_2(.din(w_dff_B_yWPTjqYi3_2),.dout(w_dff_B_XTqvdSER0_2),.clk(gclk));
	jdff dff_B_blvJ59RF3_2(.din(w_dff_B_XTqvdSER0_2),.dout(w_dff_B_blvJ59RF3_2),.clk(gclk));
	jdff dff_B_3eWlahs43_2(.din(w_dff_B_blvJ59RF3_2),.dout(w_dff_B_3eWlahs43_2),.clk(gclk));
	jdff dff_B_kqu4Jbls1_2(.din(w_dff_B_3eWlahs43_2),.dout(w_dff_B_kqu4Jbls1_2),.clk(gclk));
	jdff dff_B_YYwiy0Yh6_2(.din(w_dff_B_kqu4Jbls1_2),.dout(w_dff_B_YYwiy0Yh6_2),.clk(gclk));
	jdff dff_B_xl5dLPUD7_2(.din(w_dff_B_YYwiy0Yh6_2),.dout(w_dff_B_xl5dLPUD7_2),.clk(gclk));
	jdff dff_B_qvUOXcKk3_2(.din(w_dff_B_xl5dLPUD7_2),.dout(w_dff_B_qvUOXcKk3_2),.clk(gclk));
	jdff dff_B_k0Ka6w7K9_2(.din(w_dff_B_qvUOXcKk3_2),.dout(w_dff_B_k0Ka6w7K9_2),.clk(gclk));
	jdff dff_B_WQwh4vy97_2(.din(w_dff_B_k0Ka6w7K9_2),.dout(w_dff_B_WQwh4vy97_2),.clk(gclk));
	jdff dff_B_R44vQg6Q5_2(.din(w_dff_B_WQwh4vy97_2),.dout(w_dff_B_R44vQg6Q5_2),.clk(gclk));
	jdff dff_B_DhdwAVrR1_2(.din(w_dff_B_R44vQg6Q5_2),.dout(w_dff_B_DhdwAVrR1_2),.clk(gclk));
	jdff dff_B_ng7MdjRo8_2(.din(w_dff_B_DhdwAVrR1_2),.dout(w_dff_B_ng7MdjRo8_2),.clk(gclk));
	jdff dff_B_CFkAHw0j4_1(.din(n1715),.dout(w_dff_B_CFkAHw0j4_1),.clk(gclk));
	jdff dff_B_wQmsM3qk1_1(.din(w_dff_B_CFkAHw0j4_1),.dout(w_dff_B_wQmsM3qk1_1),.clk(gclk));
	jdff dff_B_2HXbBIk07_2(.din(n1714),.dout(w_dff_B_2HXbBIk07_2),.clk(gclk));
	jdff dff_B_HBJaj7QS8_2(.din(w_dff_B_2HXbBIk07_2),.dout(w_dff_B_HBJaj7QS8_2),.clk(gclk));
	jdff dff_B_AHSOSasA8_2(.din(w_dff_B_HBJaj7QS8_2),.dout(w_dff_B_AHSOSasA8_2),.clk(gclk));
	jdff dff_B_kDCWsug17_2(.din(w_dff_B_AHSOSasA8_2),.dout(w_dff_B_kDCWsug17_2),.clk(gclk));
	jdff dff_B_EaZG6X1D3_2(.din(w_dff_B_kDCWsug17_2),.dout(w_dff_B_EaZG6X1D3_2),.clk(gclk));
	jdff dff_B_YvPlzF8T3_2(.din(w_dff_B_EaZG6X1D3_2),.dout(w_dff_B_YvPlzF8T3_2),.clk(gclk));
	jdff dff_B_lVGBjZCS0_2(.din(w_dff_B_YvPlzF8T3_2),.dout(w_dff_B_lVGBjZCS0_2),.clk(gclk));
	jdff dff_B_ZmA2cTQN0_2(.din(w_dff_B_lVGBjZCS0_2),.dout(w_dff_B_ZmA2cTQN0_2),.clk(gclk));
	jdff dff_B_C6pjOZAS9_2(.din(w_dff_B_ZmA2cTQN0_2),.dout(w_dff_B_C6pjOZAS9_2),.clk(gclk));
	jdff dff_B_GOdzJMOV5_2(.din(w_dff_B_C6pjOZAS9_2),.dout(w_dff_B_GOdzJMOV5_2),.clk(gclk));
	jdff dff_B_HBgPADSC2_2(.din(w_dff_B_GOdzJMOV5_2),.dout(w_dff_B_HBgPADSC2_2),.clk(gclk));
	jdff dff_B_Nbebmnft4_2(.din(w_dff_B_HBgPADSC2_2),.dout(w_dff_B_Nbebmnft4_2),.clk(gclk));
	jdff dff_B_xLOns4jM0_2(.din(w_dff_B_Nbebmnft4_2),.dout(w_dff_B_xLOns4jM0_2),.clk(gclk));
	jdff dff_B_6lmMNMfw7_2(.din(w_dff_B_xLOns4jM0_2),.dout(w_dff_B_6lmMNMfw7_2),.clk(gclk));
	jdff dff_B_PgY44oFz5_2(.din(w_dff_B_6lmMNMfw7_2),.dout(w_dff_B_PgY44oFz5_2),.clk(gclk));
	jdff dff_B_N1XXNetg8_2(.din(w_dff_B_PgY44oFz5_2),.dout(w_dff_B_N1XXNetg8_2),.clk(gclk));
	jdff dff_B_aSey69M92_2(.din(w_dff_B_N1XXNetg8_2),.dout(w_dff_B_aSey69M92_2),.clk(gclk));
	jdff dff_B_opsKTvnQ6_2(.din(w_dff_B_aSey69M92_2),.dout(w_dff_B_opsKTvnQ6_2),.clk(gclk));
	jdff dff_B_Q5gwx0sm8_2(.din(w_dff_B_opsKTvnQ6_2),.dout(w_dff_B_Q5gwx0sm8_2),.clk(gclk));
	jdff dff_B_5CLvqqWM2_2(.din(w_dff_B_Q5gwx0sm8_2),.dout(w_dff_B_5CLvqqWM2_2),.clk(gclk));
	jdff dff_B_48RxOUUx8_2(.din(w_dff_B_5CLvqqWM2_2),.dout(w_dff_B_48RxOUUx8_2),.clk(gclk));
	jdff dff_B_Cz1MBfmd8_2(.din(w_dff_B_48RxOUUx8_2),.dout(w_dff_B_Cz1MBfmd8_2),.clk(gclk));
	jdff dff_B_trv2bQy57_2(.din(w_dff_B_Cz1MBfmd8_2),.dout(w_dff_B_trv2bQy57_2),.clk(gclk));
	jdff dff_B_DRpjh5Yl3_2(.din(w_dff_B_trv2bQy57_2),.dout(w_dff_B_DRpjh5Yl3_2),.clk(gclk));
	jdff dff_B_qe0x86h46_2(.din(w_dff_B_DRpjh5Yl3_2),.dout(w_dff_B_qe0x86h46_2),.clk(gclk));
	jdff dff_B_iCjHO4bM6_2(.din(w_dff_B_qe0x86h46_2),.dout(w_dff_B_iCjHO4bM6_2),.clk(gclk));
	jdff dff_B_rPKcuSzv0_2(.din(w_dff_B_iCjHO4bM6_2),.dout(w_dff_B_rPKcuSzv0_2),.clk(gclk));
	jdff dff_B_q1QBB7zv9_2(.din(w_dff_B_rPKcuSzv0_2),.dout(w_dff_B_q1QBB7zv9_2),.clk(gclk));
	jdff dff_B_SrxSrW0G3_2(.din(w_dff_B_q1QBB7zv9_2),.dout(w_dff_B_SrxSrW0G3_2),.clk(gclk));
	jdff dff_B_wNjID34g5_2(.din(w_dff_B_SrxSrW0G3_2),.dout(w_dff_B_wNjID34g5_2),.clk(gclk));
	jdff dff_B_J7N8fnvp0_2(.din(w_dff_B_wNjID34g5_2),.dout(w_dff_B_J7N8fnvp0_2),.clk(gclk));
	jdff dff_B_nFvh7y3i3_2(.din(n1713),.dout(w_dff_B_nFvh7y3i3_2),.clk(gclk));
	jdff dff_B_i0Yvv1N56_2(.din(w_dff_B_nFvh7y3i3_2),.dout(w_dff_B_i0Yvv1N56_2),.clk(gclk));
	jdff dff_B_IQO3mTKG1_2(.din(w_dff_B_i0Yvv1N56_2),.dout(w_dff_B_IQO3mTKG1_2),.clk(gclk));
	jdff dff_B_3v0ADI9U9_2(.din(w_dff_B_IQO3mTKG1_2),.dout(w_dff_B_3v0ADI9U9_2),.clk(gclk));
	jdff dff_B_SBtpTMJZ5_2(.din(w_dff_B_3v0ADI9U9_2),.dout(w_dff_B_SBtpTMJZ5_2),.clk(gclk));
	jdff dff_B_CNvUG9B36_2(.din(w_dff_B_SBtpTMJZ5_2),.dout(w_dff_B_CNvUG9B36_2),.clk(gclk));
	jdff dff_B_XKkhD4X06_2(.din(w_dff_B_CNvUG9B36_2),.dout(w_dff_B_XKkhD4X06_2),.clk(gclk));
	jdff dff_B_U0yjbSxp9_2(.din(w_dff_B_XKkhD4X06_2),.dout(w_dff_B_U0yjbSxp9_2),.clk(gclk));
	jdff dff_B_MJHupzjb4_2(.din(w_dff_B_U0yjbSxp9_2),.dout(w_dff_B_MJHupzjb4_2),.clk(gclk));
	jdff dff_B_dNBU1pdN0_2(.din(w_dff_B_MJHupzjb4_2),.dout(w_dff_B_dNBU1pdN0_2),.clk(gclk));
	jdff dff_B_WyXfI5dU9_2(.din(w_dff_B_dNBU1pdN0_2),.dout(w_dff_B_WyXfI5dU9_2),.clk(gclk));
	jdff dff_B_qyILnLYn9_2(.din(w_dff_B_WyXfI5dU9_2),.dout(w_dff_B_qyILnLYn9_2),.clk(gclk));
	jdff dff_B_DEw2b6Ni3_2(.din(w_dff_B_qyILnLYn9_2),.dout(w_dff_B_DEw2b6Ni3_2),.clk(gclk));
	jdff dff_B_CcSxBsZl0_2(.din(w_dff_B_DEw2b6Ni3_2),.dout(w_dff_B_CcSxBsZl0_2),.clk(gclk));
	jdff dff_B_mfXXv0Vv0_2(.din(w_dff_B_CcSxBsZl0_2),.dout(w_dff_B_mfXXv0Vv0_2),.clk(gclk));
	jdff dff_B_Ze9ugTDp0_2(.din(w_dff_B_mfXXv0Vv0_2),.dout(w_dff_B_Ze9ugTDp0_2),.clk(gclk));
	jdff dff_B_fpkHUbGs2_2(.din(w_dff_B_Ze9ugTDp0_2),.dout(w_dff_B_fpkHUbGs2_2),.clk(gclk));
	jdff dff_B_DLqJCdGJ9_2(.din(w_dff_B_fpkHUbGs2_2),.dout(w_dff_B_DLqJCdGJ9_2),.clk(gclk));
	jdff dff_B_eysHXuh48_2(.din(w_dff_B_DLqJCdGJ9_2),.dout(w_dff_B_eysHXuh48_2),.clk(gclk));
	jdff dff_B_NrQ5MYUw1_2(.din(w_dff_B_eysHXuh48_2),.dout(w_dff_B_NrQ5MYUw1_2),.clk(gclk));
	jdff dff_B_DKVkEJvC0_2(.din(w_dff_B_NrQ5MYUw1_2),.dout(w_dff_B_DKVkEJvC0_2),.clk(gclk));
	jdff dff_B_LCT4YpCV1_2(.din(w_dff_B_DKVkEJvC0_2),.dout(w_dff_B_LCT4YpCV1_2),.clk(gclk));
	jdff dff_B_VHjWto203_2(.din(w_dff_B_LCT4YpCV1_2),.dout(w_dff_B_VHjWto203_2),.clk(gclk));
	jdff dff_B_C9jrjA3o5_2(.din(w_dff_B_VHjWto203_2),.dout(w_dff_B_C9jrjA3o5_2),.clk(gclk));
	jdff dff_B_26Q163G92_2(.din(w_dff_B_C9jrjA3o5_2),.dout(w_dff_B_26Q163G92_2),.clk(gclk));
	jdff dff_B_uuzQMzJQ0_2(.din(w_dff_B_26Q163G92_2),.dout(w_dff_B_uuzQMzJQ0_2),.clk(gclk));
	jdff dff_B_Io0IbmwZ1_2(.din(w_dff_B_uuzQMzJQ0_2),.dout(w_dff_B_Io0IbmwZ1_2),.clk(gclk));
	jdff dff_B_aBRr0VjG5_2(.din(w_dff_B_Io0IbmwZ1_2),.dout(w_dff_B_aBRr0VjG5_2),.clk(gclk));
	jdff dff_B_xgmijSJq7_2(.din(w_dff_B_aBRr0VjG5_2),.dout(w_dff_B_xgmijSJq7_2),.clk(gclk));
	jdff dff_B_z7L8DSGO5_2(.din(w_dff_B_xgmijSJq7_2),.dout(w_dff_B_z7L8DSGO5_2),.clk(gclk));
	jdff dff_B_11QQPtNf5_2(.din(w_dff_B_z7L8DSGO5_2),.dout(w_dff_B_11QQPtNf5_2),.clk(gclk));
	jdff dff_B_D8krU0Ys7_2(.din(w_dff_B_11QQPtNf5_2),.dout(w_dff_B_D8krU0Ys7_2),.clk(gclk));
	jdff dff_B_5MEgAAAv1_2(.din(w_dff_B_D8krU0Ys7_2),.dout(w_dff_B_5MEgAAAv1_2),.clk(gclk));
	jdff dff_B_FwikrSQf0_2(.din(n1712),.dout(w_dff_B_FwikrSQf0_2),.clk(gclk));
	jdff dff_B_sTlKSnnr0_1(.din(n1710),.dout(w_dff_B_sTlKSnnr0_1),.clk(gclk));
	jdff dff_B_UWIdUfXK9_2(.din(n1668),.dout(w_dff_B_UWIdUfXK9_2),.clk(gclk));
	jdff dff_B_qWDmvnZ22_2(.din(w_dff_B_UWIdUfXK9_2),.dout(w_dff_B_qWDmvnZ22_2),.clk(gclk));
	jdff dff_B_KxwnxxyK8_2(.din(w_dff_B_qWDmvnZ22_2),.dout(w_dff_B_KxwnxxyK8_2),.clk(gclk));
	jdff dff_B_ctu5O80e3_2(.din(w_dff_B_KxwnxxyK8_2),.dout(w_dff_B_ctu5O80e3_2),.clk(gclk));
	jdff dff_B_ybng71f38_2(.din(w_dff_B_ctu5O80e3_2),.dout(w_dff_B_ybng71f38_2),.clk(gclk));
	jdff dff_B_aVfBNds87_2(.din(w_dff_B_ybng71f38_2),.dout(w_dff_B_aVfBNds87_2),.clk(gclk));
	jdff dff_B_T3Kn75uS2_2(.din(w_dff_B_aVfBNds87_2),.dout(w_dff_B_T3Kn75uS2_2),.clk(gclk));
	jdff dff_B_JIrNpzIs4_2(.din(w_dff_B_T3Kn75uS2_2),.dout(w_dff_B_JIrNpzIs4_2),.clk(gclk));
	jdff dff_B_q1fXV2007_2(.din(w_dff_B_JIrNpzIs4_2),.dout(w_dff_B_q1fXV2007_2),.clk(gclk));
	jdff dff_B_lfstOxSI8_2(.din(w_dff_B_q1fXV2007_2),.dout(w_dff_B_lfstOxSI8_2),.clk(gclk));
	jdff dff_B_Yw8iH4jl4_2(.din(w_dff_B_lfstOxSI8_2),.dout(w_dff_B_Yw8iH4jl4_2),.clk(gclk));
	jdff dff_B_6i0tAEd47_2(.din(w_dff_B_Yw8iH4jl4_2),.dout(w_dff_B_6i0tAEd47_2),.clk(gclk));
	jdff dff_B_Rl8xE0iy2_2(.din(w_dff_B_6i0tAEd47_2),.dout(w_dff_B_Rl8xE0iy2_2),.clk(gclk));
	jdff dff_B_PE1WyJXc6_2(.din(w_dff_B_Rl8xE0iy2_2),.dout(w_dff_B_PE1WyJXc6_2),.clk(gclk));
	jdff dff_B_fwnWuWeg8_2(.din(w_dff_B_PE1WyJXc6_2),.dout(w_dff_B_fwnWuWeg8_2),.clk(gclk));
	jdff dff_B_RwL3Twf68_2(.din(w_dff_B_fwnWuWeg8_2),.dout(w_dff_B_RwL3Twf68_2),.clk(gclk));
	jdff dff_B_NQRY5bSM3_2(.din(w_dff_B_RwL3Twf68_2),.dout(w_dff_B_NQRY5bSM3_2),.clk(gclk));
	jdff dff_B_oD7Naomz3_2(.din(w_dff_B_NQRY5bSM3_2),.dout(w_dff_B_oD7Naomz3_2),.clk(gclk));
	jdff dff_B_CqULvryu6_2(.din(w_dff_B_oD7Naomz3_2),.dout(w_dff_B_CqULvryu6_2),.clk(gclk));
	jdff dff_B_OPL3znrp7_2(.din(w_dff_B_CqULvryu6_2),.dout(w_dff_B_OPL3znrp7_2),.clk(gclk));
	jdff dff_B_JLRnP7sD5_2(.din(w_dff_B_OPL3znrp7_2),.dout(w_dff_B_JLRnP7sD5_2),.clk(gclk));
	jdff dff_B_uZBsouB98_2(.din(w_dff_B_JLRnP7sD5_2),.dout(w_dff_B_uZBsouB98_2),.clk(gclk));
	jdff dff_B_Zg290EZQ2_2(.din(w_dff_B_uZBsouB98_2),.dout(w_dff_B_Zg290EZQ2_2),.clk(gclk));
	jdff dff_B_PixasGwK6_2(.din(w_dff_B_Zg290EZQ2_2),.dout(w_dff_B_PixasGwK6_2),.clk(gclk));
	jdff dff_B_DyJhSiRb9_2(.din(w_dff_B_PixasGwK6_2),.dout(w_dff_B_DyJhSiRb9_2),.clk(gclk));
	jdff dff_B_KcHzvtVe1_2(.din(w_dff_B_DyJhSiRb9_2),.dout(w_dff_B_KcHzvtVe1_2),.clk(gclk));
	jdff dff_B_wBXmdGKi8_2(.din(w_dff_B_KcHzvtVe1_2),.dout(w_dff_B_wBXmdGKi8_2),.clk(gclk));
	jdff dff_B_j8eaVuxS5_2(.din(w_dff_B_wBXmdGKi8_2),.dout(w_dff_B_j8eaVuxS5_2),.clk(gclk));
	jdff dff_B_wa4oXp9q4_2(.din(w_dff_B_j8eaVuxS5_2),.dout(w_dff_B_wa4oXp9q4_2),.clk(gclk));
	jdff dff_B_zxwx0PPF5_2(.din(w_dff_B_wa4oXp9q4_2),.dout(w_dff_B_zxwx0PPF5_2),.clk(gclk));
	jdff dff_B_hapB8zjH4_2(.din(w_dff_B_zxwx0PPF5_2),.dout(w_dff_B_hapB8zjH4_2),.clk(gclk));
	jdff dff_B_CwM0rPiB5_1(.din(n1674),.dout(w_dff_B_CwM0rPiB5_1),.clk(gclk));
	jdff dff_B_OLhctYmw4_1(.din(w_dff_B_CwM0rPiB5_1),.dout(w_dff_B_OLhctYmw4_1),.clk(gclk));
	jdff dff_B_aKCpI4W40_2(.din(n1673),.dout(w_dff_B_aKCpI4W40_2),.clk(gclk));
	jdff dff_B_vg6D0js49_2(.din(w_dff_B_aKCpI4W40_2),.dout(w_dff_B_vg6D0js49_2),.clk(gclk));
	jdff dff_B_fKiiRoqR3_2(.din(w_dff_B_vg6D0js49_2),.dout(w_dff_B_fKiiRoqR3_2),.clk(gclk));
	jdff dff_B_6IGJbsmP9_2(.din(w_dff_B_fKiiRoqR3_2),.dout(w_dff_B_6IGJbsmP9_2),.clk(gclk));
	jdff dff_B_NbgeeVgi4_2(.din(w_dff_B_6IGJbsmP9_2),.dout(w_dff_B_NbgeeVgi4_2),.clk(gclk));
	jdff dff_B_f3PwT8SZ4_2(.din(w_dff_B_NbgeeVgi4_2),.dout(w_dff_B_f3PwT8SZ4_2),.clk(gclk));
	jdff dff_B_g0Si6Fu99_2(.din(w_dff_B_f3PwT8SZ4_2),.dout(w_dff_B_g0Si6Fu99_2),.clk(gclk));
	jdff dff_B_f53rVkJu8_2(.din(w_dff_B_g0Si6Fu99_2),.dout(w_dff_B_f53rVkJu8_2),.clk(gclk));
	jdff dff_B_0115tIk78_2(.din(w_dff_B_f53rVkJu8_2),.dout(w_dff_B_0115tIk78_2),.clk(gclk));
	jdff dff_B_637iVEJW7_2(.din(w_dff_B_0115tIk78_2),.dout(w_dff_B_637iVEJW7_2),.clk(gclk));
	jdff dff_B_MuNNHNug7_2(.din(w_dff_B_637iVEJW7_2),.dout(w_dff_B_MuNNHNug7_2),.clk(gclk));
	jdff dff_B_FoGxD9Oo3_2(.din(w_dff_B_MuNNHNug7_2),.dout(w_dff_B_FoGxD9Oo3_2),.clk(gclk));
	jdff dff_B_zm6CwYB79_2(.din(w_dff_B_FoGxD9Oo3_2),.dout(w_dff_B_zm6CwYB79_2),.clk(gclk));
	jdff dff_B_wN5lUYCb0_2(.din(w_dff_B_zm6CwYB79_2),.dout(w_dff_B_wN5lUYCb0_2),.clk(gclk));
	jdff dff_B_scVsnS9Q6_2(.din(w_dff_B_wN5lUYCb0_2),.dout(w_dff_B_scVsnS9Q6_2),.clk(gclk));
	jdff dff_B_8aYoBSwx4_2(.din(w_dff_B_scVsnS9Q6_2),.dout(w_dff_B_8aYoBSwx4_2),.clk(gclk));
	jdff dff_B_Zi1D8kvU1_2(.din(w_dff_B_8aYoBSwx4_2),.dout(w_dff_B_Zi1D8kvU1_2),.clk(gclk));
	jdff dff_B_7WdZfxw69_2(.din(w_dff_B_Zi1D8kvU1_2),.dout(w_dff_B_7WdZfxw69_2),.clk(gclk));
	jdff dff_B_wXT84iJF5_2(.din(w_dff_B_7WdZfxw69_2),.dout(w_dff_B_wXT84iJF5_2),.clk(gclk));
	jdff dff_B_lyGKtdyx4_2(.din(w_dff_B_wXT84iJF5_2),.dout(w_dff_B_lyGKtdyx4_2),.clk(gclk));
	jdff dff_B_NfaMFL8B7_2(.din(w_dff_B_lyGKtdyx4_2),.dout(w_dff_B_NfaMFL8B7_2),.clk(gclk));
	jdff dff_B_G8oGNQ6C3_2(.din(w_dff_B_NfaMFL8B7_2),.dout(w_dff_B_G8oGNQ6C3_2),.clk(gclk));
	jdff dff_B_CsFmnnYz9_2(.din(w_dff_B_G8oGNQ6C3_2),.dout(w_dff_B_CsFmnnYz9_2),.clk(gclk));
	jdff dff_B_fJvYJ8zi7_2(.din(w_dff_B_CsFmnnYz9_2),.dout(w_dff_B_fJvYJ8zi7_2),.clk(gclk));
	jdff dff_B_LmyQWHIX7_2(.din(w_dff_B_fJvYJ8zi7_2),.dout(w_dff_B_LmyQWHIX7_2),.clk(gclk));
	jdff dff_B_UmN3Dyph0_2(.din(w_dff_B_LmyQWHIX7_2),.dout(w_dff_B_UmN3Dyph0_2),.clk(gclk));
	jdff dff_B_uTsoFDaG1_2(.din(w_dff_B_UmN3Dyph0_2),.dout(w_dff_B_uTsoFDaG1_2),.clk(gclk));
	jdff dff_B_FpLZbDWC4_2(.din(w_dff_B_uTsoFDaG1_2),.dout(w_dff_B_FpLZbDWC4_2),.clk(gclk));
	jdff dff_B_6dtxSjAr8_2(.din(n1672),.dout(w_dff_B_6dtxSjAr8_2),.clk(gclk));
	jdff dff_B_EuWd9ZeP3_2(.din(w_dff_B_6dtxSjAr8_2),.dout(w_dff_B_EuWd9ZeP3_2),.clk(gclk));
	jdff dff_B_qOayzeZa8_2(.din(w_dff_B_EuWd9ZeP3_2),.dout(w_dff_B_qOayzeZa8_2),.clk(gclk));
	jdff dff_B_oXfcGFna4_2(.din(w_dff_B_qOayzeZa8_2),.dout(w_dff_B_oXfcGFna4_2),.clk(gclk));
	jdff dff_B_f2F0H5Y09_2(.din(w_dff_B_oXfcGFna4_2),.dout(w_dff_B_f2F0H5Y09_2),.clk(gclk));
	jdff dff_B_BPBtebEC6_2(.din(w_dff_B_f2F0H5Y09_2),.dout(w_dff_B_BPBtebEC6_2),.clk(gclk));
	jdff dff_B_OUoVzMya5_2(.din(w_dff_B_BPBtebEC6_2),.dout(w_dff_B_OUoVzMya5_2),.clk(gclk));
	jdff dff_B_t4mGRhEk9_2(.din(w_dff_B_OUoVzMya5_2),.dout(w_dff_B_t4mGRhEk9_2),.clk(gclk));
	jdff dff_B_AmJDgoIR5_2(.din(w_dff_B_t4mGRhEk9_2),.dout(w_dff_B_AmJDgoIR5_2),.clk(gclk));
	jdff dff_B_lxgtwjMq4_2(.din(w_dff_B_AmJDgoIR5_2),.dout(w_dff_B_lxgtwjMq4_2),.clk(gclk));
	jdff dff_B_xSR5WsxF3_2(.din(w_dff_B_lxgtwjMq4_2),.dout(w_dff_B_xSR5WsxF3_2),.clk(gclk));
	jdff dff_B_oAXnSN2Q4_2(.din(w_dff_B_xSR5WsxF3_2),.dout(w_dff_B_oAXnSN2Q4_2),.clk(gclk));
	jdff dff_B_YBJjziKd2_2(.din(w_dff_B_oAXnSN2Q4_2),.dout(w_dff_B_YBJjziKd2_2),.clk(gclk));
	jdff dff_B_IUtx9uST3_2(.din(w_dff_B_YBJjziKd2_2),.dout(w_dff_B_IUtx9uST3_2),.clk(gclk));
	jdff dff_B_ynu59tw81_2(.din(w_dff_B_IUtx9uST3_2),.dout(w_dff_B_ynu59tw81_2),.clk(gclk));
	jdff dff_B_CXdOWRCV6_2(.din(w_dff_B_ynu59tw81_2),.dout(w_dff_B_CXdOWRCV6_2),.clk(gclk));
	jdff dff_B_PAc7A3W79_2(.din(w_dff_B_CXdOWRCV6_2),.dout(w_dff_B_PAc7A3W79_2),.clk(gclk));
	jdff dff_B_1oRHhMWH2_2(.din(w_dff_B_PAc7A3W79_2),.dout(w_dff_B_1oRHhMWH2_2),.clk(gclk));
	jdff dff_B_ratrjSTf6_2(.din(w_dff_B_1oRHhMWH2_2),.dout(w_dff_B_ratrjSTf6_2),.clk(gclk));
	jdff dff_B_tOKyTNL04_2(.din(w_dff_B_ratrjSTf6_2),.dout(w_dff_B_tOKyTNL04_2),.clk(gclk));
	jdff dff_B_OucVIWuq3_2(.din(w_dff_B_tOKyTNL04_2),.dout(w_dff_B_OucVIWuq3_2),.clk(gclk));
	jdff dff_B_898IZUov7_2(.din(w_dff_B_OucVIWuq3_2),.dout(w_dff_B_898IZUov7_2),.clk(gclk));
	jdff dff_B_9m1alUI77_2(.din(w_dff_B_898IZUov7_2),.dout(w_dff_B_9m1alUI77_2),.clk(gclk));
	jdff dff_B_Nx1ICzwB2_2(.din(w_dff_B_9m1alUI77_2),.dout(w_dff_B_Nx1ICzwB2_2),.clk(gclk));
	jdff dff_B_oYuSsp4l1_2(.din(w_dff_B_Nx1ICzwB2_2),.dout(w_dff_B_oYuSsp4l1_2),.clk(gclk));
	jdff dff_B_dsxpN8f92_2(.din(w_dff_B_oYuSsp4l1_2),.dout(w_dff_B_dsxpN8f92_2),.clk(gclk));
	jdff dff_B_3EZMwyX26_2(.din(w_dff_B_dsxpN8f92_2),.dout(w_dff_B_3EZMwyX26_2),.clk(gclk));
	jdff dff_B_ns77EYFo5_2(.din(w_dff_B_3EZMwyX26_2),.dout(w_dff_B_ns77EYFo5_2),.clk(gclk));
	jdff dff_B_YqiDvoCs3_2(.din(w_dff_B_ns77EYFo5_2),.dout(w_dff_B_YqiDvoCs3_2),.clk(gclk));
	jdff dff_B_oOKqRdP05_2(.din(w_dff_B_YqiDvoCs3_2),.dout(w_dff_B_oOKqRdP05_2),.clk(gclk));
	jdff dff_B_r3huhRxb0_2(.din(n1671),.dout(w_dff_B_r3huhRxb0_2),.clk(gclk));
	jdff dff_B_axwawoWk7_1(.din(n1669),.dout(w_dff_B_axwawoWk7_1),.clk(gclk));
	jdff dff_B_pP1zO1dr1_2(.din(n1617),.dout(w_dff_B_pP1zO1dr1_2),.clk(gclk));
	jdff dff_B_1jCzbY4i8_2(.din(w_dff_B_pP1zO1dr1_2),.dout(w_dff_B_1jCzbY4i8_2),.clk(gclk));
	jdff dff_B_zSpTN13E8_2(.din(w_dff_B_1jCzbY4i8_2),.dout(w_dff_B_zSpTN13E8_2),.clk(gclk));
	jdff dff_B_BCucj8Jg2_2(.din(w_dff_B_zSpTN13E8_2),.dout(w_dff_B_BCucj8Jg2_2),.clk(gclk));
	jdff dff_B_x9OfUCI92_2(.din(w_dff_B_BCucj8Jg2_2),.dout(w_dff_B_x9OfUCI92_2),.clk(gclk));
	jdff dff_B_zn8hKTYi2_2(.din(w_dff_B_x9OfUCI92_2),.dout(w_dff_B_zn8hKTYi2_2),.clk(gclk));
	jdff dff_B_WbuKOWZA5_2(.din(w_dff_B_zn8hKTYi2_2),.dout(w_dff_B_WbuKOWZA5_2),.clk(gclk));
	jdff dff_B_x5OgFASA0_2(.din(w_dff_B_WbuKOWZA5_2),.dout(w_dff_B_x5OgFASA0_2),.clk(gclk));
	jdff dff_B_OqcEM6ry9_2(.din(w_dff_B_x5OgFASA0_2),.dout(w_dff_B_OqcEM6ry9_2),.clk(gclk));
	jdff dff_B_VLBYan4f1_2(.din(w_dff_B_OqcEM6ry9_2),.dout(w_dff_B_VLBYan4f1_2),.clk(gclk));
	jdff dff_B_CVeCeV9d8_2(.din(w_dff_B_VLBYan4f1_2),.dout(w_dff_B_CVeCeV9d8_2),.clk(gclk));
	jdff dff_B_AYgZOObA1_2(.din(w_dff_B_CVeCeV9d8_2),.dout(w_dff_B_AYgZOObA1_2),.clk(gclk));
	jdff dff_B_SWGQD5jE1_2(.din(w_dff_B_AYgZOObA1_2),.dout(w_dff_B_SWGQD5jE1_2),.clk(gclk));
	jdff dff_B_8VMFlyWQ0_2(.din(w_dff_B_SWGQD5jE1_2),.dout(w_dff_B_8VMFlyWQ0_2),.clk(gclk));
	jdff dff_B_Wt2wet0t6_2(.din(w_dff_B_8VMFlyWQ0_2),.dout(w_dff_B_Wt2wet0t6_2),.clk(gclk));
	jdff dff_B_DMmIc6Li5_2(.din(w_dff_B_Wt2wet0t6_2),.dout(w_dff_B_DMmIc6Li5_2),.clk(gclk));
	jdff dff_B_17kVzHi07_2(.din(w_dff_B_DMmIc6Li5_2),.dout(w_dff_B_17kVzHi07_2),.clk(gclk));
	jdff dff_B_FWHTRLI31_2(.din(w_dff_B_17kVzHi07_2),.dout(w_dff_B_FWHTRLI31_2),.clk(gclk));
	jdff dff_B_22KYK1pL5_2(.din(w_dff_B_FWHTRLI31_2),.dout(w_dff_B_22KYK1pL5_2),.clk(gclk));
	jdff dff_B_ClQDiSsc0_2(.din(w_dff_B_22KYK1pL5_2),.dout(w_dff_B_ClQDiSsc0_2),.clk(gclk));
	jdff dff_B_yld00TSB7_2(.din(w_dff_B_ClQDiSsc0_2),.dout(w_dff_B_yld00TSB7_2),.clk(gclk));
	jdff dff_B_3sWcS0aT0_2(.din(w_dff_B_yld00TSB7_2),.dout(w_dff_B_3sWcS0aT0_2),.clk(gclk));
	jdff dff_B_32dytsvL2_2(.din(w_dff_B_3sWcS0aT0_2),.dout(w_dff_B_32dytsvL2_2),.clk(gclk));
	jdff dff_B_sRhPOV9Q7_2(.din(w_dff_B_32dytsvL2_2),.dout(w_dff_B_sRhPOV9Q7_2),.clk(gclk));
	jdff dff_B_563zx3iX4_2(.din(w_dff_B_sRhPOV9Q7_2),.dout(w_dff_B_563zx3iX4_2),.clk(gclk));
	jdff dff_B_o1oX2fjh2_2(.din(w_dff_B_563zx3iX4_2),.dout(w_dff_B_o1oX2fjh2_2),.clk(gclk));
	jdff dff_B_GG2ipBND6_2(.din(w_dff_B_o1oX2fjh2_2),.dout(w_dff_B_GG2ipBND6_2),.clk(gclk));
	jdff dff_B_NpD8YZJA9_2(.din(w_dff_B_GG2ipBND6_2),.dout(w_dff_B_NpD8YZJA9_2),.clk(gclk));
	jdff dff_B_KKo5uyzD1_1(.din(n1623),.dout(w_dff_B_KKo5uyzD1_1),.clk(gclk));
	jdff dff_B_fUp5carD2_1(.din(w_dff_B_KKo5uyzD1_1),.dout(w_dff_B_fUp5carD2_1),.clk(gclk));
	jdff dff_B_iuKMDIcm1_2(.din(n1622),.dout(w_dff_B_iuKMDIcm1_2),.clk(gclk));
	jdff dff_B_kjd9Dbyd1_2(.din(w_dff_B_iuKMDIcm1_2),.dout(w_dff_B_kjd9Dbyd1_2),.clk(gclk));
	jdff dff_B_LDfN8eSa4_2(.din(w_dff_B_kjd9Dbyd1_2),.dout(w_dff_B_LDfN8eSa4_2),.clk(gclk));
	jdff dff_B_nb5uT2GN5_2(.din(w_dff_B_LDfN8eSa4_2),.dout(w_dff_B_nb5uT2GN5_2),.clk(gclk));
	jdff dff_B_MLiRERpH6_2(.din(w_dff_B_nb5uT2GN5_2),.dout(w_dff_B_MLiRERpH6_2),.clk(gclk));
	jdff dff_B_CduGgfau2_2(.din(w_dff_B_MLiRERpH6_2),.dout(w_dff_B_CduGgfau2_2),.clk(gclk));
	jdff dff_B_NOSdq8cy0_2(.din(w_dff_B_CduGgfau2_2),.dout(w_dff_B_NOSdq8cy0_2),.clk(gclk));
	jdff dff_B_psunIQm47_2(.din(w_dff_B_NOSdq8cy0_2),.dout(w_dff_B_psunIQm47_2),.clk(gclk));
	jdff dff_B_g2p7kXZc7_2(.din(w_dff_B_psunIQm47_2),.dout(w_dff_B_g2p7kXZc7_2),.clk(gclk));
	jdff dff_B_B9lEuDsJ1_2(.din(w_dff_B_g2p7kXZc7_2),.dout(w_dff_B_B9lEuDsJ1_2),.clk(gclk));
	jdff dff_B_y8oDhhuJ9_2(.din(w_dff_B_B9lEuDsJ1_2),.dout(w_dff_B_y8oDhhuJ9_2),.clk(gclk));
	jdff dff_B_xoodPjTG1_2(.din(w_dff_B_y8oDhhuJ9_2),.dout(w_dff_B_xoodPjTG1_2),.clk(gclk));
	jdff dff_B_0Mxu5Yft5_2(.din(w_dff_B_xoodPjTG1_2),.dout(w_dff_B_0Mxu5Yft5_2),.clk(gclk));
	jdff dff_B_Iwdzmfmy4_2(.din(w_dff_B_0Mxu5Yft5_2),.dout(w_dff_B_Iwdzmfmy4_2),.clk(gclk));
	jdff dff_B_99z39qjD3_2(.din(w_dff_B_Iwdzmfmy4_2),.dout(w_dff_B_99z39qjD3_2),.clk(gclk));
	jdff dff_B_5FhJnfHY4_2(.din(w_dff_B_99z39qjD3_2),.dout(w_dff_B_5FhJnfHY4_2),.clk(gclk));
	jdff dff_B_X2idDRtj5_2(.din(w_dff_B_5FhJnfHY4_2),.dout(w_dff_B_X2idDRtj5_2),.clk(gclk));
	jdff dff_B_XmqUqcaC9_2(.din(w_dff_B_X2idDRtj5_2),.dout(w_dff_B_XmqUqcaC9_2),.clk(gclk));
	jdff dff_B_2fHsdkNh4_2(.din(w_dff_B_XmqUqcaC9_2),.dout(w_dff_B_2fHsdkNh4_2),.clk(gclk));
	jdff dff_B_qjpn0hwI8_2(.din(w_dff_B_2fHsdkNh4_2),.dout(w_dff_B_qjpn0hwI8_2),.clk(gclk));
	jdff dff_B_qObceB4j2_2(.din(w_dff_B_qjpn0hwI8_2),.dout(w_dff_B_qObceB4j2_2),.clk(gclk));
	jdff dff_B_jKouMlbX3_2(.din(w_dff_B_qObceB4j2_2),.dout(w_dff_B_jKouMlbX3_2),.clk(gclk));
	jdff dff_B_SN1cEEHf9_2(.din(w_dff_B_jKouMlbX3_2),.dout(w_dff_B_SN1cEEHf9_2),.clk(gclk));
	jdff dff_B_6h0sUWPv7_2(.din(w_dff_B_SN1cEEHf9_2),.dout(w_dff_B_6h0sUWPv7_2),.clk(gclk));
	jdff dff_B_gw1iOXXp7_2(.din(w_dff_B_6h0sUWPv7_2),.dout(w_dff_B_gw1iOXXp7_2),.clk(gclk));
	jdff dff_B_PiVM0ds34_2(.din(n1621),.dout(w_dff_B_PiVM0ds34_2),.clk(gclk));
	jdff dff_B_AeGB050M3_2(.din(w_dff_B_PiVM0ds34_2),.dout(w_dff_B_AeGB050M3_2),.clk(gclk));
	jdff dff_B_6fe1ZZT72_2(.din(w_dff_B_AeGB050M3_2),.dout(w_dff_B_6fe1ZZT72_2),.clk(gclk));
	jdff dff_B_rbQzXhv49_2(.din(w_dff_B_6fe1ZZT72_2),.dout(w_dff_B_rbQzXhv49_2),.clk(gclk));
	jdff dff_B_vpNtrClQ6_2(.din(w_dff_B_rbQzXhv49_2),.dout(w_dff_B_vpNtrClQ6_2),.clk(gclk));
	jdff dff_B_zvCYuRT76_2(.din(w_dff_B_vpNtrClQ6_2),.dout(w_dff_B_zvCYuRT76_2),.clk(gclk));
	jdff dff_B_6Wx6rueF9_2(.din(w_dff_B_zvCYuRT76_2),.dout(w_dff_B_6Wx6rueF9_2),.clk(gclk));
	jdff dff_B_KywE32Fx1_2(.din(w_dff_B_6Wx6rueF9_2),.dout(w_dff_B_KywE32Fx1_2),.clk(gclk));
	jdff dff_B_1leBmKF44_2(.din(w_dff_B_KywE32Fx1_2),.dout(w_dff_B_1leBmKF44_2),.clk(gclk));
	jdff dff_B_2CqPL4yi0_2(.din(w_dff_B_1leBmKF44_2),.dout(w_dff_B_2CqPL4yi0_2),.clk(gclk));
	jdff dff_B_bMIAaMpA3_2(.din(w_dff_B_2CqPL4yi0_2),.dout(w_dff_B_bMIAaMpA3_2),.clk(gclk));
	jdff dff_B_QnRjZRUk0_2(.din(w_dff_B_bMIAaMpA3_2),.dout(w_dff_B_QnRjZRUk0_2),.clk(gclk));
	jdff dff_B_JEyLHMLm2_2(.din(w_dff_B_QnRjZRUk0_2),.dout(w_dff_B_JEyLHMLm2_2),.clk(gclk));
	jdff dff_B_4cANnGjV0_2(.din(w_dff_B_JEyLHMLm2_2),.dout(w_dff_B_4cANnGjV0_2),.clk(gclk));
	jdff dff_B_BEziTMNN8_2(.din(w_dff_B_4cANnGjV0_2),.dout(w_dff_B_BEziTMNN8_2),.clk(gclk));
	jdff dff_B_HVJ59YLJ0_2(.din(w_dff_B_BEziTMNN8_2),.dout(w_dff_B_HVJ59YLJ0_2),.clk(gclk));
	jdff dff_B_4wvzxoic9_2(.din(w_dff_B_HVJ59YLJ0_2),.dout(w_dff_B_4wvzxoic9_2),.clk(gclk));
	jdff dff_B_BXTrh1J06_2(.din(w_dff_B_4wvzxoic9_2),.dout(w_dff_B_BXTrh1J06_2),.clk(gclk));
	jdff dff_B_xPlDu62I3_2(.din(w_dff_B_BXTrh1J06_2),.dout(w_dff_B_xPlDu62I3_2),.clk(gclk));
	jdff dff_B_Uva3JQDW0_2(.din(w_dff_B_xPlDu62I3_2),.dout(w_dff_B_Uva3JQDW0_2),.clk(gclk));
	jdff dff_B_MluYXu587_2(.din(w_dff_B_Uva3JQDW0_2),.dout(w_dff_B_MluYXu587_2),.clk(gclk));
	jdff dff_B_izJ6VbzU4_2(.din(w_dff_B_MluYXu587_2),.dout(w_dff_B_izJ6VbzU4_2),.clk(gclk));
	jdff dff_B_gvN8qU1Z6_2(.din(w_dff_B_izJ6VbzU4_2),.dout(w_dff_B_gvN8qU1Z6_2),.clk(gclk));
	jdff dff_B_YJrWGonY4_2(.din(w_dff_B_gvN8qU1Z6_2),.dout(w_dff_B_YJrWGonY4_2),.clk(gclk));
	jdff dff_B_IKiF4pOz3_2(.din(w_dff_B_YJrWGonY4_2),.dout(w_dff_B_IKiF4pOz3_2),.clk(gclk));
	jdff dff_B_h1fyl2iW6_2(.din(w_dff_B_IKiF4pOz3_2),.dout(w_dff_B_h1fyl2iW6_2),.clk(gclk));
	jdff dff_B_1PFggV3Q2_2(.din(w_dff_B_h1fyl2iW6_2),.dout(w_dff_B_1PFggV3Q2_2),.clk(gclk));
	jdff dff_B_dfw6ZqK21_2(.din(n1620),.dout(w_dff_B_dfw6ZqK21_2),.clk(gclk));
	jdff dff_B_MNUGWboP9_1(.din(n1618),.dout(w_dff_B_MNUGWboP9_1),.clk(gclk));
	jdff dff_B_0FQo1S0N8_2(.din(n1560),.dout(w_dff_B_0FQo1S0N8_2),.clk(gclk));
	jdff dff_B_0Nobq94l0_2(.din(w_dff_B_0FQo1S0N8_2),.dout(w_dff_B_0Nobq94l0_2),.clk(gclk));
	jdff dff_B_zSUR7HNA1_2(.din(w_dff_B_0Nobq94l0_2),.dout(w_dff_B_zSUR7HNA1_2),.clk(gclk));
	jdff dff_B_xKJKMDGg2_2(.din(w_dff_B_zSUR7HNA1_2),.dout(w_dff_B_xKJKMDGg2_2),.clk(gclk));
	jdff dff_B_E41MIQhv0_2(.din(w_dff_B_xKJKMDGg2_2),.dout(w_dff_B_E41MIQhv0_2),.clk(gclk));
	jdff dff_B_kQUQvBjL9_2(.din(w_dff_B_E41MIQhv0_2),.dout(w_dff_B_kQUQvBjL9_2),.clk(gclk));
	jdff dff_B_HSEdLmDn3_2(.din(w_dff_B_kQUQvBjL9_2),.dout(w_dff_B_HSEdLmDn3_2),.clk(gclk));
	jdff dff_B_kfrP14b15_2(.din(w_dff_B_HSEdLmDn3_2),.dout(w_dff_B_kfrP14b15_2),.clk(gclk));
	jdff dff_B_O4Z4dzXu5_2(.din(w_dff_B_kfrP14b15_2),.dout(w_dff_B_O4Z4dzXu5_2),.clk(gclk));
	jdff dff_B_oXCel9BL5_2(.din(w_dff_B_O4Z4dzXu5_2),.dout(w_dff_B_oXCel9BL5_2),.clk(gclk));
	jdff dff_B_Wn3kuzJG9_2(.din(w_dff_B_oXCel9BL5_2),.dout(w_dff_B_Wn3kuzJG9_2),.clk(gclk));
	jdff dff_B_23vHAYbw4_2(.din(w_dff_B_Wn3kuzJG9_2),.dout(w_dff_B_23vHAYbw4_2),.clk(gclk));
	jdff dff_B_KGTKr7ge0_2(.din(w_dff_B_23vHAYbw4_2),.dout(w_dff_B_KGTKr7ge0_2),.clk(gclk));
	jdff dff_B_BGuARwc99_2(.din(w_dff_B_KGTKr7ge0_2),.dout(w_dff_B_BGuARwc99_2),.clk(gclk));
	jdff dff_B_tfGD2nFJ5_2(.din(w_dff_B_BGuARwc99_2),.dout(w_dff_B_tfGD2nFJ5_2),.clk(gclk));
	jdff dff_B_ueNhaTmM7_2(.din(w_dff_B_tfGD2nFJ5_2),.dout(w_dff_B_ueNhaTmM7_2),.clk(gclk));
	jdff dff_B_mtdXUTWK2_2(.din(w_dff_B_ueNhaTmM7_2),.dout(w_dff_B_mtdXUTWK2_2),.clk(gclk));
	jdff dff_B_5i8l131f1_2(.din(w_dff_B_mtdXUTWK2_2),.dout(w_dff_B_5i8l131f1_2),.clk(gclk));
	jdff dff_B_YXIQprDs0_2(.din(w_dff_B_5i8l131f1_2),.dout(w_dff_B_YXIQprDs0_2),.clk(gclk));
	jdff dff_B_jhqLoEnP6_2(.din(w_dff_B_YXIQprDs0_2),.dout(w_dff_B_jhqLoEnP6_2),.clk(gclk));
	jdff dff_B_Hk8ERIAI0_2(.din(w_dff_B_jhqLoEnP6_2),.dout(w_dff_B_Hk8ERIAI0_2),.clk(gclk));
	jdff dff_B_j1tesltt5_2(.din(w_dff_B_Hk8ERIAI0_2),.dout(w_dff_B_j1tesltt5_2),.clk(gclk));
	jdff dff_B_D39jm4sr1_2(.din(w_dff_B_j1tesltt5_2),.dout(w_dff_B_D39jm4sr1_2),.clk(gclk));
	jdff dff_B_73KkxonX6_2(.din(w_dff_B_D39jm4sr1_2),.dout(w_dff_B_73KkxonX6_2),.clk(gclk));
	jdff dff_B_3is5bFk90_2(.din(w_dff_B_73KkxonX6_2),.dout(w_dff_B_3is5bFk90_2),.clk(gclk));
	jdff dff_B_7mXJf0NA4_1(.din(n1566),.dout(w_dff_B_7mXJf0NA4_1),.clk(gclk));
	jdff dff_B_rttLFnrN8_1(.din(w_dff_B_7mXJf0NA4_1),.dout(w_dff_B_rttLFnrN8_1),.clk(gclk));
	jdff dff_B_20s5XONc9_2(.din(n1565),.dout(w_dff_B_20s5XONc9_2),.clk(gclk));
	jdff dff_B_qHSG2b0c2_2(.din(w_dff_B_20s5XONc9_2),.dout(w_dff_B_qHSG2b0c2_2),.clk(gclk));
	jdff dff_B_ozevfPr46_2(.din(w_dff_B_qHSG2b0c2_2),.dout(w_dff_B_ozevfPr46_2),.clk(gclk));
	jdff dff_B_tkztgueh7_2(.din(w_dff_B_ozevfPr46_2),.dout(w_dff_B_tkztgueh7_2),.clk(gclk));
	jdff dff_B_uIfNoRPO2_2(.din(w_dff_B_tkztgueh7_2),.dout(w_dff_B_uIfNoRPO2_2),.clk(gclk));
	jdff dff_B_kRscPPRT2_2(.din(w_dff_B_uIfNoRPO2_2),.dout(w_dff_B_kRscPPRT2_2),.clk(gclk));
	jdff dff_B_KhBHrXpY8_2(.din(w_dff_B_kRscPPRT2_2),.dout(w_dff_B_KhBHrXpY8_2),.clk(gclk));
	jdff dff_B_6xGnlLq75_2(.din(w_dff_B_KhBHrXpY8_2),.dout(w_dff_B_6xGnlLq75_2),.clk(gclk));
	jdff dff_B_dY5jxuO90_2(.din(w_dff_B_6xGnlLq75_2),.dout(w_dff_B_dY5jxuO90_2),.clk(gclk));
	jdff dff_B_D9bl3EcE9_2(.din(w_dff_B_dY5jxuO90_2),.dout(w_dff_B_D9bl3EcE9_2),.clk(gclk));
	jdff dff_B_XYcQzRBz0_2(.din(w_dff_B_D9bl3EcE9_2),.dout(w_dff_B_XYcQzRBz0_2),.clk(gclk));
	jdff dff_B_URmY6v2R1_2(.din(w_dff_B_XYcQzRBz0_2),.dout(w_dff_B_URmY6v2R1_2),.clk(gclk));
	jdff dff_B_sRD6j7Au3_2(.din(w_dff_B_URmY6v2R1_2),.dout(w_dff_B_sRD6j7Au3_2),.clk(gclk));
	jdff dff_B_qvKa0wlw2_2(.din(w_dff_B_sRD6j7Au3_2),.dout(w_dff_B_qvKa0wlw2_2),.clk(gclk));
	jdff dff_B_iVO4tvig4_2(.din(w_dff_B_qvKa0wlw2_2),.dout(w_dff_B_iVO4tvig4_2),.clk(gclk));
	jdff dff_B_IndCUCZF0_2(.din(w_dff_B_iVO4tvig4_2),.dout(w_dff_B_IndCUCZF0_2),.clk(gclk));
	jdff dff_B_TUXIBF0o1_2(.din(w_dff_B_IndCUCZF0_2),.dout(w_dff_B_TUXIBF0o1_2),.clk(gclk));
	jdff dff_B_cTJkwEs64_2(.din(w_dff_B_TUXIBF0o1_2),.dout(w_dff_B_cTJkwEs64_2),.clk(gclk));
	jdff dff_B_tHwxoFyi4_2(.din(w_dff_B_cTJkwEs64_2),.dout(w_dff_B_tHwxoFyi4_2),.clk(gclk));
	jdff dff_B_UMOLD7XV5_2(.din(w_dff_B_tHwxoFyi4_2),.dout(w_dff_B_UMOLD7XV5_2),.clk(gclk));
	jdff dff_B_LxCUjF5H4_2(.din(w_dff_B_UMOLD7XV5_2),.dout(w_dff_B_LxCUjF5H4_2),.clk(gclk));
	jdff dff_B_eNP0hdtM1_2(.din(w_dff_B_LxCUjF5H4_2),.dout(w_dff_B_eNP0hdtM1_2),.clk(gclk));
	jdff dff_B_At0fZjz30_2(.din(n1564),.dout(w_dff_B_At0fZjz30_2),.clk(gclk));
	jdff dff_B_A8uaYMKH2_2(.din(w_dff_B_At0fZjz30_2),.dout(w_dff_B_A8uaYMKH2_2),.clk(gclk));
	jdff dff_B_9gSPDxPc3_2(.din(w_dff_B_A8uaYMKH2_2),.dout(w_dff_B_9gSPDxPc3_2),.clk(gclk));
	jdff dff_B_djnkdzhD1_2(.din(w_dff_B_9gSPDxPc3_2),.dout(w_dff_B_djnkdzhD1_2),.clk(gclk));
	jdff dff_B_RZ6YHp8E5_2(.din(w_dff_B_djnkdzhD1_2),.dout(w_dff_B_RZ6YHp8E5_2),.clk(gclk));
	jdff dff_B_MrqTEaHc6_2(.din(w_dff_B_RZ6YHp8E5_2),.dout(w_dff_B_MrqTEaHc6_2),.clk(gclk));
	jdff dff_B_ev7Cdmy02_2(.din(w_dff_B_MrqTEaHc6_2),.dout(w_dff_B_ev7Cdmy02_2),.clk(gclk));
	jdff dff_B_COY2pKfh3_2(.din(w_dff_B_ev7Cdmy02_2),.dout(w_dff_B_COY2pKfh3_2),.clk(gclk));
	jdff dff_B_QxQ2Sil13_2(.din(w_dff_B_COY2pKfh3_2),.dout(w_dff_B_QxQ2Sil13_2),.clk(gclk));
	jdff dff_B_aiUSp1hR8_2(.din(w_dff_B_QxQ2Sil13_2),.dout(w_dff_B_aiUSp1hR8_2),.clk(gclk));
	jdff dff_B_QHXE6YZV1_2(.din(w_dff_B_aiUSp1hR8_2),.dout(w_dff_B_QHXE6YZV1_2),.clk(gclk));
	jdff dff_B_9wZfYbvL5_2(.din(w_dff_B_QHXE6YZV1_2),.dout(w_dff_B_9wZfYbvL5_2),.clk(gclk));
	jdff dff_B_uyhzLsEX9_2(.din(w_dff_B_9wZfYbvL5_2),.dout(w_dff_B_uyhzLsEX9_2),.clk(gclk));
	jdff dff_B_sgHepmNT8_2(.din(w_dff_B_uyhzLsEX9_2),.dout(w_dff_B_sgHepmNT8_2),.clk(gclk));
	jdff dff_B_NKZjq98n6_2(.din(w_dff_B_sgHepmNT8_2),.dout(w_dff_B_NKZjq98n6_2),.clk(gclk));
	jdff dff_B_eoCahL8F1_2(.din(w_dff_B_NKZjq98n6_2),.dout(w_dff_B_eoCahL8F1_2),.clk(gclk));
	jdff dff_B_nTkXefiU5_2(.din(w_dff_B_eoCahL8F1_2),.dout(w_dff_B_nTkXefiU5_2),.clk(gclk));
	jdff dff_B_MIMdLjjW5_2(.din(w_dff_B_nTkXefiU5_2),.dout(w_dff_B_MIMdLjjW5_2),.clk(gclk));
	jdff dff_B_lqViAUl30_2(.din(w_dff_B_MIMdLjjW5_2),.dout(w_dff_B_lqViAUl30_2),.clk(gclk));
	jdff dff_B_BZLKrAKe3_2(.din(w_dff_B_lqViAUl30_2),.dout(w_dff_B_BZLKrAKe3_2),.clk(gclk));
	jdff dff_B_Vh0D3MO12_2(.din(w_dff_B_BZLKrAKe3_2),.dout(w_dff_B_Vh0D3MO12_2),.clk(gclk));
	jdff dff_B_4hr0prvr4_2(.din(w_dff_B_Vh0D3MO12_2),.dout(w_dff_B_4hr0prvr4_2),.clk(gclk));
	jdff dff_B_XSo3QIbe5_2(.din(w_dff_B_4hr0prvr4_2),.dout(w_dff_B_XSo3QIbe5_2),.clk(gclk));
	jdff dff_B_SMT7j2uL7_2(.din(w_dff_B_XSo3QIbe5_2),.dout(w_dff_B_SMT7j2uL7_2),.clk(gclk));
	jdff dff_B_Tq1QvZat2_2(.din(n1563),.dout(w_dff_B_Tq1QvZat2_2),.clk(gclk));
	jdff dff_B_UvPqCIej8_1(.din(n1561),.dout(w_dff_B_UvPqCIej8_1),.clk(gclk));
	jdff dff_B_W4KPgvEX4_2(.din(n1496),.dout(w_dff_B_W4KPgvEX4_2),.clk(gclk));
	jdff dff_B_Uj9cySuM9_2(.din(w_dff_B_W4KPgvEX4_2),.dout(w_dff_B_Uj9cySuM9_2),.clk(gclk));
	jdff dff_B_CUMaRmay7_2(.din(w_dff_B_Uj9cySuM9_2),.dout(w_dff_B_CUMaRmay7_2),.clk(gclk));
	jdff dff_B_pT4qGwsF0_2(.din(w_dff_B_CUMaRmay7_2),.dout(w_dff_B_pT4qGwsF0_2),.clk(gclk));
	jdff dff_B_TvVosUeW1_2(.din(w_dff_B_pT4qGwsF0_2),.dout(w_dff_B_TvVosUeW1_2),.clk(gclk));
	jdff dff_B_eA7Hi7LT6_2(.din(w_dff_B_TvVosUeW1_2),.dout(w_dff_B_eA7Hi7LT6_2),.clk(gclk));
	jdff dff_B_ngp5YqPy1_2(.din(w_dff_B_eA7Hi7LT6_2),.dout(w_dff_B_ngp5YqPy1_2),.clk(gclk));
	jdff dff_B_F1D5UxXN3_2(.din(w_dff_B_ngp5YqPy1_2),.dout(w_dff_B_F1D5UxXN3_2),.clk(gclk));
	jdff dff_B_JyZ1M5lM7_2(.din(w_dff_B_F1D5UxXN3_2),.dout(w_dff_B_JyZ1M5lM7_2),.clk(gclk));
	jdff dff_B_D0oT6NFZ3_2(.din(w_dff_B_JyZ1M5lM7_2),.dout(w_dff_B_D0oT6NFZ3_2),.clk(gclk));
	jdff dff_B_96Iv5nAP6_2(.din(w_dff_B_D0oT6NFZ3_2),.dout(w_dff_B_96Iv5nAP6_2),.clk(gclk));
	jdff dff_B_iiEZY4z92_2(.din(w_dff_B_96Iv5nAP6_2),.dout(w_dff_B_iiEZY4z92_2),.clk(gclk));
	jdff dff_B_74D5P7Ff4_2(.din(w_dff_B_iiEZY4z92_2),.dout(w_dff_B_74D5P7Ff4_2),.clk(gclk));
	jdff dff_B_l8YfPTvn9_2(.din(w_dff_B_74D5P7Ff4_2),.dout(w_dff_B_l8YfPTvn9_2),.clk(gclk));
	jdff dff_B_4li1DH5p5_2(.din(w_dff_B_l8YfPTvn9_2),.dout(w_dff_B_4li1DH5p5_2),.clk(gclk));
	jdff dff_B_fvkDwzAC3_2(.din(w_dff_B_4li1DH5p5_2),.dout(w_dff_B_fvkDwzAC3_2),.clk(gclk));
	jdff dff_B_qyBezgsw6_2(.din(w_dff_B_fvkDwzAC3_2),.dout(w_dff_B_qyBezgsw6_2),.clk(gclk));
	jdff dff_B_NijD4bqu9_2(.din(w_dff_B_qyBezgsw6_2),.dout(w_dff_B_NijD4bqu9_2),.clk(gclk));
	jdff dff_B_pIolcipT8_2(.din(w_dff_B_NijD4bqu9_2),.dout(w_dff_B_pIolcipT8_2),.clk(gclk));
	jdff dff_B_VJZIoWdv9_2(.din(w_dff_B_pIolcipT8_2),.dout(w_dff_B_VJZIoWdv9_2),.clk(gclk));
	jdff dff_B_XNvcYRId0_2(.din(w_dff_B_VJZIoWdv9_2),.dout(w_dff_B_XNvcYRId0_2),.clk(gclk));
	jdff dff_B_srWxmUGH1_2(.din(w_dff_B_XNvcYRId0_2),.dout(w_dff_B_srWxmUGH1_2),.clk(gclk));
	jdff dff_B_ckPjZXWm5_1(.din(n1502),.dout(w_dff_B_ckPjZXWm5_1),.clk(gclk));
	jdff dff_B_H9FA1TvV4_1(.din(w_dff_B_ckPjZXWm5_1),.dout(w_dff_B_H9FA1TvV4_1),.clk(gclk));
	jdff dff_B_tXZbOlXK6_2(.din(n1501),.dout(w_dff_B_tXZbOlXK6_2),.clk(gclk));
	jdff dff_B_Jwe3YR9W9_2(.din(w_dff_B_tXZbOlXK6_2),.dout(w_dff_B_Jwe3YR9W9_2),.clk(gclk));
	jdff dff_B_uPHo45gm7_2(.din(w_dff_B_Jwe3YR9W9_2),.dout(w_dff_B_uPHo45gm7_2),.clk(gclk));
	jdff dff_B_kY3p7xUl8_2(.din(w_dff_B_uPHo45gm7_2),.dout(w_dff_B_kY3p7xUl8_2),.clk(gclk));
	jdff dff_B_nsmmMEq34_2(.din(w_dff_B_kY3p7xUl8_2),.dout(w_dff_B_nsmmMEq34_2),.clk(gclk));
	jdff dff_B_V35ZtRIk6_2(.din(w_dff_B_nsmmMEq34_2),.dout(w_dff_B_V35ZtRIk6_2),.clk(gclk));
	jdff dff_B_l54mtnv53_2(.din(w_dff_B_V35ZtRIk6_2),.dout(w_dff_B_l54mtnv53_2),.clk(gclk));
	jdff dff_B_VWcvLOD40_2(.din(w_dff_B_l54mtnv53_2),.dout(w_dff_B_VWcvLOD40_2),.clk(gclk));
	jdff dff_B_jAqZAYch5_2(.din(w_dff_B_VWcvLOD40_2),.dout(w_dff_B_jAqZAYch5_2),.clk(gclk));
	jdff dff_B_eLy6O99I6_2(.din(w_dff_B_jAqZAYch5_2),.dout(w_dff_B_eLy6O99I6_2),.clk(gclk));
	jdff dff_B_WG0M3gtT3_2(.din(w_dff_B_eLy6O99I6_2),.dout(w_dff_B_WG0M3gtT3_2),.clk(gclk));
	jdff dff_B_znoe0lDQ7_2(.din(w_dff_B_WG0M3gtT3_2),.dout(w_dff_B_znoe0lDQ7_2),.clk(gclk));
	jdff dff_B_zGe1Xepb8_2(.din(w_dff_B_znoe0lDQ7_2),.dout(w_dff_B_zGe1Xepb8_2),.clk(gclk));
	jdff dff_B_SFrvPMuE3_2(.din(w_dff_B_zGe1Xepb8_2),.dout(w_dff_B_SFrvPMuE3_2),.clk(gclk));
	jdff dff_B_zY0wbfHt5_2(.din(w_dff_B_SFrvPMuE3_2),.dout(w_dff_B_zY0wbfHt5_2),.clk(gclk));
	jdff dff_B_bJHjr5z51_2(.din(w_dff_B_zY0wbfHt5_2),.dout(w_dff_B_bJHjr5z51_2),.clk(gclk));
	jdff dff_B_j7mYsTgd0_2(.din(w_dff_B_bJHjr5z51_2),.dout(w_dff_B_j7mYsTgd0_2),.clk(gclk));
	jdff dff_B_mA9KAMsF1_2(.din(w_dff_B_j7mYsTgd0_2),.dout(w_dff_B_mA9KAMsF1_2),.clk(gclk));
	jdff dff_B_iQjh87NT6_2(.din(w_dff_B_mA9KAMsF1_2),.dout(w_dff_B_iQjh87NT6_2),.clk(gclk));
	jdff dff_B_jvcr6p3n7_2(.din(n1500),.dout(w_dff_B_jvcr6p3n7_2),.clk(gclk));
	jdff dff_B_xNRjuCEd0_2(.din(w_dff_B_jvcr6p3n7_2),.dout(w_dff_B_xNRjuCEd0_2),.clk(gclk));
	jdff dff_B_VgK0fkjq6_2(.din(w_dff_B_xNRjuCEd0_2),.dout(w_dff_B_VgK0fkjq6_2),.clk(gclk));
	jdff dff_B_aVSHeBJJ3_2(.din(w_dff_B_VgK0fkjq6_2),.dout(w_dff_B_aVSHeBJJ3_2),.clk(gclk));
	jdff dff_B_SZCVgi9k8_2(.din(w_dff_B_aVSHeBJJ3_2),.dout(w_dff_B_SZCVgi9k8_2),.clk(gclk));
	jdff dff_B_HSgFmTUo9_2(.din(w_dff_B_SZCVgi9k8_2),.dout(w_dff_B_HSgFmTUo9_2),.clk(gclk));
	jdff dff_B_aCQJyS167_2(.din(w_dff_B_HSgFmTUo9_2),.dout(w_dff_B_aCQJyS167_2),.clk(gclk));
	jdff dff_B_EEAkD4rO9_2(.din(w_dff_B_aCQJyS167_2),.dout(w_dff_B_EEAkD4rO9_2),.clk(gclk));
	jdff dff_B_FPsrj22g8_2(.din(w_dff_B_EEAkD4rO9_2),.dout(w_dff_B_FPsrj22g8_2),.clk(gclk));
	jdff dff_B_Yvglu0PZ3_2(.din(w_dff_B_FPsrj22g8_2),.dout(w_dff_B_Yvglu0PZ3_2),.clk(gclk));
	jdff dff_B_vEj4vuNa3_2(.din(w_dff_B_Yvglu0PZ3_2),.dout(w_dff_B_vEj4vuNa3_2),.clk(gclk));
	jdff dff_B_2ck013Mi6_2(.din(w_dff_B_vEj4vuNa3_2),.dout(w_dff_B_2ck013Mi6_2),.clk(gclk));
	jdff dff_B_g1lbKyY67_2(.din(w_dff_B_2ck013Mi6_2),.dout(w_dff_B_g1lbKyY67_2),.clk(gclk));
	jdff dff_B_h71LZwRD9_2(.din(w_dff_B_g1lbKyY67_2),.dout(w_dff_B_h71LZwRD9_2),.clk(gclk));
	jdff dff_B_jfWebrkp7_2(.din(w_dff_B_h71LZwRD9_2),.dout(w_dff_B_jfWebrkp7_2),.clk(gclk));
	jdff dff_B_RB8ktwhb8_2(.din(w_dff_B_jfWebrkp7_2),.dout(w_dff_B_RB8ktwhb8_2),.clk(gclk));
	jdff dff_B_wvrPjaGA6_2(.din(w_dff_B_RB8ktwhb8_2),.dout(w_dff_B_wvrPjaGA6_2),.clk(gclk));
	jdff dff_B_dOxhdNAd2_2(.din(w_dff_B_wvrPjaGA6_2),.dout(w_dff_B_dOxhdNAd2_2),.clk(gclk));
	jdff dff_B_gC1xw0672_2(.din(w_dff_B_dOxhdNAd2_2),.dout(w_dff_B_gC1xw0672_2),.clk(gclk));
	jdff dff_B_ucxniJKP3_2(.din(w_dff_B_gC1xw0672_2),.dout(w_dff_B_ucxniJKP3_2),.clk(gclk));
	jdff dff_B_GvYE6x427_2(.din(w_dff_B_ucxniJKP3_2),.dout(w_dff_B_GvYE6x427_2),.clk(gclk));
	jdff dff_B_BdadzOvs7_2(.din(n1499),.dout(w_dff_B_BdadzOvs7_2),.clk(gclk));
	jdff dff_B_UAj1SjrY2_1(.din(n1497),.dout(w_dff_B_UAj1SjrY2_1),.clk(gclk));
	jdff dff_B_ZURcfvPQ0_2(.din(n1425),.dout(w_dff_B_ZURcfvPQ0_2),.clk(gclk));
	jdff dff_B_WkGbWWub4_2(.din(w_dff_B_ZURcfvPQ0_2),.dout(w_dff_B_WkGbWWub4_2),.clk(gclk));
	jdff dff_B_eCMV28ii0_2(.din(w_dff_B_WkGbWWub4_2),.dout(w_dff_B_eCMV28ii0_2),.clk(gclk));
	jdff dff_B_YJh8Mtet8_2(.din(w_dff_B_eCMV28ii0_2),.dout(w_dff_B_YJh8Mtet8_2),.clk(gclk));
	jdff dff_B_1GAI9xrm6_2(.din(w_dff_B_YJh8Mtet8_2),.dout(w_dff_B_1GAI9xrm6_2),.clk(gclk));
	jdff dff_B_vAw4yNn23_2(.din(w_dff_B_1GAI9xrm6_2),.dout(w_dff_B_vAw4yNn23_2),.clk(gclk));
	jdff dff_B_Zz6DcGaK2_2(.din(w_dff_B_vAw4yNn23_2),.dout(w_dff_B_Zz6DcGaK2_2),.clk(gclk));
	jdff dff_B_fqzJZH849_2(.din(w_dff_B_Zz6DcGaK2_2),.dout(w_dff_B_fqzJZH849_2),.clk(gclk));
	jdff dff_B_kwB6LRBl7_2(.din(w_dff_B_fqzJZH849_2),.dout(w_dff_B_kwB6LRBl7_2),.clk(gclk));
	jdff dff_B_GQsCX0NR3_2(.din(w_dff_B_kwB6LRBl7_2),.dout(w_dff_B_GQsCX0NR3_2),.clk(gclk));
	jdff dff_B_TipRNKVT4_2(.din(w_dff_B_GQsCX0NR3_2),.dout(w_dff_B_TipRNKVT4_2),.clk(gclk));
	jdff dff_B_2gtpBNs35_2(.din(w_dff_B_TipRNKVT4_2),.dout(w_dff_B_2gtpBNs35_2),.clk(gclk));
	jdff dff_B_Flb76xP35_2(.din(w_dff_B_2gtpBNs35_2),.dout(w_dff_B_Flb76xP35_2),.clk(gclk));
	jdff dff_B_d1ssITac7_2(.din(w_dff_B_Flb76xP35_2),.dout(w_dff_B_d1ssITac7_2),.clk(gclk));
	jdff dff_B_SlYxEG5Y8_2(.din(w_dff_B_d1ssITac7_2),.dout(w_dff_B_SlYxEG5Y8_2),.clk(gclk));
	jdff dff_B_FIf92ijf8_2(.din(w_dff_B_SlYxEG5Y8_2),.dout(w_dff_B_FIf92ijf8_2),.clk(gclk));
	jdff dff_B_S3uJgSCE1_2(.din(w_dff_B_FIf92ijf8_2),.dout(w_dff_B_S3uJgSCE1_2),.clk(gclk));
	jdff dff_B_zUWqdC8v8_2(.din(w_dff_B_S3uJgSCE1_2),.dout(w_dff_B_zUWqdC8v8_2),.clk(gclk));
	jdff dff_B_m2NcjGE91_2(.din(w_dff_B_zUWqdC8v8_2),.dout(w_dff_B_m2NcjGE91_2),.clk(gclk));
	jdff dff_B_oNuiEidf0_1(.din(n1431),.dout(w_dff_B_oNuiEidf0_1),.clk(gclk));
	jdff dff_B_vUihC5lP1_1(.din(w_dff_B_oNuiEidf0_1),.dout(w_dff_B_vUihC5lP1_1),.clk(gclk));
	jdff dff_B_6ZZjHziA1_2(.din(n1430),.dout(w_dff_B_6ZZjHziA1_2),.clk(gclk));
	jdff dff_B_G0LAQaai6_2(.din(w_dff_B_6ZZjHziA1_2),.dout(w_dff_B_G0LAQaai6_2),.clk(gclk));
	jdff dff_B_MHj26KEy0_2(.din(w_dff_B_G0LAQaai6_2),.dout(w_dff_B_MHj26KEy0_2),.clk(gclk));
	jdff dff_B_PfTNKA7O1_2(.din(w_dff_B_MHj26KEy0_2),.dout(w_dff_B_PfTNKA7O1_2),.clk(gclk));
	jdff dff_B_6n8B0bJc6_2(.din(w_dff_B_PfTNKA7O1_2),.dout(w_dff_B_6n8B0bJc6_2),.clk(gclk));
	jdff dff_B_u7Hog3wX1_2(.din(w_dff_B_6n8B0bJc6_2),.dout(w_dff_B_u7Hog3wX1_2),.clk(gclk));
	jdff dff_B_KpBUQ8wl7_2(.din(w_dff_B_u7Hog3wX1_2),.dout(w_dff_B_KpBUQ8wl7_2),.clk(gclk));
	jdff dff_B_46KAuIWD5_2(.din(w_dff_B_KpBUQ8wl7_2),.dout(w_dff_B_46KAuIWD5_2),.clk(gclk));
	jdff dff_B_rHoMFQgi8_2(.din(w_dff_B_46KAuIWD5_2),.dout(w_dff_B_rHoMFQgi8_2),.clk(gclk));
	jdff dff_B_2fW30ZPh7_2(.din(w_dff_B_rHoMFQgi8_2),.dout(w_dff_B_2fW30ZPh7_2),.clk(gclk));
	jdff dff_B_z83qEetY7_2(.din(w_dff_B_2fW30ZPh7_2),.dout(w_dff_B_z83qEetY7_2),.clk(gclk));
	jdff dff_B_vZjcRGP98_2(.din(w_dff_B_z83qEetY7_2),.dout(w_dff_B_vZjcRGP98_2),.clk(gclk));
	jdff dff_B_9XesZivJ2_2(.din(w_dff_B_vZjcRGP98_2),.dout(w_dff_B_9XesZivJ2_2),.clk(gclk));
	jdff dff_B_NMAcy3rD7_2(.din(w_dff_B_9XesZivJ2_2),.dout(w_dff_B_NMAcy3rD7_2),.clk(gclk));
	jdff dff_B_qFFFDnug7_2(.din(w_dff_B_NMAcy3rD7_2),.dout(w_dff_B_qFFFDnug7_2),.clk(gclk));
	jdff dff_B_UX6p194Y7_2(.din(w_dff_B_qFFFDnug7_2),.dout(w_dff_B_UX6p194Y7_2),.clk(gclk));
	jdff dff_B_k6kywRH35_2(.din(n1429),.dout(w_dff_B_k6kywRH35_2),.clk(gclk));
	jdff dff_B_D0jKwcVk4_2(.din(w_dff_B_k6kywRH35_2),.dout(w_dff_B_D0jKwcVk4_2),.clk(gclk));
	jdff dff_B_wzsN9kEW7_2(.din(w_dff_B_D0jKwcVk4_2),.dout(w_dff_B_wzsN9kEW7_2),.clk(gclk));
	jdff dff_B_8acDGkWu4_2(.din(w_dff_B_wzsN9kEW7_2),.dout(w_dff_B_8acDGkWu4_2),.clk(gclk));
	jdff dff_B_z7WPkZ804_2(.din(w_dff_B_8acDGkWu4_2),.dout(w_dff_B_z7WPkZ804_2),.clk(gclk));
	jdff dff_B_2ZlohMTO4_2(.din(w_dff_B_z7WPkZ804_2),.dout(w_dff_B_2ZlohMTO4_2),.clk(gclk));
	jdff dff_B_JqcmM7KS0_2(.din(w_dff_B_2ZlohMTO4_2),.dout(w_dff_B_JqcmM7KS0_2),.clk(gclk));
	jdff dff_B_vyg3BJSh4_2(.din(w_dff_B_JqcmM7KS0_2),.dout(w_dff_B_vyg3BJSh4_2),.clk(gclk));
	jdff dff_B_T23OO0co1_2(.din(w_dff_B_vyg3BJSh4_2),.dout(w_dff_B_T23OO0co1_2),.clk(gclk));
	jdff dff_B_1Ehd7qne6_2(.din(w_dff_B_T23OO0co1_2),.dout(w_dff_B_1Ehd7qne6_2),.clk(gclk));
	jdff dff_B_wqOXyipe2_2(.din(w_dff_B_1Ehd7qne6_2),.dout(w_dff_B_wqOXyipe2_2),.clk(gclk));
	jdff dff_B_g2MKs5hz6_2(.din(w_dff_B_wqOXyipe2_2),.dout(w_dff_B_g2MKs5hz6_2),.clk(gclk));
	jdff dff_B_YQ2qn2jF6_2(.din(w_dff_B_g2MKs5hz6_2),.dout(w_dff_B_YQ2qn2jF6_2),.clk(gclk));
	jdff dff_B_sQN5eiBb7_2(.din(w_dff_B_YQ2qn2jF6_2),.dout(w_dff_B_sQN5eiBb7_2),.clk(gclk));
	jdff dff_B_ZFtk1Kng5_2(.din(w_dff_B_sQN5eiBb7_2),.dout(w_dff_B_ZFtk1Kng5_2),.clk(gclk));
	jdff dff_B_fPYMB1gx9_2(.din(w_dff_B_ZFtk1Kng5_2),.dout(w_dff_B_fPYMB1gx9_2),.clk(gclk));
	jdff dff_B_YkNbzws61_2(.din(w_dff_B_fPYMB1gx9_2),.dout(w_dff_B_YkNbzws61_2),.clk(gclk));
	jdff dff_B_NZ65v4E38_2(.din(w_dff_B_YkNbzws61_2),.dout(w_dff_B_NZ65v4E38_2),.clk(gclk));
	jdff dff_B_KiPv2Y083_2(.din(n1428),.dout(w_dff_B_KiPv2Y083_2),.clk(gclk));
	jdff dff_B_JOlWKl9O1_1(.din(n1426),.dout(w_dff_B_JOlWKl9O1_1),.clk(gclk));
	jdff dff_B_XfLYnpdF6_2(.din(n1347),.dout(w_dff_B_XfLYnpdF6_2),.clk(gclk));
	jdff dff_B_hcghk9XZ7_2(.din(w_dff_B_XfLYnpdF6_2),.dout(w_dff_B_hcghk9XZ7_2),.clk(gclk));
	jdff dff_B_NsWxy5j11_2(.din(w_dff_B_hcghk9XZ7_2),.dout(w_dff_B_NsWxy5j11_2),.clk(gclk));
	jdff dff_B_6f6rUad83_2(.din(w_dff_B_NsWxy5j11_2),.dout(w_dff_B_6f6rUad83_2),.clk(gclk));
	jdff dff_B_ZicVVwmB4_2(.din(w_dff_B_6f6rUad83_2),.dout(w_dff_B_ZicVVwmB4_2),.clk(gclk));
	jdff dff_B_GQ6zQRTI9_2(.din(w_dff_B_ZicVVwmB4_2),.dout(w_dff_B_GQ6zQRTI9_2),.clk(gclk));
	jdff dff_B_iOcbgWV56_2(.din(w_dff_B_GQ6zQRTI9_2),.dout(w_dff_B_iOcbgWV56_2),.clk(gclk));
	jdff dff_B_sSVQtGts7_2(.din(w_dff_B_iOcbgWV56_2),.dout(w_dff_B_sSVQtGts7_2),.clk(gclk));
	jdff dff_B_sy4tdcVL2_2(.din(w_dff_B_sSVQtGts7_2),.dout(w_dff_B_sy4tdcVL2_2),.clk(gclk));
	jdff dff_B_UeJXBPEt6_2(.din(w_dff_B_sy4tdcVL2_2),.dout(w_dff_B_UeJXBPEt6_2),.clk(gclk));
	jdff dff_B_GS14vH2t8_2(.din(w_dff_B_UeJXBPEt6_2),.dout(w_dff_B_GS14vH2t8_2),.clk(gclk));
	jdff dff_B_xNa5kF7g2_2(.din(w_dff_B_GS14vH2t8_2),.dout(w_dff_B_xNa5kF7g2_2),.clk(gclk));
	jdff dff_B_wKKe9xNQ8_2(.din(w_dff_B_xNa5kF7g2_2),.dout(w_dff_B_wKKe9xNQ8_2),.clk(gclk));
	jdff dff_B_hfWUd8FK7_2(.din(w_dff_B_wKKe9xNQ8_2),.dout(w_dff_B_hfWUd8FK7_2),.clk(gclk));
	jdff dff_B_3fmDMV6q8_2(.din(w_dff_B_hfWUd8FK7_2),.dout(w_dff_B_3fmDMV6q8_2),.clk(gclk));
	jdff dff_B_QZg7MbcJ4_2(.din(w_dff_B_3fmDMV6q8_2),.dout(w_dff_B_QZg7MbcJ4_2),.clk(gclk));
	jdff dff_B_Fhdnx1eb8_1(.din(n1353),.dout(w_dff_B_Fhdnx1eb8_1),.clk(gclk));
	jdff dff_B_64BkNosx3_1(.din(w_dff_B_Fhdnx1eb8_1),.dout(w_dff_B_64BkNosx3_1),.clk(gclk));
	jdff dff_B_AFSW1rJM9_2(.din(n1352),.dout(w_dff_B_AFSW1rJM9_2),.clk(gclk));
	jdff dff_B_Lt57vjEl0_2(.din(w_dff_B_AFSW1rJM9_2),.dout(w_dff_B_Lt57vjEl0_2),.clk(gclk));
	jdff dff_B_snHSZHEI1_2(.din(w_dff_B_Lt57vjEl0_2),.dout(w_dff_B_snHSZHEI1_2),.clk(gclk));
	jdff dff_B_dSD9j1M32_2(.din(w_dff_B_snHSZHEI1_2),.dout(w_dff_B_dSD9j1M32_2),.clk(gclk));
	jdff dff_B_wVcQnGcO0_2(.din(w_dff_B_dSD9j1M32_2),.dout(w_dff_B_wVcQnGcO0_2),.clk(gclk));
	jdff dff_B_puNNTyc77_2(.din(w_dff_B_wVcQnGcO0_2),.dout(w_dff_B_puNNTyc77_2),.clk(gclk));
	jdff dff_B_yWjKXj6o8_2(.din(w_dff_B_puNNTyc77_2),.dout(w_dff_B_yWjKXj6o8_2),.clk(gclk));
	jdff dff_B_KDSMyLue3_2(.din(w_dff_B_yWjKXj6o8_2),.dout(w_dff_B_KDSMyLue3_2),.clk(gclk));
	jdff dff_B_CgYGKt9D4_2(.din(w_dff_B_KDSMyLue3_2),.dout(w_dff_B_CgYGKt9D4_2),.clk(gclk));
	jdff dff_B_zcbSCr4D8_2(.din(w_dff_B_CgYGKt9D4_2),.dout(w_dff_B_zcbSCr4D8_2),.clk(gclk));
	jdff dff_B_uJt3UDUC2_2(.din(w_dff_B_zcbSCr4D8_2),.dout(w_dff_B_uJt3UDUC2_2),.clk(gclk));
	jdff dff_B_l0mW5TPC9_2(.din(w_dff_B_uJt3UDUC2_2),.dout(w_dff_B_l0mW5TPC9_2),.clk(gclk));
	jdff dff_B_WYj5ns8X9_2(.din(w_dff_B_l0mW5TPC9_2),.dout(w_dff_B_WYj5ns8X9_2),.clk(gclk));
	jdff dff_B_wvtTIw738_2(.din(n1351),.dout(w_dff_B_wvtTIw738_2),.clk(gclk));
	jdff dff_B_C1YSRQ7g6_2(.din(w_dff_B_wvtTIw738_2),.dout(w_dff_B_C1YSRQ7g6_2),.clk(gclk));
	jdff dff_B_dHRuiRfN8_2(.din(w_dff_B_C1YSRQ7g6_2),.dout(w_dff_B_dHRuiRfN8_2),.clk(gclk));
	jdff dff_B_gyIJUMMZ3_2(.din(w_dff_B_dHRuiRfN8_2),.dout(w_dff_B_gyIJUMMZ3_2),.clk(gclk));
	jdff dff_B_g80eCCPX6_2(.din(w_dff_B_gyIJUMMZ3_2),.dout(w_dff_B_g80eCCPX6_2),.clk(gclk));
	jdff dff_B_qG9XMwlv3_2(.din(w_dff_B_g80eCCPX6_2),.dout(w_dff_B_qG9XMwlv3_2),.clk(gclk));
	jdff dff_B_y2pTILfZ0_2(.din(w_dff_B_qG9XMwlv3_2),.dout(w_dff_B_y2pTILfZ0_2),.clk(gclk));
	jdff dff_B_3lPSPYKv0_2(.din(w_dff_B_y2pTILfZ0_2),.dout(w_dff_B_3lPSPYKv0_2),.clk(gclk));
	jdff dff_B_n7AMVRDS9_2(.din(w_dff_B_3lPSPYKv0_2),.dout(w_dff_B_n7AMVRDS9_2),.clk(gclk));
	jdff dff_B_dC3ZPlEE3_2(.din(w_dff_B_n7AMVRDS9_2),.dout(w_dff_B_dC3ZPlEE3_2),.clk(gclk));
	jdff dff_B_efvfk0rc2_2(.din(w_dff_B_dC3ZPlEE3_2),.dout(w_dff_B_efvfk0rc2_2),.clk(gclk));
	jdff dff_B_yAhbeUEa0_2(.din(w_dff_B_efvfk0rc2_2),.dout(w_dff_B_yAhbeUEa0_2),.clk(gclk));
	jdff dff_B_dcLt4VgG0_2(.din(w_dff_B_yAhbeUEa0_2),.dout(w_dff_B_dcLt4VgG0_2),.clk(gclk));
	jdff dff_B_A9qn4Qed0_2(.din(w_dff_B_dcLt4VgG0_2),.dout(w_dff_B_A9qn4Qed0_2),.clk(gclk));
	jdff dff_B_RapIJeDF9_2(.din(w_dff_B_A9qn4Qed0_2),.dout(w_dff_B_RapIJeDF9_2),.clk(gclk));
	jdff dff_B_P6NmMIMJ3_2(.din(n1350),.dout(w_dff_B_P6NmMIMJ3_2),.clk(gclk));
	jdff dff_B_DXXp7Pxl5_1(.din(n1348),.dout(w_dff_B_DXXp7Pxl5_1),.clk(gclk));
	jdff dff_B_nRvwjuUq6_2(.din(n1262),.dout(w_dff_B_nRvwjuUq6_2),.clk(gclk));
	jdff dff_B_Y3IwIJ952_2(.din(w_dff_B_nRvwjuUq6_2),.dout(w_dff_B_Y3IwIJ952_2),.clk(gclk));
	jdff dff_B_g56VptH23_2(.din(w_dff_B_Y3IwIJ952_2),.dout(w_dff_B_g56VptH23_2),.clk(gclk));
	jdff dff_B_F4Zcur6t1_2(.din(w_dff_B_g56VptH23_2),.dout(w_dff_B_F4Zcur6t1_2),.clk(gclk));
	jdff dff_B_QpK5AMUf8_2(.din(w_dff_B_F4Zcur6t1_2),.dout(w_dff_B_QpK5AMUf8_2),.clk(gclk));
	jdff dff_B_gCNhqQai0_2(.din(w_dff_B_QpK5AMUf8_2),.dout(w_dff_B_gCNhqQai0_2),.clk(gclk));
	jdff dff_B_E5GXKQ5y1_2(.din(w_dff_B_gCNhqQai0_2),.dout(w_dff_B_E5GXKQ5y1_2),.clk(gclk));
	jdff dff_B_D4EnDcGT4_2(.din(w_dff_B_E5GXKQ5y1_2),.dout(w_dff_B_D4EnDcGT4_2),.clk(gclk));
	jdff dff_B_u8dIuvGZ8_2(.din(w_dff_B_D4EnDcGT4_2),.dout(w_dff_B_u8dIuvGZ8_2),.clk(gclk));
	jdff dff_B_sP4f4yKz7_2(.din(w_dff_B_u8dIuvGZ8_2),.dout(w_dff_B_sP4f4yKz7_2),.clk(gclk));
	jdff dff_B_SZvkzbvI6_2(.din(w_dff_B_sP4f4yKz7_2),.dout(w_dff_B_SZvkzbvI6_2),.clk(gclk));
	jdff dff_B_40f00axQ4_2(.din(w_dff_B_SZvkzbvI6_2),.dout(w_dff_B_40f00axQ4_2),.clk(gclk));
	jdff dff_B_p0tOgi460_2(.din(w_dff_B_40f00axQ4_2),.dout(w_dff_B_p0tOgi460_2),.clk(gclk));
	jdff dff_B_4yk26g6X3_1(.din(n1268),.dout(w_dff_B_4yk26g6X3_1),.clk(gclk));
	jdff dff_B_J2DV1nKB9_1(.din(w_dff_B_4yk26g6X3_1),.dout(w_dff_B_J2DV1nKB9_1),.clk(gclk));
	jdff dff_B_82hRT4OB5_2(.din(n1267),.dout(w_dff_B_82hRT4OB5_2),.clk(gclk));
	jdff dff_B_23VDLF7L9_2(.din(w_dff_B_82hRT4OB5_2),.dout(w_dff_B_23VDLF7L9_2),.clk(gclk));
	jdff dff_B_bNQIYJje6_2(.din(w_dff_B_23VDLF7L9_2),.dout(w_dff_B_bNQIYJje6_2),.clk(gclk));
	jdff dff_B_fO3eHuoT5_2(.din(w_dff_B_bNQIYJje6_2),.dout(w_dff_B_fO3eHuoT5_2),.clk(gclk));
	jdff dff_B_joOBfP5k2_2(.din(w_dff_B_fO3eHuoT5_2),.dout(w_dff_B_joOBfP5k2_2),.clk(gclk));
	jdff dff_B_wexHMndp0_2(.din(w_dff_B_joOBfP5k2_2),.dout(w_dff_B_wexHMndp0_2),.clk(gclk));
	jdff dff_B_c4S10mQb8_2(.din(w_dff_B_wexHMndp0_2),.dout(w_dff_B_c4S10mQb8_2),.clk(gclk));
	jdff dff_B_QUjYMaiX1_2(.din(w_dff_B_c4S10mQb8_2),.dout(w_dff_B_QUjYMaiX1_2),.clk(gclk));
	jdff dff_B_U4AZ5aEj3_2(.din(w_dff_B_QUjYMaiX1_2),.dout(w_dff_B_U4AZ5aEj3_2),.clk(gclk));
	jdff dff_B_rVQEiO3x4_2(.din(w_dff_B_U4AZ5aEj3_2),.dout(w_dff_B_rVQEiO3x4_2),.clk(gclk));
	jdff dff_B_7CGIm1Xs9_2(.din(n1266),.dout(w_dff_B_7CGIm1Xs9_2),.clk(gclk));
	jdff dff_B_rWU2nklD9_2(.din(w_dff_B_7CGIm1Xs9_2),.dout(w_dff_B_rWU2nklD9_2),.clk(gclk));
	jdff dff_B_5hTvil179_2(.din(w_dff_B_rWU2nklD9_2),.dout(w_dff_B_5hTvil179_2),.clk(gclk));
	jdff dff_B_ER393EM95_2(.din(w_dff_B_5hTvil179_2),.dout(w_dff_B_ER393EM95_2),.clk(gclk));
	jdff dff_B_4WCWY19K4_2(.din(w_dff_B_ER393EM95_2),.dout(w_dff_B_4WCWY19K4_2),.clk(gclk));
	jdff dff_B_9pndhanH1_2(.din(w_dff_B_4WCWY19K4_2),.dout(w_dff_B_9pndhanH1_2),.clk(gclk));
	jdff dff_B_PCUxEJIg2_2(.din(w_dff_B_9pndhanH1_2),.dout(w_dff_B_PCUxEJIg2_2),.clk(gclk));
	jdff dff_B_LrnxgylS7_2(.din(w_dff_B_PCUxEJIg2_2),.dout(w_dff_B_LrnxgylS7_2),.clk(gclk));
	jdff dff_B_s6zl5eHJ9_2(.din(w_dff_B_LrnxgylS7_2),.dout(w_dff_B_s6zl5eHJ9_2),.clk(gclk));
	jdff dff_B_awqix9DE7_2(.din(w_dff_B_s6zl5eHJ9_2),.dout(w_dff_B_awqix9DE7_2),.clk(gclk));
	jdff dff_B_RrL3WYwu1_2(.din(w_dff_B_awqix9DE7_2),.dout(w_dff_B_RrL3WYwu1_2),.clk(gclk));
	jdff dff_B_HO6FzM4K1_2(.din(w_dff_B_RrL3WYwu1_2),.dout(w_dff_B_HO6FzM4K1_2),.clk(gclk));
	jdff dff_B_9nPMHveG8_1(.din(n1263),.dout(w_dff_B_9nPMHveG8_1),.clk(gclk));
	jdff dff_B_XdtLQB7X6_2(.din(n1171),.dout(w_dff_B_XdtLQB7X6_2),.clk(gclk));
	jdff dff_B_hwKN7OCW4_2(.din(w_dff_B_XdtLQB7X6_2),.dout(w_dff_B_hwKN7OCW4_2),.clk(gclk));
	jdff dff_B_6wYcFkxl1_2(.din(w_dff_B_hwKN7OCW4_2),.dout(w_dff_B_6wYcFkxl1_2),.clk(gclk));
	jdff dff_B_eaKJy4xE4_2(.din(w_dff_B_6wYcFkxl1_2),.dout(w_dff_B_eaKJy4xE4_2),.clk(gclk));
	jdff dff_B_0fGhoOSl2_2(.din(w_dff_B_eaKJy4xE4_2),.dout(w_dff_B_0fGhoOSl2_2),.clk(gclk));
	jdff dff_B_HOwsr0M04_2(.din(w_dff_B_0fGhoOSl2_2),.dout(w_dff_B_HOwsr0M04_2),.clk(gclk));
	jdff dff_B_5KbKsbZn8_2(.din(w_dff_B_HOwsr0M04_2),.dout(w_dff_B_5KbKsbZn8_2),.clk(gclk));
	jdff dff_B_J9IEz1r19_2(.din(w_dff_B_5KbKsbZn8_2),.dout(w_dff_B_J9IEz1r19_2),.clk(gclk));
	jdff dff_B_ADuKv0yc5_2(.din(w_dff_B_J9IEz1r19_2),.dout(w_dff_B_ADuKv0yc5_2),.clk(gclk));
	jdff dff_B_LKBWQccQ1_2(.din(w_dff_B_ADuKv0yc5_2),.dout(w_dff_B_LKBWQccQ1_2),.clk(gclk));
	jdff dff_B_3LF1fFik5_2(.din(w_dff_B_LKBWQccQ1_2),.dout(w_dff_B_3LF1fFik5_2),.clk(gclk));
	jdff dff_B_KpCmnpil7_2(.din(n1182),.dout(w_dff_B_KpCmnpil7_2),.clk(gclk));
	jdff dff_B_0koEPZvE1_1(.din(n1177),.dout(w_dff_B_0koEPZvE1_1),.clk(gclk));
	jdff dff_B_mW7jJoG59_1(.din(w_dff_B_0koEPZvE1_1),.dout(w_dff_B_mW7jJoG59_1),.clk(gclk));
	jdff dff_B_bPZJas5R4_2(.din(n1176),.dout(w_dff_B_bPZJas5R4_2),.clk(gclk));
	jdff dff_B_4fhzi4Bd0_2(.din(w_dff_B_bPZJas5R4_2),.dout(w_dff_B_4fhzi4Bd0_2),.clk(gclk));
	jdff dff_B_97e0JX4Y1_2(.din(w_dff_B_4fhzi4Bd0_2),.dout(w_dff_B_97e0JX4Y1_2),.clk(gclk));
	jdff dff_B_5CtKi17v4_2(.din(w_dff_B_97e0JX4Y1_2),.dout(w_dff_B_5CtKi17v4_2),.clk(gclk));
	jdff dff_B_RHiQYOYh5_2(.din(w_dff_B_5CtKi17v4_2),.dout(w_dff_B_RHiQYOYh5_2),.clk(gclk));
	jdff dff_B_s7rXv6oG9_2(.din(w_dff_B_RHiQYOYh5_2),.dout(w_dff_B_s7rXv6oG9_2),.clk(gclk));
	jdff dff_B_1YbWHAfd8_2(.din(w_dff_B_s7rXv6oG9_2),.dout(w_dff_B_1YbWHAfd8_2),.clk(gclk));
	jdff dff_B_XpA3bmsu4_2(.din(n1175),.dout(w_dff_B_XpA3bmsu4_2),.clk(gclk));
	jdff dff_B_Un1YDpde2_2(.din(w_dff_B_XpA3bmsu4_2),.dout(w_dff_B_Un1YDpde2_2),.clk(gclk));
	jdff dff_B_BXuAESMg7_2(.din(w_dff_B_Un1YDpde2_2),.dout(w_dff_B_BXuAESMg7_2),.clk(gclk));
	jdff dff_B_IFJ7U6Uv5_2(.din(w_dff_B_BXuAESMg7_2),.dout(w_dff_B_IFJ7U6Uv5_2),.clk(gclk));
	jdff dff_B_VLnNGJHJ5_2(.din(w_dff_B_IFJ7U6Uv5_2),.dout(w_dff_B_VLnNGJHJ5_2),.clk(gclk));
	jdff dff_B_1P3xHSq93_2(.din(w_dff_B_VLnNGJHJ5_2),.dout(w_dff_B_1P3xHSq93_2),.clk(gclk));
	jdff dff_B_fp6zLPHS6_2(.din(w_dff_B_1P3xHSq93_2),.dout(w_dff_B_fp6zLPHS6_2),.clk(gclk));
	jdff dff_B_5t0S9Tc66_2(.din(w_dff_B_fp6zLPHS6_2),.dout(w_dff_B_5t0S9Tc66_2),.clk(gclk));
	jdff dff_B_ec9y6jOn3_2(.din(w_dff_B_5t0S9Tc66_2),.dout(w_dff_B_ec9y6jOn3_2),.clk(gclk));
	jdff dff_B_LvUd9uLj8_1(.din(n1172),.dout(w_dff_B_LvUd9uLj8_1),.clk(gclk));
	jdff dff_B_kmHm9Wpt5_2(.din(n1073),.dout(w_dff_B_kmHm9Wpt5_2),.clk(gclk));
	jdff dff_B_X5V6kJyn2_2(.din(w_dff_B_kmHm9Wpt5_2),.dout(w_dff_B_X5V6kJyn2_2),.clk(gclk));
	jdff dff_B_i8NYvCSz4_2(.din(w_dff_B_X5V6kJyn2_2),.dout(w_dff_B_i8NYvCSz4_2),.clk(gclk));
	jdff dff_B_gZBN4ew09_2(.din(w_dff_B_i8NYvCSz4_2),.dout(w_dff_B_gZBN4ew09_2),.clk(gclk));
	jdff dff_B_sGm4xLkU6_2(.din(w_dff_B_gZBN4ew09_2),.dout(w_dff_B_sGm4xLkU6_2),.clk(gclk));
	jdff dff_B_tYzdjnY44_2(.din(w_dff_B_sGm4xLkU6_2),.dout(w_dff_B_tYzdjnY44_2),.clk(gclk));
	jdff dff_B_DTtGETrj7_2(.din(w_dff_B_tYzdjnY44_2),.dout(w_dff_B_DTtGETrj7_2),.clk(gclk));
	jdff dff_B_XrMHkfLs9_2(.din(w_dff_B_DTtGETrj7_2),.dout(w_dff_B_XrMHkfLs9_2),.clk(gclk));
	jdff dff_B_1Wo4CiF30_2(.din(w_dff_B_XrMHkfLs9_2),.dout(w_dff_B_1Wo4CiF30_2),.clk(gclk));
	jdff dff_B_S5tqoVU85_2(.din(n1083),.dout(w_dff_B_S5tqoVU85_2),.clk(gclk));
	jdff dff_B_5RHH1Fax3_2(.din(w_dff_B_S5tqoVU85_2),.dout(w_dff_B_5RHH1Fax3_2),.clk(gclk));
	jdff dff_B_Br8rk8lT2_2(.din(n1078),.dout(w_dff_B_Br8rk8lT2_2),.clk(gclk));
	jdff dff_B_0t79R8j42_2(.din(w_dff_B_Br8rk8lT2_2),.dout(w_dff_B_0t79R8j42_2),.clk(gclk));
	jdff dff_B_O2P6ExlF7_2(.din(w_dff_B_0t79R8j42_2),.dout(w_dff_B_O2P6ExlF7_2),.clk(gclk));
	jdff dff_B_SSM5SvsX8_2(.din(w_dff_B_O2P6ExlF7_2),.dout(w_dff_B_SSM5SvsX8_2),.clk(gclk));
	jdff dff_B_fdbm5c8k8_2(.din(n1077),.dout(w_dff_B_fdbm5c8k8_2),.clk(gclk));
	jdff dff_B_BjhJC7Mp1_2(.din(w_dff_B_fdbm5c8k8_2),.dout(w_dff_B_BjhJC7Mp1_2),.clk(gclk));
	jdff dff_B_DL47iGsn1_2(.din(w_dff_B_BjhJC7Mp1_2),.dout(w_dff_B_DL47iGsn1_2),.clk(gclk));
	jdff dff_B_w74yMYTa7_2(.din(w_dff_B_DL47iGsn1_2),.dout(w_dff_B_w74yMYTa7_2),.clk(gclk));
	jdff dff_B_h0WeFLoh1_2(.din(w_dff_B_w74yMYTa7_2),.dout(w_dff_B_h0WeFLoh1_2),.clk(gclk));
	jdff dff_B_HQl7EJU00_2(.din(w_dff_B_h0WeFLoh1_2),.dout(w_dff_B_HQl7EJU00_2),.clk(gclk));
	jdff dff_B_cv0a7YUk9_1(.din(n1074),.dout(w_dff_B_cv0a7YUk9_1),.clk(gclk));
	jdff dff_B_Gz9mkbZW3_2(.din(n974),.dout(w_dff_B_Gz9mkbZW3_2),.clk(gclk));
	jdff dff_B_3j5auCwl7_2(.din(w_dff_B_Gz9mkbZW3_2),.dout(w_dff_B_3j5auCwl7_2),.clk(gclk));
	jdff dff_B_pOROb8Pk7_2(.din(w_dff_B_3j5auCwl7_2),.dout(w_dff_B_pOROb8Pk7_2),.clk(gclk));
	jdff dff_B_3R0Sen8r1_2(.din(w_dff_B_pOROb8Pk7_2),.dout(w_dff_B_3R0Sen8r1_2),.clk(gclk));
	jdff dff_B_UfCzOdpd3_2(.din(w_dff_B_3R0Sen8r1_2),.dout(w_dff_B_UfCzOdpd3_2),.clk(gclk));
	jdff dff_B_ChYkX4iW9_2(.din(w_dff_B_UfCzOdpd3_2),.dout(w_dff_B_ChYkX4iW9_2),.clk(gclk));
	jdff dff_B_wCp8FuyK2_2(.din(w_dff_B_ChYkX4iW9_2),.dout(w_dff_B_wCp8FuyK2_2),.clk(gclk));
	jdff dff_B_TyAkCYbZ4_2(.din(n984),.dout(w_dff_B_TyAkCYbZ4_2),.clk(gclk));
	jdff dff_B_ZorCzA459_2(.din(w_dff_B_TyAkCYbZ4_2),.dout(w_dff_B_ZorCzA459_2),.clk(gclk));
	jdff dff_B_drOzPVID4_2(.din(w_dff_B_ZorCzA459_2),.dout(w_dff_B_drOzPVID4_2),.clk(gclk));
	jdff dff_B_0GefHd6l8_2(.din(n983),.dout(w_dff_B_0GefHd6l8_2),.clk(gclk));
	jdff dff_B_6JgC3XOe7_2(.din(w_dff_B_0GefHd6l8_2),.dout(w_dff_B_6JgC3XOe7_2),.clk(gclk));
	jdff dff_B_PNRnO2Eg7_2(.din(w_dff_B_6JgC3XOe7_2),.dout(w_dff_B_PNRnO2Eg7_2),.clk(gclk));
	jdff dff_A_2dt4Jpqk0_0(.dout(w_n980_0[0]),.din(w_dff_A_2dt4Jpqk0_0),.clk(gclk));
	jdff dff_A_5ImTVvdP6_0(.dout(w_dff_A_2dt4Jpqk0_0),.din(w_dff_A_5ImTVvdP6_0),.clk(gclk));
	jdff dff_B_cde1KABN0_2(.din(n980),.dout(w_dff_B_cde1KABN0_2),.clk(gclk));
	jdff dff_A_9MgiCG545_0(.dout(w_n877_0[0]),.din(w_dff_A_9MgiCG545_0),.clk(gclk));
	jdff dff_A_jqTD4e0F0_0(.dout(w_dff_A_9MgiCG545_0),.din(w_dff_A_jqTD4e0F0_0),.clk(gclk));
	jdff dff_A_d5Hs080Z2_0(.dout(w_dff_A_jqTD4e0F0_0),.din(w_dff_A_d5Hs080Z2_0),.clk(gclk));
	jdff dff_B_NlKQY1ue6_2(.din(n877),.dout(w_dff_B_NlKQY1ue6_2),.clk(gclk));
	jdff dff_A_G9SnM9lB2_0(.dout(w_n875_0[0]),.din(w_dff_A_G9SnM9lB2_0),.clk(gclk));
	jdff dff_A_64J3g8NG2_0(.dout(w_dff_A_G9SnM9lB2_0),.din(w_dff_A_64J3g8NG2_0),.clk(gclk));
	jdff dff_B_ZBbanpTL9_2(.din(n874),.dout(w_dff_B_ZBbanpTL9_2),.clk(gclk));
	jdff dff_B_xjGe0H5j2_2(.din(w_dff_B_ZBbanpTL9_2),.dout(w_dff_B_xjGe0H5j2_2),.clk(gclk));
endmodule

